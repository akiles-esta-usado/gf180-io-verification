* NGSPICE file created from gf180mcu_fd_io__in_c_pex.ext - technology: gf180mcuD

.subckt gf180mcu_fd_io__in_c_pex DVSS DVDD PAD Y PD VSS VDD PU
X0 GF_NI_IN_C_BASE_0.comp018green_out_predrv_1.ENB.t0 GF_NI_IN_C_BASE_0.comp018green_out_predrv_1.EN.t1 DVDD.t194 DVDD.t193 pfet_06v0 ad=2.64p pd=12.879999u as=1.56p ps=6.52u w=6u l=0.7u
X1 GF_NI_IN_C_BASE_0.pdrive_y_<1>.t0 GF_NI_IN_C_BASE_0.comp018green_out_predrv_0.SLB.t2 GF_NI_IN_C_BASE_0.pdrive_x_<1>.t1 DVSS.t35 nfet_06v0 ad=1.56p pd=6.52u as=2.64p ps=12.879999u w=6u l=0.7u
X2 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_cms_smt_0.nmos_6p0_CDNS_4066195314540_0.S.t3 GF_NI_IN_C_BASE_0.comp018green_esd_cdm_0.IP_IN.t1 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_drv_0.A.t6 DVSS.t16 nfet_06v0 ad=1.32p pd=6.88u as=0.78p ps=3.52u w=3u l=0.7u
X3 PU.t1 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_logic_pupd_0.comp018green_std_xor2_0.nmos_6p0_CDNS_4066195314530_0.D.t1 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_logic_pupd_0.comp018green_std_nand2_0.A.t0 VSS.t46 nfet_06v0 ad=0.66p pd=3.88u as=0.66p ps=3.88u w=1.5u l=0.7u
X4 VDD.t37 PU.t2 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_logic_pupd_0.comp018green_std_xor2_0.nmos_6p0_CDNS_4066195314530_2.D.t0 VDD.t36 pfet_06v0 ad=1.32p pd=6.88u as=1.32p ps=6.88u w=3u l=0.7u
X5 VSS.t13 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.t6 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_1.nmos_6p0_CDNS_4066195314511_0.S.t0 VSS.t12 nfet_06v0 ad=1.32p pd=6.88u as=0.78p ps=3.52u w=3u l=0.7u
X6 GF_NI_IN_C_BASE_0.comp018green_out_predrv_1.nmos_6p0_CDNS_4066195314519_0.D.t0 GF_NI_IN_C_BASE_0.comp018green_out_predrv_0.A.t2 DVSS.t6 DVSS.t5 nfet_06v0 ad=2.64p pd=12.879999u as=1.56p ps=6.52u w=6u l=0.7u
X7 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_pupd_0.ppolyf_u_CDNS_4066195314532_0.PLUS PAD.t15 w_4468_53312# ppolyf_u r_width=2.5u r_length=2.8u
X8 DVSS.t192 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_1.nmos_6p0_CDNS_4066195314530_0.D.t2 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_1.Z.t0 DVSS.t191 nfet_06v0 ad=0.39p pd=2.02u as=0.39p ps=2.02u w=1.5u l=0.7u
X9 Y.t5 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_drv_0.Z.t1 VSS.t34 VSS.t33 nfet_06v0 ad=0.39p pd=2.02u as=0.39p ps=2.02u w=1.5u l=0.7u
X10 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.nmos_6p0_CDNS_4066195314511_1.S.t0 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.t7 VDD.t17 VDD.t16 pfet_06v0 ad=0.78p pd=3.52u as=1.32p ps=6.88u w=3u l=0.7u
X11 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_1.nmos_6p0_CDNS_4066195314511_0.S.t1 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.t8 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_1.nmos_6p0_CDNS_4066195314511_1.S.t0 VSS.t11 nfet_06v0 ad=0.78p pd=3.52u as=1.32p ps=6.88u w=3u l=0.7u
X12 VSS.t10 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.t9 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_a_0.nmos_6p0_CDNS_4066195314511_1.S.t0 VSS.t9 nfet_06v0 ad=1.32p pd=6.88u as=0.78p ps=3.52u w=3u l=0.7u
X13 GF_NI_IN_C_BASE_0.ndrive_Y_<1>.t4 GF_NI_IN_C_BASE_0.comp018green_out_predrv_3.nmos_6p0_CDNS_4066195314519_2.S.t2 DVDD.t57 DVDD.t56 pfet_06v0 ad=5.28p pd=24.88u as=3.12p ps=12.52u w=11.999999u l=0.7u
X14 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_drv_0.nmos_6p0_CDNS_4066195314547_0.S.t2 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_drv_0.A.t9 DVDD.t30 DVDD.t29 pfet_06v0 ad=0.88p pd=4.88u as=0.88p ps=4.88u w=2u l=0.7u
D0 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_pupd_0.ppolyf_u_CDNS_4066195314532_0.PLUS DVDD diode_pd2nw_06v0 pj=42u area=20p
X15 GF_NI_IN_C_BASE_0.comp018green_out_predrv_2.nmos_6p0_CDNS_4066195314519_2.S.t1 GF_NI_IN_C_BASE_0.comp018green_out_predrv_0.A.t3 DVDD.t6 DVDD.t5 pfet_06v0 ad=5.28p pd=24.88u as=3.12p ps=12.52u w=11.999999u l=0.7u
X16 GF_NI_IN_C_BASE_0.ndrive_x_<2>.t2 GF_NI_IN_C_BASE_0.comp018green_out_predrv_2.nmos_6p0_CDNS_4066195314519_2.S.t2 DVSS.t163 DVSS.t162 nfet_06v0 ad=1.56p pd=6.52u as=2.64p ps=12.879999u w=6u l=0.7u
X17 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_a_0.nmos_6p0_CDNS_4066195314511_1.S.t1 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.t10 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_a_0.nmos_6p0_CDNS_4066195314511_1.D.t0 VSS.t8 nfet_06v0 ad=0.78p pd=3.52u as=1.32p ps=6.88u w=3u l=0.7u
X18 PAD GF_NI_IN_C_BASE_0.ndrive_x_<0>.t3 DVSS DVSS.t25 nfet_06v0_dss d_sab=3.78u s_sab=0.28u ad=0.14364n pd=83.56u as=10.639999p ps=76.56u w=38u l=1.15u
X19 DVDD.t198 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_1.EN.t2 GF_NI_IN_C_BASE_0.comp018green_out_predrv_2.nmos_6p0_CDNS_4066195314519_2.S.t0 DVDD.t197 pfet_06v0 ad=3.12p pd=12.52u as=3.12p ps=12.52u w=11.999999u l=0.7u
X20 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_0.nmos_6p0_CDNS_4066195314530_0.D.t1 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_logic_pupd_0.PDB_OUT.t1 VDD.t21 VDD.t20 pfet_06v0 ad=1.32p pd=6.88u as=1.32p ps=6.88u w=3u l=0.7u
X21 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_pupd_0.ppolyf_u_CDNS_4066195314533_0.PLUS.t0 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_pupd_0.ppolyf_u_CDNS_4066195314533_0.MINUS.t0 DVDD.t40 ppolyf_u r_width=0.8u r_length=35.7u
X22 GF_NI_IN_C_BASE_0.comp018green_out_predrv_0.SLB.t0 GF_NI_IN_C_BASE_0.comp018green_out_predrv_0.SL.t2 DVDD.t39 DVDD.t38 pfet_06v0 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.7u
X23 DVDD GF_NI_IN_C_BASE_0.pdrive_x_<2>.t4 PAD DVDD.t157 pfet_06v0_dss d_sab=0.28u s_sab=2.78u ad=11.199999p pd=80.56u as=0.1112n ps=85.56u w=40u l=0.7u
X24 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_1.nmos_6p0_CDNS_4066195314530_0.D.t0 GF_NI_IN_C_BASE_0.ppolyf_u_CDNS_4066195314551_0.MINUS.t1 VSS.t45 VSS.t44 nfet_06v0 ad=0.66p pd=3.88u as=0.66p ps=3.88u w=1.5u l=0.7u
X25 DVSS.t153 GF_NI_IN_C_BASE_0.comp018green_out_predrv_0.nmos_6p0_CDNS_4066195314519_2.S.t2 GF_NI_IN_C_BASE_0.ndrive_y_<0>.t0 DVSS.t152 nfet_06v0 ad=1.56p pd=6.52u as=1.56p ps=6.52u w=6u l=0.7u
X26 PAD GF_NI_IN_C_BASE_0.pdrive_x_<0>.t4 DVDD DVDD.t99 pfet_06v0_dss d_sab=2.78u s_sab=0.28u ad=0.1112n pd=85.56u as=11.199999p ps=80.56u w=40u l=0.7u
X27 DVSS.t143 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_2.nmos_6p0_CDNS_4066195314530_0.D.t2 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_pupd_0.PU_B.t0 DVSS.t142 nfet_06v0 ad=0.66p pd=3.88u as=0.39p ps=2.02u w=1.5u l=0.7u
X28 DVDD.t170 GF_NI_IN_C_BASE_0.comp018green_out_predrv_0.nmos_6p0_CDNS_4066195314519_0.D.t3 GF_NI_IN_C_BASE_0.pdrive_x_<0>.t3 DVDD.t169 pfet_06v0 ad=5.28p pd=24.88u as=3.12p ps=12.52u w=11.999999u l=0.7u
X29 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_0.Z.t0 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_0.nmos_6p0_CDNS_4066195314530_0.D.t2 DVSS.t170 DVSS.t169 nfet_06v0 ad=0.39p pd=2.02u as=0.66p ps=3.88u w=1.5u l=0.7u
X30 GF_NI_IN_C_BASE_0.ndrive_y_<0>.t0 GF_NI_IN_C_BASE_0.comp018green_out_predrv_0.nmos_6p0_CDNS_4066195314519_2.S.t3 DVSS.t155 DVSS.t154 nfet_06v0 ad=1.56p pd=6.52u as=1.56p ps=6.52u w=6u l=0.7u
X31 DVDD.t81 GF_NI_IN_C_BASE_0.comp018green_out_predrv_2.nmos_6p0_CDNS_4066195314519_0.D.t3 GF_NI_IN_C_BASE_0.pdrive_y_<2>.t3 DVDD.t80 pfet_06v0 ad=3.12p pd=12.52u as=3.12p ps=12.52u w=11.999999u l=0.7u
X32 DVSS.t182 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_1.Z.t2 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_cms_smt_0.nmos_6p0_CDNS_4066195314537_0.D.t2 DVSS.t181 nfet_06v0 ad=0.832p pd=3.72u as=0.832p ps=3.72u w=3.2u l=0.7u
X33 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_cms_smt_0.nmos_6p0_CDNS_4066195314536_1.S.t2 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_3.Z.t1 DVDD.t117 DVDD.t116 pfet_06v0 ad=0.39p pd=2.02u as=0.66p ps=3.88u w=1.5u l=0.7u
X34 DVDD.t139 GF_NI_IN_C_BASE_0.comp018green_out_predrv_1.nmos_6p0_CDNS_4066195314519_2.S.t2 GF_NI_IN_C_BASE_0.ndrive_Y_<3>.t2 DVDD.t138 pfet_06v0 ad=3.12p pd=12.52u as=3.12p ps=12.52u w=11.999999u l=0.7u
X35 GF_NI_IN_C_BASE_0.comp018green_out_predrv_3.nmos_6p0_CDNS_4066195314519_2.S.t0 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_1.EN.t3 DVDD.t64 DVDD.t63 pfet_06v0 ad=3.12p pd=12.52u as=3.12p ps=12.52u w=11.999999u l=0.7u
X36 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_cms_smt_0.nmos_6p0_CDNS_4066195314537_0.D.t2 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_1.Z.t3 DVSS.t184 DVSS.t183 nfet_06v0 ad=0.832p pd=3.72u as=0.832p ps=3.72u w=3.2u l=0.7u
X37 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_drv_0.A.t4 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_3.Z.t2 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_cms_smt_0.nmos_6p0_CDNS_4066195314536_1.S.t1 DVSS.t117 nfet_06v0 ad=0.66p pd=3.88u as=0.66p ps=3.88u w=1.5u l=0.7u
X38 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_pupd_0.ppolyf_u_CDNS_4066195314533_1.PLUS.t0 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_pupd_0.ppolyf_u_CDNS_4066195314533_1.MINUS.t0 DVDD.t40 ppolyf_u r_width=0.8u r_length=35.7u
X39 DVDD.t184 GF_NI_IN_C_BASE_0.comp018green_out_predrv_3.nmos_6p0_CDNS_4066195314519_0.D.t3 GF_NI_IN_C_BASE_0.pdrive_y_<1>.t3 DVDD.t183 pfet_06v0 ad=5.28p pd=24.88u as=3.12p ps=12.52u w=11.999999u l=0.7u
X40 VDD.t19 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.t11 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_3.nmos_6p0_CDNS_4066195314530_0.D.t1 VDD.t18 pfet_06v0 ad=1.32p pd=6.88u as=1.32p ps=6.88u w=3u l=0.7u
X41 DVSS.t134 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_0.Z.t2 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_pupd_0.PD.t0 DVSS.t133 nfet_06v0 ad=0.66p pd=3.88u as=0.39p ps=2.02u w=1.5u l=0.7u
X42 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_cms_smt_0.nmos_6p0_CDNS_4066195314540_0.S.t0 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_cms_smt_0.nmos_6p0_CDNS_4066195314530_0.D.t2 DVDD.t55 DVSS.t63 nfet_06v0 ad=0.572p pd=3.48u as=0.572p ps=3.48u w=1.3u l=0.7u
X43 GF_NI_IN_C_BASE_0.ndrive_Y_<3>.t2 GF_NI_IN_C_BASE_0.comp018green_out_predrv_0.SL.t3 GF_NI_IN_C_BASE_0.ndrive_x_<3>.t2 DVDD.t52 pfet_06v0 ad=3.12p pd=12.52u as=3.12p ps=12.52u w=11.999999u l=0.7u
D1 GF_NI_IN_C_BASE_0.ppolyf_u_CDNS_4066195314551_0.MINUS.t1 VDD.t58 diode_pd2nw_06v0 pj=4u area=1p
X44 GF_NI_IN_C_BASE_0.ndrive_y_<2>.t2 GF_NI_IN_C_BASE_0.comp018green_out_predrv_0.SL.t4 GF_NI_IN_C_BASE_0.ndrive_x_<2>.t0 DVDD.t53 pfet_06v0 ad=5.28p pd=24.88u as=3.12p ps=12.52u w=11.999999u l=0.7u
X45 GF_NI_IN_C_BASE_0.ndrive_x_<3>.t1 DVSS.t204 GF_NI_IN_C_BASE_0.ndrive_Y_<3>.t3 DVDD.t201 pfet_06v0 ad=0.528p pd=3.28u as=0.528p ps=3.28u w=1.2u l=0.7u
X46 DVSS.t69 GF_NI_IN_C_BASE_0.comp018green_out_predrv_3.nmos_6p0_CDNS_4066195314519_2.S.t3 GF_NI_IN_C_BASE_0.ndrive_x_<1>.t1 DVSS.t68 nfet_06v0 ad=2.64p pd=12.879999u as=1.56p ps=6.52u w=6u l=0.7u
X47 DVSS.t24 GF_NI_IN_C_BASE_0.comp018green_out_predrv_0.A.t4 GF_NI_IN_C_BASE_0.comp018green_out_predrv_2.nmos_6p0_CDNS_4066195314519_0.D.t2 DVSS.t23 nfet_06v0 ad=1.56p pd=6.52u as=2.64p ps=12.879999u w=6u l=0.7u
X48 VDD.t15 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.t12 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_1.nmos_6p0_CDNS_4066195314511_1.S.t1 VDD.t14 pfet_06v0 ad=1.32p pd=6.88u as=0.78p ps=3.52u w=3u l=0.7u
X49 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_logic_pupd_0.comp018green_std_nand2_0.A.t1 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_logic_pupd_0.comp018green_std_xor2_0.nmos_6p0_CDNS_4066195314530_0.D.t2 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_logic_pupd_0.comp018green_std_xor2_0.nmos_6p0_CDNS_4066195314530_2.D.t3 VDD.t65 pfet_06v0 ad=1.32p pd=6.88u as=1.32p ps=6.88u w=3u l=0.7u
X50 GF_NI_IN_C_BASE_0.pdrive_y_<0>.t3 GF_NI_IN_C_BASE_0.comp018green_out_predrv_0.nmos_6p0_CDNS_4066195314519_0.D.t4 DVDD.t172 DVDD.t171 pfet_06v0 ad=3.12p pd=12.52u as=5.28p ps=24.88u w=11.999999u l=0.7u
X51 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_1.nmos_6p0_CDNS_4066195314511_1.S.t1 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.t13 VDD.t13 VDD.t12 pfet_06v0 ad=0.78p pd=3.52u as=1.32p ps=6.88u w=3u l=0.7u
X52 VDD.t11 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.t14 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_a_0.nmos_6p0_CDNS_4066195314511_1.D.t1 VDD.t10 pfet_06v0 ad=1.32p pd=6.88u as=0.78p ps=3.52u w=3u l=0.7u
X53 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_a_0.nmos_6p0_CDNS_4066195314511_1.D.t1 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.t15 VDD.t9 VDD.t8 pfet_06v0 ad=0.78p pd=3.52u as=1.32p ps=6.88u w=3u l=0.7u
X54 GF_NI_IN_C_BASE_0.ppolyf_u_CDNS_4066195314551_0.MINUS.t0 VDD.t23 VDD.t22 ppolyf_u r_width=0.8u r_length=3.9u
X55 DVDD.t188 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_1.Z.t4 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_1.ZB.t1 DVDD.t187 pfet_06v0 ad=1.32p pd=6.88u as=0.78p ps=3.52u w=3u l=0.7u
X56 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_1.ZB.t1 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_1.Z.t5 DVDD.t190 DVDD.t189 pfet_06v0 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.7u
X57 VSS.t29 PU.t3 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_logic_pupd_0.comp018green_std_nand2_1.nmos_6p0_CDNS_4066195314511_0.D.t0 VSS.t28 nfet_06v0 ad=1.32p pd=6.88u as=0.78p ps=3.52u w=3u l=0.7u
X58 GF_NI_IN_C_BASE_0.pdrive_x_<0>.t2 DVDD.t205 GF_NI_IN_C_BASE_0.pdrive_y_<0>.t1 DVSS.t34 nfet_06v0 ad=0.528p pd=3.28u as=0.528p ps=3.28u w=1.2u l=0.7u
X59 PAD GF_NI_IN_C_BASE_0.pdrive_y_<0>.t4 DVDD DVDD.t113 pfet_06v0_dss d_sab=2.78u s_sab=0.28u ad=0.1112n pd=85.56u as=11.199999p ps=80.56u w=40u l=0.7u
X60 a_5575_62984.t5 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_cms_smt_0.nmos_6p0_CDNS_4066195314536_1.S.t3 DVSS.t173 DVDD.t175 pfet_06v0 ad=0.836p pd=4.68u as=0.494p ps=2.42u w=1.9u l=0.7u
X61 GF_NI_IN_C_BASE_0.comp018green_sigbuf_1_0.nmos_6p0_CDNS_4066195314530_0.D.t1 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.t16 VDD.t7 VDD.t6 pfet_06v0 ad=1.32p pd=6.88u as=1.32p ps=6.88u w=3u l=0.7u
X62 DVSS.t161 GF_NI_IN_C_BASE_0.comp018green_out_predrv_1.ENB.t2 GF_NI_IN_C_BASE_0.comp018green_out_predrv_1.nmos_6p0_CDNS_4066195314519_0.D.t1 DVSS.t160 nfet_06v0 ad=1.56p pd=6.52u as=1.56p ps=6.52u w=6u l=0.7u
X63 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.t0 VSS.t30 VDD.t38 ppolyf_u r_width=0.8u r_length=3.9u
X64 DVSS GF_NI_IN_C_BASE_0.ndrive_Y_<3>.t5 PAD DVSS.t130 nfet_06v0_dss d_sab=0.28u s_sab=3.78u ad=10.639999p pd=76.56u as=0.14364n ps=83.56u w=38u l=1.15u
X65 DVSS.t178 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_cms_smt_0.nmos_6p0_CDNS_4066195314536_1.S.t4 a_5575_62984.t4 DVDD.t182 pfet_06v0 ad=0.494p pd=2.42u as=0.836p ps=4.68u w=1.9u l=0.7u
X66 VDD.t35 PU.t4 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_logic_pupd_0.PUB_OUT.t0 VDD.t34 pfet_06v0 ad=1.32p pd=6.88u as=0.78p ps=3.52u w=3u l=0.7u
X67 GF_NI_IN_C_BASE_0.pdrive_x_<0>.t1 GF_NI_IN_C_BASE_0.comp018green_out_predrv_0.SLB.t3 GF_NI_IN_C_BASE_0.pdrive_y_<0>.t0 DVSS.t34 nfet_06v0 ad=2.64p pd=12.879999u as=1.56p ps=6.52u w=6u l=0.7u
X68 DVDD.t8 GF_NI_IN_C_BASE_0.comp018green_out_predrv_1.nmos_6p0_CDNS_4066195314519_0.D.t3 GF_NI_IN_C_BASE_0.pdrive_x_<3>.t3 DVDD.t7 pfet_06v0 ad=3.12p pd=12.52u as=3.12p ps=12.52u w=11.999999u l=0.7u
X69 GF_NI_IN_C_BASE_0.pdrive_y_<1>.t3 GF_NI_IN_C_BASE_0.comp018green_out_predrv_3.nmos_6p0_CDNS_4066195314519_0.D.t4 DVDD.t186 DVDD.t185 pfet_06v0 ad=3.12p pd=12.52u as=3.12p ps=12.52u w=11.999999u l=0.7u
X70 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_drv_0.nmos_6p0_CDNS_4066195314547_0.S.t1 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_drv_0.A.t10 DVSS.t20 DVSS.t19 nfet_06v0 ad=1.76p pd=8.88u as=1.04p ps=4.52u w=4u l=0.7u
X71 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_pupd_0.ppolyf_u_CDNS_4066195314533_0.PLUS.t1 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_pupd_0.ppolyf_u_CDNS_4066195314533_1.MINUS.t1 DVDD.t40 ppolyf_u r_width=0.8u r_length=35.7u
X72 PAD GF_NI_IN_C_BASE_0.pdrive_x_<2>.t5 DVDD DVDD.t160 pfet_06v0_dss d_sab=2.78u s_sab=0.28u ad=0.1112n pd=85.56u as=11.199999p ps=80.56u w=40u l=0.7u
X73 GF_NI_IN_C_BASE_0.comp018green_out_predrv_1.nmos_6p0_CDNS_4066195314519_0.D.t2 GF_NI_IN_C_BASE_0.comp018green_out_predrv_1.ENB.t3 GF_NI_IN_C_BASE_0.comp018green_out_predrv_1.nmos_6p0_CDNS_4066195314519_2.S.t1 DVDD.t18 pfet_06v0 ad=5.28p pd=24.88u as=3.12p ps=12.52u w=11.999999u l=0.7u
X74 GF_NI_IN_C_BASE_0.pdrive_x_<3>.t3 GF_NI_IN_C_BASE_0.comp018green_out_predrv_1.nmos_6p0_CDNS_4066195314519_0.D.t4 DVDD.t1 DVDD.t0 pfet_06v0 ad=3.12p pd=12.52u as=5.28p ps=24.88u w=11.999999u l=0.7u
X75 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_cms_smt_0.nmos_6p0_CDNS_4066195314540_0.S.t6 GF_NI_IN_C_BASE_0.comp018green_esd_cdm_0.IP_IN.t2 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_cms_smt_0.nmos_6p0_CDNS_4066195314537_0.D.t6 DVSS.t15 nfet_06v0 ad=1.166p pd=6.18u as=0.689p ps=3.17u w=2.65u l=0.7u
X76 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_drv_0.A.t6 GF_NI_IN_C_BASE_0.comp018green_esd_cdm_0.IP_IN.t3 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_cms_smt_0.nmos_6p0_CDNS_4066195314540_0.S.t2 DVSS.t10 nfet_06v0 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.7u
X77 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_drv_0.A.t3 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_1.Z.t6 DVDD.t73 DVDD.t72 pfet_06v0 ad=0.88p pd=4.88u as=0.52p ps=2.52u w=2u l=0.7u
X78 GF_NI_IN_C_BASE_0.ndrive_x_<3>.t0 GF_NI_IN_C_BASE_0.comp018green_out_predrv_1.nmos_6p0_CDNS_4066195314519_2.S.t3 DVSS.t123 DVSS.t122 nfet_06v0 ad=1.56p pd=6.52u as=1.56p ps=6.52u w=6u l=0.7u
X79 DVSS GF_NI_IN_C_BASE_0.ndrive_y_<0>.t5 PAD DVSS.t60 nfet_06v0_dss d_sab=0.28u s_sab=3.78u ad=10.639999p pd=76.56u as=0.14364n ps=83.56u w=38u l=1.15u
X80 DVSS.t125 GF_NI_IN_C_BASE_0.comp018green_out_predrv_1.nmos_6p0_CDNS_4066195314519_2.S.t4 GF_NI_IN_C_BASE_0.ndrive_Y_<3>.t0 DVSS.t124 nfet_06v0 ad=1.56p pd=6.52u as=1.56p ps=6.52u w=6u l=0.7u
X81 DVSS.t1 GF_NI_IN_C_BASE_0.comp018green_out_predrv_1.nmos_6p0_CDNS_4066195314519_0.D.t5 GF_NI_IN_C_BASE_0.pdrive_y_<3>.t2 DVSS.t0 nfet_06v0 ad=1.56p pd=6.52u as=1.56p ps=6.52u w=6u l=0.7u
X82 DVSS.t194 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_3.nmos_6p0_CDNS_4066195314530_0.D.t2 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_3.Z.t0 DVSS.t193 nfet_06v0 ad=0.66p pd=3.88u as=0.39p ps=2.02u w=1.5u l=0.7u
X83 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_3.Z GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_3.nmos_6p0_CDNS_4066195314530_0.D.t3 DVDD.t77 DVDD.t76 pfet_06v0 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.7u
X84 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_pupd_0.PD.t1 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_0.Z.t3 DVDD.t135 DVDD.t134 pfet_06v0 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.7u
D2 VSS.t51 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.t5 diode_pd2nw_06v0 pj=1.92u area=0.2304p
X85 PAD GF_NI_IN_C_BASE_0.pdrive_x_<3>.t4 DVDD DVDD.t140 pfet_06v0_dss d_sab=2.78u s_sab=0.28u ad=0.1112n pd=85.56u as=11.199999p ps=80.56u w=40u l=0.7u
X86 DVSS.t39 GF_NI_IN_C_BASE_0.comp018green_out_predrv_2.nmos_6p0_CDNS_4066195314519_2.S.t3 GF_NI_IN_C_BASE_0.ndrive_y_<2>.t3 DVSS.t38 nfet_06v0 ad=1.56p pd=6.52u as=1.56p ps=6.52u w=6u l=0.7u
X87 DVDD.t119 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_3.Z.t3 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_3.ZB.t1 DVDD.t118 pfet_06v0 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.7u
X88 DVDD.t181 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_0.nmos_6p0_CDNS_4066195314530_0.D.t3 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_0.Z.t1 DVDD.t180 pfet_06v0 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.7u
X89 GF_NI_IN_C_BASE_0.comp018green_out_predrv_0.nmos_6p0_CDNS_4066195314519_2.S.t1 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.ENB.t2 GF_NI_IN_C_BASE_0.comp018green_out_predrv_0.nmos_6p0_CDNS_4066195314519_0.D.t1 DVDD.t128 pfet_06v0 ad=3.12p pd=12.52u as=5.28p ps=24.88u w=11.999999u l=0.7u
X90 VDD.t43 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_drv_0.Z.t2 Y.t11 VDD.t42 pfet_06v0 ad=0.91p pd=4.02u as=0.91p ps=4.02u w=3.5u l=0.7u
X91 Y.t10 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_drv_0.Z.t3 VDD.t45 VDD.t44 pfet_06v0 ad=0.91p pd=4.02u as=1.54p ps=7.88u w=3.5u l=0.7u
X92 DVDD.t206 DVSS.t59 cap_nmos_06v0 c_width=5u c_length=1.5u
X93 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_cms_smt_0.nmos_6p0_CDNS_4066195314530_0.D.t0 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_cms_smt_0.nmos_6p0_CDNS_4066195314535_0.D.t2 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_drv_0.A.t0 DVDD.t60 pfet_06v0 ad=0.88p pd=4.88u as=0.88p ps=4.88u w=2u l=0.7u
D3 DVSS.t14 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_pupd_0.ppolyf_u_CDNS_4066195314532_0.PLUS diode_nd2ps_06v0 pj=42u area=20p
X94 DVSS.t159 GF_NI_IN_C_BASE_0.comp018green_sigbuf_1_0.nmos_6p0_CDNS_4066195314530_0.D.t2 GF_NI_IN_C_BASE_0.comp018green_out_predrv_0.SL.t0 DVSS.t158 nfet_06v0 ad=0.39p pd=2.02u as=0.39p ps=2.02u w=1.5u l=0.7u
X95 GF_NI_IN_C_BASE_0.pdrive_y_<1>.t2 GF_NI_IN_C_BASE_0.comp018green_out_predrv_3.nmos_6p0_CDNS_4066195314519_0.D.t5 DVSS.t180 DVSS.t179 nfet_06v0 ad=1.56p pd=6.52u as=2.64p ps=12.879999u w=6u l=0.7u
X96 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_cms_smt_0.nmos_6p0_CDNS_4066195314537_0.D.t5 GF_NI_IN_C_BASE_0.comp018green_esd_cdm_0.IP_IN.t4 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_cms_smt_0.nmos_6p0_CDNS_4066195314540_0.S.t5 DVSS.t3 nfet_06v0 ad=0.689p pd=3.17u as=1.166p ps=6.18u w=2.65u l=0.7u
X97 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_pupd_0.ppolyf_u_CDNS_4066195314533_1.PLUS.t1 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_pupd_0.ppolyf_u_CDNS_4066195314533_2.PLUS.t0 DVDD.t40 ppolyf_u r_width=0.8u r_length=35.7u
X98 VSS.t19 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_drv_0.Z.t4 Y.t4 VSS.t18 nfet_06v0 ad=0.39p pd=2.02u as=0.39p ps=2.02u w=1.5u l=0.7u
X99 VSS.t27 PU.t5 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_logic_pupd_0.comp018green_std_xor2_0.nmos_6p0_CDNS_4066195314530_2.D.t1 VSS.t26 nfet_06v0 ad=0.66p pd=3.88u as=0.66p ps=3.88u w=1.5u l=0.7u
X100 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_pupd_0.ppolyf_u_CDNS_4066195314533_5.MINUS.t0 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_pupd_0.PU_B.t2 DVDD.t91 DVDD.t90 pfet_06v0 ad=1.32p pd=6.88u as=1.32p ps=6.88u w=3u l=0.7u
X101 DVSS.t172 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_a_0.nmos_6p0_CDNS_4066195314511_3.S.t2 GF_NI_IN_C_BASE_0.comp018green_out_predrv_0.A.t0 DVSS.t171 nfet_06v0 ad=0.78p pd=3.52u as=1.32p ps=6.88u w=3u l=0.7u
X102 GF_NI_IN_C_BASE_0.ndrive_x_<1>.t2 GF_NI_IN_C_BASE_0.comp018green_out_predrv_0.SL.t5 GF_NI_IN_C_BASE_0.ndrive_Y_<1>.t2 DVDD.t54 pfet_06v0 ad=3.12p pd=12.52u as=5.28p ps=24.88u w=11.999999u l=0.7u
X103 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_3.ZB.t0 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_3.Z.t4 DVSS.t149 DVSS.t148 nfet_06v0 ad=0.39p pd=2.02u as=0.66p ps=3.88u w=1.5u l=0.7u
X104 DVSS.t77 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_cms_smt_0.nmos_6p0_CDNS_4066195314535_0.D.t3 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_cms_smt_0.nmos_6p0_CDNS_4066195314530_0.D.t1 DVSS.t76 nfet_06v0 ad=0.66p pd=3.88u as=0.66p ps=3.88u w=1.5u l=0.7u
X105 DVSS.t127 GF_NI_IN_C_BASE_0.comp018green_out_predrv_0.nmos_6p0_CDNS_4066195314519_0.D.t5 GF_NI_IN_C_BASE_0.pdrive_y_<0>.t2 DVSS.t126 nfet_06v0 ad=2.64p pd=12.879999u as=1.56p ps=6.52u w=6u l=0.7u
X106 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_pupd_0.PU_B.t0 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_2.nmos_6p0_CDNS_4066195314530_0.D.t3 DVSS.t145 DVSS.t144 nfet_06v0 ad=0.39p pd=2.02u as=0.39p ps=2.02u w=1.5u l=0.7u
X107 Y.t3 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_drv_0.Z.t5 VSS.t21 VSS.t20 nfet_06v0 ad=0.39p pd=2.02u as=0.66p ps=3.88u w=1.5u l=0.7u
X108 DVDD.t174 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_a_0.nmos_6p0_CDNS_4066195314511_3.S.t3 GF_NI_IN_C_BASE_0.comp018green_out_predrv_0.A.t1 DVDD.t173 pfet_06v0 ad=1.56p pd=6.52u as=2.64p ps=12.879999u w=6u l=0.7u
X109 GF_NI_IN_C_BASE_0.pdrive_y_<0>.t2 GF_NI_IN_C_BASE_0.comp018green_out_predrv_0.nmos_6p0_CDNS_4066195314519_0.D.t6 DVSS.t129 DVSS.t128 nfet_06v0 ad=1.56p pd=6.52u as=1.56p ps=6.52u w=6u l=0.7u
X110 DVDD.t93 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_pupd_0.PU_B.t3 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_2.ZB.t1 DVDD.t92 pfet_06v0 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.7u
X111 GF_NI_IN_C_BASE_0.comp018green_out_predrv_0.nmos_6p0_CDNS_4066195314519_2.S GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.EN.t2 GF_NI_IN_C_BASE_0.comp018green_out_predrv_0.nmos_6p0_CDNS_4066195314519_0.D.t2 DVSS.t164 nfet_06v0 ad=2.64p pd=12.879999u as=1.56p ps=6.52u w=6u l=0.7u
X112 GF_NI_IN_C_BASE_0.pdrive_y_<2>.t3 GF_NI_IN_C_BASE_0.comp018green_out_predrv_2.nmos_6p0_CDNS_4066195314519_0.D.t4 DVDD.t106 DVDD.t105 pfet_06v0 ad=3.12p pd=12.52u as=5.28p ps=24.88u w=11.999999u l=0.7u
X113 GF_NI_IN_C_BASE_0.pdrive_y_<3>.t1 DVDD.t207 GF_NI_IN_C_BASE_0.pdrive_x_<3>.t2 DVSS.t32 nfet_06v0 ad=0.528p pd=3.28u as=0.528p ps=3.28u w=1.2u l=0.7u
X114 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_2.ZB.t1 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_pupd_0.PU_B.t4 DVDD.t95 DVDD.t94 pfet_06v0 ad=0.78p pd=3.52u as=1.32p ps=6.88u w=3u l=0.7u
X115 DVSS.t45 GF_NI_IN_C_BASE_0.comp018green_out_predrv_0.SL.t6 GF_NI_IN_C_BASE_0.comp018green_out_predrv_0.SLB.t1 DVSS.t44 nfet_06v0 ad=0.66p pd=3.88u as=0.39p ps=2.02u w=1.5u l=0.7u
X116 PAD GF_NI_IN_C_BASE_0.pdrive_y_<2>.t4 DVDD DVDD.t148 pfet_06v0_dss d_sab=2.78u s_sab=0.28u ad=0.1112n pd=85.56u as=11.199999p ps=80.56u w=40u l=0.7u
X117 GF_NI_IN_C_BASE_0.pdrive_x_<3>.t1 GF_NI_IN_C_BASE_0.comp018green_out_predrv_0.SLB.t4 GF_NI_IN_C_BASE_0.pdrive_y_<3>.t0 DVSS.t33 nfet_06v0 ad=2.64p pd=12.879999u as=1.56p ps=6.52u w=6u l=0.7u
X118 DVDD.t208 DVSS.t58 cap_nmos_06v0 c_width=5u c_length=1.5u
X119 DVDD.t209 DVSS.t57 cap_nmos_06v0 c_width=3u c_length=3u
X120 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_2.nmos_6p0_CDNS_4066195314511_1.S.t0 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.t17 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_2.nmos_6p0_CDNS_4066195314511_0.S.t0 VSS.t7 nfet_06v0 ad=1.32p pd=6.88u as=0.78p ps=3.52u w=3u l=0.7u
X121 PAD GF_NI_IN_C_BASE_0.ndrive_x_<2>.t3 DVSS DVSS.t101 nfet_06v0_dss d_sab=3.78u s_sab=0.28u ad=0.14364n pd=83.56u as=10.639999p ps=76.56u w=38u l=1.15u
X122 DVDD.t210 DVSS.t56 cap_nmos_06v0 c_width=5u c_length=1.5u
X123 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_1.Z.t0 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_1.nmos_6p0_CDNS_4066195314530_0.D.t3 DVSS.t88 DVSS.t87 nfet_06v0 ad=0.39p pd=2.02u as=0.66p ps=3.88u w=1.5u l=0.7u
X124 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_2.nmos_6p0_CDNS_4066195314511_0.S.t1 VDD.t68 VSS.t1 VSS.t0 nfet_06v0 ad=0.78p pd=3.52u as=1.32p ps=6.88u w=3u l=0.7u
X125 GF_NI_IN_C_BASE_0.pdrive_y_<3>.t0 GF_NI_IN_C_BASE_0.comp018green_out_predrv_0.SLB.t5 GF_NI_IN_C_BASE_0.pdrive_x_<3>.t0 DVSS.t32 nfet_06v0 ad=1.56p pd=6.52u as=2.64p ps=12.879999u w=6u l=0.7u
X126 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_cms_smt_0.nmos_6p0_CDNS_4066195314537_0.D.t1 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_1.Z.t7 DVSS.t90 DVSS.t89 nfet_06v0 ad=1.408p pd=7.28u as=0.832p ps=3.72u w=3.2u l=0.7u
X127 a_5575_62984.t1 GF_NI_IN_C_BASE_0.comp018green_esd_cdm_0.IP_IN.t5 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_drv_0.A.t7 DVDD.t4 pfet_06v0 ad=0.946p pd=5.18u as=0.559p ps=2.67u w=2.15u l=0.7u
X128 DVSS.t73 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_1.EN.t4 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_1.ENB.t0 DVSS.t72 nfet_06v0 ad=0.78p pd=3.52u as=1.32p ps=6.88u w=3u l=0.7u
D4 VSS.t52 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.t4 diode_pd2nw_06v0 pj=1.92u area=0.2304p
D5 VSS.t53 VDD.t39 diode_pd2nw_06v0 pj=1.92u area=0.2304p
X129 GF_NI_IN_C_BASE_0.ndrive_x_<2>.t0 GF_NI_IN_C_BASE_0.comp018green_out_predrv_0.SL.t7 GF_NI_IN_C_BASE_0.ndrive_y_<2>.t1 DVDD.t47 pfet_06v0 ad=3.12p pd=12.52u as=3.12p ps=12.52u w=11.999999u l=0.7u
X130 VSS.t43 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_logic_pupd_0.PUB_OUT.t2 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_2.nmos_6p0_CDNS_4066195314530_0.D.t0 VSS.t42 nfet_06v0 ad=0.66p pd=3.88u as=0.66p ps=3.88u w=1.5u l=0.7u
X131 DVDD.t66 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_1.EN.t5 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_1.ENB.t1 DVDD.t65 pfet_06v0 ad=1.56p pd=6.52u as=2.64p ps=12.879999u w=6u l=0.7u
X132 GF_NI_IN_C_BASE_0.ndrive_y_<2>.t0 DVSS.t205 GF_NI_IN_C_BASE_0.ndrive_x_<2>.t1 DVDD.t202 pfet_06v0 ad=0.528p pd=3.28u as=0.528p ps=3.28u w=1.2u l=0.7u
X133 GF_NI_IN_C_BASE_0.comp018green_esd_cdm_0.IP_IN.t0 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_pupd_0.ppolyf_u_CDNS_4066195314533_2.PLUS.t1 DVDD.t131 ppolyf_u r_width=0.8u r_length=22.999998u
X134 GF_NI_IN_C_BASE_0.pdrive_x_<0>.t3 GF_NI_IN_C_BASE_0.comp018green_out_predrv_0.nmos_6p0_CDNS_4066195314519_0.D.t7 DVDD.t133 DVDD.t132 pfet_06v0 ad=3.12p pd=12.52u as=3.12p ps=12.52u w=11.999999u l=0.7u
X135 DVDD.t211 DVSS.t55 cap_nmos_06v0 c_width=5u c_length=1.5u
X136 GF_NI_IN_C_BASE_0.comp018green_out_predrv_0.SL.t0 GF_NI_IN_C_BASE_0.comp018green_sigbuf_1_0.nmos_6p0_CDNS_4066195314530_0.D.t3 DVSS.t119 DVSS.t118 nfet_06v0 ad=0.39p pd=2.02u as=0.66p ps=3.88u w=1.5u l=0.7u
X137 DVDD.t212 DVSS.t54 cap_nmos_06v0 c_width=3u c_length=3u
X138 DVDD.t28 GF_NI_IN_C_BASE_0.comp018green_out_predrv_0.A.t5 GF_NI_IN_C_BASE_0.comp018green_out_predrv_3.nmos_6p0_CDNS_4066195314519_2.S.t1 DVDD.t27 pfet_06v0 ad=3.12p pd=12.52u as=5.28p ps=24.88u w=11.999999u l=0.7u
X139 DVDD GF_NI_IN_C_BASE_0.pdrive_y_<3>.t4 PAD DVDD.t96 pfet_06v0_dss d_sab=0.28u s_sab=2.78u ad=11.199999p pd=80.56u as=0.1112n ps=85.56u w=40u l=0.7u
X140 GF_NI_IN_C_BASE_0.ndrive_Y_<1>.t3 GF_NI_IN_C_BASE_0.comp018green_out_predrv_3.nmos_6p0_CDNS_4066195314519_2.S.t4 DVSS.t71 DVSS.t70 nfet_06v0 ad=1.56p pd=6.52u as=1.56p ps=6.52u w=6u l=0.7u
X141 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_drv_0.nmos_6p0_CDNS_4066195314550_0.D GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_drv_0.nmos_6p0_CDNS_4066195314547_0.S.t3 VDD.t29 VDD.t28 pfet_06v0 ad=0.65p pd=3.02u as=1.1p ps=5.88u w=2.5u l=0.7u
X142 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_logic_pupd_0.comp018green_std_xor2_0.nmos_6p0_CDNS_4066195314530_0.D.t0 PD.t0 VDD.t64 VDD.t63 pfet_06v0 ad=1.32p pd=6.88u as=1.32p ps=6.88u w=3u l=0.7u
D6 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.t18 VDD.t5 diode_pd2nw_06v0 pj=4u area=1p
X143 DVSS.t37 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_1.ENB.t2 GF_NI_IN_C_BASE_0.comp018green_out_predrv_3.nmos_6p0_CDNS_4066195314519_0.D.t0 DVSS.t36 nfet_06v0 ad=1.56p pd=6.52u as=1.56p ps=6.52u w=6u l=0.7u
X144 DVDD.t108 GF_NI_IN_C_BASE_0.comp018green_out_predrv_2.nmos_6p0_CDNS_4066195314519_0.D.t5 GF_NI_IN_C_BASE_0.pdrive_x_<2>.t3 DVDD.t107 pfet_06v0 ad=5.28p pd=24.88u as=3.12p ps=12.52u w=11.999999u l=0.7u
X145 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_1.nmos_6p0_CDNS_4066195314530_0.D.t1 GF_NI_IN_C_BASE_0.ppolyf_u_CDNS_4066195314551_0.MINUS.t1 VDD.t60 VDD.t59 pfet_06v0 ad=1.32p pd=6.88u as=1.32p ps=6.88u w=3u l=0.7u
X146 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.nmos_6p0_CDNS_4066195314511_1.S.t1 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.t19 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.nmos_6p0_CDNS_4066195314511_0.S.t1 VSS.t6 nfet_06v0 ad=1.32p pd=6.88u as=0.78p ps=3.52u w=3u l=0.7u
X147 DVDD.t154 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_3.Z.t5 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_cms_smt_0.nmos_6p0_CDNS_4066195314536_1.S.t2 DVDD.t153 pfet_06v0 ad=0.66p pd=3.88u as=0.39p ps=2.02u w=1.5u l=0.7u
X148 VDD.t25 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_drv_0.nmos_6p0_CDNS_4066195314547_0.S.t4 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_drv_0.nmos_6p0_CDNS_4066195314550_0.D VDD.t24 pfet_06v0 ad=1.1p pd=5.88u as=0.65p ps=3.02u w=2.5u l=0.7u
X149 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_pupd_0.ppolyf_u_CDNS_4066195314533_5.MINUS.t2 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_pupd_0.ppolyf_u_CDNS_4066195314533_4.PLUS.t1 DVDD.t40 ppolyf_u r_width=0.8u r_length=35.7u
X150 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_logic_pupd_0.comp018green_std_nand2_0.A.t0 PD.t1 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_logic_pupd_0.comp018green_std_xor2_0.nmos_6p0_CDNS_4066195314530_2.D.t2 VSS.t40 nfet_06v0 ad=0.66p pd=3.88u as=0.66p ps=3.88u w=1.5u l=0.7u
X151 GF_NI_IN_C_BASE_0.comp018green_out_predrv_1.nmos_6p0_CDNS_4066195314519_2.S.t1 GF_NI_IN_C_BASE_0.comp018green_out_predrv_1.EN.t2 DVDD.t192 DVDD.t191 pfet_06v0 ad=3.12p pd=12.52u as=3.12p ps=12.52u w=11.999999u l=0.7u
X152 DVDD.t35 GF_NI_IN_C_BASE_0.comp018green_out_predrv_1.nmos_6p0_CDNS_4066195314519_0.D.t6 GF_NI_IN_C_BASE_0.pdrive_y_<3>.t3 DVDD.t34 pfet_06v0 ad=5.28p pd=24.88u as=3.12p ps=12.52u w=11.999999u l=0.7u
X153 VDD.t4 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.t20 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_2.nmos_6p0_CDNS_4066195314511_1.S.t1 VDD.t3 pfet_06v0 ad=1.32p pd=6.88u as=0.78p ps=3.52u w=3u l=0.7u
X154 DVSS.t113 GF_NI_IN_C_BASE_0.comp018green_out_predrv_2.nmos_6p0_CDNS_4066195314519_0.D.t6 GF_NI_IN_C_BASE_0.pdrive_y_<2>.t2 DVSS.t112 nfet_06v0 ad=2.64p pd=12.879999u as=1.56p ps=6.52u w=6u l=0.7u
X155 GF_NI_IN_C_BASE_0.ndrive_y_<2>.t3 GF_NI_IN_C_BASE_0.comp018green_out_predrv_2.nmos_6p0_CDNS_4066195314519_2.S.t4 DVSS.t41 DVSS.t40 nfet_06v0 ad=1.56p pd=6.52u as=1.56p ps=6.52u w=6u l=0.7u
X156 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_2.nmos_6p0_CDNS_4066195314511_1.S.t1 VDD.t50 VDD.t52 VDD.t51 pfet_06v0 ad=0.78p pd=3.52u as=1.32p ps=6.88u w=3u l=0.7u
X157 GF_NI_IN_C_BASE_0.pdrive_y_<2>.t2 GF_NI_IN_C_BASE_0.comp018green_out_predrv_2.nmos_6p0_CDNS_4066195314519_0.D.t7 DVSS.t107 DVSS.t106 nfet_06v0 ad=1.56p pd=6.52u as=1.56p ps=6.52u w=6u l=0.7u
X158 DVDD.t196 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_1.nmos_6p0_CDNS_4066195314530_0.D.t4 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_1.Z.t1 DVDD.t195 pfet_06v0 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.7u
X159 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_cms_smt_0.nmos_6p0_CDNS_4066195314535_0.D.t0 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_3.Z.t6 DVSS.t151 DVSS.t150 nfet_06v0 ad=0.52p pd=2.52u as=0.88p ps=4.88u w=2u l=0.7u
X160 DVSS GF_NI_IN_C_BASE_0.ndrive_Y_<1>.t5 PAD DVSS.t78 nfet_06v0_dss d_sab=0.28u s_sab=3.78u ad=10.639999p pd=76.56u as=0.14364n ps=83.56u w=38u l=1.15u
X161 GF_NI_IN_C_BASE_0.ndrive_y_<0>.t2 GF_NI_IN_C_BASE_0.comp018green_out_predrv_0.nmos_6p0_CDNS_4066195314519_2.S.t4 DVDD.t125 DVDD.t124 pfet_06v0 ad=3.12p pd=12.52u as=3.12p ps=12.52u w=11.999999u l=0.7u
X162 GF_NI_IN_C_BASE_0.comp018green_out_predrv_2.nmos_6p0_CDNS_4066195314519_2.S GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_1.EN.t6 GF_NI_IN_C_BASE_0.comp018green_out_predrv_2.nmos_6p0_CDNS_4066195314519_0.D.t1 DVSS.t81 nfet_06v0 ad=2.64p pd=12.879999u as=1.56p ps=6.52u w=6u l=0.7u
D7 VSS.t54 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.t3 diode_pd2nw_06v0 pj=1.92u area=0.2304p
X163 VDD.t31 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_drv_0.Z.t6 Y.t9 VDD.t30 pfet_06v0 ad=0.91p pd=4.02u as=0.91p ps=4.02u w=3.5u l=0.7u
D8 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.t21 VDD.t5 diode_pd2nw_06v0 pj=4u area=1p
X164 GF_NI_IN_C_BASE_0.pdrive_y_<0>.t0 GF_NI_IN_C_BASE_0.comp018green_out_predrv_0.SLB.t6 GF_NI_IN_C_BASE_0.pdrive_x_<0>.t0 DVSS.t31 nfet_06v0 ad=1.56p pd=6.52u as=2.64p ps=12.879999u w=6u l=0.7u
X165 DVDD GF_NI_IN_C_BASE_0.pdrive_x_<1>.t4 PAD DVDD.t24 pfet_06v0_dss d_sab=0.28u s_sab=2.78u ad=11.199999p pd=80.56u as=0.1112n ps=85.56u w=40u l=0.7u
X166 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_cms_smt_0.nmos_6p0_CDNS_4066195314535_0.D.t1 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_3.Z.t7 DVDD.t152 DVDD.t151 pfet_06v0 ad=1.04p pd=4.52u as=1.76p ps=8.88u w=4u l=0.7u
X167 DVSS.t147 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_2.nmos_6p0_CDNS_4066195314511_1.S.t2 GF_NI_IN_C_BASE_0.comp018green_out_predrv_1.EN DVSS.t146 nfet_06v0 ad=0.78p pd=3.52u as=1.32p ps=6.88u w=3u l=0.7u
X168 DVSS.t22 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_drv_0.A.t11 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_drv_0.nmos_6p0_CDNS_4066195314547_0.S.t0 DVSS.t21 nfet_06v0 ad=1.04p pd=4.52u as=1.76p ps=8.88u w=4u l=0.7u
X169 DVDD.t213 DVSS.t53 cap_nmos_06v0 c_width=3u c_length=3u
X170 DVDD.t156 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_2.nmos_6p0_CDNS_4066195314511_1.S.t3 GF_NI_IN_C_BASE_0.comp018green_out_predrv_1.EN.t0 DVDD.t155 pfet_06v0 ad=1.56p pd=6.52u as=2.64p ps=12.879999u w=6u l=0.7u
X171 GF_NI_IN_C_BASE_0.comp018green_out_predrv_1.nmos_6p0_CDNS_4066195314519_0.D.t1 GF_NI_IN_C_BASE_0.comp018green_out_predrv_1.EN.t3 GF_NI_IN_C_BASE_0.comp018green_out_predrv_1.nmos_6p0_CDNS_4066195314519_2.S DVSS.t190 nfet_06v0 ad=1.56p pd=6.52u as=2.64p ps=12.879999u w=6u l=0.7u
X172 DVDD.t164 GF_NI_IN_C_BASE_0.comp018green_out_predrv_3.nmos_6p0_CDNS_4066195314519_0.D.t6 GF_NI_IN_C_BASE_0.pdrive_x_<1>.t3 DVDD.t163 pfet_06v0 ad=3.12p pd=12.52u as=3.12p ps=12.52u w=11.999999u l=0.7u
X173 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_0.nmos_6p0_CDNS_4066195314530_0.D.t0 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_logic_pupd_0.PDB_OUT.t2 VSS.t17 VSS.t16 nfet_06v0 ad=0.66p pd=3.88u as=0.66p ps=3.88u w=1.5u l=0.7u
X174 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_cms_smt_0.nmos_6p0_CDNS_4066195314530_0.D GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_3.Z.t8 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_drv_0.A.t8 DVSS.t139 nfet_06v0 ad=0.66p pd=3.88u as=0.66p ps=3.88u w=1.5u l=0.7u
X175 GF_NI_IN_C_BASE_0.comp018green_out_predrv_3.nmos_6p0_CDNS_4066195314519_0.D.t2 GF_NI_IN_C_BASE_0.comp018green_out_predrv_0.A.t6 DVSS.t9 DVSS.t8 nfet_06v0 ad=2.64p pd=12.879999u as=1.56p ps=6.52u w=6u l=0.7u
X176 GF_NI_IN_C_BASE_0.pdrive_x_<2>.t2 DVDD.t214 GF_NI_IN_C_BASE_0.pdrive_y_<2>.t1 DVSS.t30 nfet_06v0 ad=0.528p pd=3.28u as=0.528p ps=3.28u w=1.2u l=0.7u
X177 VSS.t23 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_drv_0.Z.t7 Y.t2 VSS.t22 nfet_06v0 ad=0.39p pd=2.02u as=0.39p ps=2.02u w=1.5u l=0.7u
X178 DVSS.t168 GF_NI_IN_C_BASE_0.comp018green_out_predrv_3.nmos_6p0_CDNS_4066195314519_0.D.t7 GF_NI_IN_C_BASE_0.pdrive_y_<1>.t2 DVSS.t167 nfet_06v0 ad=1.56p pd=6.52u as=1.56p ps=6.52u w=6u l=0.7u
X179 VDD.t33 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_drv_0.Z.t8 Y.t8 VDD.t32 pfet_06v0 ad=1.54p pd=7.88u as=0.91p ps=4.02u w=3.5u l=0.7u
X180 DVSS GF_NI_IN_C_BASE_0.ndrive_y_<2>.t5 PAD DVSS.t185 nfet_06v0_dss d_sab=0.28u s_sab=3.78u ad=10.639999p pd=76.56u as=0.14364n ps=83.56u w=38u l=1.15u
X181 GF_NI_IN_C_BASE_0.pdrive_x_<2>.t1 GF_NI_IN_C_BASE_0.comp018green_out_predrv_0.SLB.t7 GF_NI_IN_C_BASE_0.pdrive_y_<2>.t0 DVSS.t30 nfet_06v0 ad=2.64p pd=12.879999u as=1.56p ps=6.52u w=6u l=0.7u
X182 DVDD.t75 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_1.Z.t8 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_drv_0.A.t2 DVDD.t74 pfet_06v0 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=0.7u
X183 DVDD.t168 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_2.nmos_6p0_CDNS_4066195314530_0.D.t4 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_pupd_0.PU_B.t1 DVDD.t167 pfet_06v0 ad=1.32p pd=6.88u as=0.78p ps=3.52u w=3u l=0.7u
X184 DVDD.t121 GF_NI_IN_C_BASE_0.comp018green_sigbuf_1_0.nmos_6p0_CDNS_4066195314530_0.D.t4 GF_NI_IN_C_BASE_0.comp018green_out_predrv_0.SL.t1 DVDD.t120 pfet_06v0 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.7u
X185 GF_NI_IN_C_BASE_0.pdrive_y_<3>.t3 GF_NI_IN_C_BASE_0.comp018green_out_predrv_1.nmos_6p0_CDNS_4066195314519_0.D.t7 DVDD.t17 DVDD.t16 pfet_06v0 ad=3.12p pd=12.52u as=3.12p ps=12.52u w=11.999999u l=0.7u
D9 PU.t6 VDD.t0 diode_pd2nw_06v0 pj=4u area=1p
X186 DVSS.t92 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_1.Z.t9 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_1.ZB.t0 DVSS.t91 nfet_06v0 ad=0.66p pd=3.88u as=0.39p ps=2.02u w=1.5u l=0.7u
X187 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_0.Z.t1 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_0.nmos_6p0_CDNS_4066195314530_0.D.t4 DVDD.t179 DVDD.t178 pfet_06v0 ad=0.78p pd=3.52u as=1.32p ps=6.88u w=3u l=0.7u
X188 VSS.t39 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_logic_pupd_0.comp018green_std_nand2_0.A.t2 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_logic_pupd_0.comp018green_std_nand2_0.nmos_6p0_CDNS_4066195314511_0.D.t0 VSS.t38 nfet_06v0 ad=1.32p pd=6.88u as=0.78p ps=3.52u w=3u l=0.7u
X189 PU.t0 PD.t2 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_logic_pupd_0.comp018green_std_nand2_0.A.t1 VDD.t57 pfet_06v0 ad=1.32p pd=6.88u as=1.32p ps=6.88u w=3u l=0.7u
X190 GF_NI_IN_C_BASE_0.ndrive_Y_<3>.t1 GF_NI_IN_C_BASE_0.comp018green_out_predrv_1.nmos_6p0_CDNS_4066195314519_2.S.t5 DVDD.t130 DVDD.t129 pfet_06v0 ad=5.28p pd=24.88u as=3.12p ps=12.52u w=11.999999u l=0.7u
X191 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_1.ZB.t0 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_1.Z.t10 DVSS.t94 DVSS.t93 nfet_06v0 ad=0.39p pd=2.02u as=0.39p ps=2.02u w=1.5u l=0.7u
X192 VSS.t25 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_drv_0.Z.t9 Y.t1 VSS.t24 nfet_06v0 ad=0.66p pd=3.88u as=0.39p ps=2.02u w=1.5u l=0.7u
X193 VDD.t2 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.t22 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.nmos_6p0_CDNS_4066195314511_1.S.t0 VDD.t1 pfet_06v0 ad=1.32p pd=6.88u as=0.78p ps=3.52u w=3u l=0.7u
X194 VDD.t56 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_logic_pupd_0.comp018green_std_nand2_0.A.t3 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_logic_pupd_0.PDB_OUT.t0 VDD.t55 pfet_06v0 ad=1.32p pd=6.88u as=0.78p ps=3.52u w=3u l=0.7u
X195 DVDD.t137 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_0.Z.t4 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_pupd_0.PD.t1 DVDD.t136 pfet_06v0 ad=1.32p pd=6.88u as=0.78p ps=3.52u w=3u l=0.7u
X196 DVDD.t215 DVSS.t52 cap_nmos_06v0 c_width=3u c_length=3u
X197 VSS.t15 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.t23 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_3.nmos_6p0_CDNS_4066195314530_0.D.t0 VSS.t14 nfet_06v0 ad=0.66p pd=3.88u as=0.66p ps=3.88u w=1.5u l=0.7u
X198 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_pupd_0.ppolyf_u_CDNS_4066195314532_0.PLUS PAD.t21 w_4468_53312# ppolyf_u r_width=2.5u r_length=2.8u
X199 DVDD.t177 GF_NI_IN_C_BASE_0.comp018green_out_predrv_0.SL.t8 GF_NI_IN_C_BASE_0.comp018green_out_predrv_0.SLB.t0 DVDD.t176 pfet_06v0 ad=1.32p pd=6.88u as=0.78p ps=3.52u w=3u l=0.7u
X200 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.ENB.t1 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.EN.t3 DVSS.t166 DVSS.t165 nfet_06v0 ad=1.32p pd=6.88u as=0.78p ps=3.52u w=3u l=0.7u
X201 Y.t7 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_drv_0.Z.t10 VDD.t47 VDD.t46 pfet_06v0 ad=0.91p pd=4.02u as=0.91p ps=4.02u w=3.5u l=0.7u
X202 DVSS.t121 GF_NI_IN_C_BASE_0.comp018green_out_predrv_0.nmos_6p0_CDNS_4066195314519_2.S.t5 GF_NI_IN_C_BASE_0.ndrive_x_<0>.t2 DVSS.t120 nfet_06v0 ad=1.56p pd=6.52u as=1.56p ps=6.52u w=6u l=0.7u
X203 PAD GF_NI_IN_C_BASE_0.ndrive_x_<3>.t3 DVSS DVSS.t114 nfet_06v0_dss d_sab=3.78u s_sab=0.28u ad=0.14364n pd=83.56u as=10.639999p ps=76.56u w=38u l=1.15u
X204 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.ENB.t0 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.EN.t4 DVDD.t110 DVDD.t109 pfet_06v0 ad=2.64p pd=12.879999u as=1.56p ps=6.52u w=6u l=0.7u
X205 DVDD.t147 GF_NI_IN_C_BASE_0.comp018green_out_predrv_0.nmos_6p0_CDNS_4066195314519_0.D.t8 GF_NI_IN_C_BASE_0.pdrive_y_<0>.t3 DVDD.t146 pfet_06v0 ad=3.12p pd=12.52u as=3.12p ps=12.52u w=11.999999u l=0.7u
X206 DVSS.t96 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_1.Z.t11 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_cms_smt_0.nmos_6p0_CDNS_4066195314537_0.D.t0 DVSS.t95 nfet_06v0 ad=0.832p pd=3.72u as=0.832p ps=3.72u w=3.2u l=0.7u
X207 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_cms_smt_0.nmos_6p0_CDNS_4066195314540_0.S.t2 GF_NI_IN_C_BASE_0.comp018green_esd_cdm_0.IP_IN.t6 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_drv_0.A.t5 DVSS.t7 nfet_06v0 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.7u
X208 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_pupd_0.ppolyf_u_CDNS_4066195314533_3.MINUS.t0 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_pupd_0.ppolyf_u_CDNS_4066195314533_4.PLUS.t0 DVDD.t40 ppolyf_u r_width=0.8u r_length=35.7u
X209 GF_NI_IN_C_BASE_0.comp018green_out_predrv_0.SLB.t1 GF_NI_IN_C_BASE_0.comp018green_out_predrv_0.SL.t9 DVSS.t175 DVSS.t174 nfet_06v0 ad=0.39p pd=2.02u as=0.39p ps=2.02u w=1.5u l=0.7u
X210 GF_NI_IN_C_BASE_0.pdrive_y_<3>.t2 GF_NI_IN_C_BASE_0.comp018green_out_predrv_1.nmos_6p0_CDNS_4066195314519_0.D.t8 DVSS.t12 DVSS.t11 nfet_06v0 ad=1.56p pd=6.52u as=2.64p ps=12.879999u w=6u l=0.7u
X211 DVDD.t59 GF_NI_IN_C_BASE_0.comp018green_out_predrv_3.nmos_6p0_CDNS_4066195314519_2.S.t5 GF_NI_IN_C_BASE_0.ndrive_Y_<1>.t0 DVDD.t58 pfet_06v0 ad=3.12p pd=12.52u as=3.12p ps=12.52u w=11.999999u l=0.7u
X212 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_3.Z.t0 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_3.nmos_6p0_CDNS_4066195314530_0.D.t4 DVSS.t100 DVSS.t99 nfet_06v0 ad=0.39p pd=2.02u as=0.39p ps=2.02u w=1.5u l=0.7u
X213 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_pupd_0.PD.t0 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_0.Z.t5 DVSS.t136 DVSS.t135 nfet_06v0 ad=0.39p pd=2.02u as=0.39p ps=2.02u w=1.5u l=0.7u
X214 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_cms_smt_0.nmos_6p0_CDNS_4066195314537_0.D.t0 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_1.Z.t12 DVSS.t86 DVSS.t85 nfet_06v0 ad=0.832p pd=3.72u as=1.408p ps=7.28u w=3.2u l=0.7u
X215 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_drv_0.A.t5 GF_NI_IN_C_BASE_0.comp018green_esd_cdm_0.IP_IN.t7 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_cms_smt_0.nmos_6p0_CDNS_4066195314540_0.S.t1 DVSS.t13 nfet_06v0 ad=0.78p pd=3.52u as=1.32p ps=6.88u w=3u l=0.7u
D10 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_pupd_0.ppolyf_u_CDNS_4066195314532_0.PLUS DVDD diode_pd2nw_06v0 pj=42u area=20p
X216 GF_NI_IN_C_BASE_0.pdrive_x_<1>.t0 GF_NI_IN_C_BASE_0.comp018green_out_predrv_0.SLB.t8 GF_NI_IN_C_BASE_0.pdrive_y_<1>.t0 DVSS.t29 nfet_06v0 ad=2.64p pd=12.879999u as=1.56p ps=6.52u w=6u l=0.7u
X217 DVDD GF_NI_IN_C_BASE_0.pdrive_x_<0>.t5 PAD DVDD.t102 pfet_06v0_dss d_sab=0.28u s_sab=2.78u ad=11.199999p pd=80.56u as=0.1112n ps=85.56u w=40u l=0.7u
X218 GF_NI_IN_C_BASE_0.ndrive_x_<3>.t2 GF_NI_IN_C_BASE_0.comp018green_out_predrv_0.SL.t10 GF_NI_IN_C_BASE_0.ndrive_Y_<3>.t4 DVDD.t48 pfet_06v0 ad=3.12p pd=12.52u as=5.28p ps=24.88u w=11.999999u l=0.7u
X219 GF_NI_IN_C_BASE_0.ndrive_Y_<1>.t0 GF_NI_IN_C_BASE_0.comp018green_out_predrv_0.SL.t11 GF_NI_IN_C_BASE_0.ndrive_x_<1>.t2 DVDD.t49 pfet_06v0 ad=3.12p pd=12.52u as=3.12p ps=12.52u w=11.999999u l=0.7u
X220 Y.t0 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_drv_0.Z.t11 VSS.t36 VSS.t35 nfet_06v0 ad=0.39p pd=2.02u as=0.39p ps=2.02u w=1.5u l=0.7u
X221 GF_NI_IN_C_BASE_0.comp018green_out_predrv_0.nmos_6p0_CDNS_4066195314519_0.D.t2 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.ENB.t3 DVSS.t157 DVSS.t156 nfet_06v0 ad=1.56p pd=6.52u as=1.56p ps=6.52u w=6u l=0.7u
X222 DVSS.t141 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_3.Z.t9 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_3.ZB.t0 DVSS.t140 nfet_06v0 ad=0.39p pd=2.02u as=0.39p ps=2.02u w=1.5u l=0.7u
X223 DVSS.t177 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_0.nmos_6p0_CDNS_4066195314530_0.D.t5 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_0.Z.t0 DVSS.t176 nfet_06v0 ad=0.39p pd=2.02u as=0.39p ps=2.02u w=1.5u l=0.7u
X224 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_drv_0.A.t7 GF_NI_IN_C_BASE_0.comp018green_esd_cdm_0.IP_IN.t8 a_5575_62984.t0 DVDD.t13 pfet_06v0 ad=0.559p pd=2.67u as=0.946p ps=5.18u w=2.15u l=0.7u
X225 GF_NI_IN_C_BASE_0.comp018green_out_predrv_2.nmos_6p0_CDNS_4066195314519_2.S.t0 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_1.ENB.t3 GF_NI_IN_C_BASE_0.comp018green_out_predrv_2.nmos_6p0_CDNS_4066195314519_0.D.t0 DVDD.t50 pfet_06v0 ad=3.12p pd=12.52u as=5.28p ps=24.88u w=11.999999u l=0.7u
X226 GF_NI_IN_C_BASE_0.ndrive_x_<1>.t0 DVSS.t206 GF_NI_IN_C_BASE_0.ndrive_Y_<1>.t1 DVDD.t203 pfet_06v0 ad=0.528p pd=3.28u as=0.528p ps=3.28u w=1.2u l=0.7u
X227 GF_NI_IN_C_BASE_0.comp018green_out_predrv_0.SL.t1 GF_NI_IN_C_BASE_0.comp018green_sigbuf_1_0.nmos_6p0_CDNS_4066195314530_0.D.t5 DVDD.t123 DVDD.t122 pfet_06v0 ad=0.78p pd=3.52u as=1.32p ps=6.88u w=3u l=0.7u
X228 GF_NI_IN_C_BASE_0.ndrive_y_<2>.t1 GF_NI_IN_C_BASE_0.comp018green_out_predrv_2.nmos_6p0_CDNS_4066195314519_2.S.t5 DVDD.t42 DVDD.t41 pfet_06v0 ad=3.12p pd=12.52u as=3.12p ps=12.52u w=11.999999u l=0.7u
X229 DVDD.t127 GF_NI_IN_C_BASE_0.comp018green_out_predrv_0.nmos_6p0_CDNS_4066195314519_2.S.t6 GF_NI_IN_C_BASE_0.ndrive_y_<0>.t1 DVDD.t126 pfet_06v0 ad=3.12p pd=12.52u as=5.28p ps=24.88u w=11.999999u l=0.7u
X230 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_logic_pupd_0.comp018green_std_nand2_0.nmos_6p0_CDNS_4066195314511_0.D.t1 PD.t3 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_logic_pupd_0.PDB_OUT.t0 VSS.t41 nfet_06v0 ad=0.78p pd=3.52u as=1.32p ps=6.88u w=3u l=0.7u
D11 DVSS.t14 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_pupd_0.ppolyf_u_CDNS_4066195314532_0.PLUS diode_nd2ps_06v0 pj=42u area=20p
X231 PAD GF_NI_IN_C_BASE_0.pdrive_x_<1>.t5 DVDD DVDD.t21 pfet_06v0_dss d_sab=2.78u s_sab=0.28u ad=0.1112n pd=85.56u as=11.199999p ps=80.56u w=40u l=0.7u
X232 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_logic_pupd_0.PDB_OUT.t0 PD.t4 VDD.t41 VDD.t40 pfet_06v0 ad=0.78p pd=3.52u as=1.32p ps=6.88u w=3u l=0.7u
X233 DVSS.t201 GF_NI_IN_C_BASE_0.comp018green_out_predrv_1.nmos_6p0_CDNS_4066195314519_2.S.t6 GF_NI_IN_C_BASE_0.ndrive_x_<3>.t0 DVSS.t200 nfet_06v0 ad=2.64p pd=12.879999u as=1.56p ps=6.52u w=6u l=0.7u
X234 a_5575_62984.t3 GF_NI_IN_C_BASE_0.comp018green_esd_cdm_0.IP_IN.t9 DVDD.t12 DVDD.t11 pfet_06v0 ad=0.836p pd=4.68u as=0.494p ps=2.42u w=1.9u l=0.7u
X235 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_1.EN.t0 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_1.nmos_6p0_CDNS_4066195314511_1.S.t2 DVSS.t84 DVSS.t83 nfet_06v0 ad=1.32p pd=6.88u as=0.78p ps=3.52u w=3u l=0.7u
X236 DVDD.t79 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_3.nmos_6p0_CDNS_4066195314530_0.D.t5 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_3.Z DVDD.t78 pfet_06v0 ad=1.32p pd=6.88u as=0.78p ps=3.52u w=3u l=0.7u
X237 DVSS.t109 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_pupd_0.PU_B.t5 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_2.ZB.t0 DVSS.t108 nfet_06v0 ad=0.39p pd=2.02u as=0.39p ps=2.02u w=1.5u l=0.7u
X238 DVDD.t10 GF_NI_IN_C_BASE_0.comp018green_esd_cdm_0.IP_IN.t10 a_5575_62984.t2 DVDD.t9 pfet_06v0 ad=0.494p pd=2.42u as=0.836p ps=4.68u w=1.9u l=0.7u
X239 DVSS.t199 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.nmos_6p0_CDNS_4066195314511_1.S.t2 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.EN.t0 DVSS.t198 nfet_06v0 ad=0.78p pd=3.52u as=1.32p ps=6.88u w=3u l=0.7u
D12 VSS.t55 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.t2 diode_pd2nw_06v0 pj=1.92u area=0.2304p
X240 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_2.ZB.t0 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_pupd_0.PU_B.t6 DVSS.t111 DVSS.t110 nfet_06v0 ad=0.39p pd=2.02u as=0.66p ps=3.88u w=1.5u l=0.7u
X241 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_logic_pupd_0.comp018green_std_xor2_0.nmos_6p0_CDNS_4066195314530_0.D.t0 PD.t5 VSS.t32 VSS.t31 nfet_06v0 ad=0.66p pd=3.88u as=0.66p ps=3.88u w=1.5u l=0.7u
X242 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_pupd_0.ppolyf_u_CDNS_4066195314532_0.PLUS PAD.t4 w_4468_53312# ppolyf_u r_width=2.5u r_length=2.8u
X243 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_1.EN.t1 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_1.nmos_6p0_CDNS_4066195314511_1.S.t3 DVDD.t69 DVDD.t68 pfet_06v0 ad=2.64p pd=12.879999u as=1.56p ps=6.52u w=6u l=0.7u
X244 GF_NI_IN_C_BASE_0.comp018green_out_predrv_0.nmos_6p0_CDNS_4066195314519_2.S.t0 GF_NI_IN_C_BASE_0.comp018green_out_predrv_0.A.t7 DVDD.t20 DVDD.t19 pfet_06v0 ad=5.28p pd=24.88u as=3.12p ps=12.52u w=11.999999u l=0.7u
X245 DVDD.t200 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.nmos_6p0_CDNS_4066195314511_1.S.t3 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.EN.t1 DVDD.t199 pfet_06v0 ad=1.56p pd=6.52u as=2.64p ps=12.879999u w=6u l=0.7u
X246 GF_NI_IN_C_BASE_0.pdrive_x_<2>.t3 GF_NI_IN_C_BASE_0.comp018green_out_predrv_2.nmos_6p0_CDNS_4066195314519_0.D.t8 DVDD.t87 DVDD.t86 pfet_06v0 ad=3.12p pd=12.52u as=3.12p ps=12.52u w=11.999999u l=0.7u
X247 DVDD.t112 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.EN.t5 GF_NI_IN_C_BASE_0.comp018green_out_predrv_0.nmos_6p0_CDNS_4066195314519_2.S.t1 DVDD.t111 pfet_06v0 ad=3.12p pd=12.52u as=3.12p ps=12.52u w=11.999999u l=0.7u
X248 DVSS.t105 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_3.Z.t10 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_cms_smt_0.nmos_6p0_CDNS_4066195314535_0.D.t0 DVSS.t104 nfet_06v0 ad=0.88p pd=4.88u as=0.52p ps=2.52u w=2u l=0.7u
X249 DVDD.t216 DVSS.t51 cap_nmos_06v0 c_width=5u c_length=1.5u
X250 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_drv_0.A.t1 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_cms_smt_0.nmos_6p0_CDNS_4066195314535_0.D.t4 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_cms_smt_0.nmos_6p0_CDNS_4066195314536_1.S.t0 DVDD.t67 pfet_06v0 ad=0.88p pd=4.88u as=0.88p ps=4.88u w=2u l=0.7u
X251 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_pupd_0.ppolyf_u_CDNS_4066195314533_5.MINUS.t1 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_pupd_0.PD.t2 DVSS.t138 DVSS.t137 nfet_06v0 ad=0.66p pd=3.88u as=0.66p ps=3.88u w=1.5u l=0.7u
X252 GF_NI_IN_C_BASE_0.comp018green_out_predrv_3.nmos_6p0_CDNS_4066195314519_0.D.t1 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_1.ENB.t4 GF_NI_IN_C_BASE_0.comp018green_out_predrv_3.nmos_6p0_CDNS_4066195314519_2.S.t0 DVDD.t51 pfet_06v0 ad=5.28p pd=24.88u as=3.12p ps=12.52u w=11.999999u l=0.7u
X253 VDD.t62 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_logic_pupd_0.PUB_OUT.t3 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_2.nmos_6p0_CDNS_4066195314530_0.D.t1 VDD.t61 pfet_06v0 ad=1.32p pd=6.88u as=1.32p ps=6.88u w=3u l=0.7u
X254 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_cms_smt_0.nmos_6p0_CDNS_4066195314537_0.D.t4 GF_NI_IN_C_BASE_0.comp018green_esd_cdm_0.IP_IN.t11 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_cms_smt_0.nmos_6p0_CDNS_4066195314540_0.S.t4 DVSS.t4 nfet_06v0 ad=0.689p pd=3.17u as=0.689p ps=3.17u w=2.65u l=0.7u
X255 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.nmos_6p0_CDNS_4066195314511_0.S.t0 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.t24 VSS.t5 VSS.t4 nfet_06v0 ad=0.78p pd=3.52u as=1.32p ps=6.88u w=3u l=0.7u
X256 DVDD.t3 GF_NI_IN_C_BASE_0.comp018green_out_predrv_0.A.t8 GF_NI_IN_C_BASE_0.comp018green_out_predrv_1.nmos_6p0_CDNS_4066195314519_2.S.t0 DVDD.t2 pfet_06v0 ad=3.12p pd=12.52u as=5.28p ps=24.88u w=11.999999u l=0.7u
X257 GF_NI_IN_C_BASE_0.pdrive_x_<1>.t3 GF_NI_IN_C_BASE_0.comp018green_out_predrv_3.nmos_6p0_CDNS_4066195314519_0.D.t8 DVDD.t166 DVDD.t165 pfet_06v0 ad=3.12p pd=12.52u as=5.28p ps=24.88u w=11.999999u l=0.7u
X258 GF_NI_IN_C_BASE_0.ndrive_x_<1>.t1 GF_NI_IN_C_BASE_0.comp018green_out_predrv_3.nmos_6p0_CDNS_4066195314519_2.S.t6 DVSS.t65 DVSS.t64 nfet_06v0 ad=1.56p pd=6.52u as=1.56p ps=6.52u w=6u l=0.7u
D13 PD.t6 VDD.t58 diode_pd2nw_06v0 pj=4u area=1p
X259 DVDD.t83 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_3.Z.t11 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_cms_smt_0.nmos_6p0_CDNS_4066195314535_0.D.t1 DVDD.t82 pfet_06v0 ad=1.76p pd=8.88u as=1.04p ps=4.52u w=4u l=0.7u
X260 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_drv_0.nmos_6p0_CDNS_4066195314550_0.D GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_drv_0.nmos_6p0_CDNS_4066195314547_0.S.t5 VDD.t27 VDD.t26 pfet_06v0 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.7u
X261 DVDD GF_NI_IN_C_BASE_0.pdrive_y_<1>.t4 PAD DVDD.t31 pfet_06v0_dss d_sab=0.28u s_sab=2.78u ad=11.199999p pd=80.56u as=0.1112n ps=85.56u w=40u l=0.7u
X262 GF_NI_IN_C_BASE_0.ndrive_Y_<3>.t0 GF_NI_IN_C_BASE_0.comp018green_out_predrv_1.nmos_6p0_CDNS_4066195314519_2.S.t7 DVSS.t203 DVSS.t202 nfet_06v0 ad=1.56p pd=6.52u as=1.56p ps=6.52u w=6u l=0.7u
D14 VSS.t56 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.t1 diode_pd2nw_06v0 pj=1.92u area=0.2304p
X263 DVSS.t67 GF_NI_IN_C_BASE_0.comp018green_out_predrv_3.nmos_6p0_CDNS_4066195314519_2.S.t7 GF_NI_IN_C_BASE_0.ndrive_Y_<1>.t3 DVSS.t66 nfet_06v0 ad=1.56p pd=6.52u as=1.56p ps=6.52u w=6u l=0.7u
X264 VDD.t67 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_drv_0.nmos_6p0_CDNS_4066195314547_0.S.t6 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_drv_0.nmos_6p0_CDNS_4066195314550_0.D VDD.t66 pfet_06v0 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.7u
X265 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_a_0.nmos_6p0_CDNS_4066195314511_3.S.t0 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_a_0.nmos_6p0_CDNS_4066195314511_1.D.t2 DVSS.t43 DVSS.t42 nfet_06v0 ad=1.32p pd=6.88u as=0.78p ps=3.52u w=3u l=0.7u
X266 DVDD.t44 GF_NI_IN_C_BASE_0.comp018green_out_predrv_2.nmos_6p0_CDNS_4066195314519_2.S.t6 GF_NI_IN_C_BASE_0.ndrive_y_<2>.t4 DVDD.t43 pfet_06v0 ad=3.12p pd=12.52u as=5.28p ps=24.88u w=11.999999u l=0.7u
X267 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_3.ZB.t1 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_3.Z.t12 DVDD.t85 DVDD.t84 pfet_06v0 ad=0.78p pd=3.52u as=1.32p ps=6.88u w=3u l=0.7u
X268 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_a_0.nmos_6p0_CDNS_4066195314511_3.S.t1 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_a_0.nmos_6p0_CDNS_4066195314511_1.D.t3 DVDD.t46 DVDD.t45 pfet_06v0 ad=2.64p pd=12.879999u as=1.56p ps=6.52u w=6u l=0.7u
X269 DVSS.t75 GF_NI_IN_C_BASE_0.comp018green_out_predrv_2.nmos_6p0_CDNS_4066195314519_2.S.t7 GF_NI_IN_C_BASE_0.ndrive_x_<2>.t2 DVSS.t74 nfet_06v0 ad=1.56p pd=6.52u as=1.56p ps=6.52u w=6u l=0.7u
X270 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_pupd_0.PU_B.t1 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_2.nmos_6p0_CDNS_4066195314530_0.D.t5 DVDD.t89 DVDD.t88 pfet_06v0 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.7u
X271 GF_NI_IN_C_BASE_0.comp018green_sigbuf_1_0.nmos_6p0_CDNS_4066195314530_0.D.t0 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.t25 VSS.t3 VSS.t2 nfet_06v0 ad=0.66p pd=3.88u as=0.66p ps=3.88u w=1.5u l=0.7u
X272 GF_NI_IN_C_BASE_0.ndrive_x_<0>.t2 GF_NI_IN_C_BASE_0.comp018green_out_predrv_0.nmos_6p0_CDNS_4066195314519_2.S.t7 DVSS.t98 DVSS.t97 nfet_06v0 ad=1.56p pd=6.52u as=2.64p ps=12.879999u w=6u l=0.7u
X273 DVDD.t217 DVSS.t50 cap_nmos_06v0 c_width=5u c_length=1.5u
D15 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.t26 VDD.t0 diode_pd2nw_06v0 pj=4u area=1p
X274 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_logic_pupd_0.comp018green_std_nand2_1.nmos_6p0_CDNS_4066195314511_0.D.t1 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_logic_pupd_0.comp018green_std_nand2_0.A.t4 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_logic_pupd_0.PUB_OUT.t1 VSS.t37 nfet_06v0 ad=0.78p pd=3.52u as=1.32p ps=6.88u w=3u l=0.7u
X275 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_1.Z.t1 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_1.nmos_6p0_CDNS_4066195314530_0.D.t5 DVDD.t62 DVDD.t61 pfet_06v0 ad=0.78p pd=3.52u as=1.32p ps=6.88u w=3u l=0.7u
X276 VSS.t48 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_drv_0.nmos_6p0_CDNS_4066195314547_0.S.t7 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_drv_0.Z.t0 VSS.t47 nfet_06v0 ad=0.55p pd=3.38u as=0.325p ps=1.77u w=1.25u l=0.7u
X277 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_pupd_0.ppolyf_u_CDNS_4066195314533_3.MINUS.t1 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_pupd_0.ppolyf_u_CDNS_4066195314533_0.MINUS.t1 DVDD.t40 ppolyf_u r_width=0.8u r_length=35.7u
X278 GF_NI_IN_C_BASE_0.comp018green_out_predrv_2.nmos_6p0_CDNS_4066195314519_0.D.t1 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_1.ENB.t5 DVSS.t47 DVSS.t46 nfet_06v0 ad=1.56p pd=6.52u as=1.56p ps=6.52u w=6u l=0.7u
X279 DVDD GF_NI_IN_C_BASE_0.pdrive_x_<3>.t5 PAD DVDD.t143 pfet_06v0_dss d_sab=0.28u s_sab=2.78u ad=11.199999p pd=80.56u as=0.1112n ps=85.56u w=40u l=0.7u
X280 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_drv_0.Z.t0 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_drv_0.nmos_6p0_CDNS_4066195314547_0.S.t8 VSS.t50 VSS.t49 nfet_06v0 ad=0.325p pd=1.77u as=0.55p ps=3.38u w=1.25u l=0.7u
X281 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_logic_pupd_0.PUB_OUT.t0 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_logic_pupd_0.comp018green_std_nand2_0.A.t5 VDD.t54 VDD.t53 pfet_06v0 ad=0.78p pd=3.52u as=1.32p ps=6.88u w=3u l=0.7u
X282 GF_NI_IN_C_BASE_0.comp018green_out_predrv_3.nmos_6p0_CDNS_4066195314519_0.D.t0 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_1.EN.t7 GF_NI_IN_C_BASE_0.comp018green_out_predrv_3.nmos_6p0_CDNS_4066195314519_2.S DVSS.t82 nfet_06v0 ad=1.56p pd=6.52u as=2.64p ps=12.879999u w=6u l=0.7u
X283 GF_NI_IN_C_BASE_0.ndrive_y_<0>.t4 GF_NI_IN_C_BASE_0.comp018green_out_predrv_0.SL.t12 GF_NI_IN_C_BASE_0.ndrive_x_<0>.t0 DVDD.t36 pfet_06v0 ad=5.28p pd=24.88u as=3.12p ps=12.52u w=11.999999u l=0.7u
X284 DVSS.t18 GF_NI_IN_C_BASE_0.comp018green_out_predrv_0.A.t9 GF_NI_IN_C_BASE_0.comp018green_out_predrv_0.nmos_6p0_CDNS_4066195314519_0.D.t0 DVSS.t17 nfet_06v0 ad=1.56p pd=6.52u as=2.64p ps=12.879999u w=6u l=0.7u
X285 GF_NI_IN_C_BASE_0.ndrive_x_<0>.t0 GF_NI_IN_C_BASE_0.comp018green_out_predrv_0.SL.t13 GF_NI_IN_C_BASE_0.ndrive_y_<0>.t2 DVDD.t37 pfet_06v0 ad=3.12p pd=12.52u as=3.12p ps=12.52u w=11.999999u l=0.7u
X286 DVDD.t218 DVSS.t49 cap_nmos_06v0 c_width=5u c_length=1.5u
X287 Y.t6 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_drv_0.Z.t12 VDD.t49 VDD.t48 pfet_06v0 ad=0.91p pd=4.02u as=0.91p ps=4.02u w=3.5u l=0.7u
X288 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_pupd_0.ppolyf_u_CDNS_4066195314532_0.PLUS PAD.t6 w_4468_53312# ppolyf_u r_width=2.5u r_length=2.8u
X289 GF_NI_IN_C_BASE_0.pdrive_y_<1>.t1 DVDD.t219 GF_NI_IN_C_BASE_0.pdrive_x_<1>.t2 DVSS.t35 nfet_06v0 ad=0.528p pd=3.28u as=0.528p ps=3.28u w=1.2u l=0.7u
X290 GF_NI_IN_C_BASE_0.pdrive_y_<2>.t0 GF_NI_IN_C_BASE_0.comp018green_out_predrv_0.SLB.t9 GF_NI_IN_C_BASE_0.pdrive_x_<2>.t0 DVSS.t28 nfet_06v0 ad=1.56p pd=6.52u as=2.64p ps=12.879999u w=6u l=0.7u
X291 DVDD.t220 DVSS.t48 cap_nmos_06v0 c_width=5u c_length=1.5u
X292 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_cms_smt_0.nmos_6p0_CDNS_4066195314540_0.S.t4 GF_NI_IN_C_BASE_0.comp018green_esd_cdm_0.IP_IN.t12 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_cms_smt_0.nmos_6p0_CDNS_4066195314537_0.D.t3 DVSS.t2 nfet_06v0 ad=0.689p pd=3.17u as=0.689p ps=3.17u w=2.65u l=0.7u
X293 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_drv_0.A.t2 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_1.Z.t13 DVDD.t71 DVDD.t70 pfet_06v0 ad=0.52p pd=2.52u as=0.88p ps=4.88u w=2u l=0.7u
X294 GF_NI_IN_C_BASE_0.comp018green_out_predrv_1.ENB.t1 GF_NI_IN_C_BASE_0.comp018green_out_predrv_1.EN.t4 DVSS.t189 DVSS.t188 nfet_06v0 ad=1.32p pd=6.88u as=0.78p ps=3.52u w=3u l=0.7u
X295 GF_NI_IN_C_BASE_0.ndrive_y_<0>.t3 DVSS.t207 GF_NI_IN_C_BASE_0.ndrive_x_<0>.t1 DVDD.t204 pfet_06v0 ad=0.528p pd=3.28u as=0.528p ps=3.28u w=1.2u l=0.7u
X296 PAD GF_NI_IN_C_BASE_0.ndrive_x_<1>.t3 DVSS DVSS.t195 nfet_06v0_dss d_sab=3.78u s_sab=0.28u ad=0.14364n pd=83.56u as=10.639999p ps=76.56u w=38u l=1.15u
R0 GF_NI_IN_C_BASE_0.comp018green_out_predrv_1.EN GF_NI_IN_C_BASE_0.comp018green_out_predrv_1.EN.t2 82.1164
R1 GF_NI_IN_C_BASE_0.comp018green_out_predrv_1.EN.n0 GF_NI_IN_C_BASE_0.comp018green_out_predrv_1.EN.t1 44.3219
R2 GF_NI_IN_C_BASE_0.comp018green_out_predrv_1.EN GF_NI_IN_C_BASE_0.comp018green_out_predrv_1.EN.t3 42.2319
R3 GF_NI_IN_C_BASE_0.comp018green_out_predrv_1.EN.n0 GF_NI_IN_C_BASE_0.comp018green_out_predrv_1.EN.t4 28.0534
R4 GF_NI_IN_C_BASE_0.comp018green_out_predrv_1.EN GF_NI_IN_C_BASE_0.comp018green_out_predrv_1.EN.n0 4.00859
R5 GF_NI_IN_C_BASE_0.comp018green_out_predrv_1.EN GF_NI_IN_C_BASE_0.comp018green_out_predrv_1.EN.t0 1.33388
R6 DVDD.n1327 DVDD.n1326 13303.9
R7 DVDD.n1377 DVDD.n1327 13198.6
R8 DVDD.n1378 DVDD.n1326 10692.2
R9 DVDD.n1378 DVDD.n1377 10540.9
R10 DVDD.n3027 DVDD.t131 926.309
R11 DVDD.n4235 DVDD.t202 902.129
R12 DVDD.n4235 DVDD.t203 902.129
R13 DVDD.t116 DVDD.t82 746.523
R14 DVDD.t175 DVDD.t67 596.601
R15 DVDD.n1884 DVDD.t201 502.392
R16 DVDD.n4199 DVDD.t204 502.392
R17 DVDD.t11 DVDD.t13 482.226
R18 DVDD.t131 DVDD.t40 425.889
R19 DVDD.n3025 DVDD.n2077 359.661
R20 DVDD.t9 DVDD.t72 357.033
R21 DVDD.t60 DVDD.n2718 353.346
R22 DVDD.t70 DVDD.t153 349.305
R23 DVDD.t151 DVDD.n2790 309.892
R24 DVDD.t67 DVDD.t60 299.846
R25 DVDD.t4 DVDD.t182 299.846
R26 DVDD.n2792 DVDD.n2714 261.661
R27 DVDD.n2487 DVDD.t78 237.623
R28 DVDD.t61 DVDD.n2457 237.623
R29 DVDD.n2562 DVDD.t167 237.623
R30 DVDD.t178 DVDD.n2532 237.623
R31 DVDD.t84 DVDD.n2485 234.93
R32 DVDD.n2485 DVDD.t187 234.93
R33 DVDD.t94 DVDD.n2560 234.93
R34 DVDD.n2560 DVDD.t136 234.93
R35 DVDD.t176 DVDD.n3691 210.464
R36 DVDD.t193 DVDD.n1954 208.482
R37 DVDD.n1921 DVDD.t65 208.482
R38 DVDD.t109 DVDD.n1921 208.482
R39 DVDD.t122 DVDD.n3692 208.102
R40 DVDD.n1954 DVDD.t173 203.769
R41 DVDD.t78 DVDD.t76 188.564
R42 DVDD.t118 DVDD.t84 188.564
R43 DVDD.t189 DVDD.t187 188.564
R44 DVDD.t195 DVDD.t61 188.564
R45 DVDD.t167 DVDD.t88 188.564
R46 DVDD.t92 DVDD.t94 188.564
R47 DVDD.t134 DVDD.t136 188.564
R48 DVDD.t180 DVDD.t178 188.564
R49 DVDD.t182 DVDD.t175 188.564
R50 DVDD.t13 DVDD.t4 188.564
R51 DVDD.t72 DVDD.t74 188.564
R52 DVDD.t74 DVDD.t70 188.564
R53 DVDD.t153 DVDD.t116 188.564
R54 DVDD.t82 DVDD.t151 188.564
R55 DVDD.n2791 DVDD.t11 145.286
R56 DVDD.t38 DVDD.t176 143.698
R57 DVDD.t120 DVDD.t122 143.698
R58 DVDD.t48 DVDD.t18 139.505
R59 DVDD.t2 DVDD.t34 139.505
R60 DVDD.t105 DVDD.t5 139.505
R61 DVDD.t50 DVDD.t53 139.505
R62 DVDD.t54 DVDD.t51 139.505
R63 DVDD.t27 DVDD.t183 139.505
R64 DVDD.t19 DVDD.t171 139.505
R65 DVDD.t36 DVDD.t128 139.505
R66 DVDD.n2790 DVDD.n2789 122.816
R67 DVDD.n1885 DVDD.t129 121.04
R68 DVDD.n4200 DVDD.t126 121.04
R69 DVDD.n4236 DVDD.t0 120.725
R70 DVDD.n4236 DVDD.t107 120.725
R71 DVDD.t43 DVDD.n4235 120.725
R72 DVDD.n4235 DVDD.t56 120.725
R73 DVDD.t165 DVDD.n4234 120.725
R74 DVDD.n4234 DVDD.t169 120.725
R75 DVDD.n1372 DVDD.n1328 114.094
R76 DVDD.n1376 DVDD.n1328 113.204
R77 DVDD.t173 DVDD.n1953 108.52
R78 DVDD.t65 DVDD.n1920 103.829
R79 DVDD.n1922 DVDD.t109 103.829
R80 DVDD.n1956 DVDD.t193 103.829
R81 DVDD.n2770 DVDD.n2764 96.2887
R82 DVDD.n5485 DVDD.n260 96.0189
R83 DVDD.n5659 DVDD.n5500 95.6467
R84 DVDD.n2789 DVDD.n2719 95.5887
R85 DVDD.n2785 DVDD.n2719 95.5887
R86 DVDD.n2785 DVDD.n2784 95.5887
R87 DVDD.n2784 DVDD.n2779 95.5887
R88 DVDD.n2779 DVDD.n2778 95.5887
R89 DVDD.n2778 DVDD.n2742 95.5887
R90 DVDD.n2774 DVDD.n2742 95.5887
R91 DVDD.n2774 DVDD.n2773 95.5887
R92 DVDD.n2773 DVDD.n2772 95.5887
R93 DVDD.n2772 DVDD.n2771 95.5887
R94 DVDD.n2771 DVDD.n2770 95.5887
R95 DVDD.n2486 DVDD.t118 95.0546
R96 DVDD.n2458 DVDD.t189 95.0546
R97 DVDD.n2561 DVDD.t92 95.0546
R98 DVDD.n2533 DVDD.t134 95.0546
R99 DVDD.t76 DVDD.n2486 93.509
R100 DVDD.n2458 DVDD.t195 93.509
R101 DVDD.t88 DVDD.n2561 93.509
R102 DVDD.n2533 DVDD.t180 93.509
R103 DVDD.n3323 DVDD.n3315 87.5869
R104 DVDD.n3323 DVDD.n3238 87.546
R105 DVDD.t138 DVDD.t52 81.8248
R106 DVDD.t52 DVDD.t48 81.8248
R107 DVDD.t18 DVDD.t191 81.8248
R108 DVDD.t191 DVDD.t2 81.8248
R109 DVDD.t34 DVDD.t16 81.8248
R110 DVDD.t16 DVDD.t7 81.8248
R111 DVDD.t7 DVDD.t0 81.8248
R112 DVDD.t107 DVDD.t86 81.8248
R113 DVDD.t86 DVDD.t80 81.8248
R114 DVDD.t80 DVDD.t105 81.8248
R115 DVDD.t5 DVDD.t197 81.8248
R116 DVDD.t197 DVDD.t50 81.8248
R117 DVDD.t53 DVDD.t47 81.8248
R118 DVDD.t47 DVDD.t41 81.8248
R119 DVDD.t41 DVDD.t43 81.8248
R120 DVDD.t56 DVDD.t58 81.8248
R121 DVDD.t58 DVDD.t49 81.8248
R122 DVDD.t49 DVDD.t54 81.8248
R123 DVDD.t51 DVDD.t63 81.8248
R124 DVDD.t63 DVDD.t27 81.8248
R125 DVDD.t183 DVDD.t185 81.8248
R126 DVDD.t185 DVDD.t163 81.8248
R127 DVDD.t163 DVDD.t165 81.8248
R128 DVDD.t132 DVDD.t169 81.8248
R129 DVDD.t146 DVDD.t132 81.8248
R130 DVDD.t171 DVDD.t146 81.8248
R131 DVDD.t111 DVDD.t19 81.8248
R132 DVDD.t128 DVDD.t111 81.8248
R133 DVDD.t37 DVDD.t36 81.8248
R134 DVDD.t124 DVDD.t37 81.8248
R135 DVDD.n3693 DVDD.t120 73.0276
R136 DVDD.n3693 DVDD.t38 70.6719
R137 DVDD.n3383 DVDD.n3237 66.4038
R138 DVDD.n3337 DVDD.n3237 66.4007
R139 DVDD.n3319 DVDD.n3318 66.1618
R140 DVDD.n3331 DVDD.n3319 66.1584
R141 DVDD.n3323 DVDD.n3314 55.0525
R142 DVDD.n3323 DVDD.n3240 54.9859
R143 DVDD.n5490 DVDD.t143 52.7139
R144 DVDD.n5494 DVDD.t99 52.7139
R145 DVDD.n5492 DVDD.t160 52.4178
R146 DVDD.t24 DVDD.n5498 52.4178
R147 DVDD.n5491 DVDD.t96 51.3813
R148 DVDD.n5495 DVDD.t113 51.3813
R149 DVDD.t148 DVDD.n5491 51.0851
R150 DVDD.n5495 DVDD.t31 51.0851
R151 DVDD.n5492 DVDD.t157 50.0486
R152 DVDD.n5498 DVDD.t21 50.0486
R153 DVDD.t140 DVDD.n5490 49.7525
R154 DVDD.t102 DVDD.n5494 49.7525
R155 DVDD.t129 DVDD.n1884 46.6135
R156 DVDD.t126 DVDD.n4199 46.6135
R157 DVDD.n2669 DVDD 46.0855
R158 DVDD.n2791 DVDD.t9 43.2772
R159 DVDD.n2717 DVDD.n2715 39.6905
R160 DVDD.t40 DVDD.n3026 39.5713
R161 DVDD.n1884 DVDD.t138 35.2118
R162 DVDD.n4199 DVDD.t124 35.2118
R163 DVDD.n1956 DVDD.t155 34.7933
R164 DVDD.n1922 DVDD.t199 34.7929
R165 DVDD.n1920 DVDD.t68 34.7928
R166 DVDD.n1953 DVDD.t45 31.2268
R167 DVDD.t96 DVDD.t140 28.4302
R168 DVDD.t157 DVDD.t148 28.4302
R169 DVDD.t31 DVDD.t21 28.4302
R170 DVDD.t113 DVDD.t102 28.4302
R171 DVDD.n5487 DVDD.t143 25.0246
R172 DVDD.n5661 DVDD.t99 25.0246
R173 DVDD.n4147 DVDD.t205 21.0793
R174 DVDD.n1873 DVDD.t207 21.0793
R175 DVDD.n3959 DVDD.t214 21.0793
R176 DVDD.n4137 DVDD.t219 21.0793
R177 DVDD.n3383 DVDD.n3382 20.9305
R178 DVDD.n3337 DVDD.n3310 20.9305
R179 DVDD.n3318 DVDD.n3316 20.7205
R180 DVDD.n3332 DVDD.n3331 20.7205
R181 DVDD.n2012 DVDD 19.7447
R182 DVDD.n3660 DVDD 19.7447
R183 DVDD.n2009 DVDD 19.7447
R184 DVDD.n3657 DVDD 19.7447
R185 DVDD.n5661 DVDD.n5660 19.6523
R186 DVDD.n5487 DVDD.n5486 19.5041
R187 DVDD DVDD.t220 19.104
R188 DVDD.t220 DVDD 19.104
R189 DVDD DVDD.t210 19.104
R190 DVDD.t210 DVDD 19.104
R191 DVDD DVDD.t217 19.104
R192 DVDD.t217 DVDD 19.104
R193 DVDD DVDD.t206 19.104
R194 DVDD.t206 DVDD 19.104
R195 DVDD DVDD.t216 19.104
R196 DVDD.t216 DVDD 19.104
R197 DVDD DVDD.t211 19.104
R198 DVDD.t211 DVDD 19.104
R199 DVDD DVDD.t218 19.104
R200 DVDD.t218 DVDD 19.104
R201 DVDD.t208 DVDD 19.104
R202 DVDD DVDD.t208 19.104
R203 DVDD.n3337 DVDD.n3336 14.6999
R204 DVDD.n3383 DVDD.n3236 14.6999
R205 DVDD.n3331 DVDD.n3312 14.6413
R206 DVDD.n3318 DVDD.n3241 14.6413
R207 DVDD.n2013 DVDD 14.3168
R208 DVDD.n3661 DVDD 14.3168
R209 DVDD.n2010 DVDD 14.3168
R210 DVDD.n3658 DVDD 14.3168
R211 DVDD.n5499 DVDD.t24 14.2154
R212 DVDD.t160 DVDD.n261 12.8827
R213 DVDD.n5486 DVDD.n5485 12.4047
R214 DVDD.n5660 DVDD.n5659 12.3937
R215 DVDD.n2077 DVDD.n2076 9.73503
R216 DVDD DVDD.t215 7.42907
R217 DVDD DVDD.t212 7.42907
R218 DVDD DVDD.t213 7.42907
R219 DVDD DVDD.t209 7.42907
R220 DVDD.n3027 DVDD.n2076 7.19237
R221 DVDD.n2707 DVDD.t55 6.5562
R222 DVDD.n2769 DVDD.n2768 6.3005
R223 DVDD.n2775 DVDD.n2746 6.3005
R224 DVDD.n2777 DVDD.n2746 6.3005
R225 DVDD.n2783 DVDD.n2723 6.3005
R226 DVDD.n2786 DVDD.n2723 6.3005
R227 DVDD.n2788 DVDD.n2723 6.3005
R228 DVDD.n2769 DVDD.n2748 6.3005
R229 DVDD.n2752 DVDD.n2748 6.3005
R230 DVDD.n2755 DVDD.n2748 6.3005
R231 DVDD.n2751 DVDD.n2748 6.3005
R232 DVDD.n2775 DVDD.n2748 6.3005
R233 DVDD.n2777 DVDD.n2748 6.3005
R234 DVDD.n2737 DVDD.n2725 6.3005
R235 DVDD.n2786 DVDD.n2725 6.3005
R236 DVDD.n2788 DVDD.n2725 6.3005
R237 DVDD.n2769 DVDD.n2745 6.3005
R238 DVDD.n2752 DVDD.n2745 6.3005
R239 DVDD.n2755 DVDD.n2745 6.3005
R240 DVDD.n2751 DVDD.n2745 6.3005
R241 DVDD.n2775 DVDD.n2745 6.3005
R242 DVDD.n2777 DVDD.n2745 6.3005
R243 DVDD.n2737 DVDD.n2722 6.3005
R244 DVDD.n2788 DVDD.n2722 6.3005
R245 DVDD.n2769 DVDD.n2727 6.3005
R246 DVDD.n2752 DVDD.n2727 6.3005
R247 DVDD.n2755 DVDD.n2727 6.3005
R248 DVDD.n2751 DVDD.n2727 6.3005
R249 DVDD.n2775 DVDD.n2727 6.3005
R250 DVDD.n2777 DVDD.n2727 6.3005
R251 DVDD.n2786 DVDD.n2727 6.3005
R252 DVDD.n2788 DVDD.n2727 6.3005
R253 DVDD.n2769 DVDD.n2744 6.3005
R254 DVDD.n2752 DVDD.n2744 6.3005
R255 DVDD.n2755 DVDD.n2744 6.3005
R256 DVDD.n2751 DVDD.n2744 6.3005
R257 DVDD.n2775 DVDD.n2744 6.3005
R258 DVDD.n2777 DVDD.n2744 6.3005
R259 DVDD.n2737 DVDD.n2721 6.3005
R260 DVDD.n2786 DVDD.n2721 6.3005
R261 DVDD.n2788 DVDD.n2721 6.3005
R262 DVDD.n2769 DVDD.n2749 6.3005
R263 DVDD.n2752 DVDD.n2749 6.3005
R264 DVDD.n2755 DVDD.n2749 6.3005
R265 DVDD.n2751 DVDD.n2749 6.3005
R266 DVDD.n2775 DVDD.n2749 6.3005
R267 DVDD.n2777 DVDD.n2749 6.3005
R268 DVDD.n2737 DVDD.n2728 6.3005
R269 DVDD.n2786 DVDD.n2728 6.3005
R270 DVDD.n2788 DVDD.n2728 6.3005
R271 DVDD.n2769 DVDD.n2743 6.3005
R272 DVDD.n2752 DVDD.n2743 6.3005
R273 DVDD.n2755 DVDD.n2743 6.3005
R274 DVDD.n2751 DVDD.n2743 6.3005
R275 DVDD.n2775 DVDD.n2743 6.3005
R276 DVDD.n2777 DVDD.n2743 6.3005
R277 DVDD.n2737 DVDD.n2720 6.3005
R278 DVDD.n2786 DVDD.n2720 6.3005
R279 DVDD.n2788 DVDD.n2720 6.3005
R280 DVDD.n2776 DVDD.n2752 6.3005
R281 DVDD.n2776 DVDD.n2755 6.3005
R282 DVDD.n2776 DVDD.n2751 6.3005
R283 DVDD.n2776 DVDD.n2775 6.3005
R284 DVDD.n2777 DVDD.n2776 6.3005
R285 DVDD.n2787 DVDD.n2737 6.3005
R286 DVDD.n2787 DVDD.n2786 6.3005
R287 DVDD.n2787 DVDD.n2733 6.3005
R288 DVDD.n2788 DVDD.n2787 6.3005
R289 DVDD.n5497 DVDD.n5493 5.57024
R290 DVDD.n3241 DVDD.n3239 5.56181
R291 DVDD.n3333 DVDD.n3312 5.56181
R292 DVDD.n5489 DVDD.n262 5.41553
R293 DVDD.n5493 DVDD.n262 5.41553
R294 DVDD.n5497 DVDD.n5496 5.41553
R295 DVDD.n5496 DVDD.n256 5.41553
R296 DVDD.n3336 DVDD.n3311 5.21853
R297 DVDD.n3381 DVDD.n3236 5.21853
R298 DVDD.n3380 DVDD.n3379 4.9705
R299 DVDD.n3335 DVDD.n3334 4.9005
R300 DVDD.n2048 DVDD.n2047 4.66866
R301 DVDD.n2067 DVDD.n2065 4.66866
R302 DVDD.n2063 DVDD.n2062 4.66866
R303 DVDD.n3054 DVDD.n3053 4.66866
R304 DVDD.n1682 DVDD.n1675 4.66866
R305 DVDD.n3815 DVDD.n1836 4.66866
R306 DVDD.n4065 DVDD.n4052 4.66866
R307 DVDD.n1761 DVDD.n1730 4.66866
R308 DVDD.n2716 DVDD.t30 4.51467
R309 DVDD.n3417 DVDD.n3416 4.5005
R310 DVDD.n3416 DVDD.n3411 4.5005
R311 DVDD.n3414 DVDD.n3411 4.5005
R312 DVDD.n3416 DVDD.n3415 4.5005
R313 DVDD.n3415 DVDD.n3414 4.5005
R314 DVDD.n3113 DVDD.n3111 4.5005
R315 DVDD.n3603 DVDD.n3111 4.5005
R316 DVDD.n3604 DVDD.n3603 4.5005
R317 DVDD.n3605 DVDD.n3111 4.5005
R318 DVDD.n3605 DVDD.n3604 4.5005
R319 DVDD.n3224 DVDD.n3223 4.5005
R320 DVDD.n3353 DVDD.n3350 4.5005
R321 DVDD.n3395 DVDD.n3223 4.5005
R322 DVDD.n3352 DVDD.n3349 4.5005
R323 DVDD.n3353 DVDD.n3352 4.5005
R324 DVDD.n3396 DVDD.n3224 4.5005
R325 DVDD.n3396 DVDD.n3395 4.5005
R326 DVDD.n3350 DVDD.n3349 4.5005
R327 DVDD.n3313 DVDD.n3276 4.5005
R328 DVDD.n3378 DVDD.n3377 4.5005
R329 DVDD.n3377 DVDD.n3376 4.5005
R330 DVDD.n3326 DVDD.n3276 4.5005
R331 DVDD.n2804 DVDD.n2702 4.5005
R332 DVDD.n2804 DVDD.n2803 4.5005
R333 DVDD.n2803 DVDD.n2704 4.5005
R334 DVDD.n2802 DVDD.n2800 4.5005
R335 DVDD.n2803 DVDD.n2802 4.5005
R336 DVDD.n2842 DVDD.n2841 4.5005
R337 DVDD.n2841 DVDD.n2695 4.5005
R338 DVDD.n2844 DVDD.n2695 4.5005
R339 DVDD.n2840 DVDD.n2695 4.5005
R340 DVDD.n2840 DVDD.n2839 4.5005
R341 DVDD.n2687 DVDD.n2682 4.5005
R342 DVDD.n2864 DVDD.n2687 4.5005
R343 DVDD.n2687 DVDD.n2136 4.5005
R344 DVDD.n2689 DVDD.n2136 4.5005
R345 DVDD.n2864 DVDD.n2689 4.5005
R346 DVDD.n2689 DVDD.n2682 4.5005
R347 DVDD.n2686 DVDD.n2682 4.5005
R348 DVDD.n2864 DVDD.n2686 4.5005
R349 DVDD.n2686 DVDD.n2136 4.5005
R350 DVDD.n2690 DVDD.n2682 4.5005
R351 DVDD.n2864 DVDD.n2690 4.5005
R352 DVDD.n2690 DVDD.n2136 4.5005
R353 DVDD.n2685 DVDD.n2136 4.5005
R354 DVDD.n2864 DVDD.n2685 4.5005
R355 DVDD.n2685 DVDD.n2682 4.5005
R356 DVDD.n2691 DVDD.n2682 4.5005
R357 DVDD.n2864 DVDD.n2691 4.5005
R358 DVDD.n2691 DVDD.n2136 4.5005
R359 DVDD.n2684 DVDD.n2682 4.5005
R360 DVDD.n2864 DVDD.n2684 4.5005
R361 DVDD.n2684 DVDD.n2136 4.5005
R362 DVDD.n2692 DVDD.n2136 4.5005
R363 DVDD.n2864 DVDD.n2692 4.5005
R364 DVDD.n2692 DVDD.n2682 4.5005
R365 DVDD.n2683 DVDD.n2136 4.5005
R366 DVDD.n2864 DVDD.n2683 4.5005
R367 DVDD.n2683 DVDD.n2682 4.5005
R368 DVDD.n2863 DVDD.n2682 4.5005
R369 DVDD.n2864 DVDD.n2863 4.5005
R370 DVDD.n2863 DVDD.n2136 4.5005
R371 DVDD.n2947 DVDD.n2092 4.5005
R372 DVDD.n2097 DVDD.n2092 4.5005
R373 DVDD.n2945 DVDD.n2092 4.5005
R374 DVDD.n2947 DVDD.n2093 4.5005
R375 DVDD.n2097 DVDD.n2093 4.5005
R376 DVDD.n2945 DVDD.n2093 4.5005
R377 DVDD.n2945 DVDD.n2091 4.5005
R378 DVDD.n2097 DVDD.n2091 4.5005
R379 DVDD.n2947 DVDD.n2091 4.5005
R380 DVDD.n2947 DVDD.n2094 4.5005
R381 DVDD.n2097 DVDD.n2094 4.5005
R382 DVDD.n2945 DVDD.n2094 4.5005
R383 DVDD.n2947 DVDD.n2090 4.5005
R384 DVDD.n2097 DVDD.n2090 4.5005
R385 DVDD.n2945 DVDD.n2090 4.5005
R386 DVDD.n2945 DVDD.n2095 4.5005
R387 DVDD.n2097 DVDD.n2095 4.5005
R388 DVDD.n2947 DVDD.n2095 4.5005
R389 DVDD.n2947 DVDD.n2089 4.5005
R390 DVDD.n2097 DVDD.n2089 4.5005
R391 DVDD.n2945 DVDD.n2089 4.5005
R392 DVDD.n2946 DVDD.n2945 4.5005
R393 DVDD.n2946 DVDD.n2097 4.5005
R394 DVDD.n2947 DVDD.n2946 4.5005
R395 DVDD.n3053 DVDD.n3052 4.5005
R396 DVDD.n3036 DVDD.n3035 4.5005
R397 DVDD.n3043 DVDD.n3042 4.5005
R398 DVDD.n3040 DVDD.n2040 4.5005
R399 DVDD.n3067 DVDD.n1995 4.5005
R400 DVDD.n3069 DVDD.n3068 4.5005
R401 DVDD.n2039 DVDD.n2038 4.5005
R402 DVDD.n2062 DVDD.n2061 4.5005
R403 DVDD.n2067 DVDD.n2066 4.5005
R404 DVDD.n2069 DVDD.n2068 4.5005
R405 DVDD.n2072 DVDD.n2071 4.5005
R406 DVDD.n2073 DVDD.n2027 4.5005
R407 DVDD.n2060 DVDD.n2026 4.5005
R408 DVDD.n2059 DVDD.n2058 4.5005
R409 DVDD.n2050 DVDD.n2041 4.5005
R410 DVDD.n2049 DVDD.n2048 4.5005
R411 DVDD.n3343 DVDD.n3221 4.5005
R412 DVDD.n3371 DVDD.n3370 4.5005
R413 DVDD.n3282 DVDD.n3268 4.5005
R414 DVDD.n3293 DVDD.n3227 4.5005
R415 DVDD.n3390 DVDD.n3228 4.5005
R416 DVDD.n3391 DVDD.n3089 4.5005
R417 DVDD.n3344 DVDD.n3343 4.5005
R418 DVDD.n3370 DVDD.n3369 4.5005
R419 DVDD.n3282 DVDD.n3272 4.5005
R420 DVDD.n3294 DVDD.n3293 4.5005
R421 DVDD.n3299 DVDD.n3228 4.5005
R422 DVDD.n3340 DVDD.n3089 4.5005
R423 DVDD.n3157 DVDD.n3143 4.5005
R424 DVDD.n3160 DVDD.n3143 4.5005
R425 DVDD.n3150 DVDD.n3143 4.5005
R426 DVDD.n3167 DVDD.n3143 4.5005
R427 DVDD.n3151 DVDD.n3143 4.5005
R428 DVDD.n3166 DVDD.n3143 4.5005
R429 DVDD.n3152 DVDD.n3143 4.5005
R430 DVDD.n3165 DVDD.n3143 4.5005
R431 DVDD.n3153 DVDD.n3143 4.5005
R432 DVDD.n3164 DVDD.n3143 4.5005
R433 DVDD.n3154 DVDD.n3143 4.5005
R434 DVDD.n3163 DVDD.n3143 4.5005
R435 DVDD.n3155 DVDD.n3143 4.5005
R436 DVDD.n3162 DVDD.n3143 4.5005
R437 DVDD.n3156 DVDD.n3143 4.5005
R438 DVDD.n3161 DVDD.n3143 4.5005
R439 DVDD.n3571 DVDD.n3158 4.5005
R440 DVDD.n3571 DVDD.n3160 4.5005
R441 DVDD.n3571 DVDD.n3157 4.5005
R442 DVDD.n3568 DVDD.n3161 4.5005
R443 DVDD.n3568 DVDD.n3156 4.5005
R444 DVDD.n3568 DVDD.n3162 4.5005
R445 DVDD.n3568 DVDD.n3155 4.5005
R446 DVDD.n3568 DVDD.n3163 4.5005
R447 DVDD.n3568 DVDD.n3154 4.5005
R448 DVDD.n3568 DVDD.n3164 4.5005
R449 DVDD.n3568 DVDD.n3153 4.5005
R450 DVDD.n3568 DVDD.n3165 4.5005
R451 DVDD.n3568 DVDD.n3152 4.5005
R452 DVDD.n3568 DVDD.n3166 4.5005
R453 DVDD.n3568 DVDD.n3151 4.5005
R454 DVDD.n3568 DVDD.n3167 4.5005
R455 DVDD.n3568 DVDD.n3150 4.5005
R456 DVDD.n3570 DVDD.n3568 4.5005
R457 DVDD.n3568 DVDD.n3158 4.5005
R458 DVDD.n3568 DVDD.n3160 4.5005
R459 DVDD.n3568 DVDD.n3157 4.5005
R460 DVDD.n3571 DVDD.n3161 4.5005
R461 DVDD.n3571 DVDD.n3156 4.5005
R462 DVDD.n3571 DVDD.n3162 4.5005
R463 DVDD.n3571 DVDD.n3155 4.5005
R464 DVDD.n3571 DVDD.n3163 4.5005
R465 DVDD.n3571 DVDD.n3154 4.5005
R466 DVDD.n3571 DVDD.n3164 4.5005
R467 DVDD.n3571 DVDD.n3153 4.5005
R468 DVDD.n3571 DVDD.n3165 4.5005
R469 DVDD.n3571 DVDD.n3152 4.5005
R470 DVDD.n3571 DVDD.n3166 4.5005
R471 DVDD.n3571 DVDD.n3151 4.5005
R472 DVDD.n3571 DVDD.n3167 4.5005
R473 DVDD.n3571 DVDD.n3150 4.5005
R474 DVDD.n3571 DVDD.n3570 4.5005
R475 DVDD.n3514 DVDD.n3172 4.5005
R476 DVDD.n3174 DVDD.n3172 4.5005
R477 DVDD.n3512 DVDD.n3172 4.5005
R478 DVDD.n3175 DVDD.n3172 4.5005
R479 DVDD.n3191 DVDD.n3172 4.5005
R480 DVDD.n3176 DVDD.n3172 4.5005
R481 DVDD.n3190 DVDD.n3172 4.5005
R482 DVDD.n3177 DVDD.n3172 4.5005
R483 DVDD.n3189 DVDD.n3172 4.5005
R484 DVDD.n3178 DVDD.n3172 4.5005
R485 DVDD.n3188 DVDD.n3172 4.5005
R486 DVDD.n3179 DVDD.n3172 4.5005
R487 DVDD.n3187 DVDD.n3172 4.5005
R488 DVDD.n3180 DVDD.n3172 4.5005
R489 DVDD.n3184 DVDD.n3172 4.5005
R490 DVDD.n3182 DVDD.n3172 4.5005
R491 DVDD.n3514 DVDD.n3171 4.5005
R492 DVDD.n3174 DVDD.n3171 4.5005
R493 DVDD.n3512 DVDD.n3171 4.5005
R494 DVDD.n3175 DVDD.n3171 4.5005
R495 DVDD.n3191 DVDD.n3171 4.5005
R496 DVDD.n3176 DVDD.n3171 4.5005
R497 DVDD.n3190 DVDD.n3171 4.5005
R498 DVDD.n3177 DVDD.n3171 4.5005
R499 DVDD.n3189 DVDD.n3171 4.5005
R500 DVDD.n3178 DVDD.n3171 4.5005
R501 DVDD.n3188 DVDD.n3171 4.5005
R502 DVDD.n3179 DVDD.n3171 4.5005
R503 DVDD.n3187 DVDD.n3171 4.5005
R504 DVDD.n3180 DVDD.n3171 4.5005
R505 DVDD.n3186 DVDD.n3171 4.5005
R506 DVDD.n3181 DVDD.n3171 4.5005
R507 DVDD.n3184 DVDD.n3171 4.5005
R508 DVDD.n3182 DVDD.n3171 4.5005
R509 DVDD.n3513 DVDD.n3182 4.5005
R510 DVDD.n3513 DVDD.n3184 4.5005
R511 DVDD.n3513 DVDD.n3181 4.5005
R512 DVDD.n3513 DVDD.n3186 4.5005
R513 DVDD.n3513 DVDD.n3180 4.5005
R514 DVDD.n3513 DVDD.n3187 4.5005
R515 DVDD.n3513 DVDD.n3179 4.5005
R516 DVDD.n3513 DVDD.n3188 4.5005
R517 DVDD.n3513 DVDD.n3178 4.5005
R518 DVDD.n3513 DVDD.n3189 4.5005
R519 DVDD.n3513 DVDD.n3177 4.5005
R520 DVDD.n3513 DVDD.n3190 4.5005
R521 DVDD.n3513 DVDD.n3176 4.5005
R522 DVDD.n3513 DVDD.n3191 4.5005
R523 DVDD.n3513 DVDD.n3175 4.5005
R524 DVDD.n3513 DVDD.n3512 4.5005
R525 DVDD.n3513 DVDD.n3174 4.5005
R526 DVDD.n3514 DVDD.n3513 4.5005
R527 DVDD.n4066 DVDD.n4065 4.5005
R528 DVDD.n4064 DVDD.n4063 4.5005
R529 DVDD.n4055 DVDD.n4054 4.5005
R530 DVDD.n4056 DVDD.n1719 4.5005
R531 DVDD.n4226 DVDD.n4225 4.5005
R532 DVDD.n1728 DVDD.n1720 4.5005
R533 DVDD.n1763 DVDD.n1762 4.5005
R534 DVDD.n1761 DVDD.n1760 4.5005
R535 DVDD.n1682 DVDD.n1680 4.5005
R536 DVDD.n4265 DVDD.n4264 4.5005
R537 DVDD.n4263 DVDD.n4262 4.5005
R538 DVDD.n1684 DVDD.n1683 4.5005
R539 DVDD.n1843 DVDD.n1842 4.5005
R540 DVDD.n3813 DVDD.n3812 4.5005
R541 DVDD.n3814 DVDD.n1840 4.5005
R542 DVDD.n3816 DVDD.n3815 4.5005
R543 DVDD.n3777 DVDD.n1887 4.5005
R544 DVDD.n3777 DVDD.n1861 4.5005
R545 DVDD.n3777 DVDD.n3776 4.5005
R546 DVDD.n2618 DVDD.n2193 4.5005
R547 DVDD.n2620 DVDD.n2193 4.5005
R548 DVDD.n2620 DVDD.n2194 4.5005
R549 DVDD.n2620 DVDD.n2172 4.5005
R550 DVDD.n2620 DVDD.n2195 4.5005
R551 DVDD.n2620 DVDD.n2171 4.5005
R552 DVDD.n2620 DVDD.n2196 4.5005
R553 DVDD.n2620 DVDD.n2170 4.5005
R554 DVDD.n2620 DVDD.n2197 4.5005
R555 DVDD.n2620 DVDD.n2169 4.5005
R556 DVDD.n2619 DVDD.n2618 4.5005
R557 DVDD.n2620 DVDD.n2619 4.5005
R558 DVDD.n2602 DVDD.n2198 4.5005
R559 DVDD.n2602 DVDD.n2601 4.5005
R560 DVDD.n2601 DVDD.n2207 4.5005
R561 DVDD.n2601 DVDD.n2204 4.5005
R562 DVDD.n2601 DVDD.n2209 4.5005
R563 DVDD.n2601 DVDD.n2203 4.5005
R564 DVDD.n2601 DVDD.n2211 4.5005
R565 DVDD.n2601 DVDD.n2202 4.5005
R566 DVDD.n2601 DVDD.n2213 4.5005
R567 DVDD.n2601 DVDD.n2201 4.5005
R568 DVDD.n2600 DVDD.n2198 4.5005
R569 DVDD.n2601 DVDD.n2600 4.5005
R570 DVDD.n3776 DVDD.n3775 4.5005
R571 DVDD.n3775 DVDD.n3730 4.5005
R572 DVDD.n3775 DVDD.n3735 4.5005
R573 DVDD.n3775 DVDD.n3729 4.5005
R574 DVDD.n3775 DVDD.n3736 4.5005
R575 DVDD.n3775 DVDD.n3728 4.5005
R576 DVDD.n3775 DVDD.n3737 4.5005
R577 DVDD.n3775 DVDD.n3727 4.5005
R578 DVDD.n3775 DVDD.n3738 4.5005
R579 DVDD.n3775 DVDD.n1861 4.5005
R580 DVDD.n3775 DVDD.n1887 4.5005
R581 DVDD.n3775 DVDD.n3726 4.5005
R582 DVDD.n3775 DVDD.n3739 4.5005
R583 DVDD.n3775 DVDD.n3725 4.5005
R584 DVDD.n3775 DVDD.n3740 4.5005
R585 DVDD.n3775 DVDD.n3724 4.5005
R586 DVDD.n3775 DVDD.n3741 4.5005
R587 DVDD.n3775 DVDD.n3723 4.5005
R588 DVDD.n3775 DVDD.n3742 4.5005
R589 DVDD.n3775 DVDD.n3722 4.5005
R590 DVDD.n3774 DVDD.n3752 4.5005
R591 DVDD.n3775 DVDD.n3774 4.5005
R592 DVDD.n1323 DVDD.n1321 4.5005
R593 DVDD.n1388 DVDD.n1383 4.5005
R594 DVDD.n1388 DVDD.n1385 4.5005
R595 DVDD.n1323 DVDD.n1322 4.5005
R596 DVDD.n1388 DVDD.n1382 4.5005
R597 DVDD.n1382 DVDD.n1380 4.5005
R598 DVDD.n1325 DVDD.n1318 4.5005
R599 DVDD.n1323 DVDD.n1318 4.5005
R600 DVDD.n1388 DVDD.n1386 4.5005
R601 DVDD.n1386 DVDD.n1380 4.5005
R602 DVDD.n1325 DVDD.n1320 4.5005
R603 DVDD.n1323 DVDD.n1320 4.5005
R604 DVDD.n1325 DVDD.n1317 4.5005
R605 DVDD.n1323 DVDD.n1317 4.5005
R606 DVDD.n1381 DVDD.n1380 4.5005
R607 DVDD.n1388 DVDD.n1381 4.5005
R608 DVDD.n1325 DVDD.n1324 4.5005
R609 DVDD.n1324 DVDD.n1323 4.5005
R610 DVDD.n1387 DVDD.n1380 4.5005
R611 DVDD.n1388 DVDD.n1387 4.5005
R612 DVDD.n1365 DVDD.n1331 4.5005
R613 DVDD.n1332 DVDD.n1331 4.5005
R614 DVDD.n1369 DVDD.n1331 4.5005
R615 DVDD.n1394 DVDD.n1309 4.5005
R616 DVDD.n1394 DVDD.n1311 4.5005
R617 DVDD.n1394 DVDD.n1308 4.5005
R618 DVDD.n1312 DVDD.n1305 4.5005
R619 DVDD.n1394 DVDD.n1312 4.5005
R620 DVDD.n1307 DVDD.n1305 4.5005
R621 DVDD.n1394 DVDD.n1307 4.5005
R622 DVDD.n1313 DVDD.n1305 4.5005
R623 DVDD.n1394 DVDD.n1313 4.5005
R624 DVDD.n1306 DVDD.n1305 4.5005
R625 DVDD.n1394 DVDD.n1306 4.5005
R626 DVDD.n1308 DVDD.n1305 4.5005
R627 DVDD.n1311 DVDD.n1305 4.5005
R628 DVDD.n1309 DVDD.n1305 4.5005
R629 DVDD.n1393 DVDD.n1305 4.5005
R630 DVDD.n1394 DVDD.n1393 4.5005
R631 DVDD.n1554 DVDD.n1214 4.5005
R632 DVDD.n1554 DVDD.n1221 4.5005
R633 DVDD.n1554 DVDD.n1215 4.5005
R634 DVDD.n1556 DVDD.n1217 4.5005
R635 DVDD.n1554 DVDD.n1217 4.5005
R636 DVDD.n1556 DVDD.n1219 4.5005
R637 DVDD.n1554 DVDD.n1219 4.5005
R638 DVDD.n1556 DVDD.n1216 4.5005
R639 DVDD.n1554 DVDD.n1216 4.5005
R640 DVDD.n1556 DVDD.n1220 4.5005
R641 DVDD.n1554 DVDD.n1220 4.5005
R642 DVDD.n1556 DVDD.n1215 4.5005
R643 DVDD.n1556 DVDD.n1221 4.5005
R644 DVDD.n1556 DVDD.n1214 4.5005
R645 DVDD.n1556 DVDD.n1555 4.5005
R646 DVDD.n1555 DVDD.n1554 4.5005
R647 DVDD.n1364 DVDD.n1329 4.5005
R648 DVDD.n1364 DVDD.n1336 4.5005
R649 DVDD.n1368 DVDD.n1336 4.5005
R650 DVDD.n1368 DVDD.n1339 4.5005
R651 DVDD.n1368 DVDD.n1335 4.5005
R652 DVDD.n1368 DVDD.n1329 4.5005
R653 DVDD.n1369 DVDD.n1368 4.5005
R654 DVDD.n1368 DVDD.n1367 4.5005
R655 DVDD.n1367 DVDD.n1331 4.5005
R656 DVDD.n1195 DVDD.n1192 4.5005
R657 DVDD.n1200 DVDD.n1192 4.5005
R658 DVDD.n1577 DVDD.n1192 4.5005
R659 DVDD.n1577 DVDD.n1576 4.5005
R660 DVDD.n1576 DVDD.n1199 4.5005
R661 DVDD.n1576 DVDD.n1196 4.5005
R662 DVDD.n1576 DVDD.n1200 4.5005
R663 DVDD.n1576 DVDD.n1195 4.5005
R664 DVDD.n1576 DVDD.n1202 4.5005
R665 DVDD.n1576 DVDD.n1194 4.5005
R666 DVDD.n1576 DVDD.n1575 4.5005
R667 DVDD.n1575 DVDD.n1192 4.5005
R668 DVDD.n5422 DVDD.n341 4.5005
R669 DVDD.n5915 DVDD.n5914 4.5005
R670 DVDD.n5420 DVDD.n5417 4.5005
R671 DVDD.n5917 DVDD.n94 4.5005
R672 DVDD.n5422 DVDD.n342 4.5005
R673 DVDD.n350 DVDD.n342 4.5005
R674 DVDD.n5420 DVDD.n342 4.5005
R675 DVDD.n5915 DVDD.n95 4.5005
R676 DVDD.n105 DVDD.n95 4.5005
R677 DVDD.n5917 DVDD.n95 4.5005
R678 DVDD.n350 DVDD.n347 4.5005
R679 DVDD.n5420 DVDD.n347 4.5005
R680 DVDD.n5915 DVDD.n93 4.5005
R681 DVDD.n350 DVDD.n335 4.5005
R682 DVDD.n5420 DVDD.n335 4.5005
R683 DVDD.n5915 DVDD.n96 4.5005
R684 DVDD.n350 DVDD.n346 4.5005
R685 DVDD.n5420 DVDD.n346 4.5005
R686 DVDD.n5915 DVDD.n92 4.5005
R687 DVDD.n350 DVDD.n336 4.5005
R688 DVDD.n5420 DVDD.n336 4.5005
R689 DVDD.n5915 DVDD.n97 4.5005
R690 DVDD.n350 DVDD.n345 4.5005
R691 DVDD.n5420 DVDD.n345 4.5005
R692 DVDD.n5915 DVDD.n91 4.5005
R693 DVDD.n350 DVDD.n337 4.5005
R694 DVDD.n5915 DVDD.n98 4.5005
R695 DVDD.n350 DVDD.n344 4.5005
R696 DVDD.n5915 DVDD.n90 4.5005
R697 DVDD.n350 DVDD.n338 4.5005
R698 DVDD.n5420 DVDD.n338 4.5005
R699 DVDD.n5915 DVDD.n99 4.5005
R700 DVDD.n350 DVDD.n343 4.5005
R701 DVDD.n5420 DVDD.n343 4.5005
R702 DVDD.n5915 DVDD.n89 4.5005
R703 DVDD.n350 DVDD.n339 4.5005
R704 DVDD.n5420 DVDD.n339 4.5005
R705 DVDD.n5915 DVDD.n100 4.5005
R706 DVDD.n5422 DVDD.n339 4.5005
R707 DVDD.n5422 DVDD.n343 4.5005
R708 DVDD.n5422 DVDD.n338 4.5005
R709 DVDD.n5422 DVDD.n344 4.5005
R710 DVDD.n5422 DVDD.n337 4.5005
R711 DVDD.n5422 DVDD.n345 4.5005
R712 DVDD.n5422 DVDD.n336 4.5005
R713 DVDD.n5422 DVDD.n346 4.5005
R714 DVDD.n5422 DVDD.n335 4.5005
R715 DVDD.n5422 DVDD.n347 4.5005
R716 DVDD.n105 DVDD.n93 4.5005
R717 DVDD.n5917 DVDD.n93 4.5005
R718 DVDD.n105 DVDD.n96 4.5005
R719 DVDD.n5917 DVDD.n96 4.5005
R720 DVDD.n105 DVDD.n92 4.5005
R721 DVDD.n5917 DVDD.n92 4.5005
R722 DVDD.n105 DVDD.n97 4.5005
R723 DVDD.n5917 DVDD.n97 4.5005
R724 DVDD.n105 DVDD.n91 4.5005
R725 DVDD.n5917 DVDD.n91 4.5005
R726 DVDD.n5917 DVDD.n98 4.5005
R727 DVDD.n5917 DVDD.n90 4.5005
R728 DVDD.n105 DVDD.n99 4.5005
R729 DVDD.n5917 DVDD.n99 4.5005
R730 DVDD.n105 DVDD.n89 4.5005
R731 DVDD.n5917 DVDD.n89 4.5005
R732 DVDD.n105 DVDD.n100 4.5005
R733 DVDD.n5917 DVDD.n100 4.5005
R734 DVDD.n5917 DVDD.n88 4.5005
R735 DVDD.n5915 DVDD.n88 4.5005
R736 DVDD.n5420 DVDD.n334 4.5005
R737 DVDD.n5422 DVDD.n334 4.5005
R738 DVDD.n5917 DVDD.n5916 4.5005
R739 DVDD.n5916 DVDD.n5915 4.5005
R740 DVDD.n5421 DVDD.n5420 4.5005
R741 DVDD.n5422 DVDD.n5421 4.5005
R742 DVDD.n5427 DVDD.n327 4.5005
R743 DVDD.n327 DVDD.n321 4.5005
R744 DVDD.n5427 DVDD.n5426 4.5005
R745 DVDD.n5426 DVDD.n321 4.5005
R746 DVDD.n5427 DVDD.n326 4.5005
R747 DVDD.n326 DVDD.n321 4.5005
R748 DVDD.n5919 DVDD.n77 4.5005
R749 DVDD.n5919 DVDD.n79 4.5005
R750 DVDD.n81 DVDD.n77 4.5005
R751 DVDD.n81 DVDD.n79 4.5005
R752 DVDD.n5921 DVDD.n77 4.5005
R753 DVDD.n5921 DVDD.n79 4.5005
R754 DVDD.n1578 DVDD.n1120 4.5005
R755 DVDD.n1579 DVDD.n1578 4.5005
R756 DVDD.n1189 DVDD.n1120 4.5005
R757 DVDD.n1582 DVDD.n1134 4.5005
R758 DVDD.n1582 DVDD.n1130 4.5005
R759 DVDD.n1582 DVDD.n1136 4.5005
R760 DVDD.n1582 DVDD.n1129 4.5005
R761 DVDD.n1582 DVDD.n1138 4.5005
R762 DVDD.n1582 DVDD.n1128 4.5005
R763 DVDD.n1582 DVDD.n1140 4.5005
R764 DVDD.n1582 DVDD.n1127 4.5005
R765 DVDD.n1582 DVDD.n1142 4.5005
R766 DVDD.n1582 DVDD.n1126 4.5005
R767 DVDD.n1582 DVDD.n1144 4.5005
R768 DVDD.n1582 DVDD.n1125 4.5005
R769 DVDD.n1582 DVDD.n1146 4.5005
R770 DVDD.n1582 DVDD.n1124 4.5005
R771 DVDD.n1582 DVDD.n1148 4.5005
R772 DVDD.n1582 DVDD.n1123 4.5005
R773 DVDD.n1582 DVDD.n1581 4.5005
R774 DVDD.n1582 DVDD.n1122 4.5005
R775 DVDD.n1583 DVDD.n1120 4.5005
R776 DVDD.n1583 DVDD.n1582 4.5005
R777 DVDD.n5379 DVDD.n378 4.5005
R778 DVDD.n5381 DVDD.n378 4.5005
R779 DVDD.n5379 DVDD.n380 4.5005
R780 DVDD.n5381 DVDD.n380 4.5005
R781 DVDD.n5379 DVDD.n377 4.5005
R782 DVDD.n5381 DVDD.n377 4.5005
R783 DVDD.n5380 DVDD.n5379 4.5005
R784 DVDD.n5381 DVDD.n5380 4.5005
R785 DVDD.n5359 DVDD.n401 4.5005
R786 DVDD.n5361 DVDD.n401 4.5005
R787 DVDD.n5359 DVDD.n403 4.5005
R788 DVDD.n5361 DVDD.n403 4.5005
R789 DVDD.n5359 DVDD.n400 4.5005
R790 DVDD.n5361 DVDD.n400 4.5005
R791 DVDD.n5360 DVDD.n5359 4.5005
R792 DVDD.n5361 DVDD.n5360 4.5005
R793 DVDD.n5338 DVDD.n425 4.5005
R794 DVDD.n5340 DVDD.n425 4.5005
R795 DVDD.n5338 DVDD.n427 4.5005
R796 DVDD.n5340 DVDD.n427 4.5005
R797 DVDD.n5338 DVDD.n424 4.5005
R798 DVDD.n5340 DVDD.n424 4.5005
R799 DVDD.n5339 DVDD.n5338 4.5005
R800 DVDD.n5340 DVDD.n5339 4.5005
R801 DVDD.n5134 DVDD.n5102 4.5005
R802 DVDD.n5102 DVDD.n449 4.5005
R803 DVDD.n5139 DVDD.n5134 4.5005
R804 DVDD.n5139 DVDD.n449 4.5005
R805 DVDD.n5137 DVDD.n5134 4.5005
R806 DVDD.n5137 DVDD.n449 4.5005
R807 DVDD.n5135 DVDD.n5134 4.5005
R808 DVDD.n5135 DVDD.n449 4.5005
R809 DVDD.n136 DVDD.n130 4.5005
R810 DVDD.n5849 DVDD.n136 4.5005
R811 DVDD.n138 DVDD.n130 4.5005
R812 DVDD.n5849 DVDD.n138 4.5005
R813 DVDD.n135 DVDD.n130 4.5005
R814 DVDD.n5849 DVDD.n135 4.5005
R815 DVDD.n5848 DVDD.n130 4.5005
R816 DVDD.n5849 DVDD.n5848 4.5005
R817 DVDD.n79 DVDD.n74 4.5005
R818 DVDD.n77 DVDD.n74 4.5005
R819 DVDD.n76 DVDD.n74 4.5005
R820 DVDD.n5920 DVDD.n74 4.5005
R821 DVDD.n5921 DVDD.n76 4.5005
R822 DVDD.n5921 DVDD.n5920 4.5005
R823 DVDD.n81 DVDD.n76 4.5005
R824 DVDD.n5920 DVDD.n81 4.5005
R825 DVDD.n5919 DVDD.n76 4.5005
R826 DVDD.n5920 DVDD.n5919 4.5005
R827 DVDD.n5428 DVDD.n322 4.5005
R828 DVDD.n5428 DVDD.n324 4.5005
R829 DVDD.n5428 DVDD.n321 4.5005
R830 DVDD.n5428 DVDD.n5427 4.5005
R831 DVDD.n327 DVDD.n322 4.5005
R832 DVDD.n5426 DVDD.n322 4.5005
R833 DVDD.n326 DVDD.n322 4.5005
R834 DVDD.n326 DVDD.n324 4.5005
R835 DVDD.n5426 DVDD.n324 4.5005
R836 DVDD.n327 DVDD.n324 4.5005
R837 DVDD.n5912 DVDD.n114 4.5005
R838 DVDD.n5912 DVDD.n5908 4.5005
R839 DVDD.n5912 DVDD.n113 4.5005
R840 DVDD.n5909 DVDD.n108 4.5005
R841 DVDD.n5909 DVDD.n107 4.5005
R842 DVDD.n5912 DVDD.n5909 4.5005
R843 DVDD.n112 DVDD.n108 4.5005
R844 DVDD.n112 DVDD.n107 4.5005
R845 DVDD.n5912 DVDD.n112 4.5005
R846 DVDD.n5910 DVDD.n108 4.5005
R847 DVDD.n5910 DVDD.n107 4.5005
R848 DVDD.n5912 DVDD.n5910 4.5005
R849 DVDD.n111 DVDD.n108 4.5005
R850 DVDD.n111 DVDD.n107 4.5005
R851 DVDD.n5912 DVDD.n111 4.5005
R852 DVDD.n5912 DVDD.n5911 4.5005
R853 DVDD.n5912 DVDD.n110 4.5005
R854 DVDD.n110 DVDD.n107 4.5005
R855 DVDD.n110 DVDD.n108 4.5005
R856 DVDD.n5911 DVDD.n107 4.5005
R857 DVDD.n5911 DVDD.n108 4.5005
R858 DVDD.n113 DVDD.n107 4.5005
R859 DVDD.n113 DVDD.n108 4.5005
R860 DVDD.n5908 DVDD.n107 4.5005
R861 DVDD.n5908 DVDD.n108 4.5005
R862 DVDD.n114 DVDD.n107 4.5005
R863 DVDD.n114 DVDD.n108 4.5005
R864 DVDD.n5912 DVDD.n102 4.5005
R865 DVDD.n109 DVDD.n108 4.5005
R866 DVDD.n109 DVDD.n107 4.5005
R867 DVDD.n5912 DVDD.n109 4.5005
R868 DVDD.n5913 DVDD.n108 4.5005
R869 DVDD.n5913 DVDD.n107 4.5005
R870 DVDD.n5913 DVDD.n5912 4.5005
R871 DVDD.n108 DVDD.n102 4.5005
R872 DVDD.n107 DVDD.n102 4.5005
R873 DVDD.n5415 DVDD.n5410 4.5005
R874 DVDD.n5415 DVDD.n5411 4.5005
R875 DVDD.n5415 DVDD.n5409 4.5005
R876 DVDD.n5412 DVDD.n325 4.5005
R877 DVDD.n5412 DVDD.n353 4.5005
R878 DVDD.n5415 DVDD.n5412 4.5005
R879 DVDD.n5408 DVDD.n325 4.5005
R880 DVDD.n5408 DVDD.n353 4.5005
R881 DVDD.n5415 DVDD.n5408 4.5005
R882 DVDD.n5413 DVDD.n325 4.5005
R883 DVDD.n5413 DVDD.n353 4.5005
R884 DVDD.n5415 DVDD.n5413 4.5005
R885 DVDD.n5407 DVDD.n325 4.5005
R886 DVDD.n5407 DVDD.n353 4.5005
R887 DVDD.n5415 DVDD.n5407 4.5005
R888 DVDD.n5415 DVDD.n5414 4.5005
R889 DVDD.n5415 DVDD.n5406 4.5005
R890 DVDD.n5406 DVDD.n353 4.5005
R891 DVDD.n5406 DVDD.n325 4.5005
R892 DVDD.n5414 DVDD.n353 4.5005
R893 DVDD.n5414 DVDD.n325 4.5005
R894 DVDD.n5409 DVDD.n353 4.5005
R895 DVDD.n5409 DVDD.n325 4.5005
R896 DVDD.n5411 DVDD.n353 4.5005
R897 DVDD.n5411 DVDD.n325 4.5005
R898 DVDD.n5410 DVDD.n353 4.5005
R899 DVDD.n5410 DVDD.n325 4.5005
R900 DVDD.n5415 DVDD.n349 4.5005
R901 DVDD.n352 DVDD.n325 4.5005
R902 DVDD.n353 DVDD.n352 4.5005
R903 DVDD.n5415 DVDD.n352 4.5005
R904 DVDD.n5416 DVDD.n325 4.5005
R905 DVDD.n5416 DVDD.n353 4.5005
R906 DVDD.n5416 DVDD.n5415 4.5005
R907 DVDD.n349 DVDD.n325 4.5005
R908 DVDD.n353 DVDD.n349 4.5005
R909 DVDD.n285 DVDD.n271 4.5005
R910 DVDD.n5475 DVDD.n285 4.5005
R911 DVDD.n283 DVDD.n271 4.5005
R912 DVDD.n5475 DVDD.n283 4.5005
R913 DVDD.n286 DVDD.n271 4.5005
R914 DVDD.n5475 DVDD.n286 4.5005
R915 DVDD.n282 DVDD.n271 4.5005
R916 DVDD.n5475 DVDD.n282 4.5005
R917 DVDD.n287 DVDD.n271 4.5005
R918 DVDD.n5475 DVDD.n287 4.5005
R919 DVDD.n281 DVDD.n271 4.5005
R920 DVDD.n5475 DVDD.n281 4.5005
R921 DVDD.n288 DVDD.n271 4.5005
R922 DVDD.n5475 DVDD.n288 4.5005
R923 DVDD.n280 DVDD.n271 4.5005
R924 DVDD.n5475 DVDD.n280 4.5005
R925 DVDD.n289 DVDD.n271 4.5005
R926 DVDD.n5475 DVDD.n289 4.5005
R927 DVDD.n279 DVDD.n271 4.5005
R928 DVDD.n5475 DVDD.n279 4.5005
R929 DVDD.n290 DVDD.n271 4.5005
R930 DVDD.n5475 DVDD.n290 4.5005
R931 DVDD.n278 DVDD.n271 4.5005
R932 DVDD.n5475 DVDD.n278 4.5005
R933 DVDD.n291 DVDD.n271 4.5005
R934 DVDD.n5475 DVDD.n291 4.5005
R935 DVDD.n277 DVDD.n271 4.5005
R936 DVDD.n5475 DVDD.n277 4.5005
R937 DVDD.n292 DVDD.n271 4.5005
R938 DVDD.n5475 DVDD.n292 4.5005
R939 DVDD.n276 DVDD.n271 4.5005
R940 DVDD.n5475 DVDD.n276 4.5005
R941 DVDD.n293 DVDD.n271 4.5005
R942 DVDD.n5475 DVDD.n293 4.5005
R943 DVDD.n275 DVDD.n271 4.5005
R944 DVDD.n5475 DVDD.n275 4.5005
R945 DVDD.n5476 DVDD.n271 4.5005
R946 DVDD.n5476 DVDD.n5475 4.5005
R947 DVDD.n5563 DVDD.n69 4.5005
R948 DVDD.n5649 DVDD.n69 4.5005
R949 DVDD.n5574 DVDD.n5563 4.5005
R950 DVDD.n5649 DVDD.n5574 4.5005
R951 DVDD.n5602 DVDD.n5563 4.5005
R952 DVDD.n5649 DVDD.n5602 4.5005
R953 DVDD.n5573 DVDD.n5563 4.5005
R954 DVDD.n5649 DVDD.n5573 4.5005
R955 DVDD.n5603 DVDD.n5563 4.5005
R956 DVDD.n5649 DVDD.n5603 4.5005
R957 DVDD.n5572 DVDD.n5563 4.5005
R958 DVDD.n5649 DVDD.n5572 4.5005
R959 DVDD.n5604 DVDD.n5563 4.5005
R960 DVDD.n5649 DVDD.n5604 4.5005
R961 DVDD.n5571 DVDD.n5563 4.5005
R962 DVDD.n5649 DVDD.n5571 4.5005
R963 DVDD.n5605 DVDD.n5563 4.5005
R964 DVDD.n5649 DVDD.n5605 4.5005
R965 DVDD.n5570 DVDD.n5563 4.5005
R966 DVDD.n5649 DVDD.n5570 4.5005
R967 DVDD.n5606 DVDD.n5563 4.5005
R968 DVDD.n5649 DVDD.n5606 4.5005
R969 DVDD.n5569 DVDD.n5563 4.5005
R970 DVDD.n5649 DVDD.n5569 4.5005
R971 DVDD.n5607 DVDD.n5563 4.5005
R972 DVDD.n5649 DVDD.n5607 4.5005
R973 DVDD.n5568 DVDD.n5563 4.5005
R974 DVDD.n5649 DVDD.n5568 4.5005
R975 DVDD.n5608 DVDD.n5563 4.5005
R976 DVDD.n5649 DVDD.n5608 4.5005
R977 DVDD.n5567 DVDD.n5563 4.5005
R978 DVDD.n5649 DVDD.n5567 4.5005
R979 DVDD.n5648 DVDD.n5563 4.5005
R980 DVDD.n5649 DVDD.n5648 4.5005
R981 DVDD.n5566 DVDD.n5563 4.5005
R982 DVDD.n5649 DVDD.n5566 4.5005
R983 DVDD.n5650 DVDD.n5563 4.5005
R984 DVDD.n5650 DVDD.n5649 4.5005
R985 DVDD.n4411 DVDD.n1584 4.5005
R986 DVDD.n4414 DVDD.n1584 4.5005
R987 DVDD.n4414 DVDD.n1118 4.5005
R988 DVDD.n4414 DVDD.n1585 4.5005
R989 DVDD.n4414 DVDD.n1117 4.5005
R990 DVDD.n4414 DVDD.n1586 4.5005
R991 DVDD.n4414 DVDD.n1116 4.5005
R992 DVDD.n4414 DVDD.n1587 4.5005
R993 DVDD.n4414 DVDD.n1115 4.5005
R994 DVDD.n4414 DVDD.n1588 4.5005
R995 DVDD.n4414 DVDD.n1114 4.5005
R996 DVDD.n4414 DVDD.n1589 4.5005
R997 DVDD.n4414 DVDD.n1113 4.5005
R998 DVDD.n4414 DVDD.n1590 4.5005
R999 DVDD.n4414 DVDD.n1112 4.5005
R1000 DVDD.n4414 DVDD.n1591 4.5005
R1001 DVDD.n4414 DVDD.n1111 4.5005
R1002 DVDD.n4414 DVDD.n1592 4.5005
R1003 DVDD.n4414 DVDD.n1110 4.5005
R1004 DVDD.n4414 DVDD.n1593 4.5005
R1005 DVDD.n4414 DVDD.n1109 4.5005
R1006 DVDD.n4413 DVDD.n4398 4.5005
R1007 DVDD.n4414 DVDD.n4413 4.5005
R1008 DVDD.n4498 DVDD.n1073 4.5005
R1009 DVDD.n4560 DVDD.n4498 4.5005
R1010 DVDD.n4560 DVDD.n1084 4.5005
R1011 DVDD.n1084 DVDD.n1073 4.5005
R1012 DVDD.n4560 DVDD.n4499 4.5005
R1013 DVDD.n4499 DVDD.n1073 4.5005
R1014 DVDD.n1076 DVDD.n1073 4.5005
R1015 DVDD.n4506 DVDD.n1073 4.5005
R1016 DVDD.n1077 DVDD.n1073 4.5005
R1017 DVDD.n4560 DVDD.n1083 4.5005
R1018 DVDD.n1083 DVDD.n1073 4.5005
R1019 DVDD.n4560 DVDD.n4500 4.5005
R1020 DVDD.n4500 DVDD.n1073 4.5005
R1021 DVDD.n4560 DVDD.n1082 4.5005
R1022 DVDD.n1082 DVDD.n1073 4.5005
R1023 DVDD.n4560 DVDD.n4501 4.5005
R1024 DVDD.n4501 DVDD.n1073 4.5005
R1025 DVDD.n4505 DVDD.n1073 4.5005
R1026 DVDD.n1078 DVDD.n1073 4.5005
R1027 DVDD.n4504 DVDD.n1073 4.5005
R1028 DVDD.n4560 DVDD.n1081 4.5005
R1029 DVDD.n1081 DVDD.n1073 4.5005
R1030 DVDD.n4560 DVDD.n4502 4.5005
R1031 DVDD.n4502 DVDD.n1073 4.5005
R1032 DVDD.n4560 DVDD.n1080 4.5005
R1033 DVDD.n1080 DVDD.n1073 4.5005
R1034 DVDD.n4560 DVDD.n4503 4.5005
R1035 DVDD.n4503 DVDD.n1073 4.5005
R1036 DVDD.n1079 DVDD.n1073 4.5005
R1037 DVDD.n4561 DVDD.n1073 4.5005
R1038 DVDD.n1073 DVDD.n1071 4.5005
R1039 DVDD.n4560 DVDD.n1071 4.5005
R1040 DVDD.n4561 DVDD.n4560 4.5005
R1041 DVDD.n4560 DVDD.n1079 4.5005
R1042 DVDD.n4560 DVDD.n4504 4.5005
R1043 DVDD.n4560 DVDD.n1078 4.5005
R1044 DVDD.n4560 DVDD.n4505 4.5005
R1045 DVDD.n4560 DVDD.n1077 4.5005
R1046 DVDD.n4560 DVDD.n4506 4.5005
R1047 DVDD.n4560 DVDD.n1076 4.5005
R1048 DVDD.n4560 DVDD.n4559 4.5005
R1049 DVDD.n4559 DVDD.n1073 4.5005
R1050 DVDD.n756 DVDD.n695 4.5005
R1051 DVDD.n756 DVDD.n702 4.5005
R1052 DVDD.n771 DVDD.n702 4.5005
R1053 DVDD.n771 DVDD.n695 4.5005
R1054 DVDD.n755 DVDD.n702 4.5005
R1055 DVDD.n755 DVDD.n695 4.5005
R1056 DVDD.n777 DVDD.n695 4.5005
R1057 DVDD.n779 DVDD.n695 4.5005
R1058 DVDD.n751 DVDD.n695 4.5005
R1059 DVDD.n784 DVDD.n702 4.5005
R1060 DVDD.n784 DVDD.n695 4.5005
R1061 DVDD.n786 DVDD.n702 4.5005
R1062 DVDD.n786 DVDD.n695 4.5005
R1063 DVDD.n749 DVDD.n702 4.5005
R1064 DVDD.n749 DVDD.n695 4.5005
R1065 DVDD.n791 DVDD.n702 4.5005
R1066 DVDD.n791 DVDD.n695 4.5005
R1067 DVDD.n747 DVDD.n695 4.5005
R1068 DVDD.n797 DVDD.n695 4.5005
R1069 DVDD.n799 DVDD.n695 4.5005
R1070 DVDD.n745 DVDD.n702 4.5005
R1071 DVDD.n745 DVDD.n695 4.5005
R1072 DVDD.n804 DVDD.n702 4.5005
R1073 DVDD.n804 DVDD.n695 4.5005
R1074 DVDD.n806 DVDD.n702 4.5005
R1075 DVDD.n806 DVDD.n695 4.5005
R1076 DVDD.n744 DVDD.n702 4.5005
R1077 DVDD.n744 DVDD.n695 4.5005
R1078 DVDD.n812 DVDD.n695 4.5005
R1079 DVDD.n814 DVDD.n695 4.5005
R1080 DVDD.n740 DVDD.n695 4.5005
R1081 DVDD.n740 DVDD.n702 4.5005
R1082 DVDD.n814 DVDD.n702 4.5005
R1083 DVDD.n812 DVDD.n702 4.5005
R1084 DVDD.n799 DVDD.n702 4.5005
R1085 DVDD.n797 DVDD.n702 4.5005
R1086 DVDD.n747 DVDD.n702 4.5005
R1087 DVDD.n751 DVDD.n702 4.5005
R1088 DVDD.n779 DVDD.n702 4.5005
R1089 DVDD.n777 DVDD.n702 4.5005
R1090 DVDD.n769 DVDD.n702 4.5005
R1091 DVDD.n769 DVDD.n695 4.5005
R1092 DVDD.n4939 DVDD.n672 4.5005
R1093 DVDD.n5004 DVDD.n4939 4.5005
R1094 DVDD.n5004 DVDD.n683 4.5005
R1095 DVDD.n683 DVDD.n672 4.5005
R1096 DVDD.n5004 DVDD.n4940 4.5005
R1097 DVDD.n4940 DVDD.n672 4.5005
R1098 DVDD.n675 DVDD.n672 4.5005
R1099 DVDD.n4948 DVDD.n672 4.5005
R1100 DVDD.n676 DVDD.n672 4.5005
R1101 DVDD.n5004 DVDD.n682 4.5005
R1102 DVDD.n682 DVDD.n672 4.5005
R1103 DVDD.n5004 DVDD.n4941 4.5005
R1104 DVDD.n4941 DVDD.n672 4.5005
R1105 DVDD.n5004 DVDD.n681 4.5005
R1106 DVDD.n681 DVDD.n672 4.5005
R1107 DVDD.n5004 DVDD.n4942 4.5005
R1108 DVDD.n4942 DVDD.n672 4.5005
R1109 DVDD.n4947 DVDD.n672 4.5005
R1110 DVDD.n677 DVDD.n672 4.5005
R1111 DVDD.n4946 DVDD.n672 4.5005
R1112 DVDD.n5004 DVDD.n680 4.5005
R1113 DVDD.n680 DVDD.n672 4.5005
R1114 DVDD.n5004 DVDD.n4943 4.5005
R1115 DVDD.n4943 DVDD.n672 4.5005
R1116 DVDD.n5004 DVDD.n679 4.5005
R1117 DVDD.n679 DVDD.n672 4.5005
R1118 DVDD.n5004 DVDD.n4944 4.5005
R1119 DVDD.n4944 DVDD.n672 4.5005
R1120 DVDD.n678 DVDD.n672 4.5005
R1121 DVDD.n4945 DVDD.n672 4.5005
R1122 DVDD.n5005 DVDD.n672 4.5005
R1123 DVDD.n5005 DVDD.n5004 4.5005
R1124 DVDD.n5004 DVDD.n4945 4.5005
R1125 DVDD.n5004 DVDD.n678 4.5005
R1126 DVDD.n5004 DVDD.n4946 4.5005
R1127 DVDD.n5004 DVDD.n677 4.5005
R1128 DVDD.n5004 DVDD.n4947 4.5005
R1129 DVDD.n5004 DVDD.n676 4.5005
R1130 DVDD.n5004 DVDD.n4948 4.5005
R1131 DVDD.n5004 DVDD.n675 4.5005
R1132 DVDD.n5004 DVDD.n5003 4.5005
R1133 DVDD.n5003 DVDD.n672 4.5005
R1134 DVDD.n5316 DVDD.n463 4.5005
R1135 DVDD.n5318 DVDD.n463 4.5005
R1136 DVDD.n5318 DVDD.n461 4.5005
R1137 DVDD.n5316 DVDD.n461 4.5005
R1138 DVDD.n5318 DVDD.n464 4.5005
R1139 DVDD.n5316 DVDD.n464 4.5005
R1140 DVDD.n5316 DVDD.n452 4.5005
R1141 DVDD.n5316 DVDD.n472 4.5005
R1142 DVDD.n5316 DVDD.n453 4.5005
R1143 DVDD.n5318 DVDD.n460 4.5005
R1144 DVDD.n5316 DVDD.n460 4.5005
R1145 DVDD.n5318 DVDD.n465 4.5005
R1146 DVDD.n5316 DVDD.n465 4.5005
R1147 DVDD.n5318 DVDD.n459 4.5005
R1148 DVDD.n5316 DVDD.n459 4.5005
R1149 DVDD.n5318 DVDD.n466 4.5005
R1150 DVDD.n5316 DVDD.n466 4.5005
R1151 DVDD.n5316 DVDD.n471 4.5005
R1152 DVDD.n5316 DVDD.n454 4.5005
R1153 DVDD.n5316 DVDD.n470 4.5005
R1154 DVDD.n5318 DVDD.n458 4.5005
R1155 DVDD.n5316 DVDD.n458 4.5005
R1156 DVDD.n5318 DVDD.n467 4.5005
R1157 DVDD.n5316 DVDD.n467 4.5005
R1158 DVDD.n5318 DVDD.n457 4.5005
R1159 DVDD.n5316 DVDD.n457 4.5005
R1160 DVDD.n5318 DVDD.n468 4.5005
R1161 DVDD.n5316 DVDD.n468 4.5005
R1162 DVDD.n5316 DVDD.n455 4.5005
R1163 DVDD.n5316 DVDD.n469 4.5005
R1164 DVDD.n5316 DVDD.n456 4.5005
R1165 DVDD.n5318 DVDD.n456 4.5005
R1166 DVDD.n5318 DVDD.n469 4.5005
R1167 DVDD.n5318 DVDD.n455 4.5005
R1168 DVDD.n5318 DVDD.n470 4.5005
R1169 DVDD.n5318 DVDD.n454 4.5005
R1170 DVDD.n5318 DVDD.n471 4.5005
R1171 DVDD.n5318 DVDD.n453 4.5005
R1172 DVDD.n5318 DVDD.n472 4.5005
R1173 DVDD.n5318 DVDD.n452 4.5005
R1174 DVDD.n5318 DVDD.n5317 4.5005
R1175 DVDD.n5317 DVDD.n5316 4.5005
R1176 DVDD.n5834 DVDD.n140 4.5005
R1177 DVDD.n143 DVDD.n140 4.5005
R1178 DVDD.n154 DVDD.n143 4.5005
R1179 DVDD.n5834 DVDD.n154 4.5005
R1180 DVDD.n156 DVDD.n143 4.5005
R1181 DVDD.n5834 DVDD.n156 4.5005
R1182 DVDD.n5834 DVDD.n153 4.5005
R1183 DVDD.n5834 DVDD.n157 4.5005
R1184 DVDD.n5834 DVDD.n152 4.5005
R1185 DVDD.n158 DVDD.n143 4.5005
R1186 DVDD.n5834 DVDD.n158 4.5005
R1187 DVDD.n151 DVDD.n143 4.5005
R1188 DVDD.n5834 DVDD.n151 4.5005
R1189 DVDD.n159 DVDD.n143 4.5005
R1190 DVDD.n5834 DVDD.n159 4.5005
R1191 DVDD.n150 DVDD.n143 4.5005
R1192 DVDD.n5834 DVDD.n150 4.5005
R1193 DVDD.n5834 DVDD.n160 4.5005
R1194 DVDD.n5834 DVDD.n149 4.5005
R1195 DVDD.n5834 DVDD.n161 4.5005
R1196 DVDD.n148 DVDD.n143 4.5005
R1197 DVDD.n5834 DVDD.n148 4.5005
R1198 DVDD.n162 DVDD.n143 4.5005
R1199 DVDD.n5834 DVDD.n162 4.5005
R1200 DVDD.n147 DVDD.n143 4.5005
R1201 DVDD.n5834 DVDD.n147 4.5005
R1202 DVDD.n163 DVDD.n143 4.5005
R1203 DVDD.n5834 DVDD.n163 4.5005
R1204 DVDD.n5834 DVDD.n146 4.5005
R1205 DVDD.n5834 DVDD.n5833 4.5005
R1206 DVDD.n5834 DVDD.n145 4.5005
R1207 DVDD.n145 DVDD.n143 4.5005
R1208 DVDD.n5833 DVDD.n143 4.5005
R1209 DVDD.n146 DVDD.n143 4.5005
R1210 DVDD.n161 DVDD.n143 4.5005
R1211 DVDD.n149 DVDD.n143 4.5005
R1212 DVDD.n160 DVDD.n143 4.5005
R1213 DVDD.n152 DVDD.n143 4.5005
R1214 DVDD.n157 DVDD.n143 4.5005
R1215 DVDD.n153 DVDD.n143 4.5005
R1216 DVDD.n5835 DVDD.n143 4.5005
R1217 DVDD.n5835 DVDD.n5834 4.5005
R1218 DVDD.n59 DVDD.n43 4.5005
R1219 DVDD.n5932 DVDD.n59 4.5005
R1220 DVDD.n57 DVDD.n43 4.5005
R1221 DVDD.n5932 DVDD.n57 4.5005
R1222 DVDD.n5932 DVDD.n60 4.5005
R1223 DVDD.n5932 DVDD.n56 4.5005
R1224 DVDD.n5932 DVDD.n61 4.5005
R1225 DVDD.n55 DVDD.n43 4.5005
R1226 DVDD.n5932 DVDD.n55 4.5005
R1227 DVDD.n62 DVDD.n43 4.5005
R1228 DVDD.n5932 DVDD.n62 4.5005
R1229 DVDD.n54 DVDD.n43 4.5005
R1230 DVDD.n5932 DVDD.n54 4.5005
R1231 DVDD.n63 DVDD.n43 4.5005
R1232 DVDD.n5932 DVDD.n63 4.5005
R1233 DVDD.n5932 DVDD.n53 4.5005
R1234 DVDD.n5932 DVDD.n64 4.5005
R1235 DVDD.n5932 DVDD.n52 4.5005
R1236 DVDD.n65 DVDD.n43 4.5005
R1237 DVDD.n5932 DVDD.n65 4.5005
R1238 DVDD.n51 DVDD.n43 4.5005
R1239 DVDD.n5932 DVDD.n51 4.5005
R1240 DVDD.n66 DVDD.n43 4.5005
R1241 DVDD.n5932 DVDD.n66 4.5005
R1242 DVDD.n50 DVDD.n43 4.5005
R1243 DVDD.n5932 DVDD.n50 4.5005
R1244 DVDD.n5932 DVDD.n67 4.5005
R1245 DVDD.n5932 DVDD.n49 4.5005
R1246 DVDD.n5932 DVDD.n68 4.5005
R1247 DVDD.n5563 DVDD.n5561 4.5005
R1248 DVDD.n5649 DVDD.n5561 4.5005
R1249 DVDD.n68 DVDD.n43 4.5005
R1250 DVDD.n5649 DVDD.n70 4.5005
R1251 DVDD.n5563 DVDD.n70 4.5005
R1252 DVDD.n5932 DVDD.n48 4.5005
R1253 DVDD.n48 DVDD.n43 4.5005
R1254 DVDD.n49 DVDD.n43 4.5005
R1255 DVDD.n67 DVDD.n43 4.5005
R1256 DVDD.n52 DVDD.n43 4.5005
R1257 DVDD.n64 DVDD.n43 4.5005
R1258 DVDD.n53 DVDD.n43 4.5005
R1259 DVDD.n61 DVDD.n43 4.5005
R1260 DVDD.n56 DVDD.n43 4.5005
R1261 DVDD.n60 DVDD.n43 4.5005
R1262 DVDD.n5931 DVDD.n43 4.5005
R1263 DVDD.n5932 DVDD.n5931 4.5005
R1264 DVDD.n5475 DVDD.n268 4.5005
R1265 DVDD.n271 DVDD.n268 4.5005
R1266 DVDD.n295 DVDD.n270 4.5005
R1267 DVDD.n308 DVDD.n295 4.5005
R1268 DVDD.n5472 DVDD.n308 4.5005
R1269 DVDD.n306 DVDD.n295 4.5005
R1270 DVDD.n5472 DVDD.n306 4.5005
R1271 DVDD.n309 DVDD.n295 4.5005
R1272 DVDD.n5472 DVDD.n309 4.5005
R1273 DVDD.n5472 DVDD.n305 4.5005
R1274 DVDD.n5472 DVDD.n310 4.5005
R1275 DVDD.n5472 DVDD.n304 4.5005
R1276 DVDD.n311 DVDD.n295 4.5005
R1277 DVDD.n5472 DVDD.n311 4.5005
R1278 DVDD.n303 DVDD.n295 4.5005
R1279 DVDD.n5472 DVDD.n303 4.5005
R1280 DVDD.n312 DVDD.n295 4.5005
R1281 DVDD.n5472 DVDD.n312 4.5005
R1282 DVDD.n302 DVDD.n295 4.5005
R1283 DVDD.n5472 DVDD.n302 4.5005
R1284 DVDD.n5472 DVDD.n313 4.5005
R1285 DVDD.n5472 DVDD.n301 4.5005
R1286 DVDD.n5472 DVDD.n314 4.5005
R1287 DVDD.n300 DVDD.n295 4.5005
R1288 DVDD.n5472 DVDD.n300 4.5005
R1289 DVDD.n315 DVDD.n295 4.5005
R1290 DVDD.n5472 DVDD.n315 4.5005
R1291 DVDD.n299 DVDD.n295 4.5005
R1292 DVDD.n5472 DVDD.n299 4.5005
R1293 DVDD.n5471 DVDD.n295 4.5005
R1294 DVDD.n5472 DVDD.n5471 4.5005
R1295 DVDD.n5472 DVDD.n298 4.5005
R1296 DVDD.n5472 DVDD.n272 4.5005
R1297 DVDD.n5472 DVDD.n270 4.5005
R1298 DVDD.n295 DVDD.n272 4.5005
R1299 DVDD.n298 DVDD.n295 4.5005
R1300 DVDD.n314 DVDD.n295 4.5005
R1301 DVDD.n301 DVDD.n295 4.5005
R1302 DVDD.n313 DVDD.n295 4.5005
R1303 DVDD.n304 DVDD.n295 4.5005
R1304 DVDD.n310 DVDD.n295 4.5005
R1305 DVDD.n305 DVDD.n295 4.5005
R1306 DVDD.n5475 DVDD.n5474 4.5005
R1307 DVDD.n5474 DVDD.n271 4.5005
R1308 DVDD.n5473 DVDD.n295 4.5005
R1309 DVDD.n5473 DVDD.n5472 4.5005
R1310 DVDD.n4698 DVDD.n4645 4.5005
R1311 DVDD.n4645 DVDD.n971 4.5005
R1312 DVDD.n4698 DVDD.n984 4.5005
R1313 DVDD.n984 DVDD.n971 4.5005
R1314 DVDD.n4698 DVDD.n4646 4.5005
R1315 DVDD.n4646 DVDD.n971 4.5005
R1316 DVDD.n4698 DVDD.n983 4.5005
R1317 DVDD.n983 DVDD.n971 4.5005
R1318 DVDD.n4698 DVDD.n4647 4.5005
R1319 DVDD.n4647 DVDD.n971 4.5005
R1320 DVDD.n4698 DVDD.n982 4.5005
R1321 DVDD.n982 DVDD.n971 4.5005
R1322 DVDD.n4698 DVDD.n4648 4.5005
R1323 DVDD.n4648 DVDD.n971 4.5005
R1324 DVDD.n4698 DVDD.n981 4.5005
R1325 DVDD.n981 DVDD.n971 4.5005
R1326 DVDD.n4698 DVDD.n4649 4.5005
R1327 DVDD.n4649 DVDD.n971 4.5005
R1328 DVDD.n4698 DVDD.n980 4.5005
R1329 DVDD.n980 DVDD.n971 4.5005
R1330 DVDD.n4698 DVDD.n4650 4.5005
R1331 DVDD.n4650 DVDD.n971 4.5005
R1332 DVDD.n4698 DVDD.n979 4.5005
R1333 DVDD.n979 DVDD.n971 4.5005
R1334 DVDD.n4698 DVDD.n4651 4.5005
R1335 DVDD.n4651 DVDD.n971 4.5005
R1336 DVDD.n4698 DVDD.n978 4.5005
R1337 DVDD.n978 DVDD.n971 4.5005
R1338 DVDD.n4698 DVDD.n4652 4.5005
R1339 DVDD.n4652 DVDD.n971 4.5005
R1340 DVDD.n4698 DVDD.n977 4.5005
R1341 DVDD.n977 DVDD.n971 4.5005
R1342 DVDD.n4698 DVDD.n4653 4.5005
R1343 DVDD.n4653 DVDD.n971 4.5005
R1344 DVDD.n4698 DVDD.n976 4.5005
R1345 DVDD.n976 DVDD.n971 4.5005
R1346 DVDD.n4698 DVDD.n4697 4.5005
R1347 DVDD.n4697 DVDD.n971 4.5005
R1348 DVDD.n31 DVDD.n18 4.5005
R1349 DVDD.n5954 DVDD.n18 4.5005
R1350 DVDD.n31 DVDD.n17 4.5005
R1351 DVDD.n5954 DVDD.n17 4.5005
R1352 DVDD.n31 DVDD.n19 4.5005
R1353 DVDD.n5954 DVDD.n19 4.5005
R1354 DVDD.n31 DVDD.n16 4.5005
R1355 DVDD.n5954 DVDD.n16 4.5005
R1356 DVDD.n31 DVDD.n20 4.5005
R1357 DVDD.n5954 DVDD.n20 4.5005
R1358 DVDD.n31 DVDD.n15 4.5005
R1359 DVDD.n5954 DVDD.n15 4.5005
R1360 DVDD.n31 DVDD.n21 4.5005
R1361 DVDD.n5954 DVDD.n21 4.5005
R1362 DVDD.n31 DVDD.n14 4.5005
R1363 DVDD.n5954 DVDD.n14 4.5005
R1364 DVDD.n31 DVDD.n22 4.5005
R1365 DVDD.n5954 DVDD.n22 4.5005
R1366 DVDD.n31 DVDD.n13 4.5005
R1367 DVDD.n5954 DVDD.n13 4.5005
R1368 DVDD.n31 DVDD.n23 4.5005
R1369 DVDD.n5954 DVDD.n23 4.5005
R1370 DVDD.n31 DVDD.n12 4.5005
R1371 DVDD.n5954 DVDD.n12 4.5005
R1372 DVDD.n31 DVDD.n24 4.5005
R1373 DVDD.n5954 DVDD.n24 4.5005
R1374 DVDD.n31 DVDD.n11 4.5005
R1375 DVDD.n5954 DVDD.n11 4.5005
R1376 DVDD.n31 DVDD.n25 4.5005
R1377 DVDD.n5954 DVDD.n25 4.5005
R1378 DVDD.n31 DVDD.n10 4.5005
R1379 DVDD.n5954 DVDD.n10 4.5005
R1380 DVDD.n31 DVDD.n26 4.5005
R1381 DVDD.n5954 DVDD.n26 4.5005
R1382 DVDD.n31 DVDD.n9 4.5005
R1383 DVDD.n5954 DVDD.n9 4.5005
R1384 DVDD.n31 DVDD.n27 4.5005
R1385 DVDD.n5954 DVDD.n27 4.5005
R1386 DVDD.n4387 DVDD.n1595 4.5005
R1387 DVDD.n4387 DVDD.n4386 4.5005
R1388 DVDD.n4386 DVDD.n1606 4.5005
R1389 DVDD.n4386 DVDD.n1609 4.5005
R1390 DVDD.n4386 DVDD.n1605 4.5005
R1391 DVDD.n4386 DVDD.n1611 4.5005
R1392 DVDD.n4386 DVDD.n1604 4.5005
R1393 DVDD.n4386 DVDD.n1613 4.5005
R1394 DVDD.n4386 DVDD.n1603 4.5005
R1395 DVDD.n4386 DVDD.n1615 4.5005
R1396 DVDD.n4386 DVDD.n1602 4.5005
R1397 DVDD.n4386 DVDD.n1617 4.5005
R1398 DVDD.n4386 DVDD.n1601 4.5005
R1399 DVDD.n4386 DVDD.n1619 4.5005
R1400 DVDD.n4386 DVDD.n1600 4.5005
R1401 DVDD.n4386 DVDD.n1621 4.5005
R1402 DVDD.n4386 DVDD.n1599 4.5005
R1403 DVDD.n4386 DVDD.n1623 4.5005
R1404 DVDD.n4386 DVDD.n1598 4.5005
R1405 DVDD.n4386 DVDD.n1625 4.5005
R1406 DVDD.n4386 DVDD.n1597 4.5005
R1407 DVDD.n4385 DVDD.n4383 4.5005
R1408 DVDD.n4386 DVDD.n4385 4.5005
R1409 DVDD.n4615 DVDD.n1047 4.5005
R1410 DVDD.n4615 DVDD.n1019 4.5005
R1411 DVDD.n1048 DVDD.n1005 4.5005
R1412 DVDD.n4615 DVDD.n1048 4.5005
R1413 DVDD.n1018 DVDD.n1005 4.5005
R1414 DVDD.n4615 DVDD.n1018 4.5005
R1415 DVDD.n1049 DVDD.n1005 4.5005
R1416 DVDD.n4615 DVDD.n1049 4.5005
R1417 DVDD.n1017 DVDD.n1005 4.5005
R1418 DVDD.n4615 DVDD.n1017 4.5005
R1419 DVDD.n4615 DVDD.n1050 4.5005
R1420 DVDD.n4615 DVDD.n1016 4.5005
R1421 DVDD.n4615 DVDD.n1051 4.5005
R1422 DVDD.n1015 DVDD.n1005 4.5005
R1423 DVDD.n4615 DVDD.n1015 4.5005
R1424 DVDD.n1052 DVDD.n1005 4.5005
R1425 DVDD.n4615 DVDD.n1052 4.5005
R1426 DVDD.n1014 DVDD.n1005 4.5005
R1427 DVDD.n4615 DVDD.n1014 4.5005
R1428 DVDD.n1053 DVDD.n1005 4.5005
R1429 DVDD.n4615 DVDD.n1053 4.5005
R1430 DVDD.n4615 DVDD.n1013 4.5005
R1431 DVDD.n4615 DVDD.n1054 4.5005
R1432 DVDD.n4615 DVDD.n1012 4.5005
R1433 DVDD.n1055 DVDD.n1005 4.5005
R1434 DVDD.n4615 DVDD.n1055 4.5005
R1435 DVDD.n1011 DVDD.n1005 4.5005
R1436 DVDD.n4615 DVDD.n1011 4.5005
R1437 DVDD.n1056 DVDD.n1005 4.5005
R1438 DVDD.n4615 DVDD.n1056 4.5005
R1439 DVDD.n1010 DVDD.n1005 4.5005
R1440 DVDD.n4615 DVDD.n1010 4.5005
R1441 DVDD.n4615 DVDD.n4614 4.5005
R1442 DVDD.n4614 DVDD.n1005 4.5005
R1443 DVDD.n1012 DVDD.n1005 4.5005
R1444 DVDD.n1054 DVDD.n1005 4.5005
R1445 DVDD.n1013 DVDD.n1005 4.5005
R1446 DVDD.n1051 DVDD.n1005 4.5005
R1447 DVDD.n1016 DVDD.n1005 4.5005
R1448 DVDD.n1050 DVDD.n1005 4.5005
R1449 DVDD.n1019 DVDD.n1005 4.5005
R1450 DVDD.n1047 DVDD.n1005 4.5005
R1451 DVDD.n4877 DVDD.n716 4.5005
R1452 DVDD.n4877 DVDD.n714 4.5005
R1453 DVDD.n4875 DVDD.n717 4.5005
R1454 DVDD.n4877 DVDD.n717 4.5005
R1455 DVDD.n4875 DVDD.n713 4.5005
R1456 DVDD.n4877 DVDD.n713 4.5005
R1457 DVDD.n4875 DVDD.n718 4.5005
R1458 DVDD.n4877 DVDD.n718 4.5005
R1459 DVDD.n4875 DVDD.n712 4.5005
R1460 DVDD.n4877 DVDD.n712 4.5005
R1461 DVDD.n4877 DVDD.n719 4.5005
R1462 DVDD.n4877 DVDD.n711 4.5005
R1463 DVDD.n4877 DVDD.n720 4.5005
R1464 DVDD.n4875 DVDD.n710 4.5005
R1465 DVDD.n4877 DVDD.n710 4.5005
R1466 DVDD.n4875 DVDD.n721 4.5005
R1467 DVDD.n4877 DVDD.n721 4.5005
R1468 DVDD.n4875 DVDD.n709 4.5005
R1469 DVDD.n4877 DVDD.n709 4.5005
R1470 DVDD.n4875 DVDD.n722 4.5005
R1471 DVDD.n4877 DVDD.n722 4.5005
R1472 DVDD.n4877 DVDD.n708 4.5005
R1473 DVDD.n4877 DVDD.n723 4.5005
R1474 DVDD.n4877 DVDD.n707 4.5005
R1475 DVDD.n4875 DVDD.n724 4.5005
R1476 DVDD.n4877 DVDD.n724 4.5005
R1477 DVDD.n4875 DVDD.n706 4.5005
R1478 DVDD.n4877 DVDD.n706 4.5005
R1479 DVDD.n4875 DVDD.n725 4.5005
R1480 DVDD.n4877 DVDD.n725 4.5005
R1481 DVDD.n4875 DVDD.n705 4.5005
R1482 DVDD.n4877 DVDD.n705 4.5005
R1483 DVDD.n4877 DVDD.n4876 4.5005
R1484 DVDD.n4876 DVDD.n4875 4.5005
R1485 DVDD.n4875 DVDD.n707 4.5005
R1486 DVDD.n4875 DVDD.n723 4.5005
R1487 DVDD.n4875 DVDD.n708 4.5005
R1488 DVDD.n4875 DVDD.n720 4.5005
R1489 DVDD.n4875 DVDD.n711 4.5005
R1490 DVDD.n4875 DVDD.n719 4.5005
R1491 DVDD.n4875 DVDD.n714 4.5005
R1492 DVDD.n4875 DVDD.n716 4.5005
R1493 DVDD.n5011 DVDD.n603 4.5005
R1494 DVDD.n606 DVDD.n603 4.5005
R1495 DVDD.n5012 DVDD.n617 4.5005
R1496 DVDD.n617 DVDD.n603 4.5005
R1497 DVDD.n5012 DVDD.n615 4.5005
R1498 DVDD.n615 DVDD.n603 4.5005
R1499 DVDD.n5012 DVDD.n618 4.5005
R1500 DVDD.n618 DVDD.n603 4.5005
R1501 DVDD.n5012 DVDD.n614 4.5005
R1502 DVDD.n614 DVDD.n603 4.5005
R1503 DVDD.n625 DVDD.n603 4.5005
R1504 DVDD.n607 DVDD.n603 4.5005
R1505 DVDD.n624 DVDD.n603 4.5005
R1506 DVDD.n5012 DVDD.n619 4.5005
R1507 DVDD.n619 DVDD.n603 4.5005
R1508 DVDD.n5012 DVDD.n613 4.5005
R1509 DVDD.n613 DVDD.n603 4.5005
R1510 DVDD.n5012 DVDD.n620 4.5005
R1511 DVDD.n620 DVDD.n603 4.5005
R1512 DVDD.n5012 DVDD.n612 4.5005
R1513 DVDD.n612 DVDD.n603 4.5005
R1514 DVDD.n608 DVDD.n603 4.5005
R1515 DVDD.n623 DVDD.n603 4.5005
R1516 DVDD.n609 DVDD.n603 4.5005
R1517 DVDD.n5012 DVDD.n621 4.5005
R1518 DVDD.n621 DVDD.n603 4.5005
R1519 DVDD.n5012 DVDD.n611 4.5005
R1520 DVDD.n611 DVDD.n603 4.5005
R1521 DVDD.n5012 DVDD.n622 4.5005
R1522 DVDD.n622 DVDD.n603 4.5005
R1523 DVDD.n5012 DVDD.n610 4.5005
R1524 DVDD.n610 DVDD.n603 4.5005
R1525 DVDD.n5013 DVDD.n603 4.5005
R1526 DVDD.n5013 DVDD.n5012 4.5005
R1527 DVDD.n5012 DVDD.n609 4.5005
R1528 DVDD.n5012 DVDD.n623 4.5005
R1529 DVDD.n5012 DVDD.n608 4.5005
R1530 DVDD.n5012 DVDD.n624 4.5005
R1531 DVDD.n5012 DVDD.n607 4.5005
R1532 DVDD.n5012 DVDD.n625 4.5005
R1533 DVDD.n5012 DVDD.n606 4.5005
R1534 DVDD.n5012 DVDD.n5011 4.5005
R1535 DVDD.n5242 DVDD.n556 4.5005
R1536 DVDD.n5242 DVDD.n495 4.5005
R1537 DVDD.n557 DVDD.n485 4.5005
R1538 DVDD.n5242 DVDD.n557 4.5005
R1539 DVDD.n494 DVDD.n485 4.5005
R1540 DVDD.n5242 DVDD.n494 4.5005
R1541 DVDD.n558 DVDD.n485 4.5005
R1542 DVDD.n5242 DVDD.n558 4.5005
R1543 DVDD.n493 DVDD.n485 4.5005
R1544 DVDD.n5242 DVDD.n493 4.5005
R1545 DVDD.n5242 DVDD.n559 4.5005
R1546 DVDD.n5242 DVDD.n492 4.5005
R1547 DVDD.n5242 DVDD.n560 4.5005
R1548 DVDD.n491 DVDD.n485 4.5005
R1549 DVDD.n5242 DVDD.n491 4.5005
R1550 DVDD.n561 DVDD.n485 4.5005
R1551 DVDD.n5242 DVDD.n561 4.5005
R1552 DVDD.n490 DVDD.n485 4.5005
R1553 DVDD.n5242 DVDD.n490 4.5005
R1554 DVDD.n562 DVDD.n485 4.5005
R1555 DVDD.n5242 DVDD.n562 4.5005
R1556 DVDD.n5242 DVDD.n489 4.5005
R1557 DVDD.n5242 DVDD.n563 4.5005
R1558 DVDD.n5242 DVDD.n488 4.5005
R1559 DVDD.n564 DVDD.n485 4.5005
R1560 DVDD.n5242 DVDD.n564 4.5005
R1561 DVDD.n487 DVDD.n485 4.5005
R1562 DVDD.n5242 DVDD.n487 4.5005
R1563 DVDD.n565 DVDD.n485 4.5005
R1564 DVDD.n5242 DVDD.n565 4.5005
R1565 DVDD.n486 DVDD.n485 4.5005
R1566 DVDD.n5242 DVDD.n486 4.5005
R1567 DVDD.n5242 DVDD.n5241 4.5005
R1568 DVDD.n5241 DVDD.n485 4.5005
R1569 DVDD.n488 DVDD.n485 4.5005
R1570 DVDD.n563 DVDD.n485 4.5005
R1571 DVDD.n489 DVDD.n485 4.5005
R1572 DVDD.n560 DVDD.n485 4.5005
R1573 DVDD.n492 DVDD.n485 4.5005
R1574 DVDD.n559 DVDD.n485 4.5005
R1575 DVDD.n495 DVDD.n485 4.5005
R1576 DVDD.n556 DVDD.n485 4.5005
R1577 DVDD.n169 DVDD.n166 4.5005
R1578 DVDD.n5784 DVDD.n169 4.5005
R1579 DVDD.n5783 DVDD.n181 4.5005
R1580 DVDD.n181 DVDD.n169 4.5005
R1581 DVDD.n5783 DVDD.n179 4.5005
R1582 DVDD.n179 DVDD.n169 4.5005
R1583 DVDD.n5783 DVDD.n182 4.5005
R1584 DVDD.n182 DVDD.n169 4.5005
R1585 DVDD.n5783 DVDD.n178 4.5005
R1586 DVDD.n178 DVDD.n169 4.5005
R1587 DVDD.n5782 DVDD.n169 4.5005
R1588 DVDD.n171 DVDD.n169 4.5005
R1589 DVDD.n189 DVDD.n169 4.5005
R1590 DVDD.n5783 DVDD.n183 4.5005
R1591 DVDD.n183 DVDD.n169 4.5005
R1592 DVDD.n5783 DVDD.n177 4.5005
R1593 DVDD.n177 DVDD.n169 4.5005
R1594 DVDD.n5783 DVDD.n184 4.5005
R1595 DVDD.n184 DVDD.n169 4.5005
R1596 DVDD.n5783 DVDD.n176 4.5005
R1597 DVDD.n176 DVDD.n169 4.5005
R1598 DVDD.n172 DVDD.n169 4.5005
R1599 DVDD.n188 DVDD.n169 4.5005
R1600 DVDD.n173 DVDD.n169 4.5005
R1601 DVDD.n5783 DVDD.n185 4.5005
R1602 DVDD.n185 DVDD.n169 4.5005
R1603 DVDD.n5783 DVDD.n175 4.5005
R1604 DVDD.n175 DVDD.n169 4.5005
R1605 DVDD.n5783 DVDD.n186 4.5005
R1606 DVDD.n186 DVDD.n169 4.5005
R1607 DVDD.n5783 DVDD.n174 4.5005
R1608 DVDD.n174 DVDD.n169 4.5005
R1609 DVDD.n187 DVDD.n169 4.5005
R1610 DVDD.n5783 DVDD.n187 4.5005
R1611 DVDD.n5783 DVDD.n173 4.5005
R1612 DVDD.n5783 DVDD.n188 4.5005
R1613 DVDD.n5783 DVDD.n172 4.5005
R1614 DVDD.n5783 DVDD.n189 4.5005
R1615 DVDD.n5783 DVDD.n171 4.5005
R1616 DVDD.n5783 DVDD.n5782 4.5005
R1617 DVDD.n5784 DVDD.n5783 4.5005
R1618 DVDD.n5783 DVDD.n166 4.5005
R1619 DVDD.n29 DVDD.n8 4.5005
R1620 DVDD.n31 DVDD.n8 4.5005
R1621 DVDD.n5954 DVDD.n8 4.5005
R1622 DVDD.n5953 DVDD.n29 4.5005
R1623 DVDD.n5953 DVDD.n31 4.5005
R1624 DVDD.n5954 DVDD.n5953 4.5005
R1625 DVDD.n5953 DVDD.n5952 4.5005
R1626 DVDD.n5952 DVDD.n27 4.5005
R1627 DVDD.n29 DVDD.n27 4.5005
R1628 DVDD.n5952 DVDD.n9 4.5005
R1629 DVDD.n29 DVDD.n9 4.5005
R1630 DVDD.n5952 DVDD.n26 4.5005
R1631 DVDD.n29 DVDD.n26 4.5005
R1632 DVDD.n29 DVDD.n10 4.5005
R1633 DVDD.n5952 DVDD.n10 4.5005
R1634 DVDD.n29 DVDD.n25 4.5005
R1635 DVDD.n5952 DVDD.n25 4.5005
R1636 DVDD.n29 DVDD.n11 4.5005
R1637 DVDD.n5952 DVDD.n11 4.5005
R1638 DVDD.n29 DVDD.n24 4.5005
R1639 DVDD.n5952 DVDD.n24 4.5005
R1640 DVDD.n5952 DVDD.n12 4.5005
R1641 DVDD.n29 DVDD.n12 4.5005
R1642 DVDD.n5952 DVDD.n23 4.5005
R1643 DVDD.n29 DVDD.n23 4.5005
R1644 DVDD.n5952 DVDD.n13 4.5005
R1645 DVDD.n29 DVDD.n13 4.5005
R1646 DVDD.n29 DVDD.n22 4.5005
R1647 DVDD.n5952 DVDD.n22 4.5005
R1648 DVDD.n29 DVDD.n14 4.5005
R1649 DVDD.n5952 DVDD.n14 4.5005
R1650 DVDD.n29 DVDD.n21 4.5005
R1651 DVDD.n5952 DVDD.n21 4.5005
R1652 DVDD.n29 DVDD.n15 4.5005
R1653 DVDD.n5952 DVDD.n15 4.5005
R1654 DVDD.n5952 DVDD.n20 4.5005
R1655 DVDD.n29 DVDD.n20 4.5005
R1656 DVDD.n5952 DVDD.n16 4.5005
R1657 DVDD.n29 DVDD.n16 4.5005
R1658 DVDD.n5952 DVDD.n19 4.5005
R1659 DVDD.n29 DVDD.n19 4.5005
R1660 DVDD.n29 DVDD.n17 4.5005
R1661 DVDD.n5952 DVDD.n17 4.5005
R1662 DVDD.n29 DVDD.n18 4.5005
R1663 DVDD.n5952 DVDD.n18 4.5005
R1664 DVDD.n5952 DVDD.n8 4.5005
R1665 DVDD.n4699 DVDD.n972 4.5005
R1666 DVDD.n4699 DVDD.n974 4.5005
R1667 DVDD.n4699 DVDD.n971 4.5005
R1668 DVDD.n4699 DVDD.n4698 4.5005
R1669 DVDD.n4645 DVDD.n972 4.5005
R1670 DVDD.n984 DVDD.n974 4.5005
R1671 DVDD.n984 DVDD.n972 4.5005
R1672 DVDD.n4646 DVDD.n974 4.5005
R1673 DVDD.n4646 DVDD.n972 4.5005
R1674 DVDD.n983 DVDD.n974 4.5005
R1675 DVDD.n983 DVDD.n972 4.5005
R1676 DVDD.n4647 DVDD.n974 4.5005
R1677 DVDD.n4647 DVDD.n972 4.5005
R1678 DVDD.n982 DVDD.n972 4.5005
R1679 DVDD.n4648 DVDD.n972 4.5005
R1680 DVDD.n981 DVDD.n972 4.5005
R1681 DVDD.n4649 DVDD.n974 4.5005
R1682 DVDD.n4649 DVDD.n972 4.5005
R1683 DVDD.n980 DVDD.n974 4.5005
R1684 DVDD.n980 DVDD.n972 4.5005
R1685 DVDD.n4650 DVDD.n974 4.5005
R1686 DVDD.n4650 DVDD.n972 4.5005
R1687 DVDD.n979 DVDD.n974 4.5005
R1688 DVDD.n979 DVDD.n972 4.5005
R1689 DVDD.n4651 DVDD.n972 4.5005
R1690 DVDD.n978 DVDD.n972 4.5005
R1691 DVDD.n4652 DVDD.n972 4.5005
R1692 DVDD.n977 DVDD.n974 4.5005
R1693 DVDD.n977 DVDD.n972 4.5005
R1694 DVDD.n4653 DVDD.n974 4.5005
R1695 DVDD.n4653 DVDD.n972 4.5005
R1696 DVDD.n976 DVDD.n974 4.5005
R1697 DVDD.n976 DVDD.n972 4.5005
R1698 DVDD.n4697 DVDD.n974 4.5005
R1699 DVDD.n4697 DVDD.n972 4.5005
R1700 DVDD.n4652 DVDD.n974 4.5005
R1701 DVDD.n978 DVDD.n974 4.5005
R1702 DVDD.n4651 DVDD.n974 4.5005
R1703 DVDD.n981 DVDD.n974 4.5005
R1704 DVDD.n4648 DVDD.n974 4.5005
R1705 DVDD.n982 DVDD.n974 4.5005
R1706 DVDD.n4645 DVDD.n974 4.5005
R1707 DVDD.n972 DVDD.n267 4.5005
R1708 DVDD.n974 DVDD.n267 4.5005
R1709 DVDD.n971 DVDD.n267 4.5005
R1710 DVDD.n4698 DVDD.n267 4.5005
R1711 DVDD.n4706 DVDD.n946 4.5005
R1712 DVDD.n946 DVDD.n914 4.5005
R1713 DVDD.n4706 DVDD.n945 4.5005
R1714 DVDD.n945 DVDD.n914 4.5005
R1715 DVDD.n4706 DVDD.n947 4.5005
R1716 DVDD.n947 DVDD.n914 4.5005
R1717 DVDD.n224 DVDD.n222 4.5005
R1718 DVDD.n5705 DVDD.n222 4.5005
R1719 DVDD.n224 DVDD.n219 4.5005
R1720 DVDD.n5705 DVDD.n219 4.5005
R1721 DVDD.n224 DVDD.n221 4.5005
R1722 DVDD.n5705 DVDD.n221 4.5005
R1723 DVDD.n4344 DVDD.n1627 4.5005
R1724 DVDD.n4344 DVDD.n4343 4.5005
R1725 DVDD.n4343 DVDD.n1638 4.5005
R1726 DVDD.n4343 DVDD.n1641 4.5005
R1727 DVDD.n4343 DVDD.n1637 4.5005
R1728 DVDD.n4343 DVDD.n1643 4.5005
R1729 DVDD.n4343 DVDD.n1636 4.5005
R1730 DVDD.n4343 DVDD.n1645 4.5005
R1731 DVDD.n4343 DVDD.n1635 4.5005
R1732 DVDD.n4343 DVDD.n1647 4.5005
R1733 DVDD.n4343 DVDD.n1634 4.5005
R1734 DVDD.n4343 DVDD.n1649 4.5005
R1735 DVDD.n4343 DVDD.n1633 4.5005
R1736 DVDD.n4343 DVDD.n1651 4.5005
R1737 DVDD.n4343 DVDD.n1632 4.5005
R1738 DVDD.n4343 DVDD.n1653 4.5005
R1739 DVDD.n4343 DVDD.n1631 4.5005
R1740 DVDD.n4343 DVDD.n1655 4.5005
R1741 DVDD.n4343 DVDD.n1630 4.5005
R1742 DVDD.n4343 DVDD.n1657 4.5005
R1743 DVDD.n4343 DVDD.n1629 4.5005
R1744 DVDD.n4342 DVDD.n4340 4.5005
R1745 DVDD.n4343 DVDD.n4342 4.5005
R1746 DVDD.n4744 DVDD.n894 4.5005
R1747 DVDD.n4742 DVDD.n893 4.5005
R1748 DVDD.n4744 DVDD.n893 4.5005
R1749 DVDD.n4742 DVDD.n895 4.5005
R1750 DVDD.n4744 DVDD.n895 4.5005
R1751 DVDD.n4742 DVDD.n892 4.5005
R1752 DVDD.n4744 DVDD.n892 4.5005
R1753 DVDD.n4743 DVDD.n4742 4.5005
R1754 DVDD.n4744 DVDD.n4743 4.5005
R1755 DVDD.n4742 DVDD.n894 4.5005
R1756 DVDD.n4773 DVDD.n737 4.5005
R1757 DVDD.n4771 DVDD.n736 4.5005
R1758 DVDD.n4773 DVDD.n736 4.5005
R1759 DVDD.n4771 DVDD.n738 4.5005
R1760 DVDD.n4773 DVDD.n738 4.5005
R1761 DVDD.n4771 DVDD.n735 4.5005
R1762 DVDD.n4773 DVDD.n735 4.5005
R1763 DVDD.n4772 DVDD.n4771 4.5005
R1764 DVDD.n4773 DVDD.n4772 4.5005
R1765 DVDD.n4771 DVDD.n737 4.5005
R1766 DVDD.n5019 DVDD.n584 4.5005
R1767 DVDD.n5020 DVDD.n592 4.5005
R1768 DVDD.n592 DVDD.n584 4.5005
R1769 DVDD.n5020 DVDD.n590 4.5005
R1770 DVDD.n590 DVDD.n584 4.5005
R1771 DVDD.n5020 DVDD.n593 4.5005
R1772 DVDD.n593 DVDD.n584 4.5005
R1773 DVDD.n5020 DVDD.n589 4.5005
R1774 DVDD.n589 DVDD.n584 4.5005
R1775 DVDD.n5020 DVDD.n5019 4.5005
R1776 DVDD.n5095 DVDD.n570 4.5005
R1777 DVDD.n5094 DVDD.n5086 4.5005
R1778 DVDD.n5086 DVDD.n570 4.5005
R1779 DVDD.n5094 DVDD.n573 4.5005
R1780 DVDD.n573 DVDD.n570 4.5005
R1781 DVDD.n5094 DVDD.n5093 4.5005
R1782 DVDD.n5093 DVDD.n570 4.5005
R1783 DVDD.n5094 DVDD.n572 4.5005
R1784 DVDD.n572 DVDD.n570 4.5005
R1785 DVDD.n5095 DVDD.n5094 4.5005
R1786 DVDD.n5733 DVDD.n193 4.5005
R1787 DVDD.n5734 DVDD.n196 4.5005
R1788 DVDD.n5734 DVDD.n5733 4.5005
R1789 DVDD.n5728 DVDD.n196 4.5005
R1790 DVDD.n5733 DVDD.n5728 4.5005
R1791 DVDD.n198 DVDD.n196 4.5005
R1792 DVDD.n5733 DVDD.n198 4.5005
R1793 DVDD.n5732 DVDD.n196 4.5005
R1794 DVDD.n5733 DVDD.n5732 4.5005
R1795 DVDD.n196 DVDD.n193 4.5005
R1796 DVDD.n5704 DVDD.n233 4.5005
R1797 DVDD.n5704 DVDD.n235 4.5005
R1798 DVDD.n241 DVDD.n235 4.5005
R1799 DVDD.n5702 DVDD.n235 4.5005
R1800 DVDD.n241 DVDD.n233 4.5005
R1801 DVDD.n5702 DVDD.n233 4.5005
R1802 DVDD.n5702 DVDD.n232 4.5005
R1803 DVDD.n241 DVDD.n232 4.5005
R1804 DVDD.n5704 DVDD.n232 4.5005
R1805 DVDD.n5702 DVDD.n236 4.5005
R1806 DVDD.n241 DVDD.n236 4.5005
R1807 DVDD.n5704 DVDD.n236 4.5005
R1808 DVDD.n5702 DVDD.n231 4.5005
R1809 DVDD.n241 DVDD.n231 4.5005
R1810 DVDD.n5704 DVDD.n231 4.5005
R1811 DVDD.n5704 DVDD.n237 4.5005
R1812 DVDD.n241 DVDD.n237 4.5005
R1813 DVDD.n5702 DVDD.n237 4.5005
R1814 DVDD.n5704 DVDD.n230 4.5005
R1815 DVDD.n241 DVDD.n230 4.5005
R1816 DVDD.n5702 DVDD.n230 4.5005
R1817 DVDD.n5704 DVDD.n238 4.5005
R1818 DVDD.n241 DVDD.n238 4.5005
R1819 DVDD.n5702 DVDD.n238 4.5005
R1820 DVDD.n5704 DVDD.n229 4.5005
R1821 DVDD.n241 DVDD.n229 4.5005
R1822 DVDD.n5702 DVDD.n229 4.5005
R1823 DVDD.n5702 DVDD.n239 4.5005
R1824 DVDD.n241 DVDD.n239 4.5005
R1825 DVDD.n5704 DVDD.n239 4.5005
R1826 DVDD.n5702 DVDD.n228 4.5005
R1827 DVDD.n241 DVDD.n228 4.5005
R1828 DVDD.n5704 DVDD.n228 4.5005
R1829 DVDD.n5703 DVDD.n5702 4.5005
R1830 DVDD.n5703 DVDD.n241 4.5005
R1831 DVDD.n5704 DVDD.n5703 4.5005
R1832 DVDD.n226 DVDD.n218 4.5005
R1833 DVDD.n224 DVDD.n218 4.5005
R1834 DVDD.n5705 DVDD.n218 4.5005
R1835 DVDD.n5707 DVDD.n221 4.5005
R1836 DVDD.n226 DVDD.n221 4.5005
R1837 DVDD.n5707 DVDD.n219 4.5005
R1838 DVDD.n226 DVDD.n219 4.5005
R1839 DVDD.n226 DVDD.n222 4.5005
R1840 DVDD.n5707 DVDD.n222 4.5005
R1841 DVDD.n5707 DVDD.n218 4.5005
R1842 DVDD.n5707 DVDD.n5706 4.5005
R1843 DVDD.n5706 DVDD.n226 4.5005
R1844 DVDD.n5706 DVDD.n224 4.5005
R1845 DVDD.n5706 DVDD.n5705 4.5005
R1846 DVDD.n943 DVDD.n920 4.5005
R1847 DVDD.n4708 DVDD.n920 4.5005
R1848 DVDD.n4710 DVDD.n920 4.5005
R1849 DVDD.n943 DVDD.n923 4.5005
R1850 DVDD.n4708 DVDD.n923 4.5005
R1851 DVDD.n4710 DVDD.n923 4.5005
R1852 DVDD.n4710 DVDD.n919 4.5005
R1853 DVDD.n4710 DVDD.n924 4.5005
R1854 DVDD.n4710 DVDD.n918 4.5005
R1855 DVDD.n943 DVDD.n925 4.5005
R1856 DVDD.n4708 DVDD.n925 4.5005
R1857 DVDD.n4710 DVDD.n925 4.5005
R1858 DVDD.n943 DVDD.n917 4.5005
R1859 DVDD.n4708 DVDD.n917 4.5005
R1860 DVDD.n4710 DVDD.n917 4.5005
R1861 DVDD.n943 DVDD.n926 4.5005
R1862 DVDD.n4708 DVDD.n926 4.5005
R1863 DVDD.n4710 DVDD.n926 4.5005
R1864 DVDD.n943 DVDD.n916 4.5005
R1865 DVDD.n4708 DVDD.n916 4.5005
R1866 DVDD.n4710 DVDD.n916 4.5005
R1867 DVDD.n4710 DVDD.n941 4.5005
R1868 DVDD.n4710 DVDD.n915 4.5005
R1869 DVDD.n4708 DVDD.n915 4.5005
R1870 DVDD.n943 DVDD.n915 4.5005
R1871 DVDD.n4708 DVDD.n941 4.5005
R1872 DVDD.n943 DVDD.n941 4.5005
R1873 DVDD.n4708 DVDD.n918 4.5005
R1874 DVDD.n943 DVDD.n918 4.5005
R1875 DVDD.n4708 DVDD.n924 4.5005
R1876 DVDD.n943 DVDD.n924 4.5005
R1877 DVDD.n4708 DVDD.n919 4.5005
R1878 DVDD.n943 DVDD.n919 4.5005
R1879 DVDD.n4710 DVDD.n4709 4.5005
R1880 DVDD.n4709 DVDD.n943 4.5005
R1881 DVDD.n4709 DVDD.n4708 4.5005
R1882 DVDD.n944 DVDD.n922 4.5005
R1883 DVDD.n944 DVDD.n910 4.5005
R1884 DVDD.n944 DVDD.n914 4.5005
R1885 DVDD.n4706 DVDD.n944 4.5005
R1886 DVDD.n4706 DVDD.n4705 4.5005
R1887 DVDD.n4705 DVDD.n914 4.5005
R1888 DVDD.n4705 DVDD.n922 4.5005
R1889 DVDD.n4705 DVDD.n910 4.5005
R1890 DVDD.n946 DVDD.n922 4.5005
R1891 DVDD.n946 DVDD.n910 4.5005
R1892 DVDD.n945 DVDD.n922 4.5005
R1893 DVDD.n945 DVDD.n910 4.5005
R1894 DVDD.n947 DVDD.n922 4.5005
R1895 DVDD.n947 DVDD.n910 4.5005
R1896 DVDD.n2796 DVDD.n2707 4.39376
R1897 DVDD.n3023 DVDD.n2077 4.29432
R1898 DVDD.n3314 DVDD.n3310 4.03391
R1899 DVDD.n2711 DVDD.t71 3.97738
R1900 DVDD.n3316 DVDD.n3240 3.90569
R1901 DVDD.n2712 DVDD.t154 3.75601
R1902 DVDD.n2734 DVDD.t117 3.75601
R1903 DVDD.t215 DVDD.n2013 3.6505
R1904 DVDD.t212 DVDD.n3661 3.6505
R1905 DVDD.t213 DVDD.n2010 3.6505
R1906 DVDD.t209 DVDD.n3658 3.6505
R1907 DVDD.n5489 DVDD.n5488 3.24952
R1908 DVDD.n5662 DVDD.n256 3.24952
R1909 DVDD.n3382 DVDD.n3238 3.1505
R1910 DVDD.n2767 DVDD.n2764 3.148
R1911 DVDD.n2759 DVDD.n2756 3.148
R1912 DVDD.n2764 DVDD.n2763 3.148
R1913 DVDD.n2759 DVDD.n2757 3.148
R1914 DVDD.n2764 DVDD.n2762 3.148
R1915 DVDD.n2759 DVDD.n2758 3.148
R1916 DVDD.n2764 DVDD.n2761 3.148
R1917 DVDD.n2759 DVDD.n2750 3.148
R1918 DVDD.n2739 DVDD.n2737 3.14761
R1919 DVDD.n2733 DVDD.n2732 3.14761
R1920 DVDD.n2783 DVDD.n2780 3.14761
R1921 DVDD.n2733 DVDD.n2731 3.14761
R1922 DVDD.n2783 DVDD.n2782 3.14761
R1923 DVDD.n2733 DVDD.n2730 3.14761
R1924 DVDD.n2783 DVDD.n2729 3.14761
R1925 DVDD.n2768 DVDD.n2766 2.98283
R1926 DVDD.n2768 DVDD.n2760 2.98283
R1927 DVDD.n2768 DVDD.n2747 2.98283
R1928 DVDD.n2741 DVDD.n2740 2.98283
R1929 DVDD.n2740 DVDD.n2724 2.98283
R1930 DVDD.n2765 DVDD.n2746 2.98283
R1931 DVDD.n2754 DVDD.n2746 2.98283
R1932 DVDD.n2738 DVDD.n2722 2.98283
R1933 DVDD.n2781 DVDD.n2727 2.98283
R1934 DVDD.n2776 DVDD.n2753 2.98283
R1935 DVDD.n3334 DVDD.n3315 2.94507
R1936 DVDD.n2013 DVDD.n2012 2.85774
R1937 DVDD.n3661 DVDD.n3660 2.85774
R1938 DVDD.n2010 DVDD.n2009 2.85774
R1939 DVDD.n3658 DVDD.n3657 2.85774
R1940 DVDD.n2711 DVDD.n2710 2.76877
R1941 DVDD.n3380 DVDD.n3238 2.76479
R1942 DVDD.n3332 DVDD.n3315 2.74405
R1943 DVDD.n4235 DVDD.n1710 2.69653
R1944 DVDD.n3024 DVDD.n3023 2.63997
R1945 DVDD.n2012 DVDD 2.57263
R1946 DVDD.n3660 DVDD 2.57263
R1947 DVDD.n2009 DVDD 2.57263
R1948 DVDD.n3657 DVDD 2.57263
R1949 DVDD.n3065 DVDD.n3064 2.56264
R1950 DVDD.n1936 DVDD.n1935 2.54396
R1951 DVDD.n2795 DVDD.n2794 2.52684
R1952 DVDD DVDD.n4200 2.51792
R1953 DVDD.n1885 DVDD 2.51792
R1954 DVDD.n3336 DVDD.n3335 2.42304
R1955 DVDD.n3379 DVDD.n3236 2.42304
R1956 DVDD.n3335 DVDD.n3312 2.38608
R1957 DVDD.n3379 DVDD.n3241 2.38608
R1958 DVDD.n3692 DVDD.t123 2.32044
R1959 DVDD.n3691 DVDD.t177 2.32044
R1960 DVDD.n5706 DVDD.n223 2.25251
R1961 DVDD.n961 DVDD.n944 2.25251
R1962 DVDD.n5919 DVDD.n5918 2.25174
R1963 DVDD.n5423 DVDD.n327 2.25174
R1964 DVDD.n5730 DVDD.n5729 2.2505
R1965 DVDD.n195 DVDD.n194 2.2505
R1966 DVDD.n5736 DVDD.n5735 2.2505
R1967 DVDD.n5738 DVDD.n5737 2.2505
R1968 DVDD.n5739 DVDD.n192 2.2505
R1969 DVDD.n5741 DVDD.n5740 2.2505
R1970 DVDD.n5743 DVDD.n5742 2.2505
R1971 DVDD.n5745 DVDD.n5744 2.2505
R1972 DVDD.n5747 DVDD.n5746 2.2505
R1973 DVDD.n5749 DVDD.n5748 2.2505
R1974 DVDD.n5751 DVDD.n5750 2.2505
R1975 DVDD.n5753 DVDD.n5752 2.2505
R1976 DVDD.n5755 DVDD.n5754 2.2505
R1977 DVDD.n5757 DVDD.n5756 2.2505
R1978 DVDD.n5759 DVDD.n5758 2.2505
R1979 DVDD.n5761 DVDD.n5760 2.2505
R1980 DVDD.n5763 DVDD.n5762 2.2505
R1981 DVDD.n5765 DVDD.n5764 2.2505
R1982 DVDD.n5767 DVDD.n5766 2.2505
R1983 DVDD.n5769 DVDD.n5768 2.2505
R1984 DVDD.n5771 DVDD.n5770 2.2505
R1985 DVDD.n5772 DVDD.n190 2.2505
R1986 DVDD.n5781 DVDD.n5780 2.2505
R1987 DVDD.n5779 DVDD.n191 2.2505
R1988 DVDD.n5778 DVDD.n5777 2.2505
R1989 DVDD.n5776 DVDD.n5775 2.2505
R1990 DVDD.n5774 DVDD.n5773 2.2505
R1991 DVDD.n168 DVDD.n167 2.2505
R1992 DVDD.n5786 DVDD.n5785 2.2505
R1993 DVDD.n5788 DVDD.n5787 2.2505
R1994 DVDD.n5789 DVDD.n165 2.2505
R1995 DVDD.n5791 DVDD.n5790 2.2505
R1996 DVDD.n5792 DVDD.n164 2.2505
R1997 DVDD.n5832 DVDD.n5831 2.2505
R1998 DVDD.n5830 DVDD.n5829 2.2505
R1999 DVDD.n5828 DVDD.n5827 2.2505
R2000 DVDD.n5826 DVDD.n5825 2.2505
R2001 DVDD.n5824 DVDD.n5823 2.2505
R2002 DVDD.n5822 DVDD.n5821 2.2505
R2003 DVDD.n5820 DVDD.n5819 2.2505
R2004 DVDD.n5818 DVDD.n5817 2.2505
R2005 DVDD.n5816 DVDD.n5815 2.2505
R2006 DVDD.n5814 DVDD.n5813 2.2505
R2007 DVDD.n5812 DVDD.n5811 2.2505
R2008 DVDD.n5810 DVDD.n5809 2.2505
R2009 DVDD.n5808 DVDD.n5807 2.2505
R2010 DVDD.n5806 DVDD.n5805 2.2505
R2011 DVDD.n5804 DVDD.n5803 2.2505
R2012 DVDD.n5802 DVDD.n5801 2.2505
R2013 DVDD.n5800 DVDD.n5799 2.2505
R2014 DVDD.n5798 DVDD.n5797 2.2505
R2015 DVDD.n5796 DVDD.n5795 2.2505
R2016 DVDD.n5794 DVDD.n5793 2.2505
R2017 DVDD.n142 DVDD.n141 2.2505
R2018 DVDD.n5837 DVDD.n5836 2.2505
R2019 DVDD.n5839 DVDD.n5838 2.2505
R2020 DVDD.n5840 DVDD.n139 2.2505
R2021 DVDD.n5842 DVDD.n5841 2.2505
R2022 DVDD.n5844 DVDD.n5843 2.2505
R2023 DVDD.n5846 DVDD.n5845 2.2505
R2024 DVDD.n5092 DVDD.n5091 2.2505
R2025 DVDD.n5090 DVDD.n5089 2.2505
R2026 DVDD.n5088 DVDD.n569 2.2505
R2027 DVDD.n5096 DVDD.n568 2.2505
R2028 DVDD.n5098 DVDD.n5097 2.2505
R2029 DVDD.n5099 DVDD.n566 2.2505
R2030 DVDD.n5240 DVDD.n5239 2.2505
R2031 DVDD.n5238 DVDD.n567 2.2505
R2032 DVDD.n5237 DVDD.n5236 2.2505
R2033 DVDD.n5235 DVDD.n5234 2.2505
R2034 DVDD.n5233 DVDD.n5232 2.2505
R2035 DVDD.n5231 DVDD.n5230 2.2505
R2036 DVDD.n5229 DVDD.n5228 2.2505
R2037 DVDD.n5227 DVDD.n5226 2.2505
R2038 DVDD.n5225 DVDD.n5224 2.2505
R2039 DVDD.n5223 DVDD.n5222 2.2505
R2040 DVDD.n5221 DVDD.n5220 2.2505
R2041 DVDD.n5219 DVDD.n5218 2.2505
R2042 DVDD.n5217 DVDD.n5216 2.2505
R2043 DVDD.n5215 DVDD.n5214 2.2505
R2044 DVDD.n5213 DVDD.n5212 2.2505
R2045 DVDD.n5211 DVDD.n5210 2.2505
R2046 DVDD.n5209 DVDD.n5208 2.2505
R2047 DVDD.n5207 DVDD.n5206 2.2505
R2048 DVDD.n5205 DVDD.n5204 2.2505
R2049 DVDD.n5203 DVDD.n5202 2.2505
R2050 DVDD.n5201 DVDD.n5200 2.2505
R2051 DVDD.n5199 DVDD.n5198 2.2505
R2052 DVDD.n5197 DVDD.n5196 2.2505
R2053 DVDD.n5195 DVDD.n5194 2.2505
R2054 DVDD.n5193 DVDD.n5100 2.2505
R2055 DVDD.n5192 DVDD.n5191 2.2505
R2056 DVDD.n5190 DVDD.n5189 2.2505
R2057 DVDD.n5188 DVDD.n5187 2.2505
R2058 DVDD.n5186 DVDD.n5185 2.2505
R2059 DVDD.n5184 DVDD.n5183 2.2505
R2060 DVDD.n5182 DVDD.n5181 2.2505
R2061 DVDD.n5180 DVDD.n5179 2.2505
R2062 DVDD.n5178 DVDD.n5177 2.2505
R2063 DVDD.n5176 DVDD.n5175 2.2505
R2064 DVDD.n5174 DVDD.n5173 2.2505
R2065 DVDD.n5172 DVDD.n5171 2.2505
R2066 DVDD.n5170 DVDD.n5169 2.2505
R2067 DVDD.n5168 DVDD.n5167 2.2505
R2068 DVDD.n5166 DVDD.n5165 2.2505
R2069 DVDD.n5164 DVDD.n5163 2.2505
R2070 DVDD.n5162 DVDD.n5161 2.2505
R2071 DVDD.n5160 DVDD.n5159 2.2505
R2072 DVDD.n5158 DVDD.n5157 2.2505
R2073 DVDD.n5156 DVDD.n5155 2.2505
R2074 DVDD.n5154 DVDD.n5153 2.2505
R2075 DVDD.n5152 DVDD.n5151 2.2505
R2076 DVDD.n5150 DVDD.n5149 2.2505
R2077 DVDD.n5148 DVDD.n473 2.2505
R2078 DVDD.n5147 DVDD.n474 2.2505
R2079 DVDD.n5146 DVDD.n5145 2.2505
R2080 DVDD.n5144 DVDD.n5101 2.2505
R2081 DVDD.n5143 DVDD.n5142 2.2505
R2082 DVDD.n5141 DVDD.n5140 2.2505
R2083 DVDD.n5138 DVDD.n5103 2.2505
R2084 DVDD.n598 DVDD.n597 2.2505
R2085 DVDD.n600 DVDD.n599 2.2505
R2086 DVDD.n601 DVDD.n594 2.2505
R2087 DVDD.n5018 DVDD.n5017 2.2505
R2088 DVDD.n5016 DVDD.n595 2.2505
R2089 DVDD.n5015 DVDD.n5014 2.2505
R2090 DVDD.n604 DVDD.n602 2.2505
R2091 DVDD.n629 DVDD.n628 2.2505
R2092 DVDD.n631 DVDD.n630 2.2505
R2093 DVDD.n633 DVDD.n632 2.2505
R2094 DVDD.n635 DVDD.n634 2.2505
R2095 DVDD.n637 DVDD.n636 2.2505
R2096 DVDD.n639 DVDD.n638 2.2505
R2097 DVDD.n641 DVDD.n640 2.2505
R2098 DVDD.n643 DVDD.n642 2.2505
R2099 DVDD.n645 DVDD.n644 2.2505
R2100 DVDD.n647 DVDD.n646 2.2505
R2101 DVDD.n649 DVDD.n648 2.2505
R2102 DVDD.n651 DVDD.n650 2.2505
R2103 DVDD.n653 DVDD.n652 2.2505
R2104 DVDD.n655 DVDD.n654 2.2505
R2105 DVDD.n657 DVDD.n656 2.2505
R2106 DVDD.n659 DVDD.n658 2.2505
R2107 DVDD.n661 DVDD.n660 2.2505
R2108 DVDD.n663 DVDD.n662 2.2505
R2109 DVDD.n665 DVDD.n664 2.2505
R2110 DVDD.n667 DVDD.n666 2.2505
R2111 DVDD.n669 DVDD.n668 2.2505
R2112 DVDD.n670 DVDD.n626 2.2505
R2113 DVDD.n5010 DVDD.n5009 2.2505
R2114 DVDD.n5008 DVDD.n627 2.2505
R2115 DVDD.n5007 DVDD.n5006 2.2505
R2116 DVDD.n673 DVDD.n671 2.2505
R2117 DVDD.n4951 DVDD.n4950 2.2505
R2118 DVDD.n4953 DVDD.n4952 2.2505
R2119 DVDD.n4955 DVDD.n4954 2.2505
R2120 DVDD.n4957 DVDD.n4956 2.2505
R2121 DVDD.n4959 DVDD.n4958 2.2505
R2122 DVDD.n4961 DVDD.n4960 2.2505
R2123 DVDD.n4963 DVDD.n4962 2.2505
R2124 DVDD.n4965 DVDD.n4964 2.2505
R2125 DVDD.n4967 DVDD.n4966 2.2505
R2126 DVDD.n4969 DVDD.n4968 2.2505
R2127 DVDD.n4971 DVDD.n4970 2.2505
R2128 DVDD.n4973 DVDD.n4972 2.2505
R2129 DVDD.n4975 DVDD.n4974 2.2505
R2130 DVDD.n4977 DVDD.n4976 2.2505
R2131 DVDD.n4979 DVDD.n4978 2.2505
R2132 DVDD.n4981 DVDD.n4980 2.2505
R2133 DVDD.n4983 DVDD.n4982 2.2505
R2134 DVDD.n4985 DVDD.n4984 2.2505
R2135 DVDD.n4987 DVDD.n4986 2.2505
R2136 DVDD.n4989 DVDD.n4988 2.2505
R2137 DVDD.n4990 DVDD.n4949 2.2505
R2138 DVDD.n5002 DVDD.n5001 2.2505
R2139 DVDD.n5000 DVDD.n4999 2.2505
R2140 DVDD.n4998 DVDD.n4991 2.2505
R2141 DVDD.n4997 DVDD.n4996 2.2505
R2142 DVDD.n4995 DVDD.n4994 2.2505
R2143 DVDD.n4993 DVDD.n4992 2.2505
R2144 DVDD.n877 DVDD.n876 2.2505
R2145 DVDD.n875 DVDD.n874 2.2505
R2146 DVDD.n873 DVDD.n872 2.2505
R2147 DVDD.n871 DVDD.n870 2.2505
R2148 DVDD.n869 DVDD.n868 2.2505
R2149 DVDD.n867 DVDD.n726 2.2505
R2150 DVDD.n866 DVDD.n727 2.2505
R2151 DVDD.n865 DVDD.n864 2.2505
R2152 DVDD.n863 DVDD.n862 2.2505
R2153 DVDD.n861 DVDD.n860 2.2505
R2154 DVDD.n859 DVDD.n858 2.2505
R2155 DVDD.n857 DVDD.n856 2.2505
R2156 DVDD.n855 DVDD.n854 2.2505
R2157 DVDD.n853 DVDD.n852 2.2505
R2158 DVDD.n851 DVDD.n850 2.2505
R2159 DVDD.n849 DVDD.n848 2.2505
R2160 DVDD.n847 DVDD.n846 2.2505
R2161 DVDD.n845 DVDD.n844 2.2505
R2162 DVDD.n843 DVDD.n842 2.2505
R2163 DVDD.n841 DVDD.n840 2.2505
R2164 DVDD.n839 DVDD.n838 2.2505
R2165 DVDD.n837 DVDD.n836 2.2505
R2166 DVDD.n835 DVDD.n834 2.2505
R2167 DVDD.n833 DVDD.n832 2.2505
R2168 DVDD.n831 DVDD.n830 2.2505
R2169 DVDD.n829 DVDD.n828 2.2505
R2170 DVDD.n827 DVDD.n826 2.2505
R2171 DVDD.n825 DVDD.n824 2.2505
R2172 DVDD.n823 DVDD.n822 2.2505
R2173 DVDD.n821 DVDD.n820 2.2505
R2174 DVDD.n819 DVDD.n739 2.2505
R2175 DVDD.n818 DVDD.n817 2.2505
R2176 DVDD.n816 DVDD.n815 2.2505
R2177 DVDD.n813 DVDD.n741 2.2505
R2178 DVDD.n811 DVDD.n810 2.2505
R2179 DVDD.n809 DVDD.n742 2.2505
R2180 DVDD.n808 DVDD.n807 2.2505
R2181 DVDD.n805 DVDD.n743 2.2505
R2182 DVDD.n803 DVDD.n802 2.2505
R2183 DVDD.n801 DVDD.n800 2.2505
R2184 DVDD.n798 DVDD.n746 2.2505
R2185 DVDD.n796 DVDD.n795 2.2505
R2186 DVDD.n794 DVDD.n793 2.2505
R2187 DVDD.n792 DVDD.n748 2.2505
R2188 DVDD.n790 DVDD.n789 2.2505
R2189 DVDD.n788 DVDD.n787 2.2505
R2190 DVDD.n785 DVDD.n750 2.2505
R2191 DVDD.n783 DVDD.n782 2.2505
R2192 DVDD.n781 DVDD.n780 2.2505
R2193 DVDD.n778 DVDD.n752 2.2505
R2194 DVDD.n776 DVDD.n775 2.2505
R2195 DVDD.n774 DVDD.n753 2.2505
R2196 DVDD.n773 DVDD.n772 2.2505
R2197 DVDD.n770 DVDD.n754 2.2505
R2198 DVDD.n768 DVDD.n767 2.2505
R2199 DVDD.n766 DVDD.n765 2.2505
R2200 DVDD.n764 DVDD.n757 2.2505
R2201 DVDD.n763 DVDD.n762 2.2505
R2202 DVDD.n761 DVDD.n760 2.2505
R2203 DVDD.n759 DVDD.n758 2.2505
R2204 DVDD.n1060 DVDD.n1059 2.2505
R2205 DVDD.n1062 DVDD.n1061 2.2505
R2206 DVDD.n1064 DVDD.n1063 2.2505
R2207 DVDD.n1066 DVDD.n1065 2.2505
R2208 DVDD.n1068 DVDD.n1067 2.2505
R2209 DVDD.n1069 DVDD.n1057 2.2505
R2210 DVDD.n4613 DVDD.n4612 2.2505
R2211 DVDD.n4611 DVDD.n1058 2.2505
R2212 DVDD.n4610 DVDD.n4609 2.2505
R2213 DVDD.n4608 DVDD.n4607 2.2505
R2214 DVDD.n4606 DVDD.n4605 2.2505
R2215 DVDD.n4604 DVDD.n4603 2.2505
R2216 DVDD.n4602 DVDD.n4601 2.2505
R2217 DVDD.n4600 DVDD.n4599 2.2505
R2218 DVDD.n4598 DVDD.n4597 2.2505
R2219 DVDD.n4596 DVDD.n4595 2.2505
R2220 DVDD.n4594 DVDD.n4593 2.2505
R2221 DVDD.n4592 DVDD.n4591 2.2505
R2222 DVDD.n4590 DVDD.n4589 2.2505
R2223 DVDD.n4588 DVDD.n4587 2.2505
R2224 DVDD.n4586 DVDD.n4585 2.2505
R2225 DVDD.n4584 DVDD.n4583 2.2505
R2226 DVDD.n4582 DVDD.n4581 2.2505
R2227 DVDD.n4580 DVDD.n4579 2.2505
R2228 DVDD.n4578 DVDD.n4577 2.2505
R2229 DVDD.n4576 DVDD.n4575 2.2505
R2230 DVDD.n4574 DVDD.n4573 2.2505
R2231 DVDD.n4572 DVDD.n4571 2.2505
R2232 DVDD.n4570 DVDD.n4569 2.2505
R2233 DVDD.n4568 DVDD.n4567 2.2505
R2234 DVDD.n4566 DVDD.n1070 2.2505
R2235 DVDD.n4565 DVDD.n4564 2.2505
R2236 DVDD.n4563 DVDD.n4562 2.2505
R2237 DVDD.n1074 DVDD.n1072 2.2505
R2238 DVDD.n4509 DVDD.n4508 2.2505
R2239 DVDD.n4511 DVDD.n4510 2.2505
R2240 DVDD.n4513 DVDD.n4512 2.2505
R2241 DVDD.n4515 DVDD.n4514 2.2505
R2242 DVDD.n4517 DVDD.n4516 2.2505
R2243 DVDD.n4519 DVDD.n4518 2.2505
R2244 DVDD.n4521 DVDD.n4520 2.2505
R2245 DVDD.n4523 DVDD.n4522 2.2505
R2246 DVDD.n4525 DVDD.n4524 2.2505
R2247 DVDD.n4527 DVDD.n4526 2.2505
R2248 DVDD.n4529 DVDD.n4528 2.2505
R2249 DVDD.n4531 DVDD.n4530 2.2505
R2250 DVDD.n4533 DVDD.n4532 2.2505
R2251 DVDD.n4535 DVDD.n4534 2.2505
R2252 DVDD.n4537 DVDD.n4536 2.2505
R2253 DVDD.n4539 DVDD.n4538 2.2505
R2254 DVDD.n4541 DVDD.n4540 2.2505
R2255 DVDD.n4543 DVDD.n4542 2.2505
R2256 DVDD.n4545 DVDD.n4544 2.2505
R2257 DVDD.n4546 DVDD.n4507 2.2505
R2258 DVDD.n4558 DVDD.n4557 2.2505
R2259 DVDD.n4556 DVDD.n4555 2.2505
R2260 DVDD.n4554 DVDD.n4547 2.2505
R2261 DVDD.n4553 DVDD.n4552 2.2505
R2262 DVDD.n4551 DVDD.n4550 2.2505
R2263 DVDD.n4549 DVDD.n4548 2.2505
R2264 DVDD.n3663 DVDD.n3659 2.2505
R2265 DVDD.n2015 DVDD.n2011 2.2505
R2266 DVDD.n3663 DVDD.n3662 2.2505
R2267 DVDD.n2015 DVDD.n2014 2.2505
R2268 DVDD.n3263 DVDD.n3258 2.2505
R2269 DVDD.n3387 DVDD.n3386 2.2505
R2270 DVDD.n3385 DVDD.n3233 2.2505
R2271 DVDD.n3259 DVDD.n3235 2.2505
R2272 DVDD.n3265 DVDD.n3264 2.2505
R2273 DVDD.n3356 DVDD.n3355 2.2505
R2274 DVDD.n3339 DVDD.n3308 2.2505
R2275 DVDD.n3280 DVDD.n3279 2.2505
R2276 DVDD.n3364 DVDD.n3363 2.2505
R2277 DVDD.n3366 DVDD.n3365 2.2505
R2278 DVDD.n3344 DVDD.n3099 2.2505
R2279 DVDD.n3369 DVDD.n3368 2.2505
R2280 DVDD.n3296 DVDD.n3272 2.2505
R2281 DVDD.n3361 DVDD.n3294 2.2505
R2282 DVDD.n3358 DVDD.n3299 2.2505
R2283 DVDD.n3340 DVDD.n3098 2.2505
R2284 DVDD.n3351 DVDD.n3099 2.2505
R2285 DVDD.n3358 DVDD.n3357 2.2505
R2286 DVDD.n3368 DVDD.n3367 2.2505
R2287 DVDD.n3296 DVDD.n3277 2.2505
R2288 DVDD.n3362 DVDD.n3361 2.2505
R2289 DVDD.n3309 DVDD.n3098 2.2505
R2290 DVDD.n3398 DVDD.n3221 2.2505
R2291 DVDD.n3372 DVDD.n3371 2.2505
R2292 DVDD.n3268 DVDD.n3267 2.2505
R2293 DVDD.n3261 DVDD.n3227 2.2505
R2294 DVDD.n3390 DVDD.n3389 2.2505
R2295 DVDD.n3391 DVDD.n3096 2.2505
R2296 DVDD.n3267 DVDD.n3266 2.2505
R2297 DVDD.n3262 DVDD.n3261 2.2505
R2298 DVDD.n3389 DVDD.n3388 2.2505
R2299 DVDD.n3234 DVDD.n3096 2.2505
R2300 DVDD.n3398 DVDD.n3397 2.2505
R2301 DVDD.n3372 DVDD.n3243 2.2505
R2302 DVDD.n1391 DVDD.n1390 2.2505
R2303 DVDD.n1315 DVDD.n1314 2.2505
R2304 DVDD.n5501 DVDD.n225 2.2505
R2305 DVDD.n5503 DVDD.n5502 2.2505
R2306 DVDD.n5506 DVDD.n5505 2.2505
R2307 DVDD.n5508 DVDD.n5507 2.2505
R2308 DVDD.n5510 DVDD.n5509 2.2505
R2309 DVDD.n5512 DVDD.n5511 2.2505
R2310 DVDD.n5513 DVDD.n28 2.2505
R2311 DVDD.n5514 DVDD.n30 2.2505
R2312 DVDD.n5516 DVDD.n5515 2.2505
R2313 DVDD.n5518 DVDD.n5517 2.2505
R2314 DVDD.n5520 DVDD.n5519 2.2505
R2315 DVDD.n5522 DVDD.n5521 2.2505
R2316 DVDD.n5524 DVDD.n5523 2.2505
R2317 DVDD.n5526 DVDD.n5525 2.2505
R2318 DVDD.n5528 DVDD.n5527 2.2505
R2319 DVDD.n5530 DVDD.n5529 2.2505
R2320 DVDD.n5532 DVDD.n5531 2.2505
R2321 DVDD.n5534 DVDD.n5533 2.2505
R2322 DVDD.n5536 DVDD.n5535 2.2505
R2323 DVDD.n5539 DVDD.n5538 2.2505
R2324 DVDD.n5541 DVDD.n5540 2.2505
R2325 DVDD.n5543 DVDD.n5542 2.2505
R2326 DVDD.n5545 DVDD.n5544 2.2505
R2327 DVDD.n5547 DVDD.n5546 2.2505
R2328 DVDD.n5549 DVDD.n5548 2.2505
R2329 DVDD.n5551 DVDD.n5550 2.2505
R2330 DVDD.n5553 DVDD.n5552 2.2505
R2331 DVDD.n5555 DVDD.n5554 2.2505
R2332 DVDD.n5557 DVDD.n5556 2.2505
R2333 DVDD.n5559 DVDD.n5558 2.2505
R2334 DVDD.n5657 DVDD.n5656 2.2505
R2335 DVDD.n5655 DVDD.n5560 2.2505
R2336 DVDD.n5654 DVDD.n5653 2.2505
R2337 DVDD.n5652 DVDD.n5651 2.2505
R2338 DVDD.n5565 DVDD.n5562 2.2505
R2339 DVDD.n5610 DVDD.n5609 2.2505
R2340 DVDD.n5647 DVDD.n5646 2.2505
R2341 DVDD.n5645 DVDD.n5644 2.2505
R2342 DVDD.n5643 DVDD.n5642 2.2505
R2343 DVDD.n5641 DVDD.n5640 2.2505
R2344 DVDD.n5639 DVDD.n5638 2.2505
R2345 DVDD.n5637 DVDD.n5636 2.2505
R2346 DVDD.n5635 DVDD.n5634 2.2505
R2347 DVDD.n5633 DVDD.n5632 2.2505
R2348 DVDD.n5629 DVDD.n5570 2.2505
R2349 DVDD.n5628 DVDD.n5627 2.2505
R2350 DVDD.n5626 DVDD.n5625 2.2505
R2351 DVDD.n5624 DVDD.n5623 2.2505
R2352 DVDD.n5622 DVDD.n5621 2.2505
R2353 DVDD.n5620 DVDD.n5619 2.2505
R2354 DVDD.n5618 DVDD.n5617 2.2505
R2355 DVDD.n5616 DVDD.n5615 2.2505
R2356 DVDD.n5614 DVDD.n5613 2.2505
R2357 DVDD.n5612 DVDD.n5611 2.2505
R2358 DVDD.n72 DVDD.n71 2.2505
R2359 DVDD.n5930 DVDD.n5929 2.2505
R2360 DVDD.n5928 DVDD.n5927 2.2505
R2361 DVDD.n5926 DVDD.n73 2.2505
R2362 DVDD.n5925 DVDD.n5924 2.2505
R2363 DVDD.n5923 DVDD.n5922 2.2505
R2364 DVDD.n78 DVDD.n75 2.2505
R2365 DVDD.n86 DVDD.n83 2.2505
R2366 DVDD.n4704 DVDD.n4703 2.2505
R2367 DVDD.n969 DVDD.n948 2.2505
R2368 DVDD.n968 DVDD.n967 2.2505
R2369 DVDD.n965 DVDD.n964 2.2505
R2370 DVDD.n963 DVDD.n962 2.2505
R2371 DVDD.n4702 DVDD.n949 2.2505
R2372 DVDD.n4701 DVDD.n4700 2.2505
R2373 DVDD.n973 DVDD.n970 2.2505
R2374 DVDD.n5483 DVDD.n5482 2.2505
R2375 DVDD.n4644 DVDD.n265 2.2505
R2376 DVDD.n4657 DVDD.n4656 2.2505
R2377 DVDD.n4659 DVDD.n4658 2.2505
R2378 DVDD.n4661 DVDD.n4660 2.2505
R2379 DVDD.n4663 DVDD.n4662 2.2505
R2380 DVDD.n4665 DVDD.n4664 2.2505
R2381 DVDD.n4667 DVDD.n4666 2.2505
R2382 DVDD.n4669 DVDD.n4668 2.2505
R2383 DVDD.n4671 DVDD.n4670 2.2505
R2384 DVDD.n4673 DVDD.n4672 2.2505
R2385 DVDD.n4675 DVDD.n4674 2.2505
R2386 DVDD.n4678 DVDD.n4677 2.2505
R2387 DVDD.n4680 DVDD.n4679 2.2505
R2388 DVDD.n4682 DVDD.n4681 2.2505
R2389 DVDD.n4684 DVDD.n4683 2.2505
R2390 DVDD.n4686 DVDD.n4685 2.2505
R2391 DVDD.n4688 DVDD.n4687 2.2505
R2392 DVDD.n4690 DVDD.n4689 2.2505
R2393 DVDD.n4692 DVDD.n4691 2.2505
R2394 DVDD.n4694 DVDD.n4693 2.2505
R2395 DVDD.n4696 DVDD.n4695 2.2505
R2396 DVDD.n4655 DVDD.n4654 2.2505
R2397 DVDD.n5481 DVDD.n266 2.2505
R2398 DVDD.n5480 DVDD.n5479 2.2505
R2399 DVDD.n5478 DVDD.n5477 2.2505
R2400 DVDD.n5433 DVDD.n294 2.2505
R2401 DVDD.n5432 DVDD.n296 2.2505
R2402 DVDD.n5435 DVDD.n5434 2.2505
R2403 DVDD.n5437 DVDD.n5436 2.2505
R2404 DVDD.n5439 DVDD.n5438 2.2505
R2405 DVDD.n5441 DVDD.n5440 2.2505
R2406 DVDD.n5443 DVDD.n5442 2.2505
R2407 DVDD.n5445 DVDD.n5444 2.2505
R2408 DVDD.n5447 DVDD.n5446 2.2505
R2409 DVDD.n5449 DVDD.n5448 2.2505
R2410 DVDD.n5451 DVDD.n5450 2.2505
R2411 DVDD.n5453 DVDD.n5452 2.2505
R2412 DVDD.n5454 DVDD.n279 2.2505
R2413 DVDD.n5458 DVDD.n5457 2.2505
R2414 DVDD.n5460 DVDD.n5459 2.2505
R2415 DVDD.n5462 DVDD.n5461 2.2505
R2416 DVDD.n5464 DVDD.n5463 2.2505
R2417 DVDD.n5466 DVDD.n5465 2.2505
R2418 DVDD.n5468 DVDD.n5467 2.2505
R2419 DVDD.n5470 DVDD.n5469 2.2505
R2420 DVDD.n319 DVDD.n316 2.2505
R2421 DVDD.n318 DVDD.n317 2.2505
R2422 DVDD.n274 DVDD.n269 2.2505
R2423 DVDD.n5431 DVDD.n5430 2.2505
R2424 DVDD.n5429 DVDD.n320 2.2505
R2425 DVDD.n5425 DVDD.n5424 2.2505
R2426 DVDD.n332 DVDD.n331 2.2505
R2427 DVDD.n330 DVDD.n323 2.2505
R2428 DVDD.n351 DVDD.n341 2.24971
R2429 DVDD.n5914 DVDD.n87 2.24971
R2430 DVDD.n5417 DVDD.n340 2.24971
R2431 DVDD.n106 DVDD.n94 2.24971
R2432 DVDD.n1573 DVDD.n1204 2.24621
R2433 DVDD.n1573 DVDD.n1203 2.24621
R2434 DVDD.n1573 DVDD.n1191 2.24621
R2435 DVDD.n1574 DVDD.n1573 2.24621
R2436 DVDD.n1201 DVDD.n1192 2.24621
R2437 DVDD.n1198 DVDD.n1192 2.24621
R2438 DVDD.n3417 DVDD.n3412 2.24442
R2439 DVDD.n3413 DVDD.n3209 2.24442
R2440 DVDD.n3113 DVDD.n3112 2.24442
R2441 DVDD.n3123 DVDD.n3110 2.24442
R2442 DVDD.n2843 DVDD.n2842 2.24442
R2443 DVDD.n2839 DVDD.n2694 2.24442
R2444 DVDD.n2800 DVDD.n2701 2.24405
R2445 DVDD.n2801 DVDD.n2702 2.24405
R2446 DVDD.n1582 DVDD.n1132 2.24398
R2447 DVDD.n1579 DVDD.n1190 2.24398
R2448 DVDD.n1133 DVDD.n1120 2.24398
R2449 DVDD.n1579 DVDD.n1188 2.24398
R2450 DVDD.n1135 DVDD.n1120 2.24398
R2451 DVDD.n1579 DVDD.n1187 2.24398
R2452 DVDD.n1137 DVDD.n1120 2.24398
R2453 DVDD.n1579 DVDD.n1186 2.24398
R2454 DVDD.n1139 DVDD.n1120 2.24398
R2455 DVDD.n1579 DVDD.n1185 2.24398
R2456 DVDD.n1141 DVDD.n1120 2.24398
R2457 DVDD.n1579 DVDD.n1184 2.24398
R2458 DVDD.n1143 DVDD.n1120 2.24398
R2459 DVDD.n1579 DVDD.n1183 2.24398
R2460 DVDD.n1145 DVDD.n1120 2.24398
R2461 DVDD.n1579 DVDD.n1182 2.24398
R2462 DVDD.n1147 DVDD.n1120 2.24398
R2463 DVDD.n1580 DVDD.n1579 2.24398
R2464 DVDD.n1149 DVDD.n1120 2.24398
R2465 DVDD.n1579 DVDD.n1119 2.24398
R2466 DVDD.n5420 DVDD.n5419 2.24383
R2467 DVDD.n105 DVDD.n104 2.24383
R2468 DVDD.n105 DVDD.n101 2.24383
R2469 DVDD.n350 DVDD.n348 2.24383
R2470 DVDD.n3777 DVDD.n1866 2.24304
R2471 DVDD.n3777 DVDD.n1865 2.24304
R2472 DVDD.n3777 DVDD.n1864 2.24304
R2473 DVDD.n3777 DVDD.n1863 2.24304
R2474 DVDD.n3777 DVDD.n1862 2.24304
R2475 DVDD.n3777 DVDD.n1860 2.24304
R2476 DVDD.n3777 DVDD.n1859 2.24304
R2477 DVDD.n3777 DVDD.n1858 2.24304
R2478 DVDD.n3777 DVDD.n1857 2.24304
R2479 DVDD.n2609 DVDD.n2608 2.24304
R2480 DVDD.n2618 DVDD.n2614 2.24304
R2481 DVDD.n2609 DVDD.n2607 2.24304
R2482 DVDD.n2618 DVDD.n2615 2.24304
R2483 DVDD.n2609 DVDD.n2606 2.24304
R2484 DVDD.n2618 DVDD.n2616 2.24304
R2485 DVDD.n2609 DVDD.n2605 2.24304
R2486 DVDD.n2618 DVDD.n2617 2.24304
R2487 DVDD.n2609 DVDD.n2603 2.24304
R2488 DVDD.n2598 DVDD.n2199 2.24304
R2489 DVDD.n2206 DVDD.n2198 2.24304
R2490 DVDD.n2598 DVDD.n2243 2.24304
R2491 DVDD.n2208 DVDD.n2198 2.24304
R2492 DVDD.n2598 DVDD.n2242 2.24304
R2493 DVDD.n2210 DVDD.n2198 2.24304
R2494 DVDD.n2598 DVDD.n2241 2.24304
R2495 DVDD.n2212 DVDD.n2198 2.24304
R2496 DVDD.n2599 DVDD.n2598 2.24304
R2497 DVDD.n3752 DVDD.n3720 2.24304
R2498 DVDD.n3752 DVDD.n3751 2.24304
R2499 DVDD.n3752 DVDD.n3750 2.24304
R2500 DVDD.n3752 DVDD.n3749 2.24304
R2501 DVDD.n3752 DVDD.n3748 2.24304
R2502 DVDD.n3752 DVDD.n3747 2.24304
R2503 DVDD.n3752 DVDD.n3746 2.24304
R2504 DVDD.n3752 DVDD.n3745 2.24304
R2505 DVDD.n3752 DVDD.n3744 2.24304
R2506 DVDD.n3752 DVDD.n3743 2.24304
R2507 DVDD.n4398 DVDD.n4388 2.24304
R2508 DVDD.n4411 DVDD.n4408 2.24304
R2509 DVDD.n4398 DVDD.n4389 2.24304
R2510 DVDD.n4411 DVDD.n4407 2.24304
R2511 DVDD.n4398 DVDD.n4390 2.24304
R2512 DVDD.n4411 DVDD.n4406 2.24304
R2513 DVDD.n4398 DVDD.n4391 2.24304
R2514 DVDD.n4411 DVDD.n4405 2.24304
R2515 DVDD.n4398 DVDD.n4392 2.24304
R2516 DVDD.n4411 DVDD.n4404 2.24304
R2517 DVDD.n4398 DVDD.n4393 2.24304
R2518 DVDD.n4411 DVDD.n4403 2.24304
R2519 DVDD.n4398 DVDD.n4394 2.24304
R2520 DVDD.n4411 DVDD.n4402 2.24304
R2521 DVDD.n4398 DVDD.n4395 2.24304
R2522 DVDD.n4411 DVDD.n4401 2.24304
R2523 DVDD.n4398 DVDD.n4396 2.24304
R2524 DVDD.n4411 DVDD.n4400 2.24304
R2525 DVDD.n4398 DVDD.n4397 2.24304
R2526 DVDD.n4412 DVDD.n4411 2.24304
R2527 DVDD.n4383 DVDD.n1594 2.24304
R2528 DVDD.n1608 DVDD.n1595 2.24304
R2529 DVDD.n4383 DVDD.n4374 2.24304
R2530 DVDD.n1610 DVDD.n1595 2.24304
R2531 DVDD.n4383 DVDD.n4375 2.24304
R2532 DVDD.n1612 DVDD.n1595 2.24304
R2533 DVDD.n4383 DVDD.n4376 2.24304
R2534 DVDD.n1614 DVDD.n1595 2.24304
R2535 DVDD.n4383 DVDD.n4377 2.24304
R2536 DVDD.n1616 DVDD.n1595 2.24304
R2537 DVDD.n4383 DVDD.n4378 2.24304
R2538 DVDD.n1618 DVDD.n1595 2.24304
R2539 DVDD.n4383 DVDD.n4379 2.24304
R2540 DVDD.n1620 DVDD.n1595 2.24304
R2541 DVDD.n4383 DVDD.n4380 2.24304
R2542 DVDD.n1622 DVDD.n1595 2.24304
R2543 DVDD.n4383 DVDD.n4381 2.24304
R2544 DVDD.n1624 DVDD.n1595 2.24304
R2545 DVDD.n4383 DVDD.n4382 2.24304
R2546 DVDD.n4384 DVDD.n1595 2.24304
R2547 DVDD.n4340 DVDD.n1626 2.24304
R2548 DVDD.n1640 DVDD.n1627 2.24304
R2549 DVDD.n4340 DVDD.n4331 2.24304
R2550 DVDD.n1642 DVDD.n1627 2.24304
R2551 DVDD.n4340 DVDD.n4332 2.24304
R2552 DVDD.n1644 DVDD.n1627 2.24304
R2553 DVDD.n4340 DVDD.n4333 2.24304
R2554 DVDD.n1646 DVDD.n1627 2.24304
R2555 DVDD.n4340 DVDD.n4334 2.24304
R2556 DVDD.n1648 DVDD.n1627 2.24304
R2557 DVDD.n4340 DVDD.n4335 2.24304
R2558 DVDD.n1650 DVDD.n1627 2.24304
R2559 DVDD.n4340 DVDD.n4336 2.24304
R2560 DVDD.n1652 DVDD.n1627 2.24304
R2561 DVDD.n4340 DVDD.n4337 2.24304
R2562 DVDD.n1654 DVDD.n1627 2.24304
R2563 DVDD.n4340 DVDD.n4338 2.24304
R2564 DVDD.n1656 DVDD.n1627 2.24304
R2565 DVDD.n4340 DVDD.n4339 2.24304
R2566 DVDD.n4341 DVDD.n1627 2.24304
R2567 DVDD.n3569 DVDD.n3143 2.24235
R2568 DVDD.n3185 DVDD.n3172 2.24235
R2569 DVDD.n1334 DVDD.n1331 2.24216
R2570 DVDD.n1338 DVDD.n1331 2.24216
R2571 DVDD.n1364 DVDD.n1330 2.24216
R2572 DVDD.n1364 DVDD.n1341 2.24216
R2573 DVDD.n1368 DVDD.n1333 2.24216
R2574 DVDD.n1366 DVDD.n1364 2.24216
R2575 DVDD.n1384 DVDD.n1380 2.23827
R2576 DVDD.n1325 DVDD.n1319 2.23827
R2577 DVDD.n1935 DVDD.n1915 2.20973
R2578 DVDD.n3316 DVDD.n3239 2.1705
R2579 DVDD.n3333 DVDD.n3332 2.1705
R2580 DVDD.n2735 DVDD.t83 2.09436
R2581 DVDD.n2736 DVDD.t152 2.09436
R2582 DVDD.n3380 DVDD.n3239 2.05485
R2583 DVDD.n3334 DVDD.n3333 1.98637
R2584 DVDD.n3382 DVDD.n3381 1.9605
R2585 DVDD.n3311 DVDD.n3310 1.9605
R2586 DVDD.n2715 DVDD.t29 1.95886
R2587 DVDD.n3065 DVDD.n2075 1.93369
R2588 DVDD.n3381 DVDD.n3380 1.92907
R2589 DVDD.n3334 DVDD.n3311 1.86479
R2590 DVDD.n3380 DVDD.n3240 1.8504
R2591 DVDD.n2794 DVDD.n2709 1.81438
R2592 DVDD.n2669 DVDD.t90 1.75468
R2593 DVDD.n2672 DVDD.n2671 1.74881
R2594 DVDD.n3334 DVDD.n3314 1.73846
R2595 DVDD.n2708 DVDD.n2706 1.71988
R2596 DVDD.n1375 DVDD.n1374 1.7146
R2597 DVDD.n3690 DVDD.n3689 1.71444
R2598 DVDD.n1374 DVDD.n1373 1.71412
R2599 DVDD.n2670 DVDD.n2669 1.70307
R2600 DVDD.n4237 DVDD.n1708 1.6972
R2601 DVDD.n4233 DVDD.n4232 1.6972
R2602 DVDD.n4203 DVDD.n4201 1.688
R2603 DVDD.n4136 DVDD.n1713 1.688
R2604 DVDD.n4126 DVDD.n4124 1.688
R2605 DVDD.n4123 DVDD.n1785 1.688
R2606 DVDD.n4122 DVDD.n4121 1.688
R2607 DVDD.n4013 DVDD.n4011 1.688
R2608 DVDD.n3994 DVDD.n3992 1.688
R2609 DVDD.n3930 DVDD.n3929 1.688
R2610 DVDD.n3964 DVDD.n3963 1.688
R2611 DVDD.n3962 DVDD.n3932 1.688
R2612 DVDD.n3961 DVDD.n3960 1.688
R2613 DVDD.n1875 DVDD.n1874 1.688
R2614 DVDD.n1878 DVDD.n1877 1.688
R2615 DVDD.n1869 DVDD.n1868 1.688
R2616 DVDD.n4231 DVDD.n1714 1.688
R2617 DVDD.n1958 DVDD.n1954 1.67609
R2618 DVDD.n1921 DVDD.n1916 1.67609
R2619 DVDD.n1882 DVDD.n1871 1.63826
R2620 DVDD.n1879 DVDD.n1872 1.63826
R2621 DVDD.n4230 DVDD.n1716 1.63826
R2622 DVDD.n4229 DVDD.n1717 1.63826
R2623 DVDD.n4174 DVDD.n1718 1.63826
R2624 DVDD.n4011 DVDD.n1711 1.63109
R2625 DVDD.n3992 DVDD.n1709 1.63109
R2626 DVDD.n3024 DVDD.n2075 1.62357
R2627 DVDD.n4201 DVDD.n4188 1.59264
R2628 DVDD.n2716 DVDD.n2715 1.58954
R2629 DVDD.n1883 DVDD.n1869 1.56519
R2630 DVDD.n2671 DVDD.t91 1.54008
R2631 DVDD.n3370 DVDD.n3269 1.52457
R2632 DVDD.n3628 DVDD.n3627 1.52019
R2633 DVDD.n2619 DVDD.n2602 1.5195
R2634 DVDD.n3515 DVDD.n3514 1.51933
R2635 DVDD.n3516 DVDD.n3161 1.51933
R2636 DVDD.n3776 DVDD.n3719 1.51565
R2637 DVDD.n2838 DVDD.n2089 1.50841
R2638 DVDD.n3663 DVDD.n1975 1.50806
R2639 DVDD.n2352 DVDD.t85 1.50625
R2640 DVDD.n2461 DVDD.t188 1.50625
R2641 DVDD.n2489 DVDD.t79 1.50625
R2642 DVDD.n2286 DVDD.t95 1.50625
R2643 DVDD.n2540 DVDD.t179 1.50625
R2644 DVDD.n2536 DVDD.t137 1.50625
R2645 DVDD.n2564 DVDD.t168 1.50625
R2646 DVDD.n3606 DVDD.n3605 1.50588
R2647 DVDD.n3415 DVDD.n3408 1.50588
R2648 DVDD.n3347 DVDD.n3099 1.50474
R2649 DVDD.n3398 DVDD.n3222 1.50474
R2650 DVDD.n2863 DVDD.n2693 1.50441
R2651 DVDD.n3719 DVDD.n3718 1.50165
R2652 DVDD.n3773 DVDD.n3772 1.50092
R2653 DVDD.n3555 DVDD.n3554 1.5005
R2654 DVDD.n3553 DVDD.n3552 1.5005
R2655 DVDD.n3140 DVDD.n3139 1.5005
R2656 DVDD.n3579 DVDD.n3578 1.5005
R2657 DVDD.n3581 DVDD.n3580 1.5005
R2658 DVDD.n3582 DVDD.n3137 1.5005
R2659 DVDD.n3136 DVDD.n3135 1.5005
R2660 DVDD.n3127 DVDD.n3125 1.5005
R2661 DVDD.n3591 DVDD.n3590 1.5005
R2662 DVDD.n3592 DVDD.n3122 1.5005
R2663 DVDD.n3594 DVDD.n3593 1.5005
R2664 DVDD.n3124 DVDD.n3121 1.5005
R2665 DVDD.n3472 DVDD.n3471 1.5005
R2666 DVDD.n3470 DVDD.n3193 1.5005
R2667 DVDD.n3469 DVDD.n3468 1.5005
R2668 DVDD.n3467 DVDD.n3466 1.5005
R2669 DVDD.n3196 DVDD.n3195 1.5005
R2670 DVDD.n3445 DVDD.n3444 1.5005
R2671 DVDD.n3443 DVDD.n3206 1.5005
R2672 DVDD.n3442 DVDD.n3441 1.5005
R2673 DVDD.n3436 DVDD.n3207 1.5005
R2674 DVDD.n3434 DVDD.n3433 1.5005
R2675 DVDD.n3432 DVDD.n3208 1.5005
R2676 DVDD.n3431 DVDD.n3430 1.5005
R2677 DVDD.n3476 DVDD.n3475 1.5005
R2678 DVDD.n3480 DVDD.n3479 1.5005
R2679 DVDD.n3482 DVDD.n3481 1.5005
R2680 DVDD.n3484 DVDD.n3483 1.5005
R2681 DVDD.n3486 DVDD.n3485 1.5005
R2682 DVDD.n3488 DVDD.n3487 1.5005
R2683 DVDD.n3490 DVDD.n3489 1.5005
R2684 DVDD.n3492 DVDD.n3491 1.5005
R2685 DVDD.n3494 DVDD.n3493 1.5005
R2686 DVDD.n3496 DVDD.n3495 1.5005
R2687 DVDD.n3498 DVDD.n3497 1.5005
R2688 DVDD.n3500 DVDD.n3499 1.5005
R2689 DVDD.n3502 DVDD.n3501 1.5005
R2690 DVDD.n3504 DVDD.n3503 1.5005
R2691 DVDD.n3506 DVDD.n3505 1.5005
R2692 DVDD.n3507 DVDD.n3192 1.5005
R2693 DVDD.n3511 DVDD.n3510 1.5005
R2694 DVDD.n3509 DVDD.n3508 1.5005
R2695 DVDD.n3170 DVDD.n3169 1.5005
R2696 DVDD.n3478 DVDD.n3477 1.5005
R2697 DVDD.n3518 DVDD.n3517 1.5005
R2698 DVDD.n3520 DVDD.n3519 1.5005
R2699 DVDD.n3522 DVDD.n3521 1.5005
R2700 DVDD.n3524 DVDD.n3523 1.5005
R2701 DVDD.n3526 DVDD.n3525 1.5005
R2702 DVDD.n3528 DVDD.n3527 1.5005
R2703 DVDD.n3530 DVDD.n3529 1.5005
R2704 DVDD.n3532 DVDD.n3531 1.5005
R2705 DVDD.n3534 DVDD.n3533 1.5005
R2706 DVDD.n3536 DVDD.n3535 1.5005
R2707 DVDD.n3538 DVDD.n3537 1.5005
R2708 DVDD.n3540 DVDD.n3539 1.5005
R2709 DVDD.n3542 DVDD.n3541 1.5005
R2710 DVDD.n3544 DVDD.n3543 1.5005
R2711 DVDD.n3546 DVDD.n3545 1.5005
R2712 DVDD.n3548 DVDD.n3547 1.5005
R2713 DVDD.n3550 DVDD.n3549 1.5005
R2714 DVDD.n3551 DVDD.n3168 1.5005
R2715 DVDD.n3559 DVDD.n3558 1.5005
R2716 DVDD.n3561 DVDD.n3560 1.5005
R2717 DVDD.n2837 DVDD.n2836 1.5005
R2718 DVDD.n2835 DVDD.n2834 1.5005
R2719 DVDD.n2833 DVDD.n2832 1.5005
R2720 DVDD.n2831 DVDD.n2830 1.5005
R2721 DVDD.n2829 DVDD.n2828 1.5005
R2722 DVDD.n2827 DVDD.n2826 1.5005
R2723 DVDD.n2825 DVDD.n2824 1.5005
R2724 DVDD.n2823 DVDD.n2822 1.5005
R2725 DVDD.n2821 DVDD.n2098 1.5005
R2726 DVDD.n2820 DVDD.n2096 1.5005
R2727 DVDD.n2819 DVDD.n2818 1.5005
R2728 DVDD.n2817 DVDD.n2696 1.5005
R2729 DVDD.n2816 DVDD.n2815 1.5005
R2730 DVDD.n2814 DVDD.n2697 1.5005
R2731 DVDD.n2813 DVDD.n2812 1.5005
R2732 DVDD.n2811 DVDD.n2698 1.5005
R2733 DVDD.n2810 DVDD.n2809 1.5005
R2734 DVDD.n2808 DVDD.n2699 1.5005
R2735 DVDD.n2807 DVDD.n2806 1.5005
R2736 DVDD.n2805 DVDD.n2700 1.5005
R2737 DVDD.n2846 DVDD.n2845 1.5005
R2738 DVDD.n2848 DVDD.n2847 1.5005
R2739 DVDD.n2850 DVDD.n2849 1.5005
R2740 DVDD.n2852 DVDD.n2851 1.5005
R2741 DVDD.n2854 DVDD.n2853 1.5005
R2742 DVDD.n2856 DVDD.n2855 1.5005
R2743 DVDD.n2858 DVDD.n2857 1.5005
R2744 DVDD.n2860 DVDD.n2859 1.5005
R2745 DVDD.n2862 DVDD.n2861 1.5005
R2746 DVDD.n1909 DVDD.n1903 1.5005
R2747 DVDD.n1912 DVDD.n1908 1.5005
R2748 DVDD.n3290 DVDD.n3288 1.5005
R2749 DVDD.n3291 DVDD.n3287 1.5005
R2750 DVDD.n3286 DVDD.n3285 1.5005
R2751 DVDD.n1910 DVDD.n1909 1.5005
R2752 DVDD.n1912 DVDD.n1911 1.5005
R2753 DVDD.n1913 DVDD.n1907 1.5005
R2754 DVDD.n3284 DVDD.n3270 1.5005
R2755 DVDD.n3285 DVDD.n3283 1.5005
R2756 DVDD.n3292 DVDD.n3291 1.5005
R2757 DVDD.n3290 DVDD.n3289 1.5005
R2758 DVDD.n3341 DVDD.n3097 1.5005
R2759 DVDD.n3368 DVDD.n3275 1.5005
R2760 DVDD.n3297 DVDD.n3296 1.5005
R2761 DVDD.n3361 DVDD.n3360 1.5005
R2762 DVDD.n3359 DVDD.n3358 1.5005
R2763 DVDD.n3298 DVDD.n3098 1.5005
R2764 DVDD.n3141 DVDD.n3138 1.5005
R2765 DVDD.n3583 DVDD.n3582 1.5005
R2766 DVDD.n3589 DVDD.n3588 1.5005
R2767 DVDD.n3126 DVDD.n1993 1.5005
R2768 DVDD.n3120 DVDD.n3114 1.5005
R2769 DVDD.n3602 DVDD.n3601 1.5005
R2770 DVDD.n3596 DVDD.n3595 1.5005
R2771 DVDD.n3134 DVDD.n3128 1.5005
R2772 DVDD.n3577 DVDD.n3576 1.5005
R2773 DVDD.n3373 DVDD.n3372 1.5005
R2774 DVDD.n3267 DVDD.n3246 1.5005
R2775 DVDD.n3261 DVDD.n3260 1.5005
R2776 DVDD.n3389 DVDD.n3232 1.5005
R2777 DVDD.n3231 DVDD.n3096 1.5005
R2778 DVDD.n3409 DVDD.n3210 1.5005
R2779 DVDD.n3429 DVDD.n3428 1.5005
R2780 DVDD.n3435 DVDD.n1991 1.5005
R2781 DVDD.n3439 DVDD.n3438 1.5005
R2782 DVDD.n3440 DVDD.n3205 1.5005
R2783 DVDD.n3446 DVDD.n3445 1.5005
R2784 DVDD.n3465 DVDD.n3464 1.5005
R2785 DVDD.n3198 DVDD.n3194 1.5005
R2786 DVDD.n3419 DVDD.n3418 1.5005
R2787 DVDD.n3639 DVDD.n3638 1.5005
R2788 DVDD.n3627 DVDD.n2016 1.5005
R2789 DVDD.n3640 DVDD.n2007 1.5005
R2790 DVDD.n3642 DVDD.n3641 1.5005
R2791 DVDD.n2008 DVDD.n1981 1.5005
R2792 DVDD.n3655 DVDD.n3654 1.5005
R2793 DVDD.n3656 DVDD.n1979 1.5005
R2794 DVDD.n3667 DVDD.n3666 1.5005
R2795 DVDD.n3665 DVDD.n3664 1.5005
R2796 DVDD.n4299 DVDD.n4298 1.5005
R2797 DVDD.n4293 DVDD.n1658 1.5005
R2798 DVDD.n4292 DVDD.n4291 1.5005
R2799 DVDD.n4290 DVDD.n4289 1.5005
R2800 DVDD.n1665 DVDD.n1664 1.5005
R2801 DVDD.n3765 DVDD.n3764 1.5005
R2802 DVDD.n3767 DVDD.n3766 1.5005
R2803 DVDD.n3761 DVDD.n3759 1.5005
R2804 DVDD.n3754 DVDD.n3753 1.5005
R2805 DVDD.n1889 DVDD.n1888 1.5005
R2806 DVDD.n3713 DVDD.n3712 1.5005
R2807 DVDD.n3711 DVDD.n1893 1.5005
R2808 DVDD.n3710 DVDD.n3709 1.5005
R2809 DVDD.n2180 DVDD.n1895 1.5005
R2810 DVDD.n2184 DVDD.n2183 1.5005
R2811 DVDD.n2186 DVDD.n2185 1.5005
R2812 DVDD.n2175 DVDD.n2173 1.5005
R2813 DVDD.n2192 DVDD.n2191 1.5005
R2814 DVDD.n960 DVDD.n942 1.5005
R2815 DVDD.n928 DVDD.n927 1.5005
R2816 DVDD.n940 DVDD.n939 1.5005
R2817 DVDD.n938 DVDD.n937 1.5005
R2818 DVDD.n936 DVDD.n935 1.5005
R2819 DVDD.n934 DVDD.n933 1.5005
R2820 DVDD.n932 DVDD.n931 1.5005
R2821 DVDD.n930 DVDD.n929 1.5005
R2822 DVDD.n951 DVDD.n950 1.5005
R2823 DVDD.n953 DVDD.n952 1.5005
R2824 DVDD.n955 DVDD.n954 1.5005
R2825 DVDD.n957 DVDD.n956 1.5005
R2826 DVDD.n959 DVDD.n958 1.5005
R2827 DVDD.n245 DVDD.n244 1.5005
R2828 DVDD.n258 DVDD.n257 1.5005
R2829 DVDD.n247 DVDD.n246 1.5005
R2830 DVDD.n249 DVDD.n248 1.5005
R2831 DVDD.n251 DVDD.n250 1.5005
R2832 DVDD.n253 DVDD.n252 1.5005
R2833 DVDD.n255 DVDD.n254 1.5005
R2834 DVDD.n5665 DVDD.n5664 1.5005
R2835 DVDD.n5667 DVDD.n5666 1.5005
R2836 DVDD.n5669 DVDD.n5668 1.5005
R2837 DVDD.n5670 DVDD.n242 1.5005
R2838 DVDD.n5672 DVDD.n5671 1.5005
R2839 DVDD.n243 DVDD.n240 1.5005
R2840 DVDD.n2465 DVDD.t62 1.49967
R2841 DVDD.n2466 DVDD.n2465 1.45483
R2842 DVDD.n2276 DVDD.n2275 1.4515
R2843 DVDD.n2535 DVDD.n2295 1.4515
R2844 DVDD.n2342 DVDD.n2341 1.4515
R2845 DVDD.n2460 DVDD.n2361 1.4515
R2846 DVDD.n2565 DVDD.n2564 1.45148
R2847 DVDD.n2287 DVDD.n2286 1.45148
R2848 DVDD.n2536 DVDD.n2264 1.45148
R2849 DVDD.n2541 DVDD.n2540 1.45148
R2850 DVDD.n2490 DVDD.n2489 1.45148
R2851 DVDD.n2353 DVDD.n2352 1.45148
R2852 DVDD.n2461 DVDD.n2328 1.45148
R2853 DVDD.n2600 DVDD 1.39172
R2854 DVDD.n2239 DVDD.n2238 1.33383
R2855 DVDD.n5499 DVDD.n261 1.33314
R2856 DVDD.n2793 DVDD.n2713 1.33037
R2857 DVDD.n4238 DVDD.n4237 1.3141
R2858 DVDD.n4233 DVDD.n1712 1.3141
R2859 DVDD.n2840 DVDD.n2838 1.31276
R2860 DVDD.n1953 DVDD.n1952 1.31159
R2861 DVDD.n2484 DVDD.n2483 1.2972
R2862 DVDD.n2457 DVDD.n2456 1.2972
R2863 DVDD.n2487 DVDD.n2323 1.2972
R2864 DVDD.n2559 DVDD.n2558 1.2972
R2865 DVDD.n2532 DVDD.n2531 1.2972
R2866 DVDD.n2562 DVDD.n2255 1.2972
R2867 DVDD.n3414 DVDD.n3111 1.29474
R2868 DVDD.n1957 DVDD.n1956 1.28124
R2869 DVDD.n1923 DVDD.n1922 1.28123
R2870 DVDD.n1920 DVDD.n1919 1.28123
R2871 DVDD.n4157 DVDD.n1716 1.26907
R2872 DVDD.n1877 DVDD.n1695 1.26907
R2873 DVDD.n3952 DVDD.n3932 1.26907
R2874 DVDD.n3965 DVDD.n3964 1.26907
R2875 DVDD.n3929 DVDD.n3923 1.26907
R2876 DVDD.n4121 DVDD.n4119 1.26907
R2877 DVDD.n4113 DVDD.n1785 1.26907
R2878 DVDD.n4127 DVDD.n4126 1.26907
R2879 DVDD.n1392 DVDD.n1391 1.18293
R2880 DVDD.n1315 DVDD.n1222 1.18293
R2881 DVDD.n5731 DVDD.n5730 1.17409
R2882 DVDD.n5091 DVDD.n5087 1.17409
R2883 DVDD.n598 DVDD.n596 1.17409
R2884 DVDD.n878 DVDD.n877 1.17409
R2885 DVDD.n1060 DVDD.n896 1.17409
R2886 DVDD.n5847 DVDD.n5846 1.17318
R2887 DVDD.n5136 DVDD.n5103 1.17318
R2888 DVDD.n4993 DVDD.n428 1.17318
R2889 DVDD.n759 DVDD.n404 1.17318
R2890 DVDD.n4549 DVDD.n381 1.17318
R2891 DVDD.n2193 DVDD.n2192 1.15295
R2892 DVDD.n2485 DVDD.n2484 1.14595
R2893 DVDD.n2560 DVDD.n2559 1.14595
R2894 DVDD.n3696 DVDD.n3695 1.1282
R2895 DVDD.n2236 DVDD.n2235 1.1255
R2896 DVDD.n2238 DVDD.n2237 1.1255
R2897 DVDD.n2232 DVDD.n2231 1.1255
R2898 DVDD.n2234 DVDD.n2233 1.1255
R2899 DVDD.n2228 DVDD.n2227 1.1255
R2900 DVDD.n2230 DVDD.n2229 1.1255
R2901 DVDD.n2224 DVDD.n2223 1.1255
R2902 DVDD.n2226 DVDD.n2225 1.1255
R2903 DVDD.n2220 DVDD.n2219 1.1255
R2904 DVDD.n2222 DVDD.n2221 1.1255
R2905 DVDD.n2216 DVDD.n2215 1.1255
R2906 DVDD.n2218 DVDD.n2217 1.1255
R2907 DVDD.n2796 DVDD.n2795 1.1255
R2908 DVDD.n1957 DVDD.n1955 1.11867
R2909 DVDD.n1952 DVDD.n1951 1.11867
R2910 DVDD.n1923 DVDD.n1917 1.11867
R2911 DVDD.n1919 DVDD.n1918 1.11867
R2912 DVDD.n3023 DVDD.n3022 1.08635
R2913 DVDD.n2463 DVDD.n2458 1.0505
R2914 DVDD.n2486 DVDD.n2325 1.0505
R2915 DVDD.n2538 DVDD.n2533 1.0505
R2916 DVDD.n2561 DVDD.n2261 1.0505
R2917 DVDD.n3694 DVDD.n3693 0.969731
R2918 DVDD.n1578 DVDD.n1577 0.969652
R2919 DVDD.n2799 DVDD.n2798 0.968342
R2920 DVDD.n2709 DVDD.t12 0.958395
R2921 DVDD.n2709 DVDD.t10 0.958395
R2922 DVDD.n2710 DVDD.t73 0.9105
R2923 DVDD.n2710 DVDD.t75 0.9105
R2924 DVDD.n2191 DVDD.n2174 0.909532
R2925 DVDD.n4298 DVDD.n4297 0.908802
R2926 DVDD.n3718 DVDD.n3717 0.908384
R2927 DVDD.n3772 DVDD.n3771 0.908384
R2928 DVDD.n4137 DVDD.n4136 0.904312
R2929 DVDD.n3960 DVDD.n3959 0.904312
R2930 DVDD.n1874 DVDD.n1873 0.904312
R2931 DVDD.n4147 DVDD.n1714 0.904312
R2932 DVDD.n3384 DVDD.n3383 0.9005
R2933 DVDD.n3331 DVDD.n3330 0.9005
R2934 DVDD.n3338 DVDD.n3337 0.9005
R2935 DVDD.n3318 DVDD.n3317 0.9005
R2936 DVDD.n2188 DVDD.n2176 0.9005
R2937 DVDD.n2178 DVDD.n2177 0.9005
R2938 DVDD.n2181 DVDD.n1968 0.9005
R2939 DVDD.n3706 DVDD.n3705 0.9005
R2940 DVDD.n1892 DVDD.n1891 0.9005
R2941 DVDD.n3716 DVDD.n3715 0.9005
R2942 DVDD.n2190 DVDD.n2189 0.9005
R2943 DVDD.n2188 DVDD.n2187 0.9005
R2944 DVDD.n2179 DVDD.n2178 0.9005
R2945 DVDD.n2182 DVDD.n2181 0.9005
R2946 DVDD.n3707 DVDD.n3706 0.9005
R2947 DVDD.n3708 DVDD.n1892 0.9005
R2948 DVDD.n3715 DVDD.n3714 0.9005
R2949 DVDD.n1894 DVDD.n1890 0.9005
R2950 DVDD.n3770 DVDD.n3769 0.9005
R2951 DVDD.n3757 DVDD.n3756 0.9005
R2952 DVDD.n3762 DVDD.n1667 0.9005
R2953 DVDD.n4287 DVDD.n4286 0.9005
R2954 DVDD.n1662 DVDD.n1661 0.9005
R2955 DVDD.n4296 DVDD.n4295 0.9005
R2956 DVDD.n3758 DVDD.n3755 0.9005
R2957 DVDD.n3769 DVDD.n3768 0.9005
R2958 DVDD.n3760 DVDD.n3757 0.9005
R2959 DVDD.n3763 DVDD.n3762 0.9005
R2960 DVDD.n4288 DVDD.n4287 0.9005
R2961 DVDD.n1663 DVDD.n1662 0.9005
R2962 DVDD.n4295 DVDD.n4294 0.9005
R2963 DVDD.n1660 DVDD.n1659 0.9005
R2964 DVDD.n2460 DVDD.n2459 0.899883
R2965 DVDD.n2341 DVDD.n2340 0.899883
R2966 DVDD.n2535 DVDD.n2534 0.899883
R2967 DVDD.n2275 DVDD.n2274 0.899883
R2968 DVDD.n1375 DVDD.n1370 0.886656
R2969 DVDD.n2795 DVDD.n2708 0.875562
R2970 DVDD.n1373 DVDD.n1371 0.87516
R2971 DVDD.n2735 DVDD.n2734 0.8555
R2972 DVDD.n5662 DVDD.n259 0.82049
R2973 DVDD.n5488 DVDD.n263 0.814302
R2974 DVDD.n1915 DVDD.n1914 0.791147
R2975 DVDD.n1868 DVDD.n1852 0.773058
R2976 DVDD.n1871 DVDD.n1690 0.773058
R2977 DVDD.n1872 DVDD.n1691 0.773058
R2978 DVDD.n3995 DVDD.n3994 0.773058
R2979 DVDD.n4014 DVDD.n4013 0.773058
R2980 DVDD.n1769 DVDD.n1717 0.773058
R2981 DVDD.n4175 DVDD.n4174 0.773058
R2982 DVDD.n4204 DVDD.n4203 0.773058
R2983 DVDD.n2215 DVDD.n2214 0.771833
R2984 DVDD.n1960 DVDD.n1959 0.769687
R2985 DVDD.n3286 DVDD.n3269 0.769684
R2986 DVDD.n3064 DVDD.n3063 0.755277
R2987 DVDD.n3474 DVDD.n3473 0.751
R2988 DVDD.n3557 DVDD.n3556 0.751
R2989 DVDD.n3651 DVDD.n3650 0.7505
R2990 DVDD.n3650 DVDD.n3649 0.7505
R2991 DVDD.n3329 DVDD.n3328 0.735937
R2992 DVDD.n3322 DVDD.n3271 0.735937
R2993 DVDD.n3374 DVDD.n3245 0.735937
R2994 DVDD.n3320 DVDD.n3249 0.735937
R2995 DVDD.n2706 DVDD.n2693 0.734685
R2996 DVDD.n2464 DVDD.n2457 0.714509
R2997 DVDD.n2488 DVDD.n2487 0.714509
R2998 DVDD.n2539 DVDD.n2532 0.714509
R2999 DVDD.n2563 DVDD.n2562 0.714509
R3000 DVDD.n2777 DVDD.n2737 0.711129
R3001 DVDD.n2775 DVDD.n2759 0.711129
R3002 DVDD.n2770 DVDD.n2769 0.7005
R3003 DVDD.n2771 DVDD.n2752 0.7005
R3004 DVDD.n2772 DVDD.n2755 0.7005
R3005 DVDD.n2773 DVDD.n2751 0.7005
R3006 DVDD.n2775 DVDD.n2774 0.7005
R3007 DVDD.n2759 DVDD.n2742 0.7005
R3008 DVDD.n2778 DVDD.n2777 0.7005
R3009 DVDD.n2779 DVDD.n2737 0.7005
R3010 DVDD.n2784 DVDD.n2783 0.7005
R3011 DVDD.n2786 DVDD.n2785 0.7005
R3012 DVDD.n2733 DVDD.n2719 0.7005
R3013 DVDD.n2789 DVDD.n2788 0.7005
R3014 DVDD.n2718 DVDD.n2717 0.668882
R3015 DVDD.n2713 DVDD.n2711 0.666798
R3016 DVDD.n3692 DVDD.n3690 0.646382
R3017 DVDD.n2718 DVDD.n2708 0.645825
R3018 DVDD.n4200 DVDD.n4198 0.634998
R3019 DVDD.n1935 DVDD.n1934 0.634532
R3020 DVDD.n1379 DVDD.n1325 0.634344
R3021 DVDD.n1380 DVDD.n1379 0.632309
R3022 DVDD.n2459 DVDD.t190 0.607167
R3023 DVDD.n2459 DVDD.t196 0.607167
R3024 DVDD.n2340 DVDD.t77 0.607167
R3025 DVDD.n2340 DVDD.t119 0.607167
R3026 DVDD.n2534 DVDD.t135 0.607167
R3027 DVDD.n2534 DVDD.t181 0.607167
R3028 DVDD.n2274 DVDD.t89 0.607167
R3029 DVDD.n2274 DVDD.t93 0.607167
R3030 DVDD.n3689 DVDD.t39 0.607167
R3031 DVDD.n3689 DVDD.t121 0.607167
R3032 DVDD.n2797 DVDD.n2796 0.594875
R3033 DVDD.n4231 DVDD.n4230 0.590794
R3034 DVDD.n4230 DVDD.n4229 0.578395
R3035 DVDD.n2726 DVDD.n2714 0.573227
R3036 DVDD.n2790 DVDD.n2714 0.573227
R3037 DVDD.n2736 DVDD 0.565368
R3038 DVDD.n3394 DVDD.n3222 0.563
R3039 DVDD.n3346 DVDD.n3345 0.563
R3040 DVDD.n3348 DVDD.n3347 0.563
R3041 DVDD.n3393 DVDD.n3392 0.563
R3042 DVDD.n3064 DVDD.n3027 0.563
R3043 DVDD.n2484 DVDD.n2326 0.557079
R3044 DVDD.n2559 DVDD.n2262 0.557079
R3045 DVDD.n1879 DVDD.n1878 0.552481
R3046 DVDD.n2464 DVDD.n2463 0.545794
R3047 DVDD.n2488 DVDD.n2325 0.545794
R3048 DVDD.n2539 DVDD.n2538 0.545794
R3049 DVDD.n2563 DVDD.n2261 0.545794
R3050 DVDD.n4124 DVDD.n1713 0.545794
R3051 DVDD.n4124 DVDD.n4123 0.545794
R3052 DVDD.n3963 DVDD.n3962 0.545794
R3053 DVDD.n3962 DVDD.n3961 0.545794
R3054 DVDD.n1878 DVDD.n1875 0.545794
R3055 DVDD.n3330 DVDD.n3329 0.527932
R3056 DVDD.n3317 DVDD.n3245 0.527932
R3057 DVDD.n1914 DVDD.n1908 0.525612
R3058 DVDD.n3695 DVDD 0.471676
R3059 DVDD.n2465 DVDD.n2464 0.463605
R3060 DVDD.n2598 DVDD.n2240 0.463585
R3061 DVDD.n2618 DVDD.n2604 0.463585
R3062 DVDD.n2176 DVDD.n2174 0.459655
R3063 DVDD.n3717 DVDD.n3716 0.459655
R3064 DVDD.n3771 DVDD.n3770 0.459655
R3065 DVDD.n4297 DVDD.n4296 0.459655
R3066 DVDD.n2352 DVDD.n2351 0.457026
R3067 DVDD.n2462 DVDD.n2461 0.457026
R3068 DVDD.n2489 DVDD.n2488 0.457026
R3069 DVDD.n2286 DVDD.n2285 0.457026
R3070 DVDD.n2540 DVDD.n2539 0.457026
R3071 DVDD.n2537 DVDD.n2536 0.457026
R3072 DVDD.n2564 DVDD.n2563 0.457026
R3073 DVDD.n2463 DVDD.n2460 0.457011
R3074 DVDD.n2341 DVDD.n2325 0.457011
R3075 DVDD.n2538 DVDD.n2535 0.457011
R3076 DVDD.n2275 DVDD.n2261 0.457011
R3077 DVDD.n1958 DVDD 0.455237
R3078 DVDD DVDD.n1916 0.455237
R3079 DVDD.n2595 DVDD.n2594 0.4505
R3080 DVDD.n2593 DVDD.n2244 0.4505
R3081 DVDD.n2592 DVDD.n2591 0.4505
R3082 DVDD.n2246 DVDD.n2245 0.4505
R3083 DVDD.n2587 DVDD.n2586 0.4505
R3084 DVDD.n2585 DVDD.n2248 0.4505
R3085 DVDD.n2584 DVDD.n2583 0.4505
R3086 DVDD.n2250 DVDD.n2249 0.4505
R3087 DVDD.n2579 DVDD.n2578 0.4505
R3088 DVDD.n2577 DVDD.n2252 0.4505
R3089 DVDD.n2576 DVDD.n2575 0.4505
R3090 DVDD.n2254 DVDD.n2253 0.4505
R3091 DVDD.n2571 DVDD.n2570 0.4505
R3092 DVDD.n2569 DVDD.n2256 0.4505
R3093 DVDD.n2568 DVDD.n2567 0.4505
R3094 DVDD.n2258 DVDD.n2257 0.4505
R3095 DVDD.n2272 DVDD.n2271 0.4505
R3096 DVDD.n2279 DVDD.n2278 0.4505
R3097 DVDD.n2280 DVDD.n2270 0.4505
R3098 DVDD.n2282 DVDD.n2281 0.4505
R3099 DVDD.n2268 DVDD.n2267 0.4505
R3100 DVDD.n2290 DVDD.n2289 0.4505
R3101 DVDD.n2291 DVDD.n2265 0.4505
R3102 DVDD.n2556 DVDD.n2555 0.4505
R3103 DVDD.n2554 DVDD.n2266 0.4505
R3104 DVDD.n2553 DVDD.n2552 0.4505
R3105 DVDD.n2293 DVDD.n2292 0.4505
R3106 DVDD.n2548 DVDD.n2547 0.4505
R3107 DVDD.n2546 DVDD.n2296 0.4505
R3108 DVDD.n2545 DVDD.n2544 0.4505
R3109 DVDD.n2298 DVDD.n2297 0.4505
R3110 DVDD.n2304 DVDD.n2302 0.4505
R3111 DVDD.n2529 DVDD.n2528 0.4505
R3112 DVDD.n2527 DVDD.n2303 0.4505
R3113 DVDD.n2526 DVDD.n2525 0.4505
R3114 DVDD.n2306 DVDD.n2305 0.4505
R3115 DVDD.n2521 DVDD.n2520 0.4505
R3116 DVDD.n2519 DVDD.n2308 0.4505
R3117 DVDD.n2518 DVDD.n2517 0.4505
R3118 DVDD.n2310 DVDD.n2309 0.4505
R3119 DVDD.n2513 DVDD.n2512 0.4505
R3120 DVDD.n2511 DVDD.n2312 0.4505
R3121 DVDD.n2510 DVDD.n2509 0.4505
R3122 DVDD.n2314 DVDD.n2313 0.4505
R3123 DVDD.n2505 DVDD.n2504 0.4505
R3124 DVDD.n2503 DVDD.n2316 0.4505
R3125 DVDD.n2502 DVDD.n2501 0.4505
R3126 DVDD.n2318 DVDD.n2317 0.4505
R3127 DVDD.n2497 DVDD.n2496 0.4505
R3128 DVDD.n2495 DVDD.n2320 0.4505
R3129 DVDD.n2494 DVDD.n2493 0.4505
R3130 DVDD.n2322 DVDD.n2321 0.4505
R3131 DVDD.n2337 DVDD.n2336 0.4505
R3132 DVDD.n2338 DVDD.n2335 0.4505
R3133 DVDD.n2345 DVDD.n2344 0.4505
R3134 DVDD.n2346 DVDD.n2334 0.4505
R3135 DVDD.n2348 DVDD.n2347 0.4505
R3136 DVDD.n2332 DVDD.n2331 0.4505
R3137 DVDD.n2356 DVDD.n2355 0.4505
R3138 DVDD.n2357 DVDD.n2329 0.4505
R3139 DVDD.n2481 DVDD.n2480 0.4505
R3140 DVDD.n2479 DVDD.n2330 0.4505
R3141 DVDD.n2478 DVDD.n2477 0.4505
R3142 DVDD.n2359 DVDD.n2358 0.4505
R3143 DVDD.n2473 DVDD.n2472 0.4505
R3144 DVDD.n2471 DVDD.n2362 0.4505
R3145 DVDD.n2470 DVDD.n2469 0.4505
R3146 DVDD.n2364 DVDD.n2363 0.4505
R3147 DVDD.n2370 DVDD.n2368 0.4505
R3148 DVDD.n2454 DVDD.n2453 0.4505
R3149 DVDD.n2452 DVDD.n2369 0.4505
R3150 DVDD.n2451 DVDD.n2450 0.4505
R3151 DVDD.n2372 DVDD.n2371 0.4505
R3152 DVDD.n2446 DVDD.n2445 0.4505
R3153 DVDD.n2444 DVDD.n2374 0.4505
R3154 DVDD.n2443 DVDD.n2442 0.4505
R3155 DVDD.n2376 DVDD.n2375 0.4505
R3156 DVDD.n2438 DVDD.n2437 0.4505
R3157 DVDD.n2436 DVDD.n2378 0.4505
R3158 DVDD.n2435 DVDD.n2434 0.4505
R3159 DVDD.n2380 DVDD.n2379 0.4505
R3160 DVDD.n2430 DVDD.n2429 0.4505
R3161 DVDD.n2428 DVDD.n2382 0.4505
R3162 DVDD.n2427 DVDD.n2426 0.4505
R3163 DVDD.n2384 DVDD.n2383 0.4505
R3164 DVDD.n2422 DVDD.n2421 0.4505
R3165 DVDD.n2420 DVDD.n2386 0.4505
R3166 DVDD.n2419 DVDD.n2418 0.4505
R3167 DVDD.n2388 DVDD.n2387 0.4505
R3168 DVDD.n2414 DVDD.n2413 0.4505
R3169 DVDD.n2412 DVDD.n2390 0.4505
R3170 DVDD.n2411 DVDD.n2410 0.4505
R3171 DVDD.n2392 DVDD.n2391 0.4505
R3172 DVDD.n2406 DVDD.n2405 0.4505
R3173 DVDD.n2404 DVDD.n2394 0.4505
R3174 DVDD.n2403 DVDD.n2402 0.4505
R3175 DVDD.n2396 DVDD.n2395 0.4505
R3176 DVDD.n2398 DVDD.n2397 0.4505
R3177 DVDD.n2400 DVDD.n2396 0.4505
R3178 DVDD.n2402 DVDD.n2401 0.4505
R3179 DVDD.n2394 DVDD.n2393 0.4505
R3180 DVDD.n2407 DVDD.n2406 0.4505
R3181 DVDD.n2408 DVDD.n2392 0.4505
R3182 DVDD.n2410 DVDD.n2409 0.4505
R3183 DVDD.n2390 DVDD.n2389 0.4505
R3184 DVDD.n2415 DVDD.n2414 0.4505
R3185 DVDD.n2416 DVDD.n2388 0.4505
R3186 DVDD.n2418 DVDD.n2417 0.4505
R3187 DVDD.n2386 DVDD.n2385 0.4505
R3188 DVDD.n2423 DVDD.n2422 0.4505
R3189 DVDD.n2424 DVDD.n2384 0.4505
R3190 DVDD.n2426 DVDD.n2425 0.4505
R3191 DVDD.n2382 DVDD.n2381 0.4505
R3192 DVDD.n2431 DVDD.n2430 0.4505
R3193 DVDD.n2432 DVDD.n2380 0.4505
R3194 DVDD.n2434 DVDD.n2433 0.4505
R3195 DVDD.n2378 DVDD.n2377 0.4505
R3196 DVDD.n2439 DVDD.n2438 0.4505
R3197 DVDD.n2440 DVDD.n2376 0.4505
R3198 DVDD.n2442 DVDD.n2441 0.4505
R3199 DVDD.n2374 DVDD.n2373 0.4505
R3200 DVDD.n2447 DVDD.n2446 0.4505
R3201 DVDD.n2448 DVDD.n2372 0.4505
R3202 DVDD.n2450 DVDD.n2449 0.4505
R3203 DVDD.n2369 DVDD.n2367 0.4505
R3204 DVDD.n2455 DVDD.n2454 0.4505
R3205 DVDD.n2368 DVDD.n2366 0.4505
R3206 DVDD.n2467 DVDD.n2364 0.4505
R3207 DVDD.n2469 DVDD.n2468 0.4505
R3208 DVDD.n2365 DVDD.n2362 0.4505
R3209 DVDD.n2474 DVDD.n2473 0.4505
R3210 DVDD.n2475 DVDD.n2359 0.4505
R3211 DVDD.n2477 DVDD.n2476 0.4505
R3212 DVDD.n2360 DVDD.n2330 0.4505
R3213 DVDD.n2482 DVDD.n2481 0.4505
R3214 DVDD.n2329 DVDD.n2327 0.4505
R3215 DVDD.n2355 DVDD.n2354 0.4505
R3216 DVDD.n2350 DVDD.n2332 0.4505
R3217 DVDD.n2349 DVDD.n2348 0.4505
R3218 DVDD.n2334 DVDD.n2333 0.4505
R3219 DVDD.n2344 DVDD.n2343 0.4505
R3220 DVDD.n2339 DVDD.n2338 0.4505
R3221 DVDD.n2337 DVDD.n2324 0.4505
R3222 DVDD.n2491 DVDD.n2322 0.4505
R3223 DVDD.n2493 DVDD.n2492 0.4505
R3224 DVDD.n2320 DVDD.n2319 0.4505
R3225 DVDD.n2498 DVDD.n2497 0.4505
R3226 DVDD.n2499 DVDD.n2318 0.4505
R3227 DVDD.n2501 DVDD.n2500 0.4505
R3228 DVDD.n2316 DVDD.n2315 0.4505
R3229 DVDD.n2506 DVDD.n2505 0.4505
R3230 DVDD.n2507 DVDD.n2314 0.4505
R3231 DVDD.n2509 DVDD.n2508 0.4505
R3232 DVDD.n2312 DVDD.n2311 0.4505
R3233 DVDD.n2514 DVDD.n2513 0.4505
R3234 DVDD.n2515 DVDD.n2310 0.4505
R3235 DVDD.n2517 DVDD.n2516 0.4505
R3236 DVDD.n2308 DVDD.n2307 0.4505
R3237 DVDD.n2522 DVDD.n2521 0.4505
R3238 DVDD.n2523 DVDD.n2306 0.4505
R3239 DVDD.n2525 DVDD.n2524 0.4505
R3240 DVDD.n2303 DVDD.n2301 0.4505
R3241 DVDD.n2530 DVDD.n2529 0.4505
R3242 DVDD.n2302 DVDD.n2300 0.4505
R3243 DVDD.n2542 DVDD.n2298 0.4505
R3244 DVDD.n2544 DVDD.n2543 0.4505
R3245 DVDD.n2299 DVDD.n2296 0.4505
R3246 DVDD.n2549 DVDD.n2548 0.4505
R3247 DVDD.n2550 DVDD.n2293 0.4505
R3248 DVDD.n2552 DVDD.n2551 0.4505
R3249 DVDD.n2294 DVDD.n2266 0.4505
R3250 DVDD.n2557 DVDD.n2556 0.4505
R3251 DVDD.n2265 DVDD.n2263 0.4505
R3252 DVDD.n2289 DVDD.n2288 0.4505
R3253 DVDD.n2284 DVDD.n2268 0.4505
R3254 DVDD.n2283 DVDD.n2282 0.4505
R3255 DVDD.n2270 DVDD.n2269 0.4505
R3256 DVDD.n2278 DVDD.n2277 0.4505
R3257 DVDD.n2273 DVDD.n2272 0.4505
R3258 DVDD.n2260 DVDD.n2258 0.4505
R3259 DVDD.n2567 DVDD.n2566 0.4505
R3260 DVDD.n2259 DVDD.n2256 0.4505
R3261 DVDD.n2572 DVDD.n2571 0.4505
R3262 DVDD.n2573 DVDD.n2254 0.4505
R3263 DVDD.n2575 DVDD.n2574 0.4505
R3264 DVDD.n2252 DVDD.n2251 0.4505
R3265 DVDD.n2580 DVDD.n2579 0.4505
R3266 DVDD.n2581 DVDD.n2250 0.4505
R3267 DVDD.n2583 DVDD.n2582 0.4505
R3268 DVDD.n2248 DVDD.n2247 0.4505
R3269 DVDD.n2588 DVDD.n2587 0.4505
R3270 DVDD.n2589 DVDD.n2246 0.4505
R3271 DVDD.n2591 DVDD.n2590 0.4505
R3272 DVDD.n2244 DVDD.n2205 0.4505
R3273 DVDD.n2595 DVDD.n2200 0.4505
R3274 DVDD.n2597 DVDD.n2596 0.4505
R3275 DVDD.n2611 DVDD.n2610 0.4505
R3276 DVDD.n2167 DVDD.n2166 0.4505
R3277 DVDD.n2624 DVDD.n2623 0.4505
R3278 DVDD.n2625 DVDD.n2165 0.4505
R3279 DVDD.n2627 DVDD.n2626 0.4505
R3280 DVDD.n2163 DVDD.n2162 0.4505
R3281 DVDD.n2632 DVDD.n2631 0.4505
R3282 DVDD.n2633 DVDD.n2161 0.4505
R3283 DVDD.n2635 DVDD.n2634 0.4505
R3284 DVDD.n2159 DVDD.n2158 0.4505
R3285 DVDD.n2640 DVDD.n2639 0.4505
R3286 DVDD.n2641 DVDD.n2157 0.4505
R3287 DVDD.n2643 DVDD.n2642 0.4505
R3288 DVDD.n2155 DVDD.n2154 0.4505
R3289 DVDD.n2648 DVDD.n2647 0.4505
R3290 DVDD.n2649 DVDD.n2153 0.4505
R3291 DVDD.n2651 DVDD.n2650 0.4505
R3292 DVDD.n2151 DVDD.n2150 0.4505
R3293 DVDD.n2656 DVDD.n2655 0.4505
R3294 DVDD.n2657 DVDD.n2149 0.4505
R3295 DVDD.n2659 DVDD.n2658 0.4505
R3296 DVDD.n2147 DVDD.n2146 0.4505
R3297 DVDD.n2664 DVDD.n2663 0.4505
R3298 DVDD.n2665 DVDD.n2145 0.4505
R3299 DVDD.n2667 DVDD.n2666 0.4505
R3300 DVDD.n2143 DVDD.n2142 0.4505
R3301 DVDD.n2676 DVDD.n2675 0.4505
R3302 DVDD.n2677 DVDD.n2141 0.4505
R3303 DVDD.n2679 DVDD.n2678 0.4505
R3304 DVDD.n2139 DVDD.n2138 0.4505
R3305 DVDD.n2867 DVDD.n2866 0.4505
R3306 DVDD.n2868 DVDD.n2137 0.4505
R3307 DVDD.n2870 DVDD.n2869 0.4505
R3308 DVDD.n2135 DVDD.n2134 0.4505
R3309 DVDD.n2875 DVDD.n2874 0.4505
R3310 DVDD.n2876 DVDD.n2133 0.4505
R3311 DVDD.n2878 DVDD.n2877 0.4505
R3312 DVDD.n2131 DVDD.n2130 0.4505
R3313 DVDD.n2883 DVDD.n2882 0.4505
R3314 DVDD.n2884 DVDD.n2129 0.4505
R3315 DVDD.n2886 DVDD.n2885 0.4505
R3316 DVDD.n2127 DVDD.n2126 0.4505
R3317 DVDD.n2891 DVDD.n2890 0.4505
R3318 DVDD.n2892 DVDD.n2125 0.4505
R3319 DVDD.n2894 DVDD.n2893 0.4505
R3320 DVDD.n2123 DVDD.n2122 0.4505
R3321 DVDD.n2899 DVDD.n2898 0.4505
R3322 DVDD.n2900 DVDD.n2121 0.4505
R3323 DVDD.n2902 DVDD.n2901 0.4505
R3324 DVDD.n2119 DVDD.n2118 0.4505
R3325 DVDD.n2907 DVDD.n2906 0.4505
R3326 DVDD.n2908 DVDD.n2117 0.4505
R3327 DVDD.n2910 DVDD.n2909 0.4505
R3328 DVDD.n2115 DVDD.n2114 0.4505
R3329 DVDD.n2915 DVDD.n2914 0.4505
R3330 DVDD.n2916 DVDD.n2113 0.4505
R3331 DVDD.n2918 DVDD.n2917 0.4505
R3332 DVDD.n2111 DVDD.n2110 0.4505
R3333 DVDD.n2923 DVDD.n2922 0.4505
R3334 DVDD.n2924 DVDD.n2109 0.4505
R3335 DVDD.n2926 DVDD.n2925 0.4505
R3336 DVDD.n2107 DVDD.n2106 0.4505
R3337 DVDD.n2931 DVDD.n2930 0.4505
R3338 DVDD.n2932 DVDD.n2105 0.4505
R3339 DVDD.n2934 DVDD.n2933 0.4505
R3340 DVDD.n2103 DVDD.n2102 0.4505
R3341 DVDD.n2939 DVDD.n2938 0.4505
R3342 DVDD.n2940 DVDD.n2100 0.4505
R3343 DVDD.n2943 DVDD.n2942 0.4505
R3344 DVDD.n2941 DVDD.n2101 0.4505
R3345 DVDD.n2087 DVDD.n2086 0.4505
R3346 DVDD.n2951 DVDD.n2950 0.4505
R3347 DVDD.n2952 DVDD.n2085 0.4505
R3348 DVDD.n2954 DVDD.n2953 0.4505
R3349 DVDD.n2083 DVDD.n2082 0.4505
R3350 DVDD.n2959 DVDD.n2958 0.4505
R3351 DVDD.n2960 DVDD.n2080 0.4505
R3352 DVDD.n3020 DVDD.n3019 0.4505
R3353 DVDD.n3018 DVDD.n2081 0.4505
R3354 DVDD.n3017 DVDD.n3016 0.4505
R3355 DVDD.n2962 DVDD.n2961 0.4505
R3356 DVDD.n3012 DVDD.n3011 0.4505
R3357 DVDD.n3010 DVDD.n2964 0.4505
R3358 DVDD.n3009 DVDD.n3008 0.4505
R3359 DVDD.n2966 DVDD.n2965 0.4505
R3360 DVDD.n3004 DVDD.n3003 0.4505
R3361 DVDD.n3002 DVDD.n2968 0.4505
R3362 DVDD.n3001 DVDD.n3000 0.4505
R3363 DVDD.n2970 DVDD.n2969 0.4505
R3364 DVDD.n2996 DVDD.n2995 0.4505
R3365 DVDD.n2994 DVDD.n2972 0.4505
R3366 DVDD.n2993 DVDD.n2992 0.4505
R3367 DVDD.n2974 DVDD.n2973 0.4505
R3368 DVDD.n2988 DVDD.n2987 0.4505
R3369 DVDD.n2986 DVDD.n2976 0.4505
R3370 DVDD.n2985 DVDD.n2984 0.4505
R3371 DVDD.n2978 DVDD.n2977 0.4505
R3372 DVDD.n2980 DVDD.n2979 0.4505
R3373 DVDD.n2982 DVDD.n2978 0.4505
R3374 DVDD.n2984 DVDD.n2983 0.4505
R3375 DVDD.n2976 DVDD.n2975 0.4505
R3376 DVDD.n2989 DVDD.n2988 0.4505
R3377 DVDD.n2990 DVDD.n2974 0.4505
R3378 DVDD.n2992 DVDD.n2991 0.4505
R3379 DVDD.n2972 DVDD.n2971 0.4505
R3380 DVDD.n2997 DVDD.n2996 0.4505
R3381 DVDD.n2998 DVDD.n2970 0.4505
R3382 DVDD.n3000 DVDD.n2999 0.4505
R3383 DVDD.n2968 DVDD.n2967 0.4505
R3384 DVDD.n3005 DVDD.n3004 0.4505
R3385 DVDD.n3006 DVDD.n2966 0.4505
R3386 DVDD.n3008 DVDD.n3007 0.4505
R3387 DVDD.n2964 DVDD.n2963 0.4505
R3388 DVDD.n3013 DVDD.n3012 0.4505
R3389 DVDD.n3014 DVDD.n2962 0.4505
R3390 DVDD.n3016 DVDD.n3015 0.4505
R3391 DVDD.n2081 DVDD.n2079 0.4505
R3392 DVDD.n3021 DVDD.n3020 0.4505
R3393 DVDD.n2080 DVDD.n2078 0.4505
R3394 DVDD.n2958 DVDD.n2957 0.4505
R3395 DVDD.n2956 DVDD.n2083 0.4505
R3396 DVDD.n2955 DVDD.n2954 0.4505
R3397 DVDD.n2085 DVDD.n2084 0.4505
R3398 DVDD.n2950 DVDD.n2949 0.4505
R3399 DVDD.n2948 DVDD.n2087 0.4505
R3400 DVDD.n2101 DVDD.n2088 0.4505
R3401 DVDD.n2944 DVDD.n2943 0.4505
R3402 DVDD.n2100 DVDD.n2099 0.4505
R3403 DVDD.n2938 DVDD.n2937 0.4505
R3404 DVDD.n2936 DVDD.n2103 0.4505
R3405 DVDD.n2935 DVDD.n2934 0.4505
R3406 DVDD.n2105 DVDD.n2104 0.4505
R3407 DVDD.n2930 DVDD.n2929 0.4505
R3408 DVDD.n2928 DVDD.n2107 0.4505
R3409 DVDD.n2927 DVDD.n2926 0.4505
R3410 DVDD.n2109 DVDD.n2108 0.4505
R3411 DVDD.n2922 DVDD.n2921 0.4505
R3412 DVDD.n2920 DVDD.n2111 0.4505
R3413 DVDD.n2919 DVDD.n2918 0.4505
R3414 DVDD.n2113 DVDD.n2112 0.4505
R3415 DVDD.n2914 DVDD.n2913 0.4505
R3416 DVDD.n2912 DVDD.n2115 0.4505
R3417 DVDD.n2911 DVDD.n2910 0.4505
R3418 DVDD.n2117 DVDD.n2116 0.4505
R3419 DVDD.n2906 DVDD.n2905 0.4505
R3420 DVDD.n2904 DVDD.n2119 0.4505
R3421 DVDD.n2903 DVDD.n2902 0.4505
R3422 DVDD.n2121 DVDD.n2120 0.4505
R3423 DVDD.n2898 DVDD.n2897 0.4505
R3424 DVDD.n2896 DVDD.n2123 0.4505
R3425 DVDD.n2895 DVDD.n2894 0.4505
R3426 DVDD.n2125 DVDD.n2124 0.4505
R3427 DVDD.n2890 DVDD.n2889 0.4505
R3428 DVDD.n2888 DVDD.n2127 0.4505
R3429 DVDD.n2887 DVDD.n2886 0.4505
R3430 DVDD.n2129 DVDD.n2128 0.4505
R3431 DVDD.n2882 DVDD.n2881 0.4505
R3432 DVDD.n2880 DVDD.n2131 0.4505
R3433 DVDD.n2879 DVDD.n2878 0.4505
R3434 DVDD.n2133 DVDD.n2132 0.4505
R3435 DVDD.n2874 DVDD.n2873 0.4505
R3436 DVDD.n2872 DVDD.n2135 0.4505
R3437 DVDD.n2871 DVDD.n2870 0.4505
R3438 DVDD.n2688 DVDD.n2137 0.4505
R3439 DVDD.n2866 DVDD.n2865 0.4505
R3440 DVDD.n2681 DVDD.n2139 0.4505
R3441 DVDD.n2680 DVDD.n2679 0.4505
R3442 DVDD.n2141 DVDD.n2140 0.4505
R3443 DVDD.n2675 DVDD.n2674 0.4505
R3444 DVDD.n2673 DVDD.n2143 0.4505
R3445 DVDD.n2668 DVDD.n2667 0.4505
R3446 DVDD.n2145 DVDD.n2144 0.4505
R3447 DVDD.n2663 DVDD.n2662 0.4505
R3448 DVDD.n2661 DVDD.n2147 0.4505
R3449 DVDD.n2660 DVDD.n2659 0.4505
R3450 DVDD.n2149 DVDD.n2148 0.4505
R3451 DVDD.n2655 DVDD.n2654 0.4505
R3452 DVDD.n2653 DVDD.n2151 0.4505
R3453 DVDD.n2652 DVDD.n2651 0.4505
R3454 DVDD.n2153 DVDD.n2152 0.4505
R3455 DVDD.n2647 DVDD.n2646 0.4505
R3456 DVDD.n2645 DVDD.n2155 0.4505
R3457 DVDD.n2644 DVDD.n2643 0.4505
R3458 DVDD.n2157 DVDD.n2156 0.4505
R3459 DVDD.n2639 DVDD.n2638 0.4505
R3460 DVDD.n2637 DVDD.n2159 0.4505
R3461 DVDD.n2636 DVDD.n2635 0.4505
R3462 DVDD.n2161 DVDD.n2160 0.4505
R3463 DVDD.n2631 DVDD.n2630 0.4505
R3464 DVDD.n2629 DVDD.n2163 0.4505
R3465 DVDD.n2628 DVDD.n2627 0.4505
R3466 DVDD.n2165 DVDD.n2164 0.4505
R3467 DVDD.n2623 DVDD.n2622 0.4505
R3468 DVDD.n2621 DVDD.n2167 0.4505
R3469 DVDD.n2611 DVDD.n2168 0.4505
R3470 DVDD.n2613 DVDD.n2612 0.4505
R3471 DVDD.n4123 DVDD.n4122 0.4505
R3472 DVDD.n3963 DVDD.n3930 0.4505
R3473 DVDD.n4077 DVDD.n4042 0.4505
R3474 DVDD.n4076 DVDD.n4075 0.4505
R3475 DVDD.n4074 DVDD.n4046 0.4505
R3476 DVDD.n4073 DVDD.n4072 0.4505
R3477 DVDD.n4048 DVDD.n4047 0.4505
R3478 DVDD.n4068 DVDD.n4067 0.4505
R3479 DVDD.n4053 DVDD.n4051 0.4505
R3480 DVDD.n4062 DVDD.n4061 0.4505
R3481 DVDD.n4058 DVDD.n4057 0.4505
R3482 DVDD.n1723 DVDD.n1721 0.4505
R3483 DVDD.n4224 DVDD.n4223 0.4505
R3484 DVDD.n1765 DVDD.n1764 0.4505
R3485 DVDD.n1729 DVDD.n1727 0.4505
R3486 DVDD.n1759 DVDD.n1758 0.4505
R3487 DVDD.n1734 DVDD.n1731 0.4505
R3488 DVDD.n1754 DVDD.n1753 0.4505
R3489 DVDD.n1752 DVDD.n1733 0.4505
R3490 DVDD.n1751 DVDD.n1750 0.4505
R3491 DVDD.n1736 DVDD.n1735 0.4505
R3492 DVDD.n1746 DVDD.n1745 0.4505
R3493 DVDD.n1744 DVDD.n1738 0.4505
R3494 DVDD.n1738 DVDD.n1737 0.4505
R3495 DVDD.n1747 DVDD.n1746 0.4505
R3496 DVDD.n1748 DVDD.n1736 0.4505
R3497 DVDD.n1750 DVDD.n1749 0.4505
R3498 DVDD.n1733 DVDD.n1732 0.4505
R3499 DVDD.n1755 DVDD.n1754 0.4505
R3500 DVDD.n1756 DVDD.n1731 0.4505
R3501 DVDD.n1758 DVDD.n1757 0.4505
R3502 DVDD.n1727 DVDD.n1726 0.4505
R3503 DVDD.n1766 DVDD.n1765 0.4505
R3504 DVDD.n4223 DVDD.n4222 0.4505
R3505 DVDD.n1725 DVDD.n1723 0.4505
R3506 DVDD.n4059 DVDD.n4058 0.4505
R3507 DVDD.n4061 DVDD.n4060 0.4505
R3508 DVDD.n4051 DVDD.n4050 0.4505
R3509 DVDD.n4069 DVDD.n4068 0.4505
R3510 DVDD.n4070 DVDD.n4048 0.4505
R3511 DVDD.n4072 DVDD.n4071 0.4505
R3512 DVDD.n4049 DVDD.n4046 0.4505
R3513 DVDD.n4076 DVDD.n4045 0.4505
R3514 DVDD.n4078 DVDD.n4077 0.4505
R3515 DVDD.n3899 DVDD.n3898 0.4505
R3516 DVDD.n3897 DVDD.n3870 0.4505
R3517 DVDD.n3896 DVDD.n3895 0.4505
R3518 DVDD.n3872 DVDD.n3871 0.4505
R3519 DVDD.n3891 DVDD.n3890 0.4505
R3520 DVDD.n3889 DVDD.n3875 0.4505
R3521 DVDD.n3888 DVDD.n3887 0.4505
R3522 DVDD.n3877 DVDD.n3876 0.4505
R3523 DVDD.n3883 DVDD.n3882 0.4505
R3524 DVDD.n3881 DVDD.n3880 0.4505
R3525 DVDD.n3879 DVDD.n1794 0.4505
R3526 DVDD.n4100 DVDD.n4099 0.4505
R3527 DVDD.n4098 DVDD.n1793 0.4505
R3528 DVDD.n4097 DVDD.n4096 0.4505
R3529 DVDD.n4035 DVDD.n4034 0.4505
R3530 DVDD.n4092 DVDD.n4091 0.4505
R3531 DVDD.n4090 DVDD.n4037 0.4505
R3532 DVDD.n4089 DVDD.n4088 0.4505
R3533 DVDD.n4039 DVDD.n4038 0.4505
R3534 DVDD.n4084 DVDD.n4083 0.4505
R3535 DVDD.n4082 DVDD.n4041 0.4505
R3536 DVDD.n4041 DVDD.n4040 0.4505
R3537 DVDD.n4085 DVDD.n4084 0.4505
R3538 DVDD.n4086 DVDD.n4039 0.4505
R3539 DVDD.n4088 DVDD.n4087 0.4505
R3540 DVDD.n4037 DVDD.n4036 0.4505
R3541 DVDD.n4093 DVDD.n4092 0.4505
R3542 DVDD.n4094 DVDD.n4035 0.4505
R3543 DVDD.n4096 DVDD.n4095 0.4505
R3544 DVDD.n1793 DVDD.n1791 0.4505
R3545 DVDD.n4101 DVDD.n4100 0.4505
R3546 DVDD.n3879 DVDD.n1790 0.4505
R3547 DVDD.n3880 DVDD.n3878 0.4505
R3548 DVDD.n3884 DVDD.n3883 0.4505
R3549 DVDD.n3885 DVDD.n3877 0.4505
R3550 DVDD.n3887 DVDD.n3886 0.4505
R3551 DVDD.n3875 DVDD.n3874 0.4505
R3552 DVDD.n3892 DVDD.n3891 0.4505
R3553 DVDD.n3893 DVDD.n3872 0.4505
R3554 DVDD.n3895 DVDD.n3894 0.4505
R3555 DVDD.n3873 DVDD.n3870 0.4505
R3556 DVDD.n3899 DVDD.n3867 0.4505
R3557 DVDD.n3903 DVDD.n3866 0.4505
R3558 DVDD.n3905 DVDD.n3904 0.4505
R3559 DVDD.n3864 DVDD.n3863 0.4505
R3560 DVDD.n3910 DVDD.n3909 0.4505
R3561 DVDD.n3911 DVDD.n3862 0.4505
R3562 DVDD.n3913 DVDD.n3912 0.4505
R3563 DVDD.n3860 DVDD.n3859 0.4505
R3564 DVDD.n3918 DVDD.n3917 0.4505
R3565 DVDD.n3919 DVDD.n3858 0.4505
R3566 DVDD.n3921 DVDD.n3920 0.4505
R3567 DVDD.n3855 DVDD.n3854 0.4505
R3568 DVDD.n3853 DVDD.n1820 0.4505
R3569 DVDD.n3852 DVDD.n3851 0.4505
R3570 DVDD.n1822 DVDD.n1821 0.4505
R3571 DVDD.n3847 DVDD.n3846 0.4505
R3572 DVDD.n3845 DVDD.n1824 0.4505
R3573 DVDD.n3844 DVDD.n3843 0.4505
R3574 DVDD.n1826 DVDD.n1825 0.4505
R3575 DVDD.n3839 DVDD.n3838 0.4505
R3576 DVDD.n3837 DVDD.n1828 0.4505
R3577 DVDD.n3836 DVDD.n3835 0.4505
R3578 DVDD.n3830 DVDD.n3829 0.4505
R3579 DVDD.n3828 DVDD.n1833 0.4505
R3580 DVDD.n3827 DVDD.n3826 0.4505
R3581 DVDD.n1835 DVDD.n1834 0.4505
R3582 DVDD.n3822 DVDD.n3821 0.4505
R3583 DVDD.n3820 DVDD.n1837 0.4505
R3584 DVDD.n3819 DVDD.n3818 0.4505
R3585 DVDD.n1839 DVDD.n1838 0.4505
R3586 DVDD.n3809 DVDD.n3808 0.4505
R3587 DVDD.n3807 DVDD.n1686 0.4505
R3588 DVDD.n4260 DVDD.n4259 0.4505
R3589 DVDD.n1678 DVDD.n1677 0.4505
R3590 DVDD.n4268 DVDD.n4267 0.4505
R3591 DVDD.n4269 DVDD.n1676 0.4505
R3592 DVDD.n4271 DVDD.n4270 0.4505
R3593 DVDD.n1674 DVDD.n1673 0.4505
R3594 DVDD.n4276 DVDD.n4275 0.4505
R3595 DVDD.n4277 DVDD.n1672 0.4505
R3596 DVDD.n4279 DVDD.n4278 0.4505
R3597 DVDD.n1669 DVDD.n1668 0.4505
R3598 DVDD.n4284 DVDD.n4283 0.4505
R3599 DVDD.n3835 DVDD.n3834 0.4505
R3600 DVDD.n1828 DVDD.n1827 0.4505
R3601 DVDD.n3840 DVDD.n3839 0.4505
R3602 DVDD.n3841 DVDD.n1826 0.4505
R3603 DVDD.n3843 DVDD.n3842 0.4505
R3604 DVDD.n1824 DVDD.n1823 0.4505
R3605 DVDD.n3848 DVDD.n3847 0.4505
R3606 DVDD.n3849 DVDD.n1822 0.4505
R3607 DVDD.n3851 DVDD.n3850 0.4505
R3608 DVDD.n1820 DVDD.n1819 0.4505
R3609 DVDD.n3856 DVDD.n3855 0.4505
R3610 DVDD.n3922 DVDD.n3921 0.4505
R3611 DVDD.n3858 DVDD.n3857 0.4505
R3612 DVDD.n3917 DVDD.n3916 0.4505
R3613 DVDD.n3915 DVDD.n3860 0.4505
R3614 DVDD.n3914 DVDD.n3913 0.4505
R3615 DVDD.n3862 DVDD.n3861 0.4505
R3616 DVDD.n3909 DVDD.n3908 0.4505
R3617 DVDD.n3907 DVDD.n3864 0.4505
R3618 DVDD.n3906 DVDD.n3905 0.4505
R3619 DVDD.n3866 DVDD.n3865 0.4505
R3620 DVDD.n4283 DVDD.n4282 0.4505
R3621 DVDD.n4281 DVDD.n1669 0.4505
R3622 DVDD.n4280 DVDD.n4279 0.4505
R3623 DVDD.n1672 DVDD.n1671 0.4505
R3624 DVDD.n4275 DVDD.n4274 0.4505
R3625 DVDD.n4273 DVDD.n1674 0.4505
R3626 DVDD.n4272 DVDD.n4271 0.4505
R3627 DVDD.n1679 DVDD.n1676 0.4505
R3628 DVDD.n4267 DVDD.n4266 0.4505
R3629 DVDD.n1681 DVDD.n1678 0.4505
R3630 DVDD.n4261 DVDD.n4260 0.4505
R3631 DVDD.n3807 DVDD.n3806 0.4505
R3632 DVDD.n3810 DVDD.n3809 0.4505
R3633 DVDD.n3811 DVDD.n1839 0.4505
R3634 DVDD.n3818 DVDD.n3817 0.4505
R3635 DVDD.n1841 DVDD.n1837 0.4505
R3636 DVDD.n3823 DVDD.n3822 0.4505
R3637 DVDD.n3824 DVDD.n1835 0.4505
R3638 DVDD.n3826 DVDD.n3825 0.4505
R3639 DVDD.n1833 DVDD.n1832 0.4505
R3640 DVDD.n3831 DVDD.n3830 0.4505
R3641 DVDD.n1571 DVDD.n1570 0.4505
R3642 DVDD.n1569 DVDD.n1206 0.4505
R3643 DVDD.n1568 DVDD.n1567 0.4505
R3644 DVDD.n1208 DVDD.n1207 0.4505
R3645 DVDD.n1563 DVDD.n1562 0.4505
R3646 DVDD.n1561 DVDD.n1211 0.4505
R3647 DVDD.n1560 DVDD.n1559 0.4505
R3648 DVDD.n1213 DVDD.n1212 0.4505
R3649 DVDD.n1226 DVDD.n1224 0.4505
R3650 DVDD.n1552 DVDD.n1551 0.4505
R3651 DVDD.n1550 DVDD.n1225 0.4505
R3652 DVDD.n1549 DVDD.n1548 0.4505
R3653 DVDD.n1228 DVDD.n1227 0.4505
R3654 DVDD.n1544 DVDD.n1543 0.4505
R3655 DVDD.n1542 DVDD.n1230 0.4505
R3656 DVDD.n1541 DVDD.n1540 0.4505
R3657 DVDD.n1232 DVDD.n1231 0.4505
R3658 DVDD.n1536 DVDD.n1535 0.4505
R3659 DVDD.n1534 DVDD.n1234 0.4505
R3660 DVDD.n1533 DVDD.n1532 0.4505
R3661 DVDD.n1236 DVDD.n1235 0.4505
R3662 DVDD.n1528 DVDD.n1527 0.4505
R3663 DVDD.n1526 DVDD.n1238 0.4505
R3664 DVDD.n1525 DVDD.n1524 0.4505
R3665 DVDD.n1240 DVDD.n1239 0.4505
R3666 DVDD.n1520 DVDD.n1519 0.4505
R3667 DVDD.n1518 DVDD.n1242 0.4505
R3668 DVDD.n1517 DVDD.n1516 0.4505
R3669 DVDD.n1244 DVDD.n1243 0.4505
R3670 DVDD.n1512 DVDD.n1511 0.4505
R3671 DVDD.n1510 DVDD.n1246 0.4505
R3672 DVDD.n1509 DVDD.n1508 0.4505
R3673 DVDD.n1248 DVDD.n1247 0.4505
R3674 DVDD.n1504 DVDD.n1503 0.4505
R3675 DVDD.n1502 DVDD.n1250 0.4505
R3676 DVDD.n1501 DVDD.n1500 0.4505
R3677 DVDD.n1252 DVDD.n1251 0.4505
R3678 DVDD.n1496 DVDD.n1495 0.4505
R3679 DVDD.n1494 DVDD.n1254 0.4505
R3680 DVDD.n1493 DVDD.n1492 0.4505
R3681 DVDD.n1256 DVDD.n1255 0.4505
R3682 DVDD.n1488 DVDD.n1487 0.4505
R3683 DVDD.n1486 DVDD.n1258 0.4505
R3684 DVDD.n1485 DVDD.n1484 0.4505
R3685 DVDD.n1260 DVDD.n1259 0.4505
R3686 DVDD.n1480 DVDD.n1479 0.4505
R3687 DVDD.n1478 DVDD.n1262 0.4505
R3688 DVDD.n1477 DVDD.n1476 0.4505
R3689 DVDD.n1264 DVDD.n1263 0.4505
R3690 DVDD.n1472 DVDD.n1471 0.4505
R3691 DVDD.n1470 DVDD.n1266 0.4505
R3692 DVDD.n1469 DVDD.n1468 0.4505
R3693 DVDD.n1268 DVDD.n1267 0.4505
R3694 DVDD.n1464 DVDD.n1463 0.4505
R3695 DVDD.n1462 DVDD.n1270 0.4505
R3696 DVDD.n1461 DVDD.n1460 0.4505
R3697 DVDD.n1272 DVDD.n1271 0.4505
R3698 DVDD.n1456 DVDD.n1455 0.4505
R3699 DVDD.n1454 DVDD.n1274 0.4505
R3700 DVDD.n1453 DVDD.n1452 0.4505
R3701 DVDD.n1276 DVDD.n1275 0.4505
R3702 DVDD.n1448 DVDD.n1447 0.4505
R3703 DVDD.n1446 DVDD.n1278 0.4505
R3704 DVDD.n1445 DVDD.n1444 0.4505
R3705 DVDD.n1280 DVDD.n1279 0.4505
R3706 DVDD.n1440 DVDD.n1439 0.4505
R3707 DVDD.n1438 DVDD.n1282 0.4505
R3708 DVDD.n1437 DVDD.n1436 0.4505
R3709 DVDD.n1284 DVDD.n1283 0.4505
R3710 DVDD.n1432 DVDD.n1431 0.4505
R3711 DVDD.n1430 DVDD.n1286 0.4505
R3712 DVDD.n1429 DVDD.n1428 0.4505
R3713 DVDD.n1288 DVDD.n1287 0.4505
R3714 DVDD.n1424 DVDD.n1423 0.4505
R3715 DVDD.n1422 DVDD.n1290 0.4505
R3716 DVDD.n1421 DVDD.n1420 0.4505
R3717 DVDD.n1292 DVDD.n1291 0.4505
R3718 DVDD.n1416 DVDD.n1415 0.4505
R3719 DVDD.n1414 DVDD.n1294 0.4505
R3720 DVDD.n1413 DVDD.n1412 0.4505
R3721 DVDD.n1296 DVDD.n1295 0.4505
R3722 DVDD.n1408 DVDD.n1407 0.4505
R3723 DVDD.n1406 DVDD.n1298 0.4505
R3724 DVDD.n1405 DVDD.n1404 0.4505
R3725 DVDD.n1300 DVDD.n1299 0.4505
R3726 DVDD.n1400 DVDD.n1399 0.4505
R3727 DVDD.n1398 DVDD.n1302 0.4505
R3728 DVDD.n1397 DVDD.n1396 0.4505
R3729 DVDD.n1304 DVDD.n1303 0.4505
R3730 DVDD.n1347 DVDD.n1346 0.4505
R3731 DVDD.n1351 DVDD.n1350 0.4505
R3732 DVDD.n1352 DVDD.n1345 0.4505
R3733 DVDD.n1354 DVDD.n1353 0.4505
R3734 DVDD.n1343 DVDD.n1342 0.4505
R3735 DVDD.n1359 DVDD.n1358 0.4505
R3736 DVDD.n1361 DVDD.n1360 0.4505
R3737 DVDD.n1205 DVDD.n1197 0.4505
R3738 DVDD.n1572 DVDD.n1571 0.4505
R3739 DVDD.n1209 DVDD.n1206 0.4505
R3740 DVDD.n1567 DVDD.n1566 0.4505
R3741 DVDD.n1565 DVDD.n1208 0.4505
R3742 DVDD.n1564 DVDD.n1563 0.4505
R3743 DVDD.n1211 DVDD.n1210 0.4505
R3744 DVDD.n1559 DVDD.n1558 0.4505
R3745 DVDD.n1557 DVDD.n1213 0.4505
R3746 DVDD.n1224 DVDD.n1218 0.4505
R3747 DVDD.n1553 DVDD.n1552 0.4505
R3748 DVDD.n1225 DVDD.n1223 0.4505
R3749 DVDD.n1548 DVDD.n1547 0.4505
R3750 DVDD.n1546 DVDD.n1228 0.4505
R3751 DVDD.n1545 DVDD.n1544 0.4505
R3752 DVDD.n1230 DVDD.n1229 0.4505
R3753 DVDD.n1540 DVDD.n1539 0.4505
R3754 DVDD.n1538 DVDD.n1232 0.4505
R3755 DVDD.n1537 DVDD.n1536 0.4505
R3756 DVDD.n1234 DVDD.n1233 0.4505
R3757 DVDD.n1532 DVDD.n1531 0.4505
R3758 DVDD.n1530 DVDD.n1236 0.4505
R3759 DVDD.n1529 DVDD.n1528 0.4505
R3760 DVDD.n1238 DVDD.n1237 0.4505
R3761 DVDD.n1524 DVDD.n1523 0.4505
R3762 DVDD.n1522 DVDD.n1240 0.4505
R3763 DVDD.n1521 DVDD.n1520 0.4505
R3764 DVDD.n1242 DVDD.n1241 0.4505
R3765 DVDD.n1516 DVDD.n1515 0.4505
R3766 DVDD.n1514 DVDD.n1244 0.4505
R3767 DVDD.n1513 DVDD.n1512 0.4505
R3768 DVDD.n1246 DVDD.n1245 0.4505
R3769 DVDD.n1508 DVDD.n1507 0.4505
R3770 DVDD.n1506 DVDD.n1248 0.4505
R3771 DVDD.n1505 DVDD.n1504 0.4505
R3772 DVDD.n1250 DVDD.n1249 0.4505
R3773 DVDD.n1500 DVDD.n1499 0.4505
R3774 DVDD.n1498 DVDD.n1252 0.4505
R3775 DVDD.n1497 DVDD.n1496 0.4505
R3776 DVDD.n1254 DVDD.n1253 0.4505
R3777 DVDD.n1492 DVDD.n1491 0.4505
R3778 DVDD.n1490 DVDD.n1256 0.4505
R3779 DVDD.n1489 DVDD.n1488 0.4505
R3780 DVDD.n1258 DVDD.n1257 0.4505
R3781 DVDD.n1484 DVDD.n1483 0.4505
R3782 DVDD.n1482 DVDD.n1260 0.4505
R3783 DVDD.n1481 DVDD.n1480 0.4505
R3784 DVDD.n1262 DVDD.n1261 0.4505
R3785 DVDD.n1476 DVDD.n1475 0.4505
R3786 DVDD.n1474 DVDD.n1264 0.4505
R3787 DVDD.n1473 DVDD.n1472 0.4505
R3788 DVDD.n1266 DVDD.n1265 0.4505
R3789 DVDD.n1468 DVDD.n1467 0.4505
R3790 DVDD.n1466 DVDD.n1268 0.4505
R3791 DVDD.n1465 DVDD.n1464 0.4505
R3792 DVDD.n1270 DVDD.n1269 0.4505
R3793 DVDD.n1460 DVDD.n1459 0.4505
R3794 DVDD.n1458 DVDD.n1272 0.4505
R3795 DVDD.n1457 DVDD.n1456 0.4505
R3796 DVDD.n1274 DVDD.n1273 0.4505
R3797 DVDD.n1452 DVDD.n1451 0.4505
R3798 DVDD.n1450 DVDD.n1276 0.4505
R3799 DVDD.n1449 DVDD.n1448 0.4505
R3800 DVDD.n1278 DVDD.n1277 0.4505
R3801 DVDD.n1444 DVDD.n1443 0.4505
R3802 DVDD.n1442 DVDD.n1280 0.4505
R3803 DVDD.n1441 DVDD.n1440 0.4505
R3804 DVDD.n1282 DVDD.n1281 0.4505
R3805 DVDD.n1436 DVDD.n1435 0.4505
R3806 DVDD.n1434 DVDD.n1284 0.4505
R3807 DVDD.n1433 DVDD.n1432 0.4505
R3808 DVDD.n1286 DVDD.n1285 0.4505
R3809 DVDD.n1428 DVDD.n1427 0.4505
R3810 DVDD.n1426 DVDD.n1288 0.4505
R3811 DVDD.n1425 DVDD.n1424 0.4505
R3812 DVDD.n1290 DVDD.n1289 0.4505
R3813 DVDD.n1420 DVDD.n1419 0.4505
R3814 DVDD.n1418 DVDD.n1292 0.4505
R3815 DVDD.n1417 DVDD.n1416 0.4505
R3816 DVDD.n1294 DVDD.n1293 0.4505
R3817 DVDD.n1412 DVDD.n1411 0.4505
R3818 DVDD.n1410 DVDD.n1296 0.4505
R3819 DVDD.n1409 DVDD.n1408 0.4505
R3820 DVDD.n1298 DVDD.n1297 0.4505
R3821 DVDD.n1404 DVDD.n1403 0.4505
R3822 DVDD.n1402 DVDD.n1300 0.4505
R3823 DVDD.n1401 DVDD.n1400 0.4505
R3824 DVDD.n1302 DVDD.n1301 0.4505
R3825 DVDD.n1396 DVDD.n1395 0.4505
R3826 DVDD.n1310 DVDD.n1304 0.4505
R3827 DVDD.n1348 DVDD.n1347 0.4505
R3828 DVDD.n1350 DVDD.n1349 0.4505
R3829 DVDD.n1345 DVDD.n1344 0.4505
R3830 DVDD.n1355 DVDD.n1354 0.4505
R3831 DVDD.n1356 DVDD.n1343 0.4505
R3832 DVDD.n1358 DVDD.n1357 0.4505
R3833 DVDD.n1361 DVDD.n1337 0.4505
R3834 DVDD.n1362 DVDD.n1340 0.4505
R3835 DVDD.n2798 DVDD.n2797 0.449506
R3836 DVDD.n1924 DVDD 0.448132
R3837 DVDD.n3343 DVDD.n3342 0.440554
R3838 DVDD DVDD.n2239 0.4405
R3839 DVDD.n4342 DVDD.n4299 0.437225
R3840 DVDD.n1934 DVDD.n1933 0.427206
R3841 DVDD.n2671 DVDD.n2670 0.423396
R3842 DVDD.n4237 DVDD.n4236 0.4205
R3843 DVDD.n4234 DVDD.n4233 0.4205
R3844 DVDD.n2217 DVDD.n2216 0.417167
R3845 DVDD.n2221 DVDD.n2220 0.417167
R3846 DVDD.n2225 DVDD.n2224 0.417167
R3847 DVDD.n2229 DVDD.n2228 0.417167
R3848 DVDD.n2233 DVDD.n2232 0.417167
R3849 DVDD.n2237 DVDD.n2236 0.417167
R3850 DVDD.n2238 DVDD.n2235 0.417167
R3851 DVDD.n2234 DVDD.n2231 0.417167
R3852 DVDD.n2230 DVDD.n2227 0.417167
R3853 DVDD.n2226 DVDD.n2223 0.417167
R3854 DVDD.n2222 DVDD.n2219 0.417167
R3855 DVDD.n2218 DVDD.n2215 0.417167
R3856 DVDD DVDD.n2325 0.414765
R3857 DVDD.n2463 DVDD 0.414765
R3858 DVDD DVDD.n2261 0.414765
R3859 DVDD.n2538 DVDD 0.414765
R3860 DVDD.n1881 DVDD.n1879 0.413789
R3861 DVDD.n3394 DVDD.n3393 0.41077
R3862 DVDD.n3348 DVDD.n3346 0.41077
R3863 DVDD.n3320 DVDD.n3245 0.41077
R3864 DVDD.n3329 DVDD.n3322 0.41077
R3865 DVDD.n2799 DVDD.n2705 0.402145
R3866 DVDD.n2734 DVDD.n2705 0.399579
R3867 DVDD DVDD.n1710 0.397559
R3868 DVDD DVDD.n1710 0.397559
R3869 DVDD.n3395 DVDD.n3394 0.391716
R3870 DVDD.n3349 DVDD.n3348 0.391716
R3871 DVDD.n3379 DVDD.n3378 0.376594
R3872 DVDD.n3335 DVDD.n3313 0.376594
R3873 DVDD.n3375 DVDD.n3374 0.3755
R3874 DVDD.n3325 DVDD.n3271 0.3755
R3875 DVDD.n3328 DVDD.n3327 0.3755
R3876 DVDD.n3249 DVDD.n3244 0.3755
R3877 DVDD.n1934 DVDD.n1924 0.36126
R3878 DVDD.t191 DVDD.n1883 0.3605
R3879 DVDD.t197 DVDD.n1709 0.3605
R3880 DVDD.t63 DVDD.n1711 0.3605
R3881 DVDD.t111 DVDD.n4188 0.3605
R3882 DVDD.n4136 DVDD.t166 0.360167
R3883 DVDD.n1785 DVDD.t184 0.360167
R3884 DVDD.n3964 DVDD.t106 0.360167
R3885 DVDD.n3960 DVDD.t108 0.360167
R3886 DVDD.n1874 DVDD.t1 0.360167
R3887 DVDD.n1872 DVDD.t35 0.360167
R3888 DVDD.n1714 DVDD.t170 0.360167
R3889 DVDD.n1717 DVDD.t172 0.360167
R3890 DVDD.n1904 DVDD.n1896 0.356801
R3891 DVDD.n1946 DVDD.n1896 0.356801
R3892 DVDD.n3652 DVDD.n1986 0.35585
R3893 DVDD.n3652 DVDD.n1994 0.35585
R3894 DVDD.n3652 DVDD.n1988 0.35585
R3895 DVDD.n4081 DVDD.n4080 0.35585
R3896 DVDD.n3901 DVDD.n3869 0.35585
R3897 DVDD.n4081 DVDD.n4043 0.355001
R3898 DVDD.n1898 DVDD.n1896 0.35492
R3899 DVDD.n3617 DVDD.n3087 0.35492
R3900 DVDD.n3617 DVDD.n3094 0.35492
R3901 DVDD.n3833 DVDD.n3832 0.35492
R3902 DVDD.n3869 DVDD.n3868 0.354416
R3903 DVDD.n1945 DVDD.n1896 0.35405
R3904 DVDD.n1967 DVDD.n1896 0.35405
R3905 DVDD.n3652 DVDD.n1982 0.353477
R3906 DVDD.n3652 DVDD.n1987 0.353477
R3907 DVDD.n3652 DVDD.n1989 0.353477
R3908 DVDD.n3617 DVDD.n3088 0.35312
R3909 DVDD.n3617 DVDD.n3093 0.35312
R3910 DVDD.n3833 DVDD.n1831 0.35312
R3911 DVDD.n2075 DVDD.n2074 0.346654
R3912 DVDD.n3066 DVDD.n3065 0.346654
R3913 DVDD.n1881 DVDD.n1880 0.346654
R3914 DVDD.n4228 DVDD.n4227 0.346654
R3915 DVDD.n3704 DVDD.n1904 0.340118
R3916 DVDD.n3704 DVDD.n1946 0.340118
R3917 DVDD.n3704 DVDD.n1898 0.339393
R3918 DVDD.n3094 DVDD.n2022 0.339393
R3919 DVDD.n3087 DVDD.n2022 0.339393
R3920 DVDD.n3832 DVDD.n1829 0.339393
R3921 DVDD.n4079 DVDD.n4043 0.338918
R3922 DVDD.n3902 DVDD.n3868 0.33857
R3923 DVDD.n3647 DVDD.n1986 0.338454
R3924 DVDD.n3647 DVDD.n1994 0.338454
R3925 DVDD.n3647 DVDD.n1988 0.338454
R3926 DVDD.n4080 DVDD.n4079 0.338454
R3927 DVDD.n3902 DVDD.n3901 0.338454
R3928 DVDD.n1831 DVDD.n1829 0.338193
R3929 DVDD.n3093 DVDD.n2022 0.338193
R3930 DVDD.n3088 DVDD.n2022 0.338193
R3931 DVDD.n3647 DVDD.n1987 0.337829
R3932 DVDD.n3647 DVDD.n1989 0.337829
R3933 DVDD.n3647 DVDD.n1982 0.337829
R3934 DVDD.n2788 DVDD.n2724 0.337345
R3935 DVDD.n2738 DVDD.n2733 0.337345
R3936 DVDD.n2786 DVDD.n2741 0.337345
R3937 DVDD.n2783 DVDD.n2781 0.337345
R3938 DVDD.n2777 DVDD.n2747 0.337345
R3939 DVDD.n2775 DVDD.n2760 0.337345
R3940 DVDD.n2754 DVDD.n2751 0.337345
R3941 DVDD.n2766 DVDD.n2755 0.337345
R3942 DVDD.n2765 DVDD.n2752 0.337345
R3943 DVDD.n2764 DVDD.n2753 0.337345
R3944 DVDD.n2766 DVDD.n2752 0.337345
R3945 DVDD.n2760 DVDD.n2751 0.337345
R3946 DVDD.n2759 DVDD.n2747 0.337345
R3947 DVDD.n2783 DVDD.n2741 0.337345
R3948 DVDD.n2733 DVDD.n2724 0.337345
R3949 DVDD.n2769 DVDD.n2765 0.337345
R3950 DVDD.n2755 DVDD.n2754 0.337345
R3951 DVDD.n2786 DVDD.n2738 0.337345
R3952 DVDD.n2781 DVDD.n2737 0.337345
R3953 DVDD.n2769 DVDD.n2753 0.337345
R3954 DVDD.n3704 DVDD.n1945 0.337254
R3955 DVDD.n3704 DVDD.n1967 0.337254
R3956 DVDD.n3342 DVDD.n2022 0.327632
R3957 DVDD.n4228 DVDD.n1718 0.313132
R3958 DVDD.n4148 DVDD.n4147 0.306049
R3959 DVDD.n1873 DVDD.n1706 0.306049
R3960 DVDD.n3959 DVDD.n3958 0.306049
R3961 DVDD.n4138 DVDD.n4137 0.306049
R3962 DVDD.n1955 DVDD.t194 0.303833
R3963 DVDD.n1955 DVDD.t156 0.303833
R3964 DVDD.n1951 DVDD.t46 0.303833
R3965 DVDD.n1951 DVDD.t174 0.303833
R3966 DVDD.n1917 DVDD.t110 0.303833
R3967 DVDD.n1917 DVDD.t200 0.303833
R3968 DVDD.n1918 DVDD.t69 0.303833
R3969 DVDD.n1918 DVDD.t66 0.303833
R3970 DVDD.n85 DVDD.n84 0.3005
R3971 DVDD.n333 DVDD.n329 0.3005
R3972 DVDD.n2787 DVDD.n2736 0.291153
R3973 DVDD.n1875 DVDD.n1708 0.265206
R3974 DVDD.n3961 DVDD.n1708 0.265206
R3975 DVDD.n4232 DVDD.n1713 0.265206
R3976 DVDD.n4232 DVDD.n4231 0.265206
R3977 DVDD.n2798 DVDD.n2702 0.260889
R3978 DVDD.n1959 DVDD 0.258658
R3979 DVDD.n2713 DVDD.n2712 0.252737
R3980 DVDD.n5504 DVDD.n219 0.2505
R3981 DVDD.n966 DVDD.n945 0.2505
R3982 DVDD.n3375 DVDD.n3244 0.242734
R3983 DVDD.n3327 DVDD.n3325 0.242734
R3984 DVDD.n2214 DVDD 0.232667
R3985 DVDD.n3376 DVDD.n3375 0.231484
R3986 DVDD.n3327 DVDD.n3326 0.231484
R3987 DVDD.n2594 DVDD.n2240 0.231338
R3988 DVDD.n2610 DVDD.n2604 0.231338
R3989 DVDD.n5915 DVDD.n103 0.22706
R3990 DVDD.n5420 DVDD.n5418 0.225937
R3991 DVDD.n928 DVDD.n263 0.224497
R3992 DVDD.n259 DVDD.n258 0.224242
R3993 DVDD.n2670 DVDD 0.224176
R3994 DVDD.n3775 DVDD.n3721 0.221159
R3995 DVDD.n1150 DVDD.n1120 0.221159
R3996 DVDD.n4411 DVDD.n4399 0.221159
R3997 DVDD.n4345 DVDD.n1595 0.221159
R3998 DVDD.n4300 DVDD.n1627 0.221159
R3999 DVDD.n3368 DVDD.n3273 0.218429
R4000 DVDD.n3372 DVDD.n3247 0.218429
R4001 DVDD.n2047 DVDD.n2044 0.217739
R4002 DVDD.n5687 DVDD.n5686 0.214786
R4003 DVDD.n5685 DVDD.n5684 0.214786
R4004 DVDD.n5691 DVDD.n5683 0.214786
R4005 DVDD.n5692 DVDD.n5682 0.214786
R4006 DVDD.n5693 DVDD.n5681 0.214786
R4007 DVDD.n5680 DVDD.n5678 0.214786
R4008 DVDD.n5697 DVDD.n5677 0.214786
R4009 DVDD.n5698 DVDD.n5676 0.214786
R4010 DVDD.n5699 DVDD.n5675 0.214786
R4011 DVDD.n5700 DVDD.n5674 0.214786
R4012 DVDD.n5673 DVDD.n217 0.214786
R4013 DVDD.n5709 DVDD.n216 0.214786
R4014 DVDD.n5712 DVDD.n215 0.214786
R4015 DVDD.n5713 DVDD.n214 0.214786
R4016 DVDD.n5714 DVDD.n213 0.214786
R4017 DVDD.n212 DVDD.n210 0.214786
R4018 DVDD.n5718 DVDD.n209 0.214786
R4019 DVDD.n5719 DVDD.n208 0.214786
R4020 DVDD.n5720 DVDD.n207 0.214786
R4021 DVDD.n206 DVDD.n204 0.214786
R4022 DVDD.n5724 DVDD.n203 0.214786
R4023 DVDD.n5725 DVDD.n202 0.214786
R4024 DVDD.n5726 DVDD.n201 0.214786
R4025 DVDD.n5065 DVDD.n200 0.214786
R4026 DVDD.n5067 DVDD.n5066 0.214786
R4027 DVDD.n5064 DVDD.n5063 0.214786
R4028 DVDD.n5071 DVDD.n5062 0.214786
R4029 DVDD.n5072 DVDD.n5061 0.214786
R4030 DVDD.n5073 DVDD.n5060 0.214786
R4031 DVDD.n5059 DVDD.n5057 0.214786
R4032 DVDD.n5077 DVDD.n5056 0.214786
R4033 DVDD.n5078 DVDD.n5055 0.214786
R4034 DVDD.n5079 DVDD.n5054 0.214786
R4035 DVDD.n5053 DVDD.n5051 0.214786
R4036 DVDD.n5083 DVDD.n5050 0.214786
R4037 DVDD.n5084 DVDD.n5049 0.214786
R4038 DVDD.n5047 DVDD.n5046 0.214786
R4039 DVDD.n575 DVDD.n574 0.214786
R4040 DVDD.n5042 DVDD.n5041 0.214786
R4041 DVDD.n5040 DVDD.n577 0.214786
R4042 DVDD.n5039 DVDD.n5038 0.214786
R4043 DVDD.n579 DVDD.n578 0.214786
R4044 DVDD.n5034 DVDD.n5033 0.214786
R4045 DVDD.n5032 DVDD.n581 0.214786
R4046 DVDD.n5031 DVDD.n5030 0.214786
R4047 DVDD.n583 DVDD.n582 0.214786
R4048 DVDD.n5026 DVDD.n5025 0.214786
R4049 DVDD.n5024 DVDD.n585 0.214786
R4050 DVDD.n5023 DVDD.n5022 0.214786
R4051 DVDD.n587 DVDD.n586 0.214786
R4052 DVDD.n4786 DVDD.n4785 0.214786
R4053 DVDD.n4789 DVDD.n4784 0.214786
R4054 DVDD.n4790 DVDD.n4783 0.214786
R4055 DVDD.n4791 DVDD.n4782 0.214786
R4056 DVDD.n4781 DVDD.n4779 0.214786
R4057 DVDD.n4795 DVDD.n4778 0.214786
R4058 DVDD.n4796 DVDD.n4777 0.214786
R4059 DVDD.n4797 DVDD.n4776 0.214786
R4060 DVDD.n4775 DVDD.n734 0.214786
R4061 DVDD.n4801 DVDD.n733 0.214786
R4062 DVDD.n4766 DVDD.n732 0.214786
R4063 DVDD.n4768 DVDD.n4767 0.214786
R4064 DVDD.n4764 DVDD.n880 0.214786
R4065 DVDD.n4763 DVDD.n4762 0.214786
R4066 DVDD.n882 DVDD.n881 0.214786
R4067 DVDD.n4758 DVDD.n4757 0.214786
R4068 DVDD.n4756 DVDD.n884 0.214786
R4069 DVDD.n4755 DVDD.n4754 0.214786
R4070 DVDD.n886 DVDD.n885 0.214786
R4071 DVDD.n4750 DVDD.n4749 0.214786
R4072 DVDD.n4748 DVDD.n888 0.214786
R4073 DVDD.n4747 DVDD.n4746 0.214786
R4074 DVDD.n890 DVDD.n889 0.214786
R4075 DVDD.n4740 DVDD.n4739 0.214786
R4076 DVDD.n4738 DVDD.n898 0.214786
R4077 DVDD.n4737 DVDD.n4736 0.214786
R4078 DVDD.n900 DVDD.n899 0.214786
R4079 DVDD.n4732 DVDD.n4731 0.214786
R4080 DVDD.n4730 DVDD.n902 0.214786
R4081 DVDD.n4729 DVDD.n4728 0.214786
R4082 DVDD.n904 DVDD.n903 0.214786
R4083 DVDD.n4724 DVDD.n4723 0.214786
R4084 DVDD.n4722 DVDD.n906 0.214786
R4085 DVDD.n4721 DVDD.n4720 0.214786
R4086 DVDD.n4328 DVDD.n4301 0.214786
R4087 DVDD.n4327 DVDD.n4302 0.214786
R4088 DVDD.n4326 DVDD.n4303 0.214786
R4089 DVDD.n4306 DVDD.n4304 0.214786
R4090 DVDD.n4322 DVDD.n4307 0.214786
R4091 DVDD.n4321 DVDD.n4308 0.214786
R4092 DVDD.n4320 DVDD.n4309 0.214786
R4093 DVDD.n4312 DVDD.n4310 0.214786
R4094 DVDD.n4316 DVDD.n4313 0.214786
R4095 DVDD.n4315 DVDD.n4314 0.214786
R4096 DVDD.n913 DVDD.n912 0.214786
R4097 DVDD.n4713 DVDD.n4712 0.214786
R4098 DVDD.n4714 DVDD.n911 0.214786
R4099 DVDD.n4716 DVDD.n4715 0.214786
R4100 DVDD.n5970 DVDD.n5969 0.214786
R4101 DVDD.n5968 DVDD.n5967 0.214786
R4102 DVDD.n5966 DVDD.n1 0.214786
R4103 DVDD.n5960 DVDD.n2 0.214786
R4104 DVDD.n5962 DVDD.n5961 0.214786
R4105 DVDD.n5959 DVDD.n4 0.214786
R4106 DVDD.n5958 DVDD.n5957 0.214786
R4107 DVDD.n6 DVDD.n5 0.214786
R4108 DVDD.n5947 DVDD.n5946 0.214786
R4109 DVDD.n5949 DVDD.n5945 0.214786
R4110 DVDD.n5950 DVDD.n5944 0.214786
R4111 DVDD.n5943 DVDD.n33 0.214786
R4112 DVDD.n5941 DVDD.n5940 0.214786
R4113 DVDD.n37 DVDD.n36 0.214786
R4114 DVDD.n526 DVDD.n524 0.214786
R4115 DVDD.n527 DVDD.n523 0.214786
R4116 DVDD.n528 DVDD.n522 0.214786
R4117 DVDD.n521 DVDD.n519 0.214786
R4118 DVDD.n532 DVDD.n518 0.214786
R4119 DVDD.n533 DVDD.n517 0.214786
R4120 DVDD.n534 DVDD.n516 0.214786
R4121 DVDD.n515 DVDD.n513 0.214786
R4122 DVDD.n538 DVDD.n512 0.214786
R4123 DVDD.n539 DVDD.n511 0.214786
R4124 DVDD.n540 DVDD.n510 0.214786
R4125 DVDD.n541 DVDD.n509 0.214786
R4126 DVDD.n508 DVDD.n507 0.214786
R4127 DVDD.n545 DVDD.n506 0.214786
R4128 DVDD.n546 DVDD.n505 0.214786
R4129 DVDD.n547 DVDD.n504 0.214786
R4130 DVDD.n503 DVDD.n501 0.214786
R4131 DVDD.n551 DVDD.n500 0.214786
R4132 DVDD.n552 DVDD.n499 0.214786
R4133 DVDD.n553 DVDD.n498 0.214786
R4134 DVDD.n497 DVDD.n484 0.214786
R4135 DVDD.n5244 DVDD.n483 0.214786
R4136 DVDD.n4833 DVDD.n482 0.214786
R4137 DVDD.n4835 DVDD.n4834 0.214786
R4138 DVDD.n4839 DVDD.n4832 0.214786
R4139 DVDD.n4840 DVDD.n4831 0.214786
R4140 DVDD.n4841 DVDD.n4830 0.214786
R4141 DVDD.n4829 DVDD.n4827 0.214786
R4142 DVDD.n4845 DVDD.n4826 0.214786
R4143 DVDD.n4846 DVDD.n4825 0.214786
R4144 DVDD.n4847 DVDD.n4824 0.214786
R4145 DVDD.n4823 DVDD.n4821 0.214786
R4146 DVDD.n4851 DVDD.n4820 0.214786
R4147 DVDD.n4852 DVDD.n4819 0.214786
R4148 DVDD.n4853 DVDD.n4818 0.214786
R4149 DVDD.n4854 DVDD.n4817 0.214786
R4150 DVDD.n4857 DVDD.n4816 0.214786
R4151 DVDD.n4858 DVDD.n4815 0.214786
R4152 DVDD.n4859 DVDD.n4814 0.214786
R4153 DVDD.n4813 DVDD.n4811 0.214786
R4154 DVDD.n4863 DVDD.n4810 0.214786
R4155 DVDD.n4864 DVDD.n4809 0.214786
R4156 DVDD.n4865 DVDD.n4808 0.214786
R4157 DVDD.n4807 DVDD.n4805 0.214786
R4158 DVDD.n4869 DVDD.n4804 0.214786
R4159 DVDD.n4870 DVDD.n4803 0.214786
R4160 DVDD.n4872 DVDD.n731 0.214786
R4161 DVDD.n4873 DVDD.n730 0.214786
R4162 DVDD.n1031 DVDD.n729 0.214786
R4163 DVDD.n1033 DVDD.n1032 0.214786
R4164 DVDD.n1036 DVDD.n1030 0.214786
R4165 DVDD.n1037 DVDD.n1029 0.214786
R4166 DVDD.n1038 DVDD.n1028 0.214786
R4167 DVDD.n1027 DVDD.n1025 0.214786
R4168 DVDD.n1042 DVDD.n1024 0.214786
R4169 DVDD.n1043 DVDD.n1023 0.214786
R4170 DVDD.n1044 DVDD.n1022 0.214786
R4171 DVDD.n1021 DVDD.n1009 0.214786
R4172 DVDD.n4617 DVDD.n1008 0.214786
R4173 DVDD.n4618 DVDD.n1007 0.214786
R4174 DVDD.n1006 DVDD.n1004 0.214786
R4175 DVDD.n4622 DVDD.n1003 0.214786
R4176 DVDD.n4623 DVDD.n1002 0.214786
R4177 DVDD.n4624 DVDD.n1001 0.214786
R4178 DVDD.n1000 DVDD.n998 0.214786
R4179 DVDD.n4628 DVDD.n997 0.214786
R4180 DVDD.n4629 DVDD.n996 0.214786
R4181 DVDD.n4630 DVDD.n995 0.214786
R4182 DVDD.n994 DVDD.n992 0.214786
R4183 DVDD.n4634 DVDD.n991 0.214786
R4184 DVDD.n4637 DVDD.n989 0.214786
R4185 DVDD.n4639 DVDD.n988 0.214786
R4186 DVDD.n4641 DVDD.n987 0.214786
R4187 DVDD.n4642 DVDD.n986 0.214786
R4188 DVDD.n4357 DVDD.n985 0.214786
R4189 DVDD.n4359 DVDD.n4358 0.214786
R4190 DVDD.n4356 DVDD.n4355 0.214786
R4191 DVDD.n4363 DVDD.n4354 0.214786
R4192 DVDD.n4364 DVDD.n4353 0.214786
R4193 DVDD.n4365 DVDD.n4352 0.214786
R4194 DVDD.n4351 DVDD.n4349 0.214786
R4195 DVDD.n4369 DVDD.n4348 0.214786
R4196 DVDD.n4370 DVDD.n4347 0.214786
R4197 DVDD.n4371 DVDD.n4346 0.214786
R4198 DVDD.n5589 DVDD.n5588 0.214786
R4199 DVDD.n5592 DVDD.n5587 0.214786
R4200 DVDD.n5593 DVDD.n5586 0.214786
R4201 DVDD.n5594 DVDD.n5585 0.214786
R4202 DVDD.n5584 DVDD.n5582 0.214786
R4203 DVDD.n5598 DVDD.n5581 0.214786
R4204 DVDD.n5599 DVDD.n5580 0.214786
R4205 DVDD.n5600 DVDD.n5579 0.214786
R4206 DVDD.n5578 DVDD.n5576 0.214786
R4207 DVDD.n5577 DVDD.n47 0.214786
R4208 DVDD.n5934 DVDD.n46 0.214786
R4209 DVDD.n5935 DVDD.n45 0.214786
R4210 DVDD.n5282 DVDD.n5281 0.214786
R4211 DVDD.n5284 DVDD.n5280 0.214786
R4212 DVDD.n5285 DVDD.n5279 0.214786
R4213 DVDD.n5286 DVDD.n5278 0.214786
R4214 DVDD.n5277 DVDD.n5275 0.214786
R4215 DVDD.n5290 DVDD.n5274 0.214786
R4216 DVDD.n5291 DVDD.n5273 0.214786
R4217 DVDD.n5292 DVDD.n5272 0.214786
R4218 DVDD.n5271 DVDD.n5269 0.214786
R4219 DVDD.n5296 DVDD.n5268 0.214786
R4220 DVDD.n5297 DVDD.n5267 0.214786
R4221 DVDD.n5298 DVDD.n5266 0.214786
R4222 DVDD.n5300 DVDD.n5265 0.214786
R4223 DVDD.n5301 DVDD.n5264 0.214786
R4224 DVDD.n5302 DVDD.n5263 0.214786
R4225 DVDD.n5262 DVDD.n5260 0.214786
R4226 DVDD.n5306 DVDD.n5259 0.214786
R4227 DVDD.n5307 DVDD.n5258 0.214786
R4228 DVDD.n5308 DVDD.n5257 0.214786
R4229 DVDD.n5256 DVDD.n5254 0.214786
R4230 DVDD.n5312 DVDD.n5253 0.214786
R4231 DVDD.n5313 DVDD.n5252 0.214786
R4232 DVDD.n5314 DVDD.n5251 0.214786
R4233 DVDD.n5250 DVDD.n476 0.214786
R4234 DVDD.n5248 DVDD.n5247 0.214786
R4235 DVDD.n480 DVDD.n479 0.214786
R4236 DVDD.n4924 DVDD.n4921 0.214786
R4237 DVDD.n4925 DVDD.n4920 0.214786
R4238 DVDD.n4926 DVDD.n4919 0.214786
R4239 DVDD.n4918 DVDD.n4916 0.214786
R4240 DVDD.n4930 DVDD.n4915 0.214786
R4241 DVDD.n4931 DVDD.n4914 0.214786
R4242 DVDD.n4932 DVDD.n4913 0.214786
R4243 DVDD.n4912 DVDD.n4910 0.214786
R4244 DVDD.n4936 DVDD.n4909 0.214786
R4245 DVDD.n4937 DVDD.n4908 0.214786
R4246 DVDD.n4907 DVDD.n684 0.214786
R4247 DVDD.n4906 DVDD.n4905 0.214786
R4248 DVDD.n686 DVDD.n685 0.214786
R4249 DVDD.n4901 DVDD.n4900 0.214786
R4250 DVDD.n4899 DVDD.n688 0.214786
R4251 DVDD.n4898 DVDD.n4897 0.214786
R4252 DVDD.n690 DVDD.n689 0.214786
R4253 DVDD.n4893 DVDD.n4892 0.214786
R4254 DVDD.n4891 DVDD.n692 0.214786
R4255 DVDD.n4890 DVDD.n4889 0.214786
R4256 DVDD.n694 DVDD.n693 0.214786
R4257 DVDD.n4885 DVDD.n4884 0.214786
R4258 DVDD.n4882 DVDD.n4881 0.214786
R4259 DVDD.n701 DVDD.n700 0.214786
R4260 DVDD.n4479 DVDD.n4478 0.214786
R4261 DVDD.n4483 DVDD.n4477 0.214786
R4262 DVDD.n4484 DVDD.n4476 0.214786
R4263 DVDD.n4485 DVDD.n4475 0.214786
R4264 DVDD.n4474 DVDD.n4472 0.214786
R4265 DVDD.n4489 DVDD.n4471 0.214786
R4266 DVDD.n4490 DVDD.n4470 0.214786
R4267 DVDD.n4491 DVDD.n4469 0.214786
R4268 DVDD.n4468 DVDD.n4466 0.214786
R4269 DVDD.n4495 DVDD.n4465 0.214786
R4270 DVDD.n4496 DVDD.n4464 0.214786
R4271 DVDD.n4463 DVDD.n1085 0.214786
R4272 DVDD.n4462 DVDD.n4461 0.214786
R4273 DVDD.n1087 DVDD.n1086 0.214786
R4274 DVDD.n4457 DVDD.n4456 0.214786
R4275 DVDD.n4455 DVDD.n1089 0.214786
R4276 DVDD.n4454 DVDD.n4453 0.214786
R4277 DVDD.n1091 DVDD.n1090 0.214786
R4278 DVDD.n4449 DVDD.n4448 0.214786
R4279 DVDD.n4447 DVDD.n1093 0.214786
R4280 DVDD.n4446 DVDD.n4445 0.214786
R4281 DVDD.n4442 DVDD.n4441 0.214786
R4282 DVDD.n4439 DVDD.n4438 0.214786
R4283 DVDD.n4437 DVDD.n1096 0.214786
R4284 DVDD.n4436 DVDD.n4435 0.214786
R4285 DVDD.n4434 DVDD.n1097 0.214786
R4286 DVDD.n4433 DVDD.n4432 0.214786
R4287 DVDD.n1099 DVDD.n1098 0.214786
R4288 DVDD.n4428 DVDD.n4427 0.214786
R4289 DVDD.n4426 DVDD.n1101 0.214786
R4290 DVDD.n4425 DVDD.n4424 0.214786
R4291 DVDD.n1103 DVDD.n1102 0.214786
R4292 DVDD.n4420 DVDD.n4419 0.214786
R4293 DVDD.n4418 DVDD.n1105 0.214786
R4294 DVDD.n4417 DVDD.n4416 0.214786
R4295 DVDD.n1107 DVDD.n1106 0.214786
R4296 DVDD.n5895 DVDD.n5894 0.214786
R4297 DVDD.n5898 DVDD.n5893 0.214786
R4298 DVDD.n5899 DVDD.n5892 0.214786
R4299 DVDD.n5900 DVDD.n5891 0.214786
R4300 DVDD.n5890 DVDD.n5888 0.214786
R4301 DVDD.n5904 DVDD.n5887 0.214786
R4302 DVDD.n5905 DVDD.n5886 0.214786
R4303 DVDD.n5906 DVDD.n5885 0.214786
R4304 DVDD.n5884 DVDD.n117 0.214786
R4305 DVDD.n5883 DVDD.n5882 0.214786
R4306 DVDD.n5880 DVDD.n118 0.214786
R4307 DVDD.n5879 DVDD.n5878 0.214786
R4308 DVDD.n5876 DVDD.n5875 0.214786
R4309 DVDD.n121 DVDD.n120 0.214786
R4310 DVDD.n5871 DVDD.n5870 0.214786
R4311 DVDD.n5869 DVDD.n123 0.214786
R4312 DVDD.n5868 DVDD.n5867 0.214786
R4313 DVDD.n125 DVDD.n124 0.214786
R4314 DVDD.n5863 DVDD.n5862 0.214786
R4315 DVDD.n5861 DVDD.n127 0.214786
R4316 DVDD.n5860 DVDD.n5859 0.214786
R4317 DVDD.n129 DVDD.n128 0.214786
R4318 DVDD.n5855 DVDD.n5854 0.214786
R4319 DVDD.n5853 DVDD.n131 0.214786
R4320 DVDD.n5852 DVDD.n5851 0.214786
R4321 DVDD.n133 DVDD.n132 0.214786
R4322 DVDD.n5120 DVDD.n5119 0.214786
R4323 DVDD.n5118 DVDD.n5117 0.214786
R4324 DVDD.n5124 DVDD.n5116 0.214786
R4325 DVDD.n5125 DVDD.n5115 0.214786
R4326 DVDD.n5126 DVDD.n5114 0.214786
R4327 DVDD.n5113 DVDD.n5111 0.214786
R4328 DVDD.n5130 DVDD.n5110 0.214786
R4329 DVDD.n5131 DVDD.n5109 0.214786
R4330 DVDD.n5132 DVDD.n5108 0.214786
R4331 DVDD.n5107 DVDD.n5106 0.214786
R4332 DVDD.n5322 DVDD.n447 0.214786
R4333 DVDD.n5323 DVDD.n446 0.214786
R4334 DVDD.n5324 DVDD.n445 0.214786
R4335 DVDD.n444 DVDD.n442 0.214786
R4336 DVDD.n5328 DVDD.n441 0.214786
R4337 DVDD.n5329 DVDD.n440 0.214786
R4338 DVDD.n5330 DVDD.n439 0.214786
R4339 DVDD.n438 DVDD.n436 0.214786
R4340 DVDD.n5334 DVDD.n435 0.214786
R4341 DVDD.n5335 DVDD.n434 0.214786
R4342 DVDD.n5336 DVDD.n433 0.214786
R4343 DVDD.n432 DVDD.n430 0.214786
R4344 DVDD.n431 DVDD.n423 0.214786
R4345 DVDD.n5343 DVDD.n422 0.214786
R4346 DVDD.n5344 DVDD.n421 0.214786
R4347 DVDD.n5345 DVDD.n420 0.214786
R4348 DVDD.n419 DVDD.n417 0.214786
R4349 DVDD.n5349 DVDD.n416 0.214786
R4350 DVDD.n5350 DVDD.n415 0.214786
R4351 DVDD.n5351 DVDD.n414 0.214786
R4352 DVDD.n413 DVDD.n411 0.214786
R4353 DVDD.n5355 DVDD.n410 0.214786
R4354 DVDD.n5356 DVDD.n409 0.214786
R4355 DVDD.n5357 DVDD.n408 0.214786
R4356 DVDD.n698 DVDD.n399 0.214786
R4357 DVDD.n5363 DVDD.n398 0.214786
R4358 DVDD.n5364 DVDD.n397 0.214786
R4359 DVDD.n5365 DVDD.n396 0.214786
R4360 DVDD.n395 DVDD.n393 0.214786
R4361 DVDD.n5369 DVDD.n392 0.214786
R4362 DVDD.n5370 DVDD.n391 0.214786
R4363 DVDD.n5371 DVDD.n390 0.214786
R4364 DVDD.n389 DVDD.n387 0.214786
R4365 DVDD.n5375 DVDD.n386 0.214786
R4366 DVDD.n5376 DVDD.n385 0.214786
R4367 DVDD.n5377 DVDD.n384 0.214786
R4368 DVDD.n383 DVDD.n376 0.214786
R4369 DVDD.n5383 DVDD.n375 0.214786
R4370 DVDD.n5384 DVDD.n374 0.214786
R4371 DVDD.n5385 DVDD.n373 0.214786
R4372 DVDD.n372 DVDD.n370 0.214786
R4373 DVDD.n5389 DVDD.n369 0.214786
R4374 DVDD.n5390 DVDD.n368 0.214786
R4375 DVDD.n5391 DVDD.n367 0.214786
R4376 DVDD.n366 DVDD.n364 0.214786
R4377 DVDD.n5395 DVDD.n363 0.214786
R4378 DVDD.n5396 DVDD.n362 0.214786
R4379 DVDD.n5397 DVDD.n361 0.214786
R4380 DVDD.n5401 DVDD.n357 0.214786
R4381 DVDD.n5403 DVDD.n356 0.214786
R4382 DVDD.n5404 DVDD.n355 0.214786
R4383 DVDD.n1164 DVDD.n354 0.214786
R4384 DVDD.n1166 DVDD.n1165 0.214786
R4385 DVDD.n1167 DVDD.n1163 0.214786
R4386 DVDD.n1162 DVDD.n1160 0.214786
R4387 DVDD.n1171 DVDD.n1159 0.214786
R4388 DVDD.n1172 DVDD.n1158 0.214786
R4389 DVDD.n1173 DVDD.n1157 0.214786
R4390 DVDD.n1156 DVDD.n1154 0.214786
R4391 DVDD.n1177 DVDD.n1153 0.214786
R4392 DVDD.n1178 DVDD.n1152 0.214786
R4393 DVDD.n1179 DVDD.n1151 0.214786
R4394 DVDD.n2046 DVDD.n2045 0.214786
R4395 DVDD.n2052 DVDD.n2051 0.214786
R4396 DVDD.n2043 DVDD.n2042 0.214786
R4397 DVDD.n2057 DVDD.n2056 0.214786
R4398 DVDD.n3086 DVDD.n3085 0.214786
R4399 DVDD.n2070 DVDD.n2028 0.214786
R4400 DVDD.n3081 DVDD.n2030 0.214786
R4401 DVDD.n3080 DVDD.n2031 0.214786
R4402 DVDD.n3079 DVDD.n2032 0.214786
R4403 DVDD.n2064 DVDD.n2033 0.214786
R4404 DVDD.n3075 DVDD.n2035 0.214786
R4405 DVDD.n3074 DVDD.n2036 0.214786
R4406 DVDD.n3073 DVDD.n2037 0.214786
R4407 DVDD.n3071 DVDD.n3070 0.214786
R4408 DVDD.n3039 DVDD.n1996 0.214786
R4409 DVDD.n3045 DVDD.n3044 0.214786
R4410 DVDD.n3041 DVDD.n3037 0.214786
R4411 DVDD.n3051 DVDD.n3050 0.214786
R4412 DVDD.n3038 DVDD.n3034 0.214786
R4413 DVDD.n3055 DVDD.n3033 0.214786
R4414 DVDD.n3057 DVDD.n3056 0.214786
R4415 DVDD.n3030 DVDD.n3028 0.214786
R4416 DVDD.n3062 DVDD.n3061 0.214786
R4417 DVDD.n3031 DVDD.n3029 0.214786
R4418 DVDD.n1928 DVDD.n1927 0.214786
R4419 DVDD.n1930 DVDD.n1929 0.214786
R4420 DVDD.n1931 DVDD.n1925 0.214786
R4421 DVDD.n3047 DVDD.n3037 0.214786
R4422 DVDD.n3046 DVDD.n3045 0.214786
R4423 DVDD.n3039 DVDD.n2002 0.214786
R4424 DVDD.n3071 DVDD.n2001 0.214786
R4425 DVDD.n3073 DVDD.n3072 0.214786
R4426 DVDD.n3074 DVDD.n2034 0.214786
R4427 DVDD.n3076 DVDD.n3075 0.214786
R4428 DVDD.n3077 DVDD.n2033 0.214786
R4429 DVDD.n3079 DVDD.n3078 0.214786
R4430 DVDD.n3080 DVDD.n2029 0.214786
R4431 DVDD.n3082 DVDD.n3081 0.214786
R4432 DVDD.n3083 DVDD.n2028 0.214786
R4433 DVDD.n3085 DVDD.n3084 0.214786
R4434 DVDD.n2056 DVDD.n2055 0.214786
R4435 DVDD.n2054 DVDD.n2043 0.214786
R4436 DVDD.n2053 DVDD.n2052 0.214786
R4437 DVDD.n3050 DVDD.n3049 0.214786
R4438 DVDD.n3048 DVDD.n3038 0.214786
R4439 DVDD.n3033 DVDD.n3032 0.214786
R4440 DVDD.n3058 DVDD.n3057 0.214786
R4441 DVDD.n3059 DVDD.n3030 0.214786
R4442 DVDD.n3061 DVDD.n3060 0.214786
R4443 DVDD.n3031 DVDD.n1902 0.214786
R4444 DVDD.n1927 DVDD.n1901 0.214786
R4445 DVDD.n1930 DVDD.n1926 0.214786
R4446 DVDD.n3585 DVDD.n3131 0.214786
R4447 DVDD.n3586 DVDD.n3130 0.214786
R4448 DVDD.n3129 DVDD.n1999 0.214786
R4449 DVDD.n3118 DVDD.n2000 0.214786
R4450 DVDD.n3598 DVDD.n3117 0.214786
R4451 DVDD.n3599 DVDD.n3116 0.214786
R4452 DVDD.n3115 DVDD.n3108 0.214786
R4453 DVDD.n3608 DVDD.n3107 0.214786
R4454 DVDD.n3609 DVDD.n3106 0.214786
R4455 DVDD.n3610 DVDD.n3105 0.214786
R4456 DVDD.n3104 DVDD.n3102 0.214786
R4457 DVDD.n3614 DVDD.n3101 0.214786
R4458 DVDD.n3615 DVDD.n3100 0.214786
R4459 DVDD.n3306 DVDD.n3305 0.214786
R4460 DVDD.n3304 DVDD.n3300 0.214786
R4461 DVDD.n3303 DVDD.n3302 0.214786
R4462 DVDD.n3145 DVDD.n3132 0.214786
R4463 DVDD.n3146 DVDD.n3144 0.214786
R4464 DVDD.n3574 DVDD.n3147 0.214786
R4465 DVDD.n3573 DVDD.n3148 0.214786
R4466 DVDD.n3563 DVDD.n3149 0.214786
R4467 DVDD.n3566 DVDD.n3564 0.214786
R4468 DVDD.n3565 DVDD.n1944 0.214786
R4469 DVDD.n1943 DVDD.n1942 0.214786
R4470 DVDD.n1906 DVDD.n1905 0.214786
R4471 DVDD.n3301 DVDD.n3274 0.214786
R4472 DVDD.n3302 DVDD.n3281 0.214786
R4473 DVDD.n3300 DVDD.n3295 0.214786
R4474 DVDD.n3307 DVDD.n3306 0.214786
R4475 DVDD.n3616 DVDD.n3615 0.214786
R4476 DVDD.n3614 DVDD.n3613 0.214786
R4477 DVDD.n3612 DVDD.n3102 0.214786
R4478 DVDD.n3611 DVDD.n3610 0.214786
R4479 DVDD.n3609 DVDD.n3103 0.214786
R4480 DVDD.n3608 DVDD.n3607 0.214786
R4481 DVDD.n3109 DVDD.n3108 0.214786
R4482 DVDD.n3600 DVDD.n3599 0.214786
R4483 DVDD.n3598 DVDD.n3597 0.214786
R4484 DVDD.n3119 DVDD.n3118 0.214786
R4485 DVDD.n3129 DVDD.n1992 0.214786
R4486 DVDD.n3587 DVDD.n3586 0.214786
R4487 DVDD.n3585 DVDD.n3584 0.214786
R4488 DVDD.n3133 DVDD.n3132 0.214786
R4489 DVDD.n3144 DVDD.n3142 0.214786
R4490 DVDD.n3575 DVDD.n3574 0.214786
R4491 DVDD.n3573 DVDD.n3572 0.214786
R4492 DVDD.n3159 DVDD.n3149 0.214786
R4493 DVDD.n3567 DVDD.n3566 0.214786
R4494 DVDD.n3565 DVDD.n3562 0.214786
R4495 DVDD.n1942 DVDD.n1941 0.214786
R4496 DVDD.n1940 DVDD.n1906 0.214786
R4497 DVDD.n1939 DVDD.n1938 0.214786
R4498 DVDD.n3250 DVDD.n3248 0.214786
R4499 DVDD.n3257 DVDD.n3256 0.214786
R4500 DVDD.n3251 DVDD.n3229 0.214786
R4501 DVDD.n3252 DVDD.n3230 0.214786
R4502 DVDD.n3219 DVDD.n3095 0.214786
R4503 DVDD.n3399 DVDD.n3220 0.214786
R4504 DVDD.n3401 DVDD.n3400 0.214786
R4505 DVDD.n3216 DVDD.n3215 0.214786
R4506 DVDD.n3406 DVDD.n3405 0.214786
R4507 DVDD.n3407 DVDD.n3214 0.214786
R4508 DVDD.n3421 DVDD.n3420 0.214786
R4509 DVDD.n3410 DVDD.n3212 0.214786
R4510 DVDD.n3425 DVDD.n3211 0.214786
R4511 DVDD.n3427 DVDD.n3426 0.214786
R4512 DVDD.n3203 DVDD.n1990 0.214786
R4513 DVDD.n3437 DVDD.n3204 0.214786
R4514 DVDD.n3448 DVDD.n3447 0.214786
R4515 DVDD.n3463 DVDD.n3462 0.214786
R4516 DVDD.n3201 DVDD.n3200 0.214786
R4517 DVDD.n3458 DVDD.n3452 0.214786
R4518 DVDD.n3457 DVDD.n3173 0.214786
R4519 DVDD.n3456 DVDD.n3183 0.214786
R4520 DVDD.n3454 DVDD.n3453 0.214786
R4521 DVDD.n1964 DVDD.n1948 0.214786
R4522 DVDD.n1963 DVDD.n1949 0.214786
R4523 DVDD.n1962 DVDD.n1950 0.214786
R4524 DVDD.n3199 DVDD.n3197 0.214786
R4525 DVDD.n3449 DVDD.n3448 0.214786
R4526 DVDD.n3204 DVDD.n3202 0.214786
R4527 DVDD.n3203 DVDD.n2003 0.214786
R4528 DVDD.n3426 DVDD.n2004 0.214786
R4529 DVDD.n3425 DVDD.n3424 0.214786
R4530 DVDD.n3423 DVDD.n3212 0.214786
R4531 DVDD.n3422 DVDD.n3421 0.214786
R4532 DVDD.n3214 DVDD.n3213 0.214786
R4533 DVDD.n3405 DVDD.n3404 0.214786
R4534 DVDD.n3403 DVDD.n3216 0.214786
R4535 DVDD.n3402 DVDD.n3401 0.214786
R4536 DVDD.n3220 DVDD.n3217 0.214786
R4537 DVDD.n3219 DVDD.n3218 0.214786
R4538 DVDD.n3253 DVDD.n3252 0.214786
R4539 DVDD.n3254 DVDD.n3251 0.214786
R4540 DVDD.n3256 DVDD.n3255 0.214786
R4541 DVDD.n3450 DVDD.n3199 0.214786
R4542 DVDD.n3462 DVDD.n3461 0.214786
R4543 DVDD.n3460 DVDD.n3201 0.214786
R4544 DVDD.n3459 DVDD.n3458 0.214786
R4545 DVDD.n3457 DVDD.n3451 0.214786
R4546 DVDD.n3456 DVDD.n3455 0.214786
R4547 DVDD.n3454 DVDD.n1966 0.214786
R4548 DVDD.n1965 DVDD.n1964 0.214786
R4549 DVDD.n1963 DVDD.n1947 0.214786
R4550 DVDD.n3671 DVDD.n1976 0.214786
R4551 DVDD.n3670 DVDD.n3669 0.214786
R4552 DVDD.n1978 DVDD.n1977 0.214786
R4553 DVDD.n3646 DVDD.n3645 0.214786
R4554 DVDD.n3644 DVDD.n2005 0.214786
R4555 DVDD.n3633 DVDD.n2006 0.214786
R4556 DVDD.n3635 DVDD.n3634 0.214786
R4557 DVDD.n3632 DVDD.n2017 0.214786
R4558 DVDD.n3631 DVDD.n3630 0.214786
R4559 DVDD.n2019 DVDD.n2018 0.214786
R4560 DVDD.n3623 DVDD.n3622 0.214786
R4561 DVDD.n3621 DVDD.n2021 0.214786
R4562 DVDD.n3620 DVDD.n3619 0.214786
R4563 DVDD.n1974 DVDD.n1973 0.214786
R4564 DVDD.n3678 DVDD.n3677 0.214786
R4565 DVDD.n3679 DVDD.n1972 0.214786
R4566 DVDD.n3681 DVDD.n3680 0.214786
R4567 DVDD.n1970 DVDD.n1969 0.214786
R4568 DVDD.n3686 DVDD.n3685 0.214786
R4569 DVDD.n3703 DVDD.n3702 0.214786
R4570 DVDD.n3688 DVDD.n3687 0.214786
R4571 DVDD.n3673 DVDD.n3672 0.214786
R4572 DVDD.n3619 DVDD.n3618 0.214786
R4573 DVDD.n2021 DVDD.n2020 0.214786
R4574 DVDD.n3624 DVDD.n3623 0.214786
R4575 DVDD.n3625 DVDD.n2019 0.214786
R4576 DVDD.n3630 DVDD.n3629 0.214786
R4577 DVDD.n3626 DVDD.n2017 0.214786
R4578 DVDD.n3636 DVDD.n3635 0.214786
R4579 DVDD.n3637 DVDD.n2006 0.214786
R4580 DVDD.n3644 DVDD.n3643 0.214786
R4581 DVDD.n3645 DVDD.n1983 0.214786
R4582 DVDD.n3653 DVDD.n1978 0.214786
R4583 DVDD.n3669 DVDD.n3668 0.214786
R4584 DVDD.n1980 DVDD.n1976 0.214786
R4585 DVDD.n3675 DVDD.n1974 0.214786
R4586 DVDD.n3677 DVDD.n3676 0.214786
R4587 DVDD.n1972 DVDD.n1971 0.214786
R4588 DVDD.n3682 DVDD.n3681 0.214786
R4589 DVDD.n3683 DVDD.n1970 0.214786
R4590 DVDD.n3685 DVDD.n3684 0.214786
R4591 DVDD.n3702 DVDD.n3701 0.214786
R4592 DVDD.n3700 DVDD.n3688 0.214786
R4593 DVDD.n3699 DVDD.n3698 0.214786
R4594 DVDD.n3674 DVDD.n3673 0.214786
R4595 DVDD.n4196 DVDD.n4195 0.214786
R4596 DVDD.n4193 DVDD.n4192 0.214786
R4597 DVDD.n4191 DVDD.n4186 0.214786
R4598 DVDD.n4207 DVDD.n4185 0.214786
R4599 DVDD.n4208 DVDD.n4184 0.214786
R4600 DVDD.n4209 DVDD.n4183 0.214786
R4601 DVDD.n4182 DVDD.n4180 0.214786
R4602 DVDD.n4213 DVDD.n4179 0.214786
R4603 DVDD.n4214 DVDD.n4178 0.214786
R4604 DVDD.n4215 DVDD.n4177 0.214786
R4605 DVDD.n4172 DVDD.n4171 0.214786
R4606 DVDD.n4220 DVDD.n4219 0.214786
R4607 DVDD.n4170 DVDD.n4169 0.214786
R4608 DVDD.n1768 DVDD.n1767 0.214786
R4609 DVDD.n4165 DVDD.n4164 0.214786
R4610 DVDD.n4163 DVDD.n1770 0.214786
R4611 DVDD.n4162 DVDD.n4161 0.214786
R4612 DVDD.n1772 DVDD.n1771 0.214786
R4613 DVDD.n4155 DVDD.n4154 0.214786
R4614 DVDD.n4153 DVDD.n1774 0.214786
R4615 DVDD.n4152 DVDD.n4151 0.214786
R4616 DVDD.n3732 DVDD.n3731 0.214786
R4617 DVDD.n1855 DVDD.n1854 0.214786
R4618 DVDD.n3782 DVDD.n3781 0.214786
R4619 DVDD.n3783 DVDD.n1853 0.214786
R4620 DVDD.n3785 DVDD.n3784 0.214786
R4621 DVDD.n1851 DVDD.n1850 0.214786
R4622 DVDD.n3790 DVDD.n3789 0.214786
R4623 DVDD.n3791 DVDD.n1849 0.214786
R4624 DVDD.n3793 DVDD.n3792 0.214786
R4625 DVDD.n1847 DVDD.n1846 0.214786
R4626 DVDD.n3799 DVDD.n3798 0.214786
R4627 DVDD.n3800 DVDD.n1845 0.214786
R4628 DVDD.n3802 DVDD.n3801 0.214786
R4629 DVDD.n3803 DVDD.n1687 0.214786
R4630 DVDD.n4257 DVDD.n4256 0.214786
R4631 DVDD.n1689 DVDD.n1688 0.214786
R4632 DVDD.n4252 DVDD.n1692 0.214786
R4633 DVDD.n4251 DVDD.n1693 0.214786
R4634 DVDD.n1696 DVDD.n1694 0.214786
R4635 DVDD.n4247 DVDD.n1697 0.214786
R4636 DVDD.n4246 DVDD.n1698 0.214786
R4637 DVDD.n1701 DVDD.n1699 0.214786
R4638 DVDD.n4242 DVDD.n1702 0.214786
R4639 DVDD.n4241 DVDD.n1703 0.214786
R4640 DVDD.n4240 DVDD.n1704 0.214786
R4641 DVDD.n3936 DVDD.n1705 0.214786
R4642 DVDD.n3937 DVDD.n3935 0.214786
R4643 DVDD.n3956 DVDD.n3938 0.214786
R4644 DVDD.n3955 DVDD.n3939 0.214786
R4645 DVDD.n3954 DVDD.n3940 0.214786
R4646 DVDD.n3943 DVDD.n3941 0.214786
R4647 DVDD.n3949 DVDD.n3944 0.214786
R4648 DVDD.n3948 DVDD.n3945 0.214786
R4649 DVDD.n3947 DVDD.n3946 0.214786
R4650 DVDD.n3926 DVDD.n3925 0.214786
R4651 DVDD.n3970 DVDD.n3969 0.214786
R4652 DVDD.n3971 DVDD.n3924 0.214786
R4653 DVDD.n3973 DVDD.n3972 0.214786
R4654 DVDD.n3978 DVDD.n3977 0.214786
R4655 DVDD.n3979 DVDD.n1816 0.214786
R4656 DVDD.n3981 DVDD.n3980 0.214786
R4657 DVDD.n1814 DVDD.n1813 0.214786
R4658 DVDD.n3986 DVDD.n3985 0.214786
R4659 DVDD.n3987 DVDD.n1812 0.214786
R4660 DVDD.n3989 DVDD.n3988 0.214786
R4661 DVDD.n1810 DVDD.n1809 0.214786
R4662 DVDD.n3998 DVDD.n3997 0.214786
R4663 DVDD.n3999 DVDD.n1808 0.214786
R4664 DVDD.n4001 DVDD.n4000 0.214786
R4665 DVDD.n1806 DVDD.n1805 0.214786
R4666 DVDD.n4006 DVDD.n4005 0.214786
R4667 DVDD.n4007 DVDD.n1804 0.214786
R4668 DVDD.n4009 DVDD.n4008 0.214786
R4669 DVDD.n1802 DVDD.n1801 0.214786
R4670 DVDD.n4018 DVDD.n4017 0.214786
R4671 DVDD.n4019 DVDD.n1800 0.214786
R4672 DVDD.n4021 DVDD.n4020 0.214786
R4673 DVDD.n1798 DVDD.n1797 0.214786
R4674 DVDD.n4027 DVDD.n4026 0.214786
R4675 DVDD.n4028 DVDD.n1796 0.214786
R4676 DVDD.n4030 DVDD.n4029 0.214786
R4677 DVDD.n4031 DVDD.n1789 0.214786
R4678 DVDD.n4103 DVDD.n1788 0.214786
R4679 DVDD.n4117 DVDD.n4104 0.214786
R4680 DVDD.n4116 DVDD.n4105 0.214786
R4681 DVDD.n4115 DVDD.n4106 0.214786
R4682 DVDD.n4108 DVDD.n4107 0.214786
R4683 DVDD.n4110 DVDD.n4109 0.214786
R4684 DVDD.n1783 DVDD.n1782 0.214786
R4685 DVDD.n4130 DVDD.n4129 0.214786
R4686 DVDD.n4131 DVDD.n1781 0.214786
R4687 DVDD.n4133 DVDD.n4132 0.214786
R4688 DVDD.n1779 DVDD.n1778 0.214786
R4689 DVDD.n4142 DVDD.n4141 0.214786
R4690 DVDD.n4143 DVDD.n1777 0.214786
R4691 DVDD.n4145 DVDD.n4144 0.214786
R4692 DVDD.n1776 DVDD.n1775 0.214786
R4693 DVDD.n4151 DVDD.n4150 0.214786
R4694 DVDD.n1774 DVDD.n1773 0.214786
R4695 DVDD.n4156 DVDD.n4155 0.214786
R4696 DVDD.n4158 DVDD.n1772 0.214786
R4697 DVDD.n4161 DVDD.n4160 0.214786
R4698 DVDD.n4159 DVDD.n1770 0.214786
R4699 DVDD.n4166 DVDD.n4165 0.214786
R4700 DVDD.n4167 DVDD.n1768 0.214786
R4701 DVDD.n4169 DVDD.n4168 0.214786
R4702 DVDD.n4219 DVDD.n4218 0.214786
R4703 DVDD.n4217 DVDD.n4172 0.214786
R4704 DVDD.n4216 DVDD.n4215 0.214786
R4705 DVDD.n4214 DVDD.n4176 0.214786
R4706 DVDD.n4213 DVDD.n4212 0.214786
R4707 DVDD.n4211 DVDD.n4180 0.214786
R4708 DVDD.n4210 DVDD.n4209 0.214786
R4709 DVDD.n4208 DVDD.n4181 0.214786
R4710 DVDD.n4207 DVDD.n4206 0.214786
R4711 DVDD.n4205 DVDD.n4186 0.214786
R4712 DVDD.n4193 DVDD.n4187 0.214786
R4713 DVDD.n4195 DVDD.n4194 0.214786
R4714 DVDD.n4190 DVDD.n4189 0.214786
R4715 DVDD.n3734 DVDD.n3733 0.214786
R4716 DVDD.n3732 DVDD.n1856 0.214786
R4717 DVDD.n3778 DVDD.n1855 0.214786
R4718 DVDD.n3781 DVDD.n3780 0.214786
R4719 DVDD.n3779 DVDD.n1853 0.214786
R4720 DVDD.n3786 DVDD.n3785 0.214786
R4721 DVDD.n3787 DVDD.n1851 0.214786
R4722 DVDD.n3789 DVDD.n3788 0.214786
R4723 DVDD.n1849 DVDD.n1848 0.214786
R4724 DVDD.n3794 DVDD.n3793 0.214786
R4725 DVDD.n3795 DVDD.n1847 0.214786
R4726 DVDD.n3798 DVDD.n3797 0.214786
R4727 DVDD.n3796 DVDD.n1845 0.214786
R4728 DVDD.n3802 DVDD.n1844 0.214786
R4729 DVDD.n3804 DVDD.n3803 0.214786
R4730 DVDD.n4256 DVDD.n4255 0.214786
R4731 DVDD.n4254 DVDD.n1689 0.214786
R4732 DVDD.n4253 DVDD.n4252 0.214786
R4733 DVDD.n4251 DVDD.n4250 0.214786
R4734 DVDD.n4249 DVDD.n1694 0.214786
R4735 DVDD.n4248 DVDD.n4247 0.214786
R4736 DVDD.n4246 DVDD.n4245 0.214786
R4737 DVDD.n4244 DVDD.n1699 0.214786
R4738 DVDD.n4243 DVDD.n4242 0.214786
R4739 DVDD.n4241 DVDD.n1700 0.214786
R4740 DVDD.n4240 DVDD.n4239 0.214786
R4741 DVDD.n1707 DVDD.n1705 0.214786
R4742 DVDD.n3935 DVDD.n3933 0.214786
R4743 DVDD.n3957 DVDD.n3956 0.214786
R4744 DVDD.n3955 DVDD.n3934 0.214786
R4745 DVDD.n3954 DVDD.n3953 0.214786
R4746 DVDD.n3951 DVDD.n3941 0.214786
R4747 DVDD.n3950 DVDD.n3949 0.214786
R4748 DVDD.n3948 DVDD.n3942 0.214786
R4749 DVDD.n3947 DVDD.n3927 0.214786
R4750 DVDD.n3966 DVDD.n3926 0.214786
R4751 DVDD.n3969 DVDD.n3968 0.214786
R4752 DVDD.n3967 DVDD.n3924 0.214786
R4753 DVDD.n3974 DVDD.n3973 0.214786
R4754 DVDD.n3977 DVDD.n3976 0.214786
R4755 DVDD.n1816 DVDD.n1815 0.214786
R4756 DVDD.n3982 DVDD.n3981 0.214786
R4757 DVDD.n3983 DVDD.n1814 0.214786
R4758 DVDD.n3985 DVDD.n3984 0.214786
R4759 DVDD.n1812 DVDD.n1811 0.214786
R4760 DVDD.n3990 DVDD.n3989 0.214786
R4761 DVDD.n3991 DVDD.n1810 0.214786
R4762 DVDD.n3997 DVDD.n3996 0.214786
R4763 DVDD.n1808 DVDD.n1807 0.214786
R4764 DVDD.n4002 DVDD.n4001 0.214786
R4765 DVDD.n4003 DVDD.n1806 0.214786
R4766 DVDD.n4005 DVDD.n4004 0.214786
R4767 DVDD.n1804 DVDD.n1803 0.214786
R4768 DVDD.n4010 DVDD.n4009 0.214786
R4769 DVDD.n4015 DVDD.n1802 0.214786
R4770 DVDD.n4017 DVDD.n4016 0.214786
R4771 DVDD.n1800 DVDD.n1799 0.214786
R4772 DVDD.n4022 DVDD.n4021 0.214786
R4773 DVDD.n4023 DVDD.n1798 0.214786
R4774 DVDD.n4026 DVDD.n4025 0.214786
R4775 DVDD.n4024 DVDD.n1796 0.214786
R4776 DVDD.n4030 DVDD.n1795 0.214786
R4777 DVDD.n4032 DVDD.n4031 0.214786
R4778 DVDD.n1788 DVDD.n1786 0.214786
R4779 DVDD.n4118 DVDD.n4117 0.214786
R4780 DVDD.n4116 DVDD.n1787 0.214786
R4781 DVDD.n4115 DVDD.n4114 0.214786
R4782 DVDD.n4112 DVDD.n4107 0.214786
R4783 DVDD.n4111 DVDD.n4110 0.214786
R4784 DVDD.n1784 DVDD.n1783 0.214786
R4785 DVDD.n4129 DVDD.n4128 0.214786
R4786 DVDD.n1781 DVDD.n1780 0.214786
R4787 DVDD.n4134 DVDD.n4133 0.214786
R4788 DVDD.n4135 DVDD.n1779 0.214786
R4789 DVDD.n4141 DVDD.n4140 0.214786
R4790 DVDD.n4139 DVDD.n1777 0.214786
R4791 DVDD.n4146 DVDD.n4145 0.214786
R4792 DVDD.n4149 DVDD.n1776 0.214786
R4793 DVDD.n1181 DVDD.n1180 0.214786
R4794 DVDD.n1179 DVDD.n1121 0.214786
R4795 DVDD.n1178 DVDD.n1131 0.214786
R4796 DVDD.n1177 DVDD.n1176 0.214786
R4797 DVDD.n1175 DVDD.n1154 0.214786
R4798 DVDD.n1174 DVDD.n1173 0.214786
R4799 DVDD.n1172 DVDD.n1155 0.214786
R4800 DVDD.n1171 DVDD.n1170 0.214786
R4801 DVDD.n1169 DVDD.n1160 0.214786
R4802 DVDD.n1168 DVDD.n1167 0.214786
R4803 DVDD.n1166 DVDD.n1161 0.214786
R4804 DVDD.n354 DVDD.n328 0.214786
R4805 DVDD.n5405 DVDD.n5404 0.214786
R4806 DVDD.n5403 DVDD.n5402 0.214786
R4807 DVDD.n5401 DVDD.n5400 0.214786
R4808 DVDD.n5398 DVDD.n5397 0.214786
R4809 DVDD.n5396 DVDD.n360 0.214786
R4810 DVDD.n5395 DVDD.n5394 0.214786
R4811 DVDD.n5393 DVDD.n364 0.214786
R4812 DVDD.n5392 DVDD.n5391 0.214786
R4813 DVDD.n5390 DVDD.n365 0.214786
R4814 DVDD.n5389 DVDD.n5388 0.214786
R4815 DVDD.n5387 DVDD.n370 0.214786
R4816 DVDD.n5386 DVDD.n5385 0.214786
R4817 DVDD.n5384 DVDD.n371 0.214786
R4818 DVDD.n5383 DVDD.n5382 0.214786
R4819 DVDD.n379 DVDD.n376 0.214786
R4820 DVDD.n5378 DVDD.n5377 0.214786
R4821 DVDD.n5376 DVDD.n382 0.214786
R4822 DVDD.n5375 DVDD.n5374 0.214786
R4823 DVDD.n5373 DVDD.n387 0.214786
R4824 DVDD.n5372 DVDD.n5371 0.214786
R4825 DVDD.n5370 DVDD.n388 0.214786
R4826 DVDD.n5369 DVDD.n5368 0.214786
R4827 DVDD.n5367 DVDD.n393 0.214786
R4828 DVDD.n5366 DVDD.n5365 0.214786
R4829 DVDD.n5364 DVDD.n394 0.214786
R4830 DVDD.n5363 DVDD.n5362 0.214786
R4831 DVDD.n402 DVDD.n399 0.214786
R4832 DVDD.n5358 DVDD.n5357 0.214786
R4833 DVDD.n5356 DVDD.n406 0.214786
R4834 DVDD.n5355 DVDD.n5354 0.214786
R4835 DVDD.n5353 DVDD.n411 0.214786
R4836 DVDD.n5352 DVDD.n5351 0.214786
R4837 DVDD.n5350 DVDD.n412 0.214786
R4838 DVDD.n5349 DVDD.n5348 0.214786
R4839 DVDD.n5347 DVDD.n417 0.214786
R4840 DVDD.n5346 DVDD.n5345 0.214786
R4841 DVDD.n5344 DVDD.n418 0.214786
R4842 DVDD.n5343 DVDD.n5342 0.214786
R4843 DVDD.n5341 DVDD.n423 0.214786
R4844 DVDD.n430 DVDD.n426 0.214786
R4845 DVDD.n5337 DVDD.n5336 0.214786
R4846 DVDD.n5335 DVDD.n429 0.214786
R4847 DVDD.n5334 DVDD.n5333 0.214786
R4848 DVDD.n5332 DVDD.n436 0.214786
R4849 DVDD.n5331 DVDD.n5330 0.214786
R4850 DVDD.n5329 DVDD.n437 0.214786
R4851 DVDD.n5328 DVDD.n5327 0.214786
R4852 DVDD.n5326 DVDD.n442 0.214786
R4853 DVDD.n5325 DVDD.n5324 0.214786
R4854 DVDD.n5323 DVDD.n443 0.214786
R4855 DVDD.n5322 DVDD.n5321 0.214786
R4856 DVDD.n5106 DVDD.n5104 0.214786
R4857 DVDD.n5133 DVDD.n5132 0.214786
R4858 DVDD.n5131 DVDD.n5105 0.214786
R4859 DVDD.n5130 DVDD.n5129 0.214786
R4860 DVDD.n5128 DVDD.n5111 0.214786
R4861 DVDD.n5127 DVDD.n5126 0.214786
R4862 DVDD.n5125 DVDD.n5112 0.214786
R4863 DVDD.n5124 DVDD.n5123 0.214786
R4864 DVDD.n5122 DVDD.n5117 0.214786
R4865 DVDD.n5121 DVDD.n5120 0.214786
R4866 DVDD.n134 DVDD.n133 0.214786
R4867 DVDD.n5851 DVDD.n5850 0.214786
R4868 DVDD.n137 DVDD.n131 0.214786
R4869 DVDD.n5856 DVDD.n5855 0.214786
R4870 DVDD.n5857 DVDD.n129 0.214786
R4871 DVDD.n5859 DVDD.n5858 0.214786
R4872 DVDD.n127 DVDD.n126 0.214786
R4873 DVDD.n5864 DVDD.n5863 0.214786
R4874 DVDD.n5865 DVDD.n125 0.214786
R4875 DVDD.n5867 DVDD.n5866 0.214786
R4876 DVDD.n123 DVDD.n122 0.214786
R4877 DVDD.n5872 DVDD.n5871 0.214786
R4878 DVDD.n5873 DVDD.n121 0.214786
R4879 DVDD.n5875 DVDD.n5874 0.214786
R4880 DVDD.n5879 DVDD.n80 0.214786
R4881 DVDD.n5880 DVDD.n82 0.214786
R4882 DVDD.n5882 DVDD.n5881 0.214786
R4883 DVDD.n117 DVDD.n116 0.214786
R4884 DVDD.n5907 DVDD.n5906 0.214786
R4885 DVDD.n5905 DVDD.n115 0.214786
R4886 DVDD.n5904 DVDD.n5903 0.214786
R4887 DVDD.n5902 DVDD.n5888 0.214786
R4888 DVDD.n5901 DVDD.n5900 0.214786
R4889 DVDD.n5899 DVDD.n5889 0.214786
R4890 DVDD.n5898 DVDD.n5897 0.214786
R4891 DVDD.n4410 DVDD.n4409 0.214786
R4892 DVDD.n1108 DVDD.n1107 0.214786
R4893 DVDD.n4416 DVDD.n4415 0.214786
R4894 DVDD.n1105 DVDD.n1104 0.214786
R4895 DVDD.n4421 DVDD.n4420 0.214786
R4896 DVDD.n4422 DVDD.n1103 0.214786
R4897 DVDD.n4424 DVDD.n4423 0.214786
R4898 DVDD.n1101 DVDD.n1100 0.214786
R4899 DVDD.n4429 DVDD.n4428 0.214786
R4900 DVDD.n4430 DVDD.n1099 0.214786
R4901 DVDD.n4432 DVDD.n4431 0.214786
R4902 DVDD.n1097 DVDD.n273 0.214786
R4903 DVDD.n4436 DVDD.n284 0.214786
R4904 DVDD.n4437 DVDD.n297 0.214786
R4905 DVDD.n4438 DVDD.n307 0.214786
R4906 DVDD.n4443 DVDD.n4442 0.214786
R4907 DVDD.n4445 DVDD.n4444 0.214786
R4908 DVDD.n1093 DVDD.n1092 0.214786
R4909 DVDD.n4450 DVDD.n4449 0.214786
R4910 DVDD.n4451 DVDD.n1091 0.214786
R4911 DVDD.n4453 DVDD.n4452 0.214786
R4912 DVDD.n1089 DVDD.n1088 0.214786
R4913 DVDD.n4458 DVDD.n4457 0.214786
R4914 DVDD.n4459 DVDD.n1087 0.214786
R4915 DVDD.n4461 DVDD.n4460 0.214786
R4916 DVDD.n1085 DVDD.n1075 0.214786
R4917 DVDD.n4497 DVDD.n4496 0.214786
R4918 DVDD.n4495 DVDD.n4494 0.214786
R4919 DVDD.n4493 DVDD.n4466 0.214786
R4920 DVDD.n4492 DVDD.n4491 0.214786
R4921 DVDD.n4490 DVDD.n4467 0.214786
R4922 DVDD.n4489 DVDD.n4488 0.214786
R4923 DVDD.n4487 DVDD.n4472 0.214786
R4924 DVDD.n4486 DVDD.n4485 0.214786
R4925 DVDD.n4484 DVDD.n4473 0.214786
R4926 DVDD.n4483 DVDD.n4482 0.214786
R4927 DVDD.n4481 DVDD.n4479 0.214786
R4928 DVDD.n4480 DVDD.n701 0.214786
R4929 DVDD.n4881 DVDD.n4880 0.214786
R4930 DVDD.n4886 DVDD.n4885 0.214786
R4931 DVDD.n4887 DVDD.n694 0.214786
R4932 DVDD.n4889 DVDD.n4888 0.214786
R4933 DVDD.n692 DVDD.n691 0.214786
R4934 DVDD.n4894 DVDD.n4893 0.214786
R4935 DVDD.n4895 DVDD.n690 0.214786
R4936 DVDD.n4897 DVDD.n4896 0.214786
R4937 DVDD.n688 DVDD.n687 0.214786
R4938 DVDD.n4902 DVDD.n4901 0.214786
R4939 DVDD.n4903 DVDD.n686 0.214786
R4940 DVDD.n4905 DVDD.n4904 0.214786
R4941 DVDD.n684 DVDD.n674 0.214786
R4942 DVDD.n4938 DVDD.n4937 0.214786
R4943 DVDD.n4936 DVDD.n4935 0.214786
R4944 DVDD.n4934 DVDD.n4910 0.214786
R4945 DVDD.n4933 DVDD.n4932 0.214786
R4946 DVDD.n4931 DVDD.n4911 0.214786
R4947 DVDD.n4930 DVDD.n4929 0.214786
R4948 DVDD.n4928 DVDD.n4916 0.214786
R4949 DVDD.n4927 DVDD.n4926 0.214786
R4950 DVDD.n4925 DVDD.n4917 0.214786
R4951 DVDD.n4924 DVDD.n4923 0.214786
R4952 DVDD.n4922 DVDD.n480 0.214786
R4953 DVDD.n5247 DVDD.n451 0.214786
R4954 DVDD.n476 DVDD.n462 0.214786
R4955 DVDD.n5315 DVDD.n5314 0.214786
R4956 DVDD.n5313 DVDD.n475 0.214786
R4957 DVDD.n5312 DVDD.n5311 0.214786
R4958 DVDD.n5310 DVDD.n5254 0.214786
R4959 DVDD.n5309 DVDD.n5308 0.214786
R4960 DVDD.n5307 DVDD.n5255 0.214786
R4961 DVDD.n5306 DVDD.n5305 0.214786
R4962 DVDD.n5304 DVDD.n5260 0.214786
R4963 DVDD.n5303 DVDD.n5302 0.214786
R4964 DVDD.n5301 DVDD.n5261 0.214786
R4965 DVDD.n5300 DVDD.n5299 0.214786
R4966 DVDD.n5298 DVDD.n144 0.214786
R4967 DVDD.n5297 DVDD.n155 0.214786
R4968 DVDD.n5296 DVDD.n5295 0.214786
R4969 DVDD.n5294 DVDD.n5269 0.214786
R4970 DVDD.n5293 DVDD.n5292 0.214786
R4971 DVDD.n5291 DVDD.n5270 0.214786
R4972 DVDD.n5290 DVDD.n5289 0.214786
R4973 DVDD.n5288 DVDD.n5275 0.214786
R4974 DVDD.n5287 DVDD.n5286 0.214786
R4975 DVDD.n5285 DVDD.n5276 0.214786
R4976 DVDD.n5284 DVDD.n5283 0.214786
R4977 DVDD.n5282 DVDD.n42 0.214786
R4978 DVDD.n5936 DVDD.n5935 0.214786
R4979 DVDD.n5934 DVDD.n5933 0.214786
R4980 DVDD.n58 DVDD.n47 0.214786
R4981 DVDD.n5576 DVDD.n5564 0.214786
R4982 DVDD.n5601 DVDD.n5600 0.214786
R4983 DVDD.n5599 DVDD.n5575 0.214786
R4984 DVDD.n5598 DVDD.n5597 0.214786
R4985 DVDD.n5596 DVDD.n5582 0.214786
R4986 DVDD.n5595 DVDD.n5594 0.214786
R4987 DVDD.n5593 DVDD.n5583 0.214786
R4988 DVDD.n5592 DVDD.n5591 0.214786
R4989 DVDD.n4373 DVDD.n4372 0.214786
R4990 DVDD.n4371 DVDD.n1596 0.214786
R4991 DVDD.n4370 DVDD.n1607 0.214786
R4992 DVDD.n4369 DVDD.n4368 0.214786
R4993 DVDD.n4367 DVDD.n4349 0.214786
R4994 DVDD.n4366 DVDD.n4365 0.214786
R4995 DVDD.n4364 DVDD.n4350 0.214786
R4996 DVDD.n4363 DVDD.n4362 0.214786
R4997 DVDD.n4361 DVDD.n4355 0.214786
R4998 DVDD.n4360 DVDD.n4359 0.214786
R4999 DVDD.n985 DVDD.n975 0.214786
R5000 DVDD.n4643 DVDD.n4642 0.214786
R5001 DVDD.n4641 DVDD.n4640 0.214786
R5002 DVDD.n4639 DVDD.n4638 0.214786
R5003 DVDD.n4637 DVDD.n4636 0.214786
R5004 DVDD.n4634 DVDD.n4633 0.214786
R5005 DVDD.n4632 DVDD.n992 0.214786
R5006 DVDD.n4631 DVDD.n4630 0.214786
R5007 DVDD.n4629 DVDD.n993 0.214786
R5008 DVDD.n4628 DVDD.n4627 0.214786
R5009 DVDD.n4626 DVDD.n998 0.214786
R5010 DVDD.n4625 DVDD.n4624 0.214786
R5011 DVDD.n4623 DVDD.n999 0.214786
R5012 DVDD.n4622 DVDD.n4621 0.214786
R5013 DVDD.n4620 DVDD.n1004 0.214786
R5014 DVDD.n4619 DVDD.n4618 0.214786
R5015 DVDD.n4617 DVDD.n4616 0.214786
R5016 DVDD.n1046 DVDD.n1009 0.214786
R5017 DVDD.n1045 DVDD.n1044 0.214786
R5018 DVDD.n1043 DVDD.n1020 0.214786
R5019 DVDD.n1042 DVDD.n1041 0.214786
R5020 DVDD.n1040 DVDD.n1025 0.214786
R5021 DVDD.n1039 DVDD.n1038 0.214786
R5022 DVDD.n1037 DVDD.n1026 0.214786
R5023 DVDD.n1036 DVDD.n1035 0.214786
R5024 DVDD.n1034 DVDD.n1033 0.214786
R5025 DVDD.n729 DVDD.n728 0.214786
R5026 DVDD.n4874 DVDD.n4873 0.214786
R5027 DVDD.n4872 DVDD.n704 0.214786
R5028 DVDD.n4870 DVDD.n715 0.214786
R5029 DVDD.n4869 DVDD.n4868 0.214786
R5030 DVDD.n4867 DVDD.n4805 0.214786
R5031 DVDD.n4866 DVDD.n4865 0.214786
R5032 DVDD.n4864 DVDD.n4806 0.214786
R5033 DVDD.n4863 DVDD.n4862 0.214786
R5034 DVDD.n4861 DVDD.n4811 0.214786
R5035 DVDD.n4860 DVDD.n4859 0.214786
R5036 DVDD.n4858 DVDD.n4812 0.214786
R5037 DVDD.n4857 DVDD.n4856 0.214786
R5038 DVDD.n4855 DVDD.n4854 0.214786
R5039 DVDD.n4853 DVDD.n605 0.214786
R5040 DVDD.n4852 DVDD.n616 0.214786
R5041 DVDD.n4851 DVDD.n4850 0.214786
R5042 DVDD.n4849 DVDD.n4821 0.214786
R5043 DVDD.n4848 DVDD.n4847 0.214786
R5044 DVDD.n4846 DVDD.n4822 0.214786
R5045 DVDD.n4845 DVDD.n4844 0.214786
R5046 DVDD.n4843 DVDD.n4827 0.214786
R5047 DVDD.n4842 DVDD.n4841 0.214786
R5048 DVDD.n4840 DVDD.n4828 0.214786
R5049 DVDD.n4839 DVDD.n4838 0.214786
R5050 DVDD.n4837 DVDD.n4835 0.214786
R5051 DVDD.n4836 DVDD.n482 0.214786
R5052 DVDD.n5244 DVDD.n5243 0.214786
R5053 DVDD.n555 DVDD.n484 0.214786
R5054 DVDD.n554 DVDD.n553 0.214786
R5055 DVDD.n552 DVDD.n496 0.214786
R5056 DVDD.n551 DVDD.n550 0.214786
R5057 DVDD.n549 DVDD.n501 0.214786
R5058 DVDD.n548 DVDD.n547 0.214786
R5059 DVDD.n546 DVDD.n502 0.214786
R5060 DVDD.n545 DVDD.n544 0.214786
R5061 DVDD.n543 DVDD.n507 0.214786
R5062 DVDD.n542 DVDD.n541 0.214786
R5063 DVDD.n540 DVDD.n170 0.214786
R5064 DVDD.n539 DVDD.n180 0.214786
R5065 DVDD.n538 DVDD.n537 0.214786
R5066 DVDD.n536 DVDD.n513 0.214786
R5067 DVDD.n535 DVDD.n534 0.214786
R5068 DVDD.n533 DVDD.n514 0.214786
R5069 DVDD.n532 DVDD.n531 0.214786
R5070 DVDD.n530 DVDD.n519 0.214786
R5071 DVDD.n529 DVDD.n528 0.214786
R5072 DVDD.n527 DVDD.n520 0.214786
R5073 DVDD.n526 DVDD.n525 0.214786
R5074 DVDD.n39 DVDD.n37 0.214786
R5075 DVDD.n5940 DVDD.n5939 0.214786
R5076 DVDD.n33 DVDD.n32 0.214786
R5077 DVDD.n5951 DVDD.n5950 0.214786
R5078 DVDD.n5949 DVDD.n5948 0.214786
R5079 DVDD.n5947 DVDD.n7 0.214786
R5080 DVDD.n5955 DVDD.n6 0.214786
R5081 DVDD.n5957 DVDD.n5956 0.214786
R5082 DVDD.n4 DVDD.n3 0.214786
R5083 DVDD.n5963 DVDD.n5962 0.214786
R5084 DVDD.n5964 DVDD.n2 0.214786
R5085 DVDD.n5966 DVDD.n5965 0.214786
R5086 DVDD.n5967 DVDD.n0 0.214786
R5087 DVDD.n5689 DVDD.n5684 0.214786
R5088 DVDD.n5691 DVDD.n5690 0.214786
R5089 DVDD.n5692 DVDD.n5679 0.214786
R5090 DVDD.n5694 DVDD.n5693 0.214786
R5091 DVDD.n5695 DVDD.n5678 0.214786
R5092 DVDD.n5697 DVDD.n5696 0.214786
R5093 DVDD.n5698 DVDD.n234 0.214786
R5094 DVDD.n5699 DVDD.n227 0.214786
R5095 DVDD.n5701 DVDD.n5700 0.214786
R5096 DVDD.n220 DVDD.n217 0.214786
R5097 DVDD.n5709 DVDD.n5708 0.214786
R5098 DVDD.n5712 DVDD.n5711 0.214786
R5099 DVDD.n5713 DVDD.n211 0.214786
R5100 DVDD.n5715 DVDD.n5714 0.214786
R5101 DVDD.n5716 DVDD.n210 0.214786
R5102 DVDD.n5718 DVDD.n5717 0.214786
R5103 DVDD.n5719 DVDD.n205 0.214786
R5104 DVDD.n5721 DVDD.n5720 0.214786
R5105 DVDD.n5722 DVDD.n204 0.214786
R5106 DVDD.n5724 DVDD.n5723 0.214786
R5107 DVDD.n5725 DVDD.n199 0.214786
R5108 DVDD.n5727 DVDD.n5726 0.214786
R5109 DVDD.n200 DVDD.n197 0.214786
R5110 DVDD.n5068 DVDD.n5067 0.214786
R5111 DVDD.n5069 DVDD.n5063 0.214786
R5112 DVDD.n5071 DVDD.n5070 0.214786
R5113 DVDD.n5072 DVDD.n5058 0.214786
R5114 DVDD.n5074 DVDD.n5073 0.214786
R5115 DVDD.n5075 DVDD.n5057 0.214786
R5116 DVDD.n5077 DVDD.n5076 0.214786
R5117 DVDD.n5078 DVDD.n5052 0.214786
R5118 DVDD.n5080 DVDD.n5079 0.214786
R5119 DVDD.n5081 DVDD.n5051 0.214786
R5120 DVDD.n5083 DVDD.n5082 0.214786
R5121 DVDD.n5085 DVDD.n5084 0.214786
R5122 DVDD.n5046 DVDD.n5045 0.214786
R5123 DVDD.n5044 DVDD.n575 0.214786
R5124 DVDD.n5043 DVDD.n5042 0.214786
R5125 DVDD.n577 DVDD.n576 0.214786
R5126 DVDD.n5038 DVDD.n5037 0.214786
R5127 DVDD.n5036 DVDD.n579 0.214786
R5128 DVDD.n5035 DVDD.n5034 0.214786
R5129 DVDD.n581 DVDD.n580 0.214786
R5130 DVDD.n5030 DVDD.n5029 0.214786
R5131 DVDD.n5028 DVDD.n583 0.214786
R5132 DVDD.n5027 DVDD.n5026 0.214786
R5133 DVDD.n591 DVDD.n585 0.214786
R5134 DVDD.n5022 DVDD.n5021 0.214786
R5135 DVDD.n588 DVDD.n587 0.214786
R5136 DVDD.n4787 DVDD.n4786 0.214786
R5137 DVDD.n4789 DVDD.n4788 0.214786
R5138 DVDD.n4790 DVDD.n4780 0.214786
R5139 DVDD.n4792 DVDD.n4791 0.214786
R5140 DVDD.n4793 DVDD.n4779 0.214786
R5141 DVDD.n4795 DVDD.n4794 0.214786
R5142 DVDD.n4796 DVDD.n4774 0.214786
R5143 DVDD.n4798 DVDD.n4797 0.214786
R5144 DVDD.n4799 DVDD.n734 0.214786
R5145 DVDD.n4801 DVDD.n4800 0.214786
R5146 DVDD.n4770 DVDD.n732 0.214786
R5147 DVDD.n4769 DVDD.n4768 0.214786
R5148 DVDD.n880 DVDD.n879 0.214786
R5149 DVDD.n4762 DVDD.n4761 0.214786
R5150 DVDD.n4760 DVDD.n882 0.214786
R5151 DVDD.n4759 DVDD.n4758 0.214786
R5152 DVDD.n884 DVDD.n883 0.214786
R5153 DVDD.n4754 DVDD.n4753 0.214786
R5154 DVDD.n4752 DVDD.n886 0.214786
R5155 DVDD.n4751 DVDD.n4750 0.214786
R5156 DVDD.n888 DVDD.n887 0.214786
R5157 DVDD.n4746 DVDD.n4745 0.214786
R5158 DVDD.n891 DVDD.n890 0.214786
R5159 DVDD.n4720 DVDD.n4719 0.214786
R5160 DVDD.n906 DVDD.n905 0.214786
R5161 DVDD.n4725 DVDD.n4724 0.214786
R5162 DVDD.n4726 DVDD.n904 0.214786
R5163 DVDD.n4728 DVDD.n4727 0.214786
R5164 DVDD.n902 DVDD.n901 0.214786
R5165 DVDD.n4733 DVDD.n4732 0.214786
R5166 DVDD.n4734 DVDD.n900 0.214786
R5167 DVDD.n4736 DVDD.n4735 0.214786
R5168 DVDD.n898 DVDD.n897 0.214786
R5169 DVDD.n4741 DVDD.n4740 0.214786
R5170 DVDD.n4330 DVDD.n4329 0.214786
R5171 DVDD.n4328 DVDD.n1628 0.214786
R5172 DVDD.n4327 DVDD.n1639 0.214786
R5173 DVDD.n4326 DVDD.n4325 0.214786
R5174 DVDD.n4324 DVDD.n4304 0.214786
R5175 DVDD.n4323 DVDD.n4322 0.214786
R5176 DVDD.n4321 DVDD.n4305 0.214786
R5177 DVDD.n4320 DVDD.n4319 0.214786
R5178 DVDD.n4318 DVDD.n4310 0.214786
R5179 DVDD.n4317 DVDD.n4316 0.214786
R5180 DVDD.n4315 DVDD.n4311 0.214786
R5181 DVDD.n4707 DVDD.n913 0.214786
R5182 DVDD.n4712 DVDD.n4711 0.214786
R5183 DVDD.n921 DVDD.n911 0.214786
R5184 DVDD.n4717 DVDD.n4716 0.214786
R5185 DVDD.n3648 DVDD 0.209823
R5186 DVDD.n961 DVDD.n960 0.208983
R5187 DVDD.n245 DVDD.n223 0.208899
R5188 DVDD.n2235 DVDD.n2234 0.208833
R5189 DVDD.n2231 DVDD.n2230 0.208833
R5190 DVDD.n2227 DVDD.n2226 0.208833
R5191 DVDD.n2223 DVDD.n2222 0.208833
R5192 DVDD.n2219 DVDD.n2218 0.208833
R5193 DVDD.n4203 DVDD.n4202 0.2085
R5194 DVDD.n4126 DVDD.n4125 0.2085
R5195 DVDD.n4121 DVDD.n4120 0.2085
R5196 DVDD.n4013 DVDD.n4012 0.2085
R5197 DVDD.n3994 DVDD.n3993 0.2085
R5198 DVDD.n3929 DVDD.n3928 0.2085
R5199 DVDD.n3932 DVDD.n3931 0.2085
R5200 DVDD.n1877 DVDD.n1876 0.2085
R5201 DVDD.n1868 DVDD.n1867 0.2085
R5202 DVDD.n1871 DVDD.n1870 0.2085
R5203 DVDD.n1716 DVDD.n1715 0.2085
R5204 DVDD.n4174 DVDD.n4173 0.2085
R5205 DVDD.n3652 DVDD.n1984 0.207972
R5206 DVDD.n3617 DVDD.n3092 0.2067
R5207 DVDD.n3652 DVDD.n1985 0.206229
R5208 DVDD.n3617 DVDD.n3091 0.205865
R5209 DVDD.n5423 DVDD.n5422 0.204558
R5210 DVDD.n5918 DVDD.n5917 0.204245
R5211 DVDD DVDD.n3648 0.202555
R5212 DVDD.n3092 DVDD.n2022 0.19985
R5213 DVDD.n3091 DVDD.n2022 0.199294
R5214 DVDD.n3647 DVDD.n1984 0.199041
R5215 DVDD.n3647 DVDD.n1985 0.198923
R5216 DVDD.n3516 DVDD.n3515 0.198598
R5217 DVDD.n4201 DVDD 0.191088
R5218 DVDD.n3992 DVDD 0.191088
R5219 DVDD.n4011 DVDD 0.191088
R5220 DVDD.n1869 DVDD 0.191088
R5221 DVDD.n2802 DVDD.n2799 0.190625
R5222 DVDD.n4229 DVDD.n4228 0.1805
R5223 DVDD.n2712 DVDD.n2705 0.179316
R5224 DVDD.n1952 DVDD 0.176947
R5225 DVDD.n2214 DVDD 0.17636
R5226 DVDD.n3652 DVDD.n1997 0.174559
R5227 DVDD.n1899 DVDD.n1896 0.174162
R5228 DVDD.n1743 DVDD.n1739 0.174048
R5229 DVDD.n3617 DVDD.n2025 0.173987
R5230 DVDD DVDD.n1742 0.173778
R5231 DVDD.n1886 DVDD.n1885 0.173043
R5232 DVDD.n2797 DVDD.n2706 0.172185
R5233 DVDD DVDD.n2024 0.172062
R5234 DVDD.n1900 DVDD 0.171551
R5235 DVDD.n2048 DVDD.n2041 0.168658
R5236 DVDD.n2059 DVDD.n2041 0.168658
R5237 DVDD.n2060 DVDD.n2059 0.168658
R5238 DVDD.n2073 DVDD.n2072 0.168658
R5239 DVDD.n2072 DVDD.n2069 0.168658
R5240 DVDD.n2069 DVDD.n2067 0.168658
R5241 DVDD.n2062 DVDD.n2039 0.168658
R5242 DVDD.n3068 DVDD.n2039 0.168658
R5243 DVDD.n3068 DVDD.n3067 0.168658
R5244 DVDD.n3042 DVDD.n2040 0.168658
R5245 DVDD.n3042 DVDD.n3035 0.168658
R5246 DVDD.n3053 DVDD.n3035 0.168658
R5247 DVDD.n4264 DVDD.n1682 0.168658
R5248 DVDD.n4264 DVDD.n4263 0.168658
R5249 DVDD.n4263 DVDD.n1683 0.168658
R5250 DVDD.n3813 DVDD.n1842 0.168658
R5251 DVDD.n3814 DVDD.n3813 0.168658
R5252 DVDD.n3815 DVDD.n3814 0.168658
R5253 DVDD.n4065 DVDD.n4064 0.168658
R5254 DVDD.n4064 DVDD.n4054 0.168658
R5255 DVDD.n4054 DVDD.n1719 0.168658
R5256 DVDD.n4226 DVDD.n1720 0.168658
R5257 DVDD.n1762 DVDD.n1720 0.168658
R5258 DVDD.n1762 DVDD.n1761 0.168658
R5259 DVDD.n1740 DVDD.n1739 0.16842
R5260 DVDD.n2025 DVDD.n2022 0.167884
R5261 DVDD.n3704 DVDD.n1899 0.16771
R5262 DVDD.n1742 DVDD 0.167454
R5263 DVDD.n3647 DVDD.n1997 0.16731
R5264 DVDD DVDD.n1900 0.166755
R5265 DVDD.n5486 DVDD.n263 0.165735
R5266 DVDD.n2024 DVDD 0.165645
R5267 DVDD.n5660 DVDD.n259 0.165589
R5268 DVDD.n1364 DVDD.n1363 0.164191
R5269 DVDD.n1576 DVDD.n1193 0.163126
R5270 DVDD.n2717 DVDD 0.160647
R5271 DVDD.n4202 DVDD.t125 0.152167
R5272 DVDD.n4202 DVDD.t127 0.152167
R5273 DVDD.n4125 DVDD.t186 0.152167
R5274 DVDD.n4125 DVDD.t164 0.152167
R5275 DVDD.n4120 DVDD.t64 0.152167
R5276 DVDD.n4120 DVDD.t28 0.152167
R5277 DVDD.n4012 DVDD.t57 0.152167
R5278 DVDD.n4012 DVDD.t59 0.152167
R5279 DVDD.n3993 DVDD.t42 0.152167
R5280 DVDD.n3993 DVDD.t44 0.152167
R5281 DVDD.n3928 DVDD.t6 0.152167
R5282 DVDD.n3928 DVDD.t198 0.152167
R5283 DVDD.n3931 DVDD.t87 0.152167
R5284 DVDD.n3931 DVDD.t81 0.152167
R5285 DVDD.n1876 DVDD.t17 0.152167
R5286 DVDD.n1876 DVDD.t8 0.152167
R5287 DVDD.n1867 DVDD.t130 0.152167
R5288 DVDD.n1867 DVDD.t139 0.152167
R5289 DVDD.n1870 DVDD.t192 0.152167
R5290 DVDD.n1870 DVDD.t3 0.152167
R5291 DVDD.n1715 DVDD.t133 0.152167
R5292 DVDD.n1715 DVDD.t147 0.152167
R5293 DVDD.n4173 DVDD.t20 0.152167
R5294 DVDD.n4173 DVDD.t112 0.152167
R5295 DVDD.n3026 DVDD.n2076 0.145128
R5296 DVDD.n1883 DVDD.n1882 0.144974
R5297 DVDD.n4188 DVDD.n1718 0.144974
R5298 DVDD.n2462 DVDD.n2326 0.140794
R5299 DVDD.n2351 DVDD.n2326 0.140794
R5300 DVDD.n2537 DVDD.n2262 0.140794
R5301 DVDD.n2285 DVDD.n2262 0.140794
R5302 DVDD.n5488 DVDD.n264 0.1405
R5303 DVDD.n5488 DVDD.n5487 0.1405
R5304 DVDD.n5663 DVDD.n5662 0.1405
R5305 DVDD.n5662 DVDD.n5661 0.1405
R5306 DVDD.n2351 DVDD 0.131529
R5307 DVDD DVDD.n2462 0.131529
R5308 DVDD.n2285 DVDD 0.131529
R5309 DVDD DVDD.n2537 0.131529
R5310 DVDD.n2399 DVDD 0.130618
R5311 DVDD.n2981 DVDD 0.130618
R5312 DVDD.n1363 DVDD 0.124869
R5313 DVDD.n2014 DVDD 0.123988
R5314 DVDD.n3662 DVDD 0.123988
R5315 DVDD.n2011 DVDD 0.123988
R5316 DVDD.n3659 DVDD 0.123988
R5317 DVDD.n1570 DVDD.n1193 0.122916
R5318 DVDD.n1959 DVDD.n1958 0.120105
R5319 DVDD.n3691 DVDD 0.115647
R5320 DVDD.n1961 DVDD.n1960 0.114898
R5321 DVDD.n1933 DVDD.n1932 0.114898
R5322 DVDD.n1937 DVDD.n1936 0.114153
R5323 DVDD.n3697 DVDD.n3696 0.114153
R5324 DVDD.n3330 DVDD.n3278 0.112392
R5325 DVDD.n3317 DVDD.n3242 0.112392
R5326 DVDD.n4122 DVDD.n1711 0.111676
R5327 DVDD.n3930 DVDD.n1709 0.111676
R5328 DVDD.n1151 DVDD.n1150 0.110634
R5329 DVDD.n4399 DVDD.n1106 0.110634
R5330 DVDD.n4346 DVDD.n4345 0.110634
R5331 DVDD.n4301 DVDD.n4300 0.110634
R5332 DVDD.n3255 DVDD.n3247 0.110634
R5333 DVDD.n3303 DVDD.n3273 0.110634
R5334 DVDD.n2053 DVDD.n2044 0.110634
R5335 DVDD.n3731 DVDD.n3721 0.110634
R5336 DVDD DVDD.n1957 0.109447
R5337 DVDD.n1919 DVDD 0.109447
R5338 DVDD DVDD.n1923 0.109447
R5339 DVDD.n3393 DVDD.n3226 0.1055
R5340 DVDD.n3346 DVDD.n3226 0.1055
R5341 DVDD.n3321 DVDD.n3320 0.1055
R5342 DVDD.n3322 DVDD.n3321 0.1055
R5343 DVDD DVDD.n2399 0.10093
R5344 DVDD DVDD.n2981 0.10093
R5345 DVDD.n2793 DVDD.n2792 0.0931471
R5346 DVDD.n2792 DVDD.n2791 0.0931471
R5347 DVDD.n2074 DVDD.n2060 0.084579
R5348 DVDD.n2074 DVDD.n2073 0.084579
R5349 DVDD.n3067 DVDD.n3066 0.084579
R5350 DVDD.n3066 DVDD.n2040 0.084579
R5351 DVDD.n1880 DVDD.n1683 0.084579
R5352 DVDD.n1880 DVDD.n1842 0.084579
R5353 DVDD.n4227 DVDD.n1719 0.084579
R5354 DVDD.n4227 DVDD.n4226 0.084579
R5355 DVDD.n4385 DVDD.n4344 0.0815
R5356 DVDD.n4413 DVDD.n4387 0.0815
R5357 DVDD DVDD.n2716 0.0799118
R5358 DVDD.n1882 DVDD.n1881 0.0798421
R5359 DVDD.n1584 DVDD.n1583 0.079359
R5360 DVDD.n2794 DVDD.n2793 0.0786579
R5361 DVDD.n4198 DVDD.n4197 0.0780879
R5362 DVDD.n3774 DVDD.n3773 0.077225
R5363 DVDD.n3697 DVDD.n3687 0.0760366
R5364 DVDD.n1937 DVDD.n1905 0.0760366
R5365 DVDD.n1961 DVDD.n1947 0.0757132
R5366 DVDD.n1932 DVDD.n1926 0.0757132
R5367 DVDD.n3025 DVDD.n3024 0.0737558
R5368 DVDD.n3026 DVDD.n3025 0.0737558
R5369 DVDD.n3237 DVDD.n3226 0.066125
R5370 DVDD.n3321 DVDD.n3319 0.066125
R5371 DVDD.n5896 DVDD 0.0638222
R5372 DVDD.n5590 DVDD 0.0638222
R5373 DVDD.n5971 DVDD 0.0638222
R5374 DVDD.n5688 DVDD 0.0638222
R5375 DVDD.n3324 DVDD.n3244 0.0624947
R5376 DVDD.n3325 DVDD.n3324 0.0624947
R5377 DVDD.n4197 DVDD 0.0592637
R5378 DVDD.n3695 DVDD.n3694 0.0574118
R5379 DVDD.n5631 DVDD.n5630 0.0560556
R5380 DVDD.n5537 DVDD.n13 0.0560556
R5381 DVDD.n4676 DVDD.n980 0.0560556
R5382 DVDD.n5456 DVDD.n5455 0.0560556
R5383 DVDD.n1904 DVDD.n1897 0.0527336
R5384 DVDD.n1946 DVDD.n1897 0.0527336
R5385 DVDD.n5500 DVDD.n260 0.0523993
R5386 DVDD.n3617 DVDD.n3090 0.0518309
R5387 DVDD.n1998 DVDD.n1994 0.0515891
R5388 DVDD.n1998 DVDD.n1988 0.0515891
R5389 DVDD.n1998 DVDD.n1986 0.0515891
R5390 DVDD.n4080 DVDD.n4044 0.0515891
R5391 DVDD.n3901 DVDD.n3900 0.0515891
R5392 DVDD.n1898 DVDD.n1897 0.0515834
R5393 DVDD.n3087 DVDD.n2023 0.0515834
R5394 DVDD.n3094 DVDD.n2023 0.0515834
R5395 DVDD.n3832 DVDD.n1830 0.0515834
R5396 DVDD.n4044 DVDD.n4043 0.0509336
R5397 DVDD.n3090 DVDD.n2022 0.0505959
R5398 DVDD.n3900 DVDD.n3868 0.0503876
R5399 DVDD.n1945 DVDD.n1897 0.0497891
R5400 DVDD.n1967 DVDD.n1897 0.0497891
R5401 DVDD.n1998 DVDD.n1987 0.0497849
R5402 DVDD.n1998 DVDD.n1989 0.0497849
R5403 DVDD.n1998 DVDD.n1982 0.0497849
R5404 DVDD.n1831 DVDD.n1830 0.0497834
R5405 DVDD.n3088 DVDD.n2023 0.0497834
R5406 DVDD.n3093 DVDD.n2023 0.0497834
R5407 DVDD DVDD.n5896 0.0487259
R5408 DVDD DVDD.n5590 0.0487259
R5409 DVDD DVDD.n5971 0.0487259
R5410 DVDD DVDD.n5688 0.0487259
R5411 DVDD.n3477 DVDD.n3476 0.0467228
R5412 DVDD.n3560 DVDD.n3559 0.0467228
R5413 DVDD.n5730 DVDD.n194 0.0462377
R5414 DVDD.n5736 DVDD.n194 0.0462377
R5415 DVDD.n5737 DVDD.n5736 0.0462377
R5416 DVDD.n5737 DVDD.n192 0.0462377
R5417 DVDD.n5741 DVDD.n192 0.0462377
R5418 DVDD.n5742 DVDD.n5741 0.0462377
R5419 DVDD.n5745 DVDD.n5742 0.0462377
R5420 DVDD.n5747 DVDD.n5745 0.0462377
R5421 DVDD.n5749 DVDD.n5747 0.0462377
R5422 DVDD.n5751 DVDD.n5749 0.0462377
R5423 DVDD.n5753 DVDD.n5751 0.0462377
R5424 DVDD.n5755 DVDD.n5753 0.0462377
R5425 DVDD.n5757 DVDD.n5755 0.0462377
R5426 DVDD.n5758 DVDD.n5757 0.0462377
R5427 DVDD.n5761 DVDD.n5758 0.0462377
R5428 DVDD.n5763 DVDD.n5761 0.0462377
R5429 DVDD.n5765 DVDD.n5763 0.0462377
R5430 DVDD.n5767 DVDD.n5765 0.0462377
R5431 DVDD.n5769 DVDD.n5767 0.0462377
R5432 DVDD.n5771 DVDD.n5769 0.0462377
R5433 DVDD.n5772 DVDD.n5771 0.0462377
R5434 DVDD.n5780 DVDD.n5772 0.0462377
R5435 DVDD.n5780 DVDD.n5779 0.0462377
R5436 DVDD.n5779 DVDD.n5778 0.0462377
R5437 DVDD.n5778 DVDD.n5776 0.0462377
R5438 DVDD.n5776 DVDD.n5774 0.0462377
R5439 DVDD.n5774 DVDD.n167 0.0462377
R5440 DVDD.n5786 DVDD.n167 0.0462377
R5441 DVDD.n5787 DVDD.n5786 0.0462377
R5442 DVDD.n5791 DVDD.n165 0.0462377
R5443 DVDD.n5792 DVDD.n5791 0.0462377
R5444 DVDD.n5831 DVDD.n5792 0.0462377
R5445 DVDD.n5831 DVDD.n5830 0.0462377
R5446 DVDD.n5830 DVDD.n5827 0.0462377
R5447 DVDD.n5827 DVDD.n5826 0.0462377
R5448 DVDD.n5826 DVDD.n5824 0.0462377
R5449 DVDD.n5824 DVDD.n5822 0.0462377
R5450 DVDD.n5822 DVDD.n5820 0.0462377
R5451 DVDD.n5820 DVDD.n5818 0.0462377
R5452 DVDD.n5818 DVDD.n5816 0.0462377
R5453 DVDD.n5816 DVDD.n5814 0.0462377
R5454 DVDD.n5814 DVDD.n5811 0.0462377
R5455 DVDD.n5811 DVDD.n5810 0.0462377
R5456 DVDD.n5810 DVDD.n5808 0.0462377
R5457 DVDD.n5808 DVDD.n5806 0.0462377
R5458 DVDD.n5806 DVDD.n5804 0.0462377
R5459 DVDD.n5804 DVDD.n5802 0.0462377
R5460 DVDD.n5802 DVDD.n5800 0.0462377
R5461 DVDD.n5800 DVDD.n5798 0.0462377
R5462 DVDD.n5798 DVDD.n5795 0.0462377
R5463 DVDD.n5795 DVDD.n5794 0.0462377
R5464 DVDD.n5794 DVDD.n141 0.0462377
R5465 DVDD.n5837 DVDD.n141 0.0462377
R5466 DVDD.n5838 DVDD.n5837 0.0462377
R5467 DVDD.n5838 DVDD.n139 0.0462377
R5468 DVDD.n5842 DVDD.n139 0.0462377
R5469 DVDD.n5844 DVDD.n5842 0.0462377
R5470 DVDD.n5846 DVDD.n5844 0.0462377
R5471 DVDD.n5739 DVDD.n5738 0.0462377
R5472 DVDD.n5740 DVDD.n5739 0.0462377
R5473 DVDD.n5744 DVDD.n5743 0.0462377
R5474 DVDD.n5760 DVDD.n5759 0.0462377
R5475 DVDD.n5781 DVDD.n191 0.0462377
R5476 DVDD.n5789 DVDD.n5788 0.0462377
R5477 DVDD.n5790 DVDD.n5789 0.0462377
R5478 DVDD.n5829 DVDD.n5828 0.0462377
R5479 DVDD.n5813 DVDD.n5812 0.0462377
R5480 DVDD.n5797 DVDD.n5796 0.0462377
R5481 DVDD.n5840 DVDD.n5839 0.0462377
R5482 DVDD.n5841 DVDD.n5840 0.0462377
R5483 DVDD.n5091 DVDD.n5090 0.0462377
R5484 DVDD.n5090 DVDD.n5088 0.0462377
R5485 DVDD.n5088 DVDD.n568 0.0462377
R5486 DVDD.n5098 DVDD.n568 0.0462377
R5487 DVDD.n5099 DVDD.n5098 0.0462377
R5488 DVDD.n5239 DVDD.n5099 0.0462377
R5489 DVDD.n5239 DVDD.n5238 0.0462377
R5490 DVDD.n5238 DVDD.n5237 0.0462377
R5491 DVDD.n5237 DVDD.n5235 0.0462377
R5492 DVDD.n5235 DVDD.n5233 0.0462377
R5493 DVDD.n5233 DVDD.n5231 0.0462377
R5494 DVDD.n5231 DVDD.n5229 0.0462377
R5495 DVDD.n5229 DVDD.n5227 0.0462377
R5496 DVDD.n5227 DVDD.n5225 0.0462377
R5497 DVDD.n5225 DVDD.n5222 0.0462377
R5498 DVDD.n5222 DVDD.n5221 0.0462377
R5499 DVDD.n5221 DVDD.n5219 0.0462377
R5500 DVDD.n5219 DVDD.n5217 0.0462377
R5501 DVDD.n5217 DVDD.n5215 0.0462377
R5502 DVDD.n5215 DVDD.n5213 0.0462377
R5503 DVDD.n5213 DVDD.n5211 0.0462377
R5504 DVDD.n5211 DVDD.n5209 0.0462377
R5505 DVDD.n5209 DVDD.n5206 0.0462377
R5506 DVDD.n5206 DVDD.n5205 0.0462377
R5507 DVDD.n5205 DVDD.n5203 0.0462377
R5508 DVDD.n5203 DVDD.n5201 0.0462377
R5509 DVDD.n5201 DVDD.n5199 0.0462377
R5510 DVDD.n5199 DVDD.n5197 0.0462377
R5511 DVDD.n5197 DVDD.n5195 0.0462377
R5512 DVDD.n5191 DVDD.n5100 0.0462377
R5513 DVDD.n5191 DVDD.n5190 0.0462377
R5514 DVDD.n5190 DVDD.n5188 0.0462377
R5515 DVDD.n5188 DVDD.n5186 0.0462377
R5516 DVDD.n5186 DVDD.n5183 0.0462377
R5517 DVDD.n5183 DVDD.n5182 0.0462377
R5518 DVDD.n5182 DVDD.n5180 0.0462377
R5519 DVDD.n5180 DVDD.n5178 0.0462377
R5520 DVDD.n5178 DVDD.n5176 0.0462377
R5521 DVDD.n5176 DVDD.n5174 0.0462377
R5522 DVDD.n5174 DVDD.n5172 0.0462377
R5523 DVDD.n5172 DVDD.n5170 0.0462377
R5524 DVDD.n5170 DVDD.n5167 0.0462377
R5525 DVDD.n5167 DVDD.n5166 0.0462377
R5526 DVDD.n5166 DVDD.n5164 0.0462377
R5527 DVDD.n5164 DVDD.n5162 0.0462377
R5528 DVDD.n5162 DVDD.n5160 0.0462377
R5529 DVDD.n5160 DVDD.n5158 0.0462377
R5530 DVDD.n5158 DVDD.n5156 0.0462377
R5531 DVDD.n5156 DVDD.n5154 0.0462377
R5532 DVDD.n5154 DVDD.n5151 0.0462377
R5533 DVDD.n5151 DVDD.n5150 0.0462377
R5534 DVDD.n5150 DVDD.n5148 0.0462377
R5535 DVDD.n5148 DVDD.n5147 0.0462377
R5536 DVDD.n5147 DVDD.n5146 0.0462377
R5537 DVDD.n5146 DVDD.n5101 0.0462377
R5538 DVDD.n5142 DVDD.n5101 0.0462377
R5539 DVDD.n5142 DVDD.n5141 0.0462377
R5540 DVDD.n5141 DVDD.n5103 0.0462377
R5541 DVDD.n5097 DVDD.n5096 0.0462377
R5542 DVDD.n5097 DVDD.n566 0.0462377
R5543 DVDD.n5240 DVDD.n567 0.0462377
R5544 DVDD.n5224 DVDD.n5223 0.0462377
R5545 DVDD.n5208 DVDD.n5207 0.0462377
R5546 DVDD.n5194 DVDD.n5193 0.0462377
R5547 DVDD.n5193 DVDD.n5192 0.0462377
R5548 DVDD.n5185 DVDD.n5184 0.0462377
R5549 DVDD.n5169 DVDD.n5168 0.0462377
R5550 DVDD.n5153 DVDD.n5152 0.0462377
R5551 DVDD.n5145 DVDD.n5144 0.0462377
R5552 DVDD.n5144 DVDD.n5143 0.0462377
R5553 DVDD.n600 DVDD.n598 0.0462377
R5554 DVDD.n601 DVDD.n600 0.0462377
R5555 DVDD.n5017 DVDD.n601 0.0462377
R5556 DVDD.n5017 DVDD.n5016 0.0462377
R5557 DVDD.n5016 DVDD.n5015 0.0462377
R5558 DVDD.n5015 DVDD.n602 0.0462377
R5559 DVDD.n629 DVDD.n602 0.0462377
R5560 DVDD.n631 DVDD.n629 0.0462377
R5561 DVDD.n633 DVDD.n631 0.0462377
R5562 DVDD.n635 DVDD.n633 0.0462377
R5563 DVDD.n637 DVDD.n635 0.0462377
R5564 DVDD.n639 DVDD.n637 0.0462377
R5565 DVDD.n641 DVDD.n639 0.0462377
R5566 DVDD.n642 DVDD.n641 0.0462377
R5567 DVDD.n645 DVDD.n642 0.0462377
R5568 DVDD.n647 DVDD.n645 0.0462377
R5569 DVDD.n649 DVDD.n647 0.0462377
R5570 DVDD.n651 DVDD.n649 0.0462377
R5571 DVDD.n653 DVDD.n651 0.0462377
R5572 DVDD.n655 DVDD.n653 0.0462377
R5573 DVDD.n657 DVDD.n655 0.0462377
R5574 DVDD.n658 DVDD.n657 0.0462377
R5575 DVDD.n661 DVDD.n658 0.0462377
R5576 DVDD.n663 DVDD.n661 0.0462377
R5577 DVDD.n665 DVDD.n663 0.0462377
R5578 DVDD.n667 DVDD.n665 0.0462377
R5579 DVDD.n669 DVDD.n667 0.0462377
R5580 DVDD.n670 DVDD.n669 0.0462377
R5581 DVDD.n5009 DVDD.n670 0.0462377
R5582 DVDD.n5008 DVDD.n5007 0.0462377
R5583 DVDD.n5007 DVDD.n671 0.0462377
R5584 DVDD.n4951 DVDD.n671 0.0462377
R5585 DVDD.n4952 DVDD.n4951 0.0462377
R5586 DVDD.n4955 DVDD.n4952 0.0462377
R5587 DVDD.n4957 DVDD.n4955 0.0462377
R5588 DVDD.n4959 DVDD.n4957 0.0462377
R5589 DVDD.n4961 DVDD.n4959 0.0462377
R5590 DVDD.n4963 DVDD.n4961 0.0462377
R5591 DVDD.n4965 DVDD.n4963 0.0462377
R5592 DVDD.n4967 DVDD.n4965 0.0462377
R5593 DVDD.n4968 DVDD.n4967 0.0462377
R5594 DVDD.n4971 DVDD.n4968 0.0462377
R5595 DVDD.n4973 DVDD.n4971 0.0462377
R5596 DVDD.n4975 DVDD.n4973 0.0462377
R5597 DVDD.n4977 DVDD.n4975 0.0462377
R5598 DVDD.n4979 DVDD.n4977 0.0462377
R5599 DVDD.n4981 DVDD.n4979 0.0462377
R5600 DVDD.n4983 DVDD.n4981 0.0462377
R5601 DVDD.n4984 DVDD.n4983 0.0462377
R5602 DVDD.n4987 DVDD.n4984 0.0462377
R5603 DVDD.n4989 DVDD.n4987 0.0462377
R5604 DVDD.n4990 DVDD.n4989 0.0462377
R5605 DVDD.n5001 DVDD.n4990 0.0462377
R5606 DVDD.n5001 DVDD.n5000 0.0462377
R5607 DVDD.n5000 DVDD.n4991 0.0462377
R5608 DVDD.n4996 DVDD.n4991 0.0462377
R5609 DVDD.n4996 DVDD.n4995 0.0462377
R5610 DVDD.n4995 DVDD.n4993 0.0462377
R5611 DVDD.n5018 DVDD.n595 0.0462377
R5612 DVDD.n5014 DVDD.n595 0.0462377
R5613 DVDD.n628 DVDD.n604 0.0462377
R5614 DVDD.n644 DVDD.n643 0.0462377
R5615 DVDD.n660 DVDD.n659 0.0462377
R5616 DVDD.n5010 DVDD.n627 0.0462377
R5617 DVDD.n5006 DVDD.n627 0.0462377
R5618 DVDD.n4954 DVDD.n4953 0.0462377
R5619 DVDD.n4970 DVDD.n4969 0.0462377
R5620 DVDD.n4986 DVDD.n4985 0.0462377
R5621 DVDD.n4999 DVDD.n4998 0.0462377
R5622 DVDD.n4998 DVDD.n4997 0.0462377
R5623 DVDD.n877 DVDD.n875 0.0462377
R5624 DVDD.n875 DVDD.n873 0.0462377
R5625 DVDD.n873 DVDD.n871 0.0462377
R5626 DVDD.n871 DVDD.n868 0.0462377
R5627 DVDD.n868 DVDD.n867 0.0462377
R5628 DVDD.n867 DVDD.n866 0.0462377
R5629 DVDD.n866 DVDD.n865 0.0462377
R5630 DVDD.n865 DVDD.n863 0.0462377
R5631 DVDD.n863 DVDD.n861 0.0462377
R5632 DVDD.n861 DVDD.n859 0.0462377
R5633 DVDD.n859 DVDD.n857 0.0462377
R5634 DVDD.n857 DVDD.n855 0.0462377
R5635 DVDD.n855 DVDD.n853 0.0462377
R5636 DVDD.n853 DVDD.n851 0.0462377
R5637 DVDD.n851 DVDD.n848 0.0462377
R5638 DVDD.n848 DVDD.n847 0.0462377
R5639 DVDD.n847 DVDD.n845 0.0462377
R5640 DVDD.n845 DVDD.n843 0.0462377
R5641 DVDD.n843 DVDD.n841 0.0462377
R5642 DVDD.n841 DVDD.n839 0.0462377
R5643 DVDD.n839 DVDD.n837 0.0462377
R5644 DVDD.n837 DVDD.n835 0.0462377
R5645 DVDD.n835 DVDD.n832 0.0462377
R5646 DVDD.n832 DVDD.n831 0.0462377
R5647 DVDD.n831 DVDD.n829 0.0462377
R5648 DVDD.n829 DVDD.n827 0.0462377
R5649 DVDD.n827 DVDD.n825 0.0462377
R5650 DVDD.n825 DVDD.n823 0.0462377
R5651 DVDD.n823 DVDD.n821 0.0462377
R5652 DVDD.n817 DVDD.n739 0.0462377
R5653 DVDD.n817 DVDD.n816 0.0462377
R5654 DVDD.n816 DVDD.n741 0.0462377
R5655 DVDD.n810 DVDD.n741 0.0462377
R5656 DVDD.n810 DVDD.n809 0.0462377
R5657 DVDD.n809 DVDD.n808 0.0462377
R5658 DVDD.n808 DVDD.n743 0.0462377
R5659 DVDD.n802 DVDD.n743 0.0462377
R5660 DVDD.n802 DVDD.n801 0.0462377
R5661 DVDD.n801 DVDD.n746 0.0462377
R5662 DVDD.n795 DVDD.n746 0.0462377
R5663 DVDD.n795 DVDD.n794 0.0462377
R5664 DVDD.n794 DVDD.n748 0.0462377
R5665 DVDD.n789 DVDD.n748 0.0462377
R5666 DVDD.n789 DVDD.n788 0.0462377
R5667 DVDD.n788 DVDD.n750 0.0462377
R5668 DVDD.n782 DVDD.n750 0.0462377
R5669 DVDD.n782 DVDD.n781 0.0462377
R5670 DVDD.n781 DVDD.n752 0.0462377
R5671 DVDD.n775 DVDD.n752 0.0462377
R5672 DVDD.n775 DVDD.n774 0.0462377
R5673 DVDD.n774 DVDD.n773 0.0462377
R5674 DVDD.n773 DVDD.n754 0.0462377
R5675 DVDD.n767 DVDD.n754 0.0462377
R5676 DVDD.n767 DVDD.n766 0.0462377
R5677 DVDD.n766 DVDD.n757 0.0462377
R5678 DVDD.n762 DVDD.n757 0.0462377
R5679 DVDD.n762 DVDD.n761 0.0462377
R5680 DVDD.n761 DVDD.n759 0.0462377
R5681 DVDD.n870 DVDD.n869 0.0462377
R5682 DVDD.n869 DVDD.n726 0.0462377
R5683 DVDD.n864 DVDD.n727 0.0462377
R5684 DVDD.n850 DVDD.n849 0.0462377
R5685 DVDD.n834 DVDD.n833 0.0462377
R5686 DVDD.n820 DVDD.n819 0.0462377
R5687 DVDD.n819 DVDD.n818 0.0462377
R5688 DVDD.n811 DVDD.n742 0.0462377
R5689 DVDD.n793 DVDD.n792 0.0462377
R5690 DVDD.n776 DVDD.n753 0.0462377
R5691 DVDD.n765 DVDD.n764 0.0462377
R5692 DVDD.n764 DVDD.n763 0.0462377
R5693 DVDD.n1062 DVDD.n1060 0.0462377
R5694 DVDD.n1064 DVDD.n1062 0.0462377
R5695 DVDD.n1065 DVDD.n1064 0.0462377
R5696 DVDD.n1068 DVDD.n1065 0.0462377
R5697 DVDD.n1069 DVDD.n1068 0.0462377
R5698 DVDD.n4612 DVDD.n1069 0.0462377
R5699 DVDD.n4612 DVDD.n4611 0.0462377
R5700 DVDD.n4611 DVDD.n4610 0.0462377
R5701 DVDD.n4610 DVDD.n4608 0.0462377
R5702 DVDD.n4608 DVDD.n4606 0.0462377
R5703 DVDD.n4606 DVDD.n4604 0.0462377
R5704 DVDD.n4604 DVDD.n4602 0.0462377
R5705 DVDD.n4602 DVDD.n4600 0.0462377
R5706 DVDD.n4600 DVDD.n4598 0.0462377
R5707 DVDD.n4598 DVDD.n4595 0.0462377
R5708 DVDD.n4595 DVDD.n4594 0.0462377
R5709 DVDD.n4594 DVDD.n4592 0.0462377
R5710 DVDD.n4592 DVDD.n4590 0.0462377
R5711 DVDD.n4590 DVDD.n4588 0.0462377
R5712 DVDD.n4588 DVDD.n4586 0.0462377
R5713 DVDD.n4586 DVDD.n4584 0.0462377
R5714 DVDD.n4584 DVDD.n4582 0.0462377
R5715 DVDD.n4582 DVDD.n4579 0.0462377
R5716 DVDD.n4579 DVDD.n4578 0.0462377
R5717 DVDD.n4578 DVDD.n4576 0.0462377
R5718 DVDD.n4576 DVDD.n4574 0.0462377
R5719 DVDD.n4574 DVDD.n4572 0.0462377
R5720 DVDD.n4572 DVDD.n4570 0.0462377
R5721 DVDD.n4570 DVDD.n4568 0.0462377
R5722 DVDD.n4564 DVDD.n1070 0.0462377
R5723 DVDD.n4564 DVDD.n4563 0.0462377
R5724 DVDD.n4563 DVDD.n1072 0.0462377
R5725 DVDD.n4508 DVDD.n1072 0.0462377
R5726 DVDD.n4511 DVDD.n4508 0.0462377
R5727 DVDD.n4513 DVDD.n4511 0.0462377
R5728 DVDD.n4515 DVDD.n4513 0.0462377
R5729 DVDD.n4517 DVDD.n4515 0.0462377
R5730 DVDD.n4519 DVDD.n4517 0.0462377
R5731 DVDD.n4521 DVDD.n4519 0.0462377
R5732 DVDD.n4523 DVDD.n4521 0.0462377
R5733 DVDD.n4524 DVDD.n4523 0.0462377
R5734 DVDD.n4527 DVDD.n4524 0.0462377
R5735 DVDD.n4529 DVDD.n4527 0.0462377
R5736 DVDD.n4531 DVDD.n4529 0.0462377
R5737 DVDD.n4533 DVDD.n4531 0.0462377
R5738 DVDD.n4535 DVDD.n4533 0.0462377
R5739 DVDD.n4537 DVDD.n4535 0.0462377
R5740 DVDD.n4539 DVDD.n4537 0.0462377
R5741 DVDD.n4540 DVDD.n4539 0.0462377
R5742 DVDD.n4543 DVDD.n4540 0.0462377
R5743 DVDD.n4545 DVDD.n4543 0.0462377
R5744 DVDD.n4546 DVDD.n4545 0.0462377
R5745 DVDD.n4557 DVDD.n4546 0.0462377
R5746 DVDD.n4557 DVDD.n4556 0.0462377
R5747 DVDD.n4556 DVDD.n4547 0.0462377
R5748 DVDD.n4552 DVDD.n4547 0.0462377
R5749 DVDD.n4552 DVDD.n4551 0.0462377
R5750 DVDD.n4551 DVDD.n4549 0.0462377
R5751 DVDD.n1067 DVDD.n1066 0.0462377
R5752 DVDD.n1067 DVDD.n1057 0.0462377
R5753 DVDD.n4613 DVDD.n1058 0.0462377
R5754 DVDD.n4597 DVDD.n4596 0.0462377
R5755 DVDD.n4581 DVDD.n4580 0.0462377
R5756 DVDD.n4567 DVDD.n4566 0.0462377
R5757 DVDD.n4566 DVDD.n4565 0.0462377
R5758 DVDD.n4510 DVDD.n4509 0.0462377
R5759 DVDD.n4526 DVDD.n4525 0.0462377
R5760 DVDD.n4542 DVDD.n4541 0.0462377
R5761 DVDD.n4555 DVDD.n4554 0.0462377
R5762 DVDD.n4554 DVDD.n4553 0.0462377
R5763 DVDD.n5511 DVDD.n28 0.0462377
R5764 DVDD.n4700 DVDD.n949 0.0462377
R5765 DVDD.n5787 DVDD.n165 0.0462377
R5766 DVDD.n5195 DVDD.n5100 0.0462377
R5767 DVDD.n5009 DVDD.n5008 0.0462377
R5768 DVDD.n821 DVDD.n739 0.0462377
R5769 DVDD.n4568 DVDD.n1070 0.0462377
R5770 DVDD.n3324 DVDD.n3323 0.0461522
R5771 DVDD.n3342 DVDD.n3341 0.0452755
R5772 DVDD.n5825 DVDD.n163 0.0451311
R5773 DVDD.n5181 DVDD.n468 0.0451311
R5774 DVDD.n4956 DVDD.n4944 0.0451311
R5775 DVDD.n807 DVDD.n744 0.0451311
R5776 DVDD.n4512 DVDD.n4503 0.0451311
R5777 DVDD.n5746 DVDD.n174 0.0447623
R5778 DVDD.n5236 DVDD.n486 0.0447623
R5779 DVDD.n630 DVDD.n610 0.0447623
R5780 DVDD.n862 DVDD.n705 0.0447623
R5781 DVDD.n4609 DVDD.n1010 0.0447623
R5782 DVDD.n1382 DVDD.n1313 0.0446743
R5783 DVDD.n1390 DVDD.n1309 0.0446743
R5784 DVDD.n1318 DVDD.n1216 0.0446743
R5785 DVDD.n1314 DVDD.n1214 0.0446743
R5786 DVDD.n5655 DVDD.n5654 0.0445261
R5787 DVDD.n5481 DVDD.n5480 0.0445261
R5788 DVDD.n5809 DVDD.n150 0.0443934
R5789 DVDD.n5165 DVDD.n466 0.0443934
R5790 DVDD.n4972 DVDD.n4942 0.0443934
R5791 DVDD.n791 DVDD.n790 0.0443934
R5792 DVDD.n4528 DVDD.n4501 0.0443934
R5793 DVDD.n3308 DVDD.n3280 0.0442838
R5794 DVDD.n3259 DVDD.n3233 0.0442838
R5795 DVDD.n3264 DVDD.n3263 0.0442838
R5796 DVDD.n3264 DVDD.n3235 0.0442838
R5797 DVDD.n3386 DVDD.n3385 0.0442838
R5798 DVDD.n3365 DVDD.n3364 0.0442838
R5799 DVDD.n3364 DVDD.n3279 0.0442838
R5800 DVDD.n3355 DVDD.n3339 0.0442838
R5801 DVDD.n5762 DVDD.n176 0.0440246
R5802 DVDD.n5220 DVDD.n562 0.0440246
R5803 DVDD.n646 DVDD.n612 0.0440246
R5804 DVDD.n846 DVDD.n722 0.0440246
R5805 DVDD.n4593 DVDD.n1053 0.0440246
R5806 DVDD.n5793 DVDD.n156 0.0436557
R5807 DVDD.n5149 DVDD.n464 0.0436557
R5808 DVDD.n4988 DVDD.n4940 0.0436557
R5809 DVDD.n772 DVDD.n755 0.0436557
R5810 DVDD.n4544 DVDD.n4499 0.0436557
R5811 DVDD.n3385 DVDD.n3384 0.043473
R5812 DVDD.n3339 DVDD.n3338 0.043473
R5813 DVDD.n5777 DVDD.n178 0.0432869
R5814 DVDD.n5204 DVDD.n493 0.0432869
R5815 DVDD.n662 DVDD.n614 0.0432869
R5816 DVDD.n830 DVDD.n712 0.0432869
R5817 DVDD.n4577 DVDD.n1017 0.0432869
R5818 DVDD.n5927 DVDD.n5926 0.0428146
R5819 DVDD.n5430 DVDD.n296 0.0428146
R5820 DVDD.n5782 DVDD.n190 0.0425492
R5821 DVDD.n5210 DVDD.n559 0.0425492
R5822 DVDD.n656 DVDD.n625 0.0425492
R5823 DVDD.n836 DVDD.n719 0.0425492
R5824 DVDD.n4583 DVDD.n1050 0.0425492
R5825 DVDD.n5799 DVDD.n153 0.0421803
R5826 DVDD.n5155 DVDD.n452 0.0421803
R5827 DVDD.n4982 DVDD.n675 0.0421803
R5828 DVDD.n778 DVDD.n777 0.0421803
R5829 DVDD.n4538 DVDD.n1076 0.0421803
R5830 DVDD.n5756 DVDD.n172 0.0418115
R5831 DVDD.n5226 DVDD.n489 0.0418115
R5832 DVDD.n640 DVDD.n608 0.0418115
R5833 DVDD.n852 DVDD.n708 0.0418115
R5834 DVDD.n4599 DVDD.n1013 0.0418115
R5835 DVDD.n5815 DVDD.n160 0.0414426
R5836 DVDD.n5171 DVDD.n471 0.0414426
R5837 DVDD.n4966 DVDD.n4947 0.0414426
R5838 DVDD.n796 DVDD.n747 0.0414426
R5839 DVDD.n4522 DVDD.n4505 0.0414426
R5840 DVDD.n2820 DVDD.n2819 0.0410978
R5841 DVDD.n5740 DVDD.n187 0.0410738
R5842 DVDD.n5241 DVDD.n566 0.0410738
R5843 DVDD.n5014 DVDD.n5013 0.0410738
R5844 DVDD.n4876 DVDD.n726 0.0410738
R5845 DVDD.n4614 DVDD.n1057 0.0410738
R5846 DVDD.n5832 DVDD.n146 0.0407049
R5847 DVDD.n5187 DVDD.n455 0.0407049
R5848 DVDD.n4950 DVDD.n678 0.0407049
R5849 DVDD.n813 DVDD.n812 0.0407049
R5850 DVDD.n1079 DVDD.n1074 0.0407049
R5851 DVDD.n5926 DVDD.n5925 0.0393914
R5852 DVDD.n5430 DVDD.n5429 0.0393914
R5853 DVDD.n5823 DVDD.n147 0.0384918
R5854 DVDD.n5179 DVDD.n457 0.0384918
R5855 DVDD.n4958 DVDD.n679 0.0384918
R5856 DVDD.n806 DVDD.n805 0.0384918
R5857 DVDD.n4514 DVDD.n1080 0.0384918
R5858 DVDD.n5748 DVDD.n186 0.038123
R5859 DVDD.n5234 DVDD.n565 0.038123
R5860 DVDD.n632 DVDD.n622 0.038123
R5861 DVDD.n860 DVDD.n725 0.038123
R5862 DVDD.n4607 DVDD.n1056 0.038123
R5863 DVDD.n2818 DVDD.n2096 0.03785
R5864 DVDD.n3363 DVDD.n3362 0.0377973
R5865 DVDD.n3265 DVDD.n3262 0.0377973
R5866 DVDD.n5807 DVDD.n159 0.0377541
R5867 DVDD.n5163 DVDD.n459 0.0377541
R5868 DVDD.n4974 DVDD.n681 0.0377541
R5869 DVDD.n787 DVDD.n749 0.0377541
R5870 DVDD.n4530 DVDD.n1082 0.0377541
R5871 DVDD.n5656 DVDD.n5655 0.0376798
R5872 DVDD.n5482 DVDD.n5481 0.0376798
R5873 DVDD.n5764 DVDD.n184 0.0373852
R5874 DVDD.n5218 DVDD.n490 0.0373852
R5875 DVDD.n648 DVDD.n620 0.0373852
R5876 DVDD.n844 DVDD.n709 0.0373852
R5877 DVDD.n4591 DVDD.n1014 0.0373852
R5878 DVDD.n1386 DVDD.n1307 0.0372431
R5879 DVDD.n1387 DVDD.n1311 0.0372431
R5880 DVDD.n1320 DVDD.n1219 0.0372431
R5881 DVDD.n1324 DVDD.n1221 0.0372431
R5882 DVDD.n154 DVDD.n142 0.0370164
R5883 DVDD.n473 DVDD.n461 0.0370164
R5884 DVDD.n4949 DVDD.n683 0.0370164
R5885 DVDD.n771 DVDD.n770 0.0370164
R5886 DVDD.n4507 DVDD.n1084 0.0370164
R5887 DVDD.n3357 DVDD.n3356 0.0369865
R5888 DVDD.n3388 DVDD.n3387 0.0369865
R5889 DVDD.n5775 DVDD.n182 0.0366475
R5890 DVDD.n5785 DVDD.n166 0.0366475
R5891 DVDD.n5845 DVDD.n135 0.0366475
R5892 DVDD.n5202 DVDD.n558 0.0366475
R5893 DVDD.n5196 DVDD.n556 0.0366475
R5894 DVDD.n5138 DVDD.n5137 0.0366475
R5895 DVDD.n664 DVDD.n618 0.0366475
R5896 DVDD.n5011 DVDD.n626 0.0366475
R5897 DVDD.n4992 DVDD.n424 0.0366475
R5898 DVDD.n828 DVDD.n718 0.0366475
R5899 DVDD.n822 DVDD.n716 0.0366475
R5900 DVDD.n758 DVDD.n400 0.0366475
R5901 DVDD.n4575 DVDD.n1049 0.0366475
R5902 DVDD.n4569 DVDD.n1047 0.0366475
R5903 DVDD.n4548 DVDD.n377 0.0366475
R5904 DVDD.n5770 DVDD.n171 0.0359098
R5905 DVDD.n5212 DVDD.n492 0.0359098
R5906 DVDD.n654 DVDD.n607 0.0359098
R5907 DVDD.n838 DVDD.n711 0.0359098
R5908 DVDD.n4585 DVDD.n1016 0.0359098
R5909 DVDD.n5801 DVDD.n157 0.035541
R5910 DVDD.n5157 DVDD.n472 0.035541
R5911 DVDD.n4980 DVDD.n4948 0.035541
R5912 DVDD.n780 DVDD.n779 0.035541
R5913 DVDD.n4536 DVDD.n4506 0.035541
R5914 DVDD.n3351 DVDD.n3350 0.0353649
R5915 DVDD.n3397 DVDD.n3223 0.0353649
R5916 DVDD.n5754 DVDD.n188 0.0351721
R5917 DVDD.n5228 DVDD.n563 0.0351721
R5918 DVDD.n638 DVDD.n623 0.0351721
R5919 DVDD.n854 DVDD.n723 0.0351721
R5920 DVDD.n4601 DVDD.n1054 0.0351721
R5921 DVDD.n5729 DVDD.n198 0.0348033
R5922 DVDD.n5817 DVDD.n149 0.0348033
R5923 DVDD.n5093 DVDD.n5092 0.0348033
R5924 DVDD.n5173 DVDD.n454 0.0348033
R5925 DVDD.n597 DVDD.n593 0.0348033
R5926 DVDD.n4964 DVDD.n677 0.0348033
R5927 DVDD.n876 DVDD.n735 0.0348033
R5928 DVDD.n798 DVDD.n797 0.0348033
R5929 DVDD.n1059 DVDD.n892 0.0348033
R5930 DVDD.n4520 DVDD.n1078 0.0348033
R5931 DVDD.n3367 DVDD.n3366 0.0345541
R5932 DVDD.n3258 DVDD.n3243 0.0345541
R5933 DVDD.n3328 DVDD.n3275 0.0344013
R5934 DVDD.n3369 DVDD.n3271 0.0344013
R5935 DVDD.n3374 DVDD.n3373 0.0344013
R5936 DVDD.n3371 DVDD.n3249 0.0344013
R5937 DVDD.n5833 DVDD.n164 0.0340656
R5938 DVDD.n5189 DVDD.n469 0.0340656
R5939 DVDD.n4945 DVDD.n673 0.0340656
R5940 DVDD.n815 DVDD.n814 0.0340656
R5941 DVDD.n4562 DVDD.n4561 0.0340656
R5942 DVDD.n1392 DVDD.n1309 0.0330202
R5943 DVDD.n1222 DVDD.n1214 0.0330202
R5944 DVDD.n5511 DVDD.n5510 0.0325451
R5945 DVDD.n4704 DVDD.n949 0.0325451
R5946 DVDD.n5731 DVDD.n198 0.0324979
R5947 DVDD.n5093 DVDD.n5087 0.0324979
R5948 DVDD.n596 DVDD.n593 0.0324979
R5949 DVDD.n878 DVDD.n735 0.0324979
R5950 DVDD.n896 DVDD.n892 0.0324979
R5951 DVDD.n1912 DVDD.n1909 0.03245
R5952 DVDD.n1913 DVDD.n1912 0.03245
R5953 DVDD.n3285 DVDD.n3284 0.03245
R5954 DVDD.n3291 DVDD.n3285 0.03245
R5955 DVDD.n3291 DVDD.n3290 0.03245
R5956 DVDD.n1911 DVDD.n1910 0.03245
R5957 DVDD.n1911 DVDD.n1907 0.03245
R5958 DVDD.n2192 DVDD.n2173 0.03245
R5959 DVDD.n2185 DVDD.n2173 0.03245
R5960 DVDD.n2185 DVDD.n2184 0.03245
R5961 DVDD.n2184 DVDD.n1895 0.03245
R5962 DVDD.n3710 DVDD.n1895 0.03245
R5963 DVDD.n3711 DVDD.n3710 0.03245
R5964 DVDD.n3712 DVDD.n3711 0.03245
R5965 DVDD.n3712 DVDD.n1888 0.03245
R5966 DVDD.n3719 DVDD.n1888 0.03245
R5967 DVDD.n3773 DVDD.n3753 0.03245
R5968 DVDD.n3761 DVDD.n3753 0.03245
R5969 DVDD.n3766 DVDD.n3761 0.03245
R5970 DVDD.n3766 DVDD.n3765 0.03245
R5971 DVDD.n3765 DVDD.n1664 0.03245
R5972 DVDD.n4290 DVDD.n1664 0.03245
R5973 DVDD.n4291 DVDD.n4290 0.03245
R5974 DVDD.n4291 DVDD.n1658 0.03245
R5975 DVDD.n4299 DVDD.n1658 0.03245
R5976 DVDD.n5735 DVDD.n193 0.0318525
R5977 DVDD.n5821 DVDD.n162 0.0318525
R5978 DVDD.n5095 DVDD.n569 0.0318525
R5979 DVDD.n5177 DVDD.n467 0.0318525
R5980 DVDD.n5019 DVDD.n594 0.0318525
R5981 DVDD.n4960 DVDD.n4943 0.0318525
R5982 DVDD.n872 DVDD.n737 0.0318525
R5983 DVDD.n804 DVDD.n803 0.0318525
R5984 DVDD.n1063 DVDD.n894 0.0318525
R5985 DVDD.n4516 DVDD.n4502 0.0318525
R5986 DVDD.n5847 DVDD.n135 0.0315574
R5987 DVDD.n5137 DVDD.n5136 0.0315574
R5988 DVDD.n428 DVDD.n424 0.0315574
R5989 DVDD.n404 DVDD.n400 0.0315574
R5990 DVDD.n381 DVDD.n377 0.0315574
R5991 DVDD.n5750 DVDD.n175 0.0314836
R5992 DVDD.n5232 DVDD.n487 0.0314836
R5993 DVDD.n634 DVDD.n611 0.0314836
R5994 DVDD.n858 DVDD.n706 0.0314836
R5995 DVDD.n4605 DVDD.n1011 0.0314836
R5996 DVDD.n5805 DVDD.n151 0.0311148
R5997 DVDD.n5161 DVDD.n465 0.0311148
R5998 DVDD.n4976 DVDD.n4941 0.0311148
R5999 DVDD.n786 DVDD.n785 0.0311148
R6000 DVDD.n4532 DVDD.n4500 0.0311148
R6001 DVDD.n2807 DVDD.n2700 0.0308261
R6002 DVDD.n2808 DVDD.n2807 0.0308261
R6003 DVDD.n2809 DVDD.n2808 0.0308261
R6004 DVDD.n2809 DVDD.n2698 0.0308261
R6005 DVDD.n2813 DVDD.n2698 0.0308261
R6006 DVDD.n2814 DVDD.n2813 0.0308261
R6007 DVDD.n2815 DVDD.n2814 0.0308261
R6008 DVDD.n2815 DVDD.n2696 0.0308261
R6009 DVDD.n2819 DVDD.n2696 0.0308261
R6010 DVDD.n2800 DVDD.n2702 0.0308261
R6011 DVDD.n5766 DVDD.n177 0.0307459
R6012 DVDD.n5216 DVDD.n561 0.0307459
R6013 DVDD.n650 DVDD.n613 0.0307459
R6014 DVDD.n842 DVDD.n721 0.0307459
R6015 DVDD.n4589 DVDD.n1052 0.0307459
R6016 DVDD.n5494 DVDD.n256 0.0305
R6017 DVDD.n5498 DVDD.n5497 0.0305
R6018 DVDD.n5493 DVDD.n5492 0.0305
R6019 DVDD.n5490 DVDD.n5489 0.0305
R6020 DVDD.n5836 DVDD.n5835 0.030377
R6021 DVDD.n5317 DVDD.n474 0.030377
R6022 DVDD.n5003 DVDD.n5002 0.030377
R6023 DVDD.n769 DVDD.n768 0.030377
R6024 DVDD.n4559 DVDD.n4558 0.030377
R6025 DVDD.n5773 DVDD.n179 0.0300082
R6026 DVDD.n5784 DVDD.n168 0.0300082
R6027 DVDD.n5843 DVDD.n138 0.0300082
R6028 DVDD.n5200 DVDD.n494 0.0300082
R6029 DVDD.n5198 DVDD.n495 0.0300082
R6030 DVDD.n5140 DVDD.n5139 0.0300082
R6031 DVDD.n666 DVDD.n615 0.0300082
R6032 DVDD.n668 DVDD.n606 0.0300082
R6033 DVDD.n4994 DVDD.n427 0.0300082
R6034 DVDD.n826 DVDD.n713 0.0300082
R6035 DVDD.n824 DVDD.n714 0.0300082
R6036 DVDD.n760 DVDD.n403 0.0300082
R6037 DVDD.n4573 DVDD.n1018 0.0300082
R6038 DVDD.n4571 DVDD.n1019 0.0300082
R6039 DVDD.n4550 DVDD.n380 0.0300082
R6040 DVDD.n1381 DVDD.n1312 0.0298119
R6041 DVDD.n1381 DVDD.n1308 0.0298119
R6042 DVDD.n1317 DVDD.n1217 0.0298119
R6043 DVDD.n1317 DVDD.n1215 0.0298119
R6044 DVDD.n5768 DVDD.n189 0.0292705
R6045 DVDD.n5214 DVDD.n560 0.0292705
R6046 DVDD.n652 DVDD.n624 0.0292705
R6047 DVDD.n840 DVDD.n720 0.0292705
R6048 DVDD.n4587 DVDD.n1051 0.0292705
R6049 DVDD.n937 DVDD.n936 0.0292629
R6050 DVDD.n956 DVDD.n955 0.0292629
R6051 DVDD.n5672 DVDD.n242 0.0292629
R6052 DVDD.n250 DVDD.n249 0.0292629
R6053 DVDD.n3297 DVDD.n3275 0.0291547
R6054 DVDD.n3360 DVDD.n3297 0.0291547
R6055 DVDD.n3360 DVDD.n3359 0.0291547
R6056 DVDD.n3359 DVDD.n3298 0.0291547
R6057 DVDD.n3369 DVDD.n3272 0.0291547
R6058 DVDD.n3294 DVDD.n3272 0.0291547
R6059 DVDD.n3299 DVDD.n3294 0.0291547
R6060 DVDD.n3340 DVDD.n3299 0.0291547
R6061 DVDD.n3373 DVDD.n3246 0.0291547
R6062 DVDD.n3260 DVDD.n3246 0.0291547
R6063 DVDD.n3260 DVDD.n3232 0.0291547
R6064 DVDD.n3232 DVDD.n3231 0.0291547
R6065 DVDD.n3371 DVDD.n3268 0.0291547
R6066 DVDD.n3268 DVDD.n3227 0.0291547
R6067 DVDD.n3390 DVDD.n3227 0.0291547
R6068 DVDD.n3391 DVDD.n3390 0.0291547
R6069 DVDD.n111 DVDD.n99 0.0290309
R6070 DVDD.n102 DVDD.n95 0.0290309
R6071 DVDD.n5407 DVDD.n338 0.0290309
R6072 DVDD.n349 DVDD.n342 0.0290309
R6073 DVDD.n940 DVDD.n916 0.0290309
R6074 DVDD.n958 DVDD.n923 0.0290309
R6075 DVDD.n5703 DVDD.n240 0.0290309
R6076 DVDD.n246 DVDD.n229 0.0290309
R6077 DVDD.n5803 DVDD.n152 0.0289016
R6078 DVDD.n5159 DVDD.n453 0.0289016
R6079 DVDD.n4978 DVDD.n676 0.0289016
R6080 DVDD.n783 DVDD.n751 0.0289016
R6081 DVDD.n4534 DVDD.n1077 0.0289016
R6082 DVDD.n5752 DVDD.n173 0.0285328
R6083 DVDD.n5230 DVDD.n488 0.0285328
R6084 DVDD.n636 DVDD.n609 0.0285328
R6085 DVDD.n856 DVDD.n707 0.0285328
R6086 DVDD.n4603 DVDD.n1012 0.0285328
R6087 DVDD.n2805 DVDD.n2804 0.0284
R6088 DVDD.n2806 DVDD.n2805 0.0284
R6089 DVDD.n2806 DVDD.n2699 0.0284
R6090 DVDD.n2810 DVDD.n2699 0.0284
R6091 DVDD.n2811 DVDD.n2810 0.0284
R6092 DVDD.n2812 DVDD.n2811 0.0284
R6093 DVDD.n2812 DVDD.n2697 0.0284
R6094 DVDD.n2816 DVDD.n2697 0.0284
R6095 DVDD.n2817 DVDD.n2816 0.0284
R6096 DVDD.n2818 DVDD.n2817 0.0284
R6097 DVDD.n5728 DVDD.n195 0.0281639
R6098 DVDD.n5819 DVDD.n161 0.0281639
R6099 DVDD.n5089 DVDD.n573 0.0281639
R6100 DVDD.n5175 DVDD.n470 0.0281639
R6101 DVDD.n599 DVDD.n590 0.0281639
R6102 DVDD.n4962 DVDD.n4946 0.0281639
R6103 DVDD.n874 DVDD.n738 0.0281639
R6104 DVDD.n800 DVDD.n799 0.0281639
R6105 DVDD.n1061 DVDD.n895 0.0281639
R6106 DVDD.n4518 DVDD.n4504 0.0281639
R6107 DVDD.n5496 DVDD.n5495 0.0277727
R6108 DVDD.n5491 DVDD.n262 0.0277727
R6109 DVDD.n5790 DVDD.n145 0.0274262
R6110 DVDD.n5192 DVDD.n456 0.0274262
R6111 DVDD.n5006 DVDD.n5005 0.0274262
R6112 DVDD.n818 DVDD.n740 0.0274262
R6113 DVDD.n4565 DVDD.n1071 0.0274262
R6114 DVDD.n1914 DVDD.n1913 0.027126
R6115 DVDD.n1393 DVDD.n1392 0.0270348
R6116 DVDD.n1555 DVDD.n1222 0.0270348
R6117 DVDD.n3593 DVDD.n3124 0.026913
R6118 DVDD.n3593 DVDD.n3592 0.026913
R6119 DVDD.n3592 DVDD.n3591 0.026913
R6120 DVDD.n3591 DVDD.n3125 0.026913
R6121 DVDD.n3136 DVDD.n3125 0.026913
R6122 DVDD.n3137 DVDD.n3136 0.026913
R6123 DVDD.n3580 DVDD.n3137 0.026913
R6124 DVDD.n3580 DVDD.n3579 0.026913
R6125 DVDD.n3579 DVDD.n3139 0.026913
R6126 DVDD.n3552 DVDD.n3139 0.026913
R6127 DVDD.n3555 DVDD.n3552 0.026913
R6128 DVDD.n3594 DVDD.n3122 0.026913
R6129 DVDD.n3582 DVDD.n3135 0.026913
R6130 DVDD.n3582 DVDD.n3581 0.026913
R6131 DVDD.n3553 DVDD.n3140 0.026913
R6132 DVDD.n3554 DVDD.n3553 0.026913
R6133 DVDD.n3434 DVDD.n3208 0.026913
R6134 DVDD.n3445 DVDD.n3206 0.026913
R6135 DVDD.n3445 DVDD.n3196 0.026913
R6136 DVDD.n3470 DVDD.n3469 0.026913
R6137 DVDD.n3471 DVDD.n3470 0.026913
R6138 DVDD.n3416 DVDD.n3209 0.026913
R6139 DVDD.n3123 DVDD.n3111 0.026913
R6140 DVDD.n3432 DVDD.n3431 0.026913
R6141 DVDD.n3433 DVDD.n3432 0.026913
R6142 DVDD.n3433 DVDD.n3207 0.026913
R6143 DVDD.n3442 DVDD.n3207 0.026913
R6144 DVDD.n3443 DVDD.n3442 0.026913
R6145 DVDD.n3444 DVDD.n3443 0.026913
R6146 DVDD.n3444 DVDD.n3195 0.026913
R6147 DVDD.n3467 DVDD.n3195 0.026913
R6148 DVDD.n3468 DVDD.n3467 0.026913
R6149 DVDD.n3468 DVDD.n3193 0.026913
R6150 DVDD.n3472 DVDD.n3193 0.026913
R6151 DVDD.n3475 DVDD.n3184 0.026913
R6152 DVDD.n3479 DVDD.n3478 0.026913
R6153 DVDD.n3487 DVDD.n3486 0.026913
R6154 DVDD.n3495 DVDD.n3494 0.026913
R6155 DVDD.n3503 DVDD.n3502 0.026913
R6156 DVDD.n3508 DVDD.n3170 0.026913
R6157 DVDD.n3476 DVDD.n3474 0.026913
R6158 DVDD.n3480 DVDD.n3477 0.026913
R6159 DVDD.n3482 DVDD.n3480 0.026913
R6160 DVDD.n3484 DVDD.n3482 0.026913
R6161 DVDD.n3485 DVDD.n3484 0.026913
R6162 DVDD.n3488 DVDD.n3485 0.026913
R6163 DVDD.n3490 DVDD.n3488 0.026913
R6164 DVDD.n3492 DVDD.n3490 0.026913
R6165 DVDD.n3493 DVDD.n3492 0.026913
R6166 DVDD.n3496 DVDD.n3493 0.026913
R6167 DVDD.n3498 DVDD.n3496 0.026913
R6168 DVDD.n3500 DVDD.n3498 0.026913
R6169 DVDD.n3501 DVDD.n3500 0.026913
R6170 DVDD.n3504 DVDD.n3501 0.026913
R6171 DVDD.n3506 DVDD.n3504 0.026913
R6172 DVDD.n3507 DVDD.n3506 0.026913
R6173 DVDD.n3510 DVDD.n3507 0.026913
R6174 DVDD.n3510 DVDD.n3509 0.026913
R6175 DVDD.n3509 DVDD.n3169 0.026913
R6176 DVDD.n3515 DVDD.n3169 0.026913
R6177 DVDD.n3517 DVDD.n3516 0.026913
R6178 DVDD.n3520 DVDD.n3517 0.026913
R6179 DVDD.n3522 DVDD.n3520 0.026913
R6180 DVDD.n3524 DVDD.n3522 0.026913
R6181 DVDD.n3526 DVDD.n3524 0.026913
R6182 DVDD.n3527 DVDD.n3526 0.026913
R6183 DVDD.n3530 DVDD.n3527 0.026913
R6184 DVDD.n3532 DVDD.n3530 0.026913
R6185 DVDD.n3534 DVDD.n3532 0.026913
R6186 DVDD.n3535 DVDD.n3534 0.026913
R6187 DVDD.n3538 DVDD.n3535 0.026913
R6188 DVDD.n3540 DVDD.n3538 0.026913
R6189 DVDD.n3542 DVDD.n3540 0.026913
R6190 DVDD.n3543 DVDD.n3542 0.026913
R6191 DVDD.n3546 DVDD.n3543 0.026913
R6192 DVDD.n3548 DVDD.n3546 0.026913
R6193 DVDD.n3550 DVDD.n3548 0.026913
R6194 DVDD.n3551 DVDD.n3550 0.026913
R6195 DVDD.n3559 DVDD.n3557 0.026913
R6196 DVDD.n3519 DVDD.n3518 0.026913
R6197 DVDD.n3529 DVDD.n3528 0.026913
R6198 DVDD.n3537 DVDD.n3536 0.026913
R6199 DVDD.n3545 DVDD.n3544 0.026913
R6200 DVDD.n3561 DVDD.n3168 0.026913
R6201 DVDD.n3558 DVDD.n3160 0.026913
R6202 DVDD.n2821 DVDD.n2820 0.026913
R6203 DVDD.n2822 DVDD.n2821 0.026913
R6204 DVDD.n2825 DVDD.n2822 0.026913
R6205 DVDD.n2827 DVDD.n2825 0.026913
R6206 DVDD.n2829 DVDD.n2827 0.026913
R6207 DVDD.n2831 DVDD.n2829 0.026913
R6208 DVDD.n2832 DVDD.n2831 0.026913
R6209 DVDD.n2835 DVDD.n2832 0.026913
R6210 DVDD.n2837 DVDD.n2835 0.026913
R6211 DVDD.n2861 DVDD.n2693 0.026913
R6212 DVDD.n2861 DVDD.n2860 0.026913
R6213 DVDD.n2860 DVDD.n2858 0.026913
R6214 DVDD.n2858 DVDD.n2855 0.026913
R6215 DVDD.n2855 DVDD.n2854 0.026913
R6216 DVDD.n2854 DVDD.n2852 0.026913
R6217 DVDD.n2852 DVDD.n2850 0.026913
R6218 DVDD.n2850 DVDD.n2847 0.026913
R6219 DVDD.n2847 DVDD.n2846 0.026913
R6220 DVDD.n2803 DVDD.n2703 0.026913
R6221 DVDD.n2857 DVDD.n2856 0.026913
R6222 DVDD.n2849 DVDD.n2848 0.026913
R6223 DVDD.n1385 DVDD.n1384 0.0264516
R6224 DVDD.n1322 DVDD.n1319 0.0264516
R6225 DVDD.n1321 DVDD.n1319 0.0264516
R6226 DVDD.n1384 DVDD.n1383 0.0264516
R6227 DVDD.n3263 DVDD.n3242 0.0264459
R6228 DVDD.n3365 DVDD.n3278 0.0264459
R6229 DVDD DVDD.n3551 0.0264239
R6230 DVDD.n2695 DVDD.n2683 0.0264239
R6231 DVDD.n3505 DVDD.n3191 0.0261793
R6232 DVDD.n3511 DVDD.n3174 0.0261793
R6233 DVDD.n3521 DVDD.n3156 0.0261793
R6234 DVDD.n3525 DVDD.n3163 0.0261793
R6235 DVDD.n2845 DVDD.n2691 0.0259348
R6236 DVDD.n1998 DVDD.n1984 0.025745
R6237 DVDD.n3386 DVDD.n3225 0.0256351
R6238 DVDD.n3355 DVDD.n3354 0.0256351
R6239 DVDD.n3092 DVDD.n2023 0.0255952
R6240 DVDD.n3590 DVDD.n3126 0.0254457
R6241 DVDD.n3436 DVDD.n3435 0.0254457
R6242 DVDD.n5910 DVDD.n91 0.0253196
R6243 DVDD.n114 DVDD.n93 0.0253196
R6244 DVDD.n5413 DVDD.n345 0.0253196
R6245 DVDD.n5410 DVDD.n347 0.0253196
R6246 DVDD.n933 DVDD.n926 0.0253196
R6247 DVDD.n952 DVDD.n919 0.0253196
R6248 DVDD.n5668 DVDD.n232 0.0253196
R6249 DVDD.n252 DVDD.n238 0.0253196
R6250 DVDD.n5734 DVDD.n195 0.0252131
R6251 DVDD.n5819 DVDD.n148 0.0252131
R6252 DVDD.n5089 DVDD.n5086 0.0252131
R6253 DVDD.n5175 DVDD.n458 0.0252131
R6254 DVDD.n599 DVDD.n592 0.0252131
R6255 DVDD.n4962 DVDD.n680 0.0252131
R6256 DVDD.n874 DVDD.n736 0.0252131
R6257 DVDD.n800 DVDD.n745 0.0252131
R6258 DVDD.n1061 DVDD.n893 0.0252131
R6259 DVDD.n4518 DVDD.n1081 0.0252131
R6260 DVDD.n3347 DVDD.n3298 0.024917
R6261 DVDD.n3345 DVDD.n3340 0.024917
R6262 DVDD.n3231 DVDD.n3222 0.024917
R6263 DVDD.n3392 DVDD.n3391 0.024917
R6264 DVDD.n5911 DVDD.n89 0.0248557
R6265 DVDD.n109 DVDD.n94 0.0248557
R6266 DVDD.n5414 DVDD.n343 0.0248557
R6267 DVDD.n5417 DVDD.n352 0.0248557
R6268 DVDD.n941 DVDD.n927 0.0248557
R6269 DVDD.n942 DVDD.n920 0.0248557
R6270 DVDD.n257 DVDD.n233 0.0248557
R6271 DVDD.n244 DVDD.n239 0.0248557
R6272 DVDD.n5752 DVDD.n185 0.0248443
R6273 DVDD.n5230 DVDD.n564 0.0248443
R6274 DVDD.n636 DVDD.n621 0.0248443
R6275 DVDD.n856 DVDD.n724 0.0248443
R6276 DVDD.n4603 DVDD.n1055 0.0248443
R6277 DVDD.n2824 DVDD.n2823 0.0248
R6278 DVDD.n2834 DVDD.n2833 0.0248
R6279 DVDD.n3370 DVDD.n3270 0.0248
R6280 DVDD.n3283 DVDD.n3282 0.0248
R6281 DVDD.n3293 DVDD.n3292 0.0248
R6282 DVDD.n3289 DVDD.n3228 0.0248
R6283 DVDD.n1998 DVDD.n1985 0.0247619
R6284 DVDD.n3091 DVDD.n2023 0.0247609
R6285 DVDD.n2707 DVDD 0.0247148
R6286 DVDD.n3497 DVDD.n3177 0.024712
R6287 DVDD.n3533 DVDD.n3153 0.024712
R6288 DVDD.n5803 DVDD.n158 0.0244754
R6289 DVDD.n5159 DVDD.n460 0.0244754
R6290 DVDD.n4978 DVDD.n682 0.0244754
R6291 DVDD.n784 DVDD.n783 0.0244754
R6292 DVDD.n4534 DVDD.n1083 0.0244754
R6293 DVDD.n2853 DVDD.n2686 0.0244674
R6294 DVDD.n2826 DVDD.n2093 0.02435
R6295 DVDD.n5768 DVDD.n183 0.0241066
R6296 DVDD.n5214 DVDD.n491 0.0241066
R6297 DVDD.n652 DVDD.n619 0.0241066
R6298 DVDD.n840 DVDD.n710 0.0241066
R6299 DVDD.n4587 DVDD.n1015 0.0241066
R6300 DVDD.n3366 DVDD.n3277 0.0240135
R6301 DVDD.n3266 DVDD.n3258 0.0240135
R6302 DVDD.n1370 DVDD.n1329 0.024
R6303 DVDD.n3602 DVDD.n3113 0.0239783
R6304 DVDD.n3418 DVDD.n3417 0.0239783
R6305 DVDD.n2830 DVDD.n2090 0.0239
R6306 DVDD.n2217 DVDD 0.0238333
R6307 DVDD.n2216 DVDD 0.0238333
R6308 DVDD.n2221 DVDD 0.0238333
R6309 DVDD.n2220 DVDD 0.0238333
R6310 DVDD.n2225 DVDD 0.0238333
R6311 DVDD.n2224 DVDD 0.0238333
R6312 DVDD.n2229 DVDD 0.0238333
R6313 DVDD.n2228 DVDD 0.0238333
R6314 DVDD.n2233 DVDD 0.0238333
R6315 DVDD.n2232 DVDD 0.0238333
R6316 DVDD.n2237 DVDD 0.0238333
R6317 DVDD.n2236 DVDD 0.0238333
R6318 DVDD DVDD.n2239 0.0238333
R6319 DVDD.n5839 DVDD.n140 0.0237377
R6320 DVDD.n5145 DVDD.n463 0.0237377
R6321 DVDD.n4999 DVDD.n4939 0.0237377
R6322 DVDD.n765 DVDD.n756 0.0237377
R6323 DVDD.n4555 DVDD.n4498 0.0237377
R6324 DVDD.n5773 DVDD.n181 0.0233689
R6325 DVDD.n181 DVDD.n168 0.0233689
R6326 DVDD.n5841 DVDD.n136 0.0233689
R6327 DVDD.n5843 DVDD.n136 0.0233689
R6328 DVDD.n5200 DVDD.n557 0.0233689
R6329 DVDD.n5198 DVDD.n557 0.0233689
R6330 DVDD.n5143 DVDD.n5102 0.0233689
R6331 DVDD.n5140 DVDD.n5102 0.0233689
R6332 DVDD.n666 DVDD.n617 0.0233689
R6333 DVDD.n668 DVDD.n617 0.0233689
R6334 DVDD.n4997 DVDD.n425 0.0233689
R6335 DVDD.n4994 DVDD.n425 0.0233689
R6336 DVDD.n826 DVDD.n717 0.0233689
R6337 DVDD.n824 DVDD.n717 0.0233689
R6338 DVDD.n763 DVDD.n401 0.0233689
R6339 DVDD.n760 DVDD.n401 0.0233689
R6340 DVDD.n4573 DVDD.n1048 0.0233689
R6341 DVDD.n4571 DVDD.n1048 0.0233689
R6342 DVDD.n4553 DVDD.n378 0.0233689
R6343 DVDD.n4550 DVDD.n378 0.0233689
R6344 DVDD.n3489 DVDD.n3188 0.0232446
R6345 DVDD.n3541 DVDD.n3166 0.0232446
R6346 DVDD.n3350 DVDD.n3309 0.0232027
R6347 DVDD.n3234 DVDD.n3223 0.0232027
R6348 DVDD.n5836 DVDD.n140 0.023
R6349 DVDD.n474 DVDD.n463 0.023
R6350 DVDD.n5002 DVDD.n4939 0.023
R6351 DVDD.n768 DVDD.n756 0.023
R6352 DVDD.n4558 DVDD.n4498 0.023
R6353 DVDD.n2863 DVDD.n2862 0.023
R6354 DVDD.n1741 DVDD.n1739 0.0229381
R6355 DVDD.n1998 DVDD.n1997 0.0227712
R6356 DVDD.n1899 DVDD.n1897 0.0227688
R6357 DVDD.n2025 DVDD.n2023 0.0227678
R6358 DVDD.n5766 DVDD.n183 0.0226311
R6359 DVDD.n5216 DVDD.n491 0.0226311
R6360 DVDD.n650 DVDD.n619 0.0226311
R6361 DVDD.n842 DVDD.n710 0.0226311
R6362 DVDD.n4589 DVDD.n1015 0.0226311
R6363 DVDD.n3473 DVDD.n3182 0.0225217
R6364 DVDD.n3556 DVDD.n3157 0.0225217
R6365 DVDD.n5848 DVDD.n5847 0.0224209
R6366 DVDD.n5136 DVDD.n5135 0.0224209
R6367 DVDD.n5339 DVDD.n428 0.0224209
R6368 DVDD.n5360 DVDD.n404 0.0224209
R6369 DVDD.n5380 DVDD.n381 0.0224209
R6370 DVDD.n3225 DVDD.n3224 0.0223919
R6371 DVDD.n3395 DVDD.n3225 0.0223919
R6372 DVDD.n3354 DVDD.n3349 0.0223919
R6373 DVDD.n3354 DVDD.n3353 0.0223919
R6374 DVDD.n1742 DVDD 0.0223846
R6375 DVDD.n1386 DVDD.n1312 0.0223807
R6376 DVDD.n1387 DVDD.n1308 0.0223807
R6377 DVDD.n1320 DVDD.n1217 0.0223807
R6378 DVDD.n1324 DVDD.n1215 0.0223807
R6379 DVDD.n3483 DVDD.n3179 0.0222663
R6380 DVDD.n3547 DVDD.n3151 0.0222663
R6381 DVDD.n5805 DVDD.n158 0.0222623
R6382 DVDD.n5161 DVDD.n460 0.0222623
R6383 DVDD.n4976 DVDD.n682 0.0222623
R6384 DVDD.n785 DVDD.n784 0.0222623
R6385 DVDD.n4532 DVDD.n1083 0.0222623
R6386 DVDD.n5750 DVDD.n185 0.0218934
R6387 DVDD.n5232 DVDD.n564 0.0218934
R6388 DVDD.n634 DVDD.n621 0.0218934
R6389 DVDD.n858 DVDD.n724 0.0218934
R6390 DVDD.n4605 DVDD.n1055 0.0218934
R6391 DVDD.n1908 DVDD.n1903 0.0218
R6392 DVDD.n3287 DVDD.n3286 0.0218
R6393 DVDD.n3288 DVDD.n3287 0.0218
R6394 DVDD.n3481 DVDD.n3180 0.0217772
R6395 DVDD.n3549 DVDD.n3150 0.0217772
R6396 DVDD.n3356 DVDD.n3309 0.0215811
R6397 DVDD.n3387 DVDD.n3234 0.0215811
R6398 DVDD.n5735 DVDD.n5734 0.0215246
R6399 DVDD.n5821 DVDD.n148 0.0215246
R6400 DVDD.n5086 DVDD.n569 0.0215246
R6401 DVDD.n5177 DVDD.n458 0.0215246
R6402 DVDD.n594 DVDD.n592 0.0215246
R6403 DVDD.n4960 DVDD.n680 0.0215246
R6404 DVDD.n872 DVDD.n736 0.0215246
R6405 DVDD.n803 DVDD.n745 0.0215246
R6406 DVDD.n1063 DVDD.n893 0.0215246
R6407 DVDD.n4516 DVDD.n1081 0.0215246
R6408 DVDD.n5732 DVDD.n5731 0.0215141
R6409 DVDD.n5087 DVDD.n572 0.0215141
R6410 DVDD.n596 DVDD.n589 0.0215141
R6411 DVDD.n4772 DVDD.n878 0.0215141
R6412 DVDD.n4743 DVDD.n896 0.0215141
R6413 DVDD.n112 DVDD.n97 0.0211443
R6414 DVDD.n5908 DVDD.n96 0.0211443
R6415 DVDD.n5408 DVDD.n336 0.0211443
R6416 DVDD.n5411 DVDD.n335 0.0211443
R6417 DVDD.n931 DVDD.n917 0.0211443
R6418 DVDD.n950 DVDD.n924 0.0211443
R6419 DVDD.n5666 DVDD.n236 0.0211443
R6420 DVDD.n254 DVDD.n230 0.0211443
R6421 DVDD.n2859 DVDD.n2689 0.0210435
R6422 DVDD.n3648 DVDD 0.020979
R6423 DVDD.n5953 DVDD.n28 0.0209627
R6424 DVDD.n4700 DVDD.n4699 0.0209627
R6425 DVDD.n3491 DVDD.n3189 0.0207989
R6426 DVDD.n3539 DVDD.n3165 0.0207989
R6427 DVDD.n3363 DVDD.n3277 0.0207703
R6428 DVDD.n3266 DVDD.n3265 0.0207703
R6429 DVDD.n110 DVDD.n100 0.0206804
R6430 DVDD.n5914 DVDD.n5913 0.0206804
R6431 DVDD.n5406 DVDD.n339 0.0206804
R6432 DVDD.n5416 DVDD.n341 0.0206804
R6433 DVDD.n1886 DVDD.n1861 0.020525
R6434 DVDD.n1900 DVDD 0.0204408
R6435 DVDD.n2024 DVDD 0.0202739
R6436 DVDD.n3640 DVDD.n3639 0.0201875
R6437 DVDD.n3641 DVDD.n3640 0.0201875
R6438 DVDD.n3641 DVDD.n1981 0.0201875
R6439 DVDD.n3655 DVDD.n1981 0.0201875
R6440 DVDD.n3656 DVDD.n3655 0.0201875
R6441 DVDD.n3666 DVDD.n3656 0.0201875
R6442 DVDD.n3666 DVDD.n3665 0.0201875
R6443 DVDD.n3595 DVDD.n3121 0.0200652
R6444 DVDD.n3430 DVDD.n3429 0.0200652
R6445 DVDD.n5615 DVDD.n5614 0.0197083
R6446 DVDD.n5515 DVDD.n30 0.0197083
R6447 DVDD.n5531 DVDD.n5530 0.0197083
R6448 DVDD.n5548 DVDD.n5547 0.0197083
R6449 DVDD.n4654 DVDD.n973 0.0197083
R6450 DVDD.n4683 DVDD.n4682 0.0197083
R6451 DVDD.n4666 DVDD.n4665 0.0197083
R6452 DVDD.n5440 DVDD.n5439 0.0197083
R6453 DVDD.n2851 DVDD.n2685 0.0195761
R6454 DVDD.n5648 DVDD.n5609 0.0193985
R6455 DVDD.n317 DVDD.n293 0.0193985
R6456 DVDD.n3499 DVDD.n3176 0.0193315
R6457 DVDD.n3531 DVDD.n3154 0.0193315
R6458 DVDD.n164 DVDD.n145 0.0193115
R6459 DVDD.n5189 DVDD.n456 0.0193115
R6460 DVDD.n5005 DVDD.n673 0.0193115
R6461 DVDD.n815 DVDD.n740 0.0193115
R6462 DVDD.n4562 DVDD.n1071 0.0193115
R6463 DVDD.n5644 DVDD.n50 0.0192435
R6464 DVDD.n5471 DVDD.n5470 0.0192435
R6465 DVDD.n5517 DVDD.n27 0.0190886
R6466 DVDD.n4697 DVDD.n4696 0.0190886
R6467 DVDD.n5627 DVDD.n63 0.0189337
R6468 DVDD.n5452 DVDD.n302 0.0189337
R6469 DVDD.n5533 DVDD.n12 0.0187788
R6470 DVDD.n4679 DVDD.n979 0.0187788
R6471 DVDD.n1339 DVDD.n1338 0.0186803
R6472 DVDD.n1341 DVDD.n1335 0.0186803
R6473 DVDD.n1335 DVDD.n1334 0.0186803
R6474 DVDD.n1332 DVDD.n1330 0.0186803
R6475 DVDD.n1365 DVDD.n1333 0.0186803
R6476 DVDD.n1367 DVDD.n1366 0.0186803
R6477 DVDD.n1334 DVDD.n1329 0.0186803
R6478 DVDD.n1366 DVDD.n1365 0.0186803
R6479 DVDD.n1369 DVDD.n1330 0.0186803
R6480 DVDD.n1341 DVDD.n1339 0.0186803
R6481 DVDD.n1338 DVDD.n1336 0.0186803
R6482 DVDD.n1333 DVDD.n1332 0.0186803
R6483 DVDD.n5611 DVDD.n57 0.0186239
R6484 DVDD.n5436 DVDD.n309 0.0186239
R6485 DVDD.n3134 DVDD.n3127 0.0185978
R6486 DVDD.n3578 DVDD.n3138 0.0185978
R6487 DVDD.n3441 DVDD.n3440 0.0185978
R6488 DVDD.n3466 DVDD.n3465 0.0185978
R6489 DVDD.n5729 DVDD.n5728 0.0185738
R6490 DVDD.n5817 DVDD.n161 0.0185738
R6491 DVDD.n5092 DVDD.n573 0.0185738
R6492 DVDD.n5173 DVDD.n470 0.0185738
R6493 DVDD.n597 DVDD.n590 0.0185738
R6494 DVDD.n4964 DVDD.n4946 0.0185738
R6495 DVDD.n876 DVDD.n738 0.0185738
R6496 DVDD.n799 DVDD.n798 0.0185738
R6497 DVDD.n1059 DVDD.n895 0.0185738
R6498 DVDD.n4520 DVDD.n4504 0.0185738
R6499 DVDD.n5919 DVDD.n83 0.018469
R6500 DVDD.n5550 DVDD.n20 0.018469
R6501 DVDD.n4662 DVDD.n4647 0.018469
R6502 DVDD.n5425 DVDD.n327 0.018469
R6503 DVDD.n3186 DVDD.n3185 0.0182974
R6504 DVDD.n3569 DVDD.n3158 0.0182974
R6505 DVDD.n3570 DVDD.n3569 0.0182974
R6506 DVDD.n3185 DVDD.n3181 0.0182974
R6507 DVDD.n5754 DVDD.n173 0.0182049
R6508 DVDD.n5228 DVDD.n488 0.0182049
R6509 DVDD.n638 DVDD.n609 0.0182049
R6510 DVDD.n854 DVDD.n707 0.0182049
R6511 DVDD.n4601 DVDD.n1012 0.0182049
R6512 DVDD.n5544 DVDD.n15 0.0181592
R6513 DVDD.n4668 DVDD.n982 0.0181592
R6514 DVDD.n2839 DVDD.n2692 0.0181087
R6515 DVDD.n2836 DVDD.n2095 0.01805
R6516 DVDD.n3192 DVDD.n3175 0.0178641
R6517 DVDD.n3512 DVDD.n3192 0.0178641
R6518 DVDD.n3523 DVDD.n3162 0.0178641
R6519 DVDD.n3523 DVDD.n3155 0.0178641
R6520 DVDD.n5632 DVDD.n5631 0.0178494
R6521 DVDD.n5527 DVDD.n24 0.0178494
R6522 DVDD.n4685 DVDD.n4651 0.0178494
R6523 DVDD.n5457 DVDD.n5456 0.0178494
R6524 DVDD.n5801 DVDD.n152 0.0178361
R6525 DVDD.n5157 DVDD.n453 0.0178361
R6526 DVDD.n4980 DVDD.n676 0.0178361
R6527 DVDD.n780 DVDD.n751 0.0178361
R6528 DVDD.n4536 DVDD.n1077 0.0178361
R6529 DVDD.n5706 DVDD.n225 0.0176945
R6530 DVDD.n962 DVDD.n944 0.0176945
R6531 DVDD.n1379 DVDD.n1378 0.0176362
R6532 DVDD.n2839 DVDD.n2684 0.0176196
R6533 DVDD.n2098 DVDD.n2092 0.0176
R6534 DVDD.n5770 DVDD.n189 0.0174672
R6535 DVDD.n5212 DVDD.n560 0.0174672
R6536 DVDD.n654 DVDD.n624 0.0174672
R6537 DVDD.n838 DVDD.n720 0.0174672
R6538 DVDD.n4585 DVDD.n1051 0.0174672
R6539 DVDD.n3290 DVDD.n2023 0.017375
R6540 DVDD.n5617 DVDD.n5573 0.0172298
R6541 DVDD.n5442 DVDD.n282 0.0172298
R6542 DVDD.n3589 DVDD.n3127 0.0171304
R6543 DVDD.n3578 DVDD.n3577 0.0171304
R6544 DVDD.n3441 DVDD.n3439 0.0171304
R6545 DVDD.n3466 DVDD.n3194 0.0171304
R6546 DVDD.n5659 DVDD.n5658 0.0170354
R6547 DVDD.n5485 DVDD.n5484 0.0170354
R6548 DVDD.n5909 DVDD.n92 0.0169691
R6549 DVDD.n113 DVDD.n92 0.0169691
R6550 DVDD.n5412 DVDD.n346 0.0169691
R6551 DVDD.n5409 DVDD.n346 0.0169691
R6552 DVDD.n929 DVDD.n925 0.0169691
R6553 DVDD.n929 DVDD.n918 0.0169691
R6554 DVDD.n5664 DVDD.n231 0.0169691
R6555 DVDD.n5664 DVDD.n237 0.0169691
R6556 DVDD.n5634 DVDD.n5606 0.01692
R6557 DVDD.n5459 DVDD.n290 0.01692
R6558 DVDD.n2600 DVDD.n2599 0.0169185
R6559 DVDD.n2213 DVDD.n2212 0.0169185
R6560 DVDD.n2241 DVDD.n2213 0.0169185
R6561 DVDD.n2211 DVDD.n2210 0.0169185
R6562 DVDD.n2242 DVDD.n2211 0.0169185
R6563 DVDD.n2209 DVDD.n2208 0.0169185
R6564 DVDD.n2243 DVDD.n2209 0.0169185
R6565 DVDD.n2207 DVDD.n2206 0.0169185
R6566 DVDD.n2207 DVDD.n2199 0.0169185
R6567 DVDD.n2603 DVDD.n2169 0.0169185
R6568 DVDD.n2617 DVDD.n2197 0.0169185
R6569 DVDD.n2605 DVDD.n2170 0.0169185
R6570 DVDD.n2616 DVDD.n2196 0.0169185
R6571 DVDD.n2606 DVDD.n2171 0.0169185
R6572 DVDD.n2615 DVDD.n2195 0.0169185
R6573 DVDD.n2607 DVDD.n2172 0.0169185
R6574 DVDD.n2614 DVDD.n2194 0.0169185
R6575 DVDD.n2608 DVDD.n2193 0.0169185
R6576 DVDD.n3730 DVDD.n3720 0.0169185
R6577 DVDD.n3730 DVDD.n1857 0.0169185
R6578 DVDD.n3751 DVDD.n3729 0.0169185
R6579 DVDD.n3729 DVDD.n1858 0.0169185
R6580 DVDD.n3750 DVDD.n3728 0.0169185
R6581 DVDD.n3728 DVDD.n1859 0.0169185
R6582 DVDD.n3749 DVDD.n3727 0.0169185
R6583 DVDD.n3727 DVDD.n1860 0.0169185
R6584 DVDD.n3748 DVDD.n1861 0.0169185
R6585 DVDD.n3747 DVDD.n3726 0.0169185
R6586 DVDD.n3726 DVDD.n1862 0.0169185
R6587 DVDD.n3746 DVDD.n3725 0.0169185
R6588 DVDD.n3725 DVDD.n1863 0.0169185
R6589 DVDD.n3745 DVDD.n3724 0.0169185
R6590 DVDD.n3724 DVDD.n1864 0.0169185
R6591 DVDD.n3744 DVDD.n3723 0.0169185
R6592 DVDD.n3723 DVDD.n1865 0.0169185
R6593 DVDD.n3743 DVDD.n3722 0.0169185
R6594 DVDD.n3722 DVDD.n1866 0.0169185
R6595 DVDD.n4341 DVDD.n1629 0.0169185
R6596 DVDD.n4339 DVDD.n1657 0.0169185
R6597 DVDD.n1656 DVDD.n1630 0.0169185
R6598 DVDD.n4338 DVDD.n1655 0.0169185
R6599 DVDD.n1654 DVDD.n1631 0.0169185
R6600 DVDD.n4337 DVDD.n1653 0.0169185
R6601 DVDD.n1652 DVDD.n1632 0.0169185
R6602 DVDD.n4336 DVDD.n1651 0.0169185
R6603 DVDD.n1650 DVDD.n1633 0.0169185
R6604 DVDD.n4335 DVDD.n1649 0.0169185
R6605 DVDD.n1648 DVDD.n1634 0.0169185
R6606 DVDD.n4334 DVDD.n1647 0.0169185
R6607 DVDD.n1646 DVDD.n1635 0.0169185
R6608 DVDD.n4333 DVDD.n1645 0.0169185
R6609 DVDD.n1644 DVDD.n1636 0.0169185
R6610 DVDD.n4332 DVDD.n1643 0.0169185
R6611 DVDD.n1642 DVDD.n1637 0.0169185
R6612 DVDD.n4331 DVDD.n1641 0.0169185
R6613 DVDD.n1640 DVDD.n1638 0.0169185
R6614 DVDD.n4344 DVDD.n1626 0.0169185
R6615 DVDD.n4384 DVDD.n1597 0.0169185
R6616 DVDD.n4382 DVDD.n1625 0.0169185
R6617 DVDD.n1624 DVDD.n1598 0.0169185
R6618 DVDD.n4381 DVDD.n1623 0.0169185
R6619 DVDD.n1622 DVDD.n1599 0.0169185
R6620 DVDD.n4380 DVDD.n1621 0.0169185
R6621 DVDD.n1620 DVDD.n1600 0.0169185
R6622 DVDD.n4379 DVDD.n1619 0.0169185
R6623 DVDD.n1618 DVDD.n1601 0.0169185
R6624 DVDD.n4378 DVDD.n1617 0.0169185
R6625 DVDD.n1616 DVDD.n1602 0.0169185
R6626 DVDD.n4377 DVDD.n1615 0.0169185
R6627 DVDD.n1614 DVDD.n1603 0.0169185
R6628 DVDD.n4376 DVDD.n1613 0.0169185
R6629 DVDD.n1612 DVDD.n1604 0.0169185
R6630 DVDD.n4375 DVDD.n1611 0.0169185
R6631 DVDD.n1610 DVDD.n1605 0.0169185
R6632 DVDD.n4374 DVDD.n1609 0.0169185
R6633 DVDD.n1608 DVDD.n1606 0.0169185
R6634 DVDD.n4387 DVDD.n1594 0.0169185
R6635 DVDD.n4412 DVDD.n1109 0.0169185
R6636 DVDD.n4397 DVDD.n1593 0.0169185
R6637 DVDD.n4400 DVDD.n1110 0.0169185
R6638 DVDD.n4396 DVDD.n1592 0.0169185
R6639 DVDD.n4401 DVDD.n1111 0.0169185
R6640 DVDD.n4395 DVDD.n1591 0.0169185
R6641 DVDD.n4402 DVDD.n1112 0.0169185
R6642 DVDD.n4394 DVDD.n1590 0.0169185
R6643 DVDD.n4403 DVDD.n1113 0.0169185
R6644 DVDD.n4393 DVDD.n1589 0.0169185
R6645 DVDD.n4404 DVDD.n1114 0.0169185
R6646 DVDD.n4392 DVDD.n1588 0.0169185
R6647 DVDD.n4405 DVDD.n1115 0.0169185
R6648 DVDD.n4391 DVDD.n1587 0.0169185
R6649 DVDD.n4406 DVDD.n1116 0.0169185
R6650 DVDD.n4390 DVDD.n1586 0.0169185
R6651 DVDD.n4407 DVDD.n1117 0.0169185
R6652 DVDD.n4389 DVDD.n1585 0.0169185
R6653 DVDD.n4408 DVDD.n1118 0.0169185
R6654 DVDD.n4388 DVDD.n1584 0.0169185
R6655 DVDD.n3774 DVDD.n1866 0.0169185
R6656 DVDD.n3742 DVDD.n1865 0.0169185
R6657 DVDD.n3741 DVDD.n1864 0.0169185
R6658 DVDD.n3740 DVDD.n1863 0.0169185
R6659 DVDD.n3739 DVDD.n1862 0.0169185
R6660 DVDD.n3738 DVDD.n1860 0.0169185
R6661 DVDD.n3737 DVDD.n1859 0.0169185
R6662 DVDD.n3736 DVDD.n1858 0.0169185
R6663 DVDD.n3735 DVDD.n1857 0.0169185
R6664 DVDD.n2608 DVDD.n2194 0.0169185
R6665 DVDD.n2614 DVDD.n2172 0.0169185
R6666 DVDD.n2607 DVDD.n2195 0.0169185
R6667 DVDD.n2615 DVDD.n2171 0.0169185
R6668 DVDD.n2606 DVDD.n2196 0.0169185
R6669 DVDD.n2616 DVDD.n2170 0.0169185
R6670 DVDD.n2605 DVDD.n2197 0.0169185
R6671 DVDD.n2617 DVDD.n2169 0.0169185
R6672 DVDD.n2619 DVDD.n2603 0.0169185
R6673 DVDD.n2602 DVDD.n2199 0.0169185
R6674 DVDD.n2243 DVDD.n2204 0.0169185
R6675 DVDD.n2206 DVDD.n2204 0.0169185
R6676 DVDD.n2242 DVDD.n2203 0.0169185
R6677 DVDD.n2208 DVDD.n2203 0.0169185
R6678 DVDD.n2241 DVDD.n2202 0.0169185
R6679 DVDD.n2210 DVDD.n2202 0.0169185
R6680 DVDD.n2599 DVDD.n2201 0.0169185
R6681 DVDD.n2212 DVDD.n2201 0.0169185
R6682 DVDD.n3776 DVDD.n3720 0.0169185
R6683 DVDD.n3751 DVDD.n3735 0.0169185
R6684 DVDD.n3750 DVDD.n3736 0.0169185
R6685 DVDD.n3749 DVDD.n3737 0.0169185
R6686 DVDD.n3748 DVDD.n3738 0.0169185
R6687 DVDD.n3747 DVDD.n1887 0.0169185
R6688 DVDD.n3746 DVDD.n3739 0.0169185
R6689 DVDD.n3745 DVDD.n3740 0.0169185
R6690 DVDD.n3744 DVDD.n3741 0.0169185
R6691 DVDD.n3743 DVDD.n3742 0.0169185
R6692 DVDD.n4388 DVDD.n1118 0.0169185
R6693 DVDD.n4408 DVDD.n1585 0.0169185
R6694 DVDD.n4389 DVDD.n1117 0.0169185
R6695 DVDD.n4407 DVDD.n1586 0.0169185
R6696 DVDD.n4390 DVDD.n1116 0.0169185
R6697 DVDD.n4406 DVDD.n1587 0.0169185
R6698 DVDD.n4391 DVDD.n1115 0.0169185
R6699 DVDD.n4405 DVDD.n1588 0.0169185
R6700 DVDD.n4392 DVDD.n1114 0.0169185
R6701 DVDD.n4404 DVDD.n1589 0.0169185
R6702 DVDD.n4393 DVDD.n1113 0.0169185
R6703 DVDD.n4403 DVDD.n1590 0.0169185
R6704 DVDD.n4394 DVDD.n1112 0.0169185
R6705 DVDD.n4402 DVDD.n1591 0.0169185
R6706 DVDD.n4395 DVDD.n1111 0.0169185
R6707 DVDD.n4401 DVDD.n1592 0.0169185
R6708 DVDD.n4396 DVDD.n1110 0.0169185
R6709 DVDD.n4400 DVDD.n1593 0.0169185
R6710 DVDD.n4397 DVDD.n1109 0.0169185
R6711 DVDD.n4413 DVDD.n4412 0.0169185
R6712 DVDD.n1606 DVDD.n1594 0.0169185
R6713 DVDD.n1609 DVDD.n1608 0.0169185
R6714 DVDD.n4374 DVDD.n1605 0.0169185
R6715 DVDD.n1611 DVDD.n1610 0.0169185
R6716 DVDD.n4375 DVDD.n1604 0.0169185
R6717 DVDD.n1613 DVDD.n1612 0.0169185
R6718 DVDD.n4376 DVDD.n1603 0.0169185
R6719 DVDD.n1615 DVDD.n1614 0.0169185
R6720 DVDD.n4377 DVDD.n1602 0.0169185
R6721 DVDD.n1617 DVDD.n1616 0.0169185
R6722 DVDD.n4378 DVDD.n1601 0.0169185
R6723 DVDD.n1619 DVDD.n1618 0.0169185
R6724 DVDD.n4379 DVDD.n1600 0.0169185
R6725 DVDD.n1621 DVDD.n1620 0.0169185
R6726 DVDD.n4380 DVDD.n1599 0.0169185
R6727 DVDD.n1623 DVDD.n1622 0.0169185
R6728 DVDD.n4381 DVDD.n1598 0.0169185
R6729 DVDD.n1625 DVDD.n1624 0.0169185
R6730 DVDD.n4382 DVDD.n1597 0.0169185
R6731 DVDD.n4385 DVDD.n4384 0.0169185
R6732 DVDD.n1638 DVDD.n1626 0.0169185
R6733 DVDD.n1641 DVDD.n1640 0.0169185
R6734 DVDD.n4331 DVDD.n1637 0.0169185
R6735 DVDD.n1643 DVDD.n1642 0.0169185
R6736 DVDD.n4332 DVDD.n1636 0.0169185
R6737 DVDD.n1645 DVDD.n1644 0.0169185
R6738 DVDD.n4333 DVDD.n1635 0.0169185
R6739 DVDD.n1647 DVDD.n1646 0.0169185
R6740 DVDD.n4334 DVDD.n1634 0.0169185
R6741 DVDD.n1649 DVDD.n1648 0.0169185
R6742 DVDD.n4335 DVDD.n1633 0.0169185
R6743 DVDD.n1651 DVDD.n1650 0.0169185
R6744 DVDD.n4336 DVDD.n1632 0.0169185
R6745 DVDD.n1653 DVDD.n1652 0.0169185
R6746 DVDD.n4337 DVDD.n1631 0.0169185
R6747 DVDD.n1655 DVDD.n1654 0.0169185
R6748 DVDD.n4338 DVDD.n1630 0.0169185
R6749 DVDD.n1657 DVDD.n1656 0.0169185
R6750 DVDD.n4339 DVDD.n1629 0.0169185
R6751 DVDD.n4342 DVDD.n4341 0.0169185
R6752 DVDD.n5775 DVDD.n179 0.0167295
R6753 DVDD.n5785 DVDD.n5784 0.0167295
R6754 DVDD.n5845 DVDD.n138 0.0167295
R6755 DVDD.n5202 DVDD.n494 0.0167295
R6756 DVDD.n5196 DVDD.n495 0.0167295
R6757 DVDD.n5139 DVDD.n5138 0.0167295
R6758 DVDD.n664 DVDD.n615 0.0167295
R6759 DVDD.n626 DVDD.n606 0.0167295
R6760 DVDD.n4992 DVDD.n427 0.0167295
R6761 DVDD.n828 DVDD.n713 0.0167295
R6762 DVDD.n822 DVDD.n714 0.0167295
R6763 DVDD.n758 DVDD.n403 0.0167295
R6764 DVDD.n4575 DVDD.n1018 0.0167295
R6765 DVDD.n4569 DVDD.n1019 0.0167295
R6766 DVDD.n4548 DVDD.n380 0.0167295
R6767 DVDD.n2828 DVDD.n2091 0.0167
R6768 DVDD.n3284 DVDD.n3269 0.0166964
R6769 DVDD.n5566 DVDD.n5565 0.0166102
R6770 DVDD.n275 DVDD.n274 0.0166102
R6771 DVDD.n5642 DVDD.n66 0.0164553
R6772 DVDD.n5467 DVDD.n299 0.0164553
R6773 DVDD.n3499 DVDD.n3190 0.0163967
R6774 DVDD.n3531 DVDD.n3164 0.0163967
R6775 DVDD.n5835 DVDD.n142 0.0163607
R6776 DVDD.n5317 DVDD.n473 0.0163607
R6777 DVDD.n5003 DVDD.n4949 0.0163607
R6778 DVDD.n770 DVDD.n769 0.0163607
R6779 DVDD.n4559 DVDD.n4507 0.0163607
R6780 DVDD.n5519 DVDD.n9 0.0163003
R6781 DVDD.n4693 DVDD.n976 0.0163003
R6782 DVDD.n2828 DVDD.n2094 0.01625
R6783 DVDD.n2851 DVDD.n2690 0.0161522
R6784 DVDD.n5625 DVDD.n54 0.0161454
R6785 DVDD.n5450 DVDD.n312 0.0161454
R6786 DVDD.n5764 DVDD.n177 0.0159918
R6787 DVDD.n5218 DVDD.n561 0.0159918
R6788 DVDD.n648 DVDD.n613 0.0159918
R6789 DVDD.n844 DVDD.n721 0.0159918
R6790 DVDD.n4591 DVDD.n1052 0.0159918
R6791 DVDD.n5535 DVDD.n23 0.0159905
R6792 DVDD.n4677 DVDD.n4650 0.0159905
R6793 DVDD.n71 DVDD.n59 0.0158356
R6794 DVDD.n5434 DVDD.n306 0.0158356
R6795 DVDD.n5552 DVDD.n16 0.0156807
R6796 DVDD.n5558 DVDD.n8 0.0156807
R6797 DVDD.n4660 DVDD.n983 0.0156807
R6798 DVDD.n4644 DVDD.n267 0.0156807
R6799 DVDD.n3121 DVDD.n3120 0.015663
R6800 DVDD.n3430 DVDD.n3210 0.015663
R6801 DVDD.n2838 DVDD.n2837 0.0156593
R6802 DVDD.n5807 DVDD.n151 0.015623
R6803 DVDD.n5163 DVDD.n465 0.015623
R6804 DVDD.n4974 DVDD.n4941 0.015623
R6805 DVDD.n787 DVDD.n786 0.015623
R6806 DVDD.n4530 DVDD.n4500 0.015623
R6807 DVDD.n939 DVDD.n928 0.0155811
R6808 DVDD.n939 DVDD.n938 0.0155811
R6809 DVDD.n938 DVDD.n935 0.0155811
R6810 DVDD.n935 DVDD.n934 0.0155811
R6811 DVDD.n934 DVDD.n932 0.0155811
R6812 DVDD.n932 DVDD.n930 0.0155811
R6813 DVDD.n953 DVDD.n951 0.0155811
R6814 DVDD.n954 DVDD.n953 0.0155811
R6815 DVDD.n957 DVDD.n954 0.0155811
R6816 DVDD.n959 DVDD.n957 0.0155811
R6817 DVDD.n960 DVDD.n959 0.0155811
R6818 DVDD.n1909 DVDD.n1897 0.015575
R6819 DVDD.n3341 DVDD.n2023 0.015575
R6820 DVDD.n1910 DVDD.n1896 0.015575
R6821 DVDD.n3617 DVDD.n3097 0.015575
R6822 DVDD.n258 DVDD.n243 0.0154398
R6823 DVDD.n5671 DVDD.n243 0.0154398
R6824 DVDD.n5671 DVDD.n5670 0.0154398
R6825 DVDD.n5670 DVDD.n5669 0.0154398
R6826 DVDD.n5669 DVDD.n5667 0.0154398
R6827 DVDD.n5667 DVDD.n5665 0.0154398
R6828 DVDD.n255 DVDD.n253 0.0154398
R6829 DVDD.n253 DVDD.n251 0.0154398
R6830 DVDD.n251 DVDD.n248 0.0154398
R6831 DVDD.n248 DVDD.n247 0.0154398
R6832 DVDD.n247 DVDD.n245 0.0154398
R6833 DVDD.n5542 DVDD.n21 0.0153709
R6834 DVDD.n4670 DVDD.n4648 0.0153709
R6835 DVDD.n2946 DVDD.n2098 0.01535
R6836 DVDD.n104 DVDD.n98 0.0153356
R6837 DVDD.n5916 DVDD.n101 0.0153356
R6838 DVDD.n5419 DVDD.n337 0.0153356
R6839 DVDD.n5421 DVDD.n348 0.0153356
R6840 DVDD.n5419 DVDD.n344 0.0153356
R6841 DVDD.n104 DVDD.n90 0.0153356
R6842 DVDD.n101 DVDD.n88 0.0153356
R6843 DVDD.n348 DVDD.n334 0.0153356
R6844 DVDD.n2189 DVDD.n2188 0.0153088
R6845 DVDD.n2188 DVDD.n2178 0.0153088
R6846 DVDD.n2181 DVDD.n2178 0.0153088
R6847 DVDD.n3706 DVDD.n1892 0.0153088
R6848 DVDD.n3715 DVDD.n1892 0.0153088
R6849 DVDD.n3715 DVDD.n1890 0.0153088
R6850 DVDD.n3769 DVDD.n3755 0.0153088
R6851 DVDD.n3769 DVDD.n3757 0.0153088
R6852 DVDD.n3762 DVDD.n3757 0.0153088
R6853 DVDD.n4287 DVDD.n1662 0.0153088
R6854 DVDD.n4295 DVDD.n1662 0.0153088
R6855 DVDD.n4295 DVDD.n1660 0.0153088
R6856 DVDD.n5748 DVDD.n175 0.0152541
R6857 DVDD.n5234 DVDD.n487 0.0152541
R6858 DVDD.n632 DVDD.n611 0.0152541
R6859 DVDD.n860 DVDD.n706 0.0152541
R6860 DVDD.n4607 DVDD.n1011 0.0152541
R6861 DVDD.n5525 DVDD.n11 0.0150611
R6862 DVDD.n4687 DVDD.n978 0.0150611
R6863 DVDD.n1122 DVDD.n1119 0.015031
R6864 DVDD.n1581 DVDD.n1149 0.015031
R6865 DVDD.n1580 DVDD.n1123 0.015031
R6866 DVDD.n1148 DVDD.n1147 0.015031
R6867 DVDD.n1182 DVDD.n1124 0.015031
R6868 DVDD.n1146 DVDD.n1145 0.015031
R6869 DVDD.n1183 DVDD.n1125 0.015031
R6870 DVDD.n1144 DVDD.n1143 0.015031
R6871 DVDD.n1184 DVDD.n1126 0.015031
R6872 DVDD.n1142 DVDD.n1141 0.015031
R6873 DVDD.n1185 DVDD.n1127 0.015031
R6874 DVDD.n1140 DVDD.n1139 0.015031
R6875 DVDD.n1186 DVDD.n1128 0.015031
R6876 DVDD.n1138 DVDD.n1137 0.015031
R6877 DVDD.n1187 DVDD.n1129 0.015031
R6878 DVDD.n1136 DVDD.n1135 0.015031
R6879 DVDD.n1188 DVDD.n1130 0.015031
R6880 DVDD.n1134 DVDD.n1133 0.015031
R6881 DVDD.n1190 DVDD.n1189 0.015031
R6882 DVDD.n1578 DVDD.n1132 0.015031
R6883 DVDD.n1189 DVDD.n1132 0.015031
R6884 DVDD.n1190 DVDD.n1134 0.015031
R6885 DVDD.n1133 DVDD.n1130 0.015031
R6886 DVDD.n1188 DVDD.n1136 0.015031
R6887 DVDD.n1135 DVDD.n1129 0.015031
R6888 DVDD.n1187 DVDD.n1138 0.015031
R6889 DVDD.n1137 DVDD.n1128 0.015031
R6890 DVDD.n1186 DVDD.n1140 0.015031
R6891 DVDD.n1139 DVDD.n1127 0.015031
R6892 DVDD.n1185 DVDD.n1142 0.015031
R6893 DVDD.n1141 DVDD.n1126 0.015031
R6894 DVDD.n1184 DVDD.n1144 0.015031
R6895 DVDD.n1143 DVDD.n1125 0.015031
R6896 DVDD.n1183 DVDD.n1146 0.015031
R6897 DVDD.n1145 DVDD.n1124 0.015031
R6898 DVDD.n1182 DVDD.n1148 0.015031
R6899 DVDD.n1147 DVDD.n1123 0.015031
R6900 DVDD.n1581 DVDD.n1580 0.015031
R6901 DVDD.n1149 DVDD.n1122 0.015031
R6902 DVDD.n1583 DVDD.n1119 0.015031
R6903 DVDD.n1382 DVDD.n1307 0.0149495
R6904 DVDD.n1390 DVDD.n1311 0.0149495
R6905 DVDD.n1318 DVDD.n1219 0.0149495
R6906 DVDD.n1314 DVDD.n1221 0.0149495
R6907 DVDD.n3491 DVDD.n3178 0.0149293
R6908 DVDD.n3539 DVDD.n3152 0.0149293
R6909 DVDD.n2801 DVDD.n2704 0.0149069
R6910 DVDD.n2804 DVDD.n2701 0.0149069
R6911 DVDD.n2704 DVDD.n2701 0.0149069
R6912 DVDD.n2802 DVDD.n2801 0.0149069
R6913 DVDD.n5502 DVDD.n221 0.0149062
R6914 DVDD.n964 DVDD.n947 0.0149062
R6915 DVDD.n2836 DVDD.n2089 0.0149
R6916 DVDD.n3772 DVDD.n3754 0.0148917
R6917 DVDD.n3759 DVDD.n3758 0.0148917
R6918 DVDD.n3768 DVDD.n3767 0.0148917
R6919 DVDD.n3764 DVDD.n3760 0.0148917
R6920 DVDD.n4289 DVDD.n4288 0.0148917
R6921 DVDD.n4292 DVDD.n1663 0.0148917
R6922 DVDD.n4294 DVDD.n4293 0.0148917
R6923 DVDD.n4298 DVDD.n1659 0.0148917
R6924 DVDD.n5738 DVDD.n193 0.0148852
R6925 DVDD.n5823 DVDD.n162 0.0148852
R6926 DVDD.n5096 DVDD.n5095 0.0148852
R6927 DVDD.n5179 DVDD.n467 0.0148852
R6928 DVDD.n5019 DVDD.n5018 0.0148852
R6929 DVDD.n4958 DVDD.n4943 0.0148852
R6930 DVDD.n870 DVDD.n737 0.0148852
R6931 DVDD.n805 DVDD.n804 0.0148852
R6932 DVDD.n1066 DVDD.n894 0.0148852
R6933 DVDD.n4514 DVDD.n4502 0.0148852
R6934 DVDD.n2859 DVDD.n2687 0.0146848
R6935 DVDD.n5619 DVDD.n5603 0.0144415
R6936 DVDD.n5444 DVDD.n287 0.0144415
R6937 DVDD.n2399 DVDD.n2398 0.0142903
R6938 DVDD.n2981 DVDD.n2980 0.0142903
R6939 DVDD.n1915 DVDD.n1907 0.014225
R6940 DVDD.n1363 DVDD.n1362 0.0141845
R6941 DVDD.n3603 DVDD.n3110 0.0141679
R6942 DVDD.n3413 DVDD.n3411 0.0141679
R6943 DVDD.n3414 DVDD.n3412 0.0141679
R6944 DVDD.n3604 DVDD.n3112 0.0141679
R6945 DVDD.n3412 DVDD.n3209 0.0141679
R6946 DVDD.n3415 DVDD.n3413 0.0141679
R6947 DVDD.n3123 DVDD.n3112 0.0141679
R6948 DVDD.n3605 DVDD.n3110 0.0141679
R6949 DVDD.n2844 DVDD.n2694 0.0141679
R6950 DVDD.n2844 DVDD.n2843 0.0141679
R6951 DVDD.n2843 DVDD.n2840 0.0141679
R6952 DVDD.n2841 DVDD.n2694 0.0141679
R6953 DVDD.n2191 DVDD.n2190 0.0141616
R6954 DVDD.n2187 DVDD.n2175 0.0141616
R6955 DVDD.n2186 DVDD.n2179 0.0141616
R6956 DVDD.n2183 DVDD.n2182 0.0141616
R6957 DVDD.n3709 DVDD.n3708 0.0141616
R6958 DVDD.n3714 DVDD.n1893 0.0141616
R6959 DVDD.n3713 DVDD.n1894 0.0141616
R6960 DVDD.n3718 DVDD.n1889 0.0141616
R6961 DVDD.n5636 DVDD.n5569 0.0141317
R6962 DVDD.n5461 DVDD.n278 0.0141317
R6963 DVDD.n1374 DVDD.n1328 0.0140776
R6964 DVDD.n1328 DVDD.n1327 0.0140776
R6965 DVDD.n3473 DVDD.n3184 0.013978
R6966 DVDD.n3556 DVDD.n3160 0.013978
R6967 DVDD.n3481 DVDD.n3187 0.0139511
R6968 DVDD.n3549 DVDD.n3167 0.0139511
R6969 DVDD.n5651 DVDD.n5650 0.0138219
R6970 DVDD.n5477 DVDD.n5476 0.0138219
R6971 DVDD.n2703 DVDD.n2700 0.0137065
R6972 DVDD.n5640 DVDD.n51 0.013667
R6973 DVDD.n5507 DVDD.n218 0.013667
R6974 DVDD.n4705 DVDD.n948 0.013667
R6975 DVDD.n5465 DVDD.n315 0.013667
R6976 DVDD DVDD.n2735 0.0135263
R6977 DVDD.n5521 DVDD.n26 0.013512
R6978 DVDD.n4691 DVDD.n4653 0.013512
R6979 DVDD.n3639 DVDD.n2015 0.0135078
R6980 DVDD.n3483 DVDD.n3187 0.013462
R6981 DVDD.n3547 DVDD.n3167 0.013462
R6982 DVDD.n3378 DVDD.n3242 0.0134255
R6983 DVDD.n3376 DVDD.n3242 0.0134255
R6984 DVDD.n3326 DVDD.n3278 0.0134255
R6985 DVDD.n3313 DVDD.n3278 0.0134255
R6986 DVDD.n963 DVDD.n961 0.0134017
R6987 DVDD.n965 DVDD.n963 0.0134017
R6988 DVDD.n969 DVDD.n968 0.0134017
R6989 DVDD.n4703 DVDD.n969 0.0134017
R6990 DVDD.n4703 DVDD.n4702 0.0134017
R6991 DVDD.n4702 DVDD.n4701 0.0134017
R6992 DVDD.n4701 DVDD.n970 0.0134017
R6993 DVDD.n4655 DVDD.n970 0.0134017
R6994 DVDD.n4695 DVDD.n4655 0.0134017
R6995 DVDD.n4695 DVDD.n4694 0.0134017
R6996 DVDD.n4694 DVDD.n4692 0.0134017
R6997 DVDD.n4692 DVDD.n4690 0.0134017
R6998 DVDD.n4690 DVDD.n4688 0.0134017
R6999 DVDD.n4688 DVDD.n4686 0.0134017
R7000 DVDD.n4686 DVDD.n4684 0.0134017
R7001 DVDD.n4684 DVDD.n4681 0.0134017
R7002 DVDD.n4681 DVDD.n4680 0.0134017
R7003 DVDD.n4680 DVDD.n4678 0.0134017
R7004 DVDD.n4675 DVDD.n4673 0.0134017
R7005 DVDD.n4673 DVDD.n4671 0.0134017
R7006 DVDD.n4671 DVDD.n4669 0.0134017
R7007 DVDD.n4669 DVDD.n4667 0.0134017
R7008 DVDD.n4667 DVDD.n4664 0.0134017
R7009 DVDD.n4664 DVDD.n4663 0.0134017
R7010 DVDD.n4663 DVDD.n4661 0.0134017
R7011 DVDD.n4661 DVDD.n4659 0.0134017
R7012 DVDD.n4659 DVDD.n4657 0.0134017
R7013 DVDD.n4657 DVDD.n265 0.0134017
R7014 DVDD.n5479 DVDD.n266 0.0134017
R7015 DVDD.n5479 DVDD.n5478 0.0134017
R7016 DVDD.n5478 DVDD.n269 0.0134017
R7017 DVDD.n318 DVDD.n269 0.0134017
R7018 DVDD.n319 DVDD.n318 0.0134017
R7019 DVDD.n5469 DVDD.n319 0.0134017
R7020 DVDD.n5469 DVDD.n5468 0.0134017
R7021 DVDD.n5468 DVDD.n5466 0.0134017
R7022 DVDD.n5466 DVDD.n5464 0.0134017
R7023 DVDD.n5464 DVDD.n5462 0.0134017
R7024 DVDD.n5462 DVDD.n5460 0.0134017
R7025 DVDD.n5460 DVDD.n5458 0.0134017
R7026 DVDD.n5454 DVDD.n5453 0.0134017
R7027 DVDD.n5453 DVDD.n5451 0.0134017
R7028 DVDD.n5451 DVDD.n5449 0.0134017
R7029 DVDD.n5449 DVDD.n5447 0.0134017
R7030 DVDD.n5447 DVDD.n5445 0.0134017
R7031 DVDD.n5445 DVDD.n5443 0.0134017
R7032 DVDD.n5443 DVDD.n5441 0.0134017
R7033 DVDD.n5441 DVDD.n5438 0.0134017
R7034 DVDD.n5438 DVDD.n5437 0.0134017
R7035 DVDD.n5437 DVDD.n5435 0.0134017
R7036 DVDD.n5435 DVDD.n5433 0.0134017
R7037 DVDD.n5433 DVDD.n5432 0.0134017
R7038 DVDD.n5432 DVDD.n5431 0.0134017
R7039 DVDD.n5431 DVDD.n320 0.0134017
R7040 DVDD.n330 DVDD.n320 0.0134017
R7041 DVDD.n332 DVDD.n330 0.0134017
R7042 DVDD.n5424 DVDD.n5423 0.0134017
R7043 DVDD.n5483 DVDD.n266 0.0134017
R7044 DVDD.n5657 DVDD.n5560 0.013372
R7045 DVDD.n5501 DVDD.n223 0.013372
R7046 DVDD.n5503 DVDD.n5501 0.013372
R7047 DVDD.n5508 DVDD.n5506 0.013372
R7048 DVDD.n5509 DVDD.n5508 0.013372
R7049 DVDD.n5512 DVDD.n5509 0.013372
R7050 DVDD.n5513 DVDD.n5512 0.013372
R7051 DVDD.n5514 DVDD.n5513 0.013372
R7052 DVDD.n5516 DVDD.n5514 0.013372
R7053 DVDD.n5518 DVDD.n5516 0.013372
R7054 DVDD.n5520 DVDD.n5518 0.013372
R7055 DVDD.n5522 DVDD.n5520 0.013372
R7056 DVDD.n5524 DVDD.n5522 0.013372
R7057 DVDD.n5526 DVDD.n5524 0.013372
R7058 DVDD.n5528 DVDD.n5526 0.013372
R7059 DVDD.n5529 DVDD.n5528 0.013372
R7060 DVDD.n5532 DVDD.n5529 0.013372
R7061 DVDD.n5534 DVDD.n5532 0.013372
R7062 DVDD.n5536 DVDD.n5534 0.013372
R7063 DVDD.n5541 DVDD.n5539 0.013372
R7064 DVDD.n5543 DVDD.n5541 0.013372
R7065 DVDD.n5545 DVDD.n5543 0.013372
R7066 DVDD.n5546 DVDD.n5545 0.013372
R7067 DVDD.n5549 DVDD.n5546 0.013372
R7068 DVDD.n5551 DVDD.n5549 0.013372
R7069 DVDD.n5553 DVDD.n5551 0.013372
R7070 DVDD.n5555 DVDD.n5553 0.013372
R7071 DVDD.n5557 DVDD.n5555 0.013372
R7072 DVDD.n5559 DVDD.n5557 0.013372
R7073 DVDD.n5653 DVDD.n5560 0.013372
R7074 DVDD.n5653 DVDD.n5652 0.013372
R7075 DVDD.n5652 DVDD.n5562 0.013372
R7076 DVDD.n5610 DVDD.n5562 0.013372
R7077 DVDD.n5646 DVDD.n5610 0.013372
R7078 DVDD.n5646 DVDD.n5645 0.013372
R7079 DVDD.n5645 DVDD.n5643 0.013372
R7080 DVDD.n5643 DVDD.n5641 0.013372
R7081 DVDD.n5641 DVDD.n5639 0.013372
R7082 DVDD.n5639 DVDD.n5637 0.013372
R7083 DVDD.n5637 DVDD.n5635 0.013372
R7084 DVDD.n5635 DVDD.n5633 0.013372
R7085 DVDD.n5629 DVDD.n5628 0.013372
R7086 DVDD.n5628 DVDD.n5626 0.013372
R7087 DVDD.n5626 DVDD.n5624 0.013372
R7088 DVDD.n5624 DVDD.n5622 0.013372
R7089 DVDD.n5622 DVDD.n5620 0.013372
R7090 DVDD.n5620 DVDD.n5618 0.013372
R7091 DVDD.n5618 DVDD.n5616 0.013372
R7092 DVDD.n5616 DVDD.n5613 0.013372
R7093 DVDD.n5613 DVDD.n5612 0.013372
R7094 DVDD.n5612 DVDD.n72 0.013372
R7095 DVDD.n5929 DVDD.n72 0.013372
R7096 DVDD.n5929 DVDD.n5928 0.013372
R7097 DVDD.n5928 DVDD.n73 0.013372
R7098 DVDD.n5924 DVDD.n73 0.013372
R7099 DVDD.n5924 DVDD.n5923 0.013372
R7100 DVDD.n5923 DVDD.n75 0.013372
R7101 DVDD.n5918 DVDD.n86 0.013372
R7102 DVDD.n5623 DVDD.n62 0.0133571
R7103 DVDD.n5448 DVDD.n303 0.0133571
R7104 DVDD.n1371 DVDD.n1200 0.0132218
R7105 DVDD.n5538 DVDD.n13 0.0132022
R7106 DVDD.n4674 DVDD.n980 0.0132022
R7107 DVDD.n5931 DVDD.n5930 0.0130473
R7108 DVDD.n308 DVDD.n294 0.0130473
R7109 DVDD.n5922 DVDD.n5921 0.0128924
R7110 DVDD.n5554 DVDD.n19 0.0128924
R7111 DVDD.n5556 DVDD.n18 0.0128924
R7112 DVDD.n4658 DVDD.n4646 0.0128924
R7113 DVDD.n4656 DVDD.n4645 0.0128924
R7114 DVDD.n326 DVDD.n323 0.0128924
R7115 DVDD.n5909 DVDD.n97 0.0127938
R7116 DVDD.n113 DVDD.n96 0.0127938
R7117 DVDD.n5412 DVDD.n336 0.0127938
R7118 DVDD.n5409 DVDD.n335 0.0127938
R7119 DVDD.n931 DVDD.n925 0.0127938
R7120 DVDD.n950 DVDD.n918 0.0127938
R7121 DVDD.n5666 DVDD.n231 0.0127938
R7122 DVDD.n254 DVDD.n237 0.0127938
R7123 DVDD.n2862 DVDD.n2687 0.0127283
R7124 DVDD.n5833 DVDD.n5832 0.0126721
R7125 DVDD.n5187 DVDD.n469 0.0126721
R7126 DVDD.n4950 DVDD.n4945 0.0126721
R7127 DVDD.n814 DVDD.n813 0.0126721
R7128 DVDD.n4561 DVDD.n1074 0.0126721
R7129 DVDD.n3665 DVDD.n3663 0.0126289
R7130 DVDD.n5540 DVDD.n14 0.0125826
R7131 DVDD.n4672 DVDD.n981 0.0125826
R7132 DVDD.n1370 DVDD.n1369 0.0125
R7133 DVDD.n3489 DVDD.n3178 0.0124837
R7134 DVDD.n3541 DVDD.n3152 0.0124837
R7135 DVDD.n1887 DVDD.n1886 0.012425
R7136 DVDD.n5523 DVDD.n25 0.0122728
R7137 DVDD.n4689 DVDD.n4652 0.0122728
R7138 DVDD.n5458 DVDD.n5455 0.0121532
R7139 DVDD.n5633 DVDD.n5630 0.0121263
R7140 DVDD.n5505 DVDD.n219 0.0121179
R7141 DVDD.n967 DVDD.n945 0.0121179
R7142 DVDD.n5815 DVDD.n149 0.0119344
R7143 DVDD.n5171 DVDD.n454 0.0119344
R7144 DVDD.n4966 DVDD.n677 0.0119344
R7145 DVDD.n797 DVDD.n796 0.0119344
R7146 DVDD.n4522 DVDD.n1078 0.0119344
R7147 DVDD.n1205 DVDD.n1193 0.0117585
R7148 DVDD.n3120 DVDD.n3113 0.01175
R7149 DVDD.n3417 DVDD.n3210 0.01175
R7150 DVDD.n3288 DVDD.n2022 0.01175
R7151 DVDD.n5621 DVDD.n5572 0.0116532
R7152 DVDD.n5446 DVDD.n281 0.0116532
R7153 DVDD.n5484 DVDD.n265 0.0116329
R7154 DVDD.n5658 DVDD.n5559 0.0116073
R7155 DVDD.n5756 DVDD.n188 0.0115656
R7156 DVDD.n5226 DVDD.n563 0.0115656
R7157 DVDD.n640 DVDD.n623 0.0115656
R7158 DVDD.n852 DVDD.n723 0.0115656
R7159 DVDD.n4599 DVDD.n1054 0.0115656
R7160 DVDD.n5638 DVDD.n5607 0.0113434
R7161 DVDD.n5463 DVDD.n291 0.0113434
R7162 DVDD.n2853 DVDD.n2690 0.0112609
R7163 DVDD.n5799 DVDD.n157 0.0111967
R7164 DVDD.n5155 DVDD.n472 0.0111967
R7165 DVDD.n4982 DVDD.n4948 0.0111967
R7166 DVDD.n779 DVDD.n778 0.0111967
R7167 DVDD.n4538 DVDD.n4506 0.0111967
R7168 DVDD.n5654 DVDD.n5561 0.0110336
R7169 DVDD.n5480 DVDD.n268 0.0110336
R7170 DVDD.n3497 DVDD.n3190 0.0110163
R7171 DVDD.n3533 DVDD.n3164 0.0110163
R7172 DVDD.n5638 DVDD.n65 0.0108787
R7173 DVDD.n5505 DVDD.n222 0.0108787
R7174 DVDD.n967 DVDD.n946 0.0108787
R7175 DVDD.n5463 DVDD.n300 0.0108787
R7176 DVDD.n190 DVDD.n171 0.0108279
R7177 DVDD.n5210 DVDD.n492 0.0108279
R7178 DVDD.n656 DVDD.n607 0.0108279
R7179 DVDD.n836 DVDD.n711 0.0108279
R7180 DVDD.n4583 DVDD.n1016 0.0108279
R7181 DVDD.n5523 DVDD.n10 0.0107238
R7182 DVDD.n4689 DVDD.n977 0.0107238
R7183 DVDD.n1577 DVDD.n1191 0.0105885
R7184 DVDD.n1203 DVDD.n1196 0.0105885
R7185 DVDD.n1204 DVDD.n1195 0.0105885
R7186 DVDD.n1575 DVDD.n1574 0.0105885
R7187 DVDD.n1574 DVDD.n1194 0.0105885
R7188 DVDD.n1204 DVDD.n1202 0.0105885
R7189 DVDD.n1203 DVDD.n1200 0.0105885
R7190 DVDD.n1199 DVDD.n1191 0.0105885
R7191 DVDD.n1198 DVDD.n1196 0.0105885
R7192 DVDD.n1201 DVDD.n1194 0.0105885
R7193 DVDD.n1202 DVDD.n1201 0.0105885
R7194 DVDD.n1199 DVDD.n1198 0.0105885
R7195 DVDD.n5621 DVDD.n55 0.0105688
R7196 DVDD.n5446 DVDD.n311 0.0105688
R7197 DVDD.n3704 DVDD.n1903 0.01055
R7198 DVDD.n5540 DVDD.n22 0.0104139
R7199 DVDD.n4672 DVDD.n4649 0.0104139
R7200 DVDD.n3079 DVDD.n2033 0.0104
R7201 DVDD.n3609 DVDD.n3608 0.0104
R7202 DVDD.n3607 DVDD.n3103 0.0104
R7203 DVDD.n3407 DVDD.n3406 0.0104
R7204 DVDD.n3405 DVDD.n3214 0.0104
R7205 DVDD.n3630 DVDD.n2017 0.0104
R7206 DVDD.n2177 DVDD.n2176 0.0103725
R7207 DVDD.n2177 DVDD.n1968 0.0103725
R7208 DVDD.n3705 DVDD.n1891 0.0103725
R7209 DVDD.n3716 DVDD.n1891 0.0103725
R7210 DVDD.n3770 DVDD.n3756 0.0103725
R7211 DVDD.n3756 DVDD.n1667 0.0103725
R7212 DVDD.n4286 DVDD.n1661 0.0103725
R7213 DVDD.n4296 DVDD.n1661 0.0103725
R7214 DVDD.n3590 DVDD.n3589 0.0102826
R7215 DVDD.n3577 DVDD.n3140 0.0102826
R7216 DVDD.n3439 DVDD.n3436 0.0102826
R7217 DVDD.n3469 DVDD.n3194 0.0102826
R7218 DVDD.n5927 DVDD.n48 0.010259
R7219 DVDD.n5473 DVDD.n296 0.010259
R7220 DVDD.n3629 DVDD.n3628 0.01025
R7221 DVDD.n3367 DVDD.n3276 0.0102297
R7222 DVDD.n3377 DVDD.n3243 0.0102297
R7223 DVDD.n5925 DVDD.n74 0.0101041
R7224 DVDD.n5922 DVDD.n74 0.0101041
R7225 DVDD.n5554 DVDD.n17 0.0101041
R7226 DVDD.n5556 DVDD.n17 0.0101041
R7227 DVDD.n4658 DVDD.n984 0.0101041
R7228 DVDD.n4656 DVDD.n984 0.0101041
R7229 DVDD.n5429 DVDD.n5428 0.0101041
R7230 DVDD.n5428 DVDD.n323 0.0101041
R7231 DVDD.n5777 DVDD.n182 0.0100902
R7232 DVDD.n5788 DVDD.n166 0.0100902
R7233 DVDD.n5204 DVDD.n558 0.0100902
R7234 DVDD.n5194 DVDD.n556 0.0100902
R7235 DVDD.n662 DVDD.n618 0.0100902
R7236 DVDD.n5011 DVDD.n5010 0.0100902
R7237 DVDD.n830 DVDD.n718 0.0100902
R7238 DVDD.n820 DVDD.n716 0.0100902
R7239 DVDD.n4577 DVDD.n1049 0.0100902
R7240 DVDD.n4567 DVDD.n1047 0.0100902
R7241 DVDD.n2065 DVDD.n2064 0.01007
R7242 DVDD.n2946 DVDD.n2096 0.00995
R7243 DVDD.n84 DVDD.n81 0.00994923
R7244 DVDD.n5426 DVDD.n329 0.00994923
R7245 DVDD.n3038 DVDD.n3033 0.00992
R7246 DVDD.n3574 DVDD.n3144 0.00992
R7247 DVDD.n3462 DVDD.n3201 0.00992
R7248 DVDD.n3677 DVDD.n1974 0.00992
R7249 DVDD.n3676 DVDD.n3675 0.00992
R7250 DVDD.n3055 DVDD.n3054 0.00983
R7251 DVDD.n5538 DVDD.n22 0.00979432
R7252 DVDD.n4674 DVDD.n4649 0.00979432
R7253 DVDD.n2845 DVDD.n2684 0.00979348
R7254 DVDD.n3576 DVDD.n3575 0.00977
R7255 DVDD.n3200 DVDD.n3198 0.00977
R7256 DVDD.n3617 DVDD.n3089 0.009725
R7257 DVDD.n5793 DVDD.n154 0.00972131
R7258 DVDD.n5149 DVDD.n461 0.00972131
R7259 DVDD.n4988 DVDD.n683 0.00972131
R7260 DVDD.n772 DVDD.n771 0.00972131
R7261 DVDD.n4544 DVDD.n1084 0.00972131
R7262 DVDD.n2596 DVDD.n2595 0.00962857
R7263 DVDD.n2595 DVDD.n2244 0.00962857
R7264 DVDD.n2591 DVDD.n2244 0.00962857
R7265 DVDD.n2591 DVDD.n2246 0.00962857
R7266 DVDD.n2587 DVDD.n2246 0.00962857
R7267 DVDD.n2587 DVDD.n2248 0.00962857
R7268 DVDD.n2583 DVDD.n2248 0.00962857
R7269 DVDD.n2583 DVDD.n2250 0.00962857
R7270 DVDD.n2579 DVDD.n2250 0.00962857
R7271 DVDD.n2579 DVDD.n2252 0.00962857
R7272 DVDD.n2575 DVDD.n2252 0.00962857
R7273 DVDD.n2575 DVDD.n2254 0.00962857
R7274 DVDD.n2571 DVDD.n2254 0.00962857
R7275 DVDD.n2571 DVDD.n2256 0.00962857
R7276 DVDD.n2567 DVDD.n2256 0.00962857
R7277 DVDD.n2567 DVDD.n2258 0.00962857
R7278 DVDD.n2272 DVDD.n2258 0.00962857
R7279 DVDD.n2278 DVDD.n2272 0.00962857
R7280 DVDD.n2278 DVDD.n2270 0.00962857
R7281 DVDD.n2282 DVDD.n2270 0.00962857
R7282 DVDD.n2282 DVDD.n2268 0.00962857
R7283 DVDD.n2289 DVDD.n2268 0.00962857
R7284 DVDD.n2289 DVDD.n2265 0.00962857
R7285 DVDD.n2556 DVDD.n2265 0.00962857
R7286 DVDD.n2556 DVDD.n2266 0.00962857
R7287 DVDD.n2552 DVDD.n2266 0.00962857
R7288 DVDD.n2552 DVDD.n2293 0.00962857
R7289 DVDD.n2548 DVDD.n2293 0.00962857
R7290 DVDD.n2548 DVDD.n2296 0.00962857
R7291 DVDD.n2544 DVDD.n2296 0.00962857
R7292 DVDD.n2544 DVDD.n2298 0.00962857
R7293 DVDD.n2302 DVDD.n2298 0.00962857
R7294 DVDD.n2529 DVDD.n2302 0.00962857
R7295 DVDD.n2529 DVDD.n2303 0.00962857
R7296 DVDD.n2525 DVDD.n2303 0.00962857
R7297 DVDD.n2525 DVDD.n2306 0.00962857
R7298 DVDD.n2521 DVDD.n2306 0.00962857
R7299 DVDD.n2521 DVDD.n2308 0.00962857
R7300 DVDD.n2517 DVDD.n2308 0.00962857
R7301 DVDD.n2517 DVDD.n2310 0.00962857
R7302 DVDD.n2513 DVDD.n2310 0.00962857
R7303 DVDD.n2513 DVDD.n2312 0.00962857
R7304 DVDD.n2509 DVDD.n2312 0.00962857
R7305 DVDD.n2509 DVDD.n2314 0.00962857
R7306 DVDD.n2505 DVDD.n2314 0.00962857
R7307 DVDD.n2505 DVDD.n2316 0.00962857
R7308 DVDD.n2501 DVDD.n2316 0.00962857
R7309 DVDD.n2501 DVDD.n2318 0.00962857
R7310 DVDD.n2497 DVDD.n2318 0.00962857
R7311 DVDD.n2497 DVDD.n2320 0.00962857
R7312 DVDD.n2493 DVDD.n2320 0.00962857
R7313 DVDD.n2493 DVDD.n2322 0.00962857
R7314 DVDD.n2337 DVDD.n2322 0.00962857
R7315 DVDD.n2338 DVDD.n2337 0.00962857
R7316 DVDD.n2344 DVDD.n2338 0.00962857
R7317 DVDD.n2344 DVDD.n2334 0.00962857
R7318 DVDD.n2348 DVDD.n2334 0.00962857
R7319 DVDD.n2348 DVDD.n2332 0.00962857
R7320 DVDD.n2355 DVDD.n2332 0.00962857
R7321 DVDD.n2355 DVDD.n2329 0.00962857
R7322 DVDD.n2481 DVDD.n2329 0.00962857
R7323 DVDD.n2481 DVDD.n2330 0.00962857
R7324 DVDD.n2477 DVDD.n2330 0.00962857
R7325 DVDD.n2477 DVDD.n2359 0.00962857
R7326 DVDD.n2473 DVDD.n2359 0.00962857
R7327 DVDD.n2473 DVDD.n2362 0.00962857
R7328 DVDD.n2469 DVDD.n2362 0.00962857
R7329 DVDD.n2469 DVDD.n2364 0.00962857
R7330 DVDD.n2368 DVDD.n2364 0.00962857
R7331 DVDD.n2454 DVDD.n2368 0.00962857
R7332 DVDD.n2454 DVDD.n2369 0.00962857
R7333 DVDD.n2450 DVDD.n2369 0.00962857
R7334 DVDD.n2450 DVDD.n2372 0.00962857
R7335 DVDD.n2446 DVDD.n2372 0.00962857
R7336 DVDD.n2446 DVDD.n2374 0.00962857
R7337 DVDD.n2442 DVDD.n2374 0.00962857
R7338 DVDD.n2442 DVDD.n2376 0.00962857
R7339 DVDD.n2438 DVDD.n2376 0.00962857
R7340 DVDD.n2438 DVDD.n2378 0.00962857
R7341 DVDD.n2434 DVDD.n2378 0.00962857
R7342 DVDD.n2434 DVDD.n2380 0.00962857
R7343 DVDD.n2430 DVDD.n2380 0.00962857
R7344 DVDD.n2430 DVDD.n2382 0.00962857
R7345 DVDD.n2426 DVDD.n2382 0.00962857
R7346 DVDD.n2426 DVDD.n2384 0.00962857
R7347 DVDD.n2422 DVDD.n2384 0.00962857
R7348 DVDD.n2422 DVDD.n2386 0.00962857
R7349 DVDD.n2418 DVDD.n2386 0.00962857
R7350 DVDD.n2418 DVDD.n2388 0.00962857
R7351 DVDD.n2414 DVDD.n2388 0.00962857
R7352 DVDD.n2414 DVDD.n2390 0.00962857
R7353 DVDD.n2410 DVDD.n2390 0.00962857
R7354 DVDD.n2410 DVDD.n2392 0.00962857
R7355 DVDD.n2406 DVDD.n2392 0.00962857
R7356 DVDD.n2406 DVDD.n2394 0.00962857
R7357 DVDD.n2402 DVDD.n2394 0.00962857
R7358 DVDD.n2402 DVDD.n2396 0.00962857
R7359 DVDD.n2590 DVDD.n2205 0.00962857
R7360 DVDD.n2590 DVDD.n2589 0.00962857
R7361 DVDD.n2589 DVDD.n2588 0.00962857
R7362 DVDD.n2588 DVDD.n2247 0.00962857
R7363 DVDD.n2582 DVDD.n2247 0.00962857
R7364 DVDD.n2582 DVDD.n2581 0.00962857
R7365 DVDD.n2581 DVDD.n2580 0.00962857
R7366 DVDD.n2580 DVDD.n2251 0.00962857
R7367 DVDD.n2574 DVDD.n2251 0.00962857
R7368 DVDD.n2574 DVDD.n2573 0.00962857
R7369 DVDD.n2573 DVDD.n2572 0.00962857
R7370 DVDD.n2566 DVDD.n2259 0.00962857
R7371 DVDD.n2273 DVDD.n2260 0.00962857
R7372 DVDD.n2277 DVDD.n2273 0.00962857
R7373 DVDD.n2283 DVDD.n2269 0.00962857
R7374 DVDD.n2284 DVDD.n2283 0.00962857
R7375 DVDD.n2288 DVDD.n2284 0.00962857
R7376 DVDD.n2551 DVDD.n2294 0.00962857
R7377 DVDD.n2551 DVDD.n2550 0.00962857
R7378 DVDD.n2550 DVDD.n2549 0.00962857
R7379 DVDD.n2543 DVDD.n2299 0.00962857
R7380 DVDD.n2543 DVDD.n2542 0.00962857
R7381 DVDD.n2530 DVDD.n2301 0.00962857
R7382 DVDD.n2524 DVDD.n2301 0.00962857
R7383 DVDD.n2524 DVDD.n2523 0.00962857
R7384 DVDD.n2523 DVDD.n2522 0.00962857
R7385 DVDD.n2522 DVDD.n2307 0.00962857
R7386 DVDD.n2516 DVDD.n2307 0.00962857
R7387 DVDD.n2516 DVDD.n2515 0.00962857
R7388 DVDD.n2515 DVDD.n2514 0.00962857
R7389 DVDD.n2514 DVDD.n2311 0.00962857
R7390 DVDD.n2508 DVDD.n2311 0.00962857
R7391 DVDD.n2508 DVDD.n2507 0.00962857
R7392 DVDD.n2507 DVDD.n2506 0.00962857
R7393 DVDD.n2506 DVDD.n2315 0.00962857
R7394 DVDD.n2500 DVDD.n2315 0.00962857
R7395 DVDD.n2500 DVDD.n2499 0.00962857
R7396 DVDD.n2499 DVDD.n2498 0.00962857
R7397 DVDD.n2498 DVDD.n2319 0.00962857
R7398 DVDD.n2492 DVDD.n2491 0.00962857
R7399 DVDD.n2339 DVDD.n2324 0.00962857
R7400 DVDD.n2343 DVDD.n2339 0.00962857
R7401 DVDD.n2349 DVDD.n2333 0.00962857
R7402 DVDD.n2350 DVDD.n2349 0.00962857
R7403 DVDD.n2354 DVDD.n2350 0.00962857
R7404 DVDD.n2476 DVDD.n2360 0.00962857
R7405 DVDD.n2476 DVDD.n2475 0.00962857
R7406 DVDD.n2475 DVDD.n2474 0.00962857
R7407 DVDD.n2468 DVDD.n2365 0.00962857
R7408 DVDD.n2468 DVDD.n2467 0.00962857
R7409 DVDD.n2455 DVDD.n2367 0.00962857
R7410 DVDD.n2449 DVDD.n2367 0.00962857
R7411 DVDD.n2449 DVDD.n2448 0.00962857
R7412 DVDD.n2448 DVDD.n2447 0.00962857
R7413 DVDD.n2447 DVDD.n2373 0.00962857
R7414 DVDD.n2441 DVDD.n2373 0.00962857
R7415 DVDD.n2441 DVDD.n2440 0.00962857
R7416 DVDD.n2440 DVDD.n2439 0.00962857
R7417 DVDD.n2439 DVDD.n2377 0.00962857
R7418 DVDD.n2433 DVDD.n2377 0.00962857
R7419 DVDD.n2433 DVDD.n2432 0.00962857
R7420 DVDD.n2432 DVDD.n2431 0.00962857
R7421 DVDD.n2431 DVDD.n2381 0.00962857
R7422 DVDD.n2425 DVDD.n2381 0.00962857
R7423 DVDD.n2425 DVDD.n2424 0.00962857
R7424 DVDD.n2424 DVDD.n2423 0.00962857
R7425 DVDD.n2423 DVDD.n2385 0.00962857
R7426 DVDD.n2417 DVDD.n2385 0.00962857
R7427 DVDD.n2417 DVDD.n2416 0.00962857
R7428 DVDD.n2416 DVDD.n2415 0.00962857
R7429 DVDD.n2415 DVDD.n2389 0.00962857
R7430 DVDD.n2409 DVDD.n2389 0.00962857
R7431 DVDD.n2409 DVDD.n2408 0.00962857
R7432 DVDD.n2408 DVDD.n2407 0.00962857
R7433 DVDD.n2407 DVDD.n2393 0.00962857
R7434 DVDD.n2401 DVDD.n2393 0.00962857
R7435 DVDD.n2401 DVDD.n2400 0.00962857
R7436 DVDD.n2612 DVDD.n2611 0.00962857
R7437 DVDD.n2611 DVDD.n2167 0.00962857
R7438 DVDD.n2623 DVDD.n2167 0.00962857
R7439 DVDD.n2623 DVDD.n2165 0.00962857
R7440 DVDD.n2627 DVDD.n2165 0.00962857
R7441 DVDD.n2627 DVDD.n2163 0.00962857
R7442 DVDD.n2631 DVDD.n2163 0.00962857
R7443 DVDD.n2631 DVDD.n2161 0.00962857
R7444 DVDD.n2635 DVDD.n2161 0.00962857
R7445 DVDD.n2635 DVDD.n2159 0.00962857
R7446 DVDD.n2639 DVDD.n2159 0.00962857
R7447 DVDD.n2639 DVDD.n2157 0.00962857
R7448 DVDD.n2643 DVDD.n2157 0.00962857
R7449 DVDD.n2643 DVDD.n2155 0.00962857
R7450 DVDD.n2647 DVDD.n2155 0.00962857
R7451 DVDD.n2647 DVDD.n2153 0.00962857
R7452 DVDD.n2651 DVDD.n2153 0.00962857
R7453 DVDD.n2651 DVDD.n2151 0.00962857
R7454 DVDD.n2655 DVDD.n2151 0.00962857
R7455 DVDD.n2655 DVDD.n2149 0.00962857
R7456 DVDD.n2659 DVDD.n2149 0.00962857
R7457 DVDD.n2659 DVDD.n2147 0.00962857
R7458 DVDD.n2663 DVDD.n2147 0.00962857
R7459 DVDD.n2663 DVDD.n2145 0.00962857
R7460 DVDD.n2667 DVDD.n2145 0.00962857
R7461 DVDD.n2667 DVDD.n2143 0.00962857
R7462 DVDD.n2675 DVDD.n2143 0.00962857
R7463 DVDD.n2675 DVDD.n2141 0.00962857
R7464 DVDD.n2679 DVDD.n2141 0.00962857
R7465 DVDD.n2679 DVDD.n2139 0.00962857
R7466 DVDD.n2866 DVDD.n2139 0.00962857
R7467 DVDD.n2866 DVDD.n2137 0.00962857
R7468 DVDD.n2870 DVDD.n2137 0.00962857
R7469 DVDD.n2870 DVDD.n2135 0.00962857
R7470 DVDD.n2874 DVDD.n2135 0.00962857
R7471 DVDD.n2874 DVDD.n2133 0.00962857
R7472 DVDD.n2878 DVDD.n2133 0.00962857
R7473 DVDD.n2878 DVDD.n2131 0.00962857
R7474 DVDD.n2882 DVDD.n2131 0.00962857
R7475 DVDD.n2882 DVDD.n2129 0.00962857
R7476 DVDD.n2886 DVDD.n2129 0.00962857
R7477 DVDD.n2886 DVDD.n2127 0.00962857
R7478 DVDD.n2890 DVDD.n2127 0.00962857
R7479 DVDD.n2890 DVDD.n2125 0.00962857
R7480 DVDD.n2894 DVDD.n2125 0.00962857
R7481 DVDD.n2894 DVDD.n2123 0.00962857
R7482 DVDD.n2898 DVDD.n2123 0.00962857
R7483 DVDD.n2898 DVDD.n2121 0.00962857
R7484 DVDD.n2902 DVDD.n2121 0.00962857
R7485 DVDD.n2902 DVDD.n2119 0.00962857
R7486 DVDD.n2906 DVDD.n2119 0.00962857
R7487 DVDD.n2906 DVDD.n2117 0.00962857
R7488 DVDD.n2910 DVDD.n2117 0.00962857
R7489 DVDD.n2910 DVDD.n2115 0.00962857
R7490 DVDD.n2914 DVDD.n2115 0.00962857
R7491 DVDD.n2914 DVDD.n2113 0.00962857
R7492 DVDD.n2918 DVDD.n2113 0.00962857
R7493 DVDD.n2918 DVDD.n2111 0.00962857
R7494 DVDD.n2922 DVDD.n2111 0.00962857
R7495 DVDD.n2922 DVDD.n2109 0.00962857
R7496 DVDD.n2926 DVDD.n2109 0.00962857
R7497 DVDD.n2926 DVDD.n2107 0.00962857
R7498 DVDD.n2930 DVDD.n2107 0.00962857
R7499 DVDD.n2930 DVDD.n2105 0.00962857
R7500 DVDD.n2934 DVDD.n2105 0.00962857
R7501 DVDD.n2934 DVDD.n2103 0.00962857
R7502 DVDD.n2938 DVDD.n2103 0.00962857
R7503 DVDD.n2938 DVDD.n2100 0.00962857
R7504 DVDD.n2943 DVDD.n2100 0.00962857
R7505 DVDD.n2943 DVDD.n2101 0.00962857
R7506 DVDD.n2101 DVDD.n2087 0.00962857
R7507 DVDD.n2950 DVDD.n2087 0.00962857
R7508 DVDD.n2950 DVDD.n2085 0.00962857
R7509 DVDD.n2954 DVDD.n2085 0.00962857
R7510 DVDD.n2954 DVDD.n2083 0.00962857
R7511 DVDD.n2958 DVDD.n2083 0.00962857
R7512 DVDD.n2958 DVDD.n2080 0.00962857
R7513 DVDD.n3020 DVDD.n2080 0.00962857
R7514 DVDD.n3020 DVDD.n2081 0.00962857
R7515 DVDD.n3016 DVDD.n2081 0.00962857
R7516 DVDD.n3016 DVDD.n2962 0.00962857
R7517 DVDD.n3012 DVDD.n2962 0.00962857
R7518 DVDD.n3012 DVDD.n2964 0.00962857
R7519 DVDD.n3008 DVDD.n2964 0.00962857
R7520 DVDD.n3008 DVDD.n2966 0.00962857
R7521 DVDD.n3004 DVDD.n2966 0.00962857
R7522 DVDD.n3004 DVDD.n2968 0.00962857
R7523 DVDD.n3000 DVDD.n2968 0.00962857
R7524 DVDD.n3000 DVDD.n2970 0.00962857
R7525 DVDD.n2996 DVDD.n2970 0.00962857
R7526 DVDD.n2996 DVDD.n2972 0.00962857
R7527 DVDD.n2992 DVDD.n2972 0.00962857
R7528 DVDD.n2992 DVDD.n2974 0.00962857
R7529 DVDD.n2988 DVDD.n2974 0.00962857
R7530 DVDD.n2988 DVDD.n2976 0.00962857
R7531 DVDD.n2984 DVDD.n2976 0.00962857
R7532 DVDD.n2984 DVDD.n2978 0.00962857
R7533 DVDD.n2622 DVDD.n2621 0.00962857
R7534 DVDD.n2622 DVDD.n2164 0.00962857
R7535 DVDD.n2628 DVDD.n2164 0.00962857
R7536 DVDD.n2629 DVDD.n2628 0.00962857
R7537 DVDD.n2630 DVDD.n2629 0.00962857
R7538 DVDD.n2630 DVDD.n2160 0.00962857
R7539 DVDD.n2636 DVDD.n2160 0.00962857
R7540 DVDD.n2637 DVDD.n2636 0.00962857
R7541 DVDD.n2638 DVDD.n2637 0.00962857
R7542 DVDD.n2638 DVDD.n2156 0.00962857
R7543 DVDD.n2644 DVDD.n2156 0.00962857
R7544 DVDD.n2645 DVDD.n2644 0.00962857
R7545 DVDD.n2646 DVDD.n2645 0.00962857
R7546 DVDD.n2646 DVDD.n2152 0.00962857
R7547 DVDD.n2652 DVDD.n2152 0.00962857
R7548 DVDD.n2653 DVDD.n2652 0.00962857
R7549 DVDD.n2654 DVDD.n2653 0.00962857
R7550 DVDD.n2654 DVDD.n2148 0.00962857
R7551 DVDD.n2660 DVDD.n2148 0.00962857
R7552 DVDD.n2661 DVDD.n2660 0.00962857
R7553 DVDD.n2662 DVDD.n2661 0.00962857
R7554 DVDD.n2662 DVDD.n2144 0.00962857
R7555 DVDD.n2668 DVDD.n2144 0.00962857
R7556 DVDD.n2674 DVDD.n2673 0.00962857
R7557 DVDD.n2674 DVDD.n2140 0.00962857
R7558 DVDD.n2680 DVDD.n2140 0.00962857
R7559 DVDD.n2681 DVDD.n2680 0.00962857
R7560 DVDD.n2872 DVDD.n2871 0.00962857
R7561 DVDD.n2873 DVDD.n2872 0.00962857
R7562 DVDD.n2873 DVDD.n2132 0.00962857
R7563 DVDD.n2879 DVDD.n2132 0.00962857
R7564 DVDD.n2880 DVDD.n2879 0.00962857
R7565 DVDD.n2881 DVDD.n2880 0.00962857
R7566 DVDD.n2881 DVDD.n2128 0.00962857
R7567 DVDD.n2887 DVDD.n2128 0.00962857
R7568 DVDD.n2888 DVDD.n2887 0.00962857
R7569 DVDD.n2889 DVDD.n2888 0.00962857
R7570 DVDD.n2889 DVDD.n2124 0.00962857
R7571 DVDD.n2895 DVDD.n2124 0.00962857
R7572 DVDD.n2896 DVDD.n2895 0.00962857
R7573 DVDD.n2897 DVDD.n2896 0.00962857
R7574 DVDD.n2897 DVDD.n2120 0.00962857
R7575 DVDD.n2903 DVDD.n2120 0.00962857
R7576 DVDD.n2904 DVDD.n2903 0.00962857
R7577 DVDD.n2905 DVDD.n2904 0.00962857
R7578 DVDD.n2905 DVDD.n2116 0.00962857
R7579 DVDD.n2911 DVDD.n2116 0.00962857
R7580 DVDD.n2912 DVDD.n2911 0.00962857
R7581 DVDD.n2913 DVDD.n2912 0.00962857
R7582 DVDD.n2913 DVDD.n2112 0.00962857
R7583 DVDD.n2919 DVDD.n2112 0.00962857
R7584 DVDD.n2920 DVDD.n2919 0.00962857
R7585 DVDD.n2921 DVDD.n2920 0.00962857
R7586 DVDD.n2921 DVDD.n2108 0.00962857
R7587 DVDD.n2927 DVDD.n2108 0.00962857
R7588 DVDD.n2928 DVDD.n2927 0.00962857
R7589 DVDD.n2929 DVDD.n2928 0.00962857
R7590 DVDD.n2929 DVDD.n2104 0.00962857
R7591 DVDD.n2935 DVDD.n2104 0.00962857
R7592 DVDD.n2936 DVDD.n2935 0.00962857
R7593 DVDD.n2937 DVDD.n2936 0.00962857
R7594 DVDD.n2937 DVDD.n2099 0.00962857
R7595 DVDD.n2949 DVDD.n2948 0.00962857
R7596 DVDD.n2949 DVDD.n2084 0.00962857
R7597 DVDD.n2955 DVDD.n2084 0.00962857
R7598 DVDD.n2956 DVDD.n2955 0.00962857
R7599 DVDD.n2957 DVDD.n2956 0.00962857
R7600 DVDD.n2957 DVDD.n2078 0.00962857
R7601 DVDD.n3021 DVDD.n2079 0.00962857
R7602 DVDD.n3015 DVDD.n2079 0.00962857
R7603 DVDD.n3015 DVDD.n3014 0.00962857
R7604 DVDD.n3014 DVDD.n3013 0.00962857
R7605 DVDD.n3013 DVDD.n2963 0.00962857
R7606 DVDD.n3007 DVDD.n2963 0.00962857
R7607 DVDD.n3007 DVDD.n3006 0.00962857
R7608 DVDD.n3006 DVDD.n3005 0.00962857
R7609 DVDD.n3005 DVDD.n2967 0.00962857
R7610 DVDD.n2999 DVDD.n2967 0.00962857
R7611 DVDD.n2999 DVDD.n2998 0.00962857
R7612 DVDD.n2998 DVDD.n2997 0.00962857
R7613 DVDD.n2997 DVDD.n2971 0.00962857
R7614 DVDD.n2991 DVDD.n2971 0.00962857
R7615 DVDD.n2991 DVDD.n2990 0.00962857
R7616 DVDD.n2990 DVDD.n2989 0.00962857
R7617 DVDD.n2989 DVDD.n2975 0.00962857
R7618 DVDD.n2983 DVDD.n2975 0.00962857
R7619 DVDD.n2983 DVDD.n2982 0.00962857
R7620 DVDD.n1571 DVDD.n1205 0.00962857
R7621 DVDD.n1571 DVDD.n1206 0.00962857
R7622 DVDD.n1567 DVDD.n1206 0.00962857
R7623 DVDD.n1567 DVDD.n1208 0.00962857
R7624 DVDD.n1563 DVDD.n1208 0.00962857
R7625 DVDD.n1563 DVDD.n1211 0.00962857
R7626 DVDD.n1559 DVDD.n1211 0.00962857
R7627 DVDD.n1559 DVDD.n1213 0.00962857
R7628 DVDD.n1224 DVDD.n1213 0.00962857
R7629 DVDD.n1552 DVDD.n1224 0.00962857
R7630 DVDD.n1552 DVDD.n1225 0.00962857
R7631 DVDD.n1548 DVDD.n1225 0.00962857
R7632 DVDD.n1548 DVDD.n1228 0.00962857
R7633 DVDD.n1544 DVDD.n1228 0.00962857
R7634 DVDD.n1544 DVDD.n1230 0.00962857
R7635 DVDD.n1540 DVDD.n1230 0.00962857
R7636 DVDD.n1540 DVDD.n1232 0.00962857
R7637 DVDD.n1536 DVDD.n1232 0.00962857
R7638 DVDD.n1536 DVDD.n1234 0.00962857
R7639 DVDD.n1532 DVDD.n1234 0.00962857
R7640 DVDD.n1532 DVDD.n1236 0.00962857
R7641 DVDD.n1528 DVDD.n1236 0.00962857
R7642 DVDD.n1528 DVDD.n1238 0.00962857
R7643 DVDD.n1524 DVDD.n1238 0.00962857
R7644 DVDD.n1524 DVDD.n1240 0.00962857
R7645 DVDD.n1520 DVDD.n1240 0.00962857
R7646 DVDD.n1520 DVDD.n1242 0.00962857
R7647 DVDD.n1516 DVDD.n1242 0.00962857
R7648 DVDD.n1516 DVDD.n1244 0.00962857
R7649 DVDD.n1512 DVDD.n1244 0.00962857
R7650 DVDD.n1512 DVDD.n1246 0.00962857
R7651 DVDD.n1508 DVDD.n1246 0.00962857
R7652 DVDD.n1508 DVDD.n1248 0.00962857
R7653 DVDD.n1504 DVDD.n1248 0.00962857
R7654 DVDD.n1504 DVDD.n1250 0.00962857
R7655 DVDD.n1500 DVDD.n1250 0.00962857
R7656 DVDD.n1500 DVDD.n1252 0.00962857
R7657 DVDD.n1496 DVDD.n1252 0.00962857
R7658 DVDD.n1496 DVDD.n1254 0.00962857
R7659 DVDD.n1492 DVDD.n1254 0.00962857
R7660 DVDD.n1492 DVDD.n1256 0.00962857
R7661 DVDD.n1488 DVDD.n1256 0.00962857
R7662 DVDD.n1488 DVDD.n1258 0.00962857
R7663 DVDD.n1484 DVDD.n1258 0.00962857
R7664 DVDD.n1484 DVDD.n1260 0.00962857
R7665 DVDD.n1480 DVDD.n1260 0.00962857
R7666 DVDD.n1480 DVDD.n1262 0.00962857
R7667 DVDD.n1476 DVDD.n1262 0.00962857
R7668 DVDD.n1476 DVDD.n1264 0.00962857
R7669 DVDD.n1472 DVDD.n1264 0.00962857
R7670 DVDD.n1472 DVDD.n1266 0.00962857
R7671 DVDD.n1468 DVDD.n1266 0.00962857
R7672 DVDD.n1468 DVDD.n1268 0.00962857
R7673 DVDD.n1464 DVDD.n1268 0.00962857
R7674 DVDD.n1464 DVDD.n1270 0.00962857
R7675 DVDD.n1460 DVDD.n1270 0.00962857
R7676 DVDD.n1460 DVDD.n1272 0.00962857
R7677 DVDD.n1456 DVDD.n1272 0.00962857
R7678 DVDD.n1456 DVDD.n1274 0.00962857
R7679 DVDD.n1452 DVDD.n1274 0.00962857
R7680 DVDD.n1452 DVDD.n1276 0.00962857
R7681 DVDD.n1448 DVDD.n1276 0.00962857
R7682 DVDD.n1448 DVDD.n1278 0.00962857
R7683 DVDD.n1444 DVDD.n1278 0.00962857
R7684 DVDD.n1444 DVDD.n1280 0.00962857
R7685 DVDD.n1440 DVDD.n1280 0.00962857
R7686 DVDD.n1440 DVDD.n1282 0.00962857
R7687 DVDD.n1436 DVDD.n1282 0.00962857
R7688 DVDD.n1436 DVDD.n1284 0.00962857
R7689 DVDD.n1432 DVDD.n1284 0.00962857
R7690 DVDD.n1432 DVDD.n1286 0.00962857
R7691 DVDD.n1428 DVDD.n1286 0.00962857
R7692 DVDD.n1428 DVDD.n1288 0.00962857
R7693 DVDD.n1424 DVDD.n1288 0.00962857
R7694 DVDD.n1424 DVDD.n1290 0.00962857
R7695 DVDD.n1420 DVDD.n1290 0.00962857
R7696 DVDD.n1420 DVDD.n1292 0.00962857
R7697 DVDD.n1416 DVDD.n1292 0.00962857
R7698 DVDD.n1416 DVDD.n1294 0.00962857
R7699 DVDD.n1412 DVDD.n1294 0.00962857
R7700 DVDD.n1412 DVDD.n1296 0.00962857
R7701 DVDD.n1408 DVDD.n1296 0.00962857
R7702 DVDD.n1408 DVDD.n1298 0.00962857
R7703 DVDD.n1404 DVDD.n1298 0.00962857
R7704 DVDD.n1404 DVDD.n1300 0.00962857
R7705 DVDD.n1400 DVDD.n1300 0.00962857
R7706 DVDD.n1400 DVDD.n1302 0.00962857
R7707 DVDD.n1396 DVDD.n1302 0.00962857
R7708 DVDD.n1396 DVDD.n1304 0.00962857
R7709 DVDD.n1347 DVDD.n1304 0.00962857
R7710 DVDD.n1350 DVDD.n1347 0.00962857
R7711 DVDD.n1350 DVDD.n1345 0.00962857
R7712 DVDD.n1354 DVDD.n1345 0.00962857
R7713 DVDD.n1354 DVDD.n1343 0.00962857
R7714 DVDD.n1358 DVDD.n1343 0.00962857
R7715 DVDD.n1362 DVDD.n1361 0.00962857
R7716 DVDD.n1566 DVDD.n1209 0.00962857
R7717 DVDD.n1566 DVDD.n1565 0.00962857
R7718 DVDD.n1565 DVDD.n1564 0.00962857
R7719 DVDD.n1564 DVDD.n1210 0.00962857
R7720 DVDD.n1558 DVDD.n1210 0.00962857
R7721 DVDD.n1558 DVDD.n1557 0.00962857
R7722 DVDD.n1553 DVDD.n1223 0.00962857
R7723 DVDD.n1547 DVDD.n1223 0.00962857
R7724 DVDD.n1547 DVDD.n1546 0.00962857
R7725 DVDD.n1546 DVDD.n1545 0.00962857
R7726 DVDD.n1545 DVDD.n1229 0.00962857
R7727 DVDD.n1539 DVDD.n1229 0.00962857
R7728 DVDD.n1539 DVDD.n1538 0.00962857
R7729 DVDD.n1538 DVDD.n1537 0.00962857
R7730 DVDD.n1537 DVDD.n1233 0.00962857
R7731 DVDD.n1531 DVDD.n1233 0.00962857
R7732 DVDD.n1531 DVDD.n1530 0.00962857
R7733 DVDD.n1530 DVDD.n1529 0.00962857
R7734 DVDD.n1529 DVDD.n1237 0.00962857
R7735 DVDD.n1523 DVDD.n1237 0.00962857
R7736 DVDD.n1523 DVDD.n1522 0.00962857
R7737 DVDD.n1522 DVDD.n1521 0.00962857
R7738 DVDD.n1521 DVDD.n1241 0.00962857
R7739 DVDD.n1515 DVDD.n1241 0.00962857
R7740 DVDD.n1515 DVDD.n1514 0.00962857
R7741 DVDD.n1514 DVDD.n1513 0.00962857
R7742 DVDD.n1513 DVDD.n1245 0.00962857
R7743 DVDD.n1507 DVDD.n1245 0.00962857
R7744 DVDD.n1507 DVDD.n1506 0.00962857
R7745 DVDD.n1506 DVDD.n1505 0.00962857
R7746 DVDD.n1505 DVDD.n1249 0.00962857
R7747 DVDD.n1499 DVDD.n1249 0.00962857
R7748 DVDD.n1499 DVDD.n1498 0.00962857
R7749 DVDD.n1498 DVDD.n1497 0.00962857
R7750 DVDD.n1497 DVDD.n1253 0.00962857
R7751 DVDD.n1491 DVDD.n1253 0.00962857
R7752 DVDD.n1491 DVDD.n1490 0.00962857
R7753 DVDD.n1490 DVDD.n1489 0.00962857
R7754 DVDD.n1489 DVDD.n1257 0.00962857
R7755 DVDD.n1483 DVDD.n1257 0.00962857
R7756 DVDD.n1483 DVDD.n1482 0.00962857
R7757 DVDD.n1482 DVDD.n1481 0.00962857
R7758 DVDD.n1481 DVDD.n1261 0.00962857
R7759 DVDD.n1475 DVDD.n1261 0.00962857
R7760 DVDD.n1475 DVDD.n1474 0.00962857
R7761 DVDD.n1474 DVDD.n1473 0.00962857
R7762 DVDD.n1473 DVDD.n1265 0.00962857
R7763 DVDD.n1467 DVDD.n1265 0.00962857
R7764 DVDD.n1467 DVDD.n1466 0.00962857
R7765 DVDD.n1466 DVDD.n1465 0.00962857
R7766 DVDD.n1465 DVDD.n1269 0.00962857
R7767 DVDD.n1459 DVDD.n1269 0.00962857
R7768 DVDD.n1459 DVDD.n1458 0.00962857
R7769 DVDD.n1458 DVDD.n1457 0.00962857
R7770 DVDD.n1457 DVDD.n1273 0.00962857
R7771 DVDD.n1451 DVDD.n1273 0.00962857
R7772 DVDD.n1451 DVDD.n1450 0.00962857
R7773 DVDD.n1450 DVDD.n1449 0.00962857
R7774 DVDD.n1449 DVDD.n1277 0.00962857
R7775 DVDD.n1443 DVDD.n1277 0.00962857
R7776 DVDD.n1443 DVDD.n1442 0.00962857
R7777 DVDD.n1442 DVDD.n1441 0.00962857
R7778 DVDD.n1441 DVDD.n1281 0.00962857
R7779 DVDD.n1435 DVDD.n1281 0.00962857
R7780 DVDD.n1435 DVDD.n1434 0.00962857
R7781 DVDD.n1434 DVDD.n1433 0.00962857
R7782 DVDD.n1433 DVDD.n1285 0.00962857
R7783 DVDD.n1427 DVDD.n1285 0.00962857
R7784 DVDD.n1427 DVDD.n1426 0.00962857
R7785 DVDD.n1426 DVDD.n1425 0.00962857
R7786 DVDD.n1425 DVDD.n1289 0.00962857
R7787 DVDD.n1419 DVDD.n1289 0.00962857
R7788 DVDD.n1419 DVDD.n1418 0.00962857
R7789 DVDD.n1418 DVDD.n1417 0.00962857
R7790 DVDD.n1417 DVDD.n1293 0.00962857
R7791 DVDD.n1411 DVDD.n1293 0.00962857
R7792 DVDD.n1411 DVDD.n1410 0.00962857
R7793 DVDD.n1410 DVDD.n1409 0.00962857
R7794 DVDD.n1409 DVDD.n1297 0.00962857
R7795 DVDD.n1403 DVDD.n1297 0.00962857
R7796 DVDD.n1403 DVDD.n1402 0.00962857
R7797 DVDD.n1402 DVDD.n1401 0.00962857
R7798 DVDD.n1401 DVDD.n1301 0.00962857
R7799 DVDD.n1348 DVDD.n1310 0.00962857
R7800 DVDD.n1349 DVDD.n1348 0.00962857
R7801 DVDD.n1349 DVDD.n1344 0.00962857
R7802 DVDD.n1355 DVDD.n1344 0.00962857
R7803 DVDD.n1356 DVDD.n1355 0.00962857
R7804 DVDD.n1357 DVDD.n1356 0.00962857
R7805 DVDD.n1337 DVDD.n1331 0.00956429
R7806 DVDD.n1364 DVDD.n1340 0.00956429
R7807 DVDD.n5424 DVDD.n333 0.00955202
R7808 DVDD.n3505 DVDD.n3175 0.00954891
R7809 DVDD.n3512 DVDD.n3511 0.00954891
R7810 DVDD.n3521 DVDD.n3162 0.00954891
R7811 DVDD.n3525 DVDD.n3155 0.00954891
R7812 DVDD.n86 DVDD.n85 0.00953114
R7813 DVDD.n5521 DVDD.n10 0.00948451
R7814 DVDD.n4691 DVDD.n977 0.00948451
R7815 DVDD.n3352 DVDD.n3351 0.00941892
R7816 DVDD.n3397 DVDD.n3396 0.00941892
R7817 DVDD.n5762 DVDD.n184 0.00935246
R7818 DVDD.n5220 DVDD.n490 0.00935246
R7819 DVDD.n646 DVDD.n620 0.00935246
R7820 DVDD.n846 DVDD.n709 0.00935246
R7821 DVDD.n4593 DVDD.n1014 0.00935246
R7822 DVDD.n5507 DVDD.n222 0.0093296
R7823 DVDD.n948 DVDD.n946 0.0093296
R7824 DVDD.n2695 DVDD.n2692 0.00930435
R7825 DVDD.n2572 DVDD.n2255 0.00917857
R7826 DVDD.n5930 DVDD.n70 0.0091747
R7827 DVDD.n5474 DVDD.n294 0.0091747
R7828 DVDD.n110 DVDD.n89 0.00908247
R7829 DVDD.n5913 DVDD.n94 0.00908247
R7830 DVDD.n5406 DVDD.n343 0.00908247
R7831 DVDD.n5417 DVDD.n5416 0.00908247
R7832 DVDD.n927 DVDD.n915 0.00908247
R7833 DVDD.n4709 DVDD.n942 0.00908247
R7834 DVDD.n257 DVDD.n235 0.00908247
R7835 DVDD.n244 DVDD.n228 0.00908247
R7836 DVDD.n2830 DVDD.n2094 0.00905
R7837 DVDD.n4676 DVDD.n4675 0.00903179
R7838 DVDD.n5539 DVDD.n5537 0.00901211
R7839 DVDD.n5809 DVDD.n159 0.00898361
R7840 DVDD.n5165 DVDD.n459 0.00898361
R7841 DVDD.n4972 DVDD.n681 0.00898361
R7842 DVDD.n790 DVDD.n749 0.00898361
R7843 DVDD.n4528 DVDD.n1082 0.00898361
R7844 DVDD.n2353 DVDD.n2327 0.00892143
R7845 DVDD.n2365 DVDD.n2361 0.00892143
R7846 DVDD.n5623 DVDD.n5604 0.00886489
R7847 DVDD.n5448 DVDD.n288 0.00886489
R7848 DVDD.n3135 DVDD.n3134 0.00881522
R7849 DVDD.n3581 DVDD.n3138 0.00881522
R7850 DVDD.n3440 DVDD.n3206 0.00881522
R7851 DVDD.n3465 DVDD.n3196 0.00881522
R7852 DVDD.n3475 DVDD.n3181 0.00881522
R7853 DVDD.n3558 DVDD.n3158 0.00881522
R7854 DVDD.n2531 DVDD.n2300 0.00879286
R7855 DVDD.n2945 DVDD.n2099 0.00879286
R7856 DVDD.n2944 DVDD.n2097 0.00879286
R7857 DVDD.n2947 DVDD.n2088 0.00879286
R7858 DVDD.n1556 DVDD.n1218 0.00879286
R7859 DVDD.n1554 DVDD.n1553 0.00879286
R7860 DVDD.n3090 DVDD.n2023 0.00868173
R7861 DVDD.n112 DVDD.n91 0.00861856
R7862 DVDD.n5908 DVDD.n93 0.00861856
R7863 DVDD.n5408 DVDD.n345 0.00861856
R7864 DVDD.n5411 DVDD.n347 0.00861856
R7865 DVDD.n933 DVDD.n917 0.00861856
R7866 DVDD.n952 DVDD.n924 0.00861856
R7867 DVDD.n5668 DVDD.n236 0.00861856
R7868 DVDD.n252 DVDD.n230 0.00861856
R7869 DVDD.n5746 DVDD.n186 0.00861475
R7870 DVDD.n5236 DVDD.n565 0.00861475
R7871 DVDD.n630 DVDD.n622 0.00861475
R7872 DVDD.n862 DVDD.n725 0.00861475
R7873 DVDD.n4609 DVDD.n1056 0.00861475
R7874 DVDD.n2826 DVDD.n2091 0.0086
R7875 DVDD.n5640 DVDD.n5568 0.00855508
R7876 DVDD.n5465 DVDD.n277 0.00855508
R7877 DVDD.n2597 DVDD.n2198 0.00853571
R7878 DVDD.n2601 DVDD.n2200 0.00853571
R7879 DVDD.n2323 DVDD.n2319 0.00853571
R7880 DVDD.n2613 DVDD.n2609 0.00853571
R7881 DVDD.n2620 DVDD.n2168 0.00853571
R7882 DVDD.n2865 DVDD.n2682 0.00853571
R7883 DVDD.n2864 DVDD.n2688 0.00853571
R7884 DVDD.n2871 DVDD.n2136 0.00853571
R7885 DVDD.n3022 DVDD.n2078 0.00853571
R7886 DVDD.n4077 DVDD.n4076 0.0084875
R7887 DVDD.n4076 DVDD.n4046 0.0084875
R7888 DVDD.n4072 DVDD.n4046 0.0084875
R7889 DVDD.n4072 DVDD.n4048 0.0084875
R7890 DVDD.n4068 DVDD.n4048 0.0084875
R7891 DVDD.n4068 DVDD.n4051 0.0084875
R7892 DVDD.n4061 DVDD.n4051 0.0084875
R7893 DVDD.n4061 DVDD.n4058 0.0084875
R7894 DVDD.n4058 DVDD.n1723 0.0084875
R7895 DVDD.n4223 DVDD.n1723 0.0084875
R7896 DVDD.n1765 DVDD.n1727 0.0084875
R7897 DVDD.n1758 DVDD.n1727 0.0084875
R7898 DVDD.n1758 DVDD.n1731 0.0084875
R7899 DVDD.n1754 DVDD.n1731 0.0084875
R7900 DVDD.n1754 DVDD.n1733 0.0084875
R7901 DVDD.n1750 DVDD.n1733 0.0084875
R7902 DVDD.n1750 DVDD.n1736 0.0084875
R7903 DVDD.n1746 DVDD.n1736 0.0084875
R7904 DVDD.n1746 DVDD.n1738 0.0084875
R7905 DVDD.n4075 DVDD.n4042 0.0084875
R7906 DVDD.n4075 DVDD.n4074 0.0084875
R7907 DVDD.n4074 DVDD.n4073 0.0084875
R7908 DVDD.n4073 DVDD.n4047 0.0084875
R7909 DVDD.n1753 DVDD.n1734 0.0084875
R7910 DVDD.n1753 DVDD.n1752 0.0084875
R7911 DVDD.n1752 DVDD.n1751 0.0084875
R7912 DVDD.n1751 DVDD.n1735 0.0084875
R7913 DVDD.n1745 DVDD.n1735 0.0084875
R7914 DVDD.n1745 DVDD.n1744 0.0084875
R7915 DVDD.n3898 DVDD.n3897 0.0084875
R7916 DVDD.n3897 DVDD.n3896 0.0084875
R7917 DVDD.n3896 DVDD.n3871 0.0084875
R7918 DVDD.n3890 DVDD.n3871 0.0084875
R7919 DVDD.n3890 DVDD.n3889 0.0084875
R7920 DVDD.n3889 DVDD.n3888 0.0084875
R7921 DVDD.n3888 DVDD.n3876 0.0084875
R7922 DVDD.n3882 DVDD.n3876 0.0084875
R7923 DVDD.n3882 DVDD.n3881 0.0084875
R7924 DVDD.n3881 DVDD.n1794 0.0084875
R7925 DVDD.n4099 DVDD.n4098 0.0084875
R7926 DVDD.n4098 DVDD.n4097 0.0084875
R7927 DVDD.n4097 DVDD.n4034 0.0084875
R7928 DVDD.n4091 DVDD.n4034 0.0084875
R7929 DVDD.n4091 DVDD.n4090 0.0084875
R7930 DVDD.n4090 DVDD.n4089 0.0084875
R7931 DVDD.n4089 DVDD.n4038 0.0084875
R7932 DVDD.n4083 DVDD.n4038 0.0084875
R7933 DVDD.n4083 DVDD.n4082 0.0084875
R7934 DVDD.n3899 DVDD.n3870 0.0084875
R7935 DVDD.n3895 DVDD.n3870 0.0084875
R7936 DVDD.n3895 DVDD.n3872 0.0084875
R7937 DVDD.n3891 DVDD.n3872 0.0084875
R7938 DVDD.n3891 DVDD.n3875 0.0084875
R7939 DVDD.n3887 DVDD.n3875 0.0084875
R7940 DVDD.n3887 DVDD.n3877 0.0084875
R7941 DVDD.n3883 DVDD.n3877 0.0084875
R7942 DVDD.n3883 DVDD.n3880 0.0084875
R7943 DVDD.n3880 DVDD.n3879 0.0084875
R7944 DVDD.n4100 DVDD.n1793 0.0084875
R7945 DVDD.n4096 DVDD.n1793 0.0084875
R7946 DVDD.n4096 DVDD.n4035 0.0084875
R7947 DVDD.n4092 DVDD.n4035 0.0084875
R7948 DVDD.n4092 DVDD.n4037 0.0084875
R7949 DVDD.n4088 DVDD.n4037 0.0084875
R7950 DVDD.n4088 DVDD.n4039 0.0084875
R7951 DVDD.n4084 DVDD.n4039 0.0084875
R7952 DVDD.n4084 DVDD.n4041 0.0084875
R7953 DVDD.n3835 DVDD.n1828 0.0084875
R7954 DVDD.n3839 DVDD.n1828 0.0084875
R7955 DVDD.n3839 DVDD.n1826 0.0084875
R7956 DVDD.n3843 DVDD.n1826 0.0084875
R7957 DVDD.n3843 DVDD.n1824 0.0084875
R7958 DVDD.n3847 DVDD.n1824 0.0084875
R7959 DVDD.n3847 DVDD.n1822 0.0084875
R7960 DVDD.n3851 DVDD.n1822 0.0084875
R7961 DVDD.n3851 DVDD.n1820 0.0084875
R7962 DVDD.n3855 DVDD.n1820 0.0084875
R7963 DVDD.n3921 DVDD.n3858 0.0084875
R7964 DVDD.n3917 DVDD.n3858 0.0084875
R7965 DVDD.n3917 DVDD.n3860 0.0084875
R7966 DVDD.n3913 DVDD.n3860 0.0084875
R7967 DVDD.n3913 DVDD.n3862 0.0084875
R7968 DVDD.n3909 DVDD.n3862 0.0084875
R7969 DVDD.n3909 DVDD.n3864 0.0084875
R7970 DVDD.n3905 DVDD.n3864 0.0084875
R7971 DVDD.n3905 DVDD.n3866 0.0084875
R7972 DVDD.n4283 DVDD.n1669 0.0084875
R7973 DVDD.n4279 DVDD.n1669 0.0084875
R7974 DVDD.n4279 DVDD.n1672 0.0084875
R7975 DVDD.n4275 DVDD.n1672 0.0084875
R7976 DVDD.n4275 DVDD.n1674 0.0084875
R7977 DVDD.n4271 DVDD.n1674 0.0084875
R7978 DVDD.n4271 DVDD.n1676 0.0084875
R7979 DVDD.n4267 DVDD.n1676 0.0084875
R7980 DVDD.n4267 DVDD.n1678 0.0084875
R7981 DVDD.n4260 DVDD.n1678 0.0084875
R7982 DVDD.n3809 DVDD.n3807 0.0084875
R7983 DVDD.n3809 DVDD.n1839 0.0084875
R7984 DVDD.n3818 DVDD.n1839 0.0084875
R7985 DVDD.n3818 DVDD.n1837 0.0084875
R7986 DVDD.n3822 DVDD.n1837 0.0084875
R7987 DVDD.n3822 DVDD.n1835 0.0084875
R7988 DVDD.n3826 DVDD.n1835 0.0084875
R7989 DVDD.n3826 DVDD.n1833 0.0084875
R7990 DVDD.n3830 DVDD.n1833 0.0084875
R7991 DVDD.n3834 DVDD.n1827 0.0084875
R7992 DVDD.n3840 DVDD.n1827 0.0084875
R7993 DVDD.n3841 DVDD.n3840 0.0084875
R7994 DVDD.n3842 DVDD.n3841 0.0084875
R7995 DVDD.n3842 DVDD.n1823 0.0084875
R7996 DVDD.n3848 DVDD.n1823 0.0084875
R7997 DVDD.n3849 DVDD.n3848 0.0084875
R7998 DVDD.n3850 DVDD.n3849 0.0084875
R7999 DVDD.n3850 DVDD.n1819 0.0084875
R8000 DVDD.n3856 DVDD.n1819 0.0084875
R8001 DVDD.n3922 DVDD.n3857 0.0084875
R8002 DVDD.n3916 DVDD.n3857 0.0084875
R8003 DVDD.n3916 DVDD.n3915 0.0084875
R8004 DVDD.n3915 DVDD.n3914 0.0084875
R8005 DVDD.n3914 DVDD.n3861 0.0084875
R8006 DVDD.n3908 DVDD.n3861 0.0084875
R8007 DVDD.n3908 DVDD.n3907 0.0084875
R8008 DVDD.n3907 DVDD.n3906 0.0084875
R8009 DVDD.n3906 DVDD.n3865 0.0084875
R8010 DVDD.n4282 DVDD.n4281 0.0084875
R8011 DVDD.n4281 DVDD.n4280 0.0084875
R8012 DVDD.n4280 DVDD.n1671 0.0084875
R8013 DVDD.n4274 DVDD.n1671 0.0084875
R8014 DVDD.n4274 DVDD.n4273 0.0084875
R8015 DVDD.n4273 DVDD.n4272 0.0084875
R8016 DVDD.n3824 DVDD.n3823 0.0084875
R8017 DVDD.n3825 DVDD.n3824 0.0084875
R8018 DVDD.n3825 DVDD.n1832 0.0084875
R8019 DVDD.n3831 DVDD.n1832 0.0084875
R8020 DVDD.n5651 DVDD.n68 0.00840017
R8021 DVDD.n5477 DVDD.n270 0.00840017
R8022 DVDD.n2181 DVDD.n1897 0.00832155
R8023 DVDD.n4287 DVDD.n1666 0.00832155
R8024 DVDD.n2189 DVDD.n2174 0.00830425
R8025 DVDD.n3717 DVDD.n1890 0.00830425
R8026 DVDD.n3771 DVDD.n3755 0.00830425
R8027 DVDD.n4297 DVDD.n1660 0.00830425
R8028 DVDD.n968 DVDD.n966 0.00830347
R8029 DVDD.n5506 DVDD.n5504 0.00828547
R8030 DVDD.n2287 DVDD.n2263 0.00827857
R8031 DVDD.n2299 DVDD.n2295 0.00827857
R8032 DVDD.n5825 DVDD.n147 0.0082459
R8033 DVDD.n5181 DVDD.n457 0.0082459
R8034 DVDD.n4956 DVDD.n679 0.0082459
R8035 DVDD.n807 DVDD.n806 0.0082459
R8036 DVDD.n4512 DVDD.n1080 0.0082459
R8037 DVDD.n2456 DVDD.n2366 0.00815
R8038 DVDD.n3282 DVDD.n3270 0.00815
R8039 DVDD.n3293 DVDD.n3283 0.00815
R8040 DVDD.n3292 DVDD.n3228 0.00815
R8041 DVDD.n3289 DVDD.n3089 0.00815
R8042 DVDD.n3343 DVDD.n3097 0.00815
R8043 DVDD.n5636 DVDD.n52 0.00809036
R8044 DVDD.n5502 DVDD.n219 0.00809036
R8045 DVDD.n964 DVDD.n945 0.00809036
R8046 DVDD.n5461 DVDD.n314 0.00809036
R8047 DVDD.n3502 DVDD.n3176 0.00808152
R8048 DVDD.n3514 DVDD.n3170 0.00808152
R8049 DVDD.n3518 DVDD.n3161 0.00808152
R8050 DVDD.n3529 DVDD.n3154 0.00808152
R8051 DVDD.n930 DVDD.n264 0.00804054
R8052 DVDD.n951 DVDD.n264 0.00804054
R8053 DVDD.n5665 DVDD.n5663 0.00796988
R8054 DVDD.n5663 DVDD.n255 0.00796988
R8055 DVDD.n2672 DVDD.n2668 0.00795714
R8056 DVDD.n5525 DVDD.n25 0.00793546
R8057 DVDD.n4687 DVDD.n4652 0.00793546
R8058 DVDD.n1670 DVDD.n1665 0.0079044
R8059 DVDD.n2849 DVDD.n2685 0.00783696
R8060 DVDD DVDD.n2396 0.00782857
R8061 DVDD.n2400 DVDD 0.00782857
R8062 DVDD DVDD.n2978 0.00782857
R8063 DVDD.n2982 DVDD 0.00782857
R8064 DVDD.n1358 DVDD 0.00782857
R8065 DVDD.n1357 DVDD 0.00782857
R8066 DVDD.n3357 DVDD.n3308 0.0077973
R8067 DVDD.n3388 DVDD.n3233 0.0077973
R8068 DVDD.n5619 DVDD.n61 0.00778055
R8069 DVDD.n5444 DVDD.n304 0.00778055
R8070 DVDD.n2740 DVDD.n2739 0.00777531
R8071 DVDD.n2732 DVDD.n2725 0.00777531
R8072 DVDD.n2780 DVDD.n2722 0.00777531
R8073 DVDD.n2731 DVDD.n2721 0.00777531
R8074 DVDD.n2782 DVDD.n2728 0.00777531
R8075 DVDD.n2730 DVDD.n2720 0.00777531
R8076 DVDD.n2787 DVDD.n2729 0.00777531
R8077 DVDD.n2739 DVDD.n2723 0.00777531
R8078 DVDD.n2732 DVDD.n2723 0.00777531
R8079 DVDD.n2780 DVDD.n2725 0.00777531
R8080 DVDD.n2731 DVDD.n2727 0.00777531
R8081 DVDD.n2782 DVDD.n2721 0.00777531
R8082 DVDD.n2730 DVDD.n2728 0.00777531
R8083 DVDD.n2729 DVDD.n2720 0.00777531
R8084 DVDD.n2490 DVDD.n2324 0.00776429
R8085 DVDD.n1305 DVDD.n1301 0.00776429
R8086 DVDD.n1395 DVDD.n1394 0.00776429
R8087 DVDD.n5688 DVDD.n5687 0.00772462
R8088 DVDD.n5971 DVDD.n5970 0.00772462
R8089 DVDD.n5590 DVDD.n5589 0.00772462
R8090 DVDD.n5896 DVDD.n5895 0.00772462
R8091 DVDD.n3652 DVDD.n3651 0.00770384
R8092 DVDD.n3650 DVDD.n1998 0.00770384
R8093 DVDD.n2823 DVDD.n2092 0.0077
R8094 DVDD.n3830 DVDD.n1830 0.0077
R8095 DVDD.n3833 DVDD.n3831 0.0077
R8096 DVDD.n5542 DVDD.n14 0.00762565
R8097 DVDD.n4670 DVDD.n981 0.00762565
R8098 DVDD.n1924 DVDD.n1916 0.00760526
R8099 DVDD.n2727 DVDD.n2726 0.00754348
R8100 DVDD.n1385 DVDD.n1313 0.00751835
R8101 DVDD.n1322 DVDD.n1216 0.00751835
R8102 DVDD.n1323 DVDD.n1316 0.00751005
R8103 DVDD.n1325 DVDD.n1316 0.00751005
R8104 DVDD.n1389 DVDD.n1380 0.00751005
R8105 DVDD.n1389 DVDD.n1388 0.00751005
R8106 DVDD.n3706 DVDD.n1897 0.00748725
R8107 DVDD.n3707 DVDD.n1896 0.00748725
R8108 DVDD.n3762 DVDD.n1666 0.00748725
R8109 DVDD.n3763 DVDD.n1670 0.00748725
R8110 DVDD.n3595 DVDD.n3594 0.00734783
R8111 DVDD.n3429 DVDD.n3208 0.00734783
R8112 DVDD.n2846 DVDD.n2844 0.00734783
R8113 DVDD.n5921 DVDD.n78 0.00731583
R8114 DVDD.n5552 DVDD.n19 0.00731583
R8115 DVDD.n5558 DVDD.n18 0.00731583
R8116 DVDD.n4660 DVDD.n4646 0.00731583
R8117 DVDD.n4645 DVDD.n4644 0.00731583
R8118 DVDD.n331 DVDD.n326 0.00731583
R8119 DVDD.n2834 DVDD.n2095 0.00725
R8120 DVDD.n3900 DVDD.n3866 0.00725
R8121 DVDD.n3869 DVDD.n3865 0.00725
R8122 DVDD.n1373 DVDD.n1372 0.00720213
R8123 DVDD.n1372 DVDD.n1326 0.00720213
R8124 DVDD.n1376 DVDD.n1375 0.00720213
R8125 DVDD.n1377 DVDD.n1376 0.00720213
R8126 DVDD.n3627 DVDD.n2015 0.00717969
R8127 DVDD.n2180 DVDD.n1896 0.00717439
R8128 DVDD.n1765 DVDD.n1724 0.0071375
R8129 DVDD.n2565 DVDD.n2260 0.00712143
R8130 DVDD.n1576 DVDD.n1197 0.00712143
R8131 DVDD.n1573 DVDD.n1572 0.00712143
R8132 DVDD.n1209 DVDD.n1192 0.00712143
R8133 DVDD.n3632 DVDD.n3631 0.0071
R8134 DVDD.n3404 DVDD.n3213 0.0071
R8135 DVDD.n3107 DVDD.n3106 0.0071
R8136 DVDD.n3078 DVDD.n3077 0.0071
R8137 DVDD.n2726 DVDD.n2722 0.00702174
R8138 DVDD.n5535 DVDD.n13 0.00700602
R8139 DVDD.n4677 DVDD.n980 0.00700602
R8140 DVDD.n1371 DVDD.n1195 0.00699624
R8141 DVDD.n2767 DVDD.n2746 0.00699429
R8142 DVDD.n2756 DVDD.n2748 0.00699429
R8143 DVDD.n2763 DVDD.n2745 0.00699429
R8144 DVDD.n2757 DVDD.n2727 0.00699429
R8145 DVDD.n2762 DVDD.n2744 0.00699429
R8146 DVDD.n2758 DVDD.n2749 0.00699429
R8147 DVDD.n2761 DVDD.n2743 0.00699429
R8148 DVDD.n2776 DVDD.n2750 0.00699429
R8149 DVDD.n2768 DVDD.n2767 0.00699429
R8150 DVDD.n2756 DVDD.n2746 0.00699429
R8151 DVDD.n2763 DVDD.n2748 0.00699429
R8152 DVDD.n2757 DVDD.n2745 0.00699429
R8153 DVDD.n2762 DVDD.n2727 0.00699429
R8154 DVDD.n2758 DVDD.n2744 0.00699429
R8155 DVDD.n2761 DVDD.n2749 0.00699429
R8156 DVDD.n2750 DVDD.n2743 0.00699429
R8157 DVDD.n2277 DVDD.n2276 0.00699286
R8158 DVDD.n2557 DVDD.n2264 0.00699286
R8159 DVDD.n3362 DVDD.n3280 0.00698649
R8160 DVDD.n3262 DVDD.n3259 0.00698649
R8161 DVDD.n4082 DVDD.n4081 0.0068
R8162 DVDD.n4044 DVDD.n4041 0.0068
R8163 DVDD.n3678 DVDD.n1973 0.00678
R8164 DVDD.n3461 DVDD.n3460 0.00678
R8165 DVDD.n3147 DVDD.n3146 0.00678
R8166 DVDD.n3048 DVDD.n3032 0.00678
R8167 DVDD.n5519 DVDD.n26 0.00669621
R8168 DVDD.n4693 DVDD.n4653 0.00669621
R8169 DVDD.n4099 DVDD.n4033 0.0066875
R8170 DVDD.n4100 DVDD.n1792 0.0066875
R8171 DVDD.n3494 DVDD.n3189 0.00661413
R8172 DVDD.n3537 DVDD.n3165 0.00661413
R8173 DVDD.n5500 DVDD.n103 0.00660465
R8174 DVDD.n5500 DVDD.n5499 0.00660465
R8175 DVDD.n2594 DVDD.n2593 0.00658571
R8176 DVDD.n2593 DVDD.n2592 0.00658571
R8177 DVDD.n2592 DVDD.n2245 0.00658571
R8178 DVDD.n2586 DVDD.n2245 0.00658571
R8179 DVDD.n2586 DVDD.n2585 0.00658571
R8180 DVDD.n2585 DVDD.n2584 0.00658571
R8181 DVDD.n2584 DVDD.n2249 0.00658571
R8182 DVDD.n2578 DVDD.n2249 0.00658571
R8183 DVDD.n2578 DVDD.n2577 0.00658571
R8184 DVDD.n2577 DVDD.n2576 0.00658571
R8185 DVDD.n2576 DVDD.n2253 0.00658571
R8186 DVDD.n2570 DVDD.n2253 0.00658571
R8187 DVDD.n2570 DVDD.n2569 0.00658571
R8188 DVDD.n2569 DVDD.n2568 0.00658571
R8189 DVDD.n2568 DVDD.n2257 0.00658571
R8190 DVDD.n2271 DVDD.n2257 0.00658571
R8191 DVDD.n2279 DVDD.n2271 0.00658571
R8192 DVDD.n2280 DVDD.n2279 0.00658571
R8193 DVDD.n2281 DVDD.n2280 0.00658571
R8194 DVDD.n2281 DVDD.n2267 0.00658571
R8195 DVDD.n2290 DVDD.n2267 0.00658571
R8196 DVDD.n2291 DVDD.n2290 0.00658571
R8197 DVDD.n2555 DVDD.n2291 0.00658571
R8198 DVDD.n2555 DVDD.n2554 0.00658571
R8199 DVDD.n2554 DVDD.n2553 0.00658571
R8200 DVDD.n2553 DVDD.n2292 0.00658571
R8201 DVDD.n2547 DVDD.n2292 0.00658571
R8202 DVDD.n2547 DVDD.n2546 0.00658571
R8203 DVDD.n2546 DVDD.n2545 0.00658571
R8204 DVDD.n2545 DVDD.n2297 0.00658571
R8205 DVDD.n2304 DVDD.n2297 0.00658571
R8206 DVDD.n2528 DVDD.n2304 0.00658571
R8207 DVDD.n2528 DVDD.n2527 0.00658571
R8208 DVDD.n2527 DVDD.n2526 0.00658571
R8209 DVDD.n2526 DVDD.n2305 0.00658571
R8210 DVDD.n2520 DVDD.n2305 0.00658571
R8211 DVDD.n2520 DVDD.n2519 0.00658571
R8212 DVDD.n2519 DVDD.n2518 0.00658571
R8213 DVDD.n2518 DVDD.n2309 0.00658571
R8214 DVDD.n2512 DVDD.n2309 0.00658571
R8215 DVDD.n2512 DVDD.n2511 0.00658571
R8216 DVDD.n2511 DVDD.n2510 0.00658571
R8217 DVDD.n2510 DVDD.n2313 0.00658571
R8218 DVDD.n2504 DVDD.n2313 0.00658571
R8219 DVDD.n2504 DVDD.n2503 0.00658571
R8220 DVDD.n2503 DVDD.n2502 0.00658571
R8221 DVDD.n2502 DVDD.n2317 0.00658571
R8222 DVDD.n2496 DVDD.n2317 0.00658571
R8223 DVDD.n2496 DVDD.n2495 0.00658571
R8224 DVDD.n2495 DVDD.n2494 0.00658571
R8225 DVDD.n2494 DVDD.n2321 0.00658571
R8226 DVDD.n2336 DVDD.n2321 0.00658571
R8227 DVDD.n2336 DVDD.n2335 0.00658571
R8228 DVDD.n2345 DVDD.n2335 0.00658571
R8229 DVDD.n2346 DVDD.n2345 0.00658571
R8230 DVDD.n2347 DVDD.n2346 0.00658571
R8231 DVDD.n2347 DVDD.n2331 0.00658571
R8232 DVDD.n2356 DVDD.n2331 0.00658571
R8233 DVDD.n2357 DVDD.n2356 0.00658571
R8234 DVDD.n2480 DVDD.n2357 0.00658571
R8235 DVDD.n2480 DVDD.n2479 0.00658571
R8236 DVDD.n2479 DVDD.n2478 0.00658571
R8237 DVDD.n2478 DVDD.n2358 0.00658571
R8238 DVDD.n2472 DVDD.n2358 0.00658571
R8239 DVDD.n2472 DVDD.n2471 0.00658571
R8240 DVDD.n2471 DVDD.n2470 0.00658571
R8241 DVDD.n2470 DVDD.n2363 0.00658571
R8242 DVDD.n2370 DVDD.n2363 0.00658571
R8243 DVDD.n2453 DVDD.n2370 0.00658571
R8244 DVDD.n2453 DVDD.n2452 0.00658571
R8245 DVDD.n2452 DVDD.n2451 0.00658571
R8246 DVDD.n2451 DVDD.n2371 0.00658571
R8247 DVDD.n2445 DVDD.n2371 0.00658571
R8248 DVDD.n2445 DVDD.n2444 0.00658571
R8249 DVDD.n2444 DVDD.n2443 0.00658571
R8250 DVDD.n2443 DVDD.n2375 0.00658571
R8251 DVDD.n2437 DVDD.n2375 0.00658571
R8252 DVDD.n2437 DVDD.n2436 0.00658571
R8253 DVDD.n2436 DVDD.n2435 0.00658571
R8254 DVDD.n2435 DVDD.n2379 0.00658571
R8255 DVDD.n2429 DVDD.n2379 0.00658571
R8256 DVDD.n2429 DVDD.n2428 0.00658571
R8257 DVDD.n2428 DVDD.n2427 0.00658571
R8258 DVDD.n2427 DVDD.n2383 0.00658571
R8259 DVDD.n2421 DVDD.n2383 0.00658571
R8260 DVDD.n2421 DVDD.n2420 0.00658571
R8261 DVDD.n2420 DVDD.n2419 0.00658571
R8262 DVDD.n2419 DVDD.n2387 0.00658571
R8263 DVDD.n2413 DVDD.n2387 0.00658571
R8264 DVDD.n2413 DVDD.n2412 0.00658571
R8265 DVDD.n2412 DVDD.n2411 0.00658571
R8266 DVDD.n2411 DVDD.n2391 0.00658571
R8267 DVDD.n2405 DVDD.n2391 0.00658571
R8268 DVDD.n2405 DVDD.n2404 0.00658571
R8269 DVDD.n2404 DVDD.n2403 0.00658571
R8270 DVDD.n2403 DVDD.n2395 0.00658571
R8271 DVDD.n2610 DVDD.n2166 0.00658571
R8272 DVDD.n2624 DVDD.n2166 0.00658571
R8273 DVDD.n2625 DVDD.n2624 0.00658571
R8274 DVDD.n2626 DVDD.n2625 0.00658571
R8275 DVDD.n2626 DVDD.n2162 0.00658571
R8276 DVDD.n2632 DVDD.n2162 0.00658571
R8277 DVDD.n2633 DVDD.n2632 0.00658571
R8278 DVDD.n2634 DVDD.n2633 0.00658571
R8279 DVDD.n2634 DVDD.n2158 0.00658571
R8280 DVDD.n2640 DVDD.n2158 0.00658571
R8281 DVDD.n2641 DVDD.n2640 0.00658571
R8282 DVDD.n2642 DVDD.n2641 0.00658571
R8283 DVDD.n2642 DVDD.n2154 0.00658571
R8284 DVDD.n2648 DVDD.n2154 0.00658571
R8285 DVDD.n2649 DVDD.n2648 0.00658571
R8286 DVDD.n2650 DVDD.n2649 0.00658571
R8287 DVDD.n2650 DVDD.n2150 0.00658571
R8288 DVDD.n2656 DVDD.n2150 0.00658571
R8289 DVDD.n2657 DVDD.n2656 0.00658571
R8290 DVDD.n2658 DVDD.n2657 0.00658571
R8291 DVDD.n2658 DVDD.n2146 0.00658571
R8292 DVDD.n2664 DVDD.n2146 0.00658571
R8293 DVDD.n2665 DVDD.n2664 0.00658571
R8294 DVDD.n2666 DVDD.n2665 0.00658571
R8295 DVDD.n2666 DVDD.n2142 0.00658571
R8296 DVDD.n2676 DVDD.n2142 0.00658571
R8297 DVDD.n2677 DVDD.n2676 0.00658571
R8298 DVDD.n2678 DVDD.n2677 0.00658571
R8299 DVDD.n2678 DVDD.n2138 0.00658571
R8300 DVDD.n2867 DVDD.n2138 0.00658571
R8301 DVDD.n2868 DVDD.n2867 0.00658571
R8302 DVDD.n2869 DVDD.n2868 0.00658571
R8303 DVDD.n2869 DVDD.n2134 0.00658571
R8304 DVDD.n2875 DVDD.n2134 0.00658571
R8305 DVDD.n2876 DVDD.n2875 0.00658571
R8306 DVDD.n2877 DVDD.n2876 0.00658571
R8307 DVDD.n2877 DVDD.n2130 0.00658571
R8308 DVDD.n2883 DVDD.n2130 0.00658571
R8309 DVDD.n2884 DVDD.n2883 0.00658571
R8310 DVDD.n2885 DVDD.n2884 0.00658571
R8311 DVDD.n2885 DVDD.n2126 0.00658571
R8312 DVDD.n2891 DVDD.n2126 0.00658571
R8313 DVDD.n2892 DVDD.n2891 0.00658571
R8314 DVDD.n2893 DVDD.n2892 0.00658571
R8315 DVDD.n2893 DVDD.n2122 0.00658571
R8316 DVDD.n2899 DVDD.n2122 0.00658571
R8317 DVDD.n2900 DVDD.n2899 0.00658571
R8318 DVDD.n2901 DVDD.n2900 0.00658571
R8319 DVDD.n2901 DVDD.n2118 0.00658571
R8320 DVDD.n2907 DVDD.n2118 0.00658571
R8321 DVDD.n2908 DVDD.n2907 0.00658571
R8322 DVDD.n2909 DVDD.n2908 0.00658571
R8323 DVDD.n2909 DVDD.n2114 0.00658571
R8324 DVDD.n2915 DVDD.n2114 0.00658571
R8325 DVDD.n2916 DVDD.n2915 0.00658571
R8326 DVDD.n2917 DVDD.n2916 0.00658571
R8327 DVDD.n2917 DVDD.n2110 0.00658571
R8328 DVDD.n2923 DVDD.n2110 0.00658571
R8329 DVDD.n2924 DVDD.n2923 0.00658571
R8330 DVDD.n2925 DVDD.n2924 0.00658571
R8331 DVDD.n2925 DVDD.n2106 0.00658571
R8332 DVDD.n2931 DVDD.n2106 0.00658571
R8333 DVDD.n2932 DVDD.n2931 0.00658571
R8334 DVDD.n2933 DVDD.n2932 0.00658571
R8335 DVDD.n2933 DVDD.n2102 0.00658571
R8336 DVDD.n2939 DVDD.n2102 0.00658571
R8337 DVDD.n2940 DVDD.n2939 0.00658571
R8338 DVDD.n2942 DVDD.n2940 0.00658571
R8339 DVDD.n2942 DVDD.n2941 0.00658571
R8340 DVDD.n2941 DVDD.n2086 0.00658571
R8341 DVDD.n2951 DVDD.n2086 0.00658571
R8342 DVDD.n2952 DVDD.n2951 0.00658571
R8343 DVDD.n2953 DVDD.n2952 0.00658571
R8344 DVDD.n2953 DVDD.n2082 0.00658571
R8345 DVDD.n2959 DVDD.n2082 0.00658571
R8346 DVDD.n2960 DVDD.n2959 0.00658571
R8347 DVDD.n3019 DVDD.n2960 0.00658571
R8348 DVDD.n3019 DVDD.n3018 0.00658571
R8349 DVDD.n3018 DVDD.n3017 0.00658571
R8350 DVDD.n3017 DVDD.n2961 0.00658571
R8351 DVDD.n3011 DVDD.n2961 0.00658571
R8352 DVDD.n3011 DVDD.n3010 0.00658571
R8353 DVDD.n3010 DVDD.n3009 0.00658571
R8354 DVDD.n3009 DVDD.n2965 0.00658571
R8355 DVDD.n3003 DVDD.n2965 0.00658571
R8356 DVDD.n3003 DVDD.n3002 0.00658571
R8357 DVDD.n3002 DVDD.n3001 0.00658571
R8358 DVDD.n3001 DVDD.n2969 0.00658571
R8359 DVDD.n2995 DVDD.n2969 0.00658571
R8360 DVDD.n2995 DVDD.n2994 0.00658571
R8361 DVDD.n2994 DVDD.n2993 0.00658571
R8362 DVDD.n2993 DVDD.n2973 0.00658571
R8363 DVDD.n2987 DVDD.n2973 0.00658571
R8364 DVDD.n2987 DVDD.n2986 0.00658571
R8365 DVDD.n2986 DVDD.n2985 0.00658571
R8366 DVDD.n2985 DVDD.n2977 0.00658571
R8367 DVDD.n2979 DVDD.n2977 0.00658571
R8368 DVDD.n1570 DVDD.n1569 0.00658571
R8369 DVDD.n1569 DVDD.n1568 0.00658571
R8370 DVDD.n1568 DVDD.n1207 0.00658571
R8371 DVDD.n1562 DVDD.n1207 0.00658571
R8372 DVDD.n1562 DVDD.n1561 0.00658571
R8373 DVDD.n1561 DVDD.n1560 0.00658571
R8374 DVDD.n1560 DVDD.n1212 0.00658571
R8375 DVDD.n1226 DVDD.n1212 0.00658571
R8376 DVDD.n1551 DVDD.n1226 0.00658571
R8377 DVDD.n1551 DVDD.n1550 0.00658571
R8378 DVDD.n1550 DVDD.n1549 0.00658571
R8379 DVDD.n1549 DVDD.n1227 0.00658571
R8380 DVDD.n1543 DVDD.n1227 0.00658571
R8381 DVDD.n1543 DVDD.n1542 0.00658571
R8382 DVDD.n1542 DVDD.n1541 0.00658571
R8383 DVDD.n1541 DVDD.n1231 0.00658571
R8384 DVDD.n1535 DVDD.n1231 0.00658571
R8385 DVDD.n1535 DVDD.n1534 0.00658571
R8386 DVDD.n1534 DVDD.n1533 0.00658571
R8387 DVDD.n1533 DVDD.n1235 0.00658571
R8388 DVDD.n1527 DVDD.n1235 0.00658571
R8389 DVDD.n1527 DVDD.n1526 0.00658571
R8390 DVDD.n1526 DVDD.n1525 0.00658571
R8391 DVDD.n1525 DVDD.n1239 0.00658571
R8392 DVDD.n1519 DVDD.n1239 0.00658571
R8393 DVDD.n1519 DVDD.n1518 0.00658571
R8394 DVDD.n1518 DVDD.n1517 0.00658571
R8395 DVDD.n1517 DVDD.n1243 0.00658571
R8396 DVDD.n1511 DVDD.n1243 0.00658571
R8397 DVDD.n1511 DVDD.n1510 0.00658571
R8398 DVDD.n1510 DVDD.n1509 0.00658571
R8399 DVDD.n1509 DVDD.n1247 0.00658571
R8400 DVDD.n1503 DVDD.n1247 0.00658571
R8401 DVDD.n1503 DVDD.n1502 0.00658571
R8402 DVDD.n1502 DVDD.n1501 0.00658571
R8403 DVDD.n1501 DVDD.n1251 0.00658571
R8404 DVDD.n1495 DVDD.n1251 0.00658571
R8405 DVDD.n1495 DVDD.n1494 0.00658571
R8406 DVDD.n1494 DVDD.n1493 0.00658571
R8407 DVDD.n1493 DVDD.n1255 0.00658571
R8408 DVDD.n1487 DVDD.n1255 0.00658571
R8409 DVDD.n1487 DVDD.n1486 0.00658571
R8410 DVDD.n1486 DVDD.n1485 0.00658571
R8411 DVDD.n1485 DVDD.n1259 0.00658571
R8412 DVDD.n1479 DVDD.n1259 0.00658571
R8413 DVDD.n1479 DVDD.n1478 0.00658571
R8414 DVDD.n1478 DVDD.n1477 0.00658571
R8415 DVDD.n1477 DVDD.n1263 0.00658571
R8416 DVDD.n1471 DVDD.n1263 0.00658571
R8417 DVDD.n1471 DVDD.n1470 0.00658571
R8418 DVDD.n1470 DVDD.n1469 0.00658571
R8419 DVDD.n1469 DVDD.n1267 0.00658571
R8420 DVDD.n1463 DVDD.n1267 0.00658571
R8421 DVDD.n1463 DVDD.n1462 0.00658571
R8422 DVDD.n1462 DVDD.n1461 0.00658571
R8423 DVDD.n1461 DVDD.n1271 0.00658571
R8424 DVDD.n1455 DVDD.n1271 0.00658571
R8425 DVDD.n1455 DVDD.n1454 0.00658571
R8426 DVDD.n1454 DVDD.n1453 0.00658571
R8427 DVDD.n1453 DVDD.n1275 0.00658571
R8428 DVDD.n1447 DVDD.n1275 0.00658571
R8429 DVDD.n1447 DVDD.n1446 0.00658571
R8430 DVDD.n1446 DVDD.n1445 0.00658571
R8431 DVDD.n1445 DVDD.n1279 0.00658571
R8432 DVDD.n1439 DVDD.n1279 0.00658571
R8433 DVDD.n1439 DVDD.n1438 0.00658571
R8434 DVDD.n1438 DVDD.n1437 0.00658571
R8435 DVDD.n1437 DVDD.n1283 0.00658571
R8436 DVDD.n1431 DVDD.n1283 0.00658571
R8437 DVDD.n1431 DVDD.n1430 0.00658571
R8438 DVDD.n1430 DVDD.n1429 0.00658571
R8439 DVDD.n1429 DVDD.n1287 0.00658571
R8440 DVDD.n1423 DVDD.n1287 0.00658571
R8441 DVDD.n1423 DVDD.n1422 0.00658571
R8442 DVDD.n1422 DVDD.n1421 0.00658571
R8443 DVDD.n1421 DVDD.n1291 0.00658571
R8444 DVDD.n1415 DVDD.n1291 0.00658571
R8445 DVDD.n1415 DVDD.n1414 0.00658571
R8446 DVDD.n1414 DVDD.n1413 0.00658571
R8447 DVDD.n1413 DVDD.n1295 0.00658571
R8448 DVDD.n1407 DVDD.n1295 0.00658571
R8449 DVDD.n1407 DVDD.n1406 0.00658571
R8450 DVDD.n1406 DVDD.n1405 0.00658571
R8451 DVDD.n1405 DVDD.n1299 0.00658571
R8452 DVDD.n1399 DVDD.n1299 0.00658571
R8453 DVDD.n1399 DVDD.n1398 0.00658571
R8454 DVDD.n1398 DVDD.n1397 0.00658571
R8455 DVDD.n1397 DVDD.n1303 0.00658571
R8456 DVDD.n1346 DVDD.n1303 0.00658571
R8457 DVDD.n1351 DVDD.n1346 0.00658571
R8458 DVDD.n1352 DVDD.n1351 0.00658571
R8459 DVDD.n1353 DVDD.n1352 0.00658571
R8460 DVDD.n1353 DVDD.n1342 0.00658571
R8461 DVDD.n1359 DVDD.n1342 0.00658571
R8462 DVDD.n1360 DVDD.n1359 0.00658571
R8463 DVDD.n5510 DVDD.n218 0.00654131
R8464 DVDD.n4705 DVDD.n4704 0.00654131
R8465 DVDD.n4878 DVDD.n703 0.0065
R8466 DVDD.n571 DVDD.n450 0.0065
R8467 DVDD.n909 DVDD.n359 0.0065
R8468 DVDD.n4879 DVDD.n4878 0.0065
R8469 DVDD.n990 DVDD.n358 0.0065
R8470 DVDD.n696 DVDD.n407 0.0065
R8471 DVDD.n4635 DVDD.n990 0.0065
R8472 DVDD.n4871 DVDD.n696 0.0065
R8473 DVDD.n5245 DVDD.n481 0.0065
R8474 DVDD.n4871 DVDD.n4802 0.0065
R8475 DVDD.n4635 DVDD.n908 0.0065
R8476 DVDD.n5710 DVDD.n38 0.0065
R8477 DVDD.n44 DVDD.n38 0.0065
R8478 DVDD.n5246 DVDD.n5245 0.0065
R8479 DVDD.n5246 DVDD.n448 0.0065
R8480 DVDD.n119 DVDD.n44 0.0065
R8481 DVDD.n5399 DVDD.n359 0.0065
R8482 DVDD.n4879 DVDD.n405 0.0065
R8483 DVDD.n5937 DVDD.n41 0.0065
R8484 DVDD.n5319 DVDD.n450 0.0065
R8485 DVDD.n5320 DVDD.n5319 0.0065
R8486 DVDD.n5938 DVDD.n40 0.0065
R8487 DVDD.n5938 DVDD.n5937 0.0065
R8488 DVDD.n4718 DVDD.n909 0.0065
R8489 DVDD.n4197 DVDD.n4190 0.00642084
R8490 DVDD.n71 DVDD.n69 0.0063864
R8491 DVDD.n5434 DVDD.n285 0.0063864
R8492 DVDD.n2857 DVDD.n2689 0.00636957
R8493 DVDD.n2343 DVDD.n2342 0.00635
R8494 DVDD.n2483 DVDD.n2482 0.00635
R8495 DVDD.n2482 DVDD.n2328 0.00635
R8496 DVDD.n1741 DVDD.n1738 0.00635
R8497 DVDD.n1744 DVDD.n1743 0.00635
R8498 DVDD.n1391 DVDD.n1389 0.00635
R8499 DVDD.n1316 DVDD.n1315 0.00635
R8500 DVDD.n3921 DVDD.n1818 0.0062375
R8501 DVDD.n3975 DVDD.n3922 0.0062375
R8502 DVDD.n84 DVDD.n78 0.0062315
R8503 DVDD.n331 DVDD.n329 0.0062315
R8504 DVDD.n5625 DVDD.n5571 0.00607659
R8505 DVDD.n5450 DVDD.n280 0.00607659
R8506 DVDD.n5829 DVDD.n146 0.00603279
R8507 DVDD.n5185 DVDD.n455 0.00603279
R8508 DVDD.n4953 DVDD.n678 0.00603279
R8509 DVDD.n812 DVDD.n811 0.00603279
R8510 DVDD.n4509 DVDD.n1079 0.00603279
R8511 DVDD.n4067 DVDD.n4052 0.0060125
R8512 DVDD.n4066 DVDD.n4053 0.0060125
R8513 DVDD.n4063 DVDD.n4062 0.0060125
R8514 DVDD.n4057 DVDD.n4055 0.0060125
R8515 DVDD.n4056 DVDD.n1721 0.0060125
R8516 DVDD.n4225 DVDD.n4224 0.0060125
R8517 DVDD.n1764 DVDD.n1728 0.0060125
R8518 DVDD.n1763 DVDD.n1729 0.0060125
R8519 DVDD.n1760 DVDD.n1759 0.0060125
R8520 DVDD.n1734 DVDD.n1730 0.0060125
R8521 DVDD.n3124 DVDD.n3123 0.00588043
R8522 DVDD.n3557 DVDD.n3555 0.00588043
R8523 DVDD.n3554 DVDD.n3160 0.00588043
R8524 DVDD.n3471 DVDD.n3184 0.00588043
R8525 DVDD.n3431 DVDD.n3209 0.00588043
R8526 DVDD.n3474 DVDD.n3472 0.00588043
R8527 DVDD.n3651 DVDD 0.00587887
R8528 DVDD.n3650 DVDD 0.00587887
R8529 DVDD.n1679 DVDD.n1675 0.00584375
R8530 DVDD.n4266 DVDD.n1680 0.00584375
R8531 DVDD.n4265 DVDD.n1681 0.00584375
R8532 DVDD.n4262 DVDD.n4261 0.00584375
R8533 DVDD.n3810 DVDD.n1843 0.00584375
R8534 DVDD.n3812 DVDD.n3811 0.00584375
R8535 DVDD.n3817 DVDD.n1840 0.00584375
R8536 DVDD.n3816 DVDD.n1841 0.00584375
R8537 DVDD.n3823 DVDD.n1836 0.00584375
R8538 DVDD.n2542 DVDD.n2541 0.00583571
R8539 DVDD.n4078 DVDD.n4045 0.005825
R8540 DVDD.n4049 DVDD.n4045 0.005825
R8541 DVDD.n4071 DVDD.n4049 0.005825
R8542 DVDD.n4071 DVDD.n4070 0.005825
R8543 DVDD.n4070 DVDD.n4069 0.005825
R8544 DVDD.n4069 DVDD.n4050 0.005825
R8545 DVDD.n4060 DVDD.n4050 0.005825
R8546 DVDD.n4060 DVDD.n4059 0.005825
R8547 DVDD.n4059 DVDD.n1725 0.005825
R8548 DVDD.n4222 DVDD.n1725 0.005825
R8549 DVDD.n1766 DVDD.n1726 0.005825
R8550 DVDD.n1757 DVDD.n1726 0.005825
R8551 DVDD.n1757 DVDD.n1756 0.005825
R8552 DVDD.n1756 DVDD.n1755 0.005825
R8553 DVDD.n1755 DVDD.n1732 0.005825
R8554 DVDD.n1749 DVDD.n1732 0.005825
R8555 DVDD.n1749 DVDD.n1748 0.005825
R8556 DVDD.n1748 DVDD.n1747 0.005825
R8557 DVDD.n1747 DVDD.n1737 0.005825
R8558 DVDD.n4284 DVDD.n1668 0.005825
R8559 DVDD.n4278 DVDD.n1668 0.005825
R8560 DVDD.n4278 DVDD.n4277 0.005825
R8561 DVDD.n4277 DVDD.n4276 0.005825
R8562 DVDD.n4276 DVDD.n1673 0.005825
R8563 DVDD.n4270 DVDD.n1673 0.005825
R8564 DVDD.n4270 DVDD.n4269 0.005825
R8565 DVDD.n4269 DVDD.n4268 0.005825
R8566 DVDD.n4268 DVDD.n1677 0.005825
R8567 DVDD.n4259 DVDD.n1677 0.005825
R8568 DVDD.n3808 DVDD.n1686 0.005825
R8569 DVDD.n3808 DVDD.n1838 0.005825
R8570 DVDD.n3819 DVDD.n1838 0.005825
R8571 DVDD.n3820 DVDD.n3819 0.005825
R8572 DVDD.n3821 DVDD.n3820 0.005825
R8573 DVDD.n3821 DVDD.n1834 0.005825
R8574 DVDD.n3827 DVDD.n1834 0.005825
R8575 DVDD.n3828 DVDD.n3827 0.005825
R8576 DVDD.n3829 DVDD.n3828 0.005825
R8577 DVDD.n3873 DVDD.n3867 0.005825
R8578 DVDD.n3894 DVDD.n3873 0.005825
R8579 DVDD.n3894 DVDD.n3893 0.005825
R8580 DVDD.n3893 DVDD.n3892 0.005825
R8581 DVDD.n3892 DVDD.n3874 0.005825
R8582 DVDD.n3886 DVDD.n3874 0.005825
R8583 DVDD.n3886 DVDD.n3885 0.005825
R8584 DVDD.n3885 DVDD.n3884 0.005825
R8585 DVDD.n3884 DVDD.n3878 0.005825
R8586 DVDD.n3878 DVDD.n1790 0.005825
R8587 DVDD.n4101 DVDD.n1791 0.005825
R8588 DVDD.n4095 DVDD.n1791 0.005825
R8589 DVDD.n4095 DVDD.n4094 0.005825
R8590 DVDD.n4094 DVDD.n4093 0.005825
R8591 DVDD.n4093 DVDD.n4036 0.005825
R8592 DVDD.n4087 DVDD.n4036 0.005825
R8593 DVDD.n4087 DVDD.n4086 0.005825
R8594 DVDD.n4086 DVDD.n4085 0.005825
R8595 DVDD.n4085 DVDD.n4040 0.005825
R8596 DVDD.n3837 DVDD.n3836 0.005825
R8597 DVDD.n3838 DVDD.n3837 0.005825
R8598 DVDD.n3838 DVDD.n1825 0.005825
R8599 DVDD.n3844 DVDD.n1825 0.005825
R8600 DVDD.n3845 DVDD.n3844 0.005825
R8601 DVDD.n3846 DVDD.n3845 0.005825
R8602 DVDD.n3846 DVDD.n1821 0.005825
R8603 DVDD.n3852 DVDD.n1821 0.005825
R8604 DVDD.n3853 DVDD.n3852 0.005825
R8605 DVDD.n3854 DVDD.n3853 0.005825
R8606 DVDD.n3920 DVDD.n3919 0.005825
R8607 DVDD.n3919 DVDD.n3918 0.005825
R8608 DVDD.n3918 DVDD.n3859 0.005825
R8609 DVDD.n3912 DVDD.n3859 0.005825
R8610 DVDD.n3912 DVDD.n3911 0.005825
R8611 DVDD.n3911 DVDD.n3910 0.005825
R8612 DVDD.n3910 DVDD.n3863 0.005825
R8613 DVDD.n3904 DVDD.n3863 0.005825
R8614 DVDD.n3904 DVDD.n3903 0.005825
R8615 DVDD.n3807 DVDD.n1685 0.0057875
R8616 DVDD.n3806 DVDD.n3805 0.0057875
R8617 DVDD.n5642 DVDD.n5608 0.00576678
R8618 DVDD.n5467 DVDD.n292 0.00576678
R8619 DVDD.n3704 DVDD.n1968 0.00571437
R8620 DVDD.n4286 DVDD.n4285 0.00571437
R8621 DVDD.n2558 DVDD.n2557 0.00570714
R8622 DVDD.n5743 DVDD.n187 0.00566393
R8623 DVDD.n5241 DVDD.n5240 0.00566393
R8624 DVDD.n5013 DVDD.n604 0.00566393
R8625 DVDD.n4876 DVDD.n727 0.00566393
R8626 DVDD.n4614 DVDD.n4613 0.00566393
R8627 DVDD.n3479 DVDD.n3180 0.00563587
R8628 DVDD.n3168 DVDD.n3150 0.00563587
R8629 DVDD.n5565 DVDD.n49 0.00561188
R8630 DVDD.n274 DVDD.n272 0.00561188
R8631 DVDD.n966 DVDD.n965 0.00559827
R8632 DVDD.n5504 DVDD.n5503 0.00558651
R8633 DVDD.n2596 DVDD.n2240 0.00548841
R8634 DVDD.n2612 DVDD.n2604 0.00548841
R8635 DVDD DVDD.n2395 0.00538571
R8636 DVDD.n3649 DVDD.n3647 0.00530256
R8637 DVDD.n5634 DVDD.n64 0.00530207
R8638 DVDD.n225 DVDD.n221 0.00530207
R8639 DVDD.n962 DVDD.n947 0.00530207
R8640 DVDD.n5459 DVDD.n301 0.00530207
R8641 DVDD.n3829 DVDD.n1829 0.0053
R8642 DVDD.n5813 DVDD.n160 0.00529508
R8643 DVDD.n5169 DVDD.n471 0.00529508
R8644 DVDD.n4969 DVDD.n4947 0.00529508
R8645 DVDD.n793 DVDD.n747 0.00529508
R8646 DVDD.n4525 DVDD.n4505 0.00529508
R8647 DVDD.n2467 DVDD.n2466 0.00519286
R8648 DVDD.n3705 DVDD.n3704 0.00515817
R8649 DVDD.n4285 DVDD.n1667 0.00515817
R8650 DVDD.n5527 DVDD.n11 0.00514716
R8651 DVDD.n4685 DVDD.n978 0.00514716
R8652 DVDD.n3486 DVDD.n3179 0.00514674
R8653 DVDD.n3545 DVDD.n3151 0.00514674
R8654 DVDD.n3903 DVDD.n3902 0.005
R8655 DVDD.n5617 DVDD.n56 0.00499225
R8656 DVDD.n5442 DVDD.n310 0.00499225
R8657 DVDD.n2466 DVDD.n2366 0.00493571
R8658 DVDD.n5759 DVDD.n172 0.00492623
R8659 DVDD.n5224 DVDD.n489 0.00492623
R8660 DVDD.n643 DVDD.n608 0.00492623
R8661 DVDD.n850 DVDD.n708 0.00492623
R8662 DVDD.n4597 DVDD.n1013 0.00492623
R8663 DVDD.n4221 DVDD.n1766 0.004925
R8664 DVDD.n5911 DVDD.n99 0.00490722
R8665 DVDD.n109 DVDD.n95 0.00490722
R8666 DVDD.n5414 DVDD.n338 0.00490722
R8667 DVDD.n352 DVDD.n342 0.00490722
R8668 DVDD.n941 DVDD.n940 0.00490722
R8669 DVDD.n958 DVDD.n920 0.00490722
R8670 DVDD.n240 DVDD.n233 0.00490722
R8671 DVDD.n246 DVDD.n239 0.00490722
R8672 DVDD.n1932 DVDD.n1931 0.00489803
R8673 DVDD.n1962 DVDD.n1961 0.00489803
R8674 DVDD.n1938 DVDD.n1937 0.00488868
R8675 DVDD.n3698 DVDD.n3697 0.00488868
R8676 DVDD.n4678 DVDD.n4676 0.00486994
R8677 DVDD.n5537 DVDD.n5536 0.00485986
R8678 DVDD.n5544 DVDD.n21 0.00483735
R8679 DVDD.n4668 DVDD.n4648 0.00483735
R8680 DVDD.n4329 DVDD.n4328 0.00476
R8681 DVDD.n4328 DVDD.n4327 0.00476
R8682 DVDD.n4327 DVDD.n4326 0.00476
R8683 DVDD.n4326 DVDD.n4304 0.00476
R8684 DVDD.n4322 DVDD.n4304 0.00476
R8685 DVDD.n4322 DVDD.n4321 0.00476
R8686 DVDD.n4321 DVDD.n4320 0.00476
R8687 DVDD.n4320 DVDD.n4310 0.00476
R8688 DVDD.n4316 DVDD.n4310 0.00476
R8689 DVDD.n4316 DVDD.n4315 0.00476
R8690 DVDD.n4315 DVDD.n913 0.00476
R8691 DVDD.n4712 DVDD.n913 0.00476
R8692 DVDD.n4712 DVDD.n911 0.00476
R8693 DVDD.n4716 DVDD.n911 0.00476
R8694 DVDD.n4720 DVDD.n906 0.00476
R8695 DVDD.n4724 DVDD.n906 0.00476
R8696 DVDD.n4724 DVDD.n904 0.00476
R8697 DVDD.n4728 DVDD.n904 0.00476
R8698 DVDD.n4728 DVDD.n902 0.00476
R8699 DVDD.n4732 DVDD.n902 0.00476
R8700 DVDD.n4732 DVDD.n900 0.00476
R8701 DVDD.n4736 DVDD.n900 0.00476
R8702 DVDD.n4736 DVDD.n898 0.00476
R8703 DVDD.n4740 DVDD.n898 0.00476
R8704 DVDD.n4740 DVDD.n890 0.00476
R8705 DVDD.n4746 DVDD.n890 0.00476
R8706 DVDD.n4746 DVDD.n888 0.00476
R8707 DVDD.n4750 DVDD.n888 0.00476
R8708 DVDD.n4750 DVDD.n886 0.00476
R8709 DVDD.n4754 DVDD.n886 0.00476
R8710 DVDD.n4754 DVDD.n884 0.00476
R8711 DVDD.n4758 DVDD.n884 0.00476
R8712 DVDD.n4758 DVDD.n882 0.00476
R8713 DVDD.n4762 DVDD.n882 0.00476
R8714 DVDD.n4762 DVDD.n880 0.00476
R8715 DVDD.n4768 DVDD.n880 0.00476
R8716 DVDD.n4768 DVDD.n732 0.00476
R8717 DVDD.n4801 DVDD.n734 0.00476
R8718 DVDD.n4797 DVDD.n734 0.00476
R8719 DVDD.n4797 DVDD.n4796 0.00476
R8720 DVDD.n4796 DVDD.n4795 0.00476
R8721 DVDD.n4795 DVDD.n4779 0.00476
R8722 DVDD.n4791 DVDD.n4779 0.00476
R8723 DVDD.n4791 DVDD.n4790 0.00476
R8724 DVDD.n4790 DVDD.n4789 0.00476
R8725 DVDD.n4789 DVDD.n4786 0.00476
R8726 DVDD.n4786 DVDD.n587 0.00476
R8727 DVDD.n5022 DVDD.n587 0.00476
R8728 DVDD.n5022 DVDD.n585 0.00476
R8729 DVDD.n5026 DVDD.n585 0.00476
R8730 DVDD.n5026 DVDD.n583 0.00476
R8731 DVDD.n5030 DVDD.n583 0.00476
R8732 DVDD.n5030 DVDD.n581 0.00476
R8733 DVDD.n5034 DVDD.n581 0.00476
R8734 DVDD.n5034 DVDD.n579 0.00476
R8735 DVDD.n5038 DVDD.n579 0.00476
R8736 DVDD.n5038 DVDD.n577 0.00476
R8737 DVDD.n5042 DVDD.n577 0.00476
R8738 DVDD.n5042 DVDD.n575 0.00476
R8739 DVDD.n5046 DVDD.n575 0.00476
R8740 DVDD.n5084 DVDD.n5083 0.00476
R8741 DVDD.n5083 DVDD.n5051 0.00476
R8742 DVDD.n5079 DVDD.n5051 0.00476
R8743 DVDD.n5079 DVDD.n5078 0.00476
R8744 DVDD.n5078 DVDD.n5077 0.00476
R8745 DVDD.n5077 DVDD.n5057 0.00476
R8746 DVDD.n5073 DVDD.n5057 0.00476
R8747 DVDD.n5073 DVDD.n5072 0.00476
R8748 DVDD.n5072 DVDD.n5071 0.00476
R8749 DVDD.n5071 DVDD.n5063 0.00476
R8750 DVDD.n5067 DVDD.n5063 0.00476
R8751 DVDD.n5067 DVDD.n200 0.00476
R8752 DVDD.n5726 DVDD.n200 0.00476
R8753 DVDD.n5726 DVDD.n5725 0.00476
R8754 DVDD.n5725 DVDD.n5724 0.00476
R8755 DVDD.n5724 DVDD.n204 0.00476
R8756 DVDD.n5720 DVDD.n204 0.00476
R8757 DVDD.n5720 DVDD.n5719 0.00476
R8758 DVDD.n5719 DVDD.n5718 0.00476
R8759 DVDD.n5718 DVDD.n210 0.00476
R8760 DVDD.n5714 DVDD.n210 0.00476
R8761 DVDD.n5714 DVDD.n5713 0.00476
R8762 DVDD.n5713 DVDD.n5712 0.00476
R8763 DVDD.n5709 DVDD.n217 0.00476
R8764 DVDD.n5700 DVDD.n217 0.00476
R8765 DVDD.n5700 DVDD.n5699 0.00476
R8766 DVDD.n5699 DVDD.n5698 0.00476
R8767 DVDD.n5698 DVDD.n5697 0.00476
R8768 DVDD.n5697 DVDD.n5678 0.00476
R8769 DVDD.n5693 DVDD.n5678 0.00476
R8770 DVDD.n5693 DVDD.n5692 0.00476
R8771 DVDD.n5692 DVDD.n5691 0.00476
R8772 DVDD.n5691 DVDD.n5684 0.00476
R8773 DVDD.n4372 DVDD.n4371 0.00476
R8774 DVDD.n4371 DVDD.n4370 0.00476
R8775 DVDD.n4370 DVDD.n4369 0.00476
R8776 DVDD.n4369 DVDD.n4349 0.00476
R8777 DVDD.n4365 DVDD.n4349 0.00476
R8778 DVDD.n4365 DVDD.n4364 0.00476
R8779 DVDD.n4364 DVDD.n4363 0.00476
R8780 DVDD.n4363 DVDD.n4355 0.00476
R8781 DVDD.n4359 DVDD.n4355 0.00476
R8782 DVDD.n4359 DVDD.n985 0.00476
R8783 DVDD.n4642 DVDD.n985 0.00476
R8784 DVDD.n4642 DVDD.n4641 0.00476
R8785 DVDD.n4641 DVDD.n4639 0.00476
R8786 DVDD.n4639 DVDD.n4637 0.00476
R8787 DVDD.n4634 DVDD.n992 0.00476
R8788 DVDD.n4630 DVDD.n992 0.00476
R8789 DVDD.n4630 DVDD.n4629 0.00476
R8790 DVDD.n4629 DVDD.n4628 0.00476
R8791 DVDD.n4628 DVDD.n998 0.00476
R8792 DVDD.n4624 DVDD.n998 0.00476
R8793 DVDD.n4624 DVDD.n4623 0.00476
R8794 DVDD.n4623 DVDD.n4622 0.00476
R8795 DVDD.n4622 DVDD.n1004 0.00476
R8796 DVDD.n4618 DVDD.n1004 0.00476
R8797 DVDD.n4618 DVDD.n4617 0.00476
R8798 DVDD.n4617 DVDD.n1009 0.00476
R8799 DVDD.n1044 DVDD.n1009 0.00476
R8800 DVDD.n1044 DVDD.n1043 0.00476
R8801 DVDD.n1043 DVDD.n1042 0.00476
R8802 DVDD.n1042 DVDD.n1025 0.00476
R8803 DVDD.n1038 DVDD.n1025 0.00476
R8804 DVDD.n1038 DVDD.n1037 0.00476
R8805 DVDD.n1037 DVDD.n1036 0.00476
R8806 DVDD.n1036 DVDD.n1033 0.00476
R8807 DVDD.n1033 DVDD.n729 0.00476
R8808 DVDD.n4873 DVDD.n729 0.00476
R8809 DVDD.n4873 DVDD.n4872 0.00476
R8810 DVDD.n4870 DVDD.n4869 0.00476
R8811 DVDD.n4869 DVDD.n4805 0.00476
R8812 DVDD.n4865 DVDD.n4805 0.00476
R8813 DVDD.n4865 DVDD.n4864 0.00476
R8814 DVDD.n4864 DVDD.n4863 0.00476
R8815 DVDD.n4863 DVDD.n4811 0.00476
R8816 DVDD.n4859 DVDD.n4811 0.00476
R8817 DVDD.n4859 DVDD.n4858 0.00476
R8818 DVDD.n4858 DVDD.n4857 0.00476
R8819 DVDD.n4857 DVDD.n4854 0.00476
R8820 DVDD.n4854 DVDD.n4853 0.00476
R8821 DVDD.n4853 DVDD.n4852 0.00476
R8822 DVDD.n4852 DVDD.n4851 0.00476
R8823 DVDD.n4851 DVDD.n4821 0.00476
R8824 DVDD.n4847 DVDD.n4821 0.00476
R8825 DVDD.n4847 DVDD.n4846 0.00476
R8826 DVDD.n4846 DVDD.n4845 0.00476
R8827 DVDD.n4845 DVDD.n4827 0.00476
R8828 DVDD.n4841 DVDD.n4827 0.00476
R8829 DVDD.n4841 DVDD.n4840 0.00476
R8830 DVDD.n4840 DVDD.n4839 0.00476
R8831 DVDD.n4839 DVDD.n4835 0.00476
R8832 DVDD.n4835 DVDD.n482 0.00476
R8833 DVDD.n5244 DVDD.n484 0.00476
R8834 DVDD.n553 DVDD.n484 0.00476
R8835 DVDD.n553 DVDD.n552 0.00476
R8836 DVDD.n552 DVDD.n551 0.00476
R8837 DVDD.n551 DVDD.n501 0.00476
R8838 DVDD.n547 DVDD.n501 0.00476
R8839 DVDD.n547 DVDD.n546 0.00476
R8840 DVDD.n546 DVDD.n545 0.00476
R8841 DVDD.n545 DVDD.n507 0.00476
R8842 DVDD.n541 DVDD.n507 0.00476
R8843 DVDD.n541 DVDD.n540 0.00476
R8844 DVDD.n540 DVDD.n539 0.00476
R8845 DVDD.n539 DVDD.n538 0.00476
R8846 DVDD.n538 DVDD.n513 0.00476
R8847 DVDD.n534 DVDD.n513 0.00476
R8848 DVDD.n534 DVDD.n533 0.00476
R8849 DVDD.n533 DVDD.n532 0.00476
R8850 DVDD.n532 DVDD.n519 0.00476
R8851 DVDD.n528 DVDD.n519 0.00476
R8852 DVDD.n528 DVDD.n527 0.00476
R8853 DVDD.n527 DVDD.n526 0.00476
R8854 DVDD.n526 DVDD.n37 0.00476
R8855 DVDD.n5940 DVDD.n37 0.00476
R8856 DVDD.n5950 DVDD.n33 0.00476
R8857 DVDD.n5950 DVDD.n5949 0.00476
R8858 DVDD.n5949 DVDD.n5947 0.00476
R8859 DVDD.n5947 DVDD.n6 0.00476
R8860 DVDD.n5957 DVDD.n6 0.00476
R8861 DVDD.n5957 DVDD.n4 0.00476
R8862 DVDD.n5962 DVDD.n4 0.00476
R8863 DVDD.n5962 DVDD.n2 0.00476
R8864 DVDD.n5966 DVDD.n2 0.00476
R8865 DVDD.n5967 DVDD.n5966 0.00476
R8866 DVDD.n4409 DVDD.n1107 0.00476
R8867 DVDD.n4416 DVDD.n1107 0.00476
R8868 DVDD.n4416 DVDD.n1105 0.00476
R8869 DVDD.n4420 DVDD.n1105 0.00476
R8870 DVDD.n4420 DVDD.n1103 0.00476
R8871 DVDD.n4424 DVDD.n1103 0.00476
R8872 DVDD.n4424 DVDD.n1101 0.00476
R8873 DVDD.n4428 DVDD.n1101 0.00476
R8874 DVDD.n4428 DVDD.n1099 0.00476
R8875 DVDD.n4432 DVDD.n1099 0.00476
R8876 DVDD.n4432 DVDD.n1097 0.00476
R8877 DVDD.n4436 DVDD.n1097 0.00476
R8878 DVDD.n4437 DVDD.n4436 0.00476
R8879 DVDD.n4438 DVDD.n4437 0.00476
R8880 DVDD.n4445 DVDD.n4442 0.00476
R8881 DVDD.n4445 DVDD.n1093 0.00476
R8882 DVDD.n4449 DVDD.n1093 0.00476
R8883 DVDD.n4449 DVDD.n1091 0.00476
R8884 DVDD.n4453 DVDD.n1091 0.00476
R8885 DVDD.n4453 DVDD.n1089 0.00476
R8886 DVDD.n4457 DVDD.n1089 0.00476
R8887 DVDD.n4457 DVDD.n1087 0.00476
R8888 DVDD.n4461 DVDD.n1087 0.00476
R8889 DVDD.n4461 DVDD.n1085 0.00476
R8890 DVDD.n4496 DVDD.n1085 0.00476
R8891 DVDD.n4496 DVDD.n4495 0.00476
R8892 DVDD.n4495 DVDD.n4466 0.00476
R8893 DVDD.n4491 DVDD.n4466 0.00476
R8894 DVDD.n4491 DVDD.n4490 0.00476
R8895 DVDD.n4490 DVDD.n4489 0.00476
R8896 DVDD.n4489 DVDD.n4472 0.00476
R8897 DVDD.n4485 DVDD.n4472 0.00476
R8898 DVDD.n4485 DVDD.n4484 0.00476
R8899 DVDD.n4484 DVDD.n4483 0.00476
R8900 DVDD.n4483 DVDD.n4479 0.00476
R8901 DVDD.n4479 DVDD.n701 0.00476
R8902 DVDD.n4881 DVDD.n701 0.00476
R8903 DVDD.n4885 DVDD.n694 0.00476
R8904 DVDD.n4889 DVDD.n694 0.00476
R8905 DVDD.n4889 DVDD.n692 0.00476
R8906 DVDD.n4893 DVDD.n692 0.00476
R8907 DVDD.n4893 DVDD.n690 0.00476
R8908 DVDD.n4897 DVDD.n690 0.00476
R8909 DVDD.n4897 DVDD.n688 0.00476
R8910 DVDD.n4901 DVDD.n688 0.00476
R8911 DVDD.n4901 DVDD.n686 0.00476
R8912 DVDD.n4905 DVDD.n686 0.00476
R8913 DVDD.n4905 DVDD.n684 0.00476
R8914 DVDD.n4937 DVDD.n684 0.00476
R8915 DVDD.n4937 DVDD.n4936 0.00476
R8916 DVDD.n4936 DVDD.n4910 0.00476
R8917 DVDD.n4932 DVDD.n4910 0.00476
R8918 DVDD.n4932 DVDD.n4931 0.00476
R8919 DVDD.n4931 DVDD.n4930 0.00476
R8920 DVDD.n4930 DVDD.n4916 0.00476
R8921 DVDD.n4926 DVDD.n4916 0.00476
R8922 DVDD.n4926 DVDD.n4925 0.00476
R8923 DVDD.n4925 DVDD.n4924 0.00476
R8924 DVDD.n4924 DVDD.n480 0.00476
R8925 DVDD.n5247 DVDD.n480 0.00476
R8926 DVDD.n5314 DVDD.n476 0.00476
R8927 DVDD.n5314 DVDD.n5313 0.00476
R8928 DVDD.n5313 DVDD.n5312 0.00476
R8929 DVDD.n5312 DVDD.n5254 0.00476
R8930 DVDD.n5308 DVDD.n5254 0.00476
R8931 DVDD.n5308 DVDD.n5307 0.00476
R8932 DVDD.n5307 DVDD.n5306 0.00476
R8933 DVDD.n5306 DVDD.n5260 0.00476
R8934 DVDD.n5302 DVDD.n5260 0.00476
R8935 DVDD.n5302 DVDD.n5301 0.00476
R8936 DVDD.n5301 DVDD.n5300 0.00476
R8937 DVDD.n5300 DVDD.n5298 0.00476
R8938 DVDD.n5298 DVDD.n5297 0.00476
R8939 DVDD.n5297 DVDD.n5296 0.00476
R8940 DVDD.n5296 DVDD.n5269 0.00476
R8941 DVDD.n5292 DVDD.n5269 0.00476
R8942 DVDD.n5292 DVDD.n5291 0.00476
R8943 DVDD.n5291 DVDD.n5290 0.00476
R8944 DVDD.n5290 DVDD.n5275 0.00476
R8945 DVDD.n5286 DVDD.n5275 0.00476
R8946 DVDD.n5286 DVDD.n5285 0.00476
R8947 DVDD.n5285 DVDD.n5284 0.00476
R8948 DVDD.n5284 DVDD.n5282 0.00476
R8949 DVDD.n5935 DVDD.n5934 0.00476
R8950 DVDD.n5934 DVDD.n47 0.00476
R8951 DVDD.n5576 DVDD.n47 0.00476
R8952 DVDD.n5600 DVDD.n5576 0.00476
R8953 DVDD.n5600 DVDD.n5599 0.00476
R8954 DVDD.n5599 DVDD.n5598 0.00476
R8955 DVDD.n5598 DVDD.n5582 0.00476
R8956 DVDD.n5594 DVDD.n5582 0.00476
R8957 DVDD.n5594 DVDD.n5593 0.00476
R8958 DVDD.n5593 DVDD.n5592 0.00476
R8959 DVDD.n1180 DVDD.n1179 0.00476
R8960 DVDD.n1179 DVDD.n1178 0.00476
R8961 DVDD.n1178 DVDD.n1177 0.00476
R8962 DVDD.n1177 DVDD.n1154 0.00476
R8963 DVDD.n1173 DVDD.n1154 0.00476
R8964 DVDD.n1173 DVDD.n1172 0.00476
R8965 DVDD.n1172 DVDD.n1171 0.00476
R8966 DVDD.n1171 DVDD.n1160 0.00476
R8967 DVDD.n1167 DVDD.n1160 0.00476
R8968 DVDD.n1167 DVDD.n1166 0.00476
R8969 DVDD.n1166 DVDD.n354 0.00476
R8970 DVDD.n5404 DVDD.n354 0.00476
R8971 DVDD.n5404 DVDD.n5403 0.00476
R8972 DVDD.n5403 DVDD.n5401 0.00476
R8973 DVDD.n5397 DVDD.n5396 0.00476
R8974 DVDD.n5396 DVDD.n5395 0.00476
R8975 DVDD.n5395 DVDD.n364 0.00476
R8976 DVDD.n5391 DVDD.n364 0.00476
R8977 DVDD.n5391 DVDD.n5390 0.00476
R8978 DVDD.n5390 DVDD.n5389 0.00476
R8979 DVDD.n5389 DVDD.n370 0.00476
R8980 DVDD.n5385 DVDD.n370 0.00476
R8981 DVDD.n5385 DVDD.n5384 0.00476
R8982 DVDD.n5384 DVDD.n5383 0.00476
R8983 DVDD.n5383 DVDD.n376 0.00476
R8984 DVDD.n5377 DVDD.n376 0.00476
R8985 DVDD.n5377 DVDD.n5376 0.00476
R8986 DVDD.n5376 DVDD.n5375 0.00476
R8987 DVDD.n5375 DVDD.n387 0.00476
R8988 DVDD.n5371 DVDD.n387 0.00476
R8989 DVDD.n5371 DVDD.n5370 0.00476
R8990 DVDD.n5370 DVDD.n5369 0.00476
R8991 DVDD.n5369 DVDD.n393 0.00476
R8992 DVDD.n5365 DVDD.n393 0.00476
R8993 DVDD.n5365 DVDD.n5364 0.00476
R8994 DVDD.n5364 DVDD.n5363 0.00476
R8995 DVDD.n5363 DVDD.n399 0.00476
R8996 DVDD.n5357 DVDD.n5356 0.00476
R8997 DVDD.n5356 DVDD.n5355 0.00476
R8998 DVDD.n5355 DVDD.n411 0.00476
R8999 DVDD.n5351 DVDD.n411 0.00476
R9000 DVDD.n5351 DVDD.n5350 0.00476
R9001 DVDD.n5350 DVDD.n5349 0.00476
R9002 DVDD.n5349 DVDD.n417 0.00476
R9003 DVDD.n5345 DVDD.n417 0.00476
R9004 DVDD.n5345 DVDD.n5344 0.00476
R9005 DVDD.n5344 DVDD.n5343 0.00476
R9006 DVDD.n5343 DVDD.n423 0.00476
R9007 DVDD.n430 DVDD.n423 0.00476
R9008 DVDD.n5336 DVDD.n430 0.00476
R9009 DVDD.n5336 DVDD.n5335 0.00476
R9010 DVDD.n5335 DVDD.n5334 0.00476
R9011 DVDD.n5334 DVDD.n436 0.00476
R9012 DVDD.n5330 DVDD.n436 0.00476
R9013 DVDD.n5330 DVDD.n5329 0.00476
R9014 DVDD.n5329 DVDD.n5328 0.00476
R9015 DVDD.n5328 DVDD.n442 0.00476
R9016 DVDD.n5324 DVDD.n442 0.00476
R9017 DVDD.n5324 DVDD.n5323 0.00476
R9018 DVDD.n5323 DVDD.n5322 0.00476
R9019 DVDD.n5132 DVDD.n5106 0.00476
R9020 DVDD.n5132 DVDD.n5131 0.00476
R9021 DVDD.n5131 DVDD.n5130 0.00476
R9022 DVDD.n5130 DVDD.n5111 0.00476
R9023 DVDD.n5126 DVDD.n5111 0.00476
R9024 DVDD.n5126 DVDD.n5125 0.00476
R9025 DVDD.n5125 DVDD.n5124 0.00476
R9026 DVDD.n5124 DVDD.n5117 0.00476
R9027 DVDD.n5120 DVDD.n5117 0.00476
R9028 DVDD.n5120 DVDD.n133 0.00476
R9029 DVDD.n5851 DVDD.n133 0.00476
R9030 DVDD.n5851 DVDD.n131 0.00476
R9031 DVDD.n5855 DVDD.n131 0.00476
R9032 DVDD.n5855 DVDD.n129 0.00476
R9033 DVDD.n5859 DVDD.n129 0.00476
R9034 DVDD.n5859 DVDD.n127 0.00476
R9035 DVDD.n5863 DVDD.n127 0.00476
R9036 DVDD.n5863 DVDD.n125 0.00476
R9037 DVDD.n5867 DVDD.n125 0.00476
R9038 DVDD.n5867 DVDD.n123 0.00476
R9039 DVDD.n5871 DVDD.n123 0.00476
R9040 DVDD.n5871 DVDD.n121 0.00476
R9041 DVDD.n5875 DVDD.n121 0.00476
R9042 DVDD.n5880 DVDD.n5879 0.00476
R9043 DVDD.n5882 DVDD.n5880 0.00476
R9044 DVDD.n5882 DVDD.n117 0.00476
R9045 DVDD.n5906 DVDD.n117 0.00476
R9046 DVDD.n5906 DVDD.n5905 0.00476
R9047 DVDD.n5905 DVDD.n5904 0.00476
R9048 DVDD.n5904 DVDD.n5888 0.00476
R9049 DVDD.n5900 DVDD.n5888 0.00476
R9050 DVDD.n5900 DVDD.n5899 0.00476
R9051 DVDD.n5899 DVDD.n5898 0.00476
R9052 DVDD.n3056 DVDD.n3055 0.00476
R9053 DVDD.n3056 DVDD.n3028 0.00476
R9054 DVDD.n3062 DVDD.n3029 0.00476
R9055 DVDD.n1929 DVDD.n1928 0.00476
R9056 DVDD.n1929 DVDD.n1925 0.00476
R9057 DVDD.n2052 DVDD.n2045 0.00476
R9058 DVDD.n2052 DVDD.n2043 0.00476
R9059 DVDD.n2056 DVDD.n2043 0.00476
R9060 DVDD.n3085 DVDD.n2028 0.00476
R9061 DVDD.n3081 DVDD.n2028 0.00476
R9062 DVDD.n3081 DVDD.n3080 0.00476
R9063 DVDD.n3080 DVDD.n3079 0.00476
R9064 DVDD.n3075 DVDD.n2033 0.00476
R9065 DVDD.n3075 DVDD.n3074 0.00476
R9066 DVDD.n3074 DVDD.n3073 0.00476
R9067 DVDD.n3073 DVDD.n3071 0.00476
R9068 DVDD.n3045 DVDD.n3039 0.00476
R9069 DVDD.n3045 DVDD.n3037 0.00476
R9070 DVDD.n3050 DVDD.n3037 0.00476
R9071 DVDD.n3050 DVDD.n3038 0.00476
R9072 DVDD.n3057 DVDD.n3033 0.00476
R9073 DVDD.n3057 DVDD.n3030 0.00476
R9074 DVDD.n3061 DVDD.n3030 0.00476
R9075 DVDD.n3061 DVDD.n3031 0.00476
R9076 DVDD.n1930 DVDD.n1927 0.00476
R9077 DVDD.n1931 DVDD.n1930 0.00476
R9078 DVDD.n3302 DVDD.n3301 0.00476
R9079 DVDD.n3302 DVDD.n3300 0.00476
R9080 DVDD.n3306 DVDD.n3300 0.00476
R9081 DVDD.n3615 DVDD.n3614 0.00476
R9082 DVDD.n3614 DVDD.n3102 0.00476
R9083 DVDD.n3610 DVDD.n3102 0.00476
R9084 DVDD.n3610 DVDD.n3609 0.00476
R9085 DVDD.n3608 DVDD.n3108 0.00476
R9086 DVDD.n3599 DVDD.n3108 0.00476
R9087 DVDD.n3599 DVDD.n3598 0.00476
R9088 DVDD.n3598 DVDD.n3118 0.00476
R9089 DVDD.n3586 DVDD.n3129 0.00476
R9090 DVDD.n3586 DVDD.n3585 0.00476
R9091 DVDD.n3585 DVDD.n3132 0.00476
R9092 DVDD.n3144 DVDD.n3132 0.00476
R9093 DVDD.n3574 DVDD.n3573 0.00476
R9094 DVDD.n3573 DVDD.n3149 0.00476
R9095 DVDD.n3566 DVDD.n3149 0.00476
R9096 DVDD.n3566 DVDD.n3565 0.00476
R9097 DVDD.n1942 DVDD.n1906 0.00476
R9098 DVDD.n1938 DVDD.n1906 0.00476
R9099 DVDD.n3613 DVDD.n3612 0.00476
R9100 DVDD.n3612 DVDD.n3611 0.00476
R9101 DVDD.n3611 DVDD.n3103 0.00476
R9102 DVDD.n3567 DVDD.n3562 0.00476
R9103 DVDD.n1941 DVDD.n1940 0.00476
R9104 DVDD.n1940 DVDD.n1939 0.00476
R9105 DVDD.n3400 DVDD.n3399 0.00476
R9106 DVDD.n3400 DVDD.n3215 0.00476
R9107 DVDD.n3406 DVDD.n3215 0.00476
R9108 DVDD.n3453 DVDD.n3183 0.00476
R9109 DVDD.n1949 DVDD.n1948 0.00476
R9110 DVDD.n1950 DVDD.n1949 0.00476
R9111 DVDD.n3256 DVDD.n3250 0.00476
R9112 DVDD.n3256 DVDD.n3251 0.00476
R9113 DVDD.n3252 DVDD.n3251 0.00476
R9114 DVDD.n3220 DVDD.n3219 0.00476
R9115 DVDD.n3401 DVDD.n3220 0.00476
R9116 DVDD.n3401 DVDD.n3216 0.00476
R9117 DVDD.n3405 DVDD.n3216 0.00476
R9118 DVDD.n3421 DVDD.n3214 0.00476
R9119 DVDD.n3421 DVDD.n3212 0.00476
R9120 DVDD.n3425 DVDD.n3212 0.00476
R9121 DVDD.n3426 DVDD.n3425 0.00476
R9122 DVDD.n3204 DVDD.n3203 0.00476
R9123 DVDD.n3448 DVDD.n3204 0.00476
R9124 DVDD.n3448 DVDD.n3199 0.00476
R9125 DVDD.n3462 DVDD.n3199 0.00476
R9126 DVDD.n3458 DVDD.n3201 0.00476
R9127 DVDD.n3458 DVDD.n3457 0.00476
R9128 DVDD.n3457 DVDD.n3456 0.00476
R9129 DVDD.n3456 DVDD.n3454 0.00476
R9130 DVDD.n1964 DVDD.n1963 0.00476
R9131 DVDD.n1963 DVDD.n1962 0.00476
R9132 DVDD.n3619 DVDD.n2021 0.00476
R9133 DVDD.n3623 DVDD.n2021 0.00476
R9134 DVDD.n3623 DVDD.n2019 0.00476
R9135 DVDD.n3630 DVDD.n2019 0.00476
R9136 DVDD.n3635 DVDD.n2017 0.00476
R9137 DVDD.n3635 DVDD.n2006 0.00476
R9138 DVDD.n3644 DVDD.n2006 0.00476
R9139 DVDD.n3645 DVDD.n3644 0.00476
R9140 DVDD.n3669 DVDD.n1978 0.00476
R9141 DVDD.n3669 DVDD.n1976 0.00476
R9142 DVDD.n3673 DVDD.n1976 0.00476
R9143 DVDD.n3673 DVDD.n1974 0.00476
R9144 DVDD.n3677 DVDD.n1972 0.00476
R9145 DVDD.n3681 DVDD.n1972 0.00476
R9146 DVDD.n3681 DVDD.n1970 0.00476
R9147 DVDD.n3685 DVDD.n1970 0.00476
R9148 DVDD.n3702 DVDD.n3688 0.00476
R9149 DVDD.n3698 DVDD.n3688 0.00476
R9150 DVDD.n3618 DVDD.n2020 0.00476
R9151 DVDD.n3624 DVDD.n2020 0.00476
R9152 DVDD.n3625 DVDD.n3624 0.00476
R9153 DVDD.n3629 DVDD.n3625 0.00476
R9154 DVDD.n3675 DVDD.n3674 0.00476
R9155 DVDD.n3676 DVDD.n1971 0.00476
R9156 DVDD.n3682 DVDD.n1971 0.00476
R9157 DVDD.n3683 DVDD.n3682 0.00476
R9158 DVDD.n3684 DVDD.n3683 0.00476
R9159 DVDD.n3701 DVDD.n3700 0.00476
R9160 DVDD.n3700 DVDD.n3699 0.00476
R9161 DVDD.n3733 DVDD.n3732 0.00476
R9162 DVDD.n3732 DVDD.n1855 0.00476
R9163 DVDD.n3781 DVDD.n1855 0.00476
R9164 DVDD.n3781 DVDD.n1853 0.00476
R9165 DVDD.n3785 DVDD.n1853 0.00476
R9166 DVDD.n3785 DVDD.n1851 0.00476
R9167 DVDD.n3789 DVDD.n1851 0.00476
R9168 DVDD.n3789 DVDD.n1849 0.00476
R9169 DVDD.n3793 DVDD.n1849 0.00476
R9170 DVDD.n3793 DVDD.n1847 0.00476
R9171 DVDD.n3798 DVDD.n1847 0.00476
R9172 DVDD.n3798 DVDD.n1845 0.00476
R9173 DVDD.n3802 DVDD.n1845 0.00476
R9174 DVDD.n3803 DVDD.n3802 0.00476
R9175 DVDD.n4256 DVDD.n1689 0.00476
R9176 DVDD.n4252 DVDD.n1689 0.00476
R9177 DVDD.n4252 DVDD.n4251 0.00476
R9178 DVDD.n4251 DVDD.n1694 0.00476
R9179 DVDD.n4247 DVDD.n1694 0.00476
R9180 DVDD.n4247 DVDD.n4246 0.00476
R9181 DVDD.n4246 DVDD.n1699 0.00476
R9182 DVDD.n4242 DVDD.n1699 0.00476
R9183 DVDD.n4242 DVDD.n4241 0.00476
R9184 DVDD.n4241 DVDD.n4240 0.00476
R9185 DVDD.n4240 DVDD.n1705 0.00476
R9186 DVDD.n3935 DVDD.n1705 0.00476
R9187 DVDD.n3956 DVDD.n3935 0.00476
R9188 DVDD.n3956 DVDD.n3955 0.00476
R9189 DVDD.n3955 DVDD.n3954 0.00476
R9190 DVDD.n3954 DVDD.n3941 0.00476
R9191 DVDD.n3949 DVDD.n3941 0.00476
R9192 DVDD.n3949 DVDD.n3948 0.00476
R9193 DVDD.n3948 DVDD.n3947 0.00476
R9194 DVDD.n3947 DVDD.n3926 0.00476
R9195 DVDD.n3969 DVDD.n3926 0.00476
R9196 DVDD.n3969 DVDD.n3924 0.00476
R9197 DVDD.n3973 DVDD.n3924 0.00476
R9198 DVDD.n3977 DVDD.n1816 0.00476
R9199 DVDD.n3981 DVDD.n1816 0.00476
R9200 DVDD.n3981 DVDD.n1814 0.00476
R9201 DVDD.n3985 DVDD.n1814 0.00476
R9202 DVDD.n3985 DVDD.n1812 0.00476
R9203 DVDD.n3989 DVDD.n1812 0.00476
R9204 DVDD.n3989 DVDD.n1810 0.00476
R9205 DVDD.n3997 DVDD.n1810 0.00476
R9206 DVDD.n3997 DVDD.n1808 0.00476
R9207 DVDD.n4001 DVDD.n1808 0.00476
R9208 DVDD.n4001 DVDD.n1806 0.00476
R9209 DVDD.n4005 DVDD.n1806 0.00476
R9210 DVDD.n4005 DVDD.n1804 0.00476
R9211 DVDD.n4009 DVDD.n1804 0.00476
R9212 DVDD.n4009 DVDD.n1802 0.00476
R9213 DVDD.n4017 DVDD.n1802 0.00476
R9214 DVDD.n4017 DVDD.n1800 0.00476
R9215 DVDD.n4021 DVDD.n1800 0.00476
R9216 DVDD.n4021 DVDD.n1798 0.00476
R9217 DVDD.n4026 DVDD.n1798 0.00476
R9218 DVDD.n4026 DVDD.n1796 0.00476
R9219 DVDD.n4030 DVDD.n1796 0.00476
R9220 DVDD.n4031 DVDD.n4030 0.00476
R9221 DVDD.n4117 DVDD.n1788 0.00476
R9222 DVDD.n4117 DVDD.n4116 0.00476
R9223 DVDD.n4116 DVDD.n4115 0.00476
R9224 DVDD.n4115 DVDD.n4107 0.00476
R9225 DVDD.n4110 DVDD.n4107 0.00476
R9226 DVDD.n4110 DVDD.n1783 0.00476
R9227 DVDD.n4129 DVDD.n1783 0.00476
R9228 DVDD.n4129 DVDD.n1781 0.00476
R9229 DVDD.n4133 DVDD.n1781 0.00476
R9230 DVDD.n4133 DVDD.n1779 0.00476
R9231 DVDD.n4141 DVDD.n1779 0.00476
R9232 DVDD.n4141 DVDD.n1777 0.00476
R9233 DVDD.n4145 DVDD.n1777 0.00476
R9234 DVDD.n4145 DVDD.n1776 0.00476
R9235 DVDD.n4151 DVDD.n1776 0.00476
R9236 DVDD.n4151 DVDD.n1774 0.00476
R9237 DVDD.n4155 DVDD.n1774 0.00476
R9238 DVDD.n4155 DVDD.n1772 0.00476
R9239 DVDD.n4161 DVDD.n1772 0.00476
R9240 DVDD.n4161 DVDD.n1770 0.00476
R9241 DVDD.n4165 DVDD.n1770 0.00476
R9242 DVDD.n4165 DVDD.n1768 0.00476
R9243 DVDD.n4169 DVDD.n1768 0.00476
R9244 DVDD.n4219 DVDD.n4172 0.00476
R9245 DVDD.n4215 DVDD.n4172 0.00476
R9246 DVDD.n4215 DVDD.n4214 0.00476
R9247 DVDD.n4214 DVDD.n4213 0.00476
R9248 DVDD.n4213 DVDD.n4180 0.00476
R9249 DVDD.n4209 DVDD.n4180 0.00476
R9250 DVDD.n4209 DVDD.n4208 0.00476
R9251 DVDD.n4208 DVDD.n4207 0.00476
R9252 DVDD.n4207 DVDD.n4186 0.00476
R9253 DVDD.n4193 DVDD.n4186 0.00476
R9254 DVDD.n4195 DVDD.n4190 0.00476
R9255 DVDD.n3780 DVDD.n3778 0.00476
R9256 DVDD.n3780 DVDD.n3779 0.00476
R9257 DVDD.n3787 DVDD.n3786 0.00476
R9258 DVDD.n3788 DVDD.n3787 0.00476
R9259 DVDD.n3788 DVDD.n1848 0.00476
R9260 DVDD.n3794 DVDD.n1848 0.00476
R9261 DVDD.n3795 DVDD.n3794 0.00476
R9262 DVDD.n3797 DVDD.n3795 0.00476
R9263 DVDD.n3797 DVDD.n3796 0.00476
R9264 DVDD.n3796 DVDD.n1844 0.00476
R9265 DVDD.n3804 DVDD.n1844 0.00476
R9266 DVDD.n4255 DVDD.n4254 0.00476
R9267 DVDD.n4254 DVDD.n4253 0.00476
R9268 DVDD.n4250 DVDD.n4249 0.00476
R9269 DVDD.n4249 DVDD.n4248 0.00476
R9270 DVDD.n4245 DVDD.n4244 0.00476
R9271 DVDD.n4244 DVDD.n4243 0.00476
R9272 DVDD.n4243 DVDD.n1700 0.00476
R9273 DVDD.n3933 DVDD.n1707 0.00476
R9274 DVDD.n3957 DVDD.n3934 0.00476
R9275 DVDD.n3953 DVDD.n3934 0.00476
R9276 DVDD.n3951 DVDD.n3950 0.00476
R9277 DVDD.n3950 DVDD.n3942 0.00476
R9278 DVDD.n3942 DVDD.n3927 0.00476
R9279 DVDD.n3968 DVDD.n3966 0.00476
R9280 DVDD.n3968 DVDD.n3967 0.00476
R9281 DVDD.n3976 DVDD.n1815 0.00476
R9282 DVDD.n3982 DVDD.n1815 0.00476
R9283 DVDD.n3983 DVDD.n3982 0.00476
R9284 DVDD.n3984 DVDD.n3983 0.00476
R9285 DVDD.n3984 DVDD.n1811 0.00476
R9286 DVDD.n3990 DVDD.n1811 0.00476
R9287 DVDD.n3991 DVDD.n3990 0.00476
R9288 DVDD.n3996 DVDD.n3991 0.00476
R9289 DVDD.n4002 DVDD.n1807 0.00476
R9290 DVDD.n4003 DVDD.n4002 0.00476
R9291 DVDD.n4004 DVDD.n4003 0.00476
R9292 DVDD.n4004 DVDD.n1803 0.00476
R9293 DVDD.n4010 DVDD.n1803 0.00476
R9294 DVDD.n4016 DVDD.n4015 0.00476
R9295 DVDD.n4016 DVDD.n1799 0.00476
R9296 DVDD.n4022 DVDD.n1799 0.00476
R9297 DVDD.n4023 DVDD.n4022 0.00476
R9298 DVDD.n4025 DVDD.n4023 0.00476
R9299 DVDD.n4025 DVDD.n4024 0.00476
R9300 DVDD.n4024 DVDD.n1795 0.00476
R9301 DVDD.n4032 DVDD.n1795 0.00476
R9302 DVDD.n4118 DVDD.n1787 0.00476
R9303 DVDD.n4114 DVDD.n1787 0.00476
R9304 DVDD.n4112 DVDD.n4111 0.00476
R9305 DVDD.n4111 DVDD.n1784 0.00476
R9306 DVDD.n4128 DVDD.n1784 0.00476
R9307 DVDD.n4134 DVDD.n1780 0.00476
R9308 DVDD.n4135 DVDD.n4134 0.00476
R9309 DVDD.n4140 DVDD.n4139 0.00476
R9310 DVDD.n4150 DVDD.n4149 0.00476
R9311 DVDD.n4150 DVDD.n1773 0.00476
R9312 DVDD.n4156 DVDD.n1773 0.00476
R9313 DVDD.n4160 DVDD.n4158 0.00476
R9314 DVDD.n4160 DVDD.n4159 0.00476
R9315 DVDD.n4167 DVDD.n4166 0.00476
R9316 DVDD.n4168 DVDD.n4167 0.00476
R9317 DVDD.n4218 DVDD.n4217 0.00476
R9318 DVDD.n4217 DVDD.n4216 0.00476
R9319 DVDD.n4216 DVDD.n4176 0.00476
R9320 DVDD.n4212 DVDD.n4176 0.00476
R9321 DVDD.n4212 DVDD.n4211 0.00476
R9322 DVDD.n4211 DVDD.n4210 0.00476
R9323 DVDD.n4210 DVDD.n4181 0.00476
R9324 DVDD.n4206 DVDD.n4181 0.00476
R9325 DVDD.n4206 DVDD.n4205 0.00476
R9326 DVDD.n4194 DVDD.n4189 0.00476
R9327 DVDD.n1176 DVDD.n1131 0.00476
R9328 DVDD.n1176 DVDD.n1175 0.00476
R9329 DVDD.n1175 DVDD.n1174 0.00476
R9330 DVDD.n1174 DVDD.n1155 0.00476
R9331 DVDD.n1170 DVDD.n1155 0.00476
R9332 DVDD.n1170 DVDD.n1169 0.00476
R9333 DVDD.n1169 DVDD.n1168 0.00476
R9334 DVDD.n1168 DVDD.n1161 0.00476
R9335 DVDD.n5398 DVDD.n360 0.00476
R9336 DVDD.n5394 DVDD.n360 0.00476
R9337 DVDD.n5394 DVDD.n5393 0.00476
R9338 DVDD.n5393 DVDD.n5392 0.00476
R9339 DVDD.n5392 DVDD.n365 0.00476
R9340 DVDD.n5388 DVDD.n365 0.00476
R9341 DVDD.n5388 DVDD.n5387 0.00476
R9342 DVDD.n5387 DVDD.n5386 0.00476
R9343 DVDD.n5386 DVDD.n371 0.00476
R9344 DVDD.n5382 DVDD.n371 0.00476
R9345 DVDD.n5378 DVDD.n382 0.00476
R9346 DVDD.n5374 DVDD.n382 0.00476
R9347 DVDD.n5374 DVDD.n5373 0.00476
R9348 DVDD.n5373 DVDD.n5372 0.00476
R9349 DVDD.n5372 DVDD.n388 0.00476
R9350 DVDD.n5368 DVDD.n388 0.00476
R9351 DVDD.n5368 DVDD.n5367 0.00476
R9352 DVDD.n5367 DVDD.n5366 0.00476
R9353 DVDD.n5366 DVDD.n394 0.00476
R9354 DVDD.n5362 DVDD.n394 0.00476
R9355 DVDD.n5358 DVDD.n406 0.00476
R9356 DVDD.n5354 DVDD.n406 0.00476
R9357 DVDD.n5354 DVDD.n5353 0.00476
R9358 DVDD.n5353 DVDD.n5352 0.00476
R9359 DVDD.n5352 DVDD.n412 0.00476
R9360 DVDD.n5348 DVDD.n412 0.00476
R9361 DVDD.n5348 DVDD.n5347 0.00476
R9362 DVDD.n5347 DVDD.n5346 0.00476
R9363 DVDD.n5346 DVDD.n418 0.00476
R9364 DVDD.n5342 DVDD.n418 0.00476
R9365 DVDD.n5342 DVDD.n5341 0.00476
R9366 DVDD.n5337 DVDD.n429 0.00476
R9367 DVDD.n5333 DVDD.n429 0.00476
R9368 DVDD.n5333 DVDD.n5332 0.00476
R9369 DVDD.n5332 DVDD.n5331 0.00476
R9370 DVDD.n5331 DVDD.n437 0.00476
R9371 DVDD.n5327 DVDD.n437 0.00476
R9372 DVDD.n5327 DVDD.n5326 0.00476
R9373 DVDD.n5326 DVDD.n5325 0.00476
R9374 DVDD.n5325 DVDD.n443 0.00476
R9375 DVDD.n5321 DVDD.n443 0.00476
R9376 DVDD.n5133 DVDD.n5105 0.00476
R9377 DVDD.n5129 DVDD.n5105 0.00476
R9378 DVDD.n5129 DVDD.n5128 0.00476
R9379 DVDD.n5128 DVDD.n5127 0.00476
R9380 DVDD.n5127 DVDD.n5112 0.00476
R9381 DVDD.n5123 DVDD.n5112 0.00476
R9382 DVDD.n5123 DVDD.n5122 0.00476
R9383 DVDD.n5122 DVDD.n5121 0.00476
R9384 DVDD.n5121 DVDD.n134 0.00476
R9385 DVDD.n5850 DVDD.n134 0.00476
R9386 DVDD.n5857 DVDD.n5856 0.00476
R9387 DVDD.n5858 DVDD.n5857 0.00476
R9388 DVDD.n5858 DVDD.n126 0.00476
R9389 DVDD.n5864 DVDD.n126 0.00476
R9390 DVDD.n5865 DVDD.n5864 0.00476
R9391 DVDD.n5866 DVDD.n5865 0.00476
R9392 DVDD.n5866 DVDD.n122 0.00476
R9393 DVDD.n5872 DVDD.n122 0.00476
R9394 DVDD.n5873 DVDD.n5872 0.00476
R9395 DVDD.n5874 DVDD.n5873 0.00476
R9396 DVDD.n5907 DVDD.n115 0.00476
R9397 DVDD.n5903 DVDD.n115 0.00476
R9398 DVDD.n5903 DVDD.n5902 0.00476
R9399 DVDD.n5902 DVDD.n5901 0.00476
R9400 DVDD.n5901 DVDD.n5889 0.00476
R9401 DVDD.n5897 DVDD.n5889 0.00476
R9402 DVDD.n4415 DVDD.n1104 0.00476
R9403 DVDD.n4421 DVDD.n1104 0.00476
R9404 DVDD.n4422 DVDD.n4421 0.00476
R9405 DVDD.n4423 DVDD.n4422 0.00476
R9406 DVDD.n4423 DVDD.n1100 0.00476
R9407 DVDD.n4429 DVDD.n1100 0.00476
R9408 DVDD.n4430 DVDD.n4429 0.00476
R9409 DVDD.n4431 DVDD.n4430 0.00476
R9410 DVDD.n4444 DVDD.n4443 0.00476
R9411 DVDD.n4444 DVDD.n1092 0.00476
R9412 DVDD.n4450 DVDD.n1092 0.00476
R9413 DVDD.n4451 DVDD.n4450 0.00476
R9414 DVDD.n4452 DVDD.n4451 0.00476
R9415 DVDD.n4452 DVDD.n1088 0.00476
R9416 DVDD.n4458 DVDD.n1088 0.00476
R9417 DVDD.n4459 DVDD.n4458 0.00476
R9418 DVDD.n4460 DVDD.n4459 0.00476
R9419 DVDD.n4460 DVDD.n1075 0.00476
R9420 DVDD.n4494 DVDD.n4493 0.00476
R9421 DVDD.n4493 DVDD.n4492 0.00476
R9422 DVDD.n4492 DVDD.n4467 0.00476
R9423 DVDD.n4488 DVDD.n4467 0.00476
R9424 DVDD.n4488 DVDD.n4487 0.00476
R9425 DVDD.n4487 DVDD.n4486 0.00476
R9426 DVDD.n4486 DVDD.n4473 0.00476
R9427 DVDD.n4482 DVDD.n4473 0.00476
R9428 DVDD.n4482 DVDD.n4481 0.00476
R9429 DVDD.n4481 DVDD.n4480 0.00476
R9430 DVDD.n4887 DVDD.n4886 0.00476
R9431 DVDD.n4888 DVDD.n4887 0.00476
R9432 DVDD.n4888 DVDD.n691 0.00476
R9433 DVDD.n4894 DVDD.n691 0.00476
R9434 DVDD.n4895 DVDD.n4894 0.00476
R9435 DVDD.n4896 DVDD.n4895 0.00476
R9436 DVDD.n4896 DVDD.n687 0.00476
R9437 DVDD.n4902 DVDD.n687 0.00476
R9438 DVDD.n4903 DVDD.n4902 0.00476
R9439 DVDD.n4904 DVDD.n4903 0.00476
R9440 DVDD.n4904 DVDD.n674 0.00476
R9441 DVDD.n4935 DVDD.n4934 0.00476
R9442 DVDD.n4934 DVDD.n4933 0.00476
R9443 DVDD.n4933 DVDD.n4911 0.00476
R9444 DVDD.n4929 DVDD.n4911 0.00476
R9445 DVDD.n4929 DVDD.n4928 0.00476
R9446 DVDD.n4928 DVDD.n4927 0.00476
R9447 DVDD.n4927 DVDD.n4917 0.00476
R9448 DVDD.n4923 DVDD.n4917 0.00476
R9449 DVDD.n4923 DVDD.n4922 0.00476
R9450 DVDD.n4922 DVDD.n451 0.00476
R9451 DVDD.n5315 DVDD.n475 0.00476
R9452 DVDD.n5311 DVDD.n475 0.00476
R9453 DVDD.n5311 DVDD.n5310 0.00476
R9454 DVDD.n5310 DVDD.n5309 0.00476
R9455 DVDD.n5309 DVDD.n5255 0.00476
R9456 DVDD.n5305 DVDD.n5255 0.00476
R9457 DVDD.n5305 DVDD.n5304 0.00476
R9458 DVDD.n5304 DVDD.n5303 0.00476
R9459 DVDD.n5303 DVDD.n5261 0.00476
R9460 DVDD.n5299 DVDD.n5261 0.00476
R9461 DVDD.n5295 DVDD.n155 0.00476
R9462 DVDD.n5295 DVDD.n5294 0.00476
R9463 DVDD.n5294 DVDD.n5293 0.00476
R9464 DVDD.n5293 DVDD.n5270 0.00476
R9465 DVDD.n5289 DVDD.n5270 0.00476
R9466 DVDD.n5289 DVDD.n5288 0.00476
R9467 DVDD.n5288 DVDD.n5287 0.00476
R9468 DVDD.n5287 DVDD.n5276 0.00476
R9469 DVDD.n5283 DVDD.n5276 0.00476
R9470 DVDD.n5283 DVDD.n42 0.00476
R9471 DVDD.n5601 DVDD.n5575 0.00476
R9472 DVDD.n5597 DVDD.n5575 0.00476
R9473 DVDD.n5597 DVDD.n5596 0.00476
R9474 DVDD.n5596 DVDD.n5595 0.00476
R9475 DVDD.n5595 DVDD.n5583 0.00476
R9476 DVDD.n5591 DVDD.n5583 0.00476
R9477 DVDD.n4368 DVDD.n1607 0.00476
R9478 DVDD.n4368 DVDD.n4367 0.00476
R9479 DVDD.n4367 DVDD.n4366 0.00476
R9480 DVDD.n4366 DVDD.n4350 0.00476
R9481 DVDD.n4362 DVDD.n4350 0.00476
R9482 DVDD.n4362 DVDD.n4361 0.00476
R9483 DVDD.n4361 DVDD.n4360 0.00476
R9484 DVDD.n4360 DVDD.n975 0.00476
R9485 DVDD.n4633 DVDD.n4632 0.00476
R9486 DVDD.n4632 DVDD.n4631 0.00476
R9487 DVDD.n4631 DVDD.n993 0.00476
R9488 DVDD.n4627 DVDD.n993 0.00476
R9489 DVDD.n4627 DVDD.n4626 0.00476
R9490 DVDD.n4626 DVDD.n4625 0.00476
R9491 DVDD.n4625 DVDD.n999 0.00476
R9492 DVDD.n4621 DVDD.n999 0.00476
R9493 DVDD.n4621 DVDD.n4620 0.00476
R9494 DVDD.n4620 DVDD.n4619 0.00476
R9495 DVDD.n1046 DVDD.n1045 0.00476
R9496 DVDD.n1045 DVDD.n1020 0.00476
R9497 DVDD.n1041 DVDD.n1020 0.00476
R9498 DVDD.n1041 DVDD.n1040 0.00476
R9499 DVDD.n1040 DVDD.n1039 0.00476
R9500 DVDD.n1039 DVDD.n1026 0.00476
R9501 DVDD.n1035 DVDD.n1026 0.00476
R9502 DVDD.n1035 DVDD.n1034 0.00476
R9503 DVDD.n1034 DVDD.n728 0.00476
R9504 DVDD.n4874 DVDD.n728 0.00476
R9505 DVDD.n4868 DVDD.n715 0.00476
R9506 DVDD.n4868 DVDD.n4867 0.00476
R9507 DVDD.n4867 DVDD.n4866 0.00476
R9508 DVDD.n4866 DVDD.n4806 0.00476
R9509 DVDD.n4862 DVDD.n4806 0.00476
R9510 DVDD.n4862 DVDD.n4861 0.00476
R9511 DVDD.n4861 DVDD.n4860 0.00476
R9512 DVDD.n4860 DVDD.n4812 0.00476
R9513 DVDD.n4856 DVDD.n4812 0.00476
R9514 DVDD.n4856 DVDD.n4855 0.00476
R9515 DVDD.n4855 DVDD.n605 0.00476
R9516 DVDD.n4850 DVDD.n4849 0.00476
R9517 DVDD.n4849 DVDD.n4848 0.00476
R9518 DVDD.n4848 DVDD.n4822 0.00476
R9519 DVDD.n4844 DVDD.n4822 0.00476
R9520 DVDD.n4844 DVDD.n4843 0.00476
R9521 DVDD.n4843 DVDD.n4842 0.00476
R9522 DVDD.n4842 DVDD.n4828 0.00476
R9523 DVDD.n4838 DVDD.n4828 0.00476
R9524 DVDD.n4838 DVDD.n4837 0.00476
R9525 DVDD.n4837 DVDD.n4836 0.00476
R9526 DVDD.n555 DVDD.n554 0.00476
R9527 DVDD.n554 DVDD.n496 0.00476
R9528 DVDD.n550 DVDD.n496 0.00476
R9529 DVDD.n550 DVDD.n549 0.00476
R9530 DVDD.n549 DVDD.n548 0.00476
R9531 DVDD.n548 DVDD.n502 0.00476
R9532 DVDD.n544 DVDD.n502 0.00476
R9533 DVDD.n544 DVDD.n543 0.00476
R9534 DVDD.n543 DVDD.n542 0.00476
R9535 DVDD.n542 DVDD.n170 0.00476
R9536 DVDD.n537 DVDD.n536 0.00476
R9537 DVDD.n536 DVDD.n535 0.00476
R9538 DVDD.n535 DVDD.n514 0.00476
R9539 DVDD.n531 DVDD.n514 0.00476
R9540 DVDD.n531 DVDD.n530 0.00476
R9541 DVDD.n530 DVDD.n529 0.00476
R9542 DVDD.n529 DVDD.n520 0.00476
R9543 DVDD.n525 DVDD.n520 0.00476
R9544 DVDD.n525 DVDD.n39 0.00476
R9545 DVDD.n5939 DVDD.n39 0.00476
R9546 DVDD.n5956 DVDD.n5955 0.00476
R9547 DVDD.n5956 DVDD.n3 0.00476
R9548 DVDD.n5963 DVDD.n3 0.00476
R9549 DVDD.n5964 DVDD.n5963 0.00476
R9550 DVDD.n5965 DVDD.n5964 0.00476
R9551 DVDD.n5965 DVDD.n0 0.00476
R9552 DVDD.n4325 DVDD.n1639 0.00476
R9553 DVDD.n4325 DVDD.n4324 0.00476
R9554 DVDD.n4324 DVDD.n4323 0.00476
R9555 DVDD.n4323 DVDD.n4305 0.00476
R9556 DVDD.n4319 DVDD.n4305 0.00476
R9557 DVDD.n4319 DVDD.n4318 0.00476
R9558 DVDD.n4318 DVDD.n4317 0.00476
R9559 DVDD.n4317 DVDD.n4311 0.00476
R9560 DVDD.n4719 DVDD.n905 0.00476
R9561 DVDD.n4725 DVDD.n905 0.00476
R9562 DVDD.n4726 DVDD.n4725 0.00476
R9563 DVDD.n4727 DVDD.n4726 0.00476
R9564 DVDD.n4727 DVDD.n901 0.00476
R9565 DVDD.n4733 DVDD.n901 0.00476
R9566 DVDD.n4734 DVDD.n4733 0.00476
R9567 DVDD.n4735 DVDD.n4734 0.00476
R9568 DVDD.n4735 DVDD.n897 0.00476
R9569 DVDD.n4741 DVDD.n897 0.00476
R9570 DVDD.n4745 DVDD.n887 0.00476
R9571 DVDD.n4751 DVDD.n887 0.00476
R9572 DVDD.n4752 DVDD.n4751 0.00476
R9573 DVDD.n4753 DVDD.n4752 0.00476
R9574 DVDD.n4753 DVDD.n883 0.00476
R9575 DVDD.n4759 DVDD.n883 0.00476
R9576 DVDD.n4760 DVDD.n4759 0.00476
R9577 DVDD.n4761 DVDD.n4760 0.00476
R9578 DVDD.n4761 DVDD.n879 0.00476
R9579 DVDD.n4769 DVDD.n879 0.00476
R9580 DVDD.n4800 DVDD.n4799 0.00476
R9581 DVDD.n4799 DVDD.n4798 0.00476
R9582 DVDD.n4798 DVDD.n4774 0.00476
R9583 DVDD.n4794 DVDD.n4774 0.00476
R9584 DVDD.n4794 DVDD.n4793 0.00476
R9585 DVDD.n4793 DVDD.n4792 0.00476
R9586 DVDD.n4792 DVDD.n4780 0.00476
R9587 DVDD.n4788 DVDD.n4780 0.00476
R9588 DVDD.n4788 DVDD.n4787 0.00476
R9589 DVDD.n4787 DVDD.n588 0.00476
R9590 DVDD.n5021 DVDD.n588 0.00476
R9591 DVDD.n5028 DVDD.n5027 0.00476
R9592 DVDD.n5029 DVDD.n5028 0.00476
R9593 DVDD.n5029 DVDD.n580 0.00476
R9594 DVDD.n5035 DVDD.n580 0.00476
R9595 DVDD.n5036 DVDD.n5035 0.00476
R9596 DVDD.n5037 DVDD.n5036 0.00476
R9597 DVDD.n5037 DVDD.n576 0.00476
R9598 DVDD.n5043 DVDD.n576 0.00476
R9599 DVDD.n5044 DVDD.n5043 0.00476
R9600 DVDD.n5045 DVDD.n5044 0.00476
R9601 DVDD.n5082 DVDD.n5081 0.00476
R9602 DVDD.n5081 DVDD.n5080 0.00476
R9603 DVDD.n5080 DVDD.n5052 0.00476
R9604 DVDD.n5076 DVDD.n5052 0.00476
R9605 DVDD.n5076 DVDD.n5075 0.00476
R9606 DVDD.n5075 DVDD.n5074 0.00476
R9607 DVDD.n5074 DVDD.n5058 0.00476
R9608 DVDD.n5070 DVDD.n5058 0.00476
R9609 DVDD.n5070 DVDD.n5069 0.00476
R9610 DVDD.n5069 DVDD.n5068 0.00476
R9611 DVDD.n5727 DVDD.n199 0.00476
R9612 DVDD.n5723 DVDD.n199 0.00476
R9613 DVDD.n5723 DVDD.n5722 0.00476
R9614 DVDD.n5722 DVDD.n5721 0.00476
R9615 DVDD.n5721 DVDD.n205 0.00476
R9616 DVDD.n5717 DVDD.n205 0.00476
R9617 DVDD.n5717 DVDD.n5716 0.00476
R9618 DVDD.n5716 DVDD.n5715 0.00476
R9619 DVDD.n5715 DVDD.n211 0.00476
R9620 DVDD.n5711 DVDD.n211 0.00476
R9621 DVDD.n5696 DVDD.n234 0.00476
R9622 DVDD.n5696 DVDD.n5695 0.00476
R9623 DVDD.n5695 DVDD.n5694 0.00476
R9624 DVDD.n5694 DVDD.n5679 0.00476
R9625 DVDD.n5690 DVDD.n5679 0.00476
R9626 DVDD.n5690 DVDD.n5689 0.00476
R9627 DVDD.n3345 DVDD.n3344 0.00473767
R9628 DVDD.n3392 DVDD.n3221 0.00473767
R9629 DVDD.n5340 DVDD.n426 0.00473
R9630 DVDD.n5338 DVDD.n5337 0.00473
R9631 DVDD.n5004 DVDD.n4938 0.00473
R9632 DVDD.n4935 DVDD.n672 0.00473
R9633 DVDD.n5012 DVDD.n616 0.00473
R9634 DVDD.n4850 DVDD.n603 0.00473
R9635 DVDD.n5020 DVDD.n591 0.00473
R9636 DVDD.n5027 DVDD.n584 0.00473
R9637 DVDD.n4079 DVDD.n4040 0.0047
R9638 DVDD.n2063 DVDD.n2035 0.00467
R9639 DVDD.n2061 DVDD.n2036 0.00467
R9640 DVDD.n2038 DVDD.n2037 0.00467
R9641 DVDD.n3070 DVDD.n3069 0.00467
R9642 DVDD.n3044 DVDD.n3040 0.00467
R9643 DVDD.n3043 DVDD.n3041 0.00467
R9644 DVDD.n3051 DVDD.n3036 0.00467
R9645 DVDD.n3052 DVDD.n3034 0.00467
R9646 DVDD.n4102 DVDD.n4101 0.004625
R9647 DVDD.n3606 DVDD.n3109 0.00461
R9648 DVDD.n3601 DVDD.n3600 0.00461
R9649 DVDD.n3597 DVDD.n3114 0.00461
R9650 DVDD.n3596 DVDD.n3119 0.00461
R9651 DVDD.n3588 DVDD.n3587 0.00461
R9652 DVDD.n3584 DVDD.n3128 0.00461
R9653 DVDD.n3583 DVDD.n3133 0.00461
R9654 DVDD.n3142 DVDD.n3141 0.00461
R9655 DVDD.n3420 DVDD.n3408 0.00461
R9656 DVDD.n3419 DVDD.n3410 0.00461
R9657 DVDD.n3409 DVDD.n3211 0.00461
R9658 DVDD.n3428 DVDD.n3427 0.00461
R9659 DVDD.n3438 DVDD.n3437 0.00461
R9660 DVDD.n3447 DVDD.n3205 0.00461
R9661 DVDD.n3446 DVDD.n3197 0.00461
R9662 DVDD.n3464 DVDD.n3463 0.00461
R9663 DVDD.n5418 DVDD.n260 0.0045724
R9664 DVDD.n261 DVDD.n260 0.0045724
R9665 DVDD.n5797 DVDD.n153 0.00455738
R9666 DVDD.n5153 DVDD.n452 0.00455738
R9667 DVDD.n4985 DVDD.n675 0.00455738
R9668 DVDD.n777 DVDD.n776 0.00455738
R9669 DVDD.n4541 DVDD.n1076 0.00455738
R9670 DVDD.n3953 DVDD.n3952 0.00455
R9671 DVDD.n83 DVDD.n81 0.00452754
R9672 DVDD.n5550 DVDD.n16 0.00452754
R9673 DVDD.n5656 DVDD.n8 0.00452754
R9674 DVDD.n4662 DVDD.n983 0.00452754
R9675 DVDD.n5482 DVDD.n267 0.00452754
R9676 DVDD.n5426 DVDD.n5425 0.00452754
R9677 DVDD.n4765 DVDD.n697 0.0045
R9678 DVDD.n5048 DVDD.n477 0.0045
R9679 DVDD.n4440 DVDD.n1094 0.0045
R9680 DVDD.n4883 DVDD.n697 0.0045
R9681 DVDD.n4440 DVDD.n1095 0.0045
R9682 DVDD.n4883 DVDD.n699 0.0045
R9683 DVDD.n5877 DVDD.n35 0.0045
R9684 DVDD.n5249 DVDD.n477 0.0045
R9685 DVDD.n5249 DVDD.n478 0.0045
R9686 DVDD.n5942 DVDD.n34 0.0045
R9687 DVDD.n5942 DVDD.n35 0.0045
R9688 DVDD.n1094 DVDD.n907 0.0045
R9689 DVDD.n5910 DVDD.n98 0.0044433
R9690 DVDD.n114 DVDD.n88 0.0044433
R9691 DVDD.n5413 DVDD.n337 0.0044433
R9692 DVDD.n5410 DVDD.n334 0.0044433
R9693 DVDD.n936 DVDD.n926 0.0044433
R9694 DVDD.n955 DVDD.n919 0.0044433
R9695 DVDD.n242 DVDD.n232 0.0044433
R9696 DVDD.n250 DVDD.n238 0.0044433
R9697 DVDD.n2047 DVDD.n2046 0.00443
R9698 DVDD.n2051 DVDD.n2049 0.00443
R9699 DVDD.n2050 DVDD.n2042 0.00443
R9700 DVDD.n2058 DVDD.n2057 0.00443
R9701 DVDD.n2070 DVDD.n2027 0.00443
R9702 DVDD.n2071 DVDD.n2030 0.00443
R9703 DVDD.n2068 DVDD.n2031 0.00443
R9704 DVDD.n2066 DVDD.n2032 0.00443
R9705 DVDD.n3572 DVDD.n3143 0.00443
R9706 DVDD.n3571 DVDD.n3159 0.00443
R9707 DVDD.n3568 DVDD.n3567 0.00443
R9708 DVDD.n3452 DVDD.n3172 0.00443
R9709 DVDD.n3173 DVDD.n3171 0.00443
R9710 DVDD.n3513 DVDD.n3183 0.00443
R9711 DVDD.n4127 DVDD.n1780 0.00443
R9712 DVDD.n2558 DVDD.n2263 0.00442143
R9713 DVDD.n2800 DVDD.n2703 0.00441304
R9714 DVDD.n1740 DVDD.n1737 0.0044
R9715 DVDD.n4014 DVDD.n4010 0.00437
R9716 DVDD.n5850 DVDD.n5849 0.00437
R9717 DVDD.n137 DVDD.n130 0.00437
R9718 DVDD.n5299 DVDD.n143 0.00437
R9719 DVDD.n5834 DVDD.n144 0.00437
R9720 DVDD.n5783 DVDD.n170 0.00437
R9721 DVDD.n180 DVDD.n169 0.00437
R9722 DVDD.n5068 DVDD.n196 0.00437
R9723 DVDD.n5733 DVDD.n197 0.00437
R9724 DVDD.n333 DVDD.n332 0.00434971
R9725 DVDD.n85 DVDD.n75 0.00434083
R9726 DVDD.n3920 DVDD.n1817 0.004325
R9727 DVDD.n3063 DVDD.n3062 0.00431
R9728 DVDD.n5381 DVDD.n379 0.00431
R9729 DVDD.n5379 DVDD.n5378 0.00431
R9730 DVDD.n4560 DVDD.n4497 0.00431
R9731 DVDD.n4494 DVDD.n1073 0.00431
R9732 DVDD.n4616 DVDD.n1005 0.00431
R9733 DVDD.n4615 DVDD.n1046 0.00431
R9734 DVDD.n4742 DVDD.n891 0.00431
R9735 DVDD.n4745 DVDD.n4744 0.00431
R9736 DVDD.n2541 DVDD.n2300 0.00429286
R9737 DVDD.n3752 DVDD.n3734 0.00425
R9738 DVDD.n3777 DVDD.n1856 0.00425
R9739 DVDD.n3995 DVDD.n1807 0.00425
R9740 DVDD.n1579 DVDD.n1181 0.00425
R9741 DVDD.n1582 DVDD.n1121 0.00425
R9742 DVDD.n4410 DVDD.n4398 0.00425
R9743 DVDD.n4414 DVDD.n1108 0.00425
R9744 DVDD.n4383 DVDD.n4373 0.00425
R9745 DVDD.n4386 DVDD.n1596 0.00425
R9746 DVDD.n4340 DVDD.n4330 0.00425
R9747 DVDD.n4343 DVDD.n1628 0.00425
R9748 DVDD.n5533 DVDD.n23 0.00421773
R9749 DVDD.n4679 DVDD.n4650 0.00421773
R9750 DVDD.n4148 DVDD.n4146 0.00419
R9751 DVDD.n4198 DVDD.n4189 0.00419
R9752 DVDD.n5782 DVDD.n5781 0.00418852
R9753 DVDD.n5208 DVDD.n559 0.00418852
R9754 DVDD.n659 DVDD.n625 0.00418852
R9755 DVDD.n834 DVDD.n719 0.00418852
R9756 DVDD.n4581 DVDD.n1050 0.00418852
R9757 DVDD.n3487 DVDD.n3188 0.00416848
R9758 DVDD.n3544 DVDD.n3166 0.00416848
R9759 DVDD.n3649 DVDD 0.00408591
R9760 DVDD.n4239 DVDD.n1706 0.00407
R9761 DVDD.n4239 DVDD.n4238 0.00407
R9762 DVDD.n5710 DVDD.n5709 0.00404
R9763 DVDD.n38 DVDD.n33 0.00404
R9764 DVDD.n5935 DVDD.n44 0.00404
R9765 DVDD.n5879 DVDD.n119 0.00404
R9766 DVDD.n4219 DVDD.n1724 0.00404
R9767 DVDD.n80 DVDD.n41 0.00404
R9768 DVDD.n5937 DVDD.n5936 0.00404
R9769 DVDD.n5938 DVDD.n32 0.00404
R9770 DVDD.n5708 DVDD.n40 0.00404
R9771 DVDD.n4258 DVDD.n1686 0.004025
R9772 DVDD.n4146 DVDD.n1712 0.00395
R9773 DVDD DVDD.n5684 0.00392
R9774 DVDD.n5967 DVDD 0.00392
R9775 DVDD.n5592 DVDD 0.00392
R9776 DVDD.n5898 DVDD 0.00392
R9777 DVDD DVDD.n4193 0.00392
R9778 DVDD DVDD.n4187 0.00392
R9779 DVDD.n5897 DVDD 0.00392
R9780 DVDD.n5591 DVDD 0.00392
R9781 DVDD DVDD.n0 0.00392
R9782 DVDD.n5689 DVDD 0.00392
R9783 DVDD.n5517 DVDD.n9 0.00390792
R9784 DVDD.n4696 DVDD.n976 0.00390792
R9785 DVDD.n3642 DVDD.n2008 0.00386
R9786 DVDD.n3664 DVDD.n1975 0.00386
R9787 DVDD.n5084 DVDD.n481 0.0038
R9788 DVDD.n5245 DVDD.n5244 0.0038
R9789 DVDD.n5246 DVDD.n476 0.0038
R9790 DVDD.n5106 DVDD.n448 0.0038
R9791 DVDD.n1792 DVDD.n1788 0.0038
R9792 DVDD.n4033 DVDD.n1786 0.0038
R9793 DVDD.n2342 DVDD.n2333 0.00377857
R9794 DVDD.n2483 DVDD.n2327 0.00377857
R9795 DVDD.n2360 DVDD.n2328 0.00377857
R9796 DVDD.n3617 DVDD 0.00376574
R9797 DVDD DVDD.n2023 0.00376574
R9798 DVDD DVDD.n1897 0.00376574
R9799 DVDD DVDD.n1896 0.00376574
R9800 DVDD.n3368 DVDD.n3274 0.00374
R9801 DVDD.n3296 DVDD.n3281 0.00374
R9802 DVDD.n3361 DVDD.n3295 0.00374
R9803 DVDD.n3358 DVDD.n3307 0.00374
R9804 DVDD.n3613 DVDD.n3099 0.00374
R9805 DVDD.n3372 DVDD.n3248 0.00374
R9806 DVDD.n3267 DVDD.n3257 0.00374
R9807 DVDD.n3261 DVDD.n3229 0.00374
R9808 DVDD.n3389 DVDD.n3230 0.00374
R9809 DVDD.n3399 DVDD.n3398 0.00374
R9810 DVDD.n3626 DVDD.n2016 0.00371
R9811 DVDD.n3478 DVDD.n3186 0.00367935
R9812 DVDD.n3570 DVDD.n3561 0.00367935
R9813 DVDD.n4077 DVDD.n4044 0.00365
R9814 DVDD.n4081 DVDD.n4042 0.00365
R9815 DVDD.n4159 DVDD.n1769 0.00365
R9816 DVDD.n5611 DVDD.n5574 0.00359811
R9817 DVDD.n5436 DVDD.n283 0.00359811
R9818 DVDD.n3667 DVDD.n1980 0.00359
R9819 DVDD.n4248 DVDD.n1695 0.00359
R9820 DVDD.n350 DVDD.n340 0.00357827
R9821 DVDD.n5420 DVDD.n351 0.00357827
R9822 DVDD.n106 DVDD.n105 0.00357827
R9823 DVDD.n5917 DVDD.n87 0.00357827
R9824 DVDD.n351 DVDD.n350 0.00357827
R9825 DVDD.n105 DVDD.n87 0.00357827
R9826 DVDD.n5422 DVDD.n340 0.00357827
R9827 DVDD.n5915 DVDD.n106 0.00357827
R9828 DVDD.n4802 DVDD.n4801 0.00356
R9829 DVDD.n4871 DVDD.n4870 0.00356
R9830 DVDD.n4885 DVDD.n696 0.00356
R9831 DVDD.n5357 DVDD.n407 0.00356
R9832 DVDD.n3977 DVDD.n1818 0.00356
R9833 DVDD.n3976 DVDD.n3975 0.00356
R9834 DVDD.n4250 DVDD.n1691 0.00353
R9835 DVDD.n4119 DVDD.n1786 0.00353
R9836 DVDD.n4158 DVDD.n4157 0.00347
R9837 DVDD.n191 DVDD.n178 0.00345082
R9838 DVDD.n5207 DVDD.n493 0.00345082
R9839 DVDD.n660 DVDD.n614 0.00345082
R9840 DVDD.n833 DVDD.n712 0.00345082
R9841 DVDD.n4580 DVDD.n1017 0.00345082
R9842 DVDD.n3603 DVDD.n3602 0.00343478
R9843 DVDD.n3418 DVDD.n3411 0.00343478
R9844 DVDD.n3974 DVDD.n3923 0.00341
R9845 DVDD.n3643 DVDD.n2007 0.00335
R9846 DVDD.n1152 DVDD.n1151 0.00334
R9847 DVDD.n1153 DVDD.n1152 0.00334
R9848 DVDD.n1156 DVDD.n1153 0.00334
R9849 DVDD.n1157 DVDD.n1156 0.00334
R9850 DVDD.n1158 DVDD.n1157 0.00334
R9851 DVDD.n1159 DVDD.n1158 0.00334
R9852 DVDD.n1162 DVDD.n1159 0.00334
R9853 DVDD.n1163 DVDD.n1162 0.00334
R9854 DVDD.n1165 DVDD.n1163 0.00334
R9855 DVDD.n1165 DVDD.n1164 0.00334
R9856 DVDD.n1164 DVDD.n355 0.00334
R9857 DVDD.n356 DVDD.n355 0.00334
R9858 DVDD.n357 DVDD.n356 0.00334
R9859 DVDD.n362 DVDD.n361 0.00334
R9860 DVDD.n363 DVDD.n362 0.00334
R9861 DVDD.n366 DVDD.n363 0.00334
R9862 DVDD.n367 DVDD.n366 0.00334
R9863 DVDD.n368 DVDD.n367 0.00334
R9864 DVDD.n369 DVDD.n368 0.00334
R9865 DVDD.n372 DVDD.n369 0.00334
R9866 DVDD.n373 DVDD.n372 0.00334
R9867 DVDD.n374 DVDD.n373 0.00334
R9868 DVDD.n375 DVDD.n374 0.00334
R9869 DVDD.n383 DVDD.n375 0.00334
R9870 DVDD.n384 DVDD.n383 0.00334
R9871 DVDD.n385 DVDD.n384 0.00334
R9872 DVDD.n386 DVDD.n385 0.00334
R9873 DVDD.n389 DVDD.n386 0.00334
R9874 DVDD.n390 DVDD.n389 0.00334
R9875 DVDD.n391 DVDD.n390 0.00334
R9876 DVDD.n392 DVDD.n391 0.00334
R9877 DVDD.n395 DVDD.n392 0.00334
R9878 DVDD.n396 DVDD.n395 0.00334
R9879 DVDD.n397 DVDD.n396 0.00334
R9880 DVDD.n398 DVDD.n397 0.00334
R9881 DVDD.n698 DVDD.n398 0.00334
R9882 DVDD.n409 DVDD.n408 0.00334
R9883 DVDD.n410 DVDD.n409 0.00334
R9884 DVDD.n413 DVDD.n410 0.00334
R9885 DVDD.n414 DVDD.n413 0.00334
R9886 DVDD.n415 DVDD.n414 0.00334
R9887 DVDD.n416 DVDD.n415 0.00334
R9888 DVDD.n419 DVDD.n416 0.00334
R9889 DVDD.n420 DVDD.n419 0.00334
R9890 DVDD.n421 DVDD.n420 0.00334
R9891 DVDD.n422 DVDD.n421 0.00334
R9892 DVDD.n431 DVDD.n422 0.00334
R9893 DVDD.n432 DVDD.n431 0.00334
R9894 DVDD.n433 DVDD.n432 0.00334
R9895 DVDD.n434 DVDD.n433 0.00334
R9896 DVDD.n435 DVDD.n434 0.00334
R9897 DVDD.n438 DVDD.n435 0.00334
R9898 DVDD.n439 DVDD.n438 0.00334
R9899 DVDD.n440 DVDD.n439 0.00334
R9900 DVDD.n441 DVDD.n440 0.00334
R9901 DVDD.n444 DVDD.n441 0.00334
R9902 DVDD.n445 DVDD.n444 0.00334
R9903 DVDD.n446 DVDD.n445 0.00334
R9904 DVDD.n447 DVDD.n446 0.00334
R9905 DVDD.n5108 DVDD.n5107 0.00334
R9906 DVDD.n5109 DVDD.n5108 0.00334
R9907 DVDD.n5110 DVDD.n5109 0.00334
R9908 DVDD.n5113 DVDD.n5110 0.00334
R9909 DVDD.n5114 DVDD.n5113 0.00334
R9910 DVDD.n5115 DVDD.n5114 0.00334
R9911 DVDD.n5116 DVDD.n5115 0.00334
R9912 DVDD.n5118 DVDD.n5116 0.00334
R9913 DVDD.n5119 DVDD.n5118 0.00334
R9914 DVDD.n5119 DVDD.n132 0.00334
R9915 DVDD.n5852 DVDD.n132 0.00334
R9916 DVDD.n5853 DVDD.n5852 0.00334
R9917 DVDD.n5854 DVDD.n5853 0.00334
R9918 DVDD.n5854 DVDD.n128 0.00334
R9919 DVDD.n5860 DVDD.n128 0.00334
R9920 DVDD.n5861 DVDD.n5860 0.00334
R9921 DVDD.n5862 DVDD.n5861 0.00334
R9922 DVDD.n5862 DVDD.n124 0.00334
R9923 DVDD.n5868 DVDD.n124 0.00334
R9924 DVDD.n5869 DVDD.n5868 0.00334
R9925 DVDD.n5870 DVDD.n5869 0.00334
R9926 DVDD.n5870 DVDD.n120 0.00334
R9927 DVDD.n5876 DVDD.n120 0.00334
R9928 DVDD.n5878 DVDD.n118 0.00334
R9929 DVDD.n5883 DVDD.n118 0.00334
R9930 DVDD.n5884 DVDD.n5883 0.00334
R9931 DVDD.n5885 DVDD.n5884 0.00334
R9932 DVDD.n5886 DVDD.n5885 0.00334
R9933 DVDD.n5887 DVDD.n5886 0.00334
R9934 DVDD.n5890 DVDD.n5887 0.00334
R9935 DVDD.n5891 DVDD.n5890 0.00334
R9936 DVDD.n5892 DVDD.n5891 0.00334
R9937 DVDD.n5893 DVDD.n5892 0.00334
R9938 DVDD.n4417 DVDD.n1106 0.00334
R9939 DVDD.n4418 DVDD.n4417 0.00334
R9940 DVDD.n4419 DVDD.n4418 0.00334
R9941 DVDD.n4419 DVDD.n1102 0.00334
R9942 DVDD.n4425 DVDD.n1102 0.00334
R9943 DVDD.n4426 DVDD.n4425 0.00334
R9944 DVDD.n4427 DVDD.n4426 0.00334
R9945 DVDD.n4427 DVDD.n1098 0.00334
R9946 DVDD.n4433 DVDD.n1098 0.00334
R9947 DVDD.n4434 DVDD.n4433 0.00334
R9948 DVDD.n4435 DVDD.n4434 0.00334
R9949 DVDD.n4435 DVDD.n1096 0.00334
R9950 DVDD.n4439 DVDD.n1096 0.00334
R9951 DVDD.n4446 DVDD.n4441 0.00334
R9952 DVDD.n4447 DVDD.n4446 0.00334
R9953 DVDD.n4448 DVDD.n4447 0.00334
R9954 DVDD.n4448 DVDD.n1090 0.00334
R9955 DVDD.n4454 DVDD.n1090 0.00334
R9956 DVDD.n4455 DVDD.n4454 0.00334
R9957 DVDD.n4456 DVDD.n4455 0.00334
R9958 DVDD.n4456 DVDD.n1086 0.00334
R9959 DVDD.n4462 DVDD.n1086 0.00334
R9960 DVDD.n4463 DVDD.n4462 0.00334
R9961 DVDD.n4464 DVDD.n4463 0.00334
R9962 DVDD.n4465 DVDD.n4464 0.00334
R9963 DVDD.n4468 DVDD.n4465 0.00334
R9964 DVDD.n4469 DVDD.n4468 0.00334
R9965 DVDD.n4470 DVDD.n4469 0.00334
R9966 DVDD.n4471 DVDD.n4470 0.00334
R9967 DVDD.n4474 DVDD.n4471 0.00334
R9968 DVDD.n4475 DVDD.n4474 0.00334
R9969 DVDD.n4476 DVDD.n4475 0.00334
R9970 DVDD.n4477 DVDD.n4476 0.00334
R9971 DVDD.n4478 DVDD.n4477 0.00334
R9972 DVDD.n4478 DVDD.n700 0.00334
R9973 DVDD.n4882 DVDD.n700 0.00334
R9974 DVDD.n4884 DVDD.n693 0.00334
R9975 DVDD.n4890 DVDD.n693 0.00334
R9976 DVDD.n4891 DVDD.n4890 0.00334
R9977 DVDD.n4892 DVDD.n4891 0.00334
R9978 DVDD.n4892 DVDD.n689 0.00334
R9979 DVDD.n4898 DVDD.n689 0.00334
R9980 DVDD.n4899 DVDD.n4898 0.00334
R9981 DVDD.n4900 DVDD.n4899 0.00334
R9982 DVDD.n4900 DVDD.n685 0.00334
R9983 DVDD.n4906 DVDD.n685 0.00334
R9984 DVDD.n4907 DVDD.n4906 0.00334
R9985 DVDD.n4908 DVDD.n4907 0.00334
R9986 DVDD.n4909 DVDD.n4908 0.00334
R9987 DVDD.n4912 DVDD.n4909 0.00334
R9988 DVDD.n4913 DVDD.n4912 0.00334
R9989 DVDD.n4914 DVDD.n4913 0.00334
R9990 DVDD.n4915 DVDD.n4914 0.00334
R9991 DVDD.n4918 DVDD.n4915 0.00334
R9992 DVDD.n4919 DVDD.n4918 0.00334
R9993 DVDD.n4920 DVDD.n4919 0.00334
R9994 DVDD.n4921 DVDD.n4920 0.00334
R9995 DVDD.n4921 DVDD.n479 0.00334
R9996 DVDD.n5248 DVDD.n479 0.00334
R9997 DVDD.n5251 DVDD.n5250 0.00334
R9998 DVDD.n5252 DVDD.n5251 0.00334
R9999 DVDD.n5253 DVDD.n5252 0.00334
R10000 DVDD.n5256 DVDD.n5253 0.00334
R10001 DVDD.n5257 DVDD.n5256 0.00334
R10002 DVDD.n5258 DVDD.n5257 0.00334
R10003 DVDD.n5259 DVDD.n5258 0.00334
R10004 DVDD.n5262 DVDD.n5259 0.00334
R10005 DVDD.n5263 DVDD.n5262 0.00334
R10006 DVDD.n5264 DVDD.n5263 0.00334
R10007 DVDD.n5265 DVDD.n5264 0.00334
R10008 DVDD.n5266 DVDD.n5265 0.00334
R10009 DVDD.n5267 DVDD.n5266 0.00334
R10010 DVDD.n5268 DVDD.n5267 0.00334
R10011 DVDD.n5271 DVDD.n5268 0.00334
R10012 DVDD.n5272 DVDD.n5271 0.00334
R10013 DVDD.n5273 DVDD.n5272 0.00334
R10014 DVDD.n5274 DVDD.n5273 0.00334
R10015 DVDD.n5277 DVDD.n5274 0.00334
R10016 DVDD.n5278 DVDD.n5277 0.00334
R10017 DVDD.n5279 DVDD.n5278 0.00334
R10018 DVDD.n5280 DVDD.n5279 0.00334
R10019 DVDD.n5281 DVDD.n5280 0.00334
R10020 DVDD.n46 DVDD.n45 0.00334
R10021 DVDD.n5577 DVDD.n46 0.00334
R10022 DVDD.n5578 DVDD.n5577 0.00334
R10023 DVDD.n5579 DVDD.n5578 0.00334
R10024 DVDD.n5580 DVDD.n5579 0.00334
R10025 DVDD.n5581 DVDD.n5580 0.00334
R10026 DVDD.n5584 DVDD.n5581 0.00334
R10027 DVDD.n5585 DVDD.n5584 0.00334
R10028 DVDD.n5586 DVDD.n5585 0.00334
R10029 DVDD.n5587 DVDD.n5586 0.00334
R10030 DVDD.n4347 DVDD.n4346 0.00334
R10031 DVDD.n4348 DVDD.n4347 0.00334
R10032 DVDD.n4351 DVDD.n4348 0.00334
R10033 DVDD.n4352 DVDD.n4351 0.00334
R10034 DVDD.n4353 DVDD.n4352 0.00334
R10035 DVDD.n4354 DVDD.n4353 0.00334
R10036 DVDD.n4356 DVDD.n4354 0.00334
R10037 DVDD.n4358 DVDD.n4356 0.00334
R10038 DVDD.n4358 DVDD.n4357 0.00334
R10039 DVDD.n4357 DVDD.n986 0.00334
R10040 DVDD.n987 DVDD.n986 0.00334
R10041 DVDD.n988 DVDD.n987 0.00334
R10042 DVDD.n989 DVDD.n988 0.00334
R10043 DVDD.n994 DVDD.n991 0.00334
R10044 DVDD.n995 DVDD.n994 0.00334
R10045 DVDD.n996 DVDD.n995 0.00334
R10046 DVDD.n997 DVDD.n996 0.00334
R10047 DVDD.n1000 DVDD.n997 0.00334
R10048 DVDD.n1001 DVDD.n1000 0.00334
R10049 DVDD.n1002 DVDD.n1001 0.00334
R10050 DVDD.n1003 DVDD.n1002 0.00334
R10051 DVDD.n1006 DVDD.n1003 0.00334
R10052 DVDD.n1007 DVDD.n1006 0.00334
R10053 DVDD.n1008 DVDD.n1007 0.00334
R10054 DVDD.n1021 DVDD.n1008 0.00334
R10055 DVDD.n1022 DVDD.n1021 0.00334
R10056 DVDD.n1023 DVDD.n1022 0.00334
R10057 DVDD.n1024 DVDD.n1023 0.00334
R10058 DVDD.n1027 DVDD.n1024 0.00334
R10059 DVDD.n1028 DVDD.n1027 0.00334
R10060 DVDD.n1029 DVDD.n1028 0.00334
R10061 DVDD.n1030 DVDD.n1029 0.00334
R10062 DVDD.n1032 DVDD.n1030 0.00334
R10063 DVDD.n1032 DVDD.n1031 0.00334
R10064 DVDD.n1031 DVDD.n730 0.00334
R10065 DVDD.n731 DVDD.n730 0.00334
R10066 DVDD.n4804 DVDD.n4803 0.00334
R10067 DVDD.n4807 DVDD.n4804 0.00334
R10068 DVDD.n4808 DVDD.n4807 0.00334
R10069 DVDD.n4809 DVDD.n4808 0.00334
R10070 DVDD.n4810 DVDD.n4809 0.00334
R10071 DVDD.n4813 DVDD.n4810 0.00334
R10072 DVDD.n4814 DVDD.n4813 0.00334
R10073 DVDD.n4815 DVDD.n4814 0.00334
R10074 DVDD.n4816 DVDD.n4815 0.00334
R10075 DVDD.n4817 DVDD.n4816 0.00334
R10076 DVDD.n4818 DVDD.n4817 0.00334
R10077 DVDD.n4819 DVDD.n4818 0.00334
R10078 DVDD.n4820 DVDD.n4819 0.00334
R10079 DVDD.n4823 DVDD.n4820 0.00334
R10080 DVDD.n4824 DVDD.n4823 0.00334
R10081 DVDD.n4825 DVDD.n4824 0.00334
R10082 DVDD.n4826 DVDD.n4825 0.00334
R10083 DVDD.n4829 DVDD.n4826 0.00334
R10084 DVDD.n4830 DVDD.n4829 0.00334
R10085 DVDD.n4831 DVDD.n4830 0.00334
R10086 DVDD.n4832 DVDD.n4831 0.00334
R10087 DVDD.n4834 DVDD.n4832 0.00334
R10088 DVDD.n4834 DVDD.n4833 0.00334
R10089 DVDD.n497 DVDD.n483 0.00334
R10090 DVDD.n498 DVDD.n497 0.00334
R10091 DVDD.n499 DVDD.n498 0.00334
R10092 DVDD.n500 DVDD.n499 0.00334
R10093 DVDD.n503 DVDD.n500 0.00334
R10094 DVDD.n504 DVDD.n503 0.00334
R10095 DVDD.n505 DVDD.n504 0.00334
R10096 DVDD.n506 DVDD.n505 0.00334
R10097 DVDD.n508 DVDD.n506 0.00334
R10098 DVDD.n509 DVDD.n508 0.00334
R10099 DVDD.n510 DVDD.n509 0.00334
R10100 DVDD.n511 DVDD.n510 0.00334
R10101 DVDD.n512 DVDD.n511 0.00334
R10102 DVDD.n515 DVDD.n512 0.00334
R10103 DVDD.n516 DVDD.n515 0.00334
R10104 DVDD.n517 DVDD.n516 0.00334
R10105 DVDD.n518 DVDD.n517 0.00334
R10106 DVDD.n521 DVDD.n518 0.00334
R10107 DVDD.n522 DVDD.n521 0.00334
R10108 DVDD.n523 DVDD.n522 0.00334
R10109 DVDD.n524 DVDD.n523 0.00334
R10110 DVDD.n524 DVDD.n36 0.00334
R10111 DVDD.n5941 DVDD.n36 0.00334
R10112 DVDD.n5944 DVDD.n5943 0.00334
R10113 DVDD.n5945 DVDD.n5944 0.00334
R10114 DVDD.n5946 DVDD.n5945 0.00334
R10115 DVDD.n5946 DVDD.n5 0.00334
R10116 DVDD.n5958 DVDD.n5 0.00334
R10117 DVDD.n5959 DVDD.n5958 0.00334
R10118 DVDD.n5961 DVDD.n5959 0.00334
R10119 DVDD.n5961 DVDD.n5960 0.00334
R10120 DVDD.n5960 DVDD.n1 0.00334
R10121 DVDD.n5968 DVDD.n1 0.00334
R10122 DVDD.n5969 DVDD.n5968 0.00334
R10123 DVDD.n4302 DVDD.n4301 0.00334
R10124 DVDD.n4303 DVDD.n4302 0.00334
R10125 DVDD.n4306 DVDD.n4303 0.00334
R10126 DVDD.n4307 DVDD.n4306 0.00334
R10127 DVDD.n4308 DVDD.n4307 0.00334
R10128 DVDD.n4309 DVDD.n4308 0.00334
R10129 DVDD.n4312 DVDD.n4309 0.00334
R10130 DVDD.n4313 DVDD.n4312 0.00334
R10131 DVDD.n4314 DVDD.n4313 0.00334
R10132 DVDD.n4314 DVDD.n912 0.00334
R10133 DVDD.n4713 DVDD.n912 0.00334
R10134 DVDD.n4714 DVDD.n4713 0.00334
R10135 DVDD.n4715 DVDD.n4714 0.00334
R10136 DVDD.n4722 DVDD.n4721 0.00334
R10137 DVDD.n4723 DVDD.n4722 0.00334
R10138 DVDD.n4723 DVDD.n903 0.00334
R10139 DVDD.n4729 DVDD.n903 0.00334
R10140 DVDD.n4730 DVDD.n4729 0.00334
R10141 DVDD.n4731 DVDD.n4730 0.00334
R10142 DVDD.n4731 DVDD.n899 0.00334
R10143 DVDD.n4737 DVDD.n899 0.00334
R10144 DVDD.n4738 DVDD.n4737 0.00334
R10145 DVDD.n4739 DVDD.n4738 0.00334
R10146 DVDD.n4739 DVDD.n889 0.00334
R10147 DVDD.n4747 DVDD.n889 0.00334
R10148 DVDD.n4748 DVDD.n4747 0.00334
R10149 DVDD.n4749 DVDD.n4748 0.00334
R10150 DVDD.n4749 DVDD.n885 0.00334
R10151 DVDD.n4755 DVDD.n885 0.00334
R10152 DVDD.n4756 DVDD.n4755 0.00334
R10153 DVDD.n4757 DVDD.n4756 0.00334
R10154 DVDD.n4757 DVDD.n881 0.00334
R10155 DVDD.n4763 DVDD.n881 0.00334
R10156 DVDD.n4764 DVDD.n4763 0.00334
R10157 DVDD.n4767 DVDD.n4764 0.00334
R10158 DVDD.n4767 DVDD.n4766 0.00334
R10159 DVDD.n4775 DVDD.n733 0.00334
R10160 DVDD.n4776 DVDD.n4775 0.00334
R10161 DVDD.n4777 DVDD.n4776 0.00334
R10162 DVDD.n4778 DVDD.n4777 0.00334
R10163 DVDD.n4781 DVDD.n4778 0.00334
R10164 DVDD.n4782 DVDD.n4781 0.00334
R10165 DVDD.n4783 DVDD.n4782 0.00334
R10166 DVDD.n4784 DVDD.n4783 0.00334
R10167 DVDD.n4785 DVDD.n4784 0.00334
R10168 DVDD.n4785 DVDD.n586 0.00334
R10169 DVDD.n5023 DVDD.n586 0.00334
R10170 DVDD.n5024 DVDD.n5023 0.00334
R10171 DVDD.n5025 DVDD.n5024 0.00334
R10172 DVDD.n5025 DVDD.n582 0.00334
R10173 DVDD.n5031 DVDD.n582 0.00334
R10174 DVDD.n5032 DVDD.n5031 0.00334
R10175 DVDD.n5033 DVDD.n5032 0.00334
R10176 DVDD.n5033 DVDD.n578 0.00334
R10177 DVDD.n5039 DVDD.n578 0.00334
R10178 DVDD.n5040 DVDD.n5039 0.00334
R10179 DVDD.n5041 DVDD.n5040 0.00334
R10180 DVDD.n5041 DVDD.n574 0.00334
R10181 DVDD.n5047 DVDD.n574 0.00334
R10182 DVDD.n5050 DVDD.n5049 0.00334
R10183 DVDD.n5053 DVDD.n5050 0.00334
R10184 DVDD.n5054 DVDD.n5053 0.00334
R10185 DVDD.n5055 DVDD.n5054 0.00334
R10186 DVDD.n5056 DVDD.n5055 0.00334
R10187 DVDD.n5059 DVDD.n5056 0.00334
R10188 DVDD.n5060 DVDD.n5059 0.00334
R10189 DVDD.n5061 DVDD.n5060 0.00334
R10190 DVDD.n5062 DVDD.n5061 0.00334
R10191 DVDD.n5064 DVDD.n5062 0.00334
R10192 DVDD.n5066 DVDD.n5064 0.00334
R10193 DVDD.n5066 DVDD.n5065 0.00334
R10194 DVDD.n5065 DVDD.n201 0.00334
R10195 DVDD.n202 DVDD.n201 0.00334
R10196 DVDD.n203 DVDD.n202 0.00334
R10197 DVDD.n206 DVDD.n203 0.00334
R10198 DVDD.n207 DVDD.n206 0.00334
R10199 DVDD.n208 DVDD.n207 0.00334
R10200 DVDD.n209 DVDD.n208 0.00334
R10201 DVDD.n212 DVDD.n209 0.00334
R10202 DVDD.n213 DVDD.n212 0.00334
R10203 DVDD.n214 DVDD.n213 0.00334
R10204 DVDD.n215 DVDD.n214 0.00334
R10205 DVDD.n5673 DVDD.n216 0.00334
R10206 DVDD.n5674 DVDD.n5673 0.00334
R10207 DVDD.n5675 DVDD.n5674 0.00334
R10208 DVDD.n5676 DVDD.n5675 0.00334
R10209 DVDD.n5677 DVDD.n5676 0.00334
R10210 DVDD.n5680 DVDD.n5677 0.00334
R10211 DVDD.n5681 DVDD.n5680 0.00334
R10212 DVDD.n5682 DVDD.n5681 0.00334
R10213 DVDD.n5683 DVDD.n5682 0.00334
R10214 DVDD.n5685 DVDD.n5683 0.00334
R10215 DVDD.n5686 DVDD.n5685 0.00334
R10216 DVDD.n3621 DVDD.n3620 0.00334
R10217 DVDD.n3622 DVDD.n3621 0.00334
R10218 DVDD.n3622 DVDD.n2018 0.00334
R10219 DVDD.n3631 DVDD.n2018 0.00334
R10220 DVDD.n3634 DVDD.n3632 0.00334
R10221 DVDD.n3634 DVDD.n3633 0.00334
R10222 DVDD.n3633 DVDD.n2005 0.00334
R10223 DVDD.n3646 DVDD.n2005 0.00334
R10224 DVDD.n3670 DVDD.n1977 0.00334
R10225 DVDD.n3671 DVDD.n3670 0.00334
R10226 DVDD.n3672 DVDD.n3671 0.00334
R10227 DVDD.n3672 DVDD.n1973 0.00334
R10228 DVDD.n3679 DVDD.n3678 0.00334
R10229 DVDD.n3680 DVDD.n3679 0.00334
R10230 DVDD.n3680 DVDD.n1969 0.00334
R10231 DVDD.n3686 DVDD.n1969 0.00334
R10232 DVDD.n3703 DVDD.n3687 0.00334
R10233 DVDD.n3255 DVDD.n3254 0.00334
R10234 DVDD.n3254 DVDD.n3253 0.00334
R10235 DVDD.n3218 DVDD.n3217 0.00334
R10236 DVDD.n3402 DVDD.n3217 0.00334
R10237 DVDD.n3403 DVDD.n3402 0.00334
R10238 DVDD.n3404 DVDD.n3403 0.00334
R10239 DVDD.n3422 DVDD.n3213 0.00334
R10240 DVDD.n3423 DVDD.n3422 0.00334
R10241 DVDD.n3424 DVDD.n3423 0.00334
R10242 DVDD.n3424 DVDD.n2004 0.00334
R10243 DVDD.n3202 DVDD.n2003 0.00334
R10244 DVDD.n3449 DVDD.n3202 0.00334
R10245 DVDD.n3450 DVDD.n3449 0.00334
R10246 DVDD.n3461 DVDD.n3450 0.00334
R10247 DVDD.n3460 DVDD.n3459 0.00334
R10248 DVDD.n3459 DVDD.n3451 0.00334
R10249 DVDD.n3455 DVDD.n3451 0.00334
R10250 DVDD.n3455 DVDD.n1966 0.00334
R10251 DVDD.n1965 DVDD.n1947 0.00334
R10252 DVDD.n3304 DVDD.n3303 0.00334
R10253 DVDD.n3305 DVDD.n3304 0.00334
R10254 DVDD.n3101 DVDD.n3100 0.00334
R10255 DVDD.n3104 DVDD.n3101 0.00334
R10256 DVDD.n3105 DVDD.n3104 0.00334
R10257 DVDD.n3106 DVDD.n3105 0.00334
R10258 DVDD.n3115 DVDD.n3107 0.00334
R10259 DVDD.n3116 DVDD.n3115 0.00334
R10260 DVDD.n3117 DVDD.n3116 0.00334
R10261 DVDD.n3117 DVDD.n2000 0.00334
R10262 DVDD.n3130 DVDD.n1999 0.00334
R10263 DVDD.n3131 DVDD.n3130 0.00334
R10264 DVDD.n3145 DVDD.n3131 0.00334
R10265 DVDD.n3146 DVDD.n3145 0.00334
R10266 DVDD.n3148 DVDD.n3147 0.00334
R10267 DVDD.n3563 DVDD.n3148 0.00334
R10268 DVDD.n3564 DVDD.n3563 0.00334
R10269 DVDD.n3564 DVDD.n1944 0.00334
R10270 DVDD.n1943 DVDD.n1905 0.00334
R10271 DVDD.n2054 DVDD.n2053 0.00334
R10272 DVDD.n2055 DVDD.n2054 0.00334
R10273 DVDD.n3084 DVDD.n3083 0.00334
R10274 DVDD.n3083 DVDD.n3082 0.00334
R10275 DVDD.n3082 DVDD.n2029 0.00334
R10276 DVDD.n3078 DVDD.n2029 0.00334
R10277 DVDD.n3077 DVDD.n3076 0.00334
R10278 DVDD.n3076 DVDD.n2034 0.00334
R10279 DVDD.n3072 DVDD.n2034 0.00334
R10280 DVDD.n3072 DVDD.n2001 0.00334
R10281 DVDD.n3046 DVDD.n2002 0.00334
R10282 DVDD.n3047 DVDD.n3046 0.00334
R10283 DVDD.n3049 DVDD.n3047 0.00334
R10284 DVDD.n3049 DVDD.n3048 0.00334
R10285 DVDD.n3058 DVDD.n3032 0.00334
R10286 DVDD.n3059 DVDD.n3058 0.00334
R10287 DVDD.n3060 DVDD.n3059 0.00334
R10288 DVDD.n3060 DVDD.n1902 0.00334
R10289 DVDD.n1926 DVDD.n1901 0.00334
R10290 DVDD.n3731 DVDD.n1854 0.00334
R10291 DVDD.n3782 DVDD.n1854 0.00334
R10292 DVDD.n3783 DVDD.n3782 0.00334
R10293 DVDD.n3784 DVDD.n3783 0.00334
R10294 DVDD.n3784 DVDD.n1850 0.00334
R10295 DVDD.n3790 DVDD.n1850 0.00334
R10296 DVDD.n3791 DVDD.n3790 0.00334
R10297 DVDD.n3792 DVDD.n3791 0.00334
R10298 DVDD.n3792 DVDD.n1846 0.00334
R10299 DVDD.n3799 DVDD.n1846 0.00334
R10300 DVDD.n3800 DVDD.n3799 0.00334
R10301 DVDD.n3801 DVDD.n3800 0.00334
R10302 DVDD.n3801 DVDD.n1687 0.00334
R10303 DVDD.n4257 DVDD.n1688 0.00334
R10304 DVDD.n1692 DVDD.n1688 0.00334
R10305 DVDD.n1693 DVDD.n1692 0.00334
R10306 DVDD.n1696 DVDD.n1693 0.00334
R10307 DVDD.n1697 DVDD.n1696 0.00334
R10308 DVDD.n1698 DVDD.n1697 0.00334
R10309 DVDD.n1701 DVDD.n1698 0.00334
R10310 DVDD.n1702 DVDD.n1701 0.00334
R10311 DVDD.n1703 DVDD.n1702 0.00334
R10312 DVDD.n1704 DVDD.n1703 0.00334
R10313 DVDD.n3936 DVDD.n1704 0.00334
R10314 DVDD.n3937 DVDD.n3936 0.00334
R10315 DVDD.n3938 DVDD.n3937 0.00334
R10316 DVDD.n3939 DVDD.n3938 0.00334
R10317 DVDD.n3940 DVDD.n3939 0.00334
R10318 DVDD.n3943 DVDD.n3940 0.00334
R10319 DVDD.n3944 DVDD.n3943 0.00334
R10320 DVDD.n3945 DVDD.n3944 0.00334
R10321 DVDD.n3946 DVDD.n3945 0.00334
R10322 DVDD.n3946 DVDD.n3925 0.00334
R10323 DVDD.n3970 DVDD.n3925 0.00334
R10324 DVDD.n3971 DVDD.n3970 0.00334
R10325 DVDD.n3972 DVDD.n3971 0.00334
R10326 DVDD.n3979 DVDD.n3978 0.00334
R10327 DVDD.n3980 DVDD.n3979 0.00334
R10328 DVDD.n3980 DVDD.n1813 0.00334
R10329 DVDD.n3986 DVDD.n1813 0.00334
R10330 DVDD.n3987 DVDD.n3986 0.00334
R10331 DVDD.n3988 DVDD.n3987 0.00334
R10332 DVDD.n3988 DVDD.n1809 0.00334
R10333 DVDD.n3998 DVDD.n1809 0.00334
R10334 DVDD.n3999 DVDD.n3998 0.00334
R10335 DVDD.n4000 DVDD.n3999 0.00334
R10336 DVDD.n4000 DVDD.n1805 0.00334
R10337 DVDD.n4006 DVDD.n1805 0.00334
R10338 DVDD.n4007 DVDD.n4006 0.00334
R10339 DVDD.n4008 DVDD.n4007 0.00334
R10340 DVDD.n4008 DVDD.n1801 0.00334
R10341 DVDD.n4018 DVDD.n1801 0.00334
R10342 DVDD.n4019 DVDD.n4018 0.00334
R10343 DVDD.n4020 DVDD.n4019 0.00334
R10344 DVDD.n4020 DVDD.n1797 0.00334
R10345 DVDD.n4027 DVDD.n1797 0.00334
R10346 DVDD.n4028 DVDD.n4027 0.00334
R10347 DVDD.n4029 DVDD.n4028 0.00334
R10348 DVDD.n4029 DVDD.n1789 0.00334
R10349 DVDD.n4104 DVDD.n4103 0.00334
R10350 DVDD.n4105 DVDD.n4104 0.00334
R10351 DVDD.n4106 DVDD.n4105 0.00334
R10352 DVDD.n4108 DVDD.n4106 0.00334
R10353 DVDD.n4109 DVDD.n4108 0.00334
R10354 DVDD.n4109 DVDD.n1782 0.00334
R10355 DVDD.n4130 DVDD.n1782 0.00334
R10356 DVDD.n4131 DVDD.n4130 0.00334
R10357 DVDD.n4132 DVDD.n4131 0.00334
R10358 DVDD.n4132 DVDD.n1778 0.00334
R10359 DVDD.n4142 DVDD.n1778 0.00334
R10360 DVDD.n4143 DVDD.n4142 0.00334
R10361 DVDD.n4144 DVDD.n4143 0.00334
R10362 DVDD.n4144 DVDD.n1775 0.00334
R10363 DVDD.n4152 DVDD.n1775 0.00334
R10364 DVDD.n4153 DVDD.n4152 0.00334
R10365 DVDD.n4154 DVDD.n4153 0.00334
R10366 DVDD.n4154 DVDD.n1771 0.00334
R10367 DVDD.n4162 DVDD.n1771 0.00334
R10368 DVDD.n4163 DVDD.n4162 0.00334
R10369 DVDD.n4164 DVDD.n4163 0.00334
R10370 DVDD.n4164 DVDD.n1767 0.00334
R10371 DVDD.n4170 DVDD.n1767 0.00334
R10372 DVDD.n4220 DVDD.n4171 0.00334
R10373 DVDD.n4177 DVDD.n4171 0.00334
R10374 DVDD.n4178 DVDD.n4177 0.00334
R10375 DVDD.n4179 DVDD.n4178 0.00334
R10376 DVDD.n4182 DVDD.n4179 0.00334
R10377 DVDD.n4183 DVDD.n4182 0.00334
R10378 DVDD.n4184 DVDD.n4183 0.00334
R10379 DVDD.n4185 DVDD.n4184 0.00334
R10380 DVDD.n4191 DVDD.n4185 0.00334
R10381 DVDD.n4192 DVDD.n4191 0.00334
R10382 DVDD.n4196 DVDD.n4192 0.00334
R10383 DVDD.n4720 DVDD.n908 0.00332
R10384 DVDD.n4635 DVDD.n4634 0.00332
R10385 DVDD.n4442 DVDD.n990 0.00332
R10386 DVDD.n5397 DVDD.n358 0.00332
R10387 DVDD.n4256 DVDD.n1685 0.00332
R10388 DVDD.n5399 DVDD.n5398 0.00332
R10389 DVDD.n4443 DVDD.n359 0.00332
R10390 DVDD.n4633 DVDD.n909 0.00332
R10391 DVDD.n4719 DVDD.n4718 0.00332
R10392 DVDD.n5402 DVDD.n322 0.00329
R10393 DVDD.n295 DVDD.n284 0.00329
R10394 DVDD.n5472 DVDD.n297 0.00329
R10395 DVDD.n4640 DVDD.n974 0.00329
R10396 DVDD.n4638 DVDD.n972 0.00329
R10397 DVDD.n921 DVDD.n910 0.00329
R10398 DVDD.n5627 DVDD.n5605 0.0032883
R10399 DVDD.n5452 DVDD.n289 0.0032883
R10400 DVDD.n4255 DVDD.n1690 0.00323
R10401 DVDD.n4114 DVDD.n4113 0.00323
R10402 DVDD.n5920 DVDD.n82 0.00323
R10403 DVDD.n5933 DVDD.n43 0.00323
R10404 DVDD.n5932 DVDD.n58 0.00323
R10405 DVDD.n5952 DVDD.n5951 0.00323
R10406 DVDD.n5948 DVDD.n29 0.00323
R10407 DVDD.n5707 DVDD.n220 0.00323
R10408 DVDD.n3898 DVDD.n3869 0.0032
R10409 DVDD.n3900 DVDD.n3899 0.0032
R10410 DVDD.n4260 DVDD.n1685 0.0032
R10411 DVDD.n3694 DVDD.n3690 0.00314706
R10412 DVDD.n4272 DVDD.n1675 0.00314375
R10413 DVDD.n1680 DVDD.n1679 0.00314375
R10414 DVDD.n4266 DVDD.n4265 0.00314375
R10415 DVDD.n4262 DVDD.n1681 0.00314375
R10416 DVDD.n4261 DVDD.n1684 0.00314375
R10417 DVDD.n3806 DVDD.n1843 0.00314375
R10418 DVDD.n3812 DVDD.n3810 0.00314375
R10419 DVDD.n3811 DVDD.n1840 0.00314375
R10420 DVDD.n3817 DVDD.n3816 0.00314375
R10421 DVDD.n1841 DVDD.n1836 0.00314375
R10422 DVDD.n2276 DVDD.n2269 0.00313571
R10423 DVDD.n2294 DVDD.n2264 0.00313571
R10424 DVDD.n3966 DVDD.n3965 0.00311
R10425 DVDD.n4329 DVDD.n4300 0.00309529
R10426 DVDD.n4372 DVDD.n4345 0.00309529
R10427 DVDD.n4409 DVDD.n4399 0.00309529
R10428 DVDD.n1180 DVDD.n1150 0.00309529
R10429 DVDD.n2045 DVDD.n2044 0.00309529
R10430 DVDD.n3301 DVDD.n3273 0.00309529
R10431 DVDD.n3250 DVDD.n3247 0.00309529
R10432 DVDD.n3733 DVDD.n3721 0.00309529
R10433 DVDD.n5796 DVDD.n156 0.00308197
R10434 DVDD.n5152 DVDD.n464 0.00308197
R10435 DVDD.n4986 DVDD.n4940 0.00308197
R10436 DVDD.n755 DVDD.n753 0.00308197
R10437 DVDD.n4542 DVDD.n4499 0.00308197
R10438 DVDD.n5881 DVDD.n77 0.00302
R10439 DVDD.n116 DVDD.n79 0.00302
R10440 DVDD.n5563 DVDD.n58 0.00302
R10441 DVDD.n5649 DVDD.n5564 0.00302
R10442 DVDD.n5948 DVDD.n31 0.00302
R10443 DVDD.n5954 DVDD.n7 0.00302
R10444 DVDD.n5701 DVDD.n224 0.00302
R10445 DVDD.n5705 DVDD.n227 0.00302
R10446 DVDD.n2566 DVDD.n2565 0.00300714
R10447 DVDD.n1573 DVDD.n1197 0.00300714
R10448 DVDD.n1572 DVDD.n1192 0.00300714
R10449 DVDD.n5644 DVDD.n5567 0.00297849
R10450 DVDD.n5470 DVDD.n276 0.00297849
R10451 DVDD.n4052 DVDD.n4047 0.002975
R10452 DVDD.n4067 DVDD.n4066 0.002975
R10453 DVDD.n4063 DVDD.n4053 0.002975
R10454 DVDD.n4062 DVDD.n4055 0.002975
R10455 DVDD.n4057 DVDD.n4056 0.002975
R10456 DVDD.n4225 DVDD.n1721 0.002975
R10457 DVDD.n1764 DVDD.n1763 0.002975
R10458 DVDD.n1760 DVDD.n1729 0.002975
R10459 DVDD.n1759 DVDD.n1730 0.002975
R10460 DVDD.n5427 DVDD.n328 0.00296
R10461 DVDD.n5405 DVDD.n321 0.00296
R10462 DVDD.n273 DVDD.n271 0.00296
R10463 DVDD.n5475 DVDD.n284 0.00296
R10464 DVDD.n4698 DVDD.n4643 0.00296
R10465 DVDD.n4640 DVDD.n971 0.00296
R10466 DVDD.n4707 DVDD.n4706 0.00296
R10467 DVDD.n4711 DVDD.n914 0.00296
R10468 DVDD.n2856 DVDD.n2686 0.00294565
R10469 DVDD.n3779 DVDD.n1852 0.00287
R10470 DVDD.n5362 DVDD.n5361 0.00287
R10471 DVDD.n4480 DVDD.n702 0.00287
R10472 DVDD.n4875 DVDD.n4874 0.00287
R10473 DVDD.n4771 DVDD.n4769 0.00287
R10474 DVDD.n5878 DVDD.n5877 0.00286
R10475 DVDD.n45 DVDD.n35 0.00286
R10476 DVDD.n5943 DVDD.n5942 0.00286
R10477 DVDD.n216 DVDD.n34 0.00286
R10478 DVDD.n4221 DVDD.n4220 0.00286
R10479 DVDD.n5609 DVDD.n67 0.00282358
R10480 DVDD.n317 DVDD.n298 0.00282358
R10481 DVDD.n3638 DVDD.n3636 0.00281
R10482 DVDD.n5104 DVDD.n449 0.00281
R10483 DVDD.n5134 DVDD.n5133 0.00281
R10484 DVDD.n5318 DVDD.n462 0.00281
R10485 DVDD.n5316 DVDD.n5315 0.00281
R10486 DVDD.n5243 DVDD.n485 0.00281
R10487 DVDD.n5242 DVDD.n555 0.00281
R10488 DVDD.n5094 DVDD.n5085 0.00281
R10489 DVDD.n5082 DVDD.n570 0.00281
R10490 DVDD DVDD.n5893 0.00278
R10491 DVDD DVDD.n5587 0.00278
R10492 DVDD.n3652 DVDD.n1996 0.00275
R10493 DVDD.n3029 DVDD.n1896 0.00275
R10494 DVDD.n2056 DVDD.n2023 0.00275
R10495 DVDD.n3039 DVDD.n1998 0.00275
R10496 DVDD.n3031 DVDD.n1897 0.00275
R10497 DVDD.n3306 DVDD.n2023 0.00275
R10498 DVDD.n3129 DVDD.n1998 0.00275
R10499 DVDD.n3565 DVDD.n1897 0.00275
R10500 DVDD.n3652 DVDD.n1992 0.00275
R10501 DVDD.n3562 DVDD.n1896 0.00275
R10502 DVDD.n3652 DVDD.n1990 0.00275
R10503 DVDD.n3453 DVDD.n1896 0.00275
R10504 DVDD.n3252 DVDD.n2023 0.00275
R10505 DVDD.n3203 DVDD.n1998 0.00275
R10506 DVDD.n3454 DVDD.n1897 0.00275
R10507 DVDD.n1998 DVDD.n1978 0.00275
R10508 DVDD.n3685 DVDD.n1897 0.00275
R10509 DVDD.n3684 DVDD.n1896 0.00275
R10510 DVDD.n3835 DVDD.n1830 0.00275
R10511 DVDD.n3855 DVDD.n1818 0.00275
R10512 DVDD.n3834 DVDD.n3833 0.00275
R10513 DVDD.n3975 DVDD.n3856 0.00275
R10514 DVDD.n4204 DVDD.n4187 0.00275
R10515 DVDD.n5760 DVDD.n176 0.00271311
R10516 DVDD.n5223 DVDD.n562 0.00271311
R10517 DVDD.n644 DVDD.n612 0.00271311
R10518 DVDD.n849 DVDD.n722 0.00271311
R10519 DVDD.n4596 DVDD.n1053 0.00271311
R10520 DVDD.n3495 DVDD.n3177 0.00270109
R10521 DVDD.n3536 DVDD.n3153 0.00270109
R10522 DVDD.n5107 DVDD.n478 0.0027
R10523 DVDD.n5250 DVDD.n5249 0.0027
R10524 DVDD.n483 DVDD.n477 0.0027
R10525 DVDD.n5049 DVDD.n5048 0.0027
R10526 DVDD.n4103 DVDD.n4102 0.0027
R10527 DVDD.n3668 DVDD.n1979 0.00269
R10528 DVDD.n3958 DVDD.n3933 0.00269
R10529 DVDD.n4138 DVDD.n4135 0.00269
R10530 DVDD DVDD.n2022 0.00267716
R10531 DVDD.n3704 DVDD 0.00267716
R10532 DVDD.n5953 DVDD.n30 0.00266867
R10533 DVDD.n4699 DVDD.n973 0.00266867
R10534 DVDD.n4175 DVDD.n1722 0.00263
R10535 DVDD.n4079 DVDD.n4078 0.0026
R10536 DVDD.n3653 DVDD.n1979 0.00257
R10537 DVDD.n3958 DVDD.n3957 0.00257
R10538 DVDD.n4140 DVDD.n4138 0.00257
R10539 DVDD.n699 DVDD.n408 0.00254
R10540 DVDD.n4884 DVDD.n4883 0.00254
R10541 DVDD.n4803 DVDD.n697 0.00254
R10542 DVDD.n4765 DVDD.n733 0.00254
R10543 DVDD.n3978 DVDD.n1817 0.00254
R10544 DVDD.n5632 DVDD.n53 0.00251377
R10545 DVDD.n5457 DVDD.n313 0.00251377
R10546 DVDD.n3617 DVDD.n3086 0.00251
R10547 DVDD.n1928 DVDD.n1896 0.00251
R10548 DVDD.n3085 DVDD.n2023 0.00251
R10549 DVDD.n3071 DVDD.n1998 0.00251
R10550 DVDD.n1927 DVDD.n1897 0.00251
R10551 DVDD.n3615 DVDD.n2023 0.00251
R10552 DVDD.n3118 DVDD.n1998 0.00251
R10553 DVDD.n1942 DVDD.n1897 0.00251
R10554 DVDD.n3617 DVDD.n3616 0.00251
R10555 DVDD.n1941 DVDD.n1896 0.00251
R10556 DVDD.n3617 DVDD.n3095 0.00251
R10557 DVDD.n1948 DVDD.n1896 0.00251
R10558 DVDD.n3219 DVDD.n2023 0.00251
R10559 DVDD.n3426 DVDD.n1998 0.00251
R10560 DVDD.n1964 DVDD.n1897 0.00251
R10561 DVDD.n3619 DVDD.n2023 0.00251
R10562 DVDD.n3645 DVDD.n1998 0.00251
R10563 DVDD.n3702 DVDD.n1897 0.00251
R10564 DVDD.n3618 DVDD.n3617 0.00251
R10565 DVDD.n3652 DVDD.n1983 0.00251
R10566 DVDD.n3701 DVDD.n1896 0.00251
R10567 DVDD.n4205 DVDD.n4204 0.00251
R10568 DVDD.n3638 DVDD.n3637 0.00245
R10569 DVDD.n5134 DVDD.n5104 0.00245
R10570 DVDD.n5316 DVDD.n462 0.00245
R10571 DVDD.n5243 DVDD.n5242 0.00245
R10572 DVDD.n5085 DVDD.n570 0.00245
R10573 DVDD.n3617 DVDD.n2026 0.00242
R10574 DVDD.n3652 DVDD.n1995 0.00242
R10575 DVDD.n3786 DVDD.n1852 0.00239
R10576 DVDD.n5361 DVDD.n402 0.00239
R10577 DVDD.n5359 DVDD.n5358 0.00239
R10578 DVDD.n4880 DVDD.n702 0.00239
R10579 DVDD.n4886 DVDD.n695 0.00239
R10580 DVDD.n4875 DVDD.n704 0.00239
R10581 DVDD.n4877 DVDD.n715 0.00239
R10582 DVDD.n4771 DVDD.n4770 0.00239
R10583 DVDD.n4800 DVDD.n4773 0.00239
R10584 DVDD.n1095 DVDD.n361 0.00238
R10585 DVDD.n4441 DVDD.n4440 0.00238
R10586 DVDD.n1094 DVDD.n991 0.00238
R10587 DVDD.n4721 DVDD.n907 0.00238
R10588 DVDD.n4258 DVDD.n4257 0.00238
R10589 DVDD.n2491 DVDD.n2490 0.00236429
R10590 DVDD.n1395 DVDD.n1305 0.00236429
R10591 DVDD.n1394 DVDD.n1310 0.00236429
R10592 DVDD.n3652 DVDD.n1993 0.00236
R10593 DVDD.n3652 DVDD.n1991 0.00236
R10594 DVDD.n5631 DVDD.n5570 0.00235886
R10595 DVDD.n5530 DVDD.n24 0.00235886
R10596 DVDD.n4683 DVDD.n4651 0.00235886
R10597 DVDD.n5456 DVDD.n279 0.00235886
R10598 DVDD.n5812 DVDD.n150 0.00234426
R10599 DVDD.n5168 DVDD.n466 0.00234426
R10600 DVDD.n4970 DVDD.n4942 0.00234426
R10601 DVDD.n792 DVDD.n791 0.00234426
R10602 DVDD.n4526 DVDD.n4501 0.00234426
R10603 DVDD.n1933 DVDD.n1925 0.00233
R10604 DVDD.n1939 DVDD.n1936 0.00233
R10605 DVDD.n1960 DVDD.n1950 0.00233
R10606 DVDD.n3699 DVDD.n3696 0.00233
R10607 DVDD.n2398 DVDD 0.0023
R10608 DVDD.n2980 DVDD 0.0023
R10609 DVDD.n4033 DVDD.n1794 0.0023
R10610 DVDD.n4259 DVDD.n4258 0.0023
R10611 DVDD.n3902 DVDD.n3867 0.0023
R10612 DVDD.n3879 DVDD.n1792 0.0023
R10613 DVDD.n4283 DVDD.n1666 0.0023
R10614 DVDD.n4282 DVDD.n1670 0.0023
R10615 DVDD.n1361 DVDD 0.0023
R10616 DVDD.n4431 DVDD.n271 0.0023
R10617 DVDD.n5475 DVDD.n273 0.0023
R10618 DVDD.n4698 DVDD.n975 0.0023
R10619 DVDD.n4643 DVDD.n971 0.0023
R10620 DVDD.n5484 DVDD.n5483 0.00226879
R10621 DVDD.n5658 DVDD.n5657 0.00226471
R10622 DVDD.n5564 DVDD.n5563 0.00224
R10623 DVDD.n5649 DVDD.n5601 0.00224
R10624 DVDD.n31 DVDD.n7 0.00224
R10625 DVDD.n5955 DVDD.n5954 0.00224
R10626 DVDD.n1368 DVDD 0.00223571
R10627 DVDD.n5615 DVDD.n60 0.00220396
R10628 DVDD.n5440 DVDD.n305 0.00220396
R10629 DVDD.n2673 DVDD.n2672 0.00217143
R10630 DVDD.n3965 DVDD.n3927 0.00215
R10631 DVDD.n108 DVDD.n76 0.00206
R10632 DVDD.n5702 DVDD.n226 0.00206
R10633 DVDD.n5547 DVDD.n15 0.00204905
R10634 DVDD.n4666 DVDD.n982 0.00204905
R10635 DVDD.n4113 DVDD.n4112 0.00203
R10636 DVDD.n5920 DVDD.n80 0.00203
R10637 DVDD.n82 DVDD.n76 0.00203
R10638 DVDD.n5936 DVDD.n43 0.00203
R10639 DVDD.n5933 DVDD.n5932 0.00203
R10640 DVDD.n5952 DVDD.n32 0.00203
R10641 DVDD.n5951 DVDD.n29 0.00203
R10642 DVDD.n5708 DVDD.n5707 0.00203
R10643 DVDD.n226 DVDD.n220 0.00203
R10644 DVDD.n3647 DVDD.n1977 0.002
R10645 DVDD.n3704 DVDD.n3686 0.002
R10646 DVDD.n3253 DVDD.n2022 0.002
R10647 DVDD.n3647 DVDD.n2003 0.002
R10648 DVDD.n3704 DVDD.n1966 0.002
R10649 DVDD.n3305 DVDD.n2022 0.002
R10650 DVDD.n3647 DVDD.n1999 0.002
R10651 DVDD.n3704 DVDD.n1944 0.002
R10652 DVDD.n2055 DVDD.n2022 0.002
R10653 DVDD.n3647 DVDD.n2002 0.002
R10654 DVDD.n3704 DVDD.n1902 0.002
R10655 DVDD.n3836 DVDD.n1829 0.002
R10656 DVDD.n3854 DVDD.n1817 0.002
R10657 DVDD.n1161 DVDD.n325 0.002
R10658 DVDD.n353 DVDD.n328 0.002
R10659 DVDD.n5415 DVDD.n5405 0.002
R10660 DVDD.n4311 DVDD.n943 0.002
R10661 DVDD.n4708 DVDD.n4707 0.002
R10662 DVDD.n4711 DVDD.n4710 0.002
R10663 DVDD.n2456 DVDD.n2455 0.00197857
R10664 DVDD.n5744 DVDD.n174 0.00197541
R10665 DVDD.n567 DVDD.n486 0.00197541
R10666 DVDD.n628 DVDD.n610 0.00197541
R10667 DVDD.n864 DVDD.n705 0.00197541
R10668 DVDD.n1058 DVDD.n1010 0.00197541
R10669 DVDD.n5402 DVDD.n324 0.00197
R10670 DVDD.n5400 DVDD.n322 0.00197
R10671 DVDD.n297 DVDD.n295 0.00197
R10672 DVDD.n5472 DVDD.n307 0.00197
R10673 DVDD.n4638 DVDD.n974 0.00197
R10674 DVDD.n4636 DVDD.n972 0.00197
R10675 DVDD.n922 DVDD.n921 0.00197
R10676 DVDD.n4717 DVDD.n910 0.00197
R10677 DVDD.n3126 DVDD.n3122 0.00196739
R10678 DVDD.n3435 DVDD.n3434 0.00196739
R10679 DVDD.n4716 DVDD.n908 0.00194
R10680 DVDD.n4637 DVDD.n4635 0.00194
R10681 DVDD.n4438 DVDD.n990 0.00194
R10682 DVDD.n5401 DVDD.n358 0.00194
R10683 DVDD.n3803 DVDD.n1685 0.00194
R10684 DVDD.n3805 DVDD.n3804 0.00194
R10685 DVDD.n5400 DVDD.n5399 0.00194
R10686 DVDD.n359 DVDD.n307 0.00194
R10687 DVDD.n4636 DVDD.n909 0.00194
R10688 DVDD.n4718 DVDD.n4717 0.00194
R10689 DVDD.n3637 DVDD.n2007 0.00191
R10690 DVDD.n4218 DVDD.n4175 0.00191
R10691 DVDD.n2288 DVDD.n2287 0.00185
R10692 DVDD.n2549 DVDD.n2295 0.00185
R10693 DVDD.n4223 DVDD.n1724 0.00185
R10694 DVDD.n4224 DVDD.n1722 0.00185
R10695 DVDD.n3967 DVDD.n3923 0.00185
R10696 DVDD.n3620 DVDD.n2022 0.00184
R10697 DVDD.n3647 DVDD.n3646 0.00184
R10698 DVDD.n3704 DVDD.n3703 0.00184
R10699 DVDD.n3218 DVDD.n2022 0.00184
R10700 DVDD.n3647 DVDD.n2004 0.00184
R10701 DVDD.n3704 DVDD.n1965 0.00184
R10702 DVDD.n3100 DVDD.n2022 0.00184
R10703 DVDD.n3647 DVDD.n2000 0.00184
R10704 DVDD.n3704 DVDD.n1943 0.00184
R10705 DVDD.n3084 DVDD.n2022 0.00184
R10706 DVDD.n3647 DVDD.n2001 0.00184
R10707 DVDD.n3704 DVDD.n1901 0.00184
R10708 DVDD.n3654 DVDD.n3653 0.00179
R10709 DVDD.n4157 DVDD.n4156 0.00179
R10710 DVDD.n5415 DVDD.n324 0.00179
R10711 DVDD.n4710 DVDD.n922 0.00179
R10712 DVDD.n5455 DVDD.n5454 0.00174855
R10713 DVDD.n5630 DVDD.n5629 0.00174567
R10714 DVDD.n5548 DVDD.n20 0.00173924
R10715 DVDD.n4665 DVDD.n4647 0.00173924
R10716 DVDD.n3617 DVDD.n3098 0.00173
R10717 DVDD.n3617 DVDD.n3096 0.00173
R10718 DVDD.n4253 DVDD.n1691 0.00173
R10719 DVDD.n4119 DVDD.n4118 0.00173
R10720 DVDD.n4802 DVDD.n732 0.0017
R10721 DVDD.n4872 DVDD.n4871 0.0017
R10722 DVDD.n4881 DVDD.n696 0.0017
R10723 DVDD.n407 DVDD.n399 0.0017
R10724 DVDD.n2397 DVDD 0.0017
R10725 DVDD.n4285 DVDD.n4284 0.0017
R10726 DVDD.n4102 DVDD.n1790 0.0017
R10727 DVDD.n3973 DVDD.n1818 0.0017
R10728 DVDD.n3975 DVDD.n3974 0.0017
R10729 DVDD.n405 DVDD.n402 0.0017
R10730 DVDD.n4880 DVDD.n4879 0.0017
R10731 DVDD.n4878 DVDD.n704 0.0017
R10732 DVDD.n4770 DVDD.n703 0.0017
R10733 DVDD.n3668 DVDD.n3667 0.00167
R10734 DVDD.n4245 DVDD.n1695 0.00167
R10735 DVDD.n5359 DVDD.n405 0.00167
R10736 DVDD.n5881 DVDD.n108 0.00167
R10737 DVDD.n116 DVDD.n107 0.00167
R10738 DVDD.n5912 DVDD.n5907 0.00167
R10739 DVDD.n4879 DVDD.n695 0.00167
R10740 DVDD.n4878 DVDD.n4877 0.00167
R10741 DVDD.n4773 DVDD.n703 0.00167
R10742 DVDD.n5702 DVDD.n5701 0.00167
R10743 DVDD.n241 DVDD.n227 0.00167
R10744 DVDD.n5704 DVDD.n234 0.00167
R10745 DVDD DVDD.n1741 0.00165261
R10746 DVDD.n1743 DVDD 0.00165261
R10747 DVDD.n2190 DVDD.n2175 0.00164716
R10748 DVDD.n2187 DVDD.n2186 0.00164716
R10749 DVDD.n2183 DVDD.n2179 0.00164716
R10750 DVDD.n2182 DVDD.n2180 0.00164716
R10751 DVDD.n3709 DVDD.n3707 0.00164716
R10752 DVDD.n3708 DVDD.n1893 0.00164716
R10753 DVDD.n3714 DVDD.n3713 0.00164716
R10754 DVDD.n1894 DVDD.n1889 0.00164716
R10755 DVDD.n1728 DVDD.n1722 0.001625
R10756 DVDD.n4166 DVDD.n1769 0.00161
R10757 DVDD.n5828 DVDD.n163 0.00160656
R10758 DVDD.n5184 DVDD.n468 0.00160656
R10759 DVDD.n4954 DVDD.n4944 0.00160656
R10760 DVDD.n744 DVDD.n742 0.00160656
R10761 DVDD.n4510 DVDD.n4503 0.00160656
R10762 DVDD.n2598 DVDD.n2597 0.00159286
R10763 DVDD.n2200 DVDD.n2198 0.00159286
R10764 DVDD.n2601 DVDD.n2205 0.00159286
R10765 DVDD.n2492 DVDD.n2323 0.00159286
R10766 DVDD.n2618 DVDD.n2613 0.00159286
R10767 DVDD.n2609 DVDD.n2168 0.00159286
R10768 DVDD.n2621 DVDD.n2620 0.00159286
R10769 DVDD.n2682 DVDD.n2681 0.00159286
R10770 DVDD.n2865 DVDD.n2864 0.00159286
R10771 DVDD.n2688 DVDD.n2136 0.00159286
R10772 DVDD.n3022 DVDD.n3021 0.00159286
R10773 DVDD.n3636 DVDD.n2016 0.00155
R10774 DVDD.n3296 DVDD.n3274 0.00152
R10775 DVDD.n3361 DVDD.n3281 0.00152
R10776 DVDD.n3358 DVDD.n3295 0.00152
R10777 DVDD.n3307 DVDD.n3098 0.00152
R10778 DVDD.n3616 DVDD.n3099 0.00152
R10779 DVDD.n3267 DVDD.n3248 0.00152
R10780 DVDD.n3261 DVDD.n3257 0.00152
R10781 DVDD.n3389 DVDD.n3229 0.00152
R10782 DVDD.n3230 DVDD.n3096 0.00152
R10783 DVDD.n3398 DVDD.n3095 0.00152
R10784 DVDD.n5320 DVDD.n449 0.00149
R10785 DVDD.n5319 DVDD.n5318 0.00149
R10786 DVDD.n485 DVDD.n450 0.00149
R10787 DVDD.n5094 DVDD.n571 0.00149
R10788 DVDD.n2848 DVDD.n2691 0.00147826
R10789 DVDD.n1095 DVDD.n357 0.00146
R10790 DVDD.n4440 DVDD.n4439 0.00146
R10791 DVDD.n1094 DVDD.n989 0.00146
R10792 DVDD.n4715 DVDD.n907 0.00146
R10793 DVDD.n5046 DVDD.n481 0.00146
R10794 DVDD.n5245 DVDD.n482 0.00146
R10795 DVDD.n5247 DVDD.n5246 0.00146
R10796 DVDD.n5322 DVDD.n448 0.00146
R10797 DVDD.n3654 DVDD.n3652 0.00146
R10798 DVDD.n4258 DVDD.n1687 0.00146
R10799 DVDD.n4031 DVDD.n1792 0.00146
R10800 DVDD.n4033 DVDD.n4032 0.00146
R10801 DVDD.n5321 DVDD.n5320 0.00146
R10802 DVDD.n5319 DVDD.n451 0.00146
R10803 DVDD.n4836 DVDD.n450 0.00146
R10804 DVDD.n5045 DVDD.n571 0.00146
R10805 DVDD.n5531 DVDD.n12 0.00142943
R10806 DVDD.n4682 DVDD.n979 0.00142943
R10807 DVDD.n2833 DVDD.n2090 0.0014
R10808 DVDD.n4222 DVDD.n4221 0.0014
R10809 DVDD.n5687 DVDD 0.00134
R10810 DVDD.n5970 DVDD 0.00134
R10811 DVDD.n5589 DVDD 0.00134
R10812 DVDD.n5895 DVDD 0.00134
R10813 DVDD.n4195 DVDD 0.00134
R10814 DVDD.n4194 DVDD 0.00134
R10815 DVDD.n2531 DVDD.n2530 0.00133571
R10816 DVDD.n2945 DVDD.n2944 0.00133571
R10817 DVDD.n2097 DVDD.n2088 0.00133571
R10818 DVDD.n2948 DVDD.n2947 0.00133571
R10819 DVDD.n1557 DVDD.n1556 0.00133571
R10820 DVDD.n1554 DVDD.n1218 0.00133571
R10821 DVDD.n3384 DVDD.n3235 0.00131081
R10822 DVDD.n3338 DVDD.n3279 0.00131081
R10823 DVDD.n4139 DVDD.n1712 0.00131
R10824 DVDD.n699 DVDD.n698 0.0013
R10825 DVDD.n4883 DVDD.n4882 0.0013
R10826 DVDD.n731 DVDD.n697 0.0013
R10827 DVDD.n4766 DVDD.n4765 0.0013
R10828 DVDD.n3972 DVDD.n1817 0.0013
R10829 DVDD.n5561 DVDD.n68 0.00127453
R10830 DVDD.n5650 DVDD.n49 0.00127453
R10831 DVDD.n5566 DVDD.n67 0.00127453
R10832 DVDD.n5567 DVDD.n66 0.00127453
R10833 DVDD.n5608 DVDD.n51 0.00127453
R10834 DVDD.n5568 DVDD.n65 0.00127453
R10835 DVDD.n5607 DVDD.n52 0.00127453
R10836 DVDD.n5569 DVDD.n64 0.00127453
R10837 DVDD.n5606 DVDD.n53 0.00127453
R10838 DVDD.n5570 DVDD.n63 0.00127453
R10839 DVDD.n5605 DVDD.n54 0.00127453
R10840 DVDD.n5571 DVDD.n62 0.00127453
R10841 DVDD.n5604 DVDD.n55 0.00127453
R10842 DVDD.n5572 DVDD.n61 0.00127453
R10843 DVDD.n5603 DVDD.n56 0.00127453
R10844 DVDD.n5573 DVDD.n60 0.00127453
R10845 DVDD.n5602 DVDD.n57 0.00127453
R10846 DVDD.n5574 DVDD.n59 0.00127453
R10847 DVDD.n5931 DVDD.n69 0.00127453
R10848 DVDD.n70 DVDD.n48 0.00127453
R10849 DVDD.n270 DVDD.n268 0.00127453
R10850 DVDD.n5476 DVDD.n272 0.00127453
R10851 DVDD.n298 DVDD.n275 0.00127453
R10852 DVDD.n299 DVDD.n276 0.00127453
R10853 DVDD.n315 DVDD.n292 0.00127453
R10854 DVDD.n300 DVDD.n277 0.00127453
R10855 DVDD.n314 DVDD.n291 0.00127453
R10856 DVDD.n301 DVDD.n278 0.00127453
R10857 DVDD.n313 DVDD.n290 0.00127453
R10858 DVDD.n302 DVDD.n279 0.00127453
R10859 DVDD.n312 DVDD.n289 0.00127453
R10860 DVDD.n303 DVDD.n280 0.00127453
R10861 DVDD.n311 DVDD.n288 0.00127453
R10862 DVDD.n304 DVDD.n281 0.00127453
R10863 DVDD.n310 DVDD.n287 0.00127453
R10864 DVDD.n305 DVDD.n282 0.00127453
R10865 DVDD.n309 DVDD.n286 0.00127453
R10866 DVDD.n306 DVDD.n283 0.00127453
R10867 DVDD.n308 DVDD.n285 0.00127453
R10868 DVDD.n5474 DVDD.n5473 0.00127453
R10869 DVDD DVDD.n1740 0.00126841
R10870 DVDD.n5418 DVDD.n103 0.00124896
R10871 DVDD.n3503 DVDD.n3191 0.0012337
R10872 DVDD.n3508 DVDD.n3174 0.0012337
R10873 DVDD.n3519 DVDD.n3156 0.0012337
R10874 DVDD.n3528 DVDD.n3163 0.0012337
R10875 DVDD.n5712 DVDD.n5710 0.00122
R10876 DVDD.n5940 DVDD.n38 0.00122
R10877 DVDD.n5282 DVDD.n44 0.00122
R10878 DVDD.n5875 DVDD.n119 0.00122
R10879 DVDD.n4169 DVDD.n1724 0.00122
R10880 DVDD.n4168 DVDD.n1722 0.00122
R10881 DVDD.n5874 DVDD.n41 0.00122
R10882 DVDD.n5937 DVDD.n42 0.00122
R10883 DVDD.n5939 DVDD.n5938 0.00122
R10884 DVDD.n5711 DVDD.n40 0.00122
R10885 DVDD.n2354 DVDD.n2353 0.00120714
R10886 DVDD.n2474 DVDD.n2361 0.00120714
R10887 DVDD.n2014 DVDD 0.00119767
R10888 DVDD.n3662 DVDD 0.00119767
R10889 DVDD.n2011 DVDD 0.00119767
R10890 DVDD.n3659 DVDD 0.00119767
R10891 DVDD.n1706 DVDD.n1700 0.00119
R10892 DVDD.n4238 DVDD.n1707 0.00119
R10893 DVDD.n478 DVDD.n447 0.00114
R10894 DVDD.n5249 DVDD.n5248 0.00114
R10895 DVDD.n4833 DVDD.n477 0.00114
R10896 DVDD.n5048 DVDD.n5047 0.00114
R10897 DVDD.n4102 DVDD.n1789 0.00114
R10898 DVDD.n3674 DVDD.n1975 0.00113
R10899 DVDD.n5515 DVDD.n27 0.00111962
R10900 DVDD.n4697 DVDD.n4654 0.00111962
R10901 DVDD.n4149 DVDD.n4148 0.00107
R10902 DVDD.n107 DVDD.n77 0.00107
R10903 DVDD.n5912 DVDD.n79 0.00107
R10904 DVDD.n241 DVDD.n224 0.00107
R10905 DVDD.n5705 DVDD.n5704 0.00107
R10906 DVDD.n5894 DVDD 0.00106
R10907 DVDD.n5588 DVDD 0.00106
R10908 DVDD.n3643 DVDD.n3642 0.00101
R10909 DVDD.n3775 DVDD.n3734 0.00101
R10910 DVDD.n3752 DVDD.n1856 0.00101
R10911 DVDD.n3778 DVDD.n3777 0.00101
R10912 DVDD.n3996 DVDD.n3995 0.00101
R10913 DVDD.n1181 DVDD.n1120 0.00101
R10914 DVDD.n1579 DVDD.n1121 0.00101
R10915 DVDD.n1582 DVDD.n1131 0.00101
R10916 DVDD.n4411 DVDD.n4410 0.00101
R10917 DVDD.n4398 DVDD.n1108 0.00101
R10918 DVDD.n4415 DVDD.n4414 0.00101
R10919 DVDD.n4373 DVDD.n1595 0.00101
R10920 DVDD.n4383 DVDD.n1596 0.00101
R10921 DVDD.n4386 DVDD.n1607 0.00101
R10922 DVDD.n4330 DVDD.n1627 0.00101
R10923 DVDD.n4340 DVDD.n1628 0.00101
R10924 DVDD.n4343 DVDD.n1639 0.00101
R10925 DVDD.n3560 DVDD 0.00098913
R10926 DVDD.n2842 DVDD.n2683 0.00098913
R10927 DVDD.n5877 DVDD.n5876 0.00098
R10928 DVDD.n5281 DVDD.n35 0.00098
R10929 DVDD.n5942 DVDD.n5941 0.00098
R10930 DVDD.n215 DVDD.n34 0.00098
R10931 DVDD.n4221 DVDD.n4170 0.00098
R10932 DVDD.n5647 DVDD.n50 0.000964716
R10933 DVDD.n5471 DVDD.n316 0.000964716
R10934 DVDD.n2259 DVDD.n2255 0.00095
R10935 DVDD.n2824 DVDD.n2093 0.00095
R10936 DVDD.n3063 DVDD.n3028 0.00095
R10937 DVDD.n5382 DVDD.n5381 0.00095
R10938 DVDD.n5379 DVDD.n379 0.00095
R10939 DVDD.n4560 DVDD.n1075 0.00095
R10940 DVDD.n4497 DVDD.n1073 0.00095
R10941 DVDD.n4619 DVDD.n1005 0.00095
R10942 DVDD.n4616 DVDD.n4615 0.00095
R10943 DVDD.n4742 DVDD.n4741 0.00095
R10944 DVDD.n4744 DVDD.n891 0.00095
R10945 DVDD.n3758 DVDD.n3754 0.000917149
R10946 DVDD.n3768 DVDD.n3759 0.000917149
R10947 DVDD.n3767 DVDD.n3760 0.000917149
R10948 DVDD.n3764 DVDD.n3763 0.000917149
R10949 DVDD.n4288 DVDD.n1665 0.000917149
R10950 DVDD.n4289 DVDD.n1663 0.000917149
R10951 DVDD.n4294 DVDD.n4292 0.000917149
R10952 DVDD.n4293 DVDD.n1659 0.000917149
R10953 DVDD.n1383 DVDD.n1306 0.000912844
R10954 DVDD.n1321 DVDD.n1220 0.000912844
R10955 DVDD.n2008 DVDD.n1983 0.00089
R10956 DVDD.n4015 DVDD.n4014 0.00089
R10957 DVDD.n5849 DVDD.n137 0.00089
R10958 DVDD.n5856 DVDD.n130 0.00089
R10959 DVDD.n144 DVDD.n143 0.00089
R10960 DVDD.n5834 DVDD.n155 0.00089
R10961 DVDD.n5783 DVDD.n180 0.00089
R10962 DVDD.n537 DVDD.n169 0.00089
R10963 DVDD.n197 DVDD.n196 0.00089
R10964 DVDD.n5733 DVDD.n5727 0.00089
R10965 DVDD.n2049 DVDD.n2046 0.00083
R10966 DVDD.n2051 DVDD.n2050 0.00083
R10967 DVDD.n2058 DVDD.n2042 0.00083
R10968 DVDD.n2057 DVDD.n2026 0.00083
R10969 DVDD.n3086 DVDD.n2027 0.00083
R10970 DVDD.n2071 DVDD.n2070 0.00083
R10971 DVDD.n2068 DVDD.n2030 0.00083
R10972 DVDD.n2066 DVDD.n2031 0.00083
R10973 DVDD.n2065 DVDD.n2032 0.00083
R10974 DVDD.n3575 DVDD.n3143 0.00083
R10975 DVDD.n3572 DVDD.n3571 0.00083
R10976 DVDD.n3568 DVDD.n3159 0.00083
R10977 DVDD.n3200 DVDD.n3172 0.00083
R10978 DVDD.n3452 DVDD.n3171 0.00083
R10979 DVDD.n3513 DVDD.n3173 0.00083
R10980 DVDD.n4128 DVDD.n4127 0.00083
R10981 DVDD.n5648 DVDD.n5647 0.000809811
R10982 DVDD.n5614 DVDD.n5602 0.000809811
R10983 DVDD.n316 DVDD.n293 0.000809811
R10984 DVDD.n5439 DVDD.n286 0.000809811
R10985 DVDD.n5427 DVDD.n325 0.0008
R10986 DVDD.n353 DVDD.n321 0.0008
R10987 DVDD.n4706 DVDD.n943 0.0008
R10988 DVDD.n4708 DVDD.n914 0.0008
R10989 DVDD.n3664 DVDD.n1980 0.00077
R10990 DVDD.n111 DVDD.n90 0.000731959
R10991 DVDD.n5916 DVDD.n102 0.000731959
R10992 DVDD.n5407 DVDD.n344 0.000731959
R10993 DVDD.n5421 DVDD.n349 0.000731959
R10994 DVDD.n937 DVDD.n916 0.000731959
R10995 DVDD.n956 DVDD.n923 0.000731959
R10996 DVDD.n5703 DVDD.n5672 0.000731959
R10997 DVDD.n249 DVDD.n229 0.000731959
R10998 DVDD.n3952 DVDD.n3951 0.00071
R10999 DVDD.n2397 DVDD 0.000671429
R11000 DVDD.n2979 DVDD 0.000671429
R11001 DVDD.n1360 DVDD 0.000671429
R11002 DVDD.n3607 DVDD.n3606 0.00065
R11003 DVDD.n3601 DVDD.n3109 0.00065
R11004 DVDD.n3600 DVDD.n3114 0.00065
R11005 DVDD.n3597 DVDD.n3596 0.00065
R11006 DVDD.n3119 DVDD.n1993 0.00065
R11007 DVDD.n3588 DVDD.n1992 0.00065
R11008 DVDD.n3587 DVDD.n3128 0.00065
R11009 DVDD.n3584 DVDD.n3583 0.00065
R11010 DVDD.n3141 DVDD.n3133 0.00065
R11011 DVDD.n3576 DVDD.n3142 0.00065
R11012 DVDD.n3408 DVDD.n3407 0.00065
R11013 DVDD.n3420 DVDD.n3419 0.00065
R11014 DVDD.n3410 DVDD.n3409 0.00065
R11015 DVDD.n3428 DVDD.n3211 0.00065
R11016 DVDD.n3427 DVDD.n1991 0.00065
R11017 DVDD.n3438 DVDD.n1990 0.00065
R11018 DVDD.n3437 DVDD.n3205 0.00065
R11019 DVDD.n3447 DVDD.n3446 0.00065
R11020 DVDD.n3464 DVDD.n3197 0.00065
R11021 DVDD.n3463 DVDD.n3198 0.00065
R11022 DVDD.n3628 DVDD.n3626 0.00065
R11023 DVDD.n2064 DVDD.n2063 0.00059
R11024 DVDD.n2061 DVDD.n2035 0.00059
R11025 DVDD.n2038 DVDD.n2036 0.00059
R11026 DVDD.n3069 DVDD.n2037 0.00059
R11027 DVDD.n3070 DVDD.n1995 0.00059
R11028 DVDD.n3040 DVDD.n1996 0.00059
R11029 DVDD.n3044 DVDD.n3043 0.00059
R11030 DVDD.n3041 DVDD.n3036 0.00059
R11031 DVDD.n3052 DVDD.n3051 0.00059
R11032 DVDD.n3054 DVDD.n3034 0.00059
R11033 DVDD.n3805 DVDD.n1690 0.00059
R11034 DVDD.n5894 DVDD 0.00058
R11035 DVDD.n5588 DVDD 0.00058
R11036 DVDD.n5969 DVDD 0.00058
R11037 DVDD.n5686 DVDD 0.00058
R11038 DVDD DVDD.n4196 0.00058
R11039 DVDD.n1368 DVDD.n1337 0.000564286
R11040 DVDD.n1340 DVDD.n1331 0.000564286
R11041 DVDD.n3805 DVDD.n1684 0.00055625
R11042 DVDD.n5341 DVDD.n5340 0.00053
R11043 DVDD.n5338 DVDD.n426 0.00053
R11044 DVDD.n5004 DVDD.n674 0.00053
R11045 DVDD.n4938 DVDD.n672 0.00053
R11046 DVDD.n5012 DVDD.n605 0.00053
R11047 DVDD.n616 DVDD.n603 0.00053
R11048 DVDD.n5021 DVDD.n5020 0.00053
R11049 DVDD.n591 DVDD.n584 0.00053
R11050 GF_NI_IN_C_BASE_0.comp018green_out_predrv_1.ENB GF_NI_IN_C_BASE_0.comp018green_out_predrv_1.ENB.t3 82.1164
R11051 GF_NI_IN_C_BASE_0.comp018green_out_predrv_1.ENB GF_NI_IN_C_BASE_0.comp018green_out_predrv_1.ENB.t2 42.2319
R11052 GF_NI_IN_C_BASE_0.comp018green_out_predrv_1.ENB GF_NI_IN_C_BASE_0.comp018green_out_predrv_1.ENB.t0 2.04837
R11053 GF_NI_IN_C_BASE_0.comp018green_out_predrv_1.ENB GF_NI_IN_C_BASE_0.comp018green_out_predrv_1.ENB.t1 1.49421
R11054 GF_NI_IN_C_BASE_0.comp018green_out_predrv_0.SLB.n5 GF_NI_IN_C_BASE_0.comp018green_out_predrv_0.SLB.t5 45.4098
R11055 GF_NI_IN_C_BASE_0.comp018green_out_predrv_0.SLB.n4 GF_NI_IN_C_BASE_0.comp018green_out_predrv_0.SLB.t7 45.4098
R11056 GF_NI_IN_C_BASE_0.comp018green_out_predrv_0.SLB.n2 GF_NI_IN_C_BASE_0.comp018green_out_predrv_0.SLB.t2 45.4098
R11057 GF_NI_IN_C_BASE_0.comp018green_out_predrv_0.SLB.n1 GF_NI_IN_C_BASE_0.comp018green_out_predrv_0.SLB.t3 45.4098
R11058 GF_NI_IN_C_BASE_0.comp018green_out_predrv_0.SLB.n5 GF_NI_IN_C_BASE_0.comp018green_out_predrv_0.SLB.t4 34.4148
R11059 GF_NI_IN_C_BASE_0.comp018green_out_predrv_0.SLB.n4 GF_NI_IN_C_BASE_0.comp018green_out_predrv_0.SLB.t9 34.4148
R11060 GF_NI_IN_C_BASE_0.comp018green_out_predrv_0.SLB.n2 GF_NI_IN_C_BASE_0.comp018green_out_predrv_0.SLB.t8 34.4148
R11061 GF_NI_IN_C_BASE_0.comp018green_out_predrv_0.SLB.n1 GF_NI_IN_C_BASE_0.comp018green_out_predrv_0.SLB.t6 34.4148
R11062 GF_NI_IN_C_BASE_0.comp018green_out_predrv_0.SLB.t1 GF_NI_IN_C_BASE_0.comp018green_out_predrv_0.SLB.n0 9.02147
R11063 GF_NI_IN_C_BASE_0.comp018green_out_predrv_0.SLB.n0 GF_NI_IN_C_BASE_0.comp018green_out_predrv_0.SLB.n3 6.99208
R11064 GF_NI_IN_C_BASE_0.comp018green_out_predrv_0.SLB GF_NI_IN_C_BASE_0.comp018green_out_predrv_0.SLB.n5 6.273
R11065 GF_NI_IN_C_BASE_0.comp018green_out_predrv_0.SLB GF_NI_IN_C_BASE_0.comp018green_out_predrv_0.SLB.n4 6.273
R11066 GF_NI_IN_C_BASE_0.comp018green_out_predrv_0.SLB GF_NI_IN_C_BASE_0.comp018green_out_predrv_0.SLB.n2 6.273
R11067 GF_NI_IN_C_BASE_0.comp018green_out_predrv_0.SLB GF_NI_IN_C_BASE_0.comp018green_out_predrv_0.SLB.n1 6.273
R11068 GF_NI_IN_C_BASE_0.comp018green_out_predrv_0.SLB.n3 GF_NI_IN_C_BASE_0.comp018green_out_predrv_0.SLB 5.57458
R11069 GF_NI_IN_C_BASE_0.comp018green_out_predrv_0.SLB.n0 GF_NI_IN_C_BASE_0.comp018green_out_predrv_0.SLB 5.57458
R11070 GF_NI_IN_C_BASE_0.comp018green_out_predrv_0.SLB.n0 GF_NI_IN_C_BASE_0.comp018green_out_predrv_0.SLB 4.26721
R11071 GF_NI_IN_C_BASE_0.comp018green_out_predrv_0.SLB.n3 GF_NI_IN_C_BASE_0.comp018green_out_predrv_0.SLB 4.26721
R11072 GF_NI_IN_C_BASE_0.comp018green_out_predrv_0.SLB.t0 GF_NI_IN_C_BASE_0.comp018green_out_predrv_0.SLB.t1 2.99904
R11073 GF_NI_IN_C_BASE_0.pdrive_x_<1>.n1 GF_NI_IN_C_BASE_0.pdrive_x_<1>.t4 113.415
R11074 GF_NI_IN_C_BASE_0.pdrive_x_<1>.n1 GF_NI_IN_C_BASE_0.pdrive_x_<1>.t5 112.626
R11075 GF_NI_IN_C_BASE_0.pdrive_x_<1>.t2 GF_NI_IN_C_BASE_0.pdrive_x_<1>.n0 6.12025
R11076 GF_NI_IN_C_BASE_0.pdrive_x_<1> GF_NI_IN_C_BASE_0.pdrive_x_<1>.n1 2.40503
R11077 GF_NI_IN_C_BASE_0.pdrive_x_<1>.t3 GF_NI_IN_C_BASE_0.pdrive_x_<1>.n0 2.26404
R11078 GF_NI_IN_C_BASE_0.pdrive_x_<1>.t1 GF_NI_IN_C_BASE_0.pdrive_x_<1> 1.43572
R11079 GF_NI_IN_C_BASE_0.pdrive_x_<1>.n0 GF_NI_IN_C_BASE_0.pdrive_x_<1>.t1 1.0357
R11080 GF_NI_IN_C_BASE_0.pdrive_x_<1> GF_NI_IN_C_BASE_0.pdrive_x_<1>.t0 0.779435
R11081 GF_NI_IN_C_BASE_0.pdrive_x_<1> GF_NI_IN_C_BASE_0.pdrive_x_<1>.t3 0.7439
R11082 GF_NI_IN_C_BASE_0.pdrive_y_<1> GF_NI_IN_C_BASE_0.pdrive_y_<1>.t4 115.45
R11083 GF_NI_IN_C_BASE_0.pdrive_y_<1>.t1 GF_NI_IN_C_BASE_0.pdrive_y_<1>.n0 6.10848
R11084 GF_NI_IN_C_BASE_0.pdrive_y_<1>.t3 GF_NI_IN_C_BASE_0.pdrive_y_<1>.n0 2.68197
R11085 GF_NI_IN_C_BASE_0.pdrive_y_<1>.n0 GF_NI_IN_C_BASE_0.pdrive_y_<1> 1.59857
R11086 GF_NI_IN_C_BASE_0.pdrive_y_<1>.n0 GF_NI_IN_C_BASE_0.pdrive_y_<1> 1.11715
R11087 GF_NI_IN_C_BASE_0.pdrive_y_<1> GF_NI_IN_C_BASE_0.pdrive_y_<1>.t2 0.773875
R11088 GF_NI_IN_C_BASE_0.pdrive_y_<1> GF_NI_IN_C_BASE_0.pdrive_y_<1>.t0 0.766858
R11089 GF_NI_IN_C_BASE_0.pdrive_y_<1> GF_NI_IN_C_BASE_0.pdrive_y_<1>.t3 0.7304
R11090 DVSS.n1845 DVSS.n1540 196056
R11091 DVSS.n3802 DVSS.n1202 37210.9
R11092 DVSS.n4760 DVSS.n4759 32551.1
R11093 DVSS.n4320 DVSS.n4319 32385.4
R11094 DVSS.n3801 DVSS.n3800 30893.3
R11095 DVSS.n1822 DVSS.n1794 30469.2
R11096 DVSS.n5337 DVSS.n5336 27088.7
R11097 DVSS.n5096 DVSS.n960 25861.7
R11098 DVSS.n4097 DVSS.n1540 21519.5
R11099 DVSS.n5336 DVSS.n962 20471.6
R11100 DVSS.n4163 DVSS.n1523 19823.1
R11101 DVSS.n5097 DVSS.n5096 19552.7
R11102 DVSS.n4172 DVSS.n1217 17654
R11103 DVSS.n4761 DVSS.n961 16516.8
R11104 DVSS.n4321 DVSS.n1450 16516.8
R11105 DVSS.n1217 DVSS.n1214 16432
R11106 DVSS.n3801 DVSS.n1524 16400
R11107 DVSS.n4138 DVSS.n4137 16252.3
R11108 DVSS.n5337 DVSS.n961 16242.7
R11109 DVSS.n1450 DVSS.n960 16242.7
R11110 DVSS.n4862 DVSS.n1204 16230.9
R11111 DVSS.n4849 DVSS.n1214 16230.9
R11112 DVSS.n4830 DVSS.n1217 16230.9
R11113 DVSS.n4173 DVSS.n4172 16230.9
R11114 DVSS.n4299 DVSS.n1463 16230.9
R11115 DVSS.n3800 DVSS.n2622 15030.2
R11116 DVSS.n2664 DVSS.n2622 14984.7
R11117 DVSS.n4163 DVSS.n4162 14824
R11118 DVSS.n4138 DVSS.n1524 14824
R11119 DVSS.n5338 DVSS.n5337 14769.2
R11120 DVSS.n5339 DVSS.n960 14767.1
R11121 DVSS.n3802 DVSS.n3801 13915.8
R11122 DVSS.n3513 DVSS.n2645 12369.1
R11123 DVSS.n3511 DVSS.n2625 12369.1
R11124 DVSS.n3510 DVSS.n2653 12369.1
R11125 DVSS.n3775 DVSS.n3772 12369.1
R11126 DVSS.n4162 DVSS.n4161 11473.2
R11127 DVSS.n4161 DVSS.n1204 10835.5
R11128 DVSS.n4870 DVSS.n1202 10290.4
R11129 DVSS.n1204 DVSS.n1202 8547.5
R11130 DVSS.n3800 DVSS.n3799 7940.47
R11131 DVSS.n4319 DVSS.n1451 7811.82
R11132 DVSS.n4097 DVSS.n4096 7328.63
R11133 DVSS.n4137 DVSS.n4136 6651.3
R11134 DVSS.n4171 DVSS.n4170 6538.35
R11135 DVSS.n3511 DVSS.n3510 6402.4
R11136 DVSS.n3772 DVSS.n3771 5994.44
R11137 DVSS.n3819 DVSS.n3802 5387.7
R11138 DVSS.n4850 DVSS.n1213 4902.86
R11139 DVSS.n4861 DVSS.n1205 4902.86
R11140 DVSS.n4829 DVSS.n1218 4902.86
R11141 DVSS.n4171 DVSS.n1463 4526.71
R11142 DVSS.n3509 DVSS.n2664 4493.06
R11143 DVSS.n3825 DVSS.n3824 4399.95
R11144 DVSS.n4137 DVSS.n1540 3491.91
R11145 DVSS.n4162 DVSS.n4160 3437.85
R11146 DVSS.n4160 DVSS.n1524 3435.27
R11147 DVSS.n2309 DVSS.t14 3354.59
R11148 DVSS.n2548 DVSS.t14 3354.59
R11149 DVSS.n4172 DVSS.n4171 3311.99
R11150 DVSS.n4098 DVSS.n4097 3307.91
R11151 DVSS.n4136 DVSS.n1523 3086.59
R11152 DVSS.n3510 DVSS.n3509 3080.18
R11153 DVSS.n4096 DVSS.n1554 2507.4
R11154 DVSS.n3770 DVSS.n1024 2402.48
R11155 DVSS.n5215 DVSS.n1024 2401.2
R11156 DVSS.n3770 DVSS.n1023 2400.01
R11157 DVSS.n5215 DVSS.n1023 2398.73
R11158 DVSS.n3512 DVSS.n3511 2352.1
R11159 DVSS.n4756 DVSS.n4755 2286.22
R11160 DVSS.n4509 DVSS.n4508 2282.35
R11161 DVSS.n4509 DVSS.n1393 2282.35
R11162 DVSS.n4508 DVSS.n4507 2278.48
R11163 DVSS.n4755 DVSS.n1393 2277.19
R11164 DVSS.n4104 DVSS.n1463 2219.8
R11165 DVSS.n4762 DVSS.n4756 2185.59
R11166 DVSS.n4507 DVSS.n4322 2179.14
R11167 DVSS.n3772 DVSS.n1794 2166.67
R11168 DVSS.n4161 DVSS.n1214 2099.5
R11169 DVSS.n4137 DVSS.n4135 1819.86
R11170 DVSS.n2622 DVSS.n2621 1783.15
R11171 DVSS.n4758 DVSS.n1203 1674.85
R11172 DVSS.n3513 DVSS.n3512 1481.53
R11173 DVSS.n1257 DVSS.t35 1472.87
R11174 DVSS.n1261 DVSS.t34 1472.87
R11175 DVSS.t32 DVSS.n1509 1472.87
R11176 DVSS.t30 DVSS.n1505 1472.87
R11177 DVSS.n4857 DVSS.n1209 1449.32
R11178 DVSS.n4839 DVSS.n1216 1375
R11179 DVSS.n2621 DVSS.n2620 1219.32
R11180 DVSS.n4838 DVSS.n4831 1124.46
R11181 DVSS.n4839 DVSS.n4838 1124.46
R11182 DVSS.n4839 DVSS.n1215 1124.46
R11183 DVSS.n4848 DVSS.n1215 1124.46
R11184 DVSS.n4828 DVSS.t146 1075.57
R11185 DVSS.t83 DVSS.n4851 1075.57
R11186 DVSS.n4860 DVSS.t198 1075.57
R11187 DVSS.n4870 DVSS.n1203 1041.24
R11188 DVSS.n4322 DVSS.n4321 967.646
R11189 DVSS.n4762 DVSS.n4761 967.646
R11190 DVSS.n4098 DVSS.n1553 835.686
R11191 DVSS.n4857 DVSS.t72 824.14
R11192 DVSS.t165 DVSS.n4857 824.14
R11193 DVSS.n4870 DVSS.n4869 796.203
R11194 DVSS.n2617 DVSS.t137 782.032
R11195 DVSS.n2622 DVSS.n1554 724.26
R11196 DVSS.n4831 DVSS.n4830 693.769
R11197 DVSS.n4849 DVSS.n4848 693.769
R11198 DVSS.n4869 DVSS.n4862 693.769
R11199 DVSS.t130 DVSS.t114 640.298
R11200 DVSS.t185 DVSS.t101 640.298
R11201 DVSS.t195 DVSS.t78 640.298
R11202 DVSS.t25 DVSS.t60 640.298
R11203 DVSS.n2620 DVSS.n1845 614.245
R11204 DVSS.n4321 DVSS.n4320 608.972
R11205 DVSS.n4761 DVSS.n4760 608.972
R11206 DVSS.t150 DVSS.n3823 587.904
R11207 DVSS.n2664 DVSS.n2663 562.811
R11208 DVSS.n4829 DVSS.n4828 547.1
R11209 DVSS.n4851 DVSS.n4850 547.1
R11210 DVSS.n4861 DVSS.n4860 547.1
R11211 DVSS.n3508 DVSS.n1792 517.379
R11212 DVSS.n3826 DVSS.n1792 517.379
R11213 DVSS.n3508 DVSS.n1793 517.379
R11214 DVSS.n3826 DVSS.n1793 517.379
R11215 DVSS.n1257 DVSS.n1230 488.243
R11216 DVSS.n1262 DVSS.n1261 488.243
R11217 DVSS.n1509 DVSS.n1464 488.243
R11218 DVSS.n1505 DVSS.n1472 488.243
R11219 DVSS.n4112 DVSS.n1549 486.896
R11220 DVSS.n1549 DVSS.n1548 472.783
R11221 DVSS.t126 DVSS.t31 463.173
R11222 DVSS.n4852 DVSS.t72 409.743
R11223 DVSS.n4858 DVSS.t165 409.743
R11224 DVSS.n3771 DVSS.n3513 407.959
R11225 DVSS.t162 DVSS.n4824 400.822
R11226 DVSS.n3777 DVSS.t104 367.289
R11227 DVSS.n2660 DVSS.n2654 344.332
R11228 DVSS.n2655 DVSS.n2654 344.332
R11229 DVSS.n3791 DVSS.n2631 344.332
R11230 DVSS.n3778 DVSS.n3776 344.332
R11231 DVSS.t179 DVSS.n1213 320.659
R11232 DVSS.t110 DVSS.n1623 306.072
R11233 DVSS.n1623 DVSS.t133 306.072
R11234 DVSS.t35 DVSS.n1256 303.188
R11235 DVSS.n1256 DVSS.t34 303.188
R11236 DVSS.n2655 DVSS.n2653 300.031
R11237 DVSS.n2653 DVSS.n2652 300.031
R11238 DVSS.n275 DVSS.t130 298.296
R11239 DVSS.n3938 DVSS.n1696 290.733
R11240 DVSS.n2633 DVSS.t21 287.95
R11241 DVSS.n4112 DVSS.n4111 285.283
R11242 DVSS.n5710 DVSS.t25 282.926
R11243 DVSS.n2628 DVSS.n2624 278.889
R11244 DVSS.n4120 DVSS.n4118 273.185
R11245 DVSS.t154 DVSS.t152 271.668
R11246 DVSS.t97 DVSS.t120 271.668
R11247 DVSS.t64 DVSS.t68 271.668
R11248 DVSS.t66 DVSS.t70 271.668
R11249 DVSS.t70 DVSS.t36 271.668
R11250 DVSS.t8 DVSS.n4809 271.668
R11251 DVSS.t167 DVSS.t8 271.668
R11252 DVSS.t35 DVSS.t29 271.668
R11253 DVSS.t128 DVSS.t17 271.668
R11254 DVSS.t17 DVSS.n4783 271.668
R11255 DVSS.t156 DVSS.t164 271.668
R11256 DVSS.n4104 DVSS.n1451 271
R11257 DVSS.n2645 DVSS.t16 270.834
R11258 DVSS.t68 DVSS.n1218 269.442
R11259 DVSS.n2641 DVSS.t139 256.738
R11260 DVSS.n4099 DVSS.n4098 255.427
R11261 DVSS.t152 DVSS.t156 252.742
R11262 DVSS.n4825 DVSS.t162 250.514
R11263 DVSS.n2652 DVSS.n2651 248.684
R11264 DVSS.t142 DVSS.t144 245.663
R11265 DVSS.t108 DVSS.t110 245.663
R11266 DVSS.t169 DVSS.t176 245.663
R11267 DVSS.t148 DVSS.t140 245.663
R11268 DVSS.t4 DVSS.t15 245.663
R11269 DVSS.t85 DVSS.t95 245.663
R11270 DVSS.n4318 DVSS.t200 241.587
R11271 DVSS.n3825 DVSS.n1794 239.081
R11272 DVSS.n1704 DVSS.t2 238.615
R11273 DVSS.n3778 DVSS.t76 235.595
R11274 DVSS.n2309 DVSS.n2308 233.749
R11275 DVSS.n2548 DVSS.n2547 233.749
R11276 DVSS.n4759 DVSS.n4758 232.701
R11277 DVSS.n3792 DVSS.n2630 227.541
R11278 DVSS.t34 DVSS.n1209 226.019
R11279 DVSS.n1523 DVSS.n1518 224.798
R11280 DVSS.n3823 DVSS.n3822 219.064
R11281 DVSS.t10 DVSS.n1683 216.465
R11282 DVSS.n2644 DVSS.t117 210.424
R11283 DVSS.n4174 DVSS.n4173 199.98
R11284 DVSS.n3775 DVSS.t183 192.303
R11285 DVSS.n4809 DVSS.t82 191.505
R11286 DVSS.t33 DVSS.n1507 188.571
R11287 DVSS.n3509 DVSS.n3508 184.061
R11288 DVSS.t63 DVSS.n2644 180.22
R11289 DVSS.t89 DVSS.t191 170.153
R11290 DVSS.t181 DVSS.t87 170.153
R11291 DVSS.n2616 DVSS.n1845 169.606
R11292 DVSS.n3937 DVSS.t3 169.145
R11293 DVSS.n4758 DVSS.t97 168.124
R11294 DVSS.n4057 DVSS.t133 166.125
R11295 DVSS.n4810 DVSS.t167 165.897
R11296 DVSS.n4784 DVSS.t128 165.897
R11297 DVSS.n3824 DVSS.t150 164.453
R11298 DVSS.n4311 DVSS.t5 163.742
R11299 DVSS.t28 DVSS.t30 163.742
R11300 DVSS.t38 DVSS.t40 163.742
R11301 DVSS.t114 DVSS.t185 161.953
R11302 DVSS.t60 DVSS.t195 161.953
R11303 DVSS.n4289 DVSS.t23 161.728
R11304 DVSS.n4852 DVSS.t83 158.31
R11305 DVSS.n4858 DVSS.t198 158.31
R11306 DVSS.t7 DVSS.t193 154.043
R11307 DVSS.t42 DVSS.t23 153.675
R11308 DVSS.n4303 DVSS.t200 152.333
R11309 DVSS.n4320 DVSS.n1023 152.252
R11310 DVSS.n4760 DVSS.n1024 152.252
R11311 DVSS.t19 DVSS.n3798 151.023
R11312 DVSS.t82 DVSS.n1216 150.309
R11313 DVSS.n4830 DVSS.n4829 146.669
R11314 DVSS.n4850 DVSS.n4849 146.669
R11315 DVSS.n4862 DVSS.n4861 146.669
R11316 DVSS.n4310 DVSS.t0 145.624
R11317 DVSS.t29 DVSS.n1213 142.516
R11318 DVSS.n3774 DVSS.t181 137.935
R11319 DVSS.n4111 DVSS.n1451 137.097
R11320 DVSS.n4757 DVSS.t154 135.834
R11321 DVSS.t120 DVSS.n4757 135.834
R11322 DVSS.n4812 DVSS.t64 135.834
R11323 DVSS.n4812 DVSS.t66 135.834
R11324 DVSS.n2641 DVSS.t117 133.906
R11325 DVSS.n4177 DVSS.n4176 132.07
R11326 DVSS.n4824 DVSS.n1218 131.381
R11327 DVSS.n4297 DVSS.n1452 129.345
R11328 DVSS.n4785 DVSS.n1263 129.345
R11329 DVSS.n4291 DVSS.n1473 129.345
R11330 DVSS.n4813 DVSS.n4811 129.345
R11331 DVSS.n4317 DVSS.n1452 128.957
R11332 DVSS.n1275 DVSS.n1263 128.957
R11333 DVSS.t171 DVSS.t46 125.49
R11334 DVSS.n1624 DVSS.t108 123.838
R11335 DVSS.t135 DVSS.n4056 123.838
R11336 DVSS.t93 DVSS.n3936 123.838
R11337 DVSS.n1510 DVSS.t32 122.806
R11338 DVSS.t144 DVSS.n1624 121.826
R11339 DVSS.n4056 DVSS.t176 121.826
R11340 DVSS.n1703 DVSS.t99 121.826
R11341 DVSS.n3936 DVSS.t191 121.826
R11342 DVSS.t36 DVSS.n1216 121.361
R11343 DVSS.n2645 DVSS.t63 119.811
R11344 DVSS.n4783 DVSS.n1205 118.02
R11345 DVSS.n4120 DVSS.n4119 114.919
R11346 DVSS.n4127 DVSS.n4126 114.919
R11347 DVSS.n4128 DVSS.n4127 114.919
R11348 DVSS.n4128 DVSS.n1541 114.919
R11349 DVSS.n4134 DVSS.n1541 114.919
R11350 DVSS.n4169 DVSS.n1518 114.919
R11351 DVSS.n4177 DVSS.n1503 112.962
R11352 DVSS.n4170 DVSS.n1517 112.903
R11353 DVSS.n4135 DVSS.n4134 111.895
R11354 DVSS.t76 DVSS.n3777 108.737
R11355 DVSS.t183 DVSS.n3774 107.73
R11356 DVSS.t46 DVSS.n4286 106.701
R11357 DVSS.n4810 DVSS.t179 105.773
R11358 DVSS.n4784 DVSS.t126 105.773
R11359 DVSS.n3822 DVSS.n1795 102.416
R11360 DVSS.n1259 DVSS.n1254 102.356
R11361 DVSS.n4178 DVSS.n1502 102.356
R11362 DVSS.t202 DVSS.t44 101.332
R11363 DVSS.t158 DVSS.t190 101.332
R11364 DVSS.n4290 DVSS.t106 99.9902
R11365 DVSS.n4764 DVSS.n959 99.728
R11366 DVSS.n5340 DVSS.n958 99.7229
R11367 DVSS.n4119 DVSS.n1545 98.7908
R11368 DVSS.t193 DVSS.t10 91.6207
R11369 DVSS.t99 DVSS.t7 91.6207
R11370 DVSS.t140 DVSS.t13 91.6207
R11371 DVSS.n2633 DVSS.n2630 90.6139
R11372 DVSS.n1507 DVSS.t11 90.5952
R11373 DVSS.t32 DVSS.n1503 89.3577
R11374 DVSS.t78 DVSS.n5709 87.8106
R11375 DVSS.t139 DVSS.n2631 87.5934
R11376 DVSS.n3824 DVSS.t104 86.3383
R11377 DVSS.n5710 DVSS.n59 86.0408
R11378 DVSS.n4287 DVSS.t81 85.2266
R11379 DVSS.n3798 DVSS.n2625 82.5594
R11380 DVSS.n4304 DVSS.t122 81.8712
R11381 DVSS.t124 DVSS.n4304 81.8712
R11382 DVSS.n275 DVSS.n59 80.8661
R11383 DVSS.n4305 DVSS.t174 80.5291
R11384 DVSS.n4057 DVSS.t135 79.5389
R11385 DVSS.t87 DVSS.t89 75.5117
R11386 DVSS.n5709 DVSS.t101 74.1437
R11387 DVSS.t164 DVSS.n1205 73.4846
R11388 DVSS.n2550 DVSS.n1918 73.4718
R11389 DVSS.n2550 DVSS.n2549 73.4718
R11390 DVSS.n2311 DVSS.n1921 73.2997
R11391 DVSS.n2311 DVSS.n2310 73.2997
R11392 DVSS.n4823 DVSS.n1223 72.4894
R11393 DVSS.n4176 DVSS.t30 70.25
R11394 DVSS.n4323 DVSS.n958 69.3341
R11395 DVSS.n4764 DVSS.n4763 69.3341
R11396 DVSS.t2 DVSS.t91 67.4571
R11397 DVSS.t3 DVSS.t93 67.4571
R11398 DVSS.t188 DVSS.n1222 65.0944
R11399 DVSS.n1553 DVSS.n1451 64.5166
R11400 DVSS.n4298 DVSS.t11 63.7523
R11401 DVSS.n4290 DVSS.t112 63.7523
R11402 DVSS.t44 DVSS.t124 62.4102
R11403 DVSS.t174 DVSS.t202 62.4102
R11404 DVSS.t160 DVSS.t158 62.4102
R11405 DVSS.t190 DVSS.t118 62.4102
R11406 DVSS.n1259 DVSS.n1258 61.1338
R11407 DVSS.n1260 DVSS.n1259 61.1338
R11408 DVSS.n1508 DVSS.n1502 61.1338
R11409 DVSS.n1504 DVSS.n1502 61.1338
R11410 DVSS.n1511 DVSS.n1506 59.6561
R11411 DVSS.n2617 DVSS.n1846 59.6561
R11412 DVSS.n3779 DVSS.n2639 59.6561
R11413 DVSS.n2659 DVSS.n2657 59.6561
R11414 DVSS.n2651 DVSS.t142 59.4026
R11415 DVSS.n5708 DVSS.n59 58.4662
R11416 DVSS.n4286 DVSS.t38 57.0416
R11417 DVSS.n1473 DVSS.n1223 56.4672
R11418 DVSS.n4813 DVSS.n1223 56.4672
R11419 DVSS.n3779 DVSS.n2637 56.0005
R11420 DVSS.n2643 DVSS.n2642 56.0005
R11421 DVSS.n2657 DVSS.n2656 56.0005
R11422 DVSS.t0 DVSS.n4299 54.3573
R11423 DVSS.t15 DVSS.t148 53.3617
R11424 DVSS.t95 DVSS.n3775 53.3617
R11425 DVSS.n4311 DVSS.t118 53.0152
R11426 DVSS.n4826 DVSS.n1222 53.0152
R11427 DVSS.n3799 DVSS.t19 46.314
R11428 DVSS.t31 DVSS.n1209 45.6497
R11429 DVSS.n4299 DVSS.n4298 45.6334
R11430 DVSS.n4174 DVSS.t28 44.9623
R11431 DVSS.n1510 DVSS.t33 40.9359
R11432 DVSS.n4297 DVSS.n1464 40.8338
R11433 DVSS.n4785 DVSS.n1262 40.8338
R11434 DVSS.n4811 DVSS.n1230 40.8338
R11435 DVSS.n4291 DVSS.n1472 40.8338
R11436 DVSS.n2254 DVSS.n1929 40.2769
R11437 DVSS.n2254 DVSS.n1919 40.2769
R11438 DVSS.n3822 DVSS.n3821 39.6013
R11439 DVSS.t81 DVSS.t171 38.2516
R11440 DVSS.n2663 DVSS.n2660 37.2527
R11441 DVSS.n4173 DVSS.t112 34.2252
R11442 DVSS.n3786 DVSS.n2632 33.0561
R11443 DVSS.t13 DVSS.n1703 32.2186
R11444 DVSS.n4287 DVSS.n1477 30.1987
R11445 DVSS.n5103 DVSS.n1079 29.3117
R11446 DVSS.n5104 DVSS.n5103 29.3117
R11447 DVSS.n5105 DVSS.n5104 29.3117
R11448 DVSS.n5105 DVSS.n1075 29.3117
R11449 DVSS.n5111 DVSS.n1075 29.3117
R11450 DVSS.n5112 DVSS.n5111 29.3117
R11451 DVSS.n5113 DVSS.n5112 29.3117
R11452 DVSS.n5113 DVSS.n1071 29.3117
R11453 DVSS.n5119 DVSS.n1071 29.3117
R11454 DVSS.n5120 DVSS.n5119 29.3117
R11455 DVSS.n5121 DVSS.n5120 29.3117
R11456 DVSS.n5121 DVSS.n1067 29.3117
R11457 DVSS.n5127 DVSS.n1067 29.3117
R11458 DVSS.n5128 DVSS.n5127 29.3117
R11459 DVSS.n5129 DVSS.n5128 29.3117
R11460 DVSS.n5129 DVSS.n1063 29.3117
R11461 DVSS.n5135 DVSS.n1063 29.3117
R11462 DVSS.n5136 DVSS.n5135 29.3117
R11463 DVSS.n5137 DVSS.n5136 29.3117
R11464 DVSS.n5137 DVSS.n1059 29.3117
R11465 DVSS.n5143 DVSS.n1059 29.3117
R11466 DVSS.n5144 DVSS.n5143 29.3117
R11467 DVSS.n5145 DVSS.n5144 29.3117
R11468 DVSS.n5145 DVSS.n1055 29.3117
R11469 DVSS.n5151 DVSS.n1055 29.3117
R11470 DVSS.n5152 DVSS.n5151 29.3117
R11471 DVSS.n5153 DVSS.n5152 29.3117
R11472 DVSS.n5153 DVSS.n1051 29.3117
R11473 DVSS.n5159 DVSS.n1051 29.3117
R11474 DVSS.n5160 DVSS.n5159 29.3117
R11475 DVSS.n5161 DVSS.n5160 29.3117
R11476 DVSS.n5161 DVSS.n1047 29.3117
R11477 DVSS.n5167 DVSS.n1047 29.3117
R11478 DVSS.n5168 DVSS.n5167 29.3117
R11479 DVSS.n5169 DVSS.n5168 29.3117
R11480 DVSS.n5169 DVSS.n1043 29.3117
R11481 DVSS.n5175 DVSS.n1043 29.3117
R11482 DVSS.n5176 DVSS.n5175 29.3117
R11483 DVSS.n5177 DVSS.n5176 29.3117
R11484 DVSS.n5177 DVSS.n1039 29.3117
R11485 DVSS.n5183 DVSS.n1039 29.3117
R11486 DVSS.n5184 DVSS.n5183 29.3117
R11487 DVSS.n5185 DVSS.n5184 29.3117
R11488 DVSS.n5185 DVSS.n1035 29.3117
R11489 DVSS.n5191 DVSS.n1035 29.3117
R11490 DVSS.n5192 DVSS.n5191 29.3117
R11491 DVSS.n5193 DVSS.n5192 29.3117
R11492 DVSS.n5193 DVSS.n1031 29.3117
R11493 DVSS.n5199 DVSS.n1031 29.3117
R11494 DVSS.n5200 DVSS.n5199 29.3117
R11495 DVSS.n5201 DVSS.n5200 29.3117
R11496 DVSS.n5201 DVSS.n1027 29.3117
R11497 DVSS.n5208 DVSS.n1027 29.3117
R11498 DVSS.n5209 DVSS.n5208 29.3117
R11499 DVSS.n5210 DVSS.n5209 29.3117
R11500 DVSS.n5210 DVSS.n1022 29.3117
R11501 DVSS.n5218 DVSS.n5217 29.3117
R11502 DVSS.n5218 DVSS.n1018 29.3117
R11503 DVSS.n5224 DVSS.n1018 29.3117
R11504 DVSS.n5225 DVSS.n5224 29.3117
R11505 DVSS.n5226 DVSS.n5225 29.3117
R11506 DVSS.n5226 DVSS.n1014 29.3117
R11507 DVSS.n5232 DVSS.n1014 29.3117
R11508 DVSS.n5233 DVSS.n5232 29.3117
R11509 DVSS.n5234 DVSS.n5233 29.3117
R11510 DVSS.n5234 DVSS.n1010 29.3117
R11511 DVSS.n5240 DVSS.n1010 29.3117
R11512 DVSS.n5241 DVSS.n5240 29.3117
R11513 DVSS.n5242 DVSS.n5241 29.3117
R11514 DVSS.n5242 DVSS.n1006 29.3117
R11515 DVSS.n5248 DVSS.n1006 29.3117
R11516 DVSS.n5249 DVSS.n5248 29.3117
R11517 DVSS.n5250 DVSS.n5249 29.3117
R11518 DVSS.n5250 DVSS.n1002 29.3117
R11519 DVSS.n5256 DVSS.n1002 29.3117
R11520 DVSS.n5257 DVSS.n5256 29.3117
R11521 DVSS.n5258 DVSS.n5257 29.3117
R11522 DVSS.n5258 DVSS.n998 29.3117
R11523 DVSS.n5264 DVSS.n998 29.3117
R11524 DVSS.n5265 DVSS.n5264 29.3117
R11525 DVSS.n5266 DVSS.n5265 29.3117
R11526 DVSS.n5266 DVSS.n994 29.3117
R11527 DVSS.n5272 DVSS.n994 29.3117
R11528 DVSS.n5273 DVSS.n5272 29.3117
R11529 DVSS.n5274 DVSS.n5273 29.3117
R11530 DVSS.n5274 DVSS.n990 29.3117
R11531 DVSS.n5280 DVSS.n990 29.3117
R11532 DVSS.n5281 DVSS.n5280 29.3117
R11533 DVSS.n5282 DVSS.n5281 29.3117
R11534 DVSS.n5282 DVSS.n986 29.3117
R11535 DVSS.n5288 DVSS.n986 29.3117
R11536 DVSS.n5289 DVSS.n5288 29.3117
R11537 DVSS.n5290 DVSS.n5289 29.3117
R11538 DVSS.n5290 DVSS.n982 29.3117
R11539 DVSS.n5296 DVSS.n982 29.3117
R11540 DVSS.n5297 DVSS.n5296 29.3117
R11541 DVSS.n5298 DVSS.n5297 29.3117
R11542 DVSS.n5298 DVSS.n978 29.3117
R11543 DVSS.n5304 DVSS.n978 29.3117
R11544 DVSS.n5305 DVSS.n5304 29.3117
R11545 DVSS.n5306 DVSS.n5305 29.3117
R11546 DVSS.n5306 DVSS.n974 29.3117
R11547 DVSS.n5312 DVSS.n974 29.3117
R11548 DVSS.n5313 DVSS.n5312 29.3117
R11549 DVSS.n5314 DVSS.n5313 29.3117
R11550 DVSS.n5314 DVSS.n970 29.3117
R11551 DVSS.n5320 DVSS.n970 29.3117
R11552 DVSS.n5321 DVSS.n5320 29.3117
R11553 DVSS.n5322 DVSS.n5321 29.3117
R11554 DVSS.n5322 DVSS.n966 29.3117
R11555 DVSS.n5329 DVSS.n966 29.3117
R11556 DVSS.n5330 DVSS.n5329 29.3117
R11557 DVSS.n5331 DVSS.n5330 29.3117
R11558 DVSS.n2628 DVSS.t169 29.1981
R11559 DVSS.t16 DVSS.n1683 29.1981
R11560 DVSS.n4826 DVSS.t74 28.8566
R11561 DVSS.n3790 DVSS.n2632 26.6005
R11562 DVSS.n2642 DVSS.n2632 26.6005
R11563 DVSS.n3792 DVSS.n3791 26.1777
R11564 DVSS.n5097 DVSS.n1079 21.9839
R11565 DVSS.n4319 DVSS.n4318 21.4748
R11566 DVSS.n4305 DVSS.t160 20.8037
R11567 DVSS.n3799 DVSS.n2624 20.1368
R11568 DVSS.n5333 DVSS.n962 19.8563
R11569 DVSS.t5 DVSS.n4310 18.1194
R11570 DVSS.t40 DVSS.t188 16.7773
R11571 DVSS.n4126 DVSS.n1545 16.1295
R11572 DVSS.n1456 DVSS.t204 15.9461
R11573 DVSS.n4814 DVSS.t206 15.9461
R11574 DVSS.n1478 DVSS.t205 15.9461
R11575 DVSS.n1271 DVSS.t207 15.9461
R11576 DVSS.n5335 DVSS.n963 14.9905
R11577 DVSS.n5217 DVSS.n5216 14.8925
R11578 DVSS.n5095 DVSS.n5094 14.6859
R11579 DVSS.n5216 DVSS.n1022 14.4197
R11580 DVSS.n4118 DVSS.n1548 14.1134
R11581 DVSS.n2016 DVSS.n2015 12.4433
R11582 DVSS.t21 DVSS.n2625 12.0823
R11583 DVSS.n5331 DVSS.n962 12.0559
R11584 DVSS.n3794 DVSS.n3793 11.7115
R11585 DVSS.t122 DVSS.n4303 11.4087
R11586 DVSS.n4834 VSS 10.8266
R11587 DVSS.n4846 VSS 10.8266
R11588 DVSS.n4867 VSS 10.8266
R11589 DVSS.n3768 DVSS.n3522 10.6235
R11590 DVSS.n5093 DVSS.n1081 10.6235
R11591 DVSS.n4176 DVSS.n4175 10.3873
R11592 DVSS.n1506 DVSS.n1503 10.1573
R11593 DVSS.n1477 DVSS.t42 10.0666
R11594 DVSS.n5098 DVSS.n5097 9.92831
R11595 DVSS.n3937 DVSS.t91 9.06184
R11596 DVSS.n1836 DVSS.t86 8.35531
R11597 DVSS.n1837 DVSS.t86 8.13558
R11598 DVSS.n3769 DVSS.n3768 8.07493
R11599 DVSS.n3769 DVSS.n1081 8.03957
R11600 DVSS.t74 DVSS.n4825 7.95592
R11601 DVSS.n1921 DVSS.n1919 7.77509
R11602 DVSS.n2310 DVSS.n1929 7.77509
R11603 DVSS.n4754 DVSS.n1371 7.61966
R11604 DVSS.n4510 DVSS.n1449 7.60677
R11605 DVSS.n4510 DVSS.n1394 7.60677
R11606 DVSS.n1929 DVSS.n1918 7.60296
R11607 DVSS.n2549 DVSS.n1919 7.60296
R11608 DVSS.n4506 DVSS.n1449 7.59387
R11609 DVSS.n4754 DVSS.n1394 7.58957
R11610 DVSS.n4763 DVSS.n1371 7.28428
R11611 DVSS.n4506 DVSS.n4323 7.26279
R11612 DVSS.n1704 DVSS.t4 7.04821
R11613 DVSS.n3785 DVSS.n2634 6.95655
R11614 DVSS.n3783 VSS 6.91517
R11615 DVSS.n1848 DVSS.n1847 6.3005
R11616 DVSS.n4805 DVSS.n4804 6.3005
R11617 DVSS.n4184 DVSS.n4183 6.3005
R11618 DVSS.n1975 DVSS.n1974 6.3005
R11619 DVSS.n1830 DVSS.n1829 6.3005
R11620 DVSS.n1266 DVSS.n1265 6.3005
R11621 DVSS.n1346 DVSS.n1345 6.3005
R11622 DVSS.n3522 DVSS.n963 6.17435
R11623 DVSS.n5094 DVSS.n5093 6.17435
R11624 DVSS.n4769 DVSS.n4768 5.42247
R11625 VSS DVSS.n4833 5.2005
R11626 VSS DVSS.n4832 5.2005
R11627 VSS DVSS.n4845 5.2005
R11628 VSS DVSS.n4844 5.2005
R11629 VSS DVSS.n4866 5.2005
R11630 VSS DVSS.n4865 5.2005
R11631 DVSS.n1822 DVSS.n1801 5.2005
R11632 DVSS.n3820 DVSS.n1822 5.2005
R11633 DVSS.n3821 DVSS.n1801 5.2005
R11634 DVSS.n3821 DVSS.n1804 5.2005
R11635 DVSS.n3821 DVSS.n1800 5.2005
R11636 DVSS.n3821 DVSS.n1806 5.2005
R11637 DVSS.n3821 DVSS.n1799 5.2005
R11638 DVSS.n3821 DVSS.n1808 5.2005
R11639 DVSS.n3821 DVSS.n1798 5.2005
R11640 DVSS.n3821 DVSS.n1810 5.2005
R11641 DVSS.n3821 DVSS.n1797 5.2005
R11642 DVSS.n3821 DVSS.n1812 5.2005
R11643 DVSS.n3821 DVSS.n1796 5.2005
R11644 DVSS.n3821 DVSS.n3820 5.2005
R11645 DVSS.n1815 DVSS.n1801 5.2005
R11646 DVSS.n1815 DVSS.n1804 5.2005
R11647 DVSS.n1815 DVSS.n1800 5.2005
R11648 DVSS.n1815 DVSS.n1806 5.2005
R11649 DVSS.n1815 DVSS.n1799 5.2005
R11650 DVSS.n1815 DVSS.n1808 5.2005
R11651 DVSS.n1815 DVSS.n1798 5.2005
R11652 DVSS.n1815 DVSS.n1810 5.2005
R11653 DVSS.n1815 DVSS.n1797 5.2005
R11654 DVSS.n1815 DVSS.n1812 5.2005
R11655 DVSS.n3820 DVSS.n1815 5.2005
R11656 DVSS.n1824 DVSS.n1801 5.2005
R11657 DVSS.n1824 DVSS.n1804 5.2005
R11658 DVSS.n1824 DVSS.n1800 5.2005
R11659 DVSS.n1824 DVSS.n1806 5.2005
R11660 DVSS.n1824 DVSS.n1799 5.2005
R11661 DVSS.n1824 DVSS.n1808 5.2005
R11662 DVSS.n1824 DVSS.n1798 5.2005
R11663 DVSS.n1824 DVSS.n1810 5.2005
R11664 DVSS.n1824 DVSS.n1797 5.2005
R11665 DVSS.n1824 DVSS.n1812 5.2005
R11666 DVSS.n3820 DVSS.n1824 5.2005
R11667 DVSS.n1814 DVSS.n1801 5.2005
R11668 DVSS.n1814 DVSS.n1804 5.2005
R11669 DVSS.n1814 DVSS.n1800 5.2005
R11670 DVSS.n1814 DVSS.n1806 5.2005
R11671 DVSS.n1814 DVSS.n1799 5.2005
R11672 DVSS.n1814 DVSS.n1808 5.2005
R11673 DVSS.n1814 DVSS.n1798 5.2005
R11674 DVSS.n1814 DVSS.n1810 5.2005
R11675 DVSS.n1814 DVSS.n1797 5.2005
R11676 DVSS.n1814 DVSS.n1812 5.2005
R11677 DVSS.n3820 DVSS.n1814 5.2005
R11678 DVSS.n1826 DVSS.n1801 5.2005
R11679 DVSS.n1826 DVSS.n1804 5.2005
R11680 DVSS.n1826 DVSS.n1800 5.2005
R11681 DVSS.n1826 DVSS.n1806 5.2005
R11682 DVSS.n1826 DVSS.n1799 5.2005
R11683 DVSS.n1826 DVSS.n1808 5.2005
R11684 DVSS.n1826 DVSS.n1798 5.2005
R11685 DVSS.n1826 DVSS.n1810 5.2005
R11686 DVSS.n1826 DVSS.n1797 5.2005
R11687 DVSS.n1826 DVSS.n1812 5.2005
R11688 DVSS.n3820 DVSS.n1826 5.2005
R11689 DVSS.n1813 DVSS.n1801 5.2005
R11690 DVSS.n1813 DVSS.n1804 5.2005
R11691 DVSS.n1813 DVSS.n1800 5.2005
R11692 DVSS.n1813 DVSS.n1806 5.2005
R11693 DVSS.n1813 DVSS.n1799 5.2005
R11694 DVSS.n1813 DVSS.n1808 5.2005
R11695 DVSS.n1813 DVSS.n1798 5.2005
R11696 DVSS.n1813 DVSS.n1810 5.2005
R11697 DVSS.n1813 DVSS.n1797 5.2005
R11698 DVSS.n1813 DVSS.n1812 5.2005
R11699 DVSS.n3820 DVSS.n1813 5.2005
R11700 DVSS.n3819 DVSS.n1804 5.2005
R11701 DVSS.n3819 DVSS.n1800 5.2005
R11702 DVSS.n3819 DVSS.n1806 5.2005
R11703 DVSS.n3819 DVSS.n1799 5.2005
R11704 DVSS.n3819 DVSS.n1808 5.2005
R11705 DVSS.n3819 DVSS.n1798 5.2005
R11706 DVSS.n3819 DVSS.n1810 5.2005
R11707 DVSS.n3819 DVSS.n1797 5.2005
R11708 DVSS.n3819 DVSS.n1812 5.2005
R11709 DVSS.n3820 DVSS.n3819 5.2005
R11710 DVSS.n2016 DVSS.n1972 5.08553
R11711 DVSS.n3805 DVSS.n1795 4.84618
R11712 DVSS.n1815 DVSS.n1802 4.84618
R11713 DVSS.n1824 DVSS.n1823 4.84618
R11714 DVSS.n3804 DVSS.n1814 4.84618
R11715 DVSS.n1826 DVSS.n1825 4.84618
R11716 DVSS.n3803 DVSS.n1813 4.84618
R11717 DVSS.n3819 DVSS.n1844 4.84618
R11718 DVSS.n3805 DVSS.n1822 4.84618
R11719 DVSS.n3821 DVSS.n1802 4.84618
R11720 DVSS.n1823 DVSS.n1815 4.84618
R11721 DVSS.n3804 DVSS.n1824 4.84618
R11722 DVSS.n1825 DVSS.n1814 4.84618
R11723 DVSS.n3803 DVSS.n1826 4.84618
R11724 DVSS.n1844 DVSS.n1813 4.84618
R11725 DVSS.n4115 DVSS.n1098 4.82802
R11726 DVSS.n5045 DVSS.n5044 4.66866
R11727 DVSS.n1127 DVSS.n1121 4.66866
R11728 DVSS.n3784 DVSS.n3783 4.58103
R11729 DVSS.n4653 DVSS.n4652 4.5005
R11730 DVSS.n4652 DVSS.n4644 4.5005
R11731 DVSS.n4652 DVSS.n4642 4.5005
R11732 DVSS.n4651 DVSS.n4646 4.5005
R11733 DVSS.n4652 DVSS.n4651 4.5005
R11734 DVSS.n4704 DVSS.n4639 4.5005
R11735 DVSS.n4662 DVSS.n4639 4.5005
R11736 DVSS.n4707 DVSS.n4639 4.5005
R11737 DVSS.n4704 DVSS.n4654 4.5005
R11738 DVSS.n4707 DVSS.n4654 4.5005
R11739 DVSS.n4707 DVSS.n4638 4.5005
R11740 DVSS.n4707 DVSS.n4655 4.5005
R11741 DVSS.n4707 DVSS.n4637 4.5005
R11742 DVSS.n4707 DVSS.n4656 4.5005
R11743 DVSS.n4707 DVSS.n4636 4.5005
R11744 DVSS.n4707 DVSS.n4657 4.5005
R11745 DVSS.n4707 DVSS.n4635 4.5005
R11746 DVSS.n4706 DVSS.n4662 4.5005
R11747 DVSS.n4707 DVSS.n4706 4.5005
R11748 DVSS.n4371 DVSS.n4341 4.5005
R11749 DVSS.n4376 DVSS.n4371 4.5005
R11750 DVSS.n4371 DVSS.n4343 4.5005
R11751 DVSS.n4359 DVSS.n4341 4.5005
R11752 DVSS.n4359 DVSS.n4343 4.5005
R11753 DVSS.n4355 DVSS.n4343 4.5005
R11754 DVSS.n4353 DVSS.n4343 4.5005
R11755 DVSS.n4351 DVSS.n4343 4.5005
R11756 DVSS.n4349 DVSS.n4343 4.5005
R11757 DVSS.n4347 DVSS.n4343 4.5005
R11758 DVSS.n4345 DVSS.n4343 4.5005
R11759 DVSS.n4373 DVSS.n4343 4.5005
R11760 DVSS.n4376 DVSS.n4375 4.5005
R11761 DVSS.n4375 DVSS.n4343 4.5005
R11762 DVSS.n4370 DVSS.n4369 4.5005
R11763 DVSS.n4369 DVSS.n4357 4.5005
R11764 DVSS.n4367 DVSS.n4357 4.5005
R11765 DVSS.n4367 DVSS.n4366 4.5005
R11766 DVSS.n4367 DVSS.n4364 4.5005
R11767 DVSS.n4369 DVSS.n4368 4.5005
R11768 DVSS.n4368 DVSS.n4367 4.5005
R11769 DVSS.n2252 DVSS.n2251 4.5005
R11770 DVSS.n1954 DVSS.n1539 4.5005
R11771 DVSS.n2253 DVSS.n2252 4.5005
R11772 DVSS.n2253 DVSS.n1951 4.5005
R11773 DVSS.n2253 DVSS.n1539 4.5005
R11774 DVSS.n4155 DVSS.n1533 4.5005
R11775 DVSS.n1533 DVSS.n1527 4.5005
R11776 DVSS.n1533 DVSS.n1528 4.5005
R11777 DVSS.n4155 DVSS.n1535 4.5005
R11778 DVSS.n1535 DVSS.n1527 4.5005
R11779 DVSS.n1535 DVSS.n1528 4.5005
R11780 DVSS.n1532 DVSS.n1528 4.5005
R11781 DVSS.n1532 DVSS.n1527 4.5005
R11782 DVSS.n4155 DVSS.n1532 4.5005
R11783 DVSS.n1536 DVSS.n1528 4.5005
R11784 DVSS.n1536 DVSS.n1527 4.5005
R11785 DVSS.n4155 DVSS.n1536 4.5005
R11786 DVSS.n4155 DVSS.n1531 4.5005
R11787 DVSS.n1531 DVSS.n1527 4.5005
R11788 DVSS.n1531 DVSS.n1528 4.5005
R11789 DVSS.n4156 DVSS.n1528 4.5005
R11790 DVSS.n4156 DVSS.n1527 4.5005
R11791 DVSS.n4156 DVSS.n4155 4.5005
R11792 DVSS.n4155 DVSS.n1530 4.5005
R11793 DVSS.n1530 DVSS.n1527 4.5005
R11794 DVSS.n1530 DVSS.n1528 4.5005
R11795 DVSS.n4154 DVSS.n1528 4.5005
R11796 DVSS.n4154 DVSS.n1527 4.5005
R11797 DVSS.n4155 DVSS.n4154 4.5005
R11798 DVSS.n2249 DVSS.n1952 4.5005
R11799 DVSS.n1957 DVSS.n1952 4.5005
R11800 DVSS.n1959 DVSS.n1952 4.5005
R11801 DVSS.n2249 DVSS.n1955 4.5005
R11802 DVSS.n1957 DVSS.n1955 4.5005
R11803 DVSS.n1959 DVSS.n1955 4.5005
R11804 DVSS.n2250 DVSS.n1959 4.5005
R11805 DVSS.n2250 DVSS.n1957 4.5005
R11806 DVSS.n2250 DVSS.n2249 4.5005
R11807 DVSS.n2249 DVSS.n2227 4.5005
R11808 DVSS.n2227 DVSS.n1957 4.5005
R11809 DVSS.n2227 DVSS.n1959 4.5005
R11810 DVSS.n2249 DVSS.n1963 4.5005
R11811 DVSS.n1963 DVSS.n1957 4.5005
R11812 DVSS.n1963 DVSS.n1959 4.5005
R11813 DVSS.n2228 DVSS.n1959 4.5005
R11814 DVSS.n2228 DVSS.n1957 4.5005
R11815 DVSS.n2249 DVSS.n2228 4.5005
R11816 DVSS.n1962 DVSS.n1959 4.5005
R11817 DVSS.n1962 DVSS.n1957 4.5005
R11818 DVSS.n2249 DVSS.n1962 4.5005
R11819 DVSS.n2249 DVSS.n2229 4.5005
R11820 DVSS.n2229 DVSS.n1957 4.5005
R11821 DVSS.n2229 DVSS.n1959 4.5005
R11822 DVSS.n1961 DVSS.n1959 4.5005
R11823 DVSS.n1961 DVSS.n1957 4.5005
R11824 DVSS.n2249 DVSS.n1961 4.5005
R11825 DVSS.n2248 DVSS.n1959 4.5005
R11826 DVSS.n2248 DVSS.n1957 4.5005
R11827 DVSS.n2249 DVSS.n2248 4.5005
R11828 DVSS.n2557 DVSS.n1911 4.5005
R11829 DVSS.n1914 DVSS.n1911 4.5005
R11830 DVSS.n2556 DVSS.n1914 4.5005
R11831 DVSS.n2557 DVSS.n2556 4.5005
R11832 DVSS.n2533 DVSS.n1912 4.5005
R11833 DVSS.n2537 DVSS.n1912 4.5005
R11834 DVSS.n1932 DVSS.n1859 4.5005
R11835 DVSS.n1946 DVSS.n1855 4.5005
R11836 DVSS.n1946 DVSS.n1859 4.5005
R11837 DVSS.n1934 DVSS.n1855 4.5005
R11838 DVSS.n1934 DVSS.n1859 4.5005
R11839 DVSS.n1932 DVSS.n1855 4.5005
R11840 DVSS.n2306 DVSS.n1855 4.5005
R11841 DVSS.n2306 DVSS.n1859 4.5005
R11842 DVSS.n2567 DVSS.n1902 4.5005
R11843 DVSS.n2567 DVSS.n2566 4.5005
R11844 DVSS.n2566 DVSS.n2565 4.5005
R11845 DVSS.n2565 DVSS.n1902 4.5005
R11846 DVSS.n2264 DVSS.n1903 4.5005
R11847 DVSS.n2265 DVSS.n2264 4.5005
R11848 DVSS.n2368 DVSS.n2346 4.5005
R11849 DVSS.n2347 DVSS.n2346 4.5005
R11850 DVSS.n2348 DVSS.n2346 4.5005
R11851 DVSS.n2370 DVSS.n2346 4.5005
R11852 DVSS.n2370 DVSS.n2369 4.5005
R11853 DVSS.n2369 DVSS.n2348 4.5005
R11854 DVSS.n2369 DVSS.n2347 4.5005
R11855 DVSS.n2369 DVSS.n2368 4.5005
R11856 DVSS.n2364 DVSS.n2352 4.5005
R11857 DVSS.n2367 DVSS.n2352 4.5005
R11858 DVSS.n2367 DVSS.n2366 4.5005
R11859 DVSS.n2367 DVSS.n2351 4.5005
R11860 DVSS.n2364 DVSS.n1927 4.5005
R11861 DVSS.n2367 DVSS.n1927 4.5005
R11862 DVSS.n2488 DVSS.n1924 4.5005
R11863 DVSS.n2488 DVSS.n1925 4.5005
R11864 DVSS.n2545 DVSS.n1924 4.5005
R11865 DVSS.n2545 DVSS.n1925 4.5005
R11866 DVSS.n2494 DVSS.n1925 4.5005
R11867 DVSS.n2494 DVSS.n1924 4.5005
R11868 DVSS.n2503 DVSS.n2473 4.5005
R11869 DVSS.n2475 DVSS.n2473 4.5005
R11870 DVSS.n2502 DVSS.n2475 4.5005
R11871 DVSS.n2503 DVSS.n2502 4.5005
R11872 DVSS.n2492 DVSS.n1925 4.5005
R11873 DVSS.n2492 DVSS.n1924 4.5005
R11874 DVSS.n2546 DVSS.n2545 4.5005
R11875 DVSS.n2307 DVSS.n2306 4.5005
R11876 DVSS.n2306 DVSS.n2305 4.5005
R11877 DVSS.n2545 DVSS.n2544 4.5005
R11878 DVSS.n2499 DVSS.n2476 4.5005
R11879 DVSS.n2500 DVSS.n2499 4.5005
R11880 DVSS.n2330 DVSS.n2328 4.5005
R11881 DVSS.n2336 DVSS.n2330 4.5005
R11882 DVSS.n2501 DVSS.n2476 4.5005
R11883 DVSS.n2501 DVSS.n2500 4.5005
R11884 DVSS.n2553 DVSS.n1917 4.5005
R11885 DVSS.n2553 DVSS.n2552 4.5005
R11886 DVSS.n2568 DVSS.n1901 4.5005
R11887 DVSS.n2568 DVSS.n1898 4.5005
R11888 DVSS.n1869 DVSS.n1866 4.5005
R11889 DVSS.n1889 DVSS.n1869 4.5005
R11890 DVSS.n2585 DVSS.n1874 4.5005
R11891 DVSS.n2585 DVSS.n1876 4.5005
R11892 DVSS.n2585 DVSS.n1873 4.5005
R11893 DVSS.n2585 DVSS.n2584 4.5005
R11894 DVSS.n2584 DVSS.n2583 4.5005
R11895 DVSS.n2583 DVSS.n1873 4.5005
R11896 DVSS.n2583 DVSS.n1876 4.5005
R11897 DVSS.n2583 DVSS.n1874 4.5005
R11898 DVSS.n2269 DVSS.n1875 4.5005
R11899 DVSS.n2300 DVSS.n1875 4.5005
R11900 DVSS.n2300 DVSS.n2299 4.5005
R11901 DVSS.n2300 DVSS.n2270 4.5005
R11902 DVSS.n2301 DVSS.n2269 4.5005
R11903 DVSS.n2301 DVSS.n2300 4.5005
R11904 DVSS.n2594 DVSS.n1864 4.5005
R11905 DVSS.n2590 DVSS.n1864 4.5005
R11906 DVSS.n2286 DVSS.n2276 4.5005
R11907 DVSS.n2278 DVSS.n2276 4.5005
R11908 DVSS.n2288 DVSS.n2276 4.5005
R11909 DVSS.n2288 DVSS.n2287 4.5005
R11910 DVSS.n2287 DVSS.n2278 4.5005
R11911 DVSS.n2287 DVSS.n2286 4.5005
R11912 DVSS.n2277 DVSS.n1657 4.5005
R11913 DVSS.n2277 DVSS.n1662 4.5005
R11914 DVSS.n1668 DVSS.n1657 4.5005
R11915 DVSS.n3994 DVSS.n1666 4.5005
R11916 DVSS.n3994 DVSS.n3985 4.5005
R11917 DVSS.n3994 DVSS.n1665 4.5005
R11918 DVSS.n3994 DVSS.n3988 4.5005
R11919 DVSS.n3994 DVSS.n1664 4.5005
R11920 DVSS.n3994 DVSS.n3991 4.5005
R11921 DVSS.n3994 DVSS.n1663 4.5005
R11922 DVSS.n3993 DVSS.n1662 4.5005
R11923 DVSS.n3994 DVSS.n3993 4.5005
R11924 DVSS.n4834 VSS 4.5005
R11925 DVSS.n4846 VSS 4.5005
R11926 DVSS.n1122 DVSS.n1121 4.5005
R11927 DVSS.n5033 DVSS.n5032 4.5005
R11928 DVSS.n5035 DVSS.n5034 4.5005
R11929 DVSS.n1119 DVSS.n1117 4.5005
R11930 DVSS.n1110 DVSS.n1109 4.5005
R11931 DVSS.n5044 DVSS.n5043 4.5005
R11932 DVSS.n4885 DVSS.n1196 4.5005
R11933 DVSS.n1196 DVSS.n1193 4.5005
R11934 DVSS.n4885 DVSS.n4874 4.5005
R11935 DVSS.n4888 DVSS.n1198 4.5005
R11936 DVSS.n4888 DVSS.n1201 4.5005
R11937 DVSS.n4888 DVSS.n1197 4.5005
R11938 DVSS.n4888 DVSS.n4874 4.5005
R11939 DVSS.n4888 DVSS.n1196 4.5005
R11940 DVSS.n4882 DVSS.n1193 4.5005
R11941 DVSS.n4880 DVSS.n1193 4.5005
R11942 DVSS.n4879 DVSS.n1193 4.5005
R11943 DVSS.n4877 DVSS.n1193 4.5005
R11944 DVSS.n4888 DVSS.n4887 4.5005
R11945 DVSS.n4887 DVSS.n1193 4.5005
R11946 DVSS.n4867 VSS 4.5005
R11947 DVSS.n3761 DVSS.n3528 4.5005
R11948 DVSS.n3759 DVSS.n3528 4.5005
R11949 DVSS.n3759 DVSS.n3750 4.5005
R11950 DVSS.n3759 DVSS.n3538 4.5005
R11951 DVSS.n3759 DVSS.n3751 4.5005
R11952 DVSS.n3759 DVSS.n3537 4.5005
R11953 DVSS.n3759 DVSS.n3752 4.5005
R11954 DVSS.n3759 DVSS.n3536 4.5005
R11955 DVSS.n3759 DVSS.n3758 4.5005
R11956 DVSS.n3759 DVSS.n3535 4.5005
R11957 DVSS.n3761 DVSS.n3760 4.5005
R11958 DVSS.n3760 DVSS.n3759 4.5005
R11959 DVSS.n4770 DVSS.n1362 4.5005
R11960 DVSS.n1362 DVSS.n1354 4.5005
R11961 DVSS.n1362 DVSS.n1355 4.5005
R11962 DVSS.n1362 DVSS.n1357 4.5005
R11963 DVSS.n1359 DVSS.n1355 4.5005
R11964 DVSS.n1359 DVSS.n1357 4.5005
R11965 DVSS.n4770 DVSS.n1363 4.5005
R11966 DVSS.n1363 DVSS.n1354 4.5005
R11967 DVSS.n1363 DVSS.n1355 4.5005
R11968 DVSS.n1363 DVSS.n1357 4.5005
R11969 DVSS.n4770 DVSS.n1361 4.5005
R11970 DVSS.n1361 DVSS.n1354 4.5005
R11971 DVSS.n1361 DVSS.n1355 4.5005
R11972 DVSS.n1361 DVSS.n1357 4.5005
R11973 DVSS.n1366 DVSS.n1355 4.5005
R11974 DVSS.n1366 DVSS.n1357 4.5005
R11975 DVSS.n1360 DVSS.n1355 4.5005
R11976 DVSS.n1360 DVSS.n1357 4.5005
R11977 DVSS.n4770 DVSS.n1364 4.5005
R11978 DVSS.n1364 DVSS.n1354 4.5005
R11979 DVSS.n1364 DVSS.n1355 4.5005
R11980 DVSS.n1364 DVSS.n1357 4.5005
R11981 DVSS.n1365 DVSS.n1355 4.5005
R11982 DVSS.n1365 DVSS.n1357 4.5005
R11983 DVSS.n4771 DVSS.n1355 4.5005
R11984 DVSS.n4771 DVSS.n1357 4.5005
R11985 DVSS.n4771 DVSS.n1354 4.5005
R11986 DVSS.n4771 DVSS.n4770 4.5005
R11987 DVSS.n1365 DVSS.n1354 4.5005
R11988 DVSS.n4770 DVSS.n1365 4.5005
R11989 DVSS.n1360 DVSS.n1354 4.5005
R11990 DVSS.n4770 DVSS.n1360 4.5005
R11991 DVSS.n1366 DVSS.n1354 4.5005
R11992 DVSS.n4770 DVSS.n1366 4.5005
R11993 DVSS.n1359 DVSS.n1354 4.5005
R11994 DVSS.n4770 DVSS.n1359 4.5005
R11995 DVSS.n4769 DVSS.n1357 4.5005
R11996 DVSS.n4769 DVSS.n1355 4.5005
R11997 DVSS.n4769 DVSS.n1354 4.5005
R11998 DVSS.n4770 DVSS.n4769 4.5005
R11999 DVSS.n5538 DVSS.n5537 4.5005
R12000 DVSS.n4768 DVSS.n855 4.5005
R12001 DVSS.n5541 DVSS.n6 4.5005
R12002 DVSS.n5796 DVSS.n5795 4.5005
R12003 DVSS.n5539 DVSS.n829 4.5005
R12004 DVSS.n5544 DVSS.n5543 4.5005
R12005 DVSS.n3528 DVSS.n2636 4.24863
R12006 DVSS.n1827 DVSS.t151 4.10856
R12007 DVSS.n1828 DVSS.t105 4.10856
R12008 DVSS.n5098 DVSS.n1080 4.05657
R12009 DVSS.n5102 DVSS.n1080 4.05657
R12010 DVSS.n5102 DVSS.n1078 4.05657
R12011 DVSS.n5106 DVSS.n1078 4.05657
R12012 DVSS.n5106 DVSS.n1076 4.05657
R12013 DVSS.n5110 DVSS.n1076 4.05657
R12014 DVSS.n5110 DVSS.n1074 4.05657
R12015 DVSS.n5114 DVSS.n1074 4.05657
R12016 DVSS.n5114 DVSS.n1072 4.05657
R12017 DVSS.n5118 DVSS.n1072 4.05657
R12018 DVSS.n5118 DVSS.n1070 4.05657
R12019 DVSS.n5122 DVSS.n1070 4.05657
R12020 DVSS.n5122 DVSS.n1068 4.05657
R12021 DVSS.n5126 DVSS.n1068 4.05657
R12022 DVSS.n5126 DVSS.n1066 4.05657
R12023 DVSS.n5130 DVSS.n1066 4.05657
R12024 DVSS.n5130 DVSS.n1064 4.05657
R12025 DVSS.n5134 DVSS.n1064 4.05657
R12026 DVSS.n5134 DVSS.n1062 4.05657
R12027 DVSS.n5138 DVSS.n1062 4.05657
R12028 DVSS.n5138 DVSS.n1060 4.05657
R12029 DVSS.n5142 DVSS.n1060 4.05657
R12030 DVSS.n5142 DVSS.n1058 4.05657
R12031 DVSS.n5146 DVSS.n1058 4.05657
R12032 DVSS.n5146 DVSS.n1056 4.05657
R12033 DVSS.n5150 DVSS.n1056 4.05657
R12034 DVSS.n5150 DVSS.n1054 4.05657
R12035 DVSS.n5154 DVSS.n1054 4.05657
R12036 DVSS.n5154 DVSS.n1052 4.05657
R12037 DVSS.n5158 DVSS.n1052 4.05657
R12038 DVSS.n5158 DVSS.n1050 4.05657
R12039 DVSS.n5162 DVSS.n1050 4.05657
R12040 DVSS.n5162 DVSS.n1048 4.05657
R12041 DVSS.n5166 DVSS.n1048 4.05657
R12042 DVSS.n5166 DVSS.n1046 4.05657
R12043 DVSS.n5170 DVSS.n1046 4.05657
R12044 DVSS.n5170 DVSS.n1044 4.05657
R12045 DVSS.n5174 DVSS.n1044 4.05657
R12046 DVSS.n5174 DVSS.n1042 4.05657
R12047 DVSS.n5178 DVSS.n1042 4.05657
R12048 DVSS.n5178 DVSS.n1040 4.05657
R12049 DVSS.n5182 DVSS.n1040 4.05657
R12050 DVSS.n5182 DVSS.n1038 4.05657
R12051 DVSS.n5186 DVSS.n1038 4.05657
R12052 DVSS.n5186 DVSS.n1036 4.05657
R12053 DVSS.n5190 DVSS.n1036 4.05657
R12054 DVSS.n5190 DVSS.n1034 4.05657
R12055 DVSS.n5194 DVSS.n1034 4.05657
R12056 DVSS.n5194 DVSS.n1032 4.05657
R12057 DVSS.n5198 DVSS.n1032 4.05657
R12058 DVSS.n5198 DVSS.n1030 4.05657
R12059 DVSS.n5202 DVSS.n1030 4.05657
R12060 DVSS.n5202 DVSS.n1028 4.05657
R12061 DVSS.n5207 DVSS.n1028 4.05657
R12062 DVSS.n5207 DVSS.n1026 4.05657
R12063 DVSS.n5211 DVSS.n1026 4.05657
R12064 DVSS.n5212 DVSS.n5211 4.05657
R12065 DVSS.n5212 DVSS.n1021 4.05657
R12066 DVSS.n5219 DVSS.n1021 4.05657
R12067 DVSS.n5219 DVSS.n1019 4.05657
R12068 DVSS.n5223 DVSS.n1019 4.05657
R12069 DVSS.n5223 DVSS.n1017 4.05657
R12070 DVSS.n5227 DVSS.n1017 4.05657
R12071 DVSS.n5227 DVSS.n1015 4.05657
R12072 DVSS.n5231 DVSS.n1015 4.05657
R12073 DVSS.n5231 DVSS.n1013 4.05657
R12074 DVSS.n5235 DVSS.n1013 4.05657
R12075 DVSS.n5235 DVSS.n1011 4.05657
R12076 DVSS.n5239 DVSS.n1011 4.05657
R12077 DVSS.n5239 DVSS.n1009 4.05657
R12078 DVSS.n5243 DVSS.n1009 4.05657
R12079 DVSS.n5243 DVSS.n1007 4.05657
R12080 DVSS.n5247 DVSS.n1007 4.05657
R12081 DVSS.n5247 DVSS.n1005 4.05657
R12082 DVSS.n5251 DVSS.n1005 4.05657
R12083 DVSS.n5251 DVSS.n1003 4.05657
R12084 DVSS.n5255 DVSS.n1003 4.05657
R12085 DVSS.n5255 DVSS.n1001 4.05657
R12086 DVSS.n5259 DVSS.n1001 4.05657
R12087 DVSS.n5259 DVSS.n999 4.05657
R12088 DVSS.n5263 DVSS.n999 4.05657
R12089 DVSS.n5263 DVSS.n997 4.05657
R12090 DVSS.n5267 DVSS.n997 4.05657
R12091 DVSS.n5267 DVSS.n995 4.05657
R12092 DVSS.n5271 DVSS.n995 4.05657
R12093 DVSS.n5271 DVSS.n993 4.05657
R12094 DVSS.n5275 DVSS.n993 4.05657
R12095 DVSS.n5275 DVSS.n991 4.05657
R12096 DVSS.n5279 DVSS.n991 4.05657
R12097 DVSS.n5279 DVSS.n989 4.05657
R12098 DVSS.n5283 DVSS.n989 4.05657
R12099 DVSS.n5283 DVSS.n987 4.05657
R12100 DVSS.n5287 DVSS.n987 4.05657
R12101 DVSS.n5287 DVSS.n985 4.05657
R12102 DVSS.n5291 DVSS.n985 4.05657
R12103 DVSS.n5291 DVSS.n983 4.05657
R12104 DVSS.n5295 DVSS.n983 4.05657
R12105 DVSS.n5295 DVSS.n981 4.05657
R12106 DVSS.n5299 DVSS.n981 4.05657
R12107 DVSS.n5299 DVSS.n979 4.05657
R12108 DVSS.n5303 DVSS.n979 4.05657
R12109 DVSS.n5303 DVSS.n977 4.05657
R12110 DVSS.n5307 DVSS.n977 4.05657
R12111 DVSS.n5307 DVSS.n975 4.05657
R12112 DVSS.n5311 DVSS.n975 4.05657
R12113 DVSS.n5311 DVSS.n973 4.05657
R12114 DVSS.n5315 DVSS.n973 4.05657
R12115 DVSS.n5315 DVSS.n971 4.05657
R12116 DVSS.n5319 DVSS.n971 4.05657
R12117 DVSS.n5319 DVSS.n969 4.05657
R12118 DVSS.n5323 DVSS.n969 4.05657
R12119 DVSS.n5323 DVSS.n967 4.05657
R12120 DVSS.n5328 DVSS.n967 4.05657
R12121 DVSS.n5328 DVSS.n965 4.05657
R12122 DVSS.n5332 DVSS.n965 4.05657
R12123 DVSS.n5333 DVSS.n5332 4.05657
R12124 DVSS.n3866 DVSS.n3865 3.98035
R12125 DVSS.n4093 DVSS.n4092 3.8345
R12126 DVSS.n2638 DVSS.n2636 3.7805
R12127 DVSS.n3782 DVSS.n2636 3.77031
R12128 DVSS.n4856 DVSS.n1210 3.68022
R12129 DVSS.n3954 DVSS.n1686 3.3741
R12130 DVSS.n1829 DVSS 3.20629
R12131 DVSS.n1847 DVSS 3.18489
R12132 DVSS.n4300 DVSS.t119 3.17811
R12133 DVSS.n4306 DVSS.t45 3.17811
R12134 DVSS.n1685 DVSS.t194 3.17811
R12135 DVSS.n1706 DVSS.t149 3.17811
R12136 DVSS.n1727 DVSS.t88 3.17811
R12137 DVSS.n1701 DVSS.t92 3.17811
R12138 DVSS.n1626 DVSS.t143 3.17811
R12139 DVSS.n4010 DVSS.t170 3.17811
R12140 DVSS.n1615 DVSS.t134 3.17811
R12141 DVSS.n1618 DVSS.t111 3.17811
R12142 DVSS.n4825 DVSS.t146 3.126
R12143 DVSS.n4135 DVSS.n1517 3.02469
R12144 DVSS.n3760 DVSS.n1196 2.95295
R12145 DVSS.n4285 DVSS.n4283 2.90887
R12146 DVSS.n4835 DVSS.n4834 2.81187
R12147 DVSS.n4847 DVSS.n4846 2.81187
R12148 DVSS.n4868 DVSS.n4867 2.81187
R12149 DVSS.n5334 DVSS.n5333 2.6005
R12150 DVSS.n5332 DVSS.n964 2.6005
R12151 DVSS.n5332 DVSS.n5331 2.6005
R12152 DVSS.n5326 DVSS.n965 2.6005
R12153 DVSS.n5330 DVSS.n965 2.6005
R12154 DVSS.n5328 DVSS.n5327 2.6005
R12155 DVSS.n5329 DVSS.n5328 2.6005
R12156 DVSS.n5325 DVSS.n967 2.6005
R12157 DVSS.n967 DVSS.n966 2.6005
R12158 DVSS.n5324 DVSS.n5323 2.6005
R12159 DVSS.n5323 DVSS.n5322 2.6005
R12160 DVSS.n969 DVSS.n968 2.6005
R12161 DVSS.n5321 DVSS.n969 2.6005
R12162 DVSS.n5319 DVSS.n5318 2.6005
R12163 DVSS.n5320 DVSS.n5319 2.6005
R12164 DVSS.n5317 DVSS.n971 2.6005
R12165 DVSS.n971 DVSS.n970 2.6005
R12166 DVSS.n5316 DVSS.n5315 2.6005
R12167 DVSS.n5315 DVSS.n5314 2.6005
R12168 DVSS.n973 DVSS.n972 2.6005
R12169 DVSS.n5313 DVSS.n973 2.6005
R12170 DVSS.n5311 DVSS.n5310 2.6005
R12171 DVSS.n5312 DVSS.n5311 2.6005
R12172 DVSS.n5309 DVSS.n975 2.6005
R12173 DVSS.n975 DVSS.n974 2.6005
R12174 DVSS.n5308 DVSS.n5307 2.6005
R12175 DVSS.n5307 DVSS.n5306 2.6005
R12176 DVSS.n977 DVSS.n976 2.6005
R12177 DVSS.n5305 DVSS.n977 2.6005
R12178 DVSS.n5303 DVSS.n5302 2.6005
R12179 DVSS.n5304 DVSS.n5303 2.6005
R12180 DVSS.n5301 DVSS.n979 2.6005
R12181 DVSS.n979 DVSS.n978 2.6005
R12182 DVSS.n5300 DVSS.n5299 2.6005
R12183 DVSS.n5299 DVSS.n5298 2.6005
R12184 DVSS.n981 DVSS.n980 2.6005
R12185 DVSS.n5297 DVSS.n981 2.6005
R12186 DVSS.n5295 DVSS.n5294 2.6005
R12187 DVSS.n5296 DVSS.n5295 2.6005
R12188 DVSS.n5293 DVSS.n983 2.6005
R12189 DVSS.n983 DVSS.n982 2.6005
R12190 DVSS.n5292 DVSS.n5291 2.6005
R12191 DVSS.n5291 DVSS.n5290 2.6005
R12192 DVSS.n985 DVSS.n984 2.6005
R12193 DVSS.n5289 DVSS.n985 2.6005
R12194 DVSS.n5287 DVSS.n5286 2.6005
R12195 DVSS.n5288 DVSS.n5287 2.6005
R12196 DVSS.n5285 DVSS.n987 2.6005
R12197 DVSS.n987 DVSS.n986 2.6005
R12198 DVSS.n5284 DVSS.n5283 2.6005
R12199 DVSS.n5283 DVSS.n5282 2.6005
R12200 DVSS.n989 DVSS.n988 2.6005
R12201 DVSS.n5281 DVSS.n989 2.6005
R12202 DVSS.n5279 DVSS.n5278 2.6005
R12203 DVSS.n5280 DVSS.n5279 2.6005
R12204 DVSS.n5277 DVSS.n991 2.6005
R12205 DVSS.n991 DVSS.n990 2.6005
R12206 DVSS.n5276 DVSS.n5275 2.6005
R12207 DVSS.n5275 DVSS.n5274 2.6005
R12208 DVSS.n993 DVSS.n992 2.6005
R12209 DVSS.n5273 DVSS.n993 2.6005
R12210 DVSS.n5271 DVSS.n5270 2.6005
R12211 DVSS.n5272 DVSS.n5271 2.6005
R12212 DVSS.n5269 DVSS.n995 2.6005
R12213 DVSS.n995 DVSS.n994 2.6005
R12214 DVSS.n5268 DVSS.n5267 2.6005
R12215 DVSS.n5267 DVSS.n5266 2.6005
R12216 DVSS.n997 DVSS.n996 2.6005
R12217 DVSS.n5265 DVSS.n997 2.6005
R12218 DVSS.n5263 DVSS.n5262 2.6005
R12219 DVSS.n5264 DVSS.n5263 2.6005
R12220 DVSS.n5261 DVSS.n999 2.6005
R12221 DVSS.n999 DVSS.n998 2.6005
R12222 DVSS.n5260 DVSS.n5259 2.6005
R12223 DVSS.n5259 DVSS.n5258 2.6005
R12224 DVSS.n1001 DVSS.n1000 2.6005
R12225 DVSS.n5257 DVSS.n1001 2.6005
R12226 DVSS.n5255 DVSS.n5254 2.6005
R12227 DVSS.n5256 DVSS.n5255 2.6005
R12228 DVSS.n5253 DVSS.n1003 2.6005
R12229 DVSS.n1003 DVSS.n1002 2.6005
R12230 DVSS.n5252 DVSS.n5251 2.6005
R12231 DVSS.n5251 DVSS.n5250 2.6005
R12232 DVSS.n1005 DVSS.n1004 2.6005
R12233 DVSS.n5249 DVSS.n1005 2.6005
R12234 DVSS.n5247 DVSS.n5246 2.6005
R12235 DVSS.n5248 DVSS.n5247 2.6005
R12236 DVSS.n5245 DVSS.n1007 2.6005
R12237 DVSS.n1007 DVSS.n1006 2.6005
R12238 DVSS.n5244 DVSS.n5243 2.6005
R12239 DVSS.n5243 DVSS.n5242 2.6005
R12240 DVSS.n1009 DVSS.n1008 2.6005
R12241 DVSS.n5241 DVSS.n1009 2.6005
R12242 DVSS.n5239 DVSS.n5238 2.6005
R12243 DVSS.n5240 DVSS.n5239 2.6005
R12244 DVSS.n5237 DVSS.n1011 2.6005
R12245 DVSS.n1011 DVSS.n1010 2.6005
R12246 DVSS.n5236 DVSS.n5235 2.6005
R12247 DVSS.n5235 DVSS.n5234 2.6005
R12248 DVSS.n1013 DVSS.n1012 2.6005
R12249 DVSS.n5233 DVSS.n1013 2.6005
R12250 DVSS.n5231 DVSS.n5230 2.6005
R12251 DVSS.n5232 DVSS.n5231 2.6005
R12252 DVSS.n5229 DVSS.n1015 2.6005
R12253 DVSS.n1015 DVSS.n1014 2.6005
R12254 DVSS.n5228 DVSS.n5227 2.6005
R12255 DVSS.n5227 DVSS.n5226 2.6005
R12256 DVSS.n1017 DVSS.n1016 2.6005
R12257 DVSS.n5225 DVSS.n1017 2.6005
R12258 DVSS.n5223 DVSS.n5222 2.6005
R12259 DVSS.n5224 DVSS.n5223 2.6005
R12260 DVSS.n5221 DVSS.n1019 2.6005
R12261 DVSS.n1019 DVSS.n1018 2.6005
R12262 DVSS.n5220 DVSS.n5219 2.6005
R12263 DVSS.n5219 DVSS.n5218 2.6005
R12264 DVSS.n1021 DVSS.n1020 2.6005
R12265 DVSS.n5217 DVSS.n1021 2.6005
R12266 DVSS.n5213 DVSS.n5212 2.6005
R12267 DVSS.n5212 DVSS.n1022 2.6005
R12268 DVSS.n5211 DVSS.n1025 2.6005
R12269 DVSS.n5211 DVSS.n5210 2.6005
R12270 DVSS.n5205 DVSS.n1026 2.6005
R12271 DVSS.n5209 DVSS.n1026 2.6005
R12272 DVSS.n5207 DVSS.n5206 2.6005
R12273 DVSS.n5208 DVSS.n5207 2.6005
R12274 DVSS.n5204 DVSS.n1028 2.6005
R12275 DVSS.n1028 DVSS.n1027 2.6005
R12276 DVSS.n5203 DVSS.n5202 2.6005
R12277 DVSS.n5202 DVSS.n5201 2.6005
R12278 DVSS.n1030 DVSS.n1029 2.6005
R12279 DVSS.n5200 DVSS.n1030 2.6005
R12280 DVSS.n5198 DVSS.n5197 2.6005
R12281 DVSS.n5199 DVSS.n5198 2.6005
R12282 DVSS.n5196 DVSS.n1032 2.6005
R12283 DVSS.n1032 DVSS.n1031 2.6005
R12284 DVSS.n5195 DVSS.n5194 2.6005
R12285 DVSS.n5194 DVSS.n5193 2.6005
R12286 DVSS.n1034 DVSS.n1033 2.6005
R12287 DVSS.n5192 DVSS.n1034 2.6005
R12288 DVSS.n5190 DVSS.n5189 2.6005
R12289 DVSS.n5191 DVSS.n5190 2.6005
R12290 DVSS.n5188 DVSS.n1036 2.6005
R12291 DVSS.n1036 DVSS.n1035 2.6005
R12292 DVSS.n5187 DVSS.n5186 2.6005
R12293 DVSS.n5186 DVSS.n5185 2.6005
R12294 DVSS.n1038 DVSS.n1037 2.6005
R12295 DVSS.n5184 DVSS.n1038 2.6005
R12296 DVSS.n5182 DVSS.n5181 2.6005
R12297 DVSS.n5183 DVSS.n5182 2.6005
R12298 DVSS.n5180 DVSS.n1040 2.6005
R12299 DVSS.n1040 DVSS.n1039 2.6005
R12300 DVSS.n5179 DVSS.n5178 2.6005
R12301 DVSS.n5178 DVSS.n5177 2.6005
R12302 DVSS.n1042 DVSS.n1041 2.6005
R12303 DVSS.n5176 DVSS.n1042 2.6005
R12304 DVSS.n5174 DVSS.n5173 2.6005
R12305 DVSS.n5175 DVSS.n5174 2.6005
R12306 DVSS.n5172 DVSS.n1044 2.6005
R12307 DVSS.n1044 DVSS.n1043 2.6005
R12308 DVSS.n5171 DVSS.n5170 2.6005
R12309 DVSS.n5170 DVSS.n5169 2.6005
R12310 DVSS.n1046 DVSS.n1045 2.6005
R12311 DVSS.n5168 DVSS.n1046 2.6005
R12312 DVSS.n5166 DVSS.n5165 2.6005
R12313 DVSS.n5167 DVSS.n5166 2.6005
R12314 DVSS.n5164 DVSS.n1048 2.6005
R12315 DVSS.n1048 DVSS.n1047 2.6005
R12316 DVSS.n5163 DVSS.n5162 2.6005
R12317 DVSS.n5162 DVSS.n5161 2.6005
R12318 DVSS.n1050 DVSS.n1049 2.6005
R12319 DVSS.n5160 DVSS.n1050 2.6005
R12320 DVSS.n5158 DVSS.n5157 2.6005
R12321 DVSS.n5159 DVSS.n5158 2.6005
R12322 DVSS.n5156 DVSS.n1052 2.6005
R12323 DVSS.n1052 DVSS.n1051 2.6005
R12324 DVSS.n5155 DVSS.n5154 2.6005
R12325 DVSS.n5154 DVSS.n5153 2.6005
R12326 DVSS.n1054 DVSS.n1053 2.6005
R12327 DVSS.n5152 DVSS.n1054 2.6005
R12328 DVSS.n5150 DVSS.n5149 2.6005
R12329 DVSS.n5151 DVSS.n5150 2.6005
R12330 DVSS.n5148 DVSS.n1056 2.6005
R12331 DVSS.n1056 DVSS.n1055 2.6005
R12332 DVSS.n5147 DVSS.n5146 2.6005
R12333 DVSS.n5146 DVSS.n5145 2.6005
R12334 DVSS.n1058 DVSS.n1057 2.6005
R12335 DVSS.n5144 DVSS.n1058 2.6005
R12336 DVSS.n5142 DVSS.n5141 2.6005
R12337 DVSS.n5143 DVSS.n5142 2.6005
R12338 DVSS.n5140 DVSS.n1060 2.6005
R12339 DVSS.n1060 DVSS.n1059 2.6005
R12340 DVSS.n5139 DVSS.n5138 2.6005
R12341 DVSS.n5138 DVSS.n5137 2.6005
R12342 DVSS.n1062 DVSS.n1061 2.6005
R12343 DVSS.n5136 DVSS.n1062 2.6005
R12344 DVSS.n5134 DVSS.n5133 2.6005
R12345 DVSS.n5135 DVSS.n5134 2.6005
R12346 DVSS.n5132 DVSS.n1064 2.6005
R12347 DVSS.n1064 DVSS.n1063 2.6005
R12348 DVSS.n5131 DVSS.n5130 2.6005
R12349 DVSS.n5130 DVSS.n5129 2.6005
R12350 DVSS.n1066 DVSS.n1065 2.6005
R12351 DVSS.n5128 DVSS.n1066 2.6005
R12352 DVSS.n5126 DVSS.n5125 2.6005
R12353 DVSS.n5127 DVSS.n5126 2.6005
R12354 DVSS.n5124 DVSS.n1068 2.6005
R12355 DVSS.n1068 DVSS.n1067 2.6005
R12356 DVSS.n5123 DVSS.n5122 2.6005
R12357 DVSS.n5122 DVSS.n5121 2.6005
R12358 DVSS.n1070 DVSS.n1069 2.6005
R12359 DVSS.n5120 DVSS.n1070 2.6005
R12360 DVSS.n5118 DVSS.n5117 2.6005
R12361 DVSS.n5119 DVSS.n5118 2.6005
R12362 DVSS.n5116 DVSS.n1072 2.6005
R12363 DVSS.n1072 DVSS.n1071 2.6005
R12364 DVSS.n5115 DVSS.n5114 2.6005
R12365 DVSS.n5114 DVSS.n5113 2.6005
R12366 DVSS.n1074 DVSS.n1073 2.6005
R12367 DVSS.n5112 DVSS.n1074 2.6005
R12368 DVSS.n5110 DVSS.n5109 2.6005
R12369 DVSS.n5111 DVSS.n5110 2.6005
R12370 DVSS.n5108 DVSS.n1076 2.6005
R12371 DVSS.n1076 DVSS.n1075 2.6005
R12372 DVSS.n5107 DVSS.n5106 2.6005
R12373 DVSS.n5106 DVSS.n5105 2.6005
R12374 DVSS.n1078 DVSS.n1077 2.6005
R12375 DVSS.n5104 DVSS.n1078 2.6005
R12376 DVSS.n5102 DVSS.n5101 2.6005
R12377 DVSS.n5103 DVSS.n5102 2.6005
R12378 DVSS.n5100 DVSS.n1080 2.6005
R12379 DVSS.n1080 DVSS.n1079 2.6005
R12380 DVSS.n5099 DVSS.n5098 2.6005
R12381 DVSS.n1836 DVSS.n1835 2.49974
R12382 DVSS.n1835 DVSS.n1832 2.49796
R12383 DVSS.n4772 DVSS.n4771 2.43717
R12384 DVSS.n1822 DVSS.n1821 2.41753
R12385 DVSS.n1822 DVSS.n1820 2.41753
R12386 DVSS.n1822 DVSS.n1819 2.41753
R12387 DVSS.n1822 DVSS.n1818 2.41753
R12388 DVSS.n1822 DVSS.n1817 2.41753
R12389 DVSS.n1803 DVSS.n1795 2.41753
R12390 DVSS.n1805 DVSS.n1795 2.41753
R12391 DVSS.n1807 DVSS.n1795 2.41753
R12392 DVSS.n1809 DVSS.n1795 2.41753
R12393 DVSS.n1811 DVSS.n1795 2.41753
R12394 DVSS.n1816 DVSS.n1795 2.41753
R12395 DVSS.n3819 DVSS.n3818 2.41753
R12396 DVSS.n4788 DVSS.n1250 2.41274
R12397 DVSS.n4788 DVSS.n4787 2.41274
R12398 DVSS.n4295 DVSS.n4294 2.41274
R12399 DVSS.n4294 DVSS.n4293 2.41274
R12400 DVSS.n4092 DVSS.n1556 2.311
R12401 DVSS.n1833 DVSS 2.30994
R12402 DVSS.n1831 DVSS 2.30994
R12403 DVSS.t137 DVSS.n2616 2.29246
R12404 DVSS.n1939 DVSS.n1936 2.2728
R12405 DVSS.n4853 DVSS.n4851 2.25682
R12406 DVSS.n4289 DVSS.n4288 2.25682
R12407 DVSS.n4828 DVSS.n4827 2.25682
R12408 DVSS.n4860 DVSS.n4859 2.25682
R12409 DVSS.n4283 DVSS.n1483 2.25392
R12410 DVSS.n1835 DVSS.n1834 2.25346
R12411 DVSS.n2349 DVSS.n2329 2.2505
R12412 DVSS.n2524 DVSS.n2523 2.2505
R12413 DVSS.n2324 DVSS.n2318 2.2505
R12414 DVSS.n2323 DVSS.n2313 2.2505
R12415 DVSS.n1892 DVSS.n1878 2.2505
R12416 DVSS.n2257 DVSS.n1888 2.2505
R12417 DVSS.n2575 DVSS.n2574 2.2505
R12418 DVSS.n1894 DVSS.n1885 2.2505
R12419 DVSS.n2477 DVSS.n2472 2.2505
R12420 DVSS.n2480 DVSS.n2340 2.2505
R12421 DVSS.n2512 DVSS.n2511 2.2505
R12422 DVSS.n2371 DVSS.n2332 2.2505
R12423 DVSS.n2497 DVSS.n2486 2.2505
R12424 DVSS.n2489 DVSS.n1923 2.2505
R12425 DVSS.n2491 DVSS.n2490 2.2505
R12426 DVSS.n2493 DVSS.n2487 2.2505
R12427 DVSS.n2496 DVSS.n2495 2.2505
R12428 DVSS.n1950 DVSS.n1949 2.2505
R12429 DVSS.n1948 DVSS.n1947 2.2505
R12430 DVSS.n1945 DVSS.n1944 2.2505
R12431 DVSS.n1943 DVSS.n1942 2.2505
R12432 DVSS.n1941 DVSS.n1935 2.2505
R12433 DVSS.n2484 DVSS.n2483 2.2505
R12434 DVSS.n2482 DVSS.n2481 2.2505
R12435 DVSS.n2479 DVSS.n2478 2.2505
R12436 DVSS.n2338 DVSS.n2337 2.2505
R12437 DVSS.n2514 DVSS.n2513 2.2505
R12438 DVSS.n2516 DVSS.n2515 2.2505
R12439 DVSS.n2519 DVSS.n2518 2.2505
R12440 DVSS.n2520 DVSS.n2321 2.2505
R12441 DVSS.n2522 DVSS.n2521 2.2505
R12442 DVSS.n2327 DVSS.n2320 2.2505
R12443 DVSS.n2326 DVSS.n2325 2.2505
R12444 DVSS.n2322 DVSS.n1916 2.2505
R12445 DVSS.n2571 DVSS.n2570 2.2505
R12446 DVSS.n2573 DVSS.n2572 2.2505
R12447 DVSS.n1897 DVSS.n1887 2.2505
R12448 DVSS.n1896 DVSS.n1895 2.2505
R12449 DVSS.n1893 DVSS.n1891 2.2505
R12450 DVSS.n1890 DVSS.n1868 2.2505
R12451 DVSS.n2589 DVSS.n2588 2.2505
R12452 DVSS.n1863 DVSS.n1861 2.2505
R12453 DVSS.n2596 DVSS.n2595 2.2505
R12454 DVSS.n2279 DVSS.n1862 2.2505
R12455 DVSS.n2598 DVSS.n2597 2.2505
R12456 DVSS.n1939 DVSS.n1938 2.2505
R12457 DVSS.n4092 DVSS.n4091 2.2505
R12458 DVSS.n294 DVSS.n265 2.2505
R12459 DVSS.n293 DVSS.n292 2.2505
R12460 DVSS.n291 DVSS.n266 2.2505
R12461 DVSS.n290 DVSS.n289 2.2505
R12462 DVSS.n288 DVSS.n267 2.2505
R12463 DVSS.n287 DVSS.n286 2.2505
R12464 DVSS.n285 DVSS.n268 2.2505
R12465 DVSS.n284 DVSS.n283 2.2505
R12466 DVSS.n282 DVSS.n269 2.2505
R12467 DVSS.n281 DVSS.n280 2.2505
R12468 DVSS.n279 DVSS.n270 2.2505
R12469 DVSS.n278 DVSS.n277 2.2505
R12470 DVSS.n274 DVSS.n271 2.2505
R12471 DVSS.n273 DVSS.n272 2.2505
R12472 DVSS.n429 DVSS.n428 2.2505
R12473 DVSS.n430 DVSS.n240 2.2505
R12474 DVSS.n432 DVSS.n431 2.2505
R12475 DVSS.n433 DVSS.n239 2.2505
R12476 DVSS.n435 DVSS.n434 2.2505
R12477 DVSS.n436 DVSS.n238 2.2505
R12478 DVSS.n438 DVSS.n437 2.2505
R12479 DVSS.n439 DVSS.n237 2.2505
R12480 DVSS.n441 DVSS.n440 2.2505
R12481 DVSS.n442 DVSS.n236 2.2505
R12482 DVSS.n444 DVSS.n443 2.2505
R12483 DVSS.n445 DVSS.n235 2.2505
R12484 DVSS.n447 DVSS.n446 2.2505
R12485 DVSS.n448 DVSS.n234 2.2505
R12486 DVSS.n450 DVSS.n449 2.2505
R12487 DVSS.n451 DVSS.n233 2.2505
R12488 DVSS.n453 DVSS.n452 2.2505
R12489 DVSS.n454 DVSS.n232 2.2505
R12490 DVSS.n456 DVSS.n455 2.2505
R12491 DVSS.n457 DVSS.n231 2.2505
R12492 DVSS.n459 DVSS.n458 2.2505
R12493 DVSS.n460 DVSS.n230 2.2505
R12494 DVSS.n462 DVSS.n461 2.2505
R12495 DVSS.n307 DVSS.n261 2.2505
R12496 DVSS.n309 DVSS.n308 2.2505
R12497 DVSS.n306 DVSS.n259 2.2505
R12498 DVSS.n305 DVSS.n304 2.2505
R12499 DVSS.n303 DVSS.n262 2.2505
R12500 DVSS.n302 DVSS.n301 2.2505
R12501 DVSS.n300 DVSS.n263 2.2505
R12502 DVSS.n299 DVSS.n298 2.2505
R12503 DVSS.n297 DVSS.n264 2.2505
R12504 DVSS.n296 DVSS.n295 2.2505
R12505 DVSS.n800 DVSS.n754 2.2505
R12506 DVSS.n799 DVSS.n798 2.2505
R12507 DVSS.n797 DVSS.n755 2.2505
R12508 DVSS.n796 DVSS.n795 2.2505
R12509 DVSS.n794 DVSS.n756 2.2505
R12510 DVSS.n793 DVSS.n792 2.2505
R12511 DVSS.n791 DVSS.n757 2.2505
R12512 DVSS.n790 DVSS.n789 2.2505
R12513 DVSS.n787 DVSS.n786 2.2505
R12514 DVSS.n785 DVSS.n759 2.2505
R12515 DVSS.n784 DVSS.n783 2.2505
R12516 DVSS.n782 DVSS.n760 2.2505
R12517 DVSS.n781 DVSS.n780 2.2505
R12518 DVSS.n779 DVSS.n761 2.2505
R12519 DVSS.n778 DVSS.n777 2.2505
R12520 DVSS.n776 DVSS.n762 2.2505
R12521 DVSS.n775 DVSS.n774 2.2505
R12522 DVSS.n773 DVSS.n763 2.2505
R12523 DVSS.n772 DVSS.n771 2.2505
R12524 DVSS.n770 DVSS.n764 2.2505
R12525 DVSS.n769 DVSS.n768 2.2505
R12526 DVSS.n767 DVSS.n766 2.2505
R12527 DVSS.n5714 DVSS.n5713 2.2505
R12528 DVSS.n5712 DVSS.n56 2.2505
R12529 DVSS.n72 DVSS.n58 2.2505
R12530 DVSS.n74 DVSS.n73 2.2505
R12531 DVSS.n75 DVSS.n71 2.2505
R12532 DVSS.n77 DVSS.n76 2.2505
R12533 DVSS.n78 DVSS.n70 2.2505
R12534 DVSS.n80 DVSS.n79 2.2505
R12535 DVSS.n81 DVSS.n69 2.2505
R12536 DVSS.n83 DVSS.n82 2.2505
R12537 DVSS.n84 DVSS.n68 2.2505
R12538 DVSS.n86 DVSS.n85 2.2505
R12539 DVSS.n87 DVSS.n67 2.2505
R12540 DVSS.n89 DVSS.n88 2.2505
R12541 DVSS.n90 DVSS.n66 2.2505
R12542 DVSS.n92 DVSS.n91 2.2505
R12543 DVSS.n93 DVSS.n65 2.2505
R12544 DVSS.n95 DVSS.n94 2.2505
R12545 DVSS.n96 DVSS.n64 2.2505
R12546 DVSS.n98 DVSS.n97 2.2505
R12547 DVSS.n99 DVSS.n63 2.2505
R12548 DVSS.n101 DVSS.n100 2.2505
R12549 DVSS.n5703 DVSS.n62 2.2505
R12550 DVSS.n5705 DVSS.n5704 2.2505
R12551 DVSS.n788 DVSS.n758 2.2505
R12552 DVSS.n4653 DVSS.n4641 2.24683
R12553 DVSS.n4647 DVSS.n4643 2.24683
R12554 DVSS.n4370 DVSS.n4358 2.24683
R12555 DVSS.n5537 DVSS.n852 2.24648
R12556 DVSS.n5537 DVSS.n851 2.24648
R12557 DVSS.n5537 DVSS.n850 2.24648
R12558 DVSS.n5537 DVSS.n849 2.24648
R12559 DVSS.n855 DVSS.n848 2.24648
R12560 DVSS.n855 DVSS.n853 2.24648
R12561 DVSS.n1368 DVSS.n855 2.24648
R12562 DVSS.n855 DVSS.n854 2.24648
R12563 DVSS.n2251 DVSS.n1956 2.24442
R12564 DVSS.n1954 DVSS.n1953 2.24442
R12565 DVSS.n4649 DVSS.n4648 2.24405
R12566 DVSS.n4646 DVSS.n4645 2.24405
R12567 DVSS.n4650 DVSS.n4649 2.24405
R12568 DVSS.n4365 DVSS.n4361 2.24405
R12569 DVSS.n4369 DVSS.n4362 2.24405
R12570 DVSS.n4363 DVSS.n4361 2.24405
R12571 DVSS.n2365 DVSS.n2364 2.24386
R12572 DVSS.n2363 DVSS.n2362 2.24386
R12573 DVSS.n2362 DVSS.n2361 2.24386
R12574 DVSS.n2298 DVSS.n2269 2.24386
R12575 DVSS.n2297 DVSS.n2296 2.24386
R12576 DVSS.n2296 DVSS.n2268 2.24386
R12577 DVSS.n4704 DVSS.n4666 2.24304
R12578 DVSS.n4662 DVSS.n4661 2.24304
R12579 DVSS.n4704 DVSS.n4665 2.24304
R12580 DVSS.n4662 DVSS.n4660 2.24304
R12581 DVSS.n4704 DVSS.n4664 2.24304
R12582 DVSS.n4662 DVSS.n4659 2.24304
R12583 DVSS.n4705 DVSS.n4704 2.24304
R12584 DVSS.n4662 DVSS.n4658 2.24304
R12585 DVSS.n4376 DVSS.n4356 2.24304
R12586 DVSS.n4354 DVSS.n4341 2.24304
R12587 DVSS.n4376 DVSS.n4352 2.24304
R12588 DVSS.n4350 DVSS.n4341 2.24304
R12589 DVSS.n4376 DVSS.n4348 2.24304
R12590 DVSS.n4346 DVSS.n4341 2.24304
R12591 DVSS.n4376 DVSS.n4344 2.24304
R12592 DVSS.n4374 DVSS.n4341 2.24304
R12593 DVSS.n3994 DVSS.n1669 2.24304
R12594 DVSS.n1667 DVSS.n1662 2.24304
R12595 DVSS.n3984 DVSS.n1657 2.24304
R12596 DVSS.n3983 DVSS.n1662 2.24304
R12597 DVSS.n3987 DVSS.n1657 2.24304
R12598 DVSS.n3986 DVSS.n1662 2.24304
R12599 DVSS.n3990 DVSS.n1657 2.24304
R12600 DVSS.n3989 DVSS.n1662 2.24304
R12601 DVSS.n3992 DVSS.n1657 2.24304
R12602 DVSS.n4873 DVSS.n1193 2.24304
R12603 DVSS.n4885 DVSS.n4884 2.24304
R12604 DVSS.n1200 DVSS.n1193 2.24304
R12605 DVSS.n4888 DVSS.n4875 2.24304
R12606 DVSS.n4885 DVSS.n4883 2.24304
R12607 DVSS.n4888 DVSS.n4876 2.24304
R12608 DVSS.n4885 DVSS.n4881 2.24304
R12609 DVSS.n4886 DVSS.n4885 2.24304
R12610 DVSS.n3761 DVSS.n3529 2.24304
R12611 DVSS.n3756 DVSS.n3753 2.24304
R12612 DVSS.n3761 DVSS.n3530 2.24304
R12613 DVSS.n3756 DVSS.n3754 2.24304
R12614 DVSS.n3761 DVSS.n3531 2.24304
R12615 DVSS.n3756 DVSS.n3755 2.24304
R12616 DVSS.n3761 DVSS.n3532 2.24304
R12617 DVSS.n3757 DVSS.n3756 2.24304
R12618 DVSS.n3756 DVSS.n3533 2.24304
R12619 DVSS.n2335 DVSS.n2331 2.24011
R12620 DVSS.n2333 DVSS.n2331 2.24011
R12621 DVSS.n2586 DVSS.n1872 2.24011
R12622 DVSS.n2586 DVSS.n1870 2.24011
R12623 DVSS.n2591 DVSS.n1865 2.24011
R12624 DVSS.n2593 DVSS.n1865 2.24011
R12625 DVSS.n1900 DVSS.n1899 2.24011
R12626 DVSS.n2555 DVSS.n1915 2.24011
R12627 DVSS.n2334 DVSS.n2330 2.24011
R12628 DVSS.n1871 DVSS.n1869 2.24011
R12629 DVSS.n2592 DVSS.n1864 2.24011
R12630 DVSS.n2534 DVSS.n2532 2.23777
R12631 DVSS.n2535 DVSS.n1912 2.23777
R12632 DVSS.n2536 DVSS.n2532 2.23777
R12633 DVSS.n2262 DVSS.n2261 2.23777
R12634 DVSS.n2264 DVSS.n2263 2.23777
R12635 DVSS.n2261 DVSS.n2256 2.23777
R12636 DVSS.n5796 DVSS.n25 2.23644
R12637 DVSS.n24 DVSS.n6 2.23644
R12638 DVSS.n5796 DVSS.n23 2.23644
R12639 DVSS.n22 DVSS.n6 2.23644
R12640 DVSS.n5796 DVSS.n21 2.23644
R12641 DVSS.n20 DVSS.n6 2.23644
R12642 DVSS.n5796 DVSS.n19 2.23644
R12643 DVSS.n18 DVSS.n6 2.23644
R12644 DVSS.n5796 DVSS.n17 2.23644
R12645 DVSS.n16 DVSS.n6 2.23644
R12646 DVSS.n5796 DVSS.n15 2.23644
R12647 DVSS.n14 DVSS.n6 2.23644
R12648 DVSS.n5796 DVSS.n13 2.23644
R12649 DVSS.n12 DVSS.n6 2.23644
R12650 DVSS.n5796 DVSS.n11 2.23644
R12651 DVSS.n10 DVSS.n6 2.23644
R12652 DVSS.n5796 DVSS.n9 2.23644
R12653 DVSS.n8 DVSS.n6 2.23644
R12654 DVSS.n5796 DVSS.n7 2.23644
R12655 DVSS.n5794 DVSS.n6 2.23644
R12656 DVSS.n5544 DVSS.n5540 2.23644
R12657 DVSS.n847 DVSS.n829 2.23644
R12658 DVSS.n5544 DVSS.n846 2.23644
R12659 DVSS.n845 DVSS.n829 2.23644
R12660 DVSS.n5544 DVSS.n844 2.23644
R12661 DVSS.n843 DVSS.n829 2.23644
R12662 DVSS.n5544 DVSS.n842 2.23644
R12663 DVSS.n841 DVSS.n829 2.23644
R12664 DVSS.n5544 DVSS.n840 2.23644
R12665 DVSS.n839 DVSS.n829 2.23644
R12666 DVSS.n5544 DVSS.n838 2.23644
R12667 DVSS.n837 DVSS.n829 2.23644
R12668 DVSS.n5544 DVSS.n836 2.23644
R12669 DVSS.n835 DVSS.n829 2.23644
R12670 DVSS.n5544 DVSS.n834 2.23644
R12671 DVSS.n833 DVSS.n829 2.23644
R12672 DVSS.n5544 DVSS.n832 2.23644
R12673 DVSS.n831 DVSS.n829 2.23644
R12674 DVSS.n5544 DVSS.n830 2.23644
R12675 DVSS.n5542 DVSS.n829 2.23644
R12676 DVSS.n1834 DVSS.n1833 2.18437
R12677 DVSS.n1832 DVSS.n1831 2.18437
R12678 DVSS.n4117 DVSS.n1545 2.16228
R12679 DVSS.n5339 DVSS.n5338 2.15282
R12680 DVSS.n4059 DVSS.n4058 2.12226
R12681 DVSS.n3944 DVSS.n3940 2.10421
R12682 DVSS.n2629 DVSS.n2628 2.10097
R12683 DVSS.n4302 DVSS.n4301 2.08611
R12684 DVSS.n1699 DVSS.n1698 2.08611
R12685 DVSS.n3942 DVSS.n3941 2.08611
R12686 DVSS.n1613 DVSS.n1612 2.08611
R12687 DVSS.n1621 DVSS.n1620 2.08611
R12688 DVSS.n4175 DVSS.n4174 2.07167
R12689 DVSS.n3794 DVSS.n1686 2.04166
R12690 DVSS.n4170 DVSS.n4169 2.01663
R12691 DVSS.t106 DVSS.n4289 2.01372
R12692 DVSS.n1729 DVSS.n1695 1.96906
R12693 DVSS.n1512 DVSS.n1507 1.94426
R12694 DVSS.n3789 DVSS.n2633 1.94426
R12695 DVSS.n2620 DVSS.n2619 1.91475
R12696 DVSS.n2621 DVSS.n1555 1.91081
R12697 DVSS.n2663 DVSS.n2662 1.89625
R12698 DVSS.n1258 DVSS.n1255 1.81109
R12699 DVSS.n1508 DVSS.n1467 1.81109
R12700 DVSS.n1260 DVSS.n1251 1.81109
R12701 DVSS.n1504 DVSS.n1469 1.81109
R12702 DVSS.n4310 DVSS.n4309 1.80682
R12703 DVSS.n1553 VSS 1.7864
R12704 DVSS.n4096 VSS 1.7864
R12705 DVSS.n1456 DVSS.n1452 1.73383
R12706 DVSS.n4304 DVSS.n1452 1.73383
R12707 DVSS.n1271 DVSS.n1263 1.73383
R12708 DVSS.n4757 DVSS.n1263 1.73383
R12709 DVSS.n1478 DVSS.n1473 1.73383
R12710 DVSS.n1473 DVSS.n1222 1.73383
R12711 DVSS.n4814 DVSS.n4813 1.73383
R12712 DVSS.n4813 DVSS.n4812 1.73383
R12713 DVSS.n5335 DVSS.n5334 1.69628
R12714 DVSS.n5707 DVSS.n5706 1.66284
R12715 DVSS.n4317 DVSS.n4316 1.66212
R12716 DVSS.n5707 DVSS.n60 1.64846
R12717 DVSS.n4835 DVSS.n4831 1.61108
R12718 DVSS.n4848 DVSS.n4847 1.61108
R12719 DVSS.n4869 DVSS.n4868 1.61108
R12720 DVSS.n4103 DVSS.t54 1.5965
R12721 DVSS.n4100 DVSS.t57 1.5965
R12722 DVSS.n4109 DVSS.t52 1.5965
R12723 DVSS.n1552 DVSS.t53 1.5965
R12724 DVSS.n1551 DVSS.t53 1.5965
R12725 DVSS.n1551 DVSS.t57 1.5965
R12726 DVSS.n4101 DVSS.t52 1.5965
R12727 DVSS.n4101 DVSS.t54 1.5965
R12728 DVSS.n4049 DVSS.n4048 1.59033
R12729 DVSS.n4040 DVSS.n1622 1.59033
R12730 DVSS.n4031 DVSS.n1619 1.59033
R12731 DVSS.n1642 DVSS.n1616 1.59033
R12732 DVSS.n1647 DVSS.n1614 1.59033
R12733 DVSS.n4012 DVSS.n4011 1.59033
R12734 DVSS.n3931 DVSS.n3930 1.59033
R12735 DVSS.n1721 DVSS.n1702 1.59033
R12736 DVSS.n1726 DVSS.n1700 1.59033
R12737 DVSS.n3784 DVSS.n2635 1.56129
R12738 DVSS.n4114 DVSS.n1549 1.52301
R12739 DVSS.n3795 DVSS.n3792 1.51243
R12740 DVSS.n4732 DVSS.n4731 1.50734
R12741 DVSS.n4717 DVSS.n4716 1.50734
R12742 DVSS.n4586 DVSS.n4585 1.50734
R12743 DVSS.n4602 DVSS.n4601 1.50734
R12744 DVSS.n1429 DVSS.n1428 1.50734
R12745 DVSS.n4568 DVSS.n4567 1.50734
R12746 DVSS.n4452 DVSS.n4451 1.50734
R12747 DVSS.n4528 DVSS.n4527 1.50734
R12748 DVSS.n4484 DVSS.n4483 1.50734
R12749 DVSS.n4469 DVSS.n4468 1.50734
R12750 DVSS.n4393 DVSS.n4392 1.50734
R12751 DVSS.n4409 DVSS.n4408 1.50734
R12752 DVSS.n2671 DVSS.n2667 1.5055
R12753 DVSS.n3829 DVSS.n3828 1.5055
R12754 DVSS.n3504 DVSS.n2667 1.5055
R12755 DVSS.n3829 DVSS.n1788 1.5055
R12756 DVSS.n1249 DVSS.n1234 1.50326
R12757 DVSS.n4180 DVSS.n4179 1.50326
R12758 DVSS.n2248 DVSS.n2247 1.50157
R12759 DVSS.n4407 DVSS.n4329 1.5005
R12760 DVSS.n4502 DVSS.n4501 1.5005
R12761 DVSS.n4399 DVSS.n4326 1.5005
R12762 DVSS.n4398 DVSS.n4397 1.5005
R12763 DVSS.n4337 DVSS.n4335 1.5005
R12764 DVSS.n4434 DVSS.n4427 1.5005
R12765 DVSS.n4473 DVSS.n4472 1.5005
R12766 DVSS.n4429 DVSS.n4424 1.5005
R12767 DVSS.n4428 DVSS.n4417 1.5005
R12768 DVSS.n4482 DVSS.n4481 1.5005
R12769 DVSS.n1442 DVSS.n1438 1.5005
R12770 DVSS.n4524 DVSS.n4523 1.5005
R12771 DVSS.n4515 DVSS.n4514 1.5005
R12772 DVSS.n1447 DVSS.n1446 1.5005
R12773 DVSS.n4450 DVSS.n4449 1.5005
R12774 DVSS.n1421 DVSS.n1417 1.5005
R12775 DVSS.n4564 DVSS.n4563 1.5005
R12776 DVSS.n4554 DVSS.n4553 1.5005
R12777 DVSS.n1427 DVSS.n1426 1.5005
R12778 DVSS.n4547 DVSS.n4546 1.5005
R12779 DVSS.n4600 DVSS.n1400 1.5005
R12780 DVSS.n4750 DVSS.n4749 1.5005
R12781 DVSS.n4592 DVSS.n1397 1.5005
R12782 DVSS.n4591 DVSS.n4590 1.5005
R12783 DVSS.n1408 DVSS.n1406 1.5005
R12784 DVSS.n4627 DVSS.n4620 1.5005
R12785 DVSS.n4721 DVSS.n4720 1.5005
R12786 DVSS.n4622 DVSS.n4617 1.5005
R12787 DVSS.n4621 DVSS.n4610 1.5005
R12788 DVSS.n4730 DVSS.n4729 1.5005
R12789 DVSS.n2246 DVSS.n2230 1.5005
R12790 DVSS.n2245 DVSS.n2244 1.5005
R12791 DVSS.n2243 DVSS.n2242 1.5005
R12792 DVSS.n2241 DVSS.n2240 1.5005
R12793 DVSS.n2239 DVSS.n2238 1.5005
R12794 DVSS.n2237 DVSS.n2236 1.5005
R12795 DVSS.n2235 DVSS.n2234 1.5005
R12796 DVSS.n2233 DVSS.n2232 1.5005
R12797 DVSS.n2231 DVSS.n1958 1.5005
R12798 DVSS.n4158 DVSS.n4157 1.5005
R12799 DVSS.n1526 DVSS.n1525 1.5005
R12800 DVSS.n4143 DVSS.n4142 1.5005
R12801 DVSS.n4145 DVSS.n4144 1.5005
R12802 DVSS.n4147 DVSS.n4146 1.5005
R12803 DVSS.n4149 DVSS.n4148 1.5005
R12804 DVSS.n4151 DVSS.n4150 1.5005
R12805 DVSS.n4153 DVSS.n4152 1.5005
R12806 DVSS.n4141 DVSS.n1537 1.5005
R12807 DVSS.n3269 DVSS.n3268 1.5005
R12808 DVSS.n3267 DVSS.n1790 1.5005
R12809 DVSS.n3828 DVSS.n3827 1.5005
R12810 DVSS.n3271 DVSS.n3270 1.5005
R12811 DVSS.n3266 DVSS.n3000 1.5005
R12812 DVSS.n3265 DVSS.n2986 1.5005
R12813 DVSS.n3281 DVSS.n3280 1.5005
R12814 DVSS.n3283 DVSS.n3282 1.5005
R12815 DVSS.n2984 DVSS.n2980 1.5005
R12816 DVSS.n2983 DVSS.n2982 1.5005
R12817 DVSS.n2968 DVSS.n2967 1.5005
R12818 DVSS.n3293 DVSS.n3292 1.5005
R12819 DVSS.n3296 DVSS.n3295 1.5005
R12820 DVSS.n2966 DVSS.n2964 1.5005
R12821 DVSS.n2951 DVSS.n2949 1.5005
R12822 DVSS.n3306 DVSS.n3305 1.5005
R12823 DVSS.n3307 DVSS.n2946 1.5005
R12824 DVSS.n3309 DVSS.n3308 1.5005
R12825 DVSS.n2947 DVSS.n2945 1.5005
R12826 DVSS.n2932 DVSS.n2931 1.5005
R12827 DVSS.n3319 DVSS.n3318 1.5005
R12828 DVSS.n3321 DVSS.n3320 1.5005
R12829 DVSS.n2930 DVSS.n2928 1.5005
R12830 DVSS.n3007 DVSS.n2915 1.5005
R12831 DVSS.n3330 DVSS.n2914 1.5005
R12832 DVSS.n3332 DVSS.n3331 1.5005
R12833 DVSS.n3334 DVSS.n3333 1.5005
R12834 DVSS.n2913 DVSS.n2910 1.5005
R12835 DVSS.n2912 DVSS.n2897 1.5005
R12836 DVSS.n3344 DVSS.n3343 1.5005
R12837 DVSS.n3347 DVSS.n3346 1.5005
R12838 DVSS.n2896 DVSS.n2891 1.5005
R12839 DVSS.n2895 DVSS.n2894 1.5005
R12840 DVSS.n2879 DVSS.n2878 1.5005
R12841 DVSS.n3357 DVSS.n3356 1.5005
R12842 DVSS.n3359 DVSS.n3358 1.5005
R12843 DVSS.n2876 DVSS.n2874 1.5005
R12844 DVSS.n2861 DVSS.n2860 1.5005
R12845 DVSS.n3369 DVSS.n3368 1.5005
R12846 DVSS.n3371 DVSS.n3370 1.5005
R12847 DVSS.n2859 DVSS.n2853 1.5005
R12848 DVSS.n2858 DVSS.n2857 1.5005
R12849 DVSS.n2855 DVSS.n2841 1.5005
R12850 DVSS.n3381 DVSS.n3380 1.5005
R12851 DVSS.n3383 DVSS.n3382 1.5005
R12852 DVSS.n2839 DVSS.n2837 1.5005
R12853 DVSS.n2826 DVSS.n2825 1.5005
R12854 DVSS.n3393 DVSS.n3392 1.5005
R12855 DVSS.n3395 DVSS.n3394 1.5005
R12856 DVSS.n3397 DVSS.n3396 1.5005
R12857 DVSS.n3399 DVSS.n3398 1.5005
R12858 DVSS.n2821 DVSS.n2818 1.5005
R12859 DVSS.n2820 DVSS.n2805 1.5005
R12860 DVSS.n3409 DVSS.n3408 1.5005
R12861 DVSS.n3411 DVSS.n3410 1.5005
R12862 DVSS.n2803 DVSS.n2798 1.5005
R12863 DVSS.n2802 DVSS.n2801 1.5005
R12864 DVSS.n2786 DVSS.n2785 1.5005
R12865 DVSS.n3421 DVSS.n3420 1.5005
R12866 DVSS.n3423 DVSS.n3422 1.5005
R12867 DVSS.n2784 DVSS.n2782 1.5005
R12868 DVSS.n2769 DVSS.n2768 1.5005
R12869 DVSS.n3433 DVSS.n3432 1.5005
R12870 DVSS.n3435 DVSS.n3434 1.5005
R12871 DVSS.n2767 DVSS.n2761 1.5005
R12872 DVSS.n2766 DVSS.n2765 1.5005
R12873 DVSS.n2763 DVSS.n2749 1.5005
R12874 DVSS.n3445 DVSS.n3444 1.5005
R12875 DVSS.n3447 DVSS.n3446 1.5005
R12876 DVSS.n2747 DVSS.n2745 1.5005
R12877 DVSS.n2734 DVSS.n2733 1.5005
R12878 DVSS.n3457 DVSS.n3456 1.5005
R12879 DVSS.n3459 DVSS.n3458 1.5005
R12880 DVSS.n3461 DVSS.n3460 1.5005
R12881 DVSS.n3463 DVSS.n3462 1.5005
R12882 DVSS.n2730 DVSS.n2727 1.5005
R12883 DVSS.n2729 DVSS.n2714 1.5005
R12884 DVSS.n3473 DVSS.n3472 1.5005
R12885 DVSS.n3475 DVSS.n3474 1.5005
R12886 DVSS.n2712 DVSS.n2708 1.5005
R12887 DVSS.n2711 DVSS.n2710 1.5005
R12888 DVSS.n2696 DVSS.n2695 1.5005
R12889 DVSS.n3485 DVSS.n3484 1.5005
R12890 DVSS.n3487 DVSS.n3486 1.5005
R12891 DVSS.n2694 DVSS.n2692 1.5005
R12892 DVSS.n2676 DVSS.n2674 1.5005
R12893 DVSS.n3497 DVSS.n3496 1.5005
R12894 DVSS.n3498 DVSS.n2672 1.5005
R12895 DVSS.n3500 DVSS.n3499 1.5005
R12896 DVSS.n2673 DVSS.n2671 1.5005
R12897 DVSS.n3258 DVSS.n3003 1.5005
R12898 DVSS.n1791 DVSS.n1788 1.5005
R12899 DVSS.n3505 DVSS.n3504 1.5005
R12900 DVSS.n2668 DVSS.n2666 1.5005
R12901 DVSS.n3027 DVSS.n3026 1.5005
R12902 DVSS.n3031 DVSS.n3030 1.5005
R12903 DVSS.n3033 DVSS.n3032 1.5005
R12904 DVSS.n3036 DVSS.n3035 1.5005
R12905 DVSS.n3038 DVSS.n3037 1.5005
R12906 DVSS.n3042 DVSS.n3041 1.5005
R12907 DVSS.n3044 DVSS.n3043 1.5005
R12908 DVSS.n3045 DVSS.n3023 1.5005
R12909 DVSS.n3047 DVSS.n3046 1.5005
R12910 DVSS.n3050 DVSS.n3049 1.5005
R12911 DVSS.n3054 DVSS.n3053 1.5005
R12912 DVSS.n3056 DVSS.n3055 1.5005
R12913 DVSS.n3059 DVSS.n3058 1.5005
R12914 DVSS.n3060 DVSS.n3022 1.5005
R12915 DVSS.n3063 DVSS.n3062 1.5005
R12916 DVSS.n3021 DVSS.n3020 1.5005
R12917 DVSS.n3074 DVSS.n3073 1.5005
R12918 DVSS.n3076 DVSS.n3075 1.5005
R12919 DVSS.n3079 DVSS.n3078 1.5005
R12920 DVSS.n3081 DVSS.n3080 1.5005
R12921 DVSS.n3085 DVSS.n3084 1.5005
R12922 DVSS.n3088 DVSS.n3087 1.5005
R12923 DVSS.n3090 DVSS.n3089 1.5005
R12924 DVSS.n3092 DVSS.n3091 1.5005
R12925 DVSS.n3094 DVSS.n3093 1.5005
R12926 DVSS.n3098 DVSS.n3097 1.5005
R12927 DVSS.n3100 DVSS.n3099 1.5005
R12928 DVSS.n3103 DVSS.n3102 1.5005
R12929 DVSS.n3105 DVSS.n3104 1.5005
R12930 DVSS.n3109 DVSS.n3108 1.5005
R12931 DVSS.n3111 DVSS.n3110 1.5005
R12932 DVSS.n3112 DVSS.n3016 1.5005
R12933 DVSS.n3115 DVSS.n3114 1.5005
R12934 DVSS.n3118 DVSS.n3117 1.5005
R12935 DVSS.n3122 DVSS.n3121 1.5005
R12936 DVSS.n3124 DVSS.n3123 1.5005
R12937 DVSS.n3127 DVSS.n3126 1.5005
R12938 DVSS.n3128 DVSS.n3015 1.5005
R12939 DVSS.n3132 DVSS.n3131 1.5005
R12940 DVSS.n3014 DVSS.n3013 1.5005
R12941 DVSS.n3143 DVSS.n3142 1.5005
R12942 DVSS.n3145 DVSS.n3144 1.5005
R12943 DVSS.n3148 DVSS.n3147 1.5005
R12944 DVSS.n3150 DVSS.n3149 1.5005
R12945 DVSS.n3154 DVSS.n3153 1.5005
R12946 DVSS.n3157 DVSS.n3156 1.5005
R12947 DVSS.n3159 DVSS.n3158 1.5005
R12948 DVSS.n3161 DVSS.n3160 1.5005
R12949 DVSS.n3163 DVSS.n3162 1.5005
R12950 DVSS.n3167 DVSS.n3166 1.5005
R12951 DVSS.n3169 DVSS.n3168 1.5005
R12952 DVSS.n3172 DVSS.n3171 1.5005
R12953 DVSS.n3175 DVSS.n3174 1.5005
R12954 DVSS.n3179 DVSS.n3178 1.5005
R12955 DVSS.n3181 DVSS.n3180 1.5005
R12956 DVSS.n3182 DVSS.n3011 1.5005
R12957 DVSS.n3185 DVSS.n3184 1.5005
R12958 DVSS.n3187 DVSS.n3186 1.5005
R12959 DVSS.n3191 DVSS.n3190 1.5005
R12960 DVSS.n3193 DVSS.n3192 1.5005
R12961 DVSS.n3196 DVSS.n3195 1.5005
R12962 DVSS.n3198 DVSS.n3197 1.5005
R12963 DVSS.n3201 DVSS.n3009 1.5005
R12964 DVSS.n3203 DVSS.n3202 1.5005
R12965 DVSS.n3206 DVSS.n3205 1.5005
R12966 DVSS.n3209 DVSS.n3208 1.5005
R12967 DVSS.n3211 DVSS.n3210 1.5005
R12968 DVSS.n3215 DVSS.n3214 1.5005
R12969 DVSS.n3217 DVSS.n3216 1.5005
R12970 DVSS.n3220 DVSS.n3219 1.5005
R12971 DVSS.n3223 DVSS.n3222 1.5005
R12972 DVSS.n3224 DVSS.n3006 1.5005
R12973 DVSS.n3228 DVSS.n3227 1.5005
R12974 DVSS.n3230 DVSS.n3229 1.5005
R12975 DVSS.n3233 DVSS.n3232 1.5005
R12976 DVSS.n3235 DVSS.n3234 1.5005
R12977 DVSS.n3239 DVSS.n3238 1.5005
R12978 DVSS.n3241 DVSS.n3240 1.5005
R12979 DVSS.n3242 DVSS.n3004 1.5005
R12980 DVSS.n3244 DVSS.n3243 1.5005
R12981 DVSS.n3246 DVSS.n3245 1.5005
R12982 DVSS.n3250 DVSS.n3249 1.5005
R12983 DVSS.n3253 DVSS.n3252 1.5005
R12984 DVSS.n3256 DVSS.n3255 1.5005
R12985 DVSS.n3257 DVSS.n3001 1.5005
R12986 DVSS.n3260 DVSS.n3259 1.5005
R12987 DVSS.n3002 DVSS.n1787 1.5005
R12988 DVSS.n3263 DVSS.n3261 1.5005
R12989 DVSS.n3273 DVSS.n2997 1.5005
R12990 DVSS.n3254 DVSS.n2989 1.5005
R12991 DVSS.n3278 DVSS.n2988 1.5005
R12992 DVSS.n3248 DVSS.n3247 1.5005
R12993 DVSS.n3285 DVSS.n2978 1.5005
R12994 DVSS.n3242 DVSS.n2971 1.5005
R12995 DVSS.n3290 DVSS.n2970 1.5005
R12996 DVSS.n3237 DVSS.n3236 1.5005
R12997 DVSS.n3298 DVSS.n2961 1.5005
R12998 DVSS.n3231 DVSS.n2954 1.5005
R12999 DVSS.n3303 DVSS.n2953 1.5005
R13000 DVSS.n3226 DVSS.n3225 1.5005
R13001 DVSS.n3311 DVSS.n2942 1.5005
R13002 DVSS.n3218 DVSS.n2935 1.5005
R13003 DVSS.n3316 DVSS.n2934 1.5005
R13004 DVSS.n3213 DVSS.n3212 1.5005
R13005 DVSS.n3323 DVSS.n2925 1.5005
R13006 DVSS.n3207 DVSS.n2918 1.5005
R13007 DVSS.n3328 DVSS.n2917 1.5005
R13008 DVSS.n3200 DVSS.n3199 1.5005
R13009 DVSS.n3336 DVSS.n2907 1.5005
R13010 DVSS.n3194 DVSS.n2900 1.5005
R13011 DVSS.n3341 DVSS.n2899 1.5005
R13012 DVSS.n3189 DVSS.n3188 1.5005
R13013 DVSS.n3349 DVSS.n2889 1.5005
R13014 DVSS.n3183 DVSS.n2882 1.5005
R13015 DVSS.n3354 DVSS.n2881 1.5005
R13016 DVSS.n3177 DVSS.n3176 1.5005
R13017 DVSS.n3361 DVSS.n2871 1.5005
R13018 DVSS.n3170 DVSS.n2864 1.5005
R13019 DVSS.n3366 DVSS.n2863 1.5005
R13020 DVSS.n3165 DVSS.n3164 1.5005
R13021 DVSS.n3373 DVSS.n2851 1.5005
R13022 DVSS.n3012 DVSS.n2844 1.5005
R13023 DVSS.n3378 DVSS.n2843 1.5005
R13024 DVSS.n3152 DVSS.n3151 1.5005
R13025 DVSS.n3385 DVSS.n2834 1.5005
R13026 DVSS.n3146 DVSS.n2829 1.5005
R13027 DVSS.n3390 DVSS.n2828 1.5005
R13028 DVSS.n3141 DVSS.n3140 1.5005
R13029 DVSS.n3134 DVSS.n3133 1.5005
R13030 DVSS.n3401 DVSS.n2815 1.5005
R13031 DVSS.n3125 DVSS.n2808 1.5005
R13032 DVSS.n3406 DVSS.n2807 1.5005
R13033 DVSS.n3120 DVSS.n3119 1.5005
R13034 DVSS.n3413 DVSS.n2796 1.5005
R13035 DVSS.n3113 DVSS.n2789 1.5005
R13036 DVSS.n3418 DVSS.n2788 1.5005
R13037 DVSS.n3107 DVSS.n3106 1.5005
R13038 DVSS.n3425 DVSS.n2779 1.5005
R13039 DVSS.n3101 DVSS.n2772 1.5005
R13040 DVSS.n3430 DVSS.n2771 1.5005
R13041 DVSS.n3096 DVSS.n3095 1.5005
R13042 DVSS.n3437 DVSS.n2759 1.5005
R13043 DVSS.n3019 DVSS.n2752 1.5005
R13044 DVSS.n3442 DVSS.n2751 1.5005
R13045 DVSS.n3083 DVSS.n3082 1.5005
R13046 DVSS.n3449 DVSS.n2742 1.5005
R13047 DVSS.n3077 DVSS.n2737 1.5005
R13048 DVSS.n3454 DVSS.n2736 1.5005
R13049 DVSS.n3072 DVSS.n3071 1.5005
R13050 DVSS.n3065 DVSS.n3064 1.5005
R13051 DVSS.n3465 DVSS.n2724 1.5005
R13052 DVSS.n3057 DVSS.n2717 1.5005
R13053 DVSS.n3470 DVSS.n2716 1.5005
R13054 DVSS.n3052 DVSS.n3051 1.5005
R13055 DVSS.n3477 DVSS.n2706 1.5005
R13056 DVSS.n3045 DVSS.n2699 1.5005
R13057 DVSS.n3482 DVSS.n2698 1.5005
R13058 DVSS.n3040 DVSS.n3039 1.5005
R13059 DVSS.n3489 DVSS.n2689 1.5005
R13060 DVSS.n3034 DVSS.n2679 1.5005
R13061 DVSS.n3494 DVSS.n2678 1.5005
R13062 DVSS.n3029 DVSS.n3028 1.5005
R13063 DVSS.n3503 DVSS.n3502 1.5005
R13064 DVSS.n1789 DVSS.n1787 1.5005
R13065 DVSS.n3264 DVSS.n3263 1.5005
R13066 DVSS.n3273 DVSS.n3272 1.5005
R13067 DVSS.n2999 DVSS.n2989 1.5005
R13068 DVSS.n3279 DVSS.n3278 1.5005
R13069 DVSS.n3247 DVSS.n2981 1.5005
R13070 DVSS.n3285 DVSS.n3284 1.5005
R13071 DVSS.n2982 DVSS.n2971 1.5005
R13072 DVSS.n3291 DVSS.n3290 1.5005
R13073 DVSS.n3236 DVSS.n2965 1.5005
R13074 DVSS.n3298 DVSS.n3297 1.5005
R13075 DVSS.n2963 DVSS.n2954 1.5005
R13076 DVSS.n3304 DVSS.n3303 1.5005
R13077 DVSS.n3225 DVSS.n2950 1.5005
R13078 DVSS.n3311 DVSS.n3310 1.5005
R13079 DVSS.n2944 DVSS.n2935 1.5005
R13080 DVSS.n3317 DVSS.n3316 1.5005
R13081 DVSS.n3212 DVSS.n2929 1.5005
R13082 DVSS.n3323 DVSS.n3322 1.5005
R13083 DVSS.n2927 DVSS.n2918 1.5005
R13084 DVSS.n3329 DVSS.n3328 1.5005
R13085 DVSS.n3199 DVSS.n2911 1.5005
R13086 DVSS.n3336 DVSS.n3335 1.5005
R13087 DVSS.n2909 DVSS.n2900 1.5005
R13088 DVSS.n3342 DVSS.n3341 1.5005
R13089 DVSS.n3188 DVSS.n2892 1.5005
R13090 DVSS.n3349 DVSS.n3348 1.5005
R13091 DVSS.n2893 DVSS.n2882 1.5005
R13092 DVSS.n3355 DVSS.n3354 1.5005
R13093 DVSS.n3176 DVSS.n2875 1.5005
R13094 DVSS.n3361 DVSS.n3360 1.5005
R13095 DVSS.n2873 DVSS.n2864 1.5005
R13096 DVSS.n3367 DVSS.n3366 1.5005
R13097 DVSS.n3164 DVSS.n2854 1.5005
R13098 DVSS.n3373 DVSS.n3372 1.5005
R13099 DVSS.n2856 DVSS.n2844 1.5005
R13100 DVSS.n3379 DVSS.n3378 1.5005
R13101 DVSS.n3151 DVSS.n2838 1.5005
R13102 DVSS.n3385 DVSS.n3384 1.5005
R13103 DVSS.n2836 DVSS.n2829 1.5005
R13104 DVSS.n3391 DVSS.n3390 1.5005
R13105 DVSS.n3140 DVSS.n2823 1.5005
R13106 DVSS.n3134 DVSS.n2819 1.5005
R13107 DVSS.n3401 DVSS.n3400 1.5005
R13108 DVSS.n2817 DVSS.n2808 1.5005
R13109 DVSS.n3407 DVSS.n3406 1.5005
R13110 DVSS.n3119 DVSS.n2799 1.5005
R13111 DVSS.n3413 DVSS.n3412 1.5005
R13112 DVSS.n2800 DVSS.n2789 1.5005
R13113 DVSS.n3419 DVSS.n3418 1.5005
R13114 DVSS.n3106 DVSS.n2783 1.5005
R13115 DVSS.n3425 DVSS.n3424 1.5005
R13116 DVSS.n2781 DVSS.n2772 1.5005
R13117 DVSS.n3431 DVSS.n3430 1.5005
R13118 DVSS.n3095 DVSS.n2762 1.5005
R13119 DVSS.n3437 DVSS.n3436 1.5005
R13120 DVSS.n2764 DVSS.n2752 1.5005
R13121 DVSS.n3443 DVSS.n3442 1.5005
R13122 DVSS.n3082 DVSS.n2746 1.5005
R13123 DVSS.n3449 DVSS.n3448 1.5005
R13124 DVSS.n2744 DVSS.n2737 1.5005
R13125 DVSS.n3455 DVSS.n3454 1.5005
R13126 DVSS.n3071 DVSS.n2732 1.5005
R13127 DVSS.n3065 DVSS.n2728 1.5005
R13128 DVSS.n3465 DVSS.n3464 1.5005
R13129 DVSS.n2726 DVSS.n2717 1.5005
R13130 DVSS.n3471 DVSS.n3470 1.5005
R13131 DVSS.n3051 DVSS.n2709 1.5005
R13132 DVSS.n3477 DVSS.n3476 1.5005
R13133 DVSS.n2710 DVSS.n2699 1.5005
R13134 DVSS.n3483 DVSS.n3482 1.5005
R13135 DVSS.n3039 DVSS.n2693 1.5005
R13136 DVSS.n3489 DVSS.n3488 1.5005
R13137 DVSS.n2691 DVSS.n2679 1.5005
R13138 DVSS.n3495 DVSS.n3494 1.5005
R13139 DVSS.n3028 DVSS.n2675 1.5005
R13140 DVSS.n3502 DVSS.n3501 1.5005
R13141 DVSS.n1391 DVSS.n1356 1.5005
R13142 DVSS.n1390 DVSS.n1389 1.5005
R13143 DVSS.n1388 DVSS.n1387 1.5005
R13144 DVSS.n1386 DVSS.n1385 1.5005
R13145 DVSS.n1384 DVSS.n1383 1.5005
R13146 DVSS.n1382 DVSS.n1381 1.5005
R13147 DVSS.n1380 DVSS.n1379 1.5005
R13148 DVSS.n1378 DVSS.n1377 1.5005
R13149 DVSS.n1376 DVSS.n1375 1.5005
R13150 DVSS.n1374 DVSS.n1373 1.5005
R13151 DVSS.n1372 DVSS.n1367 1.5005
R13152 DVSS.n4767 DVSS.n4766 1.5005
R13153 DVSS.n4140 DVSS.n1538 1.49818
R13154 DVSS.n3796 DVSS.n2630 1.49138
R13155 DVSS.n2539 DVSS.n2538 1.44688
R13156 DVSS.n2266 DVSS.n1928 1.44688
R13157 DVSS DVSS.n1453 1.41642
R13158 DVSS.n1460 DVSS 1.41642
R13159 DVSS.n4805 DVSS 1.41642
R13160 DVSS.n1227 DVSS 1.41642
R13161 DVSS DVSS.n4819 1.41642
R13162 DVSS DVSS.n1224 1.41642
R13163 DVSS.n1498 DVSS 1.41642
R13164 DVSS.n4183 DVSS 1.41642
R13165 DVSS.n1974 DVSS 1.41642
R13166 DVSS.n1266 DVSS 1.41642
R13167 DVSS.n1269 DVSS 1.41642
R13168 DVSS.n1345 DVSS 1.41642
R13169 DVSS.n4823 DVSS.n4822 1.39741
R13170 DVSS.n5099 DVSS.n5095 1.38866
R13171 DVSS.n2308 DVSS.n1929 1.35477
R13172 DVSS.n2547 DVSS.n1919 1.35477
R13173 DVSS.n3787 DVSS.n3785 1.328
R13174 DVSS.n1631 DVSS.n1625 1.31286
R13175 DVSS.n2623 DVSS.n1652 1.31286
R13176 DVSS.n3958 DVSS.n3957 1.31286
R13177 DVSS.n3773 DVSS.n1735 1.31286
R13178 DVSS.n4864 DVSS.n1203 1.3005
R13179 DVSS.n4113 DVSS.n4112 1.3005
R13180 DVSS.n4118 DVSS.n4117 1.3005
R13181 DVSS.n4838 DVSS.n4837 1.3005
R13182 DVSS.n4843 DVSS.n1215 1.3005
R13183 DVSS.n1261 DVSS.n1260 1.3005
R13184 DVSS.n1258 DVSS.n1257 1.3005
R13185 DVSS.n1505 DVSS.n1504 1.3005
R13186 DVSS.n1509 DVSS.n1508 1.3005
R13187 DVSS.n4296 DVSS.n1466 1.29067
R13188 DVSS.n4292 DVSS.n1471 1.29067
R13189 DVSS.n4786 DVSS.n1253 1.29067
R13190 DVSS.n1233 DVSS.n1232 1.29067
R13191 DVSS.n2659 VSS 1.28985
R13192 DVSS.n4779 DVSS.n4778 1.26649
R13193 DVSS.n4029 DVSS.n1617 1.25594
R13194 DVSS.n1708 DVSS.n1705 1.25594
R13195 DVSS.n4100 DVSS.n4099 1.20054
R13196 DVSS.n4099 DVSS.n1552 1.19935
R13197 DVSS.n4840 DVSS.n1156 1.19925
R13198 DVSS.n4806 DVSS.n4805 1.16866
R13199 DVSS.n4183 DVSS.n4182 1.16866
R13200 DVSS.n1974 DVSS.n1973 1.16866
R13201 DVSS.n1267 DVSS.n1266 1.16866
R13202 DVSS.n1345 DVSS.n1344 1.16866
R13203 DVSS.n1838 DVSS.n1695 1.16402
R13204 DVSS.n4303 DVSS.n1455 1.15745
R13205 DVSS.n3798 DVSS.n3797 1.15606
R13206 DVSS.n4288 DVSS.n4287 1.15606
R13207 DVSS.n4827 DVSS.n4826 1.15606
R13208 DVSS.n4853 DVSS.n4852 1.15606
R13209 DVSS.n4859 DVSS.n4858 1.15606
R13210 DVSS.n2618 DVSS.n2615 1.13009
R13211 DVSS.n1839 DVSS.n1830 1.12941
R13212 DVSS.n3940 DVSS.n3939 1.10843
R13213 DVSS.n3957 DVSS.n1683 1.10563
R13214 DVSS.n3774 DVSS.n3773 1.10563
R13215 DVSS.n2652 DVSS.n1625 1.10563
R13216 DVSS.n2624 DVSS.n2623 1.10563
R13217 DVSS.n1847 DVSS.t138 1.0925
R13218 DVSS.n4301 DVSS.t175 1.0925
R13219 DVSS.n4301 DVSS.t159 1.0925
R13220 DVSS.n1698 DVSS.t94 1.0925
R13221 DVSS.n1698 DVSS.t192 1.0925
R13222 DVSS.n3941 DVSS.t100 1.0925
R13223 DVSS.n3941 DVSS.t141 1.0925
R13224 DVSS.n1612 DVSS.t136 1.0925
R13225 DVSS.n1612 DVSS.t177 1.0925
R13226 DVSS.n1620 DVSS.t145 1.0925
R13227 DVSS.n1620 DVSS.t109 1.0925
R13228 DVSS.n1829 DVSS.t77 1.0925
R13229 DVSS.n1268 DVSS.n1234 1.08844
R13230 DVSS.n4807 DVSS.n1234 1.08844
R13231 DVSS.n4181 DVSS.n4180 1.08844
R13232 DVSS.n4180 DVSS.n1462 1.08844
R13233 DVSS.n4808 DVSS.n4807 1.0805
R13234 DVSS.n4181 DVSS.n1501 1.0805
R13235 DVSS.n4312 DVSS.n1462 1.0805
R13236 DVSS.n4782 DVSS.n1268 1.0805
R13237 DVSS.n3939 DVSS.n1695 1.07932
R13238 DVSS.n4360 DVSS.n956 1.07349
R13239 DVSS.n2287 DVSS.n2277 1.05604
R13240 DVSS.n1458 DVSS.n1457 1.0505
R13241 DVSS.n4816 DVSS.n4815 1.0505
R13242 DVSS.n1480 DVSS.n1479 1.0505
R13243 DVSS.n1273 DVSS.n1272 1.0505
R13244 DVSS.n1514 DVSS.n1506 1.05029
R13245 DVSS.n2658 DVSS.n2657 1.0405
R13246 DVSS.n2657 DVSS.n2654 1.0405
R13247 DVSS.n3791 DVSS.n3790 1.0405
R13248 DVSS.n2642 DVSS.n2640 1.0405
R13249 DVSS.n2642 DVSS.n2641 1.0405
R13250 DVSS.n3780 DVSS.n3779 1.0405
R13251 DVSS.n3779 DVSS.n3778 1.0405
R13252 DVSS.n2616 DVSS.n1846 1.0405
R13253 DVSS.n1511 DVSS.n1510 1.0405
R13254 DVSS.n4786 DVSS.n4785 1.0405
R13255 DVSS.n4785 DVSS.n4784 1.0405
R13256 DVSS.n4292 DVSS.n4291 1.0405
R13257 DVSS.n4291 DVSS.n4290 1.0405
R13258 DVSS.n4811 DVSS.n1233 1.0405
R13259 DVSS.n4811 DVSS.n4810 1.0405
R13260 DVSS.n4297 DVSS.n4296 1.0405
R13261 DVSS.n4298 DVSS.n4297 1.0405
R13262 DVSS.n1212 DVSS.n1211 1.02439
R13263 DVSS.n1475 DVSS.n1474 1.02439
R13264 DVSS.n1220 DVSS.n1219 1.02439
R13265 DVSS.n1207 DVSS.n1206 1.02439
R13266 DVSS.n3776 DVSS.t85 1.00732
R13267 DVSS.n1705 DVSS.n1704 1.00517
R13268 DVSS.n1623 DVSS.n1617 1.00517
R13269 DVSS.n4058 VSS 1.00241
R13270 DVSS.n3783 DVSS.n3782 0.998789
R13271 DVSS.n2619 DVSS.n1846 0.998488
R13272 DVSS.n3790 DVSS.n3789 0.996088
R13273 DVSS.n1512 DVSS.n1511 0.996088
R13274 DVSS.n1571 DVSS.n1081 0.988551
R13275 DVSS.n3793 DVSS.t173 0.958395
R13276 DVSS.n3793 DVSS.t178 0.958395
R13277 DVSS.n3251 DVSS.t48 0.9581
R13278 DVSS.n3221 DVSS.t56 0.9581
R13279 DVSS.n3010 DVSS.t50 0.9581
R13280 DVSS.n3155 DVSS.t59 0.9581
R13281 DVSS.n3116 DVSS.t51 0.9581
R13282 DVSS.n3086 DVSS.t55 0.9581
R13283 DVSS.n3048 DVSS.t49 0.9581
R13284 DVSS.n3506 DVSS.t58 0.9581
R13285 DVSS.n2985 DVSS.t48 0.9581
R13286 DVSS.n2948 DVSS.t56 0.9581
R13287 DVSS.n3345 DVSS.t50 0.9581
R13288 DVSS.n2840 DVSS.t59 0.9581
R13289 DVSS.n2804 DVSS.t51 0.9581
R13290 DVSS.n2748 DVSS.t55 0.9581
R13291 DVSS.n2713 DVSS.t49 0.9581
R13292 DVSS.n2665 DVSS.t58 0.9581
R13293 DVSS.n4871 DVSS.n4870 0.945955
R13294 DVSS.n4058 DVSS.n4057 0.945955
R13295 DVSS.n4286 DVSS.n4285 0.945955
R13296 DVSS.n4840 DVSS.n4839 0.945955
R13297 DVSS.n4857 DVSS.n4856 0.945955
R13298 DVSS.n1454 DVSS.n1453 0.941532
R13299 DVSS.n4820 DVSS.n4819 0.941532
R13300 DVSS.n1225 DVSS.n1224 0.941532
R13301 DVSS.n1459 DVSS.n1458 0.941367
R13302 DVSS.n1461 DVSS.n1460 0.941367
R13303 DVSS.n1228 DVSS.n1227 0.941367
R13304 DVSS.n4817 DVSS.n4816 0.941367
R13305 DVSS.n1481 DVSS.n1480 0.941367
R13306 DVSS.n1499 DVSS.n1498 0.941367
R13307 DVSS.n1270 DVSS.n1269 0.941367
R13308 DVSS.n1274 DVSS.n1273 0.941367
R13309 DVSS.n3768 DVSS.n3767 0.922787
R13310 DVSS.n3522 DVSS.n3521 0.922694
R13311 DVSS.n5093 DVSS.n5092 0.922457
R13312 DVSS.n4095 DVSS.n4094 0.910322
R13313 DVSS.n955 DVSS.n952 0.902366
R13314 DVSS.n5345 DVSS.n952 0.902313
R13315 DVSS.n5345 DVSS.n5344 0.902282
R13316 DVSS.n5344 DVSS.n955 0.901878
R13317 DVSS.n5342 DVSS.n956 0.879171
R13318 DVSS.n4765 DVSS.n1370 0.879171
R13319 DVSS.n3944 DVSS.n3943 0.875366
R13320 DVSS.n1729 DVSS.n1728 0.875366
R13321 DVSS.n3955 DVSS.n3954 0.87493
R13322 DVSS.n4803 DVSS.n4802 0.8749
R13323 DVSS.n4186 DVSS.n4185 0.8749
R13324 DVSS.n1348 DVSS.n1347 0.8749
R13325 DVSS.n4093 DVSS.n1555 0.873402
R13326 DVSS.n1457 DVSS.n1456 0.872079
R13327 DVSS.n4815 DVSS.n4814 0.872079
R13328 DVSS.n1479 DVSS.n1478 0.872079
R13329 DVSS.n1272 DVSS.n1271 0.872079
R13330 DVSS.n4766 DVSS.n4765 0.870066
R13331 DVSS.n4051 DVSS.n1624 0.867167
R13332 DVSS.n4056 DVSS.n4055 0.867167
R13333 DVSS.n1703 DVSS.n1684 0.867167
R13334 DVSS.n3936 DVSS.n3935 0.867167
R13335 DVSS.n2640 DVSS.n2635 0.843937
R13336 DVSS.n2658 DVSS.n2634 0.843937
R13337 DVSS.n3781 DVSS.n3780 0.843937
R13338 DVSS.n3940 DVSS.n1686 0.827218
R13339 DVSS.n5539 DVSS.n5538 0.820816
R13340 DVSS.n3785 DVSS.n3784 0.815237
R13341 DVSS.n1838 DVSS.n1837 0.80914
R13342 DVSS.n4308 DVSS.n4305 0.8005
R13343 DVSS.n4121 DVSS.n1546 0.796907
R13344 DVSS.n4125 DVSS.n1546 0.796907
R13345 DVSS.n4125 DVSS.n1544 0.796907
R13346 DVSS.n4129 DVSS.n1544 0.796907
R13347 DVSS.n4129 DVSS.n1542 0.796907
R13348 DVSS.n4133 DVSS.n1542 0.796907
R13349 DVSS.n4133 DVSS.n1519 0.796907
R13350 DVSS.n4168 DVSS.n1519 0.796907
R13351 DVSS.n4168 DVSS.n1520 0.796907
R13352 DVSS.n4871 VSS 0.78605
R13353 DVSS.n2306 DVSS.n2253 0.778288
R13354 DVSS.n4283 DVSS.n4282 0.774059
R13355 DVSS.n4778 DVSS.n4777 0.752663
R13356 DVSS.n2627 DVSS.n2626 0.751952
R13357 DVSS.n2638 VSS 0.751638
R13358 DVSS.n2267 DVSS.n2266 0.7505
R13359 DVSS.n2538 DVSS.n1926 0.7505
R13360 DVSS DVSS.n2618 0.746344
R13361 DVSS.n5600 DVSS.n5599 0.745113
R13362 DVSS.n688 DVSS.n169 0.745113
R13363 DVSS.n620 DVSS.n194 0.745113
R13364 DVSS.n2310 DVSS.n1930 0.743357
R13365 DVSS.n2310 DVSS.n2309 0.743357
R13366 DVSS.n2549 DVSS.n1920 0.743357
R13367 DVSS.n2549 DVSS.n2548 0.743357
R13368 DVSS.n2540 DVSS.n1921 0.743357
R13369 DVSS.n2548 DVSS.n1921 0.743357
R13370 DVSS.n1933 DVSS.n1918 0.743357
R13371 DVSS.n2309 DVSS.n1918 0.743357
R13372 DVSS.n5600 DVSS.n123 0.736857
R13373 DVSS.n688 DVSS.n687 0.736857
R13374 DVSS.n621 DVSS.n620 0.736857
R13375 DVSS.n2542 DVSS.n2541 0.735937
R13376 DVSS.n2303 DVSS.n2302 0.735937
R13377 DVSS.n4315 DVSS.n1455 0.7304
R13378 DVSS.n3945 DVSS.n3944 0.71546
R13379 DVSS.n1730 DVSS.n1729 0.71546
R13380 DVSS.n3954 DVSS.n3953 0.71533
R13381 DVSS.n1501 DVSS.n1500 0.707265
R13382 DVSS.n1841 DVSS.n1827 0.696386
R13383 DVSS.n1840 DVSS.n1828 0.696386
R13384 DVSS.n1255 DVSS.n1230 0.693432
R13385 DVSS.n1262 DVSS.n1251 0.693432
R13386 DVSS.n1472 DVSS.n1469 0.693432
R13387 DVSS.n1467 DVSS.n1464 0.693432
R13388 DVSS.n4293 DVSS.n1469 0.682241
R13389 DVSS.n4787 DVSS.n1251 0.682241
R13390 DVSS.n1255 DVSS.n1250 0.682241
R13391 DVSS.n4295 DVSS.n1467 0.682241
R13392 DVSS.n4140 DVSS.n4139 0.666308
R13393 DVSS.n4165 DVSS.n4164 0.66242
R13394 DVSS.n4808 DVSS.n1229 0.662265
R13395 DVSS.n4313 DVSS.n4312 0.662265
R13396 DVSS.n4782 DVSS.n4781 0.662265
R13397 DVSS.n4139 DVSS.n1539 0.64762
R13398 DVSS.n1841 DVSS.n1840 0.646382
R13399 DVSS.n4609 DVSS.n4608 0.643357
R13400 DVSS.n4624 DVSS.n4623 0.643357
R13401 DVSS.n4626 DVSS.n4619 0.643357
R13402 DVSS.n4719 DVSS.n4718 0.643357
R13403 DVSS.n4588 DVSS.n4587 0.643357
R13404 DVSS.n4589 DVSS.n1395 0.643357
R13405 DVSS.n4752 DVSS.n4751 0.643357
R13406 DVSS.n1398 DVSS.n1396 0.643357
R13407 DVSS.n4549 DVSS.n4548 0.643357
R13408 DVSS.n4552 DVSS.n4551 0.643357
R13409 DVSS.n1419 DVSS.n1418 0.643357
R13410 DVSS.n4566 DVSS.n4565 0.643357
R13411 DVSS.n4447 DVSS.n1448 0.643357
R13412 DVSS.n4513 DVSS.n4512 0.643357
R13413 DVSS.n1440 DVSS.n1439 0.643357
R13414 DVSS.n4526 DVSS.n4525 0.643357
R13415 DVSS.n4416 DVSS.n4415 0.643357
R13416 DVSS.n4431 DVSS.n4430 0.643357
R13417 DVSS.n4433 DVSS.n4426 0.643357
R13418 DVSS.n4471 DVSS.n4470 0.643357
R13419 DVSS.n4395 DVSS.n4394 0.643357
R13420 DVSS.n4396 DVSS.n4324 0.643357
R13421 DVSS.n4504 DVSS.n4503 0.643357
R13422 DVSS.n4327 DVSS.n4325 0.643357
R13423 DVSS.n4114 DVSS.n4113 0.634889
R13424 DVSS.n4116 VSS 0.622069
R13425 DVSS.n1550 VSS 0.622069
R13426 DVSS.n4836 VSS 0.622069
R13427 DVSS.n4842 VSS 0.622069
R13428 DVSS.n4863 VSS 0.622069
R13429 DVSS.n1840 DVSS.n1839 0.618588
R13430 DVSS.n4164 DVSS 0.600908
R13431 DVSS.n4314 DVSS.n1459 0.597759
R13432 DVSS.n4313 DVSS.n1461 0.597759
R13433 DVSS.n1229 DVSS.n1228 0.597759
R13434 DVSS.n4818 DVSS.n4817 0.597759
R13435 DVSS.n1482 DVSS.n1481 0.597759
R13436 DVSS.n4781 DVSS.n1270 0.597759
R13437 DVSS.n4780 DVSS.n1274 0.597759
R13438 DVSS DVSS.n1454 0.595564
R13439 DVSS DVSS.n4820 0.595564
R13440 DVSS DVSS.n1225 0.595564
R13441 DVSS.n3817 DVSS.n3816 0.588678
R13442 DVSS.n2643 DVSS.n2635 0.585632
R13443 DVSS.n2656 DVSS.n2634 0.585632
R13444 DVSS.n3781 DVSS.n2637 0.585632
R13445 DVSS.n3957 DVSS.n3956 0.584525
R13446 DVSS.n3773 DVSS.n1697 0.584525
R13447 DVSS.n4050 DVSS.n1625 0.584525
R13448 DVSS.n2623 DVSS.n1611 0.584525
R13449 DVSS.n1515 VSS 0.581806
R13450 DVSS.n3816 DVSS.n1801 0.578278
R13451 DVSS.n3815 DVSS.n1804 0.578278
R13452 DVSS.n3814 DVSS.n1800 0.578278
R13453 DVSS.n3813 DVSS.n1806 0.578278
R13454 DVSS.n3812 DVSS.n1799 0.578278
R13455 DVSS.n3811 DVSS.n1808 0.578278
R13456 DVSS.n3810 DVSS.n1798 0.578278
R13457 DVSS.n3809 DVSS.n1810 0.578278
R13458 DVSS.n3808 DVSS.n1797 0.578278
R13459 DVSS.n3807 DVSS.n1812 0.578278
R13460 DVSS.n3806 DVSS.n1796 0.578278
R13461 DVSS.n3820 DVSS.n1843 0.578278
R13462 DVSS DVSS.n3826 0.578278
R13463 DVSS.n3826 DVSS.n3825 0.578278
R13464 DVSS.n3508 DVSS.n3507 0.578278
R13465 DVSS.n4166 DVSS.n1520 0.578278
R13466 DVSS.n1520 DVSS.n1518 0.578278
R13467 DVSS.n4168 DVSS.n4167 0.578278
R13468 DVSS.n4169 DVSS.n4168 0.578278
R13469 DVSS.n1521 DVSS.n1519 0.578278
R13470 DVSS.n1519 DVSS.n1517 0.578278
R13471 DVSS.n4133 DVSS.n4132 0.578278
R13472 DVSS.n4134 DVSS.n4133 0.578278
R13473 DVSS.n4131 DVSS.n1542 0.578278
R13474 DVSS.n1542 DVSS.n1541 0.578278
R13475 DVSS.n4130 DVSS.n4129 0.578278
R13476 DVSS.n4129 DVSS.n4128 0.578278
R13477 DVSS.n1544 DVSS.n1543 0.578278
R13478 DVSS.n4127 DVSS.n1544 0.578278
R13479 DVSS.n4125 DVSS.n4124 0.578278
R13480 DVSS.n4126 DVSS.n4125 0.578278
R13481 DVSS.n4123 DVSS.n1546 0.578278
R13482 DVSS.n4119 DVSS.n1546 0.578278
R13483 DVSS.n4122 DVSS.n4121 0.578278
R13484 DVSS.n4121 DVSS.n4120 0.578278
R13485 DVSS.n3782 DVSS.n3781 0.563
R13486 DVSS.n4285 DVSS.n4284 0.557079
R13487 DVSS.n3797 DVSS.n3796 0.557079
R13488 DVSS.n3788 DVSS.n3787 0.557079
R13489 DVSS.n4841 DVSS.n4840 0.557079
R13490 DVSS.n4856 DVSS.n4855 0.557079
R13491 DVSS.n4837 DVSS.n4835 0.553108
R13492 DVSS.n4847 DVSS.n4843 0.553108
R13493 DVSS.n4868 DVSS.n4864 0.553108
R13494 DVSS.n1500 DVSS.n1499 0.548022
R13495 DVSS.n1211 DVSS.t84 0.5465
R13496 DVSS.n1211 DVSS.t73 0.5465
R13497 DVSS.n1474 DVSS.t43 0.5465
R13498 DVSS.n1474 DVSS.t172 0.5465
R13499 DVSS.n1219 DVSS.t189 0.5465
R13500 DVSS.n1219 DVSS.t147 0.5465
R13501 DVSS.n1206 DVSS.t166 0.5465
R13502 DVSS.n1206 DVSS.t199 0.5465
R13503 DVSS.n2648 DVSS.n2647 0.545794
R13504 DVSS.n4309 DVSS.n4308 0.545794
R13505 DVSS.n4314 DVSS.n4313 0.545794
R13506 DVSS.n4818 DVSS.n1229 0.545794
R13507 DVSS.n4821 DVSS.n4818 0.545794
R13508 DVSS.n1482 DVSS.n1226 0.545794
R13509 DVSS.n3956 DVSS.n1684 0.545794
R13510 DVSS.n3935 DVSS.n1697 0.545794
R13511 DVSS.n4055 DVSS.n1611 0.545794
R13512 DVSS.n4051 DVSS.n4050 0.545794
R13513 DVSS.n4781 DVSS.n4780 0.545794
R13514 DVSS.n4780 DVSS.n4779 0.545794
R13515 DVSS.n4807 DVSS.n4806 0.5442
R13516 DVSS.n4182 DVSS.n4181 0.5442
R13517 DVSS.n1973 DVSS.n1462 0.5442
R13518 DVSS.n1268 DVSS.n1267 0.5442
R13519 DVSS.n1555 VSS 0.544091
R13520 DVSS.n4095 VSS 0.544091
R13521 DVSS.n2662 DVSS.n2661 0.543147
R13522 DVSS.n1344 DVSS 0.541831
R13523 DVSS.n2629 DVSS.n2627 0.536572
R13524 DVSS.n1264 DVSS.n1210 0.532494
R13525 DVSS.n2302 DVSS.n1930 0.5255
R13526 DVSS.n2541 DVSS.n2540 0.5255
R13527 DVSS.n2656 DVSS.n2655 0.5205
R13528 DVSS.n2644 DVSS.n2643 0.5205
R13529 DVSS.n3776 DVSS.n2637 0.5205
R13530 DVSS.n4854 DVSS.n1212 0.518873
R13531 DVSS.n1476 DVSS.n1475 0.518873
R13532 DVSS.n1221 DVSS.n1220 0.518873
R13533 DVSS.n1208 DVSS.n1207 0.518873
R13534 DVSS.n1833 DVSS.t184 0.512375
R13535 DVSS.n1833 DVSS.t96 0.512375
R13536 DVSS.n1831 DVSS.t90 0.512375
R13537 DVSS.n1831 DVSS.t182 0.512375
R13538 DVSS.n1513 VSS 0.50383
R13539 DVSS.n1466 DVSS.n1465 0.500875
R13540 DVSS.n1471 DVSS.n1470 0.500875
R13541 DVSS.n1253 DVSS.n1252 0.500875
R13542 DVSS.n1232 DVSS.n1231 0.500875
R13543 DVSS.n2685 DVSS.n2680 0.5005
R13544 DVSS.n3492 DVSS.n2686 0.5005
R13545 DVSS.n3491 DVSS.n2687 0.5005
R13546 DVSS.n2701 DVSS.n2688 0.5005
R13547 DVSS.n2702 DVSS.n2700 0.5005
R13548 DVSS.n3480 DVSS.n2703 0.5005
R13549 DVSS.n3479 DVSS.n2704 0.5005
R13550 DVSS.n2719 DVSS.n2705 0.5005
R13551 DVSS.n2720 DVSS.n2718 0.5005
R13552 DVSS.n3468 DVSS.n2721 0.5005
R13553 DVSS.n3467 DVSS.n2722 0.5005
R13554 DVSS.n3066 DVSS.n2723 0.5005
R13555 DVSS.n3069 DVSS.n3068 0.5005
R13556 DVSS.n3067 DVSS.n2738 0.5005
R13557 DVSS.n3452 DVSS.n2739 0.5005
R13558 DVSS.n3451 DVSS.n2740 0.5005
R13559 DVSS.n2754 DVSS.n2741 0.5005
R13560 DVSS.n2755 DVSS.n2753 0.5005
R13561 DVSS.n3440 DVSS.n2756 0.5005
R13562 DVSS.n3439 DVSS.n2757 0.5005
R13563 DVSS.n2774 DVSS.n2758 0.5005
R13564 DVSS.n2775 DVSS.n2773 0.5005
R13565 DVSS.n3428 DVSS.n2776 0.5005
R13566 DVSS.n3427 DVSS.n2777 0.5005
R13567 DVSS.n2791 DVSS.n2778 0.5005
R13568 DVSS.n2792 DVSS.n2790 0.5005
R13569 DVSS.n3416 DVSS.n2793 0.5005
R13570 DVSS.n3415 DVSS.n2794 0.5005
R13571 DVSS.n2810 DVSS.n2795 0.5005
R13572 DVSS.n2811 DVSS.n2809 0.5005
R13573 DVSS.n3404 DVSS.n2812 0.5005
R13574 DVSS.n3403 DVSS.n2813 0.5005
R13575 DVSS.n3135 DVSS.n2814 0.5005
R13576 DVSS.n3138 DVSS.n3137 0.5005
R13577 DVSS.n3136 DVSS.n2830 0.5005
R13578 DVSS.n3388 DVSS.n2831 0.5005
R13579 DVSS.n3387 DVSS.n2832 0.5005
R13580 DVSS.n2846 DVSS.n2833 0.5005
R13581 DVSS.n2847 DVSS.n2845 0.5005
R13582 DVSS.n3376 DVSS.n2848 0.5005
R13583 DVSS.n3375 DVSS.n2849 0.5005
R13584 DVSS.n2866 DVSS.n2850 0.5005
R13585 DVSS.n2867 DVSS.n2865 0.5005
R13586 DVSS.n3364 DVSS.n2868 0.5005
R13587 DVSS.n3363 DVSS.n2869 0.5005
R13588 DVSS.n2884 DVSS.n2870 0.5005
R13589 DVSS.n2885 DVSS.n2883 0.5005
R13590 DVSS.n3352 DVSS.n2886 0.5005
R13591 DVSS.n3351 DVSS.n2887 0.5005
R13592 DVSS.n2902 DVSS.n2888 0.5005
R13593 DVSS.n2903 DVSS.n2901 0.5005
R13594 DVSS.n3339 DVSS.n2904 0.5005
R13595 DVSS.n3338 DVSS.n2905 0.5005
R13596 DVSS.n2920 DVSS.n2906 0.5005
R13597 DVSS.n2921 DVSS.n2919 0.5005
R13598 DVSS.n3326 DVSS.n2922 0.5005
R13599 DVSS.n3325 DVSS.n2923 0.5005
R13600 DVSS.n2937 DVSS.n2924 0.5005
R13601 DVSS.n2938 DVSS.n2936 0.5005
R13602 DVSS.n3314 DVSS.n2939 0.5005
R13603 DVSS.n3313 DVSS.n2940 0.5005
R13604 DVSS.n2956 DVSS.n2941 0.5005
R13605 DVSS.n2957 DVSS.n2955 0.5005
R13606 DVSS.n3301 DVSS.n2958 0.5005
R13607 DVSS.n3300 DVSS.n2959 0.5005
R13608 DVSS.n2973 DVSS.n2960 0.5005
R13609 DVSS.n2974 DVSS.n2972 0.5005
R13610 DVSS.n3288 DVSS.n2975 0.5005
R13611 DVSS.n3287 DVSS.n2976 0.5005
R13612 DVSS.n2991 DVSS.n2977 0.5005
R13613 DVSS.n2992 DVSS.n2990 0.5005
R13614 DVSS.n3276 DVSS.n2993 0.5005
R13615 DVSS.n3275 DVSS.n2994 0.5005
R13616 DVSS.n2996 DVSS.n2995 0.5005
R13617 DVSS.n1786 DVSS.n1785 0.5005
R13618 DVSS.n3832 DVSS.n3831 0.5005
R13619 DVSS.n3833 DVSS.n1784 0.5005
R13620 DVSS.n3835 DVSS.n3834 0.5005
R13621 DVSS.n1782 DVSS.n1781 0.5005
R13622 DVSS.n3840 DVSS.n3839 0.5005
R13623 DVSS.n3841 DVSS.n1780 0.5005
R13624 DVSS.n3863 DVSS.n3842 0.5005
R13625 DVSS.n3862 DVSS.n3843 0.5005
R13626 DVSS.n3861 DVSS.n3844 0.5005
R13627 DVSS.n3847 DVSS.n3845 0.5005
R13628 DVSS.n3857 DVSS.n3848 0.5005
R13629 DVSS.n3856 DVSS.n3849 0.5005
R13630 DVSS.n3855 DVSS.n3850 0.5005
R13631 DVSS.n3852 DVSS.n3851 0.5005
R13632 DVSS.n2684 DVSS.n2683 0.5005
R13633 DVSS.n3864 DVSS.n3863 0.5005
R13634 DVSS.n3862 DVSS.n1779 0.5005
R13635 DVSS.n3861 DVSS.n3860 0.5005
R13636 DVSS.n3859 DVSS.n3845 0.5005
R13637 DVSS.n3858 DVSS.n3857 0.5005
R13638 DVSS.n3856 DVSS.n3846 0.5005
R13639 DVSS.n3855 DVSS.n3854 0.5005
R13640 DVSS.n1780 DVSS.n1778 0.5005
R13641 DVSS.n3839 DVSS.n3838 0.5005
R13642 DVSS.n3837 DVSS.n1782 0.5005
R13643 DVSS.n3836 DVSS.n3835 0.5005
R13644 DVSS.n1784 DVSS.n1783 0.5005
R13645 DVSS.n3831 DVSS.n3830 0.5005
R13646 DVSS.n3262 DVSS.n1786 0.5005
R13647 DVSS.n2998 DVSS.n2996 0.5005
R13648 DVSS.n3275 DVSS.n3274 0.5005
R13649 DVSS.n3277 DVSS.n3276 0.5005
R13650 DVSS.n2990 DVSS.n2987 0.5005
R13651 DVSS.n2979 DVSS.n2977 0.5005
R13652 DVSS.n3287 DVSS.n3286 0.5005
R13653 DVSS.n3289 DVSS.n3288 0.5005
R13654 DVSS.n2972 DVSS.n2969 0.5005
R13655 DVSS.n2962 DVSS.n2960 0.5005
R13656 DVSS.n3300 DVSS.n3299 0.5005
R13657 DVSS.n3302 DVSS.n3301 0.5005
R13658 DVSS.n2955 DVSS.n2952 0.5005
R13659 DVSS.n2943 DVSS.n2941 0.5005
R13660 DVSS.n3313 DVSS.n3312 0.5005
R13661 DVSS.n3315 DVSS.n3314 0.5005
R13662 DVSS.n2936 DVSS.n2933 0.5005
R13663 DVSS.n2926 DVSS.n2924 0.5005
R13664 DVSS.n3325 DVSS.n3324 0.5005
R13665 DVSS.n3327 DVSS.n3326 0.5005
R13666 DVSS.n2919 DVSS.n2916 0.5005
R13667 DVSS.n2908 DVSS.n2906 0.5005
R13668 DVSS.n3338 DVSS.n3337 0.5005
R13669 DVSS.n3340 DVSS.n3339 0.5005
R13670 DVSS.n2901 DVSS.n2898 0.5005
R13671 DVSS.n2890 DVSS.n2888 0.5005
R13672 DVSS.n3351 DVSS.n3350 0.5005
R13673 DVSS.n3353 DVSS.n3352 0.5005
R13674 DVSS.n2883 DVSS.n2880 0.5005
R13675 DVSS.n2872 DVSS.n2870 0.5005
R13676 DVSS.n3363 DVSS.n3362 0.5005
R13677 DVSS.n3365 DVSS.n3364 0.5005
R13678 DVSS.n2865 DVSS.n2862 0.5005
R13679 DVSS.n2852 DVSS.n2850 0.5005
R13680 DVSS.n3375 DVSS.n3374 0.5005
R13681 DVSS.n3377 DVSS.n3376 0.5005
R13682 DVSS.n2845 DVSS.n2842 0.5005
R13683 DVSS.n2835 DVSS.n2833 0.5005
R13684 DVSS.n3387 DVSS.n3386 0.5005
R13685 DVSS.n3389 DVSS.n3388 0.5005
R13686 DVSS.n2830 DVSS.n2827 0.5005
R13687 DVSS.n3139 DVSS.n3138 0.5005
R13688 DVSS.n2816 DVSS.n2814 0.5005
R13689 DVSS.n3403 DVSS.n3402 0.5005
R13690 DVSS.n3405 DVSS.n3404 0.5005
R13691 DVSS.n2809 DVSS.n2806 0.5005
R13692 DVSS.n2797 DVSS.n2795 0.5005
R13693 DVSS.n3415 DVSS.n3414 0.5005
R13694 DVSS.n3417 DVSS.n3416 0.5005
R13695 DVSS.n2790 DVSS.n2787 0.5005
R13696 DVSS.n2780 DVSS.n2778 0.5005
R13697 DVSS.n3427 DVSS.n3426 0.5005
R13698 DVSS.n3429 DVSS.n3428 0.5005
R13699 DVSS.n2773 DVSS.n2770 0.5005
R13700 DVSS.n2760 DVSS.n2758 0.5005
R13701 DVSS.n3439 DVSS.n3438 0.5005
R13702 DVSS.n3441 DVSS.n3440 0.5005
R13703 DVSS.n2753 DVSS.n2750 0.5005
R13704 DVSS.n2743 DVSS.n2741 0.5005
R13705 DVSS.n3451 DVSS.n3450 0.5005
R13706 DVSS.n3453 DVSS.n3452 0.5005
R13707 DVSS.n2738 DVSS.n2735 0.5005
R13708 DVSS.n3070 DVSS.n3069 0.5005
R13709 DVSS.n2725 DVSS.n2723 0.5005
R13710 DVSS.n3467 DVSS.n3466 0.5005
R13711 DVSS.n3469 DVSS.n3468 0.5005
R13712 DVSS.n2718 DVSS.n2715 0.5005
R13713 DVSS.n2707 DVSS.n2705 0.5005
R13714 DVSS.n3479 DVSS.n3478 0.5005
R13715 DVSS.n3481 DVSS.n3480 0.5005
R13716 DVSS.n2700 DVSS.n2697 0.5005
R13717 DVSS.n2690 DVSS.n2688 0.5005
R13718 DVSS.n3491 DVSS.n3490 0.5005
R13719 DVSS.n3493 DVSS.n3492 0.5005
R13720 DVSS.n2680 DVSS.n2677 0.5005
R13721 DVSS.n2682 DVSS.n2669 0.5005
R13722 DVSS.n2683 DVSS.n2670 0.5005
R13723 DVSS.n4309 DVSS.n4300 0.497977
R13724 DVSS.n4308 DVSS.n4302 0.497977
R13725 DVSS.n4307 DVSS.n4306 0.497977
R13726 DVSS.n3933 DVSS.n1705 0.497868
R13727 DVSS.n4053 DVSS.n1617 0.497868
R13728 DVSS.n4094 DVSS.n1554 0.495738
R13729 DVSS.n5795 DVSS.n5793 0.490418
R13730 DVSS.n1842 DVSS.n1696 0.477527
R13731 DVSS.n3823 DVSS.n1696 0.473227
R13732 DVSS.n2660 DVSS.n2659 0.473227
R13733 DVSS.n3787 DVSS.n3786 0.473227
R13734 DVSS.n3786 DVSS.n2631 0.473227
R13735 DVSS.n2639 DVSS.n2638 0.473227
R13736 DVSS.n3777 DVSS.n2639 0.473227
R13737 DVSS.n2618 DVSS.n2617 0.473227
R13738 DVSS.n4308 DVSS 0.469029
R13739 DVSS.n1483 DVSS.n1482 0.465755
R13740 DVSS.n4679 DVSS.n4678 0.455549
R13741 DVSS.n1572 DVSS.n1571 0.455549
R13742 DVSS.n3767 DVSS.n3766 0.455549
R13743 DVSS.n5092 DVSS.n5091 0.455549
R13744 DVSS.n3521 DVSS.n3520 0.455549
R13745 DVSS.n5062 DVSS.n1098 0.452884
R13746 DVSS.n4872 DVSS.n4871 0.452868
R13747 DVSS.n1099 DVSS.n1098 0.452744
R13748 DVSS.n950 DVSS.n949 0.4505
R13749 DVSS.n5349 DVSS.n5348 0.4505
R13750 DVSS.n5350 DVSS.n948 0.4505
R13751 DVSS.n5352 DVSS.n5351 0.4505
R13752 DVSS.n946 DVSS.n945 0.4505
R13753 DVSS.n5357 DVSS.n5356 0.4505
R13754 DVSS.n5358 DVSS.n944 0.4505
R13755 DVSS.n5360 DVSS.n5359 0.4505
R13756 DVSS.n942 DVSS.n941 0.4505
R13757 DVSS.n5365 DVSS.n5364 0.4505
R13758 DVSS.n5366 DVSS.n940 0.4505
R13759 DVSS.n5368 DVSS.n5367 0.4505
R13760 DVSS.n938 DVSS.n937 0.4505
R13761 DVSS.n5373 DVSS.n5372 0.4505
R13762 DVSS.n5374 DVSS.n936 0.4505
R13763 DVSS.n5376 DVSS.n5375 0.4505
R13764 DVSS.n934 DVSS.n933 0.4505
R13765 DVSS.n5381 DVSS.n5380 0.4505
R13766 DVSS.n5382 DVSS.n932 0.4505
R13767 DVSS.n5384 DVSS.n5383 0.4505
R13768 DVSS.n930 DVSS.n929 0.4505
R13769 DVSS.n5389 DVSS.n5388 0.4505
R13770 DVSS.n5390 DVSS.n928 0.4505
R13771 DVSS.n5392 DVSS.n5391 0.4505
R13772 DVSS.n926 DVSS.n925 0.4505
R13773 DVSS.n5397 DVSS.n5396 0.4505
R13774 DVSS.n5398 DVSS.n924 0.4505
R13775 DVSS.n5400 DVSS.n5399 0.4505
R13776 DVSS.n922 DVSS.n921 0.4505
R13777 DVSS.n5405 DVSS.n5404 0.4505
R13778 DVSS.n5406 DVSS.n920 0.4505
R13779 DVSS.n5408 DVSS.n5407 0.4505
R13780 DVSS.n918 DVSS.n917 0.4505
R13781 DVSS.n5413 DVSS.n5412 0.4505
R13782 DVSS.n5414 DVSS.n916 0.4505
R13783 DVSS.n5416 DVSS.n5415 0.4505
R13784 DVSS.n914 DVSS.n913 0.4505
R13785 DVSS.n5421 DVSS.n5420 0.4505
R13786 DVSS.n5422 DVSS.n912 0.4505
R13787 DVSS.n5424 DVSS.n5423 0.4505
R13788 DVSS.n910 DVSS.n909 0.4505
R13789 DVSS.n5429 DVSS.n5428 0.4505
R13790 DVSS.n5430 DVSS.n908 0.4505
R13791 DVSS.n5432 DVSS.n5431 0.4505
R13792 DVSS.n906 DVSS.n905 0.4505
R13793 DVSS.n5437 DVSS.n5436 0.4505
R13794 DVSS.n5438 DVSS.n904 0.4505
R13795 DVSS.n5440 DVSS.n5439 0.4505
R13796 DVSS.n902 DVSS.n901 0.4505
R13797 DVSS.n5445 DVSS.n5444 0.4505
R13798 DVSS.n5446 DVSS.n900 0.4505
R13799 DVSS.n5448 DVSS.n5447 0.4505
R13800 DVSS.n898 DVSS.n897 0.4505
R13801 DVSS.n5453 DVSS.n5452 0.4505
R13802 DVSS.n5454 DVSS.n896 0.4505
R13803 DVSS.n5456 DVSS.n5455 0.4505
R13804 DVSS.n894 DVSS.n893 0.4505
R13805 DVSS.n5461 DVSS.n5460 0.4505
R13806 DVSS.n5462 DVSS.n892 0.4505
R13807 DVSS.n5464 DVSS.n5463 0.4505
R13808 DVSS.n890 DVSS.n889 0.4505
R13809 DVSS.n5469 DVSS.n5468 0.4505
R13810 DVSS.n5470 DVSS.n888 0.4505
R13811 DVSS.n5472 DVSS.n5471 0.4505
R13812 DVSS.n886 DVSS.n885 0.4505
R13813 DVSS.n5477 DVSS.n5476 0.4505
R13814 DVSS.n5478 DVSS.n884 0.4505
R13815 DVSS.n5480 DVSS.n5479 0.4505
R13816 DVSS.n882 DVSS.n881 0.4505
R13817 DVSS.n5485 DVSS.n5484 0.4505
R13818 DVSS.n5486 DVSS.n880 0.4505
R13819 DVSS.n5488 DVSS.n5487 0.4505
R13820 DVSS.n878 DVSS.n877 0.4505
R13821 DVSS.n5493 DVSS.n5492 0.4505
R13822 DVSS.n5494 DVSS.n876 0.4505
R13823 DVSS.n5496 DVSS.n5495 0.4505
R13824 DVSS.n874 DVSS.n873 0.4505
R13825 DVSS.n5501 DVSS.n5500 0.4505
R13826 DVSS.n5502 DVSS.n872 0.4505
R13827 DVSS.n5504 DVSS.n5503 0.4505
R13828 DVSS.n870 DVSS.n869 0.4505
R13829 DVSS.n5509 DVSS.n5508 0.4505
R13830 DVSS.n5510 DVSS.n868 0.4505
R13831 DVSS.n5512 DVSS.n5511 0.4505
R13832 DVSS.n866 DVSS.n865 0.4505
R13833 DVSS.n5517 DVSS.n5516 0.4505
R13834 DVSS.n5518 DVSS.n864 0.4505
R13835 DVSS.n5520 DVSS.n5519 0.4505
R13836 DVSS.n862 DVSS.n861 0.4505
R13837 DVSS.n5525 DVSS.n5524 0.4505
R13838 DVSS.n5526 DVSS.n860 0.4505
R13839 DVSS.n5528 DVSS.n5527 0.4505
R13840 DVSS.n858 DVSS.n857 0.4505
R13841 DVSS.n5533 DVSS.n5532 0.4505
R13842 DVSS.n5535 DVSS.n5534 0.4505
R13843 DVSS.n953 DVSS.n951 0.4505
R13844 DVSS.n5346 DVSS.n950 0.4505
R13845 DVSS.n5348 DVSS.n5347 0.4505
R13846 DVSS.n948 DVSS.n947 0.4505
R13847 DVSS.n5353 DVSS.n5352 0.4505
R13848 DVSS.n5354 DVSS.n946 0.4505
R13849 DVSS.n5356 DVSS.n5355 0.4505
R13850 DVSS.n944 DVSS.n943 0.4505
R13851 DVSS.n5361 DVSS.n5360 0.4505
R13852 DVSS.n5362 DVSS.n942 0.4505
R13853 DVSS.n5364 DVSS.n5363 0.4505
R13854 DVSS.n940 DVSS.n939 0.4505
R13855 DVSS.n5369 DVSS.n5368 0.4505
R13856 DVSS.n5370 DVSS.n938 0.4505
R13857 DVSS.n5372 DVSS.n5371 0.4505
R13858 DVSS.n936 DVSS.n935 0.4505
R13859 DVSS.n5377 DVSS.n5376 0.4505
R13860 DVSS.n5378 DVSS.n934 0.4505
R13861 DVSS.n5380 DVSS.n5379 0.4505
R13862 DVSS.n932 DVSS.n931 0.4505
R13863 DVSS.n5385 DVSS.n5384 0.4505
R13864 DVSS.n5386 DVSS.n930 0.4505
R13865 DVSS.n5388 DVSS.n5387 0.4505
R13866 DVSS.n928 DVSS.n927 0.4505
R13867 DVSS.n5393 DVSS.n5392 0.4505
R13868 DVSS.n5394 DVSS.n926 0.4505
R13869 DVSS.n5396 DVSS.n5395 0.4505
R13870 DVSS.n924 DVSS.n923 0.4505
R13871 DVSS.n5401 DVSS.n5400 0.4505
R13872 DVSS.n5402 DVSS.n922 0.4505
R13873 DVSS.n5404 DVSS.n5403 0.4505
R13874 DVSS.n920 DVSS.n919 0.4505
R13875 DVSS.n5409 DVSS.n5408 0.4505
R13876 DVSS.n5410 DVSS.n918 0.4505
R13877 DVSS.n5412 DVSS.n5411 0.4505
R13878 DVSS.n916 DVSS.n915 0.4505
R13879 DVSS.n5417 DVSS.n5416 0.4505
R13880 DVSS.n5418 DVSS.n914 0.4505
R13881 DVSS.n5420 DVSS.n5419 0.4505
R13882 DVSS.n912 DVSS.n911 0.4505
R13883 DVSS.n5425 DVSS.n5424 0.4505
R13884 DVSS.n5426 DVSS.n910 0.4505
R13885 DVSS.n5428 DVSS.n5427 0.4505
R13886 DVSS.n908 DVSS.n907 0.4505
R13887 DVSS.n5433 DVSS.n5432 0.4505
R13888 DVSS.n5434 DVSS.n906 0.4505
R13889 DVSS.n5436 DVSS.n5435 0.4505
R13890 DVSS.n904 DVSS.n903 0.4505
R13891 DVSS.n5441 DVSS.n5440 0.4505
R13892 DVSS.n5442 DVSS.n902 0.4505
R13893 DVSS.n5444 DVSS.n5443 0.4505
R13894 DVSS.n900 DVSS.n899 0.4505
R13895 DVSS.n5449 DVSS.n5448 0.4505
R13896 DVSS.n5450 DVSS.n898 0.4505
R13897 DVSS.n5452 DVSS.n5451 0.4505
R13898 DVSS.n896 DVSS.n895 0.4505
R13899 DVSS.n5457 DVSS.n5456 0.4505
R13900 DVSS.n5458 DVSS.n894 0.4505
R13901 DVSS.n5460 DVSS.n5459 0.4505
R13902 DVSS.n892 DVSS.n891 0.4505
R13903 DVSS.n5465 DVSS.n5464 0.4505
R13904 DVSS.n5466 DVSS.n890 0.4505
R13905 DVSS.n5468 DVSS.n5467 0.4505
R13906 DVSS.n888 DVSS.n887 0.4505
R13907 DVSS.n5473 DVSS.n5472 0.4505
R13908 DVSS.n5474 DVSS.n886 0.4505
R13909 DVSS.n5476 DVSS.n5475 0.4505
R13910 DVSS.n884 DVSS.n883 0.4505
R13911 DVSS.n5481 DVSS.n5480 0.4505
R13912 DVSS.n5482 DVSS.n882 0.4505
R13913 DVSS.n5484 DVSS.n5483 0.4505
R13914 DVSS.n880 DVSS.n879 0.4505
R13915 DVSS.n5489 DVSS.n5488 0.4505
R13916 DVSS.n5490 DVSS.n878 0.4505
R13917 DVSS.n5492 DVSS.n5491 0.4505
R13918 DVSS.n876 DVSS.n875 0.4505
R13919 DVSS.n5497 DVSS.n5496 0.4505
R13920 DVSS.n5498 DVSS.n874 0.4505
R13921 DVSS.n5500 DVSS.n5499 0.4505
R13922 DVSS.n872 DVSS.n871 0.4505
R13923 DVSS.n5505 DVSS.n5504 0.4505
R13924 DVSS.n5506 DVSS.n870 0.4505
R13925 DVSS.n5508 DVSS.n5507 0.4505
R13926 DVSS.n868 DVSS.n867 0.4505
R13927 DVSS.n5513 DVSS.n5512 0.4505
R13928 DVSS.n5514 DVSS.n866 0.4505
R13929 DVSS.n5516 DVSS.n5515 0.4505
R13930 DVSS.n864 DVSS.n863 0.4505
R13931 DVSS.n5521 DVSS.n5520 0.4505
R13932 DVSS.n5522 DVSS.n862 0.4505
R13933 DVSS.n5524 DVSS.n5523 0.4505
R13934 DVSS.n860 DVSS.n859 0.4505
R13935 DVSS.n5529 DVSS.n5528 0.4505
R13936 DVSS.n5530 DVSS.n858 0.4505
R13937 DVSS.n5532 DVSS.n5531 0.4505
R13938 DVSS.n5536 DVSS.n5535 0.4505
R13939 DVSS.n4686 DVSS.n4677 0.4505
R13940 DVSS.n4685 DVSS.n4684 0.4505
R13941 DVSS.n4380 DVSS.n4342 0.4505
R13942 DVSS.n4382 DVSS.n4381 0.4505
R13943 DVSS.n4340 DVSS.n4339 0.4505
R13944 DVSS.n4387 DVSS.n4386 0.4505
R13945 DVSS.n4388 DVSS.n4338 0.4505
R13946 DVSS.n4390 DVSS.n4389 0.4505
R13947 DVSS.n4333 DVSS.n4332 0.4505
R13948 DVSS.n4402 DVSS.n4401 0.4505
R13949 DVSS.n4403 DVSS.n4330 0.4505
R13950 DVSS.n4499 DVSS.n4498 0.4505
R13951 DVSS.n4497 DVSS.n4331 0.4505
R13952 DVSS.n4496 DVSS.n4495 0.4505
R13953 DVSS.n4405 DVSS.n4404 0.4505
R13954 DVSS.n4491 DVSS.n4490 0.4505
R13955 DVSS.n4489 DVSS.n4411 0.4505
R13956 DVSS.n4488 DVSS.n4487 0.4505
R13957 DVSS.n4413 DVSS.n4412 0.4505
R13958 DVSS.n4420 DVSS.n4418 0.4505
R13959 DVSS.n4479 DVSS.n4478 0.4505
R13960 DVSS.n4477 DVSS.n4419 0.4505
R13961 DVSS.n4476 DVSS.n4475 0.4505
R13962 DVSS.n4422 DVSS.n4421 0.4505
R13963 DVSS.n4439 DVSS.n4437 0.4505
R13964 DVSS.n4466 DVSS.n4465 0.4505
R13965 DVSS.n4464 DVSS.n4438 0.4505
R13966 DVSS.n4463 DVSS.n4462 0.4505
R13967 DVSS.n4441 DVSS.n4440 0.4505
R13968 DVSS.n4458 DVSS.n4457 0.4505
R13969 DVSS.n4456 DVSS.n4443 0.4505
R13970 DVSS.n4455 DVSS.n4454 0.4505
R13971 DVSS.n4445 DVSS.n4444 0.4505
R13972 DVSS.n1445 DVSS.n1444 0.4505
R13973 DVSS.n4518 DVSS.n4517 0.4505
R13974 DVSS.n4519 DVSS.n1443 0.4505
R13975 DVSS.n4521 DVSS.n4520 0.4505
R13976 DVSS.n1436 DVSS.n1435 0.4505
R13977 DVSS.n4531 DVSS.n4530 0.4505
R13978 DVSS.n4532 DVSS.n1434 0.4505
R13979 DVSS.n4534 DVSS.n4533 0.4505
R13980 DVSS.n1432 DVSS.n1431 0.4505
R13981 DVSS.n4540 DVSS.n4539 0.4505
R13982 DVSS.n4541 DVSS.n1430 0.4505
R13983 DVSS.n4543 DVSS.n4542 0.4505
R13984 DVSS.n1425 DVSS.n1424 0.4505
R13985 DVSS.n4557 DVSS.n4556 0.4505
R13986 DVSS.n4558 DVSS.n1422 0.4505
R13987 DVSS.n4561 DVSS.n4560 0.4505
R13988 DVSS.n4559 DVSS.n1423 0.4505
R13989 DVSS.n1415 DVSS.n1414 0.4505
R13990 DVSS.n4572 DVSS.n4571 0.4505
R13991 DVSS.n4573 DVSS.n1413 0.4505
R13992 DVSS.n4575 DVSS.n4574 0.4505
R13993 DVSS.n1411 DVSS.n1410 0.4505
R13994 DVSS.n4580 DVSS.n4579 0.4505
R13995 DVSS.n4581 DVSS.n1409 0.4505
R13996 DVSS.n4583 DVSS.n4582 0.4505
R13997 DVSS.n1404 DVSS.n1403 0.4505
R13998 DVSS.n4595 DVSS.n4594 0.4505
R13999 DVSS.n4596 DVSS.n1401 0.4505
R14000 DVSS.n4747 DVSS.n4746 0.4505
R14001 DVSS.n4745 DVSS.n1402 0.4505
R14002 DVSS.n4744 DVSS.n4743 0.4505
R14003 DVSS.n4598 DVSS.n4597 0.4505
R14004 DVSS.n4739 DVSS.n4738 0.4505
R14005 DVSS.n4737 DVSS.n4604 0.4505
R14006 DVSS.n4736 DVSS.n4735 0.4505
R14007 DVSS.n4606 DVSS.n4605 0.4505
R14008 DVSS.n4613 DVSS.n4611 0.4505
R14009 DVSS.n4727 DVSS.n4726 0.4505
R14010 DVSS.n4725 DVSS.n4612 0.4505
R14011 DVSS.n4724 DVSS.n4723 0.4505
R14012 DVSS.n4615 DVSS.n4614 0.4505
R14013 DVSS.n4632 DVSS.n4630 0.4505
R14014 DVSS.n4714 DVSS.n4713 0.4505
R14015 DVSS.n4712 DVSS.n4631 0.4505
R14016 DVSS.n4711 DVSS.n4710 0.4505
R14017 DVSS.n4634 DVSS.n4633 0.4505
R14018 DVSS.n4671 DVSS.n4670 0.4505
R14019 DVSS.n4672 DVSS.n4668 0.4505
R14020 DVSS.n4702 DVSS.n4701 0.4505
R14021 DVSS.n4700 DVSS.n4669 0.4505
R14022 DVSS.n4699 DVSS.n4698 0.4505
R14023 DVSS.n4674 DVSS.n4673 0.4505
R14024 DVSS.n4694 DVSS.n4693 0.4505
R14025 DVSS.n4692 DVSS.n4676 0.4505
R14026 DVSS.n4691 DVSS.n4690 0.4505
R14027 DVSS.n4689 DVSS.n4687 0.4505
R14028 DVSS.n4682 DVSS.n4680 0.4505
R14029 DVSS.n4684 DVSS.n4683 0.4505
R14030 DVSS.n4681 DVSS.n4677 0.4505
R14031 DVSS.n4378 DVSS.n4377 0.4505
R14032 DVSS.n4372 DVSS.n4342 0.4505
R14033 DVSS.n4383 DVSS.n4382 0.4505
R14034 DVSS.n4384 DVSS.n4340 0.4505
R14035 DVSS.n4386 DVSS.n4385 0.4505
R14036 DVSS.n4338 DVSS.n4336 0.4505
R14037 DVSS.n4391 DVSS.n4390 0.4505
R14038 DVSS.n4334 DVSS.n4333 0.4505
R14039 DVSS.n4401 DVSS.n4400 0.4505
R14040 DVSS.n4330 DVSS.n4328 0.4505
R14041 DVSS.n4500 DVSS.n4499 0.4505
R14042 DVSS.n4406 DVSS.n4331 0.4505
R14043 DVSS.n4495 DVSS.n4494 0.4505
R14044 DVSS.n4493 DVSS.n4405 0.4505
R14045 DVSS.n4492 DVSS.n4491 0.4505
R14046 DVSS.n4411 DVSS.n4410 0.4505
R14047 DVSS.n4487 DVSS.n4486 0.4505
R14048 DVSS.n4485 DVSS.n4413 0.4505
R14049 DVSS.n4418 DVSS.n4414 0.4505
R14050 DVSS.n4480 DVSS.n4479 0.4505
R14051 DVSS.n4423 DVSS.n4419 0.4505
R14052 DVSS.n4475 DVSS.n4474 0.4505
R14053 DVSS.n4425 DVSS.n4422 0.4505
R14054 DVSS.n4437 DVSS.n4435 0.4505
R14055 DVSS.n4467 DVSS.n4466 0.4505
R14056 DVSS.n4438 DVSS.n4436 0.4505
R14057 DVSS.n4462 DVSS.n4461 0.4505
R14058 DVSS.n4460 DVSS.n4441 0.4505
R14059 DVSS.n4459 DVSS.n4458 0.4505
R14060 DVSS.n4443 DVSS.n4442 0.4505
R14061 DVSS.n4454 DVSS.n4453 0.4505
R14062 DVSS.n4446 DVSS.n4445 0.4505
R14063 DVSS.n4448 DVSS.n1445 0.4505
R14064 DVSS.n4517 DVSS.n4516 0.4505
R14065 DVSS.n1443 DVSS.n1441 0.4505
R14066 DVSS.n4522 DVSS.n4521 0.4505
R14067 DVSS.n1437 DVSS.n1436 0.4505
R14068 DVSS.n4530 DVSS.n4529 0.4505
R14069 DVSS.n1434 DVSS.n1433 0.4505
R14070 DVSS.n4535 DVSS.n4534 0.4505
R14071 DVSS.n4536 DVSS.n1432 0.4505
R14072 DVSS.n4539 DVSS.n4538 0.4505
R14073 DVSS.n4537 DVSS.n1430 0.4505
R14074 DVSS.n4544 DVSS.n4543 0.4505
R14075 DVSS.n4545 DVSS.n1425 0.4505
R14076 DVSS.n4556 DVSS.n4555 0.4505
R14077 DVSS.n1422 DVSS.n1420 0.4505
R14078 DVSS.n4562 DVSS.n4561 0.4505
R14079 DVSS.n1423 DVSS.n1416 0.4505
R14080 DVSS.n4569 DVSS.n1415 0.4505
R14081 DVSS.n4571 DVSS.n4570 0.4505
R14082 DVSS.n1413 DVSS.n1412 0.4505
R14083 DVSS.n4576 DVSS.n4575 0.4505
R14084 DVSS.n4577 DVSS.n1411 0.4505
R14085 DVSS.n4579 DVSS.n4578 0.4505
R14086 DVSS.n1409 DVSS.n1407 0.4505
R14087 DVSS.n4584 DVSS.n4583 0.4505
R14088 DVSS.n1405 DVSS.n1404 0.4505
R14089 DVSS.n4594 DVSS.n4593 0.4505
R14090 DVSS.n1401 DVSS.n1399 0.4505
R14091 DVSS.n4748 DVSS.n4747 0.4505
R14092 DVSS.n4599 DVSS.n1402 0.4505
R14093 DVSS.n4743 DVSS.n4742 0.4505
R14094 DVSS.n4741 DVSS.n4598 0.4505
R14095 DVSS.n4740 DVSS.n4739 0.4505
R14096 DVSS.n4604 DVSS.n4603 0.4505
R14097 DVSS.n4735 DVSS.n4734 0.4505
R14098 DVSS.n4733 DVSS.n4606 0.4505
R14099 DVSS.n4611 DVSS.n4607 0.4505
R14100 DVSS.n4728 DVSS.n4727 0.4505
R14101 DVSS.n4616 DVSS.n4612 0.4505
R14102 DVSS.n4723 DVSS.n4722 0.4505
R14103 DVSS.n4618 DVSS.n4615 0.4505
R14104 DVSS.n4630 DVSS.n4628 0.4505
R14105 DVSS.n4715 DVSS.n4714 0.4505
R14106 DVSS.n4631 DVSS.n4629 0.4505
R14107 DVSS.n4710 DVSS.n4709 0.4505
R14108 DVSS.n4708 DVSS.n4634 0.4505
R14109 DVSS.n4670 DVSS.n4640 0.4505
R14110 DVSS.n4668 DVSS.n4663 0.4505
R14111 DVSS.n4703 DVSS.n4702 0.4505
R14112 DVSS.n4669 DVSS.n4667 0.4505
R14113 DVSS.n4698 DVSS.n4697 0.4505
R14114 DVSS.n4696 DVSS.n4674 0.4505
R14115 DVSS.n4695 DVSS.n4694 0.4505
R14116 DVSS.n4676 DVSS.n4675 0.4505
R14117 DVSS.n4690 DVSS.n1358 0.4505
R14118 DVSS.n4689 DVSS.n4688 0.4505
R14119 DVSS.n3765 DVSS.n3764 0.4505
R14120 DVSS.n3526 DVSS.n3525 0.4505
R14121 DVSS.n3746 DVSS.n3745 0.4505
R14122 DVSS.n3748 DVSS.n3747 0.4505
R14123 DVSS.n3744 DVSS.n3539 0.4505
R14124 DVSS.n3743 DVSS.n3742 0.4505
R14125 DVSS.n3541 DVSS.n3540 0.4505
R14126 DVSS.n3738 DVSS.n3737 0.4505
R14127 DVSS.n3736 DVSS.n3543 0.4505
R14128 DVSS.n3735 DVSS.n3734 0.4505
R14129 DVSS.n3545 DVSS.n3544 0.4505
R14130 DVSS.n3730 DVSS.n3729 0.4505
R14131 DVSS.n3728 DVSS.n3547 0.4505
R14132 DVSS.n3727 DVSS.n3726 0.4505
R14133 DVSS.n3549 DVSS.n3548 0.4505
R14134 DVSS.n3722 DVSS.n3721 0.4505
R14135 DVSS.n3720 DVSS.n3551 0.4505
R14136 DVSS.n3719 DVSS.n3718 0.4505
R14137 DVSS.n3553 DVSS.n3552 0.4505
R14138 DVSS.n3714 DVSS.n3713 0.4505
R14139 DVSS.n3712 DVSS.n3555 0.4505
R14140 DVSS.n3711 DVSS.n3710 0.4505
R14141 DVSS.n3557 DVSS.n3556 0.4505
R14142 DVSS.n3706 DVSS.n3705 0.4505
R14143 DVSS.n3704 DVSS.n3559 0.4505
R14144 DVSS.n3703 DVSS.n3702 0.4505
R14145 DVSS.n3561 DVSS.n3560 0.4505
R14146 DVSS.n3698 DVSS.n3697 0.4505
R14147 DVSS.n3696 DVSS.n3563 0.4505
R14148 DVSS.n3695 DVSS.n3694 0.4505
R14149 DVSS.n3565 DVSS.n3564 0.4505
R14150 DVSS.n3690 DVSS.n3689 0.4505
R14151 DVSS.n3688 DVSS.n3567 0.4505
R14152 DVSS.n3687 DVSS.n3686 0.4505
R14153 DVSS.n3569 DVSS.n3568 0.4505
R14154 DVSS.n3682 DVSS.n3681 0.4505
R14155 DVSS.n3680 DVSS.n3571 0.4505
R14156 DVSS.n3679 DVSS.n3678 0.4505
R14157 DVSS.n3573 DVSS.n3572 0.4505
R14158 DVSS.n3674 DVSS.n3673 0.4505
R14159 DVSS.n3672 DVSS.n3575 0.4505
R14160 DVSS.n3671 DVSS.n3670 0.4505
R14161 DVSS.n3577 DVSS.n3576 0.4505
R14162 DVSS.n3666 DVSS.n3665 0.4505
R14163 DVSS.n3664 DVSS.n3579 0.4505
R14164 DVSS.n3663 DVSS.n3662 0.4505
R14165 DVSS.n3581 DVSS.n3580 0.4505
R14166 DVSS.n3658 DVSS.n3657 0.4505
R14167 DVSS.n3656 DVSS.n3583 0.4505
R14168 DVSS.n3655 DVSS.n3654 0.4505
R14169 DVSS.n3585 DVSS.n3584 0.4505
R14170 DVSS.n3650 DVSS.n3649 0.4505
R14171 DVSS.n3648 DVSS.n3587 0.4505
R14172 DVSS.n3647 DVSS.n3646 0.4505
R14173 DVSS.n3589 DVSS.n3588 0.4505
R14174 DVSS.n3642 DVSS.n3641 0.4505
R14175 DVSS.n3640 DVSS.n3591 0.4505
R14176 DVSS.n3639 DVSS.n3638 0.4505
R14177 DVSS.n3593 DVSS.n3592 0.4505
R14178 DVSS.n3634 DVSS.n3633 0.4505
R14179 DVSS.n3632 DVSS.n3595 0.4505
R14180 DVSS.n3631 DVSS.n3630 0.4505
R14181 DVSS.n3597 DVSS.n3596 0.4505
R14182 DVSS.n3626 DVSS.n3625 0.4505
R14183 DVSS.n3624 DVSS.n3599 0.4505
R14184 DVSS.n3623 DVSS.n3622 0.4505
R14185 DVSS.n3601 DVSS.n3600 0.4505
R14186 DVSS.n3618 DVSS.n3617 0.4505
R14187 DVSS.n3616 DVSS.n3603 0.4505
R14188 DVSS.n3615 DVSS.n3614 0.4505
R14189 DVSS.n3605 DVSS.n3604 0.4505
R14190 DVSS.n3610 DVSS.n3609 0.4505
R14191 DVSS.n3608 DVSS.n3607 0.4505
R14192 DVSS.n1570 DVSS.n1569 0.4505
R14193 DVSS.n1578 DVSS.n1577 0.4505
R14194 DVSS.n1579 DVSS.n1568 0.4505
R14195 DVSS.n1581 DVSS.n1580 0.4505
R14196 DVSS.n1566 DVSS.n1565 0.4505
R14197 DVSS.n1586 DVSS.n1585 0.4505
R14198 DVSS.n1587 DVSS.n1564 0.4505
R14199 DVSS.n1589 DVSS.n1588 0.4505
R14200 DVSS.n1562 DVSS.n1561 0.4505
R14201 DVSS.n1594 DVSS.n1593 0.4505
R14202 DVSS.n1595 DVSS.n1559 0.4505
R14203 DVSS.n4089 DVSS.n4088 0.4505
R14204 DVSS.n4087 DVSS.n1560 0.4505
R14205 DVSS.n4086 DVSS.n4085 0.4505
R14206 DVSS.n1597 DVSS.n1596 0.4505
R14207 DVSS.n4081 DVSS.n4080 0.4505
R14208 DVSS.n4079 DVSS.n1599 0.4505
R14209 DVSS.n4078 DVSS.n4077 0.4505
R14210 DVSS.n1601 DVSS.n1600 0.4505
R14211 DVSS.n4073 DVSS.n4072 0.4505
R14212 DVSS.n4071 DVSS.n1603 0.4505
R14213 DVSS.n4070 DVSS.n4069 0.4505
R14214 DVSS.n1605 DVSS.n1604 0.4505
R14215 DVSS.n4065 DVSS.n4064 0.4505
R14216 DVSS.n4063 DVSS.n1607 0.4505
R14217 DVSS.n4062 DVSS.n4061 0.4505
R14218 DVSS.n1609 DVSS.n1608 0.4505
R14219 DVSS.n2649 DVSS.n2648 0.4505
R14220 DVSS.n1858 DVSS.n1857 0.4505
R14221 DVSS.n2282 DVSS.n2281 0.4505
R14222 DVSS.n2284 DVSS.n2283 0.4505
R14223 DVSS.n2274 DVSS.n2273 0.4505
R14224 DVSS.n2291 DVSS.n2290 0.4505
R14225 DVSS.n2292 DVSS.n2272 0.4505
R14226 DVSS.n2294 DVSS.n2293 0.4505
R14227 DVSS.n1881 DVSS.n1879 0.4505
R14228 DVSS.n2581 DVSS.n2580 0.4505
R14229 DVSS.n2579 DVSS.n1880 0.4505
R14230 DVSS.n2578 DVSS.n2577 0.4505
R14231 DVSS.n1883 DVSS.n1882 0.4505
R14232 DVSS.n2259 DVSS.n2258 0.4505
R14233 DVSS.n1908 DVSS.n1906 0.4505
R14234 DVSS.n2563 DVSS.n2562 0.4505
R14235 DVSS.n2561 DVSS.n1907 0.4505
R14236 DVSS.n2560 DVSS.n2559 0.4505
R14237 DVSS.n1910 DVSS.n1909 0.4505
R14238 DVSS.n2530 DVSS.n2529 0.4505
R14239 DVSS.n2528 DVSS.n2314 0.4505
R14240 DVSS.n2527 DVSS.n2526 0.4505
R14241 DVSS.n2316 DVSS.n2315 0.4505
R14242 DVSS.n2356 DVSS.n2355 0.4505
R14243 DVSS.n2357 DVSS.n2354 0.4505
R14244 DVSS.n2359 DVSS.n2358 0.4505
R14245 DVSS.n2344 DVSS.n2343 0.4505
R14246 DVSS.n2374 DVSS.n2373 0.4505
R14247 DVSS.n2375 DVSS.n2341 0.4505
R14248 DVSS.n2509 DVSS.n2508 0.4505
R14249 DVSS.n2507 DVSS.n2342 0.4505
R14250 DVSS.n2506 DVSS.n2505 0.4505
R14251 DVSS.n2470 DVSS.n2376 0.4505
R14252 DVSS.n2469 DVSS.n2378 0.4505
R14253 DVSS.n2381 DVSS.n2377 0.4505
R14254 DVSS.n2465 DVSS.n2464 0.4505
R14255 DVSS.n2463 DVSS.n2380 0.4505
R14256 DVSS.n2462 DVSS.n2461 0.4505
R14257 DVSS.n2383 DVSS.n2382 0.4505
R14258 DVSS.n2457 DVSS.n2456 0.4505
R14259 DVSS.n2455 DVSS.n2385 0.4505
R14260 DVSS.n2454 DVSS.n2453 0.4505
R14261 DVSS.n2387 DVSS.n2386 0.4505
R14262 DVSS.n2449 DVSS.n2448 0.4505
R14263 DVSS.n2447 DVSS.n2389 0.4505
R14264 DVSS.n2446 DVSS.n2445 0.4505
R14265 DVSS.n2391 DVSS.n2390 0.4505
R14266 DVSS.n2441 DVSS.n2440 0.4505
R14267 DVSS.n2439 DVSS.n2393 0.4505
R14268 DVSS.n2438 DVSS.n2437 0.4505
R14269 DVSS.n2395 DVSS.n2394 0.4505
R14270 DVSS.n2433 DVSS.n2432 0.4505
R14271 DVSS.n2431 DVSS.n2397 0.4505
R14272 DVSS.n2430 DVSS.n2429 0.4505
R14273 DVSS.n2399 DVSS.n2398 0.4505
R14274 DVSS.n2425 DVSS.n2424 0.4505
R14275 DVSS.n2423 DVSS.n2401 0.4505
R14276 DVSS.n2422 DVSS.n2421 0.4505
R14277 DVSS.n2403 DVSS.n2402 0.4505
R14278 DVSS.n2417 DVSS.n2416 0.4505
R14279 DVSS.n2415 DVSS.n2405 0.4505
R14280 DVSS.n2414 DVSS.n2413 0.4505
R14281 DVSS.n2407 DVSS.n2406 0.4505
R14282 DVSS.n2409 DVSS.n2408 0.4505
R14283 DVSS.n2612 DVSS.n2611 0.4505
R14284 DVSS.n2610 DVSS.n1851 0.4505
R14285 DVSS.n2609 DVSS.n2608 0.4505
R14286 DVSS.n1853 DVSS.n1852 0.4505
R14287 DVSS.n2604 DVSS.n2603 0.4505
R14288 DVSS.n2602 DVSS.n1856 0.4505
R14289 DVSS.n2601 DVSS.n2600 0.4505
R14290 DVSS.n2091 DVSS.n2090 0.4505
R14291 DVSS.n2095 DVSS.n2094 0.4505
R14292 DVSS.n2096 DVSS.n2089 0.4505
R14293 DVSS.n2098 DVSS.n2097 0.4505
R14294 DVSS.n2087 DVSS.n2086 0.4505
R14295 DVSS.n2103 DVSS.n2102 0.4505
R14296 DVSS.n2104 DVSS.n2085 0.4505
R14297 DVSS.n2106 DVSS.n2105 0.4505
R14298 DVSS.n2083 DVSS.n2082 0.4505
R14299 DVSS.n2111 DVSS.n2110 0.4505
R14300 DVSS.n2112 DVSS.n2081 0.4505
R14301 DVSS.n2114 DVSS.n2113 0.4505
R14302 DVSS.n2079 DVSS.n2078 0.4505
R14303 DVSS.n2119 DVSS.n2118 0.4505
R14304 DVSS.n2120 DVSS.n2077 0.4505
R14305 DVSS.n2122 DVSS.n2121 0.4505
R14306 DVSS.n2075 DVSS.n2074 0.4505
R14307 DVSS.n2127 DVSS.n2126 0.4505
R14308 DVSS.n2128 DVSS.n2073 0.4505
R14309 DVSS.n2130 DVSS.n2129 0.4505
R14310 DVSS.n2071 DVSS.n2070 0.4505
R14311 DVSS.n2135 DVSS.n2134 0.4505
R14312 DVSS.n2136 DVSS.n2069 0.4505
R14313 DVSS.n2138 DVSS.n2137 0.4505
R14314 DVSS.n2066 DVSS.n2065 0.4505
R14315 DVSS.n2143 DVSS.n2142 0.4505
R14316 DVSS.n2144 DVSS.n2064 0.4505
R14317 DVSS.n2020 DVSS.n2019 0.4505
R14318 DVSS.n1968 DVSS.n1967 0.4505
R14319 DVSS.n2025 DVSS.n2024 0.4505
R14320 DVSS.n2026 DVSS.n1964 0.4505
R14321 DVSS.n2225 DVSS.n2224 0.4505
R14322 DVSS.n2223 DVSS.n1966 0.4505
R14323 DVSS.n2222 DVSS.n2221 0.4505
R14324 DVSS.n2028 DVSS.n2027 0.4505
R14325 DVSS.n2217 DVSS.n2216 0.4505
R14326 DVSS.n2215 DVSS.n2030 0.4505
R14327 DVSS.n2214 DVSS.n2213 0.4505
R14328 DVSS.n2032 DVSS.n2031 0.4505
R14329 DVSS.n2209 DVSS.n2208 0.4505
R14330 DVSS.n2207 DVSS.n2034 0.4505
R14331 DVSS.n2206 DVSS.n2205 0.4505
R14332 DVSS.n2036 DVSS.n2035 0.4505
R14333 DVSS.n2201 DVSS.n2200 0.4505
R14334 DVSS.n2199 DVSS.n2038 0.4505
R14335 DVSS.n2198 DVSS.n2197 0.4505
R14336 DVSS.n2040 DVSS.n2039 0.4505
R14337 DVSS.n2193 DVSS.n2192 0.4505
R14338 DVSS.n2191 DVSS.n2042 0.4505
R14339 DVSS.n2190 DVSS.n2189 0.4505
R14340 DVSS.n2044 DVSS.n2043 0.4505
R14341 DVSS.n2185 DVSS.n2184 0.4505
R14342 DVSS.n2183 DVSS.n2046 0.4505
R14343 DVSS.n2182 DVSS.n2181 0.4505
R14344 DVSS.n2048 DVSS.n2047 0.4505
R14345 DVSS.n2177 DVSS.n2176 0.4505
R14346 DVSS.n2175 DVSS.n2050 0.4505
R14347 DVSS.n2174 DVSS.n2173 0.4505
R14348 DVSS.n2052 DVSS.n2051 0.4505
R14349 DVSS.n2169 DVSS.n2168 0.4505
R14350 DVSS.n2167 DVSS.n2054 0.4505
R14351 DVSS.n2166 DVSS.n2165 0.4505
R14352 DVSS.n2056 DVSS.n2055 0.4505
R14353 DVSS.n2161 DVSS.n2160 0.4505
R14354 DVSS.n2159 DVSS.n2058 0.4505
R14355 DVSS.n2158 DVSS.n2157 0.4505
R14356 DVSS.n2060 DVSS.n2059 0.4505
R14357 DVSS.n2153 DVSS.n2152 0.4505
R14358 DVSS.n2151 DVSS.n2062 0.4505
R14359 DVSS.n2150 DVSS.n2149 0.4505
R14360 DVSS.n2147 DVSS.n2063 0.4505
R14361 DVSS.n2146 DVSS.n2145 0.4505
R14362 DVSS.n2067 DVSS.n2064 0.4505
R14363 DVSS.n1971 DVSS.n1970 0.4505
R14364 DVSS.n2142 DVSS.n2141 0.4505
R14365 DVSS.n2140 DVSS.n2066 0.4505
R14366 DVSS.n2139 DVSS.n2138 0.4505
R14367 DVSS.n2069 DVSS.n2068 0.4505
R14368 DVSS.n2134 DVSS.n2133 0.4505
R14369 DVSS.n2132 DVSS.n2071 0.4505
R14370 DVSS.n2131 DVSS.n2130 0.4505
R14371 DVSS.n2073 DVSS.n2072 0.4505
R14372 DVSS.n2126 DVSS.n2125 0.4505
R14373 DVSS.n2124 DVSS.n2075 0.4505
R14374 DVSS.n2123 DVSS.n2122 0.4505
R14375 DVSS.n2077 DVSS.n2076 0.4505
R14376 DVSS.n2118 DVSS.n2117 0.4505
R14377 DVSS.n2116 DVSS.n2079 0.4505
R14378 DVSS.n2115 DVSS.n2114 0.4505
R14379 DVSS.n2081 DVSS.n2080 0.4505
R14380 DVSS.n2110 DVSS.n2109 0.4505
R14381 DVSS.n2108 DVSS.n2083 0.4505
R14382 DVSS.n2107 DVSS.n2106 0.4505
R14383 DVSS.n2085 DVSS.n2084 0.4505
R14384 DVSS.n2102 DVSS.n2101 0.4505
R14385 DVSS.n2100 DVSS.n2087 0.4505
R14386 DVSS.n2099 DVSS.n2098 0.4505
R14387 DVSS.n2089 DVSS.n2088 0.4505
R14388 DVSS.n2094 DVSS.n2093 0.4505
R14389 DVSS.n2021 DVSS.n2020 0.4505
R14390 DVSS.n2022 DVSS.n1968 0.4505
R14391 DVSS.n2024 DVSS.n2023 0.4505
R14392 DVSS.n1964 DVSS.n1960 0.4505
R14393 DVSS.n2226 DVSS.n2225 0.4505
R14394 DVSS.n1966 DVSS.n1965 0.4505
R14395 DVSS.n2221 DVSS.n2220 0.4505
R14396 DVSS.n2219 DVSS.n2028 0.4505
R14397 DVSS.n2218 DVSS.n2217 0.4505
R14398 DVSS.n2030 DVSS.n2029 0.4505
R14399 DVSS.n2213 DVSS.n2212 0.4505
R14400 DVSS.n2211 DVSS.n2032 0.4505
R14401 DVSS.n2210 DVSS.n2209 0.4505
R14402 DVSS.n2034 DVSS.n2033 0.4505
R14403 DVSS.n2205 DVSS.n2204 0.4505
R14404 DVSS.n2203 DVSS.n2036 0.4505
R14405 DVSS.n2202 DVSS.n2201 0.4505
R14406 DVSS.n2038 DVSS.n2037 0.4505
R14407 DVSS.n2197 DVSS.n2196 0.4505
R14408 DVSS.n2195 DVSS.n2040 0.4505
R14409 DVSS.n2194 DVSS.n2193 0.4505
R14410 DVSS.n2042 DVSS.n2041 0.4505
R14411 DVSS.n2189 DVSS.n2188 0.4505
R14412 DVSS.n2187 DVSS.n2044 0.4505
R14413 DVSS.n2186 DVSS.n2185 0.4505
R14414 DVSS.n2046 DVSS.n2045 0.4505
R14415 DVSS.n2181 DVSS.n2180 0.4505
R14416 DVSS.n2179 DVSS.n2048 0.4505
R14417 DVSS.n2178 DVSS.n2177 0.4505
R14418 DVSS.n2050 DVSS.n2049 0.4505
R14419 DVSS.n2173 DVSS.n2172 0.4505
R14420 DVSS.n2171 DVSS.n2052 0.4505
R14421 DVSS.n2170 DVSS.n2169 0.4505
R14422 DVSS.n2054 DVSS.n2053 0.4505
R14423 DVSS.n2165 DVSS.n2164 0.4505
R14424 DVSS.n2163 DVSS.n2056 0.4505
R14425 DVSS.n2162 DVSS.n2161 0.4505
R14426 DVSS.n2058 DVSS.n2057 0.4505
R14427 DVSS.n2157 DVSS.n2156 0.4505
R14428 DVSS.n2155 DVSS.n2060 0.4505
R14429 DVSS.n2154 DVSS.n2153 0.4505
R14430 DVSS.n2062 DVSS.n2061 0.4505
R14431 DVSS.n2149 DVSS.n2148 0.4505
R14432 DVSS.n2147 DVSS.n1529 0.4505
R14433 DVSS.n2146 DVSS.n1534 0.4505
R14434 DVSS.n2411 DVSS.n2407 0.4505
R14435 DVSS.n2413 DVSS.n2412 0.4505
R14436 DVSS.n2405 DVSS.n2404 0.4505
R14437 DVSS.n2418 DVSS.n2417 0.4505
R14438 DVSS.n2419 DVSS.n2403 0.4505
R14439 DVSS.n2421 DVSS.n2420 0.4505
R14440 DVSS.n2401 DVSS.n2400 0.4505
R14441 DVSS.n2426 DVSS.n2425 0.4505
R14442 DVSS.n2427 DVSS.n2399 0.4505
R14443 DVSS.n2429 DVSS.n2428 0.4505
R14444 DVSS.n2397 DVSS.n2396 0.4505
R14445 DVSS.n2434 DVSS.n2433 0.4505
R14446 DVSS.n2435 DVSS.n2395 0.4505
R14447 DVSS.n2437 DVSS.n2436 0.4505
R14448 DVSS.n2393 DVSS.n2392 0.4505
R14449 DVSS.n2442 DVSS.n2441 0.4505
R14450 DVSS.n2443 DVSS.n2391 0.4505
R14451 DVSS.n2445 DVSS.n2444 0.4505
R14452 DVSS.n2389 DVSS.n2388 0.4505
R14453 DVSS.n2450 DVSS.n2449 0.4505
R14454 DVSS.n2451 DVSS.n2387 0.4505
R14455 DVSS.n2453 DVSS.n2452 0.4505
R14456 DVSS.n2385 DVSS.n2384 0.4505
R14457 DVSS.n2458 DVSS.n2457 0.4505
R14458 DVSS.n2459 DVSS.n2383 0.4505
R14459 DVSS.n2461 DVSS.n2460 0.4505
R14460 DVSS.n2380 DVSS.n2379 0.4505
R14461 DVSS.n2466 DVSS.n2465 0.4505
R14462 DVSS.n2467 DVSS.n2377 0.4505
R14463 DVSS.n2469 DVSS.n2468 0.4505
R14464 DVSS.n2474 DVSS.n2470 0.4505
R14465 DVSS.n2505 DVSS.n2504 0.4505
R14466 DVSS.n2471 DVSS.n2342 0.4505
R14467 DVSS.n2510 DVSS.n2509 0.4505
R14468 DVSS.n2341 DVSS.n2339 0.4505
R14469 DVSS.n2373 DVSS.n2372 0.4505
R14470 DVSS.n2345 DVSS.n2344 0.4505
R14471 DVSS.n2360 DVSS.n2359 0.4505
R14472 DVSS.n2354 DVSS.n2353 0.4505
R14473 DVSS.n2355 DVSS.n2350 0.4505
R14474 DVSS.n2319 DVSS.n2316 0.4505
R14475 DVSS.n2526 DVSS.n2525 0.4505
R14476 DVSS.n2317 DVSS.n2314 0.4505
R14477 DVSS.n2531 DVSS.n2530 0.4505
R14478 DVSS.n1913 DVSS.n1910 0.4505
R14479 DVSS.n2559 DVSS.n2558 0.4505
R14480 DVSS.n1907 DVSS.n1905 0.4505
R14481 DVSS.n2564 DVSS.n2563 0.4505
R14482 DVSS.n1906 DVSS.n1904 0.4505
R14483 DVSS.n2260 DVSS.n2259 0.4505
R14484 DVSS.n1886 DVSS.n1883 0.4505
R14485 DVSS.n2577 DVSS.n2576 0.4505
R14486 DVSS.n1884 DVSS.n1880 0.4505
R14487 DVSS.n2582 DVSS.n2581 0.4505
R14488 DVSS.n1879 DVSS.n1877 0.4505
R14489 DVSS.n2295 DVSS.n2294 0.4505
R14490 DVSS.n2272 DVSS.n2271 0.4505
R14491 DVSS.n1860 DVSS.n1858 0.4505
R14492 DVSS.n2281 DVSS.n2280 0.4505
R14493 DVSS.n2285 DVSS.n2284 0.4505
R14494 DVSS.n2275 DVSS.n2274 0.4505
R14495 DVSS.n2290 DVSS.n2289 0.4505
R14496 DVSS.n2614 DVSS.n2613 0.4505
R14497 DVSS.n2612 DVSS.n1850 0.4505
R14498 DVSS.n1854 DVSS.n1851 0.4505
R14499 DVSS.n2608 DVSS.n2607 0.4505
R14500 DVSS.n2606 DVSS.n1853 0.4505
R14501 DVSS.n2605 DVSS.n2604 0.4505
R14502 DVSS.n1937 DVSS.n1856 0.4505
R14503 DVSS.n2600 DVSS.n2599 0.4505
R14504 DVSS.n1635 DVSS.n1629 0.4505
R14505 DVSS.n4046 DVSS.n4045 0.4505
R14506 DVSS.n4044 DVSS.n1630 0.4505
R14507 DVSS.n4043 DVSS.n4042 0.4505
R14508 DVSS.n1637 DVSS.n1636 0.4505
R14509 DVSS.n4037 DVSS.n4036 0.4505
R14510 DVSS.n4035 DVSS.n1639 0.4505
R14511 DVSS.n4034 DVSS.n4033 0.4505
R14512 DVSS.n1641 DVSS.n1640 0.4505
R14513 DVSS.n4027 DVSS.n4026 0.4505
R14514 DVSS.n4025 DVSS.n1643 0.4505
R14515 DVSS.n4024 DVSS.n4023 0.4505
R14516 DVSS.n1645 DVSS.n1644 0.4505
R14517 DVSS.n4019 DVSS.n4018 0.4505
R14518 DVSS.n4017 DVSS.n1648 0.4505
R14519 DVSS.n4016 DVSS.n4015 0.4505
R14520 DVSS.n1650 DVSS.n1649 0.4505
R14521 DVSS.n4008 DVSS.n4007 0.4505
R14522 DVSS.n4006 DVSS.n1653 0.4505
R14523 DVSS.n4005 DVSS.n4004 0.4505
R14524 DVSS.n1655 DVSS.n1654 0.4505
R14525 DVSS.n4000 DVSS.n3999 0.4505
R14526 DVSS.n3998 DVSS.n1658 0.4505
R14527 DVSS.n3997 DVSS.n3996 0.4505
R14528 DVSS.n1660 DVSS.n1659 0.4505
R14529 DVSS.n3980 DVSS.n3979 0.4505
R14530 DVSS.n3978 DVSS.n1671 0.4505
R14531 DVSS.n3977 DVSS.n3976 0.4505
R14532 DVSS.n1673 DVSS.n1672 0.4505
R14533 DVSS.n3972 DVSS.n3971 0.4505
R14534 DVSS.n3970 DVSS.n1675 0.4505
R14535 DVSS.n3969 DVSS.n3968 0.4505
R14536 DVSS.n1677 DVSS.n1676 0.4505
R14537 DVSS.n3964 DVSS.n3963 0.4505
R14538 DVSS.n3962 DVSS.n1679 0.4505
R14539 DVSS.n3961 DVSS.n3960 0.4505
R14540 DVSS.n1681 DVSS.n1680 0.4505
R14541 DVSS.n1691 DVSS.n1689 0.4505
R14542 DVSS.n3951 DVSS.n3950 0.4505
R14543 DVSS.n3949 DVSS.n1690 0.4505
R14544 DVSS.n3948 DVSS.n3947 0.4505
R14545 DVSS.n1693 DVSS.n1692 0.4505
R14546 DVSS.n1712 DVSS.n1711 0.4505
R14547 DVSS.n1716 DVSS.n1715 0.4505
R14548 DVSS.n1717 DVSS.n1709 0.4505
R14549 DVSS.n3928 DVSS.n3927 0.4505
R14550 DVSS.n3926 DVSS.n1710 0.4505
R14551 DVSS.n3925 DVSS.n3924 0.4505
R14552 DVSS.n1719 DVSS.n1718 0.4505
R14553 DVSS.n3920 DVSS.n3919 0.4505
R14554 DVSS.n3918 DVSS.n1723 0.4505
R14555 DVSS.n3917 DVSS.n3916 0.4505
R14556 DVSS.n1725 DVSS.n1724 0.4505
R14557 DVSS.n3912 DVSS.n3911 0.4505
R14558 DVSS.n3910 DVSS.n1731 0.4505
R14559 DVSS.n3909 DVSS.n3908 0.4505
R14560 DVSS.n1733 DVSS.n1732 0.4505
R14561 DVSS.n3904 DVSS.n3903 0.4505
R14562 DVSS.n3902 DVSS.n1737 0.4505
R14563 DVSS.n3901 DVSS.n3900 0.4505
R14564 DVSS.n1739 DVSS.n1738 0.4505
R14565 DVSS.n3896 DVSS.n3895 0.4505
R14566 DVSS.n3894 DVSS.n1741 0.4505
R14567 DVSS.n3893 DVSS.n3892 0.4505
R14568 DVSS.n1743 DVSS.n1742 0.4505
R14569 DVSS.n3888 DVSS.n3887 0.4505
R14570 DVSS.n3886 DVSS.n1745 0.4505
R14571 DVSS.n3885 DVSS.n3884 0.4505
R14572 DVSS.n1747 DVSS.n1746 0.4505
R14573 DVSS.n3880 DVSS.n3879 0.4505
R14574 DVSS.n3878 DVSS.n1749 0.4505
R14575 DVSS.n3877 DVSS.n3876 0.4505
R14576 DVSS.n1751 DVSS.n1750 0.4505
R14577 DVSS.n3872 DVSS.n3871 0.4505
R14578 DVSS.n3870 DVSS.n1753 0.4505
R14579 DVSS.n3869 DVSS.n3868 0.4505
R14580 DVSS.n1755 DVSS.n1754 0.4505
R14581 DVSS.n1775 DVSS.n1774 0.4505
R14582 DVSS.n1773 DVSS.n1757 0.4505
R14583 DVSS.n1772 DVSS.n1771 0.4505
R14584 DVSS.n1759 DVSS.n1758 0.4505
R14585 DVSS.n1767 DVSS.n1766 0.4505
R14586 DVSS.n1765 DVSS.n1761 0.4505
R14587 DVSS.n1764 DVSS.n1763 0.4505
R14588 DVSS.n1761 DVSS.n1760 0.4505
R14589 DVSS.n1768 DVSS.n1767 0.4505
R14590 DVSS.n1769 DVSS.n1759 0.4505
R14591 DVSS.n1771 DVSS.n1770 0.4505
R14592 DVSS.n1757 DVSS.n1756 0.4505
R14593 DVSS.n1776 DVSS.n1775 0.4505
R14594 DVSS.n1777 DVSS.n1755 0.4505
R14595 DVSS.n3868 DVSS.n3867 0.4505
R14596 DVSS.n1753 DVSS.n1752 0.4505
R14597 DVSS.n3873 DVSS.n3872 0.4505
R14598 DVSS.n3874 DVSS.n1751 0.4505
R14599 DVSS.n3876 DVSS.n3875 0.4505
R14600 DVSS.n1749 DVSS.n1748 0.4505
R14601 DVSS.n3881 DVSS.n3880 0.4505
R14602 DVSS.n3882 DVSS.n1747 0.4505
R14603 DVSS.n3884 DVSS.n3883 0.4505
R14604 DVSS.n1745 DVSS.n1744 0.4505
R14605 DVSS.n3889 DVSS.n3888 0.4505
R14606 DVSS.n3890 DVSS.n1743 0.4505
R14607 DVSS.n3892 DVSS.n3891 0.4505
R14608 DVSS.n1741 DVSS.n1740 0.4505
R14609 DVSS.n3897 DVSS.n3896 0.4505
R14610 DVSS.n3898 DVSS.n1739 0.4505
R14611 DVSS.n3900 DVSS.n3899 0.4505
R14612 DVSS.n1737 DVSS.n1736 0.4505
R14613 DVSS.n3905 DVSS.n3904 0.4505
R14614 DVSS.n3906 DVSS.n1733 0.4505
R14615 DVSS.n3908 DVSS.n3907 0.4505
R14616 DVSS.n1734 DVSS.n1731 0.4505
R14617 DVSS.n3913 DVSS.n3912 0.4505
R14618 DVSS.n3914 DVSS.n1725 0.4505
R14619 DVSS.n3916 DVSS.n3915 0.4505
R14620 DVSS.n1723 DVSS.n1722 0.4505
R14621 DVSS.n3921 DVSS.n3920 0.4505
R14622 DVSS.n3922 DVSS.n1719 0.4505
R14623 DVSS.n3924 DVSS.n3923 0.4505
R14624 DVSS.n1720 DVSS.n1710 0.4505
R14625 DVSS.n3929 DVSS.n3928 0.4505
R14626 DVSS.n1709 DVSS.n1707 0.4505
R14627 DVSS.n1715 DVSS.n1714 0.4505
R14628 DVSS.n1713 DVSS.n1712 0.4505
R14629 DVSS.n1694 DVSS.n1693 0.4505
R14630 DVSS.n3947 DVSS.n3946 0.4505
R14631 DVSS.n1690 DVSS.n1688 0.4505
R14632 DVSS.n3952 DVSS.n3951 0.4505
R14633 DVSS.n1689 DVSS.n1687 0.4505
R14634 DVSS.n1682 DVSS.n1681 0.4505
R14635 DVSS.n3960 DVSS.n3959 0.4505
R14636 DVSS.n1679 DVSS.n1678 0.4505
R14637 DVSS.n3965 DVSS.n3964 0.4505
R14638 DVSS.n3966 DVSS.n1677 0.4505
R14639 DVSS.n3968 DVSS.n3967 0.4505
R14640 DVSS.n1675 DVSS.n1674 0.4505
R14641 DVSS.n3973 DVSS.n3972 0.4505
R14642 DVSS.n3974 DVSS.n1673 0.4505
R14643 DVSS.n3976 DVSS.n3975 0.4505
R14644 DVSS.n1671 DVSS.n1670 0.4505
R14645 DVSS.n3981 DVSS.n3980 0.4505
R14646 DVSS.n3982 DVSS.n1660 0.4505
R14647 DVSS.n3996 DVSS.n3995 0.4505
R14648 DVSS.n1661 DVSS.n1658 0.4505
R14649 DVSS.n4001 DVSS.n4000 0.4505
R14650 DVSS.n4002 DVSS.n1655 0.4505
R14651 DVSS.n4004 DVSS.n4003 0.4505
R14652 DVSS.n1656 DVSS.n1653 0.4505
R14653 DVSS.n4009 DVSS.n4008 0.4505
R14654 DVSS.n4013 DVSS.n1650 0.4505
R14655 DVSS.n4015 DVSS.n4014 0.4505
R14656 DVSS.n1651 DVSS.n1648 0.4505
R14657 DVSS.n4020 DVSS.n4019 0.4505
R14658 DVSS.n4021 DVSS.n1645 0.4505
R14659 DVSS.n4023 DVSS.n4022 0.4505
R14660 DVSS.n1646 DVSS.n1643 0.4505
R14661 DVSS.n4028 DVSS.n4027 0.4505
R14662 DVSS.n4030 DVSS.n1641 0.4505
R14663 DVSS.n4033 DVSS.n4032 0.4505
R14664 DVSS.n1639 DVSS.n1638 0.4505
R14665 DVSS.n4038 DVSS.n4037 0.4505
R14666 DVSS.n4039 DVSS.n1637 0.4505
R14667 DVSS.n4042 DVSS.n4041 0.4505
R14668 DVSS.n1630 DVSS.n1628 0.4505
R14669 DVSS.n4047 DVSS.n4046 0.4505
R14670 DVSS.n1629 DVSS.n1627 0.4505
R14671 DVSS.n1633 DVSS.n1632 0.4505
R14672 DVSS.n5090 DVSS.n5089 0.4505
R14673 DVSS.n1085 DVSS.n1084 0.4505
R14674 DVSS.n5085 DVSS.n5084 0.4505
R14675 DVSS.n5083 DVSS.n1087 0.4505
R14676 DVSS.n5082 DVSS.n5081 0.4505
R14677 DVSS.n1089 DVSS.n1088 0.4505
R14678 DVSS.n5077 DVSS.n5076 0.4505
R14679 DVSS.n5075 DVSS.n1091 0.4505
R14680 DVSS.n5074 DVSS.n5073 0.4505
R14681 DVSS.n1093 DVSS.n1092 0.4505
R14682 DVSS.n5069 DVSS.n5068 0.4505
R14683 DVSS.n5067 DVSS.n1095 0.4505
R14684 DVSS.n5066 DVSS.n5065 0.4505
R14685 DVSS.n1097 DVSS.n1096 0.4505
R14686 DVSS.n5060 DVSS.n5059 0.4505
R14687 DVSS.n5058 DVSS.n1100 0.4505
R14688 DVSS.n5057 DVSS.n5056 0.4505
R14689 DVSS.n1102 DVSS.n1101 0.4505
R14690 DVSS.n5052 DVSS.n5051 0.4505
R14691 DVSS.n5050 DVSS.n1105 0.4505
R14692 DVSS.n5049 DVSS.n5048 0.4505
R14693 DVSS.n1107 DVSS.n1106 0.4505
R14694 DVSS.n1113 DVSS.n1111 0.4505
R14695 DVSS.n5041 DVSS.n5040 0.4505
R14696 DVSS.n5039 DVSS.n1112 0.4505
R14697 DVSS.n5038 DVSS.n5037 0.4505
R14698 DVSS.n1115 DVSS.n1114 0.4505
R14699 DVSS.n5030 DVSS.n5029 0.4505
R14700 DVSS.n5028 DVSS.n1123 0.4505
R14701 DVSS.n5027 DVSS.n5026 0.4505
R14702 DVSS.n1125 DVSS.n1124 0.4505
R14703 DVSS.n5022 DVSS.n5021 0.4505
R14704 DVSS.n5020 DVSS.n1129 0.4505
R14705 DVSS.n5019 DVSS.n5018 0.4505
R14706 DVSS.n1131 DVSS.n1130 0.4505
R14707 DVSS.n5014 DVSS.n5013 0.4505
R14708 DVSS.n5012 DVSS.n1133 0.4505
R14709 DVSS.n5011 DVSS.n5010 0.4505
R14710 DVSS.n1135 DVSS.n1134 0.4505
R14711 DVSS.n5006 DVSS.n5005 0.4505
R14712 DVSS.n5004 DVSS.n1137 0.4505
R14713 DVSS.n5003 DVSS.n5002 0.4505
R14714 DVSS.n1139 DVSS.n1138 0.4505
R14715 DVSS.n4998 DVSS.n4997 0.4505
R14716 DVSS.n4996 DVSS.n1141 0.4505
R14717 DVSS.n4995 DVSS.n4994 0.4505
R14718 DVSS.n1143 DVSS.n1142 0.4505
R14719 DVSS.n4990 DVSS.n4989 0.4505
R14720 DVSS.n4988 DVSS.n1145 0.4505
R14721 DVSS.n4987 DVSS.n4986 0.4505
R14722 DVSS.n1147 DVSS.n1146 0.4505
R14723 DVSS.n4982 DVSS.n4981 0.4505
R14724 DVSS.n4980 DVSS.n1149 0.4505
R14725 DVSS.n4979 DVSS.n4978 0.4505
R14726 DVSS.n1151 DVSS.n1150 0.4505
R14727 DVSS.n4974 DVSS.n4973 0.4505
R14728 DVSS.n4972 DVSS.n1153 0.4505
R14729 DVSS.n4971 DVSS.n4970 0.4505
R14730 DVSS.n1155 DVSS.n1154 0.4505
R14731 DVSS.n4966 DVSS.n4965 0.4505
R14732 DVSS.n4964 DVSS.n1157 0.4505
R14733 DVSS.n4963 DVSS.n4962 0.4505
R14734 DVSS.n1159 DVSS.n1158 0.4505
R14735 DVSS.n4958 DVSS.n4957 0.4505
R14736 DVSS.n4956 DVSS.n1162 0.4505
R14737 DVSS.n4955 DVSS.n4954 0.4505
R14738 DVSS.n1164 DVSS.n1163 0.4505
R14739 DVSS.n4950 DVSS.n4949 0.4505
R14740 DVSS.n4948 DVSS.n1166 0.4505
R14741 DVSS.n4947 DVSS.n4946 0.4505
R14742 DVSS.n1168 DVSS.n1167 0.4505
R14743 DVSS.n4942 DVSS.n4941 0.4505
R14744 DVSS.n4940 DVSS.n1170 0.4505
R14745 DVSS.n4939 DVSS.n4938 0.4505
R14746 DVSS.n1172 DVSS.n1171 0.4505
R14747 DVSS.n4934 DVSS.n4933 0.4505
R14748 DVSS.n4932 DVSS.n1174 0.4505
R14749 DVSS.n4931 DVSS.n4930 0.4505
R14750 DVSS.n1176 DVSS.n1175 0.4505
R14751 DVSS.n4926 DVSS.n4925 0.4505
R14752 DVSS.n4924 DVSS.n1178 0.4505
R14753 DVSS.n4923 DVSS.n4922 0.4505
R14754 DVSS.n1180 DVSS.n1179 0.4505
R14755 DVSS.n4918 DVSS.n4917 0.4505
R14756 DVSS.n4916 DVSS.n1182 0.4505
R14757 DVSS.n4915 DVSS.n4914 0.4505
R14758 DVSS.n1184 DVSS.n1183 0.4505
R14759 DVSS.n4910 DVSS.n4909 0.4505
R14760 DVSS.n4908 DVSS.n1186 0.4505
R14761 DVSS.n4907 DVSS.n4906 0.4505
R14762 DVSS.n1188 DVSS.n1187 0.4505
R14763 DVSS.n4902 DVSS.n4901 0.4505
R14764 DVSS.n4900 DVSS.n1190 0.4505
R14765 DVSS.n4899 DVSS.n4898 0.4505
R14766 DVSS.n1192 DVSS.n1191 0.4505
R14767 DVSS.n4894 DVSS.n4893 0.4505
R14768 DVSS.n4892 DVSS.n1194 0.4505
R14769 DVSS.n4891 DVSS.n4890 0.4505
R14770 DVSS.n3516 DVSS.n1195 0.4505
R14771 DVSS.n3519 DVSS.n3518 0.4505
R14772 DVSS.n3515 DVSS.n3514 0.4505
R14773 DVSS.n3518 DVSS.n3517 0.4505
R14774 DVSS.n1199 DVSS.n1195 0.4505
R14775 DVSS.n4890 DVSS.n4889 0.4505
R14776 DVSS.n4878 DVSS.n1194 0.4505
R14777 DVSS.n4895 DVSS.n4894 0.4505
R14778 DVSS.n4896 DVSS.n1192 0.4505
R14779 DVSS.n4898 DVSS.n4897 0.4505
R14780 DVSS.n1190 DVSS.n1189 0.4505
R14781 DVSS.n4903 DVSS.n4902 0.4505
R14782 DVSS.n4904 DVSS.n1188 0.4505
R14783 DVSS.n4906 DVSS.n4905 0.4505
R14784 DVSS.n1186 DVSS.n1185 0.4505
R14785 DVSS.n4911 DVSS.n4910 0.4505
R14786 DVSS.n4912 DVSS.n1184 0.4505
R14787 DVSS.n4914 DVSS.n4913 0.4505
R14788 DVSS.n1182 DVSS.n1181 0.4505
R14789 DVSS.n4919 DVSS.n4918 0.4505
R14790 DVSS.n4920 DVSS.n1180 0.4505
R14791 DVSS.n4922 DVSS.n4921 0.4505
R14792 DVSS.n1178 DVSS.n1177 0.4505
R14793 DVSS.n4927 DVSS.n4926 0.4505
R14794 DVSS.n4928 DVSS.n1176 0.4505
R14795 DVSS.n4930 DVSS.n4929 0.4505
R14796 DVSS.n1174 DVSS.n1173 0.4505
R14797 DVSS.n4935 DVSS.n4934 0.4505
R14798 DVSS.n4936 DVSS.n1172 0.4505
R14799 DVSS.n4938 DVSS.n4937 0.4505
R14800 DVSS.n1170 DVSS.n1169 0.4505
R14801 DVSS.n4943 DVSS.n4942 0.4505
R14802 DVSS.n4944 DVSS.n1168 0.4505
R14803 DVSS.n4946 DVSS.n4945 0.4505
R14804 DVSS.n1166 DVSS.n1165 0.4505
R14805 DVSS.n4951 DVSS.n4950 0.4505
R14806 DVSS.n4952 DVSS.n1164 0.4505
R14807 DVSS.n4954 DVSS.n4953 0.4505
R14808 DVSS.n1162 DVSS.n1161 0.4505
R14809 DVSS.n4959 DVSS.n4958 0.4505
R14810 DVSS.n4960 DVSS.n1159 0.4505
R14811 DVSS.n4962 DVSS.n4961 0.4505
R14812 DVSS.n1160 DVSS.n1157 0.4505
R14813 DVSS.n4967 DVSS.n4966 0.4505
R14814 DVSS.n4968 DVSS.n1155 0.4505
R14815 DVSS.n4970 DVSS.n4969 0.4505
R14816 DVSS.n1153 DVSS.n1152 0.4505
R14817 DVSS.n4975 DVSS.n4974 0.4505
R14818 DVSS.n4976 DVSS.n1151 0.4505
R14819 DVSS.n4978 DVSS.n4977 0.4505
R14820 DVSS.n1149 DVSS.n1148 0.4505
R14821 DVSS.n4983 DVSS.n4982 0.4505
R14822 DVSS.n4984 DVSS.n1147 0.4505
R14823 DVSS.n4986 DVSS.n4985 0.4505
R14824 DVSS.n1145 DVSS.n1144 0.4505
R14825 DVSS.n4991 DVSS.n4990 0.4505
R14826 DVSS.n4992 DVSS.n1143 0.4505
R14827 DVSS.n4994 DVSS.n4993 0.4505
R14828 DVSS.n1141 DVSS.n1140 0.4505
R14829 DVSS.n4999 DVSS.n4998 0.4505
R14830 DVSS.n5000 DVSS.n1139 0.4505
R14831 DVSS.n5002 DVSS.n5001 0.4505
R14832 DVSS.n1137 DVSS.n1136 0.4505
R14833 DVSS.n5007 DVSS.n5006 0.4505
R14834 DVSS.n5008 DVSS.n1135 0.4505
R14835 DVSS.n5010 DVSS.n5009 0.4505
R14836 DVSS.n1133 DVSS.n1132 0.4505
R14837 DVSS.n5015 DVSS.n5014 0.4505
R14838 DVSS.n5016 DVSS.n1131 0.4505
R14839 DVSS.n5018 DVSS.n5017 0.4505
R14840 DVSS.n1129 DVSS.n1128 0.4505
R14841 DVSS.n5023 DVSS.n5022 0.4505
R14842 DVSS.n5024 DVSS.n1125 0.4505
R14843 DVSS.n5026 DVSS.n5025 0.4505
R14844 DVSS.n1126 DVSS.n1123 0.4505
R14845 DVSS.n5031 DVSS.n5030 0.4505
R14846 DVSS.n1118 DVSS.n1115 0.4505
R14847 DVSS.n5037 DVSS.n5036 0.4505
R14848 DVSS.n1116 DVSS.n1112 0.4505
R14849 DVSS.n5042 DVSS.n5041 0.4505
R14850 DVSS.n1111 DVSS.n1108 0.4505
R14851 DVSS.n5046 DVSS.n1107 0.4505
R14852 DVSS.n5048 DVSS.n5047 0.4505
R14853 DVSS.n1105 DVSS.n1104 0.4505
R14854 DVSS.n5053 DVSS.n5052 0.4505
R14855 DVSS.n5054 DVSS.n1102 0.4505
R14856 DVSS.n5056 DVSS.n5055 0.4505
R14857 DVSS.n1103 DVSS.n1100 0.4505
R14858 DVSS.n5061 DVSS.n5060 0.4505
R14859 DVSS.n5063 DVSS.n1097 0.4505
R14860 DVSS.n5065 DVSS.n5064 0.4505
R14861 DVSS.n1095 DVSS.n1094 0.4505
R14862 DVSS.n5070 DVSS.n5069 0.4505
R14863 DVSS.n5071 DVSS.n1093 0.4505
R14864 DVSS.n5073 DVSS.n5072 0.4505
R14865 DVSS.n1091 DVSS.n1090 0.4505
R14866 DVSS.n5078 DVSS.n5077 0.4505
R14867 DVSS.n5079 DVSS.n1089 0.4505
R14868 DVSS.n5081 DVSS.n5080 0.4505
R14869 DVSS.n1087 DVSS.n1086 0.4505
R14870 DVSS.n5086 DVSS.n5085 0.4505
R14871 DVSS.n5087 DVSS.n1085 0.4505
R14872 DVSS.n5089 DVSS.n5088 0.4505
R14873 DVSS.n1083 DVSS.n1082 0.4505
R14874 DVSS.n3607 DVSS.n3606 0.4505
R14875 DVSS.n3611 DVSS.n3610 0.4505
R14876 DVSS.n3612 DVSS.n3605 0.4505
R14877 DVSS.n3614 DVSS.n3613 0.4505
R14878 DVSS.n3603 DVSS.n3602 0.4505
R14879 DVSS.n3619 DVSS.n3618 0.4505
R14880 DVSS.n3620 DVSS.n3601 0.4505
R14881 DVSS.n3622 DVSS.n3621 0.4505
R14882 DVSS.n3599 DVSS.n3598 0.4505
R14883 DVSS.n3627 DVSS.n3626 0.4505
R14884 DVSS.n3628 DVSS.n3597 0.4505
R14885 DVSS.n3630 DVSS.n3629 0.4505
R14886 DVSS.n3595 DVSS.n3594 0.4505
R14887 DVSS.n3635 DVSS.n3634 0.4505
R14888 DVSS.n3636 DVSS.n3593 0.4505
R14889 DVSS.n3638 DVSS.n3637 0.4505
R14890 DVSS.n3591 DVSS.n3590 0.4505
R14891 DVSS.n3643 DVSS.n3642 0.4505
R14892 DVSS.n3644 DVSS.n3589 0.4505
R14893 DVSS.n3646 DVSS.n3645 0.4505
R14894 DVSS.n3587 DVSS.n3586 0.4505
R14895 DVSS.n3651 DVSS.n3650 0.4505
R14896 DVSS.n3652 DVSS.n3585 0.4505
R14897 DVSS.n3654 DVSS.n3653 0.4505
R14898 DVSS.n3583 DVSS.n3582 0.4505
R14899 DVSS.n3659 DVSS.n3658 0.4505
R14900 DVSS.n3660 DVSS.n3581 0.4505
R14901 DVSS.n3662 DVSS.n3661 0.4505
R14902 DVSS.n3579 DVSS.n3578 0.4505
R14903 DVSS.n3667 DVSS.n3666 0.4505
R14904 DVSS.n3668 DVSS.n3577 0.4505
R14905 DVSS.n3670 DVSS.n3669 0.4505
R14906 DVSS.n3575 DVSS.n3574 0.4505
R14907 DVSS.n3675 DVSS.n3674 0.4505
R14908 DVSS.n3676 DVSS.n3573 0.4505
R14909 DVSS.n3678 DVSS.n3677 0.4505
R14910 DVSS.n3571 DVSS.n3570 0.4505
R14911 DVSS.n3683 DVSS.n3682 0.4505
R14912 DVSS.n3684 DVSS.n3569 0.4505
R14913 DVSS.n3686 DVSS.n3685 0.4505
R14914 DVSS.n3567 DVSS.n3566 0.4505
R14915 DVSS.n3691 DVSS.n3690 0.4505
R14916 DVSS.n3692 DVSS.n3565 0.4505
R14917 DVSS.n3694 DVSS.n3693 0.4505
R14918 DVSS.n3563 DVSS.n3562 0.4505
R14919 DVSS.n3699 DVSS.n3698 0.4505
R14920 DVSS.n3700 DVSS.n3561 0.4505
R14921 DVSS.n3702 DVSS.n3701 0.4505
R14922 DVSS.n3559 DVSS.n3558 0.4505
R14923 DVSS.n3707 DVSS.n3706 0.4505
R14924 DVSS.n3708 DVSS.n3557 0.4505
R14925 DVSS.n3710 DVSS.n3709 0.4505
R14926 DVSS.n3555 DVSS.n3554 0.4505
R14927 DVSS.n3715 DVSS.n3714 0.4505
R14928 DVSS.n3716 DVSS.n3553 0.4505
R14929 DVSS.n3718 DVSS.n3717 0.4505
R14930 DVSS.n3551 DVSS.n3550 0.4505
R14931 DVSS.n3723 DVSS.n3722 0.4505
R14932 DVSS.n3724 DVSS.n3549 0.4505
R14933 DVSS.n3726 DVSS.n3725 0.4505
R14934 DVSS.n3547 DVSS.n3546 0.4505
R14935 DVSS.n3731 DVSS.n3730 0.4505
R14936 DVSS.n3732 DVSS.n3545 0.4505
R14937 DVSS.n3734 DVSS.n3733 0.4505
R14938 DVSS.n3543 DVSS.n3542 0.4505
R14939 DVSS.n3739 DVSS.n3738 0.4505
R14940 DVSS.n3740 DVSS.n3541 0.4505
R14941 DVSS.n3742 DVSS.n3741 0.4505
R14942 DVSS.n3539 DVSS.n3534 0.4505
R14943 DVSS.n3749 DVSS.n3748 0.4505
R14944 DVSS.n3745 DVSS.n3527 0.4505
R14945 DVSS.n3762 DVSS.n3526 0.4505
R14946 DVSS.n3764 DVSS.n3763 0.4505
R14947 DVSS.n3524 DVSS.n3523 0.4505
R14948 DVSS.n1574 DVSS.n1573 0.4505
R14949 DVSS.n1575 DVSS.n1570 0.4505
R14950 DVSS.n1577 DVSS.n1576 0.4505
R14951 DVSS.n1568 DVSS.n1567 0.4505
R14952 DVSS.n1582 DVSS.n1581 0.4505
R14953 DVSS.n1583 DVSS.n1566 0.4505
R14954 DVSS.n1585 DVSS.n1584 0.4505
R14955 DVSS.n1564 DVSS.n1563 0.4505
R14956 DVSS.n1590 DVSS.n1589 0.4505
R14957 DVSS.n1591 DVSS.n1562 0.4505
R14958 DVSS.n1593 DVSS.n1592 0.4505
R14959 DVSS.n1559 DVSS.n1557 0.4505
R14960 DVSS.n4090 DVSS.n4089 0.4505
R14961 DVSS.n1560 DVSS.n1558 0.4505
R14962 DVSS.n4085 DVSS.n4084 0.4505
R14963 DVSS.n4083 DVSS.n1597 0.4505
R14964 DVSS.n4082 DVSS.n4081 0.4505
R14965 DVSS.n1599 DVSS.n1598 0.4505
R14966 DVSS.n4077 DVSS.n4076 0.4505
R14967 DVSS.n4075 DVSS.n1601 0.4505
R14968 DVSS.n4074 DVSS.n4073 0.4505
R14969 DVSS.n1603 DVSS.n1602 0.4505
R14970 DVSS.n4069 DVSS.n4068 0.4505
R14971 DVSS.n4067 DVSS.n1605 0.4505
R14972 DVSS.n4066 DVSS.n4065 0.4505
R14973 DVSS.n1607 DVSS.n1606 0.4505
R14974 DVSS.n4061 DVSS.n4060 0.4505
R14975 DVSS.n1610 DVSS.n1609 0.4505
R14976 DVSS.n4284 DVSS 0.449176
R14977 DVSS.n4855 DVSS 0.449176
R14978 DVSS.n4855 DVSS 0.449176
R14979 DVSS.n2649 VSS 0.444617
R14980 DVSS.n2662 VSS 0.444617
R14981 DVSS.n2646 VSS 0.444542
R14982 DVSS.n2661 VSS 0.444542
R14983 DVSS.n1839 DVSS.n1838 0.441235
R14984 DVSS.n1370 DVSS.n957 0.439524
R14985 DVSS.n5342 DVSS.n5341 0.439458
R14986 DVSS.n3507 DVSS.n2665 0.429011
R14987 DVSS.n3507 DVSS.n3506 0.429011
R14988 DVSS.n4789 DVSS.n1249 0.41962
R14989 DVSS.n4179 DVSS.n1468 0.41962
R14990 DVSS.n4105 DVSS.n4104 0.4165
R14991 DVSS.n4111 DVSS.n4110 0.4165
R14992 DVSS.n2647 VSS 0.415539
R14993 DVSS.n2648 VSS 0.415539
R14994 DVSS.n4102 DVSS.n1548 0.412794
R14995 DVSS.n2626 DVSS.t20 0.41
R14996 DVSS.n2626 DVSS.t22 0.41
R14997 DVSS.n2015 DVSS.n1976 0.407769
R14998 DVSS.n3935 DVSS 0.402853
R14999 DVSS DVSS.n1684 0.402853
R15000 DVSS.n4055 DVSS 0.402853
R15001 DVSS DVSS.n4051 0.402853
R15002 DVSS.n2541 DVSS.n2539 0.388068
R15003 DVSS.n2302 DVSS.n1928 0.387662
R15004 DVSS.n4284 DVSS 0.384324
R15005 DVSS.n2015 DVSS.n2014 0.38247
R15006 DVSS.n2646 DVSS.n1556 0.375755
R15007 DVSS.n2543 DVSS.n2542 0.3755
R15008 DVSS.n2304 DVSS.n2303 0.3755
R15009 DVSS.n1516 DVSS.n1120 0.3755
R15010 DVSS.n3956 DVSS.n3955 0.368789
R15011 DVSS.n1728 DVSS.n1697 0.368789
R15012 DVSS.n3935 DVSS.n1700 0.368789
R15013 DVSS.n3934 DVSS.n1702 0.368789
R15014 DVSS.n3932 DVSS.n3931 0.368789
R15015 DVSS.n3943 DVSS.n1684 0.368789
R15016 DVSS.n4011 DVSS.n1611 0.368789
R15017 DVSS.n4055 DVSS.n1614 0.368789
R15018 DVSS.n4054 DVSS.n1616 0.368789
R15019 DVSS.n4052 DVSS.n1619 0.368789
R15020 DVSS.n4051 DVSS.n1622 0.368789
R15021 DVSS.n4050 DVSS.n4049 0.368789
R15022 DVSS.n1816 DVSS.n1796 0.367935
R15023 DVSS.n1817 DVSS.n1796 0.367935
R15024 DVSS.n1811 DVSS.n1797 0.367935
R15025 DVSS.n1818 DVSS.n1797 0.367935
R15026 DVSS.n1809 DVSS.n1798 0.367935
R15027 DVSS.n1819 DVSS.n1798 0.367935
R15028 DVSS.n1807 DVSS.n1799 0.367935
R15029 DVSS.n1820 DVSS.n1799 0.367935
R15030 DVSS.n1805 DVSS.n1800 0.367935
R15031 DVSS.n1821 DVSS.n1800 0.367935
R15032 DVSS.n1803 DVSS.n1801 0.367935
R15033 DVSS.n3818 DVSS.n3817 0.367935
R15034 DVSS.n1821 DVSS.n1804 0.367935
R15035 DVSS.n1820 DVSS.n1806 0.367935
R15036 DVSS.n1819 DVSS.n1808 0.367935
R15037 DVSS.n1818 DVSS.n1810 0.367935
R15038 DVSS.n1817 DVSS.n1812 0.367935
R15039 DVSS.n1804 DVSS.n1803 0.367935
R15040 DVSS.n1806 DVSS.n1805 0.367935
R15041 DVSS.n1808 DVSS.n1807 0.367935
R15042 DVSS.n1810 DVSS.n1809 0.367935
R15043 DVSS.n1812 DVSS.n1811 0.367935
R15044 DVSS.n3820 DVSS.n1816 0.367935
R15045 DVSS.n3818 DVSS.n1801 0.367935
R15046 DVSS.n1457 DVSS 0.366421
R15047 DVSS.n4815 DVSS 0.366421
R15048 DVSS.n1479 DVSS 0.366421
R15049 DVSS.n1272 DVSS 0.366421
R15050 DVSS.n4159 DVSS 0.358788
R15051 DVSS.n2016 DVSS.n1969 0.346654
R15052 DVSS.n2017 DVSS.n2016 0.346654
R15053 DVSS.n1459 DVSS 0.346309
R15054 DVSS.n1461 DVSS 0.346309
R15055 DVSS.n1228 DVSS 0.346309
R15056 DVSS.n4817 DVSS 0.346309
R15057 DVSS.n1481 DVSS 0.346309
R15058 DVSS.n1499 DVSS 0.346309
R15059 DVSS.n1270 DVSS 0.346309
R15060 DVSS.n1274 DVSS 0.346309
R15061 DVSS.n1454 DVSS 0.346114
R15062 DVSS.n4820 DVSS 0.346114
R15063 DVSS.n1225 DVSS 0.346114
R15064 DVSS.n1311 DVSS.n1210 0.342906
R15065 DVSS.n2651 DVSS.n2650 0.335984
R15066 DVSS.n4731 DVSS.n4608 0.328381
R15067 DVSS.n4718 DVSS.n4717 0.328381
R15068 DVSS.n4587 DVSS.n4586 0.328381
R15069 DVSS.n4601 DVSS.n1396 0.328381
R15070 DVSS.n4549 DVSS.n1428 0.328381
R15071 DVSS.n4567 DVSS.n4566 0.328381
R15072 DVSS.n4451 DVSS.n1448 0.328381
R15073 DVSS.n4527 DVSS.n4526 0.328381
R15074 DVSS.n4483 DVSS.n4415 0.328381
R15075 DVSS.n4470 DVSS.n4469 0.328381
R15076 DVSS.n4394 DVSS.n4393 0.328381
R15077 DVSS.n4408 DVSS.n4325 0.328381
R15078 DVSS.n2308 DVSS.n2307 0.311888
R15079 DVSS.n2547 DVSS.n2546 0.311888
R15080 DVSS DVSS.n1848 0.309579
R15081 DVSS.n2650 DVSS.n2646 0.307559
R15082 DVSS.n4312 DVSS.n4311 0.297643
R15083 DVSS.n1501 DVSS.n1477 0.297643
R15084 DVSS.n4809 DVSS.n4808 0.297643
R15085 DVSS.n4783 DVSS.n4782 0.297643
R15086 DVSS.n804 DVSS.n803 0.28175
R15087 DVSS.n365 DVSS.n229 0.28175
R15088 DVSS.n1842 DVSS 0.273784
R15089 DVSS.n1465 DVSS.t6 0.2735
R15090 DVSS.n1465 DVSS.t1 0.2735
R15091 DVSS.n1470 DVSS.t107 0.2735
R15092 DVSS.n1470 DVSS.t24 0.2735
R15093 DVSS.n1974 DVSS.t12 0.2735
R15094 DVSS.n1453 DVSS.t201 0.2735
R15095 DVSS.n1458 DVSS.t123 0.2735
R15096 DVSS.n1458 DVSS.t125 0.2735
R15097 DVSS.n1460 DVSS.t203 0.2735
R15098 DVSS.n1460 DVSS.t161 0.2735
R15099 DVSS.n1252 DVSS.t129 0.2735
R15100 DVSS.n1252 DVSS.t18 0.2735
R15101 DVSS.n1231 DVSS.t9 0.2735
R15102 DVSS.n1231 DVSS.t168 0.2735
R15103 DVSS.n4805 DVSS.t180 0.2735
R15104 DVSS.n1227 DVSS.t71 0.2735
R15105 DVSS.n1227 DVSS.t37 0.2735
R15106 DVSS.n4816 DVSS.t65 0.2735
R15107 DVSS.n4816 DVSS.t67 0.2735
R15108 DVSS.n4819 DVSS.t69 0.2735
R15109 DVSS.n1224 DVSS.t163 0.2735
R15110 DVSS.n1480 DVSS.t41 0.2735
R15111 DVSS.n1480 DVSS.t75 0.2735
R15112 DVSS.n1498 DVSS.t47 0.2735
R15113 DVSS.n1498 DVSS.t39 0.2735
R15114 DVSS.n4183 DVSS.t113 0.2735
R15115 DVSS.n1266 DVSS.t127 0.2735
R15116 DVSS.n1269 DVSS.t157 0.2735
R15117 DVSS.n1269 DVSS.t153 0.2735
R15118 DVSS.n1273 DVSS.t155 0.2735
R15119 DVSS.n1273 DVSS.t121 0.2735
R15120 DVSS.n1345 DVSS.t98 0.2735
R15121 DVSS.n4117 DVSS.n4116 0.273147
R15122 DVSS.n4113 DVSS.n1550 0.273147
R15123 DVSS.n4294 DVSS.n1468 0.271321
R15124 DVSS.n4789 DVSS.n4788 0.271321
R15125 DVSS.n3796 DVSS.n3795 0.268132
R15126 DVSS.n4778 DVSS.n1275 0.266421
R15127 DVSS.n4822 DVSS.n1226 0.265206
R15128 DVSS.n4822 DVSS.n4821 0.265206
R15129 DVSS.n105 DVSS.n61 0.265206
R15130 DVSS.n260 DVSS.n252 0.265206
R15131 DVSS.n1988 DVSS.n1468 0.264797
R15132 DVSS.n4790 DVSS.n4789 0.264797
R15133 DVSS.n4318 DVSS.n4317 0.2605
R15134 DVSS.n4824 DVSS.n4823 0.2605
R15135 DVSS.n4759 DVSS.n1275 0.2605
R15136 DVSS.n1514 VSS 0.258658
R15137 DVSS.n4165 DVSS.n1522 0.254359
R15138 DVSS.n4837 DVSS.n4836 0.249324
R15139 DVSS.n4843 DVSS.n4842 0.249324
R15140 DVSS.n4864 DVSS.n4863 0.249324
R15141 DVSS.n4806 DVSS.n4803 0.243385
R15142 DVSS.n4185 DVSS.n4182 0.243385
R15143 DVSS.n1976 DVSS.n1973 0.243385
R15144 DVSS.n1267 DVSS.n1264 0.243385
R15145 DVSS.n1347 DVSS.n1344 0.243385
R15146 DVSS.n3795 DVSS.n3794 0.242079
R15147 DVSS.n2650 DVSS.n2649 0.238735
R15148 DVSS.n5793 DVSS.n5792 0.232304
R15149 DVSS.n2305 DVSS.n2304 0.231484
R15150 DVSS.n2544 DVSS.n2543 0.231484
R15151 DVSS.n4685 DVSS.n4679 0.231338
R15152 DVSS.n1572 DVSS.n1569 0.231338
R15153 DVSS.n3766 DVSS.n3765 0.231338
R15154 DVSS.n5091 DVSS.n5090 0.231338
R15155 DVSS.n3520 DVSS.n3519 0.231338
R15156 DVSS.n5546 DVSS.n5545 0.229958
R15157 DVSS.n5798 DVSS.n5797 0.229958
R15158 DVSS.n2304 DVSS.n2267 0.229569
R15159 VSS DVSS.n4841 0.229471
R15160 DVSS.n4841 VSS 0.229471
R15161 DVSS.n2543 DVSS.n1926 0.228851
R15162 DVSS.n1515 DVSS.n1514 0.224316
R15163 DVSS.n1830 DVSS 0.223543
R15164 DVSS.n4773 DVSS.n4772 0.219756
R15165 DVSS.n55 DVSS.n48 0.214786
R15166 DVSS.n426 DVSS.n425 0.214786
R15167 DVSS.n4775 DVSS.n1353 0.214786
R15168 DVSS.n1352 DVSS.n1278 0.214786
R15169 DVSS.n1351 DVSS.n1350 0.214786
R15170 DVSS.n1342 DVSS.n1341 0.214786
R15171 DVSS.n1340 DVSS.n1280 0.214786
R15172 DVSS.n1339 DVSS.n1338 0.214786
R15173 DVSS.n1282 DVSS.n1281 0.214786
R15174 DVSS.n1334 DVSS.n1333 0.214786
R15175 DVSS.n1332 DVSS.n1284 0.214786
R15176 DVSS.n1331 DVSS.n1330 0.214786
R15177 DVSS.n1286 DVSS.n1285 0.214786
R15178 DVSS.n1326 DVSS.n1325 0.214786
R15179 DVSS.n1324 DVSS.n1288 0.214786
R15180 DVSS.n1323 DVSS.n1322 0.214786
R15181 DVSS.n1290 DVSS.n1289 0.214786
R15182 DVSS.n1318 DVSS.n1317 0.214786
R15183 DVSS.n1316 DVSS.n1292 0.214786
R15184 DVSS.n1315 DVSS.n1314 0.214786
R15185 DVSS.n1294 DVSS.n1293 0.214786
R15186 DVSS.n1309 DVSS.n1308 0.214786
R15187 DVSS.n1307 DVSS.n1296 0.214786
R15188 DVSS.n1306 DVSS.n1305 0.214786
R15189 DVSS.n1298 DVSS.n1297 0.214786
R15190 DVSS.n1301 DVSS.n1300 0.214786
R15191 DVSS.n1299 DVSS.n1247 0.214786
R15192 DVSS.n4792 DVSS.n1246 0.214786
R15193 DVSS.n4793 DVSS.n1245 0.214786
R15194 DVSS.n4794 DVSS.n1244 0.214786
R15195 DVSS.n1243 DVSS.n1241 0.214786
R15196 DVSS.n4798 DVSS.n1240 0.214786
R15197 DVSS.n4799 DVSS.n1239 0.214786
R15198 DVSS.n2011 DVSS.n1979 0.214786
R15199 DVSS.n2010 DVSS.n1980 0.214786
R15200 DVSS.n1983 DVSS.n1981 0.214786
R15201 DVSS.n2006 DVSS.n1984 0.214786
R15202 DVSS.n2005 DVSS.n1985 0.214786
R15203 DVSS.n2004 DVSS.n1986 0.214786
R15204 DVSS.n1990 DVSS.n1987 0.214786
R15205 DVSS.n2000 DVSS.n1991 0.214786
R15206 DVSS.n1999 DVSS.n1992 0.214786
R15207 DVSS.n1998 DVSS.n1993 0.214786
R15208 DVSS.n1995 DVSS.n1994 0.214786
R15209 DVSS.n1496 DVSS.n1495 0.214786
R15210 DVSS.n4189 DVSS.n4188 0.214786
R15211 DVSS.n4190 DVSS.n1494 0.214786
R15212 DVSS.n4192 DVSS.n4191 0.214786
R15213 DVSS.n1492 DVSS.n1491 0.214786
R15214 DVSS.n4197 DVSS.n4196 0.214786
R15215 DVSS.n4198 DVSS.n1490 0.214786
R15216 DVSS.n4200 DVSS.n4199 0.214786
R15217 DVSS.n1488 DVSS.n1487 0.214786
R15218 DVSS.n4205 DVSS.n4204 0.214786
R15219 DVSS.n4206 DVSS.n1486 0.214786
R15220 DVSS.n4280 DVSS.n4207 0.214786
R15221 DVSS.n4279 DVSS.n4208 0.214786
R15222 DVSS.n4278 DVSS.n4209 0.214786
R15223 DVSS.n4212 DVSS.n4210 0.214786
R15224 DVSS.n4274 DVSS.n4213 0.214786
R15225 DVSS.n4273 DVSS.n4214 0.214786
R15226 DVSS.n4272 DVSS.n4215 0.214786
R15227 DVSS.n4218 DVSS.n4216 0.214786
R15228 DVSS.n4268 DVSS.n4219 0.214786
R15229 DVSS.n4267 DVSS.n4220 0.214786
R15230 DVSS.n4266 DVSS.n4221 0.214786
R15231 DVSS.n4224 DVSS.n4222 0.214786
R15232 DVSS.n4262 DVSS.n4225 0.214786
R15233 DVSS.n4261 DVSS.n4226 0.214786
R15234 DVSS.n4260 DVSS.n4227 0.214786
R15235 DVSS.n4230 DVSS.n4228 0.214786
R15236 DVSS.n4256 DVSS.n4231 0.214786
R15237 DVSS.n4255 DVSS.n4232 0.214786
R15238 DVSS.n4254 DVSS.n4233 0.214786
R15239 DVSS.n4236 DVSS.n4234 0.214786
R15240 DVSS.n4250 DVSS.n4237 0.214786
R15241 DVSS.n4249 DVSS.n4238 0.214786
R15242 DVSS.n4248 DVSS.n4239 0.214786
R15243 DVSS.n4241 DVSS.n4240 0.214786
R15244 DVSS.n4244 DVSS.n4243 0.214786
R15245 DVSS.n4242 DVSS.n1237 0.214786
R15246 DVSS.n4800 DVSS.n1238 0.214786
R15247 DVSS.n1248 DVSS.n1247 0.214786
R15248 DVSS.n4774 DVSS.n1277 0.214786
R15249 DVSS.n4776 DVSS.n4775 0.214786
R15250 DVSS.n1278 DVSS.n1276 0.214786
R15251 DVSS.n1350 DVSS.n1349 0.214786
R15252 DVSS.n1343 DVSS.n1342 0.214786
R15253 DVSS.n1280 DVSS.n1279 0.214786
R15254 DVSS.n1338 DVSS.n1337 0.214786
R15255 DVSS.n1336 DVSS.n1282 0.214786
R15256 DVSS.n1335 DVSS.n1334 0.214786
R15257 DVSS.n1284 DVSS.n1283 0.214786
R15258 DVSS.n1330 DVSS.n1329 0.214786
R15259 DVSS.n1328 DVSS.n1286 0.214786
R15260 DVSS.n1327 DVSS.n1326 0.214786
R15261 DVSS.n1288 DVSS.n1287 0.214786
R15262 DVSS.n1322 DVSS.n1321 0.214786
R15263 DVSS.n1320 DVSS.n1290 0.214786
R15264 DVSS.n1319 DVSS.n1318 0.214786
R15265 DVSS.n1292 DVSS.n1291 0.214786
R15266 DVSS.n1314 DVSS.n1313 0.214786
R15267 DVSS.n1312 DVSS.n1294 0.214786
R15268 DVSS.n4799 DVSS.n1236 0.214786
R15269 DVSS.n4798 DVSS.n4797 0.214786
R15270 DVSS.n4796 DVSS.n1241 0.214786
R15271 DVSS.n4795 DVSS.n4794 0.214786
R15272 DVSS.n4793 DVSS.n1242 0.214786
R15273 DVSS.n4792 DVSS.n4791 0.214786
R15274 DVSS.n1302 DVSS.n1301 0.214786
R15275 DVSS.n1303 DVSS.n1298 0.214786
R15276 DVSS.n1305 DVSS.n1304 0.214786
R15277 DVSS.n1296 DVSS.n1295 0.214786
R15278 DVSS.n1310 DVSS.n1309 0.214786
R15279 DVSS.n2013 DVSS.n2012 0.214786
R15280 DVSS.n2011 DVSS.n1978 0.214786
R15281 DVSS.n2010 DVSS.n2009 0.214786
R15282 DVSS.n2008 DVSS.n1981 0.214786
R15283 DVSS.n2007 DVSS.n2006 0.214786
R15284 DVSS.n2005 DVSS.n1982 0.214786
R15285 DVSS.n2004 DVSS.n2003 0.214786
R15286 DVSS.n2002 DVSS.n1987 0.214786
R15287 DVSS.n2001 DVSS.n2000 0.214786
R15288 DVSS.n1999 DVSS.n1989 0.214786
R15289 DVSS.n1998 DVSS.n1997 0.214786
R15290 DVSS.n1996 DVSS.n1995 0.214786
R15291 DVSS.n1497 DVSS.n1496 0.214786
R15292 DVSS.n4188 DVSS.n4187 0.214786
R15293 DVSS.n1494 DVSS.n1493 0.214786
R15294 DVSS.n4193 DVSS.n4192 0.214786
R15295 DVSS.n4194 DVSS.n1492 0.214786
R15296 DVSS.n4196 DVSS.n4195 0.214786
R15297 DVSS.n1490 DVSS.n1489 0.214786
R15298 DVSS.n4201 DVSS.n4200 0.214786
R15299 DVSS.n4202 DVSS.n1488 0.214786
R15300 DVSS.n4204 DVSS.n4203 0.214786
R15301 DVSS.n1486 DVSS.n1484 0.214786
R15302 DVSS.n4281 DVSS.n4280 0.214786
R15303 DVSS.n4279 DVSS.n1485 0.214786
R15304 DVSS.n4278 DVSS.n4277 0.214786
R15305 DVSS.n4276 DVSS.n4210 0.214786
R15306 DVSS.n4275 DVSS.n4274 0.214786
R15307 DVSS.n4273 DVSS.n4211 0.214786
R15308 DVSS.n4272 DVSS.n4271 0.214786
R15309 DVSS.n4270 DVSS.n4216 0.214786
R15310 DVSS.n4269 DVSS.n4268 0.214786
R15311 DVSS.n4267 DVSS.n4217 0.214786
R15312 DVSS.n4266 DVSS.n4265 0.214786
R15313 DVSS.n4264 DVSS.n4222 0.214786
R15314 DVSS.n4263 DVSS.n4262 0.214786
R15315 DVSS.n4261 DVSS.n4223 0.214786
R15316 DVSS.n4260 DVSS.n4259 0.214786
R15317 DVSS.n4258 DVSS.n4228 0.214786
R15318 DVSS.n4257 DVSS.n4256 0.214786
R15319 DVSS.n4255 DVSS.n4229 0.214786
R15320 DVSS.n4254 DVSS.n4253 0.214786
R15321 DVSS.n4252 DVSS.n4234 0.214786
R15322 DVSS.n4251 DVSS.n4250 0.214786
R15323 DVSS.n4249 DVSS.n4235 0.214786
R15324 DVSS.n4248 DVSS.n4247 0.214786
R15325 DVSS.n4246 DVSS.n4240 0.214786
R15326 DVSS.n4245 DVSS.n4244 0.214786
R15327 DVSS.n1237 DVSS.n1235 0.214786
R15328 DVSS.n4801 DVSS.n4800 0.214786
R15329 DVSS.n497 DVSS.n209 0.214786
R15330 DVSS.n828 DVSS.n826 0.214786
R15331 DVSS.n827 DVSS.n825 0.214786
R15332 DVSS.n5549 DVSS.n824 0.214786
R15333 DVSS.n5550 DVSS.n823 0.214786
R15334 DVSS.n5551 DVSS.n822 0.214786
R15335 DVSS.n821 DVSS.n819 0.214786
R15336 DVSS.n5555 DVSS.n818 0.214786
R15337 DVSS.n5556 DVSS.n817 0.214786
R15338 DVSS.n5557 DVSS.n816 0.214786
R15339 DVSS.n815 DVSS.n813 0.214786
R15340 DVSS.n5561 DVSS.n812 0.214786
R15341 DVSS.n5562 DVSS.n811 0.214786
R15342 DVSS.n5563 DVSS.n810 0.214786
R15343 DVSS.n809 DVSS.n807 0.214786
R15344 DVSS.n5567 DVSS.n806 0.214786
R15345 DVSS.n5569 DVSS.n805 0.214786
R15346 DVSS.n753 DVSS.n752 0.214786
R15347 DVSS.n5573 DVSS.n751 0.214786
R15348 DVSS.n5574 DVSS.n750 0.214786
R15349 DVSS.n5575 DVSS.n749 0.214786
R15350 DVSS.n748 DVSS.n746 0.214786
R15351 DVSS.n5579 DVSS.n745 0.214786
R15352 DVSS.n5580 DVSS.n744 0.214786
R15353 DVSS.n5581 DVSS.n743 0.214786
R15354 DVSS.n742 DVSS.n740 0.214786
R15355 DVSS.n5585 DVSS.n739 0.214786
R15356 DVSS.n5586 DVSS.n738 0.214786
R15357 DVSS.n5587 DVSS.n737 0.214786
R15358 DVSS.n736 DVSS.n734 0.214786
R15359 DVSS.n5591 DVSS.n733 0.214786
R15360 DVSS.n5592 DVSS.n732 0.214786
R15361 DVSS.n5593 DVSS.n731 0.214786
R15362 DVSS.n147 DVSS.n145 0.214786
R15363 DVSS.n5598 DVSS.n5597 0.214786
R15364 DVSS.n146 DVSS.n144 0.214786
R15365 DVSS.n727 DVSS.n726 0.214786
R15366 DVSS.n725 DVSS.n149 0.214786
R15367 DVSS.n724 DVSS.n723 0.214786
R15368 DVSS.n151 DVSS.n150 0.214786
R15369 DVSS.n718 DVSS.n717 0.214786
R15370 DVSS.n154 DVSS.n153 0.214786
R15371 DVSS.n541 DVSS.n540 0.214786
R15372 DVSS.n544 DVSS.n539 0.214786
R15373 DVSS.n545 DVSS.n538 0.214786
R15374 DVSS.n546 DVSS.n537 0.214786
R15375 DVSS.n536 DVSS.n534 0.214786
R15376 DVSS.n550 DVSS.n533 0.214786
R15377 DVSS.n551 DVSS.n532 0.214786
R15378 DVSS.n552 DVSS.n531 0.214786
R15379 DVSS.n530 DVSS.n528 0.214786
R15380 DVSS.n556 DVSS.n527 0.214786
R15381 DVSS.n557 DVSS.n526 0.214786
R15382 DVSS.n558 DVSS.n525 0.214786
R15383 DVSS.n524 DVSS.n522 0.214786
R15384 DVSS.n562 DVSS.n521 0.214786
R15385 DVSS.n563 DVSS.n520 0.214786
R15386 DVSS.n564 DVSS.n519 0.214786
R15387 DVSS.n518 DVSS.n516 0.214786
R15388 DVSS.n568 DVSS.n515 0.214786
R15389 DVSS.n569 DVSS.n514 0.214786
R15390 DVSS.n570 DVSS.n513 0.214786
R15391 DVSS.n206 DVSS.n205 0.214786
R15392 DVSS.n575 DVSS.n574 0.214786
R15393 DVSS.n509 DVSS.n204 0.214786
R15394 DVSS.n508 DVSS.n507 0.214786
R15395 DVSS.n506 DVSS.n208 0.214786
R15396 DVSS.n505 DVSS.n504 0.214786
R15397 DVSS.n499 DVSS.n498 0.214786
R15398 DVSS.n496 DVSS.n211 0.214786
R15399 DVSS.n495 DVSS.n494 0.214786
R15400 DVSS.n213 DVSS.n212 0.214786
R15401 DVSS.n490 DVSS.n489 0.214786
R15402 DVSS.n488 DVSS.n215 0.214786
R15403 DVSS.n487 DVSS.n486 0.214786
R15404 DVSS.n217 DVSS.n216 0.214786
R15405 DVSS.n482 DVSS.n481 0.214786
R15406 DVSS.n480 DVSS.n219 0.214786
R15407 DVSS.n479 DVSS.n478 0.214786
R15408 DVSS.n221 DVSS.n220 0.214786
R15409 DVSS.n474 DVSS.n473 0.214786
R15410 DVSS.n472 DVSS.n223 0.214786
R15411 DVSS.n471 DVSS.n470 0.214786
R15412 DVSS.n225 DVSS.n224 0.214786
R15413 DVSS.n466 DVSS.n465 0.214786
R15414 DVSS.n367 DVSS.n366 0.214786
R15415 DVSS.n5547 DVSS.n825 0.214786
R15416 DVSS.n5549 DVSS.n5548 0.214786
R15417 DVSS.n5550 DVSS.n820 0.214786
R15418 DVSS.n5552 DVSS.n5551 0.214786
R15419 DVSS.n5553 DVSS.n819 0.214786
R15420 DVSS.n5555 DVSS.n5554 0.214786
R15421 DVSS.n5556 DVSS.n814 0.214786
R15422 DVSS.n5558 DVSS.n5557 0.214786
R15423 DVSS.n5559 DVSS.n813 0.214786
R15424 DVSS.n5561 DVSS.n5560 0.214786
R15425 DVSS.n5562 DVSS.n808 0.214786
R15426 DVSS.n5564 DVSS.n5563 0.214786
R15427 DVSS.n5565 DVSS.n807 0.214786
R15428 DVSS.n5567 DVSS.n5566 0.214786
R15429 DVSS.n5570 DVSS.n5569 0.214786
R15430 DVSS.n5571 DVSS.n752 0.214786
R15431 DVSS.n5573 DVSS.n5572 0.214786
R15432 DVSS.n5574 DVSS.n747 0.214786
R15433 DVSS.n5576 DVSS.n5575 0.214786
R15434 DVSS.n5577 DVSS.n746 0.214786
R15435 DVSS.n5579 DVSS.n5578 0.214786
R15436 DVSS.n5580 DVSS.n741 0.214786
R15437 DVSS.n5582 DVSS.n5581 0.214786
R15438 DVSS.n5583 DVSS.n740 0.214786
R15439 DVSS.n5585 DVSS.n5584 0.214786
R15440 DVSS.n5586 DVSS.n735 0.214786
R15441 DVSS.n5588 DVSS.n5587 0.214786
R15442 DVSS.n5589 DVSS.n734 0.214786
R15443 DVSS.n5591 DVSS.n5590 0.214786
R15444 DVSS.n5592 DVSS.n730 0.214786
R15445 DVSS.n5594 DVSS.n5593 0.214786
R15446 DVSS.n5595 DVSS.n147 0.214786
R15447 DVSS.n5597 DVSS.n5596 0.214786
R15448 DVSS.n729 DVSS.n146 0.214786
R15449 DVSS.n728 DVSS.n727 0.214786
R15450 DVSS.n149 DVSS.n148 0.214786
R15451 DVSS.n723 DVSS.n722 0.214786
R15452 DVSS.n721 DVSS.n151 0.214786
R15453 DVSS.n719 DVSS.n718 0.214786
R15454 DVSS.n153 DVSS.n152 0.214786
R15455 DVSS.n542 DVSS.n541 0.214786
R15456 DVSS.n544 DVSS.n543 0.214786
R15457 DVSS.n545 DVSS.n535 0.214786
R15458 DVSS.n547 DVSS.n546 0.214786
R15459 DVSS.n548 DVSS.n534 0.214786
R15460 DVSS.n550 DVSS.n549 0.214786
R15461 DVSS.n551 DVSS.n529 0.214786
R15462 DVSS.n553 DVSS.n552 0.214786
R15463 DVSS.n554 DVSS.n528 0.214786
R15464 DVSS.n556 DVSS.n555 0.214786
R15465 DVSS.n557 DVSS.n523 0.214786
R15466 DVSS.n559 DVSS.n558 0.214786
R15467 DVSS.n560 DVSS.n522 0.214786
R15468 DVSS.n562 DVSS.n561 0.214786
R15469 DVSS.n563 DVSS.n517 0.214786
R15470 DVSS.n565 DVSS.n564 0.214786
R15471 DVSS.n566 DVSS.n516 0.214786
R15472 DVSS.n568 DVSS.n567 0.214786
R15473 DVSS.n569 DVSS.n512 0.214786
R15474 DVSS.n571 DVSS.n570 0.214786
R15475 DVSS.n572 DVSS.n206 0.214786
R15476 DVSS.n574 DVSS.n573 0.214786
R15477 DVSS.n510 DVSS.n509 0.214786
R15478 DVSS.n508 DVSS.n207 0.214786
R15479 DVSS.n502 DVSS.n208 0.214786
R15480 DVSS.n504 DVSS.n503 0.214786
R15481 DVSS.n501 DVSS.n209 0.214786
R15482 DVSS.n500 DVSS.n499 0.214786
R15483 DVSS.n211 DVSS.n210 0.214786
R15484 DVSS.n494 DVSS.n493 0.214786
R15485 DVSS.n492 DVSS.n213 0.214786
R15486 DVSS.n491 DVSS.n490 0.214786
R15487 DVSS.n215 DVSS.n214 0.214786
R15488 DVSS.n486 DVSS.n485 0.214786
R15489 DVSS.n484 DVSS.n217 0.214786
R15490 DVSS.n483 DVSS.n482 0.214786
R15491 DVSS.n219 DVSS.n218 0.214786
R15492 DVSS.n478 DVSS.n477 0.214786
R15493 DVSS.n476 DVSS.n221 0.214786
R15494 DVSS.n475 DVSS.n474 0.214786
R15495 DVSS.n223 DVSS.n222 0.214786
R15496 DVSS.n470 DVSS.n469 0.214786
R15497 DVSS.n468 DVSS.n225 0.214786
R15498 DVSS.n467 DVSS.n466 0.214786
R15499 DVSS.n368 DVSS.n367 0.214786
R15500 DVSS.n227 DVSS.n226 0.214786
R15501 DVSS.n228 DVSS.n227 0.214786
R15502 DVSS.n5 DVSS.n3 0.214786
R15503 DVSS.n4 DVSS.n2 0.214786
R15504 DVSS.n5801 DVSS.n1 0.214786
R15505 DVSS.n5740 DVSS.n0 0.214786
R15506 DVSS.n5744 DVSS.n5741 0.214786
R15507 DVSS.n5745 DVSS.n5739 0.214786
R15508 DVSS.n5746 DVSS.n5738 0.214786
R15509 DVSS.n5737 DVSS.n5735 0.214786
R15510 DVSS.n5750 DVSS.n5734 0.214786
R15511 DVSS.n5751 DVSS.n5733 0.214786
R15512 DVSS.n5752 DVSS.n5732 0.214786
R15513 DVSS.n5731 DVSS.n5729 0.214786
R15514 DVSS.n5756 DVSS.n5728 0.214786
R15515 DVSS.n5757 DVSS.n5727 0.214786
R15516 DVSS.n5758 DVSS.n5726 0.214786
R15517 DVSS.n5724 DVSS.n5723 0.214786
R15518 DVSS.n5722 DVSS.n50 0.214786
R15519 DVSS.n54 DVSS.n49 0.214786
R15520 DVSS.n5718 DVSS.n5717 0.214786
R15521 DVSS.n53 DVSS.n52 0.214786
R15522 DVSS.n5621 DVSS.n5620 0.214786
R15523 DVSS.n5619 DVSS.n5618 0.214786
R15524 DVSS.n5625 DVSS.n5617 0.214786
R15525 DVSS.n5626 DVSS.n5616 0.214786
R15526 DVSS.n5627 DVSS.n5615 0.214786
R15527 DVSS.n5614 DVSS.n5612 0.214786
R15528 DVSS.n5631 DVSS.n5611 0.214786
R15529 DVSS.n5632 DVSS.n5610 0.214786
R15530 DVSS.n5633 DVSS.n5609 0.214786
R15531 DVSS.n5608 DVSS.n5606 0.214786
R15532 DVSS.n5637 DVSS.n5605 0.214786
R15533 DVSS.n5638 DVSS.n5604 0.214786
R15534 DVSS.n5639 DVSS.n5603 0.214786
R15535 DVSS.n5602 DVSS.n142 0.214786
R15536 DVSS.n5643 DVSS.n141 0.214786
R15537 DVSS.n5644 DVSS.n140 0.214786
R15538 DVSS.n5645 DVSS.n139 0.214786
R15539 DVSS.n138 DVSS.n136 0.214786
R15540 DVSS.n5649 DVSS.n135 0.214786
R15541 DVSS.n714 DVSS.n134 0.214786
R15542 DVSS.n713 DVSS.n712 0.214786
R15543 DVSS.n157 DVSS.n156 0.214786
R15544 DVSS.n707 DVSS.n706 0.214786
R15545 DVSS.n705 DVSS.n159 0.214786
R15546 DVSS.n704 DVSS.n703 0.214786
R15547 DVSS.n161 DVSS.n160 0.214786
R15548 DVSS.n699 DVSS.n698 0.214786
R15549 DVSS.n697 DVSS.n163 0.214786
R15550 DVSS.n696 DVSS.n695 0.214786
R15551 DVSS.n165 DVSS.n164 0.214786
R15552 DVSS.n691 DVSS.n690 0.214786
R15553 DVSS.n168 DVSS.n167 0.214786
R15554 DVSS.n594 DVSS.n593 0.214786
R15555 DVSS.n592 DVSS.n591 0.214786
R15556 DVSS.n598 DVSS.n590 0.214786
R15557 DVSS.n599 DVSS.n589 0.214786
R15558 DVSS.n600 DVSS.n588 0.214786
R15559 DVSS.n587 DVSS.n585 0.214786
R15560 DVSS.n604 DVSS.n584 0.214786
R15561 DVSS.n605 DVSS.n583 0.214786
R15562 DVSS.n606 DVSS.n582 0.214786
R15563 DVSS.n581 DVSS.n579 0.214786
R15564 DVSS.n610 DVSS.n578 0.214786
R15565 DVSS.n612 DVSS.n202 0.214786
R15566 DVSS.n613 DVSS.n201 0.214786
R15567 DVSS.n198 DVSS.n196 0.214786
R15568 DVSS.n618 DVSS.n617 0.214786
R15569 DVSS.n197 DVSS.n195 0.214786
R15570 DVSS.n396 DVSS.n395 0.214786
R15571 DVSS.n399 DVSS.n394 0.214786
R15572 DVSS.n400 DVSS.n393 0.214786
R15573 DVSS.n401 DVSS.n392 0.214786
R15574 DVSS.n391 DVSS.n389 0.214786
R15575 DVSS.n405 DVSS.n388 0.214786
R15576 DVSS.n406 DVSS.n387 0.214786
R15577 DVSS.n407 DVSS.n386 0.214786
R15578 DVSS.n385 DVSS.n383 0.214786
R15579 DVSS.n411 DVSS.n382 0.214786
R15580 DVSS.n412 DVSS.n381 0.214786
R15581 DVSS.n413 DVSS.n380 0.214786
R15582 DVSS.n379 DVSS.n377 0.214786
R15583 DVSS.n417 DVSS.n376 0.214786
R15584 DVSS.n418 DVSS.n375 0.214786
R15585 DVSS.n419 DVSS.n374 0.214786
R15586 DVSS.n246 DVSS.n244 0.214786
R15587 DVSS.n424 DVSS.n423 0.214786
R15588 DVSS.n245 DVSS.n243 0.214786
R15589 DVSS.n5799 DVSS.n2 0.214786
R15590 DVSS.n5801 DVSS.n5800 0.214786
R15591 DVSS.n5742 DVSS.n0 0.214786
R15592 DVSS.n5744 DVSS.n5743 0.214786
R15593 DVSS.n5745 DVSS.n5736 0.214786
R15594 DVSS.n5747 DVSS.n5746 0.214786
R15595 DVSS.n5748 DVSS.n5735 0.214786
R15596 DVSS.n5750 DVSS.n5749 0.214786
R15597 DVSS.n5751 DVSS.n5730 0.214786
R15598 DVSS.n5753 DVSS.n5752 0.214786
R15599 DVSS.n5754 DVSS.n5729 0.214786
R15600 DVSS.n5756 DVSS.n5755 0.214786
R15601 DVSS.n5757 DVSS.n45 0.214786
R15602 DVSS.n5759 DVSS.n5758 0.214786
R15603 DVSS.n5723 DVSS.n44 0.214786
R15604 DVSS.n5722 DVSS.n5721 0.214786
R15605 DVSS.n5720 DVSS.n49 0.214786
R15606 DVSS.n5719 DVSS.n5718 0.214786
R15607 DVSS.n52 DVSS.n51 0.214786
R15608 DVSS.n5622 DVSS.n5621 0.214786
R15609 DVSS.n5623 DVSS.n5618 0.214786
R15610 DVSS.n5625 DVSS.n5624 0.214786
R15611 DVSS.n5626 DVSS.n5613 0.214786
R15612 DVSS.n5628 DVSS.n5627 0.214786
R15613 DVSS.n5629 DVSS.n5612 0.214786
R15614 DVSS.n5631 DVSS.n5630 0.214786
R15615 DVSS.n5632 DVSS.n5607 0.214786
R15616 DVSS.n5634 DVSS.n5633 0.214786
R15617 DVSS.n5635 DVSS.n5606 0.214786
R15618 DVSS.n5637 DVSS.n5636 0.214786
R15619 DVSS.n5638 DVSS.n143 0.214786
R15620 DVSS.n5640 DVSS.n5639 0.214786
R15621 DVSS.n5641 DVSS.n142 0.214786
R15622 DVSS.n5643 DVSS.n5642 0.214786
R15623 DVSS.n5644 DVSS.n137 0.214786
R15624 DVSS.n5646 DVSS.n5645 0.214786
R15625 DVSS.n5647 DVSS.n136 0.214786
R15626 DVSS.n5649 DVSS.n5648 0.214786
R15627 DVSS.n710 DVSS.n134 0.214786
R15628 DVSS.n712 DVSS.n711 0.214786
R15629 DVSS.n709 DVSS.n157 0.214786
R15630 DVSS.n708 DVSS.n707 0.214786
R15631 DVSS.n159 DVSS.n158 0.214786
R15632 DVSS.n703 DVSS.n702 0.214786
R15633 DVSS.n701 DVSS.n161 0.214786
R15634 DVSS.n700 DVSS.n699 0.214786
R15635 DVSS.n163 DVSS.n162 0.214786
R15636 DVSS.n695 DVSS.n694 0.214786
R15637 DVSS.n693 DVSS.n165 0.214786
R15638 DVSS.n692 DVSS.n691 0.214786
R15639 DVSS.n167 DVSS.n166 0.214786
R15640 DVSS.n595 DVSS.n594 0.214786
R15641 DVSS.n596 DVSS.n591 0.214786
R15642 DVSS.n598 DVSS.n597 0.214786
R15643 DVSS.n599 DVSS.n586 0.214786
R15644 DVSS.n601 DVSS.n600 0.214786
R15645 DVSS.n602 DVSS.n585 0.214786
R15646 DVSS.n604 DVSS.n603 0.214786
R15647 DVSS.n605 DVSS.n580 0.214786
R15648 DVSS.n607 DVSS.n606 0.214786
R15649 DVSS.n608 DVSS.n579 0.214786
R15650 DVSS.n610 DVSS.n609 0.214786
R15651 DVSS.n612 DVSS.n200 0.214786
R15652 DVSS.n614 DVSS.n613 0.214786
R15653 DVSS.n615 DVSS.n198 0.214786
R15654 DVSS.n617 DVSS.n616 0.214786
R15655 DVSS.n199 DVSS.n197 0.214786
R15656 DVSS.n397 DVSS.n396 0.214786
R15657 DVSS.n399 DVSS.n398 0.214786
R15658 DVSS.n400 DVSS.n390 0.214786
R15659 DVSS.n402 DVSS.n401 0.214786
R15660 DVSS.n403 DVSS.n389 0.214786
R15661 DVSS.n405 DVSS.n404 0.214786
R15662 DVSS.n406 DVSS.n384 0.214786
R15663 DVSS.n408 DVSS.n407 0.214786
R15664 DVSS.n409 DVSS.n383 0.214786
R15665 DVSS.n411 DVSS.n410 0.214786
R15666 DVSS.n412 DVSS.n378 0.214786
R15667 DVSS.n414 DVSS.n413 0.214786
R15668 DVSS.n415 DVSS.n377 0.214786
R15669 DVSS.n417 DVSS.n416 0.214786
R15670 DVSS.n418 DVSS.n372 0.214786
R15671 DVSS.n420 DVSS.n419 0.214786
R15672 DVSS.n421 DVSS.n246 0.214786
R15673 DVSS.n423 DVSS.n422 0.214786
R15674 DVSS.n371 DVSS.n245 0.214786
R15675 DVSS.n27 DVSS.n26 0.214786
R15676 DVSS.n5790 DVSS.n5789 0.214786
R15677 DVSS.n5788 DVSS.n29 0.214786
R15678 DVSS.n5787 DVSS.n5786 0.214786
R15679 DVSS.n5783 DVSS.n5782 0.214786
R15680 DVSS.n5781 DVSS.n31 0.214786
R15681 DVSS.n5780 DVSS.n5779 0.214786
R15682 DVSS.n33 DVSS.n32 0.214786
R15683 DVSS.n5775 DVSS.n5774 0.214786
R15684 DVSS.n5773 DVSS.n35 0.214786
R15685 DVSS.n5772 DVSS.n5771 0.214786
R15686 DVSS.n37 DVSS.n36 0.214786
R15687 DVSS.n5767 DVSS.n5766 0.214786
R15688 DVSS.n5765 DVSS.n39 0.214786
R15689 DVSS.n5764 DVSS.n5763 0.214786
R15690 DVSS.n107 DVSS.n106 0.214786
R15691 DVSS.n108 DVSS.n103 0.214786
R15692 DVSS.n5700 DVSS.n5699 0.214786
R15693 DVSS.n104 DVSS.n102 0.214786
R15694 DVSS.n5694 DVSS.n5693 0.214786
R15695 DVSS.n5692 DVSS.n110 0.214786
R15696 DVSS.n5691 DVSS.n5690 0.214786
R15697 DVSS.n112 DVSS.n111 0.214786
R15698 DVSS.n5686 DVSS.n5685 0.214786
R15699 DVSS.n5684 DVSS.n114 0.214786
R15700 DVSS.n5683 DVSS.n5682 0.214786
R15701 DVSS.n116 DVSS.n115 0.214786
R15702 DVSS.n5678 DVSS.n5677 0.214786
R15703 DVSS.n5676 DVSS.n118 0.214786
R15704 DVSS.n5675 DVSS.n5674 0.214786
R15705 DVSS.n120 DVSS.n119 0.214786
R15706 DVSS.n5670 DVSS.n5669 0.214786
R15707 DVSS.n5668 DVSS.n122 0.214786
R15708 DVSS.n5667 DVSS.n5666 0.214786
R15709 DVSS.n5660 DVSS.n124 0.214786
R15710 DVSS.n5662 DVSS.n5661 0.214786
R15711 DVSS.n5659 DVSS.n126 0.214786
R15712 DVSS.n5658 DVSS.n5657 0.214786
R15713 DVSS.n128 DVSS.n127 0.214786
R15714 DVSS.n5652 DVSS.n132 0.214786
R15715 DVSS.n668 DVSS.n131 0.214786
R15716 DVSS.n670 DVSS.n669 0.214786
R15717 DVSS.n673 DVSS.n667 0.214786
R15718 DVSS.n674 DVSS.n666 0.214786
R15719 DVSS.n675 DVSS.n665 0.214786
R15720 DVSS.n664 DVSS.n662 0.214786
R15721 DVSS.n679 DVSS.n661 0.214786
R15722 DVSS.n680 DVSS.n660 0.214786
R15723 DVSS.n681 DVSS.n659 0.214786
R15724 DVSS.n173 DVSS.n171 0.214786
R15725 DVSS.n686 DVSS.n685 0.214786
R15726 DVSS.n172 DVSS.n170 0.214786
R15727 DVSS.n655 DVSS.n654 0.214786
R15728 DVSS.n653 DVSS.n175 0.214786
R15729 DVSS.n652 DVSS.n651 0.214786
R15730 DVSS.n177 DVSS.n176 0.214786
R15731 DVSS.n647 DVSS.n646 0.214786
R15732 DVSS.n645 DVSS.n179 0.214786
R15733 DVSS.n644 DVSS.n643 0.214786
R15734 DVSS.n181 DVSS.n180 0.214786
R15735 DVSS.n639 DVSS.n638 0.214786
R15736 DVSS.n637 DVSS.n183 0.214786
R15737 DVSS.n636 DVSS.n635 0.214786
R15738 DVSS.n631 DVSS.n630 0.214786
R15739 DVSS.n629 DVSS.n188 0.214786
R15740 DVSS.n628 DVSS.n627 0.214786
R15741 DVSS.n190 DVSS.n189 0.214786
R15742 DVSS.n623 DVSS.n622 0.214786
R15743 DVSS.n193 DVSS.n192 0.214786
R15744 DVSS.n333 DVSS.n332 0.214786
R15745 DVSS.n336 DVSS.n331 0.214786
R15746 DVSS.n337 DVSS.n330 0.214786
R15747 DVSS.n338 DVSS.n329 0.214786
R15748 DVSS.n328 DVSS.n326 0.214786
R15749 DVSS.n342 DVSS.n325 0.214786
R15750 DVSS.n343 DVSS.n324 0.214786
R15751 DVSS.n344 DVSS.n323 0.214786
R15752 DVSS.n322 DVSS.n320 0.214786
R15753 DVSS.n348 DVSS.n319 0.214786
R15754 DVSS.n349 DVSS.n318 0.214786
R15755 DVSS.n350 DVSS.n317 0.214786
R15756 DVSS.n316 DVSS.n314 0.214786
R15757 DVSS.n354 DVSS.n313 0.214786
R15758 DVSS.n355 DVSS.n312 0.214786
R15759 DVSS.n356 DVSS.n258 0.214786
R15760 DVSS.n257 DVSS.n255 0.214786
R15761 DVSS.n361 DVSS.n360 0.214786
R15762 DVSS.n5791 DVSS.n5790 0.214786
R15763 DVSS.n29 DVSS.n28 0.214786
R15764 DVSS.n5786 DVSS.n5785 0.214786
R15765 DVSS.n5784 DVSS.n5783 0.214786
R15766 DVSS.n31 DVSS.n30 0.214786
R15767 DVSS.n5779 DVSS.n5778 0.214786
R15768 DVSS.n5777 DVSS.n33 0.214786
R15769 DVSS.n5776 DVSS.n5775 0.214786
R15770 DVSS.n35 DVSS.n34 0.214786
R15771 DVSS.n5771 DVSS.n5770 0.214786
R15772 DVSS.n5769 DVSS.n37 0.214786
R15773 DVSS.n5768 DVSS.n5767 0.214786
R15774 DVSS.n39 DVSS.n38 0.214786
R15775 DVSS.n5763 DVSS.n5762 0.214786
R15776 DVSS.n107 DVSS.n42 0.214786
R15777 DVSS.n5697 DVSS.n108 0.214786
R15778 DVSS.n5699 DVSS.n5698 0.214786
R15779 DVSS.n5696 DVSS.n104 0.214786
R15780 DVSS.n5695 DVSS.n5694 0.214786
R15781 DVSS.n110 DVSS.n109 0.214786
R15782 DVSS.n5690 DVSS.n5689 0.214786
R15783 DVSS.n5688 DVSS.n112 0.214786
R15784 DVSS.n5687 DVSS.n5686 0.214786
R15785 DVSS.n114 DVSS.n113 0.214786
R15786 DVSS.n5682 DVSS.n5681 0.214786
R15787 DVSS.n5680 DVSS.n116 0.214786
R15788 DVSS.n5679 DVSS.n5678 0.214786
R15789 DVSS.n118 DVSS.n117 0.214786
R15790 DVSS.n5674 DVSS.n5673 0.214786
R15791 DVSS.n5672 DVSS.n120 0.214786
R15792 DVSS.n5671 DVSS.n5670 0.214786
R15793 DVSS.n122 DVSS.n121 0.214786
R15794 DVSS.n5666 DVSS.n5665 0.214786
R15795 DVSS.n5664 DVSS.n124 0.214786
R15796 DVSS.n5663 DVSS.n5662 0.214786
R15797 DVSS.n126 DVSS.n125 0.214786
R15798 DVSS.n5657 DVSS.n5656 0.214786
R15799 DVSS.n5655 DVSS.n128 0.214786
R15800 DVSS.n5653 DVSS.n5652 0.214786
R15801 DVSS.n131 DVSS.n130 0.214786
R15802 DVSS.n671 DVSS.n670 0.214786
R15803 DVSS.n673 DVSS.n672 0.214786
R15804 DVSS.n674 DVSS.n663 0.214786
R15805 DVSS.n676 DVSS.n675 0.214786
R15806 DVSS.n677 DVSS.n662 0.214786
R15807 DVSS.n679 DVSS.n678 0.214786
R15808 DVSS.n680 DVSS.n658 0.214786
R15809 DVSS.n682 DVSS.n681 0.214786
R15810 DVSS.n683 DVSS.n173 0.214786
R15811 DVSS.n685 DVSS.n684 0.214786
R15812 DVSS.n657 DVSS.n172 0.214786
R15813 DVSS.n656 DVSS.n655 0.214786
R15814 DVSS.n175 DVSS.n174 0.214786
R15815 DVSS.n651 DVSS.n650 0.214786
R15816 DVSS.n649 DVSS.n177 0.214786
R15817 DVSS.n648 DVSS.n647 0.214786
R15818 DVSS.n179 DVSS.n178 0.214786
R15819 DVSS.n643 DVSS.n642 0.214786
R15820 DVSS.n641 DVSS.n181 0.214786
R15821 DVSS.n640 DVSS.n639 0.214786
R15822 DVSS.n183 DVSS.n182 0.214786
R15823 DVSS.n635 DVSS.n634 0.214786
R15824 DVSS.n632 DVSS.n631 0.214786
R15825 DVSS.n188 DVSS.n187 0.214786
R15826 DVSS.n627 DVSS.n626 0.214786
R15827 DVSS.n625 DVSS.n190 0.214786
R15828 DVSS.n624 DVSS.n623 0.214786
R15829 DVSS.n192 DVSS.n191 0.214786
R15830 DVSS.n334 DVSS.n333 0.214786
R15831 DVSS.n336 DVSS.n335 0.214786
R15832 DVSS.n337 DVSS.n327 0.214786
R15833 DVSS.n339 DVSS.n338 0.214786
R15834 DVSS.n340 DVSS.n326 0.214786
R15835 DVSS.n342 DVSS.n341 0.214786
R15836 DVSS.n343 DVSS.n321 0.214786
R15837 DVSS.n345 DVSS.n344 0.214786
R15838 DVSS.n346 DVSS.n320 0.214786
R15839 DVSS.n348 DVSS.n347 0.214786
R15840 DVSS.n349 DVSS.n315 0.214786
R15841 DVSS.n351 DVSS.n350 0.214786
R15842 DVSS.n352 DVSS.n314 0.214786
R15843 DVSS.n354 DVSS.n353 0.214786
R15844 DVSS.n355 DVSS.n256 0.214786
R15845 DVSS.n357 DVSS.n356 0.214786
R15846 DVSS.n358 DVSS.n255 0.214786
R15847 DVSS.n360 DVSS.n359 0.214786
R15848 DVSS.n4307 DVSS.n1455 0.212265
R15849 DVSS.n1370 DVSS.n1369 0.201836
R15850 DVSS.n4316 DVSS.n4315 0.192412
R15851 DVSS.n3788 VSS 0.189765
R15852 VSS DVSS.n3788 0.189765
R15853 DVSS.n1837 DVSS 0.186337
R15854 DVSS.n4179 DVSS.n4178 0.186214
R15855 DVSS.n4178 DVSS.n4177 0.186214
R15856 DVSS.n1254 DVSS.n1249 0.186214
R15857 DVSS.n1256 DVSS.n1254 0.186214
R15858 DVSS.n5343 DVSS.n5342 0.185484
R15859 VSS DVSS.n4115 0.17855
R15860 DVSS.n3817 DVSS.n3805 0.178408
R15861 DVSS.n3817 DVSS.n1802 0.178408
R15862 DVSS.n1823 DVSS.n1796 0.178408
R15863 DVSS.n3817 DVSS.n3804 0.178408
R15864 DVSS.n1825 DVSS.n1796 0.178408
R15865 DVSS.n3817 DVSS.n3803 0.178408
R15866 DVSS.n1844 DVSS.n1796 0.178408
R15867 DVSS.n1513 DVSS.n1512 0.175807
R15868 DVSS.n1466 DVSS 0.175204
R15869 DVSS.n1471 DVSS 0.175204
R15870 DVSS.n1253 DVSS 0.175204
R15871 DVSS.n1232 DVSS 0.175204
R15872 DVSS.n5702 DVSS.n5701 0.173577
R15873 DVSS.n311 DVSS.n310 0.173577
R15874 VSS DVSS.n4095 0.169912
R15875 DVSS.n5044 DVSS.n1109 0.168658
R15876 DVSS.n1119 DVSS.n1109 0.168658
R15877 DVSS.n5034 DVSS.n5033 0.168658
R15878 DVSS.n5033 DVSS.n1121 0.168658
R15879 DVSS.n4175 DVSS.n1516 0.166289
R15880 DVSS.n5601 DVSS.n5600 0.163909
R15881 DVSS.n689 DVSS.n688 0.163909
R15882 DVSS.n620 DVSS.n619 0.163909
R15883 DVSS.n427 DVSS.n241 0.161214
R15884 DVSS.n765 DVSS.n57 0.161214
R15885 DVSS.n5543 DVSS.n5541 0.149124
R15886 DVSS.n2661 DVSS.n1556 0.145461
R15887 DVSS.n3853 DVSS 0.144526
R15888 DVSS.n4108 DVSS 0.1436
R15889 DVSS DVSS.n4107 0.1436
R15890 DVSS.n4107 DVSS 0.1436
R15891 DVSS DVSS.n4106 0.1436
R15892 DVSS DVSS.n3934 0.143441
R15893 DVSS.n3932 DVSS 0.143441
R15894 DVSS DVSS.n4054 0.143441
R15895 DVSS.n4052 DVSS 0.143441
R15896 DVSS.n802 DVSS.n801 0.141125
R15897 DVSS.n464 DVSS.n463 0.141125
R15898 DVSS.n3934 DVSS.n3933 0.140794
R15899 DVSS.n3933 DVSS.n3932 0.140794
R15900 DVSS.n4054 DVSS.n4053 0.140794
R15901 DVSS.n4053 DVSS.n4052 0.140794
R15902 DVSS.n3789 VSS 0.139932
R15903 DVSS.n2619 DVSS 0.138622
R15904 DVSS.n803 DVSS.n754 0.137596
R15905 DVSS.n461 DVSS.n229 0.137559
R15906 DVSS.n1848 DVSS 0.1355
R15907 DVSS DVSS.n1476 0.1355
R15908 DVSS.n5706 DVSS.n61 0.130943
R15909 DVSS.n2410 DVSS 0.130618
R15910 DVSS.n1762 DVSS 0.130618
R15911 DVSS.n260 DVSS.n60 0.130587
R15912 DVSS.n2092 DVSS 0.130161
R15913 DVSS.n3955 DVSS.n1685 0.129687
R15914 DVSS.n1728 DVSS.n1727 0.129687
R15915 DVSS.n1700 DVSS.n1699 0.129687
R15916 DVSS.n1702 DVSS.n1701 0.129687
R15917 DVSS.n3931 DVSS.n1706 0.129687
R15918 DVSS.n3943 DVSS.n3942 0.129687
R15919 DVSS.n4011 DVSS.n4010 0.129687
R15920 DVSS.n1614 DVSS.n1613 0.129687
R15921 DVSS.n1616 DVSS.n1615 0.129687
R15922 DVSS.n1619 DVSS.n1618 0.129687
R15923 DVSS.n1622 DVSS.n1621 0.129687
R15924 DVSS.n4049 DVSS.n1626 0.129687
R15925 DVSS.n955 DVSS.n954 0.129009
R15926 DVSS.n2312 DVSS.n1928 0.128608
R15927 DVSS.n2539 DVSS.n2312 0.128203
R15928 DVSS DVSS.n856 0.125798
R15929 DVSS.n856 DVSS.n855 0.12265
R15930 DVSS.n2627 DVSS 0.122025
R15931 DVSS DVSS.n1841 0.115647
R15932 DVSS.n1931 DVSS.n1930 0.114824
R15933 DVSS.n2540 DVSS.n1922 0.114824
R15934 DVSS.n5792 DVSS.n5791 0.114699
R15935 DVSS.n5799 DVSS.n5798 0.114699
R15936 DVSS.n5547 DVSS.n5546 0.114699
R15937 DVSS.n4804 DVSS.n4803 0.114184
R15938 DVSS.n4185 DVSS.n4184 0.114184
R15939 DVSS.n1976 DVSS.n1975 0.114184
R15940 DVSS.n1265 DVSS.n1264 0.114184
R15941 DVSS.n1347 DVSS.n1346 0.114184
R15942 DVSS.n2640 VSS 0.113
R15943 VSS DVSS.n2658 0.113
R15944 DVSS.n3780 VSS 0.113
R15945 DVSS DVSS.n3853 0.111845
R15946 DVSS.n4102 DVSS 0.111373
R15947 DVSS.n4773 DVSS.n1353 0.110634
R15948 DVSS.n2647 VSS 0.110353
R15949 DVSS.n2551 DVSS.n1901 0.109959
R15950 DVSS.n2552 DVSS.n2551 0.109959
R15951 DVSS.n4110 DVSS.n4109 0.109729
R15952 DVSS.n4105 DVSS.n4103 0.109572
R15953 DVSS.n5716 DVSS.n5715 0.107643
R15954 DVSS.n373 DVSS.n242 0.107643
R15955 DVSS DVSS.n4102 0.107291
R15956 DVSS.n1120 DVSS.n1119 0.107079
R15957 DVSS.n1500 DVSS.n1483 0.105895
R15958 DVSS.n954 DVSS.n949 0.102277
R15959 DVSS.n4107 DVSS 0.102157
R15960 DVSS.n5336 DVSS.n5335 0.101471
R15961 DVSS.n5096 DVSS.n5095 0.101471
R15962 DVSS DVSS.n2092 0.101206
R15963 DVSS DVSS.n2410 0.10093
R15964 DVSS.n1762 DVSS 0.10093
R15965 DVSS DVSS.n1547 0.0991804
R15966 DVSS.n5344 DVSS.n5343 0.0985668
R15967 DVSS.n5343 DVSS.n952 0.0982447
R15968 DVSS.n1212 DVSS 0.0942039
R15969 DVSS.n1475 DVSS 0.0942039
R15970 DVSS.n1220 DVSS 0.0942039
R15971 DVSS.n1207 DVSS 0.0942039
R15972 DVSS.n1516 VSS 0.0928684
R15973 DVSS.n2681 DVSS.n2667 0.0921154
R15974 DVSS.n4315 DVSS.n4314 0.0891765
R15975 DVSS.n4166 DVSS.n4165 0.0883604
R15976 DVSS.n1827 DVSS 0.0871834
R15977 DVSS.n1828 DVSS 0.0871834
R15978 DVSS.n4102 DVSS 0.0837012
R15979 DVSS.n4136 DVSS.n1522 0.08175
R15980 DVSS.n4160 DVSS.n4159 0.08175
R15981 DVSS DVSS.n1221 0.0812353
R15982 DVSS DVSS.n1208 0.0812353
R15983 DVSS DVSS.n4854 0.0812353
R15984 DVSS.n2533 DVSS.n1911 0.077375
R15985 DVSS.n2567 DVSS.n1903 0.077375
R15986 DVSS DVSS.n4307 0.0772647
R15987 DVSS.n3939 DVSS.n3938 0.0769706
R15988 DVSS.n3938 DVSS.n3937 0.0769706
R15989 DVSS.n1634 DVSS.n1631 0.0769376
R15990 DVSS.n2255 DVSS.n1926 0.0763777
R15991 DVSS.n3294 DVSS 0.0761
R15992 DVSS.n3005 DVSS 0.0761
R15993 DVSS DVSS.n3008 0.0761
R15994 DVSS.n3204 DVSS 0.0761
R15995 DVSS DVSS.n2877 0.0761
R15996 DVSS.n3173 DVSS 0.0761
R15997 DVSS DVSS.n2824 0.0761
R15998 DVSS.n3129 DVSS 0.0761
R15999 DVSS DVSS.n3017 0.0761
R16000 DVSS.n3018 DVSS 0.0761
R16001 DVSS DVSS.n2731 0.0761
R16002 DVSS.n3061 DVSS 0.0761
R16003 DVSS DVSS.n3024 0.0761
R16004 DVSS.n3025 DVSS 0.0761
R16005 DVSS.n2267 DVSS.n2255 0.0756596
R16006 DVSS.n4108 DVSS 0.0748392
R16007 DVSS.n4106 DVSS 0.0746758
R16008 DVSS.n2684 DVSS.n2681 0.0745555
R16009 DVSS.n1834 DVSS 0.0743218
R16010 DVSS.n1832 DVSS 0.0743218
R16011 DVSS.n4379 DVSS.n4343 0.0741096
R16012 DVSS.n3827 DVSS 0.0728785
R16013 DVSS DVSS.n1791 0.0728785
R16014 DVSS.n2018 DVSS.n2017 0.0728571
R16015 DVSS DVSS.n1836 0.0720477
R16016 DVSS.n2615 DVSS.n1849 0.0693638
R16017 DVSS.n4094 DVSS.n4093 0.0668158
R16018 DVSS.n4115 DVSS.n4114 0.0656316
R16019 DVSS.n4380 DVSS.n4379 0.0624601
R16020 DVSS.n5034 DVSS.n1120 0.0620789
R16021 DVSS.n1635 DVSS.n1634 0.0599397
R16022 DVSS.n5540 DVSS.n847 0.0597445
R16023 DVSS.n846 DVSS.n845 0.0597445
R16024 DVSS.n844 DVSS.n843 0.0597445
R16025 DVSS.n842 DVSS.n841 0.0597445
R16026 DVSS.n840 DVSS.n839 0.0597445
R16027 DVSS.n838 DVSS.n837 0.0597445
R16028 DVSS.n836 DVSS.n835 0.0597445
R16029 DVSS.n834 DVSS.n833 0.0597445
R16030 DVSS.n832 DVSS.n831 0.0597445
R16031 DVSS.n5542 DVSS.n830 0.0597445
R16032 DVSS.n25 DVSS.n24 0.0597445
R16033 DVSS.n23 DVSS.n22 0.0597445
R16034 DVSS.n21 DVSS.n20 0.0597445
R16035 DVSS.n19 DVSS.n18 0.0597445
R16036 DVSS.n17 DVSS.n16 0.0597445
R16037 DVSS.n15 DVSS.n14 0.0597445
R16038 DVSS.n13 DVSS.n12 0.0597445
R16039 DVSS.n11 DVSS.n10 0.0597445
R16040 DVSS.n9 DVSS.n8 0.0597445
R16041 DVSS.n5794 DVSS.n7 0.0597445
R16042 DVSS.n24 DVSS.n23 0.0597445
R16043 DVSS.n22 DVSS.n21 0.0597445
R16044 DVSS.n20 DVSS.n19 0.0597445
R16045 DVSS.n18 DVSS.n17 0.0597445
R16046 DVSS.n16 DVSS.n15 0.0597445
R16047 DVSS.n14 DVSS.n13 0.0597445
R16048 DVSS.n12 DVSS.n11 0.0597445
R16049 DVSS.n10 DVSS.n9 0.0597445
R16050 DVSS.n8 DVSS.n7 0.0597445
R16051 DVSS.n847 DVSS.n846 0.0597445
R16052 DVSS.n845 DVSS.n844 0.0597445
R16053 DVSS.n843 DVSS.n842 0.0597445
R16054 DVSS.n841 DVSS.n840 0.0597445
R16055 DVSS.n839 DVSS.n838 0.0597445
R16056 DVSS.n837 DVSS.n836 0.0597445
R16057 DVSS.n835 DVSS.n834 0.0597445
R16058 DVSS.n833 DVSS.n832 0.0597445
R16059 DVSS.n831 DVSS.n830 0.0597445
R16060 DVSS.n4369 DVSS.n4360 0.0588383
R16061 DVSS.n2538 DVSS.n2537 0.058625
R16062 DVSS.n2266 DVSS.n2265 0.058625
R16063 DVSS.n2611 DVSS.n1849 0.0585457
R16064 DVSS DVSS.n4804 0.0585263
R16065 DVSS.n4184 DVSS 0.0585263
R16066 DVSS.n1975 DVSS 0.0585263
R16067 DVSS DVSS.n1265 0.0585263
R16068 DVSS.n1346 DVSS 0.0585263
R16069 DVSS.n2019 DVSS.n2018 0.058308
R16070 DVSS DVSS.n1547 0.0574691
R16071 DVSS.n4652 DVSS.n1392 0.0562784
R16072 DVSS.n2312 DVSS.n2311 0.0546667
R16073 DVSS.n2311 DVSS.t14 0.0546667
R16074 DVSS.n2550 DVSS.t14 0.0546667
R16075 DVSS.n2551 DVSS.n2550 0.0546667
R16076 DVSS.n2535 DVSS.n2534 0.0544368
R16077 DVSS.n2536 DVSS.n2535 0.0544368
R16078 DVSS.n2263 DVSS.n2262 0.0544368
R16079 DVSS.n2263 DVSS.n2256 0.0544368
R16080 DVSS.n364 DVSS.n249 0.0532401
R16081 DVSS.n2595 DVSS.n1863 0.0532027
R16082 DVSS.n2483 DVSS.n2476 0.0532027
R16083 DVSS.n1392 DVSS.n1391 0.0500653
R16084 DVSS.n4139 DVSS.n4138 0.0495566
R16085 DVSS.n4164 DVSS.n4163 0.0495566
R16086 DVSS.n4159 DVSS.n4158 0.0486793
R16087 DVSS.n369 DVSS.n249 0.0485826
R16088 DVSS DVSS.n1551 0.0479398
R16089 DVSS DVSS.n4101 0.0479398
R16090 DVSS.n4300 DVSS 0.0456808
R16091 DVSS.n4302 DVSS 0.0456808
R16092 DVSS.n4306 DVSS 0.0456808
R16093 DVSS.n1685 DVSS 0.0456808
R16094 DVSS.n1727 DVSS 0.0456808
R16095 DVSS.n1699 DVSS 0.0456808
R16096 DVSS.n1701 DVSS 0.0456808
R16097 DVSS.n1706 DVSS 0.0456808
R16098 DVSS.n3942 DVSS 0.0456808
R16099 DVSS.n4010 DVSS 0.0456808
R16100 DVSS.n1613 DVSS 0.0456808
R16101 DVSS.n1615 DVSS 0.0456808
R16102 DVSS.n1618 DVSS 0.0456808
R16103 DVSS.n1621 DVSS 0.0456808
R16104 DVSS.n1626 DVSS 0.0456808
R16105 DVSS.n2522 DVSS.n2321 0.0450872
R16106 DVSS.n1942 DVSS.n1941 0.0450872
R16107 DVSS.n2306 DVSS.n1950 0.0450872
R16108 DVSS.n1895 DVSS.n1893 0.0450872
R16109 DVSS.n2479 DVSS.n2338 0.0450872
R16110 DVSS.n2593 DVSS.n2592 0.0450718
R16111 DVSS.n2592 DVSS.n2591 0.0450718
R16112 DVSS.n1871 DVSS.n1870 0.0450718
R16113 DVSS.n1872 DVSS.n1871 0.0450718
R16114 DVSS.n2334 DVSS.n2333 0.0450718
R16115 DVSS.n2335 DVSS.n2334 0.0450718
R16116 DVSS.n2495 DVSS.n2486 0.0442838
R16117 DVSS.n2545 DVSS.n1923 0.0442838
R16118 DVSS.n2497 DVSS.n2496 0.0442838
R16119 DVSS.n2496 DVSS.n2487 0.0442838
R16120 DVSS.n2490 DVSS.n2489 0.0442838
R16121 DVSS.n1943 DVSS.n1935 0.0442838
R16122 DVSS.n1944 DVSS.n1943 0.0442838
R16123 DVSS.n1949 DVSS.n1948 0.0442838
R16124 DVSS.n2595 DVSS.n2594 0.0442838
R16125 DVSS.n2590 DVSS.n2589 0.0442838
R16126 DVSS.n2589 DVSS.n1866 0.0442838
R16127 DVSS.n1890 DVSS.n1889 0.0442838
R16128 DVSS.n1891 DVSS.n1890 0.0442838
R16129 DVSS.n1896 DVSS.n1891 0.0442838
R16130 DVSS.n1897 DVSS.n1896 0.0442838
R16131 DVSS.n2572 DVSS.n1897 0.0442838
R16132 DVSS.n2572 DVSS.n2571 0.0442838
R16133 DVSS.n2571 DVSS.n1898 0.0442838
R16134 DVSS.n2322 DVSS.n1917 0.0442838
R16135 DVSS.n2326 DVSS.n2322 0.0442838
R16136 DVSS.n2327 DVSS.n2326 0.0442838
R16137 DVSS.n2521 DVSS.n2327 0.0442838
R16138 DVSS.n2521 DVSS.n2520 0.0442838
R16139 DVSS.n2520 DVSS.n2519 0.0442838
R16140 DVSS.n2519 DVSS.n2328 0.0442838
R16141 DVSS.n2515 DVSS.n2336 0.0442838
R16142 DVSS.n2515 DVSS.n2514 0.0442838
R16143 DVSS.n2514 DVSS.n2337 0.0442838
R16144 DVSS.n2478 DVSS.n2337 0.0442838
R16145 DVSS.n2482 DVSS.n2478 0.0442838
R16146 DVSS.n2483 DVSS.n2482 0.0442838
R16147 DVSS.n2247 DVSS.n1522 0.0432989
R16148 DVSS.n2518 DVSS.n2329 0.0430229
R16149 DVSS.n1892 DVSS.n1868 0.0430229
R16150 DVSS.n1945 DVSS.n1934 0.0426101
R16151 DVSS.n2513 DVSS.n2512 0.0421972
R16152 DVSS.n2352 DVSS.n2346 0.0418677
R16153 DVSS.n2585 DVSS.n1875 0.0418677
R16154 DVSS.n2494 DVSS.n2493 0.0418514
R16155 DVSS.n4763 DVSS.n1392 0.0417698
R16156 DVSS.n4763 DVSS.n4762 0.0417698
R16157 DVSS.n4360 DVSS.n4323 0.0417698
R16158 DVSS.n4323 DVSS.n4322 0.0417698
R16159 DVSS.n2325 DVSS.n2323 0.0405459
R16160 DVSS.n2573 DVSS.n1888 0.0405459
R16161 DVSS.n2822 DVSS.n1792 0.0398939
R16162 DVSS.n3512 DVSS.n1792 0.0398939
R16163 DVSS.n3130 DVSS.n1793 0.0398939
R16164 DVSS.n3512 DVSS.n1793 0.0398939
R16165 DVSS.n2597 DVSS.n2596 0.0397202
R16166 DVSS DVSS.n2665 0.0392931
R16167 DVSS.n3506 DVSS 0.0392931
R16168 DVSS.n2490 DVSS.n1920 0.0382027
R16169 DVSS.n1948 DVSS.n1933 0.0382027
R16170 DVSS.n2255 DVSS.n2254 0.0381812
R16171 DVSS.n2254 DVSS.t14 0.0381812
R16172 DVSS.n2486 DVSS.n2473 0.0373919
R16173 DVSS.n2014 DVSS.n1977 0.0359178
R16174 DVSS.n4141 DVSS.n4140 0.0357988
R16175 DVSS.n1552 DVSS 0.0351916
R16176 DVSS.n4109 DVSS 0.0351916
R16177 DVSS DVSS.n4100 0.0351154
R16178 DVSS.n4103 DVSS 0.0351154
R16179 VSS DVSS.n1515 0.0348421
R16180 DVSS.n2481 DVSS.n2480 0.0339404
R16181 DVSS.n363 DVSS.n248 0.033707
R16182 DVSS.n362 DVSS.n251 0.033707
R16183 DVSS.n4293 DVSS.n4292 0.0336579
R16184 DVSS.n4787 DVSS.n4786 0.0336579
R16185 DVSS.n1250 DVSS.n1233 0.0336579
R16186 DVSS.n4296 DVSS.n4295 0.0336579
R16187 DVSS.n2523 DVSS.n2320 0.0331147
R16188 DVSS.n1894 DVSS.n1887 0.0331147
R16189 DVSS.n4625 DVSS.n1371 0.033
R16190 DVSS.n4756 DVSS.n1371 0.033
R16191 DVSS.n4754 DVSS.n4753 0.033
R16192 DVSS.n4755 DVSS.n4754 0.033
R16193 DVSS.n4550 DVSS.n1394 0.033
R16194 DVSS.n1394 DVSS.n1393 0.033
R16195 DVSS.n4511 DVSS.n4510 0.033
R16196 DVSS.n4510 DVSS.n4509 0.033
R16197 DVSS.n4432 DVSS.n1449 0.033
R16198 DVSS.n4508 DVSS.n1449 0.033
R16199 DVSS.n4506 DVSS.n4505 0.033
R16200 DVSS.n4507 DVSS.n4506 0.033
R16201 DVSS.n4288 DVSS.n1476 0.0322647
R16202 DVSS.n2542 DVSS.n1927 0.031778
R16203 DVSS.n2303 DVSS.n2301 0.031778
R16204 DVSS.n3500 DVSS.n2672 0.0315
R16205 DVSS.n2710 DVSS.n2696 0.0315
R16206 DVSS.n2710 DVSS.n2708 0.0315
R16207 DVSS.n3460 DVSS.n3459 0.0315
R16208 DVSS.n2765 DVSS.n2761 0.0315
R16209 DVSS.n2801 DVSS.n2786 0.0315
R16210 DVSS.n3396 DVSS.n3395 0.0315
R16211 DVSS.n2857 DVSS.n2853 0.0315
R16212 DVSS.n2894 DVSS.n2879 0.0315
R16213 DVSS.n3331 DVSS.n3330 0.0315
R16214 DVSS.n3309 DVSS.n2946 0.0315
R16215 DVSS.n2982 DVSS.n2968 0.0315
R16216 DVSS.n2982 DVSS.n2980 0.0315
R16217 DVSS.n3268 DVSS.n3267 0.0315
R16218 DVSS.n3027 DVSS.n2668 0.0315
R16219 DVSS.n3045 DVSS.n3044 0.0315
R16220 DVSS.n3046 DVSS.n3045 0.0315
R16221 DVSS.n3063 DVSS.n3021 0.0315
R16222 DVSS.n3091 DVSS.n3090 0.0315
R16223 DVSS.n3112 DVSS.n3111 0.0315
R16224 DVSS.n3132 DVSS.n3014 0.0315
R16225 DVSS.n3160 DVSS.n3159 0.0315
R16226 DVSS.n3182 DVSS.n3181 0.0315
R16227 DVSS.n3202 DVSS.n3201 0.0315
R16228 DVSS.n3224 DVSS.n3223 0.0315
R16229 DVSS.n3242 DVSS.n3241 0.0315
R16230 DVSS.n3243 DVSS.n3242 0.0315
R16231 DVSS.n3260 DVSS.n3003 0.0315
R16232 DVSS.n1947 DVSS.n1932 0.0310505
R16233 DVSS.n3501 DVSS.n2671 0.031
R16234 DVSS.n3456 DVSS.n2732 0.031
R16235 DVSS.n3310 DVSS.n2945 0.031
R16236 DVSS.n3828 DVSS.n1789 0.031
R16237 DVSS.n3504 DVSS.n3503 0.031
R16238 DVSS.n3073 DVSS.n3072 0.031
R16239 DVSS.n3219 DVSS.n2942 0.031
R16240 DVSS.n3002 DVSS.n1788 0.031
R16241 DVSS.n2489 DVSS.n1922 0.0309054
R16242 DVSS.n1949 DVSS.n1931 0.0309054
R16243 DVSS.n2485 DVSS.n2484 0.0306376
R16244 DVSS.n2491 DVSS.n2488 0.0305
R16245 DVSS.n3436 DVSS.n3435 0.0305
R16246 DVSS.n3334 DVSS.n2911 0.0305
R16247 DVSS.n3094 DVSS.n2759 0.0305
R16248 DVSS.n3200 DVSS.n3198 0.0305
R16249 DVSS.n370 DVSS.n248 0.0304195
R16250 DVSS.n251 DVSS.n247 0.0304195
R16251 DVSS.n2517 DVSS.n2516 0.0302248
R16252 DVSS.n2588 DVSS.n2587 0.0302248
R16253 DVSS.n5541 DVSS.n25 0.0301222
R16254 DVSS.n5795 DVSS.n5794 0.0301222
R16255 DVSS.n5540 DVSS.n5539 0.0301222
R16256 DVSS.n5543 DVSS.n5542 0.0301222
R16257 DVSS.n2800 DVSS.n2798 0.03
R16258 DVSS.n3356 DVSS.n3355 0.03
R16259 DVSS.n3114 DVSS.n3113 0.03
R16260 DVSS.n3178 DVSS.n2881 0.03
R16261 DVSS.n1979 DVSS.n1977 0.0298971
R16262 DVSS.n3392 DVSS.n2823 0.0295
R16263 DVSS.n2856 DVSS.n2841 0.0295
R16264 DVSS.n3142 DVSS.n3141 0.0295
R16265 DVSS.n3156 DVSS.n3012 0.0295
R16266 DVSS.n3399 DVSS.n2819 0.029
R16267 DVSS.n3372 DVSS.n3371 0.029
R16268 DVSS.n3133 DVSS.n3015 0.029
R16269 DVSS.n3163 DVSS.n2851 0.029
R16270 DVSS.n1947 DVSS.n1946 0.0285734
R16271 DVSS.n3420 DVSS.n3419 0.0285
R16272 DVSS.n2893 DVSS.n2891 0.0285
R16273 DVSS.n3108 DVSS.n2788 0.0285
R16274 DVSS.n3184 DVSS.n3183 0.0285
R16275 DVSS.n800 DVSS.n799 0.0283304
R16276 DVSS.n799 DVSS.n755 0.0283304
R16277 DVSS.n795 DVSS.n755 0.0283304
R16278 DVSS.n795 DVSS.n794 0.0283304
R16279 DVSS.n794 DVSS.n793 0.0283304
R16280 DVSS.n793 DVSS.n757 0.0283304
R16281 DVSS.n789 DVSS.n757 0.0283304
R16282 DVSS.n789 DVSS.n788 0.0283304
R16283 DVSS.n788 DVSS.n787 0.0283304
R16284 DVSS.n787 DVSS.n759 0.0283304
R16285 DVSS.n783 DVSS.n759 0.0283304
R16286 DVSS.n783 DVSS.n782 0.0283304
R16287 DVSS.n782 DVSS.n781 0.0283304
R16288 DVSS.n781 DVSS.n761 0.0283304
R16289 DVSS.n777 DVSS.n761 0.0283304
R16290 DVSS.n777 DVSS.n776 0.0283304
R16291 DVSS.n776 DVSS.n775 0.0283304
R16292 DVSS.n775 DVSS.n763 0.0283304
R16293 DVSS.n771 DVSS.n763 0.0283304
R16294 DVSS.n771 DVSS.n770 0.0283304
R16295 DVSS.n770 DVSS.n769 0.0283304
R16296 DVSS.n769 DVSS.n766 0.0283304
R16297 DVSS.n5714 DVSS.n56 0.0283304
R16298 DVSS.n72 DVSS.n56 0.0283304
R16299 DVSS.n73 DVSS.n72 0.0283304
R16300 DVSS.n73 DVSS.n71 0.0283304
R16301 DVSS.n77 DVSS.n71 0.0283304
R16302 DVSS.n78 DVSS.n77 0.0283304
R16303 DVSS.n79 DVSS.n78 0.0283304
R16304 DVSS.n79 DVSS.n69 0.0283304
R16305 DVSS.n83 DVSS.n69 0.0283304
R16306 DVSS.n84 DVSS.n83 0.0283304
R16307 DVSS.n85 DVSS.n84 0.0283304
R16308 DVSS.n85 DVSS.n67 0.0283304
R16309 DVSS.n89 DVSS.n67 0.0283304
R16310 DVSS.n90 DVSS.n89 0.0283304
R16311 DVSS.n91 DVSS.n90 0.0283304
R16312 DVSS.n91 DVSS.n65 0.0283304
R16313 DVSS.n95 DVSS.n65 0.0283304
R16314 DVSS.n96 DVSS.n95 0.0283304
R16315 DVSS.n97 DVSS.n96 0.0283304
R16316 DVSS.n97 DVSS.n63 0.0283304
R16317 DVSS.n101 DVSS.n63 0.0283304
R16318 DVSS.n5704 DVSS.n5703 0.0283304
R16319 DVSS.n2516 DVSS.n2332 0.0281606
R16320 DVSS.n2492 DVSS.n2491 0.0280676
R16321 DVSS.n2764 DVSS.n2749 0.028
R16322 DVSS.n3329 DVSS.n2915 0.028
R16323 DVSS.n3087 DVSS.n3019 0.028
R16324 DVSS.n3206 DVSS.n2917 0.028
R16325 DVSS.n3499 DVSS.n2673 0.0279877
R16326 DVSS.n3499 DVSS.n3498 0.0279877
R16327 DVSS.n3498 DVSS.n3497 0.0279877
R16328 DVSS.n3497 DVSS.n2674 0.0279877
R16329 DVSS.n3486 DVSS.n2694 0.0279877
R16330 DVSS.n3486 DVSS.n3485 0.0279877
R16331 DVSS.n3485 DVSS.n2695 0.0279877
R16332 DVSS.n2711 DVSS.n2695 0.0279877
R16333 DVSS.n2712 DVSS.n2711 0.0279877
R16334 DVSS.n3474 DVSS.n3473 0.0279877
R16335 DVSS.n2730 DVSS.n2729 0.0279877
R16336 DVSS.n3462 DVSS.n2730 0.0279877
R16337 DVSS.n3462 DVSS.n3461 0.0279877
R16338 DVSS.n3458 DVSS.n3457 0.0279877
R16339 DVSS.n3457 DVSS.n2733 0.0279877
R16340 DVSS.n2747 DVSS.n2733 0.0279877
R16341 DVSS.n3446 DVSS.n2747 0.0279877
R16342 DVSS.n3446 DVSS.n3445 0.0279877
R16343 DVSS.n2766 DVSS.n2763 0.0279877
R16344 DVSS.n3434 DVSS.n2767 0.0279877
R16345 DVSS.n3434 DVSS.n3433 0.0279877
R16346 DVSS.n3433 DVSS.n2768 0.0279877
R16347 DVSS.n3422 DVSS.n2784 0.0279877
R16348 DVSS.n3422 DVSS.n3421 0.0279877
R16349 DVSS.n3421 DVSS.n2785 0.0279877
R16350 DVSS.n2802 DVSS.n2785 0.0279877
R16351 DVSS.n2803 DVSS.n2802 0.0279877
R16352 DVSS.n3410 DVSS.n3409 0.0279877
R16353 DVSS.n2821 DVSS.n2820 0.0279877
R16354 DVSS.n3398 DVSS.n2821 0.0279877
R16355 DVSS.n3398 DVSS.n3397 0.0279877
R16356 DVSS.n3394 DVSS.n3393 0.0279877
R16357 DVSS.n3393 DVSS.n2825 0.0279877
R16358 DVSS.n2839 DVSS.n2825 0.0279877
R16359 DVSS.n3382 DVSS.n2839 0.0279877
R16360 DVSS.n3382 DVSS.n3381 0.0279877
R16361 DVSS.n2858 DVSS.n2855 0.0279877
R16362 DVSS.n3370 DVSS.n2859 0.0279877
R16363 DVSS.n3370 DVSS.n3369 0.0279877
R16364 DVSS.n3369 DVSS.n2860 0.0279877
R16365 DVSS.n2876 DVSS.n2860 0.0279877
R16366 DVSS.n3358 DVSS.n3357 0.0279877
R16367 DVSS.n3357 DVSS.n2878 0.0279877
R16368 DVSS.n2895 DVSS.n2878 0.0279877
R16369 DVSS.n2896 DVSS.n2895 0.0279877
R16370 DVSS.n3346 DVSS.n2896 0.0279877
R16371 DVSS.n2913 DVSS.n2912 0.0279877
R16372 DVSS.n3333 DVSS.n2913 0.0279877
R16373 DVSS.n3333 DVSS.n3332 0.0279877
R16374 DVSS.n3332 DVSS.n2914 0.0279877
R16375 DVSS.n3007 DVSS.n2930 0.0279877
R16376 DVSS.n3320 DVSS.n2930 0.0279877
R16377 DVSS.n3320 DVSS.n3319 0.0279877
R16378 DVSS.n3319 DVSS.n2931 0.0279877
R16379 DVSS.n2947 DVSS.n2931 0.0279877
R16380 DVSS.n3307 DVSS.n3306 0.0279877
R16381 DVSS.n3306 DVSS.n2949 0.0279877
R16382 DVSS.n2966 DVSS.n2949 0.0279877
R16383 DVSS.n3295 DVSS.n2966 0.0279877
R16384 DVSS.n3293 DVSS.n2967 0.0279877
R16385 DVSS.n2983 DVSS.n2967 0.0279877
R16386 DVSS.n2984 DVSS.n2983 0.0279877
R16387 DVSS.n3282 DVSS.n2984 0.0279877
R16388 DVSS.n3282 DVSS.n3281 0.0279877
R16389 DVSS.n3270 DVSS.n3266 0.0279877
R16390 DVSS.n3270 DVSS.n3269 0.0279877
R16391 DVSS.n3269 DVSS.n1790 0.0279877
R16392 DVSS.n3827 DVSS.n1790 0.0279877
R16393 DVSS.n3505 DVSS.n2666 0.0279877
R16394 DVSS.n3026 DVSS.n2666 0.0279877
R16395 DVSS.n3031 DVSS.n3026 0.0279877
R16396 DVSS.n3032 DVSS.n3031 0.0279877
R16397 DVSS.n3037 DVSS.n3036 0.0279877
R16398 DVSS.n3042 DVSS.n3037 0.0279877
R16399 DVSS.n3043 DVSS.n3042 0.0279877
R16400 DVSS.n3043 DVSS.n3023 0.0279877
R16401 DVSS.n3047 DVSS.n3023 0.0279877
R16402 DVSS.n3054 DVSS.n3049 0.0279877
R16403 DVSS.n3059 DVSS.n3055 0.0279877
R16404 DVSS.n3060 DVSS.n3059 0.0279877
R16405 DVSS.n3062 DVSS.n3060 0.0279877
R16406 DVSS.n3074 DVSS.n3020 0.0279877
R16407 DVSS.n3075 DVSS.n3074 0.0279877
R16408 DVSS.n3079 DVSS.n3075 0.0279877
R16409 DVSS.n3080 DVSS.n3079 0.0279877
R16410 DVSS.n3085 DVSS.n3080 0.0279877
R16411 DVSS.n3089 DVSS.n3088 0.0279877
R16412 DVSS.n3093 DVSS.n3092 0.0279877
R16413 DVSS.n3098 DVSS.n3093 0.0279877
R16414 DVSS.n3099 DVSS.n3098 0.0279877
R16415 DVSS.n3104 DVSS.n3103 0.0279877
R16416 DVSS.n3109 DVSS.n3104 0.0279877
R16417 DVSS.n3110 DVSS.n3109 0.0279877
R16418 DVSS.n3110 DVSS.n3016 0.0279877
R16419 DVSS.n3115 DVSS.n3016 0.0279877
R16420 DVSS.n3122 DVSS.n3117 0.0279877
R16421 DVSS.n3127 DVSS.n3123 0.0279877
R16422 DVSS.n3128 DVSS.n3127 0.0279877
R16423 DVSS.n3131 DVSS.n3128 0.0279877
R16424 DVSS.n3143 DVSS.n3013 0.0279877
R16425 DVSS.n3144 DVSS.n3143 0.0279877
R16426 DVSS.n3148 DVSS.n3144 0.0279877
R16427 DVSS.n3149 DVSS.n3148 0.0279877
R16428 DVSS.n3154 DVSS.n3149 0.0279877
R16429 DVSS.n3158 DVSS.n3157 0.0279877
R16430 DVSS.n3162 DVSS.n3161 0.0279877
R16431 DVSS.n3167 DVSS.n3162 0.0279877
R16432 DVSS.n3168 DVSS.n3167 0.0279877
R16433 DVSS.n3172 DVSS.n3168 0.0279877
R16434 DVSS.n3179 DVSS.n3174 0.0279877
R16435 DVSS.n3180 DVSS.n3179 0.0279877
R16436 DVSS.n3180 DVSS.n3011 0.0279877
R16437 DVSS.n3185 DVSS.n3011 0.0279877
R16438 DVSS.n3186 DVSS.n3185 0.0279877
R16439 DVSS.n3196 DVSS.n3192 0.0279877
R16440 DVSS.n3197 DVSS.n3196 0.0279877
R16441 DVSS.n3197 DVSS.n3009 0.0279877
R16442 DVSS.n3203 DVSS.n3009 0.0279877
R16443 DVSS.n3209 DVSS.n3205 0.0279877
R16444 DVSS.n3210 DVSS.n3209 0.0279877
R16445 DVSS.n3215 DVSS.n3210 0.0279877
R16446 DVSS.n3216 DVSS.n3215 0.0279877
R16447 DVSS.n3220 DVSS.n3216 0.0279877
R16448 DVSS.n3228 DVSS.n3006 0.0279877
R16449 DVSS.n3229 DVSS.n3228 0.0279877
R16450 DVSS.n3233 DVSS.n3229 0.0279877
R16451 DVSS.n3234 DVSS.n3233 0.0279877
R16452 DVSS.n3240 DVSS.n3239 0.0279877
R16453 DVSS.n3240 DVSS.n3004 0.0279877
R16454 DVSS.n3244 DVSS.n3004 0.0279877
R16455 DVSS.n3245 DVSS.n3244 0.0279877
R16456 DVSS.n3250 DVSS.n3245 0.0279877
R16457 DVSS.n3257 DVSS.n3256 0.0279877
R16458 DVSS.n3259 DVSS.n3257 0.0279877
R16459 DVSS.n3259 DVSS.n3258 0.0279877
R16460 DVSS.n3258 DVSS.n1791 0.0279877
R16461 DVSS.n3358 DVSS.n2877 0.0275443
R16462 DVSS.n3174 DVSS.n3173 0.0275443
R16463 DVSS.n3496 DVSS.n2675 0.0275
R16464 DVSS.n3463 DVSS.n2728 0.0275
R16465 DVSS.n3305 DVSS.n2950 0.0275
R16466 DVSS.n3271 DVSS.n3264 0.0275
R16467 DVSS.n3030 DVSS.n3029 0.0275
R16468 DVSS.n3064 DVSS.n3022 0.0275
R16469 DVSS.n3227 DVSS.n3226 0.0275
R16470 DVSS.n3261 DVSS.n3001 0.0275
R16471 DVSS.n2537 DVSS.n2536 0.0274684
R16472 DVSS.n2534 DVSS.n2533 0.0274684
R16473 DVSS.n2265 DVSS.n2256 0.0274684
R16474 DVSS.n2262 DVSS.n1903 0.0274684
R16475 DVSS.n5704 DVSS.n61 0.0272082
R16476 DVSS.n3381 DVSS.n2840 0.027101
R16477 DVSS.n3155 DVSS.n3154 0.027101
R16478 DVSS.n3484 DVSS.n3483 0.027
R16479 DVSS.n3476 DVSS.n3475 0.027
R16480 DVSS.n3292 DVSS.n3291 0.027
R16481 DVSS.n3284 DVSS.n3283 0.027
R16482 DVSS.n3041 DVSS.n2698 0.027
R16483 DVSS.n3050 DVSS.n2706 0.027
R16484 DVSS.n3238 DVSS.n2970 0.027
R16485 DVSS.n3246 DVSS.n2978 0.027
R16486 DVSS.n2233 DVSS.n2231 0.026913
R16487 DVSS.n2235 DVSS.n2233 0.026913
R16488 DVSS.n2237 DVSS.n2235 0.026913
R16489 DVSS.n2239 DVSS.n2237 0.026913
R16490 DVSS.n2240 DVSS.n2239 0.026913
R16491 DVSS.n2243 DVSS.n2240 0.026913
R16492 DVSS.n2245 DVSS.n2243 0.026913
R16493 DVSS.n2246 DVSS.n2245 0.026913
R16494 DVSS.n2247 DVSS.n2246 0.026913
R16495 DVSS.n4152 DVSS.n4141 0.026913
R16496 DVSS.n4152 DVSS.n4151 0.026913
R16497 DVSS.n4151 DVSS.n4149 0.026913
R16498 DVSS.n4149 DVSS.n4146 0.026913
R16499 DVSS.n4146 DVSS.n4145 0.026913
R16500 DVSS.n4145 DVSS.n4143 0.026913
R16501 DVSS.n4143 DVSS.n1525 0.026913
R16502 DVSS.n4158 DVSS.n1525 0.026913
R16503 DVSS.n1538 DVSS.n1537 0.026913
R16504 DVSS.n4148 DVSS.n4147 0.026913
R16505 DVSS.n4157 DVSS.n1526 0.026913
R16506 DVSS.n2018 DVSS.n1970 0.0267204
R16507 DVSS.n2613 DVSS.n1849 0.0267108
R16508 DVSS.n2324 DVSS.n2320 0.0265092
R16509 DVSS.n2574 DVSS.n1887 0.0265092
R16510 DVSS.n3455 DVSS.n2734 0.0265
R16511 DVSS.n2944 DVSS.n2932 0.0265
R16512 DVSS.n3076 DVSS.n2736 0.0265
R16513 DVSS.n3218 DVSS.n3217 0.0265
R16514 DVSS.n3345 DVSS.n3344 0.0262143
R16515 DVSS.n3191 DVSS.n3010 0.0262143
R16516 DVSS.n4872 DVSS.n1196 0.02615
R16517 DVSS.n3432 DVSS.n2762 0.026
R16518 DVSS.n3335 DVSS.n2910 0.026
R16519 DVSS.n3097 DVSS.n3096 0.026
R16520 DVSS.n3195 DVSS.n2907 0.026
R16521 DVSS.n1634 DVSS.n1633 0.0259029
R16522 DVSS.n462 DVSS.n230 0.0257489
R16523 DVSS.n458 DVSS.n230 0.0257489
R16524 DVSS.n458 DVSS.n457 0.0257489
R16525 DVSS.n457 DVSS.n456 0.0257489
R16526 DVSS.n456 DVSS.n232 0.0257489
R16527 DVSS.n452 DVSS.n232 0.0257489
R16528 DVSS.n452 DVSS.n451 0.0257489
R16529 DVSS.n451 DVSS.n450 0.0257489
R16530 DVSS.n450 DVSS.n234 0.0257489
R16531 DVSS.n446 DVSS.n234 0.0257489
R16532 DVSS.n446 DVSS.n445 0.0257489
R16533 DVSS.n445 DVSS.n444 0.0257489
R16534 DVSS.n444 DVSS.n236 0.0257489
R16535 DVSS.n440 DVSS.n236 0.0257489
R16536 DVSS.n440 DVSS.n439 0.0257489
R16537 DVSS.n439 DVSS.n438 0.0257489
R16538 DVSS.n438 DVSS.n238 0.0257489
R16539 DVSS.n434 DVSS.n238 0.0257489
R16540 DVSS.n434 DVSS.n433 0.0257489
R16541 DVSS.n433 DVSS.n432 0.0257489
R16542 DVSS.n432 DVSS.n240 0.0257489
R16543 DVSS.n428 DVSS.n240 0.0257489
R16544 DVSS.n272 DVSS.n271 0.0257489
R16545 DVSS.n278 DVSS.n271 0.0257489
R16546 DVSS.n279 DVSS.n278 0.0257489
R16547 DVSS.n280 DVSS.n279 0.0257489
R16548 DVSS.n280 DVSS.n269 0.0257489
R16549 DVSS.n284 DVSS.n269 0.0257489
R16550 DVSS.n285 DVSS.n284 0.0257489
R16551 DVSS.n286 DVSS.n285 0.0257489
R16552 DVSS.n286 DVSS.n267 0.0257489
R16553 DVSS.n290 DVSS.n267 0.0257489
R16554 DVSS.n291 DVSS.n290 0.0257489
R16555 DVSS.n292 DVSS.n291 0.0257489
R16556 DVSS.n292 DVSS.n265 0.0257489
R16557 DVSS.n296 DVSS.n265 0.0257489
R16558 DVSS.n297 DVSS.n296 0.0257489
R16559 DVSS.n298 DVSS.n297 0.0257489
R16560 DVSS.n298 DVSS.n263 0.0257489
R16561 DVSS.n302 DVSS.n263 0.0257489
R16562 DVSS.n303 DVSS.n302 0.0257489
R16563 DVSS.n304 DVSS.n303 0.0257489
R16564 DVSS.n304 DVSS.n259 0.0257489
R16565 DVSS.n309 DVSS.n261 0.0257489
R16566 DVSS.n2481 DVSS.n2477 0.0256835
R16567 DVSS.n2729 DVSS 0.0255493
R16568 DVSS.n3055 DVSS 0.0255493
R16569 DVSS.n3412 DVSS.n3411 0.0255
R16570 DVSS.n3359 DVSS.n2875 0.0255
R16571 DVSS.n3118 DVSS.n2796 0.0255
R16572 DVSS.n3177 DVSS.n3175 0.0255
R16573 DVSS.n3391 DVSS.n2826 0.025
R16574 DVSS.n3380 DVSS.n3379 0.025
R16575 DVSS.n3145 DVSS.n2828 0.025
R16576 DVSS.n3153 DVSS.n2843 0.025
R16577 DVSS.n5703 DVSS.n5702 0.0249638
R16578 DVSS.n3008 DVSS.n3007 0.0248842
R16579 DVSS.n3205 DVSS.n3204 0.0248842
R16580 DVSS.n4379 DVSS.n4378 0.0248508
R16581 DVSS.n2682 DVSS.n2681 0.0247925
R16582 DVSS.n261 DVSS.n260 0.0247308
R16583 DVSS.n3400 DVSS.n2818 0.0245
R16584 DVSS.n3368 DVSS.n2854 0.0245
R16585 DVSS.n3126 DVSS.n2815 0.0245
R16586 DVSS.n3166 DVSS.n3165 0.0245
R16587 DVSS.n2804 DVSS.n2803 0.0244409
R16588 DVSS.n3116 DVSS.n3115 0.0244409
R16589 DVSS DVSS.n2629 0.0241842
R16590 DVSS.n3423 DVSS.n2783 0.024
R16591 DVSS.n3348 DVSS.n3347 0.024
R16592 DVSS.n3107 DVSS.n3105 0.024
R16593 DVSS.n3187 DVSS.n2889 0.024
R16594 DVSS.n3308 DVSS.n2948 0.0235542
R16595 DVSS.n3222 DVSS.n3221 0.0235542
R16596 DVSS.n3444 DVSS.n3443 0.0235
R16597 DVSS.n2928 DVSS.n2927 0.0235
R16598 DVSS.n3084 DVSS.n2751 0.0235
R16599 DVSS.n3208 DVSS.n3207 0.0235
R16600 DVSS.n3017 DVSS.n2768 0.0231108
R16601 DVSS.n3099 DVSS.n3018 0.0231108
R16602 DVSS.n3495 DVSS.n2676 0.023
R16603 DVSS.n3464 DVSS.n2727 0.023
R16604 DVSS.n3304 DVSS.n2951 0.023
R16605 DVSS.n3272 DVSS.n3000 0.023
R16606 DVSS.n3033 DVSS.n2678 0.023
R16607 DVSS.n3058 DVSS.n2724 0.023
R16608 DVSS.n3230 DVSS.n2953 0.023
R16609 DVSS.n3255 DVSS.n2997 0.023
R16610 DVSS.n2767 DVSS 0.0228892
R16611 DVSS.n3092 DVSS 0.0228892
R16612 DVSS.n1940 DVSS.n1861 0.0227936
R16613 DVSS.n2591 DVSS.n2590 0.0227859
R16614 DVSS.n1889 DVSS.n1872 0.0227859
R16615 DVSS.n1900 DVSS.n1898 0.0227859
R16616 DVSS.n2552 DVSS.n1915 0.0227859
R16617 DVSS.n2336 DVSS.n2335 0.0227859
R16618 DVSS.n1901 DVSS.n1900 0.0227859
R16619 DVSS.n1917 DVSS.n1915 0.0227859
R16620 DVSS.n2333 DVSS.n2328 0.0227859
R16621 DVSS.n1870 DVSS.n1866 0.0227859
R16622 DVSS.n2594 DVSS.n2593 0.0227859
R16623 DVSS.n4150 DVSS.n1535 0.0227554
R16624 DVSS.n4144 DVSS.n1532 0.0227554
R16625 DVSS.n310 DVSS.n309 0.0226946
R16626 DVSS.n250 DVSS.n249 0.0226275
R16627 DVSS.n3487 DVSS.n2693 0.0225
R16628 DVSS.n3472 DVSS.n2709 0.0225
R16629 DVSS.n3296 DVSS.n2965 0.0225
R16630 DVSS.n3280 DVSS.n2981 0.0225
R16631 DVSS.n3040 DVSS.n3038 0.0225
R16632 DVSS.n3053 DVSS.n3052 0.0225
R16633 DVSS.n3237 DVSS.n3235 0.0225
R16634 DVSS.n3249 DVSS.n3248 0.0225
R16635 DVSS.n5100 DVSS.n5099 0.0224253
R16636 DVSS.n5101 DVSS.n5100 0.0224253
R16637 DVSS.n5101 DVSS.n1077 0.0224253
R16638 DVSS.n5107 DVSS.n1077 0.0224253
R16639 DVSS.n5108 DVSS.n5107 0.0224253
R16640 DVSS.n5109 DVSS.n5108 0.0224253
R16641 DVSS.n5109 DVSS.n1073 0.0224253
R16642 DVSS.n5115 DVSS.n1073 0.0224253
R16643 DVSS.n5116 DVSS.n5115 0.0224253
R16644 DVSS.n5117 DVSS.n5116 0.0224253
R16645 DVSS.n5117 DVSS.n1069 0.0224253
R16646 DVSS.n5123 DVSS.n1069 0.0224253
R16647 DVSS.n5124 DVSS.n5123 0.0224253
R16648 DVSS.n5125 DVSS.n5124 0.0224253
R16649 DVSS.n5125 DVSS.n1065 0.0224253
R16650 DVSS.n5131 DVSS.n1065 0.0224253
R16651 DVSS.n5132 DVSS.n5131 0.0224253
R16652 DVSS.n5133 DVSS.n5132 0.0224253
R16653 DVSS.n5133 DVSS.n1061 0.0224253
R16654 DVSS.n5139 DVSS.n1061 0.0224253
R16655 DVSS.n5140 DVSS.n5139 0.0224253
R16656 DVSS.n5141 DVSS.n5140 0.0224253
R16657 DVSS.n5141 DVSS.n1057 0.0224253
R16658 DVSS.n5147 DVSS.n1057 0.0224253
R16659 DVSS.n5148 DVSS.n5147 0.0224253
R16660 DVSS.n5149 DVSS.n5148 0.0224253
R16661 DVSS.n5149 DVSS.n1053 0.0224253
R16662 DVSS.n5155 DVSS.n1053 0.0224253
R16663 DVSS.n5156 DVSS.n5155 0.0224253
R16664 DVSS.n5157 DVSS.n5156 0.0224253
R16665 DVSS.n5157 DVSS.n1049 0.0224253
R16666 DVSS.n5163 DVSS.n1049 0.0224253
R16667 DVSS.n5164 DVSS.n5163 0.0224253
R16668 DVSS.n5165 DVSS.n5164 0.0224253
R16669 DVSS.n5165 DVSS.n1045 0.0224253
R16670 DVSS.n5171 DVSS.n1045 0.0224253
R16671 DVSS.n5172 DVSS.n5171 0.0224253
R16672 DVSS.n5173 DVSS.n5172 0.0224253
R16673 DVSS.n5173 DVSS.n1041 0.0224253
R16674 DVSS.n5179 DVSS.n1041 0.0224253
R16675 DVSS.n5180 DVSS.n5179 0.0224253
R16676 DVSS.n5181 DVSS.n5180 0.0224253
R16677 DVSS.n5181 DVSS.n1037 0.0224253
R16678 DVSS.n5187 DVSS.n1037 0.0224253
R16679 DVSS.n5188 DVSS.n5187 0.0224253
R16680 DVSS.n5189 DVSS.n5188 0.0224253
R16681 DVSS.n5189 DVSS.n1033 0.0224253
R16682 DVSS.n5195 DVSS.n1033 0.0224253
R16683 DVSS.n5196 DVSS.n5195 0.0224253
R16684 DVSS.n5197 DVSS.n5196 0.0224253
R16685 DVSS.n5197 DVSS.n1029 0.0224253
R16686 DVSS.n5203 DVSS.n1029 0.0224253
R16687 DVSS.n5204 DVSS.n5203 0.0224253
R16688 DVSS.n5206 DVSS.n5204 0.0224253
R16689 DVSS.n5206 DVSS.n5205 0.0224253
R16690 DVSS.n5205 DVSS.n1025 0.0224253
R16691 DVSS.n5213 DVSS.n1025 0.0224253
R16692 DVSS.n5220 DVSS.n1020 0.0224253
R16693 DVSS.n5221 DVSS.n5220 0.0224253
R16694 DVSS.n5222 DVSS.n5221 0.0224253
R16695 DVSS.n5222 DVSS.n1016 0.0224253
R16696 DVSS.n5228 DVSS.n1016 0.0224253
R16697 DVSS.n5229 DVSS.n5228 0.0224253
R16698 DVSS.n5230 DVSS.n5229 0.0224253
R16699 DVSS.n5230 DVSS.n1012 0.0224253
R16700 DVSS.n5236 DVSS.n1012 0.0224253
R16701 DVSS.n5237 DVSS.n5236 0.0224253
R16702 DVSS.n5238 DVSS.n5237 0.0224253
R16703 DVSS.n5238 DVSS.n1008 0.0224253
R16704 DVSS.n5244 DVSS.n1008 0.0224253
R16705 DVSS.n5245 DVSS.n5244 0.0224253
R16706 DVSS.n5246 DVSS.n5245 0.0224253
R16707 DVSS.n5246 DVSS.n1004 0.0224253
R16708 DVSS.n5252 DVSS.n1004 0.0224253
R16709 DVSS.n5253 DVSS.n5252 0.0224253
R16710 DVSS.n5254 DVSS.n5253 0.0224253
R16711 DVSS.n5254 DVSS.n1000 0.0224253
R16712 DVSS.n5260 DVSS.n1000 0.0224253
R16713 DVSS.n5261 DVSS.n5260 0.0224253
R16714 DVSS.n5262 DVSS.n5261 0.0224253
R16715 DVSS.n5262 DVSS.n996 0.0224253
R16716 DVSS.n5268 DVSS.n996 0.0224253
R16717 DVSS.n5269 DVSS.n5268 0.0224253
R16718 DVSS.n5270 DVSS.n5269 0.0224253
R16719 DVSS.n5270 DVSS.n992 0.0224253
R16720 DVSS.n5276 DVSS.n992 0.0224253
R16721 DVSS.n5277 DVSS.n5276 0.0224253
R16722 DVSS.n5278 DVSS.n5277 0.0224253
R16723 DVSS.n5278 DVSS.n988 0.0224253
R16724 DVSS.n5284 DVSS.n988 0.0224253
R16725 DVSS.n5285 DVSS.n5284 0.0224253
R16726 DVSS.n5286 DVSS.n5285 0.0224253
R16727 DVSS.n5286 DVSS.n984 0.0224253
R16728 DVSS.n5292 DVSS.n984 0.0224253
R16729 DVSS.n5293 DVSS.n5292 0.0224253
R16730 DVSS.n5294 DVSS.n5293 0.0224253
R16731 DVSS.n5294 DVSS.n980 0.0224253
R16732 DVSS.n5300 DVSS.n980 0.0224253
R16733 DVSS.n5301 DVSS.n5300 0.0224253
R16734 DVSS.n5302 DVSS.n5301 0.0224253
R16735 DVSS.n5302 DVSS.n976 0.0224253
R16736 DVSS.n5308 DVSS.n976 0.0224253
R16737 DVSS.n5309 DVSS.n5308 0.0224253
R16738 DVSS.n5310 DVSS.n5309 0.0224253
R16739 DVSS.n5310 DVSS.n972 0.0224253
R16740 DVSS.n5316 DVSS.n972 0.0224253
R16741 DVSS.n5317 DVSS.n5316 0.0224253
R16742 DVSS.n5318 DVSS.n5317 0.0224253
R16743 DVSS.n5318 DVSS.n968 0.0224253
R16744 DVSS.n5324 DVSS.n968 0.0224253
R16745 DVSS.n5325 DVSS.n5324 0.0224253
R16746 DVSS.n5327 DVSS.n5325 0.0224253
R16747 DVSS.n5327 DVSS.n5326 0.0224253
R16748 DVSS.n5326 DVSS.n964 0.0224253
R16749 DVSS.n5334 DVSS.n964 0.0224253
R16750 DVSS.n2501 DVSS.n2485 0.0223919
R16751 DVSS.n2499 DVSS.n2485 0.0223919
R16752 DVSS.n1936 DVSS.n1863 0.0223919
R16753 DVSS.n2498 DVSS.n2476 0.0223919
R16754 DVSS.n2500 DVSS.n2498 0.0223919
R16755 DVSS.n1941 DVSS.n1940 0.0223807
R16756 DVSS.n1940 DVSS.n1939 0.0223807
R16757 DVSS.n3294 DVSS.n3293 0.0222241
R16758 DVSS.n3239 DVSS.n3005 0.0222241
R16759 DVSS.n2745 DVSS.n2744 0.022
R16760 DVSS.n3318 DVSS.n3317 0.022
R16761 DVSS.n3078 DVSS.n3077 0.022
R16762 DVSS.n3214 DVSS.n2934 0.022
R16763 DVSS.n3445 DVSS.n2748 0.0217808
R16764 DVSS.n3086 DVSS.n3085 0.0217808
R16765 DVSS.n4854 DVSS.n4853 0.0216765
R16766 DVSS.n4827 DVSS.n1221 0.0216765
R16767 DVSS.n4859 DVSS.n1208 0.0216765
R16768 DVSS.n2554 DVSS.n1916 0.021555
R16769 DVSS.n2588 DVSS.n1867 0.021555
R16770 DVSS.n5706 DVSS.n5705 0.0215113
R16771 DVSS.n3431 DVSS.n2769 0.0215
R16772 DVSS.n2909 DVSS.n2897 0.0215
R16773 DVSS.n3100 DVSS.n2771 0.0215
R16774 DVSS.n3194 DVSS.n3193 0.0215
R16775 DVSS.n4154 DVSS.n4153 0.021288
R16776 DVSS.n4142 DVSS.n1531 0.021288
R16777 DVSS.n2498 DVSS.n2497 0.0211757
R16778 DVSS.n1936 DVSS.n1935 0.0211757
R16779 DVSS.n2570 DVSS.n2569 0.0211422
R16780 DVSS.n3408 DVSS.n2799 0.021
R16781 DVSS.n3360 DVSS.n2874 0.021
R16782 DVSS.n3121 DVSS.n3120 0.021
R16783 DVSS.n3171 DVSS.n2871 0.021
R16784 DVSS.n3265 DVSS.n2985 0.0208941
R16785 DVSS.n3252 DVSS.n3251 0.0208941
R16786 DVSS.n2555 DVSS.n2554 0.02075
R16787 DVSS.n2554 DVSS.n2553 0.02075
R16788 DVSS.n2569 DVSS.n1899 0.02075
R16789 DVSS.n2569 DVSS.n2568 0.02075
R16790 DVSS.n3397 DVSS.n2822 0.0206724
R16791 DVSS.n3131 DVSS.n3130 0.0206724
R16792 DVSS.n307 DVSS.n60 0.0206158
R16793 DVSS.n2837 DVSS.n2836 0.0205
R16794 DVSS.n3383 DVSS.n2838 0.0205
R16795 DVSS.n3147 DVSS.n3146 0.0205
R16796 DVSS.n3152 DVSS.n3150 0.0205
R16797 DVSS.n3461 DVSS.n2731 0.0204507
R16798 DVSS.n3062 DVSS.n3061 0.0204507
R16799 DVSS.n2820 DVSS 0.0202291
R16800 DVSS.n3123 DVSS 0.0202291
R16801 DVSS.n5711 DVSS.n5710 0.020197
R16802 DVSS.n2817 DVSS.n2805 0.02
R16803 DVSS.n3367 DVSS.n2861 0.02
R16804 DVSS.n3125 DVSS.n3124 0.02
R16805 DVSS.n3169 DVSS.n2863 0.02
R16806 DVSS.n2484 DVSS.n2477 0.0199037
R16807 DVSS.n2596 DVSS.n1862 0.0199037
R16808 DVSS.n854 DVSS.n852 0.0195912
R16809 DVSS.n854 DVSS.n851 0.0195912
R16810 DVSS.n1368 DVSS.n851 0.0195912
R16811 DVSS.n853 DVSS.n850 0.0195912
R16812 DVSS.n853 DVSS.n849 0.0195912
R16813 DVSS.n849 DVSS.n848 0.0195912
R16814 DVSS.n3424 DVSS.n2782 0.0195
R16815 DVSS.n3343 DVSS.n2892 0.0195
R16816 DVSS.n3102 DVSS.n2779 0.0195
R16817 DVSS.n3190 DVSS.n3189 0.0195
R16818 DVSS.n766 DVSS.n765 0.0191284
R16819 DVSS.n2713 DVSS.n2712 0.0191207
R16820 DVSS.n3048 DVSS.n3047 0.0191207
R16821 DVSS.n2325 DVSS.n2324 0.019078
R16822 DVSS.n2574 DVSS.n2573 0.019078
R16823 DVSS.n3447 DVSS.n2746 0.019
R16824 DVSS.n3322 DVSS.n3321 0.019
R16825 DVSS.n3083 DVSS.n3081 0.019
R16826 DVSS.n3211 DVSS.n2925 0.019
R16827 DVSS DVSS.n3265 0.018899
R16828 DVSS.n3252 DVSS 0.018899
R16829 DVSS.n2692 DVSS.n2691 0.0185
R16830 DVSS.n2726 DVSS.n2714 0.0185
R16831 DVSS.n2964 DVSS.n2963 0.0185
R16832 DVSS.n2999 DVSS.n2986 0.0185
R16833 DVSS.n3035 DVSS.n3034 0.0185
R16834 DVSS.n3057 DVSS.n3056 0.0185
R16835 DVSS.n3232 DVSS.n3231 0.0185
R16836 DVSS.n3254 DVSS.n3253 0.0185
R16837 DVSS.n5535 DVSS.n856 0.018166
R16838 DVSS.n3488 DVSS.n2692 0.018
R16839 DVSS.n3471 DVSS.n2714 0.018
R16840 DVSS.n3297 DVSS.n2964 0.018
R16841 DVSS.n3279 DVSS.n2986 0.018
R16842 DVSS.n3035 DVSS.n2689 0.018
R16843 DVSS.n3056 DVSS.n2716 0.018
R16844 DVSS.n3232 DVSS.n2961 0.018
R16845 DVSS.n3253 DVSS.n2988 0.018
R16846 DVSS.n1867 DVSS.n1862 0.0178394
R16847 DVSS.n3024 DVSS.n2674 0.0177906
R16848 DVSS.n3032 DVSS.n3025 0.0177906
R16849 DVSS.n4654 DVSS.n4653 0.0176
R16850 DVSS.n4370 DVSS.n4359 0.0176
R16851 DVSS.n2859 DVSS 0.017569
R16852 DVSS.n3161 DVSS 0.017569
R16853 DVSS.n3448 DVSS.n3447 0.0175
R16854 DVSS.n3321 DVSS.n2929 0.0175
R16855 DVSS.n3081 DVSS.n2742 0.0175
R16856 DVSS.n3213 DVSS.n3211 0.0175
R16857 DVSS.n2513 DVSS.n2332 0.0174266
R16858 DVSS.n428 DVSS.n427 0.0174005
R16859 DVSS.n4369 DVSS.n4361 0.0172066
R16860 DVSS.n3770 DVSS.n3769 0.0171667
R16861 DVSS.n3771 DVSS.n3770 0.0171667
R16862 DVSS.n5215 DVSS.n5214 0.0171667
R16863 DVSS.n5216 DVSS.n5215 0.0171667
R16864 DVSS.n1946 DVSS.n1945 0.0170138
R16865 DVSS.n2782 DVSS.n2781 0.017
R16866 DVSS.n3343 DVSS.n3342 0.017
R16867 DVSS.n3102 DVSS.n3101 0.017
R16868 DVSS.n3190 DVSS.n2899 0.017
R16869 DVSS.n4661 DVSS.n4638 0.0169185
R16870 DVSS.n4666 DVSS.n4638 0.0169185
R16871 DVSS.n4660 DVSS.n4637 0.0169185
R16872 DVSS.n4665 DVSS.n4637 0.0169185
R16873 DVSS.n4659 DVSS.n4636 0.0169185
R16874 DVSS.n4664 DVSS.n4636 0.0169185
R16875 DVSS.n4658 DVSS.n4635 0.0169185
R16876 DVSS.n4705 DVSS.n4635 0.0169185
R16877 DVSS.n4661 DVSS.n4654 0.0169185
R16878 DVSS.n4666 DVSS.n4655 0.0169185
R16879 DVSS.n4660 DVSS.n4655 0.0169185
R16880 DVSS.n4665 DVSS.n4656 0.0169185
R16881 DVSS.n4659 DVSS.n4656 0.0169185
R16882 DVSS.n4664 DVSS.n4657 0.0169185
R16883 DVSS.n4658 DVSS.n4657 0.0169185
R16884 DVSS.n4706 DVSS.n4705 0.0169185
R16885 DVSS.n4356 DVSS.n4355 0.0169185
R16886 DVSS.n4354 DVSS.n4353 0.0169185
R16887 DVSS.n4352 DVSS.n4351 0.0169185
R16888 DVSS.n4350 DVSS.n4349 0.0169185
R16889 DVSS.n4348 DVSS.n4347 0.0169185
R16890 DVSS.n4346 DVSS.n4345 0.0169185
R16891 DVSS.n4373 DVSS.n4344 0.0169185
R16892 DVSS.n4375 DVSS.n4374 0.0169185
R16893 DVSS.n4359 DVSS.n4356 0.0169185
R16894 DVSS.n4355 DVSS.n4354 0.0169185
R16895 DVSS.n4353 DVSS.n4352 0.0169185
R16896 DVSS.n4351 DVSS.n4350 0.0169185
R16897 DVSS.n4349 DVSS.n4348 0.0169185
R16898 DVSS.n4347 DVSS.n4346 0.0169185
R16899 DVSS.n4345 DVSS.n4344 0.0169185
R16900 DVSS.n4374 DVSS.n4373 0.0169185
R16901 DVSS.n3992 DVSS.n1663 0.0169185
R16902 DVSS.n3991 DVSS.n3989 0.0169185
R16903 DVSS.n3990 DVSS.n1664 0.0169185
R16904 DVSS.n3988 DVSS.n3986 0.0169185
R16905 DVSS.n3987 DVSS.n1665 0.0169185
R16906 DVSS.n3985 DVSS.n3983 0.0169185
R16907 DVSS.n3984 DVSS.n1666 0.0169185
R16908 DVSS.n1668 DVSS.n1667 0.0169185
R16909 DVSS.n2277 DVSS.n1669 0.0169185
R16910 DVSS.n1669 DVSS.n1668 0.0169185
R16911 DVSS.n1667 DVSS.n1666 0.0169185
R16912 DVSS.n3985 DVSS.n3984 0.0169185
R16913 DVSS.n3983 DVSS.n1665 0.0169185
R16914 DVSS.n3988 DVSS.n3987 0.0169185
R16915 DVSS.n3986 DVSS.n1664 0.0169185
R16916 DVSS.n3991 DVSS.n3990 0.0169185
R16917 DVSS.n3989 DVSS.n1663 0.0169185
R16918 DVSS.n3993 DVSS.n3992 0.0169185
R16919 DVSS.n3753 DVSS.n3750 0.0169185
R16920 DVSS.n3750 DVSS.n3529 0.0169185
R16921 DVSS.n3754 DVSS.n3751 0.0169185
R16922 DVSS.n3751 DVSS.n3530 0.0169185
R16923 DVSS.n3755 DVSS.n3752 0.0169185
R16924 DVSS.n3752 DVSS.n3531 0.0169185
R16925 DVSS.n3758 DVSS.n3757 0.0169185
R16926 DVSS.n3758 DVSS.n3532 0.0169185
R16927 DVSS.n3760 DVSS.n3533 0.0169185
R16928 DVSS.n4873 DVSS.n1197 0.0169185
R16929 DVSS.n4884 DVSS.n1201 0.0169185
R16930 DVSS.n1200 DVSS.n1198 0.0169185
R16931 DVSS.n4883 DVSS.n4882 0.0169185
R16932 DVSS.n4882 DVSS.n4875 0.0169185
R16933 DVSS.n4881 DVSS.n4879 0.0169185
R16934 DVSS.n4879 DVSS.n4876 0.0169185
R16935 DVSS.n4887 DVSS.n4886 0.0169185
R16936 DVSS.n4874 DVSS.n4873 0.0169185
R16937 DVSS.n4884 DVSS.n1197 0.0169185
R16938 DVSS.n1201 DVSS.n1200 0.0169185
R16939 DVSS.n4883 DVSS.n1198 0.0169185
R16940 DVSS.n4880 DVSS.n4875 0.0169185
R16941 DVSS.n4881 DVSS.n4880 0.0169185
R16942 DVSS.n4877 DVSS.n4876 0.0169185
R16943 DVSS.n4886 DVSS.n4877 0.0169185
R16944 DVSS.n3753 DVSS.n3528 0.0169185
R16945 DVSS.n3538 DVSS.n3529 0.0169185
R16946 DVSS.n3754 DVSS.n3538 0.0169185
R16947 DVSS.n3537 DVSS.n3530 0.0169185
R16948 DVSS.n3755 DVSS.n3537 0.0169185
R16949 DVSS.n3536 DVSS.n3531 0.0169185
R16950 DVSS.n3757 DVSS.n3536 0.0169185
R16951 DVSS.n3535 DVSS.n3532 0.0169185
R16952 DVSS.n3535 DVSS.n3533 0.0169185
R16953 DVSS.n2493 DVSS.n2492 0.0167162
R16954 DVSS.n5708 DVSS.n5707 0.0166994
R16955 DVSS.n5709 DVSS.n5708 0.0166994
R16956 DVSS.n3407 DVSS.n2805 0.0165
R16957 DVSS.n2873 DVSS.n2861 0.0165
R16958 DVSS.n3124 DVSS.n2807 0.0165
R16959 DVSS.n3170 DVSS.n3169 0.0165
R16960 DVSS.n3308 DVSS 0.0162389
R16961 DVSS.n3222 DVSS 0.0162389
R16962 DVSS.n3384 DVSS.n2837 0.016
R16963 DVSS.n3384 DVSS.n3383 0.016
R16964 DVSS.n3147 DVSS.n2834 0.016
R16965 DVSS.n3150 DVSS.n2834 0.016
R16966 DVSS.n3408 DVSS.n3407 0.0155
R16967 DVSS.n2874 DVSS.n2873 0.0155
R16968 DVSS.n3121 DVSS.n2807 0.0155
R16969 DVSS.n3171 DVSS.n3170 0.0155
R16970 DVSS.n3853 DVSS.n3852 0.0154891
R16971 DVSS.n4653 DVSS.n4639 0.01535
R16972 DVSS.n4371 DVSS.n4370 0.01535
R16973 DVSS.n2366 DVSS.n2363 0.0152819
R16974 DVSS.n2366 DVSS.n2365 0.0152819
R16975 DVSS.n2361 DVSS.n1927 0.0152819
R16976 DVSS.n2363 DVSS.n2352 0.0152819
R16977 DVSS.n2365 DVSS.n2351 0.0152819
R16978 DVSS.n2361 DVSS.n2351 0.0152819
R16979 DVSS.n2299 DVSS.n2297 0.0152819
R16980 DVSS.n2299 DVSS.n2298 0.0152819
R16981 DVSS.n2301 DVSS.n2268 0.0152819
R16982 DVSS.n2297 DVSS.n1875 0.0152819
R16983 DVSS.n2298 DVSS.n2270 0.0152819
R16984 DVSS.n2270 DVSS.n2268 0.0152819
R16985 DVSS.n276 DVSS.n275 0.0152727
R16986 DVSS.n2781 DVSS.n2769 0.015
R16987 DVSS.n3342 DVSS.n2897 0.015
R16988 DVSS.n3101 DVSS.n3100 0.015
R16989 DVSS.n3193 DVSS.n2899 0.015
R16990 DVSS.n2597 DVSS.n1861 0.0149495
R16991 DVSS.n2912 DVSS 0.0149089
R16992 DVSS.n3192 DVSS 0.0149089
R16993 DVSS.n4651 DVSS.n4650 0.0149069
R16994 DVSS.n4645 DVSS.n4644 0.0149069
R16995 DVSS.n4648 DVSS.n4644 0.0149069
R16996 DVSS.n4648 DVSS.n4647 0.0149069
R16997 DVSS.n4650 DVSS.n4642 0.0149069
R16998 DVSS.n4645 DVSS.n4642 0.0149069
R16999 DVSS.n4364 DVSS.n4363 0.0149069
R17000 DVSS.n4366 DVSS.n4362 0.0149069
R17001 DVSS.n4365 DVSS.n4357 0.0149069
R17002 DVSS.n4366 DVSS.n4365 0.0149069
R17003 DVSS.n4364 DVSS.n4362 0.0149069
R17004 DVSS.n4368 DVSS.n4363 0.0149069
R17005 DVSS.n1391 DVSS.n1390 0.0145462
R17006 DVSS.n1390 DVSS.n1387 0.0145462
R17007 DVSS.n1387 DVSS.n1386 0.0145462
R17008 DVSS.n1386 DVSS.n1384 0.0145462
R17009 DVSS.n1384 DVSS.n1382 0.0145462
R17010 DVSS.n1382 DVSS.n1379 0.0145462
R17011 DVSS.n1379 DVSS.n1378 0.0145462
R17012 DVSS.n1378 DVSS.n1376 0.0145462
R17013 DVSS.n1376 DVSS.n1374 0.0145462
R17014 DVSS.n1374 DVSS.n1367 0.0145462
R17015 DVSS.n4766 DVSS.n1367 0.0145462
R17016 DVSS.n1950 DVSS.n1932 0.0145367
R17017 DVSS.n3448 DVSS.n2745 0.0145
R17018 DVSS.n3318 DVSS.n2929 0.0145
R17019 DVSS.n3078 DVSS.n2742 0.0145
R17020 DVSS.n3214 DVSS.n3213 0.0145
R17021 DVSS.n4153 DVSS.n1533 0.0144402
R17022 DVSS.n4142 DVSS.n1536 0.0144402
R17023 DVSS.n954 DVSS.n953 0.0144028
R17024 DVSS.n2410 DVSS.n2409 0.0142903
R17025 DVSS.n1763 DVSS.n1762 0.0142903
R17026 DVSS.n2488 DVSS.n1923 0.0142838
R17027 DVSS.n2092 DVSS.n2091 0.0142814
R17028 DVSS.n1953 DVSS.n1951 0.0141679
R17029 DVSS.n1956 DVSS.n1539 0.0141679
R17030 DVSS.n1956 DVSS.n1951 0.0141679
R17031 DVSS.n2252 DVSS.n1953 0.0141679
R17032 DVSS.n3488 DVSS.n3487 0.014
R17033 DVSS.n3472 DVSS.n3471 0.014
R17034 DVSS.n3297 DVSS.n3296 0.014
R17035 DVSS.n3280 DVSS.n3279 0.014
R17036 DVSS.n3038 DVSS.n2689 0.014
R17037 DVSS.n3053 DVSS.n2716 0.014
R17038 DVSS.n3235 DVSS.n2961 0.014
R17039 DVSS.n3249 DVSS.n2988 0.014
R17040 DVSS.n1389 DVSS.n1388 0.0136707
R17041 DVSS.n1381 DVSS.n1380 0.0136707
R17042 DVSS.n1373 DVSS.n1372 0.0136707
R17043 DVSS.n3344 DVSS 0.0135788
R17044 DVSS DVSS.n3191 0.0135788
R17045 DVSS.n4647 DVSS.n4639 0.01355
R17046 DVSS.n4371 DVSS.n4357 0.01355
R17047 DVSS.n2012 DVSS.n1977 0.0135392
R17048 DVSS.n2691 DVSS.n2676 0.0135
R17049 DVSS.n2727 DVSS.n2726 0.0135
R17050 DVSS.n2963 DVSS.n2951 0.0135
R17051 DVSS.n3000 DVSS.n2999 0.0135
R17052 DVSS.n3034 DVSS.n3033 0.0135
R17053 DVSS.n3058 DVSS.n3057 0.0135
R17054 DVSS.n3231 DVSS.n3230 0.0135
R17055 DVSS.n3255 DVSS.n3254 0.0135
R17056 DVSS.n2307 DVSS.n1931 0.0134255
R17057 DVSS.n2305 DVSS.n1931 0.0134255
R17058 DVSS.n2544 DVSS.n1922 0.0134255
R17059 DVSS.n2546 DVSS.n1922 0.0134255
R17060 DVSS.n2232 DVSS.n1958 0.0133402
R17061 DVSS.n2242 DVSS.n2241 0.0133402
R17062 DVSS.n3444 DVSS.n2746 0.013
R17063 DVSS.n3322 DVSS.n2928 0.013
R17064 DVSS.n3084 DVSS.n3083 0.013
R17065 DVSS.n3208 DVSS.n2925 0.013
R17066 DVSS.n2234 DVSS.n2227 0.0129835
R17067 DVSS.n2238 DVSS.n1962 0.0129835
R17068 DVSS.n4150 DVSS.n1533 0.0129728
R17069 DVSS.n4144 DVSS.n1536 0.0129728
R17070 DVSS.n798 DVSS.n754 0.0129415
R17071 DVSS.n798 DVSS.n797 0.0129415
R17072 DVSS.n797 DVSS.n796 0.0129415
R17073 DVSS.n796 DVSS.n756 0.0129415
R17074 DVSS.n792 DVSS.n756 0.0129415
R17075 DVSS.n792 DVSS.n791 0.0129415
R17076 DVSS.n791 DVSS.n790 0.0129415
R17077 DVSS.n790 DVSS.n758 0.0129415
R17078 DVSS.n786 DVSS.n758 0.0129415
R17079 DVSS.n786 DVSS.n785 0.0129415
R17080 DVSS.n785 DVSS.n784 0.0129415
R17081 DVSS.n784 DVSS.n760 0.0129415
R17082 DVSS.n780 DVSS.n760 0.0129415
R17083 DVSS.n780 DVSS.n779 0.0129415
R17084 DVSS.n779 DVSS.n778 0.0129415
R17085 DVSS.n778 DVSS.n762 0.0129415
R17086 DVSS.n774 DVSS.n762 0.0129415
R17087 DVSS.n774 DVSS.n773 0.0129415
R17088 DVSS.n773 DVSS.n772 0.0129415
R17089 DVSS.n772 DVSS.n764 0.0129415
R17090 DVSS.n768 DVSS.n764 0.0129415
R17091 DVSS.n768 DVSS.n767 0.0129415
R17092 DVSS.n5713 DVSS.n5712 0.0129415
R17093 DVSS.n74 DVSS.n58 0.0129415
R17094 DVSS.n75 DVSS.n74 0.0129415
R17095 DVSS.n76 DVSS.n75 0.0129415
R17096 DVSS.n76 DVSS.n70 0.0129415
R17097 DVSS.n80 DVSS.n70 0.0129415
R17098 DVSS.n81 DVSS.n80 0.0129415
R17099 DVSS.n82 DVSS.n81 0.0129415
R17100 DVSS.n82 DVSS.n68 0.0129415
R17101 DVSS.n86 DVSS.n68 0.0129415
R17102 DVSS.n87 DVSS.n86 0.0129415
R17103 DVSS.n88 DVSS.n87 0.0129415
R17104 DVSS.n88 DVSS.n66 0.0129415
R17105 DVSS.n92 DVSS.n66 0.0129415
R17106 DVSS.n93 DVSS.n92 0.0129415
R17107 DVSS.n94 DVSS.n93 0.0129415
R17108 DVSS.n94 DVSS.n64 0.0129415
R17109 DVSS.n98 DVSS.n64 0.0129415
R17110 DVSS.n99 DVSS.n98 0.0129415
R17111 DVSS.n100 DVSS.n99 0.0129415
R17112 DVSS.n100 DVSS.n62 0.0129415
R17113 DVSS.n5705 DVSS.n62 0.0129415
R17114 DVSS.n253 DVSS.n248 0.0127612
R17115 DVSS.n254 DVSS.n251 0.0127612
R17116 DVSS.n1867 DVSS.n1864 0.01265
R17117 DVSS.n1867 DVSS.n1865 0.01265
R17118 DVSS.n3424 DVSS.n3423 0.0125
R17119 DVSS.n3347 DVSS.n2892 0.0125
R17120 DVSS.n3105 DVSS.n2779 0.0125
R17121 DVSS.n3189 DVSS.n3187 0.0125
R17122 DVSS.n2523 DVSS.n2522 0.0124725
R17123 DVSS.n1895 DVSS.n1894 0.0124725
R17124 DVSS.n461 DVSS.n460 0.0123471
R17125 DVSS.n460 DVSS.n459 0.0123471
R17126 DVSS.n459 DVSS.n231 0.0123471
R17127 DVSS.n455 DVSS.n231 0.0123471
R17128 DVSS.n455 DVSS.n454 0.0123471
R17129 DVSS.n454 DVSS.n453 0.0123471
R17130 DVSS.n453 DVSS.n233 0.0123471
R17131 DVSS.n449 DVSS.n233 0.0123471
R17132 DVSS.n449 DVSS.n448 0.0123471
R17133 DVSS.n448 DVSS.n447 0.0123471
R17134 DVSS.n447 DVSS.n235 0.0123471
R17135 DVSS.n443 DVSS.n235 0.0123471
R17136 DVSS.n443 DVSS.n442 0.0123471
R17137 DVSS.n442 DVSS.n441 0.0123471
R17138 DVSS.n441 DVSS.n237 0.0123471
R17139 DVSS.n437 DVSS.n237 0.0123471
R17140 DVSS.n437 DVSS.n436 0.0123471
R17141 DVSS.n436 DVSS.n435 0.0123471
R17142 DVSS.n435 DVSS.n239 0.0123471
R17143 DVSS.n431 DVSS.n239 0.0123471
R17144 DVSS.n431 DVSS.n430 0.0123471
R17145 DVSS.n430 DVSS.n429 0.0123471
R17146 DVSS.n274 DVSS.n273 0.0123471
R17147 DVSS.n277 DVSS.n270 0.0123471
R17148 DVSS.n281 DVSS.n270 0.0123471
R17149 DVSS.n282 DVSS.n281 0.0123471
R17150 DVSS.n283 DVSS.n282 0.0123471
R17151 DVSS.n283 DVSS.n268 0.0123471
R17152 DVSS.n287 DVSS.n268 0.0123471
R17153 DVSS.n288 DVSS.n287 0.0123471
R17154 DVSS.n289 DVSS.n288 0.0123471
R17155 DVSS.n289 DVSS.n266 0.0123471
R17156 DVSS.n293 DVSS.n266 0.0123471
R17157 DVSS.n294 DVSS.n293 0.0123471
R17158 DVSS.n295 DVSS.n294 0.0123471
R17159 DVSS.n295 DVSS.n264 0.0123471
R17160 DVSS.n299 DVSS.n264 0.0123471
R17161 DVSS.n300 DVSS.n299 0.0123471
R17162 DVSS.n301 DVSS.n300 0.0123471
R17163 DVSS.n301 DVSS.n262 0.0123471
R17164 DVSS.n305 DVSS.n262 0.0123471
R17165 DVSS.n306 DVSS.n305 0.0123471
R17166 DVSS.n308 DVSS.n306 0.0123471
R17167 DVSS.n308 DVSS.n307 0.0123471
R17168 DVSS.n1365 DVSS.n1356 0.0123293
R17169 DVSS.n4767 DVSS.n1362 0.0123293
R17170 DVSS.n1954 DVSS.n1952 0.0122701
R17171 DVSS.n2248 DVSS.n2230 0.0122701
R17172 DVSS DVSS.n3307 0.0122488
R17173 DVSS DVSS.n3006 0.0122488
R17174 DVSS.n2818 DVSS.n2817 0.012
R17175 DVSS.n3368 DVSS.n3367 0.012
R17176 DVSS.n3126 DVSS.n3125 0.012
R17177 DVSS.n3166 DVSS.n2863 0.012
R17178 DVSS.n2480 DVSS.n2479 0.0116468
R17179 DVSS.n5214 DVSS.n1020 0.0116395
R17180 DVSS.n1843 DVSS.n1842 0.0116
R17181 DVSS.n1383 DVSS.n1366 0.0115976
R17182 DVSS.n1377 DVSS.n1361 0.0115976
R17183 DVSS.n2836 DVSS.n2826 0.0115
R17184 DVSS.n3380 DVSS.n2838 0.0115
R17185 DVSS.n3146 DVSS.n3145 0.0115
R17186 DVSS.n3153 DVSS.n3152 0.0115
R17187 DVSS.n2517 DVSS.n2330 0.0113969
R17188 DVSS.n2517 DVSS.n2331 0.0113969
R17189 DVSS.n2587 DVSS.n1869 0.0113969
R17190 DVSS.n2587 DVSS.n2586 0.0113969
R17191 DVSS.n5214 DVSS.n5213 0.0112859
R17192 DVSS.n4730 DVSS.n4609 0.0112561
R17193 DVSS.n4719 DVSS.n4620 0.0112561
R17194 DVSS.n4588 DVSS.n1406 0.0112561
R17195 DVSS.n4600 DVSS.n1398 0.0112561
R17196 DVSS.n4548 DVSS.n4547 0.0112561
R17197 DVSS.n4565 DVSS.n1417 0.0112561
R17198 DVSS.n4450 DVSS.n4447 0.0112561
R17199 DVSS.n4525 DVSS.n1438 0.0112561
R17200 DVSS.n4482 DVSS.n4416 0.0112561
R17201 DVSS.n4471 DVSS.n4427 0.0112561
R17202 DVSS.n4395 DVSS.n4335 0.0112561
R17203 DVSS.n4407 DVSS.n4327 0.0112561
R17204 DVSS.n4842 VSS 0.0110882
R17205 DVSS.n4836 VSS 0.0110882
R17206 DVSS.n4863 VSS 0.0110882
R17207 DVSS.n3411 DVSS.n2799 0.011
R17208 DVSS.n3360 DVSS.n3359 0.011
R17209 DVSS.n3120 DVSS.n3118 0.011
R17210 DVSS.n3175 DVSS.n2871 0.011
R17211 DVSS.n4123 DVSS.n4122 0.0109694
R17212 DVSS.n4124 DVSS.n4123 0.0109694
R17213 DVSS.n4124 DVSS.n1543 0.0109694
R17214 DVSS.n4130 DVSS.n1543 0.0109694
R17215 DVSS.n4131 DVSS.n4130 0.0109694
R17216 DVSS.n4132 DVSS.n4131 0.0109694
R17217 DVSS.n4132 DVSS.n1521 0.0109694
R17218 DVSS.n4167 DVSS.n1521 0.0109694
R17219 DVSS.n4167 DVSS.n4166 0.0109694
R17220 DVSS DVSS.n2858 0.0109187
R17221 DVSS.n3158 DVSS 0.0109187
R17222 DVSS.n3806 DVSS.n1843 0.0109
R17223 DVSS.n3807 DVSS.n3806 0.0109
R17224 DVSS.n3808 DVSS.n3807 0.0109
R17225 DVSS.n3809 DVSS.n3808 0.0109
R17226 DVSS.n3810 DVSS.n3809 0.0109
R17227 DVSS.n3811 DVSS.n3810 0.0109
R17228 DVSS.n3812 DVSS.n3811 0.0109
R17229 DVSS.n3813 DVSS.n3812 0.0109
R17230 DVSS.n3814 DVSS.n3813 0.0109
R17231 DVSS.n3815 DVSS.n3814 0.0109
R17232 DVSS.n3816 DVSS.n3815 0.0109
R17233 DVSS.n1385 DVSS.n1364 0.0108659
R17234 DVSS.n1375 DVSS.n1359 0.0108659
R17235 DVSS.n3024 DVSS.n2694 0.010697
R17236 DVSS.n3036 DVSS.n3025 0.010697
R17237 DVSS.n2683 DVSS.n2682 0.0105
R17238 DVSS.n2683 DVSS.n2680 0.0105
R17239 DVSS.n3492 DVSS.n2680 0.0105
R17240 DVSS.n3492 DVSS.n3491 0.0105
R17241 DVSS.n3491 DVSS.n2688 0.0105
R17242 DVSS.n2700 DVSS.n2688 0.0105
R17243 DVSS.n3480 DVSS.n2700 0.0105
R17244 DVSS.n3480 DVSS.n3479 0.0105
R17245 DVSS.n3479 DVSS.n2705 0.0105
R17246 DVSS.n2718 DVSS.n2705 0.0105
R17247 DVSS.n3468 DVSS.n2718 0.0105
R17248 DVSS.n3468 DVSS.n3467 0.0105
R17249 DVSS.n3467 DVSS.n2723 0.0105
R17250 DVSS.n3069 DVSS.n2723 0.0105
R17251 DVSS.n3069 DVSS.n2738 0.0105
R17252 DVSS.n3452 DVSS.n2738 0.0105
R17253 DVSS.n3452 DVSS.n3451 0.0105
R17254 DVSS.n3451 DVSS.n2741 0.0105
R17255 DVSS.n2753 DVSS.n2741 0.0105
R17256 DVSS.n3440 DVSS.n2753 0.0105
R17257 DVSS.n3440 DVSS.n3439 0.0105
R17258 DVSS.n3439 DVSS.n2758 0.0105
R17259 DVSS.n2773 DVSS.n2758 0.0105
R17260 DVSS.n3428 DVSS.n2773 0.0105
R17261 DVSS.n3428 DVSS.n3427 0.0105
R17262 DVSS.n3427 DVSS.n2778 0.0105
R17263 DVSS.n2790 DVSS.n2778 0.0105
R17264 DVSS.n3416 DVSS.n2790 0.0105
R17265 DVSS.n3416 DVSS.n3415 0.0105
R17266 DVSS.n3415 DVSS.n2795 0.0105
R17267 DVSS.n2809 DVSS.n2795 0.0105
R17268 DVSS.n3404 DVSS.n2809 0.0105
R17269 DVSS.n3404 DVSS.n3403 0.0105
R17270 DVSS.n3403 DVSS.n2814 0.0105
R17271 DVSS.n3138 DVSS.n2814 0.0105
R17272 DVSS.n3138 DVSS.n2830 0.0105
R17273 DVSS.n3388 DVSS.n2830 0.0105
R17274 DVSS.n3388 DVSS.n3387 0.0105
R17275 DVSS.n3387 DVSS.n2833 0.0105
R17276 DVSS.n2845 DVSS.n2833 0.0105
R17277 DVSS.n3376 DVSS.n2845 0.0105
R17278 DVSS.n3376 DVSS.n3375 0.0105
R17279 DVSS.n3375 DVSS.n2850 0.0105
R17280 DVSS.n2865 DVSS.n2850 0.0105
R17281 DVSS.n3364 DVSS.n2865 0.0105
R17282 DVSS.n3364 DVSS.n3363 0.0105
R17283 DVSS.n3363 DVSS.n2870 0.0105
R17284 DVSS.n2883 DVSS.n2870 0.0105
R17285 DVSS.n3352 DVSS.n2883 0.0105
R17286 DVSS.n3352 DVSS.n3351 0.0105
R17287 DVSS.n3351 DVSS.n2888 0.0105
R17288 DVSS.n2901 DVSS.n2888 0.0105
R17289 DVSS.n3339 DVSS.n2901 0.0105
R17290 DVSS.n3339 DVSS.n3338 0.0105
R17291 DVSS.n3338 DVSS.n2906 0.0105
R17292 DVSS.n2919 DVSS.n2906 0.0105
R17293 DVSS.n3326 DVSS.n2919 0.0105
R17294 DVSS.n3326 DVSS.n3325 0.0105
R17295 DVSS.n3325 DVSS.n2924 0.0105
R17296 DVSS.n2936 DVSS.n2924 0.0105
R17297 DVSS.n3314 DVSS.n2936 0.0105
R17298 DVSS.n3314 DVSS.n3313 0.0105
R17299 DVSS.n3313 DVSS.n2941 0.0105
R17300 DVSS.n2955 DVSS.n2941 0.0105
R17301 DVSS.n3301 DVSS.n2955 0.0105
R17302 DVSS.n3301 DVSS.n3300 0.0105
R17303 DVSS.n3300 DVSS.n2960 0.0105
R17304 DVSS.n2972 DVSS.n2960 0.0105
R17305 DVSS.n3288 DVSS.n2972 0.0105
R17306 DVSS.n3288 DVSS.n3287 0.0105
R17307 DVSS.n3287 DVSS.n2977 0.0105
R17308 DVSS.n2990 DVSS.n2977 0.0105
R17309 DVSS.n3276 DVSS.n2990 0.0105
R17310 DVSS.n3276 DVSS.n3275 0.0105
R17311 DVSS.n3275 DVSS.n2996 0.0105
R17312 DVSS.n2996 DVSS.n1786 0.0105
R17313 DVSS.n3831 DVSS.n1786 0.0105
R17314 DVSS.n3831 DVSS.n1784 0.0105
R17315 DVSS.n3835 DVSS.n1784 0.0105
R17316 DVSS.n3835 DVSS.n1782 0.0105
R17317 DVSS.n3839 DVSS.n1782 0.0105
R17318 DVSS.n3839 DVSS.n1780 0.0105
R17319 DVSS.n3863 DVSS.n1780 0.0105
R17320 DVSS.n3863 DVSS.n3862 0.0105
R17321 DVSS.n3862 DVSS.n3861 0.0105
R17322 DVSS.n3861 DVSS.n3845 0.0105
R17323 DVSS.n3857 DVSS.n3845 0.0105
R17324 DVSS.n3857 DVSS.n3856 0.0105
R17325 DVSS.n3856 DVSS.n3855 0.0105
R17326 DVSS.n3432 DVSS.n3431 0.0105
R17327 DVSS.n2910 DVSS.n2909 0.0105
R17328 DVSS.n3097 DVSS.n2771 0.0105
R17329 DVSS.n3195 DVSS.n3194 0.0105
R17330 DVSS.n3836 DVSS.n1783 0.0105
R17331 DVSS.n3837 DVSS.n3836 0.0105
R17332 DVSS.n3838 DVSS.n3837 0.0105
R17333 DVSS.n3838 DVSS.n1778 0.0105
R17334 DVSS.n3864 DVSS.n1779 0.0105
R17335 DVSS.n3860 DVSS.n1779 0.0105
R17336 DVSS.n3860 DVSS.n3859 0.0105
R17337 DVSS.n3859 DVSS.n3858 0.0105
R17338 DVSS.n3858 DVSS.n3846 0.0105
R17339 DVSS.n3854 DVSS.n3846 0.0105
R17340 DVSS.n3865 DVSS.n3864 0.0104296
R17341 DVSS.n5546 DVSS.n826 0.0103531
R17342 DVSS.n5798 DVSS.n3 0.0103531
R17343 DVSS.n5792 DVSS.n27 0.0103531
R17344 DVSS.n4731 DVSS.n4730 0.0101185
R17345 DVSS.n4717 DVSS.n4620 0.0101185
R17346 DVSS.n4586 DVSS.n1406 0.0101185
R17347 DVSS.n4601 DVSS.n4600 0.0101185
R17348 DVSS.n4547 DVSS.n1428 0.0101185
R17349 DVSS.n4567 DVSS.n1417 0.0101185
R17350 DVSS.n4451 DVSS.n4450 0.0101185
R17351 DVSS.n4527 DVSS.n1438 0.0101185
R17352 DVSS.n4483 DVSS.n4482 0.0101185
R17353 DVSS.n4469 DVSS.n4427 0.0101185
R17354 DVSS.n4393 DVSS.n4335 0.0101185
R17355 DVSS.n4408 DVSS.n4407 0.0101185
R17356 DVSS.n5538 DVSS.n848 0.0100456
R17357 DVSS.n1369 DVSS.n1368 0.0100456
R17358 DVSS.n4768 DVSS.n852 0.0100456
R17359 DVSS.n1369 DVSS.n850 0.0100456
R17360 DVSS.n2744 DVSS.n2734 0.01
R17361 DVSS.n3317 DVSS.n2932 0.01
R17362 DVSS.n3077 DVSS.n3076 0.01
R17363 DVSS.n3217 DVSS.n2934 0.01
R17364 DVSS.n3797 DVSS 0.00997368
R17365 DVSS.n2251 DVSS.n2250 0.00965456
R17366 DVSS.n2244 DVSS.n2229 0.00965456
R17367 DVSS.n953 DVSS.n950 0.00962857
R17368 DVSS.n5348 DVSS.n950 0.00962857
R17369 DVSS.n5348 DVSS.n948 0.00962857
R17370 DVSS.n5352 DVSS.n948 0.00962857
R17371 DVSS.n5352 DVSS.n946 0.00962857
R17372 DVSS.n5356 DVSS.n946 0.00962857
R17373 DVSS.n5356 DVSS.n944 0.00962857
R17374 DVSS.n5360 DVSS.n944 0.00962857
R17375 DVSS.n5360 DVSS.n942 0.00962857
R17376 DVSS.n5364 DVSS.n942 0.00962857
R17377 DVSS.n5364 DVSS.n940 0.00962857
R17378 DVSS.n5368 DVSS.n940 0.00962857
R17379 DVSS.n5368 DVSS.n938 0.00962857
R17380 DVSS.n5372 DVSS.n938 0.00962857
R17381 DVSS.n5372 DVSS.n936 0.00962857
R17382 DVSS.n5376 DVSS.n936 0.00962857
R17383 DVSS.n5376 DVSS.n934 0.00962857
R17384 DVSS.n5380 DVSS.n934 0.00962857
R17385 DVSS.n5380 DVSS.n932 0.00962857
R17386 DVSS.n5384 DVSS.n932 0.00962857
R17387 DVSS.n5384 DVSS.n930 0.00962857
R17388 DVSS.n5388 DVSS.n930 0.00962857
R17389 DVSS.n5388 DVSS.n928 0.00962857
R17390 DVSS.n5392 DVSS.n928 0.00962857
R17391 DVSS.n5392 DVSS.n926 0.00962857
R17392 DVSS.n5396 DVSS.n926 0.00962857
R17393 DVSS.n5396 DVSS.n924 0.00962857
R17394 DVSS.n5400 DVSS.n924 0.00962857
R17395 DVSS.n5400 DVSS.n922 0.00962857
R17396 DVSS.n5404 DVSS.n922 0.00962857
R17397 DVSS.n5404 DVSS.n920 0.00962857
R17398 DVSS.n5408 DVSS.n920 0.00962857
R17399 DVSS.n5408 DVSS.n918 0.00962857
R17400 DVSS.n5412 DVSS.n918 0.00962857
R17401 DVSS.n5412 DVSS.n916 0.00962857
R17402 DVSS.n5416 DVSS.n916 0.00962857
R17403 DVSS.n5416 DVSS.n914 0.00962857
R17404 DVSS.n5420 DVSS.n914 0.00962857
R17405 DVSS.n5420 DVSS.n912 0.00962857
R17406 DVSS.n5424 DVSS.n912 0.00962857
R17407 DVSS.n5424 DVSS.n910 0.00962857
R17408 DVSS.n5428 DVSS.n910 0.00962857
R17409 DVSS.n5428 DVSS.n908 0.00962857
R17410 DVSS.n5432 DVSS.n908 0.00962857
R17411 DVSS.n5432 DVSS.n906 0.00962857
R17412 DVSS.n5436 DVSS.n906 0.00962857
R17413 DVSS.n5436 DVSS.n904 0.00962857
R17414 DVSS.n5440 DVSS.n904 0.00962857
R17415 DVSS.n5440 DVSS.n902 0.00962857
R17416 DVSS.n5444 DVSS.n902 0.00962857
R17417 DVSS.n5444 DVSS.n900 0.00962857
R17418 DVSS.n5448 DVSS.n900 0.00962857
R17419 DVSS.n5448 DVSS.n898 0.00962857
R17420 DVSS.n5452 DVSS.n898 0.00962857
R17421 DVSS.n5452 DVSS.n896 0.00962857
R17422 DVSS.n5456 DVSS.n896 0.00962857
R17423 DVSS.n5456 DVSS.n894 0.00962857
R17424 DVSS.n5460 DVSS.n894 0.00962857
R17425 DVSS.n5460 DVSS.n892 0.00962857
R17426 DVSS.n5464 DVSS.n892 0.00962857
R17427 DVSS.n5464 DVSS.n890 0.00962857
R17428 DVSS.n5468 DVSS.n890 0.00962857
R17429 DVSS.n5468 DVSS.n888 0.00962857
R17430 DVSS.n5472 DVSS.n888 0.00962857
R17431 DVSS.n5472 DVSS.n886 0.00962857
R17432 DVSS.n5476 DVSS.n886 0.00962857
R17433 DVSS.n5476 DVSS.n884 0.00962857
R17434 DVSS.n5480 DVSS.n884 0.00962857
R17435 DVSS.n5480 DVSS.n882 0.00962857
R17436 DVSS.n5484 DVSS.n882 0.00962857
R17437 DVSS.n5484 DVSS.n880 0.00962857
R17438 DVSS.n5488 DVSS.n880 0.00962857
R17439 DVSS.n5488 DVSS.n878 0.00962857
R17440 DVSS.n5492 DVSS.n878 0.00962857
R17441 DVSS.n5492 DVSS.n876 0.00962857
R17442 DVSS.n5496 DVSS.n876 0.00962857
R17443 DVSS.n5496 DVSS.n874 0.00962857
R17444 DVSS.n5500 DVSS.n874 0.00962857
R17445 DVSS.n5500 DVSS.n872 0.00962857
R17446 DVSS.n5504 DVSS.n872 0.00962857
R17447 DVSS.n5504 DVSS.n870 0.00962857
R17448 DVSS.n5508 DVSS.n870 0.00962857
R17449 DVSS.n5508 DVSS.n868 0.00962857
R17450 DVSS.n5512 DVSS.n868 0.00962857
R17451 DVSS.n5512 DVSS.n866 0.00962857
R17452 DVSS.n5516 DVSS.n866 0.00962857
R17453 DVSS.n5516 DVSS.n864 0.00962857
R17454 DVSS.n5520 DVSS.n864 0.00962857
R17455 DVSS.n5520 DVSS.n862 0.00962857
R17456 DVSS.n5524 DVSS.n862 0.00962857
R17457 DVSS.n5524 DVSS.n860 0.00962857
R17458 DVSS.n5528 DVSS.n860 0.00962857
R17459 DVSS.n5528 DVSS.n858 0.00962857
R17460 DVSS.n5532 DVSS.n858 0.00962857
R17461 DVSS.n5347 DVSS.n5346 0.00962857
R17462 DVSS.n5347 DVSS.n947 0.00962857
R17463 DVSS.n5353 DVSS.n947 0.00962857
R17464 DVSS.n5354 DVSS.n5353 0.00962857
R17465 DVSS.n5355 DVSS.n5354 0.00962857
R17466 DVSS.n5355 DVSS.n943 0.00962857
R17467 DVSS.n5361 DVSS.n943 0.00962857
R17468 DVSS.n5362 DVSS.n5361 0.00962857
R17469 DVSS.n5363 DVSS.n5362 0.00962857
R17470 DVSS.n5363 DVSS.n939 0.00962857
R17471 DVSS.n5369 DVSS.n939 0.00962857
R17472 DVSS.n5370 DVSS.n5369 0.00962857
R17473 DVSS.n5371 DVSS.n5370 0.00962857
R17474 DVSS.n5371 DVSS.n935 0.00962857
R17475 DVSS.n5377 DVSS.n935 0.00962857
R17476 DVSS.n5378 DVSS.n5377 0.00962857
R17477 DVSS.n5379 DVSS.n5378 0.00962857
R17478 DVSS.n5379 DVSS.n931 0.00962857
R17479 DVSS.n5385 DVSS.n931 0.00962857
R17480 DVSS.n5386 DVSS.n5385 0.00962857
R17481 DVSS.n5387 DVSS.n5386 0.00962857
R17482 DVSS.n5387 DVSS.n927 0.00962857
R17483 DVSS.n5393 DVSS.n927 0.00962857
R17484 DVSS.n5394 DVSS.n5393 0.00962857
R17485 DVSS.n5395 DVSS.n5394 0.00962857
R17486 DVSS.n5395 DVSS.n923 0.00962857
R17487 DVSS.n5401 DVSS.n923 0.00962857
R17488 DVSS.n5402 DVSS.n5401 0.00962857
R17489 DVSS.n5403 DVSS.n5402 0.00962857
R17490 DVSS.n5403 DVSS.n919 0.00962857
R17491 DVSS.n5409 DVSS.n919 0.00962857
R17492 DVSS.n5410 DVSS.n5409 0.00962857
R17493 DVSS.n5411 DVSS.n5410 0.00962857
R17494 DVSS.n5411 DVSS.n915 0.00962857
R17495 DVSS.n5417 DVSS.n915 0.00962857
R17496 DVSS.n5418 DVSS.n5417 0.00962857
R17497 DVSS.n5419 DVSS.n5418 0.00962857
R17498 DVSS.n5419 DVSS.n911 0.00962857
R17499 DVSS.n5425 DVSS.n911 0.00962857
R17500 DVSS.n5426 DVSS.n5425 0.00962857
R17501 DVSS.n5427 DVSS.n5426 0.00962857
R17502 DVSS.n5427 DVSS.n907 0.00962857
R17503 DVSS.n5433 DVSS.n907 0.00962857
R17504 DVSS.n5434 DVSS.n5433 0.00962857
R17505 DVSS.n5435 DVSS.n5434 0.00962857
R17506 DVSS.n5435 DVSS.n903 0.00962857
R17507 DVSS.n5441 DVSS.n903 0.00962857
R17508 DVSS.n5442 DVSS.n5441 0.00962857
R17509 DVSS.n5443 DVSS.n5442 0.00962857
R17510 DVSS.n5443 DVSS.n899 0.00962857
R17511 DVSS.n5449 DVSS.n899 0.00962857
R17512 DVSS.n5450 DVSS.n5449 0.00962857
R17513 DVSS.n5451 DVSS.n5450 0.00962857
R17514 DVSS.n5451 DVSS.n895 0.00962857
R17515 DVSS.n5457 DVSS.n895 0.00962857
R17516 DVSS.n5458 DVSS.n5457 0.00962857
R17517 DVSS.n5459 DVSS.n5458 0.00962857
R17518 DVSS.n5459 DVSS.n891 0.00962857
R17519 DVSS.n5465 DVSS.n891 0.00962857
R17520 DVSS.n5466 DVSS.n5465 0.00962857
R17521 DVSS.n5467 DVSS.n5466 0.00962857
R17522 DVSS.n5467 DVSS.n887 0.00962857
R17523 DVSS.n5473 DVSS.n887 0.00962857
R17524 DVSS.n5474 DVSS.n5473 0.00962857
R17525 DVSS.n5475 DVSS.n5474 0.00962857
R17526 DVSS.n5475 DVSS.n883 0.00962857
R17527 DVSS.n5481 DVSS.n883 0.00962857
R17528 DVSS.n5482 DVSS.n5481 0.00962857
R17529 DVSS.n5483 DVSS.n5482 0.00962857
R17530 DVSS.n5483 DVSS.n879 0.00962857
R17531 DVSS.n5489 DVSS.n879 0.00962857
R17532 DVSS.n5490 DVSS.n5489 0.00962857
R17533 DVSS.n5491 DVSS.n5490 0.00962857
R17534 DVSS.n5491 DVSS.n875 0.00962857
R17535 DVSS.n5497 DVSS.n875 0.00962857
R17536 DVSS.n5498 DVSS.n5497 0.00962857
R17537 DVSS.n5499 DVSS.n5498 0.00962857
R17538 DVSS.n5499 DVSS.n871 0.00962857
R17539 DVSS.n5505 DVSS.n871 0.00962857
R17540 DVSS.n5506 DVSS.n5505 0.00962857
R17541 DVSS.n5507 DVSS.n5506 0.00962857
R17542 DVSS.n5507 DVSS.n867 0.00962857
R17543 DVSS.n5513 DVSS.n867 0.00962857
R17544 DVSS.n5514 DVSS.n5513 0.00962857
R17545 DVSS.n5515 DVSS.n5514 0.00962857
R17546 DVSS.n5515 DVSS.n863 0.00962857
R17547 DVSS.n5521 DVSS.n863 0.00962857
R17548 DVSS.n5522 DVSS.n5521 0.00962857
R17549 DVSS.n5523 DVSS.n5522 0.00962857
R17550 DVSS.n5523 DVSS.n859 0.00962857
R17551 DVSS.n5529 DVSS.n859 0.00962857
R17552 DVSS.n5530 DVSS.n5529 0.00962857
R17553 DVSS.n5531 DVSS.n5530 0.00962857
R17554 DVSS.n4378 DVSS.n4342 0.00962857
R17555 DVSS.n4382 DVSS.n4342 0.00962857
R17556 DVSS.n4382 DVSS.n4340 0.00962857
R17557 DVSS.n4386 DVSS.n4340 0.00962857
R17558 DVSS.n4386 DVSS.n4338 0.00962857
R17559 DVSS.n4390 DVSS.n4338 0.00962857
R17560 DVSS.n4390 DVSS.n4333 0.00962857
R17561 DVSS.n4401 DVSS.n4333 0.00962857
R17562 DVSS.n4401 DVSS.n4330 0.00962857
R17563 DVSS.n4499 DVSS.n4330 0.00962857
R17564 DVSS.n4499 DVSS.n4331 0.00962857
R17565 DVSS.n4495 DVSS.n4331 0.00962857
R17566 DVSS.n4495 DVSS.n4405 0.00962857
R17567 DVSS.n4491 DVSS.n4405 0.00962857
R17568 DVSS.n4491 DVSS.n4411 0.00962857
R17569 DVSS.n4487 DVSS.n4411 0.00962857
R17570 DVSS.n4487 DVSS.n4413 0.00962857
R17571 DVSS.n4418 DVSS.n4413 0.00962857
R17572 DVSS.n4479 DVSS.n4418 0.00962857
R17573 DVSS.n4479 DVSS.n4419 0.00962857
R17574 DVSS.n4475 DVSS.n4419 0.00962857
R17575 DVSS.n4475 DVSS.n4422 0.00962857
R17576 DVSS.n4437 DVSS.n4422 0.00962857
R17577 DVSS.n4466 DVSS.n4437 0.00962857
R17578 DVSS.n4466 DVSS.n4438 0.00962857
R17579 DVSS.n4462 DVSS.n4438 0.00962857
R17580 DVSS.n4462 DVSS.n4441 0.00962857
R17581 DVSS.n4458 DVSS.n4441 0.00962857
R17582 DVSS.n4458 DVSS.n4443 0.00962857
R17583 DVSS.n4454 DVSS.n4443 0.00962857
R17584 DVSS.n4454 DVSS.n4445 0.00962857
R17585 DVSS.n4445 DVSS.n1445 0.00962857
R17586 DVSS.n4517 DVSS.n1445 0.00962857
R17587 DVSS.n4517 DVSS.n1443 0.00962857
R17588 DVSS.n4521 DVSS.n1443 0.00962857
R17589 DVSS.n4521 DVSS.n1436 0.00962857
R17590 DVSS.n4530 DVSS.n1436 0.00962857
R17591 DVSS.n4530 DVSS.n1434 0.00962857
R17592 DVSS.n4534 DVSS.n1434 0.00962857
R17593 DVSS.n4534 DVSS.n1432 0.00962857
R17594 DVSS.n4539 DVSS.n1432 0.00962857
R17595 DVSS.n4539 DVSS.n1430 0.00962857
R17596 DVSS.n4543 DVSS.n1430 0.00962857
R17597 DVSS.n4543 DVSS.n1425 0.00962857
R17598 DVSS.n4556 DVSS.n1425 0.00962857
R17599 DVSS.n4556 DVSS.n1422 0.00962857
R17600 DVSS.n4561 DVSS.n1422 0.00962857
R17601 DVSS.n4561 DVSS.n1423 0.00962857
R17602 DVSS.n1423 DVSS.n1415 0.00962857
R17603 DVSS.n4571 DVSS.n1415 0.00962857
R17604 DVSS.n4571 DVSS.n1413 0.00962857
R17605 DVSS.n4575 DVSS.n1413 0.00962857
R17606 DVSS.n4575 DVSS.n1411 0.00962857
R17607 DVSS.n4579 DVSS.n1411 0.00962857
R17608 DVSS.n4579 DVSS.n1409 0.00962857
R17609 DVSS.n4583 DVSS.n1409 0.00962857
R17610 DVSS.n4583 DVSS.n1404 0.00962857
R17611 DVSS.n4594 DVSS.n1404 0.00962857
R17612 DVSS.n4594 DVSS.n1401 0.00962857
R17613 DVSS.n4747 DVSS.n1401 0.00962857
R17614 DVSS.n4747 DVSS.n1402 0.00962857
R17615 DVSS.n4743 DVSS.n1402 0.00962857
R17616 DVSS.n4743 DVSS.n4598 0.00962857
R17617 DVSS.n4739 DVSS.n4598 0.00962857
R17618 DVSS.n4739 DVSS.n4604 0.00962857
R17619 DVSS.n4735 DVSS.n4604 0.00962857
R17620 DVSS.n4735 DVSS.n4606 0.00962857
R17621 DVSS.n4611 DVSS.n4606 0.00962857
R17622 DVSS.n4727 DVSS.n4611 0.00962857
R17623 DVSS.n4727 DVSS.n4612 0.00962857
R17624 DVSS.n4723 DVSS.n4612 0.00962857
R17625 DVSS.n4723 DVSS.n4615 0.00962857
R17626 DVSS.n4630 DVSS.n4615 0.00962857
R17627 DVSS.n4714 DVSS.n4630 0.00962857
R17628 DVSS.n4714 DVSS.n4631 0.00962857
R17629 DVSS.n4710 DVSS.n4631 0.00962857
R17630 DVSS.n4710 DVSS.n4634 0.00962857
R17631 DVSS.n4670 DVSS.n4634 0.00962857
R17632 DVSS.n4670 DVSS.n4668 0.00962857
R17633 DVSS.n4702 DVSS.n4668 0.00962857
R17634 DVSS.n4702 DVSS.n4669 0.00962857
R17635 DVSS.n4698 DVSS.n4669 0.00962857
R17636 DVSS.n4698 DVSS.n4674 0.00962857
R17637 DVSS.n4694 DVSS.n4674 0.00962857
R17638 DVSS.n4694 DVSS.n4676 0.00962857
R17639 DVSS.n4690 DVSS.n4676 0.00962857
R17640 DVSS.n4689 DVSS.n4677 0.00962857
R17641 DVSS.n4684 DVSS.n4677 0.00962857
R17642 DVSS.n4684 DVSS.n4680 0.00962857
R17643 DVSS.n4384 DVSS.n4383 0.00962857
R17644 DVSS.n4385 DVSS.n4384 0.00962857
R17645 DVSS.n4385 DVSS.n4336 0.00962857
R17646 DVSS.n4494 DVSS.n4493 0.00962857
R17647 DVSS.n4493 DVSS.n4492 0.00962857
R17648 DVSS.n4492 DVSS.n4410 0.00962857
R17649 DVSS.n4486 DVSS.n4410 0.00962857
R17650 DVSS.n4486 DVSS.n4485 0.00962857
R17651 DVSS.n4467 DVSS.n4436 0.00962857
R17652 DVSS.n4461 DVSS.n4436 0.00962857
R17653 DVSS.n4461 DVSS.n4460 0.00962857
R17654 DVSS.n4460 DVSS.n4459 0.00962857
R17655 DVSS.n4459 DVSS.n4442 0.00962857
R17656 DVSS.n4453 DVSS.n4442 0.00962857
R17657 DVSS.n4529 DVSS.n1433 0.00962857
R17658 DVSS.n4535 DVSS.n1433 0.00962857
R17659 DVSS.n4536 DVSS.n4535 0.00962857
R17660 DVSS.n4538 DVSS.n4536 0.00962857
R17661 DVSS.n4538 DVSS.n4537 0.00962857
R17662 DVSS.n4570 DVSS.n4569 0.00962857
R17663 DVSS.n4570 DVSS.n1412 0.00962857
R17664 DVSS.n4576 DVSS.n1412 0.00962857
R17665 DVSS.n4577 DVSS.n4576 0.00962857
R17666 DVSS.n4578 DVSS.n4577 0.00962857
R17667 DVSS.n4578 DVSS.n1407 0.00962857
R17668 DVSS.n4742 DVSS.n4741 0.00962857
R17669 DVSS.n4741 DVSS.n4740 0.00962857
R17670 DVSS.n4740 DVSS.n4603 0.00962857
R17671 DVSS.n4734 DVSS.n4603 0.00962857
R17672 DVSS.n4734 DVSS.n4733 0.00962857
R17673 DVSS.n4715 DVSS.n4629 0.00962857
R17674 DVSS.n4709 DVSS.n4629 0.00962857
R17675 DVSS.n4709 DVSS.n4708 0.00962857
R17676 DVSS.n4703 DVSS.n4667 0.00962857
R17677 DVSS.n4697 DVSS.n4667 0.00962857
R17678 DVSS.n4697 DVSS.n4696 0.00962857
R17679 DVSS.n4696 DVSS.n4695 0.00962857
R17680 DVSS.n4695 DVSS.n4675 0.00962857
R17681 DVSS.n4675 DVSS.n1358 0.00962857
R17682 DVSS.n4683 DVSS.n4681 0.00962857
R17683 DVSS.n4683 DVSS.n4682 0.00962857
R17684 DVSS.n1573 DVSS.n1570 0.00962857
R17685 DVSS.n1577 DVSS.n1570 0.00962857
R17686 DVSS.n1577 DVSS.n1568 0.00962857
R17687 DVSS.n1581 DVSS.n1568 0.00962857
R17688 DVSS.n1581 DVSS.n1566 0.00962857
R17689 DVSS.n1585 DVSS.n1566 0.00962857
R17690 DVSS.n1585 DVSS.n1564 0.00962857
R17691 DVSS.n1589 DVSS.n1564 0.00962857
R17692 DVSS.n1589 DVSS.n1562 0.00962857
R17693 DVSS.n1593 DVSS.n1562 0.00962857
R17694 DVSS.n1593 DVSS.n1559 0.00962857
R17695 DVSS.n4089 DVSS.n1559 0.00962857
R17696 DVSS.n4089 DVSS.n1560 0.00962857
R17697 DVSS.n4085 DVSS.n1560 0.00962857
R17698 DVSS.n4085 DVSS.n1597 0.00962857
R17699 DVSS.n4081 DVSS.n1597 0.00962857
R17700 DVSS.n4081 DVSS.n1599 0.00962857
R17701 DVSS.n4077 DVSS.n1599 0.00962857
R17702 DVSS.n4077 DVSS.n1601 0.00962857
R17703 DVSS.n4073 DVSS.n1601 0.00962857
R17704 DVSS.n4073 DVSS.n1603 0.00962857
R17705 DVSS.n4069 DVSS.n1603 0.00962857
R17706 DVSS.n4069 DVSS.n1605 0.00962857
R17707 DVSS.n4065 DVSS.n1605 0.00962857
R17708 DVSS.n4065 DVSS.n1607 0.00962857
R17709 DVSS.n4061 DVSS.n1607 0.00962857
R17710 DVSS.n4061 DVSS.n1609 0.00962857
R17711 DVSS.n3607 DVSS.n1609 0.00962857
R17712 DVSS.n3610 DVSS.n3607 0.00962857
R17713 DVSS.n3610 DVSS.n3605 0.00962857
R17714 DVSS.n3614 DVSS.n3605 0.00962857
R17715 DVSS.n3614 DVSS.n3603 0.00962857
R17716 DVSS.n3618 DVSS.n3603 0.00962857
R17717 DVSS.n3618 DVSS.n3601 0.00962857
R17718 DVSS.n3622 DVSS.n3601 0.00962857
R17719 DVSS.n3622 DVSS.n3599 0.00962857
R17720 DVSS.n3626 DVSS.n3599 0.00962857
R17721 DVSS.n3626 DVSS.n3597 0.00962857
R17722 DVSS.n3630 DVSS.n3597 0.00962857
R17723 DVSS.n3630 DVSS.n3595 0.00962857
R17724 DVSS.n3634 DVSS.n3595 0.00962857
R17725 DVSS.n3634 DVSS.n3593 0.00962857
R17726 DVSS.n3638 DVSS.n3593 0.00962857
R17727 DVSS.n3638 DVSS.n3591 0.00962857
R17728 DVSS.n3642 DVSS.n3591 0.00962857
R17729 DVSS.n3642 DVSS.n3589 0.00962857
R17730 DVSS.n3646 DVSS.n3589 0.00962857
R17731 DVSS.n3646 DVSS.n3587 0.00962857
R17732 DVSS.n3650 DVSS.n3587 0.00962857
R17733 DVSS.n3650 DVSS.n3585 0.00962857
R17734 DVSS.n3654 DVSS.n3585 0.00962857
R17735 DVSS.n3654 DVSS.n3583 0.00962857
R17736 DVSS.n3658 DVSS.n3583 0.00962857
R17737 DVSS.n3658 DVSS.n3581 0.00962857
R17738 DVSS.n3662 DVSS.n3581 0.00962857
R17739 DVSS.n3662 DVSS.n3579 0.00962857
R17740 DVSS.n3666 DVSS.n3579 0.00962857
R17741 DVSS.n3666 DVSS.n3577 0.00962857
R17742 DVSS.n3670 DVSS.n3577 0.00962857
R17743 DVSS.n3670 DVSS.n3575 0.00962857
R17744 DVSS.n3674 DVSS.n3575 0.00962857
R17745 DVSS.n3674 DVSS.n3573 0.00962857
R17746 DVSS.n3678 DVSS.n3573 0.00962857
R17747 DVSS.n3678 DVSS.n3571 0.00962857
R17748 DVSS.n3682 DVSS.n3571 0.00962857
R17749 DVSS.n3682 DVSS.n3569 0.00962857
R17750 DVSS.n3686 DVSS.n3569 0.00962857
R17751 DVSS.n3686 DVSS.n3567 0.00962857
R17752 DVSS.n3690 DVSS.n3567 0.00962857
R17753 DVSS.n3690 DVSS.n3565 0.00962857
R17754 DVSS.n3694 DVSS.n3565 0.00962857
R17755 DVSS.n3694 DVSS.n3563 0.00962857
R17756 DVSS.n3698 DVSS.n3563 0.00962857
R17757 DVSS.n3698 DVSS.n3561 0.00962857
R17758 DVSS.n3702 DVSS.n3561 0.00962857
R17759 DVSS.n3702 DVSS.n3559 0.00962857
R17760 DVSS.n3706 DVSS.n3559 0.00962857
R17761 DVSS.n3706 DVSS.n3557 0.00962857
R17762 DVSS.n3710 DVSS.n3557 0.00962857
R17763 DVSS.n3710 DVSS.n3555 0.00962857
R17764 DVSS.n3714 DVSS.n3555 0.00962857
R17765 DVSS.n3714 DVSS.n3553 0.00962857
R17766 DVSS.n3718 DVSS.n3553 0.00962857
R17767 DVSS.n3718 DVSS.n3551 0.00962857
R17768 DVSS.n3722 DVSS.n3551 0.00962857
R17769 DVSS.n3722 DVSS.n3549 0.00962857
R17770 DVSS.n3726 DVSS.n3549 0.00962857
R17771 DVSS.n3726 DVSS.n3547 0.00962857
R17772 DVSS.n3730 DVSS.n3547 0.00962857
R17773 DVSS.n3730 DVSS.n3545 0.00962857
R17774 DVSS.n3734 DVSS.n3545 0.00962857
R17775 DVSS.n3734 DVSS.n3543 0.00962857
R17776 DVSS.n3738 DVSS.n3543 0.00962857
R17777 DVSS.n3738 DVSS.n3541 0.00962857
R17778 DVSS.n3742 DVSS.n3541 0.00962857
R17779 DVSS.n3742 DVSS.n3539 0.00962857
R17780 DVSS.n3748 DVSS.n3539 0.00962857
R17781 DVSS.n3745 DVSS.n3526 0.00962857
R17782 DVSS.n3764 DVSS.n3526 0.00962857
R17783 DVSS.n3764 DVSS.n3524 0.00962857
R17784 DVSS.n2613 DVSS.n2612 0.00962857
R17785 DVSS.n2612 DVSS.n1851 0.00962857
R17786 DVSS.n2608 DVSS.n1851 0.00962857
R17787 DVSS.n2608 DVSS.n1853 0.00962857
R17788 DVSS.n2604 DVSS.n1853 0.00962857
R17789 DVSS.n2604 DVSS.n1856 0.00962857
R17790 DVSS.n2600 DVSS.n1856 0.00962857
R17791 DVSS.n2600 DVSS.n1858 0.00962857
R17792 DVSS.n2281 DVSS.n1858 0.00962857
R17793 DVSS.n2284 DVSS.n2281 0.00962857
R17794 DVSS.n2284 DVSS.n2274 0.00962857
R17795 DVSS.n2290 DVSS.n2274 0.00962857
R17796 DVSS.n2290 DVSS.n2272 0.00962857
R17797 DVSS.n2294 DVSS.n2272 0.00962857
R17798 DVSS.n2294 DVSS.n1879 0.00962857
R17799 DVSS.n2581 DVSS.n1879 0.00962857
R17800 DVSS.n2581 DVSS.n1880 0.00962857
R17801 DVSS.n2577 DVSS.n1880 0.00962857
R17802 DVSS.n2577 DVSS.n1883 0.00962857
R17803 DVSS.n2259 DVSS.n1883 0.00962857
R17804 DVSS.n2259 DVSS.n1906 0.00962857
R17805 DVSS.n2563 DVSS.n1906 0.00962857
R17806 DVSS.n2563 DVSS.n1907 0.00962857
R17807 DVSS.n2559 DVSS.n1907 0.00962857
R17808 DVSS.n2559 DVSS.n1910 0.00962857
R17809 DVSS.n2530 DVSS.n1910 0.00962857
R17810 DVSS.n2530 DVSS.n2314 0.00962857
R17811 DVSS.n2526 DVSS.n2314 0.00962857
R17812 DVSS.n2526 DVSS.n2316 0.00962857
R17813 DVSS.n2355 DVSS.n2316 0.00962857
R17814 DVSS.n2355 DVSS.n2354 0.00962857
R17815 DVSS.n2359 DVSS.n2354 0.00962857
R17816 DVSS.n2359 DVSS.n2344 0.00962857
R17817 DVSS.n2373 DVSS.n2344 0.00962857
R17818 DVSS.n2373 DVSS.n2341 0.00962857
R17819 DVSS.n2509 DVSS.n2341 0.00962857
R17820 DVSS.n2509 DVSS.n2342 0.00962857
R17821 DVSS.n2505 DVSS.n2342 0.00962857
R17822 DVSS.n2505 DVSS.n2470 0.00962857
R17823 DVSS.n2470 DVSS.n2469 0.00962857
R17824 DVSS.n2469 DVSS.n2377 0.00962857
R17825 DVSS.n2465 DVSS.n2377 0.00962857
R17826 DVSS.n2465 DVSS.n2380 0.00962857
R17827 DVSS.n2461 DVSS.n2380 0.00962857
R17828 DVSS.n2461 DVSS.n2383 0.00962857
R17829 DVSS.n2457 DVSS.n2383 0.00962857
R17830 DVSS.n2457 DVSS.n2385 0.00962857
R17831 DVSS.n2453 DVSS.n2385 0.00962857
R17832 DVSS.n2453 DVSS.n2387 0.00962857
R17833 DVSS.n2449 DVSS.n2387 0.00962857
R17834 DVSS.n2449 DVSS.n2389 0.00962857
R17835 DVSS.n2445 DVSS.n2389 0.00962857
R17836 DVSS.n2445 DVSS.n2391 0.00962857
R17837 DVSS.n2441 DVSS.n2391 0.00962857
R17838 DVSS.n2441 DVSS.n2393 0.00962857
R17839 DVSS.n2437 DVSS.n2393 0.00962857
R17840 DVSS.n2437 DVSS.n2395 0.00962857
R17841 DVSS.n2433 DVSS.n2395 0.00962857
R17842 DVSS.n2433 DVSS.n2397 0.00962857
R17843 DVSS.n2429 DVSS.n2397 0.00962857
R17844 DVSS.n2429 DVSS.n2399 0.00962857
R17845 DVSS.n2425 DVSS.n2399 0.00962857
R17846 DVSS.n2425 DVSS.n2401 0.00962857
R17847 DVSS.n2421 DVSS.n2401 0.00962857
R17848 DVSS.n2421 DVSS.n2403 0.00962857
R17849 DVSS.n2417 DVSS.n2403 0.00962857
R17850 DVSS.n2417 DVSS.n2405 0.00962857
R17851 DVSS.n2413 DVSS.n2405 0.00962857
R17852 DVSS.n2413 DVSS.n2407 0.00962857
R17853 DVSS.n2020 DVSS.n1970 0.00962857
R17854 DVSS.n2020 DVSS.n1968 0.00962857
R17855 DVSS.n2024 DVSS.n1968 0.00962857
R17856 DVSS.n2024 DVSS.n1964 0.00962857
R17857 DVSS.n2225 DVSS.n1964 0.00962857
R17858 DVSS.n2225 DVSS.n1966 0.00962857
R17859 DVSS.n2221 DVSS.n1966 0.00962857
R17860 DVSS.n2221 DVSS.n2028 0.00962857
R17861 DVSS.n2217 DVSS.n2028 0.00962857
R17862 DVSS.n2217 DVSS.n2030 0.00962857
R17863 DVSS.n2213 DVSS.n2030 0.00962857
R17864 DVSS.n2213 DVSS.n2032 0.00962857
R17865 DVSS.n2209 DVSS.n2032 0.00962857
R17866 DVSS.n2209 DVSS.n2034 0.00962857
R17867 DVSS.n2205 DVSS.n2034 0.00962857
R17868 DVSS.n2205 DVSS.n2036 0.00962857
R17869 DVSS.n2201 DVSS.n2036 0.00962857
R17870 DVSS.n2201 DVSS.n2038 0.00962857
R17871 DVSS.n2197 DVSS.n2038 0.00962857
R17872 DVSS.n2197 DVSS.n2040 0.00962857
R17873 DVSS.n2193 DVSS.n2040 0.00962857
R17874 DVSS.n2193 DVSS.n2042 0.00962857
R17875 DVSS.n2189 DVSS.n2042 0.00962857
R17876 DVSS.n2189 DVSS.n2044 0.00962857
R17877 DVSS.n2185 DVSS.n2044 0.00962857
R17878 DVSS.n2185 DVSS.n2046 0.00962857
R17879 DVSS.n2181 DVSS.n2046 0.00962857
R17880 DVSS.n2181 DVSS.n2048 0.00962857
R17881 DVSS.n2177 DVSS.n2048 0.00962857
R17882 DVSS.n2177 DVSS.n2050 0.00962857
R17883 DVSS.n2173 DVSS.n2050 0.00962857
R17884 DVSS.n2173 DVSS.n2052 0.00962857
R17885 DVSS.n2169 DVSS.n2052 0.00962857
R17886 DVSS.n2169 DVSS.n2054 0.00962857
R17887 DVSS.n2165 DVSS.n2054 0.00962857
R17888 DVSS.n2165 DVSS.n2056 0.00962857
R17889 DVSS.n2161 DVSS.n2056 0.00962857
R17890 DVSS.n2161 DVSS.n2058 0.00962857
R17891 DVSS.n2157 DVSS.n2058 0.00962857
R17892 DVSS.n2157 DVSS.n2060 0.00962857
R17893 DVSS.n2153 DVSS.n2060 0.00962857
R17894 DVSS.n2153 DVSS.n2062 0.00962857
R17895 DVSS.n2149 DVSS.n2062 0.00962857
R17896 DVSS.n2149 DVSS.n2147 0.00962857
R17897 DVSS.n2147 DVSS.n2146 0.00962857
R17898 DVSS.n2146 DVSS.n2064 0.00962857
R17899 DVSS.n2142 DVSS.n2064 0.00962857
R17900 DVSS.n2142 DVSS.n2066 0.00962857
R17901 DVSS.n2138 DVSS.n2066 0.00962857
R17902 DVSS.n2138 DVSS.n2069 0.00962857
R17903 DVSS.n2134 DVSS.n2069 0.00962857
R17904 DVSS.n2134 DVSS.n2071 0.00962857
R17905 DVSS.n2130 DVSS.n2071 0.00962857
R17906 DVSS.n2130 DVSS.n2073 0.00962857
R17907 DVSS.n2126 DVSS.n2073 0.00962857
R17908 DVSS.n2126 DVSS.n2075 0.00962857
R17909 DVSS.n2122 DVSS.n2075 0.00962857
R17910 DVSS.n2122 DVSS.n2077 0.00962857
R17911 DVSS.n2118 DVSS.n2077 0.00962857
R17912 DVSS.n2118 DVSS.n2079 0.00962857
R17913 DVSS.n2114 DVSS.n2079 0.00962857
R17914 DVSS.n2114 DVSS.n2081 0.00962857
R17915 DVSS.n2110 DVSS.n2081 0.00962857
R17916 DVSS.n2110 DVSS.n2083 0.00962857
R17917 DVSS.n2106 DVSS.n2083 0.00962857
R17918 DVSS.n2106 DVSS.n2085 0.00962857
R17919 DVSS.n2102 DVSS.n2085 0.00962857
R17920 DVSS.n2102 DVSS.n2087 0.00962857
R17921 DVSS.n2098 DVSS.n2087 0.00962857
R17922 DVSS.n2098 DVSS.n2089 0.00962857
R17923 DVSS.n2094 DVSS.n2089 0.00962857
R17924 DVSS.n2022 DVSS.n2021 0.00962857
R17925 DVSS.n2023 DVSS.n2022 0.00962857
R17926 DVSS.n2023 DVSS.n1960 0.00962857
R17927 DVSS.n2220 DVSS.n2219 0.00962857
R17928 DVSS.n2219 DVSS.n2218 0.00962857
R17929 DVSS.n2218 DVSS.n2029 0.00962857
R17930 DVSS.n2212 DVSS.n2029 0.00962857
R17931 DVSS.n2212 DVSS.n2211 0.00962857
R17932 DVSS.n2211 DVSS.n2210 0.00962857
R17933 DVSS.n2210 DVSS.n2033 0.00962857
R17934 DVSS.n2204 DVSS.n2033 0.00962857
R17935 DVSS.n2204 DVSS.n2203 0.00962857
R17936 DVSS.n2203 DVSS.n2202 0.00962857
R17937 DVSS.n2202 DVSS.n2037 0.00962857
R17938 DVSS.n2196 DVSS.n2037 0.00962857
R17939 DVSS.n2196 DVSS.n2195 0.00962857
R17940 DVSS.n2195 DVSS.n2194 0.00962857
R17941 DVSS.n2194 DVSS.n2041 0.00962857
R17942 DVSS.n2188 DVSS.n2041 0.00962857
R17943 DVSS.n2188 DVSS.n2187 0.00962857
R17944 DVSS.n2187 DVSS.n2186 0.00962857
R17945 DVSS.n2186 DVSS.n2045 0.00962857
R17946 DVSS.n2180 DVSS.n2045 0.00962857
R17947 DVSS.n2180 DVSS.n2179 0.00962857
R17948 DVSS.n2179 DVSS.n2178 0.00962857
R17949 DVSS.n2178 DVSS.n2049 0.00962857
R17950 DVSS.n2172 DVSS.n2049 0.00962857
R17951 DVSS.n2172 DVSS.n2171 0.00962857
R17952 DVSS.n2171 DVSS.n2170 0.00962857
R17953 DVSS.n2170 DVSS.n2053 0.00962857
R17954 DVSS.n2164 DVSS.n2053 0.00962857
R17955 DVSS.n2164 DVSS.n2163 0.00962857
R17956 DVSS.n2163 DVSS.n2162 0.00962857
R17957 DVSS.n2162 DVSS.n2057 0.00962857
R17958 DVSS.n2156 DVSS.n2057 0.00962857
R17959 DVSS.n2156 DVSS.n2155 0.00962857
R17960 DVSS.n2155 DVSS.n2154 0.00962857
R17961 DVSS.n2154 DVSS.n2061 0.00962857
R17962 DVSS.n2067 DVSS.n1534 0.00962857
R17963 DVSS.n2141 DVSS.n2067 0.00962857
R17964 DVSS.n2141 DVSS.n2140 0.00962857
R17965 DVSS.n2140 DVSS.n2139 0.00962857
R17966 DVSS.n2139 DVSS.n2068 0.00962857
R17967 DVSS.n2133 DVSS.n2068 0.00962857
R17968 DVSS.n2133 DVSS.n2132 0.00962857
R17969 DVSS.n2132 DVSS.n2131 0.00962857
R17970 DVSS.n2131 DVSS.n2072 0.00962857
R17971 DVSS.n2125 DVSS.n2072 0.00962857
R17972 DVSS.n2125 DVSS.n2124 0.00962857
R17973 DVSS.n2124 DVSS.n2123 0.00962857
R17974 DVSS.n2123 DVSS.n2076 0.00962857
R17975 DVSS.n2117 DVSS.n2076 0.00962857
R17976 DVSS.n2117 DVSS.n2116 0.00962857
R17977 DVSS.n2116 DVSS.n2115 0.00962857
R17978 DVSS.n2115 DVSS.n2080 0.00962857
R17979 DVSS.n2109 DVSS.n2080 0.00962857
R17980 DVSS.n2109 DVSS.n2108 0.00962857
R17981 DVSS.n2108 DVSS.n2107 0.00962857
R17982 DVSS.n2107 DVSS.n2084 0.00962857
R17983 DVSS.n2101 DVSS.n2084 0.00962857
R17984 DVSS.n2101 DVSS.n2100 0.00962857
R17985 DVSS.n2100 DVSS.n2099 0.00962857
R17986 DVSS.n2099 DVSS.n2088 0.00962857
R17987 DVSS.n2093 DVSS.n2088 0.00962857
R17988 DVSS.n2614 DVSS.n1850 0.00962857
R17989 DVSS.n2607 DVSS.n1854 0.00962857
R17990 DVSS.n2607 DVSS.n2606 0.00962857
R17991 DVSS.n2606 DVSS.n2605 0.00962857
R17992 DVSS.n2564 DVSS.n1905 0.00962857
R17993 DVSS.n2558 DVSS.n1905 0.00962857
R17994 DVSS.n2468 DVSS.n2467 0.00962857
R17995 DVSS.n2467 DVSS.n2466 0.00962857
R17996 DVSS.n2466 DVSS.n2379 0.00962857
R17997 DVSS.n2460 DVSS.n2379 0.00962857
R17998 DVSS.n2460 DVSS.n2459 0.00962857
R17999 DVSS.n2459 DVSS.n2458 0.00962857
R18000 DVSS.n2458 DVSS.n2384 0.00962857
R18001 DVSS.n2452 DVSS.n2384 0.00962857
R18002 DVSS.n2452 DVSS.n2451 0.00962857
R18003 DVSS.n2451 DVSS.n2450 0.00962857
R18004 DVSS.n2450 DVSS.n2388 0.00962857
R18005 DVSS.n2444 DVSS.n2388 0.00962857
R18006 DVSS.n2444 DVSS.n2443 0.00962857
R18007 DVSS.n2443 DVSS.n2442 0.00962857
R18008 DVSS.n2442 DVSS.n2392 0.00962857
R18009 DVSS.n2436 DVSS.n2392 0.00962857
R18010 DVSS.n2436 DVSS.n2435 0.00962857
R18011 DVSS.n2435 DVSS.n2434 0.00962857
R18012 DVSS.n2434 DVSS.n2396 0.00962857
R18013 DVSS.n2428 DVSS.n2396 0.00962857
R18014 DVSS.n2428 DVSS.n2427 0.00962857
R18015 DVSS.n2427 DVSS.n2426 0.00962857
R18016 DVSS.n2426 DVSS.n2400 0.00962857
R18017 DVSS.n2420 DVSS.n2400 0.00962857
R18018 DVSS.n2420 DVSS.n2419 0.00962857
R18019 DVSS.n2419 DVSS.n2418 0.00962857
R18020 DVSS.n2418 DVSS.n2404 0.00962857
R18021 DVSS.n2412 DVSS.n2404 0.00962857
R18022 DVSS.n2412 DVSS.n2411 0.00962857
R18023 DVSS.n1633 DVSS.n1629 0.00962857
R18024 DVSS.n4046 DVSS.n1629 0.00962857
R18025 DVSS.n4046 DVSS.n1630 0.00962857
R18026 DVSS.n4042 DVSS.n1630 0.00962857
R18027 DVSS.n4042 DVSS.n1637 0.00962857
R18028 DVSS.n4037 DVSS.n1637 0.00962857
R18029 DVSS.n4037 DVSS.n1639 0.00962857
R18030 DVSS.n4033 DVSS.n1639 0.00962857
R18031 DVSS.n4033 DVSS.n1641 0.00962857
R18032 DVSS.n4027 DVSS.n1641 0.00962857
R18033 DVSS.n4027 DVSS.n1643 0.00962857
R18034 DVSS.n4023 DVSS.n1643 0.00962857
R18035 DVSS.n4023 DVSS.n1645 0.00962857
R18036 DVSS.n4019 DVSS.n1645 0.00962857
R18037 DVSS.n4019 DVSS.n1648 0.00962857
R18038 DVSS.n4015 DVSS.n1648 0.00962857
R18039 DVSS.n4015 DVSS.n1650 0.00962857
R18040 DVSS.n4008 DVSS.n1650 0.00962857
R18041 DVSS.n4008 DVSS.n1653 0.00962857
R18042 DVSS.n4004 DVSS.n1653 0.00962857
R18043 DVSS.n4004 DVSS.n1655 0.00962857
R18044 DVSS.n4000 DVSS.n1655 0.00962857
R18045 DVSS.n4000 DVSS.n1658 0.00962857
R18046 DVSS.n3996 DVSS.n1658 0.00962857
R18047 DVSS.n3996 DVSS.n1660 0.00962857
R18048 DVSS.n3980 DVSS.n1660 0.00962857
R18049 DVSS.n3980 DVSS.n1671 0.00962857
R18050 DVSS.n3976 DVSS.n1671 0.00962857
R18051 DVSS.n3976 DVSS.n1673 0.00962857
R18052 DVSS.n3972 DVSS.n1673 0.00962857
R18053 DVSS.n3972 DVSS.n1675 0.00962857
R18054 DVSS.n3968 DVSS.n1675 0.00962857
R18055 DVSS.n3968 DVSS.n1677 0.00962857
R18056 DVSS.n3964 DVSS.n1677 0.00962857
R18057 DVSS.n3964 DVSS.n1679 0.00962857
R18058 DVSS.n3960 DVSS.n1679 0.00962857
R18059 DVSS.n3960 DVSS.n1681 0.00962857
R18060 DVSS.n1689 DVSS.n1681 0.00962857
R18061 DVSS.n3951 DVSS.n1689 0.00962857
R18062 DVSS.n3951 DVSS.n1690 0.00962857
R18063 DVSS.n3947 DVSS.n1690 0.00962857
R18064 DVSS.n3947 DVSS.n1693 0.00962857
R18065 DVSS.n1712 DVSS.n1693 0.00962857
R18066 DVSS.n1715 DVSS.n1712 0.00962857
R18067 DVSS.n1715 DVSS.n1709 0.00962857
R18068 DVSS.n3928 DVSS.n1709 0.00962857
R18069 DVSS.n3928 DVSS.n1710 0.00962857
R18070 DVSS.n3924 DVSS.n1710 0.00962857
R18071 DVSS.n3924 DVSS.n1719 0.00962857
R18072 DVSS.n3920 DVSS.n1719 0.00962857
R18073 DVSS.n3920 DVSS.n1723 0.00962857
R18074 DVSS.n3916 DVSS.n1723 0.00962857
R18075 DVSS.n3916 DVSS.n1725 0.00962857
R18076 DVSS.n3912 DVSS.n1725 0.00962857
R18077 DVSS.n3912 DVSS.n1731 0.00962857
R18078 DVSS.n3908 DVSS.n1731 0.00962857
R18079 DVSS.n3908 DVSS.n1733 0.00962857
R18080 DVSS.n3904 DVSS.n1733 0.00962857
R18081 DVSS.n3904 DVSS.n1737 0.00962857
R18082 DVSS.n3900 DVSS.n1737 0.00962857
R18083 DVSS.n3900 DVSS.n1739 0.00962857
R18084 DVSS.n3896 DVSS.n1739 0.00962857
R18085 DVSS.n3896 DVSS.n1741 0.00962857
R18086 DVSS.n3892 DVSS.n1741 0.00962857
R18087 DVSS.n3892 DVSS.n1743 0.00962857
R18088 DVSS.n3888 DVSS.n1743 0.00962857
R18089 DVSS.n3888 DVSS.n1745 0.00962857
R18090 DVSS.n3884 DVSS.n1745 0.00962857
R18091 DVSS.n3884 DVSS.n1747 0.00962857
R18092 DVSS.n3880 DVSS.n1747 0.00962857
R18093 DVSS.n3880 DVSS.n1749 0.00962857
R18094 DVSS.n3876 DVSS.n1749 0.00962857
R18095 DVSS.n3876 DVSS.n1751 0.00962857
R18096 DVSS.n3872 DVSS.n1751 0.00962857
R18097 DVSS.n3872 DVSS.n1753 0.00962857
R18098 DVSS.n3868 DVSS.n1753 0.00962857
R18099 DVSS.n3868 DVSS.n1755 0.00962857
R18100 DVSS.n1775 DVSS.n1755 0.00962857
R18101 DVSS.n1775 DVSS.n1757 0.00962857
R18102 DVSS.n1771 DVSS.n1757 0.00962857
R18103 DVSS.n1771 DVSS.n1759 0.00962857
R18104 DVSS.n1767 DVSS.n1759 0.00962857
R18105 DVSS.n1767 DVSS.n1761 0.00962857
R18106 DVSS.n1632 DVSS.n1627 0.00962857
R18107 DVSS.n4047 DVSS.n1628 0.00962857
R18108 DVSS.n4041 DVSS.n1628 0.00962857
R18109 DVSS.n4039 DVSS.n4038 0.00962857
R18110 DVSS.n4038 DVSS.n1638 0.00962857
R18111 DVSS.n4032 DVSS.n1638 0.00962857
R18112 DVSS.n4022 DVSS.n1646 0.00962857
R18113 DVSS.n4022 DVSS.n4021 0.00962857
R18114 DVSS.n4021 DVSS.n4020 0.00962857
R18115 DVSS.n4014 DVSS.n1651 0.00962857
R18116 DVSS.n4014 DVSS.n4013 0.00962857
R18117 DVSS.n4003 DVSS.n1656 0.00962857
R18118 DVSS.n4003 DVSS.n4002 0.00962857
R18119 DVSS.n4002 DVSS.n4001 0.00962857
R18120 DVSS.n3982 DVSS.n3981 0.00962857
R18121 DVSS.n3981 DVSS.n1670 0.00962857
R18122 DVSS.n3975 DVSS.n1670 0.00962857
R18123 DVSS.n3975 DVSS.n3974 0.00962857
R18124 DVSS.n3974 DVSS.n3973 0.00962857
R18125 DVSS.n3973 DVSS.n1674 0.00962857
R18126 DVSS.n3967 DVSS.n1674 0.00962857
R18127 DVSS.n3967 DVSS.n3966 0.00962857
R18128 DVSS.n3966 DVSS.n3965 0.00962857
R18129 DVSS.n3965 DVSS.n1678 0.00962857
R18130 DVSS.n3959 DVSS.n1678 0.00962857
R18131 DVSS.n1687 DVSS.n1682 0.00962857
R18132 DVSS.n3952 DVSS.n1688 0.00962857
R18133 DVSS.n3946 DVSS.n1688 0.00962857
R18134 DVSS.n1713 DVSS.n1694 0.00962857
R18135 DVSS.n1714 DVSS.n1713 0.00962857
R18136 DVSS.n1714 DVSS.n1707 0.00962857
R18137 DVSS.n3923 DVSS.n3922 0.00962857
R18138 DVSS.n3922 DVSS.n3921 0.00962857
R18139 DVSS.n3921 DVSS.n1722 0.00962857
R18140 DVSS.n3915 DVSS.n3914 0.00962857
R18141 DVSS.n3914 DVSS.n3913 0.00962857
R18142 DVSS.n3907 DVSS.n3906 0.00962857
R18143 DVSS.n3906 DVSS.n3905 0.00962857
R18144 DVSS.n3905 DVSS.n1736 0.00962857
R18145 DVSS.n3899 DVSS.n1736 0.00962857
R18146 DVSS.n3899 DVSS.n3898 0.00962857
R18147 DVSS.n3898 DVSS.n3897 0.00962857
R18148 DVSS.n3897 DVSS.n1740 0.00962857
R18149 DVSS.n3891 DVSS.n1740 0.00962857
R18150 DVSS.n3891 DVSS.n3890 0.00962857
R18151 DVSS.n3890 DVSS.n3889 0.00962857
R18152 DVSS.n3889 DVSS.n1744 0.00962857
R18153 DVSS.n3883 DVSS.n1744 0.00962857
R18154 DVSS.n3883 DVSS.n3882 0.00962857
R18155 DVSS.n3882 DVSS.n3881 0.00962857
R18156 DVSS.n3881 DVSS.n1748 0.00962857
R18157 DVSS.n3875 DVSS.n1748 0.00962857
R18158 DVSS.n3875 DVSS.n3874 0.00962857
R18159 DVSS.n3874 DVSS.n3873 0.00962857
R18160 DVSS.n3873 DVSS.n1752 0.00962857
R18161 DVSS.n3867 DVSS.n1752 0.00962857
R18162 DVSS.n1777 DVSS.n1776 0.00962857
R18163 DVSS.n1776 DVSS.n1756 0.00962857
R18164 DVSS.n1770 DVSS.n1756 0.00962857
R18165 DVSS.n1770 DVSS.n1769 0.00962857
R18166 DVSS.n1769 DVSS.n1768 0.00962857
R18167 DVSS.n1768 DVSS.n1760 0.00962857
R18168 DVSS.n5089 DVSS.n1083 0.00962857
R18169 DVSS.n5089 DVSS.n1085 0.00962857
R18170 DVSS.n5085 DVSS.n1085 0.00962857
R18171 DVSS.n5085 DVSS.n1087 0.00962857
R18172 DVSS.n5081 DVSS.n1087 0.00962857
R18173 DVSS.n5081 DVSS.n1089 0.00962857
R18174 DVSS.n5077 DVSS.n1089 0.00962857
R18175 DVSS.n5077 DVSS.n1091 0.00962857
R18176 DVSS.n5073 DVSS.n1091 0.00962857
R18177 DVSS.n5073 DVSS.n1093 0.00962857
R18178 DVSS.n5069 DVSS.n1093 0.00962857
R18179 DVSS.n5069 DVSS.n1095 0.00962857
R18180 DVSS.n5065 DVSS.n1095 0.00962857
R18181 DVSS.n5065 DVSS.n1097 0.00962857
R18182 DVSS.n5060 DVSS.n1097 0.00962857
R18183 DVSS.n5060 DVSS.n1100 0.00962857
R18184 DVSS.n5056 DVSS.n1100 0.00962857
R18185 DVSS.n5056 DVSS.n1102 0.00962857
R18186 DVSS.n5052 DVSS.n1102 0.00962857
R18187 DVSS.n5052 DVSS.n1105 0.00962857
R18188 DVSS.n5048 DVSS.n1105 0.00962857
R18189 DVSS.n5048 DVSS.n1107 0.00962857
R18190 DVSS.n1111 DVSS.n1107 0.00962857
R18191 DVSS.n5041 DVSS.n1111 0.00962857
R18192 DVSS.n5041 DVSS.n1112 0.00962857
R18193 DVSS.n5037 DVSS.n1112 0.00962857
R18194 DVSS.n5037 DVSS.n1115 0.00962857
R18195 DVSS.n5030 DVSS.n1115 0.00962857
R18196 DVSS.n5030 DVSS.n1123 0.00962857
R18197 DVSS.n5026 DVSS.n1123 0.00962857
R18198 DVSS.n5026 DVSS.n1125 0.00962857
R18199 DVSS.n5022 DVSS.n1125 0.00962857
R18200 DVSS.n5022 DVSS.n1129 0.00962857
R18201 DVSS.n5018 DVSS.n1129 0.00962857
R18202 DVSS.n5018 DVSS.n1131 0.00962857
R18203 DVSS.n5014 DVSS.n1131 0.00962857
R18204 DVSS.n5014 DVSS.n1133 0.00962857
R18205 DVSS.n5010 DVSS.n1133 0.00962857
R18206 DVSS.n5010 DVSS.n1135 0.00962857
R18207 DVSS.n5006 DVSS.n1135 0.00962857
R18208 DVSS.n5006 DVSS.n1137 0.00962857
R18209 DVSS.n5002 DVSS.n1137 0.00962857
R18210 DVSS.n5002 DVSS.n1139 0.00962857
R18211 DVSS.n4998 DVSS.n1139 0.00962857
R18212 DVSS.n4998 DVSS.n1141 0.00962857
R18213 DVSS.n4994 DVSS.n1141 0.00962857
R18214 DVSS.n4994 DVSS.n1143 0.00962857
R18215 DVSS.n4990 DVSS.n1143 0.00962857
R18216 DVSS.n4990 DVSS.n1145 0.00962857
R18217 DVSS.n4986 DVSS.n1145 0.00962857
R18218 DVSS.n4986 DVSS.n1147 0.00962857
R18219 DVSS.n4982 DVSS.n1147 0.00962857
R18220 DVSS.n4982 DVSS.n1149 0.00962857
R18221 DVSS.n4978 DVSS.n1149 0.00962857
R18222 DVSS.n4978 DVSS.n1151 0.00962857
R18223 DVSS.n4974 DVSS.n1151 0.00962857
R18224 DVSS.n4974 DVSS.n1153 0.00962857
R18225 DVSS.n4970 DVSS.n1153 0.00962857
R18226 DVSS.n4970 DVSS.n1155 0.00962857
R18227 DVSS.n4966 DVSS.n1155 0.00962857
R18228 DVSS.n4966 DVSS.n1157 0.00962857
R18229 DVSS.n4962 DVSS.n1157 0.00962857
R18230 DVSS.n4962 DVSS.n1159 0.00962857
R18231 DVSS.n4958 DVSS.n1159 0.00962857
R18232 DVSS.n4958 DVSS.n1162 0.00962857
R18233 DVSS.n4954 DVSS.n1162 0.00962857
R18234 DVSS.n4954 DVSS.n1164 0.00962857
R18235 DVSS.n4950 DVSS.n1164 0.00962857
R18236 DVSS.n4950 DVSS.n1166 0.00962857
R18237 DVSS.n4946 DVSS.n1166 0.00962857
R18238 DVSS.n4946 DVSS.n1168 0.00962857
R18239 DVSS.n4942 DVSS.n1168 0.00962857
R18240 DVSS.n4942 DVSS.n1170 0.00962857
R18241 DVSS.n4938 DVSS.n1170 0.00962857
R18242 DVSS.n4938 DVSS.n1172 0.00962857
R18243 DVSS.n4934 DVSS.n1172 0.00962857
R18244 DVSS.n4934 DVSS.n1174 0.00962857
R18245 DVSS.n4930 DVSS.n1174 0.00962857
R18246 DVSS.n4930 DVSS.n1176 0.00962857
R18247 DVSS.n4926 DVSS.n1176 0.00962857
R18248 DVSS.n4926 DVSS.n1178 0.00962857
R18249 DVSS.n4922 DVSS.n1178 0.00962857
R18250 DVSS.n4922 DVSS.n1180 0.00962857
R18251 DVSS.n4918 DVSS.n1180 0.00962857
R18252 DVSS.n4918 DVSS.n1182 0.00962857
R18253 DVSS.n4914 DVSS.n1182 0.00962857
R18254 DVSS.n4914 DVSS.n1184 0.00962857
R18255 DVSS.n4910 DVSS.n1184 0.00962857
R18256 DVSS.n4910 DVSS.n1186 0.00962857
R18257 DVSS.n4906 DVSS.n1186 0.00962857
R18258 DVSS.n4906 DVSS.n1188 0.00962857
R18259 DVSS.n4902 DVSS.n1188 0.00962857
R18260 DVSS.n4902 DVSS.n1190 0.00962857
R18261 DVSS.n4898 DVSS.n1190 0.00962857
R18262 DVSS.n4898 DVSS.n1192 0.00962857
R18263 DVSS.n4894 DVSS.n1192 0.00962857
R18264 DVSS.n4894 DVSS.n1194 0.00962857
R18265 DVSS.n4890 DVSS.n1195 0.00962857
R18266 DVSS.n3518 DVSS.n1195 0.00962857
R18267 DVSS.n3518 DVSS.n3515 0.00962857
R18268 DVSS.n5092 DVSS.n1082 0.00962857
R18269 DVSS.n5088 DVSS.n1082 0.00962857
R18270 DVSS.n5088 DVSS.n5087 0.00962857
R18271 DVSS.n5087 DVSS.n5086 0.00962857
R18272 DVSS.n5086 DVSS.n1086 0.00962857
R18273 DVSS.n5080 DVSS.n1086 0.00962857
R18274 DVSS.n5080 DVSS.n5079 0.00962857
R18275 DVSS.n5079 DVSS.n5078 0.00962857
R18276 DVSS.n5078 DVSS.n1090 0.00962857
R18277 DVSS.n5072 DVSS.n1090 0.00962857
R18278 DVSS.n5072 DVSS.n5071 0.00962857
R18279 DVSS.n5071 DVSS.n5070 0.00962857
R18280 DVSS.n5070 DVSS.n1094 0.00962857
R18281 DVSS.n5064 DVSS.n1094 0.00962857
R18282 DVSS.n5064 DVSS.n5063 0.00962857
R18283 DVSS.n5055 DVSS.n1103 0.00962857
R18284 DVSS.n5055 DVSS.n5054 0.00962857
R18285 DVSS.n5054 DVSS.n5053 0.00962857
R18286 DVSS.n5053 DVSS.n1104 0.00962857
R18287 DVSS.n5047 DVSS.n1104 0.00962857
R18288 DVSS.n5047 DVSS.n5046 0.00962857
R18289 DVSS.n5025 DVSS.n5024 0.00962857
R18290 DVSS.n5024 DVSS.n5023 0.00962857
R18291 DVSS.n5023 DVSS.n1128 0.00962857
R18292 DVSS.n5017 DVSS.n1128 0.00962857
R18293 DVSS.n5017 DVSS.n5016 0.00962857
R18294 DVSS.n5016 DVSS.n5015 0.00962857
R18295 DVSS.n5015 DVSS.n1132 0.00962857
R18296 DVSS.n5009 DVSS.n1132 0.00962857
R18297 DVSS.n5009 DVSS.n5008 0.00962857
R18298 DVSS.n5008 DVSS.n5007 0.00962857
R18299 DVSS.n5007 DVSS.n1136 0.00962857
R18300 DVSS.n5001 DVSS.n1136 0.00962857
R18301 DVSS.n5001 DVSS.n5000 0.00962857
R18302 DVSS.n5000 DVSS.n4999 0.00962857
R18303 DVSS.n4999 DVSS.n1140 0.00962857
R18304 DVSS.n4993 DVSS.n1140 0.00962857
R18305 DVSS.n4993 DVSS.n4992 0.00962857
R18306 DVSS.n4992 DVSS.n4991 0.00962857
R18307 DVSS.n4991 DVSS.n1144 0.00962857
R18308 DVSS.n4985 DVSS.n1144 0.00962857
R18309 DVSS.n4985 DVSS.n4984 0.00962857
R18310 DVSS.n4984 DVSS.n4983 0.00962857
R18311 DVSS.n4983 DVSS.n1148 0.00962857
R18312 DVSS.n4977 DVSS.n1148 0.00962857
R18313 DVSS.n4977 DVSS.n4976 0.00962857
R18314 DVSS.n4976 DVSS.n4975 0.00962857
R18315 DVSS.n4975 DVSS.n1152 0.00962857
R18316 DVSS.n4969 DVSS.n1152 0.00962857
R18317 DVSS.n4969 DVSS.n4968 0.00962857
R18318 DVSS.n4968 DVSS.n4967 0.00962857
R18319 DVSS.n4961 DVSS.n1160 0.00962857
R18320 DVSS.n4961 DVSS.n4960 0.00962857
R18321 DVSS.n4960 DVSS.n4959 0.00962857
R18322 DVSS.n4959 DVSS.n1161 0.00962857
R18323 DVSS.n4953 DVSS.n1161 0.00962857
R18324 DVSS.n4953 DVSS.n4952 0.00962857
R18325 DVSS.n4952 DVSS.n4951 0.00962857
R18326 DVSS.n4951 DVSS.n1165 0.00962857
R18327 DVSS.n4945 DVSS.n1165 0.00962857
R18328 DVSS.n4945 DVSS.n4944 0.00962857
R18329 DVSS.n4944 DVSS.n4943 0.00962857
R18330 DVSS.n4943 DVSS.n1169 0.00962857
R18331 DVSS.n4937 DVSS.n1169 0.00962857
R18332 DVSS.n4937 DVSS.n4936 0.00962857
R18333 DVSS.n4936 DVSS.n4935 0.00962857
R18334 DVSS.n4935 DVSS.n1173 0.00962857
R18335 DVSS.n4929 DVSS.n1173 0.00962857
R18336 DVSS.n4929 DVSS.n4928 0.00962857
R18337 DVSS.n4928 DVSS.n4927 0.00962857
R18338 DVSS.n4927 DVSS.n1177 0.00962857
R18339 DVSS.n4921 DVSS.n1177 0.00962857
R18340 DVSS.n4921 DVSS.n4920 0.00962857
R18341 DVSS.n4920 DVSS.n4919 0.00962857
R18342 DVSS.n4919 DVSS.n1181 0.00962857
R18343 DVSS.n4913 DVSS.n1181 0.00962857
R18344 DVSS.n4913 DVSS.n4912 0.00962857
R18345 DVSS.n4912 DVSS.n4911 0.00962857
R18346 DVSS.n4911 DVSS.n1185 0.00962857
R18347 DVSS.n4905 DVSS.n1185 0.00962857
R18348 DVSS.n4905 DVSS.n4904 0.00962857
R18349 DVSS.n4904 DVSS.n4903 0.00962857
R18350 DVSS.n4903 DVSS.n1189 0.00962857
R18351 DVSS.n4897 DVSS.n1189 0.00962857
R18352 DVSS.n4897 DVSS.n4896 0.00962857
R18353 DVSS.n4896 DVSS.n4895 0.00962857
R18354 DVSS.n3517 DVSS.n1199 0.00962857
R18355 DVSS.n3517 DVSS.n3514 0.00962857
R18356 DVSS.n3521 DVSS.n3514 0.00962857
R18357 DVSS.n1574 DVSS.n1571 0.00962857
R18358 DVSS.n1575 DVSS.n1574 0.00962857
R18359 DVSS.n1576 DVSS.n1575 0.00962857
R18360 DVSS.n1576 DVSS.n1567 0.00962857
R18361 DVSS.n1582 DVSS.n1567 0.00962857
R18362 DVSS.n1583 DVSS.n1582 0.00962857
R18363 DVSS.n1584 DVSS.n1583 0.00962857
R18364 DVSS.n1584 DVSS.n1563 0.00962857
R18365 DVSS.n1590 DVSS.n1563 0.00962857
R18366 DVSS.n1591 DVSS.n1590 0.00962857
R18367 DVSS.n1592 DVSS.n1591 0.00962857
R18368 DVSS.n1592 DVSS.n1557 0.00962857
R18369 DVSS.n4090 DVSS.n1558 0.00962857
R18370 DVSS.n4084 DVSS.n1558 0.00962857
R18371 DVSS.n4084 DVSS.n4083 0.00962857
R18372 DVSS.n4083 DVSS.n4082 0.00962857
R18373 DVSS.n4082 DVSS.n1598 0.00962857
R18374 DVSS.n4076 DVSS.n1598 0.00962857
R18375 DVSS.n4076 DVSS.n4075 0.00962857
R18376 DVSS.n4075 DVSS.n4074 0.00962857
R18377 DVSS.n4074 DVSS.n1602 0.00962857
R18378 DVSS.n4068 DVSS.n1602 0.00962857
R18379 DVSS.n4068 DVSS.n4067 0.00962857
R18380 DVSS.n4067 DVSS.n4066 0.00962857
R18381 DVSS.n4066 DVSS.n1606 0.00962857
R18382 DVSS.n4060 DVSS.n1606 0.00962857
R18383 DVSS.n3606 DVSS.n1610 0.00962857
R18384 DVSS.n3611 DVSS.n3606 0.00962857
R18385 DVSS.n3612 DVSS.n3611 0.00962857
R18386 DVSS.n3613 DVSS.n3612 0.00962857
R18387 DVSS.n3613 DVSS.n3602 0.00962857
R18388 DVSS.n3619 DVSS.n3602 0.00962857
R18389 DVSS.n3620 DVSS.n3619 0.00962857
R18390 DVSS.n3621 DVSS.n3620 0.00962857
R18391 DVSS.n3621 DVSS.n3598 0.00962857
R18392 DVSS.n3627 DVSS.n3598 0.00962857
R18393 DVSS.n3628 DVSS.n3627 0.00962857
R18394 DVSS.n3629 DVSS.n3628 0.00962857
R18395 DVSS.n3629 DVSS.n3594 0.00962857
R18396 DVSS.n3635 DVSS.n3594 0.00962857
R18397 DVSS.n3636 DVSS.n3635 0.00962857
R18398 DVSS.n3637 DVSS.n3636 0.00962857
R18399 DVSS.n3637 DVSS.n3590 0.00962857
R18400 DVSS.n3643 DVSS.n3590 0.00962857
R18401 DVSS.n3644 DVSS.n3643 0.00962857
R18402 DVSS.n3645 DVSS.n3644 0.00962857
R18403 DVSS.n3645 DVSS.n3586 0.00962857
R18404 DVSS.n3651 DVSS.n3586 0.00962857
R18405 DVSS.n3652 DVSS.n3651 0.00962857
R18406 DVSS.n3653 DVSS.n3652 0.00962857
R18407 DVSS.n3653 DVSS.n3582 0.00962857
R18408 DVSS.n3659 DVSS.n3582 0.00962857
R18409 DVSS.n3660 DVSS.n3659 0.00962857
R18410 DVSS.n3661 DVSS.n3660 0.00962857
R18411 DVSS.n3661 DVSS.n3578 0.00962857
R18412 DVSS.n3667 DVSS.n3578 0.00962857
R18413 DVSS.n3668 DVSS.n3667 0.00962857
R18414 DVSS.n3669 DVSS.n3668 0.00962857
R18415 DVSS.n3669 DVSS.n3574 0.00962857
R18416 DVSS.n3675 DVSS.n3574 0.00962857
R18417 DVSS.n3676 DVSS.n3675 0.00962857
R18418 DVSS.n3677 DVSS.n3676 0.00962857
R18419 DVSS.n3677 DVSS.n3570 0.00962857
R18420 DVSS.n3683 DVSS.n3570 0.00962857
R18421 DVSS.n3684 DVSS.n3683 0.00962857
R18422 DVSS.n3685 DVSS.n3684 0.00962857
R18423 DVSS.n3685 DVSS.n3566 0.00962857
R18424 DVSS.n3691 DVSS.n3566 0.00962857
R18425 DVSS.n3692 DVSS.n3691 0.00962857
R18426 DVSS.n3693 DVSS.n3692 0.00962857
R18427 DVSS.n3693 DVSS.n3562 0.00962857
R18428 DVSS.n3699 DVSS.n3562 0.00962857
R18429 DVSS.n3700 DVSS.n3699 0.00962857
R18430 DVSS.n3701 DVSS.n3700 0.00962857
R18431 DVSS.n3701 DVSS.n3558 0.00962857
R18432 DVSS.n3707 DVSS.n3558 0.00962857
R18433 DVSS.n3708 DVSS.n3707 0.00962857
R18434 DVSS.n3709 DVSS.n3708 0.00962857
R18435 DVSS.n3709 DVSS.n3554 0.00962857
R18436 DVSS.n3715 DVSS.n3554 0.00962857
R18437 DVSS.n3716 DVSS.n3715 0.00962857
R18438 DVSS.n3717 DVSS.n3716 0.00962857
R18439 DVSS.n3717 DVSS.n3550 0.00962857
R18440 DVSS.n3723 DVSS.n3550 0.00962857
R18441 DVSS.n3724 DVSS.n3723 0.00962857
R18442 DVSS.n3725 DVSS.n3724 0.00962857
R18443 DVSS.n3725 DVSS.n3546 0.00962857
R18444 DVSS.n3731 DVSS.n3546 0.00962857
R18445 DVSS.n3732 DVSS.n3731 0.00962857
R18446 DVSS.n3733 DVSS.n3732 0.00962857
R18447 DVSS.n3733 DVSS.n3542 0.00962857
R18448 DVSS.n3739 DVSS.n3542 0.00962857
R18449 DVSS.n3740 DVSS.n3739 0.00962857
R18450 DVSS.n3741 DVSS.n3740 0.00962857
R18451 DVSS.n3741 DVSS.n3534 0.00962857
R18452 DVSS.n3763 DVSS.n3762 0.00962857
R18453 DVSS.n3763 DVSS.n3523 0.00962857
R18454 DVSS.n3767 DVSS.n3523 0.00962857
R18455 DVSS.n3266 DVSS 0.00958867
R18456 DVSS.n3256 DVSS 0.00958867
R18457 DVSS.n2518 DVSS.n2517 0.00958257
R18458 DVSS.n2587 DVSS.n1868 0.00958257
R18459 DVSS.n3866 DVSS.n1777 0.00956429
R18460 DVSS.n5711 DVSS.n58 0.0095301
R18461 DVSS.n2598 DVSS.n1860 0.0095
R18462 DVSS.n2280 DVSS.n2279 0.0095
R18463 DVSS.n2286 DVSS.n2285 0.0095
R18464 DVSS.n2278 DVSS.n2275 0.0095
R18465 DVSS.n2289 DVSS.n2288 0.0095
R18466 DVSS.n2584 DVSS.n2582 0.0095
R18467 DVSS.n1884 DVSS.n1878 0.0095
R18468 DVSS.n2576 DVSS.n1885 0.0095
R18469 DVSS.n2575 DVSS.n1886 0.0095
R18470 DVSS.n2566 DVSS.n2564 0.0095
R18471 DVSS.n2317 DVSS.n2313 0.0095
R18472 DVSS.n2525 DVSS.n2318 0.0095
R18473 DVSS.n2524 DVSS.n2319 0.0095
R18474 DVSS.n2350 DVSS.n2349 0.0095
R18475 DVSS.n2372 DVSS.n2370 0.0095
R18476 DVSS.n2371 DVSS.n2339 0.0095
R18477 DVSS.n2511 DVSS.n2510 0.0095
R18478 DVSS.n2471 DVSS.n2340 0.0095
R18479 DVSS.n2504 DVSS.n2472 0.0095
R18480 DVSS.n3484 DVSS.n2693 0.0095
R18481 DVSS.n3475 DVSS.n2709 0.0095
R18482 DVSS.n3292 DVSS.n2965 0.0095
R18483 DVSS.n3283 DVSS.n2981 0.0095
R18484 DVSS.n3041 DVSS.n3040 0.0095
R18485 DVSS.n3052 DVSS.n3050 0.0095
R18486 DVSS.n3238 DVSS.n3237 0.0095
R18487 DVSS.n3248 DVSS.n3246 0.0095
R18488 DVSS.n3474 DVSS.n2713 0.00936699
R18489 DVSS.n3049 DVSS.n3048 0.00936699
R18490 DVSS.n959 DVSS.n957 0.00934354
R18491 DVSS.n5338 DVSS.n959 0.00934354
R18492 DVSS.n4649 DVSS.n4641 0.00933782
R18493 DVSS.n4646 DVSS.n4643 0.00933782
R18494 DVSS.n4646 DVSS.n4641 0.00933782
R18495 DVSS.n4652 DVSS.n4643 0.00933782
R18496 DVSS.n4367 DVSS.n4358 0.00933782
R18497 DVSS.n4361 DVSS.n4358 0.00933782
R18498 DVSS.n4623 DVSS.n4621 0.00928049
R18499 DVSS.n4720 DVSS.n4619 0.00928049
R18500 DVSS.n4590 DVSS.n4589 0.00928049
R18501 DVSS.n4751 DVSS.n4750 0.00928049
R18502 DVSS.n4552 DVSS.n1427 0.00928049
R18503 DVSS.n4564 DVSS.n1419 0.00928049
R18504 DVSS.n4513 DVSS.n1447 0.00928049
R18505 DVSS.n4524 DVSS.n1440 0.00928049
R18506 DVSS.n4430 DVSS.n4428 0.00928049
R18507 DVSS.n4472 DVSS.n4426 0.00928049
R18508 DVSS.n4397 DVSS.n4396 0.00928049
R18509 DVSS.n4503 DVSS.n4502 0.00928049
R18510 DVSS.n5536 DVSS.n855 0.00924286
R18511 DVSS.n5094 DVSS.n1023 0.00910927
R18512 DVSS.n1024 DVSS.n963 0.00910927
R18513 DVSS.n277 DVSS.n276 0.00909873
R18514 DVSS.n3496 DVSS.n3495 0.009
R18515 DVSS.n3464 DVSS.n3463 0.009
R18516 DVSS.n3305 DVSS.n3304 0.009
R18517 DVSS.n3272 DVSS.n3271 0.009
R18518 DVSS.n3030 DVSS.n2678 0.009
R18519 DVSS.n3022 DVSS.n2724 0.009
R18520 DVSS.n3227 DVSS.n2953 0.009
R18521 DVSS.n3001 DVSS.n2997 0.009
R18522 DVSS.n2236 DVSS.n1963 0.00894122
R18523 DVSS.n2236 DVSS.n2228 0.00894122
R18524 DVSS.n3930 DVSS.n3929 0.00892143
R18525 DVSS.n3915 DVSS.n1726 0.00892143
R18526 DVSS.n5063 DVSS.n5062 0.00892143
R18527 DVSS.n5061 DVSS.n1099 0.00892143
R18528 DVSS.n767 DVSS.n57 0.00882776
R18529 DVSS.n2061 DVSS.n1528 0.00879286
R18530 DVSS.n2148 DVSS.n1527 0.00879286
R18531 DVSS.n4155 DVSS.n1529 0.00879286
R18532 DVSS.n4009 DVSS.n1652 0.00879286
R18533 DVSS.n2605 DVSS.n1855 0.0086
R18534 DVSS.n4585 DVSS.n4584 0.00853571
R18535 DVSS.n1408 DVSS.n1405 0.00853571
R18536 DVSS.n4593 DVSS.n4591 0.00853571
R18537 DVSS.n4592 DVSS.n1399 0.00853571
R18538 DVSS.n4749 DVSS.n4748 0.00853571
R18539 DVSS.n4599 DVSS.n1400 0.00853571
R18540 DVSS.n4742 DVSS.n4602 0.00853571
R18541 DVSS.n2249 DVSS.n2226 0.00853571
R18542 DVSS.n1965 DVSS.n1957 0.00853571
R18543 DVSS.n2220 DVSS.n1959 0.00853571
R18544 DVSS.n3959 DVSS.n3958 0.00853571
R18545 DVSS.n3855 DVSS 0.00852817
R18546 DVSS.n3854 DVSS 0.00852817
R18547 DVSS.n3443 DVSS.n2749 0.0085
R18548 DVSS.n2927 DVSS.n2915 0.0085
R18549 DVSS.n3087 DVSS.n2751 0.0085
R18550 DVSS.n3207 DVSS.n3206 0.0085
R18551 DVSS.n4678 DVSS.n1355 0.00847143
R18552 DVSS.n1938 DVSS.n1859 0.00847143
R18553 DVSS.n5046 DVSS.n5045 0.00847143
R18554 DVSS.n5043 DVSS.n1108 0.00847143
R18555 DVSS.n5042 DVSS.n1110 0.00847143
R18556 DVSS.n1117 DVSS.n1116 0.00847143
R18557 DVSS.n5036 DVSS.n5035 0.00847143
R18558 DVSS.n5032 DVSS.n1118 0.00847143
R18559 DVSS.n5031 DVSS.n1122 0.00847143
R18560 DVSS.n1127 DVSS.n1126 0.00847143
R18561 DVSS.n429 DVSS.n241 0.00842994
R18562 DVSS.n2474 DVSS.n1925 0.00834286
R18563 DVSS.n2468 DVSS.n1924 0.00834286
R18564 DVSS.n4031 DVSS.n4030 0.00827857
R18565 DVSS.n1651 DVSS.n1647 0.00827857
R18566 DVSS.n3409 DVSS 0.00825862
R18567 DVSS DVSS.n3122 0.00825862
R18568 DVSS.n4110 DVSS.n4108 0.00823128
R18569 DVSS.n2251 DVSS.n1955 0.00822787
R18570 DVSS.n2244 DVSS.n1961 0.00822787
R18571 DVSS.n4106 DVSS.n4105 0.00821429
R18572 DVSS.n1735 DVSS.n1734 0.00815
R18573 DVSS.n3458 DVSS.n2731 0.00803695
R18574 DVSS.n3061 DVSS.n3020 0.00803695
R18575 DVSS.n3502 DVSS.n2669 0.00803521
R18576 DVSS.n3028 DVSS.n2670 0.00803521
R18577 DVSS.n3494 DVSS.n2677 0.00803521
R18578 DVSS.n3493 DVSS.n2679 0.00803521
R18579 DVSS.n3490 DVSS.n3489 0.00803521
R18580 DVSS.n3039 DVSS.n2690 0.00803521
R18581 DVSS.n3482 DVSS.n2697 0.00803521
R18582 DVSS.n3481 DVSS.n2699 0.00803521
R18583 DVSS.n3478 DVSS.n3477 0.00803521
R18584 DVSS.n3051 DVSS.n2707 0.00803521
R18585 DVSS.n3470 DVSS.n2715 0.00803521
R18586 DVSS.n3469 DVSS.n2717 0.00803521
R18587 DVSS.n3466 DVSS.n3465 0.00803521
R18588 DVSS.n3065 DVSS.n2725 0.00803521
R18589 DVSS.n3071 DVSS.n3070 0.00803521
R18590 DVSS.n3454 DVSS.n2735 0.00803521
R18591 DVSS.n3453 DVSS.n2737 0.00803521
R18592 DVSS.n3450 DVSS.n3449 0.00803521
R18593 DVSS.n3082 DVSS.n2743 0.00803521
R18594 DVSS.n3442 DVSS.n2750 0.00803521
R18595 DVSS.n3441 DVSS.n2752 0.00803521
R18596 DVSS.n3438 DVSS.n3437 0.00803521
R18597 DVSS.n3095 DVSS.n2760 0.00803521
R18598 DVSS.n3430 DVSS.n2770 0.00803521
R18599 DVSS.n3429 DVSS.n2772 0.00803521
R18600 DVSS.n3426 DVSS.n3425 0.00803521
R18601 DVSS.n3106 DVSS.n2780 0.00803521
R18602 DVSS.n3418 DVSS.n2787 0.00803521
R18603 DVSS.n3417 DVSS.n2789 0.00803521
R18604 DVSS.n3414 DVSS.n3413 0.00803521
R18605 DVSS.n3119 DVSS.n2797 0.00803521
R18606 DVSS.n3406 DVSS.n2806 0.00803521
R18607 DVSS.n3405 DVSS.n2808 0.00803521
R18608 DVSS.n3402 DVSS.n3401 0.00803521
R18609 DVSS.n3134 DVSS.n2816 0.00803521
R18610 DVSS.n3140 DVSS.n3139 0.00803521
R18611 DVSS.n3390 DVSS.n2827 0.00803521
R18612 DVSS.n3389 DVSS.n2829 0.00803521
R18613 DVSS.n3386 DVSS.n3385 0.00803521
R18614 DVSS.n3151 DVSS.n2835 0.00803521
R18615 DVSS.n3378 DVSS.n2842 0.00803521
R18616 DVSS.n3377 DVSS.n2844 0.00803521
R18617 DVSS.n3374 DVSS.n3373 0.00803521
R18618 DVSS.n3164 DVSS.n2852 0.00803521
R18619 DVSS.n3366 DVSS.n2862 0.00803521
R18620 DVSS.n3365 DVSS.n2864 0.00803521
R18621 DVSS.n3362 DVSS.n3361 0.00803521
R18622 DVSS.n3176 DVSS.n2872 0.00803521
R18623 DVSS.n3354 DVSS.n2880 0.00803521
R18624 DVSS.n3353 DVSS.n2882 0.00803521
R18625 DVSS.n3350 DVSS.n3349 0.00803521
R18626 DVSS.n3188 DVSS.n2890 0.00803521
R18627 DVSS.n3341 DVSS.n2898 0.00803521
R18628 DVSS.n3340 DVSS.n2900 0.00803521
R18629 DVSS.n3337 DVSS.n3336 0.00803521
R18630 DVSS.n3199 DVSS.n2908 0.00803521
R18631 DVSS.n3328 DVSS.n2916 0.00803521
R18632 DVSS.n3327 DVSS.n2918 0.00803521
R18633 DVSS.n3324 DVSS.n3323 0.00803521
R18634 DVSS.n3212 DVSS.n2926 0.00803521
R18635 DVSS.n3316 DVSS.n2933 0.00803521
R18636 DVSS.n3315 DVSS.n2935 0.00803521
R18637 DVSS.n3312 DVSS.n3311 0.00803521
R18638 DVSS.n3225 DVSS.n2943 0.00803521
R18639 DVSS.n3303 DVSS.n2952 0.00803521
R18640 DVSS.n3302 DVSS.n2954 0.00803521
R18641 DVSS.n3299 DVSS.n3298 0.00803521
R18642 DVSS.n3236 DVSS.n2962 0.00803521
R18643 DVSS.n3290 DVSS.n2969 0.00803521
R18644 DVSS.n3289 DVSS.n2971 0.00803521
R18645 DVSS.n3286 DVSS.n3285 0.00803521
R18646 DVSS.n3247 DVSS.n2979 0.00803521
R18647 DVSS.n3278 DVSS.n2987 0.00803521
R18648 DVSS.n3277 DVSS.n2989 0.00803521
R18649 DVSS.n3274 DVSS.n3273 0.00803521
R18650 DVSS.n3263 DVSS.n2998 0.00803521
R18651 DVSS.n3262 DVSS.n1787 0.00803521
R18652 DVSS.n3830 DVSS.n3829 0.00803521
R18653 DVSS.n3420 DVSS.n2783 0.008
R18654 DVSS.n3348 DVSS.n2891 0.008
R18655 DVSS.n3108 DVSS.n3107 0.008
R18656 DVSS.n3184 DVSS.n2889 0.008
R18657 DVSS.n4878 DVSS.n1193 0.00789286
R18658 DVSS.n4888 DVSS.n1199 0.00789286
R18659 DVSS.n3759 DVSS.n3749 0.00789286
R18660 DVSS.n3762 DVSS.n3761 0.00789286
R18661 DVSS.n5532 DVSS 0.00782857
R18662 DVSS.n5531 DVSS 0.00782857
R18663 DVSS.n4690 DVSS 0.00782857
R18664 DVSS.n3748 VSS 0.00782857
R18665 DVSS DVSS.n2407 0.00782857
R18666 DVSS.n2094 DVSS 0.00782857
R18667 DVSS.n2093 DVSS 0.00782857
R18668 DVSS.n2411 DVSS 0.00782857
R18669 DVSS DVSS.n1761 0.00782857
R18670 DVSS DVSS.n1760 0.00782857
R18671 VSS DVSS.n1194 0.00782857
R18672 DVSS.n3953 DVSS.n3952 0.00776429
R18673 DVSS.n4624 DVSS.n4608 0.00761735
R18674 DVSS.n4718 DVSS.n4626 0.00761735
R18675 DVSS.n4587 DVSS.n1395 0.00761735
R18676 DVSS.n4752 DVSS.n1396 0.00761735
R18677 DVSS.n4551 DVSS.n4549 0.00761735
R18678 DVSS.n4566 DVSS.n1418 0.00761735
R18679 DVSS.n4512 DVSS.n1448 0.00761735
R18680 DVSS.n4526 DVSS.n1439 0.00761735
R18681 DVSS.n4431 DVSS.n4415 0.00761735
R18682 DVSS.n4470 DVSS.n4433 0.00761735
R18683 DVSS.n4394 DVSS.n4324 0.00761735
R18684 DVSS.n4504 DVSS.n4325 0.00761735
R18685 DVSS.n3281 DVSS.n2985 0.0075936
R18686 DVSS.n3251 DVSS.n3250 0.0075936
R18687 DVSS.n4485 DVSS.n4484 0.00757143
R18688 DVSS.n4481 DVSS.n4414 0.00757143
R18689 DVSS.n4480 DVSS.n4417 0.00757143
R18690 DVSS.n4424 DVSS.n4423 0.00757143
R18691 DVSS.n4474 DVSS.n4473 0.00757143
R18692 DVSS.n4434 DVSS.n4425 0.00757143
R18693 DVSS.n4468 DVSS.n4435 0.00757143
R18694 DVSS.n2264 DVSS.n2257 0.00757143
R18695 DVSS.n2261 DVSS.n1902 0.00757143
R18696 DVSS.n4452 DVSS.n4446 0.00750714
R18697 DVSS.n4449 DVSS.n4448 0.00750714
R18698 DVSS.n4516 DVSS.n1446 0.00750714
R18699 DVSS.n4515 DVSS.n1441 0.00750714
R18700 DVSS.n4523 DVSS.n4522 0.00750714
R18701 DVSS.n1442 DVSS.n1437 0.00750714
R18702 DVSS.n4529 DVSS.n4528 0.00750714
R18703 DVSS.n4708 DVSS.n4707 0.00750714
R18704 DVSS.n4662 DVSS.n4640 0.00750714
R18705 DVSS.n4704 DVSS.n4663 0.00750714
R18706 DVSS.n1913 DVSS.n1912 0.00750714
R18707 DVSS.n2532 DVSS.n2531 0.00750714
R18708 DVSS.n3400 DVSS.n3399 0.0075
R18709 DVSS.n3371 DVSS.n2854 0.0075
R18710 DVSS.n3015 DVSS.n2815 0.0075
R18711 DVSS.n3165 DVSS.n3163 0.0075
R18712 DVSS.n1385 DVSS.n1360 0.00745122
R18713 DVSS.n1375 DVSS.n1363 0.00745122
R18714 DVSS.n2502 DVSS.n2501 0.00739189
R18715 DVSS.n2499 DVSS.n2473 0.00739189
R18716 DVSS.n4623 DVSS.n4622 0.00730488
R18717 DVSS.n4622 DVSS.n4619 0.00730488
R18718 DVSS.n4589 DVSS.n1397 0.00730488
R18719 DVSS.n4751 DVSS.n1397 0.00730488
R18720 DVSS.n4553 DVSS.n4552 0.00730488
R18721 DVSS.n4553 DVSS.n1419 0.00730488
R18722 DVSS.n4514 DVSS.n4513 0.00730488
R18723 DVSS.n4514 DVSS.n1440 0.00730488
R18724 DVSS.n4430 DVSS.n4429 0.00730488
R18725 DVSS.n4429 DVSS.n4426 0.00730488
R18726 DVSS.n4396 DVSS.n4326 0.00730488
R18727 DVSS.n4503 DVSS.n4326 0.00730488
R18728 DVSS.n2685 DVSS.n2684 0.00716667
R18729 DVSS.n2686 DVSS.n2685 0.00716667
R18730 DVSS.n2687 DVSS.n2686 0.00716667
R18731 DVSS.n2701 DVSS.n2687 0.00716667
R18732 DVSS.n2702 DVSS.n2701 0.00716667
R18733 DVSS.n2703 DVSS.n2702 0.00716667
R18734 DVSS.n2704 DVSS.n2703 0.00716667
R18735 DVSS.n2719 DVSS.n2704 0.00716667
R18736 DVSS.n2720 DVSS.n2719 0.00716667
R18737 DVSS.n2721 DVSS.n2720 0.00716667
R18738 DVSS.n2722 DVSS.n2721 0.00716667
R18739 DVSS.n3066 DVSS.n2722 0.00716667
R18740 DVSS.n3068 DVSS.n3066 0.00716667
R18741 DVSS.n3068 DVSS.n3067 0.00716667
R18742 DVSS.n3067 DVSS.n2739 0.00716667
R18743 DVSS.n2740 DVSS.n2739 0.00716667
R18744 DVSS.n2754 DVSS.n2740 0.00716667
R18745 DVSS.n2755 DVSS.n2754 0.00716667
R18746 DVSS.n2756 DVSS.n2755 0.00716667
R18747 DVSS.n2757 DVSS.n2756 0.00716667
R18748 DVSS.n2774 DVSS.n2757 0.00716667
R18749 DVSS.n2775 DVSS.n2774 0.00716667
R18750 DVSS.n2776 DVSS.n2775 0.00716667
R18751 DVSS.n2777 DVSS.n2776 0.00716667
R18752 DVSS.n2791 DVSS.n2777 0.00716667
R18753 DVSS.n2792 DVSS.n2791 0.00716667
R18754 DVSS.n2793 DVSS.n2792 0.00716667
R18755 DVSS.n2794 DVSS.n2793 0.00716667
R18756 DVSS.n2810 DVSS.n2794 0.00716667
R18757 DVSS.n2811 DVSS.n2810 0.00716667
R18758 DVSS.n2812 DVSS.n2811 0.00716667
R18759 DVSS.n2813 DVSS.n2812 0.00716667
R18760 DVSS.n3135 DVSS.n2813 0.00716667
R18761 DVSS.n3137 DVSS.n3135 0.00716667
R18762 DVSS.n3137 DVSS.n3136 0.00716667
R18763 DVSS.n3136 DVSS.n2831 0.00716667
R18764 DVSS.n2832 DVSS.n2831 0.00716667
R18765 DVSS.n2846 DVSS.n2832 0.00716667
R18766 DVSS.n2847 DVSS.n2846 0.00716667
R18767 DVSS.n2848 DVSS.n2847 0.00716667
R18768 DVSS.n2849 DVSS.n2848 0.00716667
R18769 DVSS.n2866 DVSS.n2849 0.00716667
R18770 DVSS.n2867 DVSS.n2866 0.00716667
R18771 DVSS.n2868 DVSS.n2867 0.00716667
R18772 DVSS.n2869 DVSS.n2868 0.00716667
R18773 DVSS.n2884 DVSS.n2869 0.00716667
R18774 DVSS.n2885 DVSS.n2884 0.00716667
R18775 DVSS.n2886 DVSS.n2885 0.00716667
R18776 DVSS.n2887 DVSS.n2886 0.00716667
R18777 DVSS.n2902 DVSS.n2887 0.00716667
R18778 DVSS.n2903 DVSS.n2902 0.00716667
R18779 DVSS.n2904 DVSS.n2903 0.00716667
R18780 DVSS.n2905 DVSS.n2904 0.00716667
R18781 DVSS.n2920 DVSS.n2905 0.00716667
R18782 DVSS.n2921 DVSS.n2920 0.00716667
R18783 DVSS.n2922 DVSS.n2921 0.00716667
R18784 DVSS.n2923 DVSS.n2922 0.00716667
R18785 DVSS.n2937 DVSS.n2923 0.00716667
R18786 DVSS.n2938 DVSS.n2937 0.00716667
R18787 DVSS.n2939 DVSS.n2938 0.00716667
R18788 DVSS.n2940 DVSS.n2939 0.00716667
R18789 DVSS.n2956 DVSS.n2940 0.00716667
R18790 DVSS.n2957 DVSS.n2956 0.00716667
R18791 DVSS.n2958 DVSS.n2957 0.00716667
R18792 DVSS.n2959 DVSS.n2958 0.00716667
R18793 DVSS.n2973 DVSS.n2959 0.00716667
R18794 DVSS.n2974 DVSS.n2973 0.00716667
R18795 DVSS.n2975 DVSS.n2974 0.00716667
R18796 DVSS.n2976 DVSS.n2975 0.00716667
R18797 DVSS.n2991 DVSS.n2976 0.00716667
R18798 DVSS.n2992 DVSS.n2991 0.00716667
R18799 DVSS.n2993 DVSS.n2992 0.00716667
R18800 DVSS.n2994 DVSS.n2993 0.00716667
R18801 DVSS.n2995 DVSS.n2994 0.00716667
R18802 DVSS.n2995 DVSS.n1785 0.00716667
R18803 DVSS.n3832 DVSS.n1785 0.00716667
R18804 DVSS.n3833 DVSS.n3832 0.00716667
R18805 DVSS.n3834 DVSS.n3833 0.00716667
R18806 DVSS.n3834 DVSS.n1781 0.00716667
R18807 DVSS.n3840 DVSS.n1781 0.00716667
R18808 DVSS.n3841 DVSS.n3840 0.00716667
R18809 DVSS.n3842 DVSS.n3841 0.00716667
R18810 DVSS.n3843 DVSS.n3842 0.00716667
R18811 DVSS.n3844 DVSS.n3843 0.00716667
R18812 DVSS.n3847 DVSS.n3844 0.00716667
R18813 DVSS.n3848 DVSS.n3847 0.00716667
R18814 DVSS.n3849 DVSS.n3848 0.00716667
R18815 DVSS.n3850 DVSS.n3849 0.00716667
R18816 DVSS.n3851 DVSS.n3850 0.00716667
R18817 DVSS.n955 DVSS.n951 0.00712143
R18818 DVSS.n5346 DVSS.n5345 0.00712143
R18819 DVSS.n4770 DVSS.n1358 0.00712143
R18820 DVSS.n4688 DVSS.n1354 0.00712143
R18821 DVSS.n4048 DVSS.n4047 0.00712143
R18822 DVSS.n4001 DVSS.n1657 0.00705714
R18823 DVSS.n1662 DVSS.n1661 0.00705714
R18824 DVSS.n3995 DVSS.n3994 0.00705714
R18825 DVSS.n802 DVSS.n800 0.00700873
R18826 DVSS.n3392 DVSS.n3391 0.007
R18827 DVSS.n3379 DVSS.n2841 0.007
R18828 DVSS.n3142 DVSS.n2828 0.007
R18829 DVSS.n3156 DVSS.n2843 0.007
R18830 DVSS.n4041 DVSS.n4040 0.00699286
R18831 DVSS.n4028 DVSS.n1642 0.00699286
R18832 DVSS.n4060 DVSS.n4059 0.00692857
R18833 DVSS.n2556 DVSS.n2555 0.006875
R18834 DVSS.n2553 DVSS.n1911 0.006875
R18835 DVSS.n2565 DVSS.n1899 0.006875
R18836 DVSS.n2568 DVSS.n2567 0.006875
R18837 DVSS.n4537 DVSS.n1429 0.0068
R18838 DVSS.n4546 DVSS.n4544 0.0068
R18839 DVSS.n4545 DVSS.n1426 0.0068
R18840 DVSS.n4555 DVSS.n4554 0.0068
R18841 DVSS.n4563 DVSS.n1420 0.0068
R18842 DVSS.n4562 DVSS.n1421 0.0068
R18843 DVSS.n4568 DVSS.n1416 0.0068
R18844 DVSS.n4967 DVSS.n1156 0.0068
R18845 DVSS.n4874 DVSS.n4872 0.0068
R18846 DVSS.n1383 DVSS.n1360 0.00671951
R18847 DVSS.n1377 DVSS.n1363 0.00671951
R18848 DVSS.n2763 DVSS.n2748 0.0067069
R18849 DVSS.n3088 DVSS.n3086 0.0067069
R18850 DVSS.n5349 DVSS.n949 0.00658571
R18851 DVSS.n5350 DVSS.n5349 0.00658571
R18852 DVSS.n5351 DVSS.n5350 0.00658571
R18853 DVSS.n5351 DVSS.n945 0.00658571
R18854 DVSS.n5357 DVSS.n945 0.00658571
R18855 DVSS.n5358 DVSS.n5357 0.00658571
R18856 DVSS.n5359 DVSS.n5358 0.00658571
R18857 DVSS.n5359 DVSS.n941 0.00658571
R18858 DVSS.n5365 DVSS.n941 0.00658571
R18859 DVSS.n5366 DVSS.n5365 0.00658571
R18860 DVSS.n5367 DVSS.n5366 0.00658571
R18861 DVSS.n5367 DVSS.n937 0.00658571
R18862 DVSS.n5373 DVSS.n937 0.00658571
R18863 DVSS.n5374 DVSS.n5373 0.00658571
R18864 DVSS.n5375 DVSS.n5374 0.00658571
R18865 DVSS.n5375 DVSS.n933 0.00658571
R18866 DVSS.n5381 DVSS.n933 0.00658571
R18867 DVSS.n5382 DVSS.n5381 0.00658571
R18868 DVSS.n5383 DVSS.n5382 0.00658571
R18869 DVSS.n5383 DVSS.n929 0.00658571
R18870 DVSS.n5389 DVSS.n929 0.00658571
R18871 DVSS.n5390 DVSS.n5389 0.00658571
R18872 DVSS.n5391 DVSS.n5390 0.00658571
R18873 DVSS.n5391 DVSS.n925 0.00658571
R18874 DVSS.n5397 DVSS.n925 0.00658571
R18875 DVSS.n5398 DVSS.n5397 0.00658571
R18876 DVSS.n5399 DVSS.n5398 0.00658571
R18877 DVSS.n5399 DVSS.n921 0.00658571
R18878 DVSS.n5405 DVSS.n921 0.00658571
R18879 DVSS.n5406 DVSS.n5405 0.00658571
R18880 DVSS.n5407 DVSS.n5406 0.00658571
R18881 DVSS.n5407 DVSS.n917 0.00658571
R18882 DVSS.n5413 DVSS.n917 0.00658571
R18883 DVSS.n5414 DVSS.n5413 0.00658571
R18884 DVSS.n5415 DVSS.n5414 0.00658571
R18885 DVSS.n5415 DVSS.n913 0.00658571
R18886 DVSS.n5421 DVSS.n913 0.00658571
R18887 DVSS.n5422 DVSS.n5421 0.00658571
R18888 DVSS.n5423 DVSS.n5422 0.00658571
R18889 DVSS.n5423 DVSS.n909 0.00658571
R18890 DVSS.n5429 DVSS.n909 0.00658571
R18891 DVSS.n5430 DVSS.n5429 0.00658571
R18892 DVSS.n5431 DVSS.n5430 0.00658571
R18893 DVSS.n5431 DVSS.n905 0.00658571
R18894 DVSS.n5437 DVSS.n905 0.00658571
R18895 DVSS.n5438 DVSS.n5437 0.00658571
R18896 DVSS.n5439 DVSS.n5438 0.00658571
R18897 DVSS.n5439 DVSS.n901 0.00658571
R18898 DVSS.n5445 DVSS.n901 0.00658571
R18899 DVSS.n5446 DVSS.n5445 0.00658571
R18900 DVSS.n5447 DVSS.n5446 0.00658571
R18901 DVSS.n5447 DVSS.n897 0.00658571
R18902 DVSS.n5453 DVSS.n897 0.00658571
R18903 DVSS.n5454 DVSS.n5453 0.00658571
R18904 DVSS.n5455 DVSS.n5454 0.00658571
R18905 DVSS.n5455 DVSS.n893 0.00658571
R18906 DVSS.n5461 DVSS.n893 0.00658571
R18907 DVSS.n5462 DVSS.n5461 0.00658571
R18908 DVSS.n5463 DVSS.n5462 0.00658571
R18909 DVSS.n5463 DVSS.n889 0.00658571
R18910 DVSS.n5469 DVSS.n889 0.00658571
R18911 DVSS.n5470 DVSS.n5469 0.00658571
R18912 DVSS.n5471 DVSS.n5470 0.00658571
R18913 DVSS.n5471 DVSS.n885 0.00658571
R18914 DVSS.n5477 DVSS.n885 0.00658571
R18915 DVSS.n5478 DVSS.n5477 0.00658571
R18916 DVSS.n5479 DVSS.n5478 0.00658571
R18917 DVSS.n5479 DVSS.n881 0.00658571
R18918 DVSS.n5485 DVSS.n881 0.00658571
R18919 DVSS.n5486 DVSS.n5485 0.00658571
R18920 DVSS.n5487 DVSS.n5486 0.00658571
R18921 DVSS.n5487 DVSS.n877 0.00658571
R18922 DVSS.n5493 DVSS.n877 0.00658571
R18923 DVSS.n5494 DVSS.n5493 0.00658571
R18924 DVSS.n5495 DVSS.n5494 0.00658571
R18925 DVSS.n5495 DVSS.n873 0.00658571
R18926 DVSS.n5501 DVSS.n873 0.00658571
R18927 DVSS.n5502 DVSS.n5501 0.00658571
R18928 DVSS.n5503 DVSS.n5502 0.00658571
R18929 DVSS.n5503 DVSS.n869 0.00658571
R18930 DVSS.n5509 DVSS.n869 0.00658571
R18931 DVSS.n5510 DVSS.n5509 0.00658571
R18932 DVSS.n5511 DVSS.n5510 0.00658571
R18933 DVSS.n5511 DVSS.n865 0.00658571
R18934 DVSS.n5517 DVSS.n865 0.00658571
R18935 DVSS.n5518 DVSS.n5517 0.00658571
R18936 DVSS.n5519 DVSS.n5518 0.00658571
R18937 DVSS.n5519 DVSS.n861 0.00658571
R18938 DVSS.n5525 DVSS.n861 0.00658571
R18939 DVSS.n5526 DVSS.n5525 0.00658571
R18940 DVSS.n5527 DVSS.n5526 0.00658571
R18941 DVSS.n5527 DVSS.n857 0.00658571
R18942 DVSS.n5533 DVSS.n857 0.00658571
R18943 DVSS.n4381 DVSS.n4380 0.00658571
R18944 DVSS.n4381 DVSS.n4339 0.00658571
R18945 DVSS.n4387 DVSS.n4339 0.00658571
R18946 DVSS.n4388 DVSS.n4387 0.00658571
R18947 DVSS.n4389 DVSS.n4388 0.00658571
R18948 DVSS.n4389 DVSS.n4332 0.00658571
R18949 DVSS.n4402 DVSS.n4332 0.00658571
R18950 DVSS.n4403 DVSS.n4402 0.00658571
R18951 DVSS.n4498 DVSS.n4403 0.00658571
R18952 DVSS.n4498 DVSS.n4497 0.00658571
R18953 DVSS.n4497 DVSS.n4496 0.00658571
R18954 DVSS.n4496 DVSS.n4404 0.00658571
R18955 DVSS.n4490 DVSS.n4404 0.00658571
R18956 DVSS.n4490 DVSS.n4489 0.00658571
R18957 DVSS.n4489 DVSS.n4488 0.00658571
R18958 DVSS.n4488 DVSS.n4412 0.00658571
R18959 DVSS.n4420 DVSS.n4412 0.00658571
R18960 DVSS.n4478 DVSS.n4420 0.00658571
R18961 DVSS.n4478 DVSS.n4477 0.00658571
R18962 DVSS.n4477 DVSS.n4476 0.00658571
R18963 DVSS.n4476 DVSS.n4421 0.00658571
R18964 DVSS.n4439 DVSS.n4421 0.00658571
R18965 DVSS.n4465 DVSS.n4439 0.00658571
R18966 DVSS.n4465 DVSS.n4464 0.00658571
R18967 DVSS.n4464 DVSS.n4463 0.00658571
R18968 DVSS.n4463 DVSS.n4440 0.00658571
R18969 DVSS.n4457 DVSS.n4440 0.00658571
R18970 DVSS.n4457 DVSS.n4456 0.00658571
R18971 DVSS.n4456 DVSS.n4455 0.00658571
R18972 DVSS.n4455 DVSS.n4444 0.00658571
R18973 DVSS.n4444 DVSS.n1444 0.00658571
R18974 DVSS.n4518 DVSS.n1444 0.00658571
R18975 DVSS.n4519 DVSS.n4518 0.00658571
R18976 DVSS.n4520 DVSS.n4519 0.00658571
R18977 DVSS.n4520 DVSS.n1435 0.00658571
R18978 DVSS.n4531 DVSS.n1435 0.00658571
R18979 DVSS.n4532 DVSS.n4531 0.00658571
R18980 DVSS.n4533 DVSS.n4532 0.00658571
R18981 DVSS.n4533 DVSS.n1431 0.00658571
R18982 DVSS.n4540 DVSS.n1431 0.00658571
R18983 DVSS.n4541 DVSS.n4540 0.00658571
R18984 DVSS.n4542 DVSS.n4541 0.00658571
R18985 DVSS.n4542 DVSS.n1424 0.00658571
R18986 DVSS.n4557 DVSS.n1424 0.00658571
R18987 DVSS.n4558 DVSS.n4557 0.00658571
R18988 DVSS.n4560 DVSS.n4558 0.00658571
R18989 DVSS.n4560 DVSS.n4559 0.00658571
R18990 DVSS.n4559 DVSS.n1414 0.00658571
R18991 DVSS.n4572 DVSS.n1414 0.00658571
R18992 DVSS.n4573 DVSS.n4572 0.00658571
R18993 DVSS.n4574 DVSS.n4573 0.00658571
R18994 DVSS.n4574 DVSS.n1410 0.00658571
R18995 DVSS.n4580 DVSS.n1410 0.00658571
R18996 DVSS.n4581 DVSS.n4580 0.00658571
R18997 DVSS.n4582 DVSS.n4581 0.00658571
R18998 DVSS.n4582 DVSS.n1403 0.00658571
R18999 DVSS.n4595 DVSS.n1403 0.00658571
R19000 DVSS.n4596 DVSS.n4595 0.00658571
R19001 DVSS.n4746 DVSS.n4596 0.00658571
R19002 DVSS.n4746 DVSS.n4745 0.00658571
R19003 DVSS.n4745 DVSS.n4744 0.00658571
R19004 DVSS.n4744 DVSS.n4597 0.00658571
R19005 DVSS.n4738 DVSS.n4597 0.00658571
R19006 DVSS.n4738 DVSS.n4737 0.00658571
R19007 DVSS.n4737 DVSS.n4736 0.00658571
R19008 DVSS.n4736 DVSS.n4605 0.00658571
R19009 DVSS.n4613 DVSS.n4605 0.00658571
R19010 DVSS.n4726 DVSS.n4613 0.00658571
R19011 DVSS.n4726 DVSS.n4725 0.00658571
R19012 DVSS.n4725 DVSS.n4724 0.00658571
R19013 DVSS.n4724 DVSS.n4614 0.00658571
R19014 DVSS.n4632 DVSS.n4614 0.00658571
R19015 DVSS.n4713 DVSS.n4632 0.00658571
R19016 DVSS.n4713 DVSS.n4712 0.00658571
R19017 DVSS.n4712 DVSS.n4711 0.00658571
R19018 DVSS.n4711 DVSS.n4633 0.00658571
R19019 DVSS.n4671 DVSS.n4633 0.00658571
R19020 DVSS.n4672 DVSS.n4671 0.00658571
R19021 DVSS.n4701 DVSS.n4672 0.00658571
R19022 DVSS.n4701 DVSS.n4700 0.00658571
R19023 DVSS.n4700 DVSS.n4699 0.00658571
R19024 DVSS.n4699 DVSS.n4673 0.00658571
R19025 DVSS.n4693 DVSS.n4673 0.00658571
R19026 DVSS.n4693 DVSS.n4692 0.00658571
R19027 DVSS.n4692 DVSS.n4691 0.00658571
R19028 DVSS.n4686 DVSS.n4685 0.00658571
R19029 DVSS.n1578 DVSS.n1569 0.00658571
R19030 DVSS.n1579 DVSS.n1578 0.00658571
R19031 DVSS.n1580 DVSS.n1579 0.00658571
R19032 DVSS.n1580 DVSS.n1565 0.00658571
R19033 DVSS.n1586 DVSS.n1565 0.00658571
R19034 DVSS.n1587 DVSS.n1586 0.00658571
R19035 DVSS.n1588 DVSS.n1587 0.00658571
R19036 DVSS.n1588 DVSS.n1561 0.00658571
R19037 DVSS.n1594 DVSS.n1561 0.00658571
R19038 DVSS.n1595 DVSS.n1594 0.00658571
R19039 DVSS.n4088 DVSS.n1595 0.00658571
R19040 DVSS.n4088 DVSS.n4087 0.00658571
R19041 DVSS.n4087 DVSS.n4086 0.00658571
R19042 DVSS.n4086 DVSS.n1596 0.00658571
R19043 DVSS.n4080 DVSS.n1596 0.00658571
R19044 DVSS.n4080 DVSS.n4079 0.00658571
R19045 DVSS.n4079 DVSS.n4078 0.00658571
R19046 DVSS.n4078 DVSS.n1600 0.00658571
R19047 DVSS.n4072 DVSS.n1600 0.00658571
R19048 DVSS.n4072 DVSS.n4071 0.00658571
R19049 DVSS.n4071 DVSS.n4070 0.00658571
R19050 DVSS.n4070 DVSS.n1604 0.00658571
R19051 DVSS.n4064 DVSS.n1604 0.00658571
R19052 DVSS.n4064 DVSS.n4063 0.00658571
R19053 DVSS.n4063 DVSS.n4062 0.00658571
R19054 DVSS.n4062 DVSS.n1608 0.00658571
R19055 DVSS.n3608 DVSS.n1608 0.00658571
R19056 DVSS.n3609 DVSS.n3608 0.00658571
R19057 DVSS.n3609 DVSS.n3604 0.00658571
R19058 DVSS.n3615 DVSS.n3604 0.00658571
R19059 DVSS.n3616 DVSS.n3615 0.00658571
R19060 DVSS.n3617 DVSS.n3616 0.00658571
R19061 DVSS.n3617 DVSS.n3600 0.00658571
R19062 DVSS.n3623 DVSS.n3600 0.00658571
R19063 DVSS.n3624 DVSS.n3623 0.00658571
R19064 DVSS.n3625 DVSS.n3624 0.00658571
R19065 DVSS.n3625 DVSS.n3596 0.00658571
R19066 DVSS.n3631 DVSS.n3596 0.00658571
R19067 DVSS.n3632 DVSS.n3631 0.00658571
R19068 DVSS.n3633 DVSS.n3632 0.00658571
R19069 DVSS.n3633 DVSS.n3592 0.00658571
R19070 DVSS.n3639 DVSS.n3592 0.00658571
R19071 DVSS.n3640 DVSS.n3639 0.00658571
R19072 DVSS.n3641 DVSS.n3640 0.00658571
R19073 DVSS.n3641 DVSS.n3588 0.00658571
R19074 DVSS.n3647 DVSS.n3588 0.00658571
R19075 DVSS.n3648 DVSS.n3647 0.00658571
R19076 DVSS.n3649 DVSS.n3648 0.00658571
R19077 DVSS.n3649 DVSS.n3584 0.00658571
R19078 DVSS.n3655 DVSS.n3584 0.00658571
R19079 DVSS.n3656 DVSS.n3655 0.00658571
R19080 DVSS.n3657 DVSS.n3656 0.00658571
R19081 DVSS.n3657 DVSS.n3580 0.00658571
R19082 DVSS.n3663 DVSS.n3580 0.00658571
R19083 DVSS.n3664 DVSS.n3663 0.00658571
R19084 DVSS.n3665 DVSS.n3664 0.00658571
R19085 DVSS.n3665 DVSS.n3576 0.00658571
R19086 DVSS.n3671 DVSS.n3576 0.00658571
R19087 DVSS.n3672 DVSS.n3671 0.00658571
R19088 DVSS.n3673 DVSS.n3672 0.00658571
R19089 DVSS.n3673 DVSS.n3572 0.00658571
R19090 DVSS.n3679 DVSS.n3572 0.00658571
R19091 DVSS.n3680 DVSS.n3679 0.00658571
R19092 DVSS.n3681 DVSS.n3680 0.00658571
R19093 DVSS.n3681 DVSS.n3568 0.00658571
R19094 DVSS.n3687 DVSS.n3568 0.00658571
R19095 DVSS.n3688 DVSS.n3687 0.00658571
R19096 DVSS.n3689 DVSS.n3688 0.00658571
R19097 DVSS.n3689 DVSS.n3564 0.00658571
R19098 DVSS.n3695 DVSS.n3564 0.00658571
R19099 DVSS.n3696 DVSS.n3695 0.00658571
R19100 DVSS.n3697 DVSS.n3696 0.00658571
R19101 DVSS.n3697 DVSS.n3560 0.00658571
R19102 DVSS.n3703 DVSS.n3560 0.00658571
R19103 DVSS.n3704 DVSS.n3703 0.00658571
R19104 DVSS.n3705 DVSS.n3704 0.00658571
R19105 DVSS.n3705 DVSS.n3556 0.00658571
R19106 DVSS.n3711 DVSS.n3556 0.00658571
R19107 DVSS.n3712 DVSS.n3711 0.00658571
R19108 DVSS.n3713 DVSS.n3712 0.00658571
R19109 DVSS.n3713 DVSS.n3552 0.00658571
R19110 DVSS.n3719 DVSS.n3552 0.00658571
R19111 DVSS.n3720 DVSS.n3719 0.00658571
R19112 DVSS.n3721 DVSS.n3720 0.00658571
R19113 DVSS.n3721 DVSS.n3548 0.00658571
R19114 DVSS.n3727 DVSS.n3548 0.00658571
R19115 DVSS.n3728 DVSS.n3727 0.00658571
R19116 DVSS.n3729 DVSS.n3728 0.00658571
R19117 DVSS.n3729 DVSS.n3544 0.00658571
R19118 DVSS.n3735 DVSS.n3544 0.00658571
R19119 DVSS.n3736 DVSS.n3735 0.00658571
R19120 DVSS.n3737 DVSS.n3736 0.00658571
R19121 DVSS.n3737 DVSS.n3540 0.00658571
R19122 DVSS.n3743 DVSS.n3540 0.00658571
R19123 DVSS.n3744 DVSS.n3743 0.00658571
R19124 DVSS.n3747 DVSS.n3744 0.00658571
R19125 DVSS.n3747 DVSS.n3746 0.00658571
R19126 DVSS.n3765 DVSS.n3525 0.00658571
R19127 DVSS.n2611 DVSS.n2610 0.00658571
R19128 DVSS.n2610 DVSS.n2609 0.00658571
R19129 DVSS.n2609 DVSS.n1852 0.00658571
R19130 DVSS.n2603 DVSS.n1852 0.00658571
R19131 DVSS.n2603 DVSS.n2602 0.00658571
R19132 DVSS.n2602 DVSS.n2601 0.00658571
R19133 DVSS.n2601 DVSS.n1857 0.00658571
R19134 DVSS.n2282 DVSS.n1857 0.00658571
R19135 DVSS.n2283 DVSS.n2282 0.00658571
R19136 DVSS.n2283 DVSS.n2273 0.00658571
R19137 DVSS.n2291 DVSS.n2273 0.00658571
R19138 DVSS.n2292 DVSS.n2291 0.00658571
R19139 DVSS.n2293 DVSS.n2292 0.00658571
R19140 DVSS.n2293 DVSS.n1881 0.00658571
R19141 DVSS.n2580 DVSS.n1881 0.00658571
R19142 DVSS.n2580 DVSS.n2579 0.00658571
R19143 DVSS.n2579 DVSS.n2578 0.00658571
R19144 DVSS.n2578 DVSS.n1882 0.00658571
R19145 DVSS.n2258 DVSS.n1882 0.00658571
R19146 DVSS.n2258 DVSS.n1908 0.00658571
R19147 DVSS.n2562 DVSS.n1908 0.00658571
R19148 DVSS.n2562 DVSS.n2561 0.00658571
R19149 DVSS.n2561 DVSS.n2560 0.00658571
R19150 DVSS.n2560 DVSS.n1909 0.00658571
R19151 DVSS.n2529 DVSS.n1909 0.00658571
R19152 DVSS.n2529 DVSS.n2528 0.00658571
R19153 DVSS.n2528 DVSS.n2527 0.00658571
R19154 DVSS.n2527 DVSS.n2315 0.00658571
R19155 DVSS.n2356 DVSS.n2315 0.00658571
R19156 DVSS.n2357 DVSS.n2356 0.00658571
R19157 DVSS.n2358 DVSS.n2357 0.00658571
R19158 DVSS.n2358 DVSS.n2343 0.00658571
R19159 DVSS.n2374 DVSS.n2343 0.00658571
R19160 DVSS.n2375 DVSS.n2374 0.00658571
R19161 DVSS.n2508 DVSS.n2375 0.00658571
R19162 DVSS.n2508 DVSS.n2507 0.00658571
R19163 DVSS.n2507 DVSS.n2506 0.00658571
R19164 DVSS.n2506 DVSS.n2376 0.00658571
R19165 DVSS.n2378 DVSS.n2376 0.00658571
R19166 DVSS.n2381 DVSS.n2378 0.00658571
R19167 DVSS.n2464 DVSS.n2381 0.00658571
R19168 DVSS.n2464 DVSS.n2463 0.00658571
R19169 DVSS.n2463 DVSS.n2462 0.00658571
R19170 DVSS.n2462 DVSS.n2382 0.00658571
R19171 DVSS.n2456 DVSS.n2382 0.00658571
R19172 DVSS.n2456 DVSS.n2455 0.00658571
R19173 DVSS.n2455 DVSS.n2454 0.00658571
R19174 DVSS.n2454 DVSS.n2386 0.00658571
R19175 DVSS.n2448 DVSS.n2386 0.00658571
R19176 DVSS.n2448 DVSS.n2447 0.00658571
R19177 DVSS.n2447 DVSS.n2446 0.00658571
R19178 DVSS.n2446 DVSS.n2390 0.00658571
R19179 DVSS.n2440 DVSS.n2390 0.00658571
R19180 DVSS.n2440 DVSS.n2439 0.00658571
R19181 DVSS.n2439 DVSS.n2438 0.00658571
R19182 DVSS.n2438 DVSS.n2394 0.00658571
R19183 DVSS.n2432 DVSS.n2394 0.00658571
R19184 DVSS.n2432 DVSS.n2431 0.00658571
R19185 DVSS.n2431 DVSS.n2430 0.00658571
R19186 DVSS.n2430 DVSS.n2398 0.00658571
R19187 DVSS.n2424 DVSS.n2398 0.00658571
R19188 DVSS.n2424 DVSS.n2423 0.00658571
R19189 DVSS.n2423 DVSS.n2422 0.00658571
R19190 DVSS.n2422 DVSS.n2402 0.00658571
R19191 DVSS.n2416 DVSS.n2402 0.00658571
R19192 DVSS.n2416 DVSS.n2415 0.00658571
R19193 DVSS.n2415 DVSS.n2414 0.00658571
R19194 DVSS.n2414 DVSS.n2406 0.00658571
R19195 DVSS.n2408 DVSS.n2406 0.00658571
R19196 DVSS.n2019 DVSS.n1967 0.00658571
R19197 DVSS.n2025 DVSS.n1967 0.00658571
R19198 DVSS.n2026 DVSS.n2025 0.00658571
R19199 DVSS.n2224 DVSS.n2026 0.00658571
R19200 DVSS.n2224 DVSS.n2223 0.00658571
R19201 DVSS.n2223 DVSS.n2222 0.00658571
R19202 DVSS.n2222 DVSS.n2027 0.00658571
R19203 DVSS.n2216 DVSS.n2027 0.00658571
R19204 DVSS.n2216 DVSS.n2215 0.00658571
R19205 DVSS.n2215 DVSS.n2214 0.00658571
R19206 DVSS.n2214 DVSS.n2031 0.00658571
R19207 DVSS.n2208 DVSS.n2031 0.00658571
R19208 DVSS.n2208 DVSS.n2207 0.00658571
R19209 DVSS.n2207 DVSS.n2206 0.00658571
R19210 DVSS.n2206 DVSS.n2035 0.00658571
R19211 DVSS.n2200 DVSS.n2035 0.00658571
R19212 DVSS.n2200 DVSS.n2199 0.00658571
R19213 DVSS.n2199 DVSS.n2198 0.00658571
R19214 DVSS.n2198 DVSS.n2039 0.00658571
R19215 DVSS.n2192 DVSS.n2039 0.00658571
R19216 DVSS.n2192 DVSS.n2191 0.00658571
R19217 DVSS.n2191 DVSS.n2190 0.00658571
R19218 DVSS.n2190 DVSS.n2043 0.00658571
R19219 DVSS.n2184 DVSS.n2043 0.00658571
R19220 DVSS.n2184 DVSS.n2183 0.00658571
R19221 DVSS.n2183 DVSS.n2182 0.00658571
R19222 DVSS.n2182 DVSS.n2047 0.00658571
R19223 DVSS.n2176 DVSS.n2047 0.00658571
R19224 DVSS.n2176 DVSS.n2175 0.00658571
R19225 DVSS.n2175 DVSS.n2174 0.00658571
R19226 DVSS.n2174 DVSS.n2051 0.00658571
R19227 DVSS.n2168 DVSS.n2051 0.00658571
R19228 DVSS.n2168 DVSS.n2167 0.00658571
R19229 DVSS.n2167 DVSS.n2166 0.00658571
R19230 DVSS.n2166 DVSS.n2055 0.00658571
R19231 DVSS.n2160 DVSS.n2055 0.00658571
R19232 DVSS.n2160 DVSS.n2159 0.00658571
R19233 DVSS.n2159 DVSS.n2158 0.00658571
R19234 DVSS.n2158 DVSS.n2059 0.00658571
R19235 DVSS.n2152 DVSS.n2059 0.00658571
R19236 DVSS.n2152 DVSS.n2151 0.00658571
R19237 DVSS.n2151 DVSS.n2150 0.00658571
R19238 DVSS.n2150 DVSS.n2063 0.00658571
R19239 DVSS.n2145 DVSS.n2063 0.00658571
R19240 DVSS.n2145 DVSS.n2144 0.00658571
R19241 DVSS.n2144 DVSS.n2143 0.00658571
R19242 DVSS.n2143 DVSS.n2065 0.00658571
R19243 DVSS.n2137 DVSS.n2065 0.00658571
R19244 DVSS.n2137 DVSS.n2136 0.00658571
R19245 DVSS.n2136 DVSS.n2135 0.00658571
R19246 DVSS.n2135 DVSS.n2070 0.00658571
R19247 DVSS.n2129 DVSS.n2070 0.00658571
R19248 DVSS.n2129 DVSS.n2128 0.00658571
R19249 DVSS.n2128 DVSS.n2127 0.00658571
R19250 DVSS.n2127 DVSS.n2074 0.00658571
R19251 DVSS.n2121 DVSS.n2074 0.00658571
R19252 DVSS.n2121 DVSS.n2120 0.00658571
R19253 DVSS.n2120 DVSS.n2119 0.00658571
R19254 DVSS.n2119 DVSS.n2078 0.00658571
R19255 DVSS.n2113 DVSS.n2078 0.00658571
R19256 DVSS.n2113 DVSS.n2112 0.00658571
R19257 DVSS.n2112 DVSS.n2111 0.00658571
R19258 DVSS.n2111 DVSS.n2082 0.00658571
R19259 DVSS.n2105 DVSS.n2082 0.00658571
R19260 DVSS.n2105 DVSS.n2104 0.00658571
R19261 DVSS.n2104 DVSS.n2103 0.00658571
R19262 DVSS.n2103 DVSS.n2086 0.00658571
R19263 DVSS.n2097 DVSS.n2086 0.00658571
R19264 DVSS.n2097 DVSS.n2096 0.00658571
R19265 DVSS.n2096 DVSS.n2095 0.00658571
R19266 DVSS.n2095 DVSS.n2090 0.00658571
R19267 DVSS.n4045 DVSS.n1635 0.00658571
R19268 DVSS.n4045 DVSS.n4044 0.00658571
R19269 DVSS.n4044 DVSS.n4043 0.00658571
R19270 DVSS.n4043 DVSS.n1636 0.00658571
R19271 DVSS.n4036 DVSS.n1636 0.00658571
R19272 DVSS.n4036 DVSS.n4035 0.00658571
R19273 DVSS.n4035 DVSS.n4034 0.00658571
R19274 DVSS.n4034 DVSS.n1640 0.00658571
R19275 DVSS.n4026 DVSS.n1640 0.00658571
R19276 DVSS.n4026 DVSS.n4025 0.00658571
R19277 DVSS.n4025 DVSS.n4024 0.00658571
R19278 DVSS.n4024 DVSS.n1644 0.00658571
R19279 DVSS.n4018 DVSS.n1644 0.00658571
R19280 DVSS.n4018 DVSS.n4017 0.00658571
R19281 DVSS.n4017 DVSS.n4016 0.00658571
R19282 DVSS.n4016 DVSS.n1649 0.00658571
R19283 DVSS.n4007 DVSS.n1649 0.00658571
R19284 DVSS.n4007 DVSS.n4006 0.00658571
R19285 DVSS.n4006 DVSS.n4005 0.00658571
R19286 DVSS.n4005 DVSS.n1654 0.00658571
R19287 DVSS.n3999 DVSS.n1654 0.00658571
R19288 DVSS.n3999 DVSS.n3998 0.00658571
R19289 DVSS.n3998 DVSS.n3997 0.00658571
R19290 DVSS.n3997 DVSS.n1659 0.00658571
R19291 DVSS.n3979 DVSS.n1659 0.00658571
R19292 DVSS.n3979 DVSS.n3978 0.00658571
R19293 DVSS.n3978 DVSS.n3977 0.00658571
R19294 DVSS.n3977 DVSS.n1672 0.00658571
R19295 DVSS.n3971 DVSS.n1672 0.00658571
R19296 DVSS.n3971 DVSS.n3970 0.00658571
R19297 DVSS.n3970 DVSS.n3969 0.00658571
R19298 DVSS.n3969 DVSS.n1676 0.00658571
R19299 DVSS.n3963 DVSS.n1676 0.00658571
R19300 DVSS.n3963 DVSS.n3962 0.00658571
R19301 DVSS.n3962 DVSS.n3961 0.00658571
R19302 DVSS.n3961 DVSS.n1680 0.00658571
R19303 DVSS.n1691 DVSS.n1680 0.00658571
R19304 DVSS.n3950 DVSS.n1691 0.00658571
R19305 DVSS.n3950 DVSS.n3949 0.00658571
R19306 DVSS.n3949 DVSS.n3948 0.00658571
R19307 DVSS.n3948 DVSS.n1692 0.00658571
R19308 DVSS.n1711 DVSS.n1692 0.00658571
R19309 DVSS.n1716 DVSS.n1711 0.00658571
R19310 DVSS.n1717 DVSS.n1716 0.00658571
R19311 DVSS.n3927 DVSS.n1717 0.00658571
R19312 DVSS.n3927 DVSS.n3926 0.00658571
R19313 DVSS.n3926 DVSS.n3925 0.00658571
R19314 DVSS.n3925 DVSS.n1718 0.00658571
R19315 DVSS.n3919 DVSS.n1718 0.00658571
R19316 DVSS.n3919 DVSS.n3918 0.00658571
R19317 DVSS.n3918 DVSS.n3917 0.00658571
R19318 DVSS.n3917 DVSS.n1724 0.00658571
R19319 DVSS.n3911 DVSS.n1724 0.00658571
R19320 DVSS.n3911 DVSS.n3910 0.00658571
R19321 DVSS.n3910 DVSS.n3909 0.00658571
R19322 DVSS.n3909 DVSS.n1732 0.00658571
R19323 DVSS.n3903 DVSS.n1732 0.00658571
R19324 DVSS.n3903 DVSS.n3902 0.00658571
R19325 DVSS.n3902 DVSS.n3901 0.00658571
R19326 DVSS.n3901 DVSS.n1738 0.00658571
R19327 DVSS.n3895 DVSS.n1738 0.00658571
R19328 DVSS.n3895 DVSS.n3894 0.00658571
R19329 DVSS.n3894 DVSS.n3893 0.00658571
R19330 DVSS.n3893 DVSS.n1742 0.00658571
R19331 DVSS.n3887 DVSS.n1742 0.00658571
R19332 DVSS.n3887 DVSS.n3886 0.00658571
R19333 DVSS.n3886 DVSS.n3885 0.00658571
R19334 DVSS.n3885 DVSS.n1746 0.00658571
R19335 DVSS.n3879 DVSS.n1746 0.00658571
R19336 DVSS.n3879 DVSS.n3878 0.00658571
R19337 DVSS.n3878 DVSS.n3877 0.00658571
R19338 DVSS.n3877 DVSS.n1750 0.00658571
R19339 DVSS.n3871 DVSS.n1750 0.00658571
R19340 DVSS.n3871 DVSS.n3870 0.00658571
R19341 DVSS.n3870 DVSS.n3869 0.00658571
R19342 DVSS.n3869 DVSS.n1754 0.00658571
R19343 DVSS.n1774 DVSS.n1754 0.00658571
R19344 DVSS.n1774 DVSS.n1773 0.00658571
R19345 DVSS.n1773 DVSS.n1772 0.00658571
R19346 DVSS.n1772 DVSS.n1758 0.00658571
R19347 DVSS.n1766 DVSS.n1758 0.00658571
R19348 DVSS.n1766 DVSS.n1765 0.00658571
R19349 DVSS.n1765 DVSS.n1764 0.00658571
R19350 DVSS.n5090 DVSS.n1084 0.00658571
R19351 DVSS.n5084 DVSS.n1084 0.00658571
R19352 DVSS.n5084 DVSS.n5083 0.00658571
R19353 DVSS.n5083 DVSS.n5082 0.00658571
R19354 DVSS.n5082 DVSS.n1088 0.00658571
R19355 DVSS.n5076 DVSS.n1088 0.00658571
R19356 DVSS.n5076 DVSS.n5075 0.00658571
R19357 DVSS.n5075 DVSS.n5074 0.00658571
R19358 DVSS.n5074 DVSS.n1092 0.00658571
R19359 DVSS.n5068 DVSS.n1092 0.00658571
R19360 DVSS.n5068 DVSS.n5067 0.00658571
R19361 DVSS.n5067 DVSS.n5066 0.00658571
R19362 DVSS.n5066 DVSS.n1096 0.00658571
R19363 DVSS.n5059 DVSS.n1096 0.00658571
R19364 DVSS.n5059 DVSS.n5058 0.00658571
R19365 DVSS.n5058 DVSS.n5057 0.00658571
R19366 DVSS.n5057 DVSS.n1101 0.00658571
R19367 DVSS.n5051 DVSS.n1101 0.00658571
R19368 DVSS.n5051 DVSS.n5050 0.00658571
R19369 DVSS.n5050 DVSS.n5049 0.00658571
R19370 DVSS.n5049 DVSS.n1106 0.00658571
R19371 DVSS.n1113 DVSS.n1106 0.00658571
R19372 DVSS.n5040 DVSS.n1113 0.00658571
R19373 DVSS.n5040 DVSS.n5039 0.00658571
R19374 DVSS.n5039 DVSS.n5038 0.00658571
R19375 DVSS.n5038 DVSS.n1114 0.00658571
R19376 DVSS.n5029 DVSS.n1114 0.00658571
R19377 DVSS.n5029 DVSS.n5028 0.00658571
R19378 DVSS.n5028 DVSS.n5027 0.00658571
R19379 DVSS.n5027 DVSS.n1124 0.00658571
R19380 DVSS.n5021 DVSS.n1124 0.00658571
R19381 DVSS.n5021 DVSS.n5020 0.00658571
R19382 DVSS.n5020 DVSS.n5019 0.00658571
R19383 DVSS.n5019 DVSS.n1130 0.00658571
R19384 DVSS.n5013 DVSS.n1130 0.00658571
R19385 DVSS.n5013 DVSS.n5012 0.00658571
R19386 DVSS.n5012 DVSS.n5011 0.00658571
R19387 DVSS.n5011 DVSS.n1134 0.00658571
R19388 DVSS.n5005 DVSS.n1134 0.00658571
R19389 DVSS.n5005 DVSS.n5004 0.00658571
R19390 DVSS.n5004 DVSS.n5003 0.00658571
R19391 DVSS.n5003 DVSS.n1138 0.00658571
R19392 DVSS.n4997 DVSS.n1138 0.00658571
R19393 DVSS.n4997 DVSS.n4996 0.00658571
R19394 DVSS.n4996 DVSS.n4995 0.00658571
R19395 DVSS.n4995 DVSS.n1142 0.00658571
R19396 DVSS.n4989 DVSS.n1142 0.00658571
R19397 DVSS.n4989 DVSS.n4988 0.00658571
R19398 DVSS.n4988 DVSS.n4987 0.00658571
R19399 DVSS.n4987 DVSS.n1146 0.00658571
R19400 DVSS.n4981 DVSS.n1146 0.00658571
R19401 DVSS.n4981 DVSS.n4980 0.00658571
R19402 DVSS.n4980 DVSS.n4979 0.00658571
R19403 DVSS.n4979 DVSS.n1150 0.00658571
R19404 DVSS.n4973 DVSS.n1150 0.00658571
R19405 DVSS.n4973 DVSS.n4972 0.00658571
R19406 DVSS.n4972 DVSS.n4971 0.00658571
R19407 DVSS.n4971 DVSS.n1154 0.00658571
R19408 DVSS.n4965 DVSS.n1154 0.00658571
R19409 DVSS.n4965 DVSS.n4964 0.00658571
R19410 DVSS.n4964 DVSS.n4963 0.00658571
R19411 DVSS.n4963 DVSS.n1158 0.00658571
R19412 DVSS.n4957 DVSS.n1158 0.00658571
R19413 DVSS.n4957 DVSS.n4956 0.00658571
R19414 DVSS.n4956 DVSS.n4955 0.00658571
R19415 DVSS.n4955 DVSS.n1163 0.00658571
R19416 DVSS.n4949 DVSS.n1163 0.00658571
R19417 DVSS.n4949 DVSS.n4948 0.00658571
R19418 DVSS.n4948 DVSS.n4947 0.00658571
R19419 DVSS.n4947 DVSS.n1167 0.00658571
R19420 DVSS.n4941 DVSS.n1167 0.00658571
R19421 DVSS.n4941 DVSS.n4940 0.00658571
R19422 DVSS.n4940 DVSS.n4939 0.00658571
R19423 DVSS.n4939 DVSS.n1171 0.00658571
R19424 DVSS.n4933 DVSS.n1171 0.00658571
R19425 DVSS.n4933 DVSS.n4932 0.00658571
R19426 DVSS.n4932 DVSS.n4931 0.00658571
R19427 DVSS.n4931 DVSS.n1175 0.00658571
R19428 DVSS.n4925 DVSS.n1175 0.00658571
R19429 DVSS.n4925 DVSS.n4924 0.00658571
R19430 DVSS.n4924 DVSS.n4923 0.00658571
R19431 DVSS.n4923 DVSS.n1179 0.00658571
R19432 DVSS.n4917 DVSS.n1179 0.00658571
R19433 DVSS.n4917 DVSS.n4916 0.00658571
R19434 DVSS.n4916 DVSS.n4915 0.00658571
R19435 DVSS.n4915 DVSS.n1183 0.00658571
R19436 DVSS.n4909 DVSS.n1183 0.00658571
R19437 DVSS.n4909 DVSS.n4908 0.00658571
R19438 DVSS.n4908 DVSS.n4907 0.00658571
R19439 DVSS.n4907 DVSS.n1187 0.00658571
R19440 DVSS.n4901 DVSS.n1187 0.00658571
R19441 DVSS.n4901 DVSS.n4900 0.00658571
R19442 DVSS.n4900 DVSS.n4899 0.00658571
R19443 DVSS.n4899 DVSS.n1191 0.00658571
R19444 DVSS.n4893 DVSS.n1191 0.00658571
R19445 DVSS.n4893 DVSS.n4892 0.00658571
R19446 DVSS.n4892 DVSS.n4891 0.00658571
R19447 DVSS.n3519 DVSS.n3516 0.00658571
R19448 DVSS.n2487 DVSS.n1920 0.00658108
R19449 DVSS.n1944 DVSS.n1933 0.00658108
R19450 DVSS.n4392 DVSS.n4391 0.00654286
R19451 DVSS.n4337 DVSS.n4334 0.00654286
R19452 DVSS.n4400 DVSS.n4398 0.00654286
R19453 DVSS.n4399 DVSS.n4328 0.00654286
R19454 DVSS.n4501 DVSS.n4500 0.00654286
R19455 DVSS.n4406 DVSS.n4329 0.00654286
R19456 DVSS.n4494 DVSS.n4409 0.00654286
R19457 DVSS.n254 DVSS.n253 0.0065
R19458 DVSS.n611 DVSS.n185 0.0065
R19459 DVSS.n577 DVSS.n576 0.0065
R19460 DVSS.n716 DVSS.n715 0.0065
R19461 DVSS.n3412 DVSS.n2798 0.0065
R19462 DVSS.n3356 DVSS.n2875 0.0065
R19463 DVSS.n3114 DVSS.n2796 0.0065
R19464 DVSS.n3178 DVSS.n3177 0.0065
R19465 DVSS.n363 DVSS.n362 0.0065
R19466 DVSS.n577 DVSS.n184 0.0065
R19467 DVSS.n715 DVSS.n155 0.0065
R19468 DVSS.n5725 DVSS.n47 0.0065
R19469 DVSS.n5725 DVSS.n40 0.0065
R19470 DVSS.n364 DVSS.n363 0.0065
R19471 DVSS.n5568 DVSS.n46 0.0065
R19472 DVSS.n611 DVSS.n203 0.0065
R19473 DVSS.n253 DVSS.n250 0.0065
R19474 DVSS.n5650 DVSS.n133 0.0065
R19475 DVSS.n5651 DVSS.n5650 0.0065
R19476 DVSS.n46 DVSS.n41 0.0065
R19477 DVSS DVSS.n4686 0.00641429
R19478 VSS DVSS.n3525 0.00641429
R19479 DVSS.n3516 VSS 0.00641429
R19480 DVSS.n463 DVSS.n462 0.00640498
R19481 DVSS.n2615 DVSS.n2614 0.00635
R19482 DVSS.n3946 DVSS.n3945 0.00635
R19483 DVSS.n1720 DVSS.n1708 0.00635
R19484 DVSS.n1721 DVSS.n1720 0.00635
R19485 DVSS.n3295 DVSS.n3294 0.00626355
R19486 DVSS.n3234 DVSS.n3005 0.00626355
R19487 DVSS.n4154 DVSS.n1537 0.006125
R19488 DVSS.n1531 DVSS.n1526 0.006125
R19489 DVSS.n1971 DVSS.n1969 0.00609286
R19490 DVSS.n4885 VSS 0.00609286
R19491 DVSS.n3756 VSS 0.00609286
R19492 DVSS.n4377 DVSS.n4343 0.00602857
R19493 DVSS.n4376 DVSS.n4372 0.00602857
R19494 DVSS.n4383 DVSS.n4341 0.00602857
R19495 DVSS.n3435 DVSS.n2762 0.006
R19496 DVSS.n3335 DVSS.n3334 0.006
R19497 DVSS.n3096 DVSS.n3094 0.006
R19498 DVSS.n3198 DVSS.n2907 0.006
R19499 DVSS.n4771 DVSS.n1356 0.0059878
R19500 DVSS.n4769 DVSS.n4767 0.0059878
R19501 DVSS.n4733 DVSS.n4732 0.00596429
R19502 DVSS.n4729 DVSS.n4607 0.00596429
R19503 DVSS.n4728 DVSS.n4610 0.00596429
R19504 DVSS.n4617 DVSS.n4616 0.00596429
R19505 DVSS.n4722 DVSS.n4721 0.00596429
R19506 DVSS.n4627 DVSS.n4618 0.00596429
R19507 DVSS.n4716 DVSS.n4628 0.00596429
R19508 DVSS.n4013 DVSS.n4012 0.00583571
R19509 DVSS.n4029 DVSS.n4028 0.00570714
R19510 DVSS.n1955 DVSS.n1954 0.00561229
R19511 DVSS.n2230 DVSS.n1961 0.00561229
R19512 DVSS DVSS.n2766 0.00559852
R19513 DVSS.n2824 DVSS.n2822 0.00559852
R19514 DVSS.n3089 DVSS 0.00559852
R19515 DVSS.n3130 DVSS.n3129 0.00559852
R19516 DVSS.n5340 DVSS.n959 0.00559091
R19517 DVSS.n2300 DVSS.n1874 0.00551429
R19518 DVSS.n2296 DVSS.n1876 0.00551429
R19519 DVSS.n2269 DVSS.n1873 0.00551429
R19520 DVSS.n3456 DVSS.n3455 0.0055
R19521 DVSS.n2945 DVSS.n2944 0.0055
R19522 DVSS.n3073 DVSS.n2736 0.0055
R19523 DVSS.n3219 DVSS.n3218 0.0055
R19524 DVSS.n4680 DVSS.n4679 0.00548841
R19525 DVSS.n3766 DVSS.n3524 0.00548841
R19526 DVSS.n1573 DVSS.n1572 0.00548841
R19527 DVSS.n5091 DVSS.n1083 0.00548841
R19528 DVSS.n3520 DVSS.n3515 0.00548841
R19529 DVSS DVSS.n5533 0.00538571
R19530 DVSS.n4691 DVSS 0.00538571
R19531 DVSS.n2367 DVSS.n2353 0.00538571
R19532 DVSS.n2362 DVSS.n2360 0.00538571
R19533 DVSS.n2364 DVSS.n2345 0.00538571
R19534 DVSS.n3017 DVSS.n2784 0.00537685
R19535 DVSS.n3103 DVSS.n3018 0.00537685
R19536 DVSS.n4621 DVSS.n4609 0.00532927
R19537 DVSS.n4720 DVSS.n4719 0.00532927
R19538 DVSS.n4590 DVSS.n4588 0.00532927
R19539 DVSS.n4750 DVSS.n1398 0.00532927
R19540 DVSS.n4548 DVSS.n1427 0.00532927
R19541 DVSS.n4565 DVSS.n4564 0.00532927
R19542 DVSS.n4447 DVSS.n1447 0.00532927
R19543 DVSS.n4525 DVSS.n4524 0.00532927
R19544 DVSS.n4428 DVSS.n4416 0.00532927
R19545 DVSS.n4472 DVSS.n4471 0.00532927
R19546 DVSS.n4397 DVSS.n4395 0.00532927
R19547 DVSS.n4502 DVSS.n4327 0.00532927
R19548 DVSS.n1972 DVSS.n1850 0.00519286
R19549 DVSS.n3913 DVSS.n1730 0.00519286
R19550 DVSS.n4091 DVSS.n4090 0.00519286
R19551 DVSS.n2231 DVSS.n1951 0.00514674
R19552 DVSS.n4765 DVSS.n4764 0.00505741
R19553 DVSS.n4764 DVSS.n961 0.00505741
R19554 DVSS.n958 DVSS.n956 0.00505741
R19555 DVSS.n1450 DVSS.n958 0.00505741
R19556 DVSS.n2323 DVSS.n1916 0.00504128
R19557 DVSS.n2570 DVSS.n1888 0.00504128
R19558 DVSS.n3483 DVSS.n2696 0.005
R19559 DVSS.n3476 DVSS.n2708 0.005
R19560 DVSS.n3291 DVSS.n2968 0.005
R19561 DVSS.n3284 DVSS.n2980 0.005
R19562 DVSS.n3044 DVSS.n2698 0.005
R19563 DVSS.n3046 DVSS.n2706 0.005
R19564 DVSS.n3241 DVSS.n2970 0.005
R19565 DVSS.n3243 DVSS.n2978 0.005
R19566 DVSS.n5715 DVSS.n5714 0.00498878
R19567 DVSS.n5341 DVSS.n5340 0.0049789
R19568 DVSS.n5340 DVSS.n5339 0.0049789
R19569 DVSS.n1972 DVSS.n1854 0.00493571
R19570 DVSS.n1734 DVSS.n1730 0.00493571
R19571 DVSS.n4091 DVSS.n1557 0.00493571
R19572 DVSS.n2948 DVSS.n2947 0.0049335
R19573 DVSS.n3221 DVSS.n3220 0.0049335
R19574 DVSS.n2234 DVSS.n1963 0.00489894
R19575 DVSS.n2238 DVSS.n2228 0.00489894
R19576 DVSS.n2012 DVSS.n2011 0.00476
R19577 DVSS.n2011 DVSS.n2010 0.00476
R19578 DVSS.n2010 DVSS.n1981 0.00476
R19579 DVSS.n2006 DVSS.n1981 0.00476
R19580 DVSS.n2006 DVSS.n2005 0.00476
R19581 DVSS.n2005 DVSS.n2004 0.00476
R19582 DVSS.n2004 DVSS.n1987 0.00476
R19583 DVSS.n2000 DVSS.n1987 0.00476
R19584 DVSS.n2000 DVSS.n1999 0.00476
R19585 DVSS.n1999 DVSS.n1998 0.00476
R19586 DVSS.n1998 DVSS.n1995 0.00476
R19587 DVSS.n1995 DVSS.n1496 0.00476
R19588 DVSS.n4188 DVSS.n1496 0.00476
R19589 DVSS.n4188 DVSS.n1494 0.00476
R19590 DVSS.n4192 DVSS.n1494 0.00476
R19591 DVSS.n4192 DVSS.n1492 0.00476
R19592 DVSS.n4196 DVSS.n1492 0.00476
R19593 DVSS.n4196 DVSS.n1490 0.00476
R19594 DVSS.n4200 DVSS.n1490 0.00476
R19595 DVSS.n4200 DVSS.n1488 0.00476
R19596 DVSS.n4204 DVSS.n1488 0.00476
R19597 DVSS.n4204 DVSS.n1486 0.00476
R19598 DVSS.n4280 DVSS.n1486 0.00476
R19599 DVSS.n4280 DVSS.n4279 0.00476
R19600 DVSS.n4279 DVSS.n4278 0.00476
R19601 DVSS.n4278 DVSS.n4210 0.00476
R19602 DVSS.n4274 DVSS.n4210 0.00476
R19603 DVSS.n4274 DVSS.n4273 0.00476
R19604 DVSS.n4273 DVSS.n4272 0.00476
R19605 DVSS.n4272 DVSS.n4216 0.00476
R19606 DVSS.n4268 DVSS.n4216 0.00476
R19607 DVSS.n4268 DVSS.n4267 0.00476
R19608 DVSS.n4267 DVSS.n4266 0.00476
R19609 DVSS.n4266 DVSS.n4222 0.00476
R19610 DVSS.n4262 DVSS.n4222 0.00476
R19611 DVSS.n4262 DVSS.n4261 0.00476
R19612 DVSS.n4261 DVSS.n4260 0.00476
R19613 DVSS.n4260 DVSS.n4228 0.00476
R19614 DVSS.n4256 DVSS.n4228 0.00476
R19615 DVSS.n4256 DVSS.n4255 0.00476
R19616 DVSS.n4255 DVSS.n4254 0.00476
R19617 DVSS.n4254 DVSS.n4234 0.00476
R19618 DVSS.n4250 DVSS.n4234 0.00476
R19619 DVSS.n4250 DVSS.n4249 0.00476
R19620 DVSS.n4249 DVSS.n4248 0.00476
R19621 DVSS.n4248 DVSS.n4240 0.00476
R19622 DVSS.n4244 DVSS.n4240 0.00476
R19623 DVSS.n4244 DVSS.n1237 0.00476
R19624 DVSS.n4800 DVSS.n1237 0.00476
R19625 DVSS.n4800 DVSS.n4799 0.00476
R19626 DVSS.n4799 DVSS.n4798 0.00476
R19627 DVSS.n4798 DVSS.n1241 0.00476
R19628 DVSS.n4794 DVSS.n1241 0.00476
R19629 DVSS.n4794 DVSS.n4793 0.00476
R19630 DVSS.n4793 DVSS.n4792 0.00476
R19631 DVSS.n4792 DVSS.n1247 0.00476
R19632 DVSS.n1301 DVSS.n1247 0.00476
R19633 DVSS.n1301 DVSS.n1298 0.00476
R19634 DVSS.n1305 DVSS.n1298 0.00476
R19635 DVSS.n1305 DVSS.n1296 0.00476
R19636 DVSS.n1309 DVSS.n1296 0.00476
R19637 DVSS.n1309 DVSS.n1294 0.00476
R19638 DVSS.n1314 DVSS.n1294 0.00476
R19639 DVSS.n1314 DVSS.n1292 0.00476
R19640 DVSS.n1318 DVSS.n1292 0.00476
R19641 DVSS.n1318 DVSS.n1290 0.00476
R19642 DVSS.n1322 DVSS.n1290 0.00476
R19643 DVSS.n1322 DVSS.n1288 0.00476
R19644 DVSS.n1326 DVSS.n1288 0.00476
R19645 DVSS.n1326 DVSS.n1286 0.00476
R19646 DVSS.n1330 DVSS.n1286 0.00476
R19647 DVSS.n1330 DVSS.n1284 0.00476
R19648 DVSS.n1334 DVSS.n1284 0.00476
R19649 DVSS.n1334 DVSS.n1282 0.00476
R19650 DVSS.n1338 DVSS.n1282 0.00476
R19651 DVSS.n1338 DVSS.n1280 0.00476
R19652 DVSS.n1342 DVSS.n1280 0.00476
R19653 DVSS.n1350 DVSS.n1278 0.00476
R19654 DVSS.n4775 DVSS.n1278 0.00476
R19655 DVSS.n4775 DVSS.n4774 0.00476
R19656 DVSS.n2013 DVSS.n1978 0.00476
R19657 DVSS.n2009 DVSS.n1978 0.00476
R19658 DVSS.n2009 DVSS.n2008 0.00476
R19659 DVSS.n2008 DVSS.n2007 0.00476
R19660 DVSS.n2007 DVSS.n1982 0.00476
R19661 DVSS.n2003 DVSS.n2002 0.00476
R19662 DVSS.n2002 DVSS.n2001 0.00476
R19663 DVSS.n2001 DVSS.n1989 0.00476
R19664 DVSS.n1997 DVSS.n1989 0.00476
R19665 DVSS.n1997 DVSS.n1996 0.00476
R19666 DVSS.n1996 DVSS.n1497 0.00476
R19667 DVSS.n4187 DVSS.n1493 0.00476
R19668 DVSS.n4193 DVSS.n1493 0.00476
R19669 DVSS.n4194 DVSS.n4193 0.00476
R19670 DVSS.n4195 DVSS.n4194 0.00476
R19671 DVSS.n4195 DVSS.n1489 0.00476
R19672 DVSS.n4201 DVSS.n1489 0.00476
R19673 DVSS.n4202 DVSS.n4201 0.00476
R19674 DVSS.n4203 DVSS.n4202 0.00476
R19675 DVSS.n4203 DVSS.n1484 0.00476
R19676 DVSS.n4281 DVSS.n1485 0.00476
R19677 DVSS.n4277 DVSS.n1485 0.00476
R19678 DVSS.n4277 DVSS.n4276 0.00476
R19679 DVSS.n4276 DVSS.n4275 0.00476
R19680 DVSS.n4275 DVSS.n4211 0.00476
R19681 DVSS.n4271 DVSS.n4211 0.00476
R19682 DVSS.n4271 DVSS.n4270 0.00476
R19683 DVSS.n4270 DVSS.n4269 0.00476
R19684 DVSS.n4269 DVSS.n4217 0.00476
R19685 DVSS.n4265 DVSS.n4217 0.00476
R19686 DVSS.n4265 DVSS.n4264 0.00476
R19687 DVSS.n4264 DVSS.n4263 0.00476
R19688 DVSS.n4263 DVSS.n4223 0.00476
R19689 DVSS.n4259 DVSS.n4223 0.00476
R19690 DVSS.n4259 DVSS.n4258 0.00476
R19691 DVSS.n4258 DVSS.n4257 0.00476
R19692 DVSS.n4257 DVSS.n4229 0.00476
R19693 DVSS.n4253 DVSS.n4229 0.00476
R19694 DVSS.n4253 DVSS.n4252 0.00476
R19695 DVSS.n4252 DVSS.n4251 0.00476
R19696 DVSS.n4251 DVSS.n4235 0.00476
R19697 DVSS.n4247 DVSS.n4235 0.00476
R19698 DVSS.n4247 DVSS.n4246 0.00476
R19699 DVSS.n4246 DVSS.n4245 0.00476
R19700 DVSS.n4245 DVSS.n1235 0.00476
R19701 DVSS.n4801 DVSS.n1236 0.00476
R19702 DVSS.n4797 DVSS.n1236 0.00476
R19703 DVSS.n4797 DVSS.n4796 0.00476
R19704 DVSS.n4796 DVSS.n4795 0.00476
R19705 DVSS.n4795 DVSS.n1242 0.00476
R19706 DVSS.n4791 DVSS.n1242 0.00476
R19707 DVSS.n1302 DVSS.n1248 0.00476
R19708 DVSS.n1303 DVSS.n1302 0.00476
R19709 DVSS.n1304 DVSS.n1303 0.00476
R19710 DVSS.n1304 DVSS.n1295 0.00476
R19711 DVSS.n1310 DVSS.n1295 0.00476
R19712 DVSS.n1313 DVSS.n1312 0.00476
R19713 DVSS.n1313 DVSS.n1291 0.00476
R19714 DVSS.n1319 DVSS.n1291 0.00476
R19715 DVSS.n1320 DVSS.n1319 0.00476
R19716 DVSS.n1321 DVSS.n1320 0.00476
R19717 DVSS.n1321 DVSS.n1287 0.00476
R19718 DVSS.n1327 DVSS.n1287 0.00476
R19719 DVSS.n1328 DVSS.n1327 0.00476
R19720 DVSS.n1329 DVSS.n1328 0.00476
R19721 DVSS.n1329 DVSS.n1283 0.00476
R19722 DVSS.n1335 DVSS.n1283 0.00476
R19723 DVSS.n1336 DVSS.n1335 0.00476
R19724 DVSS.n1337 DVSS.n1336 0.00476
R19725 DVSS.n1337 DVSS.n1279 0.00476
R19726 DVSS.n1343 DVSS.n1279 0.00476
R19727 DVSS.n4776 DVSS.n1277 0.00476
R19728 DVSS.n258 DVSS.n257 0.00476
R19729 DVSS.n313 DVSS.n312 0.00476
R19730 DVSS.n316 DVSS.n313 0.00476
R19731 DVSS.n317 DVSS.n316 0.00476
R19732 DVSS.n318 DVSS.n317 0.00476
R19733 DVSS.n319 DVSS.n318 0.00476
R19734 DVSS.n322 DVSS.n319 0.00476
R19735 DVSS.n323 DVSS.n322 0.00476
R19736 DVSS.n324 DVSS.n323 0.00476
R19737 DVSS.n325 DVSS.n324 0.00476
R19738 DVSS.n328 DVSS.n325 0.00476
R19739 DVSS.n329 DVSS.n328 0.00476
R19740 DVSS.n330 DVSS.n329 0.00476
R19741 DVSS.n331 DVSS.n330 0.00476
R19742 DVSS.n332 DVSS.n331 0.00476
R19743 DVSS.n332 DVSS.n193 0.00476
R19744 DVSS.n622 DVSS.n193 0.00476
R19745 DVSS.n628 DVSS.n189 0.00476
R19746 DVSS.n629 DVSS.n628 0.00476
R19747 DVSS.n630 DVSS.n629 0.00476
R19748 DVSS.n637 DVSS.n636 0.00476
R19749 DVSS.n638 DVSS.n637 0.00476
R19750 DVSS.n638 DVSS.n180 0.00476
R19751 DVSS.n644 DVSS.n180 0.00476
R19752 DVSS.n645 DVSS.n644 0.00476
R19753 DVSS.n646 DVSS.n645 0.00476
R19754 DVSS.n646 DVSS.n176 0.00476
R19755 DVSS.n652 DVSS.n176 0.00476
R19756 DVSS.n653 DVSS.n652 0.00476
R19757 DVSS.n654 DVSS.n653 0.00476
R19758 DVSS.n654 DVSS.n170 0.00476
R19759 DVSS.n686 DVSS.n171 0.00476
R19760 DVSS.n659 DVSS.n171 0.00476
R19761 DVSS.n660 DVSS.n659 0.00476
R19762 DVSS.n661 DVSS.n660 0.00476
R19763 DVSS.n664 DVSS.n661 0.00476
R19764 DVSS.n665 DVSS.n664 0.00476
R19765 DVSS.n666 DVSS.n665 0.00476
R19766 DVSS.n667 DVSS.n666 0.00476
R19767 DVSS.n669 DVSS.n667 0.00476
R19768 DVSS.n669 DVSS.n668 0.00476
R19769 DVSS.n668 DVSS.n132 0.00476
R19770 DVSS.n5658 DVSS.n127 0.00476
R19771 DVSS.n5659 DVSS.n5658 0.00476
R19772 DVSS.n5661 DVSS.n5659 0.00476
R19773 DVSS.n5661 DVSS.n5660 0.00476
R19774 DVSS.n5668 DVSS.n5667 0.00476
R19775 DVSS.n5669 DVSS.n5668 0.00476
R19776 DVSS.n5669 DVSS.n119 0.00476
R19777 DVSS.n5675 DVSS.n119 0.00476
R19778 DVSS.n5676 DVSS.n5675 0.00476
R19779 DVSS.n5677 DVSS.n5676 0.00476
R19780 DVSS.n5677 DVSS.n115 0.00476
R19781 DVSS.n5683 DVSS.n115 0.00476
R19782 DVSS.n5684 DVSS.n5683 0.00476
R19783 DVSS.n5685 DVSS.n5684 0.00476
R19784 DVSS.n5685 DVSS.n111 0.00476
R19785 DVSS.n5691 DVSS.n111 0.00476
R19786 DVSS.n5692 DVSS.n5691 0.00476
R19787 DVSS.n5693 DVSS.n5692 0.00476
R19788 DVSS.n5693 DVSS.n102 0.00476
R19789 DVSS.n5700 DVSS.n103 0.00476
R19790 DVSS.n5765 DVSS.n5764 0.00476
R19791 DVSS.n5766 DVSS.n5765 0.00476
R19792 DVSS.n5766 DVSS.n36 0.00476
R19793 DVSS.n5772 DVSS.n36 0.00476
R19794 DVSS.n5773 DVSS.n5772 0.00476
R19795 DVSS.n5774 DVSS.n5773 0.00476
R19796 DVSS.n5774 DVSS.n32 0.00476
R19797 DVSS.n5780 DVSS.n32 0.00476
R19798 DVSS.n5781 DVSS.n5780 0.00476
R19799 DVSS.n5782 DVSS.n5781 0.00476
R19800 DVSS.n5788 DVSS.n5787 0.00476
R19801 DVSS.n5789 DVSS.n5788 0.00476
R19802 DVSS.n5789 DVSS.n26 0.00476
R19803 DVSS.n424 DVSS.n244 0.00476
R19804 DVSS.n375 DVSS.n374 0.00476
R19805 DVSS.n376 DVSS.n375 0.00476
R19806 DVSS.n379 DVSS.n376 0.00476
R19807 DVSS.n380 DVSS.n379 0.00476
R19808 DVSS.n381 DVSS.n380 0.00476
R19809 DVSS.n382 DVSS.n381 0.00476
R19810 DVSS.n385 DVSS.n382 0.00476
R19811 DVSS.n386 DVSS.n385 0.00476
R19812 DVSS.n387 DVSS.n386 0.00476
R19813 DVSS.n388 DVSS.n387 0.00476
R19814 DVSS.n391 DVSS.n388 0.00476
R19815 DVSS.n392 DVSS.n391 0.00476
R19816 DVSS.n393 DVSS.n392 0.00476
R19817 DVSS.n394 DVSS.n393 0.00476
R19818 DVSS.n395 DVSS.n394 0.00476
R19819 DVSS.n395 DVSS.n195 0.00476
R19820 DVSS.n618 DVSS.n196 0.00476
R19821 DVSS.n201 DVSS.n196 0.00476
R19822 DVSS.n202 DVSS.n201 0.00476
R19823 DVSS.n581 DVSS.n578 0.00476
R19824 DVSS.n582 DVSS.n581 0.00476
R19825 DVSS.n583 DVSS.n582 0.00476
R19826 DVSS.n584 DVSS.n583 0.00476
R19827 DVSS.n587 DVSS.n584 0.00476
R19828 DVSS.n588 DVSS.n587 0.00476
R19829 DVSS.n589 DVSS.n588 0.00476
R19830 DVSS.n590 DVSS.n589 0.00476
R19831 DVSS.n592 DVSS.n590 0.00476
R19832 DVSS.n593 DVSS.n592 0.00476
R19833 DVSS.n593 DVSS.n168 0.00476
R19834 DVSS.n690 DVSS.n164 0.00476
R19835 DVSS.n696 DVSS.n164 0.00476
R19836 DVSS.n697 DVSS.n696 0.00476
R19837 DVSS.n698 DVSS.n697 0.00476
R19838 DVSS.n698 DVSS.n160 0.00476
R19839 DVSS.n704 DVSS.n160 0.00476
R19840 DVSS.n705 DVSS.n704 0.00476
R19841 DVSS.n706 DVSS.n705 0.00476
R19842 DVSS.n706 DVSS.n156 0.00476
R19843 DVSS.n713 DVSS.n156 0.00476
R19844 DVSS.n714 DVSS.n713 0.00476
R19845 DVSS.n138 DVSS.n135 0.00476
R19846 DVSS.n139 DVSS.n138 0.00476
R19847 DVSS.n140 DVSS.n139 0.00476
R19848 DVSS.n141 DVSS.n140 0.00476
R19849 DVSS.n5603 DVSS.n5602 0.00476
R19850 DVSS.n5604 DVSS.n5603 0.00476
R19851 DVSS.n5605 DVSS.n5604 0.00476
R19852 DVSS.n5608 DVSS.n5605 0.00476
R19853 DVSS.n5609 DVSS.n5608 0.00476
R19854 DVSS.n5610 DVSS.n5609 0.00476
R19855 DVSS.n5611 DVSS.n5610 0.00476
R19856 DVSS.n5614 DVSS.n5611 0.00476
R19857 DVSS.n5615 DVSS.n5614 0.00476
R19858 DVSS.n5616 DVSS.n5615 0.00476
R19859 DVSS.n5617 DVSS.n5616 0.00476
R19860 DVSS.n5619 DVSS.n5617 0.00476
R19861 DVSS.n5620 DVSS.n5619 0.00476
R19862 DVSS.n5620 DVSS.n53 0.00476
R19863 DVSS.n5717 DVSS.n53 0.00476
R19864 DVSS.n54 DVSS.n50 0.00476
R19865 DVSS.n5727 DVSS.n5726 0.00476
R19866 DVSS.n5728 DVSS.n5727 0.00476
R19867 DVSS.n5731 DVSS.n5728 0.00476
R19868 DVSS.n5732 DVSS.n5731 0.00476
R19869 DVSS.n5733 DVSS.n5732 0.00476
R19870 DVSS.n5734 DVSS.n5733 0.00476
R19871 DVSS.n5737 DVSS.n5734 0.00476
R19872 DVSS.n5738 DVSS.n5737 0.00476
R19873 DVSS.n5739 DVSS.n5738 0.00476
R19874 DVSS.n5741 DVSS.n5739 0.00476
R19875 DVSS.n5741 DVSS.n5740 0.00476
R19876 DVSS.n4 DVSS.n1 0.00476
R19877 DVSS.n5 DVSS.n4 0.00476
R19878 DVSS.n465 DVSS.n228 0.00476
R19879 DVSS.n471 DVSS.n224 0.00476
R19880 DVSS.n472 DVSS.n471 0.00476
R19881 DVSS.n473 DVSS.n472 0.00476
R19882 DVSS.n473 DVSS.n220 0.00476
R19883 DVSS.n479 DVSS.n220 0.00476
R19884 DVSS.n480 DVSS.n479 0.00476
R19885 DVSS.n481 DVSS.n480 0.00476
R19886 DVSS.n481 DVSS.n216 0.00476
R19887 DVSS.n487 DVSS.n216 0.00476
R19888 DVSS.n488 DVSS.n487 0.00476
R19889 DVSS.n489 DVSS.n488 0.00476
R19890 DVSS.n489 DVSS.n212 0.00476
R19891 DVSS.n495 DVSS.n212 0.00476
R19892 DVSS.n496 DVSS.n495 0.00476
R19893 DVSS.n498 DVSS.n496 0.00476
R19894 DVSS.n498 DVSS.n497 0.00476
R19895 DVSS.n506 DVSS.n505 0.00476
R19896 DVSS.n507 DVSS.n506 0.00476
R19897 DVSS.n507 DVSS.n204 0.00476
R19898 DVSS.n575 DVSS.n205 0.00476
R19899 DVSS.n513 DVSS.n205 0.00476
R19900 DVSS.n514 DVSS.n513 0.00476
R19901 DVSS.n515 DVSS.n514 0.00476
R19902 DVSS.n518 DVSS.n515 0.00476
R19903 DVSS.n519 DVSS.n518 0.00476
R19904 DVSS.n520 DVSS.n519 0.00476
R19905 DVSS.n521 DVSS.n520 0.00476
R19906 DVSS.n524 DVSS.n521 0.00476
R19907 DVSS.n525 DVSS.n524 0.00476
R19908 DVSS.n526 DVSS.n525 0.00476
R19909 DVSS.n530 DVSS.n527 0.00476
R19910 DVSS.n531 DVSS.n530 0.00476
R19911 DVSS.n532 DVSS.n531 0.00476
R19912 DVSS.n533 DVSS.n532 0.00476
R19913 DVSS.n536 DVSS.n533 0.00476
R19914 DVSS.n537 DVSS.n536 0.00476
R19915 DVSS.n538 DVSS.n537 0.00476
R19916 DVSS.n539 DVSS.n538 0.00476
R19917 DVSS.n540 DVSS.n539 0.00476
R19918 DVSS.n540 DVSS.n154 0.00476
R19919 DVSS.n717 DVSS.n154 0.00476
R19920 DVSS.n724 DVSS.n150 0.00476
R19921 DVSS.n725 DVSS.n724 0.00476
R19922 DVSS.n726 DVSS.n725 0.00476
R19923 DVSS.n726 DVSS.n144 0.00476
R19924 DVSS.n5598 DVSS.n145 0.00476
R19925 DVSS.n731 DVSS.n145 0.00476
R19926 DVSS.n732 DVSS.n731 0.00476
R19927 DVSS.n733 DVSS.n732 0.00476
R19928 DVSS.n736 DVSS.n733 0.00476
R19929 DVSS.n737 DVSS.n736 0.00476
R19930 DVSS.n738 DVSS.n737 0.00476
R19931 DVSS.n739 DVSS.n738 0.00476
R19932 DVSS.n742 DVSS.n739 0.00476
R19933 DVSS.n743 DVSS.n742 0.00476
R19934 DVSS.n744 DVSS.n743 0.00476
R19935 DVSS.n745 DVSS.n744 0.00476
R19936 DVSS.n748 DVSS.n745 0.00476
R19937 DVSS.n749 DVSS.n748 0.00476
R19938 DVSS.n750 DVSS.n749 0.00476
R19939 DVSS.n753 DVSS.n751 0.00476
R19940 DVSS.n809 DVSS.n806 0.00476
R19941 DVSS.n810 DVSS.n809 0.00476
R19942 DVSS.n811 DVSS.n810 0.00476
R19943 DVSS.n812 DVSS.n811 0.00476
R19944 DVSS.n815 DVSS.n812 0.00476
R19945 DVSS.n816 DVSS.n815 0.00476
R19946 DVSS.n817 DVSS.n816 0.00476
R19947 DVSS.n818 DVSS.n817 0.00476
R19948 DVSS.n821 DVSS.n818 0.00476
R19949 DVSS.n822 DVSS.n821 0.00476
R19950 DVSS.n824 DVSS.n823 0.00476
R19951 DVSS.n827 DVSS.n824 0.00476
R19952 DVSS.n828 DVSS.n827 0.00476
R19953 DVSS.n367 DVSS.n227 0.00476
R19954 DVSS.n466 DVSS.n227 0.00476
R19955 DVSS.n466 DVSS.n225 0.00476
R19956 DVSS.n470 DVSS.n225 0.00476
R19957 DVSS.n470 DVSS.n223 0.00476
R19958 DVSS.n474 DVSS.n223 0.00476
R19959 DVSS.n474 DVSS.n221 0.00476
R19960 DVSS.n478 DVSS.n221 0.00476
R19961 DVSS.n478 DVSS.n219 0.00476
R19962 DVSS.n482 DVSS.n219 0.00476
R19963 DVSS.n482 DVSS.n217 0.00476
R19964 DVSS.n486 DVSS.n217 0.00476
R19965 DVSS.n486 DVSS.n215 0.00476
R19966 DVSS.n490 DVSS.n215 0.00476
R19967 DVSS.n490 DVSS.n213 0.00476
R19968 DVSS.n494 DVSS.n213 0.00476
R19969 DVSS.n494 DVSS.n211 0.00476
R19970 DVSS.n499 DVSS.n211 0.00476
R19971 DVSS.n499 DVSS.n209 0.00476
R19972 DVSS.n504 DVSS.n209 0.00476
R19973 DVSS.n504 DVSS.n208 0.00476
R19974 DVSS.n508 DVSS.n208 0.00476
R19975 DVSS.n509 DVSS.n508 0.00476
R19976 DVSS.n574 DVSS.n206 0.00476
R19977 DVSS.n570 DVSS.n206 0.00476
R19978 DVSS.n570 DVSS.n569 0.00476
R19979 DVSS.n569 DVSS.n568 0.00476
R19980 DVSS.n568 DVSS.n516 0.00476
R19981 DVSS.n564 DVSS.n516 0.00476
R19982 DVSS.n564 DVSS.n563 0.00476
R19983 DVSS.n563 DVSS.n562 0.00476
R19984 DVSS.n562 DVSS.n522 0.00476
R19985 DVSS.n558 DVSS.n522 0.00476
R19986 DVSS.n558 DVSS.n557 0.00476
R19987 DVSS.n557 DVSS.n556 0.00476
R19988 DVSS.n556 DVSS.n528 0.00476
R19989 DVSS.n552 DVSS.n528 0.00476
R19990 DVSS.n552 DVSS.n551 0.00476
R19991 DVSS.n551 DVSS.n550 0.00476
R19992 DVSS.n550 DVSS.n534 0.00476
R19993 DVSS.n546 DVSS.n534 0.00476
R19994 DVSS.n546 DVSS.n545 0.00476
R19995 DVSS.n545 DVSS.n544 0.00476
R19996 DVSS.n544 DVSS.n541 0.00476
R19997 DVSS.n541 DVSS.n153 0.00476
R19998 DVSS.n718 DVSS.n153 0.00476
R19999 DVSS.n723 DVSS.n151 0.00476
R20000 DVSS.n723 DVSS.n149 0.00476
R20001 DVSS.n727 DVSS.n149 0.00476
R20002 DVSS.n727 DVSS.n146 0.00476
R20003 DVSS.n5597 DVSS.n146 0.00476
R20004 DVSS.n5597 DVSS.n147 0.00476
R20005 DVSS.n5593 DVSS.n147 0.00476
R20006 DVSS.n5593 DVSS.n5592 0.00476
R20007 DVSS.n5592 DVSS.n5591 0.00476
R20008 DVSS.n5591 DVSS.n734 0.00476
R20009 DVSS.n5587 DVSS.n734 0.00476
R20010 DVSS.n5587 DVSS.n5586 0.00476
R20011 DVSS.n5586 DVSS.n5585 0.00476
R20012 DVSS.n5585 DVSS.n740 0.00476
R20013 DVSS.n5581 DVSS.n740 0.00476
R20014 DVSS.n5581 DVSS.n5580 0.00476
R20015 DVSS.n5580 DVSS.n5579 0.00476
R20016 DVSS.n5579 DVSS.n746 0.00476
R20017 DVSS.n5575 DVSS.n746 0.00476
R20018 DVSS.n5575 DVSS.n5574 0.00476
R20019 DVSS.n5574 DVSS.n5573 0.00476
R20020 DVSS.n5573 DVSS.n752 0.00476
R20021 DVSS.n5569 DVSS.n752 0.00476
R20022 DVSS.n5567 DVSS.n807 0.00476
R20023 DVSS.n5563 DVSS.n807 0.00476
R20024 DVSS.n5563 DVSS.n5562 0.00476
R20025 DVSS.n5562 DVSS.n5561 0.00476
R20026 DVSS.n5561 DVSS.n813 0.00476
R20027 DVSS.n5557 DVSS.n813 0.00476
R20028 DVSS.n5557 DVSS.n5556 0.00476
R20029 DVSS.n5556 DVSS.n5555 0.00476
R20030 DVSS.n5555 DVSS.n819 0.00476
R20031 DVSS.n5551 DVSS.n819 0.00476
R20032 DVSS.n5550 DVSS.n5549 0.00476
R20033 DVSS.n5549 DVSS.n825 0.00476
R20034 DVSS.n826 DVSS.n825 0.00476
R20035 DVSS.n423 DVSS.n245 0.00476
R20036 DVSS.n423 DVSS.n246 0.00476
R20037 DVSS.n419 DVSS.n246 0.00476
R20038 DVSS.n419 DVSS.n418 0.00476
R20039 DVSS.n418 DVSS.n417 0.00476
R20040 DVSS.n417 DVSS.n377 0.00476
R20041 DVSS.n413 DVSS.n377 0.00476
R20042 DVSS.n413 DVSS.n412 0.00476
R20043 DVSS.n412 DVSS.n411 0.00476
R20044 DVSS.n411 DVSS.n383 0.00476
R20045 DVSS.n407 DVSS.n383 0.00476
R20046 DVSS.n407 DVSS.n406 0.00476
R20047 DVSS.n406 DVSS.n405 0.00476
R20048 DVSS.n405 DVSS.n389 0.00476
R20049 DVSS.n401 DVSS.n389 0.00476
R20050 DVSS.n401 DVSS.n400 0.00476
R20051 DVSS.n400 DVSS.n399 0.00476
R20052 DVSS.n399 DVSS.n396 0.00476
R20053 DVSS.n396 DVSS.n197 0.00476
R20054 DVSS.n617 DVSS.n197 0.00476
R20055 DVSS.n617 DVSS.n198 0.00476
R20056 DVSS.n613 DVSS.n198 0.00476
R20057 DVSS.n613 DVSS.n612 0.00476
R20058 DVSS.n610 DVSS.n579 0.00476
R20059 DVSS.n606 DVSS.n579 0.00476
R20060 DVSS.n606 DVSS.n605 0.00476
R20061 DVSS.n605 DVSS.n604 0.00476
R20062 DVSS.n604 DVSS.n585 0.00476
R20063 DVSS.n600 DVSS.n585 0.00476
R20064 DVSS.n600 DVSS.n599 0.00476
R20065 DVSS.n599 DVSS.n598 0.00476
R20066 DVSS.n598 DVSS.n591 0.00476
R20067 DVSS.n594 DVSS.n591 0.00476
R20068 DVSS.n594 DVSS.n167 0.00476
R20069 DVSS.n691 DVSS.n167 0.00476
R20070 DVSS.n691 DVSS.n165 0.00476
R20071 DVSS.n695 DVSS.n165 0.00476
R20072 DVSS.n695 DVSS.n163 0.00476
R20073 DVSS.n699 DVSS.n163 0.00476
R20074 DVSS.n699 DVSS.n161 0.00476
R20075 DVSS.n703 DVSS.n161 0.00476
R20076 DVSS.n703 DVSS.n159 0.00476
R20077 DVSS.n707 DVSS.n159 0.00476
R20078 DVSS.n707 DVSS.n157 0.00476
R20079 DVSS.n712 DVSS.n157 0.00476
R20080 DVSS.n712 DVSS.n134 0.00476
R20081 DVSS.n5649 DVSS.n136 0.00476
R20082 DVSS.n5645 DVSS.n136 0.00476
R20083 DVSS.n5645 DVSS.n5644 0.00476
R20084 DVSS.n5644 DVSS.n5643 0.00476
R20085 DVSS.n5643 DVSS.n142 0.00476
R20086 DVSS.n5639 DVSS.n142 0.00476
R20087 DVSS.n5639 DVSS.n5638 0.00476
R20088 DVSS.n5638 DVSS.n5637 0.00476
R20089 DVSS.n5637 DVSS.n5606 0.00476
R20090 DVSS.n5633 DVSS.n5606 0.00476
R20091 DVSS.n5633 DVSS.n5632 0.00476
R20092 DVSS.n5632 DVSS.n5631 0.00476
R20093 DVSS.n5631 DVSS.n5612 0.00476
R20094 DVSS.n5627 DVSS.n5612 0.00476
R20095 DVSS.n5627 DVSS.n5626 0.00476
R20096 DVSS.n5626 DVSS.n5625 0.00476
R20097 DVSS.n5625 DVSS.n5618 0.00476
R20098 DVSS.n5621 DVSS.n5618 0.00476
R20099 DVSS.n5621 DVSS.n52 0.00476
R20100 DVSS.n5718 DVSS.n52 0.00476
R20101 DVSS.n5718 DVSS.n49 0.00476
R20102 DVSS.n5722 DVSS.n49 0.00476
R20103 DVSS.n5723 DVSS.n5722 0.00476
R20104 DVSS.n5758 DVSS.n5757 0.00476
R20105 DVSS.n5757 DVSS.n5756 0.00476
R20106 DVSS.n5756 DVSS.n5729 0.00476
R20107 DVSS.n5752 DVSS.n5729 0.00476
R20108 DVSS.n5752 DVSS.n5751 0.00476
R20109 DVSS.n5751 DVSS.n5750 0.00476
R20110 DVSS.n5750 DVSS.n5735 0.00476
R20111 DVSS.n5746 DVSS.n5735 0.00476
R20112 DVSS.n5746 DVSS.n5745 0.00476
R20113 DVSS.n5745 DVSS.n5744 0.00476
R20114 DVSS.n5744 DVSS.n0 0.00476
R20115 DVSS.n5801 DVSS.n2 0.00476
R20116 DVSS.n3 DVSS.n2 0.00476
R20117 DVSS.n360 DVSS.n255 0.00476
R20118 DVSS.n356 DVSS.n255 0.00476
R20119 DVSS.n356 DVSS.n355 0.00476
R20120 DVSS.n355 DVSS.n354 0.00476
R20121 DVSS.n354 DVSS.n314 0.00476
R20122 DVSS.n350 DVSS.n314 0.00476
R20123 DVSS.n350 DVSS.n349 0.00476
R20124 DVSS.n349 DVSS.n348 0.00476
R20125 DVSS.n348 DVSS.n320 0.00476
R20126 DVSS.n344 DVSS.n320 0.00476
R20127 DVSS.n344 DVSS.n343 0.00476
R20128 DVSS.n343 DVSS.n342 0.00476
R20129 DVSS.n342 DVSS.n326 0.00476
R20130 DVSS.n338 DVSS.n326 0.00476
R20131 DVSS.n338 DVSS.n337 0.00476
R20132 DVSS.n337 DVSS.n336 0.00476
R20133 DVSS.n336 DVSS.n333 0.00476
R20134 DVSS.n333 DVSS.n192 0.00476
R20135 DVSS.n623 DVSS.n192 0.00476
R20136 DVSS.n623 DVSS.n190 0.00476
R20137 DVSS.n627 DVSS.n190 0.00476
R20138 DVSS.n627 DVSS.n188 0.00476
R20139 DVSS.n631 DVSS.n188 0.00476
R20140 DVSS.n635 DVSS.n183 0.00476
R20141 DVSS.n639 DVSS.n183 0.00476
R20142 DVSS.n639 DVSS.n181 0.00476
R20143 DVSS.n643 DVSS.n181 0.00476
R20144 DVSS.n643 DVSS.n179 0.00476
R20145 DVSS.n647 DVSS.n179 0.00476
R20146 DVSS.n647 DVSS.n177 0.00476
R20147 DVSS.n651 DVSS.n177 0.00476
R20148 DVSS.n651 DVSS.n175 0.00476
R20149 DVSS.n655 DVSS.n175 0.00476
R20150 DVSS.n655 DVSS.n172 0.00476
R20151 DVSS.n685 DVSS.n172 0.00476
R20152 DVSS.n685 DVSS.n173 0.00476
R20153 DVSS.n681 DVSS.n173 0.00476
R20154 DVSS.n681 DVSS.n680 0.00476
R20155 DVSS.n680 DVSS.n679 0.00476
R20156 DVSS.n679 DVSS.n662 0.00476
R20157 DVSS.n675 DVSS.n662 0.00476
R20158 DVSS.n675 DVSS.n674 0.00476
R20159 DVSS.n674 DVSS.n673 0.00476
R20160 DVSS.n673 DVSS.n670 0.00476
R20161 DVSS.n670 DVSS.n131 0.00476
R20162 DVSS.n5652 DVSS.n131 0.00476
R20163 DVSS.n5657 DVSS.n128 0.00476
R20164 DVSS.n5657 DVSS.n126 0.00476
R20165 DVSS.n5662 DVSS.n126 0.00476
R20166 DVSS.n5662 DVSS.n124 0.00476
R20167 DVSS.n5666 DVSS.n124 0.00476
R20168 DVSS.n5666 DVSS.n122 0.00476
R20169 DVSS.n5670 DVSS.n122 0.00476
R20170 DVSS.n5670 DVSS.n120 0.00476
R20171 DVSS.n5674 DVSS.n120 0.00476
R20172 DVSS.n5674 DVSS.n118 0.00476
R20173 DVSS.n5678 DVSS.n118 0.00476
R20174 DVSS.n5678 DVSS.n116 0.00476
R20175 DVSS.n5682 DVSS.n116 0.00476
R20176 DVSS.n5682 DVSS.n114 0.00476
R20177 DVSS.n5686 DVSS.n114 0.00476
R20178 DVSS.n5686 DVSS.n112 0.00476
R20179 DVSS.n5690 DVSS.n112 0.00476
R20180 DVSS.n5690 DVSS.n110 0.00476
R20181 DVSS.n5694 DVSS.n110 0.00476
R20182 DVSS.n5694 DVSS.n104 0.00476
R20183 DVSS.n5699 DVSS.n104 0.00476
R20184 DVSS.n5699 DVSS.n108 0.00476
R20185 DVSS.n108 DVSS.n107 0.00476
R20186 DVSS.n5763 DVSS.n39 0.00476
R20187 DVSS.n5767 DVSS.n39 0.00476
R20188 DVSS.n5767 DVSS.n37 0.00476
R20189 DVSS.n5771 DVSS.n37 0.00476
R20190 DVSS.n5771 DVSS.n35 0.00476
R20191 DVSS.n5775 DVSS.n35 0.00476
R20192 DVSS.n5775 DVSS.n33 0.00476
R20193 DVSS.n5779 DVSS.n33 0.00476
R20194 DVSS.n5779 DVSS.n31 0.00476
R20195 DVSS.n5783 DVSS.n31 0.00476
R20196 DVSS.n5786 DVSS.n29 0.00476
R20197 DVSS.n5790 DVSS.n29 0.00476
R20198 DVSS.n5790 DVSS.n27 0.00476
R20199 DVSS.n4148 DVSS.n1535 0.00465761
R20200 DVSS.n4147 DVSS.n1532 0.00465761
R20201 DVSS.n2368 DVSS.n2367 0.00461429
R20202 DVSS.n2362 DVSS.n2347 0.00461429
R20203 DVSS.n2364 DVSS.n2348 0.00461429
R20204 DVSS.n5713 DVSS.n57 0.00461371
R20205 DVSS.n5782 DVSS 0.00458
R20206 DVSS.n5783 DVSS 0.00458
R20207 DVSS.n272 DVSS.n242 0.0045724
R20208 DVSS.n511 DVSS.n186 0.0045
R20209 DVSS.n720 DVSS.n129 0.0045
R20210 DVSS.n370 DVSS.n247 0.0045
R20211 DVSS.n633 DVSS.n186 0.0045
R20212 DVSS.n5654 DVSS.n129 0.0045
R20213 DVSS.n5760 DVSS.n43 0.0045
R20214 DVSS.n5761 DVSS.n5760 0.0045
R20215 DVSS.n370 DVSS.n369 0.0045
R20216 DVSS.n2675 DVSS.n2672 0.0045
R20217 DVSS.n3460 DVSS.n2728 0.0045
R20218 DVSS.n2950 DVSS.n2946 0.0045
R20219 DVSS.n3268 DVSS.n3264 0.0045
R20220 DVSS.n3029 DVSS.n3027 0.0045
R20221 DVSS.n3064 DVSS.n3063 0.0045
R20222 DVSS.n3226 DVSS.n3224 0.0045
R20223 DVSS.n3261 DVSS.n3260 0.0045
R20224 DVSS.n2300 DVSS.n2271 0.00448571
R20225 DVSS.n2296 DVSS.n2295 0.00448571
R20226 DVSS.n2269 DVSS.n1877 0.00448571
R20227 DVSS.n4030 DVSS.n4029 0.00442143
R20228 DVSS.n273 DVSS.n241 0.0044172
R20229 DVSS.n361 DVSS.n252 0.00434
R20230 DVSS.n425 DVSS.n243 0.00434
R20231 DVSS.n366 DVSS.n365 0.00434
R20232 DVSS.n2287 DVSS.n1864 0.004325
R20233 DVSS.n2276 DVSS.n1865 0.004325
R20234 DVSS.n4012 DVSS.n4009 0.00429286
R20235 DVSS.n4625 DVSS.n4624 0.00428827
R20236 DVSS.n4753 DVSS.n1395 0.00428827
R20237 DVSS.n4551 DVSS.n4550 0.00428827
R20238 DVSS.n4512 DVSS.n4511 0.00428827
R20239 DVSS.n4432 DVSS.n4431 0.00428827
R20240 DVSS.n4505 DVSS.n4324 0.00428827
R20241 DVSS.n621 DVSS.n189 0.00425
R20242 DVSS.n619 DVSS.n618 0.00425
R20243 DVSS.n505 DVSS.n194 0.00425
R20244 DVSS.n5797 DVSS.n6 0.00422
R20245 DVSS.n5545 DVSS.n829 0.00422
R20246 DVSS.n4802 DVSS.n1235 0.00419
R20247 DVSS.n4777 DVSS.n1276 0.00419
R20248 DVSS.n2250 DVSS.n1958 0.0041856
R20249 DVSS.n2242 DVSS.n2229 0.0041856
R20250 DVSS.n4732 DVSS.n4607 0.00416429
R20251 DVSS.n4729 DVSS.n4728 0.00416429
R20252 DVSS.n4616 DVSS.n4610 0.00416429
R20253 DVSS.n4722 DVSS.n4617 0.00416429
R20254 DVSS.n4721 DVSS.n4618 0.00416429
R20255 DVSS.n4628 DVSS.n4627 0.00416429
R20256 DVSS.n4716 DVSS.n4715 0.00416429
R20257 DVSS.n4377 DVSS.n4376 0.0041
R20258 DVSS.n4372 DVSS.n4341 0.0041
R20259 DVSS.n1988 DVSS.n1982 0.00407
R20260 DVSS.n4187 DVSS.n4186 0.00407
R20261 DVSS.n3410 DVSS.n2804 0.0040468
R20262 DVSS.n3117 DVSS.n3116 0.0040468
R20263 DVSS.n5764 DVSS.n40 0.00404
R20264 DVSS.n5726 DVSS.n5725 0.00404
R20265 DVSS.n806 DVSS.n47 0.00404
R20266 DVSS.n5568 DVSS.n5567 0.00404
R20267 DVSS.n5758 DVSS.n46 0.00404
R20268 DVSS.n5763 DVSS.n41 0.00404
R20269 DVSS.n2021 DVSS.n1969 0.00403571
R20270 DVSS.n2765 DVSS.n2764 0.004
R20271 DVSS.n3330 DVSS.n3329 0.004
R20272 DVSS.n3090 DVSS.n3019 0.004
R20273 DVSS.n3202 DVSS.n2917 0.004
R20274 DVSS.n4790 DVSS.n1248 0.00395
R20275 DVSS.n1348 DVSS.n1276 0.00395
R20276 DVSS.n5667 DVSS.n123 0.00395
R20277 DVSS.n5602 DVSS.n5601 0.00395
R20278 DVSS.n5599 DVSS.n5598 0.00395
R20279 DVSS.n2369 DVSS.n2330 0.00393049
R20280 DVSS.n2346 DVSS.n2331 0.00393049
R20281 DVSS.n2583 DVSS.n1869 0.00393049
R20282 DVSS.n2586 DVSS.n2585 0.00393049
R20283 DVSS.n1342 DVSS 0.00392
R20284 DVSS DVSS.n1343 0.00392
R20285 DVSS DVSS.n822 0.00392
R20286 DVSS.n5551 DVSS 0.00392
R20287 DVSS.n5712 DVSS.n5711 0.00391137
R20288 DVSS.n5702 DVSS.n101 0.00386658
R20289 DVSS.n4626 DVSS.n4625 0.00382908
R20290 DVSS.n4753 DVSS.n4752 0.00382908
R20291 DVSS.n4550 DVSS.n1418 0.00382908
R20292 DVSS.n4511 DVSS.n1439 0.00382908
R20293 DVSS.n4433 DVSS.n4432 0.00382908
R20294 DVSS.n4505 DVSS.n4504 0.00382908
R20295 DVSS.n4282 DVSS.n4281 0.0038
R20296 DVSS.n155 DVSS.n127 0.0038
R20297 DVSS.n715 DVSS.n135 0.0038
R20298 DVSS.n716 DVSS.n150 0.0038
R20299 DVSS.n151 DVSS.n133 0.0038
R20300 DVSS.n5650 DVSS.n5649 0.0038
R20301 DVSS.n5651 DVSS.n128 0.0038
R20302 DVSS.n3945 DVSS.n1694 0.00377857
R20303 DVSS.n3929 DVSS.n1708 0.00377857
R20304 DVSS.n3923 DVSS.n1721 0.00377857
R20305 DVSS.n276 DVSS.n274 0.00374841
R20306 DVSS.n4122 DVSS.n1547 0.00362245
R20307 DVSS.n3008 DVSS.n2914 0.00360345
R20308 DVSS.n3204 DVSS.n3203 0.00360345
R20309 DVSS.n5701 DVSS.n102 0.00359
R20310 DVSS.n5717 DVSS.n5716 0.00359
R20311 DVSS.n801 DVSS.n750 0.00359
R20312 DVSS.n4392 DVSS.n4336 0.00358571
R20313 DVSS.n4391 DVSS.n4337 0.00358571
R20314 DVSS.n4398 DVSS.n4334 0.00358571
R20315 DVSS.n4400 DVSS.n4399 0.00358571
R20316 DVSS.n4501 DVSS.n4328 0.00358571
R20317 DVSS.n4500 DVSS.n4329 0.00358571
R20318 DVSS.n4409 DVSS.n4406 0.00358571
R20319 DVSS.n636 DVSS.n184 0.00356
R20320 DVSS.n578 DVSS.n577 0.00356
R20321 DVSS.n576 DVSS.n575 0.00356
R20322 DVSS.n574 DVSS.n203 0.00356
R20323 DVSS.n611 DVSS.n610 0.00356
R20324 DVSS.n635 DVSS.n185 0.00356
R20325 DVSS.n310 DVSS.n259 0.0035543
R20326 DVSS DVSS.n1 0.00353
R20327 DVSS DVSS.n5801 0.00353
R20328 DVSS.n3419 DVSS.n2786 0.0035
R20329 DVSS.n2894 DVSS.n2893 0.0035
R20330 DVSS.n3111 DVSS.n2788 0.0035
R20331 DVSS.n3183 DVSS.n3182 0.0035
R20332 DVSS.n803 DVSS.n802 0.00341771
R20333 DVSS.n2512 DVSS.n2338 0.00338991
R20334 DVSS.n5793 DVSS.n26 0.0033824
R20335 DVSS.n4772 DVSS.n1277 0.00338166
R20336 DVSS.n359 DVSS.n358 0.00334
R20337 DVSS.n358 DVSS.n357 0.00334
R20338 DVSS.n357 DVSS.n256 0.00334
R20339 DVSS.n353 DVSS.n256 0.00334
R20340 DVSS.n353 DVSS.n352 0.00334
R20341 DVSS.n352 DVSS.n351 0.00334
R20342 DVSS.n351 DVSS.n315 0.00334
R20343 DVSS.n347 DVSS.n315 0.00334
R20344 DVSS.n347 DVSS.n346 0.00334
R20345 DVSS.n346 DVSS.n345 0.00334
R20346 DVSS.n345 DVSS.n321 0.00334
R20347 DVSS.n341 DVSS.n321 0.00334
R20348 DVSS.n341 DVSS.n340 0.00334
R20349 DVSS.n340 DVSS.n339 0.00334
R20350 DVSS.n339 DVSS.n327 0.00334
R20351 DVSS.n335 DVSS.n327 0.00334
R20352 DVSS.n335 DVSS.n334 0.00334
R20353 DVSS.n334 DVSS.n191 0.00334
R20354 DVSS.n624 DVSS.n191 0.00334
R20355 DVSS.n625 DVSS.n624 0.00334
R20356 DVSS.n626 DVSS.n625 0.00334
R20357 DVSS.n626 DVSS.n187 0.00334
R20358 DVSS.n632 DVSS.n187 0.00334
R20359 DVSS.n634 DVSS.n182 0.00334
R20360 DVSS.n640 DVSS.n182 0.00334
R20361 DVSS.n641 DVSS.n640 0.00334
R20362 DVSS.n642 DVSS.n641 0.00334
R20363 DVSS.n642 DVSS.n178 0.00334
R20364 DVSS.n648 DVSS.n178 0.00334
R20365 DVSS.n649 DVSS.n648 0.00334
R20366 DVSS.n650 DVSS.n649 0.00334
R20367 DVSS.n650 DVSS.n174 0.00334
R20368 DVSS.n656 DVSS.n174 0.00334
R20369 DVSS.n657 DVSS.n656 0.00334
R20370 DVSS.n684 DVSS.n657 0.00334
R20371 DVSS.n684 DVSS.n683 0.00334
R20372 DVSS.n683 DVSS.n682 0.00334
R20373 DVSS.n682 DVSS.n658 0.00334
R20374 DVSS.n678 DVSS.n658 0.00334
R20375 DVSS.n678 DVSS.n677 0.00334
R20376 DVSS.n677 DVSS.n676 0.00334
R20377 DVSS.n676 DVSS.n663 0.00334
R20378 DVSS.n672 DVSS.n663 0.00334
R20379 DVSS.n672 DVSS.n671 0.00334
R20380 DVSS.n671 DVSS.n130 0.00334
R20381 DVSS.n5653 DVSS.n130 0.00334
R20382 DVSS.n5656 DVSS.n5655 0.00334
R20383 DVSS.n5656 DVSS.n125 0.00334
R20384 DVSS.n5663 DVSS.n125 0.00334
R20385 DVSS.n5664 DVSS.n5663 0.00334
R20386 DVSS.n5665 DVSS.n5664 0.00334
R20387 DVSS.n5665 DVSS.n121 0.00334
R20388 DVSS.n5671 DVSS.n121 0.00334
R20389 DVSS.n5672 DVSS.n5671 0.00334
R20390 DVSS.n5673 DVSS.n5672 0.00334
R20391 DVSS.n5673 DVSS.n117 0.00334
R20392 DVSS.n5679 DVSS.n117 0.00334
R20393 DVSS.n5680 DVSS.n5679 0.00334
R20394 DVSS.n5681 DVSS.n5680 0.00334
R20395 DVSS.n5681 DVSS.n113 0.00334
R20396 DVSS.n5687 DVSS.n113 0.00334
R20397 DVSS.n5688 DVSS.n5687 0.00334
R20398 DVSS.n5689 DVSS.n5688 0.00334
R20399 DVSS.n5689 DVSS.n109 0.00334
R20400 DVSS.n5695 DVSS.n109 0.00334
R20401 DVSS.n5696 DVSS.n5695 0.00334
R20402 DVSS.n5698 DVSS.n5696 0.00334
R20403 DVSS.n5698 DVSS.n5697 0.00334
R20404 DVSS.n5697 DVSS.n42 0.00334
R20405 DVSS.n5762 DVSS.n38 0.00334
R20406 DVSS.n5768 DVSS.n38 0.00334
R20407 DVSS.n5769 DVSS.n5768 0.00334
R20408 DVSS.n5770 DVSS.n5769 0.00334
R20409 DVSS.n5770 DVSS.n34 0.00334
R20410 DVSS.n5776 DVSS.n34 0.00334
R20411 DVSS.n5777 DVSS.n5776 0.00334
R20412 DVSS.n5778 DVSS.n5777 0.00334
R20413 DVSS.n5778 DVSS.n30 0.00334
R20414 DVSS.n5784 DVSS.n30 0.00334
R20415 DVSS.n5785 DVSS.n5784 0.00334
R20416 DVSS.n5791 DVSS.n28 0.00334
R20417 DVSS.n422 DVSS.n371 0.00334
R20418 DVSS.n422 DVSS.n421 0.00334
R20419 DVSS.n421 DVSS.n420 0.00334
R20420 DVSS.n420 DVSS.n372 0.00334
R20421 DVSS.n416 DVSS.n372 0.00334
R20422 DVSS.n416 DVSS.n415 0.00334
R20423 DVSS.n415 DVSS.n414 0.00334
R20424 DVSS.n414 DVSS.n378 0.00334
R20425 DVSS.n410 DVSS.n378 0.00334
R20426 DVSS.n410 DVSS.n409 0.00334
R20427 DVSS.n409 DVSS.n408 0.00334
R20428 DVSS.n408 DVSS.n384 0.00334
R20429 DVSS.n404 DVSS.n384 0.00334
R20430 DVSS.n404 DVSS.n403 0.00334
R20431 DVSS.n403 DVSS.n402 0.00334
R20432 DVSS.n402 DVSS.n390 0.00334
R20433 DVSS.n398 DVSS.n390 0.00334
R20434 DVSS.n398 DVSS.n397 0.00334
R20435 DVSS.n397 DVSS.n199 0.00334
R20436 DVSS.n616 DVSS.n199 0.00334
R20437 DVSS.n616 DVSS.n615 0.00334
R20438 DVSS.n615 DVSS.n614 0.00334
R20439 DVSS.n614 DVSS.n200 0.00334
R20440 DVSS.n609 DVSS.n608 0.00334
R20441 DVSS.n608 DVSS.n607 0.00334
R20442 DVSS.n607 DVSS.n580 0.00334
R20443 DVSS.n603 DVSS.n580 0.00334
R20444 DVSS.n603 DVSS.n602 0.00334
R20445 DVSS.n602 DVSS.n601 0.00334
R20446 DVSS.n601 DVSS.n586 0.00334
R20447 DVSS.n597 DVSS.n586 0.00334
R20448 DVSS.n597 DVSS.n596 0.00334
R20449 DVSS.n596 DVSS.n595 0.00334
R20450 DVSS.n595 DVSS.n166 0.00334
R20451 DVSS.n692 DVSS.n166 0.00334
R20452 DVSS.n693 DVSS.n692 0.00334
R20453 DVSS.n694 DVSS.n693 0.00334
R20454 DVSS.n694 DVSS.n162 0.00334
R20455 DVSS.n700 DVSS.n162 0.00334
R20456 DVSS.n701 DVSS.n700 0.00334
R20457 DVSS.n702 DVSS.n701 0.00334
R20458 DVSS.n702 DVSS.n158 0.00334
R20459 DVSS.n708 DVSS.n158 0.00334
R20460 DVSS.n709 DVSS.n708 0.00334
R20461 DVSS.n711 DVSS.n709 0.00334
R20462 DVSS.n711 DVSS.n710 0.00334
R20463 DVSS.n5648 DVSS.n5647 0.00334
R20464 DVSS.n5647 DVSS.n5646 0.00334
R20465 DVSS.n5646 DVSS.n137 0.00334
R20466 DVSS.n5642 DVSS.n137 0.00334
R20467 DVSS.n5642 DVSS.n5641 0.00334
R20468 DVSS.n5641 DVSS.n5640 0.00334
R20469 DVSS.n5640 DVSS.n143 0.00334
R20470 DVSS.n5636 DVSS.n143 0.00334
R20471 DVSS.n5636 DVSS.n5635 0.00334
R20472 DVSS.n5635 DVSS.n5634 0.00334
R20473 DVSS.n5634 DVSS.n5607 0.00334
R20474 DVSS.n5630 DVSS.n5607 0.00334
R20475 DVSS.n5630 DVSS.n5629 0.00334
R20476 DVSS.n5629 DVSS.n5628 0.00334
R20477 DVSS.n5628 DVSS.n5613 0.00334
R20478 DVSS.n5624 DVSS.n5613 0.00334
R20479 DVSS.n5624 DVSS.n5623 0.00334
R20480 DVSS.n5623 DVSS.n5622 0.00334
R20481 DVSS.n5622 DVSS.n51 0.00334
R20482 DVSS.n5719 DVSS.n51 0.00334
R20483 DVSS.n5720 DVSS.n5719 0.00334
R20484 DVSS.n5721 DVSS.n5720 0.00334
R20485 DVSS.n5721 DVSS.n44 0.00334
R20486 DVSS.n5759 DVSS.n45 0.00334
R20487 DVSS.n5755 DVSS.n45 0.00334
R20488 DVSS.n5755 DVSS.n5754 0.00334
R20489 DVSS.n5754 DVSS.n5753 0.00334
R20490 DVSS.n5753 DVSS.n5730 0.00334
R20491 DVSS.n5749 DVSS.n5730 0.00334
R20492 DVSS.n5749 DVSS.n5748 0.00334
R20493 DVSS.n5748 DVSS.n5747 0.00334
R20494 DVSS.n5747 DVSS.n5736 0.00334
R20495 DVSS.n5743 DVSS.n5736 0.00334
R20496 DVSS.n5743 DVSS.n5742 0.00334
R20497 DVSS.n5800 DVSS.n5799 0.00334
R20498 DVSS.n368 DVSS.n226 0.00334
R20499 DVSS.n467 DVSS.n226 0.00334
R20500 DVSS.n468 DVSS.n467 0.00334
R20501 DVSS.n469 DVSS.n468 0.00334
R20502 DVSS.n469 DVSS.n222 0.00334
R20503 DVSS.n475 DVSS.n222 0.00334
R20504 DVSS.n476 DVSS.n475 0.00334
R20505 DVSS.n477 DVSS.n476 0.00334
R20506 DVSS.n477 DVSS.n218 0.00334
R20507 DVSS.n483 DVSS.n218 0.00334
R20508 DVSS.n484 DVSS.n483 0.00334
R20509 DVSS.n485 DVSS.n484 0.00334
R20510 DVSS.n485 DVSS.n214 0.00334
R20511 DVSS.n491 DVSS.n214 0.00334
R20512 DVSS.n492 DVSS.n491 0.00334
R20513 DVSS.n493 DVSS.n492 0.00334
R20514 DVSS.n493 DVSS.n210 0.00334
R20515 DVSS.n500 DVSS.n210 0.00334
R20516 DVSS.n501 DVSS.n500 0.00334
R20517 DVSS.n503 DVSS.n501 0.00334
R20518 DVSS.n503 DVSS.n502 0.00334
R20519 DVSS.n502 DVSS.n207 0.00334
R20520 DVSS.n510 DVSS.n207 0.00334
R20521 DVSS.n573 DVSS.n572 0.00334
R20522 DVSS.n572 DVSS.n571 0.00334
R20523 DVSS.n571 DVSS.n512 0.00334
R20524 DVSS.n567 DVSS.n512 0.00334
R20525 DVSS.n567 DVSS.n566 0.00334
R20526 DVSS.n566 DVSS.n565 0.00334
R20527 DVSS.n565 DVSS.n517 0.00334
R20528 DVSS.n561 DVSS.n517 0.00334
R20529 DVSS.n561 DVSS.n560 0.00334
R20530 DVSS.n560 DVSS.n559 0.00334
R20531 DVSS.n559 DVSS.n523 0.00334
R20532 DVSS.n555 DVSS.n523 0.00334
R20533 DVSS.n555 DVSS.n554 0.00334
R20534 DVSS.n554 DVSS.n553 0.00334
R20535 DVSS.n553 DVSS.n529 0.00334
R20536 DVSS.n549 DVSS.n529 0.00334
R20537 DVSS.n549 DVSS.n548 0.00334
R20538 DVSS.n548 DVSS.n547 0.00334
R20539 DVSS.n547 DVSS.n535 0.00334
R20540 DVSS.n543 DVSS.n535 0.00334
R20541 DVSS.n543 DVSS.n542 0.00334
R20542 DVSS.n542 DVSS.n152 0.00334
R20543 DVSS.n719 DVSS.n152 0.00334
R20544 DVSS.n722 DVSS.n721 0.00334
R20545 DVSS.n722 DVSS.n148 0.00334
R20546 DVSS.n728 DVSS.n148 0.00334
R20547 DVSS.n729 DVSS.n728 0.00334
R20548 DVSS.n5596 DVSS.n729 0.00334
R20549 DVSS.n5596 DVSS.n5595 0.00334
R20550 DVSS.n5595 DVSS.n5594 0.00334
R20551 DVSS.n5594 DVSS.n730 0.00334
R20552 DVSS.n5590 DVSS.n730 0.00334
R20553 DVSS.n5590 DVSS.n5589 0.00334
R20554 DVSS.n5589 DVSS.n5588 0.00334
R20555 DVSS.n5588 DVSS.n735 0.00334
R20556 DVSS.n5584 DVSS.n735 0.00334
R20557 DVSS.n5584 DVSS.n5583 0.00334
R20558 DVSS.n5583 DVSS.n5582 0.00334
R20559 DVSS.n5582 DVSS.n741 0.00334
R20560 DVSS.n5578 DVSS.n741 0.00334
R20561 DVSS.n5578 DVSS.n5577 0.00334
R20562 DVSS.n5577 DVSS.n5576 0.00334
R20563 DVSS.n5576 DVSS.n747 0.00334
R20564 DVSS.n5572 DVSS.n747 0.00334
R20565 DVSS.n5572 DVSS.n5571 0.00334
R20566 DVSS.n5571 DVSS.n5570 0.00334
R20567 DVSS.n5566 DVSS.n5565 0.00334
R20568 DVSS.n5565 DVSS.n5564 0.00334
R20569 DVSS.n5564 DVSS.n808 0.00334
R20570 DVSS.n5560 DVSS.n808 0.00334
R20571 DVSS.n5560 DVSS.n5559 0.00334
R20572 DVSS.n5559 DVSS.n5558 0.00334
R20573 DVSS.n5558 DVSS.n814 0.00334
R20574 DVSS.n5554 DVSS.n814 0.00334
R20575 DVSS.n5554 DVSS.n5553 0.00334
R20576 DVSS.n5553 DVSS.n5552 0.00334
R20577 DVSS.n5552 DVSS.n820 0.00334
R20578 DVSS.n5548 DVSS.n5547 0.00334
R20579 DVSS.n1980 DVSS.n1979 0.00334
R20580 DVSS.n1983 DVSS.n1980 0.00334
R20581 DVSS.n1984 DVSS.n1983 0.00334
R20582 DVSS.n1985 DVSS.n1984 0.00334
R20583 DVSS.n1986 DVSS.n1985 0.00334
R20584 DVSS.n1990 DVSS.n1986 0.00334
R20585 DVSS.n1991 DVSS.n1990 0.00334
R20586 DVSS.n1992 DVSS.n1991 0.00334
R20587 DVSS.n1993 DVSS.n1992 0.00334
R20588 DVSS.n1994 DVSS.n1993 0.00334
R20589 DVSS.n1994 DVSS.n1495 0.00334
R20590 DVSS.n4189 DVSS.n1495 0.00334
R20591 DVSS.n4190 DVSS.n4189 0.00334
R20592 DVSS.n4191 DVSS.n4190 0.00334
R20593 DVSS.n4191 DVSS.n1491 0.00334
R20594 DVSS.n4197 DVSS.n1491 0.00334
R20595 DVSS.n4198 DVSS.n4197 0.00334
R20596 DVSS.n4199 DVSS.n4198 0.00334
R20597 DVSS.n4199 DVSS.n1487 0.00334
R20598 DVSS.n4205 DVSS.n1487 0.00334
R20599 DVSS.n4206 DVSS.n4205 0.00334
R20600 DVSS.n4207 DVSS.n4206 0.00334
R20601 DVSS.n4208 DVSS.n4207 0.00334
R20602 DVSS.n4209 DVSS.n4208 0.00334
R20603 DVSS.n4212 DVSS.n4209 0.00334
R20604 DVSS.n4213 DVSS.n4212 0.00334
R20605 DVSS.n4214 DVSS.n4213 0.00334
R20606 DVSS.n4215 DVSS.n4214 0.00334
R20607 DVSS.n4218 DVSS.n4215 0.00334
R20608 DVSS.n4219 DVSS.n4218 0.00334
R20609 DVSS.n4220 DVSS.n4219 0.00334
R20610 DVSS.n4221 DVSS.n4220 0.00334
R20611 DVSS.n4224 DVSS.n4221 0.00334
R20612 DVSS.n4225 DVSS.n4224 0.00334
R20613 DVSS.n4226 DVSS.n4225 0.00334
R20614 DVSS.n4227 DVSS.n4226 0.00334
R20615 DVSS.n4230 DVSS.n4227 0.00334
R20616 DVSS.n4231 DVSS.n4230 0.00334
R20617 DVSS.n4232 DVSS.n4231 0.00334
R20618 DVSS.n4233 DVSS.n4232 0.00334
R20619 DVSS.n4236 DVSS.n4233 0.00334
R20620 DVSS.n4237 DVSS.n4236 0.00334
R20621 DVSS.n4238 DVSS.n4237 0.00334
R20622 DVSS.n4239 DVSS.n4238 0.00334
R20623 DVSS.n4241 DVSS.n4239 0.00334
R20624 DVSS.n4243 DVSS.n4241 0.00334
R20625 DVSS.n4243 DVSS.n4242 0.00334
R20626 DVSS.n4242 DVSS.n1238 0.00334
R20627 DVSS.n1239 DVSS.n1238 0.00334
R20628 DVSS.n1240 DVSS.n1239 0.00334
R20629 DVSS.n1243 DVSS.n1240 0.00334
R20630 DVSS.n1244 DVSS.n1243 0.00334
R20631 DVSS.n1245 DVSS.n1244 0.00334
R20632 DVSS.n1246 DVSS.n1245 0.00334
R20633 DVSS.n1299 DVSS.n1246 0.00334
R20634 DVSS.n1300 DVSS.n1299 0.00334
R20635 DVSS.n1300 DVSS.n1297 0.00334
R20636 DVSS.n1306 DVSS.n1297 0.00334
R20637 DVSS.n1307 DVSS.n1306 0.00334
R20638 DVSS.n1308 DVSS.n1307 0.00334
R20639 DVSS.n1308 DVSS.n1293 0.00334
R20640 DVSS.n1315 DVSS.n1293 0.00334
R20641 DVSS.n1316 DVSS.n1315 0.00334
R20642 DVSS.n1317 DVSS.n1316 0.00334
R20643 DVSS.n1317 DVSS.n1289 0.00334
R20644 DVSS.n1323 DVSS.n1289 0.00334
R20645 DVSS.n1324 DVSS.n1323 0.00334
R20646 DVSS.n1325 DVSS.n1324 0.00334
R20647 DVSS.n1325 DVSS.n1285 0.00334
R20648 DVSS.n1331 DVSS.n1285 0.00334
R20649 DVSS.n1332 DVSS.n1331 0.00334
R20650 DVSS.n1333 DVSS.n1332 0.00334
R20651 DVSS.n1333 DVSS.n1281 0.00334
R20652 DVSS.n1339 DVSS.n1281 0.00334
R20653 DVSS.n1340 DVSS.n1339 0.00334
R20654 DVSS.n1341 DVSS.n1340 0.00334
R20655 DVSS.n1353 DVSS.n1352 0.00334
R20656 DVSS.n4544 DVSS.n1429 0.00332857
R20657 DVSS.n4546 DVSS.n4545 0.00332857
R20658 DVSS.n4555 DVSS.n1426 0.00332857
R20659 DVSS.n4554 DVSS.n1420 0.00332857
R20660 DVSS.n4563 DVSS.n4562 0.00332857
R20661 DVSS.n1421 DVSS.n1416 0.00332857
R20662 DVSS.n4569 DVSS.n4568 0.00332857
R20663 DVSS.n1160 DVSS.n1156 0.00332857
R20664 DVSS.n362 DVSS.n361 0.00332
R20665 DVSS.n363 DVSS.n243 0.00332
R20666 DVSS.n366 DVSS.n364 0.00332
R20667 DVSS.n367 DVSS.n250 0.00332
R20668 DVSS.n253 DVSS.n245 0.00332
R20669 DVSS.n360 DVSS.n254 0.00332
R20670 DVSS.n1388 DVSS.n1364 0.00330488
R20671 DVSS.n1373 DVSS.n1359 0.00330488
R20672 DVSS.n687 DVSS.n170 0.00329
R20673 DVSS.n689 DVSS.n168 0.00329
R20674 DVSS.n526 DVSS.n169 0.00329
R20675 DVSS.n5548 DVSS 0.00326
R20676 DVSS.n1352 DVSS 0.00326
R20677 DVSS.n2017 DVSS.n1971 0.0032
R20678 DVSS.n4059 DVSS.n1610 0.0032
R20679 DVSS.n5715 DVSS.n55 0.00319327
R20680 DVSS.n1538 DVSS.n1530 0.00319022
R20681 DVSS.n4157 DVSS.n4156 0.00319022
R20682 DVSS.n4116 VSS 0.00314706
R20683 VSS DVSS.n1550 0.00314706
R20684 DVSS.n463 DVSS.n229 0.00314706
R20685 DVSS.n4040 DVSS.n4039 0.00313571
R20686 DVSS.n1646 DVSS.n1642 0.00313571
R20687 DVSS.n311 DVSS.n258 0.00311
R20688 DVSS.n373 DVSS.n244 0.00311
R20689 DVSS.n465 DVSS.n464 0.00311
R20690 DVSS.n4774 DVSS.n4773 0.00309529
R20691 DVSS.n1661 DVSS.n1657 0.00307143
R20692 DVSS.n3995 DVSS.n1662 0.00307143
R20693 DVSS.n3994 DVSS.n3982 0.00307143
R20694 DVSS.n5345 DVSS.n951 0.00300714
R20695 DVSS.n4681 DVSS.n1354 0.00300714
R20696 DVSS.n4048 DVSS.n1627 0.00300714
R20697 DVSS.n3396 DVSS.n2819 0.003
R20698 DVSS.n3372 DVSS.n2853 0.003
R20699 DVSS.n3133 DVSS.n3132 0.003
R20700 DVSS.n3160 DVSS.n2851 0.003
R20701 DVSS.n1942 DVSS.n1934 0.00297706
R20702 DVSS.n2669 DVSS.n2667 0.00296479
R20703 DVSS.n3502 DVSS.n2670 0.00296479
R20704 DVSS.n3028 DVSS.n2677 0.00296479
R20705 DVSS.n3494 DVSS.n3493 0.00296479
R20706 DVSS.n3490 DVSS.n2679 0.00296479
R20707 DVSS.n3489 DVSS.n2690 0.00296479
R20708 DVSS.n3039 DVSS.n2697 0.00296479
R20709 DVSS.n3482 DVSS.n3481 0.00296479
R20710 DVSS.n3478 DVSS.n2699 0.00296479
R20711 DVSS.n3477 DVSS.n2707 0.00296479
R20712 DVSS.n3051 DVSS.n2715 0.00296479
R20713 DVSS.n3470 DVSS.n3469 0.00296479
R20714 DVSS.n3466 DVSS.n2717 0.00296479
R20715 DVSS.n3465 DVSS.n2725 0.00296479
R20716 DVSS.n3070 DVSS.n3065 0.00296479
R20717 DVSS.n3071 DVSS.n2735 0.00296479
R20718 DVSS.n3454 DVSS.n3453 0.00296479
R20719 DVSS.n3450 DVSS.n2737 0.00296479
R20720 DVSS.n3449 DVSS.n2743 0.00296479
R20721 DVSS.n3082 DVSS.n2750 0.00296479
R20722 DVSS.n3442 DVSS.n3441 0.00296479
R20723 DVSS.n3438 DVSS.n2752 0.00296479
R20724 DVSS.n3437 DVSS.n2760 0.00296479
R20725 DVSS.n3095 DVSS.n2770 0.00296479
R20726 DVSS.n3430 DVSS.n3429 0.00296479
R20727 DVSS.n3426 DVSS.n2772 0.00296479
R20728 DVSS.n3425 DVSS.n2780 0.00296479
R20729 DVSS.n3106 DVSS.n2787 0.00296479
R20730 DVSS.n3418 DVSS.n3417 0.00296479
R20731 DVSS.n3414 DVSS.n2789 0.00296479
R20732 DVSS.n3413 DVSS.n2797 0.00296479
R20733 DVSS.n3119 DVSS.n2806 0.00296479
R20734 DVSS.n3406 DVSS.n3405 0.00296479
R20735 DVSS.n3402 DVSS.n2808 0.00296479
R20736 DVSS.n3401 DVSS.n2816 0.00296479
R20737 DVSS.n3139 DVSS.n3134 0.00296479
R20738 DVSS.n3140 DVSS.n2827 0.00296479
R20739 DVSS.n3390 DVSS.n3389 0.00296479
R20740 DVSS.n3386 DVSS.n2829 0.00296479
R20741 DVSS.n3385 DVSS.n2835 0.00296479
R20742 DVSS.n3151 DVSS.n2842 0.00296479
R20743 DVSS.n3378 DVSS.n3377 0.00296479
R20744 DVSS.n3374 DVSS.n2844 0.00296479
R20745 DVSS.n3373 DVSS.n2852 0.00296479
R20746 DVSS.n3164 DVSS.n2862 0.00296479
R20747 DVSS.n3366 DVSS.n3365 0.00296479
R20748 DVSS.n3362 DVSS.n2864 0.00296479
R20749 DVSS.n3361 DVSS.n2872 0.00296479
R20750 DVSS.n3176 DVSS.n2880 0.00296479
R20751 DVSS.n3354 DVSS.n3353 0.00296479
R20752 DVSS.n3350 DVSS.n2882 0.00296479
R20753 DVSS.n3349 DVSS.n2890 0.00296479
R20754 DVSS.n3188 DVSS.n2898 0.00296479
R20755 DVSS.n3341 DVSS.n3340 0.00296479
R20756 DVSS.n3337 DVSS.n2900 0.00296479
R20757 DVSS.n3336 DVSS.n2908 0.00296479
R20758 DVSS.n3199 DVSS.n2916 0.00296479
R20759 DVSS.n3328 DVSS.n3327 0.00296479
R20760 DVSS.n3324 DVSS.n2918 0.00296479
R20761 DVSS.n3323 DVSS.n2926 0.00296479
R20762 DVSS.n3212 DVSS.n2933 0.00296479
R20763 DVSS.n3316 DVSS.n3315 0.00296479
R20764 DVSS.n3312 DVSS.n2935 0.00296479
R20765 DVSS.n3311 DVSS.n2943 0.00296479
R20766 DVSS.n3225 DVSS.n2952 0.00296479
R20767 DVSS.n3303 DVSS.n3302 0.00296479
R20768 DVSS.n3299 DVSS.n2954 0.00296479
R20769 DVSS.n3298 DVSS.n2962 0.00296479
R20770 DVSS.n3236 DVSS.n2969 0.00296479
R20771 DVSS.n3290 DVSS.n3289 0.00296479
R20772 DVSS.n3286 DVSS.n2971 0.00296479
R20773 DVSS.n3285 DVSS.n2979 0.00296479
R20774 DVSS.n3247 DVSS.n2987 0.00296479
R20775 DVSS.n3278 DVSS.n3277 0.00296479
R20776 DVSS.n3274 DVSS.n2989 0.00296479
R20777 DVSS.n3273 DVSS.n2998 0.00296479
R20778 DVSS.n3263 DVSS.n3262 0.00296479
R20779 DVSS.n3830 DVSS.n1787 0.00296479
R20780 DVSS.n3829 DVSS.n1783 0.00296479
R20781 DVSS.n426 DVSS.n242 0.00294344
R20782 DVSS.n3473 DVSS 0.00293842
R20783 DVSS DVSS.n3054 0.00293842
R20784 DVSS.n2495 DVSS.n2494 0.00293243
R20785 DVSS.n106 DVSS.n105 0.0029
R20786 DVSS.n5724 DVSS.n48 0.0029
R20787 DVSS.n805 DVSS.n804 0.0029
R20788 DVSS.n4316 DVSS 0.00286842
R20789 DVSS.n4821 DVSS 0.00286842
R20790 DVSS.n1226 DVSS 0.00286842
R20791 VSS DVSS.n1513 0.00286842
R20792 DVSS.n4779 DVSS 0.00286842
R20793 DVSS.n5762 DVSS.n5761 0.00286
R20794 DVSS.n5760 DVSS.n5759 0.00286
R20795 DVSS.n5566 DVSS.n43 0.00286
R20796 DVSS DVSS.n28 0.00282
R20797 DVSS.n1341 DVSS 0.00278
R20798 DVSS.n3394 DVSS.n2824 0.00271675
R20799 DVSS.n3129 DVSS.n3013 0.00271675
R20800 DVSS.n5655 DVSS.n5654 0.0027
R20801 DVSS.n5648 DVSS.n129 0.0027
R20802 DVSS.n721 DVSS.n720 0.0027
R20803 DVSS.n1311 DVSS.n1310 0.00269
R20804 DVSS.n4453 DVSS.n4452 0.00262143
R20805 DVSS.n4449 DVSS.n4446 0.00262143
R20806 DVSS.n4448 DVSS.n1446 0.00262143
R20807 DVSS.n4516 DVSS.n4515 0.00262143
R20808 DVSS.n4523 DVSS.n1441 0.00262143
R20809 DVSS.n4522 DVSS.n1442 0.00262143
R20810 DVSS.n4528 DVSS.n1437 0.00262143
R20811 DVSS.n4707 DVSS.n4640 0.00262143
R20812 DVSS.n4663 DVSS.n4662 0.00262143
R20813 DVSS.n4704 DVSS.n4703 0.00262143
R20814 DVSS.n1381 DVSS.n1366 0.00257317
R20815 DVSS.n1380 DVSS.n1361 0.00257317
R20816 DVSS.n2014 DVSS.n2013 0.00257
R20817 DVSS.n1312 DVSS.n1311 0.00257
R20818 DVSS.n2329 DVSS.n2321 0.00256422
R20819 DVSS.n1893 DVSS.n1892 0.00256422
R20820 DVSS.n4484 DVSS.n4414 0.00255714
R20821 DVSS.n4481 DVSS.n4480 0.00255714
R20822 DVSS.n4423 DVSS.n4417 0.00255714
R20823 DVSS.n4474 DVSS.n4424 0.00255714
R20824 DVSS.n4473 DVSS.n4425 0.00255714
R20825 DVSS.n4435 DVSS.n4434 0.00255714
R20826 DVSS.n4468 DVSS.n4467 0.00255714
R20827 DVSS.n634 DVSS.n633 0.00254
R20828 DVSS.n609 DVSS.n186 0.00254
R20829 DVSS.n573 DVSS.n511 0.00254
R20830 DVSS.n765 DVSS.n55 0.00251995
R20831 DVSS.n3395 DVSS.n2823 0.0025
R20832 DVSS.n2857 DVSS.n2856 0.0025
R20833 DVSS.n3141 DVSS.n3014 0.0025
R20834 DVSS.n3159 DVSS.n3012 0.0025
R20835 DVSS.n2557 DVSS.n1912 0.00249286
R20836 DVSS.n2532 DVSS.n1914 0.00249286
R20837 DVSS.n3852 DVSS 0.00247183
R20838 DVSS.n2264 DVSS.n2260 0.00242857
R20839 DVSS.n2261 DVSS.n1904 0.00242857
R20840 DVSS.n359 DVSS.n247 0.00238
R20841 DVSS.n371 DVSS.n370 0.00238
R20842 DVSS.n369 DVSS.n368 0.00238
R20843 DVSS.n3953 DVSS.n1687 0.00236429
R20844 DVSS.n105 DVSS.n103 0.00236
R20845 DVSS.n50 DVSS.n48 0.00236
R20846 DVSS.n804 DVSS.n753 0.00236
R20847 DVSS.n427 DVSS.n426 0.00233258
R20848 DVSS.n5535 DVSS 0.0023
R20849 DVSS DVSS.n4689 0.0023
R20850 DVSS.n4688 DVSS 0.0023
R20851 DVSS.n3745 VSS 0.0023
R20852 DVSS.n2409 DVSS 0.0023
R20853 DVSS.n2091 DVSS 0.0023
R20854 DVSS.n1763 DVSS 0.0023
R20855 DVSS.n4890 VSS 0.0023
R20856 DVSS.n4889 VSS 0.0023
R20857 VSS DVSS.n3527 0.0023
R20858 DVSS.n3346 DVSS.n3345 0.0022734
R20859 DVSS.n3186 DVSS.n3010 0.0022734
R20860 DVSS.n4895 DVSS.n1193 0.00223571
R20861 DVSS.n4885 DVSS.n4878 0.00223571
R20862 DVSS.n4889 DVSS.n4888 0.00223571
R20863 DVSS.n3759 DVSS.n3534 0.00223571
R20864 DVSS.n3756 DVSS.n3749 0.00223571
R20865 DVSS.n3761 DVSS.n3527 0.00223571
R20866 DVSS.n312 DVSS.n311 0.00215
R20867 DVSS.n374 DVSS.n373 0.00215
R20868 DVSS.n464 DVSS.n224 0.00215
R20869 DVSS.n2801 DVSS.n2800 0.002
R20870 DVSS.n3355 DVSS.n2879 0.002
R20871 DVSS.n3113 DVSS.n3112 0.002
R20872 DVSS.n3181 DVSS.n2881 0.002
R20873 DVSS.n3907 DVSS.n1735 0.00197857
R20874 DVSS.n687 DVSS.n686 0.00197
R20875 DVSS.n690 DVSS.n689 0.00197
R20876 DVSS.n527 DVSS.n169 0.00197
R20877 DVSS.n5742 DVSS 0.00196
R20878 DVSS.n5537 DVSS 0.00191429
R20879 DVSS.n5800 DVSS 0.00188
R20880 DVSS.n4032 DVSS.n4031 0.00185
R20881 DVSS.n4020 DVSS.n1647 0.00185
R20882 DVSS.n1389 DVSS.n1365 0.00184146
R20883 DVSS.n1372 DVSS.n1362 0.00184146
R20884 DVSS.n5740 DVSS 0.00173
R20885 DVSS DVSS.n0 0.00173
R20886 DVSS.n5534 DVSS 0.0017
R20887 DVSS.n4687 DVSS 0.0017
R20888 DVSS.n630 DVSS.n184 0.0017
R20889 DVSS.n577 DVSS.n202 0.0017
R20890 DVSS.n576 DVSS.n204 0.0017
R20891 DVSS.n509 DVSS.n203 0.0017
R20892 DVSS.n612 DVSS.n611 0.0017
R20893 DVSS.n631 DVSS.n185 0.0017
R20894 DVSS.n5701 DVSS.n5700 0.00167
R20895 DVSS.n5716 DVSS.n54 0.00167
R20896 DVSS.n801 DVSS.n751 0.00167
R20897 DVSS.n4682 DVSS.n1355 0.00165714
R20898 DVSS.n4678 DVSS.n1357 0.00165714
R20899 DVSS.n2503 DVSS.n1925 0.00165714
R20900 DVSS.n2475 DVSS.n1924 0.00165714
R20901 DVSS.n5045 DVSS.n1108 0.00165714
R20902 DVSS.n5043 DVSS.n5042 0.00165714
R20903 DVSS.n1116 DVSS.n1110 0.00165714
R20904 DVSS.n5036 DVSS.n1117 0.00165714
R20905 DVSS.n5035 DVSS.n1118 0.00165714
R20906 DVSS.n5032 DVSS.n5031 0.00165714
R20907 DVSS.n1126 DVSS.n1122 0.00165714
R20908 DVSS.n5025 DVSS.n1127 0.00165714
R20909 DVSS.n4585 DVSS.n1407 0.00159286
R20910 DVSS.n4584 DVSS.n1408 0.00159286
R20911 DVSS.n4591 DVSS.n1405 0.00159286
R20912 DVSS.n4593 DVSS.n4592 0.00159286
R20913 DVSS.n4749 DVSS.n1399 0.00159286
R20914 DVSS.n4748 DVSS.n1400 0.00159286
R20915 DVSS.n4602 DVSS.n4599 0.00159286
R20916 DVSS.n2249 DVSS.n1960 0.00159286
R20917 DVSS.n2226 DVSS.n1957 0.00159286
R20918 DVSS.n1965 DVSS.n1959 0.00159286
R20919 DVSS.n3958 DVSS.n1682 0.00159286
R20920 DVSS.n2253 DVSS.n1952 0.00157001
R20921 DVSS.n1937 DVSS.n1855 0.00152857
R20922 DVSS.n2599 DVSS.n1859 0.00152857
R20923 DVSS.n3436 DVSS.n2761 0.0015
R20924 DVSS.n3331 DVSS.n2911 0.0015
R20925 DVSS.n3091 DVSS.n2759 0.0015
R20926 DVSS.n3201 DVSS.n3200 0.0015
R20927 DVSS.n4282 DVSS.n1484 0.00146
R20928 DVSS.n155 DVSS.n132 0.00146
R20929 DVSS.n715 DVSS.n714 0.00146
R20930 DVSS.n717 DVSS.n716 0.00146
R20931 DVSS.n718 DVSS.n133 0.00146
R20932 DVSS.n5650 DVSS.n134 0.00146
R20933 DVSS.n5652 DVSS.n5651 0.00146
R20934 DVSS.n2855 DVSS.n2840 0.0013867
R20935 DVSS.n3157 DVSS.n3155 0.0013867
R20936 DVSS.n1350 DVSS 0.00134
R20937 DVSS.n1349 DVSS 0.00134
R20938 DVSS.n823 DVSS 0.00134
R20939 DVSS DVSS.n5550 0.00134
R20940 DVSS.n2148 DVSS.n1528 0.00133571
R20941 DVSS.n1529 DVSS.n1527 0.00133571
R20942 DVSS.n4155 DVSS.n1534 0.00133571
R20943 DVSS.n1656 DVSS.n1652 0.00133571
R20944 DVSS.n4791 DVSS.n4790 0.00131
R20945 DVSS.n1349 DVSS.n1348 0.00131
R20946 DVSS.n5660 DVSS.n123 0.00131
R20947 DVSS.n5601 DVSS.n141 0.00131
R20948 DVSS.n5599 DVSS.n144 0.00131
R20949 DVSS.n633 DVSS.n632 0.0013
R20950 DVSS.n200 DVSS.n186 0.0013
R20951 DVSS.n511 DVSS.n510 0.0013
R20952 DVSS.n106 DVSS.n40 0.00122
R20953 DVSS.n5725 DVSS.n5724 0.00122
R20954 DVSS.n805 DVSS.n47 0.00122
R20955 DVSS.n5569 DVSS.n5568 0.00122
R20956 DVSS.n5723 DVSS.n46 0.00122
R20957 DVSS.n107 DVSS.n41 0.00122
R20958 DVSS.n4770 DVSS 0.00120714
R20959 DVSS.n3930 DVSS.n1707 0.00120714
R20960 DVSS.n1726 DVSS.n1722 0.00120714
R20961 DVSS.n5062 DVSS.n5061 0.00120714
R20962 DVSS.n1103 DVSS.n1099 0.00120714
R20963 DVSS.n2003 DVSS.n1988 0.00119
R20964 DVSS.n4186 DVSS.n1497 0.00119
R20965 DVSS.n5654 DVSS.n5653 0.00114
R20966 DVSS.n710 DVSS.n129 0.00114
R20967 DVSS.n720 DVSS.n719 0.00114
R20968 DVSS.n4802 DVSS.n4801 0.00107
R20969 DVSS.n4777 DVSS.n4776 0.00107
R20970 DVSS.n1351 DVSS 0.00106
R20971 DVSS.n6 DVSS.n5 0.00104
R20972 DVSS.n5797 DVSS.n5796 0.00104
R20973 DVSS.n829 DVSS.n828 0.00104
R20974 DVSS.n5545 DVSS.n5544 0.00104
R20975 DVSS.n5785 DVSS 0.00102
R20976 DVSS.n622 DVSS.n621 0.00101
R20977 DVSS.n619 DVSS.n195 0.00101
R20978 DVSS.n497 DVSS.n194 0.00101
R20979 DVSS.n3501 DVSS.n3500 0.001
R20980 DVSS.n3459 DVSS.n2732 0.001
R20981 DVSS.n3310 DVSS.n3309 0.001
R20982 DVSS.n3267 DVSS.n1789 0.001
R20983 DVSS.n3503 DVSS.n2668 0.001
R20984 DVSS.n3072 DVSS.n3021 0.001
R20985 DVSS.n3223 DVSS.n2942 0.001
R20986 DVSS.n3003 DVSS.n3002 0.001
R20987 DVSS.n5761 DVSS.n42 0.00098
R20988 DVSS.n5760 DVSS.n44 0.00098
R20989 DVSS.n5570 DVSS.n43 0.00098
R20990 DVSS.n1632 DVSS.n1631 0.00095
R20991 DVSS.n2877 DVSS.n2876 0.00094335
R20992 DVSS.n3173 DVSS.n3172 0.00094335
R20993 DVSS.n257 DVSS.n252 0.00092
R20994 DVSS.n425 DVSS.n424 0.00092
R20995 DVSS.n365 DVSS.n228 0.00092
R20996 DVSS.n5537 DVSS.n5536 0.000885714
R20997 DVSS.n2232 DVSS.n2227 0.000856671
R20998 DVSS.n2241 DVSS.n1962 0.000856671
R20999 DVSS.n2673 DVSS 0.000721675
R21000 DVSS DVSS.n3505 0.000721675
R21001 DVSS.n3851 DVSS 0.000687793
R21002 DVSS.n5787 DVSS 0.00068
R21003 DVSS.n5786 DVSS 0.00068
R21004 DVSS.n5534 DVSS 0.000671429
R21005 DVSS.n4687 DVSS 0.000671429
R21006 DVSS.n3746 VSS 0.000671429
R21007 DVSS.n2408 DVSS 0.000671429
R21008 DVSS DVSS.n2090 0.000671429
R21009 DVSS.n1764 DVSS 0.000671429
R21010 DVSS.n4891 VSS 0.000671429
R21011 DVSS.n1938 DVSS.n1937 0.000628571
R21012 DVSS.n2599 DVSS.n2598 0.000628571
R21013 DVSS.n2279 DVSS.n1860 0.000628571
R21014 DVSS.n2286 DVSS.n2280 0.000628571
R21015 DVSS.n2285 DVSS.n2278 0.000628571
R21016 DVSS.n2288 DVSS.n2275 0.000628571
R21017 DVSS.n2289 DVSS.n1874 0.000628571
R21018 DVSS.n2271 DVSS.n1876 0.000628571
R21019 DVSS.n2295 DVSS.n1873 0.000628571
R21020 DVSS.n2584 DVSS.n1877 0.000628571
R21021 DVSS.n2582 DVSS.n1878 0.000628571
R21022 DVSS.n1885 DVSS.n1884 0.000628571
R21023 DVSS.n2576 DVSS.n2575 0.000628571
R21024 DVSS.n2257 DVSS.n1886 0.000628571
R21025 DVSS.n2260 DVSS.n1902 0.000628571
R21026 DVSS.n2566 DVSS.n1904 0.000628571
R21027 DVSS.n2558 DVSS.n2557 0.000628571
R21028 DVSS.n1914 DVSS.n1913 0.000628571
R21029 DVSS.n2531 DVSS.n2313 0.000628571
R21030 DVSS.n2318 DVSS.n2317 0.000628571
R21031 DVSS.n2525 DVSS.n2524 0.000628571
R21032 DVSS.n2349 DVSS.n2319 0.000628571
R21033 DVSS.n2368 DVSS.n2350 0.000628571
R21034 DVSS.n2353 DVSS.n2347 0.000628571
R21035 DVSS.n2360 DVSS.n2348 0.000628571
R21036 DVSS.n2370 DVSS.n2345 0.000628571
R21037 DVSS.n2372 DVSS.n2371 0.000628571
R21038 DVSS.n2511 DVSS.n2339 0.000628571
R21039 DVSS.n2510 DVSS.n2340 0.000628571
R21040 DVSS.n2472 DVSS.n2471 0.000628571
R21041 DVSS.n2504 DVSS.n2503 0.000628571
R21042 DVSS.n2475 DVSS.n2474 0.000628571
R21043 DVSS DVSS.n820 0.00058
R21044 DVSS DVSS.n1351 0.00058
R21045 DVSS.n3865 DVSS.n1778 0.000570422
R21046 DVSS.n5341 DVSS.n957 0.000566519
R21047 DVSS.n3867 DVSS.n3866 0.000564286
R21048 GF_NI_IN_C_BASE_0.comp018green_esd_cdm_0.IP_IN.n0 GF_NI_IN_C_BASE_0.comp018green_esd_cdm_0.IP_IN.t7 30.5934
R21049 GF_NI_IN_C_BASE_0.comp018green_esd_cdm_0.IP_IN.n0 GF_NI_IN_C_BASE_0.comp018green_esd_cdm_0.IP_IN.t6 30.5934
R21050 GF_NI_IN_C_BASE_0.comp018green_esd_cdm_0.IP_IN.n0 GF_NI_IN_C_BASE_0.comp018green_esd_cdm_0.IP_IN.t3 30.5934
R21051 GF_NI_IN_C_BASE_0.comp018green_esd_cdm_0.IP_IN.n0 GF_NI_IN_C_BASE_0.comp018green_esd_cdm_0.IP_IN.t1 30.5934
R21052 GF_NI_IN_C_BASE_0.comp018green_esd_cdm_0.IP_IN.n0 GF_NI_IN_C_BASE_0.comp018green_esd_cdm_0.IP_IN.t4 29.0913
R21053 GF_NI_IN_C_BASE_0.comp018green_esd_cdm_0.IP_IN.n0 GF_NI_IN_C_BASE_0.comp018green_esd_cdm_0.IP_IN.t12 28.7684
R21054 GF_NI_IN_C_BASE_0.comp018green_esd_cdm_0.IP_IN.n0 GF_NI_IN_C_BASE_0.comp018green_esd_cdm_0.IP_IN.t11 28.7684
R21055 GF_NI_IN_C_BASE_0.comp018green_esd_cdm_0.IP_IN.n0 GF_NI_IN_C_BASE_0.comp018green_esd_cdm_0.IP_IN.t2 28.7684
R21056 GF_NI_IN_C_BASE_0.comp018green_esd_cdm_0.IP_IN.n0 GF_NI_IN_C_BASE_0.comp018green_esd_cdm_0.IP_IN.t5 15.5342
R21057 GF_NI_IN_C_BASE_0.comp018green_esd_cdm_0.IP_IN.n0 GF_NI_IN_C_BASE_0.comp018green_esd_cdm_0.IP_IN.t8 15.2112
R21058 GF_NI_IN_C_BASE_0.comp018green_esd_cdm_0.IP_IN.n0 GF_NI_IN_C_BASE_0.comp018green_esd_cdm_0.IP_IN.t10 14.2306
R21059 GF_NI_IN_C_BASE_0.comp018green_esd_cdm_0.IP_IN.n0 GF_NI_IN_C_BASE_0.comp018green_esd_cdm_0.IP_IN.t9 13.9076
R21060 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_pupd_0.ppolyf_u_CDNS_4066195314532_0.PLUS GF_NI_IN_C_BASE_0.comp018green_esd_cdm_0.IP_IN.n0 13.3452
R21061 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_pupd_0.ppolyf_u_CDNS_4066195314532_0.PLUS GF_NI_IN_C_BASE_0.comp018green_esd_cdm_0.IP_IN.t0 11.0117
R21062 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_drv_0.A GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_drv_0.A.t11 39.4055
R21063 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_drv_0.A.n3 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_drv_0.A.t10 35.4055
R21064 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_drv_0.A.n3 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_drv_0.A.t9 34.8841
R21065 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_drv_0.A.t0 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_drv_0.A.n1 4.05527
R21066 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_drv_0.A.t1 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_drv_0.A.n1 4.06684
R21067 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_drv_0.A.n0 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_drv_0.A.n4 6.3635
R21068 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_drv_0.A.n2 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_drv_0.A.t8 2.10166
R21069 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_drv_0.A GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_drv_0.A.n0 5.38559
R21070 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_drv_0.A.n5 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_drv_0.A.t7 4.06578
R21071 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_drv_0.A GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_drv_0.A.n3 4.0005
R21072 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_drv_0.A.n4 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_drv_0.A.t3 3.98107
R21073 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_drv_0.A.n5 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_drv_0.A 3.16412
R21074 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_drv_0.A.n4 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_drv_0.A.t2 2.94036
R21075 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_drv_0.A.n0 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_drv_0.A 2.90177
R21076 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_drv_0.A.t4 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_drv_0.A.n2 2.10189
R21077 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_drv_0.A.n1 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_drv_0.A.n2 2.7349
R21078 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_drv_0.A.n0 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_drv_0.A.n1 2.2505
R21079 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_drv_0.A.n0 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_drv_0.A.n5 2.2505
R21080 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_drv_0.A GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_drv_0.A.t5 1.57941
R21081 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_drv_0.A GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_drv_0.A.t6 1.57897
R21082 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_cms_smt_0.nmos_6p0_CDNS_4066195314540_0.S GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_cms_smt_0.nmos_6p0_CDNS_4066195314540_0.S.t0 6.51577
R21083 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_cms_smt_0.nmos_6p0_CDNS_4066195314540_0.S.t6 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_cms_smt_0.nmos_6p0_CDNS_4066195314540_0.S 3.11732
R21084 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_cms_smt_0.nmos_6p0_CDNS_4066195314540_0.S GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_cms_smt_0.nmos_6p0_CDNS_4066195314540_0.S.t6 2.17664
R21085 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_cms_smt_0.nmos_6p0_CDNS_4066195314540_0.S GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_cms_smt_0.nmos_6p0_CDNS_4066195314540_0.S.t5 1.85326
R21086 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_cms_smt_0.nmos_6p0_CDNS_4066195314540_0.S GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_cms_smt_0.nmos_6p0_CDNS_4066195314540_0.S.t1 1.57786
R21087 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_cms_smt_0.nmos_6p0_CDNS_4066195314540_0.S GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_cms_smt_0.nmos_6p0_CDNS_4066195314540_0.S.t3 1.56968
R21088 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_cms_smt_0.nmos_6p0_CDNS_4066195314540_0.S GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_cms_smt_0.nmos_6p0_CDNS_4066195314540_0.S.t4 1.23514
R21089 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_cms_smt_0.nmos_6p0_CDNS_4066195314540_0.S GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_cms_smt_0.nmos_6p0_CDNS_4066195314540_0.S.t2 1.02385
R21090 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_logic_pupd_0.comp018green_std_xor2_0.nmos_6p0_CDNS_4066195314530_0.D.t0 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_logic_pupd_0.comp018green_std_xor2_0.nmos_6p0_CDNS_4066195314530_0.D.t2 33.2287
R21091 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_logic_pupd_0.comp018green_std_xor2_0.nmos_6p0_CDNS_4066195314530_0.D.t0 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_logic_pupd_0.comp018green_std_xor2_0.nmos_6p0_CDNS_4066195314530_0.D.t1 25.193
R21092 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_logic_pupd_0.comp018green_std_nand2_0.A.n1 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_logic_pupd_0.comp018green_std_nand2_0.A.t2 35.5619
R21093 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_logic_pupd_0.comp018green_std_nand2_0.A.n0 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_logic_pupd_0.comp018green_std_nand2_0.A.t4 35.5619
R21094 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_logic_pupd_0.comp018green_std_nand2_0.A.n1 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_logic_pupd_0.comp018green_std_nand2_0.A.t3 34.9362
R21095 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_logic_pupd_0.comp018green_std_nand2_0.A.n0 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_logic_pupd_0.comp018green_std_nand2_0.A.t5 34.9362
R21096 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_logic_pupd_0.comp018green_std_xor2_0.Z GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_logic_pupd_0.comp018green_std_nand2_1.B 6.58393
R21097 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_logic_pupd_0.comp018green_std_nand2_1.B GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_logic_pupd_0.comp018green_std_nand2_0.A.n1 4.4005
R21098 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_logic_pupd_0.comp018green_std_nand2_1.B GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_logic_pupd_0.comp018green_std_nand2_0.A.n0 4.00161
R21099 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_logic_pupd_0.comp018green_std_xor2_0.Z GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_logic_pupd_0.comp018green_std_nand2_0.A.t0 3.08699
R21100 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_logic_pupd_0.comp018green_std_nand2_0.A.t1 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_logic_pupd_0.comp018green_std_xor2_0.Z 2.76118
R21101 PU.n3 PU.t2 40.5155
R21102 PU.n8 PU.n6 37.3205
R21103 PU.n0 PU.t3 35.5619
R21104 PU.n0 PU.t4 34.9362
R21105 PU.n3 PU.t5 26.3326
R21106 PU.n6 PU.n5 7.47146
R21107 PU.n1 PU.n0 4.00141
R21108 PU PU.n3 4.00106
R21109 PU.n2 PU.t1 3.17811
R21110 PU.n8 PU.n7 2.25122
R21111 PU PU.n8 1.98787
R21112 PU.n5 PU.t0 1.36552
R21113 PU.n7 PU.t6 1.31518
R21114 PU.n5 PU.n4 0.80237
R21115 PU.n4 PU.n2 0.45653
R21116 PU.n4 PU 0.163278
R21117 PU.n6 PU.n1 0.127056
R21118 PU.n2 PU 0.0456808
R21119 PU.n1 PU 0.00756793
R21120 PU.n7 PU 0.001225
R21121 VSS.n3385 VSS.n3384 196056
R21122 VSS.n5277 VSS.n5276 37210.9
R21123 VSS.n5698 VSS.n11 32548.6
R21124 VSS.n5436 VSS.n5435 32385.4
R21125 VSS.n4085 VSS.n2203 30893.3
R21126 VSS.n5128 VSS.n2223 30469.2
R21127 VSS.n5678 VSS.n5677 27088.7
R21128 VSS.n5441 VSS.n1290 25861.7
R21129 VSS.n3405 VSS.n3385 21519.5
R21130 VSS.n5677 VSS.n5676 20471.6
R21131 VSS.n5281 VSS.n2200 19823.1
R21132 VSS.n5442 VSS.n5441 19552.7
R21133 VSS.n5291 VSS.n5290 17654
R21134 VSS.n5697 VSS.n12 16516.8
R21135 VSS.n2080 VSS.n1292 16516.8
R21136 VSS.n5291 VSS.n2187 16432
R21137 VSS.n3527 VSS.n2203 16400
R21138 VSS.n3528 VSS.n3526 16252.3
R21139 VSS.n5678 VSS.n12 16242.7
R21140 VSS.n1292 VSS.n1290 16242.7
R21141 VSS.n5304 VSS.n2187 16230.9
R21142 VSS.n5278 VSS.n2202 16230.9
R21143 VSS.n5292 VSS.n5291 16230.9
R21144 VSS.n5290 VSS.n2099 16230.9
R21145 VSS.n5422 VSS.n2091 16230.9
R21146 VSS.n4085 VSS.n2291 15030.2
R21147 VSS.n4292 VSS.n2291 14984.7
R21148 VSS.n3528 VSS.n3527 14824
R21149 VSS.n5281 VSS.n5280 14824
R21150 VSS.n5679 VSS.n5678 14769.2
R21151 VSS.n1290 VSS.n1172 14767.1
R21152 VSS.n5276 VSS.n2203 13915.8
R21153 VSS.n5127 VSS.n2287 12369.1
R21154 VSS.n5125 VSS.n2288 12369.1
R21155 VSS.n5123 VSS.n2289 12369.1
R21156 VSS.n5122 VSS.n2290 12369.1
R21157 VSS.n5129 VSS.n2237 11989.7
R21158 VSS.n5280 VSS.n5279 11473.2
R21159 VSS.n5279 VSS.n5278 10835.5
R21160 VSS.n5277 VSS.n2178 9379.2
R21161 VSS.n5278 VSS.n5277 8547.5
R21162 VSS.n4088 VSS.n4085 7940.47
R21163 VSS.n5435 VSS.n2081 7811.82
R21164 VSS.n3405 VSS.n3404 7328.63
R21165 VSS.n3526 VSS.n3525 6651.3
R21166 VSS.n5289 VSS.n5288 6538.35
R21167 VSS.n5123 VSS.n5122 6402.4
R21168 VSS.n5127 VSS.n5126 5994.44
R21169 VSS.n5276 VSS.n5275 5387.7
R21170 VSS.n5305 VSS.n2186 4902.86
R21171 VSS.n5333 VSS.n2177 4902.86
R21172 VSS.n2193 VSS.n2105 4902.86
R21173 VSS.n5289 VSS.n2091 4526.71
R21174 VSS.n5121 VSS.n4292 4493.06
R21175 VSS.n5253 VSS.n2237 3620.98
R21176 VSS.n3526 VSS.n3385 3491.91
R21177 VSS.n5280 VSS.n2201 3437.85
R21178 VSS.n3527 VSS.n2201 3435.27
R21179 VSS.n3316 VSS.n2966 3354.59
R21180 VSS.n3316 VSS.n2968 3354.59
R21181 VSS.n5290 VSS.n5289 3311.99
R21182 VSS.n3406 VSS.n3405 3307.91
R21183 VSS.n3525 VSS.n2200 3086.59
R21184 VSS.n5122 VSS.n5121 3080.18
R21185 VSS.n5332 VSS.n2178 2875.76
R21186 VSS.n3871 VSS.n2781 2717.55
R21187 VSS.n3871 VSS.n2782 2717.55
R21188 VSS.n5319 VSS.n5318 2717.55
R21189 VSS.n5318 VSS.n2185 2717.55
R21190 VSS.n5699 VSS.n9 2402.48
R21191 VSS.n5699 VSS.n10 2401.2
R21192 VSS.n5437 VSS.n9 2400.01
R21193 VSS.n5437 VSS.n10 2398.73
R21194 VSS.n5124 VSS.n5123 2352.1
R21195 VSS.n1744 VSS.n13 2286.22
R21196 VSS.n1742 VSS.n1729 2282.35
R21197 VSS.n1743 VSS.n1742 2282.35
R21198 VSS.n1729 VSS.n1293 2278.48
R21199 VSS.n1744 VSS.n1743 2277.19
R21200 VSS.n3409 VSS.n2091 2219.8
R21201 VSS.n5696 VSS.n13 2185.59
R21202 VSS.n2079 VSS.n1293 2179.14
R21203 VSS.n5128 VSS.n5127 2166.67
R21204 VSS.n5279 VSS.n2187 2099.5
R21205 VSS.n5331 VSS.n11 1924.39
R21206 VSS.n3526 VSS.n3524 1819.86
R21207 VSS.n909 VSS.n220 1814.99
R21208 VSS.n910 VSS.n909 1813.28
R21209 VSS.n5125 VSS.n5124 1481.53
R21210 VSS.n5315 VSS.n5314 1449.32
R21211 VSS.n5393 VSS.n2111 1375
R21212 VSS.n5314 VSS.n5306 1235.04
R21213 VSS.n5314 VSS.n5307 1235.04
R21214 VSS.n2892 VSS.n2891 1219.32
R21215 VSS.n3404 VSS.t26 1116.18
R21216 VSS.n5403 VSS.n2104 1089.54
R21217 VSS.n2891 VSS.t31 1038.26
R21218 VSS.n2080 VSS.n2079 967.646
R21219 VSS.n5697 VSS.n5696 967.646
R21220 VSS.t46 VSS.t26 953.457
R21221 VSS.t0 VSS.n2111 882.342
R21222 VSS.t12 VSS.n2111 882.342
R21223 VSS.n3406 VSS.n3398 835.686
R21224 VSS.n5318 VSS.n2186 815.005
R21225 VSS.n5394 VSS.n5393 800.532
R21226 VSS.t7 VSS.n5293 798.532
R21227 VSS.n5303 VSS.t11 798.532
R21228 VSS.n4044 VSS.t6 797.183
R21229 VSS.t31 VSS.n2291 744.888
R21230 VSS.n5392 VSS.n2112 709.234
R21231 VSS.n5334 VSS.n2176 709.234
R21232 VSS.n5293 VSS.n5292 693.769
R21233 VSS.n5304 VSS.n5303 693.769
R21234 VSS.n4044 VSS.n2202 693.769
R21235 VSS.n5394 VSS.n2105 676.944
R21236 VSS.n2430 VSS.n2427 675.573
R21237 VSS.n2430 VSS.n2239 675.573
R21238 VSS.n5249 VSS.n2240 675.573
R21239 VSS.n5403 VSS.n5402 651.337
R21240 VSS.n4051 VSS.t4 640.203
R21241 VSS.n5318 VSS.n5315 626.841
R21242 VSS.n5315 VSS.n2176 614.595
R21243 VSS.n3384 VSS.n2892 614.245
R21244 VSS.n5436 VSS.n2080 608.972
R21245 VSS.n5698 VSS.n5697 608.972
R21246 VSS.n5332 VSS.n5331 588.939
R21247 VSS.n5333 VSS.n5332 578.966
R21248 VSS.n4292 VSS.n4291 562.811
R21249 VSS.n5306 VSS.n5305 549.35
R21250 VSS.n5307 VSS.n2177 549.35
R21251 VSS.n2193 VSS.n2104 547.1
R21252 VSS.n5120 VSS.n2285 517.379
R21253 VSS.n5130 VSS.n2285 517.379
R21254 VSS.n5130 VSS.n2286 517.379
R21255 VSS.n5120 VSS.n2286 517.379
R21256 VSS.n3401 VSS.t40 515.692
R21257 VSS.n2781 VSS.n2093 488.243
R21258 VSS.n2782 VSS.n2097 488.243
R21259 VSS.n5319 VSS.n2182 488.243
R21260 VSS.n2185 VSS.n2179 488.243
R21261 VSS.n4248 VSS.n2353 472.197
R21262 VSS.n3401 VSS.t46 437.764
R21263 VSS.n2186 VSS.n2112 426.43
R21264 VSS.n5126 VSS.n5125 407.959
R21265 VSS.n4247 VSS.n2354 396.685
R21266 VSS.n5434 VSS.n2082 393.92
R21267 VSS.n2090 VSS.n2089 388.551
R21268 VSS.t37 VSS.n3395 363.911
R21269 VSS.n3395 VSS.t38 363.911
R21270 VSS.n5250 VSS.n5249 360.44
R21271 VSS.n5410 VSS.n5409 355.668
R21272 VSS.n4075 VSS.n2459 344.332
R21273 VSS.n4065 VSS.n4063 344.332
R21274 VSS.t42 VSS.n2292 343.325
R21275 VSS.n4076 VSS.t16 343.325
R21276 VSS.n4076 VSS.t14 343.325
R21277 VSS.t44 VSS.n4064 343.325
R21278 VSS.n5393 VSS.n5392 341.812
R21279 VSS.n2361 VSS.t47 334.264
R21280 VSS.t20 VSS.n2361 330.236
R21281 VSS.n5294 VSS.t7 325.932
R21282 VSS.n5299 VSS.t11 325.932
R21283 VSS.n5412 VSS.n2100 325.471
R21284 VSS.n5250 VSS.n2239 315.134
R21285 VSS.n5409 VSS.n2102 302.654
R21286 VSS.n4081 VSS.n2289 300.031
R21287 VSS.n2459 VSS.n2288 300.031
R21288 VSS.n2427 VSS.n2288 300.031
R21289 VSS.n2287 VSS.n2240 300.031
R21290 VSS.n4063 VSS.n2287 300.031
R21291 VSS.n5427 VSS.n2090 299.969
R21292 VSS.n5252 VSS.n5251 290.733
R21293 VSS.n4087 VSS.n2354 278.889
R21294 VSS.n3409 VSS.n2081 271
R21295 VSS.n3407 VSS.n3406 255.427
R21296 VSS.t24 VSS.t33 245.663
R21297 VSS.t47 VSS.t49 245.663
R21298 VSS.n5294 VSS.t0 242.12
R21299 VSS.n5299 VSS.t12 242.12
R21300 VSS.n5129 VSS.n5128 239.081
R21301 VSS.n4050 VSS.t6 236.487
R21302 VSS.n3029 VSS.n2966 233.749
R21303 VSS.n3258 VSS.n2968 233.749
R21304 VSS.t2 VSS.n2092 229.507
R21305 VSS.n2791 VSS.t2 229.507
R21306 VSS.n4082 VSS.n2444 227.541
R21307 VSS.n2200 VSS.n2195 224.798
R21308 VSS.n5254 VSS.n5253 219.064
R21309 VSS.t8 VSS.n2780 212.731
R21310 VSS.t40 VSS.n2291 208.569
R21311 VSS.n2451 VSS.t22 208.411
R21312 VSS.n4248 VSS.n4247 203.377
R21313 VSS.n5426 VSS.n5422 199.98
R21314 VSS.n2780 VSS.n2099 199.98
R21315 VSS.n4089 VSS.n4088 197.337
R21316 VSS.n4051 VSS.n2178 185.811
R21317 VSS.n5121 VSS.n5120 184.061
R21318 VSS.n5427 VSS.n5426 181.861
R21319 VSS.t4 VSS.n4050 175.677
R21320 VSS.n3384 VSS.n3383 170.571
R21321 VSS.t28 VSS.n3415 162.298
R21322 VSS.n5421 VSS.n2092 154.346
R21323 VSS.t35 VSS.n2290 154.043
R21324 VSS.n5437 VSS.n5436 152.252
R21325 VSS.n5699 VSS.n5698 152.252
R21326 VSS.n3509 VSS.t41 150.202
R21327 VSS.t18 VSS.n2370 149.01
R21328 VSS.n5292 VSS.n2193 146.669
R21329 VSS.n5305 VSS.n5304 146.669
R21330 VSS.n2202 VSS.n2177 146.669
R21331 VSS.n2371 VSS.t35 145.988
R21332 VSS.n3415 VSS.n2081 137.097
R21333 VSS.n3871 VSS.n2791 134.886
R21334 VSS.n5402 VSS.n2105 131.381
R21335 VSS.n5420 VSS.n2083 129.345
R21336 VSS.n5329 VSS.n5326 129.345
R21337 VSS.n5414 VSS.n2098 129.345
R21338 VSS.n5395 VSS.n2110 129.345
R21339 VSS.n5433 VSS.n2083 128.957
R21340 VSS.n5330 VSS.n5329 128.957
R21341 VSS.n3416 VSS.t28 122.984
R21342 VSS.n3416 VSS.t37 122.984
R21343 VSS.t41 VSS.n3507 122.984
R21344 VSS.n5334 VSS.n5333 118.02
R21345 VSS.n3509 VSS.n3508 114.919
R21346 VSS.n3516 VSS.n3515 114.919
R21347 VSS.n3517 VSS.n3516 114.919
R21348 VSS.n3517 VSS.n3386 114.919
R21349 VSS.n3523 VSS.n3386 114.919
R21350 VSS.n5287 VSS.n2195 114.919
R21351 VSS.n5288 VSS.n2194 112.903
R21352 VSS.n3524 VSS.n3523 111.895
R21353 VSS.t38 VSS.n3393 108.871
R21354 VSS.n5255 VSS.n5254 102.416
R21355 VSS.n3870 VSS.n2794 102.356
R21356 VSS.n5317 VSS.n2183 102.356
R21357 VSS.n5413 VSS.n5412 102.004
R21358 VSS.n5680 VSS.n15 99.728
R21359 VSS.n1294 VSS.n1171 99.7229
R21360 VSS.n2371 VSS.t18 99.6752
R21361 VSS.n3508 VSS.n3390 98.7908
R21362 VSS.n5413 VSS.n2099 97.977
R21363 VSS.n2370 VSS.t20 96.6548
R21364 VSS.t49 VSS.n2353 95.648
R21365 VSS.n2089 VSS.n2082 93.2795
R21366 VSS.t22 VSS.n2290 91.6207
R21367 VSS.n4082 VSS.n4081 90.6139
R21368 VSS.n910 VSS.n219 86.0408
R21369 VSS.n3872 VSS.t9 83.8845
R21370 VSS.n4089 VSS.n2289 82.5594
R21371 VSS.n4064 VSS.n2237 81.5525
R21372 VSS.n220 VSS.n219 80.8661
R21373 VSS.n3872 VSS.t8 79.858
R21374 VSS.t9 VSS.n3871 73.8184
R21375 VSS.n3317 VSS.n2964 73.4718
R21376 VSS.n3317 VSS.n2965 73.4718
R21377 VSS.n3073 VSS.n2967 73.2997
R21378 VSS.n2974 VSS.n2967 73.2997
R21379 VSS.n5401 VSS.n2106 72.4894
R21380 VSS.n2078 VSS.n1294 69.3341
R21381 VSS.n5695 VSS.n15 69.3341
R21382 VSS.n3398 VSS.n2081 64.5166
R21383 VSS.n2452 VSS.t24 61.4162
R21384 VSS.n5320 VSS.n2183 61.1338
R21385 VSS.n2184 VSS.n2183 61.1338
R21386 VSS.n2794 VSS.n2792 61.1338
R21387 VSS.n2794 VSS.n2793 61.1338
R21388 VSS.n2790 VSS.n2783 59.6561
R21389 VSS.n4066 VSS.n4062 59.6561
R21390 VSS.n2453 VSS.n2450 59.6561
R21391 VSS.n908 VSS.n219 58.4662
R21392 VSS.n2106 VSS.n2098 56.4672
R21393 VSS.n5395 VSS.n2106 56.4672
R21394 VSS.n4066 VSS.n4059 56.0005
R21395 VSS.n4074 VSS.n2460 56.0005
R21396 VSS.n2453 VSS.n2448 56.0005
R21397 VSS.n3383 VSS.n3381 55.8444
R21398 VSS.n5404 VSS.n2102 53.0152
R21399 VSS.n5422 VSS.n5421 45.6334
R21400 VSS.n5404 VSS.n5403 41.6069
R21401 VSS.n5420 VSS.n2093 40.8338
R21402 VSS.n5326 VSS.n2179 40.8338
R21403 VSS.n2182 VSS.n2110 40.8338
R21404 VSS.n5414 VSS.n2097 40.8338
R21405 VSS.n3315 VSS.n2969 40.2769
R21406 VSS.n3315 VSS.n2970 40.2769
R21407 VSS.n5254 VSS.n2224 39.6013
R21408 VSS.n4291 VSS.n2292 37.2527
R21409 VSS.t33 VSS.n2451 37.2527
R21410 VSS.n4077 VSS.n2457 33.0561
R21411 VSS.n5410 VSS.n2100 30.1987
R21412 VSS.n5444 VSS.n5443 29.3117
R21413 VSS.n5444 VSS.n1285 29.3117
R21414 VSS.n5450 VSS.n1285 29.3117
R21415 VSS.n5451 VSS.n5450 29.3117
R21416 VSS.n5452 VSS.n5451 29.3117
R21417 VSS.n5452 VSS.n1281 29.3117
R21418 VSS.n5458 VSS.n1281 29.3117
R21419 VSS.n5459 VSS.n5458 29.3117
R21420 VSS.n5460 VSS.n5459 29.3117
R21421 VSS.n5460 VSS.n1277 29.3117
R21422 VSS.n5466 VSS.n1277 29.3117
R21423 VSS.n5467 VSS.n5466 29.3117
R21424 VSS.n5468 VSS.n5467 29.3117
R21425 VSS.n5468 VSS.n1273 29.3117
R21426 VSS.n5474 VSS.n1273 29.3117
R21427 VSS.n5475 VSS.n5474 29.3117
R21428 VSS.n5476 VSS.n5475 29.3117
R21429 VSS.n5476 VSS.n1269 29.3117
R21430 VSS.n5482 VSS.n1269 29.3117
R21431 VSS.n5483 VSS.n5482 29.3117
R21432 VSS.n5484 VSS.n5483 29.3117
R21433 VSS.n5484 VSS.n1265 29.3117
R21434 VSS.n5490 VSS.n1265 29.3117
R21435 VSS.n5491 VSS.n5490 29.3117
R21436 VSS.n5492 VSS.n5491 29.3117
R21437 VSS.n5492 VSS.n1261 29.3117
R21438 VSS.n5498 VSS.n1261 29.3117
R21439 VSS.n5499 VSS.n5498 29.3117
R21440 VSS.n5500 VSS.n5499 29.3117
R21441 VSS.n5500 VSS.n1257 29.3117
R21442 VSS.n5506 VSS.n1257 29.3117
R21443 VSS.n5507 VSS.n5506 29.3117
R21444 VSS.n5508 VSS.n5507 29.3117
R21445 VSS.n5508 VSS.n1253 29.3117
R21446 VSS.n5514 VSS.n1253 29.3117
R21447 VSS.n5515 VSS.n5514 29.3117
R21448 VSS.n5516 VSS.n5515 29.3117
R21449 VSS.n5516 VSS.n1249 29.3117
R21450 VSS.n5522 VSS.n1249 29.3117
R21451 VSS.n5523 VSS.n5522 29.3117
R21452 VSS.n5524 VSS.n5523 29.3117
R21453 VSS.n5524 VSS.n1245 29.3117
R21454 VSS.n5530 VSS.n1245 29.3117
R21455 VSS.n5531 VSS.n5530 29.3117
R21456 VSS.n5532 VSS.n5531 29.3117
R21457 VSS.n5532 VSS.n1241 29.3117
R21458 VSS.n5538 VSS.n1241 29.3117
R21459 VSS.n5539 VSS.n5538 29.3117
R21460 VSS.n5540 VSS.n5539 29.3117
R21461 VSS.n5540 VSS.n1237 29.3117
R21462 VSS.n5546 VSS.n1237 29.3117
R21463 VSS.n5547 VSS.n5546 29.3117
R21464 VSS.n5548 VSS.n5547 29.3117
R21465 VSS.n5548 VSS.n1233 29.3117
R21466 VSS.n5555 VSS.n1233 29.3117
R21467 VSS.n5556 VSS.n5555 29.3117
R21468 VSS.n5558 VSS.n1229 29.3117
R21469 VSS.n5564 VSS.n1229 29.3117
R21470 VSS.n5565 VSS.n5564 29.3117
R21471 VSS.n5566 VSS.n5565 29.3117
R21472 VSS.n5566 VSS.n1225 29.3117
R21473 VSS.n5572 VSS.n1225 29.3117
R21474 VSS.n5573 VSS.n5572 29.3117
R21475 VSS.n5574 VSS.n5573 29.3117
R21476 VSS.n5574 VSS.n1221 29.3117
R21477 VSS.n5580 VSS.n1221 29.3117
R21478 VSS.n5581 VSS.n5580 29.3117
R21479 VSS.n5582 VSS.n5581 29.3117
R21480 VSS.n5582 VSS.n1217 29.3117
R21481 VSS.n5588 VSS.n1217 29.3117
R21482 VSS.n5589 VSS.n5588 29.3117
R21483 VSS.n5590 VSS.n5589 29.3117
R21484 VSS.n5590 VSS.n1213 29.3117
R21485 VSS.n5596 VSS.n1213 29.3117
R21486 VSS.n5597 VSS.n5596 29.3117
R21487 VSS.n5598 VSS.n5597 29.3117
R21488 VSS.n5598 VSS.n1209 29.3117
R21489 VSS.n5604 VSS.n1209 29.3117
R21490 VSS.n5605 VSS.n5604 29.3117
R21491 VSS.n5606 VSS.n5605 29.3117
R21492 VSS.n5606 VSS.n1205 29.3117
R21493 VSS.n5612 VSS.n1205 29.3117
R21494 VSS.n5613 VSS.n5612 29.3117
R21495 VSS.n5614 VSS.n5613 29.3117
R21496 VSS.n5614 VSS.n1201 29.3117
R21497 VSS.n5620 VSS.n1201 29.3117
R21498 VSS.n5621 VSS.n5620 29.3117
R21499 VSS.n5622 VSS.n5621 29.3117
R21500 VSS.n5622 VSS.n1197 29.3117
R21501 VSS.n5628 VSS.n1197 29.3117
R21502 VSS.n5629 VSS.n5628 29.3117
R21503 VSS.n5630 VSS.n5629 29.3117
R21504 VSS.n5630 VSS.n1193 29.3117
R21505 VSS.n5636 VSS.n1193 29.3117
R21506 VSS.n5637 VSS.n5636 29.3117
R21507 VSS.n5638 VSS.n5637 29.3117
R21508 VSS.n5638 VSS.n1189 29.3117
R21509 VSS.n5644 VSS.n1189 29.3117
R21510 VSS.n5645 VSS.n5644 29.3117
R21511 VSS.n5646 VSS.n5645 29.3117
R21512 VSS.n5646 VSS.n1185 29.3117
R21513 VSS.n5652 VSS.n1185 29.3117
R21514 VSS.n5653 VSS.n5652 29.3117
R21515 VSS.n5654 VSS.n5653 29.3117
R21516 VSS.n5654 VSS.n1181 29.3117
R21517 VSS.n5660 VSS.n1181 29.3117
R21518 VSS.n5661 VSS.n5660 29.3117
R21519 VSS.n5662 VSS.n5661 29.3117
R21520 VSS.n5662 VSS.n1177 29.3117
R21521 VSS.n5668 VSS.n1177 29.3117
R21522 VSS.n5669 VSS.n5668 29.3117
R21523 VSS.n5670 VSS.n5669 29.3117
R21524 VSS.n5670 VSS.n1173 29.3117
R21525 VSS.n2457 VSS.n2445 26.6005
R21526 VSS.n4074 VSS.n2457 26.6005
R21527 VSS.n2458 VSS.n2444 26.1777
R21528 VSS.n5443 VSS.n5442 21.9839
R21529 VSS.n5435 VSS.n5434 21.4748
R21530 VSS.n4088 VSS.n4087 20.1368
R21531 VSS.n5676 VSS.n5675 19.8563
R21532 VSS.n3515 VSS.n3390 16.1295
R21533 VSS.n2086 VSS.n2085 15.9461
R21534 VSS.n5328 VSS.n5327 15.9461
R21535 VSS.n5396 VSS.n2109 15.9461
R21536 VSS.n2796 VSS.n2795 15.9461
R21537 VSS.n5700 VSS.n8 14.9905
R21538 VSS.n5558 VSS.n5557 14.8925
R21539 VSS.n5440 VSS.n5438 14.6859
R21540 VSS.n5557 VSS.n5556 14.4197
R21541 VSS.n4083 DVSS 14.1351
R21542 VSS.n3507 VSS.n3393 14.1134
R21543 VSS.n3731 VSS.n3729 12.4433
R21544 VSS.n5676 VSS.n1173 12.0559
R21545 VSS VSS.t30 11.0117
R21546 VSS.n5301 VSS 10.8266
R21547 VSS.n2191 VSS 10.8266
R21548 VSS.n4045 VSS 10.8266
R21549 VSS.n5701 VSS.n7 10.6235
R21550 VSS.n2312 VSS.n1291 10.6235
R21551 VSS.n5442 VSS.n1289 9.92831
R21552 VSS.n2311 VSS.n7 8.07493
R21553 VSS.n2312 VSS.n2311 8.03957
R21554 VSS.n3073 VSS.n2970 7.77509
R21555 VSS.n2974 VSS.n2969 7.77509
R21556 VSS.n1745 VSS.n14 7.61966
R21557 VSS.n1741 VSS.n1735 7.60677
R21558 VSS.n1741 VSS.n1728 7.60677
R21559 VSS.n2969 VSS.n2964 7.60296
R21560 VSS.n2970 VSS.n2965 7.60296
R21561 VSS.n1735 VSS.n1295 7.59387
R21562 VSS.n1745 VSS.n1728 7.58957
R21563 VSS.n5695 VSS.n14 7.28428
R21564 VSS.n2078 VSS.n1295 7.26279
R21565 VSS.n2456 VSS.n2455 6.95655
R21566 VSS.n4070 VSS 6.91517
R21567 VSS.n2362 VSS.t50 6.33948
R21568 VSS.n2364 VSS.t48 6.33948
R21569 VSS.n2889 VSS.n2888 6.3005
R21570 VSS.n2367 VSS.n2366 6.3005
R21571 VSS.n2294 VSS.n2293 6.3005
R21572 VSS.n4286 VSS.n4285 6.3005
R21573 VSS.n4289 VSS.n4288 6.3005
R21574 VSS.n3400 VSS.n3399 6.3005
R21575 VSS.n5701 VSS.n5700 6.17435
R21576 VSS.n5438 VSS.n1291 6.17435
R21577 VSS.n5689 VSS.n5688 5.42247
R21578 VSS VSS.t55 5.2005
R21579 VSS VSS.t52 5.2005
R21580 VSS VSS.t53 5.2005
R21581 VSS VSS.t54 5.2005
R21582 VSS VSS.t56 5.2005
R21583 VSS VSS.t51 5.2005
R21584 VSS.n5257 VSS.n2223 5.2005
R21585 VSS.n5274 VSS.n2223 5.2005
R21586 VSS.n5257 VSS.n2224 5.2005
R21587 VSS.n2224 VSS.n2210 5.2005
R21588 VSS.n2224 VSS.n2208 5.2005
R21589 VSS.n2224 VSS.n2211 5.2005
R21590 VSS.n2224 VSS.n2207 5.2005
R21591 VSS.n2224 VSS.n2212 5.2005
R21592 VSS.n2224 VSS.n2206 5.2005
R21593 VSS.n2224 VSS.n2213 5.2005
R21594 VSS.n2224 VSS.n2205 5.2005
R21595 VSS.n2224 VSS.n2214 5.2005
R21596 VSS.n5271 VSS.n2224 5.2005
R21597 VSS.n5274 VSS.n2224 5.2005
R21598 VSS.n5257 VSS.n2217 5.2005
R21599 VSS.n2217 VSS.n2210 5.2005
R21600 VSS.n2217 VSS.n2208 5.2005
R21601 VSS.n2217 VSS.n2211 5.2005
R21602 VSS.n2217 VSS.n2207 5.2005
R21603 VSS.n2217 VSS.n2212 5.2005
R21604 VSS.n2217 VSS.n2206 5.2005
R21605 VSS.n2217 VSS.n2213 5.2005
R21606 VSS.n2217 VSS.n2205 5.2005
R21607 VSS.n2217 VSS.n2214 5.2005
R21608 VSS.n5274 VSS.n2217 5.2005
R21609 VSS.n5257 VSS.n2225 5.2005
R21610 VSS.n2225 VSS.n2210 5.2005
R21611 VSS.n2225 VSS.n2208 5.2005
R21612 VSS.n2225 VSS.n2211 5.2005
R21613 VSS.n2225 VSS.n2207 5.2005
R21614 VSS.n2225 VSS.n2212 5.2005
R21615 VSS.n2225 VSS.n2206 5.2005
R21616 VSS.n2225 VSS.n2213 5.2005
R21617 VSS.n2225 VSS.n2205 5.2005
R21618 VSS.n2225 VSS.n2214 5.2005
R21619 VSS.n5274 VSS.n2225 5.2005
R21620 VSS.n5257 VSS.n2216 5.2005
R21621 VSS.n2216 VSS.n2210 5.2005
R21622 VSS.n2216 VSS.n2208 5.2005
R21623 VSS.n2216 VSS.n2211 5.2005
R21624 VSS.n2216 VSS.n2207 5.2005
R21625 VSS.n2216 VSS.n2212 5.2005
R21626 VSS.n2216 VSS.n2206 5.2005
R21627 VSS.n2216 VSS.n2213 5.2005
R21628 VSS.n2216 VSS.n2205 5.2005
R21629 VSS.n2216 VSS.n2214 5.2005
R21630 VSS.n5274 VSS.n2216 5.2005
R21631 VSS.n5257 VSS.n2226 5.2005
R21632 VSS.n2226 VSS.n2210 5.2005
R21633 VSS.n2226 VSS.n2208 5.2005
R21634 VSS.n2226 VSS.n2211 5.2005
R21635 VSS.n2226 VSS.n2207 5.2005
R21636 VSS.n2226 VSS.n2212 5.2005
R21637 VSS.n2226 VSS.n2206 5.2005
R21638 VSS.n2226 VSS.n2213 5.2005
R21639 VSS.n2226 VSS.n2205 5.2005
R21640 VSS.n2226 VSS.n2214 5.2005
R21641 VSS.n5274 VSS.n2226 5.2005
R21642 VSS.n5257 VSS.n2215 5.2005
R21643 VSS.n2215 VSS.n2210 5.2005
R21644 VSS.n2215 VSS.n2208 5.2005
R21645 VSS.n2215 VSS.n2211 5.2005
R21646 VSS.n2215 VSS.n2207 5.2005
R21647 VSS.n2215 VSS.n2212 5.2005
R21648 VSS.n2215 VSS.n2206 5.2005
R21649 VSS.n2215 VSS.n2213 5.2005
R21650 VSS.n2215 VSS.n2205 5.2005
R21651 VSS.n2215 VSS.n2214 5.2005
R21652 VSS.n5274 VSS.n2215 5.2005
R21653 VSS.n5275 VSS.n2210 5.2005
R21654 VSS.n5275 VSS.n2208 5.2005
R21655 VSS.n5275 VSS.n2211 5.2005
R21656 VSS.n5275 VSS.n2207 5.2005
R21657 VSS.n5275 VSS.n2212 5.2005
R21658 VSS.n5275 VSS.n2206 5.2005
R21659 VSS.n5275 VSS.n2213 5.2005
R21660 VSS.n5275 VSS.n2205 5.2005
R21661 VSS.n5275 VSS.n2214 5.2005
R21662 VSS.n5275 VSS.n5274 5.2005
R21663 VSS.n3729 VSS.n2817 5.08553
R21664 VSS.n5255 VSS.n2232 4.84618
R21665 VSS.n2230 VSS.n2217 4.84618
R21666 VSS.n5269 VSS.n2225 4.84618
R21667 VSS.n2229 VSS.n2216 4.84618
R21668 VSS.n5270 VSS.n2226 4.84618
R21669 VSS.n2228 VSS.n2215 4.84618
R21670 VSS.n5275 VSS.n2204 4.84618
R21671 VSS.n2232 VSS.n2223 4.84618
R21672 VSS.n2230 VSS.n2224 4.84618
R21673 VSS.n5269 VSS.n2217 4.84618
R21674 VSS.n2229 VSS.n2225 4.84618
R21675 VSS.n5270 VSS.n2216 4.84618
R21676 VSS.n2228 VSS.n2226 4.84618
R21677 VSS.n2215 VSS.n2204 4.84618
R21678 VSS.n3504 VSS.n3503 4.82802
R21679 VSS.n3486 VSS.n3485 4.66866
R21680 VSS.n3887 VSS.n3886 4.66866
R21681 VSS.n4071 VSS.n4070 4.58103
R21682 VSS.n5301 VSS 4.5005
R21683 VSS.n2191 VSS 4.5005
R21684 VSS.n4045 VSS 4.5005
R21685 VSS.n3638 VSS.n2879 4.5005
R21686 VSS.n2885 VSS.n2879 4.5005
R21687 VSS.n3640 VSS.n2879 4.5005
R21688 VSS.n3638 VSS.n2881 4.5005
R21689 VSS.n2885 VSS.n2881 4.5005
R21690 VSS.n3640 VSS.n2881 4.5005
R21691 VSS.n3640 VSS.n2878 4.5005
R21692 VSS.n2885 VSS.n2878 4.5005
R21693 VSS.n3638 VSS.n2878 4.5005
R21694 VSS.n3640 VSS.n2882 4.5005
R21695 VSS.n2885 VSS.n2882 4.5005
R21696 VSS.n3638 VSS.n2882 4.5005
R21697 VSS.n3638 VSS.n2877 4.5005
R21698 VSS.n2885 VSS.n2877 4.5005
R21699 VSS.n3640 VSS.n2877 4.5005
R21700 VSS.n3640 VSS.n2883 4.5005
R21701 VSS.n2885 VSS.n2883 4.5005
R21702 VSS.n3638 VSS.n2883 4.5005
R21703 VSS.n3638 VSS.n2876 4.5005
R21704 VSS.n2885 VSS.n2876 4.5005
R21705 VSS.n3640 VSS.n2876 4.5005
R21706 VSS.n3640 VSS.n3639 4.5005
R21707 VSS.n3639 VSS.n2885 4.5005
R21708 VSS.n3639 VSS.n3638 4.5005
R21709 VSS.n2074 VSS.n2073 4.5005
R21710 VSS.n2073 VSS.n2071 4.5005
R21711 VSS.n2073 VSS.n2067 4.5005
R21712 VSS.n2072 VSS.n1594 4.5005
R21713 VSS.n2073 VSS.n2072 4.5005
R21714 VSS.n1597 VSS.n1595 4.5005
R21715 VSS.n2062 VSS.n1595 4.5005
R21716 VSS.n2065 VSS.n1595 4.5005
R21717 VSS.n2066 VSS.n1597 4.5005
R21718 VSS.n2066 VSS.n2065 4.5005
R21719 VSS.n2065 VSS.n1602 4.5005
R21720 VSS.n2065 VSS.n1605 4.5005
R21721 VSS.n2065 VSS.n1601 4.5005
R21722 VSS.n2065 VSS.n1607 4.5005
R21723 VSS.n2065 VSS.n1600 4.5005
R21724 VSS.n2065 VSS.n1609 4.5005
R21725 VSS.n2065 VSS.n1599 4.5005
R21726 VSS.n2064 VSS.n2062 4.5005
R21727 VSS.n2065 VSS.n2064 4.5005
R21728 VSS.n1854 VSS.n1797 4.5005
R21729 VSS.n1857 VSS.n1797 4.5005
R21730 VSS.n1797 VSS.n1792 4.5005
R21731 VSS.n1854 VSS.n1820 4.5005
R21732 VSS.n1820 VSS.n1792 4.5005
R21733 VSS.n1807 VSS.n1792 4.5005
R21734 VSS.n1806 VSS.n1792 4.5005
R21735 VSS.n1804 VSS.n1792 4.5005
R21736 VSS.n1803 VSS.n1792 4.5005
R21737 VSS.n1801 VSS.n1792 4.5005
R21738 VSS.n1800 VSS.n1792 4.5005
R21739 VSS.n1799 VSS.n1792 4.5005
R21740 VSS.n1857 VSS.n1856 4.5005
R21741 VSS.n1856 VSS.n1792 4.5005
R21742 VSS.n1819 VSS.n1818 4.5005
R21743 VSS.n1818 VSS.n1810 4.5005
R21744 VSS.n1810 VSS.n16 4.5005
R21745 VSS.n1813 VSS.n16 4.5005
R21746 VSS.n1815 VSS.n16 4.5005
R21747 VSS.n1818 VSS.n1817 4.5005
R21748 VSS.n1817 VSS.n16 4.5005
R21749 VSS.n1144 VSS.n34 4.5005
R21750 VSS.n1142 VSS.n1141 4.5005
R21751 VSS.n1140 VSS.n1139 4.5005
R21752 VSS.n1078 VSS.n77 4.5005
R21753 VSS.n5688 VSS.n32 4.5005
R21754 VSS.n1145 VSS.n33 4.5005
R21755 VSS.n5690 VSS.n27 4.5005
R21756 VSS.n27 VSS.n19 4.5005
R21757 VSS.n27 VSS.n20 4.5005
R21758 VSS.n27 VSS.n22 4.5005
R21759 VSS.n24 VSS.n20 4.5005
R21760 VSS.n24 VSS.n22 4.5005
R21761 VSS.n5690 VSS.n28 4.5005
R21762 VSS.n28 VSS.n19 4.5005
R21763 VSS.n28 VSS.n20 4.5005
R21764 VSS.n28 VSS.n22 4.5005
R21765 VSS.n5690 VSS.n26 4.5005
R21766 VSS.n26 VSS.n19 4.5005
R21767 VSS.n26 VSS.n20 4.5005
R21768 VSS.n26 VSS.n22 4.5005
R21769 VSS.n30 VSS.n20 4.5005
R21770 VSS.n30 VSS.n22 4.5005
R21771 VSS.n25 VSS.n20 4.5005
R21772 VSS.n25 VSS.n22 4.5005
R21773 VSS.n5690 VSS.n29 4.5005
R21774 VSS.n29 VSS.n19 4.5005
R21775 VSS.n29 VSS.n20 4.5005
R21776 VSS.n29 VSS.n22 4.5005
R21777 VSS.n5691 VSS.n20 4.5005
R21778 VSS.n5691 VSS.n22 4.5005
R21779 VSS.n20 VSS.n18 4.5005
R21780 VSS.n22 VSS.n18 4.5005
R21781 VSS.n19 VSS.n18 4.5005
R21782 VSS.n5690 VSS.n18 4.5005
R21783 VSS.n5691 VSS.n19 4.5005
R21784 VSS.n5691 VSS.n5690 4.5005
R21785 VSS.n25 VSS.n19 4.5005
R21786 VSS.n5690 VSS.n25 4.5005
R21787 VSS.n30 VSS.n19 4.5005
R21788 VSS.n5690 VSS.n30 4.5005
R21789 VSS.n24 VSS.n19 4.5005
R21790 VSS.n5690 VSS.n24 4.5005
R21791 VSS.n5689 VSS.n22 4.5005
R21792 VSS.n5689 VSS.n20 4.5005
R21793 VSS.n5689 VSS.n19 4.5005
R21794 VSS.n5690 VSS.n5689 4.5005
R21795 VSS.n3324 VSS.n2957 4.5005
R21796 VSS.n2960 VSS.n2957 4.5005
R21797 VSS.n3323 VSS.n2960 4.5005
R21798 VSS.n3324 VSS.n3323 4.5005
R21799 VSS.n3107 VSS.n2958 4.5005
R21800 VSS.n2973 VSS.n2958 4.5005
R21801 VSS.n3334 VSS.n2948 4.5005
R21802 VSS.n3334 VSS.n3333 4.5005
R21803 VSS.n3333 VSS.n3332 4.5005
R21804 VSS.n3332 VSS.n2948 4.5005
R21805 VSS.n3068 VSS.n2949 4.5005
R21806 VSS.n3069 VSS.n3068 4.5005
R21807 VSS.n3352 VSS.n2920 4.5005
R21808 VSS.n3352 VSS.n2922 4.5005
R21809 VSS.n3352 VSS.n2919 4.5005
R21810 VSS.n3352 VSS.n3351 4.5005
R21811 VSS.n3351 VSS.n3350 4.5005
R21812 VSS.n3350 VSS.n2919 4.5005
R21813 VSS.n3350 VSS.n2922 4.5005
R21814 VSS.n3350 VSS.n2920 4.5005
R21815 VSS.n2977 VSS.n2921 4.5005
R21816 VSS.n3007 VSS.n2921 4.5005
R21817 VSS.n3007 VSS.n3006 4.5005
R21818 VSS.n3007 VSS.n2978 4.5005
R21819 VSS.n3008 VSS.n2977 4.5005
R21820 VSS.n3008 VSS.n3007 4.5005
R21821 VSS.n3137 VSS.n3077 4.5005
R21822 VSS.n3137 VSS.n3081 4.5005
R21823 VSS.n3137 VSS.n3082 4.5005
R21824 VSS.n3137 VSS.n3089 4.5005
R21825 VSS.n3094 VSS.n3089 4.5005
R21826 VSS.n3094 VSS.n3082 4.5005
R21827 VSS.n3094 VSS.n3081 4.5005
R21828 VSS.n3094 VSS.n3077 4.5005
R21829 VSS.n3079 VSS.n3076 4.5005
R21830 VSS.n3307 VSS.n3079 4.5005
R21831 VSS.n3307 VSS.n3306 4.5005
R21832 VSS.n3307 VSS.n3078 4.5005
R21833 VSS.n3308 VSS.n3076 4.5005
R21834 VSS.n3308 VSS.n3307 4.5005
R21835 VSS.n3255 VSS.n3246 4.5005
R21836 VSS.n3255 VSS.n3153 4.5005
R21837 VSS.n3261 VSS.n3246 4.5005
R21838 VSS.n3261 VSS.n3153 4.5005
R21839 VSS.n3268 VSS.n3153 4.5005
R21840 VSS.n3268 VSS.n3246 4.5005
R21841 VSS.n3277 VSS.n3154 4.5005
R21842 VSS.n3279 VSS.n3154 4.5005
R21843 VSS.n3279 VSS.n3278 4.5005
R21844 VSS.n3278 VSS.n3277 4.5005
R21845 VSS.n3266 VSS.n3153 4.5005
R21846 VSS.n3266 VSS.n3246 4.5005
R21847 VSS.n3261 VSS.n3259 4.5005
R21848 VSS.n3261 VSS.n3260 4.5005
R21849 VSS.n3273 VSS.n3247 4.5005
R21850 VSS.n3274 VSS.n3273 4.5005
R21851 VSS.n2915 VSS.n2913 4.5005
R21852 VSS.n2935 VSS.n2915 4.5005
R21853 VSS.n3140 VSS.n3096 4.5005
R21854 VSS.n3141 VSS.n3140 4.5005
R21855 VSS.n3275 VSS.n3247 4.5005
R21856 VSS.n3275 VSS.n3274 4.5005
R21857 VSS.n3320 VSS.n2963 4.5005
R21858 VSS.n3320 VSS.n3319 4.5005
R21859 VSS.n3335 VSS.n2947 4.5005
R21860 VSS.n3335 VSS.n2944 4.5005
R21861 VSS.n2413 VSS.n2408 4.5005
R21862 VSS.n4186 VSS.n2413 4.5005
R21863 VSS.n4186 VSS.n4174 4.5005
R21864 VSS.n4186 VSS.n2412 4.5005
R21865 VSS.n4186 VSS.n4177 4.5005
R21866 VSS.n4186 VSS.n2411 4.5005
R21867 VSS.n4186 VSS.n4180 4.5005
R21868 VSS.n4186 VSS.n2410 4.5005
R21869 VSS.n4186 VSS.n4183 4.5005
R21870 VSS.n4186 VSS.n2409 4.5005
R21871 VSS.n4185 VSS.n2408 4.5005
R21872 VSS.n4186 VSS.n4185 4.5005
R21873 VSS.n3359 VSS.n3358 4.5005
R21874 VSS.n3358 VSS.n3357 4.5005
R21875 VSS.n2994 VSS.n2993 4.5005
R21876 VSS.n2994 VSS.n2985 4.5005
R21877 VSS.n2995 VSS.n2994 4.5005
R21878 VSS.n2995 VSS.n2909 4.5005
R21879 VSS.n2985 VSS.n2909 4.5005
R21880 VSS.n2993 VSS.n2909 4.5005
R21881 VSS.n3055 VSS.n3030 4.5005
R21882 VSS.n3010 VSS.n2903 4.5005
R21883 VSS.n3024 VSS.n2899 4.5005
R21884 VSS.n3024 VSS.n2903 4.5005
R21885 VSS.n3012 VSS.n2899 4.5005
R21886 VSS.n3012 VSS.n2903 4.5005
R21887 VSS.n3010 VSS.n2899 4.5005
R21888 VSS.n3055 VSS.n2899 4.5005
R21889 VSS.n3055 VSS.n2903 4.5005
R21890 VSS.n3056 VSS.n3055 4.5005
R21891 VSS.n2832 VSS.n2827 4.5005
R21892 VSS.n3715 VSS.n2832 4.5005
R21893 VSS.n3713 VSS.n2832 4.5005
R21894 VSS.n2834 VSS.n2827 4.5005
R21895 VSS.n3715 VSS.n2834 4.5005
R21896 VSS.n3713 VSS.n2834 4.5005
R21897 VSS.n3713 VSS.n2831 4.5005
R21898 VSS.n3715 VSS.n2831 4.5005
R21899 VSS.n2831 VSS.n2827 4.5005
R21900 VSS.n2835 VSS.n2827 4.5005
R21901 VSS.n3715 VSS.n2835 4.5005
R21902 VSS.n3713 VSS.n2835 4.5005
R21903 VSS.n2830 VSS.n2827 4.5005
R21904 VSS.n3715 VSS.n2830 4.5005
R21905 VSS.n3713 VSS.n2830 4.5005
R21906 VSS.n3713 VSS.n2836 4.5005
R21907 VSS.n3715 VSS.n2836 4.5005
R21908 VSS.n2836 VSS.n2827 4.5005
R21909 VSS.n3713 VSS.n2829 4.5005
R21910 VSS.n3715 VSS.n2829 4.5005
R21911 VSS.n2829 VSS.n2827 4.5005
R21912 VSS.n2837 VSS.n2827 4.5005
R21913 VSS.n3715 VSS.n2837 4.5005
R21914 VSS.n3713 VSS.n2837 4.5005
R21915 VSS.n3713 VSS.n2828 4.5005
R21916 VSS.n3715 VSS.n2828 4.5005
R21917 VSS.n2828 VSS.n2827 4.5005
R21918 VSS.n3714 VSS.n3713 4.5005
R21919 VSS.n3715 VSS.n3714 4.5005
R21920 VSS.n3714 VSS.n2827 4.5005
R21921 VSS.n3053 VSS.n3052 4.5005
R21922 VSS.n3049 VSS.n2887 4.5005
R21923 VSS.n3054 VSS.n3053 4.5005
R21924 VSS.n3054 VSS.n3048 4.5005
R21925 VSS.n3054 VSS.n2887 4.5005
R21926 VSS.n4057 VSS.n2462 4.5005
R21927 VSS.n4057 VSS.n4056 4.5005
R21928 VSS.n4056 VSS.n2470 4.5005
R21929 VSS.n4056 VSS.n2467 4.5005
R21930 VSS.n4056 VSS.n2472 4.5005
R21931 VSS.n4056 VSS.n2466 4.5005
R21932 VSS.n4056 VSS.n2474 4.5005
R21933 VSS.n4056 VSS.n2465 4.5005
R21934 VSS.n4056 VSS.n2476 4.5005
R21935 VSS.n4056 VSS.n2464 4.5005
R21936 VSS.n4055 VSS.n2462 4.5005
R21937 VSS.n4056 VSS.n4055 4.5005
R21938 VSS.n3886 VSS.n3885 4.5005
R21939 VSS.n2773 VSS.n2772 4.5005
R21940 VSS.n3877 VSS.n3876 4.5005
R21941 VSS.n2779 VSS.n2777 4.5005
R21942 VSS.n3480 VSS.n3478 4.5005
R21943 VSS.n3485 VSS.n3484 4.5005
R21944 VSS.n4054 VSS.n0 4.5005
R21945 VSS.n4054 VSS.n4026 4.5005
R21946 VSS.n4043 VSS.n0 4.5005
R21947 VSS.n4037 VSS.n1 4.5005
R21948 VSS.n4039 VSS.n1 4.5005
R21949 VSS.n4041 VSS.n1 4.5005
R21950 VSS.n4043 VSS.n1 4.5005
R21951 VSS.n4054 VSS.n1 4.5005
R21952 VSS.n4035 VSS.n4026 4.5005
R21953 VSS.n4033 VSS.n4026 4.5005
R21954 VSS.n4031 VSS.n4026 4.5005
R21955 VSS.n4029 VSS.n4026 4.5005
R21956 VSS.n4027 VSS.n1 4.5005
R21957 VSS.n4027 VSS.n4026 4.5005
R21958 VSS.n4058 VSS.n4057 4.24863
R21959 VSS.n1289 VSS.n1288 4.05657
R21960 VSS.n5445 VSS.n1288 4.05657
R21961 VSS.n5445 VSS.n1286 4.05657
R21962 VSS.n5449 VSS.n1286 4.05657
R21963 VSS.n5449 VSS.n1284 4.05657
R21964 VSS.n5453 VSS.n1284 4.05657
R21965 VSS.n5453 VSS.n1282 4.05657
R21966 VSS.n5457 VSS.n1282 4.05657
R21967 VSS.n5457 VSS.n1280 4.05657
R21968 VSS.n5461 VSS.n1280 4.05657
R21969 VSS.n5461 VSS.n1278 4.05657
R21970 VSS.n5465 VSS.n1278 4.05657
R21971 VSS.n5465 VSS.n1276 4.05657
R21972 VSS.n5469 VSS.n1276 4.05657
R21973 VSS.n5469 VSS.n1274 4.05657
R21974 VSS.n5473 VSS.n1274 4.05657
R21975 VSS.n5473 VSS.n1272 4.05657
R21976 VSS.n5477 VSS.n1272 4.05657
R21977 VSS.n5477 VSS.n1270 4.05657
R21978 VSS.n5481 VSS.n1270 4.05657
R21979 VSS.n5481 VSS.n1268 4.05657
R21980 VSS.n5485 VSS.n1268 4.05657
R21981 VSS.n5485 VSS.n1266 4.05657
R21982 VSS.n5489 VSS.n1266 4.05657
R21983 VSS.n5489 VSS.n1264 4.05657
R21984 VSS.n5493 VSS.n1264 4.05657
R21985 VSS.n5493 VSS.n1262 4.05657
R21986 VSS.n5497 VSS.n1262 4.05657
R21987 VSS.n5497 VSS.n1260 4.05657
R21988 VSS.n5501 VSS.n1260 4.05657
R21989 VSS.n5501 VSS.n1258 4.05657
R21990 VSS.n5505 VSS.n1258 4.05657
R21991 VSS.n5505 VSS.n1256 4.05657
R21992 VSS.n5509 VSS.n1256 4.05657
R21993 VSS.n5509 VSS.n1254 4.05657
R21994 VSS.n5513 VSS.n1254 4.05657
R21995 VSS.n5513 VSS.n1252 4.05657
R21996 VSS.n5517 VSS.n1252 4.05657
R21997 VSS.n5517 VSS.n1250 4.05657
R21998 VSS.n5521 VSS.n1250 4.05657
R21999 VSS.n5521 VSS.n1248 4.05657
R22000 VSS.n5525 VSS.n1248 4.05657
R22001 VSS.n5525 VSS.n1246 4.05657
R22002 VSS.n5529 VSS.n1246 4.05657
R22003 VSS.n5529 VSS.n1244 4.05657
R22004 VSS.n5533 VSS.n1244 4.05657
R22005 VSS.n5533 VSS.n1242 4.05657
R22006 VSS.n5537 VSS.n1242 4.05657
R22007 VSS.n5537 VSS.n1240 4.05657
R22008 VSS.n5541 VSS.n1240 4.05657
R22009 VSS.n5541 VSS.n1238 4.05657
R22010 VSS.n5545 VSS.n1238 4.05657
R22011 VSS.n5545 VSS.n1236 4.05657
R22012 VSS.n5549 VSS.n1236 4.05657
R22013 VSS.n5549 VSS.n1234 4.05657
R22014 VSS.n5554 VSS.n1234 4.05657
R22015 VSS.n5554 VSS.n1232 4.05657
R22016 VSS.n5559 VSS.n1232 4.05657
R22017 VSS.n5559 VSS.n1230 4.05657
R22018 VSS.n5563 VSS.n1230 4.05657
R22019 VSS.n5563 VSS.n1228 4.05657
R22020 VSS.n5567 VSS.n1228 4.05657
R22021 VSS.n5567 VSS.n1226 4.05657
R22022 VSS.n5571 VSS.n1226 4.05657
R22023 VSS.n5571 VSS.n1224 4.05657
R22024 VSS.n5575 VSS.n1224 4.05657
R22025 VSS.n5575 VSS.n1222 4.05657
R22026 VSS.n5579 VSS.n1222 4.05657
R22027 VSS.n5579 VSS.n1220 4.05657
R22028 VSS.n5583 VSS.n1220 4.05657
R22029 VSS.n5583 VSS.n1218 4.05657
R22030 VSS.n5587 VSS.n1218 4.05657
R22031 VSS.n5587 VSS.n1216 4.05657
R22032 VSS.n5591 VSS.n1216 4.05657
R22033 VSS.n5591 VSS.n1214 4.05657
R22034 VSS.n5595 VSS.n1214 4.05657
R22035 VSS.n5595 VSS.n1212 4.05657
R22036 VSS.n5599 VSS.n1212 4.05657
R22037 VSS.n5599 VSS.n1210 4.05657
R22038 VSS.n5603 VSS.n1210 4.05657
R22039 VSS.n5603 VSS.n1208 4.05657
R22040 VSS.n5607 VSS.n1208 4.05657
R22041 VSS.n5607 VSS.n1206 4.05657
R22042 VSS.n5611 VSS.n1206 4.05657
R22043 VSS.n5611 VSS.n1204 4.05657
R22044 VSS.n5615 VSS.n1204 4.05657
R22045 VSS.n5615 VSS.n1202 4.05657
R22046 VSS.n5619 VSS.n1202 4.05657
R22047 VSS.n5619 VSS.n1200 4.05657
R22048 VSS.n5623 VSS.n1200 4.05657
R22049 VSS.n5623 VSS.n1198 4.05657
R22050 VSS.n5627 VSS.n1198 4.05657
R22051 VSS.n5627 VSS.n1196 4.05657
R22052 VSS.n5631 VSS.n1196 4.05657
R22053 VSS.n5631 VSS.n1194 4.05657
R22054 VSS.n5635 VSS.n1194 4.05657
R22055 VSS.n5635 VSS.n1192 4.05657
R22056 VSS.n5639 VSS.n1192 4.05657
R22057 VSS.n5639 VSS.n1190 4.05657
R22058 VSS.n5643 VSS.n1190 4.05657
R22059 VSS.n5643 VSS.n1188 4.05657
R22060 VSS.n5647 VSS.n1188 4.05657
R22061 VSS.n5647 VSS.n1186 4.05657
R22062 VSS.n5651 VSS.n1186 4.05657
R22063 VSS.n5651 VSS.n1184 4.05657
R22064 VSS.n5655 VSS.n1184 4.05657
R22065 VSS.n5655 VSS.n1182 4.05657
R22066 VSS.n5659 VSS.n1182 4.05657
R22067 VSS.n5659 VSS.n1180 4.05657
R22068 VSS.n5663 VSS.n1180 4.05657
R22069 VSS.n5663 VSS.n1178 4.05657
R22070 VSS.n5667 VSS.n1178 4.05657
R22071 VSS.n5667 VSS.n1176 4.05657
R22072 VSS.n5671 VSS.n1176 4.05657
R22073 VSS.n5671 VSS.n1174 4.05657
R22074 VSS.n5675 VSS.n1174 4.05657
R22075 VSS.n5170 VSS.n5169 3.98035
R22076 VSS.n4283 VSS.n2296 3.8345
R22077 VSS.n4061 VSS.n4058 3.7805
R22078 VSS.n4069 VSS.n4058 3.77031
R22079 VSS.n5313 VSS.n5309 3.68022
R22080 VSS.n4104 VSS.n4103 3.37368
R22081 VSS.n2888 VSS 3.18489
R22082 VSS.n2366 VSS 3.18489
R22083 VSS.n2293 VSS 3.18489
R22084 VSS.n4285 VSS 3.18489
R22085 VSS.n4288 VSS 3.18489
R22086 VSS.n3399 VSS 3.18489
R22087 VSS.n2784 VSS.t3 3.17811
R22088 VSS.n2449 VSS.t43 3.17811
R22089 VSS.n4060 VSS.t45 3.17811
R22090 VSS.n2446 VSS.t17 3.17811
R22091 VSS.n2447 VSS.t15 3.17811
R22092 VSS.n3524 VSS.n2194 3.02469
R22093 VSS.n4055 VSS.n4054 2.95295
R22094 VSS.n5408 VSS.n2103 2.90887
R22095 VSS.n5302 VSS.n5301 2.81187
R22096 VSS.n2192 VSS.n2191 2.81187
R22097 VSS.n4046 VSS.n4045 2.81187
R22098 VSS.n5675 VSS.n5674 2.6005
R22099 VSS.n5673 VSS.n1174 2.6005
R22100 VSS.n1174 VSS.n1173 2.6005
R22101 VSS.n5672 VSS.n5671 2.6005
R22102 VSS.n5671 VSS.n5670 2.6005
R22103 VSS.n1176 VSS.n1175 2.6005
R22104 VSS.n5669 VSS.n1176 2.6005
R22105 VSS.n5667 VSS.n5666 2.6005
R22106 VSS.n5668 VSS.n5667 2.6005
R22107 VSS.n5665 VSS.n1178 2.6005
R22108 VSS.n1178 VSS.n1177 2.6005
R22109 VSS.n5664 VSS.n5663 2.6005
R22110 VSS.n5663 VSS.n5662 2.6005
R22111 VSS.n1180 VSS.n1179 2.6005
R22112 VSS.n5661 VSS.n1180 2.6005
R22113 VSS.n5659 VSS.n5658 2.6005
R22114 VSS.n5660 VSS.n5659 2.6005
R22115 VSS.n5657 VSS.n1182 2.6005
R22116 VSS.n1182 VSS.n1181 2.6005
R22117 VSS.n5656 VSS.n5655 2.6005
R22118 VSS.n5655 VSS.n5654 2.6005
R22119 VSS.n1184 VSS.n1183 2.6005
R22120 VSS.n5653 VSS.n1184 2.6005
R22121 VSS.n5651 VSS.n5650 2.6005
R22122 VSS.n5652 VSS.n5651 2.6005
R22123 VSS.n5649 VSS.n1186 2.6005
R22124 VSS.n1186 VSS.n1185 2.6005
R22125 VSS.n5648 VSS.n5647 2.6005
R22126 VSS.n5647 VSS.n5646 2.6005
R22127 VSS.n1188 VSS.n1187 2.6005
R22128 VSS.n5645 VSS.n1188 2.6005
R22129 VSS.n5643 VSS.n5642 2.6005
R22130 VSS.n5644 VSS.n5643 2.6005
R22131 VSS.n5641 VSS.n1190 2.6005
R22132 VSS.n1190 VSS.n1189 2.6005
R22133 VSS.n5640 VSS.n5639 2.6005
R22134 VSS.n5639 VSS.n5638 2.6005
R22135 VSS.n1192 VSS.n1191 2.6005
R22136 VSS.n5637 VSS.n1192 2.6005
R22137 VSS.n5635 VSS.n5634 2.6005
R22138 VSS.n5636 VSS.n5635 2.6005
R22139 VSS.n5633 VSS.n1194 2.6005
R22140 VSS.n1194 VSS.n1193 2.6005
R22141 VSS.n5632 VSS.n5631 2.6005
R22142 VSS.n5631 VSS.n5630 2.6005
R22143 VSS.n1196 VSS.n1195 2.6005
R22144 VSS.n5629 VSS.n1196 2.6005
R22145 VSS.n5627 VSS.n5626 2.6005
R22146 VSS.n5628 VSS.n5627 2.6005
R22147 VSS.n5625 VSS.n1198 2.6005
R22148 VSS.n1198 VSS.n1197 2.6005
R22149 VSS.n5624 VSS.n5623 2.6005
R22150 VSS.n5623 VSS.n5622 2.6005
R22151 VSS.n1200 VSS.n1199 2.6005
R22152 VSS.n5621 VSS.n1200 2.6005
R22153 VSS.n5619 VSS.n5618 2.6005
R22154 VSS.n5620 VSS.n5619 2.6005
R22155 VSS.n5617 VSS.n1202 2.6005
R22156 VSS.n1202 VSS.n1201 2.6005
R22157 VSS.n5616 VSS.n5615 2.6005
R22158 VSS.n5615 VSS.n5614 2.6005
R22159 VSS.n1204 VSS.n1203 2.6005
R22160 VSS.n5613 VSS.n1204 2.6005
R22161 VSS.n5611 VSS.n5610 2.6005
R22162 VSS.n5612 VSS.n5611 2.6005
R22163 VSS.n5609 VSS.n1206 2.6005
R22164 VSS.n1206 VSS.n1205 2.6005
R22165 VSS.n5608 VSS.n5607 2.6005
R22166 VSS.n5607 VSS.n5606 2.6005
R22167 VSS.n1208 VSS.n1207 2.6005
R22168 VSS.n5605 VSS.n1208 2.6005
R22169 VSS.n5603 VSS.n5602 2.6005
R22170 VSS.n5604 VSS.n5603 2.6005
R22171 VSS.n5601 VSS.n1210 2.6005
R22172 VSS.n1210 VSS.n1209 2.6005
R22173 VSS.n5600 VSS.n5599 2.6005
R22174 VSS.n5599 VSS.n5598 2.6005
R22175 VSS.n1212 VSS.n1211 2.6005
R22176 VSS.n5597 VSS.n1212 2.6005
R22177 VSS.n5595 VSS.n5594 2.6005
R22178 VSS.n5596 VSS.n5595 2.6005
R22179 VSS.n5593 VSS.n1214 2.6005
R22180 VSS.n1214 VSS.n1213 2.6005
R22181 VSS.n5592 VSS.n5591 2.6005
R22182 VSS.n5591 VSS.n5590 2.6005
R22183 VSS.n1216 VSS.n1215 2.6005
R22184 VSS.n5589 VSS.n1216 2.6005
R22185 VSS.n5587 VSS.n5586 2.6005
R22186 VSS.n5588 VSS.n5587 2.6005
R22187 VSS.n5585 VSS.n1218 2.6005
R22188 VSS.n1218 VSS.n1217 2.6005
R22189 VSS.n5584 VSS.n5583 2.6005
R22190 VSS.n5583 VSS.n5582 2.6005
R22191 VSS.n1220 VSS.n1219 2.6005
R22192 VSS.n5581 VSS.n1220 2.6005
R22193 VSS.n5579 VSS.n5578 2.6005
R22194 VSS.n5580 VSS.n5579 2.6005
R22195 VSS.n5577 VSS.n1222 2.6005
R22196 VSS.n1222 VSS.n1221 2.6005
R22197 VSS.n5576 VSS.n5575 2.6005
R22198 VSS.n5575 VSS.n5574 2.6005
R22199 VSS.n1224 VSS.n1223 2.6005
R22200 VSS.n5573 VSS.n1224 2.6005
R22201 VSS.n5571 VSS.n5570 2.6005
R22202 VSS.n5572 VSS.n5571 2.6005
R22203 VSS.n5569 VSS.n1226 2.6005
R22204 VSS.n1226 VSS.n1225 2.6005
R22205 VSS.n5568 VSS.n5567 2.6005
R22206 VSS.n5567 VSS.n5566 2.6005
R22207 VSS.n1228 VSS.n1227 2.6005
R22208 VSS.n5565 VSS.n1228 2.6005
R22209 VSS.n5563 VSS.n5562 2.6005
R22210 VSS.n5564 VSS.n5563 2.6005
R22211 VSS.n5561 VSS.n1230 2.6005
R22212 VSS.n1230 VSS.n1229 2.6005
R22213 VSS.n5560 VSS.n5559 2.6005
R22214 VSS.n5559 VSS.n5558 2.6005
R22215 VSS.n5552 VSS.n1232 2.6005
R22216 VSS.n5556 VSS.n1232 2.6005
R22217 VSS.n5554 VSS.n5553 2.6005
R22218 VSS.n5555 VSS.n5554 2.6005
R22219 VSS.n5551 VSS.n1234 2.6005
R22220 VSS.n1234 VSS.n1233 2.6005
R22221 VSS.n5550 VSS.n5549 2.6005
R22222 VSS.n5549 VSS.n5548 2.6005
R22223 VSS.n1236 VSS.n1235 2.6005
R22224 VSS.n5547 VSS.n1236 2.6005
R22225 VSS.n5545 VSS.n5544 2.6005
R22226 VSS.n5546 VSS.n5545 2.6005
R22227 VSS.n5543 VSS.n1238 2.6005
R22228 VSS.n1238 VSS.n1237 2.6005
R22229 VSS.n5542 VSS.n5541 2.6005
R22230 VSS.n5541 VSS.n5540 2.6005
R22231 VSS.n1240 VSS.n1239 2.6005
R22232 VSS.n5539 VSS.n1240 2.6005
R22233 VSS.n5537 VSS.n5536 2.6005
R22234 VSS.n5538 VSS.n5537 2.6005
R22235 VSS.n5535 VSS.n1242 2.6005
R22236 VSS.n1242 VSS.n1241 2.6005
R22237 VSS.n5534 VSS.n5533 2.6005
R22238 VSS.n5533 VSS.n5532 2.6005
R22239 VSS.n1244 VSS.n1243 2.6005
R22240 VSS.n5531 VSS.n1244 2.6005
R22241 VSS.n5529 VSS.n5528 2.6005
R22242 VSS.n5530 VSS.n5529 2.6005
R22243 VSS.n5527 VSS.n1246 2.6005
R22244 VSS.n1246 VSS.n1245 2.6005
R22245 VSS.n5526 VSS.n5525 2.6005
R22246 VSS.n5525 VSS.n5524 2.6005
R22247 VSS.n1248 VSS.n1247 2.6005
R22248 VSS.n5523 VSS.n1248 2.6005
R22249 VSS.n5521 VSS.n5520 2.6005
R22250 VSS.n5522 VSS.n5521 2.6005
R22251 VSS.n5519 VSS.n1250 2.6005
R22252 VSS.n1250 VSS.n1249 2.6005
R22253 VSS.n5518 VSS.n5517 2.6005
R22254 VSS.n5517 VSS.n5516 2.6005
R22255 VSS.n1252 VSS.n1251 2.6005
R22256 VSS.n5515 VSS.n1252 2.6005
R22257 VSS.n5513 VSS.n5512 2.6005
R22258 VSS.n5514 VSS.n5513 2.6005
R22259 VSS.n5511 VSS.n1254 2.6005
R22260 VSS.n1254 VSS.n1253 2.6005
R22261 VSS.n5510 VSS.n5509 2.6005
R22262 VSS.n5509 VSS.n5508 2.6005
R22263 VSS.n1256 VSS.n1255 2.6005
R22264 VSS.n5507 VSS.n1256 2.6005
R22265 VSS.n5505 VSS.n5504 2.6005
R22266 VSS.n5506 VSS.n5505 2.6005
R22267 VSS.n5503 VSS.n1258 2.6005
R22268 VSS.n1258 VSS.n1257 2.6005
R22269 VSS.n5502 VSS.n5501 2.6005
R22270 VSS.n5501 VSS.n5500 2.6005
R22271 VSS.n1260 VSS.n1259 2.6005
R22272 VSS.n5499 VSS.n1260 2.6005
R22273 VSS.n5497 VSS.n5496 2.6005
R22274 VSS.n5498 VSS.n5497 2.6005
R22275 VSS.n5495 VSS.n1262 2.6005
R22276 VSS.n1262 VSS.n1261 2.6005
R22277 VSS.n5494 VSS.n5493 2.6005
R22278 VSS.n5493 VSS.n5492 2.6005
R22279 VSS.n1264 VSS.n1263 2.6005
R22280 VSS.n5491 VSS.n1264 2.6005
R22281 VSS.n5489 VSS.n5488 2.6005
R22282 VSS.n5490 VSS.n5489 2.6005
R22283 VSS.n5487 VSS.n1266 2.6005
R22284 VSS.n1266 VSS.n1265 2.6005
R22285 VSS.n5486 VSS.n5485 2.6005
R22286 VSS.n5485 VSS.n5484 2.6005
R22287 VSS.n1268 VSS.n1267 2.6005
R22288 VSS.n5483 VSS.n1268 2.6005
R22289 VSS.n5481 VSS.n5480 2.6005
R22290 VSS.n5482 VSS.n5481 2.6005
R22291 VSS.n5479 VSS.n1270 2.6005
R22292 VSS.n1270 VSS.n1269 2.6005
R22293 VSS.n5478 VSS.n5477 2.6005
R22294 VSS.n5477 VSS.n5476 2.6005
R22295 VSS.n1272 VSS.n1271 2.6005
R22296 VSS.n5475 VSS.n1272 2.6005
R22297 VSS.n5473 VSS.n5472 2.6005
R22298 VSS.n5474 VSS.n5473 2.6005
R22299 VSS.n5471 VSS.n1274 2.6005
R22300 VSS.n1274 VSS.n1273 2.6005
R22301 VSS.n5470 VSS.n5469 2.6005
R22302 VSS.n5469 VSS.n5468 2.6005
R22303 VSS.n1276 VSS.n1275 2.6005
R22304 VSS.n5467 VSS.n1276 2.6005
R22305 VSS.n5465 VSS.n5464 2.6005
R22306 VSS.n5466 VSS.n5465 2.6005
R22307 VSS.n5463 VSS.n1278 2.6005
R22308 VSS.n1278 VSS.n1277 2.6005
R22309 VSS.n5462 VSS.n5461 2.6005
R22310 VSS.n5461 VSS.n5460 2.6005
R22311 VSS.n1280 VSS.n1279 2.6005
R22312 VSS.n5459 VSS.n1280 2.6005
R22313 VSS.n5457 VSS.n5456 2.6005
R22314 VSS.n5458 VSS.n5457 2.6005
R22315 VSS.n5455 VSS.n1282 2.6005
R22316 VSS.n1282 VSS.n1281 2.6005
R22317 VSS.n5454 VSS.n5453 2.6005
R22318 VSS.n5453 VSS.n5452 2.6005
R22319 VSS.n1284 VSS.n1283 2.6005
R22320 VSS.n5451 VSS.n1284 2.6005
R22321 VSS.n5449 VSS.n5448 2.6005
R22322 VSS.n5450 VSS.n5449 2.6005
R22323 VSS.n5447 VSS.n1286 2.6005
R22324 VSS.n1286 VSS.n1285 2.6005
R22325 VSS.n5446 VSS.n5445 2.6005
R22326 VSS.n5445 VSS.n5444 2.6005
R22327 VSS.n1288 VSS.n1287 2.6005
R22328 VSS.n5443 VSS.n1288 2.6005
R22329 VSS.n5439 VSS.n1289 2.6005
R22330 VSS.n5238 DVSS 2.57245
R22331 VSS.n5239 VSS.n5238 2.57069
R22332 VSS.n2167 VSS.n18 2.43717
R22333 VSS.n2223 VSS.n2222 2.41753
R22334 VSS.n2223 VSS.n2221 2.41753
R22335 VSS.n2223 VSS.n2220 2.41753
R22336 VSS.n2223 VSS.n2219 2.41753
R22337 VSS.n5268 VSS.n2223 2.41753
R22338 VSS.n5256 VSS.n5255 2.41753
R22339 VSS.n5255 VSS.n2236 2.41753
R22340 VSS.n5255 VSS.n2235 2.41753
R22341 VSS.n5255 VSS.n2234 2.41753
R22342 VSS.n5255 VSS.n2233 2.41753
R22343 VSS.n5255 VSS.n2218 2.41753
R22344 VSS.n5275 VSS.n2209 2.41753
R22345 VSS.n5323 VSS.n5322 2.41274
R22346 VSS.n5324 VSS.n5323 2.41274
R22347 VSS.n5418 VSS.n5417 2.41274
R22348 VSS.n5417 VSS.n5416 2.41274
R22349 VSS.n5238 DVSS 2.32795
R22350 VSS.n4284 VSS.n4283 2.311
R22351 VSS.n4104 VSS.n4092 2.28324
R22352 VSS.n3017 VSS.n3014 2.2728
R22353 VSS.n5412 VSS.n5411 2.25682
R22354 VSS.n5405 VSS.n2104 2.25682
R22355 VSS.n2799 VSS.n2103 2.25392
R22356 VSS.n653 VSS.n358 2.2505
R22357 VSS.n652 VSS.n651 2.2505
R22358 VSS.n650 VSS.n359 2.2505
R22359 VSS.n649 VSS.n648 2.2505
R22360 VSS.n647 VSS.n360 2.2505
R22361 VSS.n646 VSS.n645 2.2505
R22362 VSS.n644 VSS.n361 2.2505
R22363 VSS.n643 VSS.n642 2.2505
R22364 VSS.n641 VSS.n362 2.2505
R22365 VSS.n640 VSS.n639 2.2505
R22366 VSS.n638 VSS.n363 2.2505
R22367 VSS.n637 VSS.n636 2.2505
R22368 VSS.n634 VSS.n364 2.2505
R22369 VSS.n633 VSS.n632 2.2505
R22370 VSS.n537 VSS.n536 2.2505
R22371 VSS.n538 VSS.n534 2.2505
R22372 VSS.n540 VSS.n539 2.2505
R22373 VSS.n541 VSS.n533 2.2505
R22374 VSS.n543 VSS.n542 2.2505
R22375 VSS.n544 VSS.n532 2.2505
R22376 VSS.n546 VSS.n545 2.2505
R22377 VSS.n547 VSS.n531 2.2505
R22378 VSS.n549 VSS.n548 2.2505
R22379 VSS.n550 VSS.n530 2.2505
R22380 VSS.n552 VSS.n551 2.2505
R22381 VSS.n553 VSS.n529 2.2505
R22382 VSS.n555 VSS.n554 2.2505
R22383 VSS.n556 VSS.n528 2.2505
R22384 VSS.n558 VSS.n557 2.2505
R22385 VSS.n559 VSS.n527 2.2505
R22386 VSS.n561 VSS.n560 2.2505
R22387 VSS.n562 VSS.n526 2.2505
R22388 VSS.n564 VSS.n563 2.2505
R22389 VSS.n565 VSS.n525 2.2505
R22390 VSS.n567 VSS.n566 2.2505
R22391 VSS.n568 VSS.n524 2.2505
R22392 VSS.n570 VSS.n569 2.2505
R22393 VSS.n666 VSS.n354 2.2505
R22394 VSS.n668 VSS.n667 2.2505
R22395 VSS.n665 VSS.n353 2.2505
R22396 VSS.n664 VSS.n663 2.2505
R22397 VSS.n662 VSS.n355 2.2505
R22398 VSS.n661 VSS.n660 2.2505
R22399 VSS.n659 VSS.n356 2.2505
R22400 VSS.n658 VSS.n657 2.2505
R22401 VSS.n656 VSS.n357 2.2505
R22402 VSS.n655 VSS.n654 2.2505
R22403 VSS.n105 VSS.n104 2.2505
R22404 VSS.n184 VSS.n183 2.2505
R22405 VSS.n185 VSS.n182 2.2505
R22406 VSS.n187 VSS.n186 2.2505
R22407 VSS.n188 VSS.n181 2.2505
R22408 VSS.n190 VSS.n189 2.2505
R22409 VSS.n191 VSS.n180 2.2505
R22410 VSS.n193 VSS.n192 2.2505
R22411 VSS.n196 VSS.n195 2.2505
R22412 VSS.n197 VSS.n178 2.2505
R22413 VSS.n199 VSS.n198 2.2505
R22414 VSS.n200 VSS.n177 2.2505
R22415 VSS.n202 VSS.n201 2.2505
R22416 VSS.n203 VSS.n176 2.2505
R22417 VSS.n205 VSS.n204 2.2505
R22418 VSS.n206 VSS.n175 2.2505
R22419 VSS.n208 VSS.n207 2.2505
R22420 VSS.n209 VSS.n174 2.2505
R22421 VSS.n211 VSS.n210 2.2505
R22422 VSS.n212 VSS.n173 2.2505
R22423 VSS.n214 VSS.n213 2.2505
R22424 VSS.n215 VSS.n172 2.2505
R22425 VSS.n914 VSS.n913 2.2505
R22426 VSS.n912 VSS.n171 2.2505
R22427 VSS.n233 VSS.n218 2.2505
R22428 VSS.n235 VSS.n234 2.2505
R22429 VSS.n236 VSS.n232 2.2505
R22430 VSS.n238 VSS.n237 2.2505
R22431 VSS.n239 VSS.n231 2.2505
R22432 VSS.n241 VSS.n240 2.2505
R22433 VSS.n242 VSS.n230 2.2505
R22434 VSS.n244 VSS.n243 2.2505
R22435 VSS.n245 VSS.n229 2.2505
R22436 VSS.n247 VSS.n246 2.2505
R22437 VSS.n248 VSS.n228 2.2505
R22438 VSS.n250 VSS.n249 2.2505
R22439 VSS.n251 VSS.n227 2.2505
R22440 VSS.n253 VSS.n252 2.2505
R22441 VSS.n254 VSS.n226 2.2505
R22442 VSS.n256 VSS.n255 2.2505
R22443 VSS.n257 VSS.n225 2.2505
R22444 VSS.n259 VSS.n258 2.2505
R22445 VSS.n260 VSS.n224 2.2505
R22446 VSS.n262 VSS.n261 2.2505
R22447 VSS.n903 VSS.n223 2.2505
R22448 VSS.n905 VSS.n904 2.2505
R22449 VSS.n194 VSS.n179 2.2505
R22450 VSS.n3101 VSS.n3097 2.2505
R22451 VSS.n3130 VSS.n3129 2.2505
R22452 VSS.n3120 VSS.n3119 2.2505
R22453 VSS.n3114 VSS.n3113 2.2505
R22454 VSS.n3061 VSS.n2934 2.2505
R22455 VSS.n3342 VSS.n3341 2.2505
R22456 VSS.n2940 VSS.n2931 2.2505
R22457 VSS.n2938 VSS.n2924 2.2505
R22458 VSS.n3248 VSS.n3147 2.2505
R22459 VSS.n3288 VSS.n3287 2.2505
R22460 VSS.n3145 VSS.n3092 2.2505
R22461 VSS.n3295 VSS.n3294 2.2505
R22462 VSS.n3271 VSS.n3253 2.2505
R22463 VSS.n3263 VSS.n3262 2.2505
R22464 VSS.n3265 VSS.n3264 2.2505
R22465 VSS.n3267 VSS.n3254 2.2505
R22466 VSS.n3270 VSS.n3269 2.2505
R22467 VSS.n3251 VSS.n3250 2.2505
R22468 VSS.n3249 VSS.n3144 2.2505
R22469 VSS.n3289 VSS.n3143 2.2505
R22470 VSS.n3291 VSS.n3290 2.2505
R22471 VSS.n3293 VSS.n3292 2.2505
R22472 VSS.n3142 VSS.n3091 2.2505
R22473 VSS.n3135 VSS.n3134 2.2505
R22474 VSS.n3133 VSS.n3132 2.2505
R22475 VSS.n3131 VSS.n3098 2.2505
R22476 VSS.n3116 VSS.n3099 2.2505
R22477 VSS.n3118 VSS.n3117 2.2505
R22478 VSS.n3115 VSS.n2962 2.2505
R22479 VSS.n3338 VSS.n3337 2.2505
R22480 VSS.n3340 VSS.n3339 2.2505
R22481 VSS.n2943 VSS.n2933 2.2505
R22482 VSS.n2942 VSS.n2941 2.2505
R22483 VSS.n2939 VSS.n2937 2.2505
R22484 VSS.n2936 VSS.n2914 2.2505
R22485 VSS.n3356 VSS.n3355 2.2505
R22486 VSS.n2907 VSS.n2905 2.2505
R22487 VSS.n3361 VSS.n3360 2.2505
R22488 VSS.n2986 VSS.n2906 2.2505
R22489 VSS.n3363 VSS.n3362 2.2505
R22490 VSS.n3017 VSS.n3016 2.2505
R22491 VSS.n3028 VSS.n3027 2.2505
R22492 VSS.n3026 VSS.n3025 2.2505
R22493 VSS.n3023 VSS.n3022 2.2505
R22494 VSS.n3021 VSS.n3020 2.2505
R22495 VSS.n3019 VSS.n3013 2.2505
R22496 VSS.n4283 VSS.n4282 2.2505
R22497 VSS.n2075 VSS.n2074 2.24683
R22498 VSS.n2069 VSS.n2068 2.24683
R22499 VSS.n1819 VSS.n1809 2.24683
R22500 VSS.n5686 VSS.n32 2.24648
R22501 VSS.n5684 VSS.n32 2.24648
R22502 VSS.n1148 VSS.n32 2.24648
R22503 VSS.n1146 VSS.n32 2.24648
R22504 VSS.n1147 VSS.n33 2.24648
R22505 VSS.n1149 VSS.n33 2.24648
R22506 VSS.n5685 VSS.n33 2.24648
R22507 VSS.n5687 VSS.n33 2.24648
R22508 VSS.n3052 VSS.n3051 2.24442
R22509 VSS.n3050 VSS.n3049 2.24442
R22510 VSS.n2076 VSS.n1593 2.24405
R22511 VSS.n2070 VSS.n1594 2.24405
R22512 VSS.n2076 VSS.n1592 2.24405
R22513 VSS.n1812 VSS.n1811 2.24405
R22514 VSS.n1818 VSS.n1814 2.24405
R22515 VSS.n1816 VSS.n1811 2.24405
R22516 VSS.n3005 VSS.n2977 2.24386
R22517 VSS.n3004 VSS.n3003 2.24386
R22518 VSS.n3003 VSS.n2976 2.24386
R22519 VSS.n3305 VSS.n3076 2.24386
R22520 VSS.n3304 VSS.n3303 2.24386
R22521 VSS.n3303 VSS.n3075 2.24386
R22522 VSS.n1604 VSS.n1597 2.24304
R22523 VSS.n2062 VSS.n1596 2.24304
R22524 VSS.n1606 VSS.n1597 2.24304
R22525 VSS.n2062 VSS.n1612 2.24304
R22526 VSS.n1608 VSS.n1597 2.24304
R22527 VSS.n2062 VSS.n1611 2.24304
R22528 VSS.n2063 VSS.n1597 2.24304
R22529 VSS.n2062 VSS.n1610 2.24304
R22530 VSS.n1857 VSS.n1796 2.24304
R22531 VSS.n1854 VSS.n1808 2.24304
R22532 VSS.n1857 VSS.n1795 2.24304
R22533 VSS.n1854 VSS.n1805 2.24304
R22534 VSS.n1857 VSS.n1794 2.24304
R22535 VSS.n1854 VSS.n1802 2.24304
R22536 VSS.n1857 VSS.n1793 2.24304
R22537 VSS.n1855 VSS.n1854 2.24304
R22538 VSS.n4173 VSS.n2403 2.24304
R22539 VSS.n4172 VSS.n2408 2.24304
R22540 VSS.n4176 VSS.n2403 2.24304
R22541 VSS.n4175 VSS.n2408 2.24304
R22542 VSS.n4179 VSS.n2403 2.24304
R22543 VSS.n4178 VSS.n2408 2.24304
R22544 VSS.n4182 VSS.n2403 2.24304
R22545 VSS.n4181 VSS.n2408 2.24304
R22546 VSS.n4184 VSS.n2403 2.24304
R22547 VSS.n2469 VSS.n2462 2.24304
R22548 VSS.n2701 VSS.n2461 2.24304
R22549 VSS.n2471 VSS.n2462 2.24304
R22550 VSS.n2701 VSS.n2698 2.24304
R22551 VSS.n2473 VSS.n2462 2.24304
R22552 VSS.n2701 VSS.n2699 2.24304
R22553 VSS.n2475 VSS.n2462 2.24304
R22554 VSS.n2701 VSS.n2700 2.24304
R22555 VSS.n2702 VSS.n2701 2.24304
R22556 VSS.n4042 VSS.n4026 2.24304
R22557 VSS.n4040 VSS.n0 2.24304
R22558 VSS.n4036 VSS.n0 2.24304
R22559 VSS.n4038 VSS.n4026 2.24304
R22560 VSS.n4034 VSS.n1 2.24304
R22561 VSS.n4030 VSS.n1 2.24304
R22562 VSS.n4032 VSS.n0 2.24304
R22563 VSS.n4028 VSS.n0 2.24304
R22564 VSS.n3138 VSS.n3093 2.24011
R22565 VSS.n3138 VSS.n3136 2.24011
R22566 VSS.n3353 VSS.n2918 2.24011
R22567 VSS.n3353 VSS.n2916 2.24011
R22568 VSS.n2984 VSS.n2912 2.24011
R22569 VSS.n2984 VSS.n2908 2.24011
R22570 VSS.n2917 VSS.n2915 2.24011
R22571 VSS.n2946 VSS.n2945 2.24011
R22572 VSS.n3322 VSS.n2961 2.24011
R22573 VSS.n3140 VSS.n3095 2.24011
R22574 VSS.n3358 VSS.n2910 2.24011
R22575 VSS.n3111 VSS.n3108 2.23777
R22576 VSS.n3109 VSS.n2958 2.23777
R22577 VSS.n3111 VSS.n3110 2.23777
R22578 VSS.n3066 VSS.n3065 2.23777
R22579 VSS.n3068 VSS.n3067 2.23777
R22580 VSS.n3065 VSS.n3060 2.23777
R22581 VSS.n1143 VSS.n1142 2.23644
R22582 VSS.n35 VSS.n34 2.23644
R22583 VSS.n1142 VSS.n38 2.23644
R22584 VSS.n39 VSS.n34 2.23644
R22585 VSS.n1142 VSS.n40 2.23644
R22586 VSS.n41 VSS.n34 2.23644
R22587 VSS.n1142 VSS.n42 2.23644
R22588 VSS.n43 VSS.n34 2.23644
R22589 VSS.n1142 VSS.n44 2.23644
R22590 VSS.n45 VSS.n34 2.23644
R22591 VSS.n1142 VSS.n46 2.23644
R22592 VSS.n47 VSS.n34 2.23644
R22593 VSS.n1142 VSS.n48 2.23644
R22594 VSS.n49 VSS.n34 2.23644
R22595 VSS.n1142 VSS.n50 2.23644
R22596 VSS.n51 VSS.n34 2.23644
R22597 VSS.n1142 VSS.n52 2.23644
R22598 VSS.n53 VSS.n34 2.23644
R22599 VSS.n1142 VSS.n54 2.23644
R22600 VSS.n55 VSS.n34 2.23644
R22601 VSS.n77 VSS.n56 2.23644
R22602 VSS.n1139 VSS.n67 2.23644
R22603 VSS.n77 VSS.n76 2.23644
R22604 VSS.n1139 VSS.n66 2.23644
R22605 VSS.n77 VSS.n75 2.23644
R22606 VSS.n1139 VSS.n65 2.23644
R22607 VSS.n77 VSS.n74 2.23644
R22608 VSS.n1139 VSS.n64 2.23644
R22609 VSS.n77 VSS.n73 2.23644
R22610 VSS.n1139 VSS.n63 2.23644
R22611 VSS.n77 VSS.n72 2.23644
R22612 VSS.n1139 VSS.n62 2.23644
R22613 VSS.n77 VSS.n71 2.23644
R22614 VSS.n1139 VSS.n61 2.23644
R22615 VSS.n77 VSS.n70 2.23644
R22616 VSS.n1139 VSS.n60 2.23644
R22617 VSS.n77 VSS.n69 2.23644
R22618 VSS.n1139 VSS.n59 2.23644
R22619 VSS.n77 VSS.n68 2.23644
R22620 VSS.n1139 VSS.n58 2.23644
R22621 VSS.n3506 VSS.n3390 2.16228
R22622 VSS.n5679 VSS.n1172 2.15282
R22623 VSS.n4250 VSS.n4249 2.12226
R22624 VSS.n4106 VSS.n4105 2.10421
R22625 VSS.n4084 VSS.n2354 2.10097
R22626 VSS.n3873 VSS.n2780 2.07167
R22627 VSS.n5288 VSS.n5287 2.01663
R22628 VSS.n5245 VSS.n5244 1.96906
R22629 VSS.n2785 VSS.n2092 1.94426
R22630 VSS.n4081 VSS.n4080 1.94426
R22631 VSS.n3382 VSS.n2892 1.91475
R22632 VSS.n2891 VSS.n2890 1.91081
R22633 VSS.n4291 VSS.n4290 1.89625
R22634 VSS.n5321 VSS.n5320 1.81109
R22635 VSS.n2792 VSS.n2094 1.81109
R22636 VSS.n2184 VSS.n2180 1.81109
R22637 VSS.n2793 VSS.n2096 1.81109
R22638 VSS.n5426 VSS.n5425 1.80682
R22639 VSS.n3398 VSS 1.7864
R22640 VSS.n3404 VSS 1.7864
R22641 VSS.n5329 VSS.n5328 1.73383
R22642 VSS.n5329 VSS.n11 1.73383
R22643 VSS.n5396 VSS.n5395 1.73383
R22644 VSS.n5395 VSS.n5394 1.73383
R22645 VSS.n2796 VSS.n2098 1.73383
R22646 VSS.n2102 VSS.n2098 1.73383
R22647 VSS.n2086 VSS.n2083 1.73383
R22648 VSS.n2089 VSS.n2083 1.73383
R22649 VSS.n5674 VSS.n8 1.69628
R22650 VSS.n907 VSS.n906 1.66284
R22651 VSS.n5433 VSS.n5432 1.66212
R22652 VSS.n907 VSS.n221 1.64846
R22653 VSS.n5303 VSS.n5302 1.61108
R22654 VSS.n5293 VSS.n2192 1.61108
R22655 VSS.n4046 VSS.n4044 1.61108
R22656 VSS.n4240 VSS.n4239 1.59033
R22657 VSS.n4231 VSS.n2360 1.59033
R22658 VSS.n4222 VSS.n2359 1.59033
R22659 VSS.n2388 VSS.n2357 1.59033
R22660 VSS.n2393 VSS.n2356 1.59033
R22661 VSS.n4203 VSS.n4202 1.59033
R22662 VSS.n4116 VSS.n2431 1.59033
R22663 VSS.n4140 VSS.n4139 1.59033
R22664 VSS.n4130 VSS.n2241 1.59033
R22665 VSS.n2787 VSS.t10 1.57022
R22666 VSS.n3394 VSS.t39 1.57022
R22667 VSS.n3396 VSS.t29 1.57022
R22668 VSS.n2188 VSS.t13 1.57022
R22669 VSS.n2190 VSS.t1 1.57022
R22670 VSS.n4047 VSS.t5 1.57022
R22671 VSS.n4072 VSS.n4071 1.56129
R22672 VSS.n3418 VSS.n3395 1.52301
R22673 VSS.n4092 VSS.n2444 1.51243
R22674 VSS.n5419 DVSS 1.50997
R22675 VSS.n5415 DVSS 1.50997
R22676 VSS.n2181 DVSS 1.50997
R22677 VSS.n5325 DVSS 1.50997
R22678 VSS.n1772 VSS.n1762 1.50734
R22679 VSS.n1787 VSS.n1786 1.50734
R22680 VSS.n1726 VSS.n1724 1.50734
R22681 VSS.n1904 VSS.n1903 1.50734
R22682 VSS.n1702 VSS.n1700 1.50734
R22683 VSS.n1942 VSS.n1941 1.50734
R22684 VSS.n1989 VSS.n1988 1.50734
R22685 VSS.n1974 VSS.n1973 1.50734
R22686 VSS.n2021 VSS.n2020 1.50734
R22687 VSS.n2006 VSS.n2005 1.50734
R22688 VSS.n1628 VSS.n1618 1.50734
R22689 VSS.n1643 VSS.n1642 1.50734
R22690 VSS.n4298 VSS.n4294 1.5055
R22691 VSS.n5133 VSS.n5132 1.5055
R22692 VSS.n5117 VSS.n4294 1.5055
R22693 VSS.n5133 VSS.n2281 1.5055
R22694 VSS.n5316 VSS.n2113 1.50326
R22695 VSS.n3869 VSS.n3868 1.50326
R22696 VSS.n3714 VSS.n2839 1.50157
R22697 VSS.n3534 VSS.n3533 1.5005
R22698 VSS.n3536 VSS.n3535 1.5005
R22699 VSS.n3538 VSS.n3537 1.5005
R22700 VSS.n3540 VSS.n3539 1.5005
R22701 VSS.n3542 VSS.n3541 1.5005
R22702 VSS.n3544 VSS.n3543 1.5005
R22703 VSS.n3546 VSS.n3545 1.5005
R22704 VSS.n3548 VSS.n3547 1.5005
R22705 VSS.n3531 VSS.n2884 1.5005
R22706 VSS.n1641 VSS.n1634 1.5005
R22707 VSS.n2039 VSS.n2038 1.5005
R22708 VSS.n1632 VSS.n1626 1.5005
R22709 VSS.n2046 VSS.n2045 1.5005
R22710 VSS.n1627 VSS.n1623 1.5005
R22711 VSS.n1663 VSS.n1661 1.5005
R22712 VSS.n2010 VSS.n2009 1.5005
R22713 VSS.n1731 VSS.n1658 1.5005
R22714 VSS.n1730 VSS.n1651 1.5005
R22715 VSS.n2019 VSS.n2018 1.5005
R22716 VSS.n1688 VSS.n1686 1.5005
R22717 VSS.n1978 VSS.n1977 1.5005
R22718 VSS.n1737 VSS.n1683 1.5005
R22719 VSS.n1736 VSS.n1678 1.5005
R22720 VSS.n1987 VSS.n1986 1.5005
R22721 VSS.n1936 VSS.n1715 1.5005
R22722 VSS.n1938 VSS.n1708 1.5005
R22723 VSS.n1951 VSS.n1950 1.5005
R22724 VSS.n1706 VSS.n1703 1.5005
R22725 VSS.n1957 VSS.n1956 1.5005
R22726 VSS.n1898 VSS.n1757 1.5005
R22727 VSS.n1900 VSS.n1750 1.5005
R22728 VSS.n1913 VSS.n1912 1.5005
R22729 VSS.n1748 VSS.n1727 1.5005
R22730 VSS.n1919 VSS.n1918 1.5005
R22731 VSS.n1785 VSS.n1778 1.5005
R22732 VSS.n1874 VSS.n1873 1.5005
R22733 VSS.n1776 VSS.n1770 1.5005
R22734 VSS.n1881 VSS.n1880 1.5005
R22735 VSS.n1771 VSS.n1767 1.5005
R22736 VSS.n5693 VSS.n5692 1.5005
R22737 VSS.n21 VSS.n17 1.5005
R22738 VSS.n1151 VSS.n1150 1.5005
R22739 VSS.n1153 VSS.n1152 1.5005
R22740 VSS.n1155 VSS.n1154 1.5005
R22741 VSS.n1157 VSS.n1156 1.5005
R22742 VSS.n1159 VSS.n1158 1.5005
R22743 VSS.n1161 VSS.n1160 1.5005
R22744 VSS.n1163 VSS.n1162 1.5005
R22745 VSS.n1165 VSS.n1164 1.5005
R22746 VSS.n1167 VSS.n1166 1.5005
R22747 VSS.n1168 VSS.n31 1.5005
R22748 VSS.n4883 VSS.n4882 1.5005
R22749 VSS.n4881 VSS.n2283 1.5005
R22750 VSS.n5132 VSS.n5131 1.5005
R22751 VSS.n4885 VSS.n4884 1.5005
R22752 VSS.n4880 VSS.n4622 1.5005
R22753 VSS.n4608 VSS.n4607 1.5005
R22754 VSS.n4895 VSS.n4894 1.5005
R22755 VSS.n4897 VSS.n4896 1.5005
R22756 VSS.n4606 VSS.n4602 1.5005
R22757 VSS.n4605 VSS.n4604 1.5005
R22758 VSS.n4590 VSS.n4589 1.5005
R22759 VSS.n4907 VSS.n4906 1.5005
R22760 VSS.n4910 VSS.n4909 1.5005
R22761 VSS.n4588 VSS.n4586 1.5005
R22762 VSS.n4573 VSS.n4571 1.5005
R22763 VSS.n4920 VSS.n4919 1.5005
R22764 VSS.n4921 VSS.n4569 1.5005
R22765 VSS.n4923 VSS.n4922 1.5005
R22766 VSS.n4570 VSS.n4568 1.5005
R22767 VSS.n4555 VSS.n4554 1.5005
R22768 VSS.n4933 VSS.n4932 1.5005
R22769 VSS.n4935 VSS.n4934 1.5005
R22770 VSS.n4553 VSS.n4551 1.5005
R22771 VSS.n4629 VSS.n4538 1.5005
R22772 VSS.n4944 VSS.n4537 1.5005
R22773 VSS.n4946 VSS.n4945 1.5005
R22774 VSS.n4948 VSS.n4947 1.5005
R22775 VSS.n4536 VSS.n4533 1.5005
R22776 VSS.n4535 VSS.n4520 1.5005
R22777 VSS.n4958 VSS.n4957 1.5005
R22778 VSS.n4960 VSS.n4959 1.5005
R22779 VSS.n4519 VSS.n4514 1.5005
R22780 VSS.n4518 VSS.n4517 1.5005
R22781 VSS.n4502 VSS.n4501 1.5005
R22782 VSS.n4970 VSS.n4969 1.5005
R22783 VSS.n4972 VSS.n4971 1.5005
R22784 VSS.n4499 VSS.n4497 1.5005
R22785 VSS.n4484 VSS.n4483 1.5005
R22786 VSS.n4982 VSS.n4981 1.5005
R22787 VSS.n4984 VSS.n4983 1.5005
R22788 VSS.n4482 VSS.n4477 1.5005
R22789 VSS.n4481 VSS.n4480 1.5005
R22790 VSS.n4465 VSS.n4464 1.5005
R22791 VSS.n4994 VSS.n4993 1.5005
R22792 VSS.n4996 VSS.n4995 1.5005
R22793 VSS.n4463 VSS.n4461 1.5005
R22794 VSS.n4450 VSS.n4449 1.5005
R22795 VSS.n5006 VSS.n5005 1.5005
R22796 VSS.n5008 VSS.n5007 1.5005
R22797 VSS.n5010 VSS.n5009 1.5005
R22798 VSS.n5012 VSS.n5011 1.5005
R22799 VSS.n4445 VSS.n4442 1.5005
R22800 VSS.n4444 VSS.n4429 1.5005
R22801 VSS.n5022 VSS.n5021 1.5005
R22802 VSS.n5024 VSS.n5023 1.5005
R22803 VSS.n4428 VSS.n4423 1.5005
R22804 VSS.n4427 VSS.n4426 1.5005
R22805 VSS.n4411 VSS.n4410 1.5005
R22806 VSS.n5034 VSS.n5033 1.5005
R22807 VSS.n5036 VSS.n5035 1.5005
R22808 VSS.n4409 VSS.n4407 1.5005
R22809 VSS.n4394 VSS.n4393 1.5005
R22810 VSS.n5046 VSS.n5045 1.5005
R22811 VSS.n5048 VSS.n5047 1.5005
R22812 VSS.n4392 VSS.n4387 1.5005
R22813 VSS.n4391 VSS.n4390 1.5005
R22814 VSS.n4375 VSS.n4374 1.5005
R22815 VSS.n5058 VSS.n5057 1.5005
R22816 VSS.n5060 VSS.n5059 1.5005
R22817 VSS.n4373 VSS.n4371 1.5005
R22818 VSS.n4360 VSS.n4359 1.5005
R22819 VSS.n5070 VSS.n5069 1.5005
R22820 VSS.n5072 VSS.n5071 1.5005
R22821 VSS.n5074 VSS.n5073 1.5005
R22822 VSS.n5076 VSS.n5075 1.5005
R22823 VSS.n4356 VSS.n4353 1.5005
R22824 VSS.n4355 VSS.n4340 1.5005
R22825 VSS.n5086 VSS.n5085 1.5005
R22826 VSS.n5088 VSS.n5087 1.5005
R22827 VSS.n4339 VSS.n4335 1.5005
R22828 VSS.n4338 VSS.n4337 1.5005
R22829 VSS.n4323 VSS.n4322 1.5005
R22830 VSS.n5098 VSS.n5097 1.5005
R22831 VSS.n5100 VSS.n5099 1.5005
R22832 VSS.n4321 VSS.n4319 1.5005
R22833 VSS.n4303 VSS.n4301 1.5005
R22834 VSS.n5110 VSS.n5109 1.5005
R22835 VSS.n5111 VSS.n4299 1.5005
R22836 VSS.n5113 VSS.n5112 1.5005
R22837 VSS.n4300 VSS.n4298 1.5005
R22838 VSS.n4873 VSS.n4625 1.5005
R22839 VSS.n2284 VSS.n2281 1.5005
R22840 VSS.n5118 VSS.n5117 1.5005
R22841 VSS.n4295 VSS.n4293 1.5005
R22842 VSS.n4648 VSS.n4647 1.5005
R22843 VSS.n4652 VSS.n4651 1.5005
R22844 VSS.n4654 VSS.n4653 1.5005
R22845 VSS.n4657 VSS.n4656 1.5005
R22846 VSS.n4659 VSS.n4658 1.5005
R22847 VSS.n4663 VSS.n4662 1.5005
R22848 VSS.n4665 VSS.n4664 1.5005
R22849 VSS.n4666 VSS.n4644 1.5005
R22850 VSS.n4668 VSS.n4667 1.5005
R22851 VSS.n4670 VSS.n4669 1.5005
R22852 VSS.n4674 VSS.n4673 1.5005
R22853 VSS.n4676 VSS.n4675 1.5005
R22854 VSS.n4679 VSS.n4678 1.5005
R22855 VSS.n4680 VSS.n4643 1.5005
R22856 VSS.n4683 VSS.n4682 1.5005
R22857 VSS.n4642 VSS.n4641 1.5005
R22858 VSS.n4694 VSS.n4693 1.5005
R22859 VSS.n4696 VSS.n4695 1.5005
R22860 VSS.n4699 VSS.n4698 1.5005
R22861 VSS.n4701 VSS.n4700 1.5005
R22862 VSS.n4705 VSS.n4704 1.5005
R22863 VSS.n4707 VSS.n4706 1.5005
R22864 VSS.n4709 VSS.n4708 1.5005
R22865 VSS.n4711 VSS.n4710 1.5005
R22866 VSS.n4713 VSS.n4712 1.5005
R22867 VSS.n4717 VSS.n4716 1.5005
R22868 VSS.n4719 VSS.n4718 1.5005
R22869 VSS.n4722 VSS.n4721 1.5005
R22870 VSS.n4724 VSS.n4723 1.5005
R22871 VSS.n4728 VSS.n4727 1.5005
R22872 VSS.n4730 VSS.n4729 1.5005
R22873 VSS.n4731 VSS.n4637 1.5005
R22874 VSS.n4734 VSS.n4733 1.5005
R22875 VSS.n4736 VSS.n4735 1.5005
R22876 VSS.n4740 VSS.n4739 1.5005
R22877 VSS.n4742 VSS.n4741 1.5005
R22878 VSS.n4745 VSS.n4744 1.5005
R22879 VSS.n4746 VSS.n4636 1.5005
R22880 VSS.n4750 VSS.n4749 1.5005
R22881 VSS.n4635 VSS.n4634 1.5005
R22882 VSS.n4761 VSS.n4760 1.5005
R22883 VSS.n4763 VSS.n4762 1.5005
R22884 VSS.n4766 VSS.n4765 1.5005
R22885 VSS.n4768 VSS.n4767 1.5005
R22886 VSS.n4772 VSS.n4771 1.5005
R22887 VSS.n4774 VSS.n4773 1.5005
R22888 VSS.n4776 VSS.n4775 1.5005
R22889 VSS.n4778 VSS.n4777 1.5005
R22890 VSS.n4780 VSS.n4779 1.5005
R22891 VSS.n4784 VSS.n4783 1.5005
R22892 VSS.n4786 VSS.n4785 1.5005
R22893 VSS.n4789 VSS.n4788 1.5005
R22894 VSS.n4792 VSS.n4791 1.5005
R22895 VSS.n4796 VSS.n4795 1.5005
R22896 VSS.n4798 VSS.n4797 1.5005
R22897 VSS.n4799 VSS.n4632 1.5005
R22898 VSS.n4802 VSS.n4801 1.5005
R22899 VSS.n4804 VSS.n4803 1.5005
R22900 VSS.n4808 VSS.n4807 1.5005
R22901 VSS.n4810 VSS.n4809 1.5005
R22902 VSS.n4813 VSS.n4812 1.5005
R22903 VSS.n4815 VSS.n4814 1.5005
R22904 VSS.n4818 VSS.n4631 1.5005
R22905 VSS.n4820 VSS.n4819 1.5005
R22906 VSS.n4823 VSS.n4822 1.5005
R22907 VSS.n4826 VSS.n4825 1.5005
R22908 VSS.n4828 VSS.n4827 1.5005
R22909 VSS.n4832 VSS.n4831 1.5005
R22910 VSS.n4834 VSS.n4833 1.5005
R22911 VSS.n4837 VSS.n4836 1.5005
R22912 VSS.n4839 VSS.n4838 1.5005
R22913 VSS.n4840 VSS.n4628 1.5005
R22914 VSS.n4844 VSS.n4843 1.5005
R22915 VSS.n4846 VSS.n4845 1.5005
R22916 VSS.n4849 VSS.n4848 1.5005
R22917 VSS.n4851 VSS.n4850 1.5005
R22918 VSS.n4855 VSS.n4854 1.5005
R22919 VSS.n4857 VSS.n4856 1.5005
R22920 VSS.n4858 VSS.n4626 1.5005
R22921 VSS.n4860 VSS.n4859 1.5005
R22922 VSS.n4862 VSS.n4861 1.5005
R22923 VSS.n4866 VSS.n4865 1.5005
R22924 VSS.n4868 VSS.n4867 1.5005
R22925 VSS.n4871 VSS.n4870 1.5005
R22926 VSS.n4872 VSS.n4623 1.5005
R22927 VSS.n4875 VSS.n4874 1.5005
R22928 VSS.n4624 VSS.n2280 1.5005
R22929 VSS.n4878 VSS.n4876 1.5005
R22930 VSS.n4887 VSS.n4619 1.5005
R22931 VSS.n4869 VSS.n4611 1.5005
R22932 VSS.n4892 VSS.n4610 1.5005
R22933 VSS.n4864 VSS.n4863 1.5005
R22934 VSS.n4899 VSS.n4600 1.5005
R22935 VSS.n4858 VSS.n4593 1.5005
R22936 VSS.n4904 VSS.n4592 1.5005
R22937 VSS.n4853 VSS.n4852 1.5005
R22938 VSS.n4912 VSS.n4583 1.5005
R22939 VSS.n4847 VSS.n4576 1.5005
R22940 VSS.n4917 VSS.n4575 1.5005
R22941 VSS.n4842 VSS.n4841 1.5005
R22942 VSS.n4925 VSS.n4565 1.5005
R22943 VSS.n4835 VSS.n4558 1.5005
R22944 VSS.n4930 VSS.n4557 1.5005
R22945 VSS.n4830 VSS.n4829 1.5005
R22946 VSS.n4937 VSS.n4548 1.5005
R22947 VSS.n4824 VSS.n4541 1.5005
R22948 VSS.n4942 VSS.n4540 1.5005
R22949 VSS.n4817 VSS.n4816 1.5005
R22950 VSS.n4950 VSS.n4530 1.5005
R22951 VSS.n4811 VSS.n4523 1.5005
R22952 VSS.n4955 VSS.n4522 1.5005
R22953 VSS.n4806 VSS.n4805 1.5005
R22954 VSS.n4962 VSS.n4512 1.5005
R22955 VSS.n4800 VSS.n4505 1.5005
R22956 VSS.n4967 VSS.n4504 1.5005
R22957 VSS.n4794 VSS.n4793 1.5005
R22958 VSS.n4974 VSS.n4494 1.5005
R22959 VSS.n4787 VSS.n4487 1.5005
R22960 VSS.n4979 VSS.n4486 1.5005
R22961 VSS.n4782 VSS.n4781 1.5005
R22962 VSS.n4986 VSS.n4475 1.5005
R22963 VSS.n4633 VSS.n4468 1.5005
R22964 VSS.n4991 VSS.n4467 1.5005
R22965 VSS.n4770 VSS.n4769 1.5005
R22966 VSS.n4998 VSS.n4458 1.5005
R22967 VSS.n4764 VSS.n4453 1.5005
R22968 VSS.n5003 VSS.n4452 1.5005
R22969 VSS.n4759 VSS.n4758 1.5005
R22970 VSS.n4752 VSS.n4751 1.5005
R22971 VSS.n5014 VSS.n4439 1.5005
R22972 VSS.n4743 VSS.n4432 1.5005
R22973 VSS.n5019 VSS.n4431 1.5005
R22974 VSS.n4738 VSS.n4737 1.5005
R22975 VSS.n5026 VSS.n4421 1.5005
R22976 VSS.n4732 VSS.n4414 1.5005
R22977 VSS.n5031 VSS.n4413 1.5005
R22978 VSS.n4726 VSS.n4725 1.5005
R22979 VSS.n5038 VSS.n4404 1.5005
R22980 VSS.n4720 VSS.n4397 1.5005
R22981 VSS.n5043 VSS.n4396 1.5005
R22982 VSS.n4715 VSS.n4714 1.5005
R22983 VSS.n5050 VSS.n4385 1.5005
R22984 VSS.n4640 VSS.n4378 1.5005
R22985 VSS.n5055 VSS.n4377 1.5005
R22986 VSS.n4703 VSS.n4702 1.5005
R22987 VSS.n5062 VSS.n4368 1.5005
R22988 VSS.n4697 VSS.n4363 1.5005
R22989 VSS.n5067 VSS.n4362 1.5005
R22990 VSS.n4692 VSS.n4691 1.5005
R22991 VSS.n4685 VSS.n4684 1.5005
R22992 VSS.n5078 VSS.n4350 1.5005
R22993 VSS.n4677 VSS.n4343 1.5005
R22994 VSS.n5083 VSS.n4342 1.5005
R22995 VSS.n4672 VSS.n4671 1.5005
R22996 VSS.n5090 VSS.n4333 1.5005
R22997 VSS.n4666 VSS.n4326 1.5005
R22998 VSS.n5095 VSS.n4325 1.5005
R22999 VSS.n4661 VSS.n4660 1.5005
R23000 VSS.n5102 VSS.n4316 1.5005
R23001 VSS.n4655 VSS.n4306 1.5005
R23002 VSS.n5107 VSS.n4305 1.5005
R23003 VSS.n4650 VSS.n4649 1.5005
R23004 VSS.n5116 VSS.n5115 1.5005
R23005 VSS.n2282 VSS.n2280 1.5005
R23006 VSS.n4879 VSS.n4878 1.5005
R23007 VSS.n4887 VSS.n4886 1.5005
R23008 VSS.n4621 VSS.n4611 1.5005
R23009 VSS.n4893 VSS.n4892 1.5005
R23010 VSS.n4863 VSS.n4603 1.5005
R23011 VSS.n4899 VSS.n4898 1.5005
R23012 VSS.n4604 VSS.n4593 1.5005
R23013 VSS.n4905 VSS.n4904 1.5005
R23014 VSS.n4852 VSS.n4587 1.5005
R23015 VSS.n4912 VSS.n4911 1.5005
R23016 VSS.n4585 VSS.n4576 1.5005
R23017 VSS.n4918 VSS.n4917 1.5005
R23018 VSS.n4841 VSS.n4572 1.5005
R23019 VSS.n4925 VSS.n4924 1.5005
R23020 VSS.n4567 VSS.n4558 1.5005
R23021 VSS.n4931 VSS.n4930 1.5005
R23022 VSS.n4829 VSS.n4552 1.5005
R23023 VSS.n4937 VSS.n4936 1.5005
R23024 VSS.n4550 VSS.n4541 1.5005
R23025 VSS.n4943 VSS.n4942 1.5005
R23026 VSS.n4816 VSS.n4534 1.5005
R23027 VSS.n4950 VSS.n4949 1.5005
R23028 VSS.n4532 VSS.n4523 1.5005
R23029 VSS.n4956 VSS.n4955 1.5005
R23030 VSS.n4805 VSS.n4515 1.5005
R23031 VSS.n4962 VSS.n4961 1.5005
R23032 VSS.n4516 VSS.n4505 1.5005
R23033 VSS.n4968 VSS.n4967 1.5005
R23034 VSS.n4793 VSS.n4498 1.5005
R23035 VSS.n4974 VSS.n4973 1.5005
R23036 VSS.n4496 VSS.n4487 1.5005
R23037 VSS.n4980 VSS.n4979 1.5005
R23038 VSS.n4781 VSS.n4478 1.5005
R23039 VSS.n4986 VSS.n4985 1.5005
R23040 VSS.n4479 VSS.n4468 1.5005
R23041 VSS.n4992 VSS.n4991 1.5005
R23042 VSS.n4769 VSS.n4462 1.5005
R23043 VSS.n4998 VSS.n4997 1.5005
R23044 VSS.n4460 VSS.n4453 1.5005
R23045 VSS.n5004 VSS.n5003 1.5005
R23046 VSS.n4758 VSS.n4447 1.5005
R23047 VSS.n4752 VSS.n4443 1.5005
R23048 VSS.n5014 VSS.n5013 1.5005
R23049 VSS.n4441 VSS.n4432 1.5005
R23050 VSS.n5020 VSS.n5019 1.5005
R23051 VSS.n4737 VSS.n4424 1.5005
R23052 VSS.n5026 VSS.n5025 1.5005
R23053 VSS.n4425 VSS.n4414 1.5005
R23054 VSS.n5032 VSS.n5031 1.5005
R23055 VSS.n4725 VSS.n4408 1.5005
R23056 VSS.n5038 VSS.n5037 1.5005
R23057 VSS.n4406 VSS.n4397 1.5005
R23058 VSS.n5044 VSS.n5043 1.5005
R23059 VSS.n4714 VSS.n4388 1.5005
R23060 VSS.n5050 VSS.n5049 1.5005
R23061 VSS.n4389 VSS.n4378 1.5005
R23062 VSS.n5056 VSS.n5055 1.5005
R23063 VSS.n4702 VSS.n4372 1.5005
R23064 VSS.n5062 VSS.n5061 1.5005
R23065 VSS.n4370 VSS.n4363 1.5005
R23066 VSS.n5068 VSS.n5067 1.5005
R23067 VSS.n4691 VSS.n4358 1.5005
R23068 VSS.n4685 VSS.n4354 1.5005
R23069 VSS.n5078 VSS.n5077 1.5005
R23070 VSS.n4352 VSS.n4343 1.5005
R23071 VSS.n5084 VSS.n5083 1.5005
R23072 VSS.n4671 VSS.n4336 1.5005
R23073 VSS.n5090 VSS.n5089 1.5005
R23074 VSS.n4337 VSS.n4326 1.5005
R23075 VSS.n5096 VSS.n5095 1.5005
R23076 VSS.n4660 VSS.n4320 1.5005
R23077 VSS.n5102 VSS.n5101 1.5005
R23078 VSS.n4318 VSS.n4306 1.5005
R23079 VSS.n5108 VSS.n5107 1.5005
R23080 VSS.n4649 VSS.n4302 1.5005
R23081 VSS.n5115 VSS.n5114 1.5005
R23082 VSS.n3031 VSS.n2838 1.5005
R23083 VSS.n3033 VSS.n3032 1.5005
R23084 VSS.n3035 VSS.n3034 1.5005
R23085 VSS.n3037 VSS.n3036 1.5005
R23086 VSS.n3039 VSS.n3038 1.5005
R23087 VSS.n3041 VSS.n3040 1.5005
R23088 VSS.n3043 VSS.n3042 1.5005
R23089 VSS.n3045 VSS.n3044 1.5005
R23090 VSS.n3047 VSS.n3046 1.5005
R23091 VSS.n3530 VSS.n2886 1.49818
R23092 VSS.n4091 VSS.n4082 1.49138
R23093 VSS.n3873 VSS.n3872 1.48621
R23094 VSS.n3312 VSS.n3311 1.44688
R23095 VSS.n3071 VSS.n3070 1.44688
R23096 VSS.n5401 VSS.n5400 1.39741
R23097 VSS.n5440 VSS.n5439 1.38866
R23098 VSS.n3029 VSS.n2969 1.35477
R23099 VSS.n3258 VSS.n2970 1.35477
R23100 VSS.n5242 DVSS 1.35085
R23101 VSS.n4078 VSS.n2456 1.328
R23102 VSS.n2377 VSS.n2372 1.31286
R23103 VSS.n4086 VSS.n2398 1.31286
R23104 VSS.n4147 VSS.n4146 1.31286
R23105 VSS.n2244 VSS.n2242 1.31286
R23106 VSS.n2185 VSS.n2184 1.3005
R23107 VSS.n5320 VSS.n5319 1.3005
R23108 VSS.n2793 VSS.n2782 1.3005
R23109 VSS.n2792 VSS.n2781 1.3005
R23110 VSS.n4050 VSS.n4049 1.3005
R23111 VSS.n5295 VSS.n5294 1.3005
R23112 VSS.n5300 VSS.n5299 1.3005
R23113 VSS.n3417 VSS.n3416 1.3005
R23114 VSS.n3507 VSS.n3506 1.3005
R23115 VSS.n2450 VSS 1.28985
R23116 VSS.n5338 VSS.n2173 1.26649
R23117 VSS.n4220 VSS.n2358 1.25594
R23118 VSS.n4117 VSS.n2432 1.25594
R23119 DVSS VSS.n3407 1.23516
R23120 VSS.n3407 DVSS 1.23404
R23121 VSS.n2087 VSS.n2086 1.23176
R23122 VSS.n5328 VSS.n2174 1.23176
R23123 VSS.n5397 VSS.n5396 1.23176
R23124 VSS.n2797 VSS.n2796 1.23176
R23125 VSS.n3951 VSS.n2189 1.19925
R23126 VSS.n5244 VSS.n5243 1.16402
R23127 VSS.n2084 VSS.n2082 1.15745
R23128 VSS.n4090 VSS.n4089 1.15606
R23129 VSS.n5411 VSS.n5410 1.15606
R23130 VSS.n5405 VSS.n5404 1.15606
R23131 VSS.n3381 VSS.n3380 1.13009
R23132 VSS.n4105 VSS.n2238 1.10843
R23133 VSS.n4146 VSS.n2427 1.10563
R23134 VSS.n2242 VSS.n2240 1.10563
R23135 VSS.n2372 VSS.n2371 1.10563
R23136 VSS.n4087 VSS.n4086 1.10563
R23137 VSS.n2888 VSS.t32 1.0925
R23138 VSS.n2366 VSS.t21 1.0925
R23139 VSS.n2293 VSS.t36 1.0925
R23140 VSS.n2293 VSS.t19 1.0925
R23141 VSS.n4285 VSS.t34 1.0925
R23142 VSS.n4285 VSS.t23 1.0925
R23143 VSS.n4288 VSS.t25 1.0925
R23144 VSS.n3399 VSS.t27 1.0925
R23145 VSS.n2175 VSS.n2113 1.08844
R23146 VSS.n5390 VSS.n2113 1.08844
R23147 VSS.n3868 VSS.n3867 1.08844
R23148 VSS.n3868 VSS.n2088 1.08844
R23149 VSS.n5428 VSS.n2088 1.0805
R23150 VSS.n5335 VSS.n2175 1.0805
R23151 VSS.n5391 VSS.n5390 1.0805
R23152 VSS.n3867 VSS.n2801 1.0805
R23153 VSS.n5244 VSS.n2238 1.07932
R23154 VSS.n2077 VSS.n1591 1.07349
R23155 VSS.n3383 VSS.n3382 1.07241
R23156 VSS.n2909 VSS.n2413 1.05604
R23157 VSS.n2790 VSS.n2789 1.05029
R23158 VSS.n2454 VSS.n2453 1.0405
R23159 VSS.n2453 VSS.n2452 1.0405
R23160 VSS.n2458 VSS.n2445 1.0405
R23161 VSS.n4074 VSS.n4073 1.0405
R23162 VSS.n4075 VSS.n4074 1.0405
R23163 VSS.n4067 VSS.n4066 1.0405
R23164 VSS.n4066 VSS.n4065 1.0405
R23165 VSS.n5326 VSS.n5325 1.0405
R23166 VSS.n5326 VSS.n2176 1.0405
R23167 VSS.n2181 VSS.n2110 1.0405
R23168 VSS.n2112 VSS.n2110 1.0405
R23169 VSS.n5415 VSS.n5414 1.0405
R23170 VSS.n5414 VSS.n5413 1.0405
R23171 VSS.n5420 VSS.n5419 1.0405
R23172 VSS.n5421 VSS.n5420 1.0405
R23173 VSS.n2783 VSS.t2 1.0405
R23174 VSS.n2452 VSS.t42 1.00732
R23175 VSS.t16 VSS.n2458 1.00732
R23176 VSS.t14 VSS.n4075 1.00732
R23177 VSS.n4065 VSS.t44 1.00732
R23178 VSS.n2432 VSS.n2239 1.00517
R23179 VSS.n2358 VSS.n2353 1.00517
R23180 VSS.n4249 VSS 1.00241
R23181 VSS.n4070 VSS.n4069 0.998789
R23182 VSS.n4080 VSS.n2445 0.996088
R23183 VSS.n2785 VSS.n2783 0.996088
R23184 VSS.n5243 VSS.n5239 0.992621
R23185 VSS.n2313 VSS.n2312 0.988551
R23186 VSS.n5429 DVSS 0.972907
R23187 VSS.n5336 DVSS 0.972907
R23188 VSS.n2108 DVSS 0.972907
R23189 VSS.n5430 VSS.n2087 0.971611
R23190 VSS.n5337 VSS.n2174 0.971611
R23191 VSS.n5398 VSS.n5397 0.971611
R23192 VSS.n2798 VSS.n2797 0.971611
R23193 VSS.n4249 VSS.n4248 0.945955
R23194 VSS.n4052 VSS.n4051 0.945955
R23195 VSS.n2189 VSS.n2111 0.945955
R23196 VSS.n5314 VSS.n5313 0.945955
R23197 VSS.n5409 VSS.n5408 0.945955
R23198 VSS.n2800 DVSS 0.92317
R23199 VSS.n2689 VSS.n7 0.922787
R23200 VSS.n5702 VSS.n5701 0.922694
R23201 VSS.n3438 VSS.n1291 0.922457
R23202 VSS.n3403 VSS.n3402 0.910322
R23203 VSS.n1587 VSS.n1296 0.902282
R23204 VSS.n1588 VSS.n1587 0.902198
R23205 VSS.n1588 VSS.n1297 0.902161
R23206 VSS.n1297 VSS.n1296 0.901878
R23207 VSS.n1591 VSS.n1590 0.879171
R23208 VSS.n5682 VSS.n1169 0.879171
R23209 VSS.n5340 VSS.n5339 0.875955
R23210 VSS.n5389 VSS.n5388 0.875955
R23211 VSS.n3866 VSS.n3865 0.875955
R23212 VSS.n4103 VSS.n2428 0.875366
R23213 VSS.n4106 VSS.n2429 0.875366
R23214 VSS.n5246 VSS.n5245 0.875366
R23215 VSS.n2890 VSS.n2296 0.873402
R23216 VSS.n1169 VSS.n1168 0.870066
R23217 VSS.n4242 VSS.n2361 0.867167
R23218 VSS.n4247 VSS.n4246 0.867167
R23219 VSS.n4144 VSS.n2430 0.867167
R23220 VSS.n5249 VSS.n5248 0.867167
R23221 VSS.n4068 VSS.n4067 0.843937
R23222 VSS.n4073 VSS.n4072 0.843937
R23223 VSS.n2455 VSS.n2454 0.843937
R23224 VSS.n4105 VSS.n4104 0.827218
R23225 VSS.n1145 VSS.n1144 0.820816
R23226 VSS.n4071 VSS.n2456 0.815237
R23227 VSS.n3730 VSS.n2088 0.803519
R23228 VSS.n5308 VSS.n2175 0.803519
R23229 VSS.n5390 VSS.n5389 0.803519
R23230 VSS.n3867 VSS.n3866 0.803519
R23231 VSS.n5339 DVSS 0.801151
R23232 VSS.n5424 VSS.n2090 0.8005
R23233 VSS.n3510 VSS.n3391 0.796907
R23234 VSS.n3514 VSS.n3391 0.796907
R23235 VSS.n3514 VSS.n3389 0.796907
R23236 VSS.n3518 VSS.n3389 0.796907
R23237 VSS.n3518 VSS.n3387 0.796907
R23238 VSS.n3522 VSS.n3387 0.796907
R23239 VSS.n3522 VSS.n2196 0.796907
R23240 VSS.n5286 VSS.n2196 0.796907
R23241 VSS.n5286 VSS.n2197 0.796907
R23242 VSS.n4052 VSS 0.78605
R23243 VSS.n5240 DVSS 0.783069
R23244 VSS.n5241 DVSS 0.783069
R23245 VSS.n3055 VSS.n3054 0.778288
R23246 VSS.n3775 VSS.n2103 0.774059
R23247 VSS.n2173 VSS.n2172 0.752663
R23248 VSS.n4061 VSS 0.751638
R23249 VSS.n3070 VSS.n2971 0.7505
R23250 VSS.n3313 VSS.n3312 0.7505
R23251 DVSS VSS.n3381 0.746344
R23252 VSS.n282 VSS.n122 0.745113
R23253 VSS.n824 VSS.n305 0.745113
R23254 VSS.n751 VSS.n330 0.745113
R23255 VSS.n2975 VSS.n2974 0.743357
R23256 VSS.n2974 VSS.n2966 0.743357
R23257 VSS.n3256 VSS.n2965 0.743357
R23258 VSS.n2968 VSS.n2965 0.743357
R23259 VSS.n3074 VSS.n3073 0.743357
R23260 VSS.n3073 VSS.n2968 0.743357
R23261 VSS.n3011 VSS.n2964 0.743357
R23262 VSS.n2966 VSS.n2964 0.743357
R23263 VSS.n283 VSS.n282 0.736857
R23264 VSS.n825 VSS.n824 0.736857
R23265 VSS.n751 VSS.n750 0.736857
R23266 VSS.n3059 VSS.n3058 0.735937
R23267 VSS.n3310 VSS.n3309 0.735937
R23268 VSS.n5431 VSS.n2084 0.7304
R23269 VSS.n4103 VSS.n4102 0.71546
R23270 VSS.n4107 VSS.n4106 0.71546
R23271 VSS.n5245 VSS.n5237 0.71546
R23272 VSS.n2801 VSS.n2800 0.707265
R23273 VSS.n5321 VSS.n2182 0.693432
R23274 VSS.n2180 VSS.n2179 0.693432
R23275 VSS.n2097 VSS.n2096 0.693432
R23276 VSS.n2094 VSS.n2093 0.693432
R23277 VSS.n5416 VSS.n2096 0.682241
R23278 VSS.n5322 VSS.n5321 0.682241
R23279 VSS.n5324 VSS.n2180 0.682241
R23280 VSS.n5418 VSS.n2094 0.682241
R23281 VSS.n3530 VSS.n3529 0.666308
R23282 VSS.n5283 VSS.n5282 0.66242
R23283 VSS.n5429 VSS.n5428 0.662265
R23284 VSS.n5336 VSS.n5335 0.662265
R23285 VSS.n5391 VSS.n2108 0.662265
R23286 VSS.n3529 VSS.n2887 0.64762
R23287 VSS.n5241 VSS.n5240 0.646382
R23288 VSS.n1773 VSS.n1769 0.643357
R23289 VSS.n1879 VSS.n1878 0.643357
R23290 VSS.n1876 VSS.n1875 0.643357
R23291 VSS.n1775 VSS.n1774 0.643357
R23292 VSS.n1917 VSS.n1916 0.643357
R23293 VSS.n1915 VSS.n1914 0.643357
R23294 VSS.n1899 VSS.n1747 0.643357
R23295 VSS.n1902 VSS.n1901 0.643357
R23296 VSS.n1955 VSS.n1954 0.643357
R23297 VSS.n1953 VSS.n1952 0.643357
R23298 VSS.n1937 VSS.n1705 0.643357
R23299 VSS.n1940 VSS.n1939 0.643357
R23300 VSS.n1677 VSS.n1676 0.643357
R23301 VSS.n1739 VSS.n1738 0.643357
R23302 VSS.n1687 VSS.n1685 0.643357
R23303 VSS.n1976 VSS.n1975 0.643357
R23304 VSS.n1650 VSS.n1649 0.643357
R23305 VSS.n1733 VSS.n1732 0.643357
R23306 VSS.n1662 VSS.n1660 0.643357
R23307 VSS.n2008 VSS.n2007 0.643357
R23308 VSS.n1629 VSS.n1625 0.643357
R23309 VSS.n2044 VSS.n2043 0.643357
R23310 VSS.n2041 VSS.n2040 0.643357
R23311 VSS.n1631 VSS.n1630 0.643357
R23312 VSS.n3418 VSS.n3417 0.634889
R23313 VSS.n2101 DVSS 0.621687
R23314 VSS.n5406 DVSS 0.621687
R23315 VSS.n5311 DVSS 0.621687
R23316 VSS.n5310 DVSS 0.621687
R23317 VSS.n5242 VSS.n5241 0.618588
R23318 VSS.n5282 DVSS 0.600908
R23319 VSS.n5258 VSS.n2231 0.588678
R23320 VSS.n4068 VSS.n4059 0.585632
R23321 VSS.n4072 VSS.n2460 0.585632
R23322 VSS.n2455 VSS.n2448 0.585632
R23323 VSS.n4146 VSS.n4145 0.584525
R23324 VSS.n5247 VSS.n2242 0.584525
R23325 VSS.n4241 VSS.n2372 0.584525
R23326 VSS.n4086 VSS.n2355 0.584525
R23327 VSS.n5120 VSS.n5119 0.578278
R23328 DVSS VSS.n5130 0.578278
R23329 VSS.n5130 VSS.n5129 0.578278
R23330 VSS.n5258 VSS.n5257 0.578278
R23331 VSS.n5259 VSS.n2210 0.578278
R23332 VSS.n5260 VSS.n2208 0.578278
R23333 VSS.n5261 VSS.n2211 0.578278
R23334 VSS.n5262 VSS.n2207 0.578278
R23335 VSS.n5263 VSS.n2212 0.578278
R23336 VSS.n5264 VSS.n2206 0.578278
R23337 VSS.n5265 VSS.n2213 0.578278
R23338 VSS.n5266 VSS.n2205 0.578278
R23339 VSS.n5267 VSS.n2214 0.578278
R23340 VSS.n5272 VSS.n5271 0.578278
R23341 VSS.n5274 VSS.n5273 0.578278
R23342 VSS.n5284 VSS.n2197 0.578278
R23343 VSS.n2197 VSS.n2195 0.578278
R23344 VSS.n5287 VSS.n5286 0.578278
R23345 VSS.n2196 VSS.n2194 0.578278
R23346 VSS.n3523 VSS.n3522 0.578278
R23347 VSS.n3387 VSS.n3386 0.578278
R23348 VSS.n3518 VSS.n3517 0.578278
R23349 VSS.n3516 VSS.n3389 0.578278
R23350 VSS.n3515 VSS.n3514 0.578278
R23351 VSS.n3508 VSS.n3391 0.578278
R23352 VSS.n3510 VSS.n3509 0.578278
R23353 VSS.n5286 VSS.n5285 0.578278
R23354 VSS.n2198 VSS.n2196 0.578278
R23355 VSS.n3522 VSS.n3521 0.578278
R23356 VSS.n3520 VSS.n3387 0.578278
R23357 VSS.n3519 VSS.n3518 0.578278
R23358 VSS.n3389 VSS.n3388 0.578278
R23359 VSS.n3514 VSS.n3513 0.578278
R23360 VSS.n3512 VSS.n3391 0.578278
R23361 VSS.n3511 VSS.n3510 0.578278
R23362 VSS.n4069 VSS.n4068 0.563
R23363 VSS.n5297 VSS.n2189 0.557079
R23364 VSS.n4079 VSS.n4078 0.557079
R23365 VSS.n5408 VSS.n5407 0.557079
R23366 VSS.n5313 VSS.n5312 0.557079
R23367 VSS.n4091 VSS.n4090 0.557079
R23368 VSS.n5302 VSS.n5300 0.553108
R23369 VSS.n5295 VSS.n2192 0.553108
R23370 VSS.n4049 VSS.n4046 0.553108
R23371 VSS.n4084 VSS.n4083 0.549281
R23372 VSS.n2365 VSS.n2363 0.545794
R23373 VSS.n5425 VSS.n5424 0.545794
R23374 VSS.n5430 VSS.n5429 0.545794
R23375 VSS.n5338 VSS.n5337 0.545794
R23376 VSS.n5337 VSS.n5336 0.545794
R23377 VSS.n5398 VSS.n2108 0.545794
R23378 VSS.n5399 VSS.n5398 0.545794
R23379 VSS.n2798 VSS.n2107 0.545794
R23380 VSS.n4145 VSS.n4144 0.545794
R23381 VSS.n5248 VSS.n5247 0.545794
R23382 VSS.n4246 VSS.n2355 0.545794
R23383 VSS.n4242 VSS.n4241 0.545794
R23384 VSS.n5425 DVSS 0.544093
R23385 VSS.n5423 DVSS 0.544093
R23386 VSS.n5424 DVSS 0.544018
R23387 VSS.n4290 VSS.n4287 0.543147
R23388 VSS.n5309 VSS.n5308 0.533549
R23389 VSS.n3059 VSS.n2975 0.5255
R23390 VSS.n3310 VSS.n3074 0.5255
R23391 VSS.n2451 VSS.n2448 0.5205
R23392 VSS.n2460 VSS.n2459 0.5205
R23393 VSS.n4063 VSS.n4059 0.5205
R23394 VSS.n3505 VSS.n3394 0.519124
R23395 VSS.n3397 VSS.n3396 0.519124
R23396 VSS.n5298 VSS.n2188 0.519124
R23397 VSS.n5296 VSS.n2190 0.519124
R23398 VSS.n4048 VSS.n4047 0.519124
R23399 VSS.n4312 VSS.n4307 0.5005
R23400 VSS.n5105 VSS.n4313 0.5005
R23401 VSS.n5104 VSS.n4314 0.5005
R23402 VSS.n4328 VSS.n4315 0.5005
R23403 VSS.n4329 VSS.n4327 0.5005
R23404 VSS.n5093 VSS.n4330 0.5005
R23405 VSS.n5092 VSS.n4331 0.5005
R23406 VSS.n4345 VSS.n4332 0.5005
R23407 VSS.n4346 VSS.n4344 0.5005
R23408 VSS.n5081 VSS.n4347 0.5005
R23409 VSS.n5080 VSS.n4348 0.5005
R23410 VSS.n4686 VSS.n4349 0.5005
R23411 VSS.n4689 VSS.n4688 0.5005
R23412 VSS.n4687 VSS.n4364 0.5005
R23413 VSS.n5065 VSS.n4365 0.5005
R23414 VSS.n5064 VSS.n4366 0.5005
R23415 VSS.n4380 VSS.n4367 0.5005
R23416 VSS.n4381 VSS.n4379 0.5005
R23417 VSS.n5053 VSS.n4382 0.5005
R23418 VSS.n5052 VSS.n4383 0.5005
R23419 VSS.n4399 VSS.n4384 0.5005
R23420 VSS.n4400 VSS.n4398 0.5005
R23421 VSS.n5041 VSS.n4401 0.5005
R23422 VSS.n5040 VSS.n4402 0.5005
R23423 VSS.n4416 VSS.n4403 0.5005
R23424 VSS.n4417 VSS.n4415 0.5005
R23425 VSS.n5029 VSS.n4418 0.5005
R23426 VSS.n5028 VSS.n4419 0.5005
R23427 VSS.n4434 VSS.n4420 0.5005
R23428 VSS.n4435 VSS.n4433 0.5005
R23429 VSS.n5017 VSS.n4436 0.5005
R23430 VSS.n5016 VSS.n4437 0.5005
R23431 VSS.n4753 VSS.n4438 0.5005
R23432 VSS.n4756 VSS.n4755 0.5005
R23433 VSS.n4754 VSS.n4454 0.5005
R23434 VSS.n5001 VSS.n4455 0.5005
R23435 VSS.n5000 VSS.n4456 0.5005
R23436 VSS.n4470 VSS.n4457 0.5005
R23437 VSS.n4471 VSS.n4469 0.5005
R23438 VSS.n4989 VSS.n4472 0.5005
R23439 VSS.n4988 VSS.n4473 0.5005
R23440 VSS.n4489 VSS.n4474 0.5005
R23441 VSS.n4490 VSS.n4488 0.5005
R23442 VSS.n4977 VSS.n4491 0.5005
R23443 VSS.n4976 VSS.n4492 0.5005
R23444 VSS.n4507 VSS.n4493 0.5005
R23445 VSS.n4508 VSS.n4506 0.5005
R23446 VSS.n4965 VSS.n4509 0.5005
R23447 VSS.n4964 VSS.n4510 0.5005
R23448 VSS.n4525 VSS.n4511 0.5005
R23449 VSS.n4526 VSS.n4524 0.5005
R23450 VSS.n4953 VSS.n4527 0.5005
R23451 VSS.n4952 VSS.n4528 0.5005
R23452 VSS.n4543 VSS.n4529 0.5005
R23453 VSS.n4544 VSS.n4542 0.5005
R23454 VSS.n4940 VSS.n4545 0.5005
R23455 VSS.n4939 VSS.n4546 0.5005
R23456 VSS.n4560 VSS.n4547 0.5005
R23457 VSS.n4561 VSS.n4559 0.5005
R23458 VSS.n4928 VSS.n4562 0.5005
R23459 VSS.n4927 VSS.n4563 0.5005
R23460 VSS.n4578 VSS.n4564 0.5005
R23461 VSS.n4579 VSS.n4577 0.5005
R23462 VSS.n4915 VSS.n4580 0.5005
R23463 VSS.n4914 VSS.n4581 0.5005
R23464 VSS.n4595 VSS.n4582 0.5005
R23465 VSS.n4596 VSS.n4594 0.5005
R23466 VSS.n4902 VSS.n4597 0.5005
R23467 VSS.n4901 VSS.n4598 0.5005
R23468 VSS.n4613 VSS.n4599 0.5005
R23469 VSS.n4614 VSS.n4612 0.5005
R23470 VSS.n4890 VSS.n4615 0.5005
R23471 VSS.n4889 VSS.n4616 0.5005
R23472 VSS.n4618 VSS.n4617 0.5005
R23473 VSS.n2279 VSS.n2278 0.5005
R23474 VSS.n5136 VSS.n5135 0.5005
R23475 VSS.n5137 VSS.n2277 0.5005
R23476 VSS.n5139 VSS.n5138 0.5005
R23477 VSS.n2275 VSS.n2274 0.5005
R23478 VSS.n5144 VSS.n5143 0.5005
R23479 VSS.n5145 VSS.n2273 0.5005
R23480 VSS.n5167 VSS.n5146 0.5005
R23481 VSS.n5166 VSS.n5147 0.5005
R23482 VSS.n5165 VSS.n5148 0.5005
R23483 VSS.n5151 VSS.n5149 0.5005
R23484 VSS.n5161 VSS.n5152 0.5005
R23485 VSS.n5160 VSS.n5153 0.5005
R23486 VSS.n5159 VSS.n5154 0.5005
R23487 VSS.n5156 VSS.n5155 0.5005
R23488 VSS.n4311 VSS.n4310 0.5005
R23489 VSS.n5168 VSS.n5167 0.5005
R23490 VSS.n5166 VSS.n2272 0.5005
R23491 VSS.n5165 VSS.n5164 0.5005
R23492 VSS.n5163 VSS.n5149 0.5005
R23493 VSS.n5162 VSS.n5161 0.5005
R23494 VSS.n5160 VSS.n5150 0.5005
R23495 VSS.n5159 VSS.n5158 0.5005
R23496 VSS.n2273 VSS.n2271 0.5005
R23497 VSS.n5143 VSS.n5142 0.5005
R23498 VSS.n5141 VSS.n2275 0.5005
R23499 VSS.n5140 VSS.n5139 0.5005
R23500 VSS.n2277 VSS.n2276 0.5005
R23501 VSS.n5135 VSS.n5134 0.5005
R23502 VSS.n4877 VSS.n2279 0.5005
R23503 VSS.n4620 VSS.n4618 0.5005
R23504 VSS.n4889 VSS.n4888 0.5005
R23505 VSS.n4891 VSS.n4890 0.5005
R23506 VSS.n4612 VSS.n4609 0.5005
R23507 VSS.n4601 VSS.n4599 0.5005
R23508 VSS.n4901 VSS.n4900 0.5005
R23509 VSS.n4903 VSS.n4902 0.5005
R23510 VSS.n4594 VSS.n4591 0.5005
R23511 VSS.n4584 VSS.n4582 0.5005
R23512 VSS.n4914 VSS.n4913 0.5005
R23513 VSS.n4916 VSS.n4915 0.5005
R23514 VSS.n4577 VSS.n4574 0.5005
R23515 VSS.n4566 VSS.n4564 0.5005
R23516 VSS.n4927 VSS.n4926 0.5005
R23517 VSS.n4929 VSS.n4928 0.5005
R23518 VSS.n4559 VSS.n4556 0.5005
R23519 VSS.n4549 VSS.n4547 0.5005
R23520 VSS.n4939 VSS.n4938 0.5005
R23521 VSS.n4941 VSS.n4940 0.5005
R23522 VSS.n4542 VSS.n4539 0.5005
R23523 VSS.n4531 VSS.n4529 0.5005
R23524 VSS.n4952 VSS.n4951 0.5005
R23525 VSS.n4954 VSS.n4953 0.5005
R23526 VSS.n4524 VSS.n4521 0.5005
R23527 VSS.n4513 VSS.n4511 0.5005
R23528 VSS.n4964 VSS.n4963 0.5005
R23529 VSS.n4966 VSS.n4965 0.5005
R23530 VSS.n4506 VSS.n4503 0.5005
R23531 VSS.n4495 VSS.n4493 0.5005
R23532 VSS.n4976 VSS.n4975 0.5005
R23533 VSS.n4978 VSS.n4977 0.5005
R23534 VSS.n4488 VSS.n4485 0.5005
R23535 VSS.n4476 VSS.n4474 0.5005
R23536 VSS.n4988 VSS.n4987 0.5005
R23537 VSS.n4990 VSS.n4989 0.5005
R23538 VSS.n4469 VSS.n4466 0.5005
R23539 VSS.n4459 VSS.n4457 0.5005
R23540 VSS.n5000 VSS.n4999 0.5005
R23541 VSS.n5002 VSS.n5001 0.5005
R23542 VSS.n4454 VSS.n4451 0.5005
R23543 VSS.n4757 VSS.n4756 0.5005
R23544 VSS.n4440 VSS.n4438 0.5005
R23545 VSS.n5016 VSS.n5015 0.5005
R23546 VSS.n5018 VSS.n5017 0.5005
R23547 VSS.n4433 VSS.n4430 0.5005
R23548 VSS.n4422 VSS.n4420 0.5005
R23549 VSS.n5028 VSS.n5027 0.5005
R23550 VSS.n5030 VSS.n5029 0.5005
R23551 VSS.n4415 VSS.n4412 0.5005
R23552 VSS.n4405 VSS.n4403 0.5005
R23553 VSS.n5040 VSS.n5039 0.5005
R23554 VSS.n5042 VSS.n5041 0.5005
R23555 VSS.n4398 VSS.n4395 0.5005
R23556 VSS.n4386 VSS.n4384 0.5005
R23557 VSS.n5052 VSS.n5051 0.5005
R23558 VSS.n5054 VSS.n5053 0.5005
R23559 VSS.n4379 VSS.n4376 0.5005
R23560 VSS.n4369 VSS.n4367 0.5005
R23561 VSS.n5064 VSS.n5063 0.5005
R23562 VSS.n5066 VSS.n5065 0.5005
R23563 VSS.n4364 VSS.n4361 0.5005
R23564 VSS.n4690 VSS.n4689 0.5005
R23565 VSS.n4351 VSS.n4349 0.5005
R23566 VSS.n5080 VSS.n5079 0.5005
R23567 VSS.n5082 VSS.n5081 0.5005
R23568 VSS.n4344 VSS.n4341 0.5005
R23569 VSS.n4334 VSS.n4332 0.5005
R23570 VSS.n5092 VSS.n5091 0.5005
R23571 VSS.n5094 VSS.n5093 0.5005
R23572 VSS.n4327 VSS.n4324 0.5005
R23573 VSS.n4317 VSS.n4315 0.5005
R23574 VSS.n5104 VSS.n5103 0.5005
R23575 VSS.n5106 VSS.n5105 0.5005
R23576 VSS.n4307 VSS.n4304 0.5005
R23577 VSS.n4309 VSS.n4296 0.5005
R23578 VSS.n4310 VSS.n4297 0.5005
R23579 VSS VSS.n4060 0.497977
R23580 VSS VSS.n2446 0.497977
R23581 VSS VSS.n2447 0.497977
R23582 VSS VSS.n2449 0.497977
R23583 VSS.n4142 VSS.n2432 0.497868
R23584 VSS.n4244 VSS.n2358 0.497868
R23585 VSS.n3402 VSS.n3401 0.495738
R23586 VSS.n1079 VSS.n1078 0.490418
R23587 VSS.n2788 VSS.n2787 0.478861
R23588 VSS.n5252 VSS.n2227 0.477527
R23589 VSS.n5253 VSS.n5252 0.473227
R23590 VSS.n2450 VSS.n2292 0.473227
R23591 VSS.n4078 VSS.n4077 0.473227
R23592 VSS.n4077 VSS.n4076 0.473227
R23593 VSS.n4062 VSS.n4061 0.473227
R23594 VSS.n4064 VSS.n4062 0.473227
R23595 VSS.n2791 VSS.n2790 0.473227
R23596 VSS.n5424 DVSS 0.469029
R23597 VSS.n5119 DVSS 0.467804
R23598 VSS.n5119 DVSS 0.467804
R23599 VSS.n2799 VSS.n2798 0.465755
R23600 VSS.n2786 VSS.n2784 0.457714
R23601 VSS.n2314 VSS.n2313 0.455549
R23602 VSS.n2689 VSS.n2686 0.455549
R23603 VSS.n1829 VSS.n1828 0.455549
R23604 VSS.n3439 VSS.n3438 0.455549
R23605 VSS.n5702 VSS.n4 0.455549
R23606 VSS.n3503 VSS.n3502 0.452884
R23607 VSS.n4053 VSS.n4052 0.452868
R23608 VSS.n3503 VSS.n3419 0.452744
R23609 VSS.n2693 VSS.n2692 0.4505
R23610 VSS.n2694 VSS.n2477 0.4505
R23611 VSS.n2696 VSS.n2695 0.4505
R23612 VSS.n2685 VSS.n2684 0.4505
R23613 VSS.n2683 VSS.n2478 0.4505
R23614 VSS.n2682 VSS.n2480 0.4505
R23615 VSS.n2676 VSS.n2479 0.4505
R23616 VSS.n2678 VSS.n2677 0.4505
R23617 VSS.n2675 VSS.n2482 0.4505
R23618 VSS.n2674 VSS.n2673 0.4505
R23619 VSS.n2484 VSS.n2483 0.4505
R23620 VSS.n2669 VSS.n2668 0.4505
R23621 VSS.n2667 VSS.n2486 0.4505
R23622 VSS.n2666 VSS.n2665 0.4505
R23623 VSS.n2488 VSS.n2487 0.4505
R23624 VSS.n2661 VSS.n2660 0.4505
R23625 VSS.n2659 VSS.n2490 0.4505
R23626 VSS.n2658 VSS.n2657 0.4505
R23627 VSS.n2492 VSS.n2491 0.4505
R23628 VSS.n2653 VSS.n2652 0.4505
R23629 VSS.n2651 VSS.n2494 0.4505
R23630 VSS.n2650 VSS.n2649 0.4505
R23631 VSS.n2496 VSS.n2495 0.4505
R23632 VSS.n2645 VSS.n2644 0.4505
R23633 VSS.n2643 VSS.n2498 0.4505
R23634 VSS.n2642 VSS.n2641 0.4505
R23635 VSS.n2500 VSS.n2499 0.4505
R23636 VSS.n2637 VSS.n2636 0.4505
R23637 VSS.n2635 VSS.n2502 0.4505
R23638 VSS.n2634 VSS.n2633 0.4505
R23639 VSS.n2504 VSS.n2503 0.4505
R23640 VSS.n2629 VSS.n2628 0.4505
R23641 VSS.n2627 VSS.n2506 0.4505
R23642 VSS.n2626 VSS.n2625 0.4505
R23643 VSS.n2508 VSS.n2507 0.4505
R23644 VSS.n2621 VSS.n2620 0.4505
R23645 VSS.n2619 VSS.n2510 0.4505
R23646 VSS.n2618 VSS.n2617 0.4505
R23647 VSS.n2512 VSS.n2511 0.4505
R23648 VSS.n2613 VSS.n2612 0.4505
R23649 VSS.n2611 VSS.n2514 0.4505
R23650 VSS.n2610 VSS.n2609 0.4505
R23651 VSS.n2516 VSS.n2515 0.4505
R23652 VSS.n2605 VSS.n2604 0.4505
R23653 VSS.n2603 VSS.n2518 0.4505
R23654 VSS.n2602 VSS.n2601 0.4505
R23655 VSS.n2520 VSS.n2519 0.4505
R23656 VSS.n2597 VSS.n2596 0.4505
R23657 VSS.n2595 VSS.n2522 0.4505
R23658 VSS.n2594 VSS.n2593 0.4505
R23659 VSS.n2524 VSS.n2523 0.4505
R23660 VSS.n2589 VSS.n2588 0.4505
R23661 VSS.n2587 VSS.n2526 0.4505
R23662 VSS.n2586 VSS.n2585 0.4505
R23663 VSS.n2528 VSS.n2527 0.4505
R23664 VSS.n2581 VSS.n2580 0.4505
R23665 VSS.n2579 VSS.n2530 0.4505
R23666 VSS.n2578 VSS.n2577 0.4505
R23667 VSS.n2532 VSS.n2531 0.4505
R23668 VSS.n2573 VSS.n2572 0.4505
R23669 VSS.n2571 VSS.n2534 0.4505
R23670 VSS.n2570 VSS.n2569 0.4505
R23671 VSS.n2536 VSS.n2535 0.4505
R23672 VSS.n2565 VSS.n2564 0.4505
R23673 VSS.n2563 VSS.n2538 0.4505
R23674 VSS.n2562 VSS.n2561 0.4505
R23675 VSS.n2540 VSS.n2539 0.4505
R23676 VSS.n2557 VSS.n2556 0.4505
R23677 VSS.n2555 VSS.n2542 0.4505
R23678 VSS.n2554 VSS.n2553 0.4505
R23679 VSS.n2544 VSS.n2543 0.4505
R23680 VSS.n2549 VSS.n2548 0.4505
R23681 VSS.n2547 VSS.n2546 0.4505
R23682 VSS.n2310 VSS.n2309 0.4505
R23683 VSS.n2320 VSS.n2319 0.4505
R23684 VSS.n2321 VSS.n2308 0.4505
R23685 VSS.n2323 VSS.n2322 0.4505
R23686 VSS.n2306 VSS.n2305 0.4505
R23687 VSS.n2328 VSS.n2327 0.4505
R23688 VSS.n2329 VSS.n2304 0.4505
R23689 VSS.n2331 VSS.n2330 0.4505
R23690 VSS.n2302 VSS.n2301 0.4505
R23691 VSS.n2336 VSS.n2335 0.4505
R23692 VSS.n2337 VSS.n2299 0.4505
R23693 VSS.n4280 VSS.n4279 0.4505
R23694 VSS.n4278 VSS.n2300 0.4505
R23695 VSS.n4277 VSS.n4276 0.4505
R23696 VSS.n2339 VSS.n2338 0.4505
R23697 VSS.n4272 VSS.n4271 0.4505
R23698 VSS.n4270 VSS.n2341 0.4505
R23699 VSS.n4269 VSS.n4268 0.4505
R23700 VSS.n2343 VSS.n2342 0.4505
R23701 VSS.n4264 VSS.n4263 0.4505
R23702 VSS.n4262 VSS.n2345 0.4505
R23703 VSS.n4261 VSS.n4260 0.4505
R23704 VSS.n2347 VSS.n2346 0.4505
R23705 VSS.n4256 VSS.n4255 0.4505
R23706 VSS.n4254 VSS.n2349 0.4505
R23707 VSS.n4253 VSS.n4252 0.4505
R23708 VSS.n2351 VSS.n2350 0.4505
R23709 VSS.n2368 VSS.n2365 0.4505
R23710 VSS.n2902 VSS.n2901 0.4505
R23711 VSS.n2989 VSS.n2988 0.4505
R23712 VSS.n2991 VSS.n2990 0.4505
R23713 VSS.n2982 VSS.n2981 0.4505
R23714 VSS.n2998 VSS.n2997 0.4505
R23715 VSS.n2999 VSS.n2980 0.4505
R23716 VSS.n3001 VSS.n3000 0.4505
R23717 VSS.n2927 VSS.n2925 0.4505
R23718 VSS.n3348 VSS.n3347 0.4505
R23719 VSS.n3346 VSS.n2926 0.4505
R23720 VSS.n3345 VSS.n3344 0.4505
R23721 VSS.n2929 VSS.n2928 0.4505
R23722 VSS.n3063 VSS.n3062 0.4505
R23723 VSS.n2954 VSS.n2952 0.4505
R23724 VSS.n3330 VSS.n3329 0.4505
R23725 VSS.n3328 VSS.n2953 0.4505
R23726 VSS.n3327 VSS.n3326 0.4505
R23727 VSS.n2956 VSS.n2955 0.4505
R23728 VSS.n3106 VSS.n3105 0.4505
R23729 VSS.n3123 VSS.n3122 0.4505
R23730 VSS.n3124 VSS.n3102 0.4505
R23731 VSS.n3127 VSS.n3126 0.4505
R23732 VSS.n3125 VSS.n3104 0.4505
R23733 VSS.n3085 VSS.n3083 0.4505
R23734 VSS.n3301 VSS.n3300 0.4505
R23735 VSS.n3299 VSS.n3084 0.4505
R23736 VSS.n3298 VSS.n3297 0.4505
R23737 VSS.n3087 VSS.n3086 0.4505
R23738 VSS.n3150 VSS.n3148 0.4505
R23739 VSS.n3285 VSS.n3284 0.4505
R23740 VSS.n3283 VSS.n3149 0.4505
R23741 VSS.n3282 VSS.n3281 0.4505
R23742 VSS.n3152 VSS.n3151 0.4505
R23743 VSS.n3243 VSS.n3242 0.4505
R23744 VSS.n3241 VSS.n3156 0.4505
R23745 VSS.n3240 VSS.n3239 0.4505
R23746 VSS.n3158 VSS.n3157 0.4505
R23747 VSS.n3235 VSS.n3234 0.4505
R23748 VSS.n3233 VSS.n3160 0.4505
R23749 VSS.n3232 VSS.n3231 0.4505
R23750 VSS.n3162 VSS.n3161 0.4505
R23751 VSS.n3227 VSS.n3226 0.4505
R23752 VSS.n3225 VSS.n3164 0.4505
R23753 VSS.n3224 VSS.n3223 0.4505
R23754 VSS.n3166 VSS.n3165 0.4505
R23755 VSS.n3219 VSS.n3218 0.4505
R23756 VSS.n3217 VSS.n3168 0.4505
R23757 VSS.n3216 VSS.n3215 0.4505
R23758 VSS.n3170 VSS.n3169 0.4505
R23759 VSS.n3211 VSS.n3210 0.4505
R23760 VSS.n3209 VSS.n3172 0.4505
R23761 VSS.n3208 VSS.n3207 0.4505
R23762 VSS.n3174 VSS.n3173 0.4505
R23763 VSS.n3203 VSS.n3202 0.4505
R23764 VSS.n3201 VSS.n3176 0.4505
R23765 VSS.n3200 VSS.n3199 0.4505
R23766 VSS.n3178 VSS.n3177 0.4505
R23767 VSS.n3195 VSS.n3194 0.4505
R23768 VSS.n3193 VSS.n3180 0.4505
R23769 VSS.n3192 VSS.n3191 0.4505
R23770 VSS.n3182 VSS.n3181 0.4505
R23771 VSS.n3187 VSS.n3186 0.4505
R23772 VSS.n3185 VSS.n3184 0.4505
R23773 VSS.n3377 VSS.n3376 0.4505
R23774 VSS.n3375 VSS.n2895 0.4505
R23775 VSS.n3374 VSS.n3373 0.4505
R23776 VSS.n2897 VSS.n2896 0.4505
R23777 VSS.n3369 VSS.n3368 0.4505
R23778 VSS.n3367 VSS.n2900 0.4505
R23779 VSS.n3366 VSS.n3365 0.4505
R23780 VSS.n3581 VSS.n3580 0.4505
R23781 VSS.n3585 VSS.n3584 0.4505
R23782 VSS.n3586 VSS.n3579 0.4505
R23783 VSS.n3588 VSS.n3587 0.4505
R23784 VSS.n3577 VSS.n3576 0.4505
R23785 VSS.n3593 VSS.n3592 0.4505
R23786 VSS.n3594 VSS.n3575 0.4505
R23787 VSS.n3596 VSS.n3595 0.4505
R23788 VSS.n3573 VSS.n3572 0.4505
R23789 VSS.n3601 VSS.n3600 0.4505
R23790 VSS.n3602 VSS.n3571 0.4505
R23791 VSS.n3604 VSS.n3603 0.4505
R23792 VSS.n3569 VSS.n3568 0.4505
R23793 VSS.n3609 VSS.n3608 0.4505
R23794 VSS.n3610 VSS.n3567 0.4505
R23795 VSS.n3612 VSS.n3611 0.4505
R23796 VSS.n3565 VSS.n3564 0.4505
R23797 VSS.n3617 VSS.n3616 0.4505
R23798 VSS.n3618 VSS.n3563 0.4505
R23799 VSS.n3620 VSS.n3619 0.4505
R23800 VSS.n3561 VSS.n3560 0.4505
R23801 VSS.n3625 VSS.n3624 0.4505
R23802 VSS.n3626 VSS.n3559 0.4505
R23803 VSS.n3628 VSS.n3627 0.4505
R23804 VSS.n3557 VSS.n3556 0.4505
R23805 VSS.n3633 VSS.n3632 0.4505
R23806 VSS.n3634 VSS.n3552 0.4505
R23807 VSS.n3725 VSS.n2821 0.4505
R23808 VSS.n2824 VSS.n2820 0.4505
R23809 VSS.n3721 VSS.n3720 0.4505
R23810 VSS.n3719 VSS.n2823 0.4505
R23811 VSS.n3718 VSS.n3717 0.4505
R23812 VSS.n2826 VSS.n2825 0.4505
R23813 VSS.n3711 VSS.n3710 0.4505
R23814 VSS.n3709 VSS.n2841 0.4505
R23815 VSS.n3708 VSS.n3707 0.4505
R23816 VSS.n2843 VSS.n2842 0.4505
R23817 VSS.n3703 VSS.n3702 0.4505
R23818 VSS.n3701 VSS.n2845 0.4505
R23819 VSS.n3700 VSS.n3699 0.4505
R23820 VSS.n2847 VSS.n2846 0.4505
R23821 VSS.n3695 VSS.n3694 0.4505
R23822 VSS.n3693 VSS.n2849 0.4505
R23823 VSS.n3692 VSS.n3691 0.4505
R23824 VSS.n2851 VSS.n2850 0.4505
R23825 VSS.n3687 VSS.n3686 0.4505
R23826 VSS.n3685 VSS.n2853 0.4505
R23827 VSS.n3684 VSS.n3683 0.4505
R23828 VSS.n2855 VSS.n2854 0.4505
R23829 VSS.n3679 VSS.n3678 0.4505
R23830 VSS.n3677 VSS.n2857 0.4505
R23831 VSS.n3676 VSS.n3675 0.4505
R23832 VSS.n2859 VSS.n2858 0.4505
R23833 VSS.n3671 VSS.n3670 0.4505
R23834 VSS.n3669 VSS.n2861 0.4505
R23835 VSS.n3668 VSS.n3667 0.4505
R23836 VSS.n2863 VSS.n2862 0.4505
R23837 VSS.n3663 VSS.n3662 0.4505
R23838 VSS.n3661 VSS.n2865 0.4505
R23839 VSS.n3660 VSS.n3659 0.4505
R23840 VSS.n2867 VSS.n2866 0.4505
R23841 VSS.n3655 VSS.n3654 0.4505
R23842 VSS.n3653 VSS.n2869 0.4505
R23843 VSS.n3652 VSS.n3651 0.4505
R23844 VSS.n2871 VSS.n2870 0.4505
R23845 VSS.n3647 VSS.n3646 0.4505
R23846 VSS.n3645 VSS.n2873 0.4505
R23847 VSS.n3644 VSS.n3643 0.4505
R23848 VSS.n2875 VSS.n2874 0.4505
R23849 VSS.n3554 VSS.n3553 0.4505
R23850 VSS.n3555 VSS.n3551 0.4505
R23851 VSS.n3636 VSS.n3635 0.4505
R23852 VSS.n3552 VSS.n3550 0.4505
R23853 VSS.n3727 VSS.n3726 0.4505
R23854 VSS.n3632 VSS.n3631 0.4505
R23855 VSS.n3630 VSS.n3557 0.4505
R23856 VSS.n3629 VSS.n3628 0.4505
R23857 VSS.n3559 VSS.n3558 0.4505
R23858 VSS.n3624 VSS.n3623 0.4505
R23859 VSS.n3622 VSS.n3561 0.4505
R23860 VSS.n3621 VSS.n3620 0.4505
R23861 VSS.n3563 VSS.n3562 0.4505
R23862 VSS.n3616 VSS.n3615 0.4505
R23863 VSS.n3614 VSS.n3565 0.4505
R23864 VSS.n3613 VSS.n3612 0.4505
R23865 VSS.n3567 VSS.n3566 0.4505
R23866 VSS.n3608 VSS.n3607 0.4505
R23867 VSS.n3606 VSS.n3569 0.4505
R23868 VSS.n3605 VSS.n3604 0.4505
R23869 VSS.n3571 VSS.n3570 0.4505
R23870 VSS.n3600 VSS.n3599 0.4505
R23871 VSS.n3598 VSS.n3573 0.4505
R23872 VSS.n3597 VSS.n3596 0.4505
R23873 VSS.n3575 VSS.n3574 0.4505
R23874 VSS.n3592 VSS.n3591 0.4505
R23875 VSS.n3590 VSS.n3577 0.4505
R23876 VSS.n3589 VSS.n3588 0.4505
R23877 VSS.n3579 VSS.n3578 0.4505
R23878 VSS.n3584 VSS.n3583 0.4505
R23879 VSS.n3725 VSS.n3724 0.4505
R23880 VSS.n3723 VSS.n2820 0.4505
R23881 VSS.n3722 VSS.n3721 0.4505
R23882 VSS.n2823 VSS.n2822 0.4505
R23883 VSS.n3717 VSS.n3716 0.4505
R23884 VSS.n2833 VSS.n2826 0.4505
R23885 VSS.n3712 VSS.n3711 0.4505
R23886 VSS.n2841 VSS.n2840 0.4505
R23887 VSS.n3707 VSS.n3706 0.4505
R23888 VSS.n3705 VSS.n2843 0.4505
R23889 VSS.n3704 VSS.n3703 0.4505
R23890 VSS.n2845 VSS.n2844 0.4505
R23891 VSS.n3699 VSS.n3698 0.4505
R23892 VSS.n3697 VSS.n2847 0.4505
R23893 VSS.n3696 VSS.n3695 0.4505
R23894 VSS.n2849 VSS.n2848 0.4505
R23895 VSS.n3691 VSS.n3690 0.4505
R23896 VSS.n3689 VSS.n2851 0.4505
R23897 VSS.n3688 VSS.n3687 0.4505
R23898 VSS.n2853 VSS.n2852 0.4505
R23899 VSS.n3683 VSS.n3682 0.4505
R23900 VSS.n3681 VSS.n2855 0.4505
R23901 VSS.n3680 VSS.n3679 0.4505
R23902 VSS.n2857 VSS.n2856 0.4505
R23903 VSS.n3675 VSS.n3674 0.4505
R23904 VSS.n3673 VSS.n2859 0.4505
R23905 VSS.n3672 VSS.n3671 0.4505
R23906 VSS.n2861 VSS.n2860 0.4505
R23907 VSS.n3667 VSS.n3666 0.4505
R23908 VSS.n3665 VSS.n2863 0.4505
R23909 VSS.n3664 VSS.n3663 0.4505
R23910 VSS.n2865 VSS.n2864 0.4505
R23911 VSS.n3659 VSS.n3658 0.4505
R23912 VSS.n3657 VSS.n2867 0.4505
R23913 VSS.n3656 VSS.n3655 0.4505
R23914 VSS.n2869 VSS.n2868 0.4505
R23915 VSS.n3651 VSS.n3650 0.4505
R23916 VSS.n3649 VSS.n2871 0.4505
R23917 VSS.n3648 VSS.n3647 0.4505
R23918 VSS.n2873 VSS.n2872 0.4505
R23919 VSS.n3643 VSS.n3642 0.4505
R23920 VSS.n3641 VSS.n2875 0.4505
R23921 VSS.n3553 VSS.n2880 0.4505
R23922 VSS.n3551 VSS.n3549 0.4505
R23923 VSS.n3637 VSS.n3636 0.4505
R23924 VSS.n1836 VSS.n1827 0.4505
R23925 VSS.n1835 VSS.n1834 0.4505
R23926 VSS.n2060 VSS.n2059 0.4505
R23927 VSS.n2058 VSS.n1614 0.4505
R23928 VSS.n2057 VSS.n2056 0.4505
R23929 VSS.n1616 VSS.n1615 0.4505
R23930 VSS.n2052 VSS.n2051 0.4505
R23931 VSS.n2050 VSS.n1619 0.4505
R23932 VSS.n2049 VSS.n2048 0.4505
R23933 VSS.n1621 VSS.n1620 0.4505
R23934 VSS.n1637 VSS.n1635 0.4505
R23935 VSS.n2036 VSS.n2035 0.4505
R23936 VSS.n2034 VSS.n1636 0.4505
R23937 VSS.n2033 VSS.n2032 0.4505
R23938 VSS.n1639 VSS.n1638 0.4505
R23939 VSS.n2028 VSS.n2027 0.4505
R23940 VSS.n2026 VSS.n1645 0.4505
R23941 VSS.n2025 VSS.n2024 0.4505
R23942 VSS.n1647 VSS.n1646 0.4505
R23943 VSS.n1654 VSS.n1652 0.4505
R23944 VSS.n2016 VSS.n2015 0.4505
R23945 VSS.n2014 VSS.n1653 0.4505
R23946 VSS.n2013 VSS.n2012 0.4505
R23947 VSS.n1656 VSS.n1655 0.4505
R23948 VSS.n1668 VSS.n1666 0.4505
R23949 VSS.n2003 VSS.n2002 0.4505
R23950 VSS.n2001 VSS.n1667 0.4505
R23951 VSS.n2000 VSS.n1999 0.4505
R23952 VSS.n1670 VSS.n1669 0.4505
R23953 VSS.n1995 VSS.n1994 0.4505
R23954 VSS.n1993 VSS.n1672 0.4505
R23955 VSS.n1992 VSS.n1991 0.4505
R23956 VSS.n1674 VSS.n1673 0.4505
R23957 VSS.n1984 VSS.n1983 0.4505
R23958 VSS.n1982 VSS.n1679 0.4505
R23959 VSS.n1981 VSS.n1980 0.4505
R23960 VSS.n1681 VSS.n1680 0.4505
R23961 VSS.n1693 VSS.n1691 0.4505
R23962 VSS.n1971 VSS.n1970 0.4505
R23963 VSS.n1969 VSS.n1692 0.4505
R23964 VSS.n1968 VSS.n1967 0.4505
R23965 VSS.n1695 VSS.n1694 0.4505
R23966 VSS.n1963 VSS.n1962 0.4505
R23967 VSS.n1961 VSS.n1697 0.4505
R23968 VSS.n1960 VSS.n1959 0.4505
R23969 VSS.n1699 VSS.n1698 0.4505
R23970 VSS.n1711 VSS.n1709 0.4505
R23971 VSS.n1948 VSS.n1947 0.4505
R23972 VSS.n1946 VSS.n1710 0.4505
R23973 VSS.n1945 VSS.n1944 0.4505
R23974 VSS.n1713 VSS.n1712 0.4505
R23975 VSS.n1933 VSS.n1932 0.4505
R23976 VSS.n1931 VSS.n1717 0.4505
R23977 VSS.n1930 VSS.n1929 0.4505
R23978 VSS.n1719 VSS.n1718 0.4505
R23979 VSS.n1925 VSS.n1924 0.4505
R23980 VSS.n1923 VSS.n1721 0.4505
R23981 VSS.n1922 VSS.n1921 0.4505
R23982 VSS.n1723 VSS.n1722 0.4505
R23983 VSS.n1753 VSS.n1751 0.4505
R23984 VSS.n1910 VSS.n1909 0.4505
R23985 VSS.n1908 VSS.n1752 0.4505
R23986 VSS.n1907 VSS.n1906 0.4505
R23987 VSS.n1755 VSS.n1754 0.4505
R23988 VSS.n1895 VSS.n1894 0.4505
R23989 VSS.n1893 VSS.n1759 0.4505
R23990 VSS.n1892 VSS.n1891 0.4505
R23991 VSS.n1761 VSS.n1760 0.4505
R23992 VSS.n1887 VSS.n1886 0.4505
R23993 VSS.n1885 VSS.n1763 0.4505
R23994 VSS.n1884 VSS.n1883 0.4505
R23995 VSS.n1765 VSS.n1764 0.4505
R23996 VSS.n1781 VSS.n1779 0.4505
R23997 VSS.n1871 VSS.n1870 0.4505
R23998 VSS.n1869 VSS.n1780 0.4505
R23999 VSS.n1868 VSS.n1867 0.4505
R24000 VSS.n1783 VSS.n1782 0.4505
R24001 VSS.n1863 VSS.n1862 0.4505
R24002 VSS.n1861 VSS.n1789 0.4505
R24003 VSS.n1860 VSS.n1859 0.4505
R24004 VSS.n1791 VSS.n1790 0.4505
R24005 VSS.n1852 VSS.n1851 0.4505
R24006 VSS.n1850 VSS.n1822 0.4505
R24007 VSS.n1849 VSS.n1848 0.4505
R24008 VSS.n1824 VSS.n1823 0.4505
R24009 VSS.n1844 VSS.n1843 0.4505
R24010 VSS.n1842 VSS.n1826 0.4505
R24011 VSS.n1841 VSS.n1840 0.4505
R24012 VSS.n1839 VSS.n1837 0.4505
R24013 VSS.n1832 VSS.n1830 0.4505
R24014 VSS.n1834 VSS.n1833 0.4505
R24015 VSS.n1831 VSS.n1827 0.4505
R24016 VSS.n1613 VSS.n1603 0.4505
R24017 VSS.n2061 VSS.n2060 0.4505
R24018 VSS.n1617 VSS.n1614 0.4505
R24019 VSS.n2056 VSS.n2055 0.4505
R24020 VSS.n2054 VSS.n1616 0.4505
R24021 VSS.n2053 VSS.n2052 0.4505
R24022 VSS.n1622 VSS.n1619 0.4505
R24023 VSS.n2048 VSS.n2047 0.4505
R24024 VSS.n1624 VSS.n1621 0.4505
R24025 VSS.n1635 VSS.n1633 0.4505
R24026 VSS.n2037 VSS.n2036 0.4505
R24027 VSS.n1640 VSS.n1636 0.4505
R24028 VSS.n2032 VSS.n2031 0.4505
R24029 VSS.n2030 VSS.n1639 0.4505
R24030 VSS.n2029 VSS.n2028 0.4505
R24031 VSS.n1645 VSS.n1644 0.4505
R24032 VSS.n2024 VSS.n2023 0.4505
R24033 VSS.n2022 VSS.n1647 0.4505
R24034 VSS.n1652 VSS.n1648 0.4505
R24035 VSS.n2017 VSS.n2016 0.4505
R24036 VSS.n1657 VSS.n1653 0.4505
R24037 VSS.n2012 VSS.n2011 0.4505
R24038 VSS.n1659 VSS.n1656 0.4505
R24039 VSS.n1666 VSS.n1664 0.4505
R24040 VSS.n2004 VSS.n2003 0.4505
R24041 VSS.n1667 VSS.n1665 0.4505
R24042 VSS.n1999 VSS.n1998 0.4505
R24043 VSS.n1997 VSS.n1670 0.4505
R24044 VSS.n1996 VSS.n1995 0.4505
R24045 VSS.n1672 VSS.n1671 0.4505
R24046 VSS.n1991 VSS.n1990 0.4505
R24047 VSS.n1675 VSS.n1674 0.4505
R24048 VSS.n1985 VSS.n1984 0.4505
R24049 VSS.n1682 VSS.n1679 0.4505
R24050 VSS.n1980 VSS.n1979 0.4505
R24051 VSS.n1684 VSS.n1681 0.4505
R24052 VSS.n1691 VSS.n1689 0.4505
R24053 VSS.n1972 VSS.n1971 0.4505
R24054 VSS.n1692 VSS.n1690 0.4505
R24055 VSS.n1967 VSS.n1966 0.4505
R24056 VSS.n1965 VSS.n1695 0.4505
R24057 VSS.n1964 VSS.n1963 0.4505
R24058 VSS.n1697 VSS.n1696 0.4505
R24059 VSS.n1959 VSS.n1958 0.4505
R24060 VSS.n1701 VSS.n1699 0.4505
R24061 VSS.n1709 VSS.n1707 0.4505
R24062 VSS.n1949 VSS.n1948 0.4505
R24063 VSS.n1714 VSS.n1710 0.4505
R24064 VSS.n1944 VSS.n1943 0.4505
R24065 VSS.n1935 VSS.n1713 0.4505
R24066 VSS.n1934 VSS.n1933 0.4505
R24067 VSS.n1717 VSS.n1716 0.4505
R24068 VSS.n1929 VSS.n1928 0.4505
R24069 VSS.n1927 VSS.n1719 0.4505
R24070 VSS.n1926 VSS.n1925 0.4505
R24071 VSS.n1721 VSS.n1720 0.4505
R24072 VSS.n1921 VSS.n1920 0.4505
R24073 VSS.n1725 VSS.n1723 0.4505
R24074 VSS.n1751 VSS.n1749 0.4505
R24075 VSS.n1911 VSS.n1910 0.4505
R24076 VSS.n1756 VSS.n1752 0.4505
R24077 VSS.n1906 VSS.n1905 0.4505
R24078 VSS.n1897 VSS.n1755 0.4505
R24079 VSS.n1896 VSS.n1895 0.4505
R24080 VSS.n1759 VSS.n1758 0.4505
R24081 VSS.n1891 VSS.n1890 0.4505
R24082 VSS.n1889 VSS.n1761 0.4505
R24083 VSS.n1888 VSS.n1887 0.4505
R24084 VSS.n1766 VSS.n1763 0.4505
R24085 VSS.n1883 VSS.n1882 0.4505
R24086 VSS.n1768 VSS.n1765 0.4505
R24087 VSS.n1779 VSS.n1777 0.4505
R24088 VSS.n1872 VSS.n1871 0.4505
R24089 VSS.n1784 VSS.n1780 0.4505
R24090 VSS.n1867 VSS.n1866 0.4505
R24091 VSS.n1865 VSS.n1783 0.4505
R24092 VSS.n1864 VSS.n1863 0.4505
R24093 VSS.n1789 VSS.n1788 0.4505
R24094 VSS.n1859 VSS.n1858 0.4505
R24095 VSS.n1798 VSS.n1791 0.4505
R24096 VSS.n1853 VSS.n1852 0.4505
R24097 VSS.n1822 VSS.n1821 0.4505
R24098 VSS.n1848 VSS.n1847 0.4505
R24099 VSS.n1846 VSS.n1824 0.4505
R24100 VSS.n1845 VSS.n1844 0.4505
R24101 VSS.n1826 VSS.n1825 0.4505
R24102 VSS.n1840 VSS.n23 0.4505
R24103 VSS.n1839 VSS.n1838 0.4505
R24104 VSS.n1585 VSS.n1584 0.4505
R24105 VSS.n1583 VSS.n1301 0.4505
R24106 VSS.n1582 VSS.n1581 0.4505
R24107 VSS.n1304 VSS.n1303 0.4505
R24108 VSS.n1577 VSS.n1576 0.4505
R24109 VSS.n1575 VSS.n1306 0.4505
R24110 VSS.n1574 VSS.n1573 0.4505
R24111 VSS.n1308 VSS.n1307 0.4505
R24112 VSS.n1569 VSS.n1568 0.4505
R24113 VSS.n1567 VSS.n1310 0.4505
R24114 VSS.n1566 VSS.n1565 0.4505
R24115 VSS.n1312 VSS.n1311 0.4505
R24116 VSS.n1561 VSS.n1560 0.4505
R24117 VSS.n1559 VSS.n1314 0.4505
R24118 VSS.n1558 VSS.n1557 0.4505
R24119 VSS.n1316 VSS.n1315 0.4505
R24120 VSS.n1553 VSS.n1552 0.4505
R24121 VSS.n1551 VSS.n1318 0.4505
R24122 VSS.n1550 VSS.n1549 0.4505
R24123 VSS.n1320 VSS.n1319 0.4505
R24124 VSS.n1545 VSS.n1544 0.4505
R24125 VSS.n1543 VSS.n1322 0.4505
R24126 VSS.n1542 VSS.n1541 0.4505
R24127 VSS.n1324 VSS.n1323 0.4505
R24128 VSS.n1537 VSS.n1536 0.4505
R24129 VSS.n1535 VSS.n1326 0.4505
R24130 VSS.n1534 VSS.n1533 0.4505
R24131 VSS.n1328 VSS.n1327 0.4505
R24132 VSS.n1529 VSS.n1528 0.4505
R24133 VSS.n1527 VSS.n1330 0.4505
R24134 VSS.n1526 VSS.n1525 0.4505
R24135 VSS.n1332 VSS.n1331 0.4505
R24136 VSS.n1521 VSS.n1520 0.4505
R24137 VSS.n1519 VSS.n1334 0.4505
R24138 VSS.n1518 VSS.n1517 0.4505
R24139 VSS.n1336 VSS.n1335 0.4505
R24140 VSS.n1513 VSS.n1512 0.4505
R24141 VSS.n1511 VSS.n1338 0.4505
R24142 VSS.n1510 VSS.n1509 0.4505
R24143 VSS.n1340 VSS.n1339 0.4505
R24144 VSS.n1505 VSS.n1504 0.4505
R24145 VSS.n1503 VSS.n1342 0.4505
R24146 VSS.n1502 VSS.n1501 0.4505
R24147 VSS.n1344 VSS.n1343 0.4505
R24148 VSS.n1497 VSS.n1496 0.4505
R24149 VSS.n1495 VSS.n1346 0.4505
R24150 VSS.n1494 VSS.n1493 0.4505
R24151 VSS.n1348 VSS.n1347 0.4505
R24152 VSS.n1489 VSS.n1488 0.4505
R24153 VSS.n1487 VSS.n1350 0.4505
R24154 VSS.n1486 VSS.n1485 0.4505
R24155 VSS.n1352 VSS.n1351 0.4505
R24156 VSS.n1481 VSS.n1480 0.4505
R24157 VSS.n1479 VSS.n1354 0.4505
R24158 VSS.n1478 VSS.n1477 0.4505
R24159 VSS.n1356 VSS.n1355 0.4505
R24160 VSS.n1473 VSS.n1472 0.4505
R24161 VSS.n1471 VSS.n1358 0.4505
R24162 VSS.n1470 VSS.n1469 0.4505
R24163 VSS.n1360 VSS.n1359 0.4505
R24164 VSS.n1465 VSS.n1464 0.4505
R24165 VSS.n1463 VSS.n1362 0.4505
R24166 VSS.n1462 VSS.n1461 0.4505
R24167 VSS.n1364 VSS.n1363 0.4505
R24168 VSS.n1457 VSS.n1456 0.4505
R24169 VSS.n1455 VSS.n1366 0.4505
R24170 VSS.n1454 VSS.n1453 0.4505
R24171 VSS.n1368 VSS.n1367 0.4505
R24172 VSS.n1449 VSS.n1448 0.4505
R24173 VSS.n1447 VSS.n1370 0.4505
R24174 VSS.n1446 VSS.n1445 0.4505
R24175 VSS.n1372 VSS.n1371 0.4505
R24176 VSS.n1441 VSS.n1440 0.4505
R24177 VSS.n1439 VSS.n1374 0.4505
R24178 VSS.n1438 VSS.n1437 0.4505
R24179 VSS.n1376 VSS.n1375 0.4505
R24180 VSS.n1433 VSS.n1432 0.4505
R24181 VSS.n1431 VSS.n1378 0.4505
R24182 VSS.n1430 VSS.n1429 0.4505
R24183 VSS.n1380 VSS.n1379 0.4505
R24184 VSS.n1425 VSS.n1424 0.4505
R24185 VSS.n1423 VSS.n1382 0.4505
R24186 VSS.n1422 VSS.n1421 0.4505
R24187 VSS.n1384 VSS.n1383 0.4505
R24188 VSS.n1417 VSS.n1416 0.4505
R24189 VSS.n1415 VSS.n1386 0.4505
R24190 VSS.n1414 VSS.n1413 0.4505
R24191 VSS.n1388 VSS.n1387 0.4505
R24192 VSS.n1409 VSS.n1408 0.4505
R24193 VSS.n1407 VSS.n1390 0.4505
R24194 VSS.n1406 VSS.n1405 0.4505
R24195 VSS.n1392 VSS.n1391 0.4505
R24196 VSS.n1401 VSS.n1400 0.4505
R24197 VSS.n1399 VSS.n1394 0.4505
R24198 VSS.n1398 VSS.n1397 0.4505
R24199 VSS.n1300 VSS.n1298 0.4505
R24200 VSS.n1586 VSS.n1585 0.4505
R24201 VSS.n1301 VSS.n1299 0.4505
R24202 VSS.n1581 VSS.n1580 0.4505
R24203 VSS.n1579 VSS.n1304 0.4505
R24204 VSS.n1578 VSS.n1577 0.4505
R24205 VSS.n1306 VSS.n1305 0.4505
R24206 VSS.n1573 VSS.n1572 0.4505
R24207 VSS.n1571 VSS.n1308 0.4505
R24208 VSS.n1570 VSS.n1569 0.4505
R24209 VSS.n1310 VSS.n1309 0.4505
R24210 VSS.n1565 VSS.n1564 0.4505
R24211 VSS.n1563 VSS.n1312 0.4505
R24212 VSS.n1562 VSS.n1561 0.4505
R24213 VSS.n1314 VSS.n1313 0.4505
R24214 VSS.n1557 VSS.n1556 0.4505
R24215 VSS.n1555 VSS.n1316 0.4505
R24216 VSS.n1554 VSS.n1553 0.4505
R24217 VSS.n1318 VSS.n1317 0.4505
R24218 VSS.n1549 VSS.n1548 0.4505
R24219 VSS.n1547 VSS.n1320 0.4505
R24220 VSS.n1546 VSS.n1545 0.4505
R24221 VSS.n1322 VSS.n1321 0.4505
R24222 VSS.n1541 VSS.n1540 0.4505
R24223 VSS.n1539 VSS.n1324 0.4505
R24224 VSS.n1538 VSS.n1537 0.4505
R24225 VSS.n1326 VSS.n1325 0.4505
R24226 VSS.n1533 VSS.n1532 0.4505
R24227 VSS.n1531 VSS.n1328 0.4505
R24228 VSS.n1530 VSS.n1529 0.4505
R24229 VSS.n1330 VSS.n1329 0.4505
R24230 VSS.n1525 VSS.n1524 0.4505
R24231 VSS.n1523 VSS.n1332 0.4505
R24232 VSS.n1522 VSS.n1521 0.4505
R24233 VSS.n1334 VSS.n1333 0.4505
R24234 VSS.n1517 VSS.n1516 0.4505
R24235 VSS.n1515 VSS.n1336 0.4505
R24236 VSS.n1514 VSS.n1513 0.4505
R24237 VSS.n1338 VSS.n1337 0.4505
R24238 VSS.n1509 VSS.n1508 0.4505
R24239 VSS.n1507 VSS.n1340 0.4505
R24240 VSS.n1506 VSS.n1505 0.4505
R24241 VSS.n1342 VSS.n1341 0.4505
R24242 VSS.n1501 VSS.n1500 0.4505
R24243 VSS.n1499 VSS.n1344 0.4505
R24244 VSS.n1498 VSS.n1497 0.4505
R24245 VSS.n1346 VSS.n1345 0.4505
R24246 VSS.n1493 VSS.n1492 0.4505
R24247 VSS.n1491 VSS.n1348 0.4505
R24248 VSS.n1490 VSS.n1489 0.4505
R24249 VSS.n1350 VSS.n1349 0.4505
R24250 VSS.n1485 VSS.n1484 0.4505
R24251 VSS.n1483 VSS.n1352 0.4505
R24252 VSS.n1482 VSS.n1481 0.4505
R24253 VSS.n1354 VSS.n1353 0.4505
R24254 VSS.n1477 VSS.n1476 0.4505
R24255 VSS.n1475 VSS.n1356 0.4505
R24256 VSS.n1474 VSS.n1473 0.4505
R24257 VSS.n1358 VSS.n1357 0.4505
R24258 VSS.n1469 VSS.n1468 0.4505
R24259 VSS.n1467 VSS.n1360 0.4505
R24260 VSS.n1466 VSS.n1465 0.4505
R24261 VSS.n1362 VSS.n1361 0.4505
R24262 VSS.n1461 VSS.n1460 0.4505
R24263 VSS.n1459 VSS.n1364 0.4505
R24264 VSS.n1458 VSS.n1457 0.4505
R24265 VSS.n1366 VSS.n1365 0.4505
R24266 VSS.n1453 VSS.n1452 0.4505
R24267 VSS.n1451 VSS.n1368 0.4505
R24268 VSS.n1450 VSS.n1449 0.4505
R24269 VSS.n1370 VSS.n1369 0.4505
R24270 VSS.n1445 VSS.n1444 0.4505
R24271 VSS.n1443 VSS.n1372 0.4505
R24272 VSS.n1442 VSS.n1441 0.4505
R24273 VSS.n1374 VSS.n1373 0.4505
R24274 VSS.n1437 VSS.n1436 0.4505
R24275 VSS.n1435 VSS.n1376 0.4505
R24276 VSS.n1434 VSS.n1433 0.4505
R24277 VSS.n1378 VSS.n1377 0.4505
R24278 VSS.n1429 VSS.n1428 0.4505
R24279 VSS.n1427 VSS.n1380 0.4505
R24280 VSS.n1426 VSS.n1425 0.4505
R24281 VSS.n1382 VSS.n1381 0.4505
R24282 VSS.n1421 VSS.n1420 0.4505
R24283 VSS.n1419 VSS.n1384 0.4505
R24284 VSS.n1418 VSS.n1417 0.4505
R24285 VSS.n1386 VSS.n1385 0.4505
R24286 VSS.n1413 VSS.n1412 0.4505
R24287 VSS.n1411 VSS.n1388 0.4505
R24288 VSS.n1410 VSS.n1409 0.4505
R24289 VSS.n1390 VSS.n1389 0.4505
R24290 VSS.n1405 VSS.n1404 0.4505
R24291 VSS.n1403 VSS.n1392 0.4505
R24292 VSS.n1402 VSS.n1401 0.4505
R24293 VSS.n1394 VSS.n1393 0.4505
R24294 VSS.n1397 VSS.n1396 0.4505
R24295 VSS.n3188 VSS.n3187 0.4505
R24296 VSS.n3189 VSS.n3182 0.4505
R24297 VSS.n3191 VSS.n3190 0.4505
R24298 VSS.n3180 VSS.n3179 0.4505
R24299 VSS.n3196 VSS.n3195 0.4505
R24300 VSS.n3197 VSS.n3178 0.4505
R24301 VSS.n3199 VSS.n3198 0.4505
R24302 VSS.n3176 VSS.n3175 0.4505
R24303 VSS.n3204 VSS.n3203 0.4505
R24304 VSS.n3205 VSS.n3174 0.4505
R24305 VSS.n3207 VSS.n3206 0.4505
R24306 VSS.n3172 VSS.n3171 0.4505
R24307 VSS.n3212 VSS.n3211 0.4505
R24308 VSS.n3213 VSS.n3170 0.4505
R24309 VSS.n3215 VSS.n3214 0.4505
R24310 VSS.n3168 VSS.n3167 0.4505
R24311 VSS.n3220 VSS.n3219 0.4505
R24312 VSS.n3221 VSS.n3166 0.4505
R24313 VSS.n3223 VSS.n3222 0.4505
R24314 VSS.n3164 VSS.n3163 0.4505
R24315 VSS.n3228 VSS.n3227 0.4505
R24316 VSS.n3229 VSS.n3162 0.4505
R24317 VSS.n3231 VSS.n3230 0.4505
R24318 VSS.n3160 VSS.n3159 0.4505
R24319 VSS.n3236 VSS.n3235 0.4505
R24320 VSS.n3237 VSS.n3158 0.4505
R24321 VSS.n3239 VSS.n3238 0.4505
R24322 VSS.n3156 VSS.n3155 0.4505
R24323 VSS.n3244 VSS.n3243 0.4505
R24324 VSS.n3245 VSS.n3152 0.4505
R24325 VSS.n3281 VSS.n3280 0.4505
R24326 VSS.n3276 VSS.n3149 0.4505
R24327 VSS.n3286 VSS.n3285 0.4505
R24328 VSS.n3148 VSS.n3146 0.4505
R24329 VSS.n3090 VSS.n3087 0.4505
R24330 VSS.n3297 VSS.n3296 0.4505
R24331 VSS.n3088 VSS.n3084 0.4505
R24332 VSS.n3302 VSS.n3301 0.4505
R24333 VSS.n3083 VSS.n3080 0.4505
R24334 VSS.n3104 VSS.n3103 0.4505
R24335 VSS.n3128 VSS.n3127 0.4505
R24336 VSS.n3102 VSS.n3100 0.4505
R24337 VSS.n3122 VSS.n3121 0.4505
R24338 VSS.n3112 VSS.n3106 0.4505
R24339 VSS.n2959 VSS.n2956 0.4505
R24340 VSS.n3326 VSS.n3325 0.4505
R24341 VSS.n2953 VSS.n2951 0.4505
R24342 VSS.n3331 VSS.n3330 0.4505
R24343 VSS.n2952 VSS.n2950 0.4505
R24344 VSS.n3064 VSS.n3063 0.4505
R24345 VSS.n2932 VSS.n2929 0.4505
R24346 VSS.n3344 VSS.n3343 0.4505
R24347 VSS.n2930 VSS.n2926 0.4505
R24348 VSS.n3349 VSS.n3348 0.4505
R24349 VSS.n2925 VSS.n2923 0.4505
R24350 VSS.n3002 VSS.n3001 0.4505
R24351 VSS.n2980 VSS.n2979 0.4505
R24352 VSS.n2904 VSS.n2902 0.4505
R24353 VSS.n2988 VSS.n2987 0.4505
R24354 VSS.n2992 VSS.n2991 0.4505
R24355 VSS.n2983 VSS.n2982 0.4505
R24356 VSS.n2997 VSS.n2996 0.4505
R24357 VSS.n3379 VSS.n3378 0.4505
R24358 VSS.n3377 VSS.n2894 0.4505
R24359 VSS.n2898 VSS.n2895 0.4505
R24360 VSS.n3373 VSS.n3372 0.4505
R24361 VSS.n3371 VSS.n2897 0.4505
R24362 VSS.n3370 VSS.n3369 0.4505
R24363 VSS.n3015 VSS.n2900 0.4505
R24364 VSS.n3365 VSS.n3364 0.4505
R24365 VSS.n2381 VSS.n2375 0.4505
R24366 VSS.n4237 VSS.n4236 0.4505
R24367 VSS.n4235 VSS.n2376 0.4505
R24368 VSS.n4234 VSS.n4233 0.4505
R24369 VSS.n2383 VSS.n2382 0.4505
R24370 VSS.n4228 VSS.n4227 0.4505
R24371 VSS.n4226 VSS.n2385 0.4505
R24372 VSS.n4225 VSS.n4224 0.4505
R24373 VSS.n2387 VSS.n2386 0.4505
R24374 VSS.n4218 VSS.n4217 0.4505
R24375 VSS.n4216 VSS.n2389 0.4505
R24376 VSS.n4215 VSS.n4214 0.4505
R24377 VSS.n2391 VSS.n2390 0.4505
R24378 VSS.n4210 VSS.n4209 0.4505
R24379 VSS.n4208 VSS.n2394 0.4505
R24380 VSS.n4207 VSS.n4206 0.4505
R24381 VSS.n2396 VSS.n2395 0.4505
R24382 VSS.n4200 VSS.n4199 0.4505
R24383 VSS.n4198 VSS.n2399 0.4505
R24384 VSS.n4197 VSS.n4196 0.4505
R24385 VSS.n2401 VSS.n2400 0.4505
R24386 VSS.n4192 VSS.n4191 0.4505
R24387 VSS.n4190 VSS.n2404 0.4505
R24388 VSS.n4189 VSS.n4188 0.4505
R24389 VSS.n2406 VSS.n2405 0.4505
R24390 VSS.n4169 VSS.n4168 0.4505
R24391 VSS.n4167 VSS.n2415 0.4505
R24392 VSS.n4166 VSS.n4165 0.4505
R24393 VSS.n2417 VSS.n2416 0.4505
R24394 VSS.n4161 VSS.n4160 0.4505
R24395 VSS.n4159 VSS.n2419 0.4505
R24396 VSS.n4158 VSS.n4157 0.4505
R24397 VSS.n2421 VSS.n2420 0.4505
R24398 VSS.n4153 VSS.n4152 0.4505
R24399 VSS.n4151 VSS.n2423 0.4505
R24400 VSS.n4150 VSS.n4149 0.4505
R24401 VSS.n2425 VSS.n2424 0.4505
R24402 VSS.n4097 VSS.n4095 0.4505
R24403 VSS.n4100 VSS.n4099 0.4505
R24404 VSS.n4098 VSS.n4096 0.4505
R24405 VSS.n2442 VSS.n2441 0.4505
R24406 VSS.n4110 VSS.n4109 0.4505
R24407 VSS.n4111 VSS.n2440 0.4505
R24408 VSS.n4113 VSS.n4112 0.4505
R24409 VSS.n2438 VSS.n2437 0.4505
R24410 VSS.n4120 VSS.n4119 0.4505
R24411 VSS.n4121 VSS.n2435 0.4505
R24412 VSS.n4137 VSS.n4136 0.4505
R24413 VSS.n4135 VSS.n2436 0.4505
R24414 VSS.n4134 VSS.n4133 0.4505
R24415 VSS.n4123 VSS.n4122 0.4505
R24416 VSS.n4128 VSS.n4127 0.4505
R24417 VSS.n4126 VSS.n4125 0.4505
R24418 VSS.n2247 VSS.n2245 0.4505
R24419 VSS.n5235 VSS.n5234 0.4505
R24420 VSS.n5233 VSS.n2246 0.4505
R24421 VSS.n5232 VSS.n5231 0.4505
R24422 VSS.n2249 VSS.n2248 0.4505
R24423 VSS.n5227 VSS.n5226 0.4505
R24424 VSS.n5225 VSS.n2252 0.4505
R24425 VSS.n5224 VSS.n5223 0.4505
R24426 VSS.n2254 VSS.n2253 0.4505
R24427 VSS.n5219 VSS.n5218 0.4505
R24428 VSS.n5217 VSS.n2256 0.4505
R24429 VSS.n5216 VSS.n5215 0.4505
R24430 VSS.n2258 VSS.n2257 0.4505
R24431 VSS.n5211 VSS.n5210 0.4505
R24432 VSS.n5209 VSS.n2260 0.4505
R24433 VSS.n5208 VSS.n5207 0.4505
R24434 VSS.n2262 VSS.n2261 0.4505
R24435 VSS.n5203 VSS.n5202 0.4505
R24436 VSS.n5201 VSS.n2264 0.4505
R24437 VSS.n5200 VSS.n5199 0.4505
R24438 VSS.n2266 VSS.n2265 0.4505
R24439 VSS.n5195 VSS.n5194 0.4505
R24440 VSS.n5193 VSS.n2268 0.4505
R24441 VSS.n5192 VSS.n5191 0.4505
R24442 VSS.n2270 VSS.n2269 0.4505
R24443 VSS.n5187 VSS.n5186 0.4505
R24444 VSS.n5185 VSS.n5172 0.4505
R24445 VSS.n5184 VSS.n5183 0.4505
R24446 VSS.n5174 VSS.n5173 0.4505
R24447 VSS.n5179 VSS.n5178 0.4505
R24448 VSS.n5177 VSS.n5176 0.4505
R24449 VSS.n5180 VSS.n5179 0.4505
R24450 VSS.n5181 VSS.n5174 0.4505
R24451 VSS.n5183 VSS.n5182 0.4505
R24452 VSS.n5172 VSS.n5171 0.4505
R24453 VSS.n5188 VSS.n5187 0.4505
R24454 VSS.n5189 VSS.n2270 0.4505
R24455 VSS.n5191 VSS.n5190 0.4505
R24456 VSS.n2268 VSS.n2267 0.4505
R24457 VSS.n5196 VSS.n5195 0.4505
R24458 VSS.n5197 VSS.n2266 0.4505
R24459 VSS.n5199 VSS.n5198 0.4505
R24460 VSS.n2264 VSS.n2263 0.4505
R24461 VSS.n5204 VSS.n5203 0.4505
R24462 VSS.n5205 VSS.n2262 0.4505
R24463 VSS.n5207 VSS.n5206 0.4505
R24464 VSS.n2260 VSS.n2259 0.4505
R24465 VSS.n5212 VSS.n5211 0.4505
R24466 VSS.n5213 VSS.n2258 0.4505
R24467 VSS.n5215 VSS.n5214 0.4505
R24468 VSS.n2256 VSS.n2255 0.4505
R24469 VSS.n5220 VSS.n5219 0.4505
R24470 VSS.n5221 VSS.n2254 0.4505
R24471 VSS.n5223 VSS.n5222 0.4505
R24472 VSS.n2252 VSS.n2251 0.4505
R24473 VSS.n5228 VSS.n5227 0.4505
R24474 VSS.n5229 VSS.n2249 0.4505
R24475 VSS.n5231 VSS.n5230 0.4505
R24476 VSS.n2250 VSS.n2246 0.4505
R24477 VSS.n5236 VSS.n5235 0.4505
R24478 VSS.n2245 VSS.n2243 0.4505
R24479 VSS.n4125 VSS.n4124 0.4505
R24480 VSS.n4129 VSS.n4128 0.4505
R24481 VSS.n4131 VSS.n4123 0.4505
R24482 VSS.n4133 VSS.n4132 0.4505
R24483 VSS.n2436 VSS.n2434 0.4505
R24484 VSS.n4138 VSS.n4137 0.4505
R24485 VSS.n2435 VSS.n2433 0.4505
R24486 VSS.n4119 VSS.n4118 0.4505
R24487 VSS.n4115 VSS.n2438 0.4505
R24488 VSS.n4114 VSS.n4113 0.4505
R24489 VSS.n2440 VSS.n2439 0.4505
R24490 VSS.n4109 VSS.n4108 0.4505
R24491 VSS.n2443 VSS.n2442 0.4505
R24492 VSS.n4096 VSS.n4094 0.4505
R24493 VSS.n4101 VSS.n4100 0.4505
R24494 VSS.n4095 VSS.n4093 0.4505
R24495 VSS.n2426 VSS.n2425 0.4505
R24496 VSS.n4149 VSS.n4148 0.4505
R24497 VSS.n2423 VSS.n2422 0.4505
R24498 VSS.n4154 VSS.n4153 0.4505
R24499 VSS.n4155 VSS.n2421 0.4505
R24500 VSS.n4157 VSS.n4156 0.4505
R24501 VSS.n2419 VSS.n2418 0.4505
R24502 VSS.n4162 VSS.n4161 0.4505
R24503 VSS.n4163 VSS.n2417 0.4505
R24504 VSS.n4165 VSS.n4164 0.4505
R24505 VSS.n2415 VSS.n2414 0.4505
R24506 VSS.n4170 VSS.n4169 0.4505
R24507 VSS.n4171 VSS.n2406 0.4505
R24508 VSS.n4188 VSS.n4187 0.4505
R24509 VSS.n2407 VSS.n2404 0.4505
R24510 VSS.n4193 VSS.n4192 0.4505
R24511 VSS.n4194 VSS.n2401 0.4505
R24512 VSS.n4196 VSS.n4195 0.4505
R24513 VSS.n2402 VSS.n2399 0.4505
R24514 VSS.n4201 VSS.n4200 0.4505
R24515 VSS.n4204 VSS.n2396 0.4505
R24516 VSS.n4206 VSS.n4205 0.4505
R24517 VSS.n2397 VSS.n2394 0.4505
R24518 VSS.n4211 VSS.n4210 0.4505
R24519 VSS.n4212 VSS.n2391 0.4505
R24520 VSS.n4214 VSS.n4213 0.4505
R24521 VSS.n2392 VSS.n2389 0.4505
R24522 VSS.n4219 VSS.n4218 0.4505
R24523 VSS.n4221 VSS.n2387 0.4505
R24524 VSS.n4224 VSS.n4223 0.4505
R24525 VSS.n2385 VSS.n2384 0.4505
R24526 VSS.n4229 VSS.n4228 0.4505
R24527 VSS.n4230 VSS.n2383 0.4505
R24528 VSS.n4233 VSS.n4232 0.4505
R24529 VSS.n2376 VSS.n2374 0.4505
R24530 VSS.n4238 VSS.n4237 0.4505
R24531 VSS.n2375 VSS.n2373 0.4505
R24532 VSS.n2379 VSS.n2378 0.4505
R24533 VSS.n2546 VSS.n2545 0.4505
R24534 VSS.n2550 VSS.n2549 0.4505
R24535 VSS.n2551 VSS.n2544 0.4505
R24536 VSS.n2553 VSS.n2552 0.4505
R24537 VSS.n2542 VSS.n2541 0.4505
R24538 VSS.n2558 VSS.n2557 0.4505
R24539 VSS.n2559 VSS.n2540 0.4505
R24540 VSS.n2561 VSS.n2560 0.4505
R24541 VSS.n2538 VSS.n2537 0.4505
R24542 VSS.n2566 VSS.n2565 0.4505
R24543 VSS.n2567 VSS.n2536 0.4505
R24544 VSS.n2569 VSS.n2568 0.4505
R24545 VSS.n2534 VSS.n2533 0.4505
R24546 VSS.n2574 VSS.n2573 0.4505
R24547 VSS.n2575 VSS.n2532 0.4505
R24548 VSS.n2577 VSS.n2576 0.4505
R24549 VSS.n2530 VSS.n2529 0.4505
R24550 VSS.n2582 VSS.n2581 0.4505
R24551 VSS.n2583 VSS.n2528 0.4505
R24552 VSS.n2585 VSS.n2584 0.4505
R24553 VSS.n2526 VSS.n2525 0.4505
R24554 VSS.n2590 VSS.n2589 0.4505
R24555 VSS.n2591 VSS.n2524 0.4505
R24556 VSS.n2593 VSS.n2592 0.4505
R24557 VSS.n2522 VSS.n2521 0.4505
R24558 VSS.n2598 VSS.n2597 0.4505
R24559 VSS.n2599 VSS.n2520 0.4505
R24560 VSS.n2601 VSS.n2600 0.4505
R24561 VSS.n2518 VSS.n2517 0.4505
R24562 VSS.n2606 VSS.n2605 0.4505
R24563 VSS.n2607 VSS.n2516 0.4505
R24564 VSS.n2609 VSS.n2608 0.4505
R24565 VSS.n2514 VSS.n2513 0.4505
R24566 VSS.n2614 VSS.n2613 0.4505
R24567 VSS.n2615 VSS.n2512 0.4505
R24568 VSS.n2617 VSS.n2616 0.4505
R24569 VSS.n2510 VSS.n2509 0.4505
R24570 VSS.n2622 VSS.n2621 0.4505
R24571 VSS.n2623 VSS.n2508 0.4505
R24572 VSS.n2625 VSS.n2624 0.4505
R24573 VSS.n2506 VSS.n2505 0.4505
R24574 VSS.n2630 VSS.n2629 0.4505
R24575 VSS.n2631 VSS.n2504 0.4505
R24576 VSS.n2633 VSS.n2632 0.4505
R24577 VSS.n2502 VSS.n2501 0.4505
R24578 VSS.n2638 VSS.n2637 0.4505
R24579 VSS.n2639 VSS.n2500 0.4505
R24580 VSS.n2641 VSS.n2640 0.4505
R24581 VSS.n2498 VSS.n2497 0.4505
R24582 VSS.n2646 VSS.n2645 0.4505
R24583 VSS.n2647 VSS.n2496 0.4505
R24584 VSS.n2649 VSS.n2648 0.4505
R24585 VSS.n2494 VSS.n2493 0.4505
R24586 VSS.n2654 VSS.n2653 0.4505
R24587 VSS.n2655 VSS.n2492 0.4505
R24588 VSS.n2657 VSS.n2656 0.4505
R24589 VSS.n2490 VSS.n2489 0.4505
R24590 VSS.n2662 VSS.n2661 0.4505
R24591 VSS.n2663 VSS.n2488 0.4505
R24592 VSS.n2665 VSS.n2664 0.4505
R24593 VSS.n2486 VSS.n2485 0.4505
R24594 VSS.n2670 VSS.n2669 0.4505
R24595 VSS.n2671 VSS.n2484 0.4505
R24596 VSS.n2673 VSS.n2672 0.4505
R24597 VSS.n2482 VSS.n2481 0.4505
R24598 VSS.n2679 VSS.n2678 0.4505
R24599 VSS.n2680 VSS.n2479 0.4505
R24600 VSS.n2682 VSS.n2681 0.4505
R24601 VSS.n2683 VSS.n2463 0.4505
R24602 VSS.n2684 VSS.n2468 0.4505
R24603 VSS.n2697 VSS.n2696 0.4505
R24604 VSS.n2688 VSS.n2477 0.4505
R24605 VSS.n2692 VSS.n2691 0.4505
R24606 VSS.n2690 VSS.n2687 0.4505
R24607 VSS.n2316 VSS.n2315 0.4505
R24608 VSS.n2317 VSS.n2310 0.4505
R24609 VSS.n2319 VSS.n2318 0.4505
R24610 VSS.n2308 VSS.n2307 0.4505
R24611 VSS.n2324 VSS.n2323 0.4505
R24612 VSS.n2325 VSS.n2306 0.4505
R24613 VSS.n2327 VSS.n2326 0.4505
R24614 VSS.n2304 VSS.n2303 0.4505
R24615 VSS.n2332 VSS.n2331 0.4505
R24616 VSS.n2333 VSS.n2302 0.4505
R24617 VSS.n2335 VSS.n2334 0.4505
R24618 VSS.n2299 VSS.n2297 0.4505
R24619 VSS.n4281 VSS.n4280 0.4505
R24620 VSS.n2300 VSS.n2298 0.4505
R24621 VSS.n4276 VSS.n4275 0.4505
R24622 VSS.n4274 VSS.n2339 0.4505
R24623 VSS.n4273 VSS.n4272 0.4505
R24624 VSS.n2341 VSS.n2340 0.4505
R24625 VSS.n4268 VSS.n4267 0.4505
R24626 VSS.n4266 VSS.n2343 0.4505
R24627 VSS.n4265 VSS.n4264 0.4505
R24628 VSS.n2345 VSS.n2344 0.4505
R24629 VSS.n4260 VSS.n4259 0.4505
R24630 VSS.n4258 VSS.n2347 0.4505
R24631 VSS.n4257 VSS.n4256 0.4505
R24632 VSS.n2349 VSS.n2348 0.4505
R24633 VSS.n4252 VSS.n4251 0.4505
R24634 VSS.n2352 VSS.n2351 0.4505
R24635 VSS.n5703 VSS.n5 0.4505
R24636 VSS.n5705 VSS.n5704 0.4505
R24637 VSS.n6 VSS.n2 0.4505
R24638 VSS.n5710 VSS.n5709 0.4505
R24639 VSS.n4025 VSS.n4024 0.4505
R24640 VSS.n4023 VSS.n2703 0.4505
R24641 VSS.n4017 VSS.n2704 0.4505
R24642 VSS.n4019 VSS.n4018 0.4505
R24643 VSS.n4016 VSS.n2706 0.4505
R24644 VSS.n4015 VSS.n4014 0.4505
R24645 VSS.n2708 VSS.n2707 0.4505
R24646 VSS.n4010 VSS.n4009 0.4505
R24647 VSS.n4008 VSS.n2710 0.4505
R24648 VSS.n4007 VSS.n4006 0.4505
R24649 VSS.n2712 VSS.n2711 0.4505
R24650 VSS.n4002 VSS.n4001 0.4505
R24651 VSS.n4000 VSS.n2714 0.4505
R24652 VSS.n3999 VSS.n3998 0.4505
R24653 VSS.n2716 VSS.n2715 0.4505
R24654 VSS.n3994 VSS.n3993 0.4505
R24655 VSS.n3992 VSS.n2718 0.4505
R24656 VSS.n3991 VSS.n3990 0.4505
R24657 VSS.n2720 VSS.n2719 0.4505
R24658 VSS.n3986 VSS.n3985 0.4505
R24659 VSS.n3984 VSS.n2722 0.4505
R24660 VSS.n3983 VSS.n3982 0.4505
R24661 VSS.n2724 VSS.n2723 0.4505
R24662 VSS.n3978 VSS.n3977 0.4505
R24663 VSS.n3976 VSS.n2726 0.4505
R24664 VSS.n3975 VSS.n3974 0.4505
R24665 VSS.n2728 VSS.n2727 0.4505
R24666 VSS.n3970 VSS.n3969 0.4505
R24667 VSS.n3968 VSS.n2730 0.4505
R24668 VSS.n3967 VSS.n3966 0.4505
R24669 VSS.n2732 VSS.n2731 0.4505
R24670 VSS.n3962 VSS.n3961 0.4505
R24671 VSS.n3960 VSS.n2734 0.4505
R24672 VSS.n3959 VSS.n3958 0.4505
R24673 VSS.n2736 VSS.n2735 0.4505
R24674 VSS.n3954 VSS.n3953 0.4505
R24675 VSS.n3952 VSS.n2738 0.4505
R24676 VSS.n3950 VSS.n3949 0.4505
R24677 VSS.n2740 VSS.n2739 0.4505
R24678 VSS.n3945 VSS.n3944 0.4505
R24679 VSS.n3943 VSS.n2742 0.4505
R24680 VSS.n3942 VSS.n3941 0.4505
R24681 VSS.n2744 VSS.n2743 0.4505
R24682 VSS.n3937 VSS.n3936 0.4505
R24683 VSS.n3935 VSS.n2746 0.4505
R24684 VSS.n3934 VSS.n3933 0.4505
R24685 VSS.n2748 VSS.n2747 0.4505
R24686 VSS.n3929 VSS.n3928 0.4505
R24687 VSS.n3927 VSS.n2750 0.4505
R24688 VSS.n3926 VSS.n3925 0.4505
R24689 VSS.n2752 VSS.n2751 0.4505
R24690 VSS.n3921 VSS.n3920 0.4505
R24691 VSS.n3919 VSS.n2754 0.4505
R24692 VSS.n3918 VSS.n3917 0.4505
R24693 VSS.n2756 VSS.n2755 0.4505
R24694 VSS.n3913 VSS.n3912 0.4505
R24695 VSS.n3911 VSS.n2758 0.4505
R24696 VSS.n3910 VSS.n3909 0.4505
R24697 VSS.n2760 VSS.n2759 0.4505
R24698 VSS.n3905 VSS.n3904 0.4505
R24699 VSS.n3903 VSS.n2762 0.4505
R24700 VSS.n3902 VSS.n3901 0.4505
R24701 VSS.n2764 VSS.n2763 0.4505
R24702 VSS.n3897 VSS.n3896 0.4505
R24703 VSS.n3895 VSS.n2766 0.4505
R24704 VSS.n3894 VSS.n3893 0.4505
R24705 VSS.n2768 VSS.n2767 0.4505
R24706 VSS.n3889 VSS.n3888 0.4505
R24707 VSS.n2771 VSS.n2770 0.4505
R24708 VSS.n3884 VSS.n3883 0.4505
R24709 VSS.n2778 VSS.n2774 0.4505
R24710 VSS.n3879 VSS.n3878 0.4505
R24711 VSS.n3479 VSS.n2776 0.4505
R24712 VSS.n3483 VSS.n3482 0.4505
R24713 VSS.n3477 VSS.n3476 0.4505
R24714 VSS.n3488 VSS.n3487 0.4505
R24715 VSS.n3474 VSS.n3473 0.4505
R24716 VSS.n3493 VSS.n3492 0.4505
R24717 VSS.n3494 VSS.n3472 0.4505
R24718 VSS.n3496 VSS.n3495 0.4505
R24719 VSS.n3423 VSS.n3421 0.4505
R24720 VSS.n3501 VSS.n3500 0.4505
R24721 VSS.n3422 VSS.n3420 0.4505
R24722 VSS.n3468 VSS.n3467 0.4505
R24723 VSS.n3466 VSS.n3425 0.4505
R24724 VSS.n3465 VSS.n3464 0.4505
R24725 VSS.n3427 VSS.n3426 0.4505
R24726 VSS.n3460 VSS.n3459 0.4505
R24727 VSS.n3458 VSS.n3429 0.4505
R24728 VSS.n3457 VSS.n3456 0.4505
R24729 VSS.n3431 VSS.n3430 0.4505
R24730 VSS.n3452 VSS.n3451 0.4505
R24731 VSS.n3450 VSS.n3433 0.4505
R24732 VSS.n3449 VSS.n3448 0.4505
R24733 VSS.n3435 VSS.n3434 0.4505
R24734 VSS.n3444 VSS.n3443 0.4505
R24735 VSS.n3442 VSS.n3437 0.4505
R24736 VSS.n3441 VSS.n3440 0.4505
R24737 VSS.n3437 VSS.n3436 0.4505
R24738 VSS.n3445 VSS.n3444 0.4505
R24739 VSS.n3446 VSS.n3435 0.4505
R24740 VSS.n3448 VSS.n3447 0.4505
R24741 VSS.n3433 VSS.n3432 0.4505
R24742 VSS.n3453 VSS.n3452 0.4505
R24743 VSS.n3454 VSS.n3431 0.4505
R24744 VSS.n3456 VSS.n3455 0.4505
R24745 VSS.n3429 VSS.n3428 0.4505
R24746 VSS.n3461 VSS.n3460 0.4505
R24747 VSS.n3462 VSS.n3427 0.4505
R24748 VSS.n3464 VSS.n3463 0.4505
R24749 VSS.n3425 VSS.n3424 0.4505
R24750 VSS.n3469 VSS.n3468 0.4505
R24751 VSS.n3470 VSS.n3422 0.4505
R24752 VSS.n3500 VSS.n3499 0.4505
R24753 VSS.n3498 VSS.n3423 0.4505
R24754 VSS.n3497 VSS.n3496 0.4505
R24755 VSS.n3472 VSS.n3471 0.4505
R24756 VSS.n3492 VSS.n3491 0.4505
R24757 VSS.n3490 VSS.n3474 0.4505
R24758 VSS.n3489 VSS.n3488 0.4505
R24759 VSS.n3476 VSS.n3475 0.4505
R24760 VSS.n3482 VSS.n3481 0.4505
R24761 VSS.n2776 VSS.n2775 0.4505
R24762 VSS.n3880 VSS.n3879 0.4505
R24763 VSS.n3881 VSS.n2774 0.4505
R24764 VSS.n3883 VSS.n3882 0.4505
R24765 VSS.n2770 VSS.n2769 0.4505
R24766 VSS.n3890 VSS.n3889 0.4505
R24767 VSS.n3891 VSS.n2768 0.4505
R24768 VSS.n3893 VSS.n3892 0.4505
R24769 VSS.n2766 VSS.n2765 0.4505
R24770 VSS.n3898 VSS.n3897 0.4505
R24771 VSS.n3899 VSS.n2764 0.4505
R24772 VSS.n3901 VSS.n3900 0.4505
R24773 VSS.n2762 VSS.n2761 0.4505
R24774 VSS.n3906 VSS.n3905 0.4505
R24775 VSS.n3907 VSS.n2760 0.4505
R24776 VSS.n3909 VSS.n3908 0.4505
R24777 VSS.n2758 VSS.n2757 0.4505
R24778 VSS.n3914 VSS.n3913 0.4505
R24779 VSS.n3915 VSS.n2756 0.4505
R24780 VSS.n3917 VSS.n3916 0.4505
R24781 VSS.n2754 VSS.n2753 0.4505
R24782 VSS.n3922 VSS.n3921 0.4505
R24783 VSS.n3923 VSS.n2752 0.4505
R24784 VSS.n3925 VSS.n3924 0.4505
R24785 VSS.n2750 VSS.n2749 0.4505
R24786 VSS.n3930 VSS.n3929 0.4505
R24787 VSS.n3931 VSS.n2748 0.4505
R24788 VSS.n3933 VSS.n3932 0.4505
R24789 VSS.n2746 VSS.n2745 0.4505
R24790 VSS.n3938 VSS.n3937 0.4505
R24791 VSS.n3939 VSS.n2744 0.4505
R24792 VSS.n3941 VSS.n3940 0.4505
R24793 VSS.n2742 VSS.n2741 0.4505
R24794 VSS.n3946 VSS.n3945 0.4505
R24795 VSS.n3947 VSS.n2740 0.4505
R24796 VSS.n3949 VSS.n3948 0.4505
R24797 VSS.n2738 VSS.n2737 0.4505
R24798 VSS.n3955 VSS.n3954 0.4505
R24799 VSS.n3956 VSS.n2736 0.4505
R24800 VSS.n3958 VSS.n3957 0.4505
R24801 VSS.n2734 VSS.n2733 0.4505
R24802 VSS.n3963 VSS.n3962 0.4505
R24803 VSS.n3964 VSS.n2732 0.4505
R24804 VSS.n3966 VSS.n3965 0.4505
R24805 VSS.n2730 VSS.n2729 0.4505
R24806 VSS.n3971 VSS.n3970 0.4505
R24807 VSS.n3972 VSS.n2728 0.4505
R24808 VSS.n3974 VSS.n3973 0.4505
R24809 VSS.n2726 VSS.n2725 0.4505
R24810 VSS.n3979 VSS.n3978 0.4505
R24811 VSS.n3980 VSS.n2724 0.4505
R24812 VSS.n3982 VSS.n3981 0.4505
R24813 VSS.n2722 VSS.n2721 0.4505
R24814 VSS.n3987 VSS.n3986 0.4505
R24815 VSS.n3988 VSS.n2720 0.4505
R24816 VSS.n3990 VSS.n3989 0.4505
R24817 VSS.n2718 VSS.n2717 0.4505
R24818 VSS.n3995 VSS.n3994 0.4505
R24819 VSS.n3996 VSS.n2716 0.4505
R24820 VSS.n3998 VSS.n3997 0.4505
R24821 VSS.n2714 VSS.n2713 0.4505
R24822 VSS.n4003 VSS.n4002 0.4505
R24823 VSS.n4004 VSS.n2712 0.4505
R24824 VSS.n4006 VSS.n4005 0.4505
R24825 VSS.n2710 VSS.n2709 0.4505
R24826 VSS.n4011 VSS.n4010 0.4505
R24827 VSS.n4012 VSS.n2708 0.4505
R24828 VSS.n4014 VSS.n4013 0.4505
R24829 VSS.n2706 VSS.n2705 0.4505
R24830 VSS.n4020 VSS.n4019 0.4505
R24831 VSS.n4021 VSS.n2704 0.4505
R24832 VSS.n4023 VSS.n4022 0.4505
R24833 VSS.n4024 VSS.n3 0.4505
R24834 VSS.n5709 VSS.n5708 0.4505
R24835 VSS.n5707 VSS.n2 0.4505
R24836 VSS.n5706 VSS.n5705 0.4505
R24837 VSS.n5407 DVSS 0.449176
R24838 VSS.n5312 DVSS 0.449176
R24839 VSS.n5312 DVSS 0.449176
R24840 VSS.n5243 VSS.n5242 0.441235
R24841 VSS.n5682 VSS.n5681 0.439524
R24842 VSS.n1590 VSS.n1170 0.439458
R24843 VSS.n5316 VSS.n2127 0.420329
R24844 VSS.n3869 VSS.n2095 0.41962
R24845 VSS.n3410 VSS.n3409 0.4165
R24846 VSS.n3415 VSS.n3414 0.4165
R24847 VSS.n3408 VSS.n3393 0.412794
R24848 VSS.n2890 VSS.n2889 0.409053
R24849 VSS.n3403 VSS.n3400 0.409053
R24850 VSS.n3731 VSS.n3730 0.40882
R24851 VSS.n4144 DVSS 0.402853
R24852 VSS.n5248 DVSS 0.402853
R24853 VSS.n4246 DVSS 0.402853
R24854 DVSS VSS.n4242 0.402853
R24855 VSS.n3311 VSS.n3310 0.388068
R24856 VSS.n3071 VSS.n3059 0.387662
R24857 VSS.n5407 DVSS 0.384324
R24858 VSS.n3732 VSS.n3731 0.382451
R24859 VSS.n4284 VSS.n2295 0.375755
R24860 VSS.n3058 VSS.n3057 0.3755
R24861 VSS.n3309 VSS.n2972 0.3755
R24862 VSS.n3875 VSS.n3874 0.3755
R24863 VSS.n4145 VSS.n2428 0.368789
R24864 VSS.n4144 VSS.n2429 0.368789
R24865 VSS.n4143 VSS.n2431 0.368789
R24866 VSS.n4141 VSS.n4140 0.368789
R24867 VSS.n5248 VSS.n2241 0.368789
R24868 VSS.n5247 VSS.n5246 0.368789
R24869 VSS.n4202 VSS.n2355 0.368789
R24870 VSS.n4246 VSS.n2356 0.368789
R24871 VSS.n4245 VSS.n2357 0.368789
R24872 VSS.n4243 VSS.n2359 0.368789
R24873 VSS.n4242 VSS.n2360 0.368789
R24874 VSS.n4241 VSS.n4240 0.368789
R24875 VSS.n5271 VSS.n2218 0.367935
R24876 VSS.n5271 VSS.n5268 0.367935
R24877 VSS.n2233 VSS.n2205 0.367935
R24878 VSS.n2219 VSS.n2205 0.367935
R24879 VSS.n2234 VSS.n2206 0.367935
R24880 VSS.n2220 VSS.n2206 0.367935
R24881 VSS.n2235 VSS.n2207 0.367935
R24882 VSS.n2221 VSS.n2207 0.367935
R24883 VSS.n2236 VSS.n2208 0.367935
R24884 VSS.n2222 VSS.n2208 0.367935
R24885 VSS.n5257 VSS.n5256 0.367935
R24886 VSS.n2231 VSS.n2209 0.367935
R24887 VSS.n2222 VSS.n2210 0.367935
R24888 VSS.n2221 VSS.n2211 0.367935
R24889 VSS.n2220 VSS.n2212 0.367935
R24890 VSS.n2219 VSS.n2213 0.367935
R24891 VSS.n5268 VSS.n2214 0.367935
R24892 VSS.n5256 VSS.n2210 0.367935
R24893 VSS.n2236 VSS.n2211 0.367935
R24894 VSS.n2235 VSS.n2212 0.367935
R24895 VSS.n2234 VSS.n2213 0.367935
R24896 VSS.n2233 VSS.n2214 0.367935
R24897 VSS.n5274 VSS.n2218 0.367935
R24898 VSS.n5257 VSS.n2209 0.367935
R24899 VSS.n2363 VSS.n2362 0.36232
R24900 VSS.n2365 VSS.n2364 0.36232
R24901 VSS.n3532 DVSS 0.358788
R24902 VSS.n3729 VSS.n2818 0.346654
R24903 VSS.n3729 VSS.n3728 0.346654
R24904 VSS.n5309 VSS.n2134 0.342906
R24905 VSS.n2370 VSS.n2369 0.335984
R24906 VSS.n1773 VSS.n1772 0.328381
R24907 VSS.n1786 VSS.n1774 0.328381
R24908 VSS.n1916 VSS.n1726 0.328381
R24909 VSS.n1903 VSS.n1902 0.328381
R24910 VSS.n1954 VSS.n1702 0.328381
R24911 VSS.n1941 VSS.n1940 0.328381
R24912 VSS.n1988 VSS.n1676 0.328381
R24913 VSS.n1975 VSS.n1974 0.328381
R24914 VSS.n2020 VSS.n1649 0.328381
R24915 VSS.n2007 VSS.n2006 0.328381
R24916 VSS.n1629 VSS.n1628 0.328381
R24917 VSS.n1642 VSS.n1630 0.328381
R24918 VSS.n3030 VSS.n3029 0.311888
R24919 VSS.n3259 VSS.n3258 0.311888
R24920 VSS.n2368 VSS.n2367 0.309579
R24921 VSS.n2295 VSS.n2294 0.309579
R24922 VSS.n4287 VSS.n4286 0.309579
R24923 VSS.n4290 VSS.n4289 0.309579
R24924 VSS.n2369 VSS.n2295 0.307559
R24925 VSS.n5392 VSS.n5391 0.297643
R24926 VSS.n5335 VSS.n5334 0.297643
R24927 VSS.n5428 VSS.n5427 0.297643
R24928 VSS.n2801 VSS.n2100 0.297643
R24929 VSS.n1006 VSS.n1005 0.28175
R24930 VSS.n523 VSS.n375 0.28175
R24931 DVSS VSS.n2227 0.273784
R24932 VSS.n3506 VSS.n3505 0.273147
R24933 VSS.n3417 VSS.n3397 0.273147
R24934 VSS.n5323 VSS.n2127 0.271399
R24935 VSS.n5417 VSS.n2095 0.271321
R24936 VSS.n4092 VSS.n4091 0.268132
R24937 VSS.n5330 VSS.n2173 0.266421
R24938 VSS.n265 VSS.n222 0.265206
R24939 VSS.n381 VSS.n380 0.265206
R24940 VSS.n5400 VSS.n2107 0.265206
R24941 VSS.n5400 VSS.n5399 0.265206
R24942 VSS.n5376 VSS.n2127 0.264882
R24943 VSS.n3745 VSS.n2095 0.264797
R24944 VSS.n5331 VSS.n5330 0.2605
R24945 VSS.n5402 VSS.n5401 0.2605
R24946 VSS.n5434 VSS.n5433 0.2605
R24947 VSS.n2789 VSS 0.258658
R24948 VSS.n5283 VSS.n2199 0.254359
R24949 VSS.n5300 VSS.n5298 0.249324
R24950 VSS.n5296 VSS.n5295 0.249324
R24951 VSS.n4049 VSS.n4048 0.249324
R24952 VSS.n2369 VSS.n2368 0.238735
R24953 VSS.n3057 VSS.n3056 0.231484
R24954 VSS.n3260 VSS.n2972 0.231484
R24955 VSS.n3439 VSS.n3436 0.231338
R24956 VSS.n5706 VSS.n4 0.231338
R24957 VSS.n2314 VSS.n2309 0.231338
R24958 VSS.n2693 VSS.n2686 0.231338
R24959 VSS.n1835 VSS.n1829 0.231338
R24960 VSS.n3057 VSS.n2971 0.229569
R24961 VSS VSS.n5297 0.229471
R24962 VSS.n5297 VSS 0.229471
R24963 VSS.n3313 VSS.n2972 0.228851
R24964 VSS.n2789 VSS.n2788 0.224316
R24965 VSS.n1080 VSS.n1079 0.219756
R24966 VSS.n2168 VSS.n2167 0.219756
R24967 VSS.n1029 VSS.n37 0.217409
R24968 VSS.n1138 VSS.n1137 0.217409
R24969 VSS.n170 VSS.n95 0.214786
R24970 VSS.n581 VSS.n366 0.214786
R24971 VSS.n2170 VSS.n2166 0.214786
R24972 VSS.n2165 VSS.n2162 0.214786
R24973 VSS.n5342 VSS.n2161 0.214786
R24974 VSS.n5343 VSS.n2160 0.214786
R24975 VSS.n5344 VSS.n2159 0.214786
R24976 VSS.n2158 VSS.n2156 0.214786
R24977 VSS.n5348 VSS.n2155 0.214786
R24978 VSS.n5349 VSS.n2154 0.214786
R24979 VSS.n5350 VSS.n2153 0.214786
R24980 VSS.n2152 VSS.n2150 0.214786
R24981 VSS.n5354 VSS.n2149 0.214786
R24982 VSS.n5355 VSS.n2148 0.214786
R24983 VSS.n5356 VSS.n2147 0.214786
R24984 VSS.n2146 VSS.n2144 0.214786
R24985 VSS.n5360 VSS.n2143 0.214786
R24986 VSS.n5361 VSS.n2142 0.214786
R24987 VSS.n5362 VSS.n2141 0.214786
R24988 VSS.n2140 VSS.n2138 0.214786
R24989 VSS.n5366 VSS.n2137 0.214786
R24990 VSS.n5367 VSS.n2136 0.214786
R24991 VSS.n2135 VSS.n2133 0.214786
R24992 VSS.n5371 VSS.n2132 0.214786
R24993 VSS.n5372 VSS.n2131 0.214786
R24994 VSS.n5373 VSS.n2130 0.214786
R24995 VSS.n2129 VSS.n2126 0.214786
R24996 VSS.n5378 VSS.n2125 0.214786
R24997 VSS.n5379 VSS.n2124 0.214786
R24998 VSS.n5380 VSS.n2123 0.214786
R24999 VSS.n2122 VSS.n2120 0.214786
R25000 VSS.n5384 VSS.n2119 0.214786
R25001 VSS.n5385 VSS.n2118 0.214786
R25002 VSS.n3735 VSS.n3734 0.214786
R25003 VSS.n2814 VSS.n2813 0.214786
R25004 VSS.n3740 VSS.n3739 0.214786
R25005 VSS.n3741 VSS.n2812 0.214786
R25006 VSS.n3743 VSS.n3742 0.214786
R25007 VSS.n2810 VSS.n2809 0.214786
R25008 VSS.n3749 VSS.n3748 0.214786
R25009 VSS.n3750 VSS.n2808 0.214786
R25010 VSS.n3752 VSS.n3751 0.214786
R25011 VSS.n2806 VSS.n2805 0.214786
R25012 VSS.n3757 VSS.n3756 0.214786
R25013 VSS.n3758 VSS.n2804 0.214786
R25014 VSS.n3863 VSS.n3759 0.214786
R25015 VSS.n3862 VSS.n3760 0.214786
R25016 VSS.n3861 VSS.n3761 0.214786
R25017 VSS.n3764 VSS.n3762 0.214786
R25018 VSS.n3857 VSS.n3765 0.214786
R25019 VSS.n3856 VSS.n3766 0.214786
R25020 VSS.n3855 VSS.n3767 0.214786
R25021 VSS.n3770 VSS.n3768 0.214786
R25022 VSS.n3851 VSS.n3771 0.214786
R25023 VSS.n3850 VSS.n3772 0.214786
R25024 VSS.n3849 VSS.n3773 0.214786
R25025 VSS.n3777 VSS.n3774 0.214786
R25026 VSS.n3845 VSS.n3778 0.214786
R25027 VSS.n3844 VSS.n3779 0.214786
R25028 VSS.n3843 VSS.n3780 0.214786
R25029 VSS.n3783 VSS.n3781 0.214786
R25030 VSS.n3839 VSS.n3784 0.214786
R25031 VSS.n3838 VSS.n3785 0.214786
R25032 VSS.n3837 VSS.n3786 0.214786
R25033 VSS.n3789 VSS.n3787 0.214786
R25034 VSS.n3833 VSS.n3790 0.214786
R25035 VSS.n3832 VSS.n3791 0.214786
R25036 VSS.n3831 VSS.n3792 0.214786
R25037 VSS.n3795 VSS.n3793 0.214786
R25038 VSS.n3827 VSS.n3796 0.214786
R25039 VSS.n3826 VSS.n3797 0.214786
R25040 VSS.n3825 VSS.n3798 0.214786
R25041 VSS.n3801 VSS.n3799 0.214786
R25042 VSS.n3821 VSS.n3802 0.214786
R25043 VSS.n3820 VSS.n3803 0.214786
R25044 VSS.n3819 VSS.n3804 0.214786
R25045 VSS.n3807 VSS.n3805 0.214786
R25046 VSS.n3815 VSS.n3808 0.214786
R25047 VSS.n3814 VSS.n3809 0.214786
R25048 VSS.n3813 VSS.n3811 0.214786
R25049 VSS.n3810 VSS.n2116 0.214786
R25050 VSS.n5386 VSS.n2117 0.214786
R25051 VSS.n1031 VSS.n1028 0.214786
R25052 VSS.n1027 VSS.n1026 0.214786
R25053 VSS.n1035 VSS.n1025 0.214786
R25054 VSS.n1036 VSS.n1024 0.214786
R25055 VSS.n1023 VSS.n1022 0.214786
R25056 VSS.n1040 VSS.n1021 0.214786
R25057 VSS.n1041 VSS.n1020 0.214786
R25058 VSS.n1042 VSS.n1019 0.214786
R25059 VSS.n1018 VSS.n1016 0.214786
R25060 VSS.n1046 VSS.n1015 0.214786
R25061 VSS.n1047 VSS.n1014 0.214786
R25062 VSS.n1048 VSS.n1013 0.214786
R25063 VSS.n1011 VSS.n1010 0.214786
R25064 VSS.n1053 VSS.n1052 0.214786
R25065 VSS.n1009 VSS.n1008 0.214786
R25066 VSS.n102 VSS.n101 0.214786
R25067 VSS.n1001 VSS.n1000 0.214786
R25068 VSS.n999 VSS.n107 0.214786
R25069 VSS.n998 VSS.n997 0.214786
R25070 VSS.n109 VSS.n108 0.214786
R25071 VSS.n993 VSS.n992 0.214786
R25072 VSS.n991 VSS.n111 0.214786
R25073 VSS.n990 VSS.n989 0.214786
R25074 VSS.n113 VSS.n112 0.214786
R25075 VSS.n985 VSS.n984 0.214786
R25076 VSS.n983 VSS.n115 0.214786
R25077 VSS.n982 VSS.n981 0.214786
R25078 VSS.n117 VSS.n116 0.214786
R25079 VSS.n977 VSS.n976 0.214786
R25080 VSS.n975 VSS.n119 0.214786
R25081 VSS.n974 VSS.n973 0.214786
R25082 VSS.n121 VSS.n120 0.214786
R25083 VSS.n969 VSS.n968 0.214786
R25084 VSS.n967 VSS.n123 0.214786
R25085 VSS.n966 VSS.n965 0.214786
R25086 VSS.n125 VSS.n124 0.214786
R25087 VSS.n960 VSS.n959 0.214786
R25088 VSS.n958 VSS.n127 0.214786
R25089 VSS.n956 VSS.n955 0.214786
R25090 VSS.n130 VSS.n129 0.214786
R25091 VSS.n456 VSS.n455 0.214786
R25092 VSS.n459 VSS.n454 0.214786
R25093 VSS.n460 VSS.n453 0.214786
R25094 VSS.n461 VSS.n452 0.214786
R25095 VSS.n451 VSS.n449 0.214786
R25096 VSS.n465 VSS.n448 0.214786
R25097 VSS.n466 VSS.n447 0.214786
R25098 VSS.n467 VSS.n446 0.214786
R25099 VSS.n445 VSS.n443 0.214786
R25100 VSS.n471 VSS.n442 0.214786
R25101 VSS.n472 VSS.n441 0.214786
R25102 VSS.n473 VSS.n440 0.214786
R25103 VSS.n439 VSS.n437 0.214786
R25104 VSS.n477 VSS.n436 0.214786
R25105 VSS.n478 VSS.n435 0.214786
R25106 VSS.n479 VSS.n434 0.214786
R25107 VSS.n433 VSS.n431 0.214786
R25108 VSS.n483 VSS.n430 0.214786
R25109 VSS.n484 VSS.n429 0.214786
R25110 VSS.n485 VSS.n428 0.214786
R25111 VSS.n427 VSS.n424 0.214786
R25112 VSS.n489 VSS.n423 0.214786
R25113 VSS.n491 VSS.n422 0.214786
R25114 VSS.n492 VSS.n421 0.214786
R25115 VSS.n420 VSS.n418 0.214786
R25116 VSS.n496 VSS.n417 0.214786
R25117 VSS.n497 VSS.n416 0.214786
R25118 VSS.n415 VSS.n414 0.214786
R25119 VSS.n501 VSS.n413 0.214786
R25120 VSS.n502 VSS.n412 0.214786
R25121 VSS.n503 VSS.n411 0.214786
R25122 VSS.n410 VSS.n408 0.214786
R25123 VSS.n507 VSS.n407 0.214786
R25124 VSS.n508 VSS.n406 0.214786
R25125 VSS.n509 VSS.n405 0.214786
R25126 VSS.n404 VSS.n402 0.214786
R25127 VSS.n513 VSS.n401 0.214786
R25128 VSS.n514 VSS.n400 0.214786
R25129 VSS.n515 VSS.n399 0.214786
R25130 VSS.n398 VSS.n396 0.214786
R25131 VSS.n519 VSS.n395 0.214786
R25132 VSS.n520 VSS.n394 0.214786
R25133 VSS.n521 VSS.n393 0.214786
R25134 VSS.n392 VSS.n390 0.214786
R25135 VSS.n576 VSS.n388 0.214786
R25136 VSS.n575 VSS.n389 0.214786
R25137 VSS.n1136 VSS.n1135 0.214786
R25138 VSS.n80 VSS.n79 0.214786
R25139 VSS.n1131 VSS.n1130 0.214786
R25140 VSS.n1129 VSS.n82 0.214786
R25141 VSS.n1128 VSS.n1127 0.214786
R25142 VSS.n84 VSS.n83 0.214786
R25143 VSS.n1123 VSS.n1122 0.214786
R25144 VSS.n1121 VSS.n86 0.214786
R25145 VSS.n1120 VSS.n1119 0.214786
R25146 VSS.n88 VSS.n87 0.214786
R25147 VSS.n1115 VSS.n1114 0.214786
R25148 VSS.n1113 VSS.n90 0.214786
R25149 VSS.n1112 VSS.n1111 0.214786
R25150 VSS.n92 VSS.n91 0.214786
R25151 VSS.n1106 VSS.n97 0.214786
R25152 VSS.n168 VSS.n96 0.214786
R25153 VSS.n919 VSS.n169 0.214786
R25154 VSS.n920 VSS.n167 0.214786
R25155 VSS.n921 VSS.n166 0.214786
R25156 VSS.n165 VSS.n163 0.214786
R25157 VSS.n925 VSS.n162 0.214786
R25158 VSS.n926 VSS.n161 0.214786
R25159 VSS.n927 VSS.n160 0.214786
R25160 VSS.n159 VSS.n157 0.214786
R25161 VSS.n931 VSS.n156 0.214786
R25162 VSS.n932 VSS.n155 0.214786
R25163 VSS.n933 VSS.n154 0.214786
R25164 VSS.n153 VSS.n151 0.214786
R25165 VSS.n937 VSS.n150 0.214786
R25166 VSS.n938 VSS.n149 0.214786
R25167 VSS.n939 VSS.n148 0.214786
R25168 VSS.n147 VSS.n145 0.214786
R25169 VSS.n943 VSS.n144 0.214786
R25170 VSS.n944 VSS.n143 0.214786
R25171 VSS.n142 VSS.n140 0.214786
R25172 VSS.n948 VSS.n139 0.214786
R25173 VSS.n949 VSS.n138 0.214786
R25174 VSS.n950 VSS.n137 0.214786
R25175 VSS.n805 VSS.n804 0.214786
R25176 VSS.n807 VSS.n803 0.214786
R25177 VSS.n808 VSS.n802 0.214786
R25178 VSS.n809 VSS.n801 0.214786
R25179 VSS.n800 VSS.n798 0.214786
R25180 VSS.n813 VSS.n797 0.214786
R25181 VSS.n814 VSS.n796 0.214786
R25182 VSS.n815 VSS.n795 0.214786
R25183 VSS.n794 VSS.n792 0.214786
R25184 VSS.n819 VSS.n791 0.214786
R25185 VSS.n820 VSS.n790 0.214786
R25186 VSS.n821 VSS.n789 0.214786
R25187 VSS.n788 VSS.n308 0.214786
R25188 VSS.n787 VSS.n786 0.214786
R25189 VSS.n310 VSS.n309 0.214786
R25190 VSS.n782 VSS.n781 0.214786
R25191 VSS.n780 VSS.n312 0.214786
R25192 VSS.n779 VSS.n778 0.214786
R25193 VSS.n314 VSS.n313 0.214786
R25194 VSS.n774 VSS.n773 0.214786
R25195 VSS.n772 VSS.n316 0.214786
R25196 VSS.n771 VSS.n770 0.214786
R25197 VSS.n318 VSS.n317 0.214786
R25198 VSS.n766 VSS.n765 0.214786
R25199 VSS.n763 VSS.n762 0.214786
R25200 VSS.n324 VSS.n323 0.214786
R25201 VSS.n758 VSS.n757 0.214786
R25202 VSS.n756 VSS.n326 0.214786
R25203 VSS.n755 VSS.n754 0.214786
R25204 VSS.n328 VSS.n327 0.214786
R25205 VSS.n608 VSS.n606 0.214786
R25206 VSS.n609 VSS.n605 0.214786
R25207 VSS.n610 VSS.n604 0.214786
R25208 VSS.n603 VSS.n601 0.214786
R25209 VSS.n614 VSS.n600 0.214786
R25210 VSS.n615 VSS.n599 0.214786
R25211 VSS.n616 VSS.n598 0.214786
R25212 VSS.n597 VSS.n595 0.214786
R25213 VSS.n620 VSS.n594 0.214786
R25214 VSS.n621 VSS.n593 0.214786
R25215 VSS.n622 VSS.n592 0.214786
R25216 VSS.n591 VSS.n589 0.214786
R25217 VSS.n626 VSS.n588 0.214786
R25218 VSS.n627 VSS.n587 0.214786
R25219 VSS.n628 VSS.n586 0.214786
R25220 VSS.n585 VSS.n369 0.214786
R25221 VSS.n584 VSS.n583 0.214786
R25222 VSS.n371 VSS.n370 0.214786
R25223 VSS.n1082 VSS.n1077 0.214786
R25224 VSS.n1076 VSS.n1074 0.214786
R25225 VSS.n1086 VSS.n1073 0.214786
R25226 VSS.n1087 VSS.n1072 0.214786
R25227 VSS.n1071 VSS.n1070 0.214786
R25228 VSS.n1091 VSS.n1069 0.214786
R25229 VSS.n1092 VSS.n1068 0.214786
R25230 VSS.n1093 VSS.n1067 0.214786
R25231 VSS.n1066 VSS.n1064 0.214786
R25232 VSS.n1097 VSS.n1063 0.214786
R25233 VSS.n1098 VSS.n1062 0.214786
R25234 VSS.n1099 VSS.n1061 0.214786
R25235 VSS.n1060 VSS.n1058 0.214786
R25236 VSS.n1103 VSS.n1057 0.214786
R25237 VSS.n100 VSS.n99 0.214786
R25238 VSS.n898 VSS.n897 0.214786
R25239 VSS.n899 VSS.n896 0.214786
R25240 VSS.n895 VSS.n267 0.214786
R25241 VSS.n894 VSS.n893 0.214786
R25242 VSS.n269 VSS.n268 0.214786
R25243 VSS.n889 VSS.n888 0.214786
R25244 VSS.n887 VSS.n271 0.214786
R25245 VSS.n886 VSS.n885 0.214786
R25246 VSS.n273 VSS.n272 0.214786
R25247 VSS.n881 VSS.n880 0.214786
R25248 VSS.n879 VSS.n275 0.214786
R25249 VSS.n878 VSS.n877 0.214786
R25250 VSS.n277 VSS.n276 0.214786
R25251 VSS.n873 VSS.n872 0.214786
R25252 VSS.n871 VSS.n279 0.214786
R25253 VSS.n870 VSS.n869 0.214786
R25254 VSS.n281 VSS.n280 0.214786
R25255 VSS.n865 VSS.n864 0.214786
R25256 VSS.n863 VSS.n284 0.214786
R25257 VSS.n862 VSS.n861 0.214786
R25258 VSS.n286 VSS.n285 0.214786
R25259 VSS.n856 VSS.n855 0.214786
R25260 VSS.n854 VSS.n288 0.214786
R25261 VSS.n852 VSS.n851 0.214786
R25262 VSS.n290 VSS.n289 0.214786
R25263 VSS.n847 VSS.n846 0.214786
R25264 VSS.n845 VSS.n293 0.214786
R25265 VSS.n844 VSS.n843 0.214786
R25266 VSS.n295 VSS.n294 0.214786
R25267 VSS.n839 VSS.n838 0.214786
R25268 VSS.n837 VSS.n297 0.214786
R25269 VSS.n836 VSS.n835 0.214786
R25270 VSS.n299 VSS.n298 0.214786
R25271 VSS.n831 VSS.n830 0.214786
R25272 VSS.n829 VSS.n301 0.214786
R25273 VSS.n828 VSS.n827 0.214786
R25274 VSS.n303 VSS.n302 0.214786
R25275 VSS.n728 VSS.n727 0.214786
R25276 VSS.n729 VSS.n726 0.214786
R25277 VSS.n725 VSS.n723 0.214786
R25278 VSS.n733 VSS.n722 0.214786
R25279 VSS.n734 VSS.n721 0.214786
R25280 VSS.n735 VSS.n720 0.214786
R25281 VSS.n719 VSS.n717 0.214786
R25282 VSS.n739 VSS.n716 0.214786
R25283 VSS.n740 VSS.n715 0.214786
R25284 VSS.n741 VSS.n714 0.214786
R25285 VSS.n711 VSS.n710 0.214786
R25286 VSS.n746 VSS.n709 0.214786
R25287 VSS.n747 VSS.n708 0.214786
R25288 VSS.n748 VSS.n707 0.214786
R25289 VSS.n706 VSS.n333 0.214786
R25290 VSS.n705 VSS.n704 0.214786
R25291 VSS.n335 VSS.n334 0.214786
R25292 VSS.n700 VSS.n699 0.214786
R25293 VSS.n698 VSS.n337 0.214786
R25294 VSS.n697 VSS.n696 0.214786
R25295 VSS.n339 VSS.n338 0.214786
R25296 VSS.n692 VSS.n691 0.214786
R25297 VSS.n690 VSS.n341 0.214786
R25298 VSS.n689 VSS.n688 0.214786
R25299 VSS.n343 VSS.n342 0.214786
R25300 VSS.n684 VSS.n683 0.214786
R25301 VSS.n682 VSS.n345 0.214786
R25302 VSS.n681 VSS.n680 0.214786
R25303 VSS.n347 VSS.n346 0.214786
R25304 VSS.n676 VSS.n675 0.214786
R25305 VSS.n674 VSS.n349 0.214786
R25306 VSS.n673 VSS.n672 0.214786
R25307 VSS.n351 VSS.n350 0.214786
R25308 VSS.n384 VSS.n383 0.214786
R25309 VSS.n333 VSS.n331 0.214786
R25310 VSS.n1081 VSS.n1075 0.214786
R25311 VSS.n1083 VSS.n1082 0.214786
R25312 VSS.n1084 VSS.n1074 0.214786
R25313 VSS.n1086 VSS.n1085 0.214786
R25314 VSS.n1088 VSS.n1087 0.214786
R25315 VSS.n1089 VSS.n1070 0.214786
R25316 VSS.n1091 VSS.n1090 0.214786
R25317 VSS.n1092 VSS.n1065 0.214786
R25318 VSS.n1094 VSS.n1093 0.214786
R25319 VSS.n1095 VSS.n1064 0.214786
R25320 VSS.n1097 VSS.n1096 0.214786
R25321 VSS.n1098 VSS.n1059 0.214786
R25322 VSS.n1100 VSS.n1099 0.214786
R25323 VSS.n1101 VSS.n1058 0.214786
R25324 VSS.n1103 VSS.n1102 0.214786
R25325 VSS.n264 VSS.n99 0.214786
R25326 VSS.n898 VSS.n266 0.214786
R25327 VSS.n900 VSS.n899 0.214786
R25328 VSS.n267 VSS.n263 0.214786
R25329 VSS.n893 VSS.n892 0.214786
R25330 VSS.n891 VSS.n269 0.214786
R25331 VSS.n890 VSS.n889 0.214786
R25332 VSS.n271 VSS.n270 0.214786
R25333 VSS.n885 VSS.n884 0.214786
R25334 VSS.n883 VSS.n273 0.214786
R25335 VSS.n882 VSS.n881 0.214786
R25336 VSS.n275 VSS.n274 0.214786
R25337 VSS.n877 VSS.n876 0.214786
R25338 VSS.n875 VSS.n277 0.214786
R25339 VSS.n874 VSS.n873 0.214786
R25340 VSS.n279 VSS.n278 0.214786
R25341 VSS.n869 VSS.n868 0.214786
R25342 VSS.n867 VSS.n281 0.214786
R25343 VSS.n866 VSS.n865 0.214786
R25344 VSS.n859 VSS.n284 0.214786
R25345 VSS.n861 VSS.n860 0.214786
R25346 VSS.n858 VSS.n286 0.214786
R25347 VSS.n857 VSS.n856 0.214786
R25348 VSS.n288 VSS.n287 0.214786
R25349 VSS.n851 VSS.n850 0.214786
R25350 VSS.n849 VSS.n290 0.214786
R25351 VSS.n848 VSS.n847 0.214786
R25352 VSS.n293 VSS.n292 0.214786
R25353 VSS.n843 VSS.n842 0.214786
R25354 VSS.n841 VSS.n295 0.214786
R25355 VSS.n840 VSS.n839 0.214786
R25356 VSS.n297 VSS.n296 0.214786
R25357 VSS.n835 VSS.n834 0.214786
R25358 VSS.n833 VSS.n299 0.214786
R25359 VSS.n832 VSS.n831 0.214786
R25360 VSS.n301 VSS.n300 0.214786
R25361 VSS.n827 VSS.n826 0.214786
R25362 VSS.n304 VSS.n303 0.214786
R25363 VSS.n728 VSS.n724 0.214786
R25364 VSS.n730 VSS.n729 0.214786
R25365 VSS.n731 VSS.n723 0.214786
R25366 VSS.n733 VSS.n732 0.214786
R25367 VSS.n734 VSS.n718 0.214786
R25368 VSS.n736 VSS.n735 0.214786
R25369 VSS.n737 VSS.n717 0.214786
R25370 VSS.n739 VSS.n738 0.214786
R25371 VSS.n740 VSS.n712 0.214786
R25372 VSS.n742 VSS.n741 0.214786
R25373 VSS.n744 VSS.n711 0.214786
R25374 VSS.n746 VSS.n745 0.214786
R25375 VSS.n747 VSS.n332 0.214786
R25376 VSS.n749 VSS.n748 0.214786
R25377 VSS.n704 VSS.n703 0.214786
R25378 VSS.n702 VSS.n335 0.214786
R25379 VSS.n701 VSS.n700 0.214786
R25380 VSS.n337 VSS.n336 0.214786
R25381 VSS.n696 VSS.n695 0.214786
R25382 VSS.n694 VSS.n339 0.214786
R25383 VSS.n693 VSS.n692 0.214786
R25384 VSS.n341 VSS.n340 0.214786
R25385 VSS.n688 VSS.n687 0.214786
R25386 VSS.n686 VSS.n343 0.214786
R25387 VSS.n685 VSS.n684 0.214786
R25388 VSS.n345 VSS.n344 0.214786
R25389 VSS.n680 VSS.n679 0.214786
R25390 VSS.n678 VSS.n347 0.214786
R25391 VSS.n677 VSS.n676 0.214786
R25392 VSS.n349 VSS.n348 0.214786
R25393 VSS.n672 VSS.n671 0.214786
R25394 VSS.n352 VSS.n351 0.214786
R25395 VSS.n383 VSS.n382 0.214786
R25396 VSS.n78 VSS.n57 0.214786
R25397 VSS.n1135 VSS.n1134 0.214786
R25398 VSS.n1133 VSS.n80 0.214786
R25399 VSS.n1132 VSS.n1131 0.214786
R25400 VSS.n82 VSS.n81 0.214786
R25401 VSS.n1127 VSS.n1126 0.214786
R25402 VSS.n1125 VSS.n84 0.214786
R25403 VSS.n1124 VSS.n1123 0.214786
R25404 VSS.n86 VSS.n85 0.214786
R25405 VSS.n1119 VSS.n1118 0.214786
R25406 VSS.n1117 VSS.n88 0.214786
R25407 VSS.n1116 VSS.n1115 0.214786
R25408 VSS.n90 VSS.n89 0.214786
R25409 VSS.n1111 VSS.n1110 0.214786
R25410 VSS.n1109 VSS.n92 0.214786
R25411 VSS.n1107 VSS.n1106 0.214786
R25412 VSS.n917 VSS.n96 0.214786
R25413 VSS.n919 VSS.n918 0.214786
R25414 VSS.n920 VSS.n164 0.214786
R25415 VSS.n922 VSS.n921 0.214786
R25416 VSS.n923 VSS.n163 0.214786
R25417 VSS.n925 VSS.n924 0.214786
R25418 VSS.n926 VSS.n158 0.214786
R25419 VSS.n928 VSS.n927 0.214786
R25420 VSS.n929 VSS.n157 0.214786
R25421 VSS.n931 VSS.n930 0.214786
R25422 VSS.n932 VSS.n152 0.214786
R25423 VSS.n934 VSS.n933 0.214786
R25424 VSS.n935 VSS.n151 0.214786
R25425 VSS.n937 VSS.n936 0.214786
R25426 VSS.n938 VSS.n146 0.214786
R25427 VSS.n940 VSS.n939 0.214786
R25428 VSS.n941 VSS.n145 0.214786
R25429 VSS.n943 VSS.n942 0.214786
R25430 VSS.n945 VSS.n944 0.214786
R25431 VSS.n946 VSS.n140 0.214786
R25432 VSS.n948 VSS.n947 0.214786
R25433 VSS.n949 VSS.n135 0.214786
R25434 VSS.n951 VSS.n950 0.214786
R25435 VSS.n805 VSS.n134 0.214786
R25436 VSS.n807 VSS.n806 0.214786
R25437 VSS.n808 VSS.n799 0.214786
R25438 VSS.n810 VSS.n809 0.214786
R25439 VSS.n811 VSS.n798 0.214786
R25440 VSS.n813 VSS.n812 0.214786
R25441 VSS.n814 VSS.n793 0.214786
R25442 VSS.n816 VSS.n815 0.214786
R25443 VSS.n817 VSS.n792 0.214786
R25444 VSS.n819 VSS.n818 0.214786
R25445 VSS.n820 VSS.n307 0.214786
R25446 VSS.n822 VSS.n821 0.214786
R25447 VSS.n308 VSS.n306 0.214786
R25448 VSS.n786 VSS.n785 0.214786
R25449 VSS.n784 VSS.n310 0.214786
R25450 VSS.n783 VSS.n782 0.214786
R25451 VSS.n312 VSS.n311 0.214786
R25452 VSS.n778 VSS.n777 0.214786
R25453 VSS.n776 VSS.n314 0.214786
R25454 VSS.n775 VSS.n774 0.214786
R25455 VSS.n316 VSS.n315 0.214786
R25456 VSS.n770 VSS.n769 0.214786
R25457 VSS.n768 VSS.n318 0.214786
R25458 VSS.n767 VSS.n766 0.214786
R25459 VSS.n762 VSS.n761 0.214786
R25460 VSS.n760 VSS.n324 0.214786
R25461 VSS.n759 VSS.n758 0.214786
R25462 VSS.n326 VSS.n325 0.214786
R25463 VSS.n754 VSS.n753 0.214786
R25464 VSS.n329 VSS.n328 0.214786
R25465 VSS.n608 VSS.n607 0.214786
R25466 VSS.n609 VSS.n602 0.214786
R25467 VSS.n611 VSS.n610 0.214786
R25468 VSS.n612 VSS.n601 0.214786
R25469 VSS.n614 VSS.n613 0.214786
R25470 VSS.n615 VSS.n596 0.214786
R25471 VSS.n617 VSS.n616 0.214786
R25472 VSS.n618 VSS.n595 0.214786
R25473 VSS.n620 VSS.n619 0.214786
R25474 VSS.n621 VSS.n590 0.214786
R25475 VSS.n623 VSS.n622 0.214786
R25476 VSS.n624 VSS.n589 0.214786
R25477 VSS.n626 VSS.n625 0.214786
R25478 VSS.n627 VSS.n368 0.214786
R25479 VSS.n629 VSS.n628 0.214786
R25480 VSS.n369 VSS.n367 0.214786
R25481 VSS.n583 VSS.n582 0.214786
R25482 VSS.n580 VSS.n371 0.214786
R25483 VSS.n1030 VSS.n36 0.214786
R25484 VSS.n1032 VSS.n1031 0.214786
R25485 VSS.n1033 VSS.n1026 0.214786
R25486 VSS.n1035 VSS.n1034 0.214786
R25487 VSS.n1037 VSS.n1036 0.214786
R25488 VSS.n1038 VSS.n1022 0.214786
R25489 VSS.n1040 VSS.n1039 0.214786
R25490 VSS.n1041 VSS.n1017 0.214786
R25491 VSS.n1043 VSS.n1042 0.214786
R25492 VSS.n1044 VSS.n1016 0.214786
R25493 VSS.n1046 VSS.n1045 0.214786
R25494 VSS.n1047 VSS.n1012 0.214786
R25495 VSS.n1049 VSS.n1048 0.214786
R25496 VSS.n1050 VSS.n1011 0.214786
R25497 VSS.n1052 VSS.n1051 0.214786
R25498 VSS.n1008 VSS.n1007 0.214786
R25499 VSS.n103 VSS.n102 0.214786
R25500 VSS.n1002 VSS.n1001 0.214786
R25501 VSS.n107 VSS.n106 0.214786
R25502 VSS.n997 VSS.n996 0.214786
R25503 VSS.n995 VSS.n109 0.214786
R25504 VSS.n994 VSS.n993 0.214786
R25505 VSS.n111 VSS.n110 0.214786
R25506 VSS.n989 VSS.n988 0.214786
R25507 VSS.n987 VSS.n113 0.214786
R25508 VSS.n986 VSS.n985 0.214786
R25509 VSS.n115 VSS.n114 0.214786
R25510 VSS.n981 VSS.n980 0.214786
R25511 VSS.n979 VSS.n117 0.214786
R25512 VSS.n978 VSS.n977 0.214786
R25513 VSS.n119 VSS.n118 0.214786
R25514 VSS.n973 VSS.n972 0.214786
R25515 VSS.n971 VSS.n121 0.214786
R25516 VSS.n970 VSS.n969 0.214786
R25517 VSS.n963 VSS.n123 0.214786
R25518 VSS.n965 VSS.n964 0.214786
R25519 VSS.n962 VSS.n125 0.214786
R25520 VSS.n961 VSS.n960 0.214786
R25521 VSS.n127 VSS.n126 0.214786
R25522 VSS.n955 VSS.n954 0.214786
R25523 VSS.n132 VSS.n130 0.214786
R25524 VSS.n457 VSS.n456 0.214786
R25525 VSS.n459 VSS.n458 0.214786
R25526 VSS.n460 VSS.n450 0.214786
R25527 VSS.n462 VSS.n461 0.214786
R25528 VSS.n463 VSS.n449 0.214786
R25529 VSS.n465 VSS.n464 0.214786
R25530 VSS.n466 VSS.n444 0.214786
R25531 VSS.n468 VSS.n467 0.214786
R25532 VSS.n469 VSS.n443 0.214786
R25533 VSS.n471 VSS.n470 0.214786
R25534 VSS.n472 VSS.n438 0.214786
R25535 VSS.n474 VSS.n473 0.214786
R25536 VSS.n475 VSS.n437 0.214786
R25537 VSS.n477 VSS.n476 0.214786
R25538 VSS.n478 VSS.n432 0.214786
R25539 VSS.n480 VSS.n479 0.214786
R25540 VSS.n481 VSS.n431 0.214786
R25541 VSS.n483 VSS.n482 0.214786
R25542 VSS.n484 VSS.n426 0.214786
R25543 VSS.n486 VSS.n485 0.214786
R25544 VSS.n487 VSS.n424 0.214786
R25545 VSS.n489 VSS.n488 0.214786
R25546 VSS.n491 VSS.n419 0.214786
R25547 VSS.n493 VSS.n492 0.214786
R25548 VSS.n494 VSS.n418 0.214786
R25549 VSS.n496 VSS.n495 0.214786
R25550 VSS.n498 VSS.n497 0.214786
R25551 VSS.n499 VSS.n414 0.214786
R25552 VSS.n501 VSS.n500 0.214786
R25553 VSS.n502 VSS.n409 0.214786
R25554 VSS.n504 VSS.n503 0.214786
R25555 VSS.n505 VSS.n408 0.214786
R25556 VSS.n507 VSS.n506 0.214786
R25557 VSS.n508 VSS.n403 0.214786
R25558 VSS.n510 VSS.n509 0.214786
R25559 VSS.n511 VSS.n402 0.214786
R25560 VSS.n513 VSS.n512 0.214786
R25561 VSS.n514 VSS.n397 0.214786
R25562 VSS.n516 VSS.n515 0.214786
R25563 VSS.n517 VSS.n396 0.214786
R25564 VSS.n519 VSS.n518 0.214786
R25565 VSS.n520 VSS.n391 0.214786
R25566 VSS.n522 VSS.n521 0.214786
R25567 VSS.n573 VSS.n390 0.214786
R25568 VSS.n577 VSS.n576 0.214786
R25569 VSS.n575 VSS.n574 0.214786
R25570 VSS.n5375 VSS.n2126 0.214786
R25571 VSS.n2169 VSS.n2164 0.214786
R25572 VSS.n2171 VSS.n2170 0.214786
R25573 VSS.n2163 VSS.n2162 0.214786
R25574 VSS.n5342 VSS.n5341 0.214786
R25575 VSS.n5343 VSS.n2157 0.214786
R25576 VSS.n5345 VSS.n5344 0.214786
R25577 VSS.n5346 VSS.n2156 0.214786
R25578 VSS.n5348 VSS.n5347 0.214786
R25579 VSS.n5349 VSS.n2151 0.214786
R25580 VSS.n5351 VSS.n5350 0.214786
R25581 VSS.n5352 VSS.n2150 0.214786
R25582 VSS.n5354 VSS.n5353 0.214786
R25583 VSS.n5355 VSS.n2145 0.214786
R25584 VSS.n5357 VSS.n5356 0.214786
R25585 VSS.n5358 VSS.n2144 0.214786
R25586 VSS.n5360 VSS.n5359 0.214786
R25587 VSS.n5361 VSS.n2139 0.214786
R25588 VSS.n5363 VSS.n5362 0.214786
R25589 VSS.n5364 VSS.n2138 0.214786
R25590 VSS.n5366 VSS.n5365 0.214786
R25591 VSS.n5385 VSS.n2115 0.214786
R25592 VSS.n5384 VSS.n5383 0.214786
R25593 VSS.n5382 VSS.n2120 0.214786
R25594 VSS.n5381 VSS.n5380 0.214786
R25595 VSS.n5379 VSS.n2121 0.214786
R25596 VSS.n5378 VSS.n5377 0.214786
R25597 VSS.n5374 VSS.n5373 0.214786
R25598 VSS.n5372 VSS.n2128 0.214786
R25599 VSS.n5371 VSS.n5370 0.214786
R25600 VSS.n5369 VSS.n2133 0.214786
R25601 VSS.n5368 VSS.n5367 0.214786
R25602 VSS.n2816 VSS.n2815 0.214786
R25603 VSS.n3736 VSS.n3735 0.214786
R25604 VSS.n3737 VSS.n2814 0.214786
R25605 VSS.n3739 VSS.n3738 0.214786
R25606 VSS.n2812 VSS.n2811 0.214786
R25607 VSS.n3744 VSS.n3743 0.214786
R25608 VSS.n3746 VSS.n2810 0.214786
R25609 VSS.n3748 VSS.n3747 0.214786
R25610 VSS.n2808 VSS.n2807 0.214786
R25611 VSS.n3753 VSS.n3752 0.214786
R25612 VSS.n3754 VSS.n2806 0.214786
R25613 VSS.n3756 VSS.n3755 0.214786
R25614 VSS.n2804 VSS.n2802 0.214786
R25615 VSS.n3864 VSS.n3863 0.214786
R25616 VSS.n3862 VSS.n2803 0.214786
R25617 VSS.n3861 VSS.n3860 0.214786
R25618 VSS.n3859 VSS.n3762 0.214786
R25619 VSS.n3858 VSS.n3857 0.214786
R25620 VSS.n3856 VSS.n3763 0.214786
R25621 VSS.n3855 VSS.n3854 0.214786
R25622 VSS.n3853 VSS.n3768 0.214786
R25623 VSS.n3852 VSS.n3851 0.214786
R25624 VSS.n3850 VSS.n3769 0.214786
R25625 VSS.n3849 VSS.n3848 0.214786
R25626 VSS.n3847 VSS.n3774 0.214786
R25627 VSS.n3846 VSS.n3845 0.214786
R25628 VSS.n3844 VSS.n3776 0.214786
R25629 VSS.n3843 VSS.n3842 0.214786
R25630 VSS.n3841 VSS.n3781 0.214786
R25631 VSS.n3840 VSS.n3839 0.214786
R25632 VSS.n3838 VSS.n3782 0.214786
R25633 VSS.n3837 VSS.n3836 0.214786
R25634 VSS.n3835 VSS.n3787 0.214786
R25635 VSS.n3834 VSS.n3833 0.214786
R25636 VSS.n3832 VSS.n3788 0.214786
R25637 VSS.n3831 VSS.n3830 0.214786
R25638 VSS.n3829 VSS.n3793 0.214786
R25639 VSS.n3828 VSS.n3827 0.214786
R25640 VSS.n3826 VSS.n3794 0.214786
R25641 VSS.n3825 VSS.n3824 0.214786
R25642 VSS.n3823 VSS.n3799 0.214786
R25643 VSS.n3822 VSS.n3821 0.214786
R25644 VSS.n3820 VSS.n3800 0.214786
R25645 VSS.n3819 VSS.n3818 0.214786
R25646 VSS.n3817 VSS.n3805 0.214786
R25647 VSS.n3816 VSS.n3815 0.214786
R25648 VSS.n3814 VSS.n3806 0.214786
R25649 VSS.n3813 VSS.n3812 0.214786
R25650 VSS.n2116 VSS.n2114 0.214786
R25651 VSS.n5387 VSS.n5386 0.214786
R25652 VSS.n5423 VSS.n2084 0.212265
R25653 VSS.n5683 VSS.n5682 0.201836
R25654 VSS.n5432 VSS.n5431 0.192412
R25655 VSS.n4079 VSS 0.189765
R25656 VSS VSS.n4079 0.189765
R25657 VSS.n5317 VSS.n5316 0.186214
R25658 VSS.n5318 VSS.n5317 0.186214
R25659 VSS.n3870 VSS.n3869 0.186214
R25660 VSS.n3871 VSS.n3870 0.186214
R25661 VSS.n1590 VSS.n1589 0.185484
R25662 VSS VSS.n3504 0.17855
R25663 VSS.n2232 VSS.n2231 0.178408
R25664 VSS.n2231 VSS.n2230 0.178408
R25665 VSS.n5271 VSS.n5269 0.178408
R25666 VSS.n2231 VSS.n2229 0.178408
R25667 VSS.n5271 VSS.n5270 0.178408
R25668 VSS.n2231 VSS.n2228 0.178408
R25669 VSS.n5271 VSS.n2204 0.178408
R25670 VSS.n2786 VSS.n2785 0.175807
R25671 VSS.n5246 DVSS 0.175804
R25672 VSS.n2428 DVSS 0.175804
R25673 VSS.n2431 DVSS 0.175804
R25674 VSS.n4140 DVSS 0.175804
R25675 VSS.n4240 DVSS 0.175804
R25676 VSS.n4202 DVSS 0.175804
R25677 VSS.n2357 DVSS 0.175804
R25678 VSS.n2359 DVSS 0.175804
R25679 VSS.n2429 DVSS 0.175729
R25680 VSS.n2241 DVSS 0.175729
R25681 VSS.n2356 DVSS 0.175729
R25682 VSS.n2360 DVSS 0.175729
R25683 VSS.n902 VSS.n901 0.173577
R25684 VSS.n670 VSS.n669 0.173577
R25685 VSS.n3730 DVSS 0.172116
R25686 VSS.n5339 DVSS 0.172116
R25687 VSS.n5308 DVSS 0.172116
R25688 VSS.n5389 DVSS 0.172116
R25689 VSS.n3866 DVSS 0.172116
R25690 VSS VSS.n3403 0.169912
R25691 VSS.n3485 VSS.n3478 0.168658
R25692 VSS.n3478 VSS.n2779 0.168658
R25693 VSS.n3876 VSS.n2772 0.168658
R25694 VSS.n3886 VSS.n2772 0.168658
R25695 VSS.n3874 VSS.n3873 0.166289
R25696 VSS.n282 VSS.n141 0.163909
R25697 VSS.n824 VSS.n823 0.163909
R25698 VSS.n752 VSS.n751 0.163909
R25699 VSS.n535 VSS.n365 0.161214
R25700 VSS.n217 VSS.n216 0.161214
R25701 VSS.n1141 VSS.n1140 0.149124
R25702 VSS.n4287 VSS.n4284 0.145461
R25703 VSS.n5157 DVSS 0.144526
R25704 VSS.n3414 DVSS 0.144421
R25705 VSS.n3410 DVSS 0.144187
R25706 VSS.n3413 DVSS 0.1436
R25707 DVSS VSS.n3412 0.1436
R25708 VSS.n3412 DVSS 0.1436
R25709 DVSS VSS.n3411 0.1436
R25710 DVSS VSS.n4143 0.143441
R25711 VSS.n4141 DVSS 0.143441
R25712 DVSS VSS.n4245 0.143441
R25713 VSS.n4243 DVSS 0.143441
R25714 VSS.n1004 VSS.n1003 0.141125
R25715 VSS.n572 VSS.n571 0.141125
R25716 VSS.n4143 VSS.n4142 0.140794
R25717 VSS.n4142 VSS.n4141 0.140794
R25718 VSS.n4245 VSS.n4244 0.140794
R25719 VSS.n4244 VSS.n4243 0.140794
R25720 VSS.n4080 VSS 0.139932
R25721 VSS.n3382 DVSS 0.138622
R25722 VSS.n1005 VSS.n104 0.137596
R25723 VSS.n569 VSS.n523 0.137559
R25724 VSS.n2889 VSS 0.1355
R25725 VSS.n2367 VSS 0.1355
R25726 VSS.n2294 VSS 0.1355
R25727 VSS.n4286 VSS 0.1355
R25728 VSS.n4289 VSS 0.1355
R25729 DVSS VSS.n2101 0.1355
R25730 VSS.n3400 VSS 0.1355
R25731 VSS.n4083 DVSS 0.132383
R25732 VSS.n906 VSS.n222 0.130943
R25733 VSS.n3183 DVSS 0.130618
R25734 VSS.n5175 DVSS 0.130618
R25735 VSS.n380 VSS.n221 0.130587
R25736 VSS.n3582 DVSS 0.130161
R25737 VSS.n1302 VSS.n1297 0.129009
R25738 VSS.n3072 VSS.n3071 0.128608
R25739 VSS.n3311 VSS.n3072 0.128203
R25740 VSS.n1395 DVSS 0.125798
R25741 VSS.n1395 VSS.n33 0.12265
R25742 VSS.n5240 DVSS 0.115647
R25743 VSS.n3009 VSS.n2975 0.114824
R25744 VSS.n3257 VSS.n3074 0.114824
R25745 VSS.n4067 VSS 0.113
R25746 VSS.n4073 VSS 0.113
R25747 VSS.n2454 VSS 0.113
R25748 DVSS VSS.n5157 0.111845
R25749 VSS.n3408 DVSS 0.111373
R25750 VSS.n2168 VSS.n2166 0.110634
R25751 VSS.n1080 VSS.n1077 0.110634
R25752 VSS.n1137 VSS.n1136 0.110634
R25753 VSS.n1029 VSS.n1028 0.110634
R25754 VSS.n2363 VSS 0.110353
R25755 VSS.n3318 VSS.n2947 0.109959
R25756 VSS.n3319 VSS.n3318 0.109959
R25757 VSS.n916 VSS.n915 0.107643
R25758 VSS.n631 VSS.n630 0.107643
R25759 DVSS VSS.n3408 0.107291
R25760 VSS.n3875 VSS.n2779 0.107079
R25761 VSS.n2800 VSS.n2799 0.105895
R25762 VSS.n1584 VSS.n1302 0.102277
R25763 VSS.n3412 DVSS 0.102157
R25764 VSS.n5677 VSS.n8 0.101471
R25765 VSS.n5441 VSS.n5440 0.101471
R25766 DVSS VSS.n3582 0.101206
R25767 VSS.n3183 DVSS 0.10093
R25768 VSS.n5175 DVSS 0.10093
R25769 DVSS VSS.n3392 0.0991804
R25770 VSS.n1589 VSS.n1296 0.0985668
R25771 VSS.n1589 VSS.n1588 0.0984658
R25772 VSS.n2787 VSS 0.0939292
R25773 VSS.n3394 VSS 0.0939292
R25774 VSS.n3396 VSS 0.0939292
R25775 VSS.n2188 VSS 0.0939292
R25776 VSS.n2190 VSS 0.0939292
R25777 VSS.n4047 VSS 0.0939292
R25778 VSS.n3874 VSS 0.0928684
R25779 VSS.n4308 VSS.n4294 0.0921154
R25780 VSS.n5431 VSS.n5430 0.0891765
R25781 VSS.n5284 VSS.n5283 0.0883604
R25782 VSS.n3408 DVSS 0.0837012
R25783 VSS.n3525 VSS.n2199 0.08175
R25784 VSS.n3532 VSS.n2201 0.08175
R25785 DVSS VSS.n5406 0.0812353
R25786 DVSS VSS.n5310 0.0812353
R25787 DVSS VSS.n5311 0.0812353
R25788 VSS.n3107 VSS.n2957 0.077375
R25789 VSS.n3334 VSS.n2949 0.077375
R25790 DVSS VSS.n5423 0.0772647
R25791 VSS.n5251 VSS.n2238 0.0769706
R25792 VSS.n5251 VSS.n5250 0.0769706
R25793 VSS.n2380 VSS.n2377 0.0769376
R25794 VSS.n3314 VSS.n3313 0.0763777
R25795 VSS.n4908 DVSS 0.0761
R25796 VSS.n4627 DVSS 0.0761
R25797 DVSS VSS.n4630 0.0761
R25798 VSS.n4821 DVSS 0.0761
R25799 DVSS VSS.n4500 0.0761
R25800 VSS.n4790 DVSS 0.0761
R25801 DVSS VSS.n4448 0.0761
R25802 VSS.n4747 DVSS 0.0761
R25803 DVSS VSS.n4638 0.0761
R25804 VSS.n4639 DVSS 0.0761
R25805 DVSS VSS.n4357 0.0761
R25806 VSS.n4681 DVSS 0.0761
R25807 DVSS VSS.n4645 0.0761
R25808 VSS.n4646 DVSS 0.0761
R25809 VSS.n3314 VSS.n2971 0.0756596
R25810 VSS.n3413 DVSS 0.0748392
R25811 VSS.n3411 DVSS 0.0746758
R25812 VSS.n4311 VSS.n4308 0.0745555
R25813 VSS.n2065 VSS.n1598 0.0741096
R25814 VSS.n5131 DVSS 0.0728785
R25815 DVSS VSS.n2284 0.0728785
R25816 VSS.n3728 VSS.n2819 0.0728571
R25817 VSS.n3380 VSS.n2893 0.0693638
R25818 VSS.n3402 VSS.n2296 0.0668158
R25819 VSS.n3504 VSS.n3418 0.0656316
R25820 VSS.n2059 VSS.n1598 0.0624601
R25821 VSS.n3876 VSS.n3875 0.0620789
R25822 VSS.n2381 VSS.n2380 0.0599397
R25823 VSS.n38 VSS.n35 0.0597445
R25824 VSS.n40 VSS.n39 0.0597445
R25825 VSS.n42 VSS.n41 0.0597445
R25826 VSS.n44 VSS.n43 0.0597445
R25827 VSS.n46 VSS.n45 0.0597445
R25828 VSS.n48 VSS.n47 0.0597445
R25829 VSS.n50 VSS.n49 0.0597445
R25830 VSS.n52 VSS.n51 0.0597445
R25831 VSS.n54 VSS.n53 0.0597445
R25832 VSS.n67 VSS.n56 0.0597445
R25833 VSS.n76 VSS.n66 0.0597445
R25834 VSS.n75 VSS.n65 0.0597445
R25835 VSS.n74 VSS.n64 0.0597445
R25836 VSS.n73 VSS.n63 0.0597445
R25837 VSS.n72 VSS.n62 0.0597445
R25838 VSS.n71 VSS.n61 0.0597445
R25839 VSS.n70 VSS.n60 0.0597445
R25840 VSS.n69 VSS.n59 0.0597445
R25841 VSS.n68 VSS.n58 0.0597445
R25842 VSS.n1143 VSS.n35 0.0597445
R25843 VSS.n39 VSS.n38 0.0597445
R25844 VSS.n41 VSS.n40 0.0597445
R25845 VSS.n43 VSS.n42 0.0597445
R25846 VSS.n45 VSS.n44 0.0597445
R25847 VSS.n47 VSS.n46 0.0597445
R25848 VSS.n49 VSS.n48 0.0597445
R25849 VSS.n51 VSS.n50 0.0597445
R25850 VSS.n53 VSS.n52 0.0597445
R25851 VSS.n55 VSS.n54 0.0597445
R25852 VSS.n76 VSS.n67 0.0597445
R25853 VSS.n75 VSS.n66 0.0597445
R25854 VSS.n74 VSS.n65 0.0597445
R25855 VSS.n73 VSS.n64 0.0597445
R25856 VSS.n72 VSS.n63 0.0597445
R25857 VSS.n71 VSS.n62 0.0597445
R25858 VSS.n70 VSS.n61 0.0597445
R25859 VSS.n69 VSS.n60 0.0597445
R25860 VSS.n68 VSS.n59 0.0597445
R25861 VSS.n2077 VSS.n2076 0.0588383
R25862 VSS.n3312 VSS.n2973 0.058625
R25863 VSS.n3070 VSS.n3069 0.058625
R25864 VSS.n3376 VSS.n2893 0.0585457
R25865 VSS.n2821 VSS.n2819 0.058308
R25866 DVSS VSS.n3392 0.0574691
R25867 VSS.n5694 VSS.n16 0.0562784
R25868 VSS.n3072 VSS.n2967 0.0546667
R25869 VSS.n3316 VSS.n2967 0.0546667
R25870 VSS.n3318 VSS.n3317 0.0546667
R25871 VSS.n3317 VSS.n3316 0.0546667
R25872 VSS.n3109 VSS.n3108 0.0544368
R25873 VSS.n3110 VSS.n3109 0.0544368
R25874 VSS.n3067 VSS.n3066 0.0544368
R25875 VSS.n3067 VSS.n3060 0.0544368
R25876 VSS.n2362 VSS 0.0537197
R25877 VSS.n2364 VSS 0.0537197
R25878 VSS.n3360 VSS.n2907 0.0532027
R25879 VSS.n3250 VSS.n3247 0.0532027
R25880 VSS.n5694 VSS.n5693 0.0500653
R25881 VSS.n3529 VSS.n3528 0.0495566
R25882 VSS.n5282 VSS.n5281 0.0495566
R25883 VSS.n3533 VSS.n3532 0.0486793
R25884 VSS.n2784 VSS 0.0456808
R25885 VSS.n4060 VSS 0.0456808
R25886 VSS.n2446 VSS 0.0456808
R25887 VSS.n2447 VSS 0.0456808
R25888 VSS.n2449 VSS 0.0456808
R25889 VSS.n3132 VSS.n3131 0.0450872
R25890 VSS.n2941 VSS.n2939 0.0450872
R25891 VSS.n3290 VSS.n3289 0.0450872
R25892 VSS.n3020 VSS.n3019 0.0450872
R25893 VSS.n3055 VSS.n3028 0.0450872
R25894 VSS.n2910 VSS.n2908 0.0450718
R25895 VSS.n2912 VSS.n2910 0.0450718
R25896 VSS.n2917 VSS.n2916 0.0450718
R25897 VSS.n2918 VSS.n2917 0.0450718
R25898 VSS.n3136 VSS.n3095 0.0450718
R25899 VSS.n3095 VSS.n3093 0.0450718
R25900 VSS.n3269 VSS.n3253 0.0442838
R25901 VSS.n3262 VSS.n3261 0.0442838
R25902 VSS.n3271 VSS.n3270 0.0442838
R25903 VSS.n3270 VSS.n3254 0.0442838
R25904 VSS.n3264 VSS.n3263 0.0442838
R25905 VSS.n3021 VSS.n3013 0.0442838
R25906 VSS.n3022 VSS.n3021 0.0442838
R25907 VSS.n3027 VSS.n3026 0.0442838
R25908 VSS.n3360 VSS.n3359 0.0442838
R25909 VSS.n3357 VSS.n3356 0.0442838
R25910 VSS.n3356 VSS.n2913 0.0442838
R25911 VSS.n2936 VSS.n2935 0.0442838
R25912 VSS.n2937 VSS.n2936 0.0442838
R25913 VSS.n2942 VSS.n2937 0.0442838
R25914 VSS.n2943 VSS.n2942 0.0442838
R25915 VSS.n3339 VSS.n2943 0.0442838
R25916 VSS.n3339 VSS.n3338 0.0442838
R25917 VSS.n3338 VSS.n2944 0.0442838
R25918 VSS.n3115 VSS.n2963 0.0442838
R25919 VSS.n3117 VSS.n3115 0.0442838
R25920 VSS.n3117 VSS.n3116 0.0442838
R25921 VSS.n3116 VSS.n3098 0.0442838
R25922 VSS.n3133 VSS.n3098 0.0442838
R25923 VSS.n3134 VSS.n3133 0.0442838
R25924 VSS.n3134 VSS.n3096 0.0442838
R25925 VSS.n3142 VSS.n3141 0.0442838
R25926 VSS.n3292 VSS.n3142 0.0442838
R25927 VSS.n3292 VSS.n3291 0.0442838
R25928 VSS.n3291 VSS.n3143 0.0442838
R25929 VSS.n3249 VSS.n3143 0.0442838
R25930 VSS.n3250 VSS.n3249 0.0442838
R25931 VSS.n2839 VSS.n2199 0.0432989
R25932 VSS.n3135 VSS.n3097 0.0430229
R25933 VSS.n2938 VSS.n2914 0.0430229
R25934 VSS.n3023 VSS.n3012 0.0426101
R25935 VSS.n3293 VSS.n3092 0.0421972
R25936 VSS.n3352 VSS.n2921 0.0418677
R25937 VSS.n3137 VSS.n3079 0.0418677
R25938 VSS.n3268 VSS.n3267 0.0418514
R25939 VSS.n5695 VSS.n5694 0.0417698
R25940 VSS.n5696 VSS.n5695 0.0417698
R25941 VSS.n2078 VSS.n2077 0.0417698
R25942 VSS.n2079 VSS.n2078 0.0417698
R25943 VSS.n3118 VSS.n3114 0.0405459
R25944 VSS.n3340 VSS.n2934 0.0405459
R25945 VSS.n4446 VSS.n2285 0.0398939
R25946 VSS.n5124 VSS.n2285 0.0398939
R25947 VSS.n4748 VSS.n2286 0.0398939
R25948 VSS.n5124 VSS.n2286 0.0398939
R25949 VSS.n3362 VSS.n3361 0.0397202
R25950 VSS.n3264 VSS.n3256 0.0382027
R25951 VSS.n3026 VSS.n3011 0.0382027
R25952 VSS.n3315 VSS.n3314 0.0381812
R25953 VSS.n3316 VSS.n3315 0.0381812
R25954 VSS.n3253 VSS.n3154 0.0373919
R25955 VSS.n3733 VSS.n3732 0.0359178
R25956 VSS.n3531 VSS.n3530 0.0357988
R25957 VSS.n2788 VSS 0.0348421
R25958 VSS.n3288 VSS.n3144 0.0339404
R25959 VSS.n377 VSS.n372 0.0336863
R25960 VSS.n579 VSS.n373 0.0336863
R25961 VSS.n5416 VSS.n5415 0.0336579
R25962 VSS.n5322 VSS.n2181 0.0336579
R25963 VSS.n5325 VSS.n5324 0.0336579
R25964 VSS.n5419 VSS.n5418 0.0336579
R25965 VSS.n578 VSS.n374 0.0332409
R25966 VSS.n3130 VSS.n3099 0.0331147
R25967 VSS.n2940 VSS.n2933 0.0331147
R25968 VSS.n1877 VSS.n14 0.033
R25969 VSS.n14 VSS.n13 0.033
R25970 VSS.n1746 VSS.n1745 0.033
R25971 VSS.n1745 VSS.n1744 0.033
R25972 VSS.n1728 VSS.n1704 0.033
R25973 VSS.n1743 VSS.n1728 0.033
R25974 VSS.n1741 VSS.n1740 0.033
R25975 VSS.n1742 VSS.n1741 0.033
R25976 VSS.n1735 VSS.n1734 0.033
R25977 VSS.n1735 VSS.n1729 0.033
R25978 VSS.n2042 VSS.n1295 0.033
R25979 VSS.n1295 VSS.n1293 0.033
R25980 VSS.n5411 VSS.n2101 0.0322647
R25981 VSS.n3058 VSS.n3008 0.031778
R25982 VSS.n3309 VSS.n3308 0.031778
R25983 VSS.n5113 VSS.n4299 0.0315
R25984 VSS.n4337 VSS.n4323 0.0315
R25985 VSS.n4337 VSS.n4335 0.0315
R25986 VSS.n5073 VSS.n5072 0.0315
R25987 VSS.n4390 VSS.n4387 0.0315
R25988 VSS.n4426 VSS.n4411 0.0315
R25989 VSS.n5009 VSS.n5008 0.0315
R25990 VSS.n4480 VSS.n4477 0.0315
R25991 VSS.n4517 VSS.n4502 0.0315
R25992 VSS.n4945 VSS.n4944 0.0315
R25993 VSS.n4923 VSS.n4569 0.0315
R25994 VSS.n4604 VSS.n4590 0.0315
R25995 VSS.n4604 VSS.n4602 0.0315
R25996 VSS.n4882 VSS.n4881 0.0315
R25997 VSS.n4648 VSS.n4295 0.0315
R25998 VSS.n4666 VSS.n4665 0.0315
R25999 VSS.n4667 VSS.n4666 0.0315
R26000 VSS.n4683 VSS.n4642 0.0315
R26001 VSS.n4710 VSS.n4709 0.0315
R26002 VSS.n4731 VSS.n4730 0.0315
R26003 VSS.n4750 VSS.n4635 0.0315
R26004 VSS.n4777 VSS.n4776 0.0315
R26005 VSS.n4799 VSS.n4798 0.0315
R26006 VSS.n4819 VSS.n4818 0.0315
R26007 VSS.n4840 VSS.n4839 0.0315
R26008 VSS.n4858 VSS.n4857 0.0315
R26009 VSS.n4859 VSS.n4858 0.0315
R26010 VSS.n4875 VSS.n4625 0.0315
R26011 VSS.n3025 VSS.n3010 0.0310505
R26012 VSS.n5114 VSS.n4298 0.031
R26013 VSS.n5069 VSS.n4358 0.031
R26014 VSS.n4924 VSS.n4568 0.031
R26015 VSS.n5132 VSS.n2282 0.031
R26016 VSS.n5117 VSS.n5116 0.031
R26017 VSS.n4693 VSS.n4692 0.031
R26018 VSS.n4836 VSS.n4565 0.031
R26019 VSS.n4624 VSS.n2281 0.031
R26020 VSS.n3263 VSS.n3257 0.0309054
R26021 VSS.n3027 VSS.n3009 0.0309054
R26022 VSS.n387 VSS.n374 0.0309017
R26023 VSS.n3252 VSS.n3251 0.0306376
R26024 VSS.n3265 VSS.n3255 0.0305
R26025 VSS.n5049 VSS.n5048 0.0305
R26026 VSS.n4948 VSS.n4534 0.0305
R26027 VSS.n4713 VSS.n4385 0.0305
R26028 VSS.n4817 VSS.n4815 0.0305
R26029 VSS.n385 VSS.n377 0.0304416
R26030 VSS.n386 VSS.n373 0.0304416
R26031 VSS.n3355 VSS.n3354 0.0302248
R26032 VSS.n3139 VSS.n3091 0.0302248
R26033 VSS.n1144 VSS.n1143 0.0301222
R26034 VSS.n1141 VSS.n55 0.0301222
R26035 VSS.n1140 VSS.n56 0.0301222
R26036 VSS.n1078 VSS.n58 0.0301222
R26037 VSS.n4425 VSS.n4423 0.03
R26038 VSS.n4969 VSS.n4968 0.03
R26039 VSS.n4733 VSS.n4732 0.03
R26040 VSS.n4795 VSS.n4504 0.03
R26041 VSS.n3734 VSS.n3733 0.0298971
R26042 VSS.n5005 VSS.n4447 0.0295
R26043 VSS.n4479 VSS.n4465 0.0295
R26044 VSS.n4760 VSS.n4759 0.0295
R26045 VSS.n4773 VSS.n4633 0.0295
R26046 VSS.n5012 VSS.n4443 0.029
R26047 VSS.n4985 VSS.n4984 0.029
R26048 VSS.n4751 VSS.n4636 0.029
R26049 VSS.n4780 VSS.n4475 0.029
R26050 VSS.n3025 VSS.n3024 0.0285734
R26051 VSS.n5033 VSS.n5032 0.0285
R26052 VSS.n4516 VSS.n4514 0.0285
R26053 VSS.n4727 VSS.n4413 0.0285
R26054 VSS.n4801 VSS.n4800 0.0285
R26055 VSS.n184 VSS.n105 0.0283304
R26056 VSS.n185 VSS.n184 0.0283304
R26057 VSS.n186 VSS.n185 0.0283304
R26058 VSS.n186 VSS.n181 0.0283304
R26059 VSS.n190 VSS.n181 0.0283304
R26060 VSS.n191 VSS.n190 0.0283304
R26061 VSS.n192 VSS.n191 0.0283304
R26062 VSS.n192 VSS.n179 0.0283304
R26063 VSS.n196 VSS.n179 0.0283304
R26064 VSS.n197 VSS.n196 0.0283304
R26065 VSS.n198 VSS.n197 0.0283304
R26066 VSS.n198 VSS.n177 0.0283304
R26067 VSS.n202 VSS.n177 0.0283304
R26068 VSS.n203 VSS.n202 0.0283304
R26069 VSS.n204 VSS.n203 0.0283304
R26070 VSS.n204 VSS.n175 0.0283304
R26071 VSS.n208 VSS.n175 0.0283304
R26072 VSS.n209 VSS.n208 0.0283304
R26073 VSS.n210 VSS.n209 0.0283304
R26074 VSS.n210 VSS.n173 0.0283304
R26075 VSS.n214 VSS.n173 0.0283304
R26076 VSS.n215 VSS.n214 0.0283304
R26077 VSS.n914 VSS.n171 0.0283304
R26078 VSS.n233 VSS.n171 0.0283304
R26079 VSS.n234 VSS.n233 0.0283304
R26080 VSS.n234 VSS.n232 0.0283304
R26081 VSS.n238 VSS.n232 0.0283304
R26082 VSS.n239 VSS.n238 0.0283304
R26083 VSS.n240 VSS.n239 0.0283304
R26084 VSS.n240 VSS.n230 0.0283304
R26085 VSS.n244 VSS.n230 0.0283304
R26086 VSS.n245 VSS.n244 0.0283304
R26087 VSS.n246 VSS.n245 0.0283304
R26088 VSS.n246 VSS.n228 0.0283304
R26089 VSS.n250 VSS.n228 0.0283304
R26090 VSS.n251 VSS.n250 0.0283304
R26091 VSS.n252 VSS.n251 0.0283304
R26092 VSS.n252 VSS.n226 0.0283304
R26093 VSS.n256 VSS.n226 0.0283304
R26094 VSS.n257 VSS.n256 0.0283304
R26095 VSS.n258 VSS.n257 0.0283304
R26096 VSS.n258 VSS.n224 0.0283304
R26097 VSS.n262 VSS.n224 0.0283304
R26098 VSS.n904 VSS.n903 0.0283304
R26099 VSS.n3294 VSS.n3091 0.0281606
R26100 VSS.n3266 VSS.n3265 0.0280676
R26101 VSS.n4389 VSS.n4375 0.028
R26102 VSS.n4943 VSS.n4538 0.028
R26103 VSS.n4706 VSS.n4640 0.028
R26104 VSS.n4823 VSS.n4540 0.028
R26105 VSS.n5058 VSS.n4374 0.0279877
R26106 VSS.n5023 VSS.n4428 0.0279877
R26107 VSS.n4922 VSS.n4570 0.0279877
R26108 VSS.n4707 VSS.n4705 0.0279877
R26109 VSS.n4735 VSS.n4734 0.0279877
R26110 VSS.n4838 VSS.n4837 0.0279877
R26111 VSS.n5112 VSS.n4300 0.0279877
R26112 VSS.n5112 VSS.n5111 0.0279877
R26113 VSS.n5111 VSS.n5110 0.0279877
R26114 VSS.n5110 VSS.n4301 0.0279877
R26115 VSS.n5099 VSS.n4321 0.0279877
R26116 VSS.n5099 VSS.n5098 0.0279877
R26117 VSS.n5098 VSS.n4322 0.0279877
R26118 VSS.n4338 VSS.n4322 0.0279877
R26119 VSS.n4339 VSS.n4338 0.0279877
R26120 VSS.n5087 VSS.n4339 0.0279877
R26121 VSS.n5087 VSS.n5086 0.0279877
R26122 VSS.n4356 VSS.n4355 0.0279877
R26123 VSS.n5075 VSS.n4356 0.0279877
R26124 VSS.n5075 VSS.n5074 0.0279877
R26125 VSS.n5071 VSS.n5070 0.0279877
R26126 VSS.n5070 VSS.n4359 0.0279877
R26127 VSS.n4373 VSS.n4359 0.0279877
R26128 VSS.n5059 VSS.n4373 0.0279877
R26129 VSS.n5059 VSS.n5058 0.0279877
R26130 VSS.n4391 VSS.n4374 0.0279877
R26131 VSS.n5047 VSS.n4392 0.0279877
R26132 VSS.n5047 VSS.n5046 0.0279877
R26133 VSS.n5046 VSS.n4393 0.0279877
R26134 VSS.n5035 VSS.n4409 0.0279877
R26135 VSS.n5035 VSS.n5034 0.0279877
R26136 VSS.n5034 VSS.n4410 0.0279877
R26137 VSS.n4427 VSS.n4410 0.0279877
R26138 VSS.n4428 VSS.n4427 0.0279877
R26139 VSS.n5023 VSS.n5022 0.0279877
R26140 VSS.n4445 VSS.n4444 0.0279877
R26141 VSS.n5011 VSS.n4445 0.0279877
R26142 VSS.n5011 VSS.n5010 0.0279877
R26143 VSS.n5007 VSS.n5006 0.0279877
R26144 VSS.n5006 VSS.n4449 0.0279877
R26145 VSS.n4463 VSS.n4449 0.0279877
R26146 VSS.n4995 VSS.n4463 0.0279877
R26147 VSS.n4995 VSS.n4994 0.0279877
R26148 VSS.n4994 VSS.n4464 0.0279877
R26149 VSS.n4481 VSS.n4464 0.0279877
R26150 VSS.n4983 VSS.n4482 0.0279877
R26151 VSS.n4983 VSS.n4982 0.0279877
R26152 VSS.n4982 VSS.n4483 0.0279877
R26153 VSS.n4499 VSS.n4483 0.0279877
R26154 VSS.n4971 VSS.n4970 0.0279877
R26155 VSS.n4970 VSS.n4501 0.0279877
R26156 VSS.n4518 VSS.n4501 0.0279877
R26157 VSS.n4519 VSS.n4518 0.0279877
R26158 VSS.n4959 VSS.n4519 0.0279877
R26159 VSS.n4959 VSS.n4958 0.0279877
R26160 VSS.n4536 VSS.n4535 0.0279877
R26161 VSS.n4947 VSS.n4536 0.0279877
R26162 VSS.n4947 VSS.n4946 0.0279877
R26163 VSS.n4946 VSS.n4537 0.0279877
R26164 VSS.n4629 VSS.n4553 0.0279877
R26165 VSS.n4934 VSS.n4553 0.0279877
R26166 VSS.n4934 VSS.n4933 0.0279877
R26167 VSS.n4933 VSS.n4554 0.0279877
R26168 VSS.n4570 VSS.n4554 0.0279877
R26169 VSS.n4921 VSS.n4920 0.0279877
R26170 VSS.n4920 VSS.n4571 0.0279877
R26171 VSS.n4588 VSS.n4571 0.0279877
R26172 VSS.n4909 VSS.n4588 0.0279877
R26173 VSS.n4907 VSS.n4589 0.0279877
R26174 VSS.n4605 VSS.n4589 0.0279877
R26175 VSS.n4606 VSS.n4605 0.0279877
R26176 VSS.n4896 VSS.n4606 0.0279877
R26177 VSS.n4896 VSS.n4895 0.0279877
R26178 VSS.n4895 VSS.n4607 0.0279877
R26179 VSS.n4884 VSS.n4880 0.0279877
R26180 VSS.n4884 VSS.n4883 0.0279877
R26181 VSS.n4883 VSS.n2283 0.0279877
R26182 VSS.n5131 VSS.n2283 0.0279877
R26183 VSS.n5118 VSS.n4293 0.0279877
R26184 VSS.n4647 VSS.n4293 0.0279877
R26185 VSS.n4652 VSS.n4647 0.0279877
R26186 VSS.n4653 VSS.n4652 0.0279877
R26187 VSS.n4658 VSS.n4657 0.0279877
R26188 VSS.n4663 VSS.n4658 0.0279877
R26189 VSS.n4664 VSS.n4663 0.0279877
R26190 VSS.n4664 VSS.n4644 0.0279877
R26191 VSS.n4668 VSS.n4644 0.0279877
R26192 VSS.n4669 VSS.n4668 0.0279877
R26193 VSS.n4674 VSS.n4669 0.0279877
R26194 VSS.n4679 VSS.n4675 0.0279877
R26195 VSS.n4680 VSS.n4679 0.0279877
R26196 VSS.n4682 VSS.n4680 0.0279877
R26197 VSS.n4694 VSS.n4641 0.0279877
R26198 VSS.n4695 VSS.n4694 0.0279877
R26199 VSS.n4699 VSS.n4695 0.0279877
R26200 VSS.n4700 VSS.n4699 0.0279877
R26201 VSS.n4705 VSS.n4700 0.0279877
R26202 VSS.n4708 VSS.n4707 0.0279877
R26203 VSS.n4712 VSS.n4711 0.0279877
R26204 VSS.n4717 VSS.n4712 0.0279877
R26205 VSS.n4718 VSS.n4717 0.0279877
R26206 VSS.n4723 VSS.n4722 0.0279877
R26207 VSS.n4728 VSS.n4723 0.0279877
R26208 VSS.n4729 VSS.n4728 0.0279877
R26209 VSS.n4729 VSS.n4637 0.0279877
R26210 VSS.n4734 VSS.n4637 0.0279877
R26211 VSS.n4740 VSS.n4735 0.0279877
R26212 VSS.n4745 VSS.n4741 0.0279877
R26213 VSS.n4746 VSS.n4745 0.0279877
R26214 VSS.n4749 VSS.n4746 0.0279877
R26215 VSS.n4761 VSS.n4634 0.0279877
R26216 VSS.n4762 VSS.n4761 0.0279877
R26217 VSS.n4766 VSS.n4762 0.0279877
R26218 VSS.n4767 VSS.n4766 0.0279877
R26219 VSS.n4772 VSS.n4767 0.0279877
R26220 VSS.n4774 VSS.n4772 0.0279877
R26221 VSS.n4775 VSS.n4774 0.0279877
R26222 VSS.n4779 VSS.n4778 0.0279877
R26223 VSS.n4784 VSS.n4779 0.0279877
R26224 VSS.n4785 VSS.n4784 0.0279877
R26225 VSS.n4789 VSS.n4785 0.0279877
R26226 VSS.n4796 VSS.n4791 0.0279877
R26227 VSS.n4797 VSS.n4796 0.0279877
R26228 VSS.n4797 VSS.n4632 0.0279877
R26229 VSS.n4802 VSS.n4632 0.0279877
R26230 VSS.n4803 VSS.n4802 0.0279877
R26231 VSS.n4808 VSS.n4803 0.0279877
R26232 VSS.n4813 VSS.n4809 0.0279877
R26233 VSS.n4814 VSS.n4813 0.0279877
R26234 VSS.n4814 VSS.n4631 0.0279877
R26235 VSS.n4820 VSS.n4631 0.0279877
R26236 VSS.n4826 VSS.n4822 0.0279877
R26237 VSS.n4827 VSS.n4826 0.0279877
R26238 VSS.n4832 VSS.n4827 0.0279877
R26239 VSS.n4833 VSS.n4832 0.0279877
R26240 VSS.n4837 VSS.n4833 0.0279877
R26241 VSS.n4844 VSS.n4628 0.0279877
R26242 VSS.n4845 VSS.n4844 0.0279877
R26243 VSS.n4849 VSS.n4845 0.0279877
R26244 VSS.n4850 VSS.n4849 0.0279877
R26245 VSS.n4856 VSS.n4855 0.0279877
R26246 VSS.n4856 VSS.n4626 0.0279877
R26247 VSS.n4860 VSS.n4626 0.0279877
R26248 VSS.n4861 VSS.n4860 0.0279877
R26249 VSS.n4866 VSS.n4861 0.0279877
R26250 VSS.n4867 VSS.n4866 0.0279877
R26251 VSS.n4872 VSS.n4871 0.0279877
R26252 VSS.n4874 VSS.n4872 0.0279877
R26253 VSS.n4874 VSS.n4873 0.0279877
R26254 VSS.n4873 VSS.n2284 0.0279877
R26255 VSS.n4971 VSS.n4500 0.0275443
R26256 VSS.n4791 VSS.n4790 0.0275443
R26257 VSS.n5109 VSS.n4302 0.0275
R26258 VSS.n5076 VSS.n4354 0.0275
R26259 VSS.n4919 VSS.n4572 0.0275
R26260 VSS.n4885 VSS.n4879 0.0275
R26261 VSS.n4651 VSS.n4650 0.0275
R26262 VSS.n4684 VSS.n4643 0.0275
R26263 VSS.n4843 VSS.n4842 0.0275
R26264 VSS.n4876 VSS.n4623 0.0275
R26265 VSS.n3110 VSS.n2973 0.0274684
R26266 VSS.n3108 VSS.n3107 0.0274684
R26267 VSS.n3069 VSS.n3060 0.0274684
R26268 VSS.n3066 VSS.n2949 0.0274684
R26269 VSS.n904 VSS.n222 0.0272082
R26270 VSS.n5097 VSS.n5096 0.027
R26271 VSS.n5089 VSS.n5088 0.027
R26272 VSS.n4906 VSS.n4905 0.027
R26273 VSS.n4898 VSS.n4897 0.027
R26274 VSS.n4662 VSS.n4325 0.027
R26275 VSS.n4670 VSS.n4333 0.027
R26276 VSS.n4854 VSS.n4592 0.027
R26277 VSS.n4862 VSS.n4600 0.027
R26278 VSS.n3047 VSS.n3044 0.026913
R26279 VSS.n3044 VSS.n3043 0.026913
R26280 VSS.n3043 VSS.n3041 0.026913
R26281 VSS.n3041 VSS.n3039 0.026913
R26282 VSS.n3039 VSS.n3037 0.026913
R26283 VSS.n3037 VSS.n3034 0.026913
R26284 VSS.n3034 VSS.n3033 0.026913
R26285 VSS.n3033 VSS.n3031 0.026913
R26286 VSS.n3031 VSS.n2839 0.026913
R26287 VSS.n3547 VSS.n3531 0.026913
R26288 VSS.n3547 VSS.n3546 0.026913
R26289 VSS.n3546 VSS.n3544 0.026913
R26290 VSS.n3544 VSS.n3541 0.026913
R26291 VSS.n3541 VSS.n3540 0.026913
R26292 VSS.n3540 VSS.n3538 0.026913
R26293 VSS.n3538 VSS.n3536 0.026913
R26294 VSS.n3536 VSS.n3533 0.026913
R26295 VSS.n2886 VSS.n2884 0.026913
R26296 VSS.n3543 VSS.n3542 0.026913
R26297 VSS.n3535 VSS.n3534 0.026913
R26298 VSS.n3726 VSS.n2819 0.0267204
R26299 VSS.n3378 VSS.n2893 0.0267108
R26300 VSS.n3119 VSS.n3099 0.0265092
R26301 VSS.n3341 VSS.n2933 0.0265092
R26302 VSS.n5068 VSS.n4360 0.0265
R26303 VSS.n4567 VSS.n4555 0.0265
R26304 VSS.n4696 VSS.n4362 0.0265
R26305 VSS.n4835 VSS.n4834 0.0265
R26306 VSS.n4054 VSS.n4053 0.02615
R26307 VSS.n5045 VSS.n4388 0.026
R26308 VSS.n4949 VSS.n4533 0.026
R26309 VSS.n4716 VSS.n4715 0.026
R26310 VSS.n4812 VSS.n4530 0.026
R26311 VSS.n2380 VSS.n2379 0.0259029
R26312 VSS.n570 VSS.n524 0.0257489
R26313 VSS.n566 VSS.n524 0.0257489
R26314 VSS.n566 VSS.n565 0.0257489
R26315 VSS.n565 VSS.n564 0.0257489
R26316 VSS.n564 VSS.n526 0.0257489
R26317 VSS.n560 VSS.n526 0.0257489
R26318 VSS.n560 VSS.n559 0.0257489
R26319 VSS.n559 VSS.n558 0.0257489
R26320 VSS.n558 VSS.n528 0.0257489
R26321 VSS.n554 VSS.n528 0.0257489
R26322 VSS.n554 VSS.n553 0.0257489
R26323 VSS.n553 VSS.n552 0.0257489
R26324 VSS.n552 VSS.n530 0.0257489
R26325 VSS.n548 VSS.n530 0.0257489
R26326 VSS.n548 VSS.n547 0.0257489
R26327 VSS.n547 VSS.n546 0.0257489
R26328 VSS.n546 VSS.n532 0.0257489
R26329 VSS.n542 VSS.n532 0.0257489
R26330 VSS.n542 VSS.n541 0.0257489
R26331 VSS.n541 VSS.n540 0.0257489
R26332 VSS.n540 VSS.n534 0.0257489
R26333 VSS.n536 VSS.n534 0.0257489
R26334 VSS.n632 VSS.n364 0.0257489
R26335 VSS.n637 VSS.n364 0.0257489
R26336 VSS.n638 VSS.n637 0.0257489
R26337 VSS.n639 VSS.n638 0.0257489
R26338 VSS.n639 VSS.n362 0.0257489
R26339 VSS.n643 VSS.n362 0.0257489
R26340 VSS.n644 VSS.n643 0.0257489
R26341 VSS.n645 VSS.n644 0.0257489
R26342 VSS.n645 VSS.n360 0.0257489
R26343 VSS.n649 VSS.n360 0.0257489
R26344 VSS.n650 VSS.n649 0.0257489
R26345 VSS.n651 VSS.n650 0.0257489
R26346 VSS.n651 VSS.n358 0.0257489
R26347 VSS.n655 VSS.n358 0.0257489
R26348 VSS.n656 VSS.n655 0.0257489
R26349 VSS.n657 VSS.n656 0.0257489
R26350 VSS.n657 VSS.n356 0.0257489
R26351 VSS.n661 VSS.n356 0.0257489
R26352 VSS.n662 VSS.n661 0.0257489
R26353 VSS.n663 VSS.n662 0.0257489
R26354 VSS.n663 VSS.n353 0.0257489
R26355 VSS.n668 VSS.n354 0.0257489
R26356 VSS.n3248 VSS.n3144 0.0256835
R26357 VSS.n4355 DVSS 0.0255493
R26358 VSS.n4675 DVSS 0.0255493
R26359 VSS.n5025 VSS.n5024 0.0255
R26360 VSS.n4972 VSS.n4498 0.0255
R26361 VSS.n4736 VSS.n4421 0.0255
R26362 VSS.n4794 VSS.n4792 0.0255
R26363 VSS.n5004 VSS.n4450 0.025
R26364 VSS.n4993 VSS.n4992 0.025
R26365 VSS.n4763 VSS.n4452 0.025
R26366 VSS.n4771 VSS.n4467 0.025
R26367 VSS.n903 VSS.n902 0.0249638
R26368 VSS.n4630 VSS.n4629 0.0248842
R26369 VSS.n4822 VSS.n4821 0.0248842
R26370 VSS.n1613 VSS.n1598 0.0248508
R26371 VSS.n4309 VSS.n4308 0.0247925
R26372 VSS.n380 VSS.n354 0.0247308
R26373 VSS.n5013 VSS.n4442 0.0245
R26374 VSS.n4981 VSS.n4478 0.0245
R26375 VSS.n4744 VSS.n4439 0.0245
R26376 VSS.n4783 VSS.n4782 0.0245
R26377 VSS.n5311 VSS.n5306 0.0242837
R26378 VSS.n5310 VSS.n5307 0.0242837
R26379 DVSS VSS.n4084 0.0241842
R26380 VSS.n5036 VSS.n4408 0.024
R26381 VSS.n4961 VSS.n4960 0.024
R26382 VSS.n4726 VSS.n4724 0.024
R26383 VSS.n4804 VSS.n4512 0.024
R26384 VSS.n5057 VSS.n5056 0.0235
R26385 VSS.n4551 VSS.n4550 0.0235
R26386 VSS.n4704 VSS.n4377 0.0235
R26387 VSS.n4825 VSS.n4824 0.0235
R26388 VSS.n4638 VSS.n4393 0.0231108
R26389 VSS.n4718 VSS.n4639 0.0231108
R26390 VSS.n5108 VSS.n4303 0.023
R26391 VSS.n5077 VSS.n4353 0.023
R26392 VSS.n4918 VSS.n4573 0.023
R26393 VSS.n4886 VSS.n4622 0.023
R26394 VSS.n4654 VSS.n4305 0.023
R26395 VSS.n4678 VSS.n4350 0.023
R26396 VSS.n4846 VSS.n4575 0.023
R26397 VSS.n4870 VSS.n4619 0.023
R26398 VSS.n4392 DVSS 0.0228892
R26399 VSS.n4711 DVSS 0.0228892
R26400 VSS.n3018 VSS.n2905 0.0227936
R26401 VSS.n3357 VSS.n2912 0.0227859
R26402 VSS.n2935 VSS.n2918 0.0227859
R26403 VSS.n2946 VSS.n2944 0.0227859
R26404 VSS.n3319 VSS.n2961 0.0227859
R26405 VSS.n3141 VSS.n3093 0.0227859
R26406 VSS.n2947 VSS.n2946 0.0227859
R26407 VSS.n2963 VSS.n2961 0.0227859
R26408 VSS.n3136 VSS.n3096 0.0227859
R26409 VSS.n2916 VSS.n2913 0.0227859
R26410 VSS.n3359 VSS.n2908 0.0227859
R26411 VSS.n3545 VSS.n2881 0.0227554
R26412 VSS.n3539 VSS.n2878 0.0227554
R26413 VSS.n669 VSS.n668 0.0226946
R26414 VSS.n5100 VSS.n4320 0.0225
R26415 VSS.n5085 VSS.n4336 0.0225
R26416 VSS.n4910 VSS.n4587 0.0225
R26417 VSS.n4894 VSS.n4603 0.0225
R26418 VSS.n4661 VSS.n4659 0.0225
R26419 VSS.n4673 VSS.n4672 0.0225
R26420 VSS.n4853 VSS.n4851 0.0225
R26421 VSS.n4865 VSS.n4864 0.0225
R26422 VSS.n5439 VSS.n1287 0.0224253
R26423 VSS.n5446 VSS.n1287 0.0224253
R26424 VSS.n5447 VSS.n5446 0.0224253
R26425 VSS.n5448 VSS.n5447 0.0224253
R26426 VSS.n5448 VSS.n1283 0.0224253
R26427 VSS.n5454 VSS.n1283 0.0224253
R26428 VSS.n5455 VSS.n5454 0.0224253
R26429 VSS.n5456 VSS.n5455 0.0224253
R26430 VSS.n5456 VSS.n1279 0.0224253
R26431 VSS.n5462 VSS.n1279 0.0224253
R26432 VSS.n5463 VSS.n5462 0.0224253
R26433 VSS.n5464 VSS.n5463 0.0224253
R26434 VSS.n5464 VSS.n1275 0.0224253
R26435 VSS.n5470 VSS.n1275 0.0224253
R26436 VSS.n5471 VSS.n5470 0.0224253
R26437 VSS.n5472 VSS.n5471 0.0224253
R26438 VSS.n5472 VSS.n1271 0.0224253
R26439 VSS.n5478 VSS.n1271 0.0224253
R26440 VSS.n5479 VSS.n5478 0.0224253
R26441 VSS.n5480 VSS.n5479 0.0224253
R26442 VSS.n5480 VSS.n1267 0.0224253
R26443 VSS.n5486 VSS.n1267 0.0224253
R26444 VSS.n5487 VSS.n5486 0.0224253
R26445 VSS.n5488 VSS.n5487 0.0224253
R26446 VSS.n5488 VSS.n1263 0.0224253
R26447 VSS.n5494 VSS.n1263 0.0224253
R26448 VSS.n5495 VSS.n5494 0.0224253
R26449 VSS.n5496 VSS.n5495 0.0224253
R26450 VSS.n5496 VSS.n1259 0.0224253
R26451 VSS.n5502 VSS.n1259 0.0224253
R26452 VSS.n5503 VSS.n5502 0.0224253
R26453 VSS.n5504 VSS.n5503 0.0224253
R26454 VSS.n5504 VSS.n1255 0.0224253
R26455 VSS.n5510 VSS.n1255 0.0224253
R26456 VSS.n5511 VSS.n5510 0.0224253
R26457 VSS.n5512 VSS.n5511 0.0224253
R26458 VSS.n5512 VSS.n1251 0.0224253
R26459 VSS.n5518 VSS.n1251 0.0224253
R26460 VSS.n5519 VSS.n5518 0.0224253
R26461 VSS.n5520 VSS.n5519 0.0224253
R26462 VSS.n5520 VSS.n1247 0.0224253
R26463 VSS.n5526 VSS.n1247 0.0224253
R26464 VSS.n5527 VSS.n5526 0.0224253
R26465 VSS.n5528 VSS.n5527 0.0224253
R26466 VSS.n5528 VSS.n1243 0.0224253
R26467 VSS.n5534 VSS.n1243 0.0224253
R26468 VSS.n5535 VSS.n5534 0.0224253
R26469 VSS.n5536 VSS.n5535 0.0224253
R26470 VSS.n5536 VSS.n1239 0.0224253
R26471 VSS.n5542 VSS.n1239 0.0224253
R26472 VSS.n5543 VSS.n5542 0.0224253
R26473 VSS.n5544 VSS.n5543 0.0224253
R26474 VSS.n5544 VSS.n1235 0.0224253
R26475 VSS.n5550 VSS.n1235 0.0224253
R26476 VSS.n5551 VSS.n5550 0.0224253
R26477 VSS.n5553 VSS.n5551 0.0224253
R26478 VSS.n5553 VSS.n5552 0.0224253
R26479 VSS.n5561 VSS.n5560 0.0224253
R26480 VSS.n5562 VSS.n5561 0.0224253
R26481 VSS.n5562 VSS.n1227 0.0224253
R26482 VSS.n5568 VSS.n1227 0.0224253
R26483 VSS.n5569 VSS.n5568 0.0224253
R26484 VSS.n5570 VSS.n5569 0.0224253
R26485 VSS.n5570 VSS.n1223 0.0224253
R26486 VSS.n5576 VSS.n1223 0.0224253
R26487 VSS.n5577 VSS.n5576 0.0224253
R26488 VSS.n5578 VSS.n5577 0.0224253
R26489 VSS.n5578 VSS.n1219 0.0224253
R26490 VSS.n5584 VSS.n1219 0.0224253
R26491 VSS.n5585 VSS.n5584 0.0224253
R26492 VSS.n5586 VSS.n5585 0.0224253
R26493 VSS.n5586 VSS.n1215 0.0224253
R26494 VSS.n5592 VSS.n1215 0.0224253
R26495 VSS.n5593 VSS.n5592 0.0224253
R26496 VSS.n5594 VSS.n5593 0.0224253
R26497 VSS.n5594 VSS.n1211 0.0224253
R26498 VSS.n5600 VSS.n1211 0.0224253
R26499 VSS.n5601 VSS.n5600 0.0224253
R26500 VSS.n5602 VSS.n5601 0.0224253
R26501 VSS.n5602 VSS.n1207 0.0224253
R26502 VSS.n5608 VSS.n1207 0.0224253
R26503 VSS.n5609 VSS.n5608 0.0224253
R26504 VSS.n5610 VSS.n5609 0.0224253
R26505 VSS.n5610 VSS.n1203 0.0224253
R26506 VSS.n5616 VSS.n1203 0.0224253
R26507 VSS.n5617 VSS.n5616 0.0224253
R26508 VSS.n5618 VSS.n5617 0.0224253
R26509 VSS.n5618 VSS.n1199 0.0224253
R26510 VSS.n5624 VSS.n1199 0.0224253
R26511 VSS.n5625 VSS.n5624 0.0224253
R26512 VSS.n5626 VSS.n5625 0.0224253
R26513 VSS.n5626 VSS.n1195 0.0224253
R26514 VSS.n5632 VSS.n1195 0.0224253
R26515 VSS.n5633 VSS.n5632 0.0224253
R26516 VSS.n5634 VSS.n5633 0.0224253
R26517 VSS.n5634 VSS.n1191 0.0224253
R26518 VSS.n5640 VSS.n1191 0.0224253
R26519 VSS.n5641 VSS.n5640 0.0224253
R26520 VSS.n5642 VSS.n5641 0.0224253
R26521 VSS.n5642 VSS.n1187 0.0224253
R26522 VSS.n5648 VSS.n1187 0.0224253
R26523 VSS.n5649 VSS.n5648 0.0224253
R26524 VSS.n5650 VSS.n5649 0.0224253
R26525 VSS.n5650 VSS.n1183 0.0224253
R26526 VSS.n5656 VSS.n1183 0.0224253
R26527 VSS.n5657 VSS.n5656 0.0224253
R26528 VSS.n5658 VSS.n5657 0.0224253
R26529 VSS.n5658 VSS.n1179 0.0224253
R26530 VSS.n5664 VSS.n1179 0.0224253
R26531 VSS.n5665 VSS.n5664 0.0224253
R26532 VSS.n5666 VSS.n5665 0.0224253
R26533 VSS.n5666 VSS.n1175 0.0224253
R26534 VSS.n5672 VSS.n1175 0.0224253
R26535 VSS.n5673 VSS.n5672 0.0224253
R26536 VSS.n5674 VSS.n5673 0.0224253
R26537 VSS.n3275 VSS.n3252 0.0223919
R26538 VSS.n3273 VSS.n3252 0.0223919
R26539 VSS.n3014 VSS.n2907 0.0223919
R26540 VSS.n3272 VSS.n3247 0.0223919
R26541 VSS.n3274 VSS.n3272 0.0223919
R26542 VSS.n3018 VSS.n3017 0.0223807
R26543 VSS.n3019 VSS.n3018 0.0223807
R26544 VSS.n4908 VSS.n4907 0.0222241
R26545 VSS.n4855 VSS.n4627 0.0222241
R26546 VSS.n4371 VSS.n4370 0.022
R26547 VSS.n4932 VSS.n4931 0.022
R26548 VSS.n4698 VSS.n4697 0.022
R26549 VSS.n4831 VSS.n4557 0.022
R26550 VSS.n5406 VSS.n5405 0.0216765
R26551 VSS.n3321 VSS.n2962 0.021555
R26552 VSS.n3355 VSS.n2911 0.021555
R26553 VSS.n906 VSS.n905 0.0215113
R26554 VSS.n5044 VSS.n4394 0.0215
R26555 VSS.n4532 VSS.n4520 0.0215
R26556 VSS.n4719 VSS.n4396 0.0215
R26557 VSS.n4811 VSS.n4810 0.0215
R26558 VSS.n3639 VSS.n3548 0.021288
R26559 VSS.n3537 VSS.n2877 0.021288
R26560 VSS.n3272 VSS.n3271 0.0211757
R26561 VSS.n3014 VSS.n3013 0.0211757
R26562 VSS.n3337 VSS.n3336 0.0211422
R26563 VSS.n5021 VSS.n4424 0.021
R26564 VSS.n4973 VSS.n4497 0.021
R26565 VSS.n4739 VSS.n4738 0.021
R26566 VSS.n4788 VSS.n4494 0.021
R26567 VSS.n3322 VSS.n3321 0.02075
R26568 VSS.n3321 VSS.n3320 0.02075
R26569 VSS.n3336 VSS.n2945 0.02075
R26570 VSS.n3336 VSS.n3335 0.02075
R26571 VSS.n5010 VSS.n4446 0.0206724
R26572 VSS.n4749 VSS.n4748 0.0206724
R26573 VSS.n666 VSS.n221 0.0206158
R26574 VSS.n4461 VSS.n4460 0.0205
R26575 VSS.n4996 VSS.n4462 0.0205
R26576 VSS.n4765 VSS.n4764 0.0205
R26577 VSS.n4770 VSS.n4768 0.0205
R26578 VSS.n5074 VSS.n4357 0.0204507
R26579 VSS.n4682 VSS.n4681 0.0204507
R26580 VSS.n4444 DVSS 0.0202291
R26581 VSS.n4741 DVSS 0.0202291
R26582 VSS.n911 VSS.n910 0.020197
R26583 VSS.n4441 VSS.n4429 0.02
R26584 VSS.n4980 VSS.n4484 0.02
R26585 VSS.n4743 VSS.n4742 0.02
R26586 VSS.n4786 VSS.n4486 0.02
R26587 VSS.n3251 VSS.n3248 0.0199037
R26588 VSS.n3361 VSS.n2906 0.0199037
R26589 VSS.n5687 VSS.n5686 0.0195912
R26590 VSS.n5686 VSS.n5685 0.0195912
R26591 VSS.n5685 VSS.n5684 0.0195912
R26592 VSS.n1149 VSS.n1148 0.0195912
R26593 VSS.n1148 VSS.n1147 0.0195912
R26594 VSS.n1147 VSS.n1146 0.0195912
R26595 VSS.n5037 VSS.n4407 0.0195
R26596 VSS.n4957 VSS.n4515 0.0195
R26597 VSS.n4721 VSS.n4404 0.0195
R26598 VSS.n4807 VSS.n4806 0.0195
R26599 VSS.n216 VSS.n215 0.0191284
R26600 VSS.n3119 VSS.n3118 0.019078
R26601 VSS.n3341 VSS.n3340 0.019078
R26602 VSS.n5060 VSS.n4372 0.019
R26603 VSS.n4936 VSS.n4935 0.019
R26604 VSS.n4703 VSS.n4701 0.019
R26605 VSS.n4828 VSS.n4548 0.019
R26606 DVSS VSS.n4607 0.018899
R26607 VSS.n4867 DVSS 0.018899
R26608 VSS.n4319 VSS.n4318 0.0185
R26609 VSS.n4352 VSS.n4340 0.0185
R26610 VSS.n4586 VSS.n4585 0.0185
R26611 VSS.n4621 VSS.n4608 0.0185
R26612 VSS.n4656 VSS.n4655 0.0185
R26613 VSS.n4677 VSS.n4676 0.0185
R26614 VSS.n4848 VSS.n4847 0.0185
R26615 VSS.n4869 VSS.n4868 0.0185
R26616 VSS.n1397 VSS.n1395 0.018166
R26617 VSS.n5101 VSS.n4319 0.018
R26618 VSS.n5084 VSS.n4340 0.018
R26619 VSS.n4911 VSS.n4586 0.018
R26620 VSS.n4893 VSS.n4608 0.018
R26621 VSS.n4656 VSS.n4316 0.018
R26622 VSS.n4676 VSS.n4342 0.018
R26623 VSS.n4848 VSS.n4583 0.018
R26624 VSS.n4868 VSS.n4610 0.018
R26625 VSS.n2911 VSS.n2906 0.0178394
R26626 VSS.n4645 VSS.n4301 0.0177906
R26627 VSS.n4653 VSS.n4646 0.0177906
R26628 VSS.n2074 VSS.n2066 0.0176
R26629 VSS.n1820 VSS.n1819 0.0176
R26630 VSS.n4482 DVSS 0.017569
R26631 VSS.n4778 DVSS 0.017569
R26632 VSS.n5061 VSS.n5060 0.0175
R26633 VSS.n4935 VSS.n4552 0.0175
R26634 VSS.n4701 VSS.n4368 0.0175
R26635 VSS.n4830 VSS.n4828 0.0175
R26636 VSS.n3294 VSS.n3293 0.0174266
R26637 VSS.n536 VSS.n535 0.0174005
R26638 VSS.n1818 VSS.n1811 0.0172066
R26639 VSS.n2311 VSS.n9 0.0171667
R26640 VSS.n5126 VSS.n9 0.0171667
R26641 VSS.n1231 VSS.n10 0.0171667
R26642 VSS.n5557 VSS.n10 0.0171667
R26643 VSS.n3024 VSS.n3023 0.0170138
R26644 VSS.n4407 VSS.n4406 0.017
R26645 VSS.n4957 VSS.n4956 0.017
R26646 VSS.n4721 VSS.n4720 0.017
R26647 VSS.n4807 VSS.n4522 0.017
R26648 VSS.n2470 VSS.n2461 0.0169185
R26649 VSS.n2470 VSS.n2469 0.0169185
R26650 VSS.n2698 VSS.n2472 0.0169185
R26651 VSS.n2472 VSS.n2471 0.0169185
R26652 VSS.n2699 VSS.n2474 0.0169185
R26653 VSS.n2474 VSS.n2473 0.0169185
R26654 VSS.n2700 VSS.n2476 0.0169185
R26655 VSS.n2476 VSS.n2475 0.0169185
R26656 VSS.n4055 VSS.n2702 0.0169185
R26657 VSS.n4042 VSS.n4041 0.0169185
R26658 VSS.n4040 VSS.n4039 0.0169185
R26659 VSS.n4038 VSS.n4037 0.0169185
R26660 VSS.n4037 VSS.n4036 0.0169185
R26661 VSS.n4035 VSS.n4034 0.0169185
R26662 VSS.n4032 VSS.n4031 0.0169185
R26663 VSS.n4031 VSS.n4030 0.0169185
R26664 VSS.n4028 VSS.n4027 0.0169185
R26665 VSS.n1602 VSS.n1596 0.0169185
R26666 VSS.n1604 VSS.n1602 0.0169185
R26667 VSS.n1612 VSS.n1601 0.0169185
R26668 VSS.n1606 VSS.n1601 0.0169185
R26669 VSS.n1611 VSS.n1600 0.0169185
R26670 VSS.n1608 VSS.n1600 0.0169185
R26671 VSS.n1610 VSS.n1599 0.0169185
R26672 VSS.n2063 VSS.n1599 0.0169185
R26673 VSS.n2066 VSS.n1596 0.0169185
R26674 VSS.n1605 VSS.n1604 0.0169185
R26675 VSS.n1612 VSS.n1605 0.0169185
R26676 VSS.n1607 VSS.n1606 0.0169185
R26677 VSS.n1611 VSS.n1607 0.0169185
R26678 VSS.n1609 VSS.n1608 0.0169185
R26679 VSS.n1610 VSS.n1609 0.0169185
R26680 VSS.n2064 VSS.n2063 0.0169185
R26681 VSS.n1807 VSS.n1796 0.0169185
R26682 VSS.n1808 VSS.n1806 0.0169185
R26683 VSS.n1804 VSS.n1795 0.0169185
R26684 VSS.n1805 VSS.n1803 0.0169185
R26685 VSS.n1801 VSS.n1794 0.0169185
R26686 VSS.n1802 VSS.n1800 0.0169185
R26687 VSS.n1799 VSS.n1793 0.0169185
R26688 VSS.n1856 VSS.n1855 0.0169185
R26689 VSS.n1820 VSS.n1796 0.0169185
R26690 VSS.n1808 VSS.n1807 0.0169185
R26691 VSS.n1806 VSS.n1795 0.0169185
R26692 VSS.n1805 VSS.n1804 0.0169185
R26693 VSS.n1803 VSS.n1794 0.0169185
R26694 VSS.n1802 VSS.n1801 0.0169185
R26695 VSS.n1800 VSS.n1793 0.0169185
R26696 VSS.n1855 VSS.n1799 0.0169185
R26697 VSS.n4185 VSS.n4184 0.0169185
R26698 VSS.n4183 VSS.n4181 0.0169185
R26699 VSS.n4183 VSS.n4182 0.0169185
R26700 VSS.n4180 VSS.n4178 0.0169185
R26701 VSS.n4180 VSS.n4179 0.0169185
R26702 VSS.n4177 VSS.n4175 0.0169185
R26703 VSS.n4177 VSS.n4176 0.0169185
R26704 VSS.n4174 VSS.n4172 0.0169185
R26705 VSS.n4174 VSS.n4173 0.0169185
R26706 VSS.n4173 VSS.n2413 0.0169185
R26707 VSS.n4176 VSS.n2412 0.0169185
R26708 VSS.n4172 VSS.n2412 0.0169185
R26709 VSS.n4179 VSS.n2411 0.0169185
R26710 VSS.n4175 VSS.n2411 0.0169185
R26711 VSS.n4182 VSS.n2410 0.0169185
R26712 VSS.n4178 VSS.n2410 0.0169185
R26713 VSS.n4184 VSS.n2409 0.0169185
R26714 VSS.n4181 VSS.n2409 0.0169185
R26715 VSS.n4057 VSS.n2461 0.0169185
R26716 VSS.n2469 VSS.n2467 0.0169185
R26717 VSS.n2698 VSS.n2467 0.0169185
R26718 VSS.n2471 VSS.n2466 0.0169185
R26719 VSS.n2699 VSS.n2466 0.0169185
R26720 VSS.n2473 VSS.n2465 0.0169185
R26721 VSS.n2700 VSS.n2465 0.0169185
R26722 VSS.n2475 VSS.n2464 0.0169185
R26723 VSS.n2702 VSS.n2464 0.0169185
R26724 VSS.n4043 VSS.n4042 0.0169185
R26725 VSS.n4041 VSS.n4040 0.0169185
R26726 VSS.n4039 VSS.n4038 0.0169185
R26727 VSS.n4036 VSS.n4035 0.0169185
R26728 VSS.n4034 VSS.n4033 0.0169185
R26729 VSS.n4033 VSS.n4032 0.0169185
R26730 VSS.n4030 VSS.n4029 0.0169185
R26731 VSS.n4029 VSS.n4028 0.0169185
R26732 VSS.n3267 VSS.n3266 0.0167162
R26733 VSS.n908 VSS.n907 0.0166994
R26734 VSS.n909 VSS.n908 0.0166994
R26735 VSS.n5020 VSS.n4429 0.0165
R26736 VSS.n4496 VSS.n4484 0.0165
R26737 VSS.n4742 VSS.n4431 0.0165
R26738 VSS.n4787 VSS.n4786 0.0165
R26739 VSS.n4922 DVSS 0.0162389
R26740 VSS.n4838 DVSS 0.0162389
R26741 VSS.n4997 VSS.n4461 0.016
R26742 VSS.n4997 VSS.n4996 0.016
R26743 VSS.n4765 VSS.n4458 0.016
R26744 VSS.n4768 VSS.n4458 0.016
R26745 VSS.n5021 VSS.n5020 0.0155
R26746 VSS.n4497 VSS.n4496 0.0155
R26747 VSS.n4739 VSS.n4431 0.0155
R26748 VSS.n4788 VSS.n4787 0.0155
R26749 VSS.n5157 VSS.n5156 0.0154891
R26750 VSS.n2074 VSS.n1595 0.01535
R26751 VSS.n1819 VSS.n1797 0.01535
R26752 VSS.n3006 VSS.n3004 0.0152819
R26753 VSS.n3006 VSS.n3005 0.0152819
R26754 VSS.n3008 VSS.n2976 0.0152819
R26755 VSS.n3004 VSS.n2921 0.0152819
R26756 VSS.n3005 VSS.n2978 0.0152819
R26757 VSS.n2978 VSS.n2976 0.0152819
R26758 VSS.n3306 VSS.n3304 0.0152819
R26759 VSS.n3306 VSS.n3305 0.0152819
R26760 VSS.n3308 VSS.n3075 0.0152819
R26761 VSS.n3304 VSS.n3079 0.0152819
R26762 VSS.n3305 VSS.n3078 0.0152819
R26763 VSS.n3078 VSS.n3075 0.0152819
R26764 VSS.n635 VSS.n220 0.0152727
R26765 VSS.n4406 VSS.n4394 0.015
R26766 VSS.n4956 VSS.n4520 0.015
R26767 VSS.n4720 VSS.n4719 0.015
R26768 VSS.n4810 VSS.n4522 0.015
R26769 VSS.n3362 VSS.n2905 0.0149495
R26770 VSS.n4535 DVSS 0.0149089
R26771 VSS.n4809 DVSS 0.0149089
R26772 VSS.n2072 VSS.n1592 0.0149069
R26773 VSS.n2071 VSS.n2070 0.0149069
R26774 VSS.n2071 VSS.n1593 0.0149069
R26775 VSS.n2068 VSS.n1593 0.0149069
R26776 VSS.n2067 VSS.n1592 0.0149069
R26777 VSS.n2070 VSS.n2067 0.0149069
R26778 VSS.n1816 VSS.n1815 0.0149069
R26779 VSS.n1814 VSS.n1813 0.0149069
R26780 VSS.n1812 VSS.n1810 0.0149069
R26781 VSS.n1813 VSS.n1812 0.0149069
R26782 VSS.n1815 VSS.n1814 0.0149069
R26783 VSS.n1817 VSS.n1816 0.0149069
R26784 VSS.n5693 VSS.n17 0.0145462
R26785 VSS.n1151 VSS.n17 0.0145462
R26786 VSS.n1153 VSS.n1151 0.0145462
R26787 VSS.n1155 VSS.n1153 0.0145462
R26788 VSS.n1156 VSS.n1155 0.0145462
R26789 VSS.n1159 VSS.n1156 0.0145462
R26790 VSS.n1161 VSS.n1159 0.0145462
R26791 VSS.n1163 VSS.n1161 0.0145462
R26792 VSS.n1164 VSS.n1163 0.0145462
R26793 VSS.n1167 VSS.n1164 0.0145462
R26794 VSS.n1168 VSS.n1167 0.0145462
R26795 VSS.n3028 VSS.n3010 0.0145367
R26796 VSS.n5061 VSS.n4371 0.0145
R26797 VSS.n4932 VSS.n4552 0.0145
R26798 VSS.n4698 VSS.n4368 0.0145
R26799 VSS.n4831 VSS.n4830 0.0145
R26800 VSS.n3548 VSS.n2879 0.0144402
R26801 VSS.n3537 VSS.n2882 0.0144402
R26802 VSS.n1302 VSS.n1300 0.0144028
R26803 VSS.n3184 VSS.n3183 0.0142903
R26804 VSS.n5176 VSS.n5175 0.0142903
R26805 VSS.n3262 VSS.n3255 0.0142838
R26806 VSS.n3582 VSS.n3581 0.0142814
R26807 VSS.n3050 VSS.n3048 0.0141679
R26808 VSS.n3051 VSS.n2887 0.0141679
R26809 VSS.n3051 VSS.n3048 0.0141679
R26810 VSS.n3053 VSS.n3050 0.0141679
R26811 VSS.n5101 VSS.n5100 0.014
R26812 VSS.n5085 VSS.n5084 0.014
R26813 VSS.n4911 VSS.n4910 0.014
R26814 VSS.n4894 VSS.n4893 0.014
R26815 VSS.n4659 VSS.n4316 0.014
R26816 VSS.n4673 VSS.n4342 0.014
R26817 VSS.n4851 VSS.n4583 0.014
R26818 VSS.n4865 VSS.n4610 0.014
R26819 VSS.n1150 VSS.n21 0.0136707
R26820 VSS.n1158 VSS.n1157 0.0136707
R26821 VSS.n1166 VSS.n1165 0.0136707
R26822 VSS.n4958 DVSS 0.0135788
R26823 DVSS VSS.n4808 0.0135788
R26824 VSS.n2068 VSS.n1595 0.01355
R26825 VSS.n1810 VSS.n1797 0.01355
R26826 VSS.n3733 VSS.n2816 0.0135392
R26827 VSS.n4318 VSS.n4303 0.0135
R26828 VSS.n4353 VSS.n4352 0.0135
R26829 VSS.n4585 VSS.n4573 0.0135
R26830 VSS.n4622 VSS.n4621 0.0135
R26831 VSS.n4655 VSS.n4654 0.0135
R26832 VSS.n4678 VSS.n4677 0.0135
R26833 VSS.n4847 VSS.n4846 0.0135
R26834 VSS.n4870 VSS.n4869 0.0135
R26835 VSS.n3030 VSS.n3009 0.0134255
R26836 VSS.n3056 VSS.n3009 0.0134255
R26837 VSS.n3260 VSS.n3257 0.0134255
R26838 VSS.n3259 VSS.n3257 0.0134255
R26839 VSS.n3046 VSS.n3045 0.0133402
R26840 VSS.n3036 VSS.n3035 0.0133402
R26841 VSS.n5057 VSS.n4372 0.013
R26842 VSS.n4936 VSS.n4551 0.013
R26843 VSS.n4704 VSS.n4703 0.013
R26844 VSS.n4825 VSS.n4548 0.013
R26845 VSS.n3042 VSS.n2835 0.0129835
R26846 VSS.n3038 VSS.n2829 0.0129835
R26847 VSS.n3545 VSS.n2879 0.0129728
R26848 VSS.n3539 VSS.n2882 0.0129728
R26849 VSS.n183 VSS.n104 0.0129415
R26850 VSS.n183 VSS.n182 0.0129415
R26851 VSS.n187 VSS.n182 0.0129415
R26852 VSS.n188 VSS.n187 0.0129415
R26853 VSS.n189 VSS.n188 0.0129415
R26854 VSS.n189 VSS.n180 0.0129415
R26855 VSS.n193 VSS.n180 0.0129415
R26856 VSS.n194 VSS.n193 0.0129415
R26857 VSS.n195 VSS.n194 0.0129415
R26858 VSS.n195 VSS.n178 0.0129415
R26859 VSS.n199 VSS.n178 0.0129415
R26860 VSS.n200 VSS.n199 0.0129415
R26861 VSS.n201 VSS.n200 0.0129415
R26862 VSS.n201 VSS.n176 0.0129415
R26863 VSS.n205 VSS.n176 0.0129415
R26864 VSS.n206 VSS.n205 0.0129415
R26865 VSS.n207 VSS.n206 0.0129415
R26866 VSS.n207 VSS.n174 0.0129415
R26867 VSS.n211 VSS.n174 0.0129415
R26868 VSS.n212 VSS.n211 0.0129415
R26869 VSS.n213 VSS.n212 0.0129415
R26870 VSS.n213 VSS.n172 0.0129415
R26871 VSS.n913 VSS.n912 0.0129415
R26872 VSS.n235 VSS.n218 0.0129415
R26873 VSS.n236 VSS.n235 0.0129415
R26874 VSS.n237 VSS.n236 0.0129415
R26875 VSS.n237 VSS.n231 0.0129415
R26876 VSS.n241 VSS.n231 0.0129415
R26877 VSS.n242 VSS.n241 0.0129415
R26878 VSS.n243 VSS.n242 0.0129415
R26879 VSS.n243 VSS.n229 0.0129415
R26880 VSS.n247 VSS.n229 0.0129415
R26881 VSS.n248 VSS.n247 0.0129415
R26882 VSS.n249 VSS.n248 0.0129415
R26883 VSS.n249 VSS.n227 0.0129415
R26884 VSS.n253 VSS.n227 0.0129415
R26885 VSS.n254 VSS.n253 0.0129415
R26886 VSS.n255 VSS.n254 0.0129415
R26887 VSS.n255 VSS.n225 0.0129415
R26888 VSS.n259 VSS.n225 0.0129415
R26889 VSS.n260 VSS.n259 0.0129415
R26890 VSS.n261 VSS.n260 0.0129415
R26891 VSS.n261 VSS.n223 0.0129415
R26892 VSS.n905 VSS.n223 0.0129415
R26893 VSS.n378 VSS.n373 0.0127609
R26894 VSS.n379 VSS.n377 0.0127609
R26895 VSS.n376 VSS.n374 0.0127528
R26896 VSS.n3358 VSS.n2911 0.01265
R26897 VSS.n2984 VSS.n2911 0.01265
R26898 VSS.n5037 VSS.n5036 0.0125
R26899 VSS.n4960 VSS.n4515 0.0125
R26900 VSS.n4724 VSS.n4404 0.0125
R26901 VSS.n4806 VSS.n4804 0.0125
R26902 VSS.n3131 VSS.n3130 0.0124725
R26903 VSS.n2941 VSS.n2940 0.0124725
R26904 VSS.n569 VSS.n568 0.0123471
R26905 VSS.n568 VSS.n567 0.0123471
R26906 VSS.n567 VSS.n525 0.0123471
R26907 VSS.n563 VSS.n525 0.0123471
R26908 VSS.n563 VSS.n562 0.0123471
R26909 VSS.n562 VSS.n561 0.0123471
R26910 VSS.n561 VSS.n527 0.0123471
R26911 VSS.n557 VSS.n527 0.0123471
R26912 VSS.n557 VSS.n556 0.0123471
R26913 VSS.n556 VSS.n555 0.0123471
R26914 VSS.n555 VSS.n529 0.0123471
R26915 VSS.n551 VSS.n529 0.0123471
R26916 VSS.n551 VSS.n550 0.0123471
R26917 VSS.n550 VSS.n549 0.0123471
R26918 VSS.n549 VSS.n531 0.0123471
R26919 VSS.n545 VSS.n531 0.0123471
R26920 VSS.n545 VSS.n544 0.0123471
R26921 VSS.n544 VSS.n543 0.0123471
R26922 VSS.n543 VSS.n533 0.0123471
R26923 VSS.n539 VSS.n533 0.0123471
R26924 VSS.n539 VSS.n538 0.0123471
R26925 VSS.n538 VSS.n537 0.0123471
R26926 VSS.n634 VSS.n633 0.0123471
R26927 VSS.n636 VSS.n363 0.0123471
R26928 VSS.n640 VSS.n363 0.0123471
R26929 VSS.n641 VSS.n640 0.0123471
R26930 VSS.n642 VSS.n641 0.0123471
R26931 VSS.n642 VSS.n361 0.0123471
R26932 VSS.n646 VSS.n361 0.0123471
R26933 VSS.n647 VSS.n646 0.0123471
R26934 VSS.n648 VSS.n647 0.0123471
R26935 VSS.n648 VSS.n359 0.0123471
R26936 VSS.n652 VSS.n359 0.0123471
R26937 VSS.n653 VSS.n652 0.0123471
R26938 VSS.n654 VSS.n653 0.0123471
R26939 VSS.n654 VSS.n357 0.0123471
R26940 VSS.n658 VSS.n357 0.0123471
R26941 VSS.n659 VSS.n658 0.0123471
R26942 VSS.n660 VSS.n659 0.0123471
R26943 VSS.n660 VSS.n355 0.0123471
R26944 VSS.n664 VSS.n355 0.0123471
R26945 VSS.n665 VSS.n664 0.0123471
R26946 VSS.n667 VSS.n665 0.0123471
R26947 VSS.n667 VSS.n666 0.0123471
R26948 VSS.n5692 VSS.n5691 0.0123293
R26949 VSS.n31 VSS.n27 0.0123293
R26950 VSS.n3049 VSS.n2832 0.0122701
R26951 VSS.n3714 VSS.n2838 0.0122701
R26952 DVSS VSS.n4921 0.0122488
R26953 DVSS VSS.n4628 0.0122488
R26954 VSS.n4442 VSS.n4441 0.012
R26955 VSS.n4981 VSS.n4980 0.012
R26956 VSS.n4744 VSS.n4743 0.012
R26957 VSS.n4783 VSS.n4486 0.012
R26958 VSS.n3289 VSS.n3288 0.0116468
R26959 VSS.n5560 VSS.n1231 0.0116395
R26960 VSS.n5273 VSS.n2227 0.0116
R26961 VSS.n1154 VSS.n30 0.0115976
R26962 VSS.n1160 VSS.n26 0.0115976
R26963 VSS.n4460 VSS.n4450 0.0115
R26964 VSS.n4993 VSS.n4462 0.0115
R26965 VSS.n4764 VSS.n4763 0.0115
R26966 VSS.n4771 VSS.n4770 0.0115
R26967 VSS.n3354 VSS.n2915 0.0113969
R26968 VSS.n3354 VSS.n3353 0.0113969
R26969 VSS.n3140 VSS.n3139 0.0113969
R26970 VSS.n3139 VSS.n3138 0.0113969
R26971 VSS.n5552 VSS.n1231 0.0112859
R26972 VSS.n1771 VSS.n1769 0.0112561
R26973 VSS.n1785 VSS.n1775 0.0112561
R26974 VSS.n1918 VSS.n1917 0.0112561
R26975 VSS.n1901 VSS.n1898 0.0112561
R26976 VSS.n1956 VSS.n1955 0.0112561
R26977 VSS.n1939 VSS.n1936 0.0112561
R26978 VSS.n1987 VSS.n1677 0.0112561
R26979 VSS.n1976 VSS.n1686 0.0112561
R26980 VSS.n2019 VSS.n1650 0.0112561
R26981 VSS.n2008 VSS.n1661 0.0112561
R26982 VSS.n1627 VSS.n1625 0.0112561
R26983 VSS.n1641 VSS.n1631 0.0112561
R26984 VSS.n5298 VSS 0.0110882
R26985 VSS VSS.n5296 0.0110882
R26986 VSS.n4048 VSS 0.0110882
R26987 VSS.n5024 VSS.n4424 0.011
R26988 VSS.n4973 VSS.n4972 0.011
R26989 VSS.n4738 VSS.n4736 0.011
R26990 VSS.n4792 VSS.n4494 0.011
R26991 VSS.n3512 VSS.n3511 0.0109694
R26992 VSS.n3513 VSS.n3512 0.0109694
R26993 VSS.n3513 VSS.n3388 0.0109694
R26994 VSS.n3519 VSS.n3388 0.0109694
R26995 VSS.n3520 VSS.n3519 0.0109694
R26996 VSS.n3521 VSS.n3520 0.0109694
R26997 VSS.n3521 VSS.n2198 0.0109694
R26998 VSS.n5285 VSS.n2198 0.0109694
R26999 VSS.n5285 VSS.n5284 0.0109694
R27000 DVSS VSS.n4481 0.0109187
R27001 VSS.n4775 DVSS 0.0109187
R27002 VSS.n5273 VSS.n5272 0.0109
R27003 VSS.n5272 VSS.n5267 0.0109
R27004 VSS.n5267 VSS.n5266 0.0109
R27005 VSS.n5266 VSS.n5265 0.0109
R27006 VSS.n5265 VSS.n5264 0.0109
R27007 VSS.n5264 VSS.n5263 0.0109
R27008 VSS.n5263 VSS.n5262 0.0109
R27009 VSS.n5262 VSS.n5261 0.0109
R27010 VSS.n5261 VSS.n5260 0.0109
R27011 VSS.n5260 VSS.n5259 0.0109
R27012 VSS.n5259 VSS.n5258 0.0109
R27013 VSS.n1152 VSS.n29 0.0108659
R27014 VSS.n1162 VSS.n24 0.0108659
R27015 VSS.n4645 VSS.n4321 0.010697
R27016 VSS.n4657 VSS.n4646 0.010697
R27017 VSS.n4310 VSS.n4309 0.0105
R27018 VSS.n4310 VSS.n4307 0.0105
R27019 VSS.n5105 VSS.n4307 0.0105
R27020 VSS.n5105 VSS.n5104 0.0105
R27021 VSS.n5104 VSS.n4315 0.0105
R27022 VSS.n4327 VSS.n4315 0.0105
R27023 VSS.n5093 VSS.n4327 0.0105
R27024 VSS.n5093 VSS.n5092 0.0105
R27025 VSS.n5092 VSS.n4332 0.0105
R27026 VSS.n4344 VSS.n4332 0.0105
R27027 VSS.n5081 VSS.n4344 0.0105
R27028 VSS.n5081 VSS.n5080 0.0105
R27029 VSS.n5080 VSS.n4349 0.0105
R27030 VSS.n4689 VSS.n4349 0.0105
R27031 VSS.n4689 VSS.n4364 0.0105
R27032 VSS.n5065 VSS.n4364 0.0105
R27033 VSS.n5065 VSS.n5064 0.0105
R27034 VSS.n5064 VSS.n4367 0.0105
R27035 VSS.n4379 VSS.n4367 0.0105
R27036 VSS.n5053 VSS.n4379 0.0105
R27037 VSS.n5053 VSS.n5052 0.0105
R27038 VSS.n5052 VSS.n4384 0.0105
R27039 VSS.n4398 VSS.n4384 0.0105
R27040 VSS.n5041 VSS.n4398 0.0105
R27041 VSS.n5041 VSS.n5040 0.0105
R27042 VSS.n5040 VSS.n4403 0.0105
R27043 VSS.n4415 VSS.n4403 0.0105
R27044 VSS.n5029 VSS.n4415 0.0105
R27045 VSS.n5029 VSS.n5028 0.0105
R27046 VSS.n5028 VSS.n4420 0.0105
R27047 VSS.n4433 VSS.n4420 0.0105
R27048 VSS.n5017 VSS.n4433 0.0105
R27049 VSS.n5017 VSS.n5016 0.0105
R27050 VSS.n5016 VSS.n4438 0.0105
R27051 VSS.n4756 VSS.n4438 0.0105
R27052 VSS.n4756 VSS.n4454 0.0105
R27053 VSS.n5001 VSS.n4454 0.0105
R27054 VSS.n5001 VSS.n5000 0.0105
R27055 VSS.n5000 VSS.n4457 0.0105
R27056 VSS.n4469 VSS.n4457 0.0105
R27057 VSS.n4989 VSS.n4469 0.0105
R27058 VSS.n4989 VSS.n4988 0.0105
R27059 VSS.n4988 VSS.n4474 0.0105
R27060 VSS.n4488 VSS.n4474 0.0105
R27061 VSS.n4977 VSS.n4488 0.0105
R27062 VSS.n4977 VSS.n4976 0.0105
R27063 VSS.n4976 VSS.n4493 0.0105
R27064 VSS.n4506 VSS.n4493 0.0105
R27065 VSS.n4965 VSS.n4506 0.0105
R27066 VSS.n4965 VSS.n4964 0.0105
R27067 VSS.n4964 VSS.n4511 0.0105
R27068 VSS.n4524 VSS.n4511 0.0105
R27069 VSS.n4953 VSS.n4524 0.0105
R27070 VSS.n4953 VSS.n4952 0.0105
R27071 VSS.n4952 VSS.n4529 0.0105
R27072 VSS.n4542 VSS.n4529 0.0105
R27073 VSS.n4940 VSS.n4542 0.0105
R27074 VSS.n4940 VSS.n4939 0.0105
R27075 VSS.n4939 VSS.n4547 0.0105
R27076 VSS.n4559 VSS.n4547 0.0105
R27077 VSS.n4928 VSS.n4559 0.0105
R27078 VSS.n4928 VSS.n4927 0.0105
R27079 VSS.n4927 VSS.n4564 0.0105
R27080 VSS.n4577 VSS.n4564 0.0105
R27081 VSS.n4915 VSS.n4577 0.0105
R27082 VSS.n4915 VSS.n4914 0.0105
R27083 VSS.n4914 VSS.n4582 0.0105
R27084 VSS.n4594 VSS.n4582 0.0105
R27085 VSS.n4902 VSS.n4594 0.0105
R27086 VSS.n4902 VSS.n4901 0.0105
R27087 VSS.n4901 VSS.n4599 0.0105
R27088 VSS.n4612 VSS.n4599 0.0105
R27089 VSS.n4890 VSS.n4612 0.0105
R27090 VSS.n4890 VSS.n4889 0.0105
R27091 VSS.n4889 VSS.n4618 0.0105
R27092 VSS.n4618 VSS.n2279 0.0105
R27093 VSS.n5135 VSS.n2279 0.0105
R27094 VSS.n5135 VSS.n2277 0.0105
R27095 VSS.n5139 VSS.n2277 0.0105
R27096 VSS.n5139 VSS.n2275 0.0105
R27097 VSS.n5143 VSS.n2275 0.0105
R27098 VSS.n5143 VSS.n2273 0.0105
R27099 VSS.n5167 VSS.n2273 0.0105
R27100 VSS.n5167 VSS.n5166 0.0105
R27101 VSS.n5166 VSS.n5165 0.0105
R27102 VSS.n5165 VSS.n5149 0.0105
R27103 VSS.n5161 VSS.n5149 0.0105
R27104 VSS.n5161 VSS.n5160 0.0105
R27105 VSS.n5160 VSS.n5159 0.0105
R27106 VSS.n5045 VSS.n5044 0.0105
R27107 VSS.n4533 VSS.n4532 0.0105
R27108 VSS.n4716 VSS.n4396 0.0105
R27109 VSS.n4812 VSS.n4811 0.0105
R27110 VSS.n5140 VSS.n2276 0.0105
R27111 VSS.n5141 VSS.n5140 0.0105
R27112 VSS.n5142 VSS.n5141 0.0105
R27113 VSS.n5142 VSS.n2271 0.0105
R27114 VSS.n5168 VSS.n2272 0.0105
R27115 VSS.n5164 VSS.n2272 0.0105
R27116 VSS.n5164 VSS.n5163 0.0105
R27117 VSS.n5163 VSS.n5162 0.0105
R27118 VSS.n5162 VSS.n5150 0.0105
R27119 VSS.n5158 VSS.n5150 0.0105
R27120 VSS.n5169 VSS.n5168 0.0104296
R27121 VSS.n1772 VSS.n1771 0.0101185
R27122 VSS.n1786 VSS.n1785 0.0101185
R27123 VSS.n1918 VSS.n1726 0.0101185
R27124 VSS.n1903 VSS.n1898 0.0101185
R27125 VSS.n1956 VSS.n1702 0.0101185
R27126 VSS.n1941 VSS.n1936 0.0101185
R27127 VSS.n1988 VSS.n1987 0.0101185
R27128 VSS.n1974 VSS.n1686 0.0101185
R27129 VSS.n2020 VSS.n2019 0.0101185
R27130 VSS.n2006 VSS.n1661 0.0101185
R27131 VSS.n1628 VSS.n1627 0.0101185
R27132 VSS.n1642 VSS.n1641 0.0101185
R27133 VSS.n5683 VSS.n1149 0.0100456
R27134 VSS.n5688 VSS.n5687 0.0100456
R27135 VSS.n5684 VSS.n5683 0.0100456
R27136 VSS.n1146 VSS.n1145 0.0100456
R27137 VSS.n4370 VSS.n4360 0.01
R27138 VSS.n4931 VSS.n4555 0.01
R27139 VSS.n4697 VSS.n4696 0.01
R27140 VSS.n4834 VSS.n4557 0.01
R27141 VSS.n4090 DVSS 0.00997368
R27142 VSS.n3052 VSS.n2831 0.00965456
R27143 VSS.n3032 VSS.n2837 0.00965456
R27144 VSS.n2315 VSS.n2310 0.00962857
R27145 VSS.n2319 VSS.n2310 0.00962857
R27146 VSS.n2319 VSS.n2308 0.00962857
R27147 VSS.n2323 VSS.n2308 0.00962857
R27148 VSS.n2323 VSS.n2306 0.00962857
R27149 VSS.n2327 VSS.n2306 0.00962857
R27150 VSS.n2327 VSS.n2304 0.00962857
R27151 VSS.n2331 VSS.n2304 0.00962857
R27152 VSS.n2331 VSS.n2302 0.00962857
R27153 VSS.n2335 VSS.n2302 0.00962857
R27154 VSS.n2335 VSS.n2299 0.00962857
R27155 VSS.n4280 VSS.n2299 0.00962857
R27156 VSS.n4280 VSS.n2300 0.00962857
R27157 VSS.n4276 VSS.n2300 0.00962857
R27158 VSS.n4276 VSS.n2339 0.00962857
R27159 VSS.n4272 VSS.n2339 0.00962857
R27160 VSS.n4272 VSS.n2341 0.00962857
R27161 VSS.n4268 VSS.n2341 0.00962857
R27162 VSS.n4268 VSS.n2343 0.00962857
R27163 VSS.n4264 VSS.n2343 0.00962857
R27164 VSS.n4264 VSS.n2345 0.00962857
R27165 VSS.n4260 VSS.n2345 0.00962857
R27166 VSS.n4260 VSS.n2347 0.00962857
R27167 VSS.n4256 VSS.n2347 0.00962857
R27168 VSS.n4256 VSS.n2349 0.00962857
R27169 VSS.n4252 VSS.n2349 0.00962857
R27170 VSS.n4252 VSS.n2351 0.00962857
R27171 VSS.n2546 VSS.n2351 0.00962857
R27172 VSS.n2549 VSS.n2546 0.00962857
R27173 VSS.n2549 VSS.n2544 0.00962857
R27174 VSS.n2553 VSS.n2544 0.00962857
R27175 VSS.n2553 VSS.n2542 0.00962857
R27176 VSS.n2557 VSS.n2542 0.00962857
R27177 VSS.n2557 VSS.n2540 0.00962857
R27178 VSS.n2561 VSS.n2540 0.00962857
R27179 VSS.n2561 VSS.n2538 0.00962857
R27180 VSS.n2565 VSS.n2538 0.00962857
R27181 VSS.n2565 VSS.n2536 0.00962857
R27182 VSS.n2569 VSS.n2536 0.00962857
R27183 VSS.n2569 VSS.n2534 0.00962857
R27184 VSS.n2573 VSS.n2534 0.00962857
R27185 VSS.n2573 VSS.n2532 0.00962857
R27186 VSS.n2577 VSS.n2532 0.00962857
R27187 VSS.n2577 VSS.n2530 0.00962857
R27188 VSS.n2581 VSS.n2530 0.00962857
R27189 VSS.n2581 VSS.n2528 0.00962857
R27190 VSS.n2585 VSS.n2528 0.00962857
R27191 VSS.n2585 VSS.n2526 0.00962857
R27192 VSS.n2589 VSS.n2526 0.00962857
R27193 VSS.n2589 VSS.n2524 0.00962857
R27194 VSS.n2593 VSS.n2524 0.00962857
R27195 VSS.n2593 VSS.n2522 0.00962857
R27196 VSS.n2597 VSS.n2522 0.00962857
R27197 VSS.n2597 VSS.n2520 0.00962857
R27198 VSS.n2601 VSS.n2520 0.00962857
R27199 VSS.n2601 VSS.n2518 0.00962857
R27200 VSS.n2605 VSS.n2518 0.00962857
R27201 VSS.n2605 VSS.n2516 0.00962857
R27202 VSS.n2609 VSS.n2516 0.00962857
R27203 VSS.n2609 VSS.n2514 0.00962857
R27204 VSS.n2613 VSS.n2514 0.00962857
R27205 VSS.n2613 VSS.n2512 0.00962857
R27206 VSS.n2617 VSS.n2512 0.00962857
R27207 VSS.n2617 VSS.n2510 0.00962857
R27208 VSS.n2621 VSS.n2510 0.00962857
R27209 VSS.n2621 VSS.n2508 0.00962857
R27210 VSS.n2625 VSS.n2508 0.00962857
R27211 VSS.n2625 VSS.n2506 0.00962857
R27212 VSS.n2629 VSS.n2506 0.00962857
R27213 VSS.n2629 VSS.n2504 0.00962857
R27214 VSS.n2633 VSS.n2504 0.00962857
R27215 VSS.n2633 VSS.n2502 0.00962857
R27216 VSS.n2637 VSS.n2502 0.00962857
R27217 VSS.n2637 VSS.n2500 0.00962857
R27218 VSS.n2641 VSS.n2500 0.00962857
R27219 VSS.n2641 VSS.n2498 0.00962857
R27220 VSS.n2645 VSS.n2498 0.00962857
R27221 VSS.n2645 VSS.n2496 0.00962857
R27222 VSS.n2649 VSS.n2496 0.00962857
R27223 VSS.n2649 VSS.n2494 0.00962857
R27224 VSS.n2653 VSS.n2494 0.00962857
R27225 VSS.n2653 VSS.n2492 0.00962857
R27226 VSS.n2657 VSS.n2492 0.00962857
R27227 VSS.n2657 VSS.n2490 0.00962857
R27228 VSS.n2661 VSS.n2490 0.00962857
R27229 VSS.n2661 VSS.n2488 0.00962857
R27230 VSS.n2665 VSS.n2488 0.00962857
R27231 VSS.n2665 VSS.n2486 0.00962857
R27232 VSS.n2669 VSS.n2486 0.00962857
R27233 VSS.n2669 VSS.n2484 0.00962857
R27234 VSS.n2673 VSS.n2484 0.00962857
R27235 VSS.n2673 VSS.n2482 0.00962857
R27236 VSS.n2678 VSS.n2482 0.00962857
R27237 VSS.n2678 VSS.n2479 0.00962857
R27238 VSS.n2682 VSS.n2479 0.00962857
R27239 VSS.n2683 VSS.n2682 0.00962857
R27240 VSS.n2684 VSS.n2683 0.00962857
R27241 VSS.n2696 VSS.n2477 0.00962857
R27242 VSS.n2692 VSS.n2477 0.00962857
R27243 VSS.n2692 VSS.n2687 0.00962857
R27244 VSS.n3378 VSS.n3377 0.00962857
R27245 VSS.n3377 VSS.n2895 0.00962857
R27246 VSS.n3373 VSS.n2895 0.00962857
R27247 VSS.n3373 VSS.n2897 0.00962857
R27248 VSS.n3369 VSS.n2897 0.00962857
R27249 VSS.n3369 VSS.n2900 0.00962857
R27250 VSS.n3365 VSS.n2900 0.00962857
R27251 VSS.n3365 VSS.n2902 0.00962857
R27252 VSS.n2988 VSS.n2902 0.00962857
R27253 VSS.n2991 VSS.n2988 0.00962857
R27254 VSS.n2991 VSS.n2982 0.00962857
R27255 VSS.n2997 VSS.n2982 0.00962857
R27256 VSS.n2997 VSS.n2980 0.00962857
R27257 VSS.n3001 VSS.n2980 0.00962857
R27258 VSS.n3001 VSS.n2925 0.00962857
R27259 VSS.n3348 VSS.n2925 0.00962857
R27260 VSS.n3348 VSS.n2926 0.00962857
R27261 VSS.n3344 VSS.n2926 0.00962857
R27262 VSS.n3344 VSS.n2929 0.00962857
R27263 VSS.n3063 VSS.n2929 0.00962857
R27264 VSS.n3063 VSS.n2952 0.00962857
R27265 VSS.n3330 VSS.n2952 0.00962857
R27266 VSS.n3330 VSS.n2953 0.00962857
R27267 VSS.n3326 VSS.n2953 0.00962857
R27268 VSS.n3326 VSS.n2956 0.00962857
R27269 VSS.n3106 VSS.n2956 0.00962857
R27270 VSS.n3122 VSS.n3106 0.00962857
R27271 VSS.n3122 VSS.n3102 0.00962857
R27272 VSS.n3127 VSS.n3102 0.00962857
R27273 VSS.n3127 VSS.n3104 0.00962857
R27274 VSS.n3104 VSS.n3083 0.00962857
R27275 VSS.n3301 VSS.n3083 0.00962857
R27276 VSS.n3301 VSS.n3084 0.00962857
R27277 VSS.n3297 VSS.n3084 0.00962857
R27278 VSS.n3297 VSS.n3087 0.00962857
R27279 VSS.n3148 VSS.n3087 0.00962857
R27280 VSS.n3285 VSS.n3148 0.00962857
R27281 VSS.n3285 VSS.n3149 0.00962857
R27282 VSS.n3281 VSS.n3149 0.00962857
R27283 VSS.n3281 VSS.n3152 0.00962857
R27284 VSS.n3243 VSS.n3152 0.00962857
R27285 VSS.n3243 VSS.n3156 0.00962857
R27286 VSS.n3239 VSS.n3156 0.00962857
R27287 VSS.n3239 VSS.n3158 0.00962857
R27288 VSS.n3235 VSS.n3158 0.00962857
R27289 VSS.n3235 VSS.n3160 0.00962857
R27290 VSS.n3231 VSS.n3160 0.00962857
R27291 VSS.n3231 VSS.n3162 0.00962857
R27292 VSS.n3227 VSS.n3162 0.00962857
R27293 VSS.n3227 VSS.n3164 0.00962857
R27294 VSS.n3223 VSS.n3164 0.00962857
R27295 VSS.n3223 VSS.n3166 0.00962857
R27296 VSS.n3219 VSS.n3166 0.00962857
R27297 VSS.n3219 VSS.n3168 0.00962857
R27298 VSS.n3215 VSS.n3168 0.00962857
R27299 VSS.n3215 VSS.n3170 0.00962857
R27300 VSS.n3211 VSS.n3170 0.00962857
R27301 VSS.n3211 VSS.n3172 0.00962857
R27302 VSS.n3207 VSS.n3172 0.00962857
R27303 VSS.n3207 VSS.n3174 0.00962857
R27304 VSS.n3203 VSS.n3174 0.00962857
R27305 VSS.n3203 VSS.n3176 0.00962857
R27306 VSS.n3199 VSS.n3176 0.00962857
R27307 VSS.n3199 VSS.n3178 0.00962857
R27308 VSS.n3195 VSS.n3178 0.00962857
R27309 VSS.n3195 VSS.n3180 0.00962857
R27310 VSS.n3191 VSS.n3180 0.00962857
R27311 VSS.n3191 VSS.n3182 0.00962857
R27312 VSS.n3187 VSS.n3182 0.00962857
R27313 VSS.n3726 VSS.n3725 0.00962857
R27314 VSS.n3725 VSS.n2820 0.00962857
R27315 VSS.n3721 VSS.n2820 0.00962857
R27316 VSS.n3721 VSS.n2823 0.00962857
R27317 VSS.n3717 VSS.n2823 0.00962857
R27318 VSS.n3717 VSS.n2826 0.00962857
R27319 VSS.n3711 VSS.n2826 0.00962857
R27320 VSS.n3711 VSS.n2841 0.00962857
R27321 VSS.n3707 VSS.n2841 0.00962857
R27322 VSS.n3707 VSS.n2843 0.00962857
R27323 VSS.n3703 VSS.n2843 0.00962857
R27324 VSS.n3703 VSS.n2845 0.00962857
R27325 VSS.n3699 VSS.n2845 0.00962857
R27326 VSS.n3699 VSS.n2847 0.00962857
R27327 VSS.n3695 VSS.n2847 0.00962857
R27328 VSS.n3695 VSS.n2849 0.00962857
R27329 VSS.n3691 VSS.n2849 0.00962857
R27330 VSS.n3691 VSS.n2851 0.00962857
R27331 VSS.n3687 VSS.n2851 0.00962857
R27332 VSS.n3687 VSS.n2853 0.00962857
R27333 VSS.n3683 VSS.n2853 0.00962857
R27334 VSS.n3683 VSS.n2855 0.00962857
R27335 VSS.n3679 VSS.n2855 0.00962857
R27336 VSS.n3679 VSS.n2857 0.00962857
R27337 VSS.n3675 VSS.n2857 0.00962857
R27338 VSS.n3675 VSS.n2859 0.00962857
R27339 VSS.n3671 VSS.n2859 0.00962857
R27340 VSS.n3671 VSS.n2861 0.00962857
R27341 VSS.n3667 VSS.n2861 0.00962857
R27342 VSS.n3667 VSS.n2863 0.00962857
R27343 VSS.n3663 VSS.n2863 0.00962857
R27344 VSS.n3663 VSS.n2865 0.00962857
R27345 VSS.n3659 VSS.n2865 0.00962857
R27346 VSS.n3659 VSS.n2867 0.00962857
R27347 VSS.n3655 VSS.n2867 0.00962857
R27348 VSS.n3655 VSS.n2869 0.00962857
R27349 VSS.n3651 VSS.n2869 0.00962857
R27350 VSS.n3651 VSS.n2871 0.00962857
R27351 VSS.n3647 VSS.n2871 0.00962857
R27352 VSS.n3647 VSS.n2873 0.00962857
R27353 VSS.n3643 VSS.n2873 0.00962857
R27354 VSS.n3643 VSS.n2875 0.00962857
R27355 VSS.n3553 VSS.n2875 0.00962857
R27356 VSS.n3553 VSS.n3551 0.00962857
R27357 VSS.n3636 VSS.n3551 0.00962857
R27358 VSS.n3636 VSS.n3552 0.00962857
R27359 VSS.n3632 VSS.n3552 0.00962857
R27360 VSS.n3632 VSS.n3557 0.00962857
R27361 VSS.n3628 VSS.n3557 0.00962857
R27362 VSS.n3628 VSS.n3559 0.00962857
R27363 VSS.n3624 VSS.n3559 0.00962857
R27364 VSS.n3624 VSS.n3561 0.00962857
R27365 VSS.n3620 VSS.n3561 0.00962857
R27366 VSS.n3620 VSS.n3563 0.00962857
R27367 VSS.n3616 VSS.n3563 0.00962857
R27368 VSS.n3616 VSS.n3565 0.00962857
R27369 VSS.n3612 VSS.n3565 0.00962857
R27370 VSS.n3612 VSS.n3567 0.00962857
R27371 VSS.n3608 VSS.n3567 0.00962857
R27372 VSS.n3608 VSS.n3569 0.00962857
R27373 VSS.n3604 VSS.n3569 0.00962857
R27374 VSS.n3604 VSS.n3571 0.00962857
R27375 VSS.n3600 VSS.n3571 0.00962857
R27376 VSS.n3600 VSS.n3573 0.00962857
R27377 VSS.n3596 VSS.n3573 0.00962857
R27378 VSS.n3596 VSS.n3575 0.00962857
R27379 VSS.n3592 VSS.n3575 0.00962857
R27380 VSS.n3592 VSS.n3577 0.00962857
R27381 VSS.n3588 VSS.n3577 0.00962857
R27382 VSS.n3588 VSS.n3579 0.00962857
R27383 VSS.n3584 VSS.n3579 0.00962857
R27384 VSS.n3724 VSS.n3723 0.00962857
R27385 VSS.n3723 VSS.n3722 0.00962857
R27386 VSS.n3722 VSS.n2822 0.00962857
R27387 VSS.n3712 VSS.n2840 0.00962857
R27388 VSS.n3706 VSS.n2840 0.00962857
R27389 VSS.n3706 VSS.n3705 0.00962857
R27390 VSS.n3705 VSS.n3704 0.00962857
R27391 VSS.n3704 VSS.n2844 0.00962857
R27392 VSS.n3698 VSS.n2844 0.00962857
R27393 VSS.n3698 VSS.n3697 0.00962857
R27394 VSS.n3697 VSS.n3696 0.00962857
R27395 VSS.n3696 VSS.n2848 0.00962857
R27396 VSS.n3690 VSS.n2848 0.00962857
R27397 VSS.n3690 VSS.n3689 0.00962857
R27398 VSS.n3689 VSS.n3688 0.00962857
R27399 VSS.n3688 VSS.n2852 0.00962857
R27400 VSS.n3682 VSS.n2852 0.00962857
R27401 VSS.n3682 VSS.n3681 0.00962857
R27402 VSS.n3681 VSS.n3680 0.00962857
R27403 VSS.n3680 VSS.n2856 0.00962857
R27404 VSS.n3674 VSS.n2856 0.00962857
R27405 VSS.n3674 VSS.n3673 0.00962857
R27406 VSS.n3673 VSS.n3672 0.00962857
R27407 VSS.n3672 VSS.n2860 0.00962857
R27408 VSS.n3666 VSS.n2860 0.00962857
R27409 VSS.n3666 VSS.n3665 0.00962857
R27410 VSS.n3665 VSS.n3664 0.00962857
R27411 VSS.n3664 VSS.n2864 0.00962857
R27412 VSS.n3658 VSS.n2864 0.00962857
R27413 VSS.n3658 VSS.n3657 0.00962857
R27414 VSS.n3657 VSS.n3656 0.00962857
R27415 VSS.n3656 VSS.n2868 0.00962857
R27416 VSS.n3650 VSS.n2868 0.00962857
R27417 VSS.n3650 VSS.n3649 0.00962857
R27418 VSS.n3649 VSS.n3648 0.00962857
R27419 VSS.n3648 VSS.n2872 0.00962857
R27420 VSS.n3642 VSS.n2872 0.00962857
R27421 VSS.n3642 VSS.n3641 0.00962857
R27422 VSS.n3637 VSS.n3550 0.00962857
R27423 VSS.n3631 VSS.n3550 0.00962857
R27424 VSS.n3631 VSS.n3630 0.00962857
R27425 VSS.n3630 VSS.n3629 0.00962857
R27426 VSS.n3629 VSS.n3558 0.00962857
R27427 VSS.n3623 VSS.n3558 0.00962857
R27428 VSS.n3623 VSS.n3622 0.00962857
R27429 VSS.n3622 VSS.n3621 0.00962857
R27430 VSS.n3621 VSS.n3562 0.00962857
R27431 VSS.n3615 VSS.n3562 0.00962857
R27432 VSS.n3615 VSS.n3614 0.00962857
R27433 VSS.n3614 VSS.n3613 0.00962857
R27434 VSS.n3613 VSS.n3566 0.00962857
R27435 VSS.n3607 VSS.n3566 0.00962857
R27436 VSS.n3607 VSS.n3606 0.00962857
R27437 VSS.n3606 VSS.n3605 0.00962857
R27438 VSS.n3605 VSS.n3570 0.00962857
R27439 VSS.n3599 VSS.n3570 0.00962857
R27440 VSS.n3599 VSS.n3598 0.00962857
R27441 VSS.n3598 VSS.n3597 0.00962857
R27442 VSS.n3597 VSS.n3574 0.00962857
R27443 VSS.n3591 VSS.n3574 0.00962857
R27444 VSS.n3591 VSS.n3590 0.00962857
R27445 VSS.n3590 VSS.n3589 0.00962857
R27446 VSS.n3589 VSS.n3578 0.00962857
R27447 VSS.n3583 VSS.n3578 0.00962857
R27448 VSS.n2060 VSS.n1613 0.00962857
R27449 VSS.n2060 VSS.n1614 0.00962857
R27450 VSS.n2056 VSS.n1614 0.00962857
R27451 VSS.n2056 VSS.n1616 0.00962857
R27452 VSS.n2052 VSS.n1616 0.00962857
R27453 VSS.n2052 VSS.n1619 0.00962857
R27454 VSS.n2048 VSS.n1619 0.00962857
R27455 VSS.n2048 VSS.n1621 0.00962857
R27456 VSS.n1635 VSS.n1621 0.00962857
R27457 VSS.n2036 VSS.n1635 0.00962857
R27458 VSS.n2036 VSS.n1636 0.00962857
R27459 VSS.n2032 VSS.n1636 0.00962857
R27460 VSS.n2032 VSS.n1639 0.00962857
R27461 VSS.n2028 VSS.n1639 0.00962857
R27462 VSS.n2028 VSS.n1645 0.00962857
R27463 VSS.n2024 VSS.n1645 0.00962857
R27464 VSS.n2024 VSS.n1647 0.00962857
R27465 VSS.n1652 VSS.n1647 0.00962857
R27466 VSS.n2016 VSS.n1652 0.00962857
R27467 VSS.n2016 VSS.n1653 0.00962857
R27468 VSS.n2012 VSS.n1653 0.00962857
R27469 VSS.n2012 VSS.n1656 0.00962857
R27470 VSS.n1666 VSS.n1656 0.00962857
R27471 VSS.n2003 VSS.n1666 0.00962857
R27472 VSS.n2003 VSS.n1667 0.00962857
R27473 VSS.n1999 VSS.n1667 0.00962857
R27474 VSS.n1999 VSS.n1670 0.00962857
R27475 VSS.n1995 VSS.n1670 0.00962857
R27476 VSS.n1995 VSS.n1672 0.00962857
R27477 VSS.n1991 VSS.n1672 0.00962857
R27478 VSS.n1991 VSS.n1674 0.00962857
R27479 VSS.n1984 VSS.n1674 0.00962857
R27480 VSS.n1984 VSS.n1679 0.00962857
R27481 VSS.n1980 VSS.n1679 0.00962857
R27482 VSS.n1980 VSS.n1681 0.00962857
R27483 VSS.n1691 VSS.n1681 0.00962857
R27484 VSS.n1971 VSS.n1691 0.00962857
R27485 VSS.n1971 VSS.n1692 0.00962857
R27486 VSS.n1967 VSS.n1692 0.00962857
R27487 VSS.n1967 VSS.n1695 0.00962857
R27488 VSS.n1963 VSS.n1695 0.00962857
R27489 VSS.n1963 VSS.n1697 0.00962857
R27490 VSS.n1959 VSS.n1697 0.00962857
R27491 VSS.n1959 VSS.n1699 0.00962857
R27492 VSS.n1709 VSS.n1699 0.00962857
R27493 VSS.n1948 VSS.n1709 0.00962857
R27494 VSS.n1948 VSS.n1710 0.00962857
R27495 VSS.n1944 VSS.n1710 0.00962857
R27496 VSS.n1944 VSS.n1713 0.00962857
R27497 VSS.n1933 VSS.n1713 0.00962857
R27498 VSS.n1933 VSS.n1717 0.00962857
R27499 VSS.n1929 VSS.n1717 0.00962857
R27500 VSS.n1929 VSS.n1719 0.00962857
R27501 VSS.n1925 VSS.n1719 0.00962857
R27502 VSS.n1925 VSS.n1721 0.00962857
R27503 VSS.n1921 VSS.n1721 0.00962857
R27504 VSS.n1921 VSS.n1723 0.00962857
R27505 VSS.n1751 VSS.n1723 0.00962857
R27506 VSS.n1910 VSS.n1751 0.00962857
R27507 VSS.n1910 VSS.n1752 0.00962857
R27508 VSS.n1906 VSS.n1752 0.00962857
R27509 VSS.n1906 VSS.n1755 0.00962857
R27510 VSS.n1895 VSS.n1755 0.00962857
R27511 VSS.n1895 VSS.n1759 0.00962857
R27512 VSS.n1891 VSS.n1759 0.00962857
R27513 VSS.n1891 VSS.n1761 0.00962857
R27514 VSS.n1887 VSS.n1761 0.00962857
R27515 VSS.n1887 VSS.n1763 0.00962857
R27516 VSS.n1883 VSS.n1763 0.00962857
R27517 VSS.n1883 VSS.n1765 0.00962857
R27518 VSS.n1779 VSS.n1765 0.00962857
R27519 VSS.n1871 VSS.n1779 0.00962857
R27520 VSS.n1871 VSS.n1780 0.00962857
R27521 VSS.n1867 VSS.n1780 0.00962857
R27522 VSS.n1867 VSS.n1783 0.00962857
R27523 VSS.n1863 VSS.n1783 0.00962857
R27524 VSS.n1863 VSS.n1789 0.00962857
R27525 VSS.n1859 VSS.n1789 0.00962857
R27526 VSS.n1859 VSS.n1791 0.00962857
R27527 VSS.n1852 VSS.n1791 0.00962857
R27528 VSS.n1852 VSS.n1822 0.00962857
R27529 VSS.n1848 VSS.n1822 0.00962857
R27530 VSS.n1848 VSS.n1824 0.00962857
R27531 VSS.n1844 VSS.n1824 0.00962857
R27532 VSS.n1844 VSS.n1826 0.00962857
R27533 VSS.n1840 VSS.n1826 0.00962857
R27534 VSS.n1839 VSS.n1827 0.00962857
R27535 VSS.n1834 VSS.n1827 0.00962857
R27536 VSS.n1834 VSS.n1830 0.00962857
R27537 VSS.n2055 VSS.n1617 0.00962857
R27538 VSS.n2055 VSS.n2054 0.00962857
R27539 VSS.n2054 VSS.n2053 0.00962857
R27540 VSS.n2031 VSS.n2030 0.00962857
R27541 VSS.n2030 VSS.n2029 0.00962857
R27542 VSS.n2029 VSS.n1644 0.00962857
R27543 VSS.n2023 VSS.n1644 0.00962857
R27544 VSS.n2023 VSS.n2022 0.00962857
R27545 VSS.n2004 VSS.n1665 0.00962857
R27546 VSS.n1998 VSS.n1665 0.00962857
R27547 VSS.n1998 VSS.n1997 0.00962857
R27548 VSS.n1997 VSS.n1996 0.00962857
R27549 VSS.n1996 VSS.n1671 0.00962857
R27550 VSS.n1990 VSS.n1671 0.00962857
R27551 VSS.n1972 VSS.n1690 0.00962857
R27552 VSS.n1966 VSS.n1690 0.00962857
R27553 VSS.n1966 VSS.n1965 0.00962857
R27554 VSS.n1965 VSS.n1964 0.00962857
R27555 VSS.n1964 VSS.n1696 0.00962857
R27556 VSS.n1935 VSS.n1934 0.00962857
R27557 VSS.n1934 VSS.n1716 0.00962857
R27558 VSS.n1928 VSS.n1716 0.00962857
R27559 VSS.n1928 VSS.n1927 0.00962857
R27560 VSS.n1927 VSS.n1926 0.00962857
R27561 VSS.n1926 VSS.n1720 0.00962857
R27562 VSS.n1897 VSS.n1896 0.00962857
R27563 VSS.n1896 VSS.n1758 0.00962857
R27564 VSS.n1890 VSS.n1758 0.00962857
R27565 VSS.n1890 VSS.n1889 0.00962857
R27566 VSS.n1889 VSS.n1888 0.00962857
R27567 VSS.n1866 VSS.n1865 0.00962857
R27568 VSS.n1865 VSS.n1864 0.00962857
R27569 VSS.n1864 VSS.n1788 0.00962857
R27570 VSS.n1853 VSS.n1821 0.00962857
R27571 VSS.n1847 VSS.n1821 0.00962857
R27572 VSS.n1847 VSS.n1846 0.00962857
R27573 VSS.n1846 VSS.n1845 0.00962857
R27574 VSS.n1845 VSS.n1825 0.00962857
R27575 VSS.n1825 VSS.n23 0.00962857
R27576 VSS.n1833 VSS.n1831 0.00962857
R27577 VSS.n1833 VSS.n1832 0.00962857
R27578 VSS.n1585 VSS.n1300 0.00962857
R27579 VSS.n1585 VSS.n1301 0.00962857
R27580 VSS.n1581 VSS.n1301 0.00962857
R27581 VSS.n1581 VSS.n1304 0.00962857
R27582 VSS.n1577 VSS.n1304 0.00962857
R27583 VSS.n1577 VSS.n1306 0.00962857
R27584 VSS.n1573 VSS.n1306 0.00962857
R27585 VSS.n1573 VSS.n1308 0.00962857
R27586 VSS.n1569 VSS.n1308 0.00962857
R27587 VSS.n1569 VSS.n1310 0.00962857
R27588 VSS.n1565 VSS.n1310 0.00962857
R27589 VSS.n1565 VSS.n1312 0.00962857
R27590 VSS.n1561 VSS.n1312 0.00962857
R27591 VSS.n1561 VSS.n1314 0.00962857
R27592 VSS.n1557 VSS.n1314 0.00962857
R27593 VSS.n1557 VSS.n1316 0.00962857
R27594 VSS.n1553 VSS.n1316 0.00962857
R27595 VSS.n1553 VSS.n1318 0.00962857
R27596 VSS.n1549 VSS.n1318 0.00962857
R27597 VSS.n1549 VSS.n1320 0.00962857
R27598 VSS.n1545 VSS.n1320 0.00962857
R27599 VSS.n1545 VSS.n1322 0.00962857
R27600 VSS.n1541 VSS.n1322 0.00962857
R27601 VSS.n1541 VSS.n1324 0.00962857
R27602 VSS.n1537 VSS.n1324 0.00962857
R27603 VSS.n1537 VSS.n1326 0.00962857
R27604 VSS.n1533 VSS.n1326 0.00962857
R27605 VSS.n1533 VSS.n1328 0.00962857
R27606 VSS.n1529 VSS.n1328 0.00962857
R27607 VSS.n1529 VSS.n1330 0.00962857
R27608 VSS.n1525 VSS.n1330 0.00962857
R27609 VSS.n1525 VSS.n1332 0.00962857
R27610 VSS.n1521 VSS.n1332 0.00962857
R27611 VSS.n1521 VSS.n1334 0.00962857
R27612 VSS.n1517 VSS.n1334 0.00962857
R27613 VSS.n1517 VSS.n1336 0.00962857
R27614 VSS.n1513 VSS.n1336 0.00962857
R27615 VSS.n1513 VSS.n1338 0.00962857
R27616 VSS.n1509 VSS.n1338 0.00962857
R27617 VSS.n1509 VSS.n1340 0.00962857
R27618 VSS.n1505 VSS.n1340 0.00962857
R27619 VSS.n1505 VSS.n1342 0.00962857
R27620 VSS.n1501 VSS.n1342 0.00962857
R27621 VSS.n1501 VSS.n1344 0.00962857
R27622 VSS.n1497 VSS.n1344 0.00962857
R27623 VSS.n1497 VSS.n1346 0.00962857
R27624 VSS.n1493 VSS.n1346 0.00962857
R27625 VSS.n1493 VSS.n1348 0.00962857
R27626 VSS.n1489 VSS.n1348 0.00962857
R27627 VSS.n1489 VSS.n1350 0.00962857
R27628 VSS.n1485 VSS.n1350 0.00962857
R27629 VSS.n1485 VSS.n1352 0.00962857
R27630 VSS.n1481 VSS.n1352 0.00962857
R27631 VSS.n1481 VSS.n1354 0.00962857
R27632 VSS.n1477 VSS.n1354 0.00962857
R27633 VSS.n1477 VSS.n1356 0.00962857
R27634 VSS.n1473 VSS.n1356 0.00962857
R27635 VSS.n1473 VSS.n1358 0.00962857
R27636 VSS.n1469 VSS.n1358 0.00962857
R27637 VSS.n1469 VSS.n1360 0.00962857
R27638 VSS.n1465 VSS.n1360 0.00962857
R27639 VSS.n1465 VSS.n1362 0.00962857
R27640 VSS.n1461 VSS.n1362 0.00962857
R27641 VSS.n1461 VSS.n1364 0.00962857
R27642 VSS.n1457 VSS.n1364 0.00962857
R27643 VSS.n1457 VSS.n1366 0.00962857
R27644 VSS.n1453 VSS.n1366 0.00962857
R27645 VSS.n1453 VSS.n1368 0.00962857
R27646 VSS.n1449 VSS.n1368 0.00962857
R27647 VSS.n1449 VSS.n1370 0.00962857
R27648 VSS.n1445 VSS.n1370 0.00962857
R27649 VSS.n1445 VSS.n1372 0.00962857
R27650 VSS.n1441 VSS.n1372 0.00962857
R27651 VSS.n1441 VSS.n1374 0.00962857
R27652 VSS.n1437 VSS.n1374 0.00962857
R27653 VSS.n1437 VSS.n1376 0.00962857
R27654 VSS.n1433 VSS.n1376 0.00962857
R27655 VSS.n1433 VSS.n1378 0.00962857
R27656 VSS.n1429 VSS.n1378 0.00962857
R27657 VSS.n1429 VSS.n1380 0.00962857
R27658 VSS.n1425 VSS.n1380 0.00962857
R27659 VSS.n1425 VSS.n1382 0.00962857
R27660 VSS.n1421 VSS.n1382 0.00962857
R27661 VSS.n1421 VSS.n1384 0.00962857
R27662 VSS.n1417 VSS.n1384 0.00962857
R27663 VSS.n1417 VSS.n1386 0.00962857
R27664 VSS.n1413 VSS.n1386 0.00962857
R27665 VSS.n1413 VSS.n1388 0.00962857
R27666 VSS.n1409 VSS.n1388 0.00962857
R27667 VSS.n1409 VSS.n1390 0.00962857
R27668 VSS.n1405 VSS.n1390 0.00962857
R27669 VSS.n1405 VSS.n1392 0.00962857
R27670 VSS.n1401 VSS.n1392 0.00962857
R27671 VSS.n1401 VSS.n1394 0.00962857
R27672 VSS.n1586 VSS.n1299 0.00962857
R27673 VSS.n1580 VSS.n1299 0.00962857
R27674 VSS.n1580 VSS.n1579 0.00962857
R27675 VSS.n1579 VSS.n1578 0.00962857
R27676 VSS.n1578 VSS.n1305 0.00962857
R27677 VSS.n1572 VSS.n1305 0.00962857
R27678 VSS.n1572 VSS.n1571 0.00962857
R27679 VSS.n1571 VSS.n1570 0.00962857
R27680 VSS.n1570 VSS.n1309 0.00962857
R27681 VSS.n1564 VSS.n1309 0.00962857
R27682 VSS.n1564 VSS.n1563 0.00962857
R27683 VSS.n1563 VSS.n1562 0.00962857
R27684 VSS.n1562 VSS.n1313 0.00962857
R27685 VSS.n1556 VSS.n1313 0.00962857
R27686 VSS.n1556 VSS.n1555 0.00962857
R27687 VSS.n1555 VSS.n1554 0.00962857
R27688 VSS.n1554 VSS.n1317 0.00962857
R27689 VSS.n1548 VSS.n1317 0.00962857
R27690 VSS.n1548 VSS.n1547 0.00962857
R27691 VSS.n1547 VSS.n1546 0.00962857
R27692 VSS.n1546 VSS.n1321 0.00962857
R27693 VSS.n1540 VSS.n1321 0.00962857
R27694 VSS.n1540 VSS.n1539 0.00962857
R27695 VSS.n1539 VSS.n1538 0.00962857
R27696 VSS.n1538 VSS.n1325 0.00962857
R27697 VSS.n1532 VSS.n1325 0.00962857
R27698 VSS.n1532 VSS.n1531 0.00962857
R27699 VSS.n1531 VSS.n1530 0.00962857
R27700 VSS.n1530 VSS.n1329 0.00962857
R27701 VSS.n1524 VSS.n1329 0.00962857
R27702 VSS.n1524 VSS.n1523 0.00962857
R27703 VSS.n1523 VSS.n1522 0.00962857
R27704 VSS.n1522 VSS.n1333 0.00962857
R27705 VSS.n1516 VSS.n1333 0.00962857
R27706 VSS.n1516 VSS.n1515 0.00962857
R27707 VSS.n1515 VSS.n1514 0.00962857
R27708 VSS.n1514 VSS.n1337 0.00962857
R27709 VSS.n1508 VSS.n1337 0.00962857
R27710 VSS.n1508 VSS.n1507 0.00962857
R27711 VSS.n1507 VSS.n1506 0.00962857
R27712 VSS.n1506 VSS.n1341 0.00962857
R27713 VSS.n1500 VSS.n1341 0.00962857
R27714 VSS.n1500 VSS.n1499 0.00962857
R27715 VSS.n1499 VSS.n1498 0.00962857
R27716 VSS.n1498 VSS.n1345 0.00962857
R27717 VSS.n1492 VSS.n1345 0.00962857
R27718 VSS.n1492 VSS.n1491 0.00962857
R27719 VSS.n1491 VSS.n1490 0.00962857
R27720 VSS.n1490 VSS.n1349 0.00962857
R27721 VSS.n1484 VSS.n1349 0.00962857
R27722 VSS.n1484 VSS.n1483 0.00962857
R27723 VSS.n1483 VSS.n1482 0.00962857
R27724 VSS.n1482 VSS.n1353 0.00962857
R27725 VSS.n1476 VSS.n1353 0.00962857
R27726 VSS.n1476 VSS.n1475 0.00962857
R27727 VSS.n1475 VSS.n1474 0.00962857
R27728 VSS.n1474 VSS.n1357 0.00962857
R27729 VSS.n1468 VSS.n1357 0.00962857
R27730 VSS.n1468 VSS.n1467 0.00962857
R27731 VSS.n1467 VSS.n1466 0.00962857
R27732 VSS.n1466 VSS.n1361 0.00962857
R27733 VSS.n1460 VSS.n1361 0.00962857
R27734 VSS.n1460 VSS.n1459 0.00962857
R27735 VSS.n1459 VSS.n1458 0.00962857
R27736 VSS.n1458 VSS.n1365 0.00962857
R27737 VSS.n1452 VSS.n1365 0.00962857
R27738 VSS.n1452 VSS.n1451 0.00962857
R27739 VSS.n1451 VSS.n1450 0.00962857
R27740 VSS.n1450 VSS.n1369 0.00962857
R27741 VSS.n1444 VSS.n1369 0.00962857
R27742 VSS.n1444 VSS.n1443 0.00962857
R27743 VSS.n1443 VSS.n1442 0.00962857
R27744 VSS.n1442 VSS.n1373 0.00962857
R27745 VSS.n1436 VSS.n1373 0.00962857
R27746 VSS.n1436 VSS.n1435 0.00962857
R27747 VSS.n1435 VSS.n1434 0.00962857
R27748 VSS.n1434 VSS.n1377 0.00962857
R27749 VSS.n1428 VSS.n1377 0.00962857
R27750 VSS.n1428 VSS.n1427 0.00962857
R27751 VSS.n1427 VSS.n1426 0.00962857
R27752 VSS.n1426 VSS.n1381 0.00962857
R27753 VSS.n1420 VSS.n1381 0.00962857
R27754 VSS.n1420 VSS.n1419 0.00962857
R27755 VSS.n1419 VSS.n1418 0.00962857
R27756 VSS.n1418 VSS.n1385 0.00962857
R27757 VSS.n1412 VSS.n1385 0.00962857
R27758 VSS.n1412 VSS.n1411 0.00962857
R27759 VSS.n1411 VSS.n1410 0.00962857
R27760 VSS.n1410 VSS.n1389 0.00962857
R27761 VSS.n1404 VSS.n1389 0.00962857
R27762 VSS.n1404 VSS.n1403 0.00962857
R27763 VSS.n1403 VSS.n1402 0.00962857
R27764 VSS.n1402 VSS.n1393 0.00962857
R27765 VSS.n3379 VSS.n2894 0.00962857
R27766 VSS.n3372 VSS.n2898 0.00962857
R27767 VSS.n3372 VSS.n3371 0.00962857
R27768 VSS.n3371 VSS.n3370 0.00962857
R27769 VSS.n3331 VSS.n2951 0.00962857
R27770 VSS.n3325 VSS.n2951 0.00962857
R27771 VSS.n3245 VSS.n3244 0.00962857
R27772 VSS.n3244 VSS.n3155 0.00962857
R27773 VSS.n3238 VSS.n3155 0.00962857
R27774 VSS.n3238 VSS.n3237 0.00962857
R27775 VSS.n3237 VSS.n3236 0.00962857
R27776 VSS.n3236 VSS.n3159 0.00962857
R27777 VSS.n3230 VSS.n3159 0.00962857
R27778 VSS.n3230 VSS.n3229 0.00962857
R27779 VSS.n3229 VSS.n3228 0.00962857
R27780 VSS.n3228 VSS.n3163 0.00962857
R27781 VSS.n3222 VSS.n3163 0.00962857
R27782 VSS.n3222 VSS.n3221 0.00962857
R27783 VSS.n3221 VSS.n3220 0.00962857
R27784 VSS.n3220 VSS.n3167 0.00962857
R27785 VSS.n3214 VSS.n3167 0.00962857
R27786 VSS.n3214 VSS.n3213 0.00962857
R27787 VSS.n3213 VSS.n3212 0.00962857
R27788 VSS.n3212 VSS.n3171 0.00962857
R27789 VSS.n3206 VSS.n3171 0.00962857
R27790 VSS.n3206 VSS.n3205 0.00962857
R27791 VSS.n3205 VSS.n3204 0.00962857
R27792 VSS.n3204 VSS.n3175 0.00962857
R27793 VSS.n3198 VSS.n3175 0.00962857
R27794 VSS.n3198 VSS.n3197 0.00962857
R27795 VSS.n3197 VSS.n3196 0.00962857
R27796 VSS.n3196 VSS.n3179 0.00962857
R27797 VSS.n3190 VSS.n3179 0.00962857
R27798 VSS.n3190 VSS.n3189 0.00962857
R27799 VSS.n3189 VSS.n3188 0.00962857
R27800 VSS.n2379 VSS.n2375 0.00962857
R27801 VSS.n4237 VSS.n2375 0.00962857
R27802 VSS.n4237 VSS.n2376 0.00962857
R27803 VSS.n4233 VSS.n2376 0.00962857
R27804 VSS.n4233 VSS.n2383 0.00962857
R27805 VSS.n4228 VSS.n2383 0.00962857
R27806 VSS.n4228 VSS.n2385 0.00962857
R27807 VSS.n4224 VSS.n2385 0.00962857
R27808 VSS.n4224 VSS.n2387 0.00962857
R27809 VSS.n4218 VSS.n2387 0.00962857
R27810 VSS.n4218 VSS.n2389 0.00962857
R27811 VSS.n4214 VSS.n2389 0.00962857
R27812 VSS.n4214 VSS.n2391 0.00962857
R27813 VSS.n4210 VSS.n2391 0.00962857
R27814 VSS.n4210 VSS.n2394 0.00962857
R27815 VSS.n4206 VSS.n2394 0.00962857
R27816 VSS.n4206 VSS.n2396 0.00962857
R27817 VSS.n4200 VSS.n2396 0.00962857
R27818 VSS.n4200 VSS.n2399 0.00962857
R27819 VSS.n4196 VSS.n2399 0.00962857
R27820 VSS.n4196 VSS.n2401 0.00962857
R27821 VSS.n4192 VSS.n2401 0.00962857
R27822 VSS.n4192 VSS.n2404 0.00962857
R27823 VSS.n4188 VSS.n2404 0.00962857
R27824 VSS.n4188 VSS.n2406 0.00962857
R27825 VSS.n4169 VSS.n2406 0.00962857
R27826 VSS.n4169 VSS.n2415 0.00962857
R27827 VSS.n4165 VSS.n2415 0.00962857
R27828 VSS.n4165 VSS.n2417 0.00962857
R27829 VSS.n4161 VSS.n2417 0.00962857
R27830 VSS.n4161 VSS.n2419 0.00962857
R27831 VSS.n4157 VSS.n2419 0.00962857
R27832 VSS.n4157 VSS.n2421 0.00962857
R27833 VSS.n4153 VSS.n2421 0.00962857
R27834 VSS.n4153 VSS.n2423 0.00962857
R27835 VSS.n4149 VSS.n2423 0.00962857
R27836 VSS.n4149 VSS.n2425 0.00962857
R27837 VSS.n4095 VSS.n2425 0.00962857
R27838 VSS.n4100 VSS.n4095 0.00962857
R27839 VSS.n4100 VSS.n4096 0.00962857
R27840 VSS.n4096 VSS.n2442 0.00962857
R27841 VSS.n4109 VSS.n2442 0.00962857
R27842 VSS.n4109 VSS.n2440 0.00962857
R27843 VSS.n4113 VSS.n2440 0.00962857
R27844 VSS.n4113 VSS.n2438 0.00962857
R27845 VSS.n4119 VSS.n2438 0.00962857
R27846 VSS.n4119 VSS.n2435 0.00962857
R27847 VSS.n4137 VSS.n2435 0.00962857
R27848 VSS.n4137 VSS.n2436 0.00962857
R27849 VSS.n4133 VSS.n2436 0.00962857
R27850 VSS.n4133 VSS.n4123 0.00962857
R27851 VSS.n4128 VSS.n4123 0.00962857
R27852 VSS.n4128 VSS.n4125 0.00962857
R27853 VSS.n4125 VSS.n2245 0.00962857
R27854 VSS.n5235 VSS.n2245 0.00962857
R27855 VSS.n5235 VSS.n2246 0.00962857
R27856 VSS.n5231 VSS.n2246 0.00962857
R27857 VSS.n5231 VSS.n2249 0.00962857
R27858 VSS.n5227 VSS.n2249 0.00962857
R27859 VSS.n5227 VSS.n2252 0.00962857
R27860 VSS.n5223 VSS.n2252 0.00962857
R27861 VSS.n5223 VSS.n2254 0.00962857
R27862 VSS.n5219 VSS.n2254 0.00962857
R27863 VSS.n5219 VSS.n2256 0.00962857
R27864 VSS.n5215 VSS.n2256 0.00962857
R27865 VSS.n5215 VSS.n2258 0.00962857
R27866 VSS.n5211 VSS.n2258 0.00962857
R27867 VSS.n5211 VSS.n2260 0.00962857
R27868 VSS.n5207 VSS.n2260 0.00962857
R27869 VSS.n5207 VSS.n2262 0.00962857
R27870 VSS.n5203 VSS.n2262 0.00962857
R27871 VSS.n5203 VSS.n2264 0.00962857
R27872 VSS.n5199 VSS.n2264 0.00962857
R27873 VSS.n5199 VSS.n2266 0.00962857
R27874 VSS.n5195 VSS.n2266 0.00962857
R27875 VSS.n5195 VSS.n2268 0.00962857
R27876 VSS.n5191 VSS.n2268 0.00962857
R27877 VSS.n5191 VSS.n2270 0.00962857
R27878 VSS.n5187 VSS.n2270 0.00962857
R27879 VSS.n5187 VSS.n5172 0.00962857
R27880 VSS.n5183 VSS.n5172 0.00962857
R27881 VSS.n5183 VSS.n5174 0.00962857
R27882 VSS.n5179 VSS.n5174 0.00962857
R27883 VSS.n2378 VSS.n2373 0.00962857
R27884 VSS.n4238 VSS.n2374 0.00962857
R27885 VSS.n4232 VSS.n2374 0.00962857
R27886 VSS.n4230 VSS.n4229 0.00962857
R27887 VSS.n4229 VSS.n2384 0.00962857
R27888 VSS.n4223 VSS.n2384 0.00962857
R27889 VSS.n4213 VSS.n2392 0.00962857
R27890 VSS.n4213 VSS.n4212 0.00962857
R27891 VSS.n4212 VSS.n4211 0.00962857
R27892 VSS.n4205 VSS.n2397 0.00962857
R27893 VSS.n4205 VSS.n4204 0.00962857
R27894 VSS.n4195 VSS.n2402 0.00962857
R27895 VSS.n4195 VSS.n4194 0.00962857
R27896 VSS.n4194 VSS.n4193 0.00962857
R27897 VSS.n4171 VSS.n4170 0.00962857
R27898 VSS.n4170 VSS.n2414 0.00962857
R27899 VSS.n4164 VSS.n2414 0.00962857
R27900 VSS.n4164 VSS.n4163 0.00962857
R27901 VSS.n4163 VSS.n4162 0.00962857
R27902 VSS.n4162 VSS.n2418 0.00962857
R27903 VSS.n4156 VSS.n2418 0.00962857
R27904 VSS.n4156 VSS.n4155 0.00962857
R27905 VSS.n4155 VSS.n4154 0.00962857
R27906 VSS.n4154 VSS.n2422 0.00962857
R27907 VSS.n4148 VSS.n2422 0.00962857
R27908 VSS.n4093 VSS.n2426 0.00962857
R27909 VSS.n4101 VSS.n4094 0.00962857
R27910 VSS.n4094 VSS.n2443 0.00962857
R27911 VSS.n4108 VSS.n2439 0.00962857
R27912 VSS.n4114 VSS.n2439 0.00962857
R27913 VSS.n4115 VSS.n4114 0.00962857
R27914 VSS.n4138 VSS.n2434 0.00962857
R27915 VSS.n4132 VSS.n2434 0.00962857
R27916 VSS.n4132 VSS.n4131 0.00962857
R27917 VSS.n4129 VSS.n4124 0.00962857
R27918 VSS.n4124 VSS.n2243 0.00962857
R27919 VSS.n5230 VSS.n2250 0.00962857
R27920 VSS.n5230 VSS.n5229 0.00962857
R27921 VSS.n5229 VSS.n5228 0.00962857
R27922 VSS.n5228 VSS.n2251 0.00962857
R27923 VSS.n5222 VSS.n2251 0.00962857
R27924 VSS.n5222 VSS.n5221 0.00962857
R27925 VSS.n5221 VSS.n5220 0.00962857
R27926 VSS.n5220 VSS.n2255 0.00962857
R27927 VSS.n5214 VSS.n2255 0.00962857
R27928 VSS.n5214 VSS.n5213 0.00962857
R27929 VSS.n5213 VSS.n5212 0.00962857
R27930 VSS.n5212 VSS.n2259 0.00962857
R27931 VSS.n5206 VSS.n2259 0.00962857
R27932 VSS.n5206 VSS.n5205 0.00962857
R27933 VSS.n5205 VSS.n5204 0.00962857
R27934 VSS.n5204 VSS.n2263 0.00962857
R27935 VSS.n5198 VSS.n2263 0.00962857
R27936 VSS.n5198 VSS.n5197 0.00962857
R27937 VSS.n5197 VSS.n5196 0.00962857
R27938 VSS.n5196 VSS.n2267 0.00962857
R27939 VSS.n5190 VSS.n5189 0.00962857
R27940 VSS.n5189 VSS.n5188 0.00962857
R27941 VSS.n5188 VSS.n5171 0.00962857
R27942 VSS.n5182 VSS.n5171 0.00962857
R27943 VSS.n5182 VSS.n5181 0.00962857
R27944 VSS.n5181 VSS.n5180 0.00962857
R27945 VSS.n2316 VSS.n2313 0.00962857
R27946 VSS.n2317 VSS.n2316 0.00962857
R27947 VSS.n2318 VSS.n2317 0.00962857
R27948 VSS.n2318 VSS.n2307 0.00962857
R27949 VSS.n2324 VSS.n2307 0.00962857
R27950 VSS.n2325 VSS.n2324 0.00962857
R27951 VSS.n2326 VSS.n2325 0.00962857
R27952 VSS.n2326 VSS.n2303 0.00962857
R27953 VSS.n2332 VSS.n2303 0.00962857
R27954 VSS.n2333 VSS.n2332 0.00962857
R27955 VSS.n2334 VSS.n2333 0.00962857
R27956 VSS.n2334 VSS.n2297 0.00962857
R27957 VSS.n4281 VSS.n2298 0.00962857
R27958 VSS.n4275 VSS.n2298 0.00962857
R27959 VSS.n4275 VSS.n4274 0.00962857
R27960 VSS.n4274 VSS.n4273 0.00962857
R27961 VSS.n4273 VSS.n2340 0.00962857
R27962 VSS.n4267 VSS.n2340 0.00962857
R27963 VSS.n4267 VSS.n4266 0.00962857
R27964 VSS.n4266 VSS.n4265 0.00962857
R27965 VSS.n4265 VSS.n2344 0.00962857
R27966 VSS.n4259 VSS.n2344 0.00962857
R27967 VSS.n4259 VSS.n4258 0.00962857
R27968 VSS.n4258 VSS.n4257 0.00962857
R27969 VSS.n4257 VSS.n2348 0.00962857
R27970 VSS.n4251 VSS.n2348 0.00962857
R27971 VSS.n2545 VSS.n2352 0.00962857
R27972 VSS.n2550 VSS.n2545 0.00962857
R27973 VSS.n2551 VSS.n2550 0.00962857
R27974 VSS.n2552 VSS.n2551 0.00962857
R27975 VSS.n2552 VSS.n2541 0.00962857
R27976 VSS.n2558 VSS.n2541 0.00962857
R27977 VSS.n2559 VSS.n2558 0.00962857
R27978 VSS.n2560 VSS.n2559 0.00962857
R27979 VSS.n2560 VSS.n2537 0.00962857
R27980 VSS.n2566 VSS.n2537 0.00962857
R27981 VSS.n2567 VSS.n2566 0.00962857
R27982 VSS.n2568 VSS.n2567 0.00962857
R27983 VSS.n2568 VSS.n2533 0.00962857
R27984 VSS.n2574 VSS.n2533 0.00962857
R27985 VSS.n2575 VSS.n2574 0.00962857
R27986 VSS.n2576 VSS.n2575 0.00962857
R27987 VSS.n2576 VSS.n2529 0.00962857
R27988 VSS.n2582 VSS.n2529 0.00962857
R27989 VSS.n2583 VSS.n2582 0.00962857
R27990 VSS.n2584 VSS.n2583 0.00962857
R27991 VSS.n2584 VSS.n2525 0.00962857
R27992 VSS.n2590 VSS.n2525 0.00962857
R27993 VSS.n2591 VSS.n2590 0.00962857
R27994 VSS.n2592 VSS.n2591 0.00962857
R27995 VSS.n2592 VSS.n2521 0.00962857
R27996 VSS.n2598 VSS.n2521 0.00962857
R27997 VSS.n2599 VSS.n2598 0.00962857
R27998 VSS.n2600 VSS.n2599 0.00962857
R27999 VSS.n2600 VSS.n2517 0.00962857
R28000 VSS.n2606 VSS.n2517 0.00962857
R28001 VSS.n2607 VSS.n2606 0.00962857
R28002 VSS.n2608 VSS.n2607 0.00962857
R28003 VSS.n2608 VSS.n2513 0.00962857
R28004 VSS.n2614 VSS.n2513 0.00962857
R28005 VSS.n2615 VSS.n2614 0.00962857
R28006 VSS.n2616 VSS.n2615 0.00962857
R28007 VSS.n2616 VSS.n2509 0.00962857
R28008 VSS.n2622 VSS.n2509 0.00962857
R28009 VSS.n2623 VSS.n2622 0.00962857
R28010 VSS.n2624 VSS.n2623 0.00962857
R28011 VSS.n2624 VSS.n2505 0.00962857
R28012 VSS.n2630 VSS.n2505 0.00962857
R28013 VSS.n2631 VSS.n2630 0.00962857
R28014 VSS.n2632 VSS.n2631 0.00962857
R28015 VSS.n2632 VSS.n2501 0.00962857
R28016 VSS.n2638 VSS.n2501 0.00962857
R28017 VSS.n2639 VSS.n2638 0.00962857
R28018 VSS.n2640 VSS.n2639 0.00962857
R28019 VSS.n2640 VSS.n2497 0.00962857
R28020 VSS.n2646 VSS.n2497 0.00962857
R28021 VSS.n2647 VSS.n2646 0.00962857
R28022 VSS.n2648 VSS.n2647 0.00962857
R28023 VSS.n2648 VSS.n2493 0.00962857
R28024 VSS.n2654 VSS.n2493 0.00962857
R28025 VSS.n2655 VSS.n2654 0.00962857
R28026 VSS.n2656 VSS.n2655 0.00962857
R28027 VSS.n2656 VSS.n2489 0.00962857
R28028 VSS.n2662 VSS.n2489 0.00962857
R28029 VSS.n2663 VSS.n2662 0.00962857
R28030 VSS.n2664 VSS.n2663 0.00962857
R28031 VSS.n2664 VSS.n2485 0.00962857
R28032 VSS.n2670 VSS.n2485 0.00962857
R28033 VSS.n2671 VSS.n2670 0.00962857
R28034 VSS.n2672 VSS.n2671 0.00962857
R28035 VSS.n2672 VSS.n2481 0.00962857
R28036 VSS.n2679 VSS.n2481 0.00962857
R28037 VSS.n2680 VSS.n2679 0.00962857
R28038 VSS.n2681 VSS.n2680 0.00962857
R28039 VSS.n2681 VSS.n2463 0.00962857
R28040 VSS.n2691 VSS.n2688 0.00962857
R28041 VSS.n2691 VSS.n2690 0.00962857
R28042 VSS.n2690 VSS.n2689 0.00962857
R28043 VSS.n3441 VSS.n3438 0.00962857
R28044 VSS.n3442 VSS.n3441 0.00962857
R28045 VSS.n3443 VSS.n3442 0.00962857
R28046 VSS.n3443 VSS.n3434 0.00962857
R28047 VSS.n3449 VSS.n3434 0.00962857
R28048 VSS.n3450 VSS.n3449 0.00962857
R28049 VSS.n3451 VSS.n3450 0.00962857
R28050 VSS.n3451 VSS.n3430 0.00962857
R28051 VSS.n3457 VSS.n3430 0.00962857
R28052 VSS.n3458 VSS.n3457 0.00962857
R28053 VSS.n3459 VSS.n3458 0.00962857
R28054 VSS.n3459 VSS.n3426 0.00962857
R28055 VSS.n3465 VSS.n3426 0.00962857
R28056 VSS.n3466 VSS.n3465 0.00962857
R28057 VSS.n3467 VSS.n3466 0.00962857
R28058 VSS.n3501 VSS.n3421 0.00962857
R28059 VSS.n3495 VSS.n3421 0.00962857
R28060 VSS.n3495 VSS.n3494 0.00962857
R28061 VSS.n3494 VSS.n3493 0.00962857
R28062 VSS.n3493 VSS.n3473 0.00962857
R28063 VSS.n3487 VSS.n3473 0.00962857
R28064 VSS.n3888 VSS.n2767 0.00962857
R28065 VSS.n3894 VSS.n2767 0.00962857
R28066 VSS.n3895 VSS.n3894 0.00962857
R28067 VSS.n3896 VSS.n3895 0.00962857
R28068 VSS.n3896 VSS.n2763 0.00962857
R28069 VSS.n3902 VSS.n2763 0.00962857
R28070 VSS.n3903 VSS.n3902 0.00962857
R28071 VSS.n3904 VSS.n3903 0.00962857
R28072 VSS.n3904 VSS.n2759 0.00962857
R28073 VSS.n3910 VSS.n2759 0.00962857
R28074 VSS.n3911 VSS.n3910 0.00962857
R28075 VSS.n3912 VSS.n3911 0.00962857
R28076 VSS.n3912 VSS.n2755 0.00962857
R28077 VSS.n3918 VSS.n2755 0.00962857
R28078 VSS.n3919 VSS.n3918 0.00962857
R28079 VSS.n3920 VSS.n3919 0.00962857
R28080 VSS.n3920 VSS.n2751 0.00962857
R28081 VSS.n3926 VSS.n2751 0.00962857
R28082 VSS.n3927 VSS.n3926 0.00962857
R28083 VSS.n3928 VSS.n3927 0.00962857
R28084 VSS.n3928 VSS.n2747 0.00962857
R28085 VSS.n3934 VSS.n2747 0.00962857
R28086 VSS.n3935 VSS.n3934 0.00962857
R28087 VSS.n3936 VSS.n3935 0.00962857
R28088 VSS.n3936 VSS.n2743 0.00962857
R28089 VSS.n3942 VSS.n2743 0.00962857
R28090 VSS.n3943 VSS.n3942 0.00962857
R28091 VSS.n3944 VSS.n3943 0.00962857
R28092 VSS.n3944 VSS.n2739 0.00962857
R28093 VSS.n3950 VSS.n2739 0.00962857
R28094 VSS.n3953 VSS.n3952 0.00962857
R28095 VSS.n3953 VSS.n2735 0.00962857
R28096 VSS.n3959 VSS.n2735 0.00962857
R28097 VSS.n3960 VSS.n3959 0.00962857
R28098 VSS.n3961 VSS.n3960 0.00962857
R28099 VSS.n3961 VSS.n2731 0.00962857
R28100 VSS.n3967 VSS.n2731 0.00962857
R28101 VSS.n3968 VSS.n3967 0.00962857
R28102 VSS.n3969 VSS.n3968 0.00962857
R28103 VSS.n3969 VSS.n2727 0.00962857
R28104 VSS.n3975 VSS.n2727 0.00962857
R28105 VSS.n3976 VSS.n3975 0.00962857
R28106 VSS.n3977 VSS.n3976 0.00962857
R28107 VSS.n3977 VSS.n2723 0.00962857
R28108 VSS.n3983 VSS.n2723 0.00962857
R28109 VSS.n3984 VSS.n3983 0.00962857
R28110 VSS.n3985 VSS.n3984 0.00962857
R28111 VSS.n3985 VSS.n2719 0.00962857
R28112 VSS.n3991 VSS.n2719 0.00962857
R28113 VSS.n3992 VSS.n3991 0.00962857
R28114 VSS.n3993 VSS.n3992 0.00962857
R28115 VSS.n3993 VSS.n2715 0.00962857
R28116 VSS.n3999 VSS.n2715 0.00962857
R28117 VSS.n4000 VSS.n3999 0.00962857
R28118 VSS.n4001 VSS.n4000 0.00962857
R28119 VSS.n4001 VSS.n2711 0.00962857
R28120 VSS.n4007 VSS.n2711 0.00962857
R28121 VSS.n4008 VSS.n4007 0.00962857
R28122 VSS.n4009 VSS.n4008 0.00962857
R28123 VSS.n4009 VSS.n2707 0.00962857
R28124 VSS.n4015 VSS.n2707 0.00962857
R28125 VSS.n4016 VSS.n4015 0.00962857
R28126 VSS.n4018 VSS.n4016 0.00962857
R28127 VSS.n4018 VSS.n4017 0.00962857
R28128 VSS.n4017 VSS.n2703 0.00962857
R28129 VSS.n5704 VSS.n6 0.00962857
R28130 VSS.n5704 VSS.n5703 0.00962857
R28131 VSS.n5703 VSS.n5702 0.00962857
R28132 VSS.n3440 VSS.n3437 0.00962857
R28133 VSS.n3444 VSS.n3437 0.00962857
R28134 VSS.n3444 VSS.n3435 0.00962857
R28135 VSS.n3448 VSS.n3435 0.00962857
R28136 VSS.n3448 VSS.n3433 0.00962857
R28137 VSS.n3452 VSS.n3433 0.00962857
R28138 VSS.n3452 VSS.n3431 0.00962857
R28139 VSS.n3456 VSS.n3431 0.00962857
R28140 VSS.n3456 VSS.n3429 0.00962857
R28141 VSS.n3460 VSS.n3429 0.00962857
R28142 VSS.n3460 VSS.n3427 0.00962857
R28143 VSS.n3464 VSS.n3427 0.00962857
R28144 VSS.n3464 VSS.n3425 0.00962857
R28145 VSS.n3468 VSS.n3425 0.00962857
R28146 VSS.n3468 VSS.n3422 0.00962857
R28147 VSS.n3500 VSS.n3422 0.00962857
R28148 VSS.n3500 VSS.n3423 0.00962857
R28149 VSS.n3496 VSS.n3423 0.00962857
R28150 VSS.n3496 VSS.n3472 0.00962857
R28151 VSS.n3492 VSS.n3472 0.00962857
R28152 VSS.n3492 VSS.n3474 0.00962857
R28153 VSS.n3488 VSS.n3474 0.00962857
R28154 VSS.n3488 VSS.n3476 0.00962857
R28155 VSS.n3482 VSS.n3476 0.00962857
R28156 VSS.n3482 VSS.n2776 0.00962857
R28157 VSS.n3879 VSS.n2776 0.00962857
R28158 VSS.n3879 VSS.n2774 0.00962857
R28159 VSS.n3883 VSS.n2774 0.00962857
R28160 VSS.n3883 VSS.n2770 0.00962857
R28161 VSS.n3889 VSS.n2770 0.00962857
R28162 VSS.n3889 VSS.n2768 0.00962857
R28163 VSS.n3893 VSS.n2768 0.00962857
R28164 VSS.n3893 VSS.n2766 0.00962857
R28165 VSS.n3897 VSS.n2766 0.00962857
R28166 VSS.n3897 VSS.n2764 0.00962857
R28167 VSS.n3901 VSS.n2764 0.00962857
R28168 VSS.n3901 VSS.n2762 0.00962857
R28169 VSS.n3905 VSS.n2762 0.00962857
R28170 VSS.n3905 VSS.n2760 0.00962857
R28171 VSS.n3909 VSS.n2760 0.00962857
R28172 VSS.n3909 VSS.n2758 0.00962857
R28173 VSS.n3913 VSS.n2758 0.00962857
R28174 VSS.n3913 VSS.n2756 0.00962857
R28175 VSS.n3917 VSS.n2756 0.00962857
R28176 VSS.n3917 VSS.n2754 0.00962857
R28177 VSS.n3921 VSS.n2754 0.00962857
R28178 VSS.n3921 VSS.n2752 0.00962857
R28179 VSS.n3925 VSS.n2752 0.00962857
R28180 VSS.n3925 VSS.n2750 0.00962857
R28181 VSS.n3929 VSS.n2750 0.00962857
R28182 VSS.n3929 VSS.n2748 0.00962857
R28183 VSS.n3933 VSS.n2748 0.00962857
R28184 VSS.n3933 VSS.n2746 0.00962857
R28185 VSS.n3937 VSS.n2746 0.00962857
R28186 VSS.n3937 VSS.n2744 0.00962857
R28187 VSS.n3941 VSS.n2744 0.00962857
R28188 VSS.n3941 VSS.n2742 0.00962857
R28189 VSS.n3945 VSS.n2742 0.00962857
R28190 VSS.n3945 VSS.n2740 0.00962857
R28191 VSS.n3949 VSS.n2740 0.00962857
R28192 VSS.n3949 VSS.n2738 0.00962857
R28193 VSS.n3954 VSS.n2738 0.00962857
R28194 VSS.n3954 VSS.n2736 0.00962857
R28195 VSS.n3958 VSS.n2736 0.00962857
R28196 VSS.n3958 VSS.n2734 0.00962857
R28197 VSS.n3962 VSS.n2734 0.00962857
R28198 VSS.n3962 VSS.n2732 0.00962857
R28199 VSS.n3966 VSS.n2732 0.00962857
R28200 VSS.n3966 VSS.n2730 0.00962857
R28201 VSS.n3970 VSS.n2730 0.00962857
R28202 VSS.n3970 VSS.n2728 0.00962857
R28203 VSS.n3974 VSS.n2728 0.00962857
R28204 VSS.n3974 VSS.n2726 0.00962857
R28205 VSS.n3978 VSS.n2726 0.00962857
R28206 VSS.n3978 VSS.n2724 0.00962857
R28207 VSS.n3982 VSS.n2724 0.00962857
R28208 VSS.n3982 VSS.n2722 0.00962857
R28209 VSS.n3986 VSS.n2722 0.00962857
R28210 VSS.n3986 VSS.n2720 0.00962857
R28211 VSS.n3990 VSS.n2720 0.00962857
R28212 VSS.n3990 VSS.n2718 0.00962857
R28213 VSS.n3994 VSS.n2718 0.00962857
R28214 VSS.n3994 VSS.n2716 0.00962857
R28215 VSS.n3998 VSS.n2716 0.00962857
R28216 VSS.n3998 VSS.n2714 0.00962857
R28217 VSS.n4002 VSS.n2714 0.00962857
R28218 VSS.n4002 VSS.n2712 0.00962857
R28219 VSS.n4006 VSS.n2712 0.00962857
R28220 VSS.n4006 VSS.n2710 0.00962857
R28221 VSS.n4010 VSS.n2710 0.00962857
R28222 VSS.n4010 VSS.n2708 0.00962857
R28223 VSS.n4014 VSS.n2708 0.00962857
R28224 VSS.n4014 VSS.n2706 0.00962857
R28225 VSS.n4019 VSS.n2706 0.00962857
R28226 VSS.n4019 VSS.n2704 0.00962857
R28227 VSS.n4023 VSS.n2704 0.00962857
R28228 VSS.n4024 VSS.n4023 0.00962857
R28229 VSS.n5709 VSS.n2 0.00962857
R28230 VSS.n5705 VSS.n2 0.00962857
R28231 VSS.n5705 VSS.n5 0.00962857
R28232 VSS.n4880 DVSS 0.00958867
R28233 VSS.n4871 DVSS 0.00958867
R28234 VSS.n3139 VSS.n3135 0.00958257
R28235 VSS.n3354 VSS.n2914 0.00958257
R28236 VSS.n5190 VSS.n5170 0.00956429
R28237 VSS.n911 VSS.n218 0.0095301
R28238 VSS.n3363 VSS.n2904 0.0095
R28239 VSS.n2987 VSS.n2986 0.0095
R28240 VSS.n2993 VSS.n2992 0.0095
R28241 VSS.n2985 VSS.n2983 0.0095
R28242 VSS.n2996 VSS.n2995 0.0095
R28243 VSS.n3351 VSS.n3349 0.0095
R28244 VSS.n2930 VSS.n2924 0.0095
R28245 VSS.n3343 VSS.n2931 0.0095
R28246 VSS.n3342 VSS.n2932 0.0095
R28247 VSS.n3333 VSS.n3331 0.0095
R28248 VSS.n3121 VSS.n3113 0.0095
R28249 VSS.n3120 VSS.n3100 0.0095
R28250 VSS.n3129 VSS.n3128 0.0095
R28251 VSS.n3103 VSS.n3101 0.0095
R28252 VSS.n3296 VSS.n3089 0.0095
R28253 VSS.n3295 VSS.n3090 0.0095
R28254 VSS.n3146 VSS.n3145 0.0095
R28255 VSS.n3287 VSS.n3286 0.0095
R28256 VSS.n3276 VSS.n3147 0.0095
R28257 VSS.n5097 VSS.n4320 0.0095
R28258 VSS.n5088 VSS.n4336 0.0095
R28259 VSS.n4906 VSS.n4587 0.0095
R28260 VSS.n4897 VSS.n4603 0.0095
R28261 VSS.n4662 VSS.n4661 0.0095
R28262 VSS.n4672 VSS.n4670 0.0095
R28263 VSS.n4854 VSS.n4853 0.0095
R28264 VSS.n4864 VSS.n4862 0.0095
R28265 VSS.n5681 VSS.n5680 0.00934354
R28266 VSS.n5680 VSS.n5679 0.00934354
R28267 VSS.n2076 VSS.n2075 0.00933782
R28268 VSS.n2069 VSS.n1594 0.00933782
R28269 VSS.n2075 VSS.n1594 0.00933782
R28270 VSS.n2073 VSS.n2069 0.00933782
R28271 VSS.n1809 VSS.n16 0.00933782
R28272 VSS.n1811 VSS.n1809 0.00933782
R28273 VSS.n1880 VSS.n1879 0.00928049
R28274 VSS.n1875 VSS.n1874 0.00928049
R28275 VSS.n1914 VSS.n1727 0.00928049
R28276 VSS.n1900 VSS.n1747 0.00928049
R28277 VSS.n1952 VSS.n1703 0.00928049
R28278 VSS.n1938 VSS.n1705 0.00928049
R28279 VSS.n1738 VSS.n1736 0.00928049
R28280 VSS.n1977 VSS.n1685 0.00928049
R28281 VSS.n1732 VSS.n1730 0.00928049
R28282 VSS.n2009 VSS.n1660 0.00928049
R28283 VSS.n2045 VSS.n2044 0.00928049
R28284 VSS.n2040 VSS.n2039 0.00928049
R28285 VSS.n1396 VSS.n33 0.00924286
R28286 VSS.n5438 VSS.n5437 0.00910927
R28287 VSS.n5700 VSS.n5699 0.00910927
R28288 VSS.n636 VSS.n635 0.00909873
R28289 VSS.n5109 VSS.n5108 0.009
R28290 VSS.n5077 VSS.n5076 0.009
R28291 VSS.n4919 VSS.n4918 0.009
R28292 VSS.n4886 VSS.n4885 0.009
R28293 VSS.n4651 VSS.n4305 0.009
R28294 VSS.n4643 VSS.n4350 0.009
R28295 VSS.n4843 VSS.n4575 0.009
R28296 VSS.n4623 VSS.n4619 0.009
R28297 VSS.n3040 VSS.n2830 0.00894122
R28298 VSS.n3040 VSS.n2836 0.00894122
R28299 VSS.n4118 VSS.n4116 0.00892143
R28300 VSS.n4130 VSS.n4129 0.00892143
R28301 VSS.n3467 VSS.n3419 0.00892143
R28302 VSS.n3502 VSS.n3420 0.00892143
R28303 VSS.n217 VSS.n172 0.00882776
R28304 VSS.n3641 VSS.n3640 0.00879286
R28305 VSS.n2885 VSS.n2880 0.00879286
R28306 VSS.n3638 VSS.n3549 0.00879286
R28307 VSS.n4201 VSS.n2398 0.00879286
R28308 VSS.n3370 VSS.n2899 0.0086
R28309 VSS.n3716 VSS.n2827 0.00853571
R28310 VSS.n3715 VSS.n2833 0.00853571
R28311 VSS.n3713 VSS.n3712 0.00853571
R28312 VSS.n1920 VSS.n1724 0.00853571
R28313 VSS.n1919 VSS.n1725 0.00853571
R28314 VSS.n1749 VSS.n1748 0.00853571
R28315 VSS.n1912 VSS.n1911 0.00853571
R28316 VSS.n1756 VSS.n1750 0.00853571
R28317 VSS.n1905 VSS.n1757 0.00853571
R28318 VSS.n1904 VSS.n1897 0.00853571
R28319 VSS.n4148 VSS.n4147 0.00853571
R28320 VSS.n5159 DVSS 0.00852817
R28321 VSS.n5158 DVSS 0.00852817
R28322 VSS.n5056 VSS.n4375 0.0085
R28323 VSS.n4550 VSS.n4538 0.0085
R28324 VSS.n4706 VSS.n4377 0.0085
R28325 VSS.n4824 VSS.n4823 0.0085
R28326 VSS.n1828 VSS.n20 0.00847143
R28327 VSS.n3016 VSS.n2903 0.00847143
R28328 VSS.n3487 VSS.n3486 0.00847143
R28329 VSS.n3484 VSS.n3477 0.00847143
R28330 VSS.n3483 VSS.n3480 0.00847143
R28331 VSS.n3479 VSS.n2777 0.00847143
R28332 VSS.n3878 VSS.n3877 0.00847143
R28333 VSS.n2778 VSS.n2773 0.00847143
R28334 VSS.n3885 VSS.n3884 0.00847143
R28335 VSS.n3887 VSS.n2771 0.00847143
R28336 VSS.n537 VSS.n365 0.00842994
R28337 VSS.n3280 VSS.n3153 0.00834286
R28338 VSS.n3246 VSS.n3245 0.00834286
R28339 VSS.n4222 VSS.n4221 0.00827857
R28340 VSS.n2397 VSS.n2393 0.00827857
R28341 VSS.n5022 DVSS 0.00825862
R28342 DVSS VSS.n4740 0.00825862
R28343 VSS.n3414 VSS.n3413 0.00823128
R28344 VSS.n3052 VSS.n2834 0.00822787
R28345 VSS.n3032 VSS.n2828 0.00822787
R28346 VSS.n3411 VSS.n3410 0.00821429
R28347 VSS.n5236 VSS.n2244 0.00815
R28348 VSS.n5071 VSS.n4357 0.00803695
R28349 VSS.n4681 VSS.n4641 0.00803695
R28350 VSS.n5115 VSS.n4296 0.00803521
R28351 VSS.n4649 VSS.n4297 0.00803521
R28352 VSS.n5107 VSS.n4304 0.00803521
R28353 VSS.n5106 VSS.n4306 0.00803521
R28354 VSS.n5103 VSS.n5102 0.00803521
R28355 VSS.n4660 VSS.n4317 0.00803521
R28356 VSS.n5095 VSS.n4324 0.00803521
R28357 VSS.n5094 VSS.n4326 0.00803521
R28358 VSS.n5091 VSS.n5090 0.00803521
R28359 VSS.n4671 VSS.n4334 0.00803521
R28360 VSS.n5083 VSS.n4341 0.00803521
R28361 VSS.n5082 VSS.n4343 0.00803521
R28362 VSS.n5079 VSS.n5078 0.00803521
R28363 VSS.n4685 VSS.n4351 0.00803521
R28364 VSS.n4691 VSS.n4690 0.00803521
R28365 VSS.n5067 VSS.n4361 0.00803521
R28366 VSS.n5066 VSS.n4363 0.00803521
R28367 VSS.n5063 VSS.n5062 0.00803521
R28368 VSS.n4702 VSS.n4369 0.00803521
R28369 VSS.n5055 VSS.n4376 0.00803521
R28370 VSS.n5054 VSS.n4378 0.00803521
R28371 VSS.n5051 VSS.n5050 0.00803521
R28372 VSS.n4714 VSS.n4386 0.00803521
R28373 VSS.n5043 VSS.n4395 0.00803521
R28374 VSS.n5042 VSS.n4397 0.00803521
R28375 VSS.n5039 VSS.n5038 0.00803521
R28376 VSS.n4725 VSS.n4405 0.00803521
R28377 VSS.n5031 VSS.n4412 0.00803521
R28378 VSS.n5030 VSS.n4414 0.00803521
R28379 VSS.n5027 VSS.n5026 0.00803521
R28380 VSS.n4737 VSS.n4422 0.00803521
R28381 VSS.n5019 VSS.n4430 0.00803521
R28382 VSS.n5018 VSS.n4432 0.00803521
R28383 VSS.n5015 VSS.n5014 0.00803521
R28384 VSS.n4752 VSS.n4440 0.00803521
R28385 VSS.n4758 VSS.n4757 0.00803521
R28386 VSS.n5003 VSS.n4451 0.00803521
R28387 VSS.n5002 VSS.n4453 0.00803521
R28388 VSS.n4999 VSS.n4998 0.00803521
R28389 VSS.n4769 VSS.n4459 0.00803521
R28390 VSS.n4991 VSS.n4466 0.00803521
R28391 VSS.n4990 VSS.n4468 0.00803521
R28392 VSS.n4987 VSS.n4986 0.00803521
R28393 VSS.n4781 VSS.n4476 0.00803521
R28394 VSS.n4979 VSS.n4485 0.00803521
R28395 VSS.n4978 VSS.n4487 0.00803521
R28396 VSS.n4975 VSS.n4974 0.00803521
R28397 VSS.n4793 VSS.n4495 0.00803521
R28398 VSS.n4967 VSS.n4503 0.00803521
R28399 VSS.n4966 VSS.n4505 0.00803521
R28400 VSS.n4963 VSS.n4962 0.00803521
R28401 VSS.n4805 VSS.n4513 0.00803521
R28402 VSS.n4955 VSS.n4521 0.00803521
R28403 VSS.n4954 VSS.n4523 0.00803521
R28404 VSS.n4951 VSS.n4950 0.00803521
R28405 VSS.n4816 VSS.n4531 0.00803521
R28406 VSS.n4942 VSS.n4539 0.00803521
R28407 VSS.n4941 VSS.n4541 0.00803521
R28408 VSS.n4938 VSS.n4937 0.00803521
R28409 VSS.n4829 VSS.n4549 0.00803521
R28410 VSS.n4930 VSS.n4556 0.00803521
R28411 VSS.n4929 VSS.n4558 0.00803521
R28412 VSS.n4926 VSS.n4925 0.00803521
R28413 VSS.n4841 VSS.n4566 0.00803521
R28414 VSS.n4917 VSS.n4574 0.00803521
R28415 VSS.n4916 VSS.n4576 0.00803521
R28416 VSS.n4913 VSS.n4912 0.00803521
R28417 VSS.n4852 VSS.n4584 0.00803521
R28418 VSS.n4904 VSS.n4591 0.00803521
R28419 VSS.n4903 VSS.n4593 0.00803521
R28420 VSS.n4900 VSS.n4899 0.00803521
R28421 VSS.n4863 VSS.n4601 0.00803521
R28422 VSS.n4892 VSS.n4609 0.00803521
R28423 VSS.n4891 VSS.n4611 0.00803521
R28424 VSS.n4888 VSS.n4887 0.00803521
R28425 VSS.n4878 VSS.n4620 0.00803521
R28426 VSS.n4877 VSS.n2280 0.00803521
R28427 VSS.n5134 VSS.n5133 0.00803521
R28428 VSS.n5033 VSS.n4408 0.008
R28429 VSS.n4961 VSS.n4514 0.008
R28430 VSS.n4727 VSS.n4726 0.008
R28431 VSS.n4801 VSS.n4512 0.008
R28432 VSS.n4056 VSS.n2468 0.00789286
R28433 VSS.n2688 VSS.n2462 0.00789286
R28434 VSS.n4026 VSS.n4025 0.00789286
R28435 VSS.n6 VSS.n1 0.00789286
R28436 VSS.n2684 VSS 0.00782857
R28437 VSS.n3187 DVSS 0.00782857
R28438 VSS.n3584 DVSS 0.00782857
R28439 VSS.n3583 DVSS 0.00782857
R28440 VSS.n1840 DVSS 0.00782857
R28441 DVSS VSS.n1394 0.00782857
R28442 VSS.n1393 DVSS 0.00782857
R28443 VSS.n3188 DVSS 0.00782857
R28444 VSS.n5179 DVSS 0.00782857
R28445 VSS.n5180 DVSS 0.00782857
R28446 VSS.n4024 VSS 0.00782857
R28447 VSS.n4102 VSS.n4101 0.00776429
R28448 VSS.n1878 VSS.n1773 0.00761735
R28449 VSS.n1876 VSS.n1774 0.00761735
R28450 VSS.n1916 VSS.n1915 0.00761735
R28451 VSS.n1902 VSS.n1899 0.00761735
R28452 VSS.n1954 VSS.n1953 0.00761735
R28453 VSS.n1940 VSS.n1937 0.00761735
R28454 VSS.n1739 VSS.n1676 0.00761735
R28455 VSS.n1975 VSS.n1687 0.00761735
R28456 VSS.n1733 VSS.n1649 0.00761735
R28457 VSS.n2007 VSS.n1662 0.00761735
R28458 VSS.n2043 VSS.n1629 0.00761735
R28459 VSS.n2041 VSS.n1630 0.00761735
R28460 VSS.n2022 VSS.n2021 0.00757143
R28461 VSS.n2018 VSS.n1648 0.00757143
R28462 VSS.n2017 VSS.n1651 0.00757143
R28463 VSS.n1658 VSS.n1657 0.00757143
R28464 VSS.n2011 VSS.n2010 0.00757143
R28465 VSS.n1663 VSS.n1659 0.00757143
R28466 VSS.n2005 VSS.n1664 0.00757143
R28467 VSS.n3068 VSS.n3061 0.00757143
R28468 VSS.n3065 VSS.n2948 0.00757143
R28469 VSS.n1989 VSS.n1675 0.00750714
R28470 VSS.n1986 VSS.n1985 0.00750714
R28471 VSS.n1682 VSS.n1678 0.00750714
R28472 VSS.n1979 VSS.n1683 0.00750714
R28473 VSS.n1978 VSS.n1684 0.00750714
R28474 VSS.n1689 VSS.n1688 0.00750714
R28475 VSS.n1973 VSS.n1972 0.00750714
R28476 VSS.n1792 VSS.n1788 0.00750714
R28477 VSS.n1858 VSS.n1857 0.00750714
R28478 VSS.n1854 VSS.n1798 0.00750714
R28479 VSS.n2959 VSS.n2958 0.00750714
R28480 VSS.n3112 VSS.n3111 0.00750714
R28481 VSS.n5013 VSS.n5012 0.0075
R28482 VSS.n4984 VSS.n4478 0.0075
R28483 VSS.n4636 VSS.n4439 0.0075
R28484 VSS.n4782 VSS.n4780 0.0075
R28485 VSS.n1152 VSS.n25 0.00745122
R28486 VSS.n1162 VSS.n28 0.00745122
R28487 VSS.n3278 VSS.n3275 0.00739189
R28488 VSS.n3273 VSS.n3154 0.00739189
R28489 VSS.n1879 VSS.n1770 0.00730488
R28490 VSS.n1875 VSS.n1770 0.00730488
R28491 VSS.n1914 VSS.n1913 0.00730488
R28492 VSS.n1913 VSS.n1747 0.00730488
R28493 VSS.n1952 VSS.n1951 0.00730488
R28494 VSS.n1951 VSS.n1705 0.00730488
R28495 VSS.n1738 VSS.n1737 0.00730488
R28496 VSS.n1737 VSS.n1685 0.00730488
R28497 VSS.n1732 VSS.n1731 0.00730488
R28498 VSS.n1731 VSS.n1660 0.00730488
R28499 VSS.n2044 VSS.n1626 0.00730488
R28500 VSS.n2040 VSS.n1626 0.00730488
R28501 VSS.n4312 VSS.n4311 0.00716667
R28502 VSS.n4313 VSS.n4312 0.00716667
R28503 VSS.n4314 VSS.n4313 0.00716667
R28504 VSS.n4328 VSS.n4314 0.00716667
R28505 VSS.n4329 VSS.n4328 0.00716667
R28506 VSS.n4330 VSS.n4329 0.00716667
R28507 VSS.n4331 VSS.n4330 0.00716667
R28508 VSS.n4345 VSS.n4331 0.00716667
R28509 VSS.n4346 VSS.n4345 0.00716667
R28510 VSS.n4347 VSS.n4346 0.00716667
R28511 VSS.n4348 VSS.n4347 0.00716667
R28512 VSS.n4686 VSS.n4348 0.00716667
R28513 VSS.n4688 VSS.n4686 0.00716667
R28514 VSS.n4688 VSS.n4687 0.00716667
R28515 VSS.n4687 VSS.n4365 0.00716667
R28516 VSS.n4366 VSS.n4365 0.00716667
R28517 VSS.n4380 VSS.n4366 0.00716667
R28518 VSS.n4381 VSS.n4380 0.00716667
R28519 VSS.n4382 VSS.n4381 0.00716667
R28520 VSS.n4383 VSS.n4382 0.00716667
R28521 VSS.n4399 VSS.n4383 0.00716667
R28522 VSS.n4400 VSS.n4399 0.00716667
R28523 VSS.n4401 VSS.n4400 0.00716667
R28524 VSS.n4402 VSS.n4401 0.00716667
R28525 VSS.n4416 VSS.n4402 0.00716667
R28526 VSS.n4417 VSS.n4416 0.00716667
R28527 VSS.n4418 VSS.n4417 0.00716667
R28528 VSS.n4419 VSS.n4418 0.00716667
R28529 VSS.n4434 VSS.n4419 0.00716667
R28530 VSS.n4435 VSS.n4434 0.00716667
R28531 VSS.n4436 VSS.n4435 0.00716667
R28532 VSS.n4437 VSS.n4436 0.00716667
R28533 VSS.n4753 VSS.n4437 0.00716667
R28534 VSS.n4755 VSS.n4753 0.00716667
R28535 VSS.n4755 VSS.n4754 0.00716667
R28536 VSS.n4754 VSS.n4455 0.00716667
R28537 VSS.n4456 VSS.n4455 0.00716667
R28538 VSS.n4470 VSS.n4456 0.00716667
R28539 VSS.n4471 VSS.n4470 0.00716667
R28540 VSS.n4472 VSS.n4471 0.00716667
R28541 VSS.n4473 VSS.n4472 0.00716667
R28542 VSS.n4489 VSS.n4473 0.00716667
R28543 VSS.n4490 VSS.n4489 0.00716667
R28544 VSS.n4491 VSS.n4490 0.00716667
R28545 VSS.n4492 VSS.n4491 0.00716667
R28546 VSS.n4507 VSS.n4492 0.00716667
R28547 VSS.n4508 VSS.n4507 0.00716667
R28548 VSS.n4509 VSS.n4508 0.00716667
R28549 VSS.n4510 VSS.n4509 0.00716667
R28550 VSS.n4525 VSS.n4510 0.00716667
R28551 VSS.n4526 VSS.n4525 0.00716667
R28552 VSS.n4527 VSS.n4526 0.00716667
R28553 VSS.n4528 VSS.n4527 0.00716667
R28554 VSS.n4543 VSS.n4528 0.00716667
R28555 VSS.n4544 VSS.n4543 0.00716667
R28556 VSS.n4545 VSS.n4544 0.00716667
R28557 VSS.n4546 VSS.n4545 0.00716667
R28558 VSS.n4560 VSS.n4546 0.00716667
R28559 VSS.n4561 VSS.n4560 0.00716667
R28560 VSS.n4562 VSS.n4561 0.00716667
R28561 VSS.n4563 VSS.n4562 0.00716667
R28562 VSS.n4578 VSS.n4563 0.00716667
R28563 VSS.n4579 VSS.n4578 0.00716667
R28564 VSS.n4580 VSS.n4579 0.00716667
R28565 VSS.n4581 VSS.n4580 0.00716667
R28566 VSS.n4595 VSS.n4581 0.00716667
R28567 VSS.n4596 VSS.n4595 0.00716667
R28568 VSS.n4597 VSS.n4596 0.00716667
R28569 VSS.n4598 VSS.n4597 0.00716667
R28570 VSS.n4613 VSS.n4598 0.00716667
R28571 VSS.n4614 VSS.n4613 0.00716667
R28572 VSS.n4615 VSS.n4614 0.00716667
R28573 VSS.n4616 VSS.n4615 0.00716667
R28574 VSS.n4617 VSS.n4616 0.00716667
R28575 VSS.n4617 VSS.n2278 0.00716667
R28576 VSS.n5136 VSS.n2278 0.00716667
R28577 VSS.n5137 VSS.n5136 0.00716667
R28578 VSS.n5138 VSS.n5137 0.00716667
R28579 VSS.n5138 VSS.n2274 0.00716667
R28580 VSS.n5144 VSS.n2274 0.00716667
R28581 VSS.n5145 VSS.n5144 0.00716667
R28582 VSS.n5146 VSS.n5145 0.00716667
R28583 VSS.n5147 VSS.n5146 0.00716667
R28584 VSS.n5148 VSS.n5147 0.00716667
R28585 VSS.n5151 VSS.n5148 0.00716667
R28586 VSS.n5152 VSS.n5151 0.00716667
R28587 VSS.n5153 VSS.n5152 0.00716667
R28588 VSS.n5154 VSS.n5153 0.00716667
R28589 VSS.n5690 VSS.n23 0.00712143
R28590 VSS.n1838 VSS.n19 0.00712143
R28591 VSS.n1298 VSS.n1297 0.00712143
R28592 VSS.n1587 VSS.n1586 0.00712143
R28593 VSS.n4239 VSS.n4238 0.00712143
R28594 VSS.n4193 VSS.n2403 0.00705714
R28595 VSS.n2408 VSS.n2407 0.00705714
R28596 VSS.n4187 VSS.n4186 0.00705714
R28597 VSS.n1004 VSS.n105 0.00700873
R28598 VSS.n5005 VSS.n5004 0.007
R28599 VSS.n4992 VSS.n4465 0.007
R28600 VSS.n4760 VSS.n4452 0.007
R28601 VSS.n4773 VSS.n4467 0.007
R28602 VSS.n4232 VSS.n4231 0.00699286
R28603 VSS.n4219 VSS.n2388 0.00699286
R28604 VSS.n4251 VSS.n4250 0.00692857
R28605 VSS.n3323 VSS.n3322 0.006875
R28606 VSS.n3320 VSS.n2957 0.006875
R28607 VSS.n3332 VSS.n2945 0.006875
R28608 VSS.n3335 VSS.n3334 0.006875
R28609 VSS.n4053 VSS.n4043 0.0068
R28610 VSS.n1700 VSS.n1696 0.0068
R28611 VSS.n1958 VSS.n1957 0.0068
R28612 VSS.n1706 VSS.n1701 0.0068
R28613 VSS.n1950 VSS.n1707 0.0068
R28614 VSS.n1949 VSS.n1708 0.0068
R28615 VSS.n1715 VSS.n1714 0.0068
R28616 VSS.n1943 VSS.n1942 0.0068
R28617 VSS.n3951 VSS.n3950 0.0068
R28618 VSS.n1154 VSS.n25 0.00671951
R28619 VSS.n1160 VSS.n28 0.00671951
R28620 VSS.n3445 VSS.n3436 0.00658571
R28621 VSS.n3446 VSS.n3445 0.00658571
R28622 VSS.n3447 VSS.n3446 0.00658571
R28623 VSS.n3447 VSS.n3432 0.00658571
R28624 VSS.n3453 VSS.n3432 0.00658571
R28625 VSS.n3454 VSS.n3453 0.00658571
R28626 VSS.n3455 VSS.n3454 0.00658571
R28627 VSS.n3455 VSS.n3428 0.00658571
R28628 VSS.n3461 VSS.n3428 0.00658571
R28629 VSS.n3462 VSS.n3461 0.00658571
R28630 VSS.n3463 VSS.n3462 0.00658571
R28631 VSS.n3463 VSS.n3424 0.00658571
R28632 VSS.n3469 VSS.n3424 0.00658571
R28633 VSS.n3470 VSS.n3469 0.00658571
R28634 VSS.n3499 VSS.n3470 0.00658571
R28635 VSS.n3499 VSS.n3498 0.00658571
R28636 VSS.n3498 VSS.n3497 0.00658571
R28637 VSS.n3497 VSS.n3471 0.00658571
R28638 VSS.n3491 VSS.n3471 0.00658571
R28639 VSS.n3491 VSS.n3490 0.00658571
R28640 VSS.n3490 VSS.n3489 0.00658571
R28641 VSS.n3489 VSS.n3475 0.00658571
R28642 VSS.n3481 VSS.n3475 0.00658571
R28643 VSS.n3481 VSS.n2775 0.00658571
R28644 VSS.n3880 VSS.n2775 0.00658571
R28645 VSS.n3881 VSS.n3880 0.00658571
R28646 VSS.n3882 VSS.n3881 0.00658571
R28647 VSS.n3882 VSS.n2769 0.00658571
R28648 VSS.n3890 VSS.n2769 0.00658571
R28649 VSS.n3891 VSS.n3890 0.00658571
R28650 VSS.n3892 VSS.n3891 0.00658571
R28651 VSS.n3892 VSS.n2765 0.00658571
R28652 VSS.n3898 VSS.n2765 0.00658571
R28653 VSS.n3899 VSS.n3898 0.00658571
R28654 VSS.n3900 VSS.n3899 0.00658571
R28655 VSS.n3900 VSS.n2761 0.00658571
R28656 VSS.n3906 VSS.n2761 0.00658571
R28657 VSS.n3907 VSS.n3906 0.00658571
R28658 VSS.n3908 VSS.n3907 0.00658571
R28659 VSS.n3908 VSS.n2757 0.00658571
R28660 VSS.n3914 VSS.n2757 0.00658571
R28661 VSS.n3915 VSS.n3914 0.00658571
R28662 VSS.n3916 VSS.n3915 0.00658571
R28663 VSS.n3916 VSS.n2753 0.00658571
R28664 VSS.n3922 VSS.n2753 0.00658571
R28665 VSS.n3923 VSS.n3922 0.00658571
R28666 VSS.n3924 VSS.n3923 0.00658571
R28667 VSS.n3924 VSS.n2749 0.00658571
R28668 VSS.n3930 VSS.n2749 0.00658571
R28669 VSS.n3931 VSS.n3930 0.00658571
R28670 VSS.n3932 VSS.n3931 0.00658571
R28671 VSS.n3932 VSS.n2745 0.00658571
R28672 VSS.n3938 VSS.n2745 0.00658571
R28673 VSS.n3939 VSS.n3938 0.00658571
R28674 VSS.n3940 VSS.n3939 0.00658571
R28675 VSS.n3940 VSS.n2741 0.00658571
R28676 VSS.n3946 VSS.n2741 0.00658571
R28677 VSS.n3947 VSS.n3946 0.00658571
R28678 VSS.n3948 VSS.n3947 0.00658571
R28679 VSS.n3948 VSS.n2737 0.00658571
R28680 VSS.n3955 VSS.n2737 0.00658571
R28681 VSS.n3956 VSS.n3955 0.00658571
R28682 VSS.n3957 VSS.n3956 0.00658571
R28683 VSS.n3957 VSS.n2733 0.00658571
R28684 VSS.n3963 VSS.n2733 0.00658571
R28685 VSS.n3964 VSS.n3963 0.00658571
R28686 VSS.n3965 VSS.n3964 0.00658571
R28687 VSS.n3965 VSS.n2729 0.00658571
R28688 VSS.n3971 VSS.n2729 0.00658571
R28689 VSS.n3972 VSS.n3971 0.00658571
R28690 VSS.n3973 VSS.n3972 0.00658571
R28691 VSS.n3973 VSS.n2725 0.00658571
R28692 VSS.n3979 VSS.n2725 0.00658571
R28693 VSS.n3980 VSS.n3979 0.00658571
R28694 VSS.n3981 VSS.n3980 0.00658571
R28695 VSS.n3981 VSS.n2721 0.00658571
R28696 VSS.n3987 VSS.n2721 0.00658571
R28697 VSS.n3988 VSS.n3987 0.00658571
R28698 VSS.n3989 VSS.n3988 0.00658571
R28699 VSS.n3989 VSS.n2717 0.00658571
R28700 VSS.n3995 VSS.n2717 0.00658571
R28701 VSS.n3996 VSS.n3995 0.00658571
R28702 VSS.n3997 VSS.n3996 0.00658571
R28703 VSS.n3997 VSS.n2713 0.00658571
R28704 VSS.n4003 VSS.n2713 0.00658571
R28705 VSS.n4004 VSS.n4003 0.00658571
R28706 VSS.n4005 VSS.n4004 0.00658571
R28707 VSS.n4005 VSS.n2709 0.00658571
R28708 VSS.n4011 VSS.n2709 0.00658571
R28709 VSS.n4012 VSS.n4011 0.00658571
R28710 VSS.n4013 VSS.n4012 0.00658571
R28711 VSS.n4013 VSS.n2705 0.00658571
R28712 VSS.n4020 VSS.n2705 0.00658571
R28713 VSS.n4021 VSS.n4020 0.00658571
R28714 VSS.n4022 VSS.n4021 0.00658571
R28715 VSS.n4022 VSS.n3 0.00658571
R28716 VSS.n5708 VSS.n3 0.00658571
R28717 VSS.n5707 VSS.n5706 0.00658571
R28718 VSS.n2320 VSS.n2309 0.00658571
R28719 VSS.n2321 VSS.n2320 0.00658571
R28720 VSS.n2322 VSS.n2321 0.00658571
R28721 VSS.n2322 VSS.n2305 0.00658571
R28722 VSS.n2328 VSS.n2305 0.00658571
R28723 VSS.n2329 VSS.n2328 0.00658571
R28724 VSS.n2330 VSS.n2329 0.00658571
R28725 VSS.n2330 VSS.n2301 0.00658571
R28726 VSS.n2336 VSS.n2301 0.00658571
R28727 VSS.n2337 VSS.n2336 0.00658571
R28728 VSS.n4279 VSS.n2337 0.00658571
R28729 VSS.n4279 VSS.n4278 0.00658571
R28730 VSS.n4278 VSS.n4277 0.00658571
R28731 VSS.n4277 VSS.n2338 0.00658571
R28732 VSS.n4271 VSS.n2338 0.00658571
R28733 VSS.n4271 VSS.n4270 0.00658571
R28734 VSS.n4270 VSS.n4269 0.00658571
R28735 VSS.n4269 VSS.n2342 0.00658571
R28736 VSS.n4263 VSS.n2342 0.00658571
R28737 VSS.n4263 VSS.n4262 0.00658571
R28738 VSS.n4262 VSS.n4261 0.00658571
R28739 VSS.n4261 VSS.n2346 0.00658571
R28740 VSS.n4255 VSS.n2346 0.00658571
R28741 VSS.n4255 VSS.n4254 0.00658571
R28742 VSS.n4254 VSS.n4253 0.00658571
R28743 VSS.n4253 VSS.n2350 0.00658571
R28744 VSS.n2547 VSS.n2350 0.00658571
R28745 VSS.n2548 VSS.n2547 0.00658571
R28746 VSS.n2548 VSS.n2543 0.00658571
R28747 VSS.n2554 VSS.n2543 0.00658571
R28748 VSS.n2555 VSS.n2554 0.00658571
R28749 VSS.n2556 VSS.n2555 0.00658571
R28750 VSS.n2556 VSS.n2539 0.00658571
R28751 VSS.n2562 VSS.n2539 0.00658571
R28752 VSS.n2563 VSS.n2562 0.00658571
R28753 VSS.n2564 VSS.n2563 0.00658571
R28754 VSS.n2564 VSS.n2535 0.00658571
R28755 VSS.n2570 VSS.n2535 0.00658571
R28756 VSS.n2571 VSS.n2570 0.00658571
R28757 VSS.n2572 VSS.n2571 0.00658571
R28758 VSS.n2572 VSS.n2531 0.00658571
R28759 VSS.n2578 VSS.n2531 0.00658571
R28760 VSS.n2579 VSS.n2578 0.00658571
R28761 VSS.n2580 VSS.n2579 0.00658571
R28762 VSS.n2580 VSS.n2527 0.00658571
R28763 VSS.n2586 VSS.n2527 0.00658571
R28764 VSS.n2587 VSS.n2586 0.00658571
R28765 VSS.n2588 VSS.n2587 0.00658571
R28766 VSS.n2588 VSS.n2523 0.00658571
R28767 VSS.n2594 VSS.n2523 0.00658571
R28768 VSS.n2595 VSS.n2594 0.00658571
R28769 VSS.n2596 VSS.n2595 0.00658571
R28770 VSS.n2596 VSS.n2519 0.00658571
R28771 VSS.n2602 VSS.n2519 0.00658571
R28772 VSS.n2603 VSS.n2602 0.00658571
R28773 VSS.n2604 VSS.n2603 0.00658571
R28774 VSS.n2604 VSS.n2515 0.00658571
R28775 VSS.n2610 VSS.n2515 0.00658571
R28776 VSS.n2611 VSS.n2610 0.00658571
R28777 VSS.n2612 VSS.n2611 0.00658571
R28778 VSS.n2612 VSS.n2511 0.00658571
R28779 VSS.n2618 VSS.n2511 0.00658571
R28780 VSS.n2619 VSS.n2618 0.00658571
R28781 VSS.n2620 VSS.n2619 0.00658571
R28782 VSS.n2620 VSS.n2507 0.00658571
R28783 VSS.n2626 VSS.n2507 0.00658571
R28784 VSS.n2627 VSS.n2626 0.00658571
R28785 VSS.n2628 VSS.n2627 0.00658571
R28786 VSS.n2628 VSS.n2503 0.00658571
R28787 VSS.n2634 VSS.n2503 0.00658571
R28788 VSS.n2635 VSS.n2634 0.00658571
R28789 VSS.n2636 VSS.n2635 0.00658571
R28790 VSS.n2636 VSS.n2499 0.00658571
R28791 VSS.n2642 VSS.n2499 0.00658571
R28792 VSS.n2643 VSS.n2642 0.00658571
R28793 VSS.n2644 VSS.n2643 0.00658571
R28794 VSS.n2644 VSS.n2495 0.00658571
R28795 VSS.n2650 VSS.n2495 0.00658571
R28796 VSS.n2651 VSS.n2650 0.00658571
R28797 VSS.n2652 VSS.n2651 0.00658571
R28798 VSS.n2652 VSS.n2491 0.00658571
R28799 VSS.n2658 VSS.n2491 0.00658571
R28800 VSS.n2659 VSS.n2658 0.00658571
R28801 VSS.n2660 VSS.n2659 0.00658571
R28802 VSS.n2660 VSS.n2487 0.00658571
R28803 VSS.n2666 VSS.n2487 0.00658571
R28804 VSS.n2667 VSS.n2666 0.00658571
R28805 VSS.n2668 VSS.n2667 0.00658571
R28806 VSS.n2668 VSS.n2483 0.00658571
R28807 VSS.n2674 VSS.n2483 0.00658571
R28808 VSS.n2675 VSS.n2674 0.00658571
R28809 VSS.n2677 VSS.n2675 0.00658571
R28810 VSS.n2677 VSS.n2676 0.00658571
R28811 VSS.n2676 VSS.n2480 0.00658571
R28812 VSS.n2480 VSS.n2478 0.00658571
R28813 VSS.n2685 VSS.n2478 0.00658571
R28814 VSS.n2694 VSS.n2693 0.00658571
R28815 VSS.n3376 VSS.n3375 0.00658571
R28816 VSS.n3375 VSS.n3374 0.00658571
R28817 VSS.n3374 VSS.n2896 0.00658571
R28818 VSS.n3368 VSS.n2896 0.00658571
R28819 VSS.n3368 VSS.n3367 0.00658571
R28820 VSS.n3367 VSS.n3366 0.00658571
R28821 VSS.n3366 VSS.n2901 0.00658571
R28822 VSS.n2989 VSS.n2901 0.00658571
R28823 VSS.n2990 VSS.n2989 0.00658571
R28824 VSS.n2990 VSS.n2981 0.00658571
R28825 VSS.n2998 VSS.n2981 0.00658571
R28826 VSS.n2999 VSS.n2998 0.00658571
R28827 VSS.n3000 VSS.n2999 0.00658571
R28828 VSS.n3000 VSS.n2927 0.00658571
R28829 VSS.n3347 VSS.n2927 0.00658571
R28830 VSS.n3347 VSS.n3346 0.00658571
R28831 VSS.n3346 VSS.n3345 0.00658571
R28832 VSS.n3345 VSS.n2928 0.00658571
R28833 VSS.n3062 VSS.n2928 0.00658571
R28834 VSS.n3062 VSS.n2954 0.00658571
R28835 VSS.n3329 VSS.n2954 0.00658571
R28836 VSS.n3329 VSS.n3328 0.00658571
R28837 VSS.n3328 VSS.n3327 0.00658571
R28838 VSS.n3327 VSS.n2955 0.00658571
R28839 VSS.n3105 VSS.n2955 0.00658571
R28840 VSS.n3123 VSS.n3105 0.00658571
R28841 VSS.n3124 VSS.n3123 0.00658571
R28842 VSS.n3126 VSS.n3124 0.00658571
R28843 VSS.n3126 VSS.n3125 0.00658571
R28844 VSS.n3125 VSS.n3085 0.00658571
R28845 VSS.n3300 VSS.n3085 0.00658571
R28846 VSS.n3300 VSS.n3299 0.00658571
R28847 VSS.n3299 VSS.n3298 0.00658571
R28848 VSS.n3298 VSS.n3086 0.00658571
R28849 VSS.n3150 VSS.n3086 0.00658571
R28850 VSS.n3284 VSS.n3150 0.00658571
R28851 VSS.n3284 VSS.n3283 0.00658571
R28852 VSS.n3283 VSS.n3282 0.00658571
R28853 VSS.n3282 VSS.n3151 0.00658571
R28854 VSS.n3242 VSS.n3151 0.00658571
R28855 VSS.n3242 VSS.n3241 0.00658571
R28856 VSS.n3241 VSS.n3240 0.00658571
R28857 VSS.n3240 VSS.n3157 0.00658571
R28858 VSS.n3234 VSS.n3157 0.00658571
R28859 VSS.n3234 VSS.n3233 0.00658571
R28860 VSS.n3233 VSS.n3232 0.00658571
R28861 VSS.n3232 VSS.n3161 0.00658571
R28862 VSS.n3226 VSS.n3161 0.00658571
R28863 VSS.n3226 VSS.n3225 0.00658571
R28864 VSS.n3225 VSS.n3224 0.00658571
R28865 VSS.n3224 VSS.n3165 0.00658571
R28866 VSS.n3218 VSS.n3165 0.00658571
R28867 VSS.n3218 VSS.n3217 0.00658571
R28868 VSS.n3217 VSS.n3216 0.00658571
R28869 VSS.n3216 VSS.n3169 0.00658571
R28870 VSS.n3210 VSS.n3169 0.00658571
R28871 VSS.n3210 VSS.n3209 0.00658571
R28872 VSS.n3209 VSS.n3208 0.00658571
R28873 VSS.n3208 VSS.n3173 0.00658571
R28874 VSS.n3202 VSS.n3173 0.00658571
R28875 VSS.n3202 VSS.n3201 0.00658571
R28876 VSS.n3201 VSS.n3200 0.00658571
R28877 VSS.n3200 VSS.n3177 0.00658571
R28878 VSS.n3194 VSS.n3177 0.00658571
R28879 VSS.n3194 VSS.n3193 0.00658571
R28880 VSS.n3193 VSS.n3192 0.00658571
R28881 VSS.n3192 VSS.n3181 0.00658571
R28882 VSS.n3186 VSS.n3181 0.00658571
R28883 VSS.n3186 VSS.n3185 0.00658571
R28884 VSS.n2824 VSS.n2821 0.00658571
R28885 VSS.n3720 VSS.n2824 0.00658571
R28886 VSS.n3720 VSS.n3719 0.00658571
R28887 VSS.n3719 VSS.n3718 0.00658571
R28888 VSS.n3718 VSS.n2825 0.00658571
R28889 VSS.n3710 VSS.n2825 0.00658571
R28890 VSS.n3710 VSS.n3709 0.00658571
R28891 VSS.n3709 VSS.n3708 0.00658571
R28892 VSS.n3708 VSS.n2842 0.00658571
R28893 VSS.n3702 VSS.n2842 0.00658571
R28894 VSS.n3702 VSS.n3701 0.00658571
R28895 VSS.n3701 VSS.n3700 0.00658571
R28896 VSS.n3700 VSS.n2846 0.00658571
R28897 VSS.n3694 VSS.n2846 0.00658571
R28898 VSS.n3694 VSS.n3693 0.00658571
R28899 VSS.n3693 VSS.n3692 0.00658571
R28900 VSS.n3692 VSS.n2850 0.00658571
R28901 VSS.n3686 VSS.n2850 0.00658571
R28902 VSS.n3686 VSS.n3685 0.00658571
R28903 VSS.n3685 VSS.n3684 0.00658571
R28904 VSS.n3684 VSS.n2854 0.00658571
R28905 VSS.n3678 VSS.n2854 0.00658571
R28906 VSS.n3678 VSS.n3677 0.00658571
R28907 VSS.n3677 VSS.n3676 0.00658571
R28908 VSS.n3676 VSS.n2858 0.00658571
R28909 VSS.n3670 VSS.n2858 0.00658571
R28910 VSS.n3670 VSS.n3669 0.00658571
R28911 VSS.n3669 VSS.n3668 0.00658571
R28912 VSS.n3668 VSS.n2862 0.00658571
R28913 VSS.n3662 VSS.n2862 0.00658571
R28914 VSS.n3662 VSS.n3661 0.00658571
R28915 VSS.n3661 VSS.n3660 0.00658571
R28916 VSS.n3660 VSS.n2866 0.00658571
R28917 VSS.n3654 VSS.n2866 0.00658571
R28918 VSS.n3654 VSS.n3653 0.00658571
R28919 VSS.n3653 VSS.n3652 0.00658571
R28920 VSS.n3652 VSS.n2870 0.00658571
R28921 VSS.n3646 VSS.n2870 0.00658571
R28922 VSS.n3646 VSS.n3645 0.00658571
R28923 VSS.n3645 VSS.n3644 0.00658571
R28924 VSS.n3644 VSS.n2874 0.00658571
R28925 VSS.n3554 VSS.n2874 0.00658571
R28926 VSS.n3555 VSS.n3554 0.00658571
R28927 VSS.n3635 VSS.n3555 0.00658571
R28928 VSS.n3635 VSS.n3634 0.00658571
R28929 VSS.n3634 VSS.n3633 0.00658571
R28930 VSS.n3633 VSS.n3556 0.00658571
R28931 VSS.n3627 VSS.n3556 0.00658571
R28932 VSS.n3627 VSS.n3626 0.00658571
R28933 VSS.n3626 VSS.n3625 0.00658571
R28934 VSS.n3625 VSS.n3560 0.00658571
R28935 VSS.n3619 VSS.n3560 0.00658571
R28936 VSS.n3619 VSS.n3618 0.00658571
R28937 VSS.n3618 VSS.n3617 0.00658571
R28938 VSS.n3617 VSS.n3564 0.00658571
R28939 VSS.n3611 VSS.n3564 0.00658571
R28940 VSS.n3611 VSS.n3610 0.00658571
R28941 VSS.n3610 VSS.n3609 0.00658571
R28942 VSS.n3609 VSS.n3568 0.00658571
R28943 VSS.n3603 VSS.n3568 0.00658571
R28944 VSS.n3603 VSS.n3602 0.00658571
R28945 VSS.n3602 VSS.n3601 0.00658571
R28946 VSS.n3601 VSS.n3572 0.00658571
R28947 VSS.n3595 VSS.n3572 0.00658571
R28948 VSS.n3595 VSS.n3594 0.00658571
R28949 VSS.n3594 VSS.n3593 0.00658571
R28950 VSS.n3593 VSS.n3576 0.00658571
R28951 VSS.n3587 VSS.n3576 0.00658571
R28952 VSS.n3587 VSS.n3586 0.00658571
R28953 VSS.n3586 VSS.n3585 0.00658571
R28954 VSS.n3585 VSS.n3580 0.00658571
R28955 VSS.n2059 VSS.n2058 0.00658571
R28956 VSS.n2058 VSS.n2057 0.00658571
R28957 VSS.n2057 VSS.n1615 0.00658571
R28958 VSS.n2051 VSS.n1615 0.00658571
R28959 VSS.n2051 VSS.n2050 0.00658571
R28960 VSS.n2050 VSS.n2049 0.00658571
R28961 VSS.n2049 VSS.n1620 0.00658571
R28962 VSS.n1637 VSS.n1620 0.00658571
R28963 VSS.n2035 VSS.n1637 0.00658571
R28964 VSS.n2035 VSS.n2034 0.00658571
R28965 VSS.n2034 VSS.n2033 0.00658571
R28966 VSS.n2033 VSS.n1638 0.00658571
R28967 VSS.n2027 VSS.n1638 0.00658571
R28968 VSS.n2027 VSS.n2026 0.00658571
R28969 VSS.n2026 VSS.n2025 0.00658571
R28970 VSS.n2025 VSS.n1646 0.00658571
R28971 VSS.n1654 VSS.n1646 0.00658571
R28972 VSS.n2015 VSS.n1654 0.00658571
R28973 VSS.n2015 VSS.n2014 0.00658571
R28974 VSS.n2014 VSS.n2013 0.00658571
R28975 VSS.n2013 VSS.n1655 0.00658571
R28976 VSS.n1668 VSS.n1655 0.00658571
R28977 VSS.n2002 VSS.n1668 0.00658571
R28978 VSS.n2002 VSS.n2001 0.00658571
R28979 VSS.n2001 VSS.n2000 0.00658571
R28980 VSS.n2000 VSS.n1669 0.00658571
R28981 VSS.n1994 VSS.n1669 0.00658571
R28982 VSS.n1994 VSS.n1993 0.00658571
R28983 VSS.n1993 VSS.n1992 0.00658571
R28984 VSS.n1992 VSS.n1673 0.00658571
R28985 VSS.n1983 VSS.n1673 0.00658571
R28986 VSS.n1983 VSS.n1982 0.00658571
R28987 VSS.n1982 VSS.n1981 0.00658571
R28988 VSS.n1981 VSS.n1680 0.00658571
R28989 VSS.n1693 VSS.n1680 0.00658571
R28990 VSS.n1970 VSS.n1693 0.00658571
R28991 VSS.n1970 VSS.n1969 0.00658571
R28992 VSS.n1969 VSS.n1968 0.00658571
R28993 VSS.n1968 VSS.n1694 0.00658571
R28994 VSS.n1962 VSS.n1694 0.00658571
R28995 VSS.n1962 VSS.n1961 0.00658571
R28996 VSS.n1961 VSS.n1960 0.00658571
R28997 VSS.n1960 VSS.n1698 0.00658571
R28998 VSS.n1711 VSS.n1698 0.00658571
R28999 VSS.n1947 VSS.n1711 0.00658571
R29000 VSS.n1947 VSS.n1946 0.00658571
R29001 VSS.n1946 VSS.n1945 0.00658571
R29002 VSS.n1945 VSS.n1712 0.00658571
R29003 VSS.n1932 VSS.n1712 0.00658571
R29004 VSS.n1932 VSS.n1931 0.00658571
R29005 VSS.n1931 VSS.n1930 0.00658571
R29006 VSS.n1930 VSS.n1718 0.00658571
R29007 VSS.n1924 VSS.n1718 0.00658571
R29008 VSS.n1924 VSS.n1923 0.00658571
R29009 VSS.n1923 VSS.n1922 0.00658571
R29010 VSS.n1922 VSS.n1722 0.00658571
R29011 VSS.n1753 VSS.n1722 0.00658571
R29012 VSS.n1909 VSS.n1753 0.00658571
R29013 VSS.n1909 VSS.n1908 0.00658571
R29014 VSS.n1908 VSS.n1907 0.00658571
R29015 VSS.n1907 VSS.n1754 0.00658571
R29016 VSS.n1894 VSS.n1754 0.00658571
R29017 VSS.n1894 VSS.n1893 0.00658571
R29018 VSS.n1893 VSS.n1892 0.00658571
R29019 VSS.n1892 VSS.n1760 0.00658571
R29020 VSS.n1886 VSS.n1760 0.00658571
R29021 VSS.n1886 VSS.n1885 0.00658571
R29022 VSS.n1885 VSS.n1884 0.00658571
R29023 VSS.n1884 VSS.n1764 0.00658571
R29024 VSS.n1781 VSS.n1764 0.00658571
R29025 VSS.n1870 VSS.n1781 0.00658571
R29026 VSS.n1870 VSS.n1869 0.00658571
R29027 VSS.n1869 VSS.n1868 0.00658571
R29028 VSS.n1868 VSS.n1782 0.00658571
R29029 VSS.n1862 VSS.n1782 0.00658571
R29030 VSS.n1862 VSS.n1861 0.00658571
R29031 VSS.n1861 VSS.n1860 0.00658571
R29032 VSS.n1860 VSS.n1790 0.00658571
R29033 VSS.n1851 VSS.n1790 0.00658571
R29034 VSS.n1851 VSS.n1850 0.00658571
R29035 VSS.n1850 VSS.n1849 0.00658571
R29036 VSS.n1849 VSS.n1823 0.00658571
R29037 VSS.n1843 VSS.n1823 0.00658571
R29038 VSS.n1843 VSS.n1842 0.00658571
R29039 VSS.n1842 VSS.n1841 0.00658571
R29040 VSS.n1836 VSS.n1835 0.00658571
R29041 VSS.n1584 VSS.n1583 0.00658571
R29042 VSS.n1583 VSS.n1582 0.00658571
R29043 VSS.n1582 VSS.n1303 0.00658571
R29044 VSS.n1576 VSS.n1303 0.00658571
R29045 VSS.n1576 VSS.n1575 0.00658571
R29046 VSS.n1575 VSS.n1574 0.00658571
R29047 VSS.n1574 VSS.n1307 0.00658571
R29048 VSS.n1568 VSS.n1307 0.00658571
R29049 VSS.n1568 VSS.n1567 0.00658571
R29050 VSS.n1567 VSS.n1566 0.00658571
R29051 VSS.n1566 VSS.n1311 0.00658571
R29052 VSS.n1560 VSS.n1311 0.00658571
R29053 VSS.n1560 VSS.n1559 0.00658571
R29054 VSS.n1559 VSS.n1558 0.00658571
R29055 VSS.n1558 VSS.n1315 0.00658571
R29056 VSS.n1552 VSS.n1315 0.00658571
R29057 VSS.n1552 VSS.n1551 0.00658571
R29058 VSS.n1551 VSS.n1550 0.00658571
R29059 VSS.n1550 VSS.n1319 0.00658571
R29060 VSS.n1544 VSS.n1319 0.00658571
R29061 VSS.n1544 VSS.n1543 0.00658571
R29062 VSS.n1543 VSS.n1542 0.00658571
R29063 VSS.n1542 VSS.n1323 0.00658571
R29064 VSS.n1536 VSS.n1323 0.00658571
R29065 VSS.n1536 VSS.n1535 0.00658571
R29066 VSS.n1535 VSS.n1534 0.00658571
R29067 VSS.n1534 VSS.n1327 0.00658571
R29068 VSS.n1528 VSS.n1327 0.00658571
R29069 VSS.n1528 VSS.n1527 0.00658571
R29070 VSS.n1527 VSS.n1526 0.00658571
R29071 VSS.n1526 VSS.n1331 0.00658571
R29072 VSS.n1520 VSS.n1331 0.00658571
R29073 VSS.n1520 VSS.n1519 0.00658571
R29074 VSS.n1519 VSS.n1518 0.00658571
R29075 VSS.n1518 VSS.n1335 0.00658571
R29076 VSS.n1512 VSS.n1335 0.00658571
R29077 VSS.n1512 VSS.n1511 0.00658571
R29078 VSS.n1511 VSS.n1510 0.00658571
R29079 VSS.n1510 VSS.n1339 0.00658571
R29080 VSS.n1504 VSS.n1339 0.00658571
R29081 VSS.n1504 VSS.n1503 0.00658571
R29082 VSS.n1503 VSS.n1502 0.00658571
R29083 VSS.n1502 VSS.n1343 0.00658571
R29084 VSS.n1496 VSS.n1343 0.00658571
R29085 VSS.n1496 VSS.n1495 0.00658571
R29086 VSS.n1495 VSS.n1494 0.00658571
R29087 VSS.n1494 VSS.n1347 0.00658571
R29088 VSS.n1488 VSS.n1347 0.00658571
R29089 VSS.n1488 VSS.n1487 0.00658571
R29090 VSS.n1487 VSS.n1486 0.00658571
R29091 VSS.n1486 VSS.n1351 0.00658571
R29092 VSS.n1480 VSS.n1351 0.00658571
R29093 VSS.n1480 VSS.n1479 0.00658571
R29094 VSS.n1479 VSS.n1478 0.00658571
R29095 VSS.n1478 VSS.n1355 0.00658571
R29096 VSS.n1472 VSS.n1355 0.00658571
R29097 VSS.n1472 VSS.n1471 0.00658571
R29098 VSS.n1471 VSS.n1470 0.00658571
R29099 VSS.n1470 VSS.n1359 0.00658571
R29100 VSS.n1464 VSS.n1359 0.00658571
R29101 VSS.n1464 VSS.n1463 0.00658571
R29102 VSS.n1463 VSS.n1462 0.00658571
R29103 VSS.n1462 VSS.n1363 0.00658571
R29104 VSS.n1456 VSS.n1363 0.00658571
R29105 VSS.n1456 VSS.n1455 0.00658571
R29106 VSS.n1455 VSS.n1454 0.00658571
R29107 VSS.n1454 VSS.n1367 0.00658571
R29108 VSS.n1448 VSS.n1367 0.00658571
R29109 VSS.n1448 VSS.n1447 0.00658571
R29110 VSS.n1447 VSS.n1446 0.00658571
R29111 VSS.n1446 VSS.n1371 0.00658571
R29112 VSS.n1440 VSS.n1371 0.00658571
R29113 VSS.n1440 VSS.n1439 0.00658571
R29114 VSS.n1439 VSS.n1438 0.00658571
R29115 VSS.n1438 VSS.n1375 0.00658571
R29116 VSS.n1432 VSS.n1375 0.00658571
R29117 VSS.n1432 VSS.n1431 0.00658571
R29118 VSS.n1431 VSS.n1430 0.00658571
R29119 VSS.n1430 VSS.n1379 0.00658571
R29120 VSS.n1424 VSS.n1379 0.00658571
R29121 VSS.n1424 VSS.n1423 0.00658571
R29122 VSS.n1423 VSS.n1422 0.00658571
R29123 VSS.n1422 VSS.n1383 0.00658571
R29124 VSS.n1416 VSS.n1383 0.00658571
R29125 VSS.n1416 VSS.n1415 0.00658571
R29126 VSS.n1415 VSS.n1414 0.00658571
R29127 VSS.n1414 VSS.n1387 0.00658571
R29128 VSS.n1408 VSS.n1387 0.00658571
R29129 VSS.n1408 VSS.n1407 0.00658571
R29130 VSS.n1407 VSS.n1406 0.00658571
R29131 VSS.n1406 VSS.n1391 0.00658571
R29132 VSS.n1400 VSS.n1391 0.00658571
R29133 VSS.n1400 VSS.n1399 0.00658571
R29134 VSS.n1399 VSS.n1398 0.00658571
R29135 VSS.n4236 VSS.n2381 0.00658571
R29136 VSS.n4236 VSS.n4235 0.00658571
R29137 VSS.n4235 VSS.n4234 0.00658571
R29138 VSS.n4234 VSS.n2382 0.00658571
R29139 VSS.n4227 VSS.n2382 0.00658571
R29140 VSS.n4227 VSS.n4226 0.00658571
R29141 VSS.n4226 VSS.n4225 0.00658571
R29142 VSS.n4225 VSS.n2386 0.00658571
R29143 VSS.n4217 VSS.n2386 0.00658571
R29144 VSS.n4217 VSS.n4216 0.00658571
R29145 VSS.n4216 VSS.n4215 0.00658571
R29146 VSS.n4215 VSS.n2390 0.00658571
R29147 VSS.n4209 VSS.n2390 0.00658571
R29148 VSS.n4209 VSS.n4208 0.00658571
R29149 VSS.n4208 VSS.n4207 0.00658571
R29150 VSS.n4207 VSS.n2395 0.00658571
R29151 VSS.n4199 VSS.n2395 0.00658571
R29152 VSS.n4199 VSS.n4198 0.00658571
R29153 VSS.n4198 VSS.n4197 0.00658571
R29154 VSS.n4197 VSS.n2400 0.00658571
R29155 VSS.n4191 VSS.n2400 0.00658571
R29156 VSS.n4191 VSS.n4190 0.00658571
R29157 VSS.n4190 VSS.n4189 0.00658571
R29158 VSS.n4189 VSS.n2405 0.00658571
R29159 VSS.n4168 VSS.n2405 0.00658571
R29160 VSS.n4168 VSS.n4167 0.00658571
R29161 VSS.n4167 VSS.n4166 0.00658571
R29162 VSS.n4166 VSS.n2416 0.00658571
R29163 VSS.n4160 VSS.n2416 0.00658571
R29164 VSS.n4160 VSS.n4159 0.00658571
R29165 VSS.n4159 VSS.n4158 0.00658571
R29166 VSS.n4158 VSS.n2420 0.00658571
R29167 VSS.n4152 VSS.n2420 0.00658571
R29168 VSS.n4152 VSS.n4151 0.00658571
R29169 VSS.n4151 VSS.n4150 0.00658571
R29170 VSS.n4150 VSS.n2424 0.00658571
R29171 VSS.n4097 VSS.n2424 0.00658571
R29172 VSS.n4099 VSS.n4097 0.00658571
R29173 VSS.n4099 VSS.n4098 0.00658571
R29174 VSS.n4098 VSS.n2441 0.00658571
R29175 VSS.n4110 VSS.n2441 0.00658571
R29176 VSS.n4111 VSS.n4110 0.00658571
R29177 VSS.n4112 VSS.n4111 0.00658571
R29178 VSS.n4112 VSS.n2437 0.00658571
R29179 VSS.n4120 VSS.n2437 0.00658571
R29180 VSS.n4121 VSS.n4120 0.00658571
R29181 VSS.n4136 VSS.n4121 0.00658571
R29182 VSS.n4136 VSS.n4135 0.00658571
R29183 VSS.n4135 VSS.n4134 0.00658571
R29184 VSS.n4134 VSS.n4122 0.00658571
R29185 VSS.n4127 VSS.n4122 0.00658571
R29186 VSS.n4127 VSS.n4126 0.00658571
R29187 VSS.n4126 VSS.n2247 0.00658571
R29188 VSS.n5234 VSS.n2247 0.00658571
R29189 VSS.n5234 VSS.n5233 0.00658571
R29190 VSS.n5233 VSS.n5232 0.00658571
R29191 VSS.n5232 VSS.n2248 0.00658571
R29192 VSS.n5226 VSS.n2248 0.00658571
R29193 VSS.n5226 VSS.n5225 0.00658571
R29194 VSS.n5225 VSS.n5224 0.00658571
R29195 VSS.n5224 VSS.n2253 0.00658571
R29196 VSS.n5218 VSS.n2253 0.00658571
R29197 VSS.n5218 VSS.n5217 0.00658571
R29198 VSS.n5217 VSS.n5216 0.00658571
R29199 VSS.n5216 VSS.n2257 0.00658571
R29200 VSS.n5210 VSS.n2257 0.00658571
R29201 VSS.n5210 VSS.n5209 0.00658571
R29202 VSS.n5209 VSS.n5208 0.00658571
R29203 VSS.n5208 VSS.n2261 0.00658571
R29204 VSS.n5202 VSS.n2261 0.00658571
R29205 VSS.n5202 VSS.n5201 0.00658571
R29206 VSS.n5201 VSS.n5200 0.00658571
R29207 VSS.n5200 VSS.n2265 0.00658571
R29208 VSS.n5194 VSS.n2265 0.00658571
R29209 VSS.n5194 VSS.n5193 0.00658571
R29210 VSS.n5193 VSS.n5192 0.00658571
R29211 VSS.n5192 VSS.n2269 0.00658571
R29212 VSS.n5186 VSS.n2269 0.00658571
R29213 VSS.n5186 VSS.n5185 0.00658571
R29214 VSS.n5185 VSS.n5184 0.00658571
R29215 VSS.n5184 VSS.n5173 0.00658571
R29216 VSS.n5178 VSS.n5173 0.00658571
R29217 VSS.n5178 VSS.n5177 0.00658571
R29218 VSS.n3256 VSS.n3254 0.00658108
R29219 VSS.n3022 VSS.n3011 0.00658108
R29220 VSS.n1622 VSS.n1618 0.00654286
R29221 VSS.n2047 VSS.n1623 0.00654286
R29222 VSS.n2046 VSS.n1624 0.00654286
R29223 VSS.n1633 VSS.n1632 0.00654286
R29224 VSS.n2038 VSS.n2037 0.00654286
R29225 VSS.n1640 VSS.n1634 0.00654286
R29226 VSS.n2031 VSS.n1643 0.00654286
R29227 VSS.n425 VSS.n319 0.0065
R29228 VSS.n953 VSS.n952 0.0065
R29229 VSS.n379 VSS.n378 0.0065
R29230 VSS.n713 VSS.n320 0.0065
R29231 VSS.n1105 VSS.n98 0.0065
R29232 VSS.n490 VSS.n320 0.0065
R29233 VSS.n378 VSS.n376 0.0065
R29234 VSS.n136 VSS.n131 0.0065
R29235 VSS.n291 VSS.n136 0.0065
R29236 VSS.n1105 VSS.n1104 0.0065
R29237 VSS.n579 VSS.n372 0.0065
R29238 VSS.n743 VSS.n319 0.0065
R29239 VSS.n952 VSS.n133 0.0065
R29240 VSS.n1108 VSS.n93 0.0065
R29241 VSS.n1108 VSS.n94 0.0065
R29242 VSS.n579 VSS.n578 0.0065
R29243 VSS.n5025 VSS.n4423 0.0065
R29244 VSS.n4969 VSS.n4498 0.0065
R29245 VSS.n4733 VSS.n4421 0.0065
R29246 VSS.n4795 VSS.n4794 0.0065
R29247 VSS VSS.n5707 0.00641429
R29248 VSS VSS.n2694 0.00641429
R29249 DVSS VSS.n1836 0.00641429
R29250 VSS.n571 VSS.n570 0.00640498
R29251 VSS.n3380 VSS.n3379 0.00635
R29252 VSS.n4107 VSS.n2443 0.00635
R29253 VSS.n4117 VSS.n2433 0.00635
R29254 VSS.n4139 VSS.n2433 0.00635
R29255 VSS.n4909 VSS.n4908 0.00626355
R29256 VSS.n4850 VSS.n4627 0.00626355
R29257 VSS.n3639 VSS.n2884 0.006125
R29258 VSS.n3535 VSS.n2877 0.006125
R29259 VSS.n3727 VSS.n2818 0.00609286
R29260 VSS.n2701 VSS 0.00609286
R29261 VSS VSS.n0 0.00609286
R29262 VSS.n2065 VSS.n1603 0.00602857
R29263 VSS.n2062 VSS.n2061 0.00602857
R29264 VSS.n1617 VSS.n1597 0.00602857
R29265 VSS.n5048 VSS.n4388 0.006
R29266 VSS.n4949 VSS.n4948 0.006
R29267 VSS.n4715 VSS.n4713 0.006
R29268 VSS.n4815 VSS.n4530 0.006
R29269 VSS.n5692 VSS.n18 0.0059878
R29270 VSS.n5689 VSS.n31 0.0059878
R29271 VSS.n1888 VSS.n1762 0.00596429
R29272 VSS.n1767 VSS.n1766 0.00596429
R29273 VSS.n1882 VSS.n1881 0.00596429
R29274 VSS.n1776 VSS.n1768 0.00596429
R29275 VSS.n1873 VSS.n1777 0.00596429
R29276 VSS.n1872 VSS.n1778 0.00596429
R29277 VSS.n1787 VSS.n1784 0.00596429
R29278 DVSS VSS.n5154 0.00585211
R29279 VSS.n4204 VSS.n4203 0.00583571
R29280 VSS.n4220 VSS.n4219 0.00570714
R29281 VSS.n3049 VSS.n2834 0.00561229
R29282 VSS.n2838 VSS.n2828 0.00561229
R29283 DVSS VSS.n4391 0.00559852
R29284 VSS.n4448 VSS.n4446 0.00559852
R29285 VSS.n4708 DVSS 0.00559852
R29286 VSS.n4748 VSS.n4747 0.00559852
R29287 VSS.n5680 VSS.n1171 0.00559091
R29288 VSS.n3007 VSS.n2920 0.00551429
R29289 VSS.n3003 VSS.n2922 0.00551429
R29290 VSS.n2977 VSS.n2919 0.00551429
R29291 VSS.n5069 VSS.n5068 0.0055
R29292 VSS.n4568 VSS.n4567 0.0055
R29293 VSS.n4693 VSS.n4362 0.0055
R29294 VSS.n4836 VSS.n4835 0.0055
R29295 VSS.n2687 VSS.n2686 0.00548841
R29296 VSS.n2315 VSS.n2314 0.00548841
R29297 VSS.n1830 VSS.n1829 0.00548841
R29298 VSS.n3440 VSS.n3439 0.00548841
R29299 VSS.n5 VSS.n4 0.00548841
R29300 VSS VSS.n2685 0.00538571
R29301 VSS.n1841 DVSS 0.00538571
R29302 VSS.n3307 VSS.n3080 0.00538571
R29303 VSS.n3303 VSS.n3302 0.00538571
R29304 VSS.n3088 VSS.n3076 0.00538571
R29305 VSS.n4638 VSS.n4409 0.00537685
R29306 VSS.n4722 VSS.n4639 0.00537685
R29307 VSS.n1880 VSS.n1769 0.00532927
R29308 VSS.n1874 VSS.n1775 0.00532927
R29309 VSS.n1917 VSS.n1727 0.00532927
R29310 VSS.n1901 VSS.n1900 0.00532927
R29311 VSS.n1955 VSS.n1703 0.00532927
R29312 VSS.n1939 VSS.n1938 0.00532927
R29313 VSS.n1736 VSS.n1677 0.00532927
R29314 VSS.n1977 VSS.n1976 0.00532927
R29315 VSS.n1730 VSS.n1650 0.00532927
R29316 VSS.n2009 VSS.n2008 0.00532927
R29317 VSS.n2045 VSS.n1625 0.00532927
R29318 VSS.n2039 VSS.n1631 0.00532927
R29319 VSS.n2894 VSS.n2817 0.00519286
R29320 VSS.n5237 VSS.n2243 0.00519286
R29321 VSS.n4282 VSS.n4281 0.00519286
R29322 VSS.n3048 VSS.n3047 0.00514674
R29323 VSS.n1169 VSS.n15 0.00505741
R29324 VSS.n15 VSS.n12 0.00505741
R29325 VSS.n1591 VSS.n1294 0.00505741
R29326 VSS.n1294 VSS.n1292 0.00505741
R29327 VSS.n3114 VSS.n2962 0.00504128
R29328 VSS.n3337 VSS.n2934 0.00504128
R29329 VSS.n5096 VSS.n4323 0.005
R29330 VSS.n5089 VSS.n4335 0.005
R29331 VSS.n4905 VSS.n4590 0.005
R29332 VSS.n4898 VSS.n4602 0.005
R29333 VSS.n4665 VSS.n4325 0.005
R29334 VSS.n4667 VSS.n4333 0.005
R29335 VSS.n4857 VSS.n4592 0.005
R29336 VSS.n4859 VSS.n4600 0.005
R29337 VSS.n915 VSS.n914 0.00498878
R29338 VSS.n1171 VSS.n1170 0.0049789
R29339 VSS.n1172 VSS.n1171 0.0049789
R29340 VSS.n2898 VSS.n2817 0.00493571
R29341 VSS.n5237 VSS.n5236 0.00493571
R29342 VSS.n4282 VSS.n2297 0.00493571
R29343 VSS.n3042 VSS.n2830 0.00489894
R29344 VSS.n3038 VSS.n2836 0.00489894
R29345 VSS.n3735 VSS.n2816 0.00476
R29346 VSS.n3735 VSS.n2814 0.00476
R29347 VSS.n3739 VSS.n2814 0.00476
R29348 VSS.n3739 VSS.n2812 0.00476
R29349 VSS.n3743 VSS.n2812 0.00476
R29350 VSS.n3743 VSS.n2810 0.00476
R29351 VSS.n3748 VSS.n2810 0.00476
R29352 VSS.n3748 VSS.n2808 0.00476
R29353 VSS.n3752 VSS.n2808 0.00476
R29354 VSS.n3752 VSS.n2806 0.00476
R29355 VSS.n3756 VSS.n2806 0.00476
R29356 VSS.n3756 VSS.n2804 0.00476
R29357 VSS.n3863 VSS.n2804 0.00476
R29358 VSS.n3863 VSS.n3862 0.00476
R29359 VSS.n3862 VSS.n3861 0.00476
R29360 VSS.n3861 VSS.n3762 0.00476
R29361 VSS.n3857 VSS.n3762 0.00476
R29362 VSS.n3857 VSS.n3856 0.00476
R29363 VSS.n3856 VSS.n3855 0.00476
R29364 VSS.n3855 VSS.n3768 0.00476
R29365 VSS.n3851 VSS.n3768 0.00476
R29366 VSS.n3851 VSS.n3850 0.00476
R29367 VSS.n3850 VSS.n3849 0.00476
R29368 VSS.n3849 VSS.n3774 0.00476
R29369 VSS.n3845 VSS.n3774 0.00476
R29370 VSS.n3845 VSS.n3844 0.00476
R29371 VSS.n3844 VSS.n3843 0.00476
R29372 VSS.n3843 VSS.n3781 0.00476
R29373 VSS.n3839 VSS.n3781 0.00476
R29374 VSS.n3839 VSS.n3838 0.00476
R29375 VSS.n3838 VSS.n3837 0.00476
R29376 VSS.n3837 VSS.n3787 0.00476
R29377 VSS.n3833 VSS.n3787 0.00476
R29378 VSS.n3833 VSS.n3832 0.00476
R29379 VSS.n3832 VSS.n3831 0.00476
R29380 VSS.n3831 VSS.n3793 0.00476
R29381 VSS.n3827 VSS.n3793 0.00476
R29382 VSS.n3827 VSS.n3826 0.00476
R29383 VSS.n3826 VSS.n3825 0.00476
R29384 VSS.n3825 VSS.n3799 0.00476
R29385 VSS.n3821 VSS.n3799 0.00476
R29386 VSS.n3821 VSS.n3820 0.00476
R29387 VSS.n3820 VSS.n3819 0.00476
R29388 VSS.n3819 VSS.n3805 0.00476
R29389 VSS.n3815 VSS.n3805 0.00476
R29390 VSS.n3815 VSS.n3814 0.00476
R29391 VSS.n3814 VSS.n3813 0.00476
R29392 VSS.n3813 VSS.n2116 0.00476
R29393 VSS.n5386 VSS.n2116 0.00476
R29394 VSS.n5386 VSS.n5385 0.00476
R29395 VSS.n5385 VSS.n5384 0.00476
R29396 VSS.n5384 VSS.n2120 0.00476
R29397 VSS.n5380 VSS.n2120 0.00476
R29398 VSS.n5380 VSS.n5379 0.00476
R29399 VSS.n5379 VSS.n5378 0.00476
R29400 VSS.n5378 VSS.n2126 0.00476
R29401 VSS.n5373 VSS.n2126 0.00476
R29402 VSS.n5373 VSS.n5372 0.00476
R29403 VSS.n5372 VSS.n5371 0.00476
R29404 VSS.n5371 VSS.n2133 0.00476
R29405 VSS.n5367 VSS.n2133 0.00476
R29406 VSS.n5367 VSS.n5366 0.00476
R29407 VSS.n5366 VSS.n2138 0.00476
R29408 VSS.n5362 VSS.n2138 0.00476
R29409 VSS.n5362 VSS.n5361 0.00476
R29410 VSS.n5361 VSS.n5360 0.00476
R29411 VSS.n5360 VSS.n2144 0.00476
R29412 VSS.n5356 VSS.n2144 0.00476
R29413 VSS.n5356 VSS.n5355 0.00476
R29414 VSS.n5355 VSS.n5354 0.00476
R29415 VSS.n5354 VSS.n2150 0.00476
R29416 VSS.n5350 VSS.n2150 0.00476
R29417 VSS.n5350 VSS.n5349 0.00476
R29418 VSS.n5349 VSS.n5348 0.00476
R29419 VSS.n5348 VSS.n2156 0.00476
R29420 VSS.n5344 VSS.n2156 0.00476
R29421 VSS.n5344 VSS.n5343 0.00476
R29422 VSS.n5342 VSS.n2162 0.00476
R29423 VSS.n2170 VSS.n2162 0.00476
R29424 VSS.n2170 VSS.n2169 0.00476
R29425 VSS.n576 VSS.n575 0.00476
R29426 VSS.n575 VSS.n390 0.00476
R29427 VSS.n521 VSS.n390 0.00476
R29428 VSS.n521 VSS.n520 0.00476
R29429 VSS.n520 VSS.n519 0.00476
R29430 VSS.n519 VSS.n396 0.00476
R29431 VSS.n515 VSS.n396 0.00476
R29432 VSS.n515 VSS.n514 0.00476
R29433 VSS.n514 VSS.n513 0.00476
R29434 VSS.n513 VSS.n402 0.00476
R29435 VSS.n509 VSS.n402 0.00476
R29436 VSS.n509 VSS.n508 0.00476
R29437 VSS.n508 VSS.n507 0.00476
R29438 VSS.n507 VSS.n408 0.00476
R29439 VSS.n503 VSS.n408 0.00476
R29440 VSS.n503 VSS.n502 0.00476
R29441 VSS.n502 VSS.n501 0.00476
R29442 VSS.n501 VSS.n414 0.00476
R29443 VSS.n497 VSS.n414 0.00476
R29444 VSS.n497 VSS.n496 0.00476
R29445 VSS.n496 VSS.n418 0.00476
R29446 VSS.n492 VSS.n418 0.00476
R29447 VSS.n492 VSS.n491 0.00476
R29448 VSS.n489 VSS.n424 0.00476
R29449 VSS.n485 VSS.n424 0.00476
R29450 VSS.n485 VSS.n484 0.00476
R29451 VSS.n484 VSS.n483 0.00476
R29452 VSS.n483 VSS.n431 0.00476
R29453 VSS.n479 VSS.n431 0.00476
R29454 VSS.n479 VSS.n478 0.00476
R29455 VSS.n478 VSS.n477 0.00476
R29456 VSS.n477 VSS.n437 0.00476
R29457 VSS.n473 VSS.n437 0.00476
R29458 VSS.n473 VSS.n472 0.00476
R29459 VSS.n472 VSS.n471 0.00476
R29460 VSS.n471 VSS.n443 0.00476
R29461 VSS.n467 VSS.n443 0.00476
R29462 VSS.n467 VSS.n466 0.00476
R29463 VSS.n466 VSS.n465 0.00476
R29464 VSS.n465 VSS.n449 0.00476
R29465 VSS.n461 VSS.n449 0.00476
R29466 VSS.n461 VSS.n460 0.00476
R29467 VSS.n460 VSS.n459 0.00476
R29468 VSS.n459 VSS.n456 0.00476
R29469 VSS.n456 VSS.n130 0.00476
R29470 VSS.n955 VSS.n130 0.00476
R29471 VSS.n960 VSS.n127 0.00476
R29472 VSS.n960 VSS.n125 0.00476
R29473 VSS.n965 VSS.n125 0.00476
R29474 VSS.n965 VSS.n123 0.00476
R29475 VSS.n969 VSS.n123 0.00476
R29476 VSS.n969 VSS.n121 0.00476
R29477 VSS.n973 VSS.n121 0.00476
R29478 VSS.n973 VSS.n119 0.00476
R29479 VSS.n977 VSS.n119 0.00476
R29480 VSS.n977 VSS.n117 0.00476
R29481 VSS.n981 VSS.n117 0.00476
R29482 VSS.n981 VSS.n115 0.00476
R29483 VSS.n985 VSS.n115 0.00476
R29484 VSS.n985 VSS.n113 0.00476
R29485 VSS.n989 VSS.n113 0.00476
R29486 VSS.n989 VSS.n111 0.00476
R29487 VSS.n993 VSS.n111 0.00476
R29488 VSS.n993 VSS.n109 0.00476
R29489 VSS.n997 VSS.n109 0.00476
R29490 VSS.n997 VSS.n107 0.00476
R29491 VSS.n1001 VSS.n107 0.00476
R29492 VSS.n1001 VSS.n102 0.00476
R29493 VSS.n1008 VSS.n102 0.00476
R29494 VSS.n1052 VSS.n1011 0.00476
R29495 VSS.n1048 VSS.n1011 0.00476
R29496 VSS.n1048 VSS.n1047 0.00476
R29497 VSS.n1047 VSS.n1046 0.00476
R29498 VSS.n1046 VSS.n1016 0.00476
R29499 VSS.n1042 VSS.n1016 0.00476
R29500 VSS.n1042 VSS.n1041 0.00476
R29501 VSS.n1041 VSS.n1040 0.00476
R29502 VSS.n1040 VSS.n1022 0.00476
R29503 VSS.n1036 VSS.n1022 0.00476
R29504 VSS.n1035 VSS.n1026 0.00476
R29505 VSS.n1031 VSS.n1026 0.00476
R29506 VSS.n1031 VSS.n1030 0.00476
R29507 VSS.n583 VSS.n371 0.00476
R29508 VSS.n583 VSS.n369 0.00476
R29509 VSS.n628 VSS.n369 0.00476
R29510 VSS.n628 VSS.n627 0.00476
R29511 VSS.n627 VSS.n626 0.00476
R29512 VSS.n626 VSS.n589 0.00476
R29513 VSS.n622 VSS.n589 0.00476
R29514 VSS.n622 VSS.n621 0.00476
R29515 VSS.n621 VSS.n620 0.00476
R29516 VSS.n620 VSS.n595 0.00476
R29517 VSS.n616 VSS.n595 0.00476
R29518 VSS.n616 VSS.n615 0.00476
R29519 VSS.n615 VSS.n614 0.00476
R29520 VSS.n614 VSS.n601 0.00476
R29521 VSS.n610 VSS.n601 0.00476
R29522 VSS.n610 VSS.n609 0.00476
R29523 VSS.n609 VSS.n608 0.00476
R29524 VSS.n608 VSS.n328 0.00476
R29525 VSS.n754 VSS.n328 0.00476
R29526 VSS.n754 VSS.n326 0.00476
R29527 VSS.n758 VSS.n326 0.00476
R29528 VSS.n758 VSS.n324 0.00476
R29529 VSS.n762 VSS.n324 0.00476
R29530 VSS.n766 VSS.n318 0.00476
R29531 VSS.n770 VSS.n318 0.00476
R29532 VSS.n770 VSS.n316 0.00476
R29533 VSS.n774 VSS.n316 0.00476
R29534 VSS.n774 VSS.n314 0.00476
R29535 VSS.n778 VSS.n314 0.00476
R29536 VSS.n778 VSS.n312 0.00476
R29537 VSS.n782 VSS.n312 0.00476
R29538 VSS.n782 VSS.n310 0.00476
R29539 VSS.n786 VSS.n310 0.00476
R29540 VSS.n786 VSS.n308 0.00476
R29541 VSS.n821 VSS.n308 0.00476
R29542 VSS.n821 VSS.n820 0.00476
R29543 VSS.n820 VSS.n819 0.00476
R29544 VSS.n819 VSS.n792 0.00476
R29545 VSS.n815 VSS.n792 0.00476
R29546 VSS.n815 VSS.n814 0.00476
R29547 VSS.n814 VSS.n813 0.00476
R29548 VSS.n813 VSS.n798 0.00476
R29549 VSS.n809 VSS.n798 0.00476
R29550 VSS.n809 VSS.n808 0.00476
R29551 VSS.n808 VSS.n807 0.00476
R29552 VSS.n807 VSS.n805 0.00476
R29553 VSS.n950 VSS.n949 0.00476
R29554 VSS.n949 VSS.n948 0.00476
R29555 VSS.n948 VSS.n140 0.00476
R29556 VSS.n944 VSS.n140 0.00476
R29557 VSS.n944 VSS.n943 0.00476
R29558 VSS.n943 VSS.n145 0.00476
R29559 VSS.n939 VSS.n145 0.00476
R29560 VSS.n939 VSS.n938 0.00476
R29561 VSS.n938 VSS.n937 0.00476
R29562 VSS.n937 VSS.n151 0.00476
R29563 VSS.n933 VSS.n151 0.00476
R29564 VSS.n933 VSS.n932 0.00476
R29565 VSS.n932 VSS.n931 0.00476
R29566 VSS.n931 VSS.n157 0.00476
R29567 VSS.n927 VSS.n157 0.00476
R29568 VSS.n927 VSS.n926 0.00476
R29569 VSS.n926 VSS.n925 0.00476
R29570 VSS.n925 VSS.n163 0.00476
R29571 VSS.n921 VSS.n163 0.00476
R29572 VSS.n921 VSS.n920 0.00476
R29573 VSS.n920 VSS.n919 0.00476
R29574 VSS.n919 VSS.n96 0.00476
R29575 VSS.n1106 VSS.n96 0.00476
R29576 VSS.n1111 VSS.n92 0.00476
R29577 VSS.n1111 VSS.n90 0.00476
R29578 VSS.n1115 VSS.n90 0.00476
R29579 VSS.n1115 VSS.n88 0.00476
R29580 VSS.n1119 VSS.n88 0.00476
R29581 VSS.n1119 VSS.n86 0.00476
R29582 VSS.n1123 VSS.n86 0.00476
R29583 VSS.n1123 VSS.n84 0.00476
R29584 VSS.n1127 VSS.n84 0.00476
R29585 VSS.n1127 VSS.n82 0.00476
R29586 VSS.n1131 VSS.n82 0.00476
R29587 VSS.n1135 VSS.n80 0.00476
R29588 VSS.n1135 VSS.n78 0.00476
R29589 VSS.n383 VSS.n351 0.00476
R29590 VSS.n672 VSS.n351 0.00476
R29591 VSS.n672 VSS.n349 0.00476
R29592 VSS.n676 VSS.n349 0.00476
R29593 VSS.n676 VSS.n347 0.00476
R29594 VSS.n680 VSS.n347 0.00476
R29595 VSS.n680 VSS.n345 0.00476
R29596 VSS.n684 VSS.n345 0.00476
R29597 VSS.n684 VSS.n343 0.00476
R29598 VSS.n688 VSS.n343 0.00476
R29599 VSS.n688 VSS.n341 0.00476
R29600 VSS.n692 VSS.n341 0.00476
R29601 VSS.n692 VSS.n339 0.00476
R29602 VSS.n696 VSS.n339 0.00476
R29603 VSS.n696 VSS.n337 0.00476
R29604 VSS.n700 VSS.n337 0.00476
R29605 VSS.n700 VSS.n335 0.00476
R29606 VSS.n704 VSS.n335 0.00476
R29607 VSS.n704 VSS.n333 0.00476
R29608 VSS.n748 VSS.n333 0.00476
R29609 VSS.n748 VSS.n747 0.00476
R29610 VSS.n747 VSS.n746 0.00476
R29611 VSS.n746 VSS.n711 0.00476
R29612 VSS.n741 VSS.n740 0.00476
R29613 VSS.n740 VSS.n739 0.00476
R29614 VSS.n739 VSS.n717 0.00476
R29615 VSS.n735 VSS.n717 0.00476
R29616 VSS.n735 VSS.n734 0.00476
R29617 VSS.n734 VSS.n733 0.00476
R29618 VSS.n733 VSS.n723 0.00476
R29619 VSS.n729 VSS.n723 0.00476
R29620 VSS.n729 VSS.n728 0.00476
R29621 VSS.n728 VSS.n303 0.00476
R29622 VSS.n827 VSS.n303 0.00476
R29623 VSS.n827 VSS.n301 0.00476
R29624 VSS.n831 VSS.n301 0.00476
R29625 VSS.n831 VSS.n299 0.00476
R29626 VSS.n835 VSS.n299 0.00476
R29627 VSS.n835 VSS.n297 0.00476
R29628 VSS.n839 VSS.n297 0.00476
R29629 VSS.n839 VSS.n295 0.00476
R29630 VSS.n843 VSS.n295 0.00476
R29631 VSS.n843 VSS.n293 0.00476
R29632 VSS.n847 VSS.n293 0.00476
R29633 VSS.n847 VSS.n290 0.00476
R29634 VSS.n851 VSS.n290 0.00476
R29635 VSS.n856 VSS.n288 0.00476
R29636 VSS.n856 VSS.n286 0.00476
R29637 VSS.n861 VSS.n286 0.00476
R29638 VSS.n861 VSS.n284 0.00476
R29639 VSS.n865 VSS.n284 0.00476
R29640 VSS.n865 VSS.n281 0.00476
R29641 VSS.n869 VSS.n281 0.00476
R29642 VSS.n869 VSS.n279 0.00476
R29643 VSS.n873 VSS.n279 0.00476
R29644 VSS.n873 VSS.n277 0.00476
R29645 VSS.n877 VSS.n277 0.00476
R29646 VSS.n877 VSS.n275 0.00476
R29647 VSS.n881 VSS.n275 0.00476
R29648 VSS.n881 VSS.n273 0.00476
R29649 VSS.n885 VSS.n273 0.00476
R29650 VSS.n885 VSS.n271 0.00476
R29651 VSS.n889 VSS.n271 0.00476
R29652 VSS.n889 VSS.n269 0.00476
R29653 VSS.n893 VSS.n269 0.00476
R29654 VSS.n893 VSS.n267 0.00476
R29655 VSS.n899 VSS.n267 0.00476
R29656 VSS.n899 VSS.n898 0.00476
R29657 VSS.n898 VSS.n99 0.00476
R29658 VSS.n1103 VSS.n1058 0.00476
R29659 VSS.n1099 VSS.n1058 0.00476
R29660 VSS.n1099 VSS.n1098 0.00476
R29661 VSS.n1098 VSS.n1097 0.00476
R29662 VSS.n1097 VSS.n1064 0.00476
R29663 VSS.n1093 VSS.n1064 0.00476
R29664 VSS.n1093 VSS.n1092 0.00476
R29665 VSS.n1092 VSS.n1091 0.00476
R29666 VSS.n1091 VSS.n1070 0.00476
R29667 VSS.n1087 VSS.n1070 0.00476
R29668 VSS.n1086 VSS.n1074 0.00476
R29669 VSS.n1082 VSS.n1074 0.00476
R29670 VSS.n1082 VSS.n1081 0.00476
R29671 VSS.n671 VSS.n352 0.00476
R29672 VSS.n677 VSS.n348 0.00476
R29673 VSS.n678 VSS.n677 0.00476
R29674 VSS.n679 VSS.n678 0.00476
R29675 VSS.n679 VSS.n344 0.00476
R29676 VSS.n685 VSS.n344 0.00476
R29677 VSS.n686 VSS.n685 0.00476
R29678 VSS.n687 VSS.n686 0.00476
R29679 VSS.n687 VSS.n340 0.00476
R29680 VSS.n693 VSS.n340 0.00476
R29681 VSS.n694 VSS.n693 0.00476
R29682 VSS.n695 VSS.n694 0.00476
R29683 VSS.n695 VSS.n336 0.00476
R29684 VSS.n701 VSS.n336 0.00476
R29685 VSS.n702 VSS.n701 0.00476
R29686 VSS.n703 VSS.n702 0.00476
R29687 VSS.n703 VSS.n331 0.00476
R29688 VSS.n749 VSS.n332 0.00476
R29689 VSS.n745 VSS.n332 0.00476
R29690 VSS.n745 VSS.n744 0.00476
R29691 VSS.n742 VSS.n712 0.00476
R29692 VSS.n738 VSS.n712 0.00476
R29693 VSS.n738 VSS.n737 0.00476
R29694 VSS.n737 VSS.n736 0.00476
R29695 VSS.n736 VSS.n718 0.00476
R29696 VSS.n732 VSS.n718 0.00476
R29697 VSS.n732 VSS.n731 0.00476
R29698 VSS.n731 VSS.n730 0.00476
R29699 VSS.n730 VSS.n724 0.00476
R29700 VSS.n724 VSS.n304 0.00476
R29701 VSS.n826 VSS.n304 0.00476
R29702 VSS.n832 VSS.n300 0.00476
R29703 VSS.n833 VSS.n832 0.00476
R29704 VSS.n834 VSS.n833 0.00476
R29705 VSS.n834 VSS.n296 0.00476
R29706 VSS.n840 VSS.n296 0.00476
R29707 VSS.n841 VSS.n840 0.00476
R29708 VSS.n842 VSS.n841 0.00476
R29709 VSS.n842 VSS.n292 0.00476
R29710 VSS.n848 VSS.n292 0.00476
R29711 VSS.n849 VSS.n848 0.00476
R29712 VSS.n850 VSS.n849 0.00476
R29713 VSS.n857 VSS.n287 0.00476
R29714 VSS.n858 VSS.n857 0.00476
R29715 VSS.n860 VSS.n858 0.00476
R29716 VSS.n860 VSS.n859 0.00476
R29717 VSS.n867 VSS.n866 0.00476
R29718 VSS.n868 VSS.n867 0.00476
R29719 VSS.n868 VSS.n278 0.00476
R29720 VSS.n874 VSS.n278 0.00476
R29721 VSS.n875 VSS.n874 0.00476
R29722 VSS.n876 VSS.n875 0.00476
R29723 VSS.n876 VSS.n274 0.00476
R29724 VSS.n882 VSS.n274 0.00476
R29725 VSS.n883 VSS.n882 0.00476
R29726 VSS.n884 VSS.n883 0.00476
R29727 VSS.n884 VSS.n270 0.00476
R29728 VSS.n890 VSS.n270 0.00476
R29729 VSS.n891 VSS.n890 0.00476
R29730 VSS.n892 VSS.n891 0.00476
R29731 VSS.n892 VSS.n263 0.00476
R29732 VSS.n900 VSS.n266 0.00476
R29733 VSS.n1102 VSS.n1101 0.00476
R29734 VSS.n1101 VSS.n1100 0.00476
R29735 VSS.n1100 VSS.n1059 0.00476
R29736 VSS.n1096 VSS.n1059 0.00476
R29737 VSS.n1096 VSS.n1095 0.00476
R29738 VSS.n1095 VSS.n1094 0.00476
R29739 VSS.n1094 VSS.n1065 0.00476
R29740 VSS.n1090 VSS.n1065 0.00476
R29741 VSS.n1090 VSS.n1089 0.00476
R29742 VSS.n1089 VSS.n1088 0.00476
R29743 VSS.n1085 VSS.n1084 0.00476
R29744 VSS.n1084 VSS.n1083 0.00476
R29745 VSS.n1083 VSS.n1075 0.00476
R29746 VSS.n582 VSS.n367 0.00476
R29747 VSS.n629 VSS.n368 0.00476
R29748 VSS.n625 VSS.n368 0.00476
R29749 VSS.n625 VSS.n624 0.00476
R29750 VSS.n624 VSS.n623 0.00476
R29751 VSS.n623 VSS.n590 0.00476
R29752 VSS.n619 VSS.n590 0.00476
R29753 VSS.n619 VSS.n618 0.00476
R29754 VSS.n618 VSS.n617 0.00476
R29755 VSS.n617 VSS.n596 0.00476
R29756 VSS.n613 VSS.n596 0.00476
R29757 VSS.n613 VSS.n612 0.00476
R29758 VSS.n612 VSS.n611 0.00476
R29759 VSS.n611 VSS.n602 0.00476
R29760 VSS.n607 VSS.n602 0.00476
R29761 VSS.n607 VSS.n329 0.00476
R29762 VSS.n753 VSS.n329 0.00476
R29763 VSS.n759 VSS.n325 0.00476
R29764 VSS.n760 VSS.n759 0.00476
R29765 VSS.n761 VSS.n760 0.00476
R29766 VSS.n768 VSS.n767 0.00476
R29767 VSS.n769 VSS.n768 0.00476
R29768 VSS.n769 VSS.n315 0.00476
R29769 VSS.n775 VSS.n315 0.00476
R29770 VSS.n776 VSS.n775 0.00476
R29771 VSS.n777 VSS.n776 0.00476
R29772 VSS.n777 VSS.n311 0.00476
R29773 VSS.n783 VSS.n311 0.00476
R29774 VSS.n784 VSS.n783 0.00476
R29775 VSS.n785 VSS.n784 0.00476
R29776 VSS.n785 VSS.n306 0.00476
R29777 VSS.n822 VSS.n307 0.00476
R29778 VSS.n818 VSS.n307 0.00476
R29779 VSS.n818 VSS.n817 0.00476
R29780 VSS.n817 VSS.n816 0.00476
R29781 VSS.n816 VSS.n793 0.00476
R29782 VSS.n812 VSS.n793 0.00476
R29783 VSS.n812 VSS.n811 0.00476
R29784 VSS.n811 VSS.n810 0.00476
R29785 VSS.n810 VSS.n799 0.00476
R29786 VSS.n806 VSS.n799 0.00476
R29787 VSS.n806 VSS.n134 0.00476
R29788 VSS.n951 VSS.n135 0.00476
R29789 VSS.n947 VSS.n135 0.00476
R29790 VSS.n947 VSS.n946 0.00476
R29791 VSS.n946 VSS.n945 0.00476
R29792 VSS.n942 VSS.n941 0.00476
R29793 VSS.n941 VSS.n940 0.00476
R29794 VSS.n940 VSS.n146 0.00476
R29795 VSS.n936 VSS.n146 0.00476
R29796 VSS.n936 VSS.n935 0.00476
R29797 VSS.n935 VSS.n934 0.00476
R29798 VSS.n934 VSS.n152 0.00476
R29799 VSS.n930 VSS.n152 0.00476
R29800 VSS.n930 VSS.n929 0.00476
R29801 VSS.n929 VSS.n928 0.00476
R29802 VSS.n928 VSS.n158 0.00476
R29803 VSS.n924 VSS.n158 0.00476
R29804 VSS.n924 VSS.n923 0.00476
R29805 VSS.n923 VSS.n922 0.00476
R29806 VSS.n922 VSS.n164 0.00476
R29807 VSS.n918 VSS.n917 0.00476
R29808 VSS.n1110 VSS.n1109 0.00476
R29809 VSS.n1110 VSS.n89 0.00476
R29810 VSS.n1116 VSS.n89 0.00476
R29811 VSS.n1117 VSS.n1116 0.00476
R29812 VSS.n1118 VSS.n1117 0.00476
R29813 VSS.n1118 VSS.n85 0.00476
R29814 VSS.n1124 VSS.n85 0.00476
R29815 VSS.n1125 VSS.n1124 0.00476
R29816 VSS.n1126 VSS.n1125 0.00476
R29817 VSS.n1126 VSS.n81 0.00476
R29818 VSS.n1132 VSS.n81 0.00476
R29819 VSS.n1134 VSS.n1133 0.00476
R29820 VSS.n1134 VSS.n57 0.00476
R29821 VSS.n574 VSS.n573 0.00476
R29822 VSS.n522 VSS.n391 0.00476
R29823 VSS.n518 VSS.n391 0.00476
R29824 VSS.n518 VSS.n517 0.00476
R29825 VSS.n517 VSS.n516 0.00476
R29826 VSS.n516 VSS.n397 0.00476
R29827 VSS.n512 VSS.n397 0.00476
R29828 VSS.n512 VSS.n511 0.00476
R29829 VSS.n511 VSS.n510 0.00476
R29830 VSS.n510 VSS.n403 0.00476
R29831 VSS.n506 VSS.n403 0.00476
R29832 VSS.n506 VSS.n505 0.00476
R29833 VSS.n505 VSS.n504 0.00476
R29834 VSS.n504 VSS.n409 0.00476
R29835 VSS.n500 VSS.n409 0.00476
R29836 VSS.n500 VSS.n499 0.00476
R29837 VSS.n499 VSS.n498 0.00476
R29838 VSS.n495 VSS.n494 0.00476
R29839 VSS.n494 VSS.n493 0.00476
R29840 VSS.n493 VSS.n419 0.00476
R29841 VSS.n488 VSS.n487 0.00476
R29842 VSS.n487 VSS.n486 0.00476
R29843 VSS.n486 VSS.n426 0.00476
R29844 VSS.n482 VSS.n426 0.00476
R29845 VSS.n482 VSS.n481 0.00476
R29846 VSS.n481 VSS.n480 0.00476
R29847 VSS.n480 VSS.n432 0.00476
R29848 VSS.n476 VSS.n432 0.00476
R29849 VSS.n476 VSS.n475 0.00476
R29850 VSS.n475 VSS.n474 0.00476
R29851 VSS.n474 VSS.n438 0.00476
R29852 VSS.n470 VSS.n469 0.00476
R29853 VSS.n469 VSS.n468 0.00476
R29854 VSS.n468 VSS.n444 0.00476
R29855 VSS.n464 VSS.n444 0.00476
R29856 VSS.n464 VSS.n463 0.00476
R29857 VSS.n463 VSS.n462 0.00476
R29858 VSS.n462 VSS.n450 0.00476
R29859 VSS.n458 VSS.n450 0.00476
R29860 VSS.n458 VSS.n457 0.00476
R29861 VSS.n457 VSS.n132 0.00476
R29862 VSS.n954 VSS.n132 0.00476
R29863 VSS.n961 VSS.n126 0.00476
R29864 VSS.n962 VSS.n961 0.00476
R29865 VSS.n964 VSS.n962 0.00476
R29866 VSS.n964 VSS.n963 0.00476
R29867 VSS.n971 VSS.n970 0.00476
R29868 VSS.n972 VSS.n971 0.00476
R29869 VSS.n972 VSS.n118 0.00476
R29870 VSS.n978 VSS.n118 0.00476
R29871 VSS.n979 VSS.n978 0.00476
R29872 VSS.n980 VSS.n979 0.00476
R29873 VSS.n980 VSS.n114 0.00476
R29874 VSS.n986 VSS.n114 0.00476
R29875 VSS.n987 VSS.n986 0.00476
R29876 VSS.n988 VSS.n987 0.00476
R29877 VSS.n988 VSS.n110 0.00476
R29878 VSS.n994 VSS.n110 0.00476
R29879 VSS.n995 VSS.n994 0.00476
R29880 VSS.n996 VSS.n995 0.00476
R29881 VSS.n996 VSS.n106 0.00476
R29882 VSS.n1002 VSS.n103 0.00476
R29883 VSS.n1051 VSS.n1050 0.00476
R29884 VSS.n1050 VSS.n1049 0.00476
R29885 VSS.n1049 VSS.n1012 0.00476
R29886 VSS.n1045 VSS.n1012 0.00476
R29887 VSS.n1045 VSS.n1044 0.00476
R29888 VSS.n1044 VSS.n1043 0.00476
R29889 VSS.n1043 VSS.n1017 0.00476
R29890 VSS.n1039 VSS.n1017 0.00476
R29891 VSS.n1039 VSS.n1038 0.00476
R29892 VSS.n1038 VSS.n1037 0.00476
R29893 VSS.n1034 VSS.n1033 0.00476
R29894 VSS.n1033 VSS.n1032 0.00476
R29895 VSS.n1032 VSS.n36 0.00476
R29896 VSS.n3736 VSS.n2815 0.00476
R29897 VSS.n3737 VSS.n3736 0.00476
R29898 VSS.n3738 VSS.n3737 0.00476
R29899 VSS.n3738 VSS.n2811 0.00476
R29900 VSS.n3744 VSS.n2811 0.00476
R29901 VSS.n3747 VSS.n3746 0.00476
R29902 VSS.n3747 VSS.n2807 0.00476
R29903 VSS.n3753 VSS.n2807 0.00476
R29904 VSS.n3754 VSS.n3753 0.00476
R29905 VSS.n3755 VSS.n3754 0.00476
R29906 VSS.n3755 VSS.n2802 0.00476
R29907 VSS.n3864 VSS.n2803 0.00476
R29908 VSS.n3860 VSS.n2803 0.00476
R29909 VSS.n3860 VSS.n3859 0.00476
R29910 VSS.n3859 VSS.n3858 0.00476
R29911 VSS.n3858 VSS.n3763 0.00476
R29912 VSS.n3854 VSS.n3763 0.00476
R29913 VSS.n3854 VSS.n3853 0.00476
R29914 VSS.n3853 VSS.n3852 0.00476
R29915 VSS.n3852 VSS.n3769 0.00476
R29916 VSS.n3848 VSS.n3847 0.00476
R29917 VSS.n3847 VSS.n3846 0.00476
R29918 VSS.n3846 VSS.n3776 0.00476
R29919 VSS.n3842 VSS.n3776 0.00476
R29920 VSS.n3842 VSS.n3841 0.00476
R29921 VSS.n3841 VSS.n3840 0.00476
R29922 VSS.n3840 VSS.n3782 0.00476
R29923 VSS.n3836 VSS.n3782 0.00476
R29924 VSS.n3836 VSS.n3835 0.00476
R29925 VSS.n3835 VSS.n3834 0.00476
R29926 VSS.n3834 VSS.n3788 0.00476
R29927 VSS.n3830 VSS.n3788 0.00476
R29928 VSS.n3830 VSS.n3829 0.00476
R29929 VSS.n3829 VSS.n3828 0.00476
R29930 VSS.n3828 VSS.n3794 0.00476
R29931 VSS.n3824 VSS.n3794 0.00476
R29932 VSS.n3824 VSS.n3823 0.00476
R29933 VSS.n3823 VSS.n3822 0.00476
R29934 VSS.n3822 VSS.n3800 0.00476
R29935 VSS.n3818 VSS.n3800 0.00476
R29936 VSS.n3818 VSS.n3817 0.00476
R29937 VSS.n3817 VSS.n3816 0.00476
R29938 VSS.n3816 VSS.n3806 0.00476
R29939 VSS.n3812 VSS.n3806 0.00476
R29940 VSS.n3812 VSS.n2114 0.00476
R29941 VSS.n5387 VSS.n2115 0.00476
R29942 VSS.n5383 VSS.n2115 0.00476
R29943 VSS.n5383 VSS.n5382 0.00476
R29944 VSS.n5382 VSS.n5381 0.00476
R29945 VSS.n5381 VSS.n2121 0.00476
R29946 VSS.n5377 VSS.n2121 0.00476
R29947 VSS.n5375 VSS.n5374 0.00476
R29948 VSS.n5374 VSS.n2128 0.00476
R29949 VSS.n5370 VSS.n2128 0.00476
R29950 VSS.n5370 VSS.n5369 0.00476
R29951 VSS.n5369 VSS.n5368 0.00476
R29952 VSS.n5365 VSS.n5364 0.00476
R29953 VSS.n5364 VSS.n5363 0.00476
R29954 VSS.n5363 VSS.n2139 0.00476
R29955 VSS.n5359 VSS.n2139 0.00476
R29956 VSS.n5359 VSS.n5358 0.00476
R29957 VSS.n5358 VSS.n5357 0.00476
R29958 VSS.n5357 VSS.n2145 0.00476
R29959 VSS.n5353 VSS.n2145 0.00476
R29960 VSS.n5353 VSS.n5352 0.00476
R29961 VSS.n5352 VSS.n5351 0.00476
R29962 VSS.n5351 VSS.n2151 0.00476
R29963 VSS.n5347 VSS.n2151 0.00476
R29964 VSS.n5347 VSS.n5346 0.00476
R29965 VSS.n5346 VSS.n5345 0.00476
R29966 VSS.n5345 VSS.n2157 0.00476
R29967 VSS.n2171 VSS.n2164 0.00476
R29968 VSS.n3543 VSS.n2881 0.00465761
R29969 VSS.n3542 VSS.n2878 0.00465761
R29970 VSS.n3307 VSS.n3077 0.00461429
R29971 VSS.n3303 VSS.n3081 0.00461429
R29972 VSS.n3082 VSS.n3076 0.00461429
R29973 VSS.n913 VSS.n217 0.00461371
R29974 VSS.n1087 DVSS 0.00458
R29975 VSS.n1088 DVSS 0.00458
R29976 VSS.n632 VSS.n631 0.0045724
R29977 VSS.n764 VSS.n321 0.0045
R29978 VSS.n957 VSS.n128 0.0045
R29979 VSS.n386 VSS.n385 0.0045
R29980 VSS.n764 VSS.n322 0.0045
R29981 VSS.n853 VSS.n128 0.0045
R29982 VSS.n1055 VSS.n1054 0.0045
R29983 VSS.n1056 VSS.n1055 0.0045
R29984 VSS.n387 VSS.n386 0.0045
R29985 VSS.n4302 VSS.n4299 0.0045
R29986 VSS.n5073 VSS.n4354 0.0045
R29987 VSS.n4572 VSS.n4569 0.0045
R29988 VSS.n4882 VSS.n4879 0.0045
R29989 VSS.n4650 VSS.n4648 0.0045
R29990 VSS.n4684 VSS.n4683 0.0045
R29991 VSS.n4842 VSS.n4840 0.0045
R29992 VSS.n4876 VSS.n4875 0.0045
R29993 VSS.n3007 VSS.n2979 0.00448571
R29994 VSS.n3003 VSS.n3002 0.00448571
R29995 VSS.n2977 VSS.n2923 0.00448571
R29996 VSS.n4221 VSS.n4220 0.00442143
R29997 VSS.n633 VSS.n365 0.0044172
R29998 VSS.n382 VSS.n381 0.00434
R29999 VSS.n581 VSS.n580 0.00434
R30000 VSS.n577 VSS.n375 0.00434
R30001 VSS.n3358 VSS.n2909 0.004325
R30002 VSS.n2994 VSS.n2984 0.004325
R30003 VSS.n4203 VSS.n4201 0.00429286
R30004 VSS.n1878 VSS.n1877 0.00428827
R30005 VSS.n1915 VSS.n1746 0.00428827
R30006 VSS.n1953 VSS.n1704 0.00428827
R30007 VSS.n1740 VSS.n1739 0.00428827
R30008 VSS.n1734 VSS.n1733 0.00428827
R30009 VSS.n2043 VSS.n2042 0.00428827
R30010 VSS.n750 VSS.n749 0.00425
R30011 VSS.n752 VSS.n325 0.00425
R30012 VSS.n495 VSS.n330 0.00425
R30013 VSS.n1139 VSS.n1138 0.00422
R30014 VSS.n1142 VSS.n37 0.00422
R30015 VSS.n5388 VSS.n2114 0.00419
R30016 VSS.n2172 VSS.n2163 0.00419
R30017 VSS.n3046 VSS.n2831 0.0041856
R30018 VSS.n3035 VSS.n2837 0.0041856
R30019 VSS.n1766 VSS.n1762 0.00416429
R30020 VSS.n1882 VSS.n1767 0.00416429
R30021 VSS.n1881 VSS.n1768 0.00416429
R30022 VSS.n1777 VSS.n1776 0.00416429
R30023 VSS.n1873 VSS.n1872 0.00416429
R30024 VSS.n1784 VSS.n1778 0.00416429
R30025 VSS.n1866 VSS.n1787 0.00416429
R30026 VSS.n2062 VSS.n1603 0.0041
R30027 VSS.n2061 VSS.n1597 0.0041
R30028 VSS.n3745 VSS.n3744 0.00407
R30029 VSS.n3865 VSS.n3864 0.00407
R30030 VSS.n1052 VSS.n98 0.00404
R30031 VSS.n1105 VSS.n92 0.00404
R30032 VSS.n1104 VSS.n1103 0.00404
R30033 VSS.n1102 VSS.n94 0.00404
R30034 VSS.n1109 VSS.n1108 0.00404
R30035 VSS.n1051 VSS.n93 0.00404
R30036 VSS.n3724 VSS.n2818 0.00403571
R30037 VSS.n4390 VSS.n4389 0.004
R30038 VSS.n4944 VSS.n4943 0.004
R30039 VSS.n4709 VSS.n4640 0.004
R30040 VSS.n4819 VSS.n4540 0.004
R30041 VSS.n866 VSS.n283 0.00395
R30042 VSS.n942 VSS.n141 0.00395
R30043 VSS.n970 VSS.n122 0.00395
R30044 VSS.n5376 VSS.n5375 0.00395
R30045 VSS.n5340 VSS.n2163 0.00395
R30046 VSS.n3350 VSS.n2915 0.00393049
R30047 VSS.n3353 VSS.n3352 0.00393049
R30048 VSS.n3140 VSS.n3094 0.00393049
R30049 VSS.n3138 VSS.n3137 0.00393049
R30050 VSS.n5343 DVSS 0.00392
R30051 VSS.n1036 DVSS 0.00392
R30052 VSS.n1037 DVSS 0.00392
R30053 DVSS VSS.n2157 0.00392
R30054 VSS.n912 VSS.n911 0.00391137
R30055 VSS.n902 VSS.n262 0.00386658
R30056 VSS.n1877 VSS.n1876 0.00382908
R30057 VSS.n1899 VSS.n1746 0.00382908
R30058 VSS.n1937 VSS.n1704 0.00382908
R30059 VSS.n1740 VSS.n1687 0.00382908
R30060 VSS.n1734 VSS.n1662 0.00382908
R30061 VSS.n2042 VSS.n2041 0.00382908
R30062 VSS.n131 VSS.n127 0.0038
R30063 VSS.n950 VSS.n136 0.0038
R30064 VSS.n291 VSS.n288 0.0038
R30065 VSS.n287 VSS.n133 0.0038
R30066 VSS.n952 VSS.n951 0.0038
R30067 VSS.n953 VSS.n126 0.0038
R30068 VSS.n3848 VSS.n3775 0.0038
R30069 VSS.n4108 VSS.n4107 0.00377857
R30070 VSS.n4118 VSS.n4117 0.00377857
R30071 VSS.n4139 VSS.n4138 0.00377857
R30072 VSS.n635 VSS.n634 0.00374841
R30073 VSS.n3511 VSS.n3392 0.00362245
R30074 VSS.n4630 VSS.n4537 0.00360345
R30075 VSS.n4821 VSS.n4820 0.00360345
R30076 VSS.n901 VSS.n263 0.00359
R30077 VSS.n916 VSS.n164 0.00359
R30078 VSS.n1003 VSS.n106 0.00359
R30079 VSS.n2053 VSS.n1618 0.00358571
R30080 VSS.n1623 VSS.n1622 0.00358571
R30081 VSS.n2047 VSS.n2046 0.00358571
R30082 VSS.n1632 VSS.n1624 0.00358571
R30083 VSS.n2038 VSS.n1633 0.00358571
R30084 VSS.n2037 VSS.n1634 0.00358571
R30085 VSS.n1643 VSS.n1640 0.00358571
R30086 VSS.n490 VSS.n489 0.00356
R30087 VSS.n766 VSS.n320 0.00356
R30088 VSS.n741 VSS.n713 0.00356
R30089 VSS.n743 VSS.n742 0.00356
R30090 VSS.n767 VSS.n319 0.00356
R30091 VSS.n488 VSS.n425 0.00356
R30092 VSS.n669 VSS.n353 0.0035543
R30093 DVSS VSS.n80 0.00353
R30094 VSS.n1133 DVSS 0.00353
R30095 VSS.n5032 VSS.n4411 0.0035
R30096 VSS.n4517 VSS.n4516 0.0035
R30097 VSS.n4730 VSS.n4413 0.0035
R30098 VSS.n4800 VSS.n4799 0.0035
R30099 VSS.n1005 VSS.n1004 0.00341771
R30100 VSS.n3290 VSS.n3092 0.00338991
R30101 VSS.n1079 VSS.n1075 0.00338166
R30102 VSS.n2167 VSS.n2164 0.00338166
R30103 VSS.n3734 VSS.n2813 0.00334
R30104 VSS.n3740 VSS.n2813 0.00334
R30105 VSS.n3741 VSS.n3740 0.00334
R30106 VSS.n3742 VSS.n3741 0.00334
R30107 VSS.n3742 VSS.n2809 0.00334
R30108 VSS.n3749 VSS.n2809 0.00334
R30109 VSS.n3750 VSS.n3749 0.00334
R30110 VSS.n3751 VSS.n3750 0.00334
R30111 VSS.n3751 VSS.n2805 0.00334
R30112 VSS.n3757 VSS.n2805 0.00334
R30113 VSS.n3758 VSS.n3757 0.00334
R30114 VSS.n3759 VSS.n3758 0.00334
R30115 VSS.n3760 VSS.n3759 0.00334
R30116 VSS.n3761 VSS.n3760 0.00334
R30117 VSS.n3764 VSS.n3761 0.00334
R30118 VSS.n3765 VSS.n3764 0.00334
R30119 VSS.n3766 VSS.n3765 0.00334
R30120 VSS.n3767 VSS.n3766 0.00334
R30121 VSS.n3770 VSS.n3767 0.00334
R30122 VSS.n3771 VSS.n3770 0.00334
R30123 VSS.n3772 VSS.n3771 0.00334
R30124 VSS.n3773 VSS.n3772 0.00334
R30125 VSS.n3777 VSS.n3773 0.00334
R30126 VSS.n3778 VSS.n3777 0.00334
R30127 VSS.n3779 VSS.n3778 0.00334
R30128 VSS.n3780 VSS.n3779 0.00334
R30129 VSS.n3783 VSS.n3780 0.00334
R30130 VSS.n3784 VSS.n3783 0.00334
R30131 VSS.n3785 VSS.n3784 0.00334
R30132 VSS.n3786 VSS.n3785 0.00334
R30133 VSS.n3789 VSS.n3786 0.00334
R30134 VSS.n3790 VSS.n3789 0.00334
R30135 VSS.n3791 VSS.n3790 0.00334
R30136 VSS.n3792 VSS.n3791 0.00334
R30137 VSS.n3795 VSS.n3792 0.00334
R30138 VSS.n3796 VSS.n3795 0.00334
R30139 VSS.n3797 VSS.n3796 0.00334
R30140 VSS.n3798 VSS.n3797 0.00334
R30141 VSS.n3801 VSS.n3798 0.00334
R30142 VSS.n3802 VSS.n3801 0.00334
R30143 VSS.n3803 VSS.n3802 0.00334
R30144 VSS.n3804 VSS.n3803 0.00334
R30145 VSS.n3807 VSS.n3804 0.00334
R30146 VSS.n3808 VSS.n3807 0.00334
R30147 VSS.n3809 VSS.n3808 0.00334
R30148 VSS.n3811 VSS.n3809 0.00334
R30149 VSS.n3811 VSS.n3810 0.00334
R30150 VSS.n3810 VSS.n2117 0.00334
R30151 VSS.n2118 VSS.n2117 0.00334
R30152 VSS.n2119 VSS.n2118 0.00334
R30153 VSS.n2122 VSS.n2119 0.00334
R30154 VSS.n2123 VSS.n2122 0.00334
R30155 VSS.n2124 VSS.n2123 0.00334
R30156 VSS.n2125 VSS.n2124 0.00334
R30157 VSS.n2129 VSS.n2125 0.00334
R30158 VSS.n2130 VSS.n2129 0.00334
R30159 VSS.n2131 VSS.n2130 0.00334
R30160 VSS.n2132 VSS.n2131 0.00334
R30161 VSS.n2135 VSS.n2132 0.00334
R30162 VSS.n2136 VSS.n2135 0.00334
R30163 VSS.n2137 VSS.n2136 0.00334
R30164 VSS.n2140 VSS.n2137 0.00334
R30165 VSS.n2141 VSS.n2140 0.00334
R30166 VSS.n2142 VSS.n2141 0.00334
R30167 VSS.n2143 VSS.n2142 0.00334
R30168 VSS.n2146 VSS.n2143 0.00334
R30169 VSS.n2147 VSS.n2146 0.00334
R30170 VSS.n2148 VSS.n2147 0.00334
R30171 VSS.n2149 VSS.n2148 0.00334
R30172 VSS.n2152 VSS.n2149 0.00334
R30173 VSS.n2153 VSS.n2152 0.00334
R30174 VSS.n2154 VSS.n2153 0.00334
R30175 VSS.n2155 VSS.n2154 0.00334
R30176 VSS.n2158 VSS.n2155 0.00334
R30177 VSS.n2159 VSS.n2158 0.00334
R30178 VSS.n2160 VSS.n2159 0.00334
R30179 VSS.n2166 VSS.n2165 0.00334
R30180 VSS.n384 VSS.n350 0.00334
R30181 VSS.n673 VSS.n350 0.00334
R30182 VSS.n674 VSS.n673 0.00334
R30183 VSS.n675 VSS.n674 0.00334
R30184 VSS.n675 VSS.n346 0.00334
R30185 VSS.n681 VSS.n346 0.00334
R30186 VSS.n682 VSS.n681 0.00334
R30187 VSS.n683 VSS.n682 0.00334
R30188 VSS.n683 VSS.n342 0.00334
R30189 VSS.n689 VSS.n342 0.00334
R30190 VSS.n690 VSS.n689 0.00334
R30191 VSS.n691 VSS.n690 0.00334
R30192 VSS.n691 VSS.n338 0.00334
R30193 VSS.n697 VSS.n338 0.00334
R30194 VSS.n698 VSS.n697 0.00334
R30195 VSS.n699 VSS.n698 0.00334
R30196 VSS.n699 VSS.n334 0.00334
R30197 VSS.n705 VSS.n334 0.00334
R30198 VSS.n706 VSS.n705 0.00334
R30199 VSS.n707 VSS.n706 0.00334
R30200 VSS.n708 VSS.n707 0.00334
R30201 VSS.n709 VSS.n708 0.00334
R30202 VSS.n710 VSS.n709 0.00334
R30203 VSS.n715 VSS.n714 0.00334
R30204 VSS.n716 VSS.n715 0.00334
R30205 VSS.n719 VSS.n716 0.00334
R30206 VSS.n720 VSS.n719 0.00334
R30207 VSS.n721 VSS.n720 0.00334
R30208 VSS.n722 VSS.n721 0.00334
R30209 VSS.n725 VSS.n722 0.00334
R30210 VSS.n726 VSS.n725 0.00334
R30211 VSS.n727 VSS.n726 0.00334
R30212 VSS.n727 VSS.n302 0.00334
R30213 VSS.n828 VSS.n302 0.00334
R30214 VSS.n829 VSS.n828 0.00334
R30215 VSS.n830 VSS.n829 0.00334
R30216 VSS.n830 VSS.n298 0.00334
R30217 VSS.n836 VSS.n298 0.00334
R30218 VSS.n837 VSS.n836 0.00334
R30219 VSS.n838 VSS.n837 0.00334
R30220 VSS.n838 VSS.n294 0.00334
R30221 VSS.n844 VSS.n294 0.00334
R30222 VSS.n845 VSS.n844 0.00334
R30223 VSS.n846 VSS.n845 0.00334
R30224 VSS.n846 VSS.n289 0.00334
R30225 VSS.n852 VSS.n289 0.00334
R30226 VSS.n855 VSS.n854 0.00334
R30227 VSS.n855 VSS.n285 0.00334
R30228 VSS.n862 VSS.n285 0.00334
R30229 VSS.n863 VSS.n862 0.00334
R30230 VSS.n864 VSS.n863 0.00334
R30231 VSS.n864 VSS.n280 0.00334
R30232 VSS.n870 VSS.n280 0.00334
R30233 VSS.n871 VSS.n870 0.00334
R30234 VSS.n872 VSS.n871 0.00334
R30235 VSS.n872 VSS.n276 0.00334
R30236 VSS.n878 VSS.n276 0.00334
R30237 VSS.n879 VSS.n878 0.00334
R30238 VSS.n880 VSS.n879 0.00334
R30239 VSS.n880 VSS.n272 0.00334
R30240 VSS.n886 VSS.n272 0.00334
R30241 VSS.n887 VSS.n886 0.00334
R30242 VSS.n888 VSS.n887 0.00334
R30243 VSS.n888 VSS.n268 0.00334
R30244 VSS.n894 VSS.n268 0.00334
R30245 VSS.n895 VSS.n894 0.00334
R30246 VSS.n896 VSS.n895 0.00334
R30247 VSS.n897 VSS.n896 0.00334
R30248 VSS.n897 VSS.n100 0.00334
R30249 VSS.n1060 VSS.n1057 0.00334
R30250 VSS.n1061 VSS.n1060 0.00334
R30251 VSS.n1062 VSS.n1061 0.00334
R30252 VSS.n1063 VSS.n1062 0.00334
R30253 VSS.n1066 VSS.n1063 0.00334
R30254 VSS.n1067 VSS.n1066 0.00334
R30255 VSS.n1068 VSS.n1067 0.00334
R30256 VSS.n1069 VSS.n1068 0.00334
R30257 VSS.n1071 VSS.n1069 0.00334
R30258 VSS.n1072 VSS.n1071 0.00334
R30259 VSS.n1073 VSS.n1072 0.00334
R30260 VSS.n1077 VSS.n1076 0.00334
R30261 VSS.n584 VSS.n370 0.00334
R30262 VSS.n585 VSS.n584 0.00334
R30263 VSS.n586 VSS.n585 0.00334
R30264 VSS.n587 VSS.n586 0.00334
R30265 VSS.n588 VSS.n587 0.00334
R30266 VSS.n591 VSS.n588 0.00334
R30267 VSS.n592 VSS.n591 0.00334
R30268 VSS.n593 VSS.n592 0.00334
R30269 VSS.n594 VSS.n593 0.00334
R30270 VSS.n597 VSS.n594 0.00334
R30271 VSS.n598 VSS.n597 0.00334
R30272 VSS.n599 VSS.n598 0.00334
R30273 VSS.n600 VSS.n599 0.00334
R30274 VSS.n603 VSS.n600 0.00334
R30275 VSS.n604 VSS.n603 0.00334
R30276 VSS.n605 VSS.n604 0.00334
R30277 VSS.n606 VSS.n605 0.00334
R30278 VSS.n606 VSS.n327 0.00334
R30279 VSS.n755 VSS.n327 0.00334
R30280 VSS.n756 VSS.n755 0.00334
R30281 VSS.n757 VSS.n756 0.00334
R30282 VSS.n757 VSS.n323 0.00334
R30283 VSS.n763 VSS.n323 0.00334
R30284 VSS.n765 VSS.n317 0.00334
R30285 VSS.n771 VSS.n317 0.00334
R30286 VSS.n772 VSS.n771 0.00334
R30287 VSS.n773 VSS.n772 0.00334
R30288 VSS.n773 VSS.n313 0.00334
R30289 VSS.n779 VSS.n313 0.00334
R30290 VSS.n780 VSS.n779 0.00334
R30291 VSS.n781 VSS.n780 0.00334
R30292 VSS.n781 VSS.n309 0.00334
R30293 VSS.n787 VSS.n309 0.00334
R30294 VSS.n788 VSS.n787 0.00334
R30295 VSS.n789 VSS.n788 0.00334
R30296 VSS.n790 VSS.n789 0.00334
R30297 VSS.n791 VSS.n790 0.00334
R30298 VSS.n794 VSS.n791 0.00334
R30299 VSS.n795 VSS.n794 0.00334
R30300 VSS.n796 VSS.n795 0.00334
R30301 VSS.n797 VSS.n796 0.00334
R30302 VSS.n800 VSS.n797 0.00334
R30303 VSS.n801 VSS.n800 0.00334
R30304 VSS.n802 VSS.n801 0.00334
R30305 VSS.n803 VSS.n802 0.00334
R30306 VSS.n804 VSS.n803 0.00334
R30307 VSS.n138 VSS.n137 0.00334
R30308 VSS.n139 VSS.n138 0.00334
R30309 VSS.n142 VSS.n139 0.00334
R30310 VSS.n143 VSS.n142 0.00334
R30311 VSS.n144 VSS.n143 0.00334
R30312 VSS.n147 VSS.n144 0.00334
R30313 VSS.n148 VSS.n147 0.00334
R30314 VSS.n149 VSS.n148 0.00334
R30315 VSS.n150 VSS.n149 0.00334
R30316 VSS.n153 VSS.n150 0.00334
R30317 VSS.n154 VSS.n153 0.00334
R30318 VSS.n155 VSS.n154 0.00334
R30319 VSS.n156 VSS.n155 0.00334
R30320 VSS.n159 VSS.n156 0.00334
R30321 VSS.n160 VSS.n159 0.00334
R30322 VSS.n161 VSS.n160 0.00334
R30323 VSS.n162 VSS.n161 0.00334
R30324 VSS.n165 VSS.n162 0.00334
R30325 VSS.n166 VSS.n165 0.00334
R30326 VSS.n167 VSS.n166 0.00334
R30327 VSS.n169 VSS.n167 0.00334
R30328 VSS.n169 VSS.n168 0.00334
R30329 VSS.n168 VSS.n97 0.00334
R30330 VSS.n1112 VSS.n91 0.00334
R30331 VSS.n1113 VSS.n1112 0.00334
R30332 VSS.n1114 VSS.n1113 0.00334
R30333 VSS.n1114 VSS.n87 0.00334
R30334 VSS.n1120 VSS.n87 0.00334
R30335 VSS.n1121 VSS.n1120 0.00334
R30336 VSS.n1122 VSS.n1121 0.00334
R30337 VSS.n1122 VSS.n83 0.00334
R30338 VSS.n1128 VSS.n83 0.00334
R30339 VSS.n1129 VSS.n1128 0.00334
R30340 VSS.n1130 VSS.n1129 0.00334
R30341 VSS.n1136 VSS.n79 0.00334
R30342 VSS.n389 VSS.n388 0.00334
R30343 VSS.n392 VSS.n389 0.00334
R30344 VSS.n393 VSS.n392 0.00334
R30345 VSS.n394 VSS.n393 0.00334
R30346 VSS.n395 VSS.n394 0.00334
R30347 VSS.n398 VSS.n395 0.00334
R30348 VSS.n399 VSS.n398 0.00334
R30349 VSS.n400 VSS.n399 0.00334
R30350 VSS.n401 VSS.n400 0.00334
R30351 VSS.n404 VSS.n401 0.00334
R30352 VSS.n405 VSS.n404 0.00334
R30353 VSS.n406 VSS.n405 0.00334
R30354 VSS.n407 VSS.n406 0.00334
R30355 VSS.n410 VSS.n407 0.00334
R30356 VSS.n411 VSS.n410 0.00334
R30357 VSS.n412 VSS.n411 0.00334
R30358 VSS.n413 VSS.n412 0.00334
R30359 VSS.n415 VSS.n413 0.00334
R30360 VSS.n416 VSS.n415 0.00334
R30361 VSS.n417 VSS.n416 0.00334
R30362 VSS.n420 VSS.n417 0.00334
R30363 VSS.n421 VSS.n420 0.00334
R30364 VSS.n422 VSS.n421 0.00334
R30365 VSS.n427 VSS.n423 0.00334
R30366 VSS.n428 VSS.n427 0.00334
R30367 VSS.n429 VSS.n428 0.00334
R30368 VSS.n430 VSS.n429 0.00334
R30369 VSS.n433 VSS.n430 0.00334
R30370 VSS.n434 VSS.n433 0.00334
R30371 VSS.n435 VSS.n434 0.00334
R30372 VSS.n436 VSS.n435 0.00334
R30373 VSS.n439 VSS.n436 0.00334
R30374 VSS.n440 VSS.n439 0.00334
R30375 VSS.n441 VSS.n440 0.00334
R30376 VSS.n442 VSS.n441 0.00334
R30377 VSS.n445 VSS.n442 0.00334
R30378 VSS.n446 VSS.n445 0.00334
R30379 VSS.n447 VSS.n446 0.00334
R30380 VSS.n448 VSS.n447 0.00334
R30381 VSS.n451 VSS.n448 0.00334
R30382 VSS.n452 VSS.n451 0.00334
R30383 VSS.n453 VSS.n452 0.00334
R30384 VSS.n454 VSS.n453 0.00334
R30385 VSS.n455 VSS.n454 0.00334
R30386 VSS.n455 VSS.n129 0.00334
R30387 VSS.n956 VSS.n129 0.00334
R30388 VSS.n959 VSS.n958 0.00334
R30389 VSS.n959 VSS.n124 0.00334
R30390 VSS.n966 VSS.n124 0.00334
R30391 VSS.n967 VSS.n966 0.00334
R30392 VSS.n968 VSS.n967 0.00334
R30393 VSS.n968 VSS.n120 0.00334
R30394 VSS.n974 VSS.n120 0.00334
R30395 VSS.n975 VSS.n974 0.00334
R30396 VSS.n976 VSS.n975 0.00334
R30397 VSS.n976 VSS.n116 0.00334
R30398 VSS.n982 VSS.n116 0.00334
R30399 VSS.n983 VSS.n982 0.00334
R30400 VSS.n984 VSS.n983 0.00334
R30401 VSS.n984 VSS.n112 0.00334
R30402 VSS.n990 VSS.n112 0.00334
R30403 VSS.n991 VSS.n990 0.00334
R30404 VSS.n992 VSS.n991 0.00334
R30405 VSS.n992 VSS.n108 0.00334
R30406 VSS.n998 VSS.n108 0.00334
R30407 VSS.n999 VSS.n998 0.00334
R30408 VSS.n1000 VSS.n999 0.00334
R30409 VSS.n1000 VSS.n101 0.00334
R30410 VSS.n1009 VSS.n101 0.00334
R30411 VSS.n1053 VSS.n1010 0.00334
R30412 VSS.n1013 VSS.n1010 0.00334
R30413 VSS.n1014 VSS.n1013 0.00334
R30414 VSS.n1015 VSS.n1014 0.00334
R30415 VSS.n1018 VSS.n1015 0.00334
R30416 VSS.n1019 VSS.n1018 0.00334
R30417 VSS.n1020 VSS.n1019 0.00334
R30418 VSS.n1021 VSS.n1020 0.00334
R30419 VSS.n1023 VSS.n1021 0.00334
R30420 VSS.n1024 VSS.n1023 0.00334
R30421 VSS.n1025 VSS.n1024 0.00334
R30422 VSS.n1028 VSS.n1027 0.00334
R30423 VSS.n1958 VSS.n1700 0.00332857
R30424 VSS.n1957 VSS.n1701 0.00332857
R30425 VSS.n1707 VSS.n1706 0.00332857
R30426 VSS.n1950 VSS.n1949 0.00332857
R30427 VSS.n1714 VSS.n1708 0.00332857
R30428 VSS.n1943 VSS.n1715 0.00332857
R30429 VSS.n1942 VSS.n1935 0.00332857
R30430 VSS.n3952 VSS.n3951 0.00332857
R30431 VSS.n576 VSS.n376 0.00332
R30432 VSS.n378 VSS.n371 0.00332
R30433 VSS.n383 VSS.n379 0.00332
R30434 VSS.n382 VSS.n372 0.00332
R30435 VSS.n580 VSS.n579 0.00332
R30436 VSS.n578 VSS.n577 0.00332
R30437 VSS.n1150 VSS.n29 0.00330488
R30438 VSS.n1165 VSS.n24 0.00330488
R30439 VSS.n826 VSS.n825 0.00329
R30440 VSS.n823 VSS.n306 0.00329
R30441 VSS.n438 VSS.n305 0.00329
R30442 VSS.n2165 DVSS 0.00326
R30443 VSS.n1027 DVSS 0.00326
R30444 VSS.n3728 VSS.n3727 0.0032
R30445 VSS.n4250 VSS.n2352 0.0032
R30446 VSS.n915 VSS.n170 0.00319327
R30447 VSS.n2886 VSS.n2876 0.00319022
R30448 VSS.n3534 VSS.n2883 0.00319022
R30449 VSS.n3505 VSS 0.00314706
R30450 VSS VSS.n3397 0.00314706
R30451 VSS.n571 VSS.n523 0.00314706
R30452 VSS.n4231 VSS.n4230 0.00313571
R30453 VSS.n2392 VSS.n2388 0.00313571
R30454 VSS.n671 VSS.n670 0.00311
R30455 VSS.n630 VSS.n367 0.00311
R30456 VSS.n573 VSS.n572 0.00311
R30457 VSS.n2169 VSS.n2168 0.00309529
R30458 VSS.n1030 VSS.n1029 0.00309529
R30459 VSS.n1137 VSS.n78 0.00309529
R30460 VSS.n1081 VSS.n1080 0.00309529
R30461 VSS.n2407 VSS.n2403 0.00307143
R30462 VSS.n4187 VSS.n2408 0.00307143
R30463 VSS.n4186 VSS.n4171 0.00307143
R30464 VSS.n1831 VSS.n19 0.00300714
R30465 VSS.n1587 VSS.n1298 0.00300714
R30466 VSS.n4239 VSS.n2373 0.00300714
R30467 VSS.n5009 VSS.n4443 0.003
R30468 VSS.n4985 VSS.n4477 0.003
R30469 VSS.n4751 VSS.n4750 0.003
R30470 VSS.n4777 VSS.n4475 0.003
R30471 VSS.n3020 VSS.n3012 0.00297706
R30472 VSS.n4296 VSS.n4294 0.00296479
R30473 VSS.n5115 VSS.n4297 0.00296479
R30474 VSS.n4649 VSS.n4304 0.00296479
R30475 VSS.n5107 VSS.n5106 0.00296479
R30476 VSS.n5103 VSS.n4306 0.00296479
R30477 VSS.n5102 VSS.n4317 0.00296479
R30478 VSS.n4660 VSS.n4324 0.00296479
R30479 VSS.n5095 VSS.n5094 0.00296479
R30480 VSS.n5091 VSS.n4326 0.00296479
R30481 VSS.n5090 VSS.n4334 0.00296479
R30482 VSS.n4671 VSS.n4341 0.00296479
R30483 VSS.n5083 VSS.n5082 0.00296479
R30484 VSS.n5079 VSS.n4343 0.00296479
R30485 VSS.n5078 VSS.n4351 0.00296479
R30486 VSS.n4690 VSS.n4685 0.00296479
R30487 VSS.n4691 VSS.n4361 0.00296479
R30488 VSS.n5067 VSS.n5066 0.00296479
R30489 VSS.n5063 VSS.n4363 0.00296479
R30490 VSS.n5062 VSS.n4369 0.00296479
R30491 VSS.n4702 VSS.n4376 0.00296479
R30492 VSS.n5055 VSS.n5054 0.00296479
R30493 VSS.n5051 VSS.n4378 0.00296479
R30494 VSS.n5050 VSS.n4386 0.00296479
R30495 VSS.n4714 VSS.n4395 0.00296479
R30496 VSS.n5043 VSS.n5042 0.00296479
R30497 VSS.n5039 VSS.n4397 0.00296479
R30498 VSS.n5038 VSS.n4405 0.00296479
R30499 VSS.n4725 VSS.n4412 0.00296479
R30500 VSS.n5031 VSS.n5030 0.00296479
R30501 VSS.n5027 VSS.n4414 0.00296479
R30502 VSS.n5026 VSS.n4422 0.00296479
R30503 VSS.n4737 VSS.n4430 0.00296479
R30504 VSS.n5019 VSS.n5018 0.00296479
R30505 VSS.n5015 VSS.n4432 0.00296479
R30506 VSS.n5014 VSS.n4440 0.00296479
R30507 VSS.n4757 VSS.n4752 0.00296479
R30508 VSS.n4758 VSS.n4451 0.00296479
R30509 VSS.n5003 VSS.n5002 0.00296479
R30510 VSS.n4999 VSS.n4453 0.00296479
R30511 VSS.n4998 VSS.n4459 0.00296479
R30512 VSS.n4769 VSS.n4466 0.00296479
R30513 VSS.n4991 VSS.n4990 0.00296479
R30514 VSS.n4987 VSS.n4468 0.00296479
R30515 VSS.n4986 VSS.n4476 0.00296479
R30516 VSS.n4781 VSS.n4485 0.00296479
R30517 VSS.n4979 VSS.n4978 0.00296479
R30518 VSS.n4975 VSS.n4487 0.00296479
R30519 VSS.n4974 VSS.n4495 0.00296479
R30520 VSS.n4793 VSS.n4503 0.00296479
R30521 VSS.n4967 VSS.n4966 0.00296479
R30522 VSS.n4963 VSS.n4505 0.00296479
R30523 VSS.n4962 VSS.n4513 0.00296479
R30524 VSS.n4805 VSS.n4521 0.00296479
R30525 VSS.n4955 VSS.n4954 0.00296479
R30526 VSS.n4951 VSS.n4523 0.00296479
R30527 VSS.n4950 VSS.n4531 0.00296479
R30528 VSS.n4816 VSS.n4539 0.00296479
R30529 VSS.n4942 VSS.n4941 0.00296479
R30530 VSS.n4938 VSS.n4541 0.00296479
R30531 VSS.n4937 VSS.n4549 0.00296479
R30532 VSS.n4829 VSS.n4556 0.00296479
R30533 VSS.n4930 VSS.n4929 0.00296479
R30534 VSS.n4926 VSS.n4558 0.00296479
R30535 VSS.n4925 VSS.n4566 0.00296479
R30536 VSS.n4841 VSS.n4574 0.00296479
R30537 VSS.n4917 VSS.n4916 0.00296479
R30538 VSS.n4913 VSS.n4576 0.00296479
R30539 VSS.n4912 VSS.n4584 0.00296479
R30540 VSS.n4852 VSS.n4591 0.00296479
R30541 VSS.n4904 VSS.n4903 0.00296479
R30542 VSS.n4900 VSS.n4593 0.00296479
R30543 VSS.n4899 VSS.n4601 0.00296479
R30544 VSS.n4863 VSS.n4609 0.00296479
R30545 VSS.n4892 VSS.n4891 0.00296479
R30546 VSS.n4888 VSS.n4611 0.00296479
R30547 VSS.n4887 VSS.n4620 0.00296479
R30548 VSS.n4878 VSS.n4877 0.00296479
R30549 VSS.n5134 VSS.n2280 0.00296479
R30550 VSS.n5133 VSS.n2276 0.00296479
R30551 VSS.n631 VSS.n366 0.00294344
R30552 VSS.n5086 DVSS 0.00293842
R30553 DVSS VSS.n4674 0.00293842
R30554 VSS.n3269 VSS.n3268 0.00293243
R30555 VSS.n265 VSS.n264 0.0029
R30556 VSS.n1107 VSS.n95 0.0029
R30557 VSS.n1007 VSS.n1006 0.0029
R30558 VSS.n5432 DVSS 0.00286842
R30559 DVSS VSS.n5338 0.00286842
R30560 VSS.n5399 DVSS 0.00286842
R30561 VSS.n2107 DVSS 0.00286842
R30562 VSS VSS.n2786 0.00286842
R30563 VSS.n1057 VSS.n1056 0.00286
R30564 VSS.n1055 VSS.n91 0.00286
R30565 VSS.n1054 VSS.n1053 0.00286
R30566 VSS.n1076 DVSS 0.00282
R30567 VSS.n2087 DVSS 0.00279616
R30568 VSS.n2174 DVSS 0.00279616
R30569 VSS.n5397 DVSS 0.00279616
R30570 VSS.n2797 DVSS 0.00279616
R30571 DVSS VSS.n2160 0.00278
R30572 VSS.n5007 VSS.n4448 0.00271675
R30573 VSS.n4747 VSS.n4634 0.00271675
R30574 VSS.n854 VSS.n853 0.0027
R30575 VSS.n137 VSS.n128 0.0027
R30576 VSS.n958 VSS.n957 0.0027
R30577 VSS.n5368 VSS.n2134 0.00269
R30578 VSS.n1990 VSS.n1989 0.00262143
R30579 VSS.n1986 VSS.n1675 0.00262143
R30580 VSS.n1985 VSS.n1678 0.00262143
R30581 VSS.n1683 VSS.n1682 0.00262143
R30582 VSS.n1979 VSS.n1978 0.00262143
R30583 VSS.n1688 VSS.n1684 0.00262143
R30584 VSS.n1973 VSS.n1689 0.00262143
R30585 VSS.n1858 VSS.n1792 0.00262143
R30586 VSS.n1857 VSS.n1798 0.00262143
R30587 VSS.n1854 VSS.n1853 0.00262143
R30588 VSS.n1157 VSS.n30 0.00257317
R30589 VSS.n1158 VSS.n26 0.00257317
R30590 VSS.n3732 VSS.n2815 0.00257
R30591 VSS.n5365 VSS.n2134 0.00257
R30592 VSS.n3132 VSS.n3097 0.00256422
R30593 VSS.n2939 VSS.n2938 0.00256422
R30594 VSS.n2021 VSS.n1648 0.00255714
R30595 VSS.n2018 VSS.n2017 0.00255714
R30596 VSS.n1657 VSS.n1651 0.00255714
R30597 VSS.n2011 VSS.n1658 0.00255714
R30598 VSS.n2010 VSS.n1659 0.00255714
R30599 VSS.n1664 VSS.n1663 0.00255714
R30600 VSS.n2005 VSS.n2004 0.00255714
R30601 VSS.n714 VSS.n322 0.00254
R30602 VSS.n765 VSS.n764 0.00254
R30603 VSS.n423 VSS.n321 0.00254
R30604 VSS.n216 VSS.n170 0.00251995
R30605 VSS.n5008 VSS.n4447 0.0025
R30606 VSS.n4480 VSS.n4479 0.0025
R30607 VSS.n4759 VSS.n4635 0.0025
R30608 VSS.n4776 VSS.n4633 0.0025
R30609 VSS.n3324 VSS.n2958 0.00249286
R30610 VSS.n3111 VSS.n2960 0.00249286
R30611 VSS.n5156 DVSS 0.00247183
R30612 VSS.n3068 VSS.n3064 0.00242857
R30613 VSS.n3065 VSS.n2950 0.00242857
R30614 VSS.n385 VSS.n384 0.00238
R30615 VSS.n386 VSS.n370 0.00238
R30616 VSS.n388 VSS.n387 0.00238
R30617 VSS.n4102 VSS.n4093 0.00236429
R30618 VSS.n266 VSS.n265 0.00236
R30619 VSS.n917 VSS.n95 0.00236
R30620 VSS.n1006 VSS.n103 0.00236
R30621 VSS.n535 VSS.n366 0.00233258
R30622 VSS.n2696 VSS 0.0023
R30623 VSS.n3184 DVSS 0.0023
R30624 VSS.n3581 DVSS 0.0023
R30625 DVSS VSS.n1839 0.0023
R30626 VSS.n1838 DVSS 0.0023
R30627 VSS.n1397 DVSS 0.0023
R30628 VSS.n5176 DVSS 0.0023
R30629 VSS VSS.n2697 0.0023
R30630 VSS VSS.n5710 0.0023
R30631 VSS.n5709 VSS 0.0023
R30632 VSS.n4056 VSS.n2463 0.00223571
R30633 VSS.n2701 VSS.n2468 0.00223571
R30634 VSS.n2697 VSS.n2462 0.00223571
R30635 VSS.n4026 VSS.n2703 0.00223571
R30636 VSS.n4025 VSS.n0 0.00223571
R30637 VSS.n5710 VSS.n1 0.00223571
R30638 VSS.n670 VSS.n348 0.00215
R30639 VSS.n630 VSS.n629 0.00215
R30640 VSS.n572 VSS.n522 0.00215
R30641 VSS.n4426 VSS.n4425 0.002
R30642 VSS.n4968 VSS.n4502 0.002
R30643 VSS.n4732 VSS.n4731 0.002
R30644 VSS.n4798 VSS.n4504 0.002
R30645 VSS.n2250 VSS.n2244 0.00197857
R30646 VSS.n825 VSS.n300 0.00197
R30647 VSS.n823 VSS.n822 0.00197
R30648 VSS.n470 VSS.n305 0.00197
R30649 VSS.n1130 DVSS 0.00196
R30650 DVSS VSS.n32 0.00191429
R30651 DVSS VSS.n79 0.00188
R30652 VSS.n4223 VSS.n4222 0.00185
R30653 VSS.n4211 VSS.n2393 0.00185
R30654 VSS.n5691 VSS.n21 0.00184146
R30655 VSS.n1166 VSS.n27 0.00184146
R30656 VSS.n5155 DVSS 0.00181455
R30657 VSS.n5239 DVSS 0.00179393
R30658 VSS.n1131 DVSS 0.00173
R30659 DVSS VSS.n1132 0.00173
R30660 VSS.n2695 VSS 0.0017
R30661 VSS.n1837 DVSS 0.0017
R30662 VSS.n491 VSS.n490 0.0017
R30663 VSS.n762 VSS.n320 0.0017
R30664 VSS.n713 VSS.n711 0.0017
R30665 VSS.n744 VSS.n743 0.0017
R30666 VSS.n761 VSS.n319 0.0017
R30667 VSS.n425 VSS.n419 0.0017
R30668 VSS.n901 VSS.n900 0.00167
R30669 VSS.n918 VSS.n916 0.00167
R30670 VSS.n1003 VSS.n1002 0.00167
R30671 VSS.n1832 VSS.n20 0.00165714
R30672 VSS.n1828 VSS.n22 0.00165714
R30673 VSS.n3277 VSS.n3153 0.00165714
R30674 VSS.n3279 VSS.n3246 0.00165714
R30675 VSS.n3486 VSS.n3477 0.00165714
R30676 VSS.n3484 VSS.n3483 0.00165714
R30677 VSS.n3480 VSS.n3479 0.00165714
R30678 VSS.n3878 VSS.n2777 0.00165714
R30679 VSS.n3877 VSS.n2778 0.00165714
R30680 VSS.n3884 VSS.n2773 0.00165714
R30681 VSS.n3885 VSS.n2771 0.00165714
R30682 VSS.n3888 VSS.n3887 0.00165714
R30683 VSS.n2827 VSS.n2822 0.00159286
R30684 VSS.n3716 VSS.n3715 0.00159286
R30685 VSS.n3713 VSS.n2833 0.00159286
R30686 VSS.n1724 VSS.n1720 0.00159286
R30687 VSS.n1920 VSS.n1919 0.00159286
R30688 VSS.n1748 VSS.n1725 0.00159286
R30689 VSS.n1912 VSS.n1749 0.00159286
R30690 VSS.n1911 VSS.n1750 0.00159286
R30691 VSS.n1757 VSS.n1756 0.00159286
R30692 VSS.n1905 VSS.n1904 0.00159286
R30693 VSS.n4147 VSS.n2426 0.00159286
R30694 VSS.n3054 VSS.n2832 0.00157001
R30695 VSS.n3015 VSS.n2899 0.00152857
R30696 VSS.n3364 VSS.n2903 0.00152857
R30697 VSS.n5049 VSS.n4387 0.0015
R30698 VSS.n4945 VSS.n4534 0.0015
R30699 VSS.n4710 VSS.n4385 0.0015
R30700 VSS.n4818 VSS.n4817 0.0015
R30701 VSS.n955 VSS.n131 0.00146
R30702 VSS.n805 VSS.n136 0.00146
R30703 VSS.n851 VSS.n291 0.00146
R30704 VSS.n850 VSS.n133 0.00146
R30705 VSS.n952 VSS.n134 0.00146
R30706 VSS.n954 VSS.n953 0.00146
R30707 VSS.n3775 VSS.n3769 0.00146
R30708 DVSS VSS.n5342 0.00134
R30709 DVSS VSS.n1035 0.00134
R30710 VSS.n1034 DVSS 0.00134
R30711 VSS.n5341 DVSS 0.00134
R30712 VSS.n3640 VSS.n2880 0.00133571
R30713 VSS.n3549 VSS.n2885 0.00133571
R30714 VSS.n3638 VSS.n3637 0.00133571
R30715 VSS.n2402 VSS.n2398 0.00133571
R30716 VSS.n859 VSS.n283 0.00131
R30717 VSS.n945 VSS.n141 0.00131
R30718 VSS.n963 VSS.n122 0.00131
R30719 VSS.n5377 VSS.n5376 0.00131
R30720 VSS.n5341 VSS.n5340 0.00131
R30721 VSS.n710 VSS.n322 0.0013
R30722 VSS.n764 VSS.n763 0.0013
R30723 VSS.n422 VSS.n321 0.0013
R30724 VSS.n1008 VSS.n98 0.00122
R30725 VSS.n1106 VSS.n1105 0.00122
R30726 VSS.n1104 VSS.n99 0.00122
R30727 VSS.n264 VSS.n94 0.00122
R30728 VSS.n1108 VSS.n1107 0.00122
R30729 VSS.n1007 VSS.n93 0.00122
R30730 VSS.n5690 DVSS 0.00120714
R30731 VSS.n4116 VSS.n4115 0.00120714
R30732 VSS.n4131 VSS.n4130 0.00120714
R30733 VSS.n3420 VSS.n3419 0.00120714
R30734 VSS.n3502 VSS.n3501 0.00120714
R30735 VSS.n3746 VSS.n3745 0.00119
R30736 VSS.n3865 VSS.n2802 0.00119
R30737 VSS.n853 VSS.n852 0.00114
R30738 VSS.n804 VSS.n128 0.00114
R30739 VSS.n957 VSS.n956 0.00114
R30740 VSS.n5388 VSS.n5387 0.00107
R30741 VSS.n2172 VSS.n2171 0.00107
R30742 VSS.n2161 DVSS 0.00106
R30743 VSS.n1139 VSS.n57 0.00104
R30744 VSS.n1138 VSS.n77 0.00104
R30745 VSS.n1142 VSS.n36 0.00104
R30746 VSS.n37 VSS.n34 0.00104
R30747 DVSS VSS.n1073 0.00102
R30748 VSS.n750 VSS.n331 0.00101
R30749 VSS.n753 VSS.n752 0.00101
R30750 VSS.n498 VSS.n330 0.00101
R30751 VSS.n5114 VSS.n5113 0.001
R30752 VSS.n5072 VSS.n4358 0.001
R30753 VSS.n4924 VSS.n4923 0.001
R30754 VSS.n4881 VSS.n2282 0.001
R30755 VSS.n5116 VSS.n4295 0.001
R30756 VSS.n4692 VSS.n4642 0.001
R30757 VSS.n4839 VSS.n4565 0.001
R30758 VSS.n4625 VSS.n4624 0.001
R30759 VSS.n1056 VSS.n100 0.00098
R30760 VSS.n1055 VSS.n97 0.00098
R30761 VSS.n1054 VSS.n1009 0.00098
R30762 VSS.n2378 VSS.n2377 0.00095
R30763 VSS.n4500 VSS.n4499 0.00094335
R30764 VSS.n4790 VSS.n4789 0.00094335
R30765 VSS.n381 VSS.n352 0.00092
R30766 VSS.n582 VSS.n581 0.00092
R30767 VSS.n574 VSS.n375 0.00092
R30768 VSS.n1396 VSS.n32 0.000885714
R30769 VSS.n3045 VSS.n2835 0.000856671
R30770 VSS.n3036 VSS.n2829 0.000856671
R30771 VSS.n4300 DVSS 0.000721675
R30772 DVSS VSS.n5118 0.000721675
R30773 VSS.n5155 DVSS 0.000687793
R30774 DVSS VSS.n1086 0.00068
R30775 VSS.n1085 DVSS 0.00068
R30776 VSS.n5708 VSS 0.000671429
R30777 VSS.n2695 VSS 0.000671429
R30778 VSS.n3185 DVSS 0.000671429
R30779 DVSS VSS.n3580 0.000671429
R30780 VSS.n1837 DVSS 0.000671429
R30781 VSS.n1398 DVSS 0.000671429
R30782 VSS.n5177 DVSS 0.000671429
R30783 VSS.n3016 VSS.n3015 0.000628571
R30784 VSS.n3364 VSS.n3363 0.000628571
R30785 VSS.n2986 VSS.n2904 0.000628571
R30786 VSS.n2993 VSS.n2987 0.000628571
R30787 VSS.n2992 VSS.n2985 0.000628571
R30788 VSS.n2995 VSS.n2983 0.000628571
R30789 VSS.n2996 VSS.n2920 0.000628571
R30790 VSS.n2979 VSS.n2922 0.000628571
R30791 VSS.n3002 VSS.n2919 0.000628571
R30792 VSS.n3351 VSS.n2923 0.000628571
R30793 VSS.n3349 VSS.n2924 0.000628571
R30794 VSS.n2931 VSS.n2930 0.000628571
R30795 VSS.n3343 VSS.n3342 0.000628571
R30796 VSS.n3061 VSS.n2932 0.000628571
R30797 VSS.n3064 VSS.n2948 0.000628571
R30798 VSS.n3333 VSS.n2950 0.000628571
R30799 VSS.n3325 VSS.n3324 0.000628571
R30800 VSS.n2960 VSS.n2959 0.000628571
R30801 VSS.n3113 VSS.n3112 0.000628571
R30802 VSS.n3121 VSS.n3120 0.000628571
R30803 VSS.n3129 VSS.n3100 0.000628571
R30804 VSS.n3128 VSS.n3101 0.000628571
R30805 VSS.n3103 VSS.n3077 0.000628571
R30806 VSS.n3081 VSS.n3080 0.000628571
R30807 VSS.n3302 VSS.n3082 0.000628571
R30808 VSS.n3089 VSS.n3088 0.000628571
R30809 VSS.n3296 VSS.n3295 0.000628571
R30810 VSS.n3145 VSS.n3090 0.000628571
R30811 VSS.n3287 VSS.n3146 0.000628571
R30812 VSS.n3286 VSS.n3147 0.000628571
R30813 VSS.n3277 VSS.n3276 0.000628571
R30814 VSS.n3280 VSS.n3279 0.000628571
R30815 DVSS VSS.n2161 0.00058
R30816 DVSS VSS.n1025 0.00058
R30817 VSS.n5169 VSS.n2271 0.000570422
R30818 VSS.n5681 VSS.n1170 0.000566519
R30819 VSS.n5170 VSS.n2267 0.000564286
R30820 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_logic_pupd_0.comp018green_std_xor2_0.nmos_6p0_CDNS_4066195314530_2.D.t0 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_logic_pupd_0.comp018green_std_xor2_0.nmos_6p0_CDNS_4066195314530_2.D 6.03467
R30821 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_logic_pupd_0.comp018green_std_xor2_0.nmos_6p0_CDNS_4066195314530_2.D GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_logic_pupd_0.comp018green_std_xor2_0.nmos_6p0_CDNS_4066195314530_2.D.t1 4.66477
R30822 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_logic_pupd_0.comp018green_std_xor2_0.nmos_6p0_CDNS_4066195314530_2.D.t0 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_logic_pupd_0.comp018green_std_xor2_0.nmos_6p0_CDNS_4066195314530_2.D.t3 3.2416
R30823 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_logic_pupd_0.comp018green_std_xor2_0.nmos_6p0_CDNS_4066195314530_2.D GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_logic_pupd_0.comp018green_std_xor2_0.nmos_6p0_CDNS_4066195314530_2.D.t2 3.17822
R30824 VDD.n176 VDD.n33 512.403
R30825 VDD VDD.t36 378.373
R30826 VDD.n332 VDD.t63 352.072
R30827 VDD.t24 VDD.t44 321.485
R30828 VDD.t36 VDD.t57 321.485
R30829 VDD.t65 VDD.t63 321.485
R30830 VDD.n388 VDD.t32 314.901
R30831 VDD.n335 VDD.t40 280.788
R30832 VDD.t34 VDD.n321 280.702
R30833 VDD.t53 VDD.n316 278.981
R30834 VDD.n316 VDD.t55 278.981
R30835 VDD.t61 VDD.n103 264.098
R30836 VDD.t20 VDD.n96 263.524
R30837 VDD.n96 VDD.t18 263.524
R30838 VDD.n400 VDD.t28 248.441
R30839 VDD.n813 VDD.n802 227.274
R30840 VDD.n819 VDD.n796 227.274
R30841 VDD.n904 VDD.t16 224.88
R30842 VDD.n828 VDD.t51 223.204
R30843 VDD.n828 VDD.t14 223.204
R30844 VDD.n138 VDD.n137 211.415
R30845 VDD.t1 VDD.n900 202.791
R30846 VDD.n790 VDD.t3 202.791
R30847 VDD.n834 VDD.t12 202.791
R30848 VDD.t6 VDD.n696 201.413
R30849 VDD.t32 VDD.t48 188.564
R30850 VDD.t48 VDD.t30 188.564
R30851 VDD.t30 VDD.t46 188.564
R30852 VDD.t46 VDD.t42 188.564
R30853 VDD.t26 VDD.t24 188.564
R30854 VDD.t66 VDD.t26 188.564
R30855 VDD.t28 VDD.t66 188.564
R30856 VDD.n703 VDD.t8 187.478
R30857 VDD.n696 VDD.t10 183.157
R30858 VDD.n318 VDD.t65 173.88
R30859 VDD.t57 VDD.n318 147.605
R30860 VDD.n399 VDD.t42 139.105
R30861 VDD.n813 VDD.t39 113.636
R30862 VDD.t39 VDD.n796 113.636
R30863 VDD.n651 VDD.n628 105.84
R30864 VDD.t5 VDD.n628 105.84
R30865 VDD.t5 VDD.n619 105.84
R30866 VDD.n670 VDD.n619 105.84
R30867 VDD.n322 VDD.t34 94.2818
R30868 VDD.n322 VDD.t53 94.2818
R30869 VDD.n334 VDD.t55 94.2818
R30870 VDD.t40 VDD.n334 94.2818
R30871 VDD.n137 VDD.n22 93.6531
R30872 VDD.n901 VDD.t1 82.4504
R30873 VDD.n827 VDD.t3 82.4504
R30874 VDD.t12 VDD.n833 82.4504
R30875 VDD.n193 VDD.t22 80.5329
R30876 VDD.n192 VDD.t38 78.388
R30877 VDD.t22 VDD.n192 78.388
R30878 VDD.n117 VDD.n50 75.7185
R30879 VDD.n117 VDD.t58 75.7185
R30880 VDD.n131 VDD.t58 75.7185
R30881 VDD.n131 VDD.n33 75.7185
R30882 VDD.n176 VDD.n38 75.7185
R30883 VDD.t0 VDD.n161 75.7185
R30884 VDD.n161 VDD.n27 75.7185
R30885 VDD.n702 VDD.t10 73.6165
R30886 VDD.n697 VDD.n695 70.1484
R30887 VDD.t8 VDD.n702 70.083
R30888 VDD.n137 VDD.t38 66.6298
R30889 VDD.n901 VDD.t16 61.249
R30890 VDD.t51 VDD.n827 61.249
R30891 VDD.n833 VDD.t14 61.249
R30892 VDD.n103 VDD.n100 53.6905
R30893 VDD.n193 VDD.n22 49.5691
R30894 VDD.t44 VDD.n399 49.4595
R30895 VDD.n792 VDD.t68 46.7726
R30896 VDD.t0 VDD.n138 45.0397
R30897 VDD.n88 VDD.n82 45.0389
R30898 VDD.n98 VDD.n97 45.0389
R30899 VDD.n105 VDD.n104 45.0389
R30900 VDD.n113 VDD.n112 44.9149
R30901 VDD.n191 VDD.n23 43.8205
R30902 VDD.n792 VDD.t50 41.2455
R30903 VDD.n138 VDD.n38 30.6794
R30904 VDD.n95 VDD.n94 29.7505
R30905 VDD.n94 VDD.n87 23.9405
R30906 VDD.n94 VDD.n93 23.9405
R30907 VDD VDD.t23 11.0117
R30908 VDD.n814 VDD.n801 10.5005
R30909 VDD.n814 VDD.n798 10.5005
R30910 VDD.n818 VDD.n798 10.5005
R30911 VDD.n808 VDD.n807 10.5005
R30912 VDD.n812 VDD.n803 10.5005
R30913 VDD.n812 VDD.n795 10.5005
R30914 VDD.n820 VDD.n795 10.5005
R30915 VDD.n23 VDD.n22 10.4028
R30916 VDD.n68 VDD.n67 10.1505
R30917 VDD.n71 VDD.n68 10.1505
R30918 VDD.n58 VDD.n52 10.1505
R30919 VDD.n55 VDD.n52 10.1505
R30920 VDD.n186 VDD.n185 10.1505
R30921 VDD.n175 VDD.n169 10.1505
R30922 VDD.n169 VDD.n167 10.1505
R30923 VDD.n167 VDD.n26 10.1505
R30924 VDD.n188 VDD.n26 10.1505
R30925 VDD.n166 VDD.n163 10.1505
R30926 VDD.n164 VDD.n28 10.1505
R30927 VDD.n172 VDD.n171 10.1505
R30928 VDD.n116 VDD.n63 10.1505
R30929 VDD.n116 VDD.n42 10.1505
R30930 VDD.n132 VDD.n42 10.1505
R30931 VDD.n133 VDD.n132 10.1505
R30932 VDD.n66 VDD.n51 10.1505
R30933 VDD.n66 VDD.n43 10.1505
R30934 VDD.n76 VDD.n75 10.1505
R30935 VDD.n178 VDD.n32 10.1505
R30936 VDD.n148 VDD.n37 10.1505
R30937 VDD.n148 VDD.n141 10.1505
R30938 VDD.n142 VDD.n141 10.1505
R30939 VDD.n151 VDD.n142 10.1505
R30940 VDD.n156 VDD.n155 10.1505
R30941 VDD.n155 VDD.n154 10.1505
R30942 VDD.n140 VDD.n139 10.1505
R30943 VDD.n160 VDD.n159 10.1505
R30944 VDD.n62 VDD.n60 10.1505
R30945 VDD.n130 VDD.n45 10.1505
R30946 VDD.n127 VDD.n46 10.1505
R30947 VDD.n118 VDD.n49 10.1505
R30948 VDD.n119 VDD.n118 10.1505
R30949 VDD.n119 VDD.n44 10.1505
R30950 VDD.n122 VDD.n44 10.1505
R30951 VDD.n639 VDD.n637 10.1505
R30952 VDD.n646 VDD.n645 10.1505
R30953 VDD.n645 VDD.n635 10.1505
R30954 VDD.n649 VDD.n627 10.1505
R30955 VDD.n665 VDD.n627 10.1505
R30956 VDD.n665 VDD.n624 10.1505
R30957 VDD.n668 VDD.n624 10.1505
R30958 VDD.n643 VDD.n638 10.1505
R30959 VDD.n638 VDD.n629 10.1505
R30960 VDD.n629 VDD.n617 10.1505
R30961 VDD.n672 VDD.n617 10.1505
R30962 VDD.n659 VDD.n618 10.1505
R30963 VDD.n623 VDD.n622 10.1505
R30964 VDD.n656 VDD.n622 10.1505
R30965 VDD.n653 VDD.n630 10.1505
R30966 VDD.n664 VDD.n630 10.1505
R30967 VDD.n664 VDD.n631 10.1505
R30968 VDD.n658 VDD.n631 10.1505
R30969 VDD.n818 VDD.n797 7.3505
R30970 VDD.n183 VDD.n28 7.0005
R30971 VDD.n175 VDD.n174 7.0005
R30972 VDD.n78 VDD.n63 7.0005
R30973 VDD.n145 VDD.n37 7.0005
R30974 VDD.n124 VDD.n122 7.0005
R30975 VDD.n653 VDD.n634 7.0005
R30976 VDD.n660 VDD.n658 7.0005
R30977 VDD.n823 VDD.n822 6.78118
R30978 VDD.n135 VDD.n23 6.45932
R30979 VDD.n159 VDD.n158 6.3005
R30980 VDD.n161 VDD.n160 6.3005
R30981 VDD.t0 VDD.n140 6.3005
R30982 VDD.n139 VDD.n38 6.3005
R30983 VDD.n179 VDD.n178 6.3005
R30984 VDD.n32 VDD 6.3005
R30985 VDD.n146 VDD.n145 6.3005
R30986 VDD.n154 VDD.n153 6.3005
R30987 VDD.n155 VDD 6.3005
R30988 VDD.n155 VDD.n27 6.3005
R30989 VDD.n157 VDD.n156 6.3005
R30990 VDD.n152 VDD.n151 6.3005
R30991 VDD.n150 VDD.n142 6.3005
R30992 VDD.n161 VDD.n142 6.3005
R30993 VDD VDD.n141 6.3005
R30994 VDD.t0 VDD.n141 6.3005
R30995 VDD.n149 VDD.n148 6.3005
R30996 VDD.n148 VDD.n38 6.3005
R30997 VDD.n147 VDD.n37 6.3005
R30998 VDD.n176 VDD.n37 6.3005
R30999 VDD.n79 VDD.n78 6.3005
R31000 VDD.n76 VDD 6.3005
R31001 VDD.n75 VDD.n74 6.3005
R31002 VDD.n174 VDD.n173 6.3005
R31003 VDD VDD.n172 6.3005
R31004 VDD.n171 VDD.n170 6.3005
R31005 VDD.n183 VDD.n182 6.3005
R31006 VDD.n185 VDD 6.3005
R31007 VDD.n186 VDD.n25 6.3005
R31008 VDD.n181 VDD.n28 6.3005
R31009 VDD.n28 VDD.n27 6.3005
R31010 VDD.n164 VDD.n161 6.3005
R31011 VDD.t0 VDD.n166 6.3005
R31012 VDD.n163 VDD.n38 6.3005
R31013 VDD.n122 VDD.n121 6.3005
R31014 VDD.n122 VDD.n33 6.3005
R31015 VDD.n120 VDD.n44 6.3005
R31016 VDD.n131 VDD.n44 6.3005
R31017 VDD VDD.n119 6.3005
R31018 VDD.n119 VDD.t58 6.3005
R31019 VDD.n118 VDD.n48 6.3005
R31020 VDD.n118 VDD.n117 6.3005
R31021 VDD.n53 VDD.n49 6.3005
R31022 VDD.n125 VDD.n124 6.3005
R31023 VDD VDD.n46 6.3005
R31024 VDD.n127 VDD.n126 6.3005
R31025 VDD.n58 VDD.n57 6.3005
R31026 VDD VDD.n52 6.3005
R31027 VDD.n52 VDD.n50 6.3005
R31028 VDD.n56 VDD.n55 6.3005
R31029 VDD.n131 VDD.n130 6.3005
R31030 VDD.n45 VDD.t58 6.3005
R31031 VDD.n117 VDD.n62 6.3005
R31032 VDD.n60 VDD 6.3005
R31033 VDD.n131 VDD.n43 6.3005
R31034 VDD VDD.n66 6.3005
R31035 VDD.n66 VDD.t58 6.3005
R31036 VDD.n117 VDD.n51 6.3005
R31037 VDD.n72 VDD.n71 6.3005
R31038 VDD.n68 VDD 6.3005
R31039 VDD.n68 VDD.n33 6.3005
R31040 VDD.n67 VDD.n39 6.3005
R31041 VDD.n134 VDD.n133 6.3005
R31042 VDD.n132 VDD.n40 6.3005
R31043 VDD.n132 VDD.n131 6.3005
R31044 VDD VDD.n42 6.3005
R31045 VDD.t58 VDD.n42 6.3005
R31046 VDD.n116 VDD.n115 6.3005
R31047 VDD.n117 VDD.n116 6.3005
R31048 VDD.n114 VDD.n63 6.3005
R31049 VDD.n63 VDD.n50 6.3005
R31050 VDD.n26 VDD.n24 6.3005
R31051 VDD.n161 VDD.n26 6.3005
R31052 VDD VDD.n167 6.3005
R31053 VDD.n167 VDD.t0 6.3005
R31054 VDD.n169 VDD.n168 6.3005
R31055 VDD.n169 VDD.n38 6.3005
R31056 VDD.n175 VDD.n136 6.3005
R31057 VDD.n176 VDD.n175 6.3005
R31058 VDD.n189 VDD.n188 6.3005
R31059 VDD.n668 VDD.n667 6.3005
R31060 VDD.n666 VDD.n624 6.3005
R31061 VDD.n624 VDD.n619 6.3005
R31062 VDD VDD.n665 6.3005
R31063 VDD.n665 VDD.t5 6.3005
R31064 VDD.n627 VDD.n626 6.3005
R31065 VDD.n628 VDD.n627 6.3005
R31066 VDD.n649 VDD.n648 6.3005
R31067 VDD.n647 VDD.n646 6.3005
R31068 VDD VDD.n645 6.3005
R31069 VDD.n651 VDD.n645 6.3005
R31070 VDD.n635 VDD.n633 6.3005
R31071 VDD.n634 VDD.n632 6.3005
R31072 VDD VDD.n639 6.3005
R31073 VDD.n640 VDD.n637 6.3005
R31074 VDD.n617 VDD.n616 6.3005
R31075 VDD.n619 VDD.n617 6.3005
R31076 VDD VDD.n629 6.3005
R31077 VDD.t5 VDD.n629 6.3005
R31078 VDD.n641 VDD.n638 6.3005
R31079 VDD.n638 VDD.n628 6.3005
R31080 VDD.n643 VDD.n642 6.3005
R31081 VDD.n657 VDD.n656 6.3005
R31082 VDD VDD.n622 6.3005
R31083 VDD.n670 VDD.n622 6.3005
R31084 VDD.n625 VDD.n623 6.3005
R31085 VDD.n662 VDD.n658 6.3005
R31086 VDD.n663 VDD.n631 6.3005
R31087 VDD.n631 VDD.n619 6.3005
R31088 VDD.n664 VDD 6.3005
R31089 VDD.t5 VDD.n664 6.3005
R31090 VDD.n655 VDD.n630 6.3005
R31091 VDD.n630 VDD.n628 6.3005
R31092 VDD.n654 VDD.n653 6.3005
R31093 VDD VDD.n659 6.3005
R31094 VDD.n661 VDD.n660 6.3005
R31095 VDD.n618 VDD.n615 6.3005
R31096 VDD.n673 VDD.n672 6.3005
R31097 VDD.n809 VDD.n808 6.3005
R31098 VDD.n807 VDD.n806 6.3005
R31099 VDD.n799 VDD.n797 6.3005
R31100 VDD.n818 VDD.n817 6.3005
R31101 VDD.n819 VDD.n818 6.3005
R31102 VDD.n816 VDD.n798 6.3005
R31103 VDD.n798 VDD.n796 6.3005
R31104 VDD.n815 VDD.n814 6.3005
R31105 VDD.n814 VDD.n813 6.3005
R31106 VDD.n801 VDD.n800 6.3005
R31107 VDD.n795 VDD.n793 6.3005
R31108 VDD.n796 VDD.n795 6.3005
R31109 VDD.n812 VDD.n811 6.3005
R31110 VDD.n813 VDD.n812 6.3005
R31111 VDD.n810 VDD.n803 6.3005
R31112 VDD.n820 VDD.n819 6.3005
R31113 VDD.n106 VDD.n105 5.80576
R31114 VDD.n111 VDD.n110 5.63063
R31115 VDD.n821 VDD.n794 5.18619
R31116 VDD.n70 VDD.n69 5.06227
R31117 VDD.n177 VDD.n30 5.06227
R31118 VDD.n162 VDD.n35 5.06227
R31119 VDD.n129 VDD.n128 5.06227
R31120 VDD.n65 VDD.n64 5.06227
R31121 VDD.n325 VDD.n315 4.62839
R31122 VDD.n331 VDD.n330 4.62839
R31123 VDD.n327 VDD.n315 4.5005
R31124 VDD.n330 VDD.n329 4.5005
R31125 VDD.n206 VDD.n8 4.5005
R31126 VDD.n555 VDD.n206 4.5005
R31127 VDD.n555 VDD.n209 4.5005
R31128 VDD.n555 VDD.n13 4.5005
R31129 VDD.n555 VDD.n211 4.5005
R31130 VDD.n555 VDD.n12 4.5005
R31131 VDD.n555 VDD.n213 4.5005
R31132 VDD.n555 VDD.n11 4.5005
R31133 VDD.n555 VDD.n554 4.5005
R31134 VDD.n555 VDD.n10 4.5005
R31135 VDD.n556 VDD.n8 4.5005
R31136 VDD.n556 VDD.n555 4.5005
R31137 VDD.n197 VDD.n196 4.5005
R31138 VDD.n196 VDD.n20 4.5005
R31139 VDD.n198 VDD.n197 4.5005
R31140 VDD.n201 VDD.n15 4.5005
R31141 VDD.n202 VDD.n201 4.5005
R31142 VDD.n203 VDD.n202 4.5005
R31143 VDD.n928 VDD.n906 4.5005
R31144 VDD.n930 VDD.n906 4.5005
R31145 VDD.n930 VDD.n908 4.5005
R31146 VDD.n930 VDD.n6 4.5005
R31147 VDD.n930 VDD.n909 4.5005
R31148 VDD.n930 VDD.n5 4.5005
R31149 VDD.n930 VDD.n910 4.5005
R31150 VDD.n930 VDD.n4 4.5005
R31151 VDD.n930 VDD.n911 4.5005
R31152 VDD.n930 VDD.n3 4.5005
R31153 VDD.n929 VDD.n928 4.5005
R31154 VDD.n930 VDD.n929 4.5005
R31155 VDD.n336 VDD.n335 4.14897
R31156 VDD.n693 VDD.n674 4.13212
R31157 VDD.n823 VDD.n792 4.0005
R31158 VDD.n797 VDD.n794 2.86464
R31159 VDD.n184 VDD.n183 2.81177
R31160 VDD.n163 VDD.n162 2.81177
R31161 VDD.n165 VDD.n164 2.81177
R31162 VDD.n174 VDD.n34 2.81177
R31163 VDD.n65 VDD.n51 2.81177
R31164 VDD.n78 VDD.n77 2.81177
R31165 VDD.n36 VDD.n32 2.81177
R31166 VDD.n139 VDD.n30 2.81177
R31167 VDD.n160 VDD.n31 2.81177
R31168 VDD.n140 VDD.n31 2.81177
R31169 VDD.n145 VDD.n36 2.81177
R31170 VDD.n77 VDD.n76 2.81177
R31171 VDD.n172 VDD.n34 2.81177
R31172 VDD.n185 VDD.n184 2.81177
R31173 VDD.n166 VDD.n165 2.81177
R31174 VDD.n61 VDD.n45 2.81177
R31175 VDD.n123 VDD.n46 2.81177
R31176 VDD.n124 VDD.n123 2.81177
R31177 VDD.n130 VDD.n129 2.81177
R31178 VDD.n62 VDD.n61 2.81177
R31179 VDD.n69 VDD.n43 2.81177
R31180 VDD.n636 VDD.n634 2.81177
R31181 VDD.n639 VDD.n636 2.81177
R31182 VDD.n660 VDD.n621 2.81177
R31183 VDD.n659 VDD.n621 2.81177
R31184 VDD.n194 VDD.n193 2.76632
R31185 VDD.n396 VDD.t25 2.46086
R31186 VDD.n294 VDD.t29 2.46086
R31187 VDD.n698 VDD.t7 2.36071
R31188 VDD.n821 VDD.n820 2.32205
R31189 VDD.n808 VDD.n804 2.32205
R31190 VDD.n807 VDD.n805 2.32205
R31191 VDD.n805 VDD.n801 2.32205
R31192 VDD.n804 VDD.n803 2.32205
R31193 VDD.n21 VDD.n19 2.25705
R31194 VDD.n133 VDD.n41 2.251
R31195 VDD.n59 VDD.n58 2.251
R31196 VDD.n54 VDD.n49 2.251
R31197 VDD.n187 VDD.n186 2.251
R31198 VDD.n171 VDD.n35 2.251
R31199 VDD.n75 VDD.n64 2.251
R31200 VDD.n159 VDD.n143 2.251
R31201 VDD.n154 VDD.n144 2.251
R31202 VDD.n178 VDD.n177 2.251
R31203 VDD.n156 VDD.n143 2.251
R31204 VDD.n151 VDD.n144 2.251
R31205 VDD.n128 VDD.n127 2.251
R31206 VDD.n55 VDD.n54 2.251
R31207 VDD.n60 VDD.n59 2.251
R31208 VDD.n71 VDD.n70 2.251
R31209 VDD.n67 VDD.n41 2.251
R31210 VDD.n188 VDD.n187 2.251
R31211 VDD.n644 VDD.n637 2.251
R31212 VDD.n650 VDD.n649 2.251
R31213 VDD.n652 VDD.n635 2.251
R31214 VDD.n650 VDD.n646 2.251
R31215 VDD.n644 VDD.n643 2.251
R31216 VDD.n671 VDD.n618 2.251
R31217 VDD.n669 VDD.n668 2.251
R31218 VDD.n656 VDD.n620 2.251
R31219 VDD.n669 VDD.n623 2.251
R31220 VDD.n658 VDD.n620 2.251
R31221 VDD.n653 VDD.n652 2.251
R31222 VDD.n672 VDD.n671 2.251
R31223 VDD.n200 VDD.n19 2.24475
R31224 VDD.n205 VDD.n14 2.24475
R31225 VDD.n199 VDD.n20 2.24405
R31226 VDD.n204 VDD.n15 2.24405
R31227 VDD.n17 VDD.n16 2.24405
R31228 VDD.n551 VDD.n217 2.24304
R31229 VDD.n208 VDD.n8 2.24304
R31230 VDD.n551 VDD.n216 2.24304
R31231 VDD.n210 VDD.n8 2.24304
R31232 VDD.n551 VDD.n215 2.24304
R31233 VDD.n212 VDD.n8 2.24304
R31234 VDD.n552 VDD.n551 2.24304
R31235 VDD.n553 VDD.n8 2.24304
R31236 VDD.n551 VDD.n7 2.24304
R31237 VDD.n928 VDD.n924 2.24304
R31238 VDD.n917 VDD.n913 2.24304
R31239 VDD.n928 VDD.n925 2.24304
R31240 VDD.n917 VDD.n914 2.24304
R31241 VDD.n928 VDD.n926 2.24304
R31242 VDD.n917 VDD.n915 2.24304
R31243 VDD.n928 VDD.n927 2.24304
R31244 VDD.n917 VDD.n916 2.24304
R31245 VDD.n917 VDD.n912 2.24304
R31246 VDD.n101 VDD.t62 2.12386
R31247 VDD.n319 VDD.t37 2.12292
R31248 VDD.n905 VDD.n556 2.10965
R31249 VDD.n328 VDD.t64 2.08373
R31250 VDD.n81 VDD.t60 2.0836
R31251 VDD.n143 VDD.n27 2.026
R31252 VDD.n177 VDD.n176 2.026
R31253 VDD.n144 VDD.n27 2.026
R31254 VDD.n64 VDD.n50 2.026
R31255 VDD.n176 VDD.n35 2.026
R31256 VDD.n187 VDD.n27 2.026
R31257 VDD.n54 VDD.n50 2.026
R31258 VDD.n59 VDD.n50 2.026
R31259 VDD.n128 VDD.n33 2.026
R31260 VDD.n70 VDD.n33 2.026
R31261 VDD.n41 VDD.n33 2.026
R31262 VDD.n670 VDD.n669 2.026
R31263 VDD.n651 VDD.n650 2.026
R31264 VDD.n652 VDD.n651 2.026
R31265 VDD.n651 VDD.n644 2.026
R31266 VDD.n670 VDD.n620 2.026
R31267 VDD.n671 VDD.n670 2.026
R31268 VDD.n804 VDD.n802 1.99047
R31269 VDD.n805 VDD.n802 1.99047
R31270 VDD.n822 VDD.n821 1.99047
R31271 VDD.n313 VDD.t41 1.96281
R31272 VDD.n903 VDD.t17 1.96281
R31273 VDD.n557 VDD.t2 1.96281
R31274 VDD.n700 VDD.t11 1.96281
R31275 VDD.n614 VDD.t9 1.96281
R31276 VDD.n585 VDD.t13 1.96281
R31277 VDD.n831 VDD.t15 1.96281
R31278 VDD.n791 VDD.t4 1.96281
R31279 VDD.n314 VDD.t56 1.92255
R31280 VDD.n324 VDD.t54 1.92255
R31281 VDD.n320 VDD.t35 1.92255
R31282 VDD.n790 VDD.n789 1.8507
R31283 VDD.n835 VDD.n834 1.8507
R31284 VDD.n900 VDD.n899 1.8228
R31285 VDD.n97 VDD.t20 1.81731
R31286 VDD.n88 VDD.t18 1.81731
R31287 VDD.n104 VDD.t61 1.81731
R31288 VDD.n401 VDD.n400 1.80879
R31289 VDD.n388 VDD.n387 1.8024
R31290 VDD.n702 VDD.n701 1.8005
R31291 VDD.n389 VDD.t33 1.78389
R31292 VDD.n397 VDD.t45 1.78389
R31293 VDD VDD.n31 1.74562
R31294 VDD VDD.n30 1.74562
R31295 VDD.n176 VDD.n36 1.74562
R31296 VDD.n77 VDD.n50 1.74562
R31297 VDD.n176 VDD.n34 1.74562
R31298 VDD.n184 VDD.n27 1.74562
R31299 VDD.n165 VDD 1.74562
R31300 VDD.n162 VDD 1.74562
R31301 VDD.n123 VDD.n33 1.74562
R31302 VDD.n129 VDD 1.74562
R31303 VDD.n61 VDD 1.74562
R31304 VDD.n69 VDD 1.74562
R31305 VDD VDD.n65 1.74562
R31306 VDD.n651 VDD.n636 1.74562
R31307 VDD.n670 VDD.n621 1.74562
R31308 VDD.n395 VDD.n394 1.73286
R31309 VDD.n326 VDD.n316 1.72301
R31310 VDD.n819 VDD.n794 1.71918
R31311 VDD.n905 VDD.n904 1.70597
R31312 VDD.n112 VDD.t59 1.67055
R31313 VDD.n112 VDD.n111 1.63706
R31314 VDD.n83 VDD.t19 1.58219
R31315 VDD.n85 VDD.t21 1.58219
R31316 VDD.n323 VDD.n322 1.5755
R31317 VDD.n334 VDD.n333 1.5755
R31318 VDD.n902 VDD.n901 1.5755
R31319 VDD.n833 VDD.n832 1.5755
R31320 VDD.n827 VDD.n826 1.5755
R31321 VDD.n337 VDD.n336 1.50189
R31322 VDD.n353 VDD.n336 1.50166
R31323 VDD.n829 VDD.n586 1.50061
R31324 VDD.n704 VDD.n703 1.46392
R31325 VDD.n824 VDD.t52 1.36414
R31326 VDD VDD.n697 1.27477
R31327 VDD.n391 VDD.n390 1.26489
R31328 VDD.n393 VDD.n392 1.26489
R31329 VDD.n93 VDD.n92 1.2605
R31330 VDD.n87 VDD.n86 1.2605
R31331 VDD.n100 VDD.n99 1.2605
R31332 VDD.n697 VDD.t6 1.24589
R31333 VDD.n103 VDD.n102 1.15029
R31334 VDD.n834 VDD.n585 1.10418
R31335 VDD.n791 VDD.n790 1.10418
R31336 VDD.n900 VDD.n557 1.1
R31337 VDD.n109 VDD.n83 1.07633
R31338 VDD.n107 VDD.n85 1.07633
R31339 VDD.n703 VDD.n614 1.06559
R31340 VDD.n110 VDD.n82 1.06155
R31341 VDD.n108 VDD.n84 1.06155
R31342 VDD.n106 VDD.n98 1.06155
R31343 VDD.n105 VDD.n99 0.973921
R31344 VDD.n92 VDD.n82 0.964726
R31345 VDD.n98 VDD.n86 0.964726
R31346 VDD.n694 VDD.n693 0.921424
R31347 VDD.n824 VDD 0.869566
R31348 VDD.n830 VDD.n829 0.861978
R31349 VDD.n699 VDD.n694 0.857799
R31350 VDD.n829 VDD.n828 0.788
R31351 VDD.n400 VDD.n294 0.756026
R31352 VDD.n394 VDD.t27 0.7285
R31353 VDD.n394 VDD.t67 0.7285
R31354 VDD.n206 VDD.n205 0.671
R31355 VDD.n389 VDD.n388 0.651808
R31356 VDD.n318 VDD.n317 0.6005
R31357 VDD.n825 VDD.n824 0.600169
R31358 VDD.n113 VDD.n80 0.577559
R31359 VDD.n95 VDD.n84 0.573227
R31360 VDD.n96 VDD.n95 0.573227
R31361 VDD.n90 VDD.n84 0.557079
R31362 VDD.n107 VDD.n106 0.555895
R31363 VDD.n110 VDD.n109 0.555895
R31364 VDD.n391 VDD.n389 0.545794
R31365 VDD.n393 VDD.n391 0.545794
R31366 VDD.n396 VDD.n395 0.545794
R31367 VDD.n395 VDD.n294 0.545794
R31368 VDD.n91 VDD.n83 0.542091
R31369 VDD.n89 VDD.n85 0.542091
R31370 VDD.n693 VDD.n692 0.541547
R31371 VDD.n191 VDD.n190 0.5255
R31372 VDD.n192 VDD.n191 0.5255
R31373 VDD.n390 VDD.t49 0.5205
R31374 VDD.n390 VDD.t31 0.5205
R31375 VDD.n392 VDD.t47 0.5205
R31376 VDD.n392 VDD.t43 0.5205
R31377 VDD.n194 VDD 0.499471
R31378 VDD.n551 VDD.n550 0.456899
R31379 VDD.n928 VDD.n923 0.456899
R31380 VDD.n384 VDD.n383 0.4505
R31381 VDD.n382 VDD.n297 0.4505
R31382 VDD.n381 VDD.n380 0.4505
R31383 VDD.n299 VDD.n298 0.4505
R31384 VDD.n376 VDD.n375 0.4505
R31385 VDD.n374 VDD.n302 0.4505
R31386 VDD.n373 VDD.n372 0.4505
R31387 VDD.n304 VDD.n303 0.4505
R31388 VDD.n368 VDD.n367 0.4505
R31389 VDD.n366 VDD.n306 0.4505
R31390 VDD.n365 VDD.n364 0.4505
R31391 VDD.n308 VDD.n307 0.4505
R31392 VDD.n360 VDD.n359 0.4505
R31393 VDD.n358 VDD.n310 0.4505
R31394 VDD.n357 VDD.n356 0.4505
R31395 VDD.n312 VDD.n311 0.4505
R31396 VDD.n351 VDD.n350 0.4505
R31397 VDD.n349 VDD.n338 0.4505
R31398 VDD.n348 VDD.n347 0.4505
R31399 VDD.n340 VDD.n339 0.4505
R31400 VDD.n343 VDD.n342 0.4505
R31401 VDD.n292 VDD.n291 0.4505
R31402 VDD.n404 VDD.n403 0.4505
R31403 VDD.n405 VDD.n290 0.4505
R31404 VDD.n407 VDD.n406 0.4505
R31405 VDD.n288 VDD.n287 0.4505
R31406 VDD.n412 VDD.n411 0.4505
R31407 VDD.n413 VDD.n286 0.4505
R31408 VDD.n415 VDD.n414 0.4505
R31409 VDD.n284 VDD.n283 0.4505
R31410 VDD.n420 VDD.n419 0.4505
R31411 VDD.n421 VDD.n282 0.4505
R31412 VDD.n423 VDD.n422 0.4505
R31413 VDD.n280 VDD.n279 0.4505
R31414 VDD.n428 VDD.n427 0.4505
R31415 VDD.n429 VDD.n278 0.4505
R31416 VDD.n431 VDD.n430 0.4505
R31417 VDD.n276 VDD.n275 0.4505
R31418 VDD.n436 VDD.n435 0.4505
R31419 VDD.n437 VDD.n274 0.4505
R31420 VDD.n439 VDD.n438 0.4505
R31421 VDD.n272 VDD.n271 0.4505
R31422 VDD.n444 VDD.n443 0.4505
R31423 VDD.n445 VDD.n270 0.4505
R31424 VDD.n447 VDD.n446 0.4505
R31425 VDD.n268 VDD.n267 0.4505
R31426 VDD.n452 VDD.n451 0.4505
R31427 VDD.n453 VDD.n266 0.4505
R31428 VDD.n455 VDD.n454 0.4505
R31429 VDD.n264 VDD.n263 0.4505
R31430 VDD.n460 VDD.n459 0.4505
R31431 VDD.n461 VDD.n262 0.4505
R31432 VDD.n463 VDD.n462 0.4505
R31433 VDD.n260 VDD.n259 0.4505
R31434 VDD.n468 VDD.n467 0.4505
R31435 VDD.n469 VDD.n258 0.4505
R31436 VDD.n471 VDD.n470 0.4505
R31437 VDD.n256 VDD.n255 0.4505
R31438 VDD.n476 VDD.n475 0.4505
R31439 VDD.n477 VDD.n254 0.4505
R31440 VDD.n479 VDD.n478 0.4505
R31441 VDD.n252 VDD.n251 0.4505
R31442 VDD.n484 VDD.n483 0.4505
R31443 VDD.n485 VDD.n250 0.4505
R31444 VDD.n487 VDD.n486 0.4505
R31445 VDD.n248 VDD.n247 0.4505
R31446 VDD.n492 VDD.n491 0.4505
R31447 VDD.n493 VDD.n246 0.4505
R31448 VDD.n495 VDD.n494 0.4505
R31449 VDD.n244 VDD.n243 0.4505
R31450 VDD.n500 VDD.n499 0.4505
R31451 VDD.n501 VDD.n242 0.4505
R31452 VDD.n503 VDD.n502 0.4505
R31453 VDD.n240 VDD.n239 0.4505
R31454 VDD.n508 VDD.n507 0.4505
R31455 VDD.n509 VDD.n238 0.4505
R31456 VDD.n511 VDD.n510 0.4505
R31457 VDD.n236 VDD.n235 0.4505
R31458 VDD.n516 VDD.n515 0.4505
R31459 VDD.n517 VDD.n234 0.4505
R31460 VDD.n519 VDD.n518 0.4505
R31461 VDD.n232 VDD.n231 0.4505
R31462 VDD.n524 VDD.n523 0.4505
R31463 VDD.n525 VDD.n230 0.4505
R31464 VDD.n527 VDD.n526 0.4505
R31465 VDD.n228 VDD.n227 0.4505
R31466 VDD.n532 VDD.n531 0.4505
R31467 VDD.n533 VDD.n226 0.4505
R31468 VDD.n535 VDD.n534 0.4505
R31469 VDD.n224 VDD.n223 0.4505
R31470 VDD.n540 VDD.n539 0.4505
R31471 VDD.n541 VDD.n222 0.4505
R31472 VDD.n543 VDD.n542 0.4505
R31473 VDD.n546 VDD.n220 0.4505
R31474 VDD.n547 VDD.n219 0.4505
R31475 VDD.n549 VDD.n548 0.4505
R31476 VDD.n218 VDD.n214 0.4505
R31477 VDD.n548 VDD.n207 0.4505
R31478 VDD.n547 VDD.n9 0.4505
R31479 VDD.n546 VDD.n545 0.4505
R31480 VDD.n544 VDD.n543 0.4505
R31481 VDD.n222 VDD.n221 0.4505
R31482 VDD.n539 VDD.n538 0.4505
R31483 VDD.n537 VDD.n224 0.4505
R31484 VDD.n536 VDD.n535 0.4505
R31485 VDD.n226 VDD.n225 0.4505
R31486 VDD.n531 VDD.n530 0.4505
R31487 VDD.n529 VDD.n228 0.4505
R31488 VDD.n528 VDD.n527 0.4505
R31489 VDD.n230 VDD.n229 0.4505
R31490 VDD.n523 VDD.n522 0.4505
R31491 VDD.n521 VDD.n232 0.4505
R31492 VDD.n520 VDD.n519 0.4505
R31493 VDD.n234 VDD.n233 0.4505
R31494 VDD.n515 VDD.n514 0.4505
R31495 VDD.n513 VDD.n236 0.4505
R31496 VDD.n512 VDD.n511 0.4505
R31497 VDD.n238 VDD.n237 0.4505
R31498 VDD.n507 VDD.n506 0.4505
R31499 VDD.n505 VDD.n240 0.4505
R31500 VDD.n504 VDD.n503 0.4505
R31501 VDD.n242 VDD.n241 0.4505
R31502 VDD.n499 VDD.n498 0.4505
R31503 VDD.n497 VDD.n244 0.4505
R31504 VDD.n496 VDD.n495 0.4505
R31505 VDD.n246 VDD.n245 0.4505
R31506 VDD.n491 VDD.n490 0.4505
R31507 VDD.n489 VDD.n248 0.4505
R31508 VDD.n488 VDD.n487 0.4505
R31509 VDD.n250 VDD.n249 0.4505
R31510 VDD.n483 VDD.n482 0.4505
R31511 VDD.n481 VDD.n252 0.4505
R31512 VDD.n480 VDD.n479 0.4505
R31513 VDD.n254 VDD.n253 0.4505
R31514 VDD.n475 VDD.n474 0.4505
R31515 VDD.n473 VDD.n256 0.4505
R31516 VDD.n472 VDD.n471 0.4505
R31517 VDD.n258 VDD.n257 0.4505
R31518 VDD.n467 VDD.n466 0.4505
R31519 VDD.n465 VDD.n260 0.4505
R31520 VDD.n464 VDD.n463 0.4505
R31521 VDD.n262 VDD.n261 0.4505
R31522 VDD.n459 VDD.n458 0.4505
R31523 VDD.n457 VDD.n264 0.4505
R31524 VDD.n456 VDD.n455 0.4505
R31525 VDD.n266 VDD.n265 0.4505
R31526 VDD.n451 VDD.n450 0.4505
R31527 VDD.n449 VDD.n268 0.4505
R31528 VDD.n448 VDD.n447 0.4505
R31529 VDD.n270 VDD.n269 0.4505
R31530 VDD.n443 VDD.n442 0.4505
R31531 VDD.n441 VDD.n272 0.4505
R31532 VDD.n440 VDD.n439 0.4505
R31533 VDD.n274 VDD.n273 0.4505
R31534 VDD.n435 VDD.n434 0.4505
R31535 VDD.n433 VDD.n276 0.4505
R31536 VDD.n432 VDD.n431 0.4505
R31537 VDD.n278 VDD.n277 0.4505
R31538 VDD.n427 VDD.n426 0.4505
R31539 VDD.n425 VDD.n280 0.4505
R31540 VDD.n424 VDD.n423 0.4505
R31541 VDD.n282 VDD.n281 0.4505
R31542 VDD.n419 VDD.n418 0.4505
R31543 VDD.n417 VDD.n284 0.4505
R31544 VDD.n416 VDD.n415 0.4505
R31545 VDD.n286 VDD.n285 0.4505
R31546 VDD.n411 VDD.n410 0.4505
R31547 VDD.n409 VDD.n288 0.4505
R31548 VDD.n408 VDD.n407 0.4505
R31549 VDD.n290 VDD.n289 0.4505
R31550 VDD.n403 VDD.n402 0.4505
R31551 VDD.n293 VDD.n292 0.4505
R31552 VDD.n344 VDD.n343 0.4505
R31553 VDD.n345 VDD.n340 0.4505
R31554 VDD.n347 VDD.n346 0.4505
R31555 VDD.n341 VDD.n338 0.4505
R31556 VDD.n352 VDD.n351 0.4505
R31557 VDD.n354 VDD.n312 0.4505
R31558 VDD.n356 VDD.n355 0.4505
R31559 VDD.n310 VDD.n309 0.4505
R31560 VDD.n361 VDD.n360 0.4505
R31561 VDD.n362 VDD.n308 0.4505
R31562 VDD.n364 VDD.n363 0.4505
R31563 VDD.n306 VDD.n305 0.4505
R31564 VDD.n369 VDD.n368 0.4505
R31565 VDD.n370 VDD.n304 0.4505
R31566 VDD.n372 VDD.n371 0.4505
R31567 VDD.n302 VDD.n301 0.4505
R31568 VDD.n377 VDD.n376 0.4505
R31569 VDD.n378 VDD.n299 0.4505
R31570 VDD.n380 VDD.n379 0.4505
R31571 VDD.n300 VDD.n297 0.4505
R31572 VDD.n384 VDD.n296 0.4505
R31573 VDD.n386 VDD.n385 0.4505
R31574 VDD.n689 VDD.n688 0.4505
R31575 VDD.n687 VDD.n677 0.4505
R31576 VDD.n686 VDD.n685 0.4505
R31577 VDD.n681 VDD.n678 0.4505
R31578 VDD.n680 VDD.n679 0.4505
R31579 VDD.n612 VDD.n611 0.4505
R31580 VDD.n708 VDD.n707 0.4505
R31581 VDD.n709 VDD.n610 0.4505
R31582 VDD.n711 VDD.n710 0.4505
R31583 VDD.n608 VDD.n607 0.4505
R31584 VDD.n716 VDD.n715 0.4505
R31585 VDD.n717 VDD.n606 0.4505
R31586 VDD.n719 VDD.n718 0.4505
R31587 VDD.n604 VDD.n603 0.4505
R31588 VDD.n724 VDD.n723 0.4505
R31589 VDD.n725 VDD.n602 0.4505
R31590 VDD.n727 VDD.n726 0.4505
R31591 VDD.n600 VDD.n599 0.4505
R31592 VDD.n732 VDD.n731 0.4505
R31593 VDD.n733 VDD.n598 0.4505
R31594 VDD.n735 VDD.n734 0.4505
R31595 VDD.n596 VDD.n595 0.4505
R31596 VDD.n740 VDD.n739 0.4505
R31597 VDD.n741 VDD.n594 0.4505
R31598 VDD.n743 VDD.n742 0.4505
R31599 VDD.n592 VDD.n591 0.4505
R31600 VDD.n748 VDD.n747 0.4505
R31601 VDD.n749 VDD.n589 0.4505
R31602 VDD.n787 VDD.n786 0.4505
R31603 VDD.n785 VDD.n590 0.4505
R31604 VDD.n784 VDD.n783 0.4505
R31605 VDD.n751 VDD.n750 0.4505
R31606 VDD.n779 VDD.n778 0.4505
R31607 VDD.n777 VDD.n753 0.4505
R31608 VDD.n776 VDD.n775 0.4505
R31609 VDD.n773 VDD.n754 0.4505
R31610 VDD.n758 VDD.n755 0.4505
R31611 VDD.n769 VDD.n768 0.4505
R31612 VDD.n767 VDD.n757 0.4505
R31613 VDD.n766 VDD.n765 0.4505
R31614 VDD.n762 VDD.n759 0.4505
R31615 VDD.n761 VDD.n760 0.4505
R31616 VDD.n583 VDD.n582 0.4505
R31617 VDD.n839 VDD.n838 0.4505
R31618 VDD.n840 VDD.n581 0.4505
R31619 VDD.n842 VDD.n841 0.4505
R31620 VDD.n579 VDD.n578 0.4505
R31621 VDD.n847 VDD.n846 0.4505
R31622 VDD.n848 VDD.n577 0.4505
R31623 VDD.n850 VDD.n849 0.4505
R31624 VDD.n575 VDD.n574 0.4505
R31625 VDD.n855 VDD.n854 0.4505
R31626 VDD.n856 VDD.n573 0.4505
R31627 VDD.n858 VDD.n857 0.4505
R31628 VDD.n571 VDD.n570 0.4505
R31629 VDD.n863 VDD.n862 0.4505
R31630 VDD.n864 VDD.n569 0.4505
R31631 VDD.n866 VDD.n865 0.4505
R31632 VDD.n567 VDD.n566 0.4505
R31633 VDD.n871 VDD.n870 0.4505
R31634 VDD.n872 VDD.n565 0.4505
R31635 VDD.n874 VDD.n873 0.4505
R31636 VDD.n563 VDD.n562 0.4505
R31637 VDD.n879 VDD.n878 0.4505
R31638 VDD.n880 VDD.n560 0.4505
R31639 VDD.n897 VDD.n896 0.4505
R31640 VDD.n895 VDD.n561 0.4505
R31641 VDD.n894 VDD.n893 0.4505
R31642 VDD.n882 VDD.n881 0.4505
R31643 VDD.n889 VDD.n888 0.4505
R31644 VDD.n887 VDD.n885 0.4505
R31645 VDD.n886 VDD.n0 0.4505
R31646 VDD.n933 VDD.n2 0.4505
R31647 VDD.n920 VDD.n1 0.4505
R31648 VDD.n922 VDD.n921 0.4505
R31649 VDD.n919 VDD.n918 0.4505
R31650 VDD.n921 VDD.n907 0.4505
R31651 VDD.n931 VDD.n1 0.4505
R31652 VDD.n933 VDD.n932 0.4505
R31653 VDD.n883 VDD.n0 0.4505
R31654 VDD.n885 VDD.n884 0.4505
R31655 VDD.n890 VDD.n889 0.4505
R31656 VDD.n891 VDD.n882 0.4505
R31657 VDD.n893 VDD.n892 0.4505
R31658 VDD.n561 VDD.n559 0.4505
R31659 VDD.n898 VDD.n897 0.4505
R31660 VDD.n560 VDD.n558 0.4505
R31661 VDD.n878 VDD.n877 0.4505
R31662 VDD.n876 VDD.n563 0.4505
R31663 VDD.n875 VDD.n874 0.4505
R31664 VDD.n565 VDD.n564 0.4505
R31665 VDD.n870 VDD.n869 0.4505
R31666 VDD.n868 VDD.n567 0.4505
R31667 VDD.n867 VDD.n866 0.4505
R31668 VDD.n569 VDD.n568 0.4505
R31669 VDD.n862 VDD.n861 0.4505
R31670 VDD.n860 VDD.n571 0.4505
R31671 VDD.n859 VDD.n858 0.4505
R31672 VDD.n573 VDD.n572 0.4505
R31673 VDD.n854 VDD.n853 0.4505
R31674 VDD.n852 VDD.n575 0.4505
R31675 VDD.n851 VDD.n850 0.4505
R31676 VDD.n577 VDD.n576 0.4505
R31677 VDD.n846 VDD.n845 0.4505
R31678 VDD.n844 VDD.n579 0.4505
R31679 VDD.n843 VDD.n842 0.4505
R31680 VDD.n581 VDD.n580 0.4505
R31681 VDD.n838 VDD.n837 0.4505
R31682 VDD.n836 VDD.n583 0.4505
R31683 VDD.n761 VDD.n584 0.4505
R31684 VDD.n763 VDD.n762 0.4505
R31685 VDD.n765 VDD.n764 0.4505
R31686 VDD.n757 VDD.n756 0.4505
R31687 VDD.n770 VDD.n769 0.4505
R31688 VDD.n771 VDD.n755 0.4505
R31689 VDD.n773 VDD.n772 0.4505
R31690 VDD.n775 VDD.n774 0.4505
R31691 VDD.n753 VDD.n752 0.4505
R31692 VDD.n780 VDD.n779 0.4505
R31693 VDD.n781 VDD.n751 0.4505
R31694 VDD.n783 VDD.n782 0.4505
R31695 VDD.n590 VDD.n588 0.4505
R31696 VDD.n788 VDD.n787 0.4505
R31697 VDD.n589 VDD.n587 0.4505
R31698 VDD.n747 VDD.n746 0.4505
R31699 VDD.n745 VDD.n592 0.4505
R31700 VDD.n744 VDD.n743 0.4505
R31701 VDD.n594 VDD.n593 0.4505
R31702 VDD.n739 VDD.n738 0.4505
R31703 VDD.n737 VDD.n596 0.4505
R31704 VDD.n736 VDD.n735 0.4505
R31705 VDD.n598 VDD.n597 0.4505
R31706 VDD.n731 VDD.n730 0.4505
R31707 VDD.n729 VDD.n600 0.4505
R31708 VDD.n728 VDD.n727 0.4505
R31709 VDD.n602 VDD.n601 0.4505
R31710 VDD.n723 VDD.n722 0.4505
R31711 VDD.n721 VDD.n604 0.4505
R31712 VDD.n720 VDD.n719 0.4505
R31713 VDD.n606 VDD.n605 0.4505
R31714 VDD.n715 VDD.n714 0.4505
R31715 VDD.n713 VDD.n608 0.4505
R31716 VDD.n712 VDD.n711 0.4505
R31717 VDD.n610 VDD.n609 0.4505
R31718 VDD.n707 VDD.n706 0.4505
R31719 VDD.n705 VDD.n612 0.4505
R31720 VDD.n680 VDD.n613 0.4505
R31721 VDD.n683 VDD.n681 0.4505
R31722 VDD.n685 VDD.n684 0.4505
R31723 VDD.n682 VDD.n677 0.4505
R31724 VDD.n689 VDD.n676 0.4505
R31725 VDD.n691 VDD.n690 0.4505
R31726 VDD.n114 VDD.n113 0.424611
R31727 VDD.n399 VDD.n398 0.406952
R31728 VDD.n695 VDD.n694 0.39425
R31729 VDD.n696 VDD.n695 0.39425
R31730 VDD.n321 VDD.n319 0.341837
R31731 VDD.n195 VDD.n194 0.310206
R31732 VDD.n902 VDD.n557 0.296971
R31733 VDD.n832 VDD.n585 0.296971
R31734 VDD.n826 VDD.n791 0.296971
R31735 VDD.n81 VDD.n80 0.290353
R31736 VDD.n701 VDD.n700 0.277118
R31737 VDD.n333 VDD.n313 0.273147
R31738 VDD.n181 VDD.n180 0.273
R31739 VDD.n701 VDD.n614 0.269176
R31740 VDD.n108 VDD.n107 0.264579
R31741 VDD.n109 VDD.n108 0.255105
R31742 VDD VDD.n903 0.250647
R31743 VDD.n825 VDD 0.250647
R31744 VDD.n831 VDD 0.250647
R31745 VDD.n903 VDD.n902 0.249324
R31746 VDD.n832 VDD.n831 0.249324
R31747 VDD.n826 VDD.n825 0.249324
R31748 VDD.n699 VDD.n698 0.241382
R31749 VDD.n102 VDD.n101 0.240059
R31750 VDD.n550 VDD.n549 0.231338
R31751 VDD.n923 VDD.n922 0.231338
R31752 VDD VDD.n393 0.226824
R31753 VDD.n158 VDD.n18 0.22175
R31754 VDD.n93 VDD.n88 0.212524
R31755 VDD.n97 VDD.n87 0.212524
R31756 VDD.n104 VDD.n100 0.212524
R31757 VDD.n333 VDD.n332 0.208294
R31758 VDD.n398 VDD.n397 0.196382
R31759 VDD.n90 VDD.n89 0.195059
R31760 VDD.n91 VDD.n90 0.184471
R31761 VDD.n335 VDD.n313 0.181824
R31762 VDD.n180 VDD.n29 0.176791
R31763 VDD.n135 VDD.n134 0.165582
R31764 VDD.n815 VDD.n800 0.1505
R31765 VDD.n817 VDD.n816 0.1505
R31766 VDD.n811 VDD.n810 0.1505
R31767 VDD.n201 VDD.n200 0.149225
R31768 VDD.n79 VDD 0.1455
R31769 VDD.n74 VDD 0.1455
R31770 VDD.n173 VDD 0.1455
R31771 VDD VDD.n170 0.1455
R31772 VDD.n179 VDD 0.1455
R31773 VDD.n146 VDD 0.1455
R31774 VDD.n149 VDD.n147 0.1455
R31775 VDD VDD.n149 0.1455
R31776 VDD.n150 VDD 0.1455
R31777 VDD.n152 VDD.n150 0.1455
R31778 VDD VDD.n25 0.1455
R31779 VDD.n182 VDD 0.1455
R31780 VDD.n182 VDD.n181 0.1455
R31781 VDD.n158 VDD.n157 0.1455
R31782 VDD.n157 VDD 0.1455
R31783 VDD.n153 VDD 0.1455
R31784 VDD.n53 VDD.n48 0.1455
R31785 VDD VDD.n48 0.1455
R31786 VDD.n120 VDD 0.1455
R31787 VDD.n121 VDD.n120 0.1455
R31788 VDD.n126 VDD 0.1455
R31789 VDD VDD.n125 0.1455
R31790 VDD.n57 VDD 0.1455
R31791 VDD VDD.n56 0.1455
R31792 VDD VDD.n39 0.1455
R31793 VDD.n72 VDD 0.1455
R31794 VDD VDD.n632 0.1455
R31795 VDD.n640 VDD 0.1455
R31796 VDD.n647 VDD 0.1455
R31797 VDD VDD.n633 0.1455
R31798 VDD VDD.n625 0.1455
R31799 VDD.n657 VDD 0.1455
R31800 VDD.n648 VDD.n626 0.1455
R31801 VDD VDD.n626 0.1455
R31802 VDD.n666 VDD 0.1455
R31803 VDD.n667 VDD.n666 0.1455
R31804 VDD.n642 VDD.n641 0.1455
R31805 VDD.n641 VDD 0.1455
R31806 VDD VDD.n616 0.1455
R31807 VDD.n655 VDD.n654 0.1455
R31808 VDD VDD.n655 0.1455
R31809 VDD VDD.n663 0.1455
R31810 VDD.n663 VDD.n662 0.1455
R31811 VDD.n661 VDD 0.1455
R31812 VDD VDD.n615 0.143658
R31813 VDD.n700 VDD 0.138147
R31814 VDD.n319 VDD 0.1355
R31815 VDD.n330 VDD.n315 0.128395
R31816 VDD.n397 VDD.n396 0.127559
R31817 VDD.n906 VDD.n905 0.1238
R31818 VDD.n398 VDD 0.123588
R31819 VDD.n822 VDD.n793 0.1235
R31820 VDD.n92 VDD.n91 0.113
R31821 VDD.n89 VDD.n86 0.113
R31822 VDD.n101 VDD.n99 0.113
R31823 VDD.n387 VDD.n295 0.107781
R31824 VDD.n170 VDD 0.107483
R31825 VDD VDD.n179 0.107483
R31826 VDD.n817 VDD.n799 0.1055
R31827 VDD.n810 VDD.n809 0.1055
R31828 VDD.n806 VDD.n800 0.1055
R31829 VDD.n114 VDD.n79 0.1005
R31830 VDD.n74 VDD.n73 0.1005
R31831 VDD.n173 VDD.n136 0.1005
R31832 VDD.n147 VDD.n146 0.1005
R31833 VDD.n189 VDD.n25 0.1005
R31834 VDD.n153 VDD.n152 0.1005
R31835 VDD.n126 VDD.n47 0.1005
R31836 VDD.n125 VDD.n121 0.1005
R31837 VDD.n57 VDD.n47 0.1005
R31838 VDD.n56 VDD.n53 0.1005
R31839 VDD.n134 VDD.n39 0.1005
R31840 VDD.n73 VDD.n72 0.1005
R31841 VDD.n654 VDD.n632 0.1005
R31842 VDD.n642 VDD.n640 0.1005
R31843 VDD.n648 VDD.n647 0.1005
R31844 VDD.n654 VDD.n633 0.1005
R31845 VDD.n667 VDD.n625 0.1005
R31846 VDD.n662 VDD.n657 0.1005
R31847 VDD.n673 VDD.n616 0.1005
R31848 VDD.n662 VDD.n661 0.1005
R31849 VDD.n189 VDD.n20 0.091309
R31850 VDD.n383 VDD.n295 0.0895132
R31851 VDD.n111 VDD.n81 0.0891765
R31852 VDD.n202 VDD.n18 0.0840281
R31853 VDD.n799 VDD 0.0755
R31854 VDD VDD.n815 0.0755
R31855 VDD.n816 VDD 0.0755
R31856 VDD.n809 VDD 0.0755
R31857 VDD.n806 VDD 0.0755
R31858 VDD.n811 VDD 0.0755
R31859 VDD VDD.n793 0.0755
R31860 VDD.n674 VDD.n615 0.0739211
R31861 VDD.n692 VDD.n675 0.0704044
R31862 VDD.n674 VDD.n673 0.0644474
R31863 VDD.n698 VDD 0.0627059
R31864 VDD VDD.n699 0.0627059
R31865 VDD.n688 VDD.n675 0.0582093
R31866 VDD.n180 VDD.n18 0.05175
R31867 VDD.n822 VDD 0.0455
R31868 VDD.n180 VDD 0.0427845
R31869 VDD.n180 VDD 0.0427845
R31870 VDD.n904 VDD 0.0402059
R31871 VDD.n830 VDD 0.0402059
R31872 VDD VDD.n830 0.0402059
R31873 VDD.n324 VDD.n323 0.037532
R31874 VDD VDD.n29 0.0371045
R31875 VDD VDD.n29 0.0371045
R31876 VDD VDD.n320 0.0322201
R31877 VDD.n325 VDD.n324 0.0284258
R31878 VDD.n690 VDD.n675 0.026721
R31879 VDD.n16 VDD.n15 0.0255787
R31880 VDD.n320 VDD.n317 0.0253904
R31881 VDD.n115 VDD.n114 0.0239607
R31882 VDD.n115 VDD 0.0239607
R31883 VDD VDD.n40 0.0239607
R31884 VDD.n134 VDD.n40 0.0239607
R31885 VDD.n168 VDD.n136 0.0239607
R31886 VDD.n168 VDD 0.0239607
R31887 VDD VDD.n24 0.0239607
R31888 VDD.n136 VDD.n135 0.0220168
R31889 VDD.n102 VDD 0.0216765
R31890 VDD.n80 VDD 0.0216765
R31891 VDD.n197 VDD.n195 0.0203202
R31892 VDD.n217 VDD.n209 0.0169185
R31893 VDD.n208 VDD.n13 0.0169185
R31894 VDD.n216 VDD.n211 0.0169185
R31895 VDD.n210 VDD.n12 0.0169185
R31896 VDD.n215 VDD.n213 0.0169185
R31897 VDD.n212 VDD.n11 0.0169185
R31898 VDD.n554 VDD.n552 0.0169185
R31899 VDD.n553 VDD.n10 0.0169185
R31900 VDD.n556 VDD.n7 0.0169185
R31901 VDD.n913 VDD.n908 0.0169185
R31902 VDD.n924 VDD.n908 0.0169185
R31903 VDD.n914 VDD.n909 0.0169185
R31904 VDD.n925 VDD.n909 0.0169185
R31905 VDD.n915 VDD.n910 0.0169185
R31906 VDD.n926 VDD.n910 0.0169185
R31907 VDD.n916 VDD.n911 0.0169185
R31908 VDD.n927 VDD.n911 0.0169185
R31909 VDD.n929 VDD.n912 0.0169185
R31910 VDD.n217 VDD.n206 0.0169185
R31911 VDD.n209 VDD.n208 0.0169185
R31912 VDD.n216 VDD.n13 0.0169185
R31913 VDD.n211 VDD.n210 0.0169185
R31914 VDD.n215 VDD.n12 0.0169185
R31915 VDD.n213 VDD.n212 0.0169185
R31916 VDD.n552 VDD.n11 0.0169185
R31917 VDD.n554 VDD.n553 0.0169185
R31918 VDD.n10 VDD.n7 0.0169185
R31919 VDD.n913 VDD.n906 0.0169185
R31920 VDD.n924 VDD.n6 0.0169185
R31921 VDD.n914 VDD.n6 0.0169185
R31922 VDD.n925 VDD.n5 0.0169185
R31923 VDD.n915 VDD.n5 0.0169185
R31924 VDD.n926 VDD.n4 0.0169185
R31925 VDD.n916 VDD.n4 0.0169185
R31926 VDD.n927 VDD.n3 0.0169185
R31927 VDD.n912 VDD.n3 0.0169185
R31928 VDD.n329 VDD.n327 0.0168912
R31929 VDD.n385 VDD.n295 0.0166957
R31930 VDD.n190 VDD.n24 0.0154663
R31931 VDD.n198 VDD.n21 0.0149069
R31932 VDD.n199 VDD.n198 0.0149069
R31933 VDD.n203 VDD.n17 0.0149069
R31934 VDD.n204 VDD.n203 0.0149069
R31935 VDD.n196 VDD.n21 0.0149069
R31936 VDD.n200 VDD.n199 0.0149069
R31937 VDD.n201 VDD.n17 0.0149069
R31938 VDD.n205 VDD.n204 0.0149069
R31939 VDD.n16 VDD.n14 0.0135045
R31940 VDD.n197 VDD.n19 0.0135045
R31941 VDD.n202 VDD.n14 0.0135045
R31942 VDD.n323 VDD.n317 0.0126417
R31943 VDD.n385 VDD.n384 0.00962857
R31944 VDD.n384 VDD.n297 0.00962857
R31945 VDD.n380 VDD.n297 0.00962857
R31946 VDD.n380 VDD.n299 0.00962857
R31947 VDD.n376 VDD.n299 0.00962857
R31948 VDD.n376 VDD.n302 0.00962857
R31949 VDD.n372 VDD.n302 0.00962857
R31950 VDD.n372 VDD.n304 0.00962857
R31951 VDD.n368 VDD.n304 0.00962857
R31952 VDD.n368 VDD.n306 0.00962857
R31953 VDD.n364 VDD.n306 0.00962857
R31954 VDD.n364 VDD.n308 0.00962857
R31955 VDD.n360 VDD.n308 0.00962857
R31956 VDD.n360 VDD.n310 0.00962857
R31957 VDD.n356 VDD.n310 0.00962857
R31958 VDD.n356 VDD.n312 0.00962857
R31959 VDD.n351 VDD.n312 0.00962857
R31960 VDD.n351 VDD.n338 0.00962857
R31961 VDD.n347 VDD.n338 0.00962857
R31962 VDD.n347 VDD.n340 0.00962857
R31963 VDD.n343 VDD.n340 0.00962857
R31964 VDD.n343 VDD.n292 0.00962857
R31965 VDD.n403 VDD.n292 0.00962857
R31966 VDD.n403 VDD.n290 0.00962857
R31967 VDD.n407 VDD.n290 0.00962857
R31968 VDD.n407 VDD.n288 0.00962857
R31969 VDD.n411 VDD.n288 0.00962857
R31970 VDD.n411 VDD.n286 0.00962857
R31971 VDD.n415 VDD.n286 0.00962857
R31972 VDD.n415 VDD.n284 0.00962857
R31973 VDD.n419 VDD.n284 0.00962857
R31974 VDD.n419 VDD.n282 0.00962857
R31975 VDD.n423 VDD.n282 0.00962857
R31976 VDD.n423 VDD.n280 0.00962857
R31977 VDD.n427 VDD.n280 0.00962857
R31978 VDD.n427 VDD.n278 0.00962857
R31979 VDD.n431 VDD.n278 0.00962857
R31980 VDD.n431 VDD.n276 0.00962857
R31981 VDD.n435 VDD.n276 0.00962857
R31982 VDD.n435 VDD.n274 0.00962857
R31983 VDD.n439 VDD.n274 0.00962857
R31984 VDD.n439 VDD.n272 0.00962857
R31985 VDD.n443 VDD.n272 0.00962857
R31986 VDD.n443 VDD.n270 0.00962857
R31987 VDD.n447 VDD.n270 0.00962857
R31988 VDD.n447 VDD.n268 0.00962857
R31989 VDD.n451 VDD.n268 0.00962857
R31990 VDD.n451 VDD.n266 0.00962857
R31991 VDD.n455 VDD.n266 0.00962857
R31992 VDD.n455 VDD.n264 0.00962857
R31993 VDD.n459 VDD.n264 0.00962857
R31994 VDD.n459 VDD.n262 0.00962857
R31995 VDD.n463 VDD.n262 0.00962857
R31996 VDD.n463 VDD.n260 0.00962857
R31997 VDD.n467 VDD.n260 0.00962857
R31998 VDD.n467 VDD.n258 0.00962857
R31999 VDD.n471 VDD.n258 0.00962857
R32000 VDD.n471 VDD.n256 0.00962857
R32001 VDD.n475 VDD.n256 0.00962857
R32002 VDD.n475 VDD.n254 0.00962857
R32003 VDD.n479 VDD.n254 0.00962857
R32004 VDD.n479 VDD.n252 0.00962857
R32005 VDD.n483 VDD.n252 0.00962857
R32006 VDD.n483 VDD.n250 0.00962857
R32007 VDD.n487 VDD.n250 0.00962857
R32008 VDD.n487 VDD.n248 0.00962857
R32009 VDD.n491 VDD.n248 0.00962857
R32010 VDD.n491 VDD.n246 0.00962857
R32011 VDD.n495 VDD.n246 0.00962857
R32012 VDD.n495 VDD.n244 0.00962857
R32013 VDD.n499 VDD.n244 0.00962857
R32014 VDD.n499 VDD.n242 0.00962857
R32015 VDD.n503 VDD.n242 0.00962857
R32016 VDD.n503 VDD.n240 0.00962857
R32017 VDD.n507 VDD.n240 0.00962857
R32018 VDD.n507 VDD.n238 0.00962857
R32019 VDD.n511 VDD.n238 0.00962857
R32020 VDD.n511 VDD.n236 0.00962857
R32021 VDD.n515 VDD.n236 0.00962857
R32022 VDD.n515 VDD.n234 0.00962857
R32023 VDD.n519 VDD.n234 0.00962857
R32024 VDD.n519 VDD.n232 0.00962857
R32025 VDD.n523 VDD.n232 0.00962857
R32026 VDD.n523 VDD.n230 0.00962857
R32027 VDD.n527 VDD.n230 0.00962857
R32028 VDD.n527 VDD.n228 0.00962857
R32029 VDD.n531 VDD.n228 0.00962857
R32030 VDD.n531 VDD.n226 0.00962857
R32031 VDD.n535 VDD.n226 0.00962857
R32032 VDD.n535 VDD.n224 0.00962857
R32033 VDD.n539 VDD.n224 0.00962857
R32034 VDD.n539 VDD.n222 0.00962857
R32035 VDD.n543 VDD.n222 0.00962857
R32036 VDD.n547 VDD.n546 0.00962857
R32037 VDD.n548 VDD.n547 0.00962857
R32038 VDD.n548 VDD.n218 0.00962857
R32039 VDD.n386 VDD.n296 0.00962857
R32040 VDD.n300 VDD.n296 0.00962857
R32041 VDD.n379 VDD.n300 0.00962857
R32042 VDD.n379 VDD.n378 0.00962857
R32043 VDD.n378 VDD.n377 0.00962857
R32044 VDD.n377 VDD.n301 0.00962857
R32045 VDD.n371 VDD.n301 0.00962857
R32046 VDD.n371 VDD.n370 0.00962857
R32047 VDD.n370 VDD.n369 0.00962857
R32048 VDD.n369 VDD.n305 0.00962857
R32049 VDD.n363 VDD.n305 0.00962857
R32050 VDD.n363 VDD.n362 0.00962857
R32051 VDD.n362 VDD.n361 0.00962857
R32052 VDD.n361 VDD.n309 0.00962857
R32053 VDD.n355 VDD.n309 0.00962857
R32054 VDD.n355 VDD.n354 0.00962857
R32055 VDD.n346 VDD.n341 0.00962857
R32056 VDD.n346 VDD.n345 0.00962857
R32057 VDD.n345 VDD.n344 0.00962857
R32058 VDD.n344 VDD.n293 0.00962857
R32059 VDD.n402 VDD.n289 0.00962857
R32060 VDD.n408 VDD.n289 0.00962857
R32061 VDD.n409 VDD.n408 0.00962857
R32062 VDD.n410 VDD.n409 0.00962857
R32063 VDD.n410 VDD.n285 0.00962857
R32064 VDD.n416 VDD.n285 0.00962857
R32065 VDD.n417 VDD.n416 0.00962857
R32066 VDD.n418 VDD.n417 0.00962857
R32067 VDD.n418 VDD.n281 0.00962857
R32068 VDD.n424 VDD.n281 0.00962857
R32069 VDD.n425 VDD.n424 0.00962857
R32070 VDD.n426 VDD.n425 0.00962857
R32071 VDD.n426 VDD.n277 0.00962857
R32072 VDD.n432 VDD.n277 0.00962857
R32073 VDD.n433 VDD.n432 0.00962857
R32074 VDD.n434 VDD.n433 0.00962857
R32075 VDD.n434 VDD.n273 0.00962857
R32076 VDD.n440 VDD.n273 0.00962857
R32077 VDD.n441 VDD.n440 0.00962857
R32078 VDD.n442 VDD.n441 0.00962857
R32079 VDD.n442 VDD.n269 0.00962857
R32080 VDD.n448 VDD.n269 0.00962857
R32081 VDD.n449 VDD.n448 0.00962857
R32082 VDD.n450 VDD.n449 0.00962857
R32083 VDD.n450 VDD.n265 0.00962857
R32084 VDD.n456 VDD.n265 0.00962857
R32085 VDD.n457 VDD.n456 0.00962857
R32086 VDD.n458 VDD.n457 0.00962857
R32087 VDD.n458 VDD.n261 0.00962857
R32088 VDD.n464 VDD.n261 0.00962857
R32089 VDD.n465 VDD.n464 0.00962857
R32090 VDD.n466 VDD.n465 0.00962857
R32091 VDD.n466 VDD.n257 0.00962857
R32092 VDD.n472 VDD.n257 0.00962857
R32093 VDD.n473 VDD.n472 0.00962857
R32094 VDD.n474 VDD.n473 0.00962857
R32095 VDD.n474 VDD.n253 0.00962857
R32096 VDD.n480 VDD.n253 0.00962857
R32097 VDD.n481 VDD.n480 0.00962857
R32098 VDD.n482 VDD.n481 0.00962857
R32099 VDD.n482 VDD.n249 0.00962857
R32100 VDD.n488 VDD.n249 0.00962857
R32101 VDD.n489 VDD.n488 0.00962857
R32102 VDD.n490 VDD.n489 0.00962857
R32103 VDD.n490 VDD.n245 0.00962857
R32104 VDD.n496 VDD.n245 0.00962857
R32105 VDD.n497 VDD.n496 0.00962857
R32106 VDD.n498 VDD.n497 0.00962857
R32107 VDD.n498 VDD.n241 0.00962857
R32108 VDD.n504 VDD.n241 0.00962857
R32109 VDD.n505 VDD.n504 0.00962857
R32110 VDD.n506 VDD.n505 0.00962857
R32111 VDD.n506 VDD.n237 0.00962857
R32112 VDD.n512 VDD.n237 0.00962857
R32113 VDD.n513 VDD.n512 0.00962857
R32114 VDD.n514 VDD.n513 0.00962857
R32115 VDD.n514 VDD.n233 0.00962857
R32116 VDD.n520 VDD.n233 0.00962857
R32117 VDD.n521 VDD.n520 0.00962857
R32118 VDD.n522 VDD.n521 0.00962857
R32119 VDD.n522 VDD.n229 0.00962857
R32120 VDD.n528 VDD.n229 0.00962857
R32121 VDD.n529 VDD.n528 0.00962857
R32122 VDD.n530 VDD.n529 0.00962857
R32123 VDD.n530 VDD.n225 0.00962857
R32124 VDD.n536 VDD.n225 0.00962857
R32125 VDD.n537 VDD.n536 0.00962857
R32126 VDD.n538 VDD.n537 0.00962857
R32127 VDD.n538 VDD.n221 0.00962857
R32128 VDD.n544 VDD.n221 0.00962857
R32129 VDD.n545 VDD.n9 0.00962857
R32130 VDD.n690 VDD.n689 0.00962857
R32131 VDD.n689 VDD.n677 0.00962857
R32132 VDD.n685 VDD.n677 0.00962857
R32133 VDD.n685 VDD.n681 0.00962857
R32134 VDD.n681 VDD.n680 0.00962857
R32135 VDD.n680 VDD.n612 0.00962857
R32136 VDD.n707 VDD.n612 0.00962857
R32137 VDD.n707 VDD.n610 0.00962857
R32138 VDD.n711 VDD.n610 0.00962857
R32139 VDD.n711 VDD.n608 0.00962857
R32140 VDD.n715 VDD.n608 0.00962857
R32141 VDD.n715 VDD.n606 0.00962857
R32142 VDD.n719 VDD.n606 0.00962857
R32143 VDD.n719 VDD.n604 0.00962857
R32144 VDD.n723 VDD.n604 0.00962857
R32145 VDD.n723 VDD.n602 0.00962857
R32146 VDD.n727 VDD.n602 0.00962857
R32147 VDD.n727 VDD.n600 0.00962857
R32148 VDD.n731 VDD.n600 0.00962857
R32149 VDD.n731 VDD.n598 0.00962857
R32150 VDD.n735 VDD.n598 0.00962857
R32151 VDD.n735 VDD.n596 0.00962857
R32152 VDD.n739 VDD.n596 0.00962857
R32153 VDD.n739 VDD.n594 0.00962857
R32154 VDD.n743 VDD.n594 0.00962857
R32155 VDD.n743 VDD.n592 0.00962857
R32156 VDD.n747 VDD.n592 0.00962857
R32157 VDD.n747 VDD.n589 0.00962857
R32158 VDD.n787 VDD.n589 0.00962857
R32159 VDD.n787 VDD.n590 0.00962857
R32160 VDD.n783 VDD.n590 0.00962857
R32161 VDD.n783 VDD.n751 0.00962857
R32162 VDD.n779 VDD.n751 0.00962857
R32163 VDD.n779 VDD.n753 0.00962857
R32164 VDD.n775 VDD.n753 0.00962857
R32165 VDD.n775 VDD.n773 0.00962857
R32166 VDD.n773 VDD.n755 0.00962857
R32167 VDD.n769 VDD.n755 0.00962857
R32168 VDD.n769 VDD.n757 0.00962857
R32169 VDD.n765 VDD.n757 0.00962857
R32170 VDD.n765 VDD.n762 0.00962857
R32171 VDD.n762 VDD.n761 0.00962857
R32172 VDD.n761 VDD.n583 0.00962857
R32173 VDD.n838 VDD.n583 0.00962857
R32174 VDD.n838 VDD.n581 0.00962857
R32175 VDD.n842 VDD.n581 0.00962857
R32176 VDD.n842 VDD.n579 0.00962857
R32177 VDD.n846 VDD.n579 0.00962857
R32178 VDD.n846 VDD.n577 0.00962857
R32179 VDD.n850 VDD.n577 0.00962857
R32180 VDD.n850 VDD.n575 0.00962857
R32181 VDD.n854 VDD.n575 0.00962857
R32182 VDD.n854 VDD.n573 0.00962857
R32183 VDD.n858 VDD.n573 0.00962857
R32184 VDD.n858 VDD.n571 0.00962857
R32185 VDD.n862 VDD.n571 0.00962857
R32186 VDD.n862 VDD.n569 0.00962857
R32187 VDD.n866 VDD.n569 0.00962857
R32188 VDD.n866 VDD.n567 0.00962857
R32189 VDD.n870 VDD.n567 0.00962857
R32190 VDD.n870 VDD.n565 0.00962857
R32191 VDD.n874 VDD.n565 0.00962857
R32192 VDD.n874 VDD.n563 0.00962857
R32193 VDD.n878 VDD.n563 0.00962857
R32194 VDD.n878 VDD.n560 0.00962857
R32195 VDD.n897 VDD.n560 0.00962857
R32196 VDD.n897 VDD.n561 0.00962857
R32197 VDD.n893 VDD.n561 0.00962857
R32198 VDD.n893 VDD.n882 0.00962857
R32199 VDD.n889 VDD.n882 0.00962857
R32200 VDD.n889 VDD.n885 0.00962857
R32201 VDD.n885 VDD.n0 0.00962857
R32202 VDD.n933 VDD.n1 0.00962857
R32203 VDD.n921 VDD.n1 0.00962857
R32204 VDD.n921 VDD.n919 0.00962857
R32205 VDD.n691 VDD.n676 0.00962857
R32206 VDD.n682 VDD.n676 0.00962857
R32207 VDD.n684 VDD.n682 0.00962857
R32208 VDD.n684 VDD.n683 0.00962857
R32209 VDD.n683 VDD.n613 0.00962857
R32210 VDD.n706 VDD.n705 0.00962857
R32211 VDD.n706 VDD.n609 0.00962857
R32212 VDD.n712 VDD.n609 0.00962857
R32213 VDD.n713 VDD.n712 0.00962857
R32214 VDD.n714 VDD.n713 0.00962857
R32215 VDD.n714 VDD.n605 0.00962857
R32216 VDD.n720 VDD.n605 0.00962857
R32217 VDD.n721 VDD.n720 0.00962857
R32218 VDD.n722 VDD.n721 0.00962857
R32219 VDD.n722 VDD.n601 0.00962857
R32220 VDD.n728 VDD.n601 0.00962857
R32221 VDD.n729 VDD.n728 0.00962857
R32222 VDD.n730 VDD.n729 0.00962857
R32223 VDD.n730 VDD.n597 0.00962857
R32224 VDD.n736 VDD.n597 0.00962857
R32225 VDD.n737 VDD.n736 0.00962857
R32226 VDD.n738 VDD.n737 0.00962857
R32227 VDD.n738 VDD.n593 0.00962857
R32228 VDD.n744 VDD.n593 0.00962857
R32229 VDD.n745 VDD.n744 0.00962857
R32230 VDD.n746 VDD.n745 0.00962857
R32231 VDD.n746 VDD.n587 0.00962857
R32232 VDD.n788 VDD.n588 0.00962857
R32233 VDD.n782 VDD.n588 0.00962857
R32234 VDD.n782 VDD.n781 0.00962857
R32235 VDD.n781 VDD.n780 0.00962857
R32236 VDD.n780 VDD.n752 0.00962857
R32237 VDD.n774 VDD.n752 0.00962857
R32238 VDD.n772 VDD.n771 0.00962857
R32239 VDD.n771 VDD.n770 0.00962857
R32240 VDD.n770 VDD.n756 0.00962857
R32241 VDD.n764 VDD.n756 0.00962857
R32242 VDD.n764 VDD.n763 0.00962857
R32243 VDD.n763 VDD.n584 0.00962857
R32244 VDD.n837 VDD.n836 0.00962857
R32245 VDD.n837 VDD.n580 0.00962857
R32246 VDD.n843 VDD.n580 0.00962857
R32247 VDD.n844 VDD.n843 0.00962857
R32248 VDD.n845 VDD.n844 0.00962857
R32249 VDD.n845 VDD.n576 0.00962857
R32250 VDD.n851 VDD.n576 0.00962857
R32251 VDD.n852 VDD.n851 0.00962857
R32252 VDD.n853 VDD.n852 0.00962857
R32253 VDD.n853 VDD.n572 0.00962857
R32254 VDD.n859 VDD.n572 0.00962857
R32255 VDD.n860 VDD.n859 0.00962857
R32256 VDD.n861 VDD.n860 0.00962857
R32257 VDD.n861 VDD.n568 0.00962857
R32258 VDD.n867 VDD.n568 0.00962857
R32259 VDD.n868 VDD.n867 0.00962857
R32260 VDD.n869 VDD.n868 0.00962857
R32261 VDD.n869 VDD.n564 0.00962857
R32262 VDD.n875 VDD.n564 0.00962857
R32263 VDD.n876 VDD.n875 0.00962857
R32264 VDD.n877 VDD.n876 0.00962857
R32265 VDD.n877 VDD.n558 0.00962857
R32266 VDD.n898 VDD.n559 0.00962857
R32267 VDD.n892 VDD.n559 0.00962857
R32268 VDD.n892 VDD.n891 0.00962857
R32269 VDD.n891 VDD.n890 0.00962857
R32270 VDD.n890 VDD.n884 0.00962857
R32271 VDD.n884 VDD.n883 0.00962857
R32272 VDD.n932 VDD.n931 0.00962857
R32273 VDD.n354 VDD.n353 0.00956429
R32274 VDD.n332 VDD.n331 0.00915093
R32275 VDD.n190 VDD.n189 0.00899438
R32276 VDD.n326 VDD.n325 0.00884739
R32277 VDD.n789 VDD.n587 0.0086
R32278 VDD.n387 VDD.n386 0.00853571
R32279 VDD.n555 VDD.n9 0.00827857
R32280 VDD.n207 VDD.n8 0.00827857
R32281 VDD.n551 VDD.n214 0.00827857
R32282 VDD.n931 VDD.n930 0.00827857
R32283 VDD.n917 VDD.n907 0.00827857
R32284 VDD.n928 VDD.n918 0.00827857
R32285 VDD.n899 VDD.n558 0.00795714
R32286 VDD.n543 VDD 0.00782857
R32287 VDD VDD.n544 0.00782857
R32288 VDD VDD.n0 0.00782857
R32289 VDD.n883 VDD 0.00782857
R32290 VDD.n352 VDD.n337 0.00763571
R32291 VDD.n401 VDD.n293 0.00692857
R32292 VDD.n774 VDD.n586 0.0068
R32293 VDD.n383 VDD.n382 0.00658571
R32294 VDD.n382 VDD.n381 0.00658571
R32295 VDD.n381 VDD.n298 0.00658571
R32296 VDD.n375 VDD.n298 0.00658571
R32297 VDD.n375 VDD.n374 0.00658571
R32298 VDD.n374 VDD.n373 0.00658571
R32299 VDD.n373 VDD.n303 0.00658571
R32300 VDD.n367 VDD.n303 0.00658571
R32301 VDD.n367 VDD.n366 0.00658571
R32302 VDD.n366 VDD.n365 0.00658571
R32303 VDD.n365 VDD.n307 0.00658571
R32304 VDD.n359 VDD.n307 0.00658571
R32305 VDD.n359 VDD.n358 0.00658571
R32306 VDD.n358 VDD.n357 0.00658571
R32307 VDD.n357 VDD.n311 0.00658571
R32308 VDD.n350 VDD.n311 0.00658571
R32309 VDD.n350 VDD.n349 0.00658571
R32310 VDD.n349 VDD.n348 0.00658571
R32311 VDD.n348 VDD.n339 0.00658571
R32312 VDD.n342 VDD.n339 0.00658571
R32313 VDD.n342 VDD.n291 0.00658571
R32314 VDD.n404 VDD.n291 0.00658571
R32315 VDD.n405 VDD.n404 0.00658571
R32316 VDD.n406 VDD.n405 0.00658571
R32317 VDD.n406 VDD.n287 0.00658571
R32318 VDD.n412 VDD.n287 0.00658571
R32319 VDD.n413 VDD.n412 0.00658571
R32320 VDD.n414 VDD.n413 0.00658571
R32321 VDD.n414 VDD.n283 0.00658571
R32322 VDD.n420 VDD.n283 0.00658571
R32323 VDD.n421 VDD.n420 0.00658571
R32324 VDD.n422 VDD.n421 0.00658571
R32325 VDD.n422 VDD.n279 0.00658571
R32326 VDD.n428 VDD.n279 0.00658571
R32327 VDD.n429 VDD.n428 0.00658571
R32328 VDD.n430 VDD.n429 0.00658571
R32329 VDD.n430 VDD.n275 0.00658571
R32330 VDD.n436 VDD.n275 0.00658571
R32331 VDD.n437 VDD.n436 0.00658571
R32332 VDD.n438 VDD.n437 0.00658571
R32333 VDD.n438 VDD.n271 0.00658571
R32334 VDD.n444 VDD.n271 0.00658571
R32335 VDD.n445 VDD.n444 0.00658571
R32336 VDD.n446 VDD.n445 0.00658571
R32337 VDD.n446 VDD.n267 0.00658571
R32338 VDD.n452 VDD.n267 0.00658571
R32339 VDD.n453 VDD.n452 0.00658571
R32340 VDD.n454 VDD.n453 0.00658571
R32341 VDD.n454 VDD.n263 0.00658571
R32342 VDD.n460 VDD.n263 0.00658571
R32343 VDD.n461 VDD.n460 0.00658571
R32344 VDD.n462 VDD.n461 0.00658571
R32345 VDD.n462 VDD.n259 0.00658571
R32346 VDD.n468 VDD.n259 0.00658571
R32347 VDD.n469 VDD.n468 0.00658571
R32348 VDD.n470 VDD.n469 0.00658571
R32349 VDD.n470 VDD.n255 0.00658571
R32350 VDD.n476 VDD.n255 0.00658571
R32351 VDD.n477 VDD.n476 0.00658571
R32352 VDD.n478 VDD.n477 0.00658571
R32353 VDD.n478 VDD.n251 0.00658571
R32354 VDD.n484 VDD.n251 0.00658571
R32355 VDD.n485 VDD.n484 0.00658571
R32356 VDD.n486 VDD.n485 0.00658571
R32357 VDD.n486 VDD.n247 0.00658571
R32358 VDD.n492 VDD.n247 0.00658571
R32359 VDD.n493 VDD.n492 0.00658571
R32360 VDD.n494 VDD.n493 0.00658571
R32361 VDD.n494 VDD.n243 0.00658571
R32362 VDD.n500 VDD.n243 0.00658571
R32363 VDD.n501 VDD.n500 0.00658571
R32364 VDD.n502 VDD.n501 0.00658571
R32365 VDD.n502 VDD.n239 0.00658571
R32366 VDD.n508 VDD.n239 0.00658571
R32367 VDD.n509 VDD.n508 0.00658571
R32368 VDD.n510 VDD.n509 0.00658571
R32369 VDD.n510 VDD.n235 0.00658571
R32370 VDD.n516 VDD.n235 0.00658571
R32371 VDD.n517 VDD.n516 0.00658571
R32372 VDD.n518 VDD.n517 0.00658571
R32373 VDD.n518 VDD.n231 0.00658571
R32374 VDD.n524 VDD.n231 0.00658571
R32375 VDD.n525 VDD.n524 0.00658571
R32376 VDD.n526 VDD.n525 0.00658571
R32377 VDD.n526 VDD.n227 0.00658571
R32378 VDD.n532 VDD.n227 0.00658571
R32379 VDD.n533 VDD.n532 0.00658571
R32380 VDD.n534 VDD.n533 0.00658571
R32381 VDD.n534 VDD.n223 0.00658571
R32382 VDD.n540 VDD.n223 0.00658571
R32383 VDD.n541 VDD.n540 0.00658571
R32384 VDD.n542 VDD.n541 0.00658571
R32385 VDD.n549 VDD.n219 0.00658571
R32386 VDD.n688 VDD.n687 0.00658571
R32387 VDD.n687 VDD.n686 0.00658571
R32388 VDD.n686 VDD.n678 0.00658571
R32389 VDD.n679 VDD.n678 0.00658571
R32390 VDD.n679 VDD.n611 0.00658571
R32391 VDD.n708 VDD.n611 0.00658571
R32392 VDD.n709 VDD.n708 0.00658571
R32393 VDD.n710 VDD.n709 0.00658571
R32394 VDD.n710 VDD.n607 0.00658571
R32395 VDD.n716 VDD.n607 0.00658571
R32396 VDD.n717 VDD.n716 0.00658571
R32397 VDD.n718 VDD.n717 0.00658571
R32398 VDD.n718 VDD.n603 0.00658571
R32399 VDD.n724 VDD.n603 0.00658571
R32400 VDD.n725 VDD.n724 0.00658571
R32401 VDD.n726 VDD.n725 0.00658571
R32402 VDD.n726 VDD.n599 0.00658571
R32403 VDD.n732 VDD.n599 0.00658571
R32404 VDD.n733 VDD.n732 0.00658571
R32405 VDD.n734 VDD.n733 0.00658571
R32406 VDD.n734 VDD.n595 0.00658571
R32407 VDD.n740 VDD.n595 0.00658571
R32408 VDD.n741 VDD.n740 0.00658571
R32409 VDD.n742 VDD.n741 0.00658571
R32410 VDD.n742 VDD.n591 0.00658571
R32411 VDD.n748 VDD.n591 0.00658571
R32412 VDD.n749 VDD.n748 0.00658571
R32413 VDD.n786 VDD.n749 0.00658571
R32414 VDD.n786 VDD.n785 0.00658571
R32415 VDD.n785 VDD.n784 0.00658571
R32416 VDD.n784 VDD.n750 0.00658571
R32417 VDD.n778 VDD.n750 0.00658571
R32418 VDD.n778 VDD.n777 0.00658571
R32419 VDD.n777 VDD.n776 0.00658571
R32420 VDD.n776 VDD.n754 0.00658571
R32421 VDD.n758 VDD.n754 0.00658571
R32422 VDD.n768 VDD.n758 0.00658571
R32423 VDD.n768 VDD.n767 0.00658571
R32424 VDD.n767 VDD.n766 0.00658571
R32425 VDD.n766 VDD.n759 0.00658571
R32426 VDD.n760 VDD.n759 0.00658571
R32427 VDD.n760 VDD.n582 0.00658571
R32428 VDD.n839 VDD.n582 0.00658571
R32429 VDD.n840 VDD.n839 0.00658571
R32430 VDD.n841 VDD.n840 0.00658571
R32431 VDD.n841 VDD.n578 0.00658571
R32432 VDD.n847 VDD.n578 0.00658571
R32433 VDD.n848 VDD.n847 0.00658571
R32434 VDD.n849 VDD.n848 0.00658571
R32435 VDD.n849 VDD.n574 0.00658571
R32436 VDD.n855 VDD.n574 0.00658571
R32437 VDD.n856 VDD.n855 0.00658571
R32438 VDD.n857 VDD.n856 0.00658571
R32439 VDD.n857 VDD.n570 0.00658571
R32440 VDD.n863 VDD.n570 0.00658571
R32441 VDD.n864 VDD.n863 0.00658571
R32442 VDD.n865 VDD.n864 0.00658571
R32443 VDD.n865 VDD.n566 0.00658571
R32444 VDD.n871 VDD.n566 0.00658571
R32445 VDD.n872 VDD.n871 0.00658571
R32446 VDD.n873 VDD.n872 0.00658571
R32447 VDD.n873 VDD.n562 0.00658571
R32448 VDD.n879 VDD.n562 0.00658571
R32449 VDD.n880 VDD.n879 0.00658571
R32450 VDD.n896 VDD.n880 0.00658571
R32451 VDD.n896 VDD.n895 0.00658571
R32452 VDD.n895 VDD.n894 0.00658571
R32453 VDD.n894 VDD.n881 0.00658571
R32454 VDD.n888 VDD.n881 0.00658571
R32455 VDD.n888 VDD.n887 0.00658571
R32456 VDD.n887 VDD.n886 0.00658571
R32457 VDD.n886 VDD.n2 0.00658571
R32458 VDD.n922 VDD.n920 0.00658571
R32459 VDD.n73 VDD 0.00654478
R32460 VDD.n47 VDD 0.00654478
R32461 VDD.n90 VDD 0.00642105
R32462 VDD.n395 VDD 0.00642105
R32463 VDD.n329 VDD.n328 0.00641906
R32464 VDD.n328 VDD.n314 0.00641906
R32465 VDD VDD.n219 0.00641429
R32466 VDD.n920 VDD 0.00641429
R32467 VDD.n692 VDD.n691 0.00583571
R32468 VDD.n195 VDD.n20 0.00575843
R32469 VDD.n704 VDD.n613 0.00564286
R32470 VDD.n550 VDD.n218 0.00548841
R32471 VDD.n923 VDD.n919 0.00548841
R32472 VDD.n542 VDD 0.00538571
R32473 VDD.n836 VDD.n835 0.00512857
R32474 VDD.n321 VDD 0.00505312
R32475 VDD VDD.n326 0.00505312
R32476 VDD.n331 VDD.n314 0.00505312
R32477 VDD.n835 VDD.n584 0.005
R32478 VDD.n705 VDD.n704 0.00448571
R32479 VDD.n327 VDD 0.00399073
R32480 VDD.n772 VDD.n586 0.00332857
R32481 VDD.n402 VDD.n401 0.0032
R32482 VDD.n341 VDD.n337 0.00249286
R32483 VDD.n546 VDD 0.0023
R32484 VDD.n545 VDD 0.0023
R32485 VDD VDD.n933 0.0023
R32486 VDD.n932 VDD 0.0023
R32487 VDD.n899 VDD.n898 0.00217143
R32488 VDD VDD.n823 0.002
R32489 VDD.n555 VDD.n207 0.00185
R32490 VDD.n214 VDD.n8 0.00185
R32491 VDD.n930 VDD.n907 0.00185
R32492 VDD.n918 VDD.n917 0.00185
R32493 VDD VDD.n220 0.0017
R32494 VDD.n789 VDD.n788 0.00152857
R32495 VDD.n220 VDD 0.000671429
R32496 VDD VDD.n2 0.000671429
R32497 VDD.n353 VDD.n352 0.000564286
R32498 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n4 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n3 1821.97
R32499 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n152 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n147 227.274
R32500 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n163 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n153 227.274
R32501 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n129 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n115 227.274
R32502 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n130 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n111 227.274
R32503 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n89 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n78 227.274
R32504 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n95 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n72 227.274
R32505 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n62 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n39 227.274
R32506 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n61 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n60 227.274
R32507 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n19 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n18 227.274
R32508 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n185 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n4 227.274
R32509 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.t4 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n152 113.636
R32510 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n163 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.t4 113.636
R32511 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.t3 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n129 113.636
R32512 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n130 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.t3 113.636
R32513 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n89 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.t1 113.636
R32514 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.t1 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n72 113.636
R32515 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n62 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.t2 113.636
R32516 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.t2 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n61 113.636
R32517 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n18 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.t5 113.636
R32518 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n185 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.t5 113.636
R32519 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n175 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.t8 46.7726
R32520 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n140 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.t17 46.7726
R32521 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n105 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.t9 46.7726
R32522 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n99 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.t24 46.7726
R32523 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n66 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.t6 46.7726
R32524 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n24 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.t10 46.7726
R32525 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n179 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.t19 46.7726
R32526 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n29 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.t16 43.0184
R32527 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n175 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.t13 41.2455
R32528 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n140 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.t20 41.2455
R32529 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n105 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.t14 41.2455
R32530 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n99 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.t7 41.2455
R32531 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n66 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.t12 41.2455
R32532 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n24 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.t15 41.2455
R32533 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n179 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.t22 41.2455
R32534 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n32 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.t11 35.9269
R32535 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n102 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n68 30.9842
R32536 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n32 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.t23 30.9212
R32537 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n29 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.t25 30.9212
R32538 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n31 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n30 27.1154
R32539 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n107 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n104 25.673
R32540 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n31 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n27 24.3538
R32541 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n102 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n101 21.9818
R32542 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n34 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE 18.5934
R32543 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n104 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n103 16.1705
R32544 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.t0 11.0117
R32545 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n16 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n11 10.5005
R32546 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n12 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n5 10.5005
R32547 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n186 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n5 10.5005
R32548 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n187 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n186 10.5005
R32549 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n189 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n2 10.5005
R32550 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n21 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n7 10.5005
R32551 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n184 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n7 10.5005
R32552 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n184 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n9 10.5005
R32553 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n171 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n170 10.5005
R32554 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n168 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n149 10.5005
R32555 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n164 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n149 10.5005
R32556 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n164 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n151 10.5005
R32557 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n173 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n146 10.5005
R32558 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n162 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n146 10.5005
R32559 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n162 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n154 10.5005
R32560 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n124 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n123 10.5005
R32561 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n128 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n116 10.5005
R32562 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n128 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n110 10.5005
R32563 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n138 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n110 10.5005
R32564 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n136 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n135 10.5005
R32565 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n120 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n114 10.5005
R32566 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n131 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n114 10.5005
R32567 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n132 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n131 10.5005
R32568 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n90 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n77 10.5005
R32569 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n90 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n74 10.5005
R32570 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n94 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n74 10.5005
R32571 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n84 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n83 10.5005
R32572 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n88 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n79 10.5005
R32573 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n88 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n71 10.5005
R32574 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n96 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n71 10.5005
R32575 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n63 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n37 10.5005
R32576 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n63 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n38 10.5005
R32577 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n52 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n38 10.5005
R32578 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n54 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n43 10.5005
R32579 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n47 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n40 10.5005
R32580 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n41 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n40 10.5005
R32581 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n58 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n41 10.5005
R32582 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n27 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n25 7.84234
R32583 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n181 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n178 7.68484
R32584 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n158 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n154 7.3505
R32585 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n156 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n151 7.3505
R32586 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n94 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n73 7.3505
R32587 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n47 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n46 7.3505
R32588 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n107 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n106 6.57761
R32589 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n160 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n154 6.3005
R32590 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n154 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n153 6.3005
R32591 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n162 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n161 6.3005
R32592 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n163 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n162 6.3005
R32593 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n146 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n144 6.3005
R32594 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n152 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n146 6.3005
R32595 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n156 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n155 6.3005
R32596 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n159 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n158 6.3005
R32597 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n151 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n150 6.3005
R32598 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n153 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n151 6.3005
R32599 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n165 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n164 6.3005
R32600 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n164 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n163 6.3005
R32601 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n166 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n149 6.3005
R32602 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n152 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n149 6.3005
R32603 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n168 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n167 6.3005
R32604 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n171 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n145 6.3005
R32605 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n170 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n148 6.3005
R32606 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n174 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n173 6.3005
R32607 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n125 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n124 6.3005
R32608 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n123 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n122 6.3005
R32609 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n110 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n108 6.3005
R32610 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n130 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n110 6.3005
R32611 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n128 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n127 6.3005
R32612 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n129 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n128 6.3005
R32613 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n126 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n116 6.3005
R32614 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n133 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n132 6.3005
R32615 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n131 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n113 6.3005
R32616 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n131 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n130 6.3005
R32617 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n119 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n114 6.3005
R32618 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n129 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n114 6.3005
R32619 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n121 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n120 6.3005
R32620 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n135 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n134 6.3005
R32621 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n136 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n109 6.3005
R32622 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n139 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n138 6.3005
R32623 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n85 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n84 6.3005
R32624 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n83 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n82 6.3005
R32625 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n75 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n73 6.3005
R32626 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n94 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n93 6.3005
R32627 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n95 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n94 6.3005
R32628 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n92 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n74 6.3005
R32629 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n74 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n72 6.3005
R32630 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n91 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n90 6.3005
R32631 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n90 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n89 6.3005
R32632 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n77 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n76 6.3005
R32633 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n71 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n69 6.3005
R32634 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n72 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n71 6.3005
R32635 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n88 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n87 6.3005
R32636 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n89 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n88 6.3005
R32637 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n86 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n79 6.3005
R32638 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n96 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n95 6.3005
R32639 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n46 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n44 6.3005
R32640 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n58 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n57 6.3005
R32641 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n50 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n41 6.3005
R32642 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n61 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n41 6.3005
R32643 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n49 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n40 6.3005
R32644 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n62 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n40 6.3005
R32645 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n48 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n47 6.3005
R32646 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n47 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n39 6.3005
R32647 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n56 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n43 6.3005
R32648 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n55 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n54 6.3005
R32649 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n53 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n52 6.3005
R32650 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n51 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n38 6.3005
R32651 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n61 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n38 6.3005
R32652 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n64 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n63 6.3005
R32653 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n63 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n62 6.3005
R32654 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n39 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n37 6.3005
R32655 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n182 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n9 6.3005
R32656 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n184 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n183 6.3005
R32657 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n185 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n184 6.3005
R32658 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n23 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n7 6.3005
R32659 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n18 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n7 6.3005
R32660 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n22 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n21 6.3005
R32661 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n11 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n10 6.3005
R32662 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n16 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n15 6.3005
R32663 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n190 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n189 6.3005
R32664 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n2 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n0 6.3005
R32665 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n187 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n1 6.3005
R32666 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n186 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n6 6.3005
R32667 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n186 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n185 6.3005
R32668 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n13 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n5 6.3005
R32669 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n18 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n5 6.3005
R32670 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n14 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n12 6.3005
R32671 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n27 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n26 5.60822
R32672 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n97 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n70 5.18619
R32673 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n45 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n36 5.18619
R32674 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n35 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE 4.92208
R32675 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n177 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n174 4.67458
R32676 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n142 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n139 4.67458
R32677 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n182 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n181 4.67458
R32678 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n30 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE 4.56015
R32679 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n143 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n107 4.54195
R32680 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n101 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n98 4.53118
R32681 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n68 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n65 4.53118
R32682 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n178 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n177 4.22221
R32683 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n143 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n142 4.22221
R32684 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n29 4.00158
R32685 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n176 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n175 4.0005
R32686 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n141 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n140 4.0005
R32687 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n106 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n105 4.0005
R32688 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n100 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n99 4.0005
R32689 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n67 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n66 4.0005
R32690 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n32 4.0005
R32691 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n25 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n24 4.0005
R32692 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n180 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n179 4.0005
R32693 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n30 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n28 3.60322
R32694 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n158 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n157 2.86464
R32695 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n157 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n156 2.86464
R32696 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n73 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n70 2.86464
R32697 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n46 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n45 2.86464
R32698 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n178 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n143 2.62471
R32699 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n177 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n176 2.49418
R32700 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n142 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n141 2.49418
R32701 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n181 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n180 2.49418
R32702 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n34 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n33 2.4573
R32703 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n21 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n20 2.32205
R32704 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n17 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n12 2.32205
R32705 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n9 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n8 2.32205
R32706 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n189 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n188 2.32205
R32707 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n172 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n171 2.32205
R32708 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n169 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n168 2.32205
R32709 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n170 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n169 2.32205
R32710 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n173 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n172 2.32205
R32711 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n124 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n117 2.32205
R32712 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n123 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n118 2.32205
R32713 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n117 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n116 2.32205
R32714 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n137 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n136 2.32205
R32715 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n135 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n112 2.32205
R32716 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n132 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n112 2.32205
R32717 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n120 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n118 2.32205
R32718 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n138 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n137 2.32205
R32719 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n97 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n96 2.32205
R32720 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n84 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n80 2.32205
R32721 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n83 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n81 2.32205
R32722 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n81 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n77 2.32205
R32723 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n80 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n79 2.32205
R32724 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n37 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n36 2.32205
R32725 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n52 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n42 2.32205
R32726 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n59 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n43 2.32205
R32727 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n59 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n58 2.32205
R32728 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n54 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n42 2.32205
R32729 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n20 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n11 2.32205
R32730 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n17 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n16 2.32205
R32731 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n8 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n2 2.32205
R32732 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n188 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n187 2.32205
R32733 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n101 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n100 2.2505
R32734 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n68 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n67 2.2505
R32735 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n103 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n102 2.2505
R32736 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n169 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n147 1.99047
R32737 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n172 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n147 1.99047
R32738 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n117 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n115 1.99047
R32739 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n118 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n115 1.99047
R32740 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n112 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n111 1.99047
R32741 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n137 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n111 1.99047
R32742 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n80 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n78 1.99047
R32743 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n81 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n78 1.99047
R32744 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n98 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n97 1.99047
R32745 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n60 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n59 1.99047
R32746 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n60 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n42 1.99047
R32747 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n65 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n36 1.99047
R32748 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n8 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n4 1.99047
R32749 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n20 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n19 1.99047
R32750 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n188 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n4 1.99047
R32751 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n19 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n17 1.99047
R32752 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n157 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n153 1.71918
R32753 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n95 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n70 1.71918
R32754 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n45 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n39 1.71918
R32755 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n28 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.t21 1.30393
R32756 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n26 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.t18 1.30393
R32757 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n33 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.t26 1.30145
R32758 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n34 0.840105
R32759 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n35 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE 0.549731
R32760 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n103 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n35 0.411421
R32761 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n23 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n22 0.1505
R32762 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n161 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n160 0.1505
R32763 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n167 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n166 0.1505
R32764 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n165 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n150 0.1505
R32765 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n127 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n126 0.1505
R32766 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n121 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n119 0.1505
R32767 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n133 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n113 0.1505
R32768 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n91 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n76 0.1505
R32769 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n93 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n92 0.1505
R32770 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n87 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n86 0.1505
R32771 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n49 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n48 0.1505
R32772 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n57 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n50 0.1505
R32773 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n53 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n51 0.1505
R32774 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n14 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n13 0.1505
R32775 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n6 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n1 0.1505
R32776 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n174 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n145 0.148132
R32777 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n139 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n109 0.148132
R32778 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n182 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n0 0.148132
R32779 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n98 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n69 0.1235
R32780 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n65 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n64 0.1235
R32781 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n22 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n10 0.1055
R32782 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n15 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n14 0.1055
R32783 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n160 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n159 0.1055
R32784 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n155 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n150 0.1055
R32785 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n167 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n148 0.1055
R32786 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n126 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n125 0.1055
R32787 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n122 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n121 0.1055
R32788 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n134 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n133 0.1055
R32789 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n93 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n75 0.1055
R32790 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n86 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n85 0.1055
R32791 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n82 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n76 0.1055
R32792 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n48 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n44 0.1055
R32793 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n55 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n53 0.1055
R32794 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n57 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n56 0.1055
R32795 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n190 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n1 0.1055
R32796 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n183 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n182 0.1005
R32797 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n174 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n144 0.1005
R32798 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n139 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n108 0.1005
R32799 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n10 0.0755
R32800 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n15 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE 0.0755
R32801 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n23 0.0755
R32802 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n183 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE 0.0755
R32803 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n144 0.0755
R32804 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n161 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE 0.0755
R32805 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n159 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE 0.0755
R32806 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n155 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE 0.0755
R32807 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n166 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE 0.0755
R32808 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n165 0.0755
R32809 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n145 0.0755
R32810 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n148 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE 0.0755
R32811 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n125 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE 0.0755
R32812 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n122 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE 0.0755
R32813 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n127 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE 0.0755
R32814 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n108 0.0755
R32815 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n119 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE 0.0755
R32816 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n113 0.0755
R32817 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n109 0.0755
R32818 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n134 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE 0.0755
R32819 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n75 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE 0.0755
R32820 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n91 0.0755
R32821 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n92 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE 0.0755
R32822 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n85 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE 0.0755
R32823 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n82 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE 0.0755
R32824 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n87 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE 0.0755
R32825 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n69 0.0755
R32826 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n44 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE 0.0755
R32827 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n49 0.0755
R32828 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n50 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE 0.0755
R32829 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n55 0.0755
R32830 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n56 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE 0.0755
R32831 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n64 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE 0.0755
R32832 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n51 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE 0.0755
R32833 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n13 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE 0.0755
R32834 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n6 0.0755
R32835 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n0 0.0755
R32836 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n190 0.0755
R32837 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n98 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE 0.0455
R32838 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n65 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE 0.0455
R32839 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n33 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE 0.01495
R32840 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n28 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE 0.012475
R32841 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n26 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE 0.012475
R32842 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n106 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE 0.004
R32843 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n104 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n31 0.00286842
R32844 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n25 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE 0.0025
R32845 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n100 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE 0.002
R32846 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n67 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE 0.002
R32847 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n176 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE 0.00168421
R32848 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n141 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE 0.00168421
R32849 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n180 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE 0.00168421
R32850 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_1.nmos_6p0_CDNS_4066195314511_1.D GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_1.nmos_6p0_CDNS_4066195314511_0.S.n0 1.15854
R32851 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_1.nmos_6p0_CDNS_4066195314511_0.S.n0 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_1.nmos_6p0_CDNS_4066195314511_0.S.t1 0.5465
R32852 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_1.nmos_6p0_CDNS_4066195314511_0.S.n0 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_1.nmos_6p0_CDNS_4066195314511_0.S.t0 0.5465
R32853 GF_NI_IN_C_BASE_0.comp018green_out_predrv_0.A GF_NI_IN_C_BASE_0.comp018green_out_predrv_0.A.t8 82.0028
R32854 GF_NI_IN_C_BASE_0.comp018green_out_predrv_0.A GF_NI_IN_C_BASE_0.comp018green_out_predrv_0.A.t5 82.0028
R32855 GF_NI_IN_C_BASE_0.comp018green_out_predrv_0.A GF_NI_IN_C_BASE_0.comp018green_out_predrv_0.A.t7 82.0028
R32856 GF_NI_IN_C_BASE_0.comp018green_out_predrv_0.A GF_NI_IN_C_BASE_0.comp018green_out_predrv_0.A.t3 82.0028
R32857 GF_NI_IN_C_BASE_0.comp018green_out_predrv_0.A GF_NI_IN_C_BASE_0.comp018green_out_predrv_0.A.t2 42.2319
R32858 GF_NI_IN_C_BASE_0.comp018green_out_predrv_0.A GF_NI_IN_C_BASE_0.comp018green_out_predrv_0.A.t6 42.2319
R32859 GF_NI_IN_C_BASE_0.comp018green_out_predrv_0.A GF_NI_IN_C_BASE_0.comp018green_out_predrv_0.A.t9 42.2319
R32860 GF_NI_IN_C_BASE_0.comp018green_out_predrv_0.A GF_NI_IN_C_BASE_0.comp018green_out_predrv_0.A.t4 42.2319
R32861 GF_NI_IN_C_BASE_0.comp018green_out_predrv_0.A.n1 GF_NI_IN_C_BASE_0.comp018green_out_predrv_0.A 10.5577
R32862 GF_NI_IN_C_BASE_0.comp018green_out_predrv_0.A.n0 GF_NI_IN_C_BASE_0.comp018green_out_predrv_0.A 10.4346
R32863 GF_NI_IN_C_BASE_0.comp018green_out_predrv_0.A.n0 GF_NI_IN_C_BASE_0.comp018green_out_predrv_0.A 6.98616
R32864 GF_NI_IN_C_BASE_0.comp018green_out_predrv_0.A.n1 GF_NI_IN_C_BASE_0.comp018green_out_predrv_0.A.n0 4.85103
R32865 GF_NI_IN_C_BASE_0.comp018green_out_predrv_0.A GF_NI_IN_C_BASE_0.comp018green_out_predrv_0.A.n2 4.69358
R32866 GF_NI_IN_C_BASE_0.comp018green_out_predrv_0.A.n2 GF_NI_IN_C_BASE_0.comp018green_out_predrv_0.A 4.47707
R32867 GF_NI_IN_C_BASE_0.comp018green_out_predrv_0.A.n2 GF_NI_IN_C_BASE_0.comp018green_out_predrv_0.A.n1 2.2505
R32868 GF_NI_IN_C_BASE_0.comp018green_out_predrv_0.A GF_NI_IN_C_BASE_0.comp018green_out_predrv_0.A.t1 2.04837
R32869 GF_NI_IN_C_BASE_0.comp018green_out_predrv_0.A GF_NI_IN_C_BASE_0.comp018green_out_predrv_0.A.t0 1.49421
R32870 GF_NI_IN_C_BASE_0.comp018green_out_predrv_1.nmos_6p0_CDNS_4066195314519_0.D.n1 GF_NI_IN_C_BASE_0.comp018green_out_predrv_1.nmos_6p0_CDNS_4066195314519_0.D.t4 80.4772
R32871 GF_NI_IN_C_BASE_0.comp018green_out_predrv_1.nmos_6p0_CDNS_4066195314519_0.D.n0 GF_NI_IN_C_BASE_0.comp018green_out_predrv_1.nmos_6p0_CDNS_4066195314519_0.D.t6 80.4772
R32872 GF_NI_IN_C_BASE_0.comp018green_out_predrv_1.nmos_6p0_CDNS_4066195314519_0.D.n1 GF_NI_IN_C_BASE_0.comp018green_out_predrv_1.nmos_6p0_CDNS_4066195314519_0.D.t3 62.5719
R32873 GF_NI_IN_C_BASE_0.comp018green_out_predrv_1.nmos_6p0_CDNS_4066195314519_0.D.n0 GF_NI_IN_C_BASE_0.comp018green_out_predrv_1.nmos_6p0_CDNS_4066195314519_0.D.t7 62.5719
R32874 GF_NI_IN_C_BASE_0.comp018green_out_predrv_1.nmos_6p0_CDNS_4066195314519_0.D.n4 GF_NI_IN_C_BASE_0.comp018green_out_predrv_1.nmos_6p0_CDNS_4066195314519_0.D.t8 45.4098
R32875 GF_NI_IN_C_BASE_0.comp018green_out_predrv_1.nmos_6p0_CDNS_4066195314519_0.D.n4 GF_NI_IN_C_BASE_0.comp018green_out_predrv_1.nmos_6p0_CDNS_4066195314519_0.D.t5 34.4148
R32876 GF_NI_IN_C_BASE_0.comp018green_out_predrv_1.nmos_6p0_CDNS_4066195314519_0.D.n2 GF_NI_IN_C_BASE_0.comp018green_out_predrv_1.nmos_6p0_CDNS_4066195314519_0.D.n1 8.06816
R32877 GF_NI_IN_C_BASE_0.comp018green_out_predrv_1.nmos_6p0_CDNS_4066195314519_0.D.n2 GF_NI_IN_C_BASE_0.comp018green_out_predrv_1.nmos_6p0_CDNS_4066195314519_0.D.n0 8.06816
R32878 GF_NI_IN_C_BASE_0.comp018green_out_predrv_1.nmos_6p0_CDNS_4066195314519_0.D.n3 GF_NI_IN_C_BASE_0.comp018green_out_predrv_1.nmos_6p0_CDNS_4066195314519_0.D.n2 6.31953
R32879 GF_NI_IN_C_BASE_0.comp018green_out_predrv_1.nmos_6p0_CDNS_4066195314519_0.D.t0 GF_NI_IN_C_BASE_0.comp018green_out_predrv_1.nmos_6p0_CDNS_4066195314519_0.D.n4 6.08116
R32880 GF_NI_IN_C_BASE_0.comp018green_out_predrv_1.nmos_6p0_CDNS_4066195314519_0.D.t1 GF_NI_IN_C_BASE_0.comp018green_out_predrv_1.nmos_6p0_CDNS_4066195314519_0.D.n3 4.80357
R32881 GF_NI_IN_C_BASE_0.comp018green_out_predrv_1.nmos_6p0_CDNS_4066195314519_0.D.n3 GF_NI_IN_C_BASE_0.comp018green_out_predrv_1.nmos_6p0_CDNS_4066195314519_0.D.t2 4.54043
R32882 GF_NI_IN_C_BASE_0.comp018green_out_predrv_1.nmos_6p0_CDNS_4066195314519_0.D.t1 GF_NI_IN_C_BASE_0.comp018green_out_predrv_1.nmos_6p0_CDNS_4066195314519_0.D.t0 1.1409
R32883 GF_NI_IN_C_BASE_0.comp018green_out_predrv_1.nmos_6p0_CDNS_4066195314519_0.D.t0 GF_NI_IN_C_BASE_0.comp018green_out_predrv_1.nmos_6p0_CDNS_4066195314519_0.D 0.702557
R32884 PAD.n6374 PAD.n6373 4.5005
R32885 PAD.n6374 PAD.n5982 4.5005
R32886 PAD.n6374 PAD.n5981 4.5005
R32887 PAD.n6374 PAD.n5980 4.5005
R32888 PAD.n11507 PAD.n11156 4.5005
R32889 PAD.n11302 PAD.n11156 4.5005
R32890 PAD.n11509 PAD.n11156 4.5005
R32891 PAD.n11156 PAD.n11100 4.5005
R32892 PAD.n6373 PAD.n6032 4.5005
R32893 PAD.n6032 PAD.n5981 4.5005
R32894 PAD.n6032 PAD.n5979 4.5005
R32895 PAD.n11507 PAD.n11154 4.5005
R32896 PAD.n11302 PAD.n11154 4.5005
R32897 PAD.n11509 PAD.n11154 4.5005
R32898 PAD.n11507 PAD.n11158 4.5005
R32899 PAD.n11509 PAD.n11158 4.5005
R32900 PAD.n11158 PAD.n11105 4.5005
R32901 PAD.n11507 PAD.n11153 4.5005
R32902 PAD.n11509 PAD.n11153 4.5005
R32903 PAD.n11153 PAD.n11105 4.5005
R32904 PAD.n11507 PAD.n11160 4.5005
R32905 PAD.n11509 PAD.n11160 4.5005
R32906 PAD.n11160 PAD.n11105 4.5005
R32907 PAD.n11507 PAD.n11152 4.5005
R32908 PAD.n11509 PAD.n11152 4.5005
R32909 PAD.n11152 PAD.n11105 4.5005
R32910 PAD.n11507 PAD.n11162 4.5005
R32911 PAD.n11509 PAD.n11162 4.5005
R32912 PAD.n11162 PAD.n11105 4.5005
R32913 PAD.n11507 PAD.n11151 4.5005
R32914 PAD.n11509 PAD.n11151 4.5005
R32915 PAD.n11151 PAD.n11105 4.5005
R32916 PAD.n11507 PAD.n11164 4.5005
R32917 PAD.n11509 PAD.n11164 4.5005
R32918 PAD.n11164 PAD.n11105 4.5005
R32919 PAD.n11507 PAD.n11150 4.5005
R32920 PAD.n11509 PAD.n11150 4.5005
R32921 PAD.n11150 PAD.n11105 4.5005
R32922 PAD.n11507 PAD.n11166 4.5005
R32923 PAD.n11509 PAD.n11166 4.5005
R32924 PAD.n11166 PAD.n11105 4.5005
R32925 PAD.n11507 PAD.n11149 4.5005
R32926 PAD.n11509 PAD.n11149 4.5005
R32927 PAD.n11149 PAD.n11105 4.5005
R32928 PAD.n11507 PAD.n11168 4.5005
R32929 PAD.n11509 PAD.n11168 4.5005
R32930 PAD.n11168 PAD.n11105 4.5005
R32931 PAD.n11507 PAD.n11148 4.5005
R32932 PAD.n11509 PAD.n11148 4.5005
R32933 PAD.n11148 PAD.n11105 4.5005
R32934 PAD.n11507 PAD.n11170 4.5005
R32935 PAD.n11509 PAD.n11170 4.5005
R32936 PAD.n11170 PAD.n11105 4.5005
R32937 PAD.n11507 PAD.n11147 4.5005
R32938 PAD.n11509 PAD.n11147 4.5005
R32939 PAD.n11147 PAD.n11105 4.5005
R32940 PAD.n11507 PAD.n11172 4.5005
R32941 PAD.n11509 PAD.n11172 4.5005
R32942 PAD.n11172 PAD.n11105 4.5005
R32943 PAD.n11507 PAD.n11146 4.5005
R32944 PAD.n11509 PAD.n11146 4.5005
R32945 PAD.n11146 PAD.n11105 4.5005
R32946 PAD.n11507 PAD.n11174 4.5005
R32947 PAD.n11509 PAD.n11174 4.5005
R32948 PAD.n11174 PAD.n11105 4.5005
R32949 PAD.n11507 PAD.n11145 4.5005
R32950 PAD.n11509 PAD.n11145 4.5005
R32951 PAD.n11145 PAD.n11105 4.5005
R32952 PAD.n11507 PAD.n11176 4.5005
R32953 PAD.n11509 PAD.n11176 4.5005
R32954 PAD.n11176 PAD.n11105 4.5005
R32955 PAD.n11507 PAD.n11144 4.5005
R32956 PAD.n11509 PAD.n11144 4.5005
R32957 PAD.n11144 PAD.n11105 4.5005
R32958 PAD.n11507 PAD.n11178 4.5005
R32959 PAD.n11509 PAD.n11178 4.5005
R32960 PAD.n11178 PAD.n11105 4.5005
R32961 PAD.n11507 PAD.n11143 4.5005
R32962 PAD.n11509 PAD.n11143 4.5005
R32963 PAD.n11143 PAD.n11105 4.5005
R32964 PAD.n11507 PAD.n11180 4.5005
R32965 PAD.n11509 PAD.n11180 4.5005
R32966 PAD.n11180 PAD.n11105 4.5005
R32967 PAD.n11507 PAD.n11142 4.5005
R32968 PAD.n11509 PAD.n11142 4.5005
R32969 PAD.n11142 PAD.n11105 4.5005
R32970 PAD.n11507 PAD.n11182 4.5005
R32971 PAD.n11509 PAD.n11182 4.5005
R32972 PAD.n11182 PAD.n11105 4.5005
R32973 PAD.n11507 PAD.n11141 4.5005
R32974 PAD.n11509 PAD.n11141 4.5005
R32975 PAD.n11141 PAD.n11105 4.5005
R32976 PAD.n11507 PAD.n11184 4.5005
R32977 PAD.n11509 PAD.n11184 4.5005
R32978 PAD.n11184 PAD.n11105 4.5005
R32979 PAD.n11507 PAD.n11140 4.5005
R32980 PAD.n11509 PAD.n11140 4.5005
R32981 PAD.n11140 PAD.n11105 4.5005
R32982 PAD.n11507 PAD.n11186 4.5005
R32983 PAD.n11509 PAD.n11186 4.5005
R32984 PAD.n11186 PAD.n11105 4.5005
R32985 PAD.n11507 PAD.n11139 4.5005
R32986 PAD.n11509 PAD.n11139 4.5005
R32987 PAD.n11139 PAD.n11105 4.5005
R32988 PAD.n11507 PAD.n11188 4.5005
R32989 PAD.n11509 PAD.n11188 4.5005
R32990 PAD.n11188 PAD.n11105 4.5005
R32991 PAD.n11507 PAD.n11138 4.5005
R32992 PAD.n11509 PAD.n11138 4.5005
R32993 PAD.n11138 PAD.n11105 4.5005
R32994 PAD.n11507 PAD.n11190 4.5005
R32995 PAD.n11509 PAD.n11190 4.5005
R32996 PAD.n11190 PAD.n11105 4.5005
R32997 PAD.n11507 PAD.n11137 4.5005
R32998 PAD.n11509 PAD.n11137 4.5005
R32999 PAD.n11137 PAD.n11105 4.5005
R33000 PAD.n11507 PAD.n11192 4.5005
R33001 PAD.n11509 PAD.n11192 4.5005
R33002 PAD.n11192 PAD.n11105 4.5005
R33003 PAD.n11507 PAD.n11136 4.5005
R33004 PAD.n11509 PAD.n11136 4.5005
R33005 PAD.n11136 PAD.n11105 4.5005
R33006 PAD.n11507 PAD.n11194 4.5005
R33007 PAD.n11509 PAD.n11194 4.5005
R33008 PAD.n11194 PAD.n11105 4.5005
R33009 PAD.n11507 PAD.n11135 4.5005
R33010 PAD.n11509 PAD.n11135 4.5005
R33011 PAD.n11135 PAD.n11105 4.5005
R33012 PAD.n11507 PAD.n11196 4.5005
R33013 PAD.n11509 PAD.n11196 4.5005
R33014 PAD.n11196 PAD.n11105 4.5005
R33015 PAD.n11507 PAD.n11134 4.5005
R33016 PAD.n11509 PAD.n11134 4.5005
R33017 PAD.n11134 PAD.n11105 4.5005
R33018 PAD.n11507 PAD.n11198 4.5005
R33019 PAD.n11509 PAD.n11198 4.5005
R33020 PAD.n11198 PAD.n11105 4.5005
R33021 PAD.n11507 PAD.n11133 4.5005
R33022 PAD.n11509 PAD.n11133 4.5005
R33023 PAD.n11133 PAD.n11105 4.5005
R33024 PAD.n11507 PAD.n11200 4.5005
R33025 PAD.n11509 PAD.n11200 4.5005
R33026 PAD.n11200 PAD.n11105 4.5005
R33027 PAD.n11507 PAD.n11132 4.5005
R33028 PAD.n11509 PAD.n11132 4.5005
R33029 PAD.n11132 PAD.n11105 4.5005
R33030 PAD.n11507 PAD.n11202 4.5005
R33031 PAD.n11509 PAD.n11202 4.5005
R33032 PAD.n11202 PAD.n11105 4.5005
R33033 PAD.n11507 PAD.n11131 4.5005
R33034 PAD.n11509 PAD.n11131 4.5005
R33035 PAD.n11131 PAD.n11105 4.5005
R33036 PAD.n11507 PAD.n11204 4.5005
R33037 PAD.n11509 PAD.n11204 4.5005
R33038 PAD.n11204 PAD.n11105 4.5005
R33039 PAD.n11507 PAD.n11130 4.5005
R33040 PAD.n11509 PAD.n11130 4.5005
R33041 PAD.n11130 PAD.n11105 4.5005
R33042 PAD.n11507 PAD.n11206 4.5005
R33043 PAD.n11509 PAD.n11206 4.5005
R33044 PAD.n11206 PAD.n11105 4.5005
R33045 PAD.n11507 PAD.n11129 4.5005
R33046 PAD.n11509 PAD.n11129 4.5005
R33047 PAD.n11129 PAD.n11105 4.5005
R33048 PAD.n11507 PAD.n11208 4.5005
R33049 PAD.n11509 PAD.n11208 4.5005
R33050 PAD.n11208 PAD.n11105 4.5005
R33051 PAD.n11507 PAD.n11128 4.5005
R33052 PAD.n11509 PAD.n11128 4.5005
R33053 PAD.n11128 PAD.n11105 4.5005
R33054 PAD.n11507 PAD.n11210 4.5005
R33055 PAD.n11509 PAD.n11210 4.5005
R33056 PAD.n11210 PAD.n11105 4.5005
R33057 PAD.n11507 PAD.n11127 4.5005
R33058 PAD.n11509 PAD.n11127 4.5005
R33059 PAD.n11127 PAD.n11105 4.5005
R33060 PAD.n11507 PAD.n11212 4.5005
R33061 PAD.n11509 PAD.n11212 4.5005
R33062 PAD.n11212 PAD.n11105 4.5005
R33063 PAD.n11507 PAD.n11126 4.5005
R33064 PAD.n11509 PAD.n11126 4.5005
R33065 PAD.n11126 PAD.n11105 4.5005
R33066 PAD.n11507 PAD.n11214 4.5005
R33067 PAD.n11509 PAD.n11214 4.5005
R33068 PAD.n11214 PAD.n11105 4.5005
R33069 PAD.n11507 PAD.n11125 4.5005
R33070 PAD.n11509 PAD.n11125 4.5005
R33071 PAD.n11125 PAD.n11105 4.5005
R33072 PAD.n11507 PAD.n11216 4.5005
R33073 PAD.n11509 PAD.n11216 4.5005
R33074 PAD.n11216 PAD.n11105 4.5005
R33075 PAD.n11507 PAD.n11124 4.5005
R33076 PAD.n11509 PAD.n11124 4.5005
R33077 PAD.n11124 PAD.n11105 4.5005
R33078 PAD.n11507 PAD.n11218 4.5005
R33079 PAD.n11509 PAD.n11218 4.5005
R33080 PAD.n11218 PAD.n11105 4.5005
R33081 PAD.n11507 PAD.n11123 4.5005
R33082 PAD.n11509 PAD.n11123 4.5005
R33083 PAD.n11123 PAD.n11105 4.5005
R33084 PAD.n11507 PAD.n11220 4.5005
R33085 PAD.n11509 PAD.n11220 4.5005
R33086 PAD.n11220 PAD.n11105 4.5005
R33087 PAD.n11507 PAD.n11122 4.5005
R33088 PAD.n11509 PAD.n11122 4.5005
R33089 PAD.n11122 PAD.n11105 4.5005
R33090 PAD.n11507 PAD.n11222 4.5005
R33091 PAD.n11509 PAD.n11222 4.5005
R33092 PAD.n11222 PAD.n11105 4.5005
R33093 PAD.n11507 PAD.n11121 4.5005
R33094 PAD.n11509 PAD.n11121 4.5005
R33095 PAD.n11121 PAD.n11105 4.5005
R33096 PAD.n11507 PAD.n11224 4.5005
R33097 PAD.n11509 PAD.n11224 4.5005
R33098 PAD.n11224 PAD.n11105 4.5005
R33099 PAD.n11507 PAD.n11120 4.5005
R33100 PAD.n11509 PAD.n11120 4.5005
R33101 PAD.n11120 PAD.n11105 4.5005
R33102 PAD.n11507 PAD.n11226 4.5005
R33103 PAD.n11509 PAD.n11226 4.5005
R33104 PAD.n11226 PAD.n11105 4.5005
R33105 PAD.n11507 PAD.n11119 4.5005
R33106 PAD.n11509 PAD.n11119 4.5005
R33107 PAD.n11119 PAD.n11105 4.5005
R33108 PAD.n11507 PAD.n11228 4.5005
R33109 PAD.n11509 PAD.n11228 4.5005
R33110 PAD.n11228 PAD.n11105 4.5005
R33111 PAD.n11507 PAD.n11118 4.5005
R33112 PAD.n11509 PAD.n11118 4.5005
R33113 PAD.n11118 PAD.n11105 4.5005
R33114 PAD.n11507 PAD.n11230 4.5005
R33115 PAD.n11509 PAD.n11230 4.5005
R33116 PAD.n11230 PAD.n11105 4.5005
R33117 PAD.n11507 PAD.n11117 4.5005
R33118 PAD.n11509 PAD.n11117 4.5005
R33119 PAD.n11117 PAD.n11105 4.5005
R33120 PAD.n11507 PAD.n11232 4.5005
R33121 PAD.n11509 PAD.n11232 4.5005
R33122 PAD.n11232 PAD.n11105 4.5005
R33123 PAD.n11507 PAD.n11116 4.5005
R33124 PAD.n11509 PAD.n11116 4.5005
R33125 PAD.n11116 PAD.n11105 4.5005
R33126 PAD.n11507 PAD.n11234 4.5005
R33127 PAD.n11509 PAD.n11234 4.5005
R33128 PAD.n11234 PAD.n11105 4.5005
R33129 PAD.n11507 PAD.n11115 4.5005
R33130 PAD.n11509 PAD.n11115 4.5005
R33131 PAD.n11115 PAD.n11105 4.5005
R33132 PAD.n11507 PAD.n11236 4.5005
R33133 PAD.n11509 PAD.n11236 4.5005
R33134 PAD.n11236 PAD.n11105 4.5005
R33135 PAD.n11507 PAD.n11114 4.5005
R33136 PAD.n11509 PAD.n11114 4.5005
R33137 PAD.n11114 PAD.n11105 4.5005
R33138 PAD.n11507 PAD.n11238 4.5005
R33139 PAD.n11509 PAD.n11238 4.5005
R33140 PAD.n11238 PAD.n11105 4.5005
R33141 PAD.n11507 PAD.n11113 4.5005
R33142 PAD.n11509 PAD.n11113 4.5005
R33143 PAD.n11113 PAD.n11105 4.5005
R33144 PAD.n11507 PAD.n11240 4.5005
R33145 PAD.n11509 PAD.n11240 4.5005
R33146 PAD.n11240 PAD.n11105 4.5005
R33147 PAD.n11507 PAD.n11112 4.5005
R33148 PAD.n11509 PAD.n11112 4.5005
R33149 PAD.n11112 PAD.n11105 4.5005
R33150 PAD.n11507 PAD.n11242 4.5005
R33151 PAD.n11509 PAD.n11242 4.5005
R33152 PAD.n11242 PAD.n11105 4.5005
R33153 PAD.n11507 PAD.n11111 4.5005
R33154 PAD.n11509 PAD.n11111 4.5005
R33155 PAD.n11111 PAD.n11105 4.5005
R33156 PAD.n11507 PAD.n11244 4.5005
R33157 PAD.n11509 PAD.n11244 4.5005
R33158 PAD.n11244 PAD.n11105 4.5005
R33159 PAD.n11507 PAD.n11110 4.5005
R33160 PAD.n11509 PAD.n11110 4.5005
R33161 PAD.n11110 PAD.n11105 4.5005
R33162 PAD.n11507 PAD.n11246 4.5005
R33163 PAD.n11509 PAD.n11246 4.5005
R33164 PAD.n11246 PAD.n11105 4.5005
R33165 PAD.n11507 PAD.n11109 4.5005
R33166 PAD.n11509 PAD.n11109 4.5005
R33167 PAD.n11109 PAD.n11105 4.5005
R33168 PAD.n11507 PAD.n11248 4.5005
R33169 PAD.n11509 PAD.n11248 4.5005
R33170 PAD.n11248 PAD.n11105 4.5005
R33171 PAD.n11507 PAD.n11108 4.5005
R33172 PAD.n11509 PAD.n11108 4.5005
R33173 PAD.n11108 PAD.n11105 4.5005
R33174 PAD.n11507 PAD.n11250 4.5005
R33175 PAD.n11509 PAD.n11250 4.5005
R33176 PAD.n11250 PAD.n11105 4.5005
R33177 PAD.n11507 PAD.n11107 4.5005
R33178 PAD.n11509 PAD.n11107 4.5005
R33179 PAD.n11107 PAD.n11105 4.5005
R33180 PAD.n11507 PAD.n11252 4.5005
R33181 PAD.n11509 PAD.n11252 4.5005
R33182 PAD.n11252 PAD.n11105 4.5005
R33183 PAD.n11507 PAD.n11106 4.5005
R33184 PAD.n11509 PAD.n11106 4.5005
R33185 PAD.n11106 PAD.n11100 4.5005
R33186 PAD.n11106 PAD.n11105 4.5005
R33187 PAD.n5969 PAD.n5963 4.5005
R33188 PAD.n5969 PAD.n5964 4.5005
R33189 PAD.n5969 PAD.n5962 4.5005
R33190 PAD.n5969 PAD.n5965 4.5005
R33191 PAD.n6386 PAD.n5969 4.5005
R33192 PAD.n11104 PAD.n11096 4.5005
R33193 PAD.n11104 PAD.n11099 4.5005
R33194 PAD.n11513 PAD.n11104 4.5005
R33195 PAD.n6387 PAD.n5963 4.5005
R33196 PAD.n6387 PAD.n5964 4.5005
R33197 PAD.n6387 PAD.n5962 4.5005
R33198 PAD.n6387 PAD.n5965 4.5005
R33199 PAD.n6387 PAD.n6386 4.5005
R33200 PAD.n11514 PAD.n11097 4.5005
R33201 PAD.n11514 PAD.n11098 4.5005
R33202 PAD.n11514 PAD.n11096 4.5005
R33203 PAD.n11514 PAD.n11099 4.5005
R33204 PAD.n11514 PAD.n11513 4.5005
R33205 PAD.n5968 PAD.n5963 4.5005
R33206 PAD.n5968 PAD.n5964 4.5005
R33207 PAD.n5968 PAD.n5962 4.5005
R33208 PAD.n5968 PAD.n5965 4.5005
R33209 PAD.n6386 PAD.n5968 4.5005
R33210 PAD.n11102 PAD.n11097 4.5005
R33211 PAD.n11102 PAD.n11098 4.5005
R33212 PAD.n11102 PAD.n11096 4.5005
R33213 PAD.n11102 PAD.n11099 4.5005
R33214 PAD.n11513 PAD.n11102 4.5005
R33215 PAD.n6385 PAD.n5963 4.5005
R33216 PAD.n6385 PAD.n5964 4.5005
R33217 PAD.n6385 PAD.n5962 4.5005
R33218 PAD.n6385 PAD.n5965 4.5005
R33219 PAD.n6386 PAD.n6385 4.5005
R33220 PAD.n11512 PAD.n11097 4.5005
R33221 PAD.n11512 PAD.n11098 4.5005
R33222 PAD.n11512 PAD.n11096 4.5005
R33223 PAD.n11512 PAD.n11099 4.5005
R33224 PAD.n11513 PAD.n11512 4.5005
R33225 PAD.n11085 PAD.n21 4.5005
R33226 PAD.n10837 PAD.n21 4.5005
R33227 PAD.n367 PAD.n74 4.5005
R33228 PAD.n367 PAD.n366 4.5005
R33229 PAD.n10716 PAD.n415 4.5005
R33230 PAD.n10716 PAD.n10715 4.5005
R33231 PAD.n523 PAD.n435 4.5005
R33232 PAD.n770 PAD.n435 4.5005
R33233 PAD.n10388 PAD.n824 4.5005
R33234 PAD.n10388 PAD.n10387 4.5005
R33235 PAD.n10106 PAD.n1132 4.5005
R33236 PAD.n10353 PAD.n1132 4.5005
R33237 PAD.n1481 PAD.n1140 4.5005
R33238 PAD.n1294 PAD.n1140 4.5005
R33239 PAD.n9998 PAD.n1531 4.5005
R33240 PAD.n9998 PAD.n9997 4.5005
R33241 PAD.n1599 PAD.n1594 4.5005
R33242 PAD.n1685 PAD.n1594 4.5005
R33243 PAD.n9712 PAD.n1984 4.5005
R33244 PAD.n9712 PAD.n9711 4.5005
R33245 PAD.n9445 PAD.n2088 4.5005
R33246 PAD.n9445 PAD.n9444 4.5005
R33247 PAD.n2151 PAD.n2139 4.5005
R33248 PAD.n2236 PAD.n2139 4.5005
R33249 PAD.n2498 PAD.n2487 4.5005
R33250 PAD.n2583 PAD.n2487 4.5005
R33251 PAD.n9140 PAD.n2876 4.5005
R33252 PAD.n9140 PAD.n9139 4.5005
R33253 PAD.n8819 PAD.n2891 4.5005
R33254 PAD.n8570 PAD.n2891 4.5005
R33255 PAD.n8517 PAD.n2994 4.5005
R33256 PAD.n8517 PAD.n8516 4.5005
R33257 PAD.n8492 PAD.n3338 4.5005
R33258 PAD.n8492 PAD.n8491 4.5005
R33259 PAD.n8468 PAD.n3683 4.5005
R33260 PAD.n8468 PAD.n8467 4.5005
R33261 PAD.n8444 PAD.n4025 4.5005
R33262 PAD.n8444 PAD.n8443 4.5005
R33263 PAD.n4420 PAD.n4333 4.5005
R33264 PAD.n4667 PAD.n4333 4.5005
R33265 PAD.n8395 PAD.n4673 4.5005
R33266 PAD.n4832 PAD.n4673 4.5005
R33267 PAD.n4847 PAD.n4843 4.5005
R33268 PAD.n4932 PAD.n4843 4.5005
R33269 PAD.n8161 PAD.n5183 4.5005
R33270 PAD.n7971 PAD.n5183 4.5005
R33271 PAD.n5211 PAD.n5197 4.5005
R33272 PAD.n5296 PAD.n5197 4.5005
R33273 PAD.n7518 PAD.n7207 4.5005
R33274 PAD.n7269 PAD.n7207 4.5005
R33275 PAD.n7780 PAD.n7105 4.5005
R33276 PAD.n7531 PAD.n7105 4.5005
R33277 PAD.n6719 PAD.n6713 4.5005
R33278 PAD.n6804 PAD.n6713 4.5005
R33279 PAD.n5892 PAD.n5551 4.5005
R33280 PAD.n5702 PAD.n5551 4.5005
R33281 PAD.n6690 PAD.n6689 4.5005
R33282 PAD.n6689 PAD.n6688 4.5005
R33283 PAD.n6034 PAD.n5979 4.5005
R33284 PAD.n6034 PAD.n5980 4.5005
R33285 PAD.n6034 PAD.n5981 4.5005
R33286 PAD.n6373 PAD.n6034 4.5005
R33287 PAD.n6030 PAD.n5979 4.5005
R33288 PAD.n6030 PAD.n5981 4.5005
R33289 PAD.n6373 PAD.n6030 4.5005
R33290 PAD.n6037 PAD.n5979 4.5005
R33291 PAD.n6037 PAD.n5981 4.5005
R33292 PAD.n6373 PAD.n6037 4.5005
R33293 PAD.n6029 PAD.n5979 4.5005
R33294 PAD.n6029 PAD.n5981 4.5005
R33295 PAD.n6373 PAD.n6029 4.5005
R33296 PAD.n6040 PAD.n5979 4.5005
R33297 PAD.n6040 PAD.n5981 4.5005
R33298 PAD.n6373 PAD.n6040 4.5005
R33299 PAD.n6028 PAD.n5979 4.5005
R33300 PAD.n6028 PAD.n5981 4.5005
R33301 PAD.n6373 PAD.n6028 4.5005
R33302 PAD.n6043 PAD.n5979 4.5005
R33303 PAD.n6043 PAD.n5981 4.5005
R33304 PAD.n6373 PAD.n6043 4.5005
R33305 PAD.n6027 PAD.n5979 4.5005
R33306 PAD.n6027 PAD.n5981 4.5005
R33307 PAD.n6373 PAD.n6027 4.5005
R33308 PAD.n6046 PAD.n5979 4.5005
R33309 PAD.n6046 PAD.n5981 4.5005
R33310 PAD.n6373 PAD.n6046 4.5005
R33311 PAD.n6026 PAD.n5979 4.5005
R33312 PAD.n6026 PAD.n5981 4.5005
R33313 PAD.n6373 PAD.n6026 4.5005
R33314 PAD.n6049 PAD.n5979 4.5005
R33315 PAD.n6049 PAD.n5981 4.5005
R33316 PAD.n6373 PAD.n6049 4.5005
R33317 PAD.n6025 PAD.n5979 4.5005
R33318 PAD.n6025 PAD.n5981 4.5005
R33319 PAD.n6373 PAD.n6025 4.5005
R33320 PAD.n6052 PAD.n5979 4.5005
R33321 PAD.n6052 PAD.n5981 4.5005
R33322 PAD.n6373 PAD.n6052 4.5005
R33323 PAD.n6024 PAD.n5979 4.5005
R33324 PAD.n6024 PAD.n5981 4.5005
R33325 PAD.n6373 PAD.n6024 4.5005
R33326 PAD.n6055 PAD.n5979 4.5005
R33327 PAD.n6055 PAD.n5981 4.5005
R33328 PAD.n6373 PAD.n6055 4.5005
R33329 PAD.n6023 PAD.n5979 4.5005
R33330 PAD.n6023 PAD.n5981 4.5005
R33331 PAD.n6373 PAD.n6023 4.5005
R33332 PAD.n6058 PAD.n5979 4.5005
R33333 PAD.n6058 PAD.n5981 4.5005
R33334 PAD.n6373 PAD.n6058 4.5005
R33335 PAD.n6022 PAD.n5979 4.5005
R33336 PAD.n6022 PAD.n5981 4.5005
R33337 PAD.n6373 PAD.n6022 4.5005
R33338 PAD.n6061 PAD.n5979 4.5005
R33339 PAD.n6061 PAD.n5981 4.5005
R33340 PAD.n6373 PAD.n6061 4.5005
R33341 PAD.n6021 PAD.n5979 4.5005
R33342 PAD.n6021 PAD.n5981 4.5005
R33343 PAD.n6373 PAD.n6021 4.5005
R33344 PAD.n6064 PAD.n5979 4.5005
R33345 PAD.n6064 PAD.n5981 4.5005
R33346 PAD.n6373 PAD.n6064 4.5005
R33347 PAD.n6020 PAD.n5979 4.5005
R33348 PAD.n6020 PAD.n5981 4.5005
R33349 PAD.n6373 PAD.n6020 4.5005
R33350 PAD.n6067 PAD.n5979 4.5005
R33351 PAD.n6067 PAD.n5981 4.5005
R33352 PAD.n6373 PAD.n6067 4.5005
R33353 PAD.n6019 PAD.n5979 4.5005
R33354 PAD.n6019 PAD.n5981 4.5005
R33355 PAD.n6373 PAD.n6019 4.5005
R33356 PAD.n6070 PAD.n5979 4.5005
R33357 PAD.n6070 PAD.n5981 4.5005
R33358 PAD.n6373 PAD.n6070 4.5005
R33359 PAD.n6018 PAD.n5979 4.5005
R33360 PAD.n6018 PAD.n5981 4.5005
R33361 PAD.n6373 PAD.n6018 4.5005
R33362 PAD.n6073 PAD.n5979 4.5005
R33363 PAD.n6073 PAD.n5981 4.5005
R33364 PAD.n6373 PAD.n6073 4.5005
R33365 PAD.n6017 PAD.n5979 4.5005
R33366 PAD.n6017 PAD.n5981 4.5005
R33367 PAD.n6373 PAD.n6017 4.5005
R33368 PAD.n6076 PAD.n5979 4.5005
R33369 PAD.n6076 PAD.n5981 4.5005
R33370 PAD.n6373 PAD.n6076 4.5005
R33371 PAD.n6016 PAD.n5979 4.5005
R33372 PAD.n6016 PAD.n5981 4.5005
R33373 PAD.n6373 PAD.n6016 4.5005
R33374 PAD.n6079 PAD.n5979 4.5005
R33375 PAD.n6079 PAD.n5981 4.5005
R33376 PAD.n6373 PAD.n6079 4.5005
R33377 PAD.n6015 PAD.n5979 4.5005
R33378 PAD.n6015 PAD.n5981 4.5005
R33379 PAD.n6373 PAD.n6015 4.5005
R33380 PAD.n6082 PAD.n5979 4.5005
R33381 PAD.n6082 PAD.n5981 4.5005
R33382 PAD.n6373 PAD.n6082 4.5005
R33383 PAD.n6014 PAD.n5979 4.5005
R33384 PAD.n6014 PAD.n5981 4.5005
R33385 PAD.n6373 PAD.n6014 4.5005
R33386 PAD.n6085 PAD.n5979 4.5005
R33387 PAD.n6085 PAD.n5981 4.5005
R33388 PAD.n6373 PAD.n6085 4.5005
R33389 PAD.n6013 PAD.n5979 4.5005
R33390 PAD.n6013 PAD.n5981 4.5005
R33391 PAD.n6373 PAD.n6013 4.5005
R33392 PAD.n6088 PAD.n5979 4.5005
R33393 PAD.n6088 PAD.n5981 4.5005
R33394 PAD.n6373 PAD.n6088 4.5005
R33395 PAD.n6012 PAD.n5979 4.5005
R33396 PAD.n6012 PAD.n5981 4.5005
R33397 PAD.n6373 PAD.n6012 4.5005
R33398 PAD.n6091 PAD.n5979 4.5005
R33399 PAD.n6091 PAD.n5981 4.5005
R33400 PAD.n6373 PAD.n6091 4.5005
R33401 PAD.n6011 PAD.n5979 4.5005
R33402 PAD.n6011 PAD.n5981 4.5005
R33403 PAD.n6373 PAD.n6011 4.5005
R33404 PAD.n6094 PAD.n5979 4.5005
R33405 PAD.n6094 PAD.n5981 4.5005
R33406 PAD.n6373 PAD.n6094 4.5005
R33407 PAD.n6010 PAD.n5979 4.5005
R33408 PAD.n6010 PAD.n5981 4.5005
R33409 PAD.n6373 PAD.n6010 4.5005
R33410 PAD.n6097 PAD.n5979 4.5005
R33411 PAD.n6097 PAD.n5981 4.5005
R33412 PAD.n6373 PAD.n6097 4.5005
R33413 PAD.n6009 PAD.n5979 4.5005
R33414 PAD.n6009 PAD.n5981 4.5005
R33415 PAD.n6373 PAD.n6009 4.5005
R33416 PAD.n6100 PAD.n5979 4.5005
R33417 PAD.n6100 PAD.n5981 4.5005
R33418 PAD.n6373 PAD.n6100 4.5005
R33419 PAD.n6008 PAD.n5979 4.5005
R33420 PAD.n6008 PAD.n5981 4.5005
R33421 PAD.n6373 PAD.n6008 4.5005
R33422 PAD.n6103 PAD.n5979 4.5005
R33423 PAD.n6103 PAD.n5981 4.5005
R33424 PAD.n6373 PAD.n6103 4.5005
R33425 PAD.n6007 PAD.n5979 4.5005
R33426 PAD.n6007 PAD.n5981 4.5005
R33427 PAD.n6373 PAD.n6007 4.5005
R33428 PAD.n6106 PAD.n5979 4.5005
R33429 PAD.n6106 PAD.n5981 4.5005
R33430 PAD.n6373 PAD.n6106 4.5005
R33431 PAD.n6006 PAD.n5979 4.5005
R33432 PAD.n6006 PAD.n5981 4.5005
R33433 PAD.n6373 PAD.n6006 4.5005
R33434 PAD.n6109 PAD.n5979 4.5005
R33435 PAD.n6109 PAD.n5981 4.5005
R33436 PAD.n6373 PAD.n6109 4.5005
R33437 PAD.n6005 PAD.n5979 4.5005
R33438 PAD.n6005 PAD.n5981 4.5005
R33439 PAD.n6373 PAD.n6005 4.5005
R33440 PAD.n6112 PAD.n5979 4.5005
R33441 PAD.n6112 PAD.n5981 4.5005
R33442 PAD.n6373 PAD.n6112 4.5005
R33443 PAD.n6004 PAD.n5979 4.5005
R33444 PAD.n6004 PAD.n5981 4.5005
R33445 PAD.n6373 PAD.n6004 4.5005
R33446 PAD.n6115 PAD.n5979 4.5005
R33447 PAD.n6115 PAD.n5981 4.5005
R33448 PAD.n6373 PAD.n6115 4.5005
R33449 PAD.n6003 PAD.n5979 4.5005
R33450 PAD.n6003 PAD.n5981 4.5005
R33451 PAD.n6373 PAD.n6003 4.5005
R33452 PAD.n6118 PAD.n5979 4.5005
R33453 PAD.n6118 PAD.n5981 4.5005
R33454 PAD.n6373 PAD.n6118 4.5005
R33455 PAD.n6002 PAD.n5979 4.5005
R33456 PAD.n6002 PAD.n5981 4.5005
R33457 PAD.n6373 PAD.n6002 4.5005
R33458 PAD.n6121 PAD.n5979 4.5005
R33459 PAD.n6121 PAD.n5981 4.5005
R33460 PAD.n6373 PAD.n6121 4.5005
R33461 PAD.n6001 PAD.n5979 4.5005
R33462 PAD.n6001 PAD.n5981 4.5005
R33463 PAD.n6373 PAD.n6001 4.5005
R33464 PAD.n6124 PAD.n5979 4.5005
R33465 PAD.n6124 PAD.n5981 4.5005
R33466 PAD.n6373 PAD.n6124 4.5005
R33467 PAD.n6000 PAD.n5979 4.5005
R33468 PAD.n6000 PAD.n5981 4.5005
R33469 PAD.n6373 PAD.n6000 4.5005
R33470 PAD.n6127 PAD.n5979 4.5005
R33471 PAD.n6127 PAD.n5981 4.5005
R33472 PAD.n6373 PAD.n6127 4.5005
R33473 PAD.n5999 PAD.n5979 4.5005
R33474 PAD.n5999 PAD.n5981 4.5005
R33475 PAD.n6373 PAD.n5999 4.5005
R33476 PAD.n6130 PAD.n5979 4.5005
R33477 PAD.n6130 PAD.n5981 4.5005
R33478 PAD.n6373 PAD.n6130 4.5005
R33479 PAD.n5998 PAD.n5979 4.5005
R33480 PAD.n5998 PAD.n5981 4.5005
R33481 PAD.n6373 PAD.n5998 4.5005
R33482 PAD.n6133 PAD.n5979 4.5005
R33483 PAD.n6133 PAD.n5981 4.5005
R33484 PAD.n6373 PAD.n6133 4.5005
R33485 PAD.n5997 PAD.n5979 4.5005
R33486 PAD.n5997 PAD.n5981 4.5005
R33487 PAD.n6373 PAD.n5997 4.5005
R33488 PAD.n6136 PAD.n5979 4.5005
R33489 PAD.n6136 PAD.n5981 4.5005
R33490 PAD.n6373 PAD.n6136 4.5005
R33491 PAD.n5996 PAD.n5979 4.5005
R33492 PAD.n5996 PAD.n5981 4.5005
R33493 PAD.n6373 PAD.n5996 4.5005
R33494 PAD.n6139 PAD.n5979 4.5005
R33495 PAD.n6139 PAD.n5981 4.5005
R33496 PAD.n6373 PAD.n6139 4.5005
R33497 PAD.n5995 PAD.n5979 4.5005
R33498 PAD.n5995 PAD.n5981 4.5005
R33499 PAD.n6373 PAD.n5995 4.5005
R33500 PAD.n6142 PAD.n5979 4.5005
R33501 PAD.n6142 PAD.n5981 4.5005
R33502 PAD.n6373 PAD.n6142 4.5005
R33503 PAD.n5994 PAD.n5979 4.5005
R33504 PAD.n5994 PAD.n5981 4.5005
R33505 PAD.n6373 PAD.n5994 4.5005
R33506 PAD.n6145 PAD.n5979 4.5005
R33507 PAD.n6145 PAD.n5981 4.5005
R33508 PAD.n6373 PAD.n6145 4.5005
R33509 PAD.n5993 PAD.n5979 4.5005
R33510 PAD.n5993 PAD.n5981 4.5005
R33511 PAD.n6373 PAD.n5993 4.5005
R33512 PAD.n6148 PAD.n5979 4.5005
R33513 PAD.n6148 PAD.n5981 4.5005
R33514 PAD.n6373 PAD.n6148 4.5005
R33515 PAD.n5992 PAD.n5979 4.5005
R33516 PAD.n5992 PAD.n5981 4.5005
R33517 PAD.n6373 PAD.n5992 4.5005
R33518 PAD.n6151 PAD.n5979 4.5005
R33519 PAD.n6151 PAD.n5981 4.5005
R33520 PAD.n6373 PAD.n6151 4.5005
R33521 PAD.n5991 PAD.n5979 4.5005
R33522 PAD.n5991 PAD.n5981 4.5005
R33523 PAD.n6373 PAD.n5991 4.5005
R33524 PAD.n6154 PAD.n5979 4.5005
R33525 PAD.n6154 PAD.n5981 4.5005
R33526 PAD.n6373 PAD.n6154 4.5005
R33527 PAD.n5990 PAD.n5979 4.5005
R33528 PAD.n5990 PAD.n5981 4.5005
R33529 PAD.n6373 PAD.n5990 4.5005
R33530 PAD.n6157 PAD.n5979 4.5005
R33531 PAD.n6157 PAD.n5981 4.5005
R33532 PAD.n6373 PAD.n6157 4.5005
R33533 PAD.n5989 PAD.n5979 4.5005
R33534 PAD.n5989 PAD.n5981 4.5005
R33535 PAD.n6373 PAD.n5989 4.5005
R33536 PAD.n6160 PAD.n5979 4.5005
R33537 PAD.n6160 PAD.n5981 4.5005
R33538 PAD.n6373 PAD.n6160 4.5005
R33539 PAD.n5988 PAD.n5979 4.5005
R33540 PAD.n5988 PAD.n5981 4.5005
R33541 PAD.n6373 PAD.n5988 4.5005
R33542 PAD.n6163 PAD.n5979 4.5005
R33543 PAD.n6163 PAD.n5981 4.5005
R33544 PAD.n6373 PAD.n6163 4.5005
R33545 PAD.n5987 PAD.n5979 4.5005
R33546 PAD.n5987 PAD.n5981 4.5005
R33547 PAD.n6373 PAD.n5987 4.5005
R33548 PAD.n6166 PAD.n5979 4.5005
R33549 PAD.n6166 PAD.n5981 4.5005
R33550 PAD.n6373 PAD.n6166 4.5005
R33551 PAD.n5986 PAD.n5979 4.5005
R33552 PAD.n5986 PAD.n5981 4.5005
R33553 PAD.n6373 PAD.n5986 4.5005
R33554 PAD.n6169 PAD.n5979 4.5005
R33555 PAD.n6169 PAD.n5981 4.5005
R33556 PAD.n6373 PAD.n6169 4.5005
R33557 PAD.n5985 PAD.n5979 4.5005
R33558 PAD.n5985 PAD.n5981 4.5005
R33559 PAD.n6373 PAD.n5985 4.5005
R33560 PAD.n6172 PAD.n5979 4.5005
R33561 PAD.n6172 PAD.n5981 4.5005
R33562 PAD.n6373 PAD.n6172 4.5005
R33563 PAD.n5984 PAD.n5979 4.5005
R33564 PAD.n5984 PAD.n5981 4.5005
R33565 PAD.n6373 PAD.n5984 4.5005
R33566 PAD.n6175 PAD.n5979 4.5005
R33567 PAD.n6175 PAD.n5981 4.5005
R33568 PAD.n6373 PAD.n6175 4.5005
R33569 PAD.n5983 PAD.n5979 4.5005
R33570 PAD.n5983 PAD.n5981 4.5005
R33571 PAD.n6373 PAD.n5983 4.5005
R33572 PAD.n6372 PAD.n5979 4.5005
R33573 PAD.n6372 PAD.n5980 4.5005
R33574 PAD.n6372 PAD.n5981 4.5005
R33575 PAD.n6373 PAD.n6372 4.5005
R33576 PAD.n11508 PAD.n11105 4.5005
R33577 PAD.n11508 PAD.n11100 4.5005
R33578 PAD.n11509 PAD.n11508 4.5005
R33579 PAD.n11508 PAD.n11302 4.5005
R33580 PAD.n11508 PAD.n11507 4.5005
R33581 PAD.n6374 PAD.n5979 4.5005
R33582 PAD.n4 PAD 4.06833
R33583 PAD.n2 PAD.n1 3.98767
R33584 PAD.n8 PAD.n7 3.98767
R33585 PAD.n7808 PAD.n7807 2.64618
R33586 PAD.n3 PAD.n2 2.64417
R33587 PAD.n7 PAD.n6 2.64417
R33588 PAD.n5 PAD.n4 2.64417
R33589 PAD.n0 PAD.t21 2.55406
R33590 PAD.n11539 PAD.n11538 2.52597
R33591 PAD.n11104 PAD.n11103 2.25086
R33592 PAD.n7518 PAD.n7517 2.2505
R33593 PAD.n7209 PAD.n7201 2.2505
R33594 PAD.n7513 PAD.n7512 2.2505
R33595 PAD.n7510 PAD.n7509 2.2505
R33596 PAD.n7507 PAD.n7506 2.2505
R33597 PAD.n7499 PAD.n7229 2.2505
R33598 PAD.n7502 PAD.n7501 2.2505
R33599 PAD.n7498 PAD.n7497 2.2505
R33600 PAD.n7495 PAD.n7494 2.2505
R33601 PAD.n7487 PAD.n7231 2.2505
R33602 PAD.n7490 PAD.n7489 2.2505
R33603 PAD.n7486 PAD.n7485 2.2505
R33604 PAD.n7483 PAD.n7482 2.2505
R33605 PAD.n7475 PAD.n7233 2.2505
R33606 PAD.n7478 PAD.n7477 2.2505
R33607 PAD.n7474 PAD.n7473 2.2505
R33608 PAD.n7471 PAD.n7470 2.2505
R33609 PAD.n7463 PAD.n7235 2.2505
R33610 PAD.n7466 PAD.n7465 2.2505
R33611 PAD.n7462 PAD.n7461 2.2505
R33612 PAD.n7459 PAD.n7458 2.2505
R33613 PAD.n7451 PAD.n7237 2.2505
R33614 PAD.n7454 PAD.n7453 2.2505
R33615 PAD.n7450 PAD.n7449 2.2505
R33616 PAD.n7447 PAD.n7446 2.2505
R33617 PAD.n7439 PAD.n7239 2.2505
R33618 PAD.n7442 PAD.n7441 2.2505
R33619 PAD.n7438 PAD.n7437 2.2505
R33620 PAD.n7435 PAD.n7434 2.2505
R33621 PAD.n7427 PAD.n7241 2.2505
R33622 PAD.n7430 PAD.n7429 2.2505
R33623 PAD.n7426 PAD.n7425 2.2505
R33624 PAD.n7423 PAD.n7422 2.2505
R33625 PAD.n7415 PAD.n7243 2.2505
R33626 PAD.n7418 PAD.n7417 2.2505
R33627 PAD.n7414 PAD.n7413 2.2505
R33628 PAD.n7411 PAD.n7410 2.2505
R33629 PAD.n7403 PAD.n7245 2.2505
R33630 PAD.n7406 PAD.n7405 2.2505
R33631 PAD.n7402 PAD.n7401 2.2505
R33632 PAD.n7399 PAD.n7398 2.2505
R33633 PAD.n7391 PAD.n7247 2.2505
R33634 PAD.n7394 PAD.n7393 2.2505
R33635 PAD.n7390 PAD.n7389 2.2505
R33636 PAD.n7387 PAD.n7386 2.2505
R33637 PAD.n7379 PAD.n7249 2.2505
R33638 PAD.n7382 PAD.n7381 2.2505
R33639 PAD.n7378 PAD.n7377 2.2505
R33640 PAD.n7375 PAD.n7374 2.2505
R33641 PAD.n7367 PAD.n7251 2.2505
R33642 PAD.n7370 PAD.n7369 2.2505
R33643 PAD.n7366 PAD.n7365 2.2505
R33644 PAD.n7363 PAD.n7362 2.2505
R33645 PAD.n7355 PAD.n7253 2.2505
R33646 PAD.n7358 PAD.n7357 2.2505
R33647 PAD.n7354 PAD.n7353 2.2505
R33648 PAD.n7351 PAD.n7350 2.2505
R33649 PAD.n7343 PAD.n7255 2.2505
R33650 PAD.n7346 PAD.n7345 2.2505
R33651 PAD.n7342 PAD.n7341 2.2505
R33652 PAD.n7339 PAD.n7338 2.2505
R33653 PAD.n7331 PAD.n7257 2.2505
R33654 PAD.n7334 PAD.n7333 2.2505
R33655 PAD.n7330 PAD.n7329 2.2505
R33656 PAD.n7327 PAD.n7326 2.2505
R33657 PAD.n7319 PAD.n7259 2.2505
R33658 PAD.n7322 PAD.n7321 2.2505
R33659 PAD.n7318 PAD.n7317 2.2505
R33660 PAD.n7315 PAD.n7314 2.2505
R33661 PAD.n7307 PAD.n7261 2.2505
R33662 PAD.n7310 PAD.n7309 2.2505
R33663 PAD.n7306 PAD.n7305 2.2505
R33664 PAD.n7303 PAD.n7302 2.2505
R33665 PAD.n7295 PAD.n7263 2.2505
R33666 PAD.n7298 PAD.n7297 2.2505
R33667 PAD.n7294 PAD.n7293 2.2505
R33668 PAD.n7291 PAD.n7290 2.2505
R33669 PAD.n7283 PAD.n7265 2.2505
R33670 PAD.n7286 PAD.n7285 2.2505
R33671 PAD.n7282 PAD.n7281 2.2505
R33672 PAD.n7279 PAD.n7278 2.2505
R33673 PAD.n7271 PAD.n7267 2.2505
R33674 PAD.n7274 PAD.n7273 2.2505
R33675 PAD.n7270 PAD.n7269 2.2505
R33676 PAD.n7270 PAD.n7268 2.2505
R33677 PAD.n7275 PAD.n7274 2.2505
R33678 PAD.n7276 PAD.n7267 2.2505
R33679 PAD.n7278 PAD.n7277 2.2505
R33680 PAD.n7282 PAD.n7266 2.2505
R33681 PAD.n7287 PAD.n7286 2.2505
R33682 PAD.n7288 PAD.n7265 2.2505
R33683 PAD.n7290 PAD.n7289 2.2505
R33684 PAD.n7294 PAD.n7264 2.2505
R33685 PAD.n7299 PAD.n7298 2.2505
R33686 PAD.n7300 PAD.n7263 2.2505
R33687 PAD.n7302 PAD.n7301 2.2505
R33688 PAD.n7306 PAD.n7262 2.2505
R33689 PAD.n7311 PAD.n7310 2.2505
R33690 PAD.n7312 PAD.n7261 2.2505
R33691 PAD.n7314 PAD.n7313 2.2505
R33692 PAD.n7318 PAD.n7260 2.2505
R33693 PAD.n7323 PAD.n7322 2.2505
R33694 PAD.n7324 PAD.n7259 2.2505
R33695 PAD.n7326 PAD.n7325 2.2505
R33696 PAD.n7330 PAD.n7258 2.2505
R33697 PAD.n7335 PAD.n7334 2.2505
R33698 PAD.n7336 PAD.n7257 2.2505
R33699 PAD.n7338 PAD.n7337 2.2505
R33700 PAD.n7342 PAD.n7256 2.2505
R33701 PAD.n7347 PAD.n7346 2.2505
R33702 PAD.n7348 PAD.n7255 2.2505
R33703 PAD.n7350 PAD.n7349 2.2505
R33704 PAD.n7354 PAD.n7254 2.2505
R33705 PAD.n7359 PAD.n7358 2.2505
R33706 PAD.n7360 PAD.n7253 2.2505
R33707 PAD.n7362 PAD.n7361 2.2505
R33708 PAD.n7366 PAD.n7252 2.2505
R33709 PAD.n7371 PAD.n7370 2.2505
R33710 PAD.n7372 PAD.n7251 2.2505
R33711 PAD.n7374 PAD.n7373 2.2505
R33712 PAD.n7378 PAD.n7250 2.2505
R33713 PAD.n7383 PAD.n7382 2.2505
R33714 PAD.n7384 PAD.n7249 2.2505
R33715 PAD.n7386 PAD.n7385 2.2505
R33716 PAD.n7390 PAD.n7248 2.2505
R33717 PAD.n7395 PAD.n7394 2.2505
R33718 PAD.n7396 PAD.n7247 2.2505
R33719 PAD.n7398 PAD.n7397 2.2505
R33720 PAD.n7402 PAD.n7246 2.2505
R33721 PAD.n7407 PAD.n7406 2.2505
R33722 PAD.n7408 PAD.n7245 2.2505
R33723 PAD.n7410 PAD.n7409 2.2505
R33724 PAD.n7414 PAD.n7244 2.2505
R33725 PAD.n7419 PAD.n7418 2.2505
R33726 PAD.n7420 PAD.n7243 2.2505
R33727 PAD.n7422 PAD.n7421 2.2505
R33728 PAD.n7426 PAD.n7242 2.2505
R33729 PAD.n7431 PAD.n7430 2.2505
R33730 PAD.n7432 PAD.n7241 2.2505
R33731 PAD.n7434 PAD.n7433 2.2505
R33732 PAD.n7438 PAD.n7240 2.2505
R33733 PAD.n7443 PAD.n7442 2.2505
R33734 PAD.n7444 PAD.n7239 2.2505
R33735 PAD.n7446 PAD.n7445 2.2505
R33736 PAD.n7450 PAD.n7238 2.2505
R33737 PAD.n7455 PAD.n7454 2.2505
R33738 PAD.n7456 PAD.n7237 2.2505
R33739 PAD.n7458 PAD.n7457 2.2505
R33740 PAD.n7462 PAD.n7236 2.2505
R33741 PAD.n7467 PAD.n7466 2.2505
R33742 PAD.n7468 PAD.n7235 2.2505
R33743 PAD.n7470 PAD.n7469 2.2505
R33744 PAD.n7474 PAD.n7234 2.2505
R33745 PAD.n7479 PAD.n7478 2.2505
R33746 PAD.n7480 PAD.n7233 2.2505
R33747 PAD.n7482 PAD.n7481 2.2505
R33748 PAD.n7486 PAD.n7232 2.2505
R33749 PAD.n7491 PAD.n7490 2.2505
R33750 PAD.n7492 PAD.n7231 2.2505
R33751 PAD.n7494 PAD.n7493 2.2505
R33752 PAD.n7498 PAD.n7230 2.2505
R33753 PAD.n7503 PAD.n7502 2.2505
R33754 PAD.n7504 PAD.n7229 2.2505
R33755 PAD.n7506 PAD.n7505 2.2505
R33756 PAD.n7510 PAD.n7228 2.2505
R33757 PAD.n7514 PAD.n7513 2.2505
R33758 PAD.n7515 PAD.n7209 2.2505
R33759 PAD.n7517 PAD.n7516 2.2505
R33760 PAD.n10695 PAD.n415 2.2505
R33761 PAD.n10694 PAD.n10693 2.2505
R33762 PAD.n10691 PAD.n10417 2.2505
R33763 PAD.n10415 PAD.n10414 2.2505
R33764 PAD.n10687 PAD.n10686 2.2505
R33765 PAD.n10684 PAD.n10683 2.2505
R33766 PAD.n10682 PAD.n10422 2.2505
R33767 PAD.n10420 PAD.n10419 2.2505
R33768 PAD.n10678 PAD.n10677 2.2505
R33769 PAD.n10675 PAD.n10674 2.2505
R33770 PAD.n10673 PAD.n10427 2.2505
R33771 PAD.n10425 PAD.n10424 2.2505
R33772 PAD.n10669 PAD.n10668 2.2505
R33773 PAD.n10666 PAD.n10665 2.2505
R33774 PAD.n10664 PAD.n10432 2.2505
R33775 PAD.n10430 PAD.n10429 2.2505
R33776 PAD.n10660 PAD.n10659 2.2505
R33777 PAD.n10657 PAD.n10656 2.2505
R33778 PAD.n10655 PAD.n10437 2.2505
R33779 PAD.n10435 PAD.n10434 2.2505
R33780 PAD.n10651 PAD.n10650 2.2505
R33781 PAD.n10648 PAD.n10647 2.2505
R33782 PAD.n10646 PAD.n10442 2.2505
R33783 PAD.n10440 PAD.n10439 2.2505
R33784 PAD.n10642 PAD.n10641 2.2505
R33785 PAD.n10639 PAD.n10638 2.2505
R33786 PAD.n10637 PAD.n10447 2.2505
R33787 PAD.n10445 PAD.n10444 2.2505
R33788 PAD.n10633 PAD.n10632 2.2505
R33789 PAD.n10630 PAD.n10629 2.2505
R33790 PAD.n10628 PAD.n10452 2.2505
R33791 PAD.n10450 PAD.n10449 2.2505
R33792 PAD.n10624 PAD.n10623 2.2505
R33793 PAD.n10621 PAD.n10620 2.2505
R33794 PAD.n10619 PAD.n10457 2.2505
R33795 PAD.n10455 PAD.n10454 2.2505
R33796 PAD.n10615 PAD.n10614 2.2505
R33797 PAD.n10612 PAD.n10611 2.2505
R33798 PAD.n10610 PAD.n10462 2.2505
R33799 PAD.n10460 PAD.n10459 2.2505
R33800 PAD.n10606 PAD.n10605 2.2505
R33801 PAD.n10603 PAD.n10602 2.2505
R33802 PAD.n10601 PAD.n10467 2.2505
R33803 PAD.n10465 PAD.n10464 2.2505
R33804 PAD.n10597 PAD.n10596 2.2505
R33805 PAD.n10594 PAD.n10593 2.2505
R33806 PAD.n10592 PAD.n10472 2.2505
R33807 PAD.n10470 PAD.n10469 2.2505
R33808 PAD.n10588 PAD.n10587 2.2505
R33809 PAD.n10585 PAD.n10584 2.2505
R33810 PAD.n10583 PAD.n10477 2.2505
R33811 PAD.n10475 PAD.n10474 2.2505
R33812 PAD.n10579 PAD.n10578 2.2505
R33813 PAD.n10576 PAD.n10575 2.2505
R33814 PAD.n10574 PAD.n10482 2.2505
R33815 PAD.n10480 PAD.n10479 2.2505
R33816 PAD.n10570 PAD.n10569 2.2505
R33817 PAD.n10567 PAD.n10566 2.2505
R33818 PAD.n10565 PAD.n10487 2.2505
R33819 PAD.n10485 PAD.n10484 2.2505
R33820 PAD.n10561 PAD.n10560 2.2505
R33821 PAD.n10558 PAD.n10557 2.2505
R33822 PAD.n10556 PAD.n10492 2.2505
R33823 PAD.n10490 PAD.n10489 2.2505
R33824 PAD.n10552 PAD.n10551 2.2505
R33825 PAD.n10549 PAD.n10548 2.2505
R33826 PAD.n10547 PAD.n10497 2.2505
R33827 PAD.n10495 PAD.n10494 2.2505
R33828 PAD.n10543 PAD.n10542 2.2505
R33829 PAD.n10540 PAD.n10539 2.2505
R33830 PAD.n10538 PAD.n10502 2.2505
R33831 PAD.n10500 PAD.n10499 2.2505
R33832 PAD.n10534 PAD.n10533 2.2505
R33833 PAD.n10531 PAD.n10530 2.2505
R33834 PAD.n10529 PAD.n10507 2.2505
R33835 PAD.n10505 PAD.n10504 2.2505
R33836 PAD.n10525 PAD.n10524 2.2505
R33837 PAD.n10522 PAD.n10521 2.2505
R33838 PAD.n10520 PAD.n10512 2.2505
R33839 PAD.n10510 PAD.n10509 2.2505
R33840 PAD.n10516 PAD.n10515 2.2505
R33841 PAD.n10513 PAD.n420 2.2505
R33842 PAD.n10713 PAD.n10712 2.2505
R33843 PAD.n10715 PAD.n416 2.2505
R33844 PAD.n10710 PAD.n416 2.2505
R33845 PAD.n10712 PAD.n10711 2.2505
R33846 PAD.n421 PAD.n420 2.2505
R33847 PAD.n10517 PAD.n10516 2.2505
R33848 PAD.n10518 PAD.n10509 2.2505
R33849 PAD.n10520 PAD.n10519 2.2505
R33850 PAD.n10521 PAD.n10508 2.2505
R33851 PAD.n10526 PAD.n10525 2.2505
R33852 PAD.n10527 PAD.n10504 2.2505
R33853 PAD.n10529 PAD.n10528 2.2505
R33854 PAD.n10530 PAD.n10503 2.2505
R33855 PAD.n10535 PAD.n10534 2.2505
R33856 PAD.n10536 PAD.n10499 2.2505
R33857 PAD.n10538 PAD.n10537 2.2505
R33858 PAD.n10539 PAD.n10498 2.2505
R33859 PAD.n10544 PAD.n10543 2.2505
R33860 PAD.n10545 PAD.n10494 2.2505
R33861 PAD.n10547 PAD.n10546 2.2505
R33862 PAD.n10548 PAD.n10493 2.2505
R33863 PAD.n10553 PAD.n10552 2.2505
R33864 PAD.n10554 PAD.n10489 2.2505
R33865 PAD.n10556 PAD.n10555 2.2505
R33866 PAD.n10557 PAD.n10488 2.2505
R33867 PAD.n10562 PAD.n10561 2.2505
R33868 PAD.n10563 PAD.n10484 2.2505
R33869 PAD.n10565 PAD.n10564 2.2505
R33870 PAD.n10566 PAD.n10483 2.2505
R33871 PAD.n10571 PAD.n10570 2.2505
R33872 PAD.n10572 PAD.n10479 2.2505
R33873 PAD.n10574 PAD.n10573 2.2505
R33874 PAD.n10575 PAD.n10478 2.2505
R33875 PAD.n10580 PAD.n10579 2.2505
R33876 PAD.n10581 PAD.n10474 2.2505
R33877 PAD.n10583 PAD.n10582 2.2505
R33878 PAD.n10584 PAD.n10473 2.2505
R33879 PAD.n10589 PAD.n10588 2.2505
R33880 PAD.n10590 PAD.n10469 2.2505
R33881 PAD.n10592 PAD.n10591 2.2505
R33882 PAD.n10593 PAD.n10468 2.2505
R33883 PAD.n10598 PAD.n10597 2.2505
R33884 PAD.n10599 PAD.n10464 2.2505
R33885 PAD.n10601 PAD.n10600 2.2505
R33886 PAD.n10602 PAD.n10463 2.2505
R33887 PAD.n10607 PAD.n10606 2.2505
R33888 PAD.n10608 PAD.n10459 2.2505
R33889 PAD.n10610 PAD.n10609 2.2505
R33890 PAD.n10611 PAD.n10458 2.2505
R33891 PAD.n10616 PAD.n10615 2.2505
R33892 PAD.n10617 PAD.n10454 2.2505
R33893 PAD.n10619 PAD.n10618 2.2505
R33894 PAD.n10620 PAD.n10453 2.2505
R33895 PAD.n10625 PAD.n10624 2.2505
R33896 PAD.n10626 PAD.n10449 2.2505
R33897 PAD.n10628 PAD.n10627 2.2505
R33898 PAD.n10629 PAD.n10448 2.2505
R33899 PAD.n10634 PAD.n10633 2.2505
R33900 PAD.n10635 PAD.n10444 2.2505
R33901 PAD.n10637 PAD.n10636 2.2505
R33902 PAD.n10638 PAD.n10443 2.2505
R33903 PAD.n10643 PAD.n10642 2.2505
R33904 PAD.n10644 PAD.n10439 2.2505
R33905 PAD.n10646 PAD.n10645 2.2505
R33906 PAD.n10647 PAD.n10438 2.2505
R33907 PAD.n10652 PAD.n10651 2.2505
R33908 PAD.n10653 PAD.n10434 2.2505
R33909 PAD.n10655 PAD.n10654 2.2505
R33910 PAD.n10656 PAD.n10433 2.2505
R33911 PAD.n10661 PAD.n10660 2.2505
R33912 PAD.n10662 PAD.n10429 2.2505
R33913 PAD.n10664 PAD.n10663 2.2505
R33914 PAD.n10665 PAD.n10428 2.2505
R33915 PAD.n10670 PAD.n10669 2.2505
R33916 PAD.n10671 PAD.n10424 2.2505
R33917 PAD.n10673 PAD.n10672 2.2505
R33918 PAD.n10674 PAD.n10423 2.2505
R33919 PAD.n10679 PAD.n10678 2.2505
R33920 PAD.n10680 PAD.n10419 2.2505
R33921 PAD.n10682 PAD.n10681 2.2505
R33922 PAD.n10683 PAD.n10418 2.2505
R33923 PAD.n10688 PAD.n10687 2.2505
R33924 PAD.n10689 PAD.n10414 2.2505
R33925 PAD.n10691 PAD.n10690 2.2505
R33926 PAD.n10694 PAD.n10413 2.2505
R33927 PAD.n10696 PAD.n10695 2.2505
R33928 PAD.n523 PAD.n522 2.2505
R33929 PAD.n525 PAD.n520 2.2505
R33930 PAD.n530 PAD.n529 2.2505
R33931 PAD.n527 PAD.n518 2.2505
R33932 PAD.n535 PAD.n534 2.2505
R33933 PAD.n537 PAD.n516 2.2505
R33934 PAD.n542 PAD.n541 2.2505
R33935 PAD.n539 PAD.n514 2.2505
R33936 PAD.n547 PAD.n546 2.2505
R33937 PAD.n549 PAD.n512 2.2505
R33938 PAD.n554 PAD.n553 2.2505
R33939 PAD.n551 PAD.n510 2.2505
R33940 PAD.n559 PAD.n558 2.2505
R33941 PAD.n561 PAD.n508 2.2505
R33942 PAD.n566 PAD.n565 2.2505
R33943 PAD.n563 PAD.n506 2.2505
R33944 PAD.n571 PAD.n570 2.2505
R33945 PAD.n573 PAD.n504 2.2505
R33946 PAD.n578 PAD.n577 2.2505
R33947 PAD.n575 PAD.n502 2.2505
R33948 PAD.n583 PAD.n582 2.2505
R33949 PAD.n585 PAD.n500 2.2505
R33950 PAD.n590 PAD.n589 2.2505
R33951 PAD.n587 PAD.n498 2.2505
R33952 PAD.n595 PAD.n594 2.2505
R33953 PAD.n597 PAD.n496 2.2505
R33954 PAD.n602 PAD.n601 2.2505
R33955 PAD.n599 PAD.n494 2.2505
R33956 PAD.n607 PAD.n606 2.2505
R33957 PAD.n609 PAD.n492 2.2505
R33958 PAD.n614 PAD.n613 2.2505
R33959 PAD.n611 PAD.n490 2.2505
R33960 PAD.n619 PAD.n618 2.2505
R33961 PAD.n621 PAD.n488 2.2505
R33962 PAD.n626 PAD.n625 2.2505
R33963 PAD.n623 PAD.n486 2.2505
R33964 PAD.n631 PAD.n630 2.2505
R33965 PAD.n633 PAD.n484 2.2505
R33966 PAD.n638 PAD.n637 2.2505
R33967 PAD.n635 PAD.n482 2.2505
R33968 PAD.n643 PAD.n642 2.2505
R33969 PAD.n645 PAD.n480 2.2505
R33970 PAD.n650 PAD.n649 2.2505
R33971 PAD.n647 PAD.n478 2.2505
R33972 PAD.n655 PAD.n654 2.2505
R33973 PAD.n657 PAD.n476 2.2505
R33974 PAD.n662 PAD.n661 2.2505
R33975 PAD.n659 PAD.n474 2.2505
R33976 PAD.n667 PAD.n666 2.2505
R33977 PAD.n669 PAD.n472 2.2505
R33978 PAD.n674 PAD.n673 2.2505
R33979 PAD.n671 PAD.n470 2.2505
R33980 PAD.n679 PAD.n678 2.2505
R33981 PAD.n681 PAD.n468 2.2505
R33982 PAD.n686 PAD.n685 2.2505
R33983 PAD.n683 PAD.n466 2.2505
R33984 PAD.n691 PAD.n690 2.2505
R33985 PAD.n693 PAD.n464 2.2505
R33986 PAD.n698 PAD.n697 2.2505
R33987 PAD.n695 PAD.n462 2.2505
R33988 PAD.n703 PAD.n702 2.2505
R33989 PAD.n705 PAD.n460 2.2505
R33990 PAD.n710 PAD.n709 2.2505
R33991 PAD.n707 PAD.n458 2.2505
R33992 PAD.n715 PAD.n714 2.2505
R33993 PAD.n717 PAD.n456 2.2505
R33994 PAD.n722 PAD.n721 2.2505
R33995 PAD.n719 PAD.n454 2.2505
R33996 PAD.n727 PAD.n726 2.2505
R33997 PAD.n729 PAD.n452 2.2505
R33998 PAD.n734 PAD.n733 2.2505
R33999 PAD.n731 PAD.n450 2.2505
R34000 PAD.n739 PAD.n738 2.2505
R34001 PAD.n741 PAD.n448 2.2505
R34002 PAD.n746 PAD.n745 2.2505
R34003 PAD.n743 PAD.n446 2.2505
R34004 PAD.n751 PAD.n750 2.2505
R34005 PAD.n753 PAD.n444 2.2505
R34006 PAD.n758 PAD.n757 2.2505
R34007 PAD.n755 PAD.n442 2.2505
R34008 PAD.n764 PAD.n763 2.2505
R34009 PAD.n766 PAD.n440 2.2505
R34010 PAD.n768 PAD.n439 2.2505
R34011 PAD.n771 PAD.n770 2.2505
R34012 PAD.n772 PAD.n771 2.2505
R34013 PAD.n439 PAD.n438 2.2505
R34014 PAD.n761 PAD.n440 2.2505
R34015 PAD.n763 PAD.n762 2.2505
R34016 PAD.n760 PAD.n442 2.2505
R34017 PAD.n759 PAD.n758 2.2505
R34018 PAD.n444 PAD.n443 2.2505
R34019 PAD.n750 PAD.n749 2.2505
R34020 PAD.n748 PAD.n446 2.2505
R34021 PAD.n747 PAD.n746 2.2505
R34022 PAD.n448 PAD.n447 2.2505
R34023 PAD.n738 PAD.n737 2.2505
R34024 PAD.n736 PAD.n450 2.2505
R34025 PAD.n735 PAD.n734 2.2505
R34026 PAD.n452 PAD.n451 2.2505
R34027 PAD.n726 PAD.n725 2.2505
R34028 PAD.n724 PAD.n454 2.2505
R34029 PAD.n723 PAD.n722 2.2505
R34030 PAD.n456 PAD.n455 2.2505
R34031 PAD.n714 PAD.n713 2.2505
R34032 PAD.n712 PAD.n458 2.2505
R34033 PAD.n711 PAD.n710 2.2505
R34034 PAD.n460 PAD.n459 2.2505
R34035 PAD.n702 PAD.n701 2.2505
R34036 PAD.n700 PAD.n462 2.2505
R34037 PAD.n699 PAD.n698 2.2505
R34038 PAD.n464 PAD.n463 2.2505
R34039 PAD.n690 PAD.n689 2.2505
R34040 PAD.n688 PAD.n466 2.2505
R34041 PAD.n687 PAD.n686 2.2505
R34042 PAD.n468 PAD.n467 2.2505
R34043 PAD.n678 PAD.n677 2.2505
R34044 PAD.n676 PAD.n470 2.2505
R34045 PAD.n675 PAD.n674 2.2505
R34046 PAD.n472 PAD.n471 2.2505
R34047 PAD.n666 PAD.n665 2.2505
R34048 PAD.n664 PAD.n474 2.2505
R34049 PAD.n663 PAD.n662 2.2505
R34050 PAD.n476 PAD.n475 2.2505
R34051 PAD.n654 PAD.n653 2.2505
R34052 PAD.n652 PAD.n478 2.2505
R34053 PAD.n651 PAD.n650 2.2505
R34054 PAD.n480 PAD.n479 2.2505
R34055 PAD.n642 PAD.n641 2.2505
R34056 PAD.n640 PAD.n482 2.2505
R34057 PAD.n639 PAD.n638 2.2505
R34058 PAD.n484 PAD.n483 2.2505
R34059 PAD.n630 PAD.n629 2.2505
R34060 PAD.n628 PAD.n486 2.2505
R34061 PAD.n627 PAD.n626 2.2505
R34062 PAD.n488 PAD.n487 2.2505
R34063 PAD.n618 PAD.n617 2.2505
R34064 PAD.n616 PAD.n490 2.2505
R34065 PAD.n615 PAD.n614 2.2505
R34066 PAD.n492 PAD.n491 2.2505
R34067 PAD.n606 PAD.n605 2.2505
R34068 PAD.n604 PAD.n494 2.2505
R34069 PAD.n603 PAD.n602 2.2505
R34070 PAD.n496 PAD.n495 2.2505
R34071 PAD.n594 PAD.n593 2.2505
R34072 PAD.n592 PAD.n498 2.2505
R34073 PAD.n591 PAD.n590 2.2505
R34074 PAD.n500 PAD.n499 2.2505
R34075 PAD.n582 PAD.n581 2.2505
R34076 PAD.n580 PAD.n502 2.2505
R34077 PAD.n579 PAD.n578 2.2505
R34078 PAD.n504 PAD.n503 2.2505
R34079 PAD.n570 PAD.n569 2.2505
R34080 PAD.n568 PAD.n506 2.2505
R34081 PAD.n567 PAD.n566 2.2505
R34082 PAD.n508 PAD.n507 2.2505
R34083 PAD.n558 PAD.n557 2.2505
R34084 PAD.n556 PAD.n510 2.2505
R34085 PAD.n555 PAD.n554 2.2505
R34086 PAD.n512 PAD.n511 2.2505
R34087 PAD.n546 PAD.n545 2.2505
R34088 PAD.n544 PAD.n514 2.2505
R34089 PAD.n543 PAD.n542 2.2505
R34090 PAD.n516 PAD.n515 2.2505
R34091 PAD.n534 PAD.n533 2.2505
R34092 PAD.n532 PAD.n518 2.2505
R34093 PAD.n531 PAD.n530 2.2505
R34094 PAD.n520 PAD.n519 2.2505
R34095 PAD.n522 PAD.n521 2.2505
R34096 PAD.n872 PAD.n824 2.2505
R34097 PAD.n871 PAD.n870 2.2505
R34098 PAD.n877 PAD.n876 2.2505
R34099 PAD.n880 PAD.n879 2.2505
R34100 PAD.n884 PAD.n883 2.2505
R34101 PAD.n881 PAD.n867 2.2505
R34102 PAD.n889 PAD.n888 2.2505
R34103 PAD.n892 PAD.n891 2.2505
R34104 PAD.n896 PAD.n895 2.2505
R34105 PAD.n893 PAD.n865 2.2505
R34106 PAD.n901 PAD.n900 2.2505
R34107 PAD.n904 PAD.n903 2.2505
R34108 PAD.n908 PAD.n907 2.2505
R34109 PAD.n905 PAD.n863 2.2505
R34110 PAD.n913 PAD.n912 2.2505
R34111 PAD.n916 PAD.n915 2.2505
R34112 PAD.n920 PAD.n919 2.2505
R34113 PAD.n917 PAD.n861 2.2505
R34114 PAD.n925 PAD.n924 2.2505
R34115 PAD.n928 PAD.n927 2.2505
R34116 PAD.n932 PAD.n931 2.2505
R34117 PAD.n929 PAD.n859 2.2505
R34118 PAD.n937 PAD.n936 2.2505
R34119 PAD.n940 PAD.n939 2.2505
R34120 PAD.n944 PAD.n943 2.2505
R34121 PAD.n941 PAD.n857 2.2505
R34122 PAD.n949 PAD.n948 2.2505
R34123 PAD.n952 PAD.n951 2.2505
R34124 PAD.n956 PAD.n955 2.2505
R34125 PAD.n953 PAD.n855 2.2505
R34126 PAD.n961 PAD.n960 2.2505
R34127 PAD.n964 PAD.n963 2.2505
R34128 PAD.n968 PAD.n967 2.2505
R34129 PAD.n965 PAD.n853 2.2505
R34130 PAD.n973 PAD.n972 2.2505
R34131 PAD.n976 PAD.n975 2.2505
R34132 PAD.n980 PAD.n979 2.2505
R34133 PAD.n977 PAD.n851 2.2505
R34134 PAD.n985 PAD.n984 2.2505
R34135 PAD.n988 PAD.n987 2.2505
R34136 PAD.n992 PAD.n991 2.2505
R34137 PAD.n989 PAD.n849 2.2505
R34138 PAD.n997 PAD.n996 2.2505
R34139 PAD.n1000 PAD.n999 2.2505
R34140 PAD.n1004 PAD.n1003 2.2505
R34141 PAD.n1001 PAD.n847 2.2505
R34142 PAD.n1009 PAD.n1008 2.2505
R34143 PAD.n1012 PAD.n1011 2.2505
R34144 PAD.n1016 PAD.n1015 2.2505
R34145 PAD.n1013 PAD.n845 2.2505
R34146 PAD.n1021 PAD.n1020 2.2505
R34147 PAD.n1024 PAD.n1023 2.2505
R34148 PAD.n1028 PAD.n1027 2.2505
R34149 PAD.n1025 PAD.n843 2.2505
R34150 PAD.n1033 PAD.n1032 2.2505
R34151 PAD.n1036 PAD.n1035 2.2505
R34152 PAD.n1040 PAD.n1039 2.2505
R34153 PAD.n1037 PAD.n841 2.2505
R34154 PAD.n1045 PAD.n1044 2.2505
R34155 PAD.n1048 PAD.n1047 2.2505
R34156 PAD.n1052 PAD.n1051 2.2505
R34157 PAD.n1049 PAD.n839 2.2505
R34158 PAD.n1057 PAD.n1056 2.2505
R34159 PAD.n1060 PAD.n1059 2.2505
R34160 PAD.n1064 PAD.n1063 2.2505
R34161 PAD.n1061 PAD.n837 2.2505
R34162 PAD.n1069 PAD.n1068 2.2505
R34163 PAD.n1072 PAD.n1071 2.2505
R34164 PAD.n1076 PAD.n1075 2.2505
R34165 PAD.n1073 PAD.n835 2.2505
R34166 PAD.n1081 PAD.n1080 2.2505
R34167 PAD.n1084 PAD.n1083 2.2505
R34168 PAD.n1088 PAD.n1087 2.2505
R34169 PAD.n1085 PAD.n833 2.2505
R34170 PAD.n1093 PAD.n1092 2.2505
R34171 PAD.n1096 PAD.n1095 2.2505
R34172 PAD.n1100 PAD.n1099 2.2505
R34173 PAD.n1097 PAD.n831 2.2505
R34174 PAD.n1105 PAD.n1104 2.2505
R34175 PAD.n1108 PAD.n1107 2.2505
R34176 PAD.n1112 PAD.n1111 2.2505
R34177 PAD.n1109 PAD.n829 2.2505
R34178 PAD.n10385 PAD.n10384 2.2505
R34179 PAD.n10387 PAD.n826 2.2505
R34180 PAD.n10382 PAD.n826 2.2505
R34181 PAD.n10384 PAD.n10383 2.2505
R34182 PAD.n1114 PAD.n829 2.2505
R34183 PAD.n1113 PAD.n1112 2.2505
R34184 PAD.n1108 PAD.n830 2.2505
R34185 PAD.n1104 PAD.n1103 2.2505
R34186 PAD.n1102 PAD.n831 2.2505
R34187 PAD.n1101 PAD.n1100 2.2505
R34188 PAD.n1096 PAD.n832 2.2505
R34189 PAD.n1092 PAD.n1091 2.2505
R34190 PAD.n1090 PAD.n833 2.2505
R34191 PAD.n1089 PAD.n1088 2.2505
R34192 PAD.n1084 PAD.n834 2.2505
R34193 PAD.n1080 PAD.n1079 2.2505
R34194 PAD.n1078 PAD.n835 2.2505
R34195 PAD.n1077 PAD.n1076 2.2505
R34196 PAD.n1072 PAD.n836 2.2505
R34197 PAD.n1068 PAD.n1067 2.2505
R34198 PAD.n1066 PAD.n837 2.2505
R34199 PAD.n1065 PAD.n1064 2.2505
R34200 PAD.n1060 PAD.n838 2.2505
R34201 PAD.n1056 PAD.n1055 2.2505
R34202 PAD.n1054 PAD.n839 2.2505
R34203 PAD.n1053 PAD.n1052 2.2505
R34204 PAD.n1048 PAD.n840 2.2505
R34205 PAD.n1044 PAD.n1043 2.2505
R34206 PAD.n1042 PAD.n841 2.2505
R34207 PAD.n1041 PAD.n1040 2.2505
R34208 PAD.n1036 PAD.n842 2.2505
R34209 PAD.n1032 PAD.n1031 2.2505
R34210 PAD.n1030 PAD.n843 2.2505
R34211 PAD.n1029 PAD.n1028 2.2505
R34212 PAD.n1024 PAD.n844 2.2505
R34213 PAD.n1020 PAD.n1019 2.2505
R34214 PAD.n1018 PAD.n845 2.2505
R34215 PAD.n1017 PAD.n1016 2.2505
R34216 PAD.n1012 PAD.n846 2.2505
R34217 PAD.n1008 PAD.n1007 2.2505
R34218 PAD.n1006 PAD.n847 2.2505
R34219 PAD.n1005 PAD.n1004 2.2505
R34220 PAD.n1000 PAD.n848 2.2505
R34221 PAD.n996 PAD.n995 2.2505
R34222 PAD.n994 PAD.n849 2.2505
R34223 PAD.n993 PAD.n992 2.2505
R34224 PAD.n988 PAD.n850 2.2505
R34225 PAD.n984 PAD.n983 2.2505
R34226 PAD.n982 PAD.n851 2.2505
R34227 PAD.n981 PAD.n980 2.2505
R34228 PAD.n976 PAD.n852 2.2505
R34229 PAD.n972 PAD.n971 2.2505
R34230 PAD.n970 PAD.n853 2.2505
R34231 PAD.n969 PAD.n968 2.2505
R34232 PAD.n964 PAD.n854 2.2505
R34233 PAD.n960 PAD.n959 2.2505
R34234 PAD.n958 PAD.n855 2.2505
R34235 PAD.n957 PAD.n956 2.2505
R34236 PAD.n952 PAD.n856 2.2505
R34237 PAD.n948 PAD.n947 2.2505
R34238 PAD.n946 PAD.n857 2.2505
R34239 PAD.n945 PAD.n944 2.2505
R34240 PAD.n940 PAD.n858 2.2505
R34241 PAD.n936 PAD.n935 2.2505
R34242 PAD.n934 PAD.n859 2.2505
R34243 PAD.n933 PAD.n932 2.2505
R34244 PAD.n928 PAD.n860 2.2505
R34245 PAD.n924 PAD.n923 2.2505
R34246 PAD.n922 PAD.n861 2.2505
R34247 PAD.n921 PAD.n920 2.2505
R34248 PAD.n916 PAD.n862 2.2505
R34249 PAD.n912 PAD.n911 2.2505
R34250 PAD.n910 PAD.n863 2.2505
R34251 PAD.n909 PAD.n908 2.2505
R34252 PAD.n904 PAD.n864 2.2505
R34253 PAD.n900 PAD.n899 2.2505
R34254 PAD.n898 PAD.n865 2.2505
R34255 PAD.n897 PAD.n896 2.2505
R34256 PAD.n892 PAD.n866 2.2505
R34257 PAD.n888 PAD.n887 2.2505
R34258 PAD.n886 PAD.n867 2.2505
R34259 PAD.n885 PAD.n884 2.2505
R34260 PAD.n880 PAD.n868 2.2505
R34261 PAD.n876 PAD.n875 2.2505
R34262 PAD.n874 PAD.n871 2.2505
R34263 PAD.n873 PAD.n872 2.2505
R34264 PAD.n10106 PAD.n10105 2.2505
R34265 PAD.n10108 PAD.n10104 2.2505
R34266 PAD.n10113 PAD.n10112 2.2505
R34267 PAD.n10110 PAD.n10102 2.2505
R34268 PAD.n10118 PAD.n10117 2.2505
R34269 PAD.n10120 PAD.n10100 2.2505
R34270 PAD.n10125 PAD.n10124 2.2505
R34271 PAD.n10122 PAD.n10098 2.2505
R34272 PAD.n10130 PAD.n10129 2.2505
R34273 PAD.n10132 PAD.n10096 2.2505
R34274 PAD.n10137 PAD.n10136 2.2505
R34275 PAD.n10134 PAD.n10094 2.2505
R34276 PAD.n10142 PAD.n10141 2.2505
R34277 PAD.n10144 PAD.n10092 2.2505
R34278 PAD.n10149 PAD.n10148 2.2505
R34279 PAD.n10146 PAD.n10090 2.2505
R34280 PAD.n10154 PAD.n10153 2.2505
R34281 PAD.n10156 PAD.n10088 2.2505
R34282 PAD.n10161 PAD.n10160 2.2505
R34283 PAD.n10158 PAD.n10086 2.2505
R34284 PAD.n10166 PAD.n10165 2.2505
R34285 PAD.n10168 PAD.n10084 2.2505
R34286 PAD.n10173 PAD.n10172 2.2505
R34287 PAD.n10170 PAD.n10082 2.2505
R34288 PAD.n10178 PAD.n10177 2.2505
R34289 PAD.n10180 PAD.n10080 2.2505
R34290 PAD.n10185 PAD.n10184 2.2505
R34291 PAD.n10182 PAD.n10078 2.2505
R34292 PAD.n10190 PAD.n10189 2.2505
R34293 PAD.n10192 PAD.n10076 2.2505
R34294 PAD.n10197 PAD.n10196 2.2505
R34295 PAD.n10194 PAD.n10074 2.2505
R34296 PAD.n10202 PAD.n10201 2.2505
R34297 PAD.n10204 PAD.n10072 2.2505
R34298 PAD.n10209 PAD.n10208 2.2505
R34299 PAD.n10206 PAD.n10070 2.2505
R34300 PAD.n10214 PAD.n10213 2.2505
R34301 PAD.n10216 PAD.n10068 2.2505
R34302 PAD.n10221 PAD.n10220 2.2505
R34303 PAD.n10218 PAD.n10066 2.2505
R34304 PAD.n10226 PAD.n10225 2.2505
R34305 PAD.n10228 PAD.n10064 2.2505
R34306 PAD.n10233 PAD.n10232 2.2505
R34307 PAD.n10230 PAD.n10062 2.2505
R34308 PAD.n10238 PAD.n10237 2.2505
R34309 PAD.n10240 PAD.n10060 2.2505
R34310 PAD.n10245 PAD.n10244 2.2505
R34311 PAD.n10242 PAD.n10058 2.2505
R34312 PAD.n10250 PAD.n10249 2.2505
R34313 PAD.n10252 PAD.n10056 2.2505
R34314 PAD.n10257 PAD.n10256 2.2505
R34315 PAD.n10254 PAD.n10054 2.2505
R34316 PAD.n10262 PAD.n10261 2.2505
R34317 PAD.n10264 PAD.n10052 2.2505
R34318 PAD.n10269 PAD.n10268 2.2505
R34319 PAD.n10266 PAD.n10050 2.2505
R34320 PAD.n10274 PAD.n10273 2.2505
R34321 PAD.n10276 PAD.n10048 2.2505
R34322 PAD.n10281 PAD.n10280 2.2505
R34323 PAD.n10278 PAD.n10046 2.2505
R34324 PAD.n10286 PAD.n10285 2.2505
R34325 PAD.n10288 PAD.n10044 2.2505
R34326 PAD.n10293 PAD.n10292 2.2505
R34327 PAD.n10290 PAD.n10042 2.2505
R34328 PAD.n10298 PAD.n10297 2.2505
R34329 PAD.n10300 PAD.n10040 2.2505
R34330 PAD.n10305 PAD.n10304 2.2505
R34331 PAD.n10302 PAD.n10038 2.2505
R34332 PAD.n10310 PAD.n10309 2.2505
R34333 PAD.n10312 PAD.n10036 2.2505
R34334 PAD.n10317 PAD.n10316 2.2505
R34335 PAD.n10314 PAD.n10034 2.2505
R34336 PAD.n10322 PAD.n10321 2.2505
R34337 PAD.n10324 PAD.n10032 2.2505
R34338 PAD.n10329 PAD.n10328 2.2505
R34339 PAD.n10326 PAD.n10030 2.2505
R34340 PAD.n10334 PAD.n10333 2.2505
R34341 PAD.n10336 PAD.n10028 2.2505
R34342 PAD.n10341 PAD.n10340 2.2505
R34343 PAD.n10338 PAD.n10026 2.2505
R34344 PAD.n10347 PAD.n10346 2.2505
R34345 PAD.n10349 PAD.n10024 2.2505
R34346 PAD.n10351 PAD.n10023 2.2505
R34347 PAD.n10354 PAD.n10353 2.2505
R34348 PAD.n10355 PAD.n10354 2.2505
R34349 PAD.n10023 PAD.n10022 2.2505
R34350 PAD.n10344 PAD.n10024 2.2505
R34351 PAD.n10346 PAD.n10345 2.2505
R34352 PAD.n10343 PAD.n10026 2.2505
R34353 PAD.n10342 PAD.n10341 2.2505
R34354 PAD.n10028 PAD.n10027 2.2505
R34355 PAD.n10333 PAD.n10332 2.2505
R34356 PAD.n10331 PAD.n10030 2.2505
R34357 PAD.n10330 PAD.n10329 2.2505
R34358 PAD.n10032 PAD.n10031 2.2505
R34359 PAD.n10321 PAD.n10320 2.2505
R34360 PAD.n10319 PAD.n10034 2.2505
R34361 PAD.n10318 PAD.n10317 2.2505
R34362 PAD.n10036 PAD.n10035 2.2505
R34363 PAD.n10309 PAD.n10308 2.2505
R34364 PAD.n10307 PAD.n10038 2.2505
R34365 PAD.n10306 PAD.n10305 2.2505
R34366 PAD.n10040 PAD.n10039 2.2505
R34367 PAD.n10297 PAD.n10296 2.2505
R34368 PAD.n10295 PAD.n10042 2.2505
R34369 PAD.n10294 PAD.n10293 2.2505
R34370 PAD.n10044 PAD.n10043 2.2505
R34371 PAD.n10285 PAD.n10284 2.2505
R34372 PAD.n10283 PAD.n10046 2.2505
R34373 PAD.n10282 PAD.n10281 2.2505
R34374 PAD.n10048 PAD.n10047 2.2505
R34375 PAD.n10273 PAD.n10272 2.2505
R34376 PAD.n10271 PAD.n10050 2.2505
R34377 PAD.n10270 PAD.n10269 2.2505
R34378 PAD.n10052 PAD.n10051 2.2505
R34379 PAD.n10261 PAD.n10260 2.2505
R34380 PAD.n10259 PAD.n10054 2.2505
R34381 PAD.n10258 PAD.n10257 2.2505
R34382 PAD.n10056 PAD.n10055 2.2505
R34383 PAD.n10249 PAD.n10248 2.2505
R34384 PAD.n10247 PAD.n10058 2.2505
R34385 PAD.n10246 PAD.n10245 2.2505
R34386 PAD.n10060 PAD.n10059 2.2505
R34387 PAD.n10237 PAD.n10236 2.2505
R34388 PAD.n10235 PAD.n10062 2.2505
R34389 PAD.n10234 PAD.n10233 2.2505
R34390 PAD.n10064 PAD.n10063 2.2505
R34391 PAD.n10225 PAD.n10224 2.2505
R34392 PAD.n10223 PAD.n10066 2.2505
R34393 PAD.n10222 PAD.n10221 2.2505
R34394 PAD.n10068 PAD.n10067 2.2505
R34395 PAD.n10213 PAD.n10212 2.2505
R34396 PAD.n10211 PAD.n10070 2.2505
R34397 PAD.n10210 PAD.n10209 2.2505
R34398 PAD.n10072 PAD.n10071 2.2505
R34399 PAD.n10201 PAD.n10200 2.2505
R34400 PAD.n10199 PAD.n10074 2.2505
R34401 PAD.n10198 PAD.n10197 2.2505
R34402 PAD.n10076 PAD.n10075 2.2505
R34403 PAD.n10189 PAD.n10188 2.2505
R34404 PAD.n10187 PAD.n10078 2.2505
R34405 PAD.n10186 PAD.n10185 2.2505
R34406 PAD.n10080 PAD.n10079 2.2505
R34407 PAD.n10177 PAD.n10176 2.2505
R34408 PAD.n10175 PAD.n10082 2.2505
R34409 PAD.n10174 PAD.n10173 2.2505
R34410 PAD.n10084 PAD.n10083 2.2505
R34411 PAD.n10165 PAD.n10164 2.2505
R34412 PAD.n10163 PAD.n10086 2.2505
R34413 PAD.n10162 PAD.n10161 2.2505
R34414 PAD.n10088 PAD.n10087 2.2505
R34415 PAD.n10153 PAD.n10152 2.2505
R34416 PAD.n10151 PAD.n10090 2.2505
R34417 PAD.n10150 PAD.n10149 2.2505
R34418 PAD.n10092 PAD.n10091 2.2505
R34419 PAD.n10141 PAD.n10140 2.2505
R34420 PAD.n10139 PAD.n10094 2.2505
R34421 PAD.n10138 PAD.n10137 2.2505
R34422 PAD.n10096 PAD.n10095 2.2505
R34423 PAD.n10129 PAD.n10128 2.2505
R34424 PAD.n10127 PAD.n10098 2.2505
R34425 PAD.n10126 PAD.n10125 2.2505
R34426 PAD.n10100 PAD.n10099 2.2505
R34427 PAD.n10117 PAD.n10116 2.2505
R34428 PAD.n10115 PAD.n10102 2.2505
R34429 PAD.n10114 PAD.n10113 2.2505
R34430 PAD.n10104 PAD.n10103 2.2505
R34431 PAD.n10105 PAD.n1124 2.2505
R34432 PAD.n1481 PAD.n1480 2.2505
R34433 PAD.n1479 PAD.n1190 2.2505
R34434 PAD.n1193 PAD.n1192 2.2505
R34435 PAD.n1475 PAD.n1474 2.2505
R34436 PAD.n1472 PAD.n1471 2.2505
R34437 PAD.n1470 PAD.n1198 2.2505
R34438 PAD.n1196 PAD.n1195 2.2505
R34439 PAD.n1466 PAD.n1465 2.2505
R34440 PAD.n1463 PAD.n1462 2.2505
R34441 PAD.n1461 PAD.n1203 2.2505
R34442 PAD.n1201 PAD.n1200 2.2505
R34443 PAD.n1457 PAD.n1456 2.2505
R34444 PAD.n1454 PAD.n1453 2.2505
R34445 PAD.n1452 PAD.n1208 2.2505
R34446 PAD.n1206 PAD.n1205 2.2505
R34447 PAD.n1448 PAD.n1447 2.2505
R34448 PAD.n1445 PAD.n1444 2.2505
R34449 PAD.n1443 PAD.n1213 2.2505
R34450 PAD.n1211 PAD.n1210 2.2505
R34451 PAD.n1439 PAD.n1438 2.2505
R34452 PAD.n1436 PAD.n1435 2.2505
R34453 PAD.n1434 PAD.n1218 2.2505
R34454 PAD.n1216 PAD.n1215 2.2505
R34455 PAD.n1430 PAD.n1429 2.2505
R34456 PAD.n1427 PAD.n1426 2.2505
R34457 PAD.n1425 PAD.n1223 2.2505
R34458 PAD.n1221 PAD.n1220 2.2505
R34459 PAD.n1421 PAD.n1420 2.2505
R34460 PAD.n1418 PAD.n1417 2.2505
R34461 PAD.n1416 PAD.n1228 2.2505
R34462 PAD.n1226 PAD.n1225 2.2505
R34463 PAD.n1412 PAD.n1411 2.2505
R34464 PAD.n1409 PAD.n1408 2.2505
R34465 PAD.n1407 PAD.n1233 2.2505
R34466 PAD.n1231 PAD.n1230 2.2505
R34467 PAD.n1403 PAD.n1402 2.2505
R34468 PAD.n1400 PAD.n1399 2.2505
R34469 PAD.n1398 PAD.n1238 2.2505
R34470 PAD.n1236 PAD.n1235 2.2505
R34471 PAD.n1394 PAD.n1393 2.2505
R34472 PAD.n1391 PAD.n1390 2.2505
R34473 PAD.n1389 PAD.n1243 2.2505
R34474 PAD.n1241 PAD.n1240 2.2505
R34475 PAD.n1385 PAD.n1384 2.2505
R34476 PAD.n1382 PAD.n1381 2.2505
R34477 PAD.n1380 PAD.n1248 2.2505
R34478 PAD.n1246 PAD.n1245 2.2505
R34479 PAD.n1376 PAD.n1375 2.2505
R34480 PAD.n1373 PAD.n1372 2.2505
R34481 PAD.n1371 PAD.n1253 2.2505
R34482 PAD.n1251 PAD.n1250 2.2505
R34483 PAD.n1367 PAD.n1366 2.2505
R34484 PAD.n1364 PAD.n1363 2.2505
R34485 PAD.n1362 PAD.n1258 2.2505
R34486 PAD.n1256 PAD.n1255 2.2505
R34487 PAD.n1358 PAD.n1357 2.2505
R34488 PAD.n1355 PAD.n1354 2.2505
R34489 PAD.n1353 PAD.n1263 2.2505
R34490 PAD.n1261 PAD.n1260 2.2505
R34491 PAD.n1349 PAD.n1348 2.2505
R34492 PAD.n1346 PAD.n1345 2.2505
R34493 PAD.n1344 PAD.n1268 2.2505
R34494 PAD.n1266 PAD.n1265 2.2505
R34495 PAD.n1340 PAD.n1339 2.2505
R34496 PAD.n1337 PAD.n1336 2.2505
R34497 PAD.n1335 PAD.n1273 2.2505
R34498 PAD.n1271 PAD.n1270 2.2505
R34499 PAD.n1331 PAD.n1330 2.2505
R34500 PAD.n1328 PAD.n1327 2.2505
R34501 PAD.n1326 PAD.n1278 2.2505
R34502 PAD.n1276 PAD.n1275 2.2505
R34503 PAD.n1322 PAD.n1321 2.2505
R34504 PAD.n1319 PAD.n1318 2.2505
R34505 PAD.n1317 PAD.n1283 2.2505
R34506 PAD.n1281 PAD.n1280 2.2505
R34507 PAD.n1313 PAD.n1312 2.2505
R34508 PAD.n1310 PAD.n1309 2.2505
R34509 PAD.n1308 PAD.n1288 2.2505
R34510 PAD.n1286 PAD.n1285 2.2505
R34511 PAD.n1304 PAD.n1303 2.2505
R34512 PAD.n1301 PAD.n1300 2.2505
R34513 PAD.n1299 PAD.n1293 2.2505
R34514 PAD.n1291 PAD.n1290 2.2505
R34515 PAD.n1295 PAD.n1294 2.2505
R34516 PAD.n1296 PAD.n1295 2.2505
R34517 PAD.n1297 PAD.n1290 2.2505
R34518 PAD.n1299 PAD.n1298 2.2505
R34519 PAD.n1300 PAD.n1289 2.2505
R34520 PAD.n1305 PAD.n1304 2.2505
R34521 PAD.n1306 PAD.n1285 2.2505
R34522 PAD.n1308 PAD.n1307 2.2505
R34523 PAD.n1309 PAD.n1284 2.2505
R34524 PAD.n1314 PAD.n1313 2.2505
R34525 PAD.n1315 PAD.n1280 2.2505
R34526 PAD.n1317 PAD.n1316 2.2505
R34527 PAD.n1318 PAD.n1279 2.2505
R34528 PAD.n1323 PAD.n1322 2.2505
R34529 PAD.n1324 PAD.n1275 2.2505
R34530 PAD.n1326 PAD.n1325 2.2505
R34531 PAD.n1327 PAD.n1274 2.2505
R34532 PAD.n1332 PAD.n1331 2.2505
R34533 PAD.n1333 PAD.n1270 2.2505
R34534 PAD.n1335 PAD.n1334 2.2505
R34535 PAD.n1336 PAD.n1269 2.2505
R34536 PAD.n1341 PAD.n1340 2.2505
R34537 PAD.n1342 PAD.n1265 2.2505
R34538 PAD.n1344 PAD.n1343 2.2505
R34539 PAD.n1345 PAD.n1264 2.2505
R34540 PAD.n1350 PAD.n1349 2.2505
R34541 PAD.n1351 PAD.n1260 2.2505
R34542 PAD.n1353 PAD.n1352 2.2505
R34543 PAD.n1354 PAD.n1259 2.2505
R34544 PAD.n1359 PAD.n1358 2.2505
R34545 PAD.n1360 PAD.n1255 2.2505
R34546 PAD.n1362 PAD.n1361 2.2505
R34547 PAD.n1363 PAD.n1254 2.2505
R34548 PAD.n1368 PAD.n1367 2.2505
R34549 PAD.n1369 PAD.n1250 2.2505
R34550 PAD.n1371 PAD.n1370 2.2505
R34551 PAD.n1372 PAD.n1249 2.2505
R34552 PAD.n1377 PAD.n1376 2.2505
R34553 PAD.n1378 PAD.n1245 2.2505
R34554 PAD.n1380 PAD.n1379 2.2505
R34555 PAD.n1381 PAD.n1244 2.2505
R34556 PAD.n1386 PAD.n1385 2.2505
R34557 PAD.n1387 PAD.n1240 2.2505
R34558 PAD.n1389 PAD.n1388 2.2505
R34559 PAD.n1390 PAD.n1239 2.2505
R34560 PAD.n1395 PAD.n1394 2.2505
R34561 PAD.n1396 PAD.n1235 2.2505
R34562 PAD.n1398 PAD.n1397 2.2505
R34563 PAD.n1399 PAD.n1234 2.2505
R34564 PAD.n1404 PAD.n1403 2.2505
R34565 PAD.n1405 PAD.n1230 2.2505
R34566 PAD.n1407 PAD.n1406 2.2505
R34567 PAD.n1408 PAD.n1229 2.2505
R34568 PAD.n1413 PAD.n1412 2.2505
R34569 PAD.n1414 PAD.n1225 2.2505
R34570 PAD.n1416 PAD.n1415 2.2505
R34571 PAD.n1417 PAD.n1224 2.2505
R34572 PAD.n1422 PAD.n1421 2.2505
R34573 PAD.n1423 PAD.n1220 2.2505
R34574 PAD.n1425 PAD.n1424 2.2505
R34575 PAD.n1426 PAD.n1219 2.2505
R34576 PAD.n1431 PAD.n1430 2.2505
R34577 PAD.n1432 PAD.n1215 2.2505
R34578 PAD.n1434 PAD.n1433 2.2505
R34579 PAD.n1435 PAD.n1214 2.2505
R34580 PAD.n1440 PAD.n1439 2.2505
R34581 PAD.n1441 PAD.n1210 2.2505
R34582 PAD.n1443 PAD.n1442 2.2505
R34583 PAD.n1444 PAD.n1209 2.2505
R34584 PAD.n1449 PAD.n1448 2.2505
R34585 PAD.n1450 PAD.n1205 2.2505
R34586 PAD.n1452 PAD.n1451 2.2505
R34587 PAD.n1453 PAD.n1204 2.2505
R34588 PAD.n1458 PAD.n1457 2.2505
R34589 PAD.n1459 PAD.n1200 2.2505
R34590 PAD.n1461 PAD.n1460 2.2505
R34591 PAD.n1462 PAD.n1199 2.2505
R34592 PAD.n1467 PAD.n1466 2.2505
R34593 PAD.n1468 PAD.n1195 2.2505
R34594 PAD.n1470 PAD.n1469 2.2505
R34595 PAD.n1471 PAD.n1194 2.2505
R34596 PAD.n1476 PAD.n1475 2.2505
R34597 PAD.n1477 PAD.n1193 2.2505
R34598 PAD.n1479 PAD.n1478 2.2505
R34599 PAD.n1480 PAD.n1145 2.2505
R34600 PAD.n9749 PAD.n1531 2.2505
R34601 PAD.n1579 PAD.n1578 2.2505
R34602 PAD.n9754 PAD.n9753 2.2505
R34603 PAD.n9757 PAD.n9756 2.2505
R34604 PAD.n9761 PAD.n9760 2.2505
R34605 PAD.n9758 PAD.n1575 2.2505
R34606 PAD.n9766 PAD.n9765 2.2505
R34607 PAD.n9769 PAD.n9768 2.2505
R34608 PAD.n9773 PAD.n9772 2.2505
R34609 PAD.n9770 PAD.n1573 2.2505
R34610 PAD.n9778 PAD.n9777 2.2505
R34611 PAD.n9781 PAD.n9780 2.2505
R34612 PAD.n9785 PAD.n9784 2.2505
R34613 PAD.n9782 PAD.n1571 2.2505
R34614 PAD.n9790 PAD.n9789 2.2505
R34615 PAD.n9793 PAD.n9792 2.2505
R34616 PAD.n9797 PAD.n9796 2.2505
R34617 PAD.n9794 PAD.n1569 2.2505
R34618 PAD.n9802 PAD.n9801 2.2505
R34619 PAD.n9805 PAD.n9804 2.2505
R34620 PAD.n9809 PAD.n9808 2.2505
R34621 PAD.n9806 PAD.n1567 2.2505
R34622 PAD.n9814 PAD.n9813 2.2505
R34623 PAD.n9817 PAD.n9816 2.2505
R34624 PAD.n9821 PAD.n9820 2.2505
R34625 PAD.n9818 PAD.n1565 2.2505
R34626 PAD.n9826 PAD.n9825 2.2505
R34627 PAD.n9829 PAD.n9828 2.2505
R34628 PAD.n9833 PAD.n9832 2.2505
R34629 PAD.n9830 PAD.n1563 2.2505
R34630 PAD.n9838 PAD.n9837 2.2505
R34631 PAD.n9841 PAD.n9840 2.2505
R34632 PAD.n9845 PAD.n9844 2.2505
R34633 PAD.n9842 PAD.n1561 2.2505
R34634 PAD.n9850 PAD.n9849 2.2505
R34635 PAD.n9853 PAD.n9852 2.2505
R34636 PAD.n9857 PAD.n9856 2.2505
R34637 PAD.n9854 PAD.n1559 2.2505
R34638 PAD.n9862 PAD.n9861 2.2505
R34639 PAD.n9865 PAD.n9864 2.2505
R34640 PAD.n9869 PAD.n9868 2.2505
R34641 PAD.n9866 PAD.n1557 2.2505
R34642 PAD.n9874 PAD.n9873 2.2505
R34643 PAD.n9877 PAD.n9876 2.2505
R34644 PAD.n9881 PAD.n9880 2.2505
R34645 PAD.n9878 PAD.n1555 2.2505
R34646 PAD.n9886 PAD.n9885 2.2505
R34647 PAD.n9889 PAD.n9888 2.2505
R34648 PAD.n9893 PAD.n9892 2.2505
R34649 PAD.n9890 PAD.n1553 2.2505
R34650 PAD.n9898 PAD.n9897 2.2505
R34651 PAD.n9901 PAD.n9900 2.2505
R34652 PAD.n9905 PAD.n9904 2.2505
R34653 PAD.n9902 PAD.n1551 2.2505
R34654 PAD.n9910 PAD.n9909 2.2505
R34655 PAD.n9913 PAD.n9912 2.2505
R34656 PAD.n9917 PAD.n9916 2.2505
R34657 PAD.n9914 PAD.n1549 2.2505
R34658 PAD.n9922 PAD.n9921 2.2505
R34659 PAD.n9925 PAD.n9924 2.2505
R34660 PAD.n9929 PAD.n9928 2.2505
R34661 PAD.n9926 PAD.n1547 2.2505
R34662 PAD.n9934 PAD.n9933 2.2505
R34663 PAD.n9937 PAD.n9936 2.2505
R34664 PAD.n9941 PAD.n9940 2.2505
R34665 PAD.n9938 PAD.n1545 2.2505
R34666 PAD.n9946 PAD.n9945 2.2505
R34667 PAD.n9949 PAD.n9948 2.2505
R34668 PAD.n9953 PAD.n9952 2.2505
R34669 PAD.n9950 PAD.n1543 2.2505
R34670 PAD.n9958 PAD.n9957 2.2505
R34671 PAD.n9961 PAD.n9960 2.2505
R34672 PAD.n9965 PAD.n9964 2.2505
R34673 PAD.n9962 PAD.n1541 2.2505
R34674 PAD.n9970 PAD.n9969 2.2505
R34675 PAD.n9973 PAD.n9972 2.2505
R34676 PAD.n9977 PAD.n9976 2.2505
R34677 PAD.n9974 PAD.n1539 2.2505
R34678 PAD.n9982 PAD.n9981 2.2505
R34679 PAD.n9985 PAD.n9984 2.2505
R34680 PAD.n9989 PAD.n9988 2.2505
R34681 PAD.n9986 PAD.n1537 2.2505
R34682 PAD.n9995 PAD.n9994 2.2505
R34683 PAD.n9997 PAD.n1535 2.2505
R34684 PAD.n9992 PAD.n1535 2.2505
R34685 PAD.n9994 PAD.n9993 2.2505
R34686 PAD.n9991 PAD.n1537 2.2505
R34687 PAD.n9990 PAD.n9989 2.2505
R34688 PAD.n9985 PAD.n1538 2.2505
R34689 PAD.n9981 PAD.n9980 2.2505
R34690 PAD.n9979 PAD.n1539 2.2505
R34691 PAD.n9978 PAD.n9977 2.2505
R34692 PAD.n9973 PAD.n1540 2.2505
R34693 PAD.n9969 PAD.n9968 2.2505
R34694 PAD.n9967 PAD.n1541 2.2505
R34695 PAD.n9966 PAD.n9965 2.2505
R34696 PAD.n9961 PAD.n1542 2.2505
R34697 PAD.n9957 PAD.n9956 2.2505
R34698 PAD.n9955 PAD.n1543 2.2505
R34699 PAD.n9954 PAD.n9953 2.2505
R34700 PAD.n9949 PAD.n1544 2.2505
R34701 PAD.n9945 PAD.n9944 2.2505
R34702 PAD.n9943 PAD.n1545 2.2505
R34703 PAD.n9942 PAD.n9941 2.2505
R34704 PAD.n9937 PAD.n1546 2.2505
R34705 PAD.n9933 PAD.n9932 2.2505
R34706 PAD.n9931 PAD.n1547 2.2505
R34707 PAD.n9930 PAD.n9929 2.2505
R34708 PAD.n9925 PAD.n1548 2.2505
R34709 PAD.n9921 PAD.n9920 2.2505
R34710 PAD.n9919 PAD.n1549 2.2505
R34711 PAD.n9918 PAD.n9917 2.2505
R34712 PAD.n9913 PAD.n1550 2.2505
R34713 PAD.n9909 PAD.n9908 2.2505
R34714 PAD.n9907 PAD.n1551 2.2505
R34715 PAD.n9906 PAD.n9905 2.2505
R34716 PAD.n9901 PAD.n1552 2.2505
R34717 PAD.n9897 PAD.n9896 2.2505
R34718 PAD.n9895 PAD.n1553 2.2505
R34719 PAD.n9894 PAD.n9893 2.2505
R34720 PAD.n9889 PAD.n1554 2.2505
R34721 PAD.n9885 PAD.n9884 2.2505
R34722 PAD.n9883 PAD.n1555 2.2505
R34723 PAD.n9882 PAD.n9881 2.2505
R34724 PAD.n9877 PAD.n1556 2.2505
R34725 PAD.n9873 PAD.n9872 2.2505
R34726 PAD.n9871 PAD.n1557 2.2505
R34727 PAD.n9870 PAD.n9869 2.2505
R34728 PAD.n9865 PAD.n1558 2.2505
R34729 PAD.n9861 PAD.n9860 2.2505
R34730 PAD.n9859 PAD.n1559 2.2505
R34731 PAD.n9858 PAD.n9857 2.2505
R34732 PAD.n9853 PAD.n1560 2.2505
R34733 PAD.n9849 PAD.n9848 2.2505
R34734 PAD.n9847 PAD.n1561 2.2505
R34735 PAD.n9846 PAD.n9845 2.2505
R34736 PAD.n9841 PAD.n1562 2.2505
R34737 PAD.n9837 PAD.n9836 2.2505
R34738 PAD.n9835 PAD.n1563 2.2505
R34739 PAD.n9834 PAD.n9833 2.2505
R34740 PAD.n9829 PAD.n1564 2.2505
R34741 PAD.n9825 PAD.n9824 2.2505
R34742 PAD.n9823 PAD.n1565 2.2505
R34743 PAD.n9822 PAD.n9821 2.2505
R34744 PAD.n9817 PAD.n1566 2.2505
R34745 PAD.n9813 PAD.n9812 2.2505
R34746 PAD.n9811 PAD.n1567 2.2505
R34747 PAD.n9810 PAD.n9809 2.2505
R34748 PAD.n9805 PAD.n1568 2.2505
R34749 PAD.n9801 PAD.n9800 2.2505
R34750 PAD.n9799 PAD.n1569 2.2505
R34751 PAD.n9798 PAD.n9797 2.2505
R34752 PAD.n9793 PAD.n1570 2.2505
R34753 PAD.n9789 PAD.n9788 2.2505
R34754 PAD.n9787 PAD.n1571 2.2505
R34755 PAD.n9786 PAD.n9785 2.2505
R34756 PAD.n9781 PAD.n1572 2.2505
R34757 PAD.n9777 PAD.n9776 2.2505
R34758 PAD.n9775 PAD.n1573 2.2505
R34759 PAD.n9774 PAD.n9773 2.2505
R34760 PAD.n9769 PAD.n1574 2.2505
R34761 PAD.n9765 PAD.n9764 2.2505
R34762 PAD.n9763 PAD.n1575 2.2505
R34763 PAD.n9762 PAD.n9761 2.2505
R34764 PAD.n9757 PAD.n1576 2.2505
R34765 PAD.n9753 PAD.n9752 2.2505
R34766 PAD.n9751 PAD.n1579 2.2505
R34767 PAD.n9750 PAD.n9749 2.2505
R34768 PAD.n1931 PAD.n1599 2.2505
R34769 PAD.n1930 PAD.n1929 2.2505
R34770 PAD.n1927 PAD.n1600 2.2505
R34771 PAD.n1925 PAD.n1924 2.2505
R34772 PAD.n1917 PAD.n1603 2.2505
R34773 PAD.n1920 PAD.n1919 2.2505
R34774 PAD.n1915 PAD.n1606 2.2505
R34775 PAD.n1913 PAD.n1912 2.2505
R34776 PAD.n1905 PAD.n1608 2.2505
R34777 PAD.n1908 PAD.n1907 2.2505
R34778 PAD.n1903 PAD.n1610 2.2505
R34779 PAD.n1901 PAD.n1900 2.2505
R34780 PAD.n1893 PAD.n1612 2.2505
R34781 PAD.n1896 PAD.n1895 2.2505
R34782 PAD.n1891 PAD.n1614 2.2505
R34783 PAD.n1889 PAD.n1888 2.2505
R34784 PAD.n1881 PAD.n1616 2.2505
R34785 PAD.n1884 PAD.n1883 2.2505
R34786 PAD.n1879 PAD.n1618 2.2505
R34787 PAD.n1877 PAD.n1876 2.2505
R34788 PAD.n1869 PAD.n1620 2.2505
R34789 PAD.n1872 PAD.n1871 2.2505
R34790 PAD.n1867 PAD.n1622 2.2505
R34791 PAD.n1865 PAD.n1864 2.2505
R34792 PAD.n1857 PAD.n1624 2.2505
R34793 PAD.n1860 PAD.n1859 2.2505
R34794 PAD.n1855 PAD.n1626 2.2505
R34795 PAD.n1853 PAD.n1852 2.2505
R34796 PAD.n1845 PAD.n1628 2.2505
R34797 PAD.n1848 PAD.n1847 2.2505
R34798 PAD.n1843 PAD.n1630 2.2505
R34799 PAD.n1841 PAD.n1840 2.2505
R34800 PAD.n1833 PAD.n1632 2.2505
R34801 PAD.n1836 PAD.n1835 2.2505
R34802 PAD.n1831 PAD.n1634 2.2505
R34803 PAD.n1829 PAD.n1828 2.2505
R34804 PAD.n1821 PAD.n1636 2.2505
R34805 PAD.n1824 PAD.n1823 2.2505
R34806 PAD.n1819 PAD.n1638 2.2505
R34807 PAD.n1817 PAD.n1816 2.2505
R34808 PAD.n1809 PAD.n1640 2.2505
R34809 PAD.n1812 PAD.n1811 2.2505
R34810 PAD.n1807 PAD.n1642 2.2505
R34811 PAD.n1805 PAD.n1804 2.2505
R34812 PAD.n1797 PAD.n1644 2.2505
R34813 PAD.n1800 PAD.n1799 2.2505
R34814 PAD.n1795 PAD.n1646 2.2505
R34815 PAD.n1793 PAD.n1792 2.2505
R34816 PAD.n1785 PAD.n1648 2.2505
R34817 PAD.n1788 PAD.n1787 2.2505
R34818 PAD.n1783 PAD.n1650 2.2505
R34819 PAD.n1781 PAD.n1780 2.2505
R34820 PAD.n1773 PAD.n1652 2.2505
R34821 PAD.n1776 PAD.n1775 2.2505
R34822 PAD.n1771 PAD.n1654 2.2505
R34823 PAD.n1769 PAD.n1768 2.2505
R34824 PAD.n1761 PAD.n1656 2.2505
R34825 PAD.n1764 PAD.n1763 2.2505
R34826 PAD.n1759 PAD.n1658 2.2505
R34827 PAD.n1757 PAD.n1756 2.2505
R34828 PAD.n1749 PAD.n1660 2.2505
R34829 PAD.n1752 PAD.n1751 2.2505
R34830 PAD.n1747 PAD.n1662 2.2505
R34831 PAD.n1745 PAD.n1744 2.2505
R34832 PAD.n1737 PAD.n1664 2.2505
R34833 PAD.n1740 PAD.n1739 2.2505
R34834 PAD.n1735 PAD.n1666 2.2505
R34835 PAD.n1733 PAD.n1732 2.2505
R34836 PAD.n1725 PAD.n1668 2.2505
R34837 PAD.n1728 PAD.n1727 2.2505
R34838 PAD.n1723 PAD.n1670 2.2505
R34839 PAD.n1721 PAD.n1720 2.2505
R34840 PAD.n1713 PAD.n1672 2.2505
R34841 PAD.n1716 PAD.n1715 2.2505
R34842 PAD.n1711 PAD.n1674 2.2505
R34843 PAD.n1709 PAD.n1708 2.2505
R34844 PAD.n1701 PAD.n1676 2.2505
R34845 PAD.n1704 PAD.n1703 2.2505
R34846 PAD.n1699 PAD.n1678 2.2505
R34847 PAD.n1697 PAD.n1696 2.2505
R34848 PAD.n1689 PAD.n1680 2.2505
R34849 PAD.n1692 PAD.n1691 2.2505
R34850 PAD.n1687 PAD.n1682 2.2505
R34851 PAD.n1685 PAD.n1684 2.2505
R34852 PAD.n1684 PAD.n1683 2.2505
R34853 PAD.n1682 PAD.n1681 2.2505
R34854 PAD.n1693 PAD.n1692 2.2505
R34855 PAD.n1694 PAD.n1680 2.2505
R34856 PAD.n1696 PAD.n1695 2.2505
R34857 PAD.n1678 PAD.n1677 2.2505
R34858 PAD.n1705 PAD.n1704 2.2505
R34859 PAD.n1706 PAD.n1676 2.2505
R34860 PAD.n1708 PAD.n1707 2.2505
R34861 PAD.n1674 PAD.n1673 2.2505
R34862 PAD.n1717 PAD.n1716 2.2505
R34863 PAD.n1718 PAD.n1672 2.2505
R34864 PAD.n1720 PAD.n1719 2.2505
R34865 PAD.n1670 PAD.n1669 2.2505
R34866 PAD.n1729 PAD.n1728 2.2505
R34867 PAD.n1730 PAD.n1668 2.2505
R34868 PAD.n1732 PAD.n1731 2.2505
R34869 PAD.n1666 PAD.n1665 2.2505
R34870 PAD.n1741 PAD.n1740 2.2505
R34871 PAD.n1742 PAD.n1664 2.2505
R34872 PAD.n1744 PAD.n1743 2.2505
R34873 PAD.n1662 PAD.n1661 2.2505
R34874 PAD.n1753 PAD.n1752 2.2505
R34875 PAD.n1754 PAD.n1660 2.2505
R34876 PAD.n1756 PAD.n1755 2.2505
R34877 PAD.n1658 PAD.n1657 2.2505
R34878 PAD.n1765 PAD.n1764 2.2505
R34879 PAD.n1766 PAD.n1656 2.2505
R34880 PAD.n1768 PAD.n1767 2.2505
R34881 PAD.n1654 PAD.n1653 2.2505
R34882 PAD.n1777 PAD.n1776 2.2505
R34883 PAD.n1778 PAD.n1652 2.2505
R34884 PAD.n1780 PAD.n1779 2.2505
R34885 PAD.n1650 PAD.n1649 2.2505
R34886 PAD.n1789 PAD.n1788 2.2505
R34887 PAD.n1790 PAD.n1648 2.2505
R34888 PAD.n1792 PAD.n1791 2.2505
R34889 PAD.n1646 PAD.n1645 2.2505
R34890 PAD.n1801 PAD.n1800 2.2505
R34891 PAD.n1802 PAD.n1644 2.2505
R34892 PAD.n1804 PAD.n1803 2.2505
R34893 PAD.n1642 PAD.n1641 2.2505
R34894 PAD.n1813 PAD.n1812 2.2505
R34895 PAD.n1814 PAD.n1640 2.2505
R34896 PAD.n1816 PAD.n1815 2.2505
R34897 PAD.n1638 PAD.n1637 2.2505
R34898 PAD.n1825 PAD.n1824 2.2505
R34899 PAD.n1826 PAD.n1636 2.2505
R34900 PAD.n1828 PAD.n1827 2.2505
R34901 PAD.n1634 PAD.n1633 2.2505
R34902 PAD.n1837 PAD.n1836 2.2505
R34903 PAD.n1838 PAD.n1632 2.2505
R34904 PAD.n1840 PAD.n1839 2.2505
R34905 PAD.n1630 PAD.n1629 2.2505
R34906 PAD.n1849 PAD.n1848 2.2505
R34907 PAD.n1850 PAD.n1628 2.2505
R34908 PAD.n1852 PAD.n1851 2.2505
R34909 PAD.n1626 PAD.n1625 2.2505
R34910 PAD.n1861 PAD.n1860 2.2505
R34911 PAD.n1862 PAD.n1624 2.2505
R34912 PAD.n1864 PAD.n1863 2.2505
R34913 PAD.n1622 PAD.n1621 2.2505
R34914 PAD.n1873 PAD.n1872 2.2505
R34915 PAD.n1874 PAD.n1620 2.2505
R34916 PAD.n1876 PAD.n1875 2.2505
R34917 PAD.n1618 PAD.n1617 2.2505
R34918 PAD.n1885 PAD.n1884 2.2505
R34919 PAD.n1886 PAD.n1616 2.2505
R34920 PAD.n1888 PAD.n1887 2.2505
R34921 PAD.n1614 PAD.n1613 2.2505
R34922 PAD.n1897 PAD.n1896 2.2505
R34923 PAD.n1898 PAD.n1612 2.2505
R34924 PAD.n1900 PAD.n1899 2.2505
R34925 PAD.n1610 PAD.n1609 2.2505
R34926 PAD.n1909 PAD.n1908 2.2505
R34927 PAD.n1910 PAD.n1608 2.2505
R34928 PAD.n1912 PAD.n1911 2.2505
R34929 PAD.n1606 PAD.n1605 2.2505
R34930 PAD.n1921 PAD.n1920 2.2505
R34931 PAD.n1922 PAD.n1603 2.2505
R34932 PAD.n1924 PAD.n1923 2.2505
R34933 PAD.n1604 PAD.n1600 2.2505
R34934 PAD.n1930 PAD.n1598 2.2505
R34935 PAD.n1932 PAD.n1931 2.2505
R34936 PAD.n9463 PAD.n1984 2.2505
R34937 PAD.n2031 PAD.n2030 2.2505
R34938 PAD.n9468 PAD.n9467 2.2505
R34939 PAD.n9471 PAD.n9470 2.2505
R34940 PAD.n9475 PAD.n9474 2.2505
R34941 PAD.n9472 PAD.n2027 2.2505
R34942 PAD.n9480 PAD.n9479 2.2505
R34943 PAD.n9483 PAD.n9482 2.2505
R34944 PAD.n9487 PAD.n9486 2.2505
R34945 PAD.n9484 PAD.n2025 2.2505
R34946 PAD.n9492 PAD.n9491 2.2505
R34947 PAD.n9495 PAD.n9494 2.2505
R34948 PAD.n9499 PAD.n9498 2.2505
R34949 PAD.n9496 PAD.n2023 2.2505
R34950 PAD.n9504 PAD.n9503 2.2505
R34951 PAD.n9507 PAD.n9506 2.2505
R34952 PAD.n9511 PAD.n9510 2.2505
R34953 PAD.n9508 PAD.n2021 2.2505
R34954 PAD.n9516 PAD.n9515 2.2505
R34955 PAD.n9519 PAD.n9518 2.2505
R34956 PAD.n9523 PAD.n9522 2.2505
R34957 PAD.n9520 PAD.n2019 2.2505
R34958 PAD.n9528 PAD.n9527 2.2505
R34959 PAD.n9531 PAD.n9530 2.2505
R34960 PAD.n9535 PAD.n9534 2.2505
R34961 PAD.n9532 PAD.n2017 2.2505
R34962 PAD.n9540 PAD.n9539 2.2505
R34963 PAD.n9543 PAD.n9542 2.2505
R34964 PAD.n9547 PAD.n9546 2.2505
R34965 PAD.n9544 PAD.n2015 2.2505
R34966 PAD.n9552 PAD.n9551 2.2505
R34967 PAD.n9555 PAD.n9554 2.2505
R34968 PAD.n9559 PAD.n9558 2.2505
R34969 PAD.n9556 PAD.n2013 2.2505
R34970 PAD.n9564 PAD.n9563 2.2505
R34971 PAD.n9567 PAD.n9566 2.2505
R34972 PAD.n9571 PAD.n9570 2.2505
R34973 PAD.n9568 PAD.n2011 2.2505
R34974 PAD.n9576 PAD.n9575 2.2505
R34975 PAD.n9579 PAD.n9578 2.2505
R34976 PAD.n9583 PAD.n9582 2.2505
R34977 PAD.n9580 PAD.n2009 2.2505
R34978 PAD.n9588 PAD.n9587 2.2505
R34979 PAD.n9591 PAD.n9590 2.2505
R34980 PAD.n9595 PAD.n9594 2.2505
R34981 PAD.n9592 PAD.n2007 2.2505
R34982 PAD.n9600 PAD.n9599 2.2505
R34983 PAD.n9603 PAD.n9602 2.2505
R34984 PAD.n9607 PAD.n9606 2.2505
R34985 PAD.n9604 PAD.n2005 2.2505
R34986 PAD.n9612 PAD.n9611 2.2505
R34987 PAD.n9615 PAD.n9614 2.2505
R34988 PAD.n9619 PAD.n9618 2.2505
R34989 PAD.n9616 PAD.n2003 2.2505
R34990 PAD.n9624 PAD.n9623 2.2505
R34991 PAD.n9627 PAD.n9626 2.2505
R34992 PAD.n9631 PAD.n9630 2.2505
R34993 PAD.n9628 PAD.n2001 2.2505
R34994 PAD.n9636 PAD.n9635 2.2505
R34995 PAD.n9639 PAD.n9638 2.2505
R34996 PAD.n9643 PAD.n9642 2.2505
R34997 PAD.n9640 PAD.n1999 2.2505
R34998 PAD.n9648 PAD.n9647 2.2505
R34999 PAD.n9651 PAD.n9650 2.2505
R35000 PAD.n9655 PAD.n9654 2.2505
R35001 PAD.n9652 PAD.n1997 2.2505
R35002 PAD.n9660 PAD.n9659 2.2505
R35003 PAD.n9663 PAD.n9662 2.2505
R35004 PAD.n9667 PAD.n9666 2.2505
R35005 PAD.n9664 PAD.n1995 2.2505
R35006 PAD.n9672 PAD.n9671 2.2505
R35007 PAD.n9675 PAD.n9674 2.2505
R35008 PAD.n9679 PAD.n9678 2.2505
R35009 PAD.n9676 PAD.n1993 2.2505
R35010 PAD.n9684 PAD.n9683 2.2505
R35011 PAD.n9687 PAD.n9686 2.2505
R35012 PAD.n9691 PAD.n9690 2.2505
R35013 PAD.n9688 PAD.n1991 2.2505
R35014 PAD.n9696 PAD.n9695 2.2505
R35015 PAD.n9699 PAD.n9698 2.2505
R35016 PAD.n9703 PAD.n9702 2.2505
R35017 PAD.n9700 PAD.n1989 2.2505
R35018 PAD.n9709 PAD.n9708 2.2505
R35019 PAD.n9711 PAD.n1987 2.2505
R35020 PAD.n9706 PAD.n1987 2.2505
R35021 PAD.n9708 PAD.n9707 2.2505
R35022 PAD.n9705 PAD.n1989 2.2505
R35023 PAD.n9704 PAD.n9703 2.2505
R35024 PAD.n9699 PAD.n1990 2.2505
R35025 PAD.n9695 PAD.n9694 2.2505
R35026 PAD.n9693 PAD.n1991 2.2505
R35027 PAD.n9692 PAD.n9691 2.2505
R35028 PAD.n9687 PAD.n1992 2.2505
R35029 PAD.n9683 PAD.n9682 2.2505
R35030 PAD.n9681 PAD.n1993 2.2505
R35031 PAD.n9680 PAD.n9679 2.2505
R35032 PAD.n9675 PAD.n1994 2.2505
R35033 PAD.n9671 PAD.n9670 2.2505
R35034 PAD.n9669 PAD.n1995 2.2505
R35035 PAD.n9668 PAD.n9667 2.2505
R35036 PAD.n9663 PAD.n1996 2.2505
R35037 PAD.n9659 PAD.n9658 2.2505
R35038 PAD.n9657 PAD.n1997 2.2505
R35039 PAD.n9656 PAD.n9655 2.2505
R35040 PAD.n9651 PAD.n1998 2.2505
R35041 PAD.n9647 PAD.n9646 2.2505
R35042 PAD.n9645 PAD.n1999 2.2505
R35043 PAD.n9644 PAD.n9643 2.2505
R35044 PAD.n9639 PAD.n2000 2.2505
R35045 PAD.n9635 PAD.n9634 2.2505
R35046 PAD.n9633 PAD.n2001 2.2505
R35047 PAD.n9632 PAD.n9631 2.2505
R35048 PAD.n9627 PAD.n2002 2.2505
R35049 PAD.n9623 PAD.n9622 2.2505
R35050 PAD.n9621 PAD.n2003 2.2505
R35051 PAD.n9620 PAD.n9619 2.2505
R35052 PAD.n9615 PAD.n2004 2.2505
R35053 PAD.n9611 PAD.n9610 2.2505
R35054 PAD.n9609 PAD.n2005 2.2505
R35055 PAD.n9608 PAD.n9607 2.2505
R35056 PAD.n9603 PAD.n2006 2.2505
R35057 PAD.n9599 PAD.n9598 2.2505
R35058 PAD.n9597 PAD.n2007 2.2505
R35059 PAD.n9596 PAD.n9595 2.2505
R35060 PAD.n9591 PAD.n2008 2.2505
R35061 PAD.n9587 PAD.n9586 2.2505
R35062 PAD.n9585 PAD.n2009 2.2505
R35063 PAD.n9584 PAD.n9583 2.2505
R35064 PAD.n9579 PAD.n2010 2.2505
R35065 PAD.n9575 PAD.n9574 2.2505
R35066 PAD.n9573 PAD.n2011 2.2505
R35067 PAD.n9572 PAD.n9571 2.2505
R35068 PAD.n9567 PAD.n2012 2.2505
R35069 PAD.n9563 PAD.n9562 2.2505
R35070 PAD.n9561 PAD.n2013 2.2505
R35071 PAD.n9560 PAD.n9559 2.2505
R35072 PAD.n9555 PAD.n2014 2.2505
R35073 PAD.n9551 PAD.n9550 2.2505
R35074 PAD.n9549 PAD.n2015 2.2505
R35075 PAD.n9548 PAD.n9547 2.2505
R35076 PAD.n9543 PAD.n2016 2.2505
R35077 PAD.n9539 PAD.n9538 2.2505
R35078 PAD.n9537 PAD.n2017 2.2505
R35079 PAD.n9536 PAD.n9535 2.2505
R35080 PAD.n9531 PAD.n2018 2.2505
R35081 PAD.n9527 PAD.n9526 2.2505
R35082 PAD.n9525 PAD.n2019 2.2505
R35083 PAD.n9524 PAD.n9523 2.2505
R35084 PAD.n9519 PAD.n2020 2.2505
R35085 PAD.n9515 PAD.n9514 2.2505
R35086 PAD.n9513 PAD.n2021 2.2505
R35087 PAD.n9512 PAD.n9511 2.2505
R35088 PAD.n9507 PAD.n2022 2.2505
R35089 PAD.n9503 PAD.n9502 2.2505
R35090 PAD.n9501 PAD.n2023 2.2505
R35091 PAD.n9500 PAD.n9499 2.2505
R35092 PAD.n9495 PAD.n2024 2.2505
R35093 PAD.n9491 PAD.n9490 2.2505
R35094 PAD.n9489 PAD.n2025 2.2505
R35095 PAD.n9488 PAD.n9487 2.2505
R35096 PAD.n9483 PAD.n2026 2.2505
R35097 PAD.n9479 PAD.n9478 2.2505
R35098 PAD.n9477 PAD.n2027 2.2505
R35099 PAD.n9476 PAD.n9475 2.2505
R35100 PAD.n9471 PAD.n2028 2.2505
R35101 PAD.n9467 PAD.n9466 2.2505
R35102 PAD.n9465 PAD.n2031 2.2505
R35103 PAD.n9464 PAD.n9463 2.2505
R35104 PAD.n9197 PAD.n2088 2.2505
R35105 PAD.n2134 PAD.n2133 2.2505
R35106 PAD.n9202 PAD.n9201 2.2505
R35107 PAD.n9205 PAD.n9204 2.2505
R35108 PAD.n9209 PAD.n9208 2.2505
R35109 PAD.n9206 PAD.n2130 2.2505
R35110 PAD.n9214 PAD.n9213 2.2505
R35111 PAD.n9217 PAD.n9216 2.2505
R35112 PAD.n9221 PAD.n9220 2.2505
R35113 PAD.n9218 PAD.n2128 2.2505
R35114 PAD.n9226 PAD.n9225 2.2505
R35115 PAD.n9229 PAD.n9228 2.2505
R35116 PAD.n9233 PAD.n9232 2.2505
R35117 PAD.n9230 PAD.n2126 2.2505
R35118 PAD.n9238 PAD.n9237 2.2505
R35119 PAD.n9241 PAD.n9240 2.2505
R35120 PAD.n9245 PAD.n9244 2.2505
R35121 PAD.n9242 PAD.n2124 2.2505
R35122 PAD.n9250 PAD.n9249 2.2505
R35123 PAD.n9253 PAD.n9252 2.2505
R35124 PAD.n9257 PAD.n9256 2.2505
R35125 PAD.n9254 PAD.n2122 2.2505
R35126 PAD.n9262 PAD.n9261 2.2505
R35127 PAD.n9265 PAD.n9264 2.2505
R35128 PAD.n9269 PAD.n9268 2.2505
R35129 PAD.n9266 PAD.n2120 2.2505
R35130 PAD.n9274 PAD.n9273 2.2505
R35131 PAD.n9277 PAD.n9276 2.2505
R35132 PAD.n9281 PAD.n9280 2.2505
R35133 PAD.n9278 PAD.n2118 2.2505
R35134 PAD.n9286 PAD.n9285 2.2505
R35135 PAD.n9289 PAD.n9288 2.2505
R35136 PAD.n9293 PAD.n9292 2.2505
R35137 PAD.n9290 PAD.n2116 2.2505
R35138 PAD.n9298 PAD.n9297 2.2505
R35139 PAD.n9301 PAD.n9300 2.2505
R35140 PAD.n9305 PAD.n9304 2.2505
R35141 PAD.n9302 PAD.n2114 2.2505
R35142 PAD.n9310 PAD.n9309 2.2505
R35143 PAD.n9313 PAD.n9312 2.2505
R35144 PAD.n9317 PAD.n9316 2.2505
R35145 PAD.n9314 PAD.n2112 2.2505
R35146 PAD.n9322 PAD.n9321 2.2505
R35147 PAD.n9325 PAD.n9324 2.2505
R35148 PAD.n9329 PAD.n9328 2.2505
R35149 PAD.n9326 PAD.n2110 2.2505
R35150 PAD.n9334 PAD.n9333 2.2505
R35151 PAD.n9337 PAD.n9336 2.2505
R35152 PAD.n9341 PAD.n9340 2.2505
R35153 PAD.n9338 PAD.n2108 2.2505
R35154 PAD.n9346 PAD.n9345 2.2505
R35155 PAD.n9349 PAD.n9348 2.2505
R35156 PAD.n9353 PAD.n9352 2.2505
R35157 PAD.n9350 PAD.n2106 2.2505
R35158 PAD.n9358 PAD.n9357 2.2505
R35159 PAD.n9361 PAD.n9360 2.2505
R35160 PAD.n9365 PAD.n9364 2.2505
R35161 PAD.n9362 PAD.n2104 2.2505
R35162 PAD.n9370 PAD.n9369 2.2505
R35163 PAD.n9373 PAD.n9372 2.2505
R35164 PAD.n9377 PAD.n9376 2.2505
R35165 PAD.n9374 PAD.n2102 2.2505
R35166 PAD.n9382 PAD.n9381 2.2505
R35167 PAD.n9385 PAD.n9384 2.2505
R35168 PAD.n9389 PAD.n9388 2.2505
R35169 PAD.n9386 PAD.n2100 2.2505
R35170 PAD.n9394 PAD.n9393 2.2505
R35171 PAD.n9397 PAD.n9396 2.2505
R35172 PAD.n9401 PAD.n9400 2.2505
R35173 PAD.n9398 PAD.n2098 2.2505
R35174 PAD.n9406 PAD.n9405 2.2505
R35175 PAD.n9409 PAD.n9408 2.2505
R35176 PAD.n9413 PAD.n9412 2.2505
R35177 PAD.n9410 PAD.n2096 2.2505
R35178 PAD.n9418 PAD.n9417 2.2505
R35179 PAD.n9421 PAD.n9420 2.2505
R35180 PAD.n9425 PAD.n9424 2.2505
R35181 PAD.n9422 PAD.n2094 2.2505
R35182 PAD.n9430 PAD.n9429 2.2505
R35183 PAD.n9433 PAD.n9432 2.2505
R35184 PAD.n9437 PAD.n9436 2.2505
R35185 PAD.n9434 PAD.n2092 2.2505
R35186 PAD.n9442 PAD.n9441 2.2505
R35187 PAD.n9444 PAD.n2090 2.2505
R35188 PAD.n2090 PAD.n2040 2.2505
R35189 PAD.n9441 PAD.n9440 2.2505
R35190 PAD.n9439 PAD.n2092 2.2505
R35191 PAD.n9438 PAD.n9437 2.2505
R35192 PAD.n9433 PAD.n2093 2.2505
R35193 PAD.n9429 PAD.n9428 2.2505
R35194 PAD.n9427 PAD.n2094 2.2505
R35195 PAD.n9426 PAD.n9425 2.2505
R35196 PAD.n9421 PAD.n2095 2.2505
R35197 PAD.n9417 PAD.n9416 2.2505
R35198 PAD.n9415 PAD.n2096 2.2505
R35199 PAD.n9414 PAD.n9413 2.2505
R35200 PAD.n9409 PAD.n2097 2.2505
R35201 PAD.n9405 PAD.n9404 2.2505
R35202 PAD.n9403 PAD.n2098 2.2505
R35203 PAD.n9402 PAD.n9401 2.2505
R35204 PAD.n9397 PAD.n2099 2.2505
R35205 PAD.n9393 PAD.n9392 2.2505
R35206 PAD.n9391 PAD.n2100 2.2505
R35207 PAD.n9390 PAD.n9389 2.2505
R35208 PAD.n9385 PAD.n2101 2.2505
R35209 PAD.n9381 PAD.n9380 2.2505
R35210 PAD.n9379 PAD.n2102 2.2505
R35211 PAD.n9378 PAD.n9377 2.2505
R35212 PAD.n9373 PAD.n2103 2.2505
R35213 PAD.n9369 PAD.n9368 2.2505
R35214 PAD.n9367 PAD.n2104 2.2505
R35215 PAD.n9366 PAD.n9365 2.2505
R35216 PAD.n9361 PAD.n2105 2.2505
R35217 PAD.n9357 PAD.n9356 2.2505
R35218 PAD.n9355 PAD.n2106 2.2505
R35219 PAD.n9354 PAD.n9353 2.2505
R35220 PAD.n9349 PAD.n2107 2.2505
R35221 PAD.n9345 PAD.n9344 2.2505
R35222 PAD.n9343 PAD.n2108 2.2505
R35223 PAD.n9342 PAD.n9341 2.2505
R35224 PAD.n9337 PAD.n2109 2.2505
R35225 PAD.n9333 PAD.n9332 2.2505
R35226 PAD.n9331 PAD.n2110 2.2505
R35227 PAD.n9330 PAD.n9329 2.2505
R35228 PAD.n9325 PAD.n2111 2.2505
R35229 PAD.n9321 PAD.n9320 2.2505
R35230 PAD.n9319 PAD.n2112 2.2505
R35231 PAD.n9318 PAD.n9317 2.2505
R35232 PAD.n9313 PAD.n2113 2.2505
R35233 PAD.n9309 PAD.n9308 2.2505
R35234 PAD.n9307 PAD.n2114 2.2505
R35235 PAD.n9306 PAD.n9305 2.2505
R35236 PAD.n9301 PAD.n2115 2.2505
R35237 PAD.n9297 PAD.n9296 2.2505
R35238 PAD.n9295 PAD.n2116 2.2505
R35239 PAD.n9294 PAD.n9293 2.2505
R35240 PAD.n9289 PAD.n2117 2.2505
R35241 PAD.n9285 PAD.n9284 2.2505
R35242 PAD.n9283 PAD.n2118 2.2505
R35243 PAD.n9282 PAD.n9281 2.2505
R35244 PAD.n9277 PAD.n2119 2.2505
R35245 PAD.n9273 PAD.n9272 2.2505
R35246 PAD.n9271 PAD.n2120 2.2505
R35247 PAD.n9270 PAD.n9269 2.2505
R35248 PAD.n9265 PAD.n2121 2.2505
R35249 PAD.n9261 PAD.n9260 2.2505
R35250 PAD.n9259 PAD.n2122 2.2505
R35251 PAD.n9258 PAD.n9257 2.2505
R35252 PAD.n9253 PAD.n2123 2.2505
R35253 PAD.n9249 PAD.n9248 2.2505
R35254 PAD.n9247 PAD.n2124 2.2505
R35255 PAD.n9246 PAD.n9245 2.2505
R35256 PAD.n9241 PAD.n2125 2.2505
R35257 PAD.n9237 PAD.n9236 2.2505
R35258 PAD.n9235 PAD.n2126 2.2505
R35259 PAD.n9234 PAD.n9233 2.2505
R35260 PAD.n9229 PAD.n2127 2.2505
R35261 PAD.n9225 PAD.n9224 2.2505
R35262 PAD.n9223 PAD.n2128 2.2505
R35263 PAD.n9222 PAD.n9221 2.2505
R35264 PAD.n9217 PAD.n2129 2.2505
R35265 PAD.n9213 PAD.n9212 2.2505
R35266 PAD.n9211 PAD.n2130 2.2505
R35267 PAD.n9210 PAD.n9209 2.2505
R35268 PAD.n9205 PAD.n2131 2.2505
R35269 PAD.n9201 PAD.n9200 2.2505
R35270 PAD.n9199 PAD.n2134 2.2505
R35271 PAD.n9198 PAD.n9197 2.2505
R35272 PAD.n2482 PAD.n2151 2.2505
R35273 PAD.n2481 PAD.n2480 2.2505
R35274 PAD.n2478 PAD.n2152 2.2505
R35275 PAD.n2476 PAD.n2475 2.2505
R35276 PAD.n2468 PAD.n2155 2.2505
R35277 PAD.n2471 PAD.n2470 2.2505
R35278 PAD.n2466 PAD.n2158 2.2505
R35279 PAD.n2464 PAD.n2463 2.2505
R35280 PAD.n2456 PAD.n2160 2.2505
R35281 PAD.n2459 PAD.n2458 2.2505
R35282 PAD.n2454 PAD.n2162 2.2505
R35283 PAD.n2452 PAD.n2451 2.2505
R35284 PAD.n2444 PAD.n2164 2.2505
R35285 PAD.n2447 PAD.n2446 2.2505
R35286 PAD.n2442 PAD.n2166 2.2505
R35287 PAD.n2440 PAD.n2439 2.2505
R35288 PAD.n2432 PAD.n2168 2.2505
R35289 PAD.n2435 PAD.n2434 2.2505
R35290 PAD.n2430 PAD.n2170 2.2505
R35291 PAD.n2428 PAD.n2427 2.2505
R35292 PAD.n2420 PAD.n2172 2.2505
R35293 PAD.n2423 PAD.n2422 2.2505
R35294 PAD.n2418 PAD.n2174 2.2505
R35295 PAD.n2416 PAD.n2415 2.2505
R35296 PAD.n2408 PAD.n2176 2.2505
R35297 PAD.n2411 PAD.n2410 2.2505
R35298 PAD.n2406 PAD.n2178 2.2505
R35299 PAD.n2404 PAD.n2403 2.2505
R35300 PAD.n2396 PAD.n2180 2.2505
R35301 PAD.n2399 PAD.n2398 2.2505
R35302 PAD.n2394 PAD.n2182 2.2505
R35303 PAD.n2392 PAD.n2391 2.2505
R35304 PAD.n2384 PAD.n2184 2.2505
R35305 PAD.n2387 PAD.n2386 2.2505
R35306 PAD.n2382 PAD.n2186 2.2505
R35307 PAD.n2380 PAD.n2379 2.2505
R35308 PAD.n2372 PAD.n2188 2.2505
R35309 PAD.n2375 PAD.n2374 2.2505
R35310 PAD.n2370 PAD.n2190 2.2505
R35311 PAD.n2368 PAD.n2367 2.2505
R35312 PAD.n2360 PAD.n2192 2.2505
R35313 PAD.n2363 PAD.n2362 2.2505
R35314 PAD.n2358 PAD.n2194 2.2505
R35315 PAD.n2356 PAD.n2355 2.2505
R35316 PAD.n2348 PAD.n2196 2.2505
R35317 PAD.n2351 PAD.n2350 2.2505
R35318 PAD.n2346 PAD.n2198 2.2505
R35319 PAD.n2344 PAD.n2343 2.2505
R35320 PAD.n2336 PAD.n2200 2.2505
R35321 PAD.n2339 PAD.n2338 2.2505
R35322 PAD.n2334 PAD.n2202 2.2505
R35323 PAD.n2332 PAD.n2331 2.2505
R35324 PAD.n2324 PAD.n2204 2.2505
R35325 PAD.n2327 PAD.n2326 2.2505
R35326 PAD.n2322 PAD.n2206 2.2505
R35327 PAD.n2320 PAD.n2319 2.2505
R35328 PAD.n2312 PAD.n2208 2.2505
R35329 PAD.n2315 PAD.n2314 2.2505
R35330 PAD.n2310 PAD.n2210 2.2505
R35331 PAD.n2308 PAD.n2307 2.2505
R35332 PAD.n2300 PAD.n2212 2.2505
R35333 PAD.n2303 PAD.n2302 2.2505
R35334 PAD.n2298 PAD.n2214 2.2505
R35335 PAD.n2296 PAD.n2295 2.2505
R35336 PAD.n2288 PAD.n2216 2.2505
R35337 PAD.n2291 PAD.n2290 2.2505
R35338 PAD.n2286 PAD.n2218 2.2505
R35339 PAD.n2284 PAD.n2283 2.2505
R35340 PAD.n2276 PAD.n2220 2.2505
R35341 PAD.n2279 PAD.n2278 2.2505
R35342 PAD.n2274 PAD.n2222 2.2505
R35343 PAD.n2272 PAD.n2271 2.2505
R35344 PAD.n2264 PAD.n2224 2.2505
R35345 PAD.n2267 PAD.n2266 2.2505
R35346 PAD.n2262 PAD.n2226 2.2505
R35347 PAD.n2260 PAD.n2259 2.2505
R35348 PAD.n2252 PAD.n2228 2.2505
R35349 PAD.n2255 PAD.n2254 2.2505
R35350 PAD.n2250 PAD.n2230 2.2505
R35351 PAD.n2248 PAD.n2247 2.2505
R35352 PAD.n2240 PAD.n2232 2.2505
R35353 PAD.n2243 PAD.n2242 2.2505
R35354 PAD.n2238 PAD.n2234 2.2505
R35355 PAD.n2236 PAD.n2235 2.2505
R35356 PAD.n2235 PAD.n2142 2.2505
R35357 PAD.n2234 PAD.n2233 2.2505
R35358 PAD.n2244 PAD.n2243 2.2505
R35359 PAD.n2245 PAD.n2232 2.2505
R35360 PAD.n2247 PAD.n2246 2.2505
R35361 PAD.n2230 PAD.n2229 2.2505
R35362 PAD.n2256 PAD.n2255 2.2505
R35363 PAD.n2257 PAD.n2228 2.2505
R35364 PAD.n2259 PAD.n2258 2.2505
R35365 PAD.n2226 PAD.n2225 2.2505
R35366 PAD.n2268 PAD.n2267 2.2505
R35367 PAD.n2269 PAD.n2224 2.2505
R35368 PAD.n2271 PAD.n2270 2.2505
R35369 PAD.n2222 PAD.n2221 2.2505
R35370 PAD.n2280 PAD.n2279 2.2505
R35371 PAD.n2281 PAD.n2220 2.2505
R35372 PAD.n2283 PAD.n2282 2.2505
R35373 PAD.n2218 PAD.n2217 2.2505
R35374 PAD.n2292 PAD.n2291 2.2505
R35375 PAD.n2293 PAD.n2216 2.2505
R35376 PAD.n2295 PAD.n2294 2.2505
R35377 PAD.n2214 PAD.n2213 2.2505
R35378 PAD.n2304 PAD.n2303 2.2505
R35379 PAD.n2305 PAD.n2212 2.2505
R35380 PAD.n2307 PAD.n2306 2.2505
R35381 PAD.n2210 PAD.n2209 2.2505
R35382 PAD.n2316 PAD.n2315 2.2505
R35383 PAD.n2317 PAD.n2208 2.2505
R35384 PAD.n2319 PAD.n2318 2.2505
R35385 PAD.n2206 PAD.n2205 2.2505
R35386 PAD.n2328 PAD.n2327 2.2505
R35387 PAD.n2329 PAD.n2204 2.2505
R35388 PAD.n2331 PAD.n2330 2.2505
R35389 PAD.n2202 PAD.n2201 2.2505
R35390 PAD.n2340 PAD.n2339 2.2505
R35391 PAD.n2341 PAD.n2200 2.2505
R35392 PAD.n2343 PAD.n2342 2.2505
R35393 PAD.n2198 PAD.n2197 2.2505
R35394 PAD.n2352 PAD.n2351 2.2505
R35395 PAD.n2353 PAD.n2196 2.2505
R35396 PAD.n2355 PAD.n2354 2.2505
R35397 PAD.n2194 PAD.n2193 2.2505
R35398 PAD.n2364 PAD.n2363 2.2505
R35399 PAD.n2365 PAD.n2192 2.2505
R35400 PAD.n2367 PAD.n2366 2.2505
R35401 PAD.n2190 PAD.n2189 2.2505
R35402 PAD.n2376 PAD.n2375 2.2505
R35403 PAD.n2377 PAD.n2188 2.2505
R35404 PAD.n2379 PAD.n2378 2.2505
R35405 PAD.n2186 PAD.n2185 2.2505
R35406 PAD.n2388 PAD.n2387 2.2505
R35407 PAD.n2389 PAD.n2184 2.2505
R35408 PAD.n2391 PAD.n2390 2.2505
R35409 PAD.n2182 PAD.n2181 2.2505
R35410 PAD.n2400 PAD.n2399 2.2505
R35411 PAD.n2401 PAD.n2180 2.2505
R35412 PAD.n2403 PAD.n2402 2.2505
R35413 PAD.n2178 PAD.n2177 2.2505
R35414 PAD.n2412 PAD.n2411 2.2505
R35415 PAD.n2413 PAD.n2176 2.2505
R35416 PAD.n2415 PAD.n2414 2.2505
R35417 PAD.n2174 PAD.n2173 2.2505
R35418 PAD.n2424 PAD.n2423 2.2505
R35419 PAD.n2425 PAD.n2172 2.2505
R35420 PAD.n2427 PAD.n2426 2.2505
R35421 PAD.n2170 PAD.n2169 2.2505
R35422 PAD.n2436 PAD.n2435 2.2505
R35423 PAD.n2437 PAD.n2168 2.2505
R35424 PAD.n2439 PAD.n2438 2.2505
R35425 PAD.n2166 PAD.n2165 2.2505
R35426 PAD.n2448 PAD.n2447 2.2505
R35427 PAD.n2449 PAD.n2164 2.2505
R35428 PAD.n2451 PAD.n2450 2.2505
R35429 PAD.n2162 PAD.n2161 2.2505
R35430 PAD.n2460 PAD.n2459 2.2505
R35431 PAD.n2461 PAD.n2160 2.2505
R35432 PAD.n2463 PAD.n2462 2.2505
R35433 PAD.n2158 PAD.n2157 2.2505
R35434 PAD.n2472 PAD.n2471 2.2505
R35435 PAD.n2473 PAD.n2155 2.2505
R35436 PAD.n2475 PAD.n2474 2.2505
R35437 PAD.n2156 PAD.n2152 2.2505
R35438 PAD.n2481 PAD.n2150 2.2505
R35439 PAD.n2483 PAD.n2482 2.2505
R35440 PAD.n2829 PAD.n2498 2.2505
R35441 PAD.n2828 PAD.n2827 2.2505
R35442 PAD.n2825 PAD.n2499 2.2505
R35443 PAD.n2823 PAD.n2822 2.2505
R35444 PAD.n2815 PAD.n2502 2.2505
R35445 PAD.n2818 PAD.n2817 2.2505
R35446 PAD.n2813 PAD.n2505 2.2505
R35447 PAD.n2811 PAD.n2810 2.2505
R35448 PAD.n2803 PAD.n2507 2.2505
R35449 PAD.n2806 PAD.n2805 2.2505
R35450 PAD.n2801 PAD.n2509 2.2505
R35451 PAD.n2799 PAD.n2798 2.2505
R35452 PAD.n2791 PAD.n2511 2.2505
R35453 PAD.n2794 PAD.n2793 2.2505
R35454 PAD.n2789 PAD.n2513 2.2505
R35455 PAD.n2787 PAD.n2786 2.2505
R35456 PAD.n2779 PAD.n2515 2.2505
R35457 PAD.n2782 PAD.n2781 2.2505
R35458 PAD.n2777 PAD.n2517 2.2505
R35459 PAD.n2775 PAD.n2774 2.2505
R35460 PAD.n2767 PAD.n2519 2.2505
R35461 PAD.n2770 PAD.n2769 2.2505
R35462 PAD.n2765 PAD.n2521 2.2505
R35463 PAD.n2763 PAD.n2762 2.2505
R35464 PAD.n2755 PAD.n2523 2.2505
R35465 PAD.n2758 PAD.n2757 2.2505
R35466 PAD.n2753 PAD.n2525 2.2505
R35467 PAD.n2751 PAD.n2750 2.2505
R35468 PAD.n2743 PAD.n2527 2.2505
R35469 PAD.n2746 PAD.n2745 2.2505
R35470 PAD.n2741 PAD.n2529 2.2505
R35471 PAD.n2739 PAD.n2738 2.2505
R35472 PAD.n2731 PAD.n2531 2.2505
R35473 PAD.n2734 PAD.n2733 2.2505
R35474 PAD.n2729 PAD.n2533 2.2505
R35475 PAD.n2727 PAD.n2726 2.2505
R35476 PAD.n2719 PAD.n2535 2.2505
R35477 PAD.n2722 PAD.n2721 2.2505
R35478 PAD.n2717 PAD.n2537 2.2505
R35479 PAD.n2715 PAD.n2714 2.2505
R35480 PAD.n2707 PAD.n2539 2.2505
R35481 PAD.n2710 PAD.n2709 2.2505
R35482 PAD.n2705 PAD.n2541 2.2505
R35483 PAD.n2703 PAD.n2702 2.2505
R35484 PAD.n2695 PAD.n2543 2.2505
R35485 PAD.n2698 PAD.n2697 2.2505
R35486 PAD.n2693 PAD.n2545 2.2505
R35487 PAD.n2691 PAD.n2690 2.2505
R35488 PAD.n2683 PAD.n2547 2.2505
R35489 PAD.n2686 PAD.n2685 2.2505
R35490 PAD.n2681 PAD.n2549 2.2505
R35491 PAD.n2679 PAD.n2678 2.2505
R35492 PAD.n2671 PAD.n2551 2.2505
R35493 PAD.n2674 PAD.n2673 2.2505
R35494 PAD.n2669 PAD.n2553 2.2505
R35495 PAD.n2667 PAD.n2666 2.2505
R35496 PAD.n2659 PAD.n2555 2.2505
R35497 PAD.n2662 PAD.n2661 2.2505
R35498 PAD.n2657 PAD.n2557 2.2505
R35499 PAD.n2655 PAD.n2654 2.2505
R35500 PAD.n2647 PAD.n2559 2.2505
R35501 PAD.n2650 PAD.n2649 2.2505
R35502 PAD.n2645 PAD.n2561 2.2505
R35503 PAD.n2643 PAD.n2642 2.2505
R35504 PAD.n2635 PAD.n2563 2.2505
R35505 PAD.n2638 PAD.n2637 2.2505
R35506 PAD.n2633 PAD.n2565 2.2505
R35507 PAD.n2631 PAD.n2630 2.2505
R35508 PAD.n2623 PAD.n2567 2.2505
R35509 PAD.n2626 PAD.n2625 2.2505
R35510 PAD.n2621 PAD.n2569 2.2505
R35511 PAD.n2619 PAD.n2618 2.2505
R35512 PAD.n2611 PAD.n2571 2.2505
R35513 PAD.n2614 PAD.n2613 2.2505
R35514 PAD.n2609 PAD.n2573 2.2505
R35515 PAD.n2607 PAD.n2606 2.2505
R35516 PAD.n2599 PAD.n2575 2.2505
R35517 PAD.n2602 PAD.n2601 2.2505
R35518 PAD.n2597 PAD.n2577 2.2505
R35519 PAD.n2595 PAD.n2594 2.2505
R35520 PAD.n2587 PAD.n2579 2.2505
R35521 PAD.n2590 PAD.n2589 2.2505
R35522 PAD.n2585 PAD.n2581 2.2505
R35523 PAD.n2583 PAD.n2582 2.2505
R35524 PAD.n2582 PAD.n2490 2.2505
R35525 PAD.n2581 PAD.n2580 2.2505
R35526 PAD.n2591 PAD.n2590 2.2505
R35527 PAD.n2592 PAD.n2579 2.2505
R35528 PAD.n2594 PAD.n2593 2.2505
R35529 PAD.n2577 PAD.n2576 2.2505
R35530 PAD.n2603 PAD.n2602 2.2505
R35531 PAD.n2604 PAD.n2575 2.2505
R35532 PAD.n2606 PAD.n2605 2.2505
R35533 PAD.n2573 PAD.n2572 2.2505
R35534 PAD.n2615 PAD.n2614 2.2505
R35535 PAD.n2616 PAD.n2571 2.2505
R35536 PAD.n2618 PAD.n2617 2.2505
R35537 PAD.n2569 PAD.n2568 2.2505
R35538 PAD.n2627 PAD.n2626 2.2505
R35539 PAD.n2628 PAD.n2567 2.2505
R35540 PAD.n2630 PAD.n2629 2.2505
R35541 PAD.n2565 PAD.n2564 2.2505
R35542 PAD.n2639 PAD.n2638 2.2505
R35543 PAD.n2640 PAD.n2563 2.2505
R35544 PAD.n2642 PAD.n2641 2.2505
R35545 PAD.n2561 PAD.n2560 2.2505
R35546 PAD.n2651 PAD.n2650 2.2505
R35547 PAD.n2652 PAD.n2559 2.2505
R35548 PAD.n2654 PAD.n2653 2.2505
R35549 PAD.n2557 PAD.n2556 2.2505
R35550 PAD.n2663 PAD.n2662 2.2505
R35551 PAD.n2664 PAD.n2555 2.2505
R35552 PAD.n2666 PAD.n2665 2.2505
R35553 PAD.n2553 PAD.n2552 2.2505
R35554 PAD.n2675 PAD.n2674 2.2505
R35555 PAD.n2676 PAD.n2551 2.2505
R35556 PAD.n2678 PAD.n2677 2.2505
R35557 PAD.n2549 PAD.n2548 2.2505
R35558 PAD.n2687 PAD.n2686 2.2505
R35559 PAD.n2688 PAD.n2547 2.2505
R35560 PAD.n2690 PAD.n2689 2.2505
R35561 PAD.n2545 PAD.n2544 2.2505
R35562 PAD.n2699 PAD.n2698 2.2505
R35563 PAD.n2700 PAD.n2543 2.2505
R35564 PAD.n2702 PAD.n2701 2.2505
R35565 PAD.n2541 PAD.n2540 2.2505
R35566 PAD.n2711 PAD.n2710 2.2505
R35567 PAD.n2712 PAD.n2539 2.2505
R35568 PAD.n2714 PAD.n2713 2.2505
R35569 PAD.n2537 PAD.n2536 2.2505
R35570 PAD.n2723 PAD.n2722 2.2505
R35571 PAD.n2724 PAD.n2535 2.2505
R35572 PAD.n2726 PAD.n2725 2.2505
R35573 PAD.n2533 PAD.n2532 2.2505
R35574 PAD.n2735 PAD.n2734 2.2505
R35575 PAD.n2736 PAD.n2531 2.2505
R35576 PAD.n2738 PAD.n2737 2.2505
R35577 PAD.n2529 PAD.n2528 2.2505
R35578 PAD.n2747 PAD.n2746 2.2505
R35579 PAD.n2748 PAD.n2527 2.2505
R35580 PAD.n2750 PAD.n2749 2.2505
R35581 PAD.n2525 PAD.n2524 2.2505
R35582 PAD.n2759 PAD.n2758 2.2505
R35583 PAD.n2760 PAD.n2523 2.2505
R35584 PAD.n2762 PAD.n2761 2.2505
R35585 PAD.n2521 PAD.n2520 2.2505
R35586 PAD.n2771 PAD.n2770 2.2505
R35587 PAD.n2772 PAD.n2519 2.2505
R35588 PAD.n2774 PAD.n2773 2.2505
R35589 PAD.n2517 PAD.n2516 2.2505
R35590 PAD.n2783 PAD.n2782 2.2505
R35591 PAD.n2784 PAD.n2515 2.2505
R35592 PAD.n2786 PAD.n2785 2.2505
R35593 PAD.n2513 PAD.n2512 2.2505
R35594 PAD.n2795 PAD.n2794 2.2505
R35595 PAD.n2796 PAD.n2511 2.2505
R35596 PAD.n2798 PAD.n2797 2.2505
R35597 PAD.n2509 PAD.n2508 2.2505
R35598 PAD.n2807 PAD.n2806 2.2505
R35599 PAD.n2808 PAD.n2507 2.2505
R35600 PAD.n2810 PAD.n2809 2.2505
R35601 PAD.n2505 PAD.n2504 2.2505
R35602 PAD.n2819 PAD.n2818 2.2505
R35603 PAD.n2820 PAD.n2502 2.2505
R35604 PAD.n2822 PAD.n2821 2.2505
R35605 PAD.n2503 PAD.n2499 2.2505
R35606 PAD.n2828 PAD.n2497 2.2505
R35607 PAD.n2830 PAD.n2829 2.2505
R35608 PAD.n9119 PAD.n2876 2.2505
R35609 PAD.n9118 PAD.n9117 2.2505
R35610 PAD.n9115 PAD.n8841 2.2505
R35611 PAD.n8839 PAD.n8838 2.2505
R35612 PAD.n9111 PAD.n9110 2.2505
R35613 PAD.n9108 PAD.n9107 2.2505
R35614 PAD.n9106 PAD.n8846 2.2505
R35615 PAD.n8844 PAD.n8843 2.2505
R35616 PAD.n9102 PAD.n9101 2.2505
R35617 PAD.n9099 PAD.n9098 2.2505
R35618 PAD.n9097 PAD.n8851 2.2505
R35619 PAD.n8849 PAD.n8848 2.2505
R35620 PAD.n9093 PAD.n9092 2.2505
R35621 PAD.n9090 PAD.n9089 2.2505
R35622 PAD.n9088 PAD.n8856 2.2505
R35623 PAD.n8854 PAD.n8853 2.2505
R35624 PAD.n9084 PAD.n9083 2.2505
R35625 PAD.n9081 PAD.n9080 2.2505
R35626 PAD.n9079 PAD.n8861 2.2505
R35627 PAD.n8859 PAD.n8858 2.2505
R35628 PAD.n9075 PAD.n9074 2.2505
R35629 PAD.n9072 PAD.n9071 2.2505
R35630 PAD.n9070 PAD.n8866 2.2505
R35631 PAD.n8864 PAD.n8863 2.2505
R35632 PAD.n9066 PAD.n9065 2.2505
R35633 PAD.n9063 PAD.n9062 2.2505
R35634 PAD.n9061 PAD.n8871 2.2505
R35635 PAD.n8869 PAD.n8868 2.2505
R35636 PAD.n9057 PAD.n9056 2.2505
R35637 PAD.n9054 PAD.n9053 2.2505
R35638 PAD.n9052 PAD.n8876 2.2505
R35639 PAD.n8874 PAD.n8873 2.2505
R35640 PAD.n9048 PAD.n9047 2.2505
R35641 PAD.n9045 PAD.n9044 2.2505
R35642 PAD.n9043 PAD.n8881 2.2505
R35643 PAD.n8879 PAD.n8878 2.2505
R35644 PAD.n9039 PAD.n9038 2.2505
R35645 PAD.n9036 PAD.n9035 2.2505
R35646 PAD.n9034 PAD.n8886 2.2505
R35647 PAD.n8884 PAD.n8883 2.2505
R35648 PAD.n9030 PAD.n9029 2.2505
R35649 PAD.n9027 PAD.n9026 2.2505
R35650 PAD.n9025 PAD.n8891 2.2505
R35651 PAD.n8889 PAD.n8888 2.2505
R35652 PAD.n9021 PAD.n9020 2.2505
R35653 PAD.n9018 PAD.n9017 2.2505
R35654 PAD.n9016 PAD.n8896 2.2505
R35655 PAD.n8894 PAD.n8893 2.2505
R35656 PAD.n9012 PAD.n9011 2.2505
R35657 PAD.n9009 PAD.n9008 2.2505
R35658 PAD.n9007 PAD.n8901 2.2505
R35659 PAD.n8899 PAD.n8898 2.2505
R35660 PAD.n9003 PAD.n9002 2.2505
R35661 PAD.n9000 PAD.n8999 2.2505
R35662 PAD.n8998 PAD.n8906 2.2505
R35663 PAD.n8904 PAD.n8903 2.2505
R35664 PAD.n8994 PAD.n8993 2.2505
R35665 PAD.n8991 PAD.n8990 2.2505
R35666 PAD.n8989 PAD.n8911 2.2505
R35667 PAD.n8909 PAD.n8908 2.2505
R35668 PAD.n8985 PAD.n8984 2.2505
R35669 PAD.n8982 PAD.n8981 2.2505
R35670 PAD.n8980 PAD.n8916 2.2505
R35671 PAD.n8914 PAD.n8913 2.2505
R35672 PAD.n8976 PAD.n8975 2.2505
R35673 PAD.n8973 PAD.n8972 2.2505
R35674 PAD.n8971 PAD.n8921 2.2505
R35675 PAD.n8919 PAD.n8918 2.2505
R35676 PAD.n8967 PAD.n8966 2.2505
R35677 PAD.n8964 PAD.n8963 2.2505
R35678 PAD.n8962 PAD.n8926 2.2505
R35679 PAD.n8924 PAD.n8923 2.2505
R35680 PAD.n8958 PAD.n8957 2.2505
R35681 PAD.n8955 PAD.n8954 2.2505
R35682 PAD.n8953 PAD.n8931 2.2505
R35683 PAD.n8929 PAD.n8928 2.2505
R35684 PAD.n8949 PAD.n8948 2.2505
R35685 PAD.n8946 PAD.n8945 2.2505
R35686 PAD.n8944 PAD.n8936 2.2505
R35687 PAD.n8934 PAD.n8933 2.2505
R35688 PAD.n8940 PAD.n8939 2.2505
R35689 PAD.n8937 PAD.n2880 2.2505
R35690 PAD.n9137 PAD.n9136 2.2505
R35691 PAD.n9139 PAD.n2877 2.2505
R35692 PAD.n9134 PAD.n2877 2.2505
R35693 PAD.n9136 PAD.n9135 2.2505
R35694 PAD.n2881 PAD.n2880 2.2505
R35695 PAD.n8941 PAD.n8940 2.2505
R35696 PAD.n8942 PAD.n8933 2.2505
R35697 PAD.n8944 PAD.n8943 2.2505
R35698 PAD.n8945 PAD.n8932 2.2505
R35699 PAD.n8950 PAD.n8949 2.2505
R35700 PAD.n8951 PAD.n8928 2.2505
R35701 PAD.n8953 PAD.n8952 2.2505
R35702 PAD.n8954 PAD.n8927 2.2505
R35703 PAD.n8959 PAD.n8958 2.2505
R35704 PAD.n8960 PAD.n8923 2.2505
R35705 PAD.n8962 PAD.n8961 2.2505
R35706 PAD.n8963 PAD.n8922 2.2505
R35707 PAD.n8968 PAD.n8967 2.2505
R35708 PAD.n8969 PAD.n8918 2.2505
R35709 PAD.n8971 PAD.n8970 2.2505
R35710 PAD.n8972 PAD.n8917 2.2505
R35711 PAD.n8977 PAD.n8976 2.2505
R35712 PAD.n8978 PAD.n8913 2.2505
R35713 PAD.n8980 PAD.n8979 2.2505
R35714 PAD.n8981 PAD.n8912 2.2505
R35715 PAD.n8986 PAD.n8985 2.2505
R35716 PAD.n8987 PAD.n8908 2.2505
R35717 PAD.n8989 PAD.n8988 2.2505
R35718 PAD.n8990 PAD.n8907 2.2505
R35719 PAD.n8995 PAD.n8994 2.2505
R35720 PAD.n8996 PAD.n8903 2.2505
R35721 PAD.n8998 PAD.n8997 2.2505
R35722 PAD.n8999 PAD.n8902 2.2505
R35723 PAD.n9004 PAD.n9003 2.2505
R35724 PAD.n9005 PAD.n8898 2.2505
R35725 PAD.n9007 PAD.n9006 2.2505
R35726 PAD.n9008 PAD.n8897 2.2505
R35727 PAD.n9013 PAD.n9012 2.2505
R35728 PAD.n9014 PAD.n8893 2.2505
R35729 PAD.n9016 PAD.n9015 2.2505
R35730 PAD.n9017 PAD.n8892 2.2505
R35731 PAD.n9022 PAD.n9021 2.2505
R35732 PAD.n9023 PAD.n8888 2.2505
R35733 PAD.n9025 PAD.n9024 2.2505
R35734 PAD.n9026 PAD.n8887 2.2505
R35735 PAD.n9031 PAD.n9030 2.2505
R35736 PAD.n9032 PAD.n8883 2.2505
R35737 PAD.n9034 PAD.n9033 2.2505
R35738 PAD.n9035 PAD.n8882 2.2505
R35739 PAD.n9040 PAD.n9039 2.2505
R35740 PAD.n9041 PAD.n8878 2.2505
R35741 PAD.n9043 PAD.n9042 2.2505
R35742 PAD.n9044 PAD.n8877 2.2505
R35743 PAD.n9049 PAD.n9048 2.2505
R35744 PAD.n9050 PAD.n8873 2.2505
R35745 PAD.n9052 PAD.n9051 2.2505
R35746 PAD.n9053 PAD.n8872 2.2505
R35747 PAD.n9058 PAD.n9057 2.2505
R35748 PAD.n9059 PAD.n8868 2.2505
R35749 PAD.n9061 PAD.n9060 2.2505
R35750 PAD.n9062 PAD.n8867 2.2505
R35751 PAD.n9067 PAD.n9066 2.2505
R35752 PAD.n9068 PAD.n8863 2.2505
R35753 PAD.n9070 PAD.n9069 2.2505
R35754 PAD.n9071 PAD.n8862 2.2505
R35755 PAD.n9076 PAD.n9075 2.2505
R35756 PAD.n9077 PAD.n8858 2.2505
R35757 PAD.n9079 PAD.n9078 2.2505
R35758 PAD.n9080 PAD.n8857 2.2505
R35759 PAD.n9085 PAD.n9084 2.2505
R35760 PAD.n9086 PAD.n8853 2.2505
R35761 PAD.n9088 PAD.n9087 2.2505
R35762 PAD.n9089 PAD.n8852 2.2505
R35763 PAD.n9094 PAD.n9093 2.2505
R35764 PAD.n9095 PAD.n8848 2.2505
R35765 PAD.n9097 PAD.n9096 2.2505
R35766 PAD.n9098 PAD.n8847 2.2505
R35767 PAD.n9103 PAD.n9102 2.2505
R35768 PAD.n9104 PAD.n8843 2.2505
R35769 PAD.n9106 PAD.n9105 2.2505
R35770 PAD.n9107 PAD.n8842 2.2505
R35771 PAD.n9112 PAD.n9111 2.2505
R35772 PAD.n9113 PAD.n8838 2.2505
R35773 PAD.n9115 PAD.n9114 2.2505
R35774 PAD.n9118 PAD.n8837 2.2505
R35775 PAD.n9120 PAD.n9119 2.2505
R35776 PAD.n8819 PAD.n8818 2.2505
R35777 PAD.n8529 PAD.n8528 2.2505
R35778 PAD.n8814 PAD.n8813 2.2505
R35779 PAD.n8811 PAD.n8810 2.2505
R35780 PAD.n8808 PAD.n8807 2.2505
R35781 PAD.n8800 PAD.n8531 2.2505
R35782 PAD.n8803 PAD.n8802 2.2505
R35783 PAD.n8799 PAD.n8798 2.2505
R35784 PAD.n8796 PAD.n8795 2.2505
R35785 PAD.n8788 PAD.n8533 2.2505
R35786 PAD.n8791 PAD.n8790 2.2505
R35787 PAD.n8787 PAD.n8786 2.2505
R35788 PAD.n8784 PAD.n8783 2.2505
R35789 PAD.n8776 PAD.n8535 2.2505
R35790 PAD.n8779 PAD.n8778 2.2505
R35791 PAD.n8775 PAD.n8774 2.2505
R35792 PAD.n8772 PAD.n8771 2.2505
R35793 PAD.n8764 PAD.n8537 2.2505
R35794 PAD.n8767 PAD.n8766 2.2505
R35795 PAD.n8763 PAD.n8762 2.2505
R35796 PAD.n8760 PAD.n8759 2.2505
R35797 PAD.n8752 PAD.n8539 2.2505
R35798 PAD.n8755 PAD.n8754 2.2505
R35799 PAD.n8751 PAD.n8750 2.2505
R35800 PAD.n8748 PAD.n8747 2.2505
R35801 PAD.n8740 PAD.n8541 2.2505
R35802 PAD.n8743 PAD.n8742 2.2505
R35803 PAD.n8739 PAD.n8738 2.2505
R35804 PAD.n8736 PAD.n8735 2.2505
R35805 PAD.n8728 PAD.n8543 2.2505
R35806 PAD.n8731 PAD.n8730 2.2505
R35807 PAD.n8727 PAD.n8726 2.2505
R35808 PAD.n8724 PAD.n8723 2.2505
R35809 PAD.n8716 PAD.n8545 2.2505
R35810 PAD.n8719 PAD.n8718 2.2505
R35811 PAD.n8715 PAD.n8714 2.2505
R35812 PAD.n8712 PAD.n8711 2.2505
R35813 PAD.n8704 PAD.n8547 2.2505
R35814 PAD.n8707 PAD.n8706 2.2505
R35815 PAD.n8703 PAD.n8702 2.2505
R35816 PAD.n8700 PAD.n8699 2.2505
R35817 PAD.n8692 PAD.n8549 2.2505
R35818 PAD.n8695 PAD.n8694 2.2505
R35819 PAD.n8691 PAD.n8690 2.2505
R35820 PAD.n8688 PAD.n8687 2.2505
R35821 PAD.n8680 PAD.n8551 2.2505
R35822 PAD.n8683 PAD.n8682 2.2505
R35823 PAD.n8679 PAD.n8678 2.2505
R35824 PAD.n8676 PAD.n8675 2.2505
R35825 PAD.n8668 PAD.n8553 2.2505
R35826 PAD.n8671 PAD.n8670 2.2505
R35827 PAD.n8667 PAD.n8666 2.2505
R35828 PAD.n8664 PAD.n8663 2.2505
R35829 PAD.n8656 PAD.n8555 2.2505
R35830 PAD.n8659 PAD.n8658 2.2505
R35831 PAD.n8655 PAD.n8654 2.2505
R35832 PAD.n8652 PAD.n8651 2.2505
R35833 PAD.n8644 PAD.n8557 2.2505
R35834 PAD.n8647 PAD.n8646 2.2505
R35835 PAD.n8643 PAD.n8642 2.2505
R35836 PAD.n8640 PAD.n8639 2.2505
R35837 PAD.n8632 PAD.n8559 2.2505
R35838 PAD.n8635 PAD.n8634 2.2505
R35839 PAD.n8631 PAD.n8630 2.2505
R35840 PAD.n8628 PAD.n8627 2.2505
R35841 PAD.n8620 PAD.n8561 2.2505
R35842 PAD.n8623 PAD.n8622 2.2505
R35843 PAD.n8619 PAD.n8618 2.2505
R35844 PAD.n8616 PAD.n8615 2.2505
R35845 PAD.n8608 PAD.n8563 2.2505
R35846 PAD.n8611 PAD.n8610 2.2505
R35847 PAD.n8607 PAD.n8606 2.2505
R35848 PAD.n8604 PAD.n8603 2.2505
R35849 PAD.n8596 PAD.n8565 2.2505
R35850 PAD.n8599 PAD.n8598 2.2505
R35851 PAD.n8595 PAD.n8594 2.2505
R35852 PAD.n8592 PAD.n8591 2.2505
R35853 PAD.n8584 PAD.n8567 2.2505
R35854 PAD.n8587 PAD.n8586 2.2505
R35855 PAD.n8583 PAD.n8582 2.2505
R35856 PAD.n8580 PAD.n8579 2.2505
R35857 PAD.n8572 PAD.n8569 2.2505
R35858 PAD.n8575 PAD.n8574 2.2505
R35859 PAD.n8571 PAD.n8570 2.2505
R35860 PAD.n8571 PAD.n2898 2.2505
R35861 PAD.n8576 PAD.n8575 2.2505
R35862 PAD.n8577 PAD.n8569 2.2505
R35863 PAD.n8579 PAD.n8578 2.2505
R35864 PAD.n8583 PAD.n8568 2.2505
R35865 PAD.n8588 PAD.n8587 2.2505
R35866 PAD.n8589 PAD.n8567 2.2505
R35867 PAD.n8591 PAD.n8590 2.2505
R35868 PAD.n8595 PAD.n8566 2.2505
R35869 PAD.n8600 PAD.n8599 2.2505
R35870 PAD.n8601 PAD.n8565 2.2505
R35871 PAD.n8603 PAD.n8602 2.2505
R35872 PAD.n8607 PAD.n8564 2.2505
R35873 PAD.n8612 PAD.n8611 2.2505
R35874 PAD.n8613 PAD.n8563 2.2505
R35875 PAD.n8615 PAD.n8614 2.2505
R35876 PAD.n8619 PAD.n8562 2.2505
R35877 PAD.n8624 PAD.n8623 2.2505
R35878 PAD.n8625 PAD.n8561 2.2505
R35879 PAD.n8627 PAD.n8626 2.2505
R35880 PAD.n8631 PAD.n8560 2.2505
R35881 PAD.n8636 PAD.n8635 2.2505
R35882 PAD.n8637 PAD.n8559 2.2505
R35883 PAD.n8639 PAD.n8638 2.2505
R35884 PAD.n8643 PAD.n8558 2.2505
R35885 PAD.n8648 PAD.n8647 2.2505
R35886 PAD.n8649 PAD.n8557 2.2505
R35887 PAD.n8651 PAD.n8650 2.2505
R35888 PAD.n8655 PAD.n8556 2.2505
R35889 PAD.n8660 PAD.n8659 2.2505
R35890 PAD.n8661 PAD.n8555 2.2505
R35891 PAD.n8663 PAD.n8662 2.2505
R35892 PAD.n8667 PAD.n8554 2.2505
R35893 PAD.n8672 PAD.n8671 2.2505
R35894 PAD.n8673 PAD.n8553 2.2505
R35895 PAD.n8675 PAD.n8674 2.2505
R35896 PAD.n8679 PAD.n8552 2.2505
R35897 PAD.n8684 PAD.n8683 2.2505
R35898 PAD.n8685 PAD.n8551 2.2505
R35899 PAD.n8687 PAD.n8686 2.2505
R35900 PAD.n8691 PAD.n8550 2.2505
R35901 PAD.n8696 PAD.n8695 2.2505
R35902 PAD.n8697 PAD.n8549 2.2505
R35903 PAD.n8699 PAD.n8698 2.2505
R35904 PAD.n8703 PAD.n8548 2.2505
R35905 PAD.n8708 PAD.n8707 2.2505
R35906 PAD.n8709 PAD.n8547 2.2505
R35907 PAD.n8711 PAD.n8710 2.2505
R35908 PAD.n8715 PAD.n8546 2.2505
R35909 PAD.n8720 PAD.n8719 2.2505
R35910 PAD.n8721 PAD.n8545 2.2505
R35911 PAD.n8723 PAD.n8722 2.2505
R35912 PAD.n8727 PAD.n8544 2.2505
R35913 PAD.n8732 PAD.n8731 2.2505
R35914 PAD.n8733 PAD.n8543 2.2505
R35915 PAD.n8735 PAD.n8734 2.2505
R35916 PAD.n8739 PAD.n8542 2.2505
R35917 PAD.n8744 PAD.n8743 2.2505
R35918 PAD.n8745 PAD.n8541 2.2505
R35919 PAD.n8747 PAD.n8746 2.2505
R35920 PAD.n8751 PAD.n8540 2.2505
R35921 PAD.n8756 PAD.n8755 2.2505
R35922 PAD.n8757 PAD.n8539 2.2505
R35923 PAD.n8759 PAD.n8758 2.2505
R35924 PAD.n8763 PAD.n8538 2.2505
R35925 PAD.n8768 PAD.n8767 2.2505
R35926 PAD.n8769 PAD.n8537 2.2505
R35927 PAD.n8771 PAD.n8770 2.2505
R35928 PAD.n8775 PAD.n8536 2.2505
R35929 PAD.n8780 PAD.n8779 2.2505
R35930 PAD.n8781 PAD.n8535 2.2505
R35931 PAD.n8783 PAD.n8782 2.2505
R35932 PAD.n8787 PAD.n8534 2.2505
R35933 PAD.n8792 PAD.n8791 2.2505
R35934 PAD.n8793 PAD.n8533 2.2505
R35935 PAD.n8795 PAD.n8794 2.2505
R35936 PAD.n8799 PAD.n8532 2.2505
R35937 PAD.n8804 PAD.n8803 2.2505
R35938 PAD.n8805 PAD.n8531 2.2505
R35939 PAD.n8807 PAD.n8806 2.2505
R35940 PAD.n8811 PAD.n8530 2.2505
R35941 PAD.n8815 PAD.n8814 2.2505
R35942 PAD.n8816 PAD.n8529 2.2505
R35943 PAD.n8818 PAD.n8817 2.2505
R35944 PAD.n3041 PAD.n2994 2.2505
R35945 PAD.n3040 PAD.n3039 2.2505
R35946 PAD.n3046 PAD.n3045 2.2505
R35947 PAD.n3049 PAD.n3048 2.2505
R35948 PAD.n3053 PAD.n3052 2.2505
R35949 PAD.n3050 PAD.n3036 2.2505
R35950 PAD.n3058 PAD.n3057 2.2505
R35951 PAD.n3061 PAD.n3060 2.2505
R35952 PAD.n3065 PAD.n3064 2.2505
R35953 PAD.n3062 PAD.n3034 2.2505
R35954 PAD.n3070 PAD.n3069 2.2505
R35955 PAD.n3073 PAD.n3072 2.2505
R35956 PAD.n3077 PAD.n3076 2.2505
R35957 PAD.n3074 PAD.n3032 2.2505
R35958 PAD.n3082 PAD.n3081 2.2505
R35959 PAD.n3085 PAD.n3084 2.2505
R35960 PAD.n3089 PAD.n3088 2.2505
R35961 PAD.n3086 PAD.n3030 2.2505
R35962 PAD.n3094 PAD.n3093 2.2505
R35963 PAD.n3097 PAD.n3096 2.2505
R35964 PAD.n3101 PAD.n3100 2.2505
R35965 PAD.n3098 PAD.n3028 2.2505
R35966 PAD.n3106 PAD.n3105 2.2505
R35967 PAD.n3109 PAD.n3108 2.2505
R35968 PAD.n3113 PAD.n3112 2.2505
R35969 PAD.n3110 PAD.n3026 2.2505
R35970 PAD.n3118 PAD.n3117 2.2505
R35971 PAD.n3121 PAD.n3120 2.2505
R35972 PAD.n3125 PAD.n3124 2.2505
R35973 PAD.n3122 PAD.n3024 2.2505
R35974 PAD.n3130 PAD.n3129 2.2505
R35975 PAD.n3133 PAD.n3132 2.2505
R35976 PAD.n3137 PAD.n3136 2.2505
R35977 PAD.n3134 PAD.n3022 2.2505
R35978 PAD.n3142 PAD.n3141 2.2505
R35979 PAD.n3145 PAD.n3144 2.2505
R35980 PAD.n3149 PAD.n3148 2.2505
R35981 PAD.n3146 PAD.n3020 2.2505
R35982 PAD.n3154 PAD.n3153 2.2505
R35983 PAD.n3157 PAD.n3156 2.2505
R35984 PAD.n3161 PAD.n3160 2.2505
R35985 PAD.n3158 PAD.n3018 2.2505
R35986 PAD.n3166 PAD.n3165 2.2505
R35987 PAD.n3169 PAD.n3168 2.2505
R35988 PAD.n3173 PAD.n3172 2.2505
R35989 PAD.n3170 PAD.n3016 2.2505
R35990 PAD.n3178 PAD.n3177 2.2505
R35991 PAD.n3181 PAD.n3180 2.2505
R35992 PAD.n3185 PAD.n3184 2.2505
R35993 PAD.n3182 PAD.n3014 2.2505
R35994 PAD.n3190 PAD.n3189 2.2505
R35995 PAD.n3193 PAD.n3192 2.2505
R35996 PAD.n3197 PAD.n3196 2.2505
R35997 PAD.n3194 PAD.n3012 2.2505
R35998 PAD.n3202 PAD.n3201 2.2505
R35999 PAD.n3205 PAD.n3204 2.2505
R36000 PAD.n3209 PAD.n3208 2.2505
R36001 PAD.n3206 PAD.n3010 2.2505
R36002 PAD.n3214 PAD.n3213 2.2505
R36003 PAD.n3217 PAD.n3216 2.2505
R36004 PAD.n3221 PAD.n3220 2.2505
R36005 PAD.n3218 PAD.n3008 2.2505
R36006 PAD.n3226 PAD.n3225 2.2505
R36007 PAD.n3229 PAD.n3228 2.2505
R36008 PAD.n3233 PAD.n3232 2.2505
R36009 PAD.n3230 PAD.n3006 2.2505
R36010 PAD.n3238 PAD.n3237 2.2505
R36011 PAD.n3241 PAD.n3240 2.2505
R36012 PAD.n3245 PAD.n3244 2.2505
R36013 PAD.n3242 PAD.n3004 2.2505
R36014 PAD.n3250 PAD.n3249 2.2505
R36015 PAD.n3253 PAD.n3252 2.2505
R36016 PAD.n3257 PAD.n3256 2.2505
R36017 PAD.n3254 PAD.n3002 2.2505
R36018 PAD.n3262 PAD.n3261 2.2505
R36019 PAD.n3265 PAD.n3264 2.2505
R36020 PAD.n3269 PAD.n3268 2.2505
R36021 PAD.n3266 PAD.n3000 2.2505
R36022 PAD.n3274 PAD.n3273 2.2505
R36023 PAD.n3277 PAD.n3276 2.2505
R36024 PAD.n3281 PAD.n3280 2.2505
R36025 PAD.n3278 PAD.n2998 2.2505
R36026 PAD.n8514 PAD.n8513 2.2505
R36027 PAD.n8516 PAD.n2995 2.2505
R36028 PAD.n8511 PAD.n2995 2.2505
R36029 PAD.n8513 PAD.n8512 2.2505
R36030 PAD.n3283 PAD.n2998 2.2505
R36031 PAD.n3282 PAD.n3281 2.2505
R36032 PAD.n3277 PAD.n2999 2.2505
R36033 PAD.n3273 PAD.n3272 2.2505
R36034 PAD.n3271 PAD.n3000 2.2505
R36035 PAD.n3270 PAD.n3269 2.2505
R36036 PAD.n3265 PAD.n3001 2.2505
R36037 PAD.n3261 PAD.n3260 2.2505
R36038 PAD.n3259 PAD.n3002 2.2505
R36039 PAD.n3258 PAD.n3257 2.2505
R36040 PAD.n3253 PAD.n3003 2.2505
R36041 PAD.n3249 PAD.n3248 2.2505
R36042 PAD.n3247 PAD.n3004 2.2505
R36043 PAD.n3246 PAD.n3245 2.2505
R36044 PAD.n3241 PAD.n3005 2.2505
R36045 PAD.n3237 PAD.n3236 2.2505
R36046 PAD.n3235 PAD.n3006 2.2505
R36047 PAD.n3234 PAD.n3233 2.2505
R36048 PAD.n3229 PAD.n3007 2.2505
R36049 PAD.n3225 PAD.n3224 2.2505
R36050 PAD.n3223 PAD.n3008 2.2505
R36051 PAD.n3222 PAD.n3221 2.2505
R36052 PAD.n3217 PAD.n3009 2.2505
R36053 PAD.n3213 PAD.n3212 2.2505
R36054 PAD.n3211 PAD.n3010 2.2505
R36055 PAD.n3210 PAD.n3209 2.2505
R36056 PAD.n3205 PAD.n3011 2.2505
R36057 PAD.n3201 PAD.n3200 2.2505
R36058 PAD.n3199 PAD.n3012 2.2505
R36059 PAD.n3198 PAD.n3197 2.2505
R36060 PAD.n3193 PAD.n3013 2.2505
R36061 PAD.n3189 PAD.n3188 2.2505
R36062 PAD.n3187 PAD.n3014 2.2505
R36063 PAD.n3186 PAD.n3185 2.2505
R36064 PAD.n3181 PAD.n3015 2.2505
R36065 PAD.n3177 PAD.n3176 2.2505
R36066 PAD.n3175 PAD.n3016 2.2505
R36067 PAD.n3174 PAD.n3173 2.2505
R36068 PAD.n3169 PAD.n3017 2.2505
R36069 PAD.n3165 PAD.n3164 2.2505
R36070 PAD.n3163 PAD.n3018 2.2505
R36071 PAD.n3162 PAD.n3161 2.2505
R36072 PAD.n3157 PAD.n3019 2.2505
R36073 PAD.n3153 PAD.n3152 2.2505
R36074 PAD.n3151 PAD.n3020 2.2505
R36075 PAD.n3150 PAD.n3149 2.2505
R36076 PAD.n3145 PAD.n3021 2.2505
R36077 PAD.n3141 PAD.n3140 2.2505
R36078 PAD.n3139 PAD.n3022 2.2505
R36079 PAD.n3138 PAD.n3137 2.2505
R36080 PAD.n3133 PAD.n3023 2.2505
R36081 PAD.n3129 PAD.n3128 2.2505
R36082 PAD.n3127 PAD.n3024 2.2505
R36083 PAD.n3126 PAD.n3125 2.2505
R36084 PAD.n3121 PAD.n3025 2.2505
R36085 PAD.n3117 PAD.n3116 2.2505
R36086 PAD.n3115 PAD.n3026 2.2505
R36087 PAD.n3114 PAD.n3113 2.2505
R36088 PAD.n3109 PAD.n3027 2.2505
R36089 PAD.n3105 PAD.n3104 2.2505
R36090 PAD.n3103 PAD.n3028 2.2505
R36091 PAD.n3102 PAD.n3101 2.2505
R36092 PAD.n3097 PAD.n3029 2.2505
R36093 PAD.n3093 PAD.n3092 2.2505
R36094 PAD.n3091 PAD.n3030 2.2505
R36095 PAD.n3090 PAD.n3089 2.2505
R36096 PAD.n3085 PAD.n3031 2.2505
R36097 PAD.n3081 PAD.n3080 2.2505
R36098 PAD.n3079 PAD.n3032 2.2505
R36099 PAD.n3078 PAD.n3077 2.2505
R36100 PAD.n3073 PAD.n3033 2.2505
R36101 PAD.n3069 PAD.n3068 2.2505
R36102 PAD.n3067 PAD.n3034 2.2505
R36103 PAD.n3066 PAD.n3065 2.2505
R36104 PAD.n3061 PAD.n3035 2.2505
R36105 PAD.n3057 PAD.n3056 2.2505
R36106 PAD.n3055 PAD.n3036 2.2505
R36107 PAD.n3054 PAD.n3053 2.2505
R36108 PAD.n3049 PAD.n3037 2.2505
R36109 PAD.n3045 PAD.n3044 2.2505
R36110 PAD.n3043 PAD.n3040 2.2505
R36111 PAD.n3042 PAD.n3041 2.2505
R36112 PAD.n3386 PAD.n3338 2.2505
R36113 PAD.n3385 PAD.n3384 2.2505
R36114 PAD.n3391 PAD.n3390 2.2505
R36115 PAD.n3394 PAD.n3393 2.2505
R36116 PAD.n3398 PAD.n3397 2.2505
R36117 PAD.n3395 PAD.n3381 2.2505
R36118 PAD.n3403 PAD.n3402 2.2505
R36119 PAD.n3406 PAD.n3405 2.2505
R36120 PAD.n3410 PAD.n3409 2.2505
R36121 PAD.n3407 PAD.n3379 2.2505
R36122 PAD.n3415 PAD.n3414 2.2505
R36123 PAD.n3418 PAD.n3417 2.2505
R36124 PAD.n3422 PAD.n3421 2.2505
R36125 PAD.n3419 PAD.n3377 2.2505
R36126 PAD.n3427 PAD.n3426 2.2505
R36127 PAD.n3430 PAD.n3429 2.2505
R36128 PAD.n3434 PAD.n3433 2.2505
R36129 PAD.n3431 PAD.n3375 2.2505
R36130 PAD.n3439 PAD.n3438 2.2505
R36131 PAD.n3442 PAD.n3441 2.2505
R36132 PAD.n3446 PAD.n3445 2.2505
R36133 PAD.n3443 PAD.n3373 2.2505
R36134 PAD.n3451 PAD.n3450 2.2505
R36135 PAD.n3454 PAD.n3453 2.2505
R36136 PAD.n3458 PAD.n3457 2.2505
R36137 PAD.n3455 PAD.n3371 2.2505
R36138 PAD.n3463 PAD.n3462 2.2505
R36139 PAD.n3466 PAD.n3465 2.2505
R36140 PAD.n3470 PAD.n3469 2.2505
R36141 PAD.n3467 PAD.n3369 2.2505
R36142 PAD.n3475 PAD.n3474 2.2505
R36143 PAD.n3478 PAD.n3477 2.2505
R36144 PAD.n3482 PAD.n3481 2.2505
R36145 PAD.n3479 PAD.n3367 2.2505
R36146 PAD.n3487 PAD.n3486 2.2505
R36147 PAD.n3490 PAD.n3489 2.2505
R36148 PAD.n3494 PAD.n3493 2.2505
R36149 PAD.n3491 PAD.n3365 2.2505
R36150 PAD.n3499 PAD.n3498 2.2505
R36151 PAD.n3502 PAD.n3501 2.2505
R36152 PAD.n3506 PAD.n3505 2.2505
R36153 PAD.n3503 PAD.n3363 2.2505
R36154 PAD.n3511 PAD.n3510 2.2505
R36155 PAD.n3514 PAD.n3513 2.2505
R36156 PAD.n3518 PAD.n3517 2.2505
R36157 PAD.n3515 PAD.n3361 2.2505
R36158 PAD.n3523 PAD.n3522 2.2505
R36159 PAD.n3526 PAD.n3525 2.2505
R36160 PAD.n3530 PAD.n3529 2.2505
R36161 PAD.n3527 PAD.n3359 2.2505
R36162 PAD.n3535 PAD.n3534 2.2505
R36163 PAD.n3538 PAD.n3537 2.2505
R36164 PAD.n3542 PAD.n3541 2.2505
R36165 PAD.n3539 PAD.n3357 2.2505
R36166 PAD.n3547 PAD.n3546 2.2505
R36167 PAD.n3550 PAD.n3549 2.2505
R36168 PAD.n3554 PAD.n3553 2.2505
R36169 PAD.n3551 PAD.n3355 2.2505
R36170 PAD.n3559 PAD.n3558 2.2505
R36171 PAD.n3562 PAD.n3561 2.2505
R36172 PAD.n3566 PAD.n3565 2.2505
R36173 PAD.n3563 PAD.n3353 2.2505
R36174 PAD.n3571 PAD.n3570 2.2505
R36175 PAD.n3574 PAD.n3573 2.2505
R36176 PAD.n3578 PAD.n3577 2.2505
R36177 PAD.n3575 PAD.n3351 2.2505
R36178 PAD.n3583 PAD.n3582 2.2505
R36179 PAD.n3586 PAD.n3585 2.2505
R36180 PAD.n3590 PAD.n3589 2.2505
R36181 PAD.n3587 PAD.n3349 2.2505
R36182 PAD.n3595 PAD.n3594 2.2505
R36183 PAD.n3598 PAD.n3597 2.2505
R36184 PAD.n3602 PAD.n3601 2.2505
R36185 PAD.n3599 PAD.n3347 2.2505
R36186 PAD.n3607 PAD.n3606 2.2505
R36187 PAD.n3610 PAD.n3609 2.2505
R36188 PAD.n3614 PAD.n3613 2.2505
R36189 PAD.n3611 PAD.n3345 2.2505
R36190 PAD.n3619 PAD.n3618 2.2505
R36191 PAD.n3622 PAD.n3621 2.2505
R36192 PAD.n3626 PAD.n3625 2.2505
R36193 PAD.n3623 PAD.n3343 2.2505
R36194 PAD.n8489 PAD.n8488 2.2505
R36195 PAD.n8491 PAD.n3340 2.2505
R36196 PAD.n8486 PAD.n3340 2.2505
R36197 PAD.n8488 PAD.n8487 2.2505
R36198 PAD.n3628 PAD.n3343 2.2505
R36199 PAD.n3627 PAD.n3626 2.2505
R36200 PAD.n3622 PAD.n3344 2.2505
R36201 PAD.n3618 PAD.n3617 2.2505
R36202 PAD.n3616 PAD.n3345 2.2505
R36203 PAD.n3615 PAD.n3614 2.2505
R36204 PAD.n3610 PAD.n3346 2.2505
R36205 PAD.n3606 PAD.n3605 2.2505
R36206 PAD.n3604 PAD.n3347 2.2505
R36207 PAD.n3603 PAD.n3602 2.2505
R36208 PAD.n3598 PAD.n3348 2.2505
R36209 PAD.n3594 PAD.n3593 2.2505
R36210 PAD.n3592 PAD.n3349 2.2505
R36211 PAD.n3591 PAD.n3590 2.2505
R36212 PAD.n3586 PAD.n3350 2.2505
R36213 PAD.n3582 PAD.n3581 2.2505
R36214 PAD.n3580 PAD.n3351 2.2505
R36215 PAD.n3579 PAD.n3578 2.2505
R36216 PAD.n3574 PAD.n3352 2.2505
R36217 PAD.n3570 PAD.n3569 2.2505
R36218 PAD.n3568 PAD.n3353 2.2505
R36219 PAD.n3567 PAD.n3566 2.2505
R36220 PAD.n3562 PAD.n3354 2.2505
R36221 PAD.n3558 PAD.n3557 2.2505
R36222 PAD.n3556 PAD.n3355 2.2505
R36223 PAD.n3555 PAD.n3554 2.2505
R36224 PAD.n3550 PAD.n3356 2.2505
R36225 PAD.n3546 PAD.n3545 2.2505
R36226 PAD.n3544 PAD.n3357 2.2505
R36227 PAD.n3543 PAD.n3542 2.2505
R36228 PAD.n3538 PAD.n3358 2.2505
R36229 PAD.n3534 PAD.n3533 2.2505
R36230 PAD.n3532 PAD.n3359 2.2505
R36231 PAD.n3531 PAD.n3530 2.2505
R36232 PAD.n3526 PAD.n3360 2.2505
R36233 PAD.n3522 PAD.n3521 2.2505
R36234 PAD.n3520 PAD.n3361 2.2505
R36235 PAD.n3519 PAD.n3518 2.2505
R36236 PAD.n3514 PAD.n3362 2.2505
R36237 PAD.n3510 PAD.n3509 2.2505
R36238 PAD.n3508 PAD.n3363 2.2505
R36239 PAD.n3507 PAD.n3506 2.2505
R36240 PAD.n3502 PAD.n3364 2.2505
R36241 PAD.n3498 PAD.n3497 2.2505
R36242 PAD.n3496 PAD.n3365 2.2505
R36243 PAD.n3495 PAD.n3494 2.2505
R36244 PAD.n3490 PAD.n3366 2.2505
R36245 PAD.n3486 PAD.n3485 2.2505
R36246 PAD.n3484 PAD.n3367 2.2505
R36247 PAD.n3483 PAD.n3482 2.2505
R36248 PAD.n3478 PAD.n3368 2.2505
R36249 PAD.n3474 PAD.n3473 2.2505
R36250 PAD.n3472 PAD.n3369 2.2505
R36251 PAD.n3471 PAD.n3470 2.2505
R36252 PAD.n3466 PAD.n3370 2.2505
R36253 PAD.n3462 PAD.n3461 2.2505
R36254 PAD.n3460 PAD.n3371 2.2505
R36255 PAD.n3459 PAD.n3458 2.2505
R36256 PAD.n3454 PAD.n3372 2.2505
R36257 PAD.n3450 PAD.n3449 2.2505
R36258 PAD.n3448 PAD.n3373 2.2505
R36259 PAD.n3447 PAD.n3446 2.2505
R36260 PAD.n3442 PAD.n3374 2.2505
R36261 PAD.n3438 PAD.n3437 2.2505
R36262 PAD.n3436 PAD.n3375 2.2505
R36263 PAD.n3435 PAD.n3434 2.2505
R36264 PAD.n3430 PAD.n3376 2.2505
R36265 PAD.n3426 PAD.n3425 2.2505
R36266 PAD.n3424 PAD.n3377 2.2505
R36267 PAD.n3423 PAD.n3422 2.2505
R36268 PAD.n3418 PAD.n3378 2.2505
R36269 PAD.n3414 PAD.n3413 2.2505
R36270 PAD.n3412 PAD.n3379 2.2505
R36271 PAD.n3411 PAD.n3410 2.2505
R36272 PAD.n3406 PAD.n3380 2.2505
R36273 PAD.n3402 PAD.n3401 2.2505
R36274 PAD.n3400 PAD.n3381 2.2505
R36275 PAD.n3399 PAD.n3398 2.2505
R36276 PAD.n3394 PAD.n3382 2.2505
R36277 PAD.n3390 PAD.n3389 2.2505
R36278 PAD.n3388 PAD.n3385 2.2505
R36279 PAD.n3387 PAD.n3386 2.2505
R36280 PAD.n3731 PAD.n3683 2.2505
R36281 PAD.n3730 PAD.n3729 2.2505
R36282 PAD.n3736 PAD.n3735 2.2505
R36283 PAD.n3739 PAD.n3738 2.2505
R36284 PAD.n3743 PAD.n3742 2.2505
R36285 PAD.n3740 PAD.n3726 2.2505
R36286 PAD.n3748 PAD.n3747 2.2505
R36287 PAD.n3751 PAD.n3750 2.2505
R36288 PAD.n3755 PAD.n3754 2.2505
R36289 PAD.n3752 PAD.n3724 2.2505
R36290 PAD.n3760 PAD.n3759 2.2505
R36291 PAD.n3763 PAD.n3762 2.2505
R36292 PAD.n3767 PAD.n3766 2.2505
R36293 PAD.n3764 PAD.n3722 2.2505
R36294 PAD.n3772 PAD.n3771 2.2505
R36295 PAD.n3775 PAD.n3774 2.2505
R36296 PAD.n3779 PAD.n3778 2.2505
R36297 PAD.n3776 PAD.n3720 2.2505
R36298 PAD.n3784 PAD.n3783 2.2505
R36299 PAD.n3787 PAD.n3786 2.2505
R36300 PAD.n3791 PAD.n3790 2.2505
R36301 PAD.n3788 PAD.n3718 2.2505
R36302 PAD.n3796 PAD.n3795 2.2505
R36303 PAD.n3799 PAD.n3798 2.2505
R36304 PAD.n3803 PAD.n3802 2.2505
R36305 PAD.n3800 PAD.n3716 2.2505
R36306 PAD.n3808 PAD.n3807 2.2505
R36307 PAD.n3811 PAD.n3810 2.2505
R36308 PAD.n3815 PAD.n3814 2.2505
R36309 PAD.n3812 PAD.n3714 2.2505
R36310 PAD.n3820 PAD.n3819 2.2505
R36311 PAD.n3823 PAD.n3822 2.2505
R36312 PAD.n3827 PAD.n3826 2.2505
R36313 PAD.n3824 PAD.n3712 2.2505
R36314 PAD.n3832 PAD.n3831 2.2505
R36315 PAD.n3835 PAD.n3834 2.2505
R36316 PAD.n3839 PAD.n3838 2.2505
R36317 PAD.n3836 PAD.n3710 2.2505
R36318 PAD.n3844 PAD.n3843 2.2505
R36319 PAD.n3847 PAD.n3846 2.2505
R36320 PAD.n3851 PAD.n3850 2.2505
R36321 PAD.n3848 PAD.n3708 2.2505
R36322 PAD.n3856 PAD.n3855 2.2505
R36323 PAD.n3859 PAD.n3858 2.2505
R36324 PAD.n3863 PAD.n3862 2.2505
R36325 PAD.n3860 PAD.n3706 2.2505
R36326 PAD.n3868 PAD.n3867 2.2505
R36327 PAD.n3871 PAD.n3870 2.2505
R36328 PAD.n3875 PAD.n3874 2.2505
R36329 PAD.n3872 PAD.n3704 2.2505
R36330 PAD.n3880 PAD.n3879 2.2505
R36331 PAD.n3883 PAD.n3882 2.2505
R36332 PAD.n3887 PAD.n3886 2.2505
R36333 PAD.n3884 PAD.n3702 2.2505
R36334 PAD.n3892 PAD.n3891 2.2505
R36335 PAD.n3895 PAD.n3894 2.2505
R36336 PAD.n3899 PAD.n3898 2.2505
R36337 PAD.n3896 PAD.n3700 2.2505
R36338 PAD.n3904 PAD.n3903 2.2505
R36339 PAD.n3907 PAD.n3906 2.2505
R36340 PAD.n3911 PAD.n3910 2.2505
R36341 PAD.n3908 PAD.n3698 2.2505
R36342 PAD.n3916 PAD.n3915 2.2505
R36343 PAD.n3919 PAD.n3918 2.2505
R36344 PAD.n3923 PAD.n3922 2.2505
R36345 PAD.n3920 PAD.n3696 2.2505
R36346 PAD.n3928 PAD.n3927 2.2505
R36347 PAD.n3931 PAD.n3930 2.2505
R36348 PAD.n3935 PAD.n3934 2.2505
R36349 PAD.n3932 PAD.n3694 2.2505
R36350 PAD.n3940 PAD.n3939 2.2505
R36351 PAD.n3943 PAD.n3942 2.2505
R36352 PAD.n3947 PAD.n3946 2.2505
R36353 PAD.n3944 PAD.n3692 2.2505
R36354 PAD.n3952 PAD.n3951 2.2505
R36355 PAD.n3955 PAD.n3954 2.2505
R36356 PAD.n3959 PAD.n3958 2.2505
R36357 PAD.n3956 PAD.n3690 2.2505
R36358 PAD.n3964 PAD.n3963 2.2505
R36359 PAD.n3967 PAD.n3966 2.2505
R36360 PAD.n3971 PAD.n3970 2.2505
R36361 PAD.n3968 PAD.n3688 2.2505
R36362 PAD.n8465 PAD.n8464 2.2505
R36363 PAD.n8467 PAD.n3685 2.2505
R36364 PAD.n8462 PAD.n3685 2.2505
R36365 PAD.n8464 PAD.n8463 2.2505
R36366 PAD.n3973 PAD.n3688 2.2505
R36367 PAD.n3972 PAD.n3971 2.2505
R36368 PAD.n3967 PAD.n3689 2.2505
R36369 PAD.n3963 PAD.n3962 2.2505
R36370 PAD.n3961 PAD.n3690 2.2505
R36371 PAD.n3960 PAD.n3959 2.2505
R36372 PAD.n3955 PAD.n3691 2.2505
R36373 PAD.n3951 PAD.n3950 2.2505
R36374 PAD.n3949 PAD.n3692 2.2505
R36375 PAD.n3948 PAD.n3947 2.2505
R36376 PAD.n3943 PAD.n3693 2.2505
R36377 PAD.n3939 PAD.n3938 2.2505
R36378 PAD.n3937 PAD.n3694 2.2505
R36379 PAD.n3936 PAD.n3935 2.2505
R36380 PAD.n3931 PAD.n3695 2.2505
R36381 PAD.n3927 PAD.n3926 2.2505
R36382 PAD.n3925 PAD.n3696 2.2505
R36383 PAD.n3924 PAD.n3923 2.2505
R36384 PAD.n3919 PAD.n3697 2.2505
R36385 PAD.n3915 PAD.n3914 2.2505
R36386 PAD.n3913 PAD.n3698 2.2505
R36387 PAD.n3912 PAD.n3911 2.2505
R36388 PAD.n3907 PAD.n3699 2.2505
R36389 PAD.n3903 PAD.n3902 2.2505
R36390 PAD.n3901 PAD.n3700 2.2505
R36391 PAD.n3900 PAD.n3899 2.2505
R36392 PAD.n3895 PAD.n3701 2.2505
R36393 PAD.n3891 PAD.n3890 2.2505
R36394 PAD.n3889 PAD.n3702 2.2505
R36395 PAD.n3888 PAD.n3887 2.2505
R36396 PAD.n3883 PAD.n3703 2.2505
R36397 PAD.n3879 PAD.n3878 2.2505
R36398 PAD.n3877 PAD.n3704 2.2505
R36399 PAD.n3876 PAD.n3875 2.2505
R36400 PAD.n3871 PAD.n3705 2.2505
R36401 PAD.n3867 PAD.n3866 2.2505
R36402 PAD.n3865 PAD.n3706 2.2505
R36403 PAD.n3864 PAD.n3863 2.2505
R36404 PAD.n3859 PAD.n3707 2.2505
R36405 PAD.n3855 PAD.n3854 2.2505
R36406 PAD.n3853 PAD.n3708 2.2505
R36407 PAD.n3852 PAD.n3851 2.2505
R36408 PAD.n3847 PAD.n3709 2.2505
R36409 PAD.n3843 PAD.n3842 2.2505
R36410 PAD.n3841 PAD.n3710 2.2505
R36411 PAD.n3840 PAD.n3839 2.2505
R36412 PAD.n3835 PAD.n3711 2.2505
R36413 PAD.n3831 PAD.n3830 2.2505
R36414 PAD.n3829 PAD.n3712 2.2505
R36415 PAD.n3828 PAD.n3827 2.2505
R36416 PAD.n3823 PAD.n3713 2.2505
R36417 PAD.n3819 PAD.n3818 2.2505
R36418 PAD.n3817 PAD.n3714 2.2505
R36419 PAD.n3816 PAD.n3815 2.2505
R36420 PAD.n3811 PAD.n3715 2.2505
R36421 PAD.n3807 PAD.n3806 2.2505
R36422 PAD.n3805 PAD.n3716 2.2505
R36423 PAD.n3804 PAD.n3803 2.2505
R36424 PAD.n3799 PAD.n3717 2.2505
R36425 PAD.n3795 PAD.n3794 2.2505
R36426 PAD.n3793 PAD.n3718 2.2505
R36427 PAD.n3792 PAD.n3791 2.2505
R36428 PAD.n3787 PAD.n3719 2.2505
R36429 PAD.n3783 PAD.n3782 2.2505
R36430 PAD.n3781 PAD.n3720 2.2505
R36431 PAD.n3780 PAD.n3779 2.2505
R36432 PAD.n3775 PAD.n3721 2.2505
R36433 PAD.n3771 PAD.n3770 2.2505
R36434 PAD.n3769 PAD.n3722 2.2505
R36435 PAD.n3768 PAD.n3767 2.2505
R36436 PAD.n3763 PAD.n3723 2.2505
R36437 PAD.n3759 PAD.n3758 2.2505
R36438 PAD.n3757 PAD.n3724 2.2505
R36439 PAD.n3756 PAD.n3755 2.2505
R36440 PAD.n3751 PAD.n3725 2.2505
R36441 PAD.n3747 PAD.n3746 2.2505
R36442 PAD.n3745 PAD.n3726 2.2505
R36443 PAD.n3744 PAD.n3743 2.2505
R36444 PAD.n3739 PAD.n3727 2.2505
R36445 PAD.n3735 PAD.n3734 2.2505
R36446 PAD.n3733 PAD.n3730 2.2505
R36447 PAD.n3732 PAD.n3731 2.2505
R36448 PAD.n4072 PAD.n4025 2.2505
R36449 PAD.n4071 PAD.n4070 2.2505
R36450 PAD.n4077 PAD.n4076 2.2505
R36451 PAD.n4080 PAD.n4079 2.2505
R36452 PAD.n4084 PAD.n4083 2.2505
R36453 PAD.n4081 PAD.n4067 2.2505
R36454 PAD.n4089 PAD.n4088 2.2505
R36455 PAD.n4092 PAD.n4091 2.2505
R36456 PAD.n4096 PAD.n4095 2.2505
R36457 PAD.n4093 PAD.n4065 2.2505
R36458 PAD.n4101 PAD.n4100 2.2505
R36459 PAD.n4104 PAD.n4103 2.2505
R36460 PAD.n4108 PAD.n4107 2.2505
R36461 PAD.n4105 PAD.n4063 2.2505
R36462 PAD.n4113 PAD.n4112 2.2505
R36463 PAD.n4116 PAD.n4115 2.2505
R36464 PAD.n4120 PAD.n4119 2.2505
R36465 PAD.n4117 PAD.n4061 2.2505
R36466 PAD.n4125 PAD.n4124 2.2505
R36467 PAD.n4128 PAD.n4127 2.2505
R36468 PAD.n4132 PAD.n4131 2.2505
R36469 PAD.n4129 PAD.n4059 2.2505
R36470 PAD.n4137 PAD.n4136 2.2505
R36471 PAD.n4140 PAD.n4139 2.2505
R36472 PAD.n4144 PAD.n4143 2.2505
R36473 PAD.n4141 PAD.n4057 2.2505
R36474 PAD.n4149 PAD.n4148 2.2505
R36475 PAD.n4152 PAD.n4151 2.2505
R36476 PAD.n4156 PAD.n4155 2.2505
R36477 PAD.n4153 PAD.n4055 2.2505
R36478 PAD.n4161 PAD.n4160 2.2505
R36479 PAD.n4164 PAD.n4163 2.2505
R36480 PAD.n4168 PAD.n4167 2.2505
R36481 PAD.n4165 PAD.n4053 2.2505
R36482 PAD.n4173 PAD.n4172 2.2505
R36483 PAD.n4176 PAD.n4175 2.2505
R36484 PAD.n4180 PAD.n4179 2.2505
R36485 PAD.n4177 PAD.n4051 2.2505
R36486 PAD.n4185 PAD.n4184 2.2505
R36487 PAD.n4188 PAD.n4187 2.2505
R36488 PAD.n4192 PAD.n4191 2.2505
R36489 PAD.n4189 PAD.n4049 2.2505
R36490 PAD.n4197 PAD.n4196 2.2505
R36491 PAD.n4200 PAD.n4199 2.2505
R36492 PAD.n4204 PAD.n4203 2.2505
R36493 PAD.n4201 PAD.n4047 2.2505
R36494 PAD.n4209 PAD.n4208 2.2505
R36495 PAD.n4212 PAD.n4211 2.2505
R36496 PAD.n4216 PAD.n4215 2.2505
R36497 PAD.n4213 PAD.n4045 2.2505
R36498 PAD.n4221 PAD.n4220 2.2505
R36499 PAD.n4224 PAD.n4223 2.2505
R36500 PAD.n4228 PAD.n4227 2.2505
R36501 PAD.n4225 PAD.n4043 2.2505
R36502 PAD.n4233 PAD.n4232 2.2505
R36503 PAD.n4236 PAD.n4235 2.2505
R36504 PAD.n4240 PAD.n4239 2.2505
R36505 PAD.n4237 PAD.n4041 2.2505
R36506 PAD.n4245 PAD.n4244 2.2505
R36507 PAD.n4248 PAD.n4247 2.2505
R36508 PAD.n4252 PAD.n4251 2.2505
R36509 PAD.n4249 PAD.n4039 2.2505
R36510 PAD.n4257 PAD.n4256 2.2505
R36511 PAD.n4260 PAD.n4259 2.2505
R36512 PAD.n4264 PAD.n4263 2.2505
R36513 PAD.n4261 PAD.n4037 2.2505
R36514 PAD.n4269 PAD.n4268 2.2505
R36515 PAD.n4272 PAD.n4271 2.2505
R36516 PAD.n4276 PAD.n4275 2.2505
R36517 PAD.n4273 PAD.n4035 2.2505
R36518 PAD.n4281 PAD.n4280 2.2505
R36519 PAD.n4284 PAD.n4283 2.2505
R36520 PAD.n4288 PAD.n4287 2.2505
R36521 PAD.n4285 PAD.n4033 2.2505
R36522 PAD.n4293 PAD.n4292 2.2505
R36523 PAD.n4296 PAD.n4295 2.2505
R36524 PAD.n4300 PAD.n4299 2.2505
R36525 PAD.n4297 PAD.n4031 2.2505
R36526 PAD.n4305 PAD.n4304 2.2505
R36527 PAD.n4308 PAD.n4307 2.2505
R36528 PAD.n4312 PAD.n4311 2.2505
R36529 PAD.n4309 PAD.n4029 2.2505
R36530 PAD.n8441 PAD.n8440 2.2505
R36531 PAD.n8443 PAD.n4026 2.2505
R36532 PAD.n8438 PAD.n4026 2.2505
R36533 PAD.n8440 PAD.n8439 2.2505
R36534 PAD.n4314 PAD.n4029 2.2505
R36535 PAD.n4313 PAD.n4312 2.2505
R36536 PAD.n4308 PAD.n4030 2.2505
R36537 PAD.n4304 PAD.n4303 2.2505
R36538 PAD.n4302 PAD.n4031 2.2505
R36539 PAD.n4301 PAD.n4300 2.2505
R36540 PAD.n4296 PAD.n4032 2.2505
R36541 PAD.n4292 PAD.n4291 2.2505
R36542 PAD.n4290 PAD.n4033 2.2505
R36543 PAD.n4289 PAD.n4288 2.2505
R36544 PAD.n4284 PAD.n4034 2.2505
R36545 PAD.n4280 PAD.n4279 2.2505
R36546 PAD.n4278 PAD.n4035 2.2505
R36547 PAD.n4277 PAD.n4276 2.2505
R36548 PAD.n4272 PAD.n4036 2.2505
R36549 PAD.n4268 PAD.n4267 2.2505
R36550 PAD.n4266 PAD.n4037 2.2505
R36551 PAD.n4265 PAD.n4264 2.2505
R36552 PAD.n4260 PAD.n4038 2.2505
R36553 PAD.n4256 PAD.n4255 2.2505
R36554 PAD.n4254 PAD.n4039 2.2505
R36555 PAD.n4253 PAD.n4252 2.2505
R36556 PAD.n4248 PAD.n4040 2.2505
R36557 PAD.n4244 PAD.n4243 2.2505
R36558 PAD.n4242 PAD.n4041 2.2505
R36559 PAD.n4241 PAD.n4240 2.2505
R36560 PAD.n4236 PAD.n4042 2.2505
R36561 PAD.n4232 PAD.n4231 2.2505
R36562 PAD.n4230 PAD.n4043 2.2505
R36563 PAD.n4229 PAD.n4228 2.2505
R36564 PAD.n4224 PAD.n4044 2.2505
R36565 PAD.n4220 PAD.n4219 2.2505
R36566 PAD.n4218 PAD.n4045 2.2505
R36567 PAD.n4217 PAD.n4216 2.2505
R36568 PAD.n4212 PAD.n4046 2.2505
R36569 PAD.n4208 PAD.n4207 2.2505
R36570 PAD.n4206 PAD.n4047 2.2505
R36571 PAD.n4205 PAD.n4204 2.2505
R36572 PAD.n4200 PAD.n4048 2.2505
R36573 PAD.n4196 PAD.n4195 2.2505
R36574 PAD.n4194 PAD.n4049 2.2505
R36575 PAD.n4193 PAD.n4192 2.2505
R36576 PAD.n4188 PAD.n4050 2.2505
R36577 PAD.n4184 PAD.n4183 2.2505
R36578 PAD.n4182 PAD.n4051 2.2505
R36579 PAD.n4181 PAD.n4180 2.2505
R36580 PAD.n4176 PAD.n4052 2.2505
R36581 PAD.n4172 PAD.n4171 2.2505
R36582 PAD.n4170 PAD.n4053 2.2505
R36583 PAD.n4169 PAD.n4168 2.2505
R36584 PAD.n4164 PAD.n4054 2.2505
R36585 PAD.n4160 PAD.n4159 2.2505
R36586 PAD.n4158 PAD.n4055 2.2505
R36587 PAD.n4157 PAD.n4156 2.2505
R36588 PAD.n4152 PAD.n4056 2.2505
R36589 PAD.n4148 PAD.n4147 2.2505
R36590 PAD.n4146 PAD.n4057 2.2505
R36591 PAD.n4145 PAD.n4144 2.2505
R36592 PAD.n4140 PAD.n4058 2.2505
R36593 PAD.n4136 PAD.n4135 2.2505
R36594 PAD.n4134 PAD.n4059 2.2505
R36595 PAD.n4133 PAD.n4132 2.2505
R36596 PAD.n4128 PAD.n4060 2.2505
R36597 PAD.n4124 PAD.n4123 2.2505
R36598 PAD.n4122 PAD.n4061 2.2505
R36599 PAD.n4121 PAD.n4120 2.2505
R36600 PAD.n4116 PAD.n4062 2.2505
R36601 PAD.n4112 PAD.n4111 2.2505
R36602 PAD.n4110 PAD.n4063 2.2505
R36603 PAD.n4109 PAD.n4108 2.2505
R36604 PAD.n4104 PAD.n4064 2.2505
R36605 PAD.n4100 PAD.n4099 2.2505
R36606 PAD.n4098 PAD.n4065 2.2505
R36607 PAD.n4097 PAD.n4096 2.2505
R36608 PAD.n4092 PAD.n4066 2.2505
R36609 PAD.n4088 PAD.n4087 2.2505
R36610 PAD.n4086 PAD.n4067 2.2505
R36611 PAD.n4085 PAD.n4084 2.2505
R36612 PAD.n4080 PAD.n4068 2.2505
R36613 PAD.n4076 PAD.n4075 2.2505
R36614 PAD.n4074 PAD.n4071 2.2505
R36615 PAD.n4073 PAD.n4072 2.2505
R36616 PAD.n4420 PAD.n4419 2.2505
R36617 PAD.n4422 PAD.n4418 2.2505
R36618 PAD.n4427 PAD.n4426 2.2505
R36619 PAD.n4424 PAD.n4416 2.2505
R36620 PAD.n4432 PAD.n4431 2.2505
R36621 PAD.n4434 PAD.n4414 2.2505
R36622 PAD.n4439 PAD.n4438 2.2505
R36623 PAD.n4436 PAD.n4412 2.2505
R36624 PAD.n4444 PAD.n4443 2.2505
R36625 PAD.n4446 PAD.n4410 2.2505
R36626 PAD.n4451 PAD.n4450 2.2505
R36627 PAD.n4448 PAD.n4408 2.2505
R36628 PAD.n4456 PAD.n4455 2.2505
R36629 PAD.n4458 PAD.n4406 2.2505
R36630 PAD.n4463 PAD.n4462 2.2505
R36631 PAD.n4460 PAD.n4404 2.2505
R36632 PAD.n4468 PAD.n4467 2.2505
R36633 PAD.n4470 PAD.n4402 2.2505
R36634 PAD.n4475 PAD.n4474 2.2505
R36635 PAD.n4472 PAD.n4400 2.2505
R36636 PAD.n4480 PAD.n4479 2.2505
R36637 PAD.n4482 PAD.n4398 2.2505
R36638 PAD.n4487 PAD.n4486 2.2505
R36639 PAD.n4484 PAD.n4396 2.2505
R36640 PAD.n4492 PAD.n4491 2.2505
R36641 PAD.n4494 PAD.n4394 2.2505
R36642 PAD.n4499 PAD.n4498 2.2505
R36643 PAD.n4496 PAD.n4392 2.2505
R36644 PAD.n4504 PAD.n4503 2.2505
R36645 PAD.n4506 PAD.n4390 2.2505
R36646 PAD.n4511 PAD.n4510 2.2505
R36647 PAD.n4508 PAD.n4388 2.2505
R36648 PAD.n4516 PAD.n4515 2.2505
R36649 PAD.n4518 PAD.n4386 2.2505
R36650 PAD.n4523 PAD.n4522 2.2505
R36651 PAD.n4520 PAD.n4384 2.2505
R36652 PAD.n4528 PAD.n4527 2.2505
R36653 PAD.n4530 PAD.n4382 2.2505
R36654 PAD.n4535 PAD.n4534 2.2505
R36655 PAD.n4532 PAD.n4380 2.2505
R36656 PAD.n4540 PAD.n4539 2.2505
R36657 PAD.n4542 PAD.n4378 2.2505
R36658 PAD.n4547 PAD.n4546 2.2505
R36659 PAD.n4544 PAD.n4376 2.2505
R36660 PAD.n4552 PAD.n4551 2.2505
R36661 PAD.n4554 PAD.n4374 2.2505
R36662 PAD.n4559 PAD.n4558 2.2505
R36663 PAD.n4556 PAD.n4372 2.2505
R36664 PAD.n4564 PAD.n4563 2.2505
R36665 PAD.n4566 PAD.n4370 2.2505
R36666 PAD.n4571 PAD.n4570 2.2505
R36667 PAD.n4568 PAD.n4368 2.2505
R36668 PAD.n4576 PAD.n4575 2.2505
R36669 PAD.n4578 PAD.n4366 2.2505
R36670 PAD.n4583 PAD.n4582 2.2505
R36671 PAD.n4580 PAD.n4364 2.2505
R36672 PAD.n4588 PAD.n4587 2.2505
R36673 PAD.n4590 PAD.n4362 2.2505
R36674 PAD.n4595 PAD.n4594 2.2505
R36675 PAD.n4592 PAD.n4360 2.2505
R36676 PAD.n4600 PAD.n4599 2.2505
R36677 PAD.n4602 PAD.n4358 2.2505
R36678 PAD.n4607 PAD.n4606 2.2505
R36679 PAD.n4604 PAD.n4356 2.2505
R36680 PAD.n4612 PAD.n4611 2.2505
R36681 PAD.n4614 PAD.n4354 2.2505
R36682 PAD.n4619 PAD.n4618 2.2505
R36683 PAD.n4616 PAD.n4352 2.2505
R36684 PAD.n4624 PAD.n4623 2.2505
R36685 PAD.n4626 PAD.n4350 2.2505
R36686 PAD.n4631 PAD.n4630 2.2505
R36687 PAD.n4628 PAD.n4348 2.2505
R36688 PAD.n4636 PAD.n4635 2.2505
R36689 PAD.n4638 PAD.n4346 2.2505
R36690 PAD.n4643 PAD.n4642 2.2505
R36691 PAD.n4640 PAD.n4344 2.2505
R36692 PAD.n4648 PAD.n4647 2.2505
R36693 PAD.n4650 PAD.n4342 2.2505
R36694 PAD.n4655 PAD.n4654 2.2505
R36695 PAD.n4652 PAD.n4340 2.2505
R36696 PAD.n4661 PAD.n4660 2.2505
R36697 PAD.n4663 PAD.n4338 2.2505
R36698 PAD.n4665 PAD.n4337 2.2505
R36699 PAD.n4668 PAD.n4667 2.2505
R36700 PAD.n4669 PAD.n4668 2.2505
R36701 PAD.n4337 PAD.n4336 2.2505
R36702 PAD.n4658 PAD.n4338 2.2505
R36703 PAD.n4660 PAD.n4659 2.2505
R36704 PAD.n4657 PAD.n4340 2.2505
R36705 PAD.n4656 PAD.n4655 2.2505
R36706 PAD.n4342 PAD.n4341 2.2505
R36707 PAD.n4647 PAD.n4646 2.2505
R36708 PAD.n4645 PAD.n4344 2.2505
R36709 PAD.n4644 PAD.n4643 2.2505
R36710 PAD.n4346 PAD.n4345 2.2505
R36711 PAD.n4635 PAD.n4634 2.2505
R36712 PAD.n4633 PAD.n4348 2.2505
R36713 PAD.n4632 PAD.n4631 2.2505
R36714 PAD.n4350 PAD.n4349 2.2505
R36715 PAD.n4623 PAD.n4622 2.2505
R36716 PAD.n4621 PAD.n4352 2.2505
R36717 PAD.n4620 PAD.n4619 2.2505
R36718 PAD.n4354 PAD.n4353 2.2505
R36719 PAD.n4611 PAD.n4610 2.2505
R36720 PAD.n4609 PAD.n4356 2.2505
R36721 PAD.n4608 PAD.n4607 2.2505
R36722 PAD.n4358 PAD.n4357 2.2505
R36723 PAD.n4599 PAD.n4598 2.2505
R36724 PAD.n4597 PAD.n4360 2.2505
R36725 PAD.n4596 PAD.n4595 2.2505
R36726 PAD.n4362 PAD.n4361 2.2505
R36727 PAD.n4587 PAD.n4586 2.2505
R36728 PAD.n4585 PAD.n4364 2.2505
R36729 PAD.n4584 PAD.n4583 2.2505
R36730 PAD.n4366 PAD.n4365 2.2505
R36731 PAD.n4575 PAD.n4574 2.2505
R36732 PAD.n4573 PAD.n4368 2.2505
R36733 PAD.n4572 PAD.n4571 2.2505
R36734 PAD.n4370 PAD.n4369 2.2505
R36735 PAD.n4563 PAD.n4562 2.2505
R36736 PAD.n4561 PAD.n4372 2.2505
R36737 PAD.n4560 PAD.n4559 2.2505
R36738 PAD.n4374 PAD.n4373 2.2505
R36739 PAD.n4551 PAD.n4550 2.2505
R36740 PAD.n4549 PAD.n4376 2.2505
R36741 PAD.n4548 PAD.n4547 2.2505
R36742 PAD.n4378 PAD.n4377 2.2505
R36743 PAD.n4539 PAD.n4538 2.2505
R36744 PAD.n4537 PAD.n4380 2.2505
R36745 PAD.n4536 PAD.n4535 2.2505
R36746 PAD.n4382 PAD.n4381 2.2505
R36747 PAD.n4527 PAD.n4526 2.2505
R36748 PAD.n4525 PAD.n4384 2.2505
R36749 PAD.n4524 PAD.n4523 2.2505
R36750 PAD.n4386 PAD.n4385 2.2505
R36751 PAD.n4515 PAD.n4514 2.2505
R36752 PAD.n4513 PAD.n4388 2.2505
R36753 PAD.n4512 PAD.n4511 2.2505
R36754 PAD.n4390 PAD.n4389 2.2505
R36755 PAD.n4503 PAD.n4502 2.2505
R36756 PAD.n4501 PAD.n4392 2.2505
R36757 PAD.n4500 PAD.n4499 2.2505
R36758 PAD.n4394 PAD.n4393 2.2505
R36759 PAD.n4491 PAD.n4490 2.2505
R36760 PAD.n4489 PAD.n4396 2.2505
R36761 PAD.n4488 PAD.n4487 2.2505
R36762 PAD.n4398 PAD.n4397 2.2505
R36763 PAD.n4479 PAD.n4478 2.2505
R36764 PAD.n4477 PAD.n4400 2.2505
R36765 PAD.n4476 PAD.n4475 2.2505
R36766 PAD.n4402 PAD.n4401 2.2505
R36767 PAD.n4467 PAD.n4466 2.2505
R36768 PAD.n4465 PAD.n4404 2.2505
R36769 PAD.n4464 PAD.n4463 2.2505
R36770 PAD.n4406 PAD.n4405 2.2505
R36771 PAD.n4455 PAD.n4454 2.2505
R36772 PAD.n4453 PAD.n4408 2.2505
R36773 PAD.n4452 PAD.n4451 2.2505
R36774 PAD.n4410 PAD.n4409 2.2505
R36775 PAD.n4443 PAD.n4442 2.2505
R36776 PAD.n4441 PAD.n4412 2.2505
R36777 PAD.n4440 PAD.n4439 2.2505
R36778 PAD.n4414 PAD.n4413 2.2505
R36779 PAD.n4431 PAD.n4430 2.2505
R36780 PAD.n4429 PAD.n4416 2.2505
R36781 PAD.n4428 PAD.n4427 2.2505
R36782 PAD.n4418 PAD.n4417 2.2505
R36783 PAD.n4419 PAD.n4325 2.2505
R36784 PAD.n8395 PAD.n8394 2.2505
R36785 PAD.n8393 PAD.n4725 2.2505
R36786 PAD.n4728 PAD.n4727 2.2505
R36787 PAD.n8389 PAD.n8388 2.2505
R36788 PAD.n8386 PAD.n8385 2.2505
R36789 PAD.n8384 PAD.n4733 2.2505
R36790 PAD.n4731 PAD.n4730 2.2505
R36791 PAD.n8380 PAD.n8379 2.2505
R36792 PAD.n8377 PAD.n8376 2.2505
R36793 PAD.n8375 PAD.n4738 2.2505
R36794 PAD.n4736 PAD.n4735 2.2505
R36795 PAD.n8371 PAD.n8370 2.2505
R36796 PAD.n8368 PAD.n8367 2.2505
R36797 PAD.n8366 PAD.n4743 2.2505
R36798 PAD.n4741 PAD.n4740 2.2505
R36799 PAD.n8362 PAD.n8361 2.2505
R36800 PAD.n8359 PAD.n8358 2.2505
R36801 PAD.n8357 PAD.n4748 2.2505
R36802 PAD.n4746 PAD.n4745 2.2505
R36803 PAD.n8353 PAD.n8352 2.2505
R36804 PAD.n8350 PAD.n8349 2.2505
R36805 PAD.n8348 PAD.n4753 2.2505
R36806 PAD.n4751 PAD.n4750 2.2505
R36807 PAD.n8344 PAD.n8343 2.2505
R36808 PAD.n8341 PAD.n8340 2.2505
R36809 PAD.n8339 PAD.n4758 2.2505
R36810 PAD.n4756 PAD.n4755 2.2505
R36811 PAD.n8335 PAD.n8334 2.2505
R36812 PAD.n8332 PAD.n8331 2.2505
R36813 PAD.n8330 PAD.n4763 2.2505
R36814 PAD.n4761 PAD.n4760 2.2505
R36815 PAD.n8326 PAD.n8325 2.2505
R36816 PAD.n8323 PAD.n8322 2.2505
R36817 PAD.n8321 PAD.n4768 2.2505
R36818 PAD.n4766 PAD.n4765 2.2505
R36819 PAD.n8317 PAD.n8316 2.2505
R36820 PAD.n8314 PAD.n8313 2.2505
R36821 PAD.n8312 PAD.n4773 2.2505
R36822 PAD.n4771 PAD.n4770 2.2505
R36823 PAD.n8308 PAD.n8307 2.2505
R36824 PAD.n8305 PAD.n8304 2.2505
R36825 PAD.n8303 PAD.n4778 2.2505
R36826 PAD.n4776 PAD.n4775 2.2505
R36827 PAD.n8299 PAD.n8298 2.2505
R36828 PAD.n8296 PAD.n8295 2.2505
R36829 PAD.n8294 PAD.n4783 2.2505
R36830 PAD.n4781 PAD.n4780 2.2505
R36831 PAD.n8290 PAD.n8289 2.2505
R36832 PAD.n8287 PAD.n8286 2.2505
R36833 PAD.n8285 PAD.n4788 2.2505
R36834 PAD.n4786 PAD.n4785 2.2505
R36835 PAD.n8281 PAD.n8280 2.2505
R36836 PAD.n8278 PAD.n8277 2.2505
R36837 PAD.n8276 PAD.n4793 2.2505
R36838 PAD.n4791 PAD.n4790 2.2505
R36839 PAD.n8272 PAD.n8271 2.2505
R36840 PAD.n8269 PAD.n8268 2.2505
R36841 PAD.n8267 PAD.n4798 2.2505
R36842 PAD.n4796 PAD.n4795 2.2505
R36843 PAD.n8263 PAD.n8262 2.2505
R36844 PAD.n8260 PAD.n8259 2.2505
R36845 PAD.n8258 PAD.n4803 2.2505
R36846 PAD.n4801 PAD.n4800 2.2505
R36847 PAD.n8254 PAD.n8253 2.2505
R36848 PAD.n8251 PAD.n8250 2.2505
R36849 PAD.n8249 PAD.n4808 2.2505
R36850 PAD.n4806 PAD.n4805 2.2505
R36851 PAD.n8245 PAD.n8244 2.2505
R36852 PAD.n8242 PAD.n8241 2.2505
R36853 PAD.n8240 PAD.n4813 2.2505
R36854 PAD.n4811 PAD.n4810 2.2505
R36855 PAD.n8236 PAD.n8235 2.2505
R36856 PAD.n8233 PAD.n8232 2.2505
R36857 PAD.n8231 PAD.n4818 2.2505
R36858 PAD.n4816 PAD.n4815 2.2505
R36859 PAD.n8227 PAD.n8226 2.2505
R36860 PAD.n8224 PAD.n8223 2.2505
R36861 PAD.n8222 PAD.n4823 2.2505
R36862 PAD.n4821 PAD.n4820 2.2505
R36863 PAD.n8218 PAD.n8217 2.2505
R36864 PAD.n8215 PAD.n8214 2.2505
R36865 PAD.n8213 PAD.n4828 2.2505
R36866 PAD.n4826 PAD.n4825 2.2505
R36867 PAD.n4832 PAD.n4829 2.2505
R36868 PAD.n8210 PAD.n4829 2.2505
R36869 PAD.n8211 PAD.n4825 2.2505
R36870 PAD.n8213 PAD.n8212 2.2505
R36871 PAD.n8214 PAD.n4824 2.2505
R36872 PAD.n8219 PAD.n8218 2.2505
R36873 PAD.n8220 PAD.n4820 2.2505
R36874 PAD.n8222 PAD.n8221 2.2505
R36875 PAD.n8223 PAD.n4819 2.2505
R36876 PAD.n8228 PAD.n8227 2.2505
R36877 PAD.n8229 PAD.n4815 2.2505
R36878 PAD.n8231 PAD.n8230 2.2505
R36879 PAD.n8232 PAD.n4814 2.2505
R36880 PAD.n8237 PAD.n8236 2.2505
R36881 PAD.n8238 PAD.n4810 2.2505
R36882 PAD.n8240 PAD.n8239 2.2505
R36883 PAD.n8241 PAD.n4809 2.2505
R36884 PAD.n8246 PAD.n8245 2.2505
R36885 PAD.n8247 PAD.n4805 2.2505
R36886 PAD.n8249 PAD.n8248 2.2505
R36887 PAD.n8250 PAD.n4804 2.2505
R36888 PAD.n8255 PAD.n8254 2.2505
R36889 PAD.n8256 PAD.n4800 2.2505
R36890 PAD.n8258 PAD.n8257 2.2505
R36891 PAD.n8259 PAD.n4799 2.2505
R36892 PAD.n8264 PAD.n8263 2.2505
R36893 PAD.n8265 PAD.n4795 2.2505
R36894 PAD.n8267 PAD.n8266 2.2505
R36895 PAD.n8268 PAD.n4794 2.2505
R36896 PAD.n8273 PAD.n8272 2.2505
R36897 PAD.n8274 PAD.n4790 2.2505
R36898 PAD.n8276 PAD.n8275 2.2505
R36899 PAD.n8277 PAD.n4789 2.2505
R36900 PAD.n8282 PAD.n8281 2.2505
R36901 PAD.n8283 PAD.n4785 2.2505
R36902 PAD.n8285 PAD.n8284 2.2505
R36903 PAD.n8286 PAD.n4784 2.2505
R36904 PAD.n8291 PAD.n8290 2.2505
R36905 PAD.n8292 PAD.n4780 2.2505
R36906 PAD.n8294 PAD.n8293 2.2505
R36907 PAD.n8295 PAD.n4779 2.2505
R36908 PAD.n8300 PAD.n8299 2.2505
R36909 PAD.n8301 PAD.n4775 2.2505
R36910 PAD.n8303 PAD.n8302 2.2505
R36911 PAD.n8304 PAD.n4774 2.2505
R36912 PAD.n8309 PAD.n8308 2.2505
R36913 PAD.n8310 PAD.n4770 2.2505
R36914 PAD.n8312 PAD.n8311 2.2505
R36915 PAD.n8313 PAD.n4769 2.2505
R36916 PAD.n8318 PAD.n8317 2.2505
R36917 PAD.n8319 PAD.n4765 2.2505
R36918 PAD.n8321 PAD.n8320 2.2505
R36919 PAD.n8322 PAD.n4764 2.2505
R36920 PAD.n8327 PAD.n8326 2.2505
R36921 PAD.n8328 PAD.n4760 2.2505
R36922 PAD.n8330 PAD.n8329 2.2505
R36923 PAD.n8331 PAD.n4759 2.2505
R36924 PAD.n8336 PAD.n8335 2.2505
R36925 PAD.n8337 PAD.n4755 2.2505
R36926 PAD.n8339 PAD.n8338 2.2505
R36927 PAD.n8340 PAD.n4754 2.2505
R36928 PAD.n8345 PAD.n8344 2.2505
R36929 PAD.n8346 PAD.n4750 2.2505
R36930 PAD.n8348 PAD.n8347 2.2505
R36931 PAD.n8349 PAD.n4749 2.2505
R36932 PAD.n8354 PAD.n8353 2.2505
R36933 PAD.n8355 PAD.n4745 2.2505
R36934 PAD.n8357 PAD.n8356 2.2505
R36935 PAD.n8358 PAD.n4744 2.2505
R36936 PAD.n8363 PAD.n8362 2.2505
R36937 PAD.n8364 PAD.n4740 2.2505
R36938 PAD.n8366 PAD.n8365 2.2505
R36939 PAD.n8367 PAD.n4739 2.2505
R36940 PAD.n8372 PAD.n8371 2.2505
R36941 PAD.n8373 PAD.n4735 2.2505
R36942 PAD.n8375 PAD.n8374 2.2505
R36943 PAD.n8376 PAD.n4734 2.2505
R36944 PAD.n8381 PAD.n8380 2.2505
R36945 PAD.n8382 PAD.n4730 2.2505
R36946 PAD.n8384 PAD.n8383 2.2505
R36947 PAD.n8385 PAD.n4729 2.2505
R36948 PAD.n8390 PAD.n8389 2.2505
R36949 PAD.n8391 PAD.n4728 2.2505
R36950 PAD.n8393 PAD.n8392 2.2505
R36951 PAD.n8394 PAD.n4676 2.2505
R36952 PAD.n5178 PAD.n4847 2.2505
R36953 PAD.n5177 PAD.n5176 2.2505
R36954 PAD.n5174 PAD.n4848 2.2505
R36955 PAD.n5172 PAD.n5171 2.2505
R36956 PAD.n5164 PAD.n4851 2.2505
R36957 PAD.n5167 PAD.n5166 2.2505
R36958 PAD.n5162 PAD.n4854 2.2505
R36959 PAD.n5160 PAD.n5159 2.2505
R36960 PAD.n5152 PAD.n4856 2.2505
R36961 PAD.n5155 PAD.n5154 2.2505
R36962 PAD.n5150 PAD.n4858 2.2505
R36963 PAD.n5148 PAD.n5147 2.2505
R36964 PAD.n5140 PAD.n4860 2.2505
R36965 PAD.n5143 PAD.n5142 2.2505
R36966 PAD.n5138 PAD.n4862 2.2505
R36967 PAD.n5136 PAD.n5135 2.2505
R36968 PAD.n5128 PAD.n4864 2.2505
R36969 PAD.n5131 PAD.n5130 2.2505
R36970 PAD.n5126 PAD.n4866 2.2505
R36971 PAD.n5124 PAD.n5123 2.2505
R36972 PAD.n5116 PAD.n4868 2.2505
R36973 PAD.n5119 PAD.n5118 2.2505
R36974 PAD.n5114 PAD.n4870 2.2505
R36975 PAD.n5112 PAD.n5111 2.2505
R36976 PAD.n5104 PAD.n4872 2.2505
R36977 PAD.n5107 PAD.n5106 2.2505
R36978 PAD.n5102 PAD.n4874 2.2505
R36979 PAD.n5100 PAD.n5099 2.2505
R36980 PAD.n5092 PAD.n4876 2.2505
R36981 PAD.n5095 PAD.n5094 2.2505
R36982 PAD.n5090 PAD.n4878 2.2505
R36983 PAD.n5088 PAD.n5087 2.2505
R36984 PAD.n5080 PAD.n4880 2.2505
R36985 PAD.n5083 PAD.n5082 2.2505
R36986 PAD.n5078 PAD.n4882 2.2505
R36987 PAD.n5076 PAD.n5075 2.2505
R36988 PAD.n5068 PAD.n4884 2.2505
R36989 PAD.n5071 PAD.n5070 2.2505
R36990 PAD.n5066 PAD.n4886 2.2505
R36991 PAD.n5064 PAD.n5063 2.2505
R36992 PAD.n5056 PAD.n4888 2.2505
R36993 PAD.n5059 PAD.n5058 2.2505
R36994 PAD.n5054 PAD.n4890 2.2505
R36995 PAD.n5052 PAD.n5051 2.2505
R36996 PAD.n5044 PAD.n4892 2.2505
R36997 PAD.n5047 PAD.n5046 2.2505
R36998 PAD.n5042 PAD.n4894 2.2505
R36999 PAD.n5040 PAD.n5039 2.2505
R37000 PAD.n5032 PAD.n4896 2.2505
R37001 PAD.n5035 PAD.n5034 2.2505
R37002 PAD.n5030 PAD.n4898 2.2505
R37003 PAD.n5028 PAD.n5027 2.2505
R37004 PAD.n5020 PAD.n4900 2.2505
R37005 PAD.n5023 PAD.n5022 2.2505
R37006 PAD.n5018 PAD.n4902 2.2505
R37007 PAD.n5016 PAD.n5015 2.2505
R37008 PAD.n5008 PAD.n4904 2.2505
R37009 PAD.n5011 PAD.n5010 2.2505
R37010 PAD.n5006 PAD.n4906 2.2505
R37011 PAD.n5004 PAD.n5003 2.2505
R37012 PAD.n4996 PAD.n4908 2.2505
R37013 PAD.n4999 PAD.n4998 2.2505
R37014 PAD.n4994 PAD.n4910 2.2505
R37015 PAD.n4992 PAD.n4991 2.2505
R37016 PAD.n4984 PAD.n4912 2.2505
R37017 PAD.n4987 PAD.n4986 2.2505
R37018 PAD.n4982 PAD.n4914 2.2505
R37019 PAD.n4980 PAD.n4979 2.2505
R37020 PAD.n4972 PAD.n4916 2.2505
R37021 PAD.n4975 PAD.n4974 2.2505
R37022 PAD.n4970 PAD.n4918 2.2505
R37023 PAD.n4968 PAD.n4967 2.2505
R37024 PAD.n4960 PAD.n4920 2.2505
R37025 PAD.n4963 PAD.n4962 2.2505
R37026 PAD.n4958 PAD.n4922 2.2505
R37027 PAD.n4956 PAD.n4955 2.2505
R37028 PAD.n4948 PAD.n4924 2.2505
R37029 PAD.n4951 PAD.n4950 2.2505
R37030 PAD.n4946 PAD.n4926 2.2505
R37031 PAD.n4944 PAD.n4943 2.2505
R37032 PAD.n4936 PAD.n4928 2.2505
R37033 PAD.n4939 PAD.n4938 2.2505
R37034 PAD.n4934 PAD.n4930 2.2505
R37035 PAD.n4932 PAD.n4931 2.2505
R37036 PAD.n4931 PAD.n4835 2.2505
R37037 PAD.n4930 PAD.n4929 2.2505
R37038 PAD.n4940 PAD.n4939 2.2505
R37039 PAD.n4941 PAD.n4928 2.2505
R37040 PAD.n4943 PAD.n4942 2.2505
R37041 PAD.n4926 PAD.n4925 2.2505
R37042 PAD.n4952 PAD.n4951 2.2505
R37043 PAD.n4953 PAD.n4924 2.2505
R37044 PAD.n4955 PAD.n4954 2.2505
R37045 PAD.n4922 PAD.n4921 2.2505
R37046 PAD.n4964 PAD.n4963 2.2505
R37047 PAD.n4965 PAD.n4920 2.2505
R37048 PAD.n4967 PAD.n4966 2.2505
R37049 PAD.n4918 PAD.n4917 2.2505
R37050 PAD.n4976 PAD.n4975 2.2505
R37051 PAD.n4977 PAD.n4916 2.2505
R37052 PAD.n4979 PAD.n4978 2.2505
R37053 PAD.n4914 PAD.n4913 2.2505
R37054 PAD.n4988 PAD.n4987 2.2505
R37055 PAD.n4989 PAD.n4912 2.2505
R37056 PAD.n4991 PAD.n4990 2.2505
R37057 PAD.n4910 PAD.n4909 2.2505
R37058 PAD.n5000 PAD.n4999 2.2505
R37059 PAD.n5001 PAD.n4908 2.2505
R37060 PAD.n5003 PAD.n5002 2.2505
R37061 PAD.n4906 PAD.n4905 2.2505
R37062 PAD.n5012 PAD.n5011 2.2505
R37063 PAD.n5013 PAD.n4904 2.2505
R37064 PAD.n5015 PAD.n5014 2.2505
R37065 PAD.n4902 PAD.n4901 2.2505
R37066 PAD.n5024 PAD.n5023 2.2505
R37067 PAD.n5025 PAD.n4900 2.2505
R37068 PAD.n5027 PAD.n5026 2.2505
R37069 PAD.n4898 PAD.n4897 2.2505
R37070 PAD.n5036 PAD.n5035 2.2505
R37071 PAD.n5037 PAD.n4896 2.2505
R37072 PAD.n5039 PAD.n5038 2.2505
R37073 PAD.n4894 PAD.n4893 2.2505
R37074 PAD.n5048 PAD.n5047 2.2505
R37075 PAD.n5049 PAD.n4892 2.2505
R37076 PAD.n5051 PAD.n5050 2.2505
R37077 PAD.n4890 PAD.n4889 2.2505
R37078 PAD.n5060 PAD.n5059 2.2505
R37079 PAD.n5061 PAD.n4888 2.2505
R37080 PAD.n5063 PAD.n5062 2.2505
R37081 PAD.n4886 PAD.n4885 2.2505
R37082 PAD.n5072 PAD.n5071 2.2505
R37083 PAD.n5073 PAD.n4884 2.2505
R37084 PAD.n5075 PAD.n5074 2.2505
R37085 PAD.n4882 PAD.n4881 2.2505
R37086 PAD.n5084 PAD.n5083 2.2505
R37087 PAD.n5085 PAD.n4880 2.2505
R37088 PAD.n5087 PAD.n5086 2.2505
R37089 PAD.n4878 PAD.n4877 2.2505
R37090 PAD.n5096 PAD.n5095 2.2505
R37091 PAD.n5097 PAD.n4876 2.2505
R37092 PAD.n5099 PAD.n5098 2.2505
R37093 PAD.n4874 PAD.n4873 2.2505
R37094 PAD.n5108 PAD.n5107 2.2505
R37095 PAD.n5109 PAD.n4872 2.2505
R37096 PAD.n5111 PAD.n5110 2.2505
R37097 PAD.n4870 PAD.n4869 2.2505
R37098 PAD.n5120 PAD.n5119 2.2505
R37099 PAD.n5121 PAD.n4868 2.2505
R37100 PAD.n5123 PAD.n5122 2.2505
R37101 PAD.n4866 PAD.n4865 2.2505
R37102 PAD.n5132 PAD.n5131 2.2505
R37103 PAD.n5133 PAD.n4864 2.2505
R37104 PAD.n5135 PAD.n5134 2.2505
R37105 PAD.n4862 PAD.n4861 2.2505
R37106 PAD.n5144 PAD.n5143 2.2505
R37107 PAD.n5145 PAD.n4860 2.2505
R37108 PAD.n5147 PAD.n5146 2.2505
R37109 PAD.n4858 PAD.n4857 2.2505
R37110 PAD.n5156 PAD.n5155 2.2505
R37111 PAD.n5157 PAD.n4856 2.2505
R37112 PAD.n5159 PAD.n5158 2.2505
R37113 PAD.n4854 PAD.n4853 2.2505
R37114 PAD.n5168 PAD.n5167 2.2505
R37115 PAD.n5169 PAD.n4851 2.2505
R37116 PAD.n5171 PAD.n5170 2.2505
R37117 PAD.n4852 PAD.n4848 2.2505
R37118 PAD.n5177 PAD.n4846 2.2505
R37119 PAD.n5179 PAD.n5178 2.2505
R37120 PAD.n8161 PAD.n8160 2.2505
R37121 PAD.n8159 PAD.n7871 2.2505
R37122 PAD.n7874 PAD.n7873 2.2505
R37123 PAD.n8155 PAD.n8154 2.2505
R37124 PAD.n8152 PAD.n8151 2.2505
R37125 PAD.n8150 PAD.n7879 2.2505
R37126 PAD.n7877 PAD.n7876 2.2505
R37127 PAD.n8146 PAD.n8145 2.2505
R37128 PAD.n8143 PAD.n8142 2.2505
R37129 PAD.n8141 PAD.n7884 2.2505
R37130 PAD.n7882 PAD.n7881 2.2505
R37131 PAD.n8137 PAD.n8136 2.2505
R37132 PAD.n8134 PAD.n8133 2.2505
R37133 PAD.n8132 PAD.n7889 2.2505
R37134 PAD.n7887 PAD.n7886 2.2505
R37135 PAD.n8128 PAD.n8127 2.2505
R37136 PAD.n8125 PAD.n8124 2.2505
R37137 PAD.n8123 PAD.n7894 2.2505
R37138 PAD.n7892 PAD.n7891 2.2505
R37139 PAD.n8119 PAD.n8118 2.2505
R37140 PAD.n8116 PAD.n8115 2.2505
R37141 PAD.n8114 PAD.n7899 2.2505
R37142 PAD.n7897 PAD.n7896 2.2505
R37143 PAD.n8110 PAD.n8109 2.2505
R37144 PAD.n8107 PAD.n8106 2.2505
R37145 PAD.n8105 PAD.n7904 2.2505
R37146 PAD.n7902 PAD.n7901 2.2505
R37147 PAD.n8101 PAD.n8100 2.2505
R37148 PAD.n8098 PAD.n8097 2.2505
R37149 PAD.n8096 PAD.n7909 2.2505
R37150 PAD.n7907 PAD.n7906 2.2505
R37151 PAD.n8092 PAD.n8091 2.2505
R37152 PAD.n8089 PAD.n8088 2.2505
R37153 PAD.n8087 PAD.n7914 2.2505
R37154 PAD.n7912 PAD.n7911 2.2505
R37155 PAD.n8083 PAD.n8082 2.2505
R37156 PAD.n8080 PAD.n8079 2.2505
R37157 PAD.n8078 PAD.n7919 2.2505
R37158 PAD.n7917 PAD.n7916 2.2505
R37159 PAD.n8074 PAD.n8073 2.2505
R37160 PAD.n8071 PAD.n8070 2.2505
R37161 PAD.n8069 PAD.n7924 2.2505
R37162 PAD.n7922 PAD.n7921 2.2505
R37163 PAD.n8065 PAD.n8064 2.2505
R37164 PAD.n8062 PAD.n8061 2.2505
R37165 PAD.n8060 PAD.n7929 2.2505
R37166 PAD.n7927 PAD.n7926 2.2505
R37167 PAD.n8056 PAD.n8055 2.2505
R37168 PAD.n8053 PAD.n8052 2.2505
R37169 PAD.n8051 PAD.n7934 2.2505
R37170 PAD.n7932 PAD.n7931 2.2505
R37171 PAD.n8047 PAD.n8046 2.2505
R37172 PAD.n8044 PAD.n8043 2.2505
R37173 PAD.n8042 PAD.n7939 2.2505
R37174 PAD.n7937 PAD.n7936 2.2505
R37175 PAD.n8038 PAD.n8037 2.2505
R37176 PAD.n8035 PAD.n8034 2.2505
R37177 PAD.n8033 PAD.n7944 2.2505
R37178 PAD.n7942 PAD.n7941 2.2505
R37179 PAD.n8029 PAD.n8028 2.2505
R37180 PAD.n8026 PAD.n8025 2.2505
R37181 PAD.n8024 PAD.n7949 2.2505
R37182 PAD.n7947 PAD.n7946 2.2505
R37183 PAD.n8020 PAD.n8019 2.2505
R37184 PAD.n8017 PAD.n8016 2.2505
R37185 PAD.n8015 PAD.n7954 2.2505
R37186 PAD.n7952 PAD.n7951 2.2505
R37187 PAD.n8011 PAD.n8010 2.2505
R37188 PAD.n8008 PAD.n8007 2.2505
R37189 PAD.n8006 PAD.n7959 2.2505
R37190 PAD.n7957 PAD.n7956 2.2505
R37191 PAD.n8002 PAD.n8001 2.2505
R37192 PAD.n7999 PAD.n7998 2.2505
R37193 PAD.n7997 PAD.n7964 2.2505
R37194 PAD.n7962 PAD.n7961 2.2505
R37195 PAD.n7993 PAD.n7992 2.2505
R37196 PAD.n7990 PAD.n7989 2.2505
R37197 PAD.n7988 PAD.n7969 2.2505
R37198 PAD.n7967 PAD.n7966 2.2505
R37199 PAD.n7984 PAD.n7983 2.2505
R37200 PAD.n7981 PAD.n7980 2.2505
R37201 PAD.n7979 PAD.n7976 2.2505
R37202 PAD.n7974 PAD.n7973 2.2505
R37203 PAD.n7972 PAD.n7971 2.2505
R37204 PAD.n7972 PAD.n5186 2.2505
R37205 PAD.n7977 PAD.n7973 2.2505
R37206 PAD.n7979 PAD.n7978 2.2505
R37207 PAD.n7980 PAD.n7970 2.2505
R37208 PAD.n7985 PAD.n7984 2.2505
R37209 PAD.n7986 PAD.n7966 2.2505
R37210 PAD.n7988 PAD.n7987 2.2505
R37211 PAD.n7989 PAD.n7965 2.2505
R37212 PAD.n7994 PAD.n7993 2.2505
R37213 PAD.n7995 PAD.n7961 2.2505
R37214 PAD.n7997 PAD.n7996 2.2505
R37215 PAD.n7998 PAD.n7960 2.2505
R37216 PAD.n8003 PAD.n8002 2.2505
R37217 PAD.n8004 PAD.n7956 2.2505
R37218 PAD.n8006 PAD.n8005 2.2505
R37219 PAD.n8007 PAD.n7955 2.2505
R37220 PAD.n8012 PAD.n8011 2.2505
R37221 PAD.n8013 PAD.n7951 2.2505
R37222 PAD.n8015 PAD.n8014 2.2505
R37223 PAD.n8016 PAD.n7950 2.2505
R37224 PAD.n8021 PAD.n8020 2.2505
R37225 PAD.n8022 PAD.n7946 2.2505
R37226 PAD.n8024 PAD.n8023 2.2505
R37227 PAD.n8025 PAD.n7945 2.2505
R37228 PAD.n8030 PAD.n8029 2.2505
R37229 PAD.n8031 PAD.n7941 2.2505
R37230 PAD.n8033 PAD.n8032 2.2505
R37231 PAD.n8034 PAD.n7940 2.2505
R37232 PAD.n8039 PAD.n8038 2.2505
R37233 PAD.n8040 PAD.n7936 2.2505
R37234 PAD.n8042 PAD.n8041 2.2505
R37235 PAD.n8043 PAD.n7935 2.2505
R37236 PAD.n8048 PAD.n8047 2.2505
R37237 PAD.n8049 PAD.n7931 2.2505
R37238 PAD.n8051 PAD.n8050 2.2505
R37239 PAD.n8052 PAD.n7930 2.2505
R37240 PAD.n8057 PAD.n8056 2.2505
R37241 PAD.n8058 PAD.n7926 2.2505
R37242 PAD.n8060 PAD.n8059 2.2505
R37243 PAD.n8061 PAD.n7925 2.2505
R37244 PAD.n8066 PAD.n8065 2.2505
R37245 PAD.n8067 PAD.n7921 2.2505
R37246 PAD.n8069 PAD.n8068 2.2505
R37247 PAD.n8070 PAD.n7920 2.2505
R37248 PAD.n8075 PAD.n8074 2.2505
R37249 PAD.n8076 PAD.n7916 2.2505
R37250 PAD.n8078 PAD.n8077 2.2505
R37251 PAD.n8079 PAD.n7915 2.2505
R37252 PAD.n8084 PAD.n8083 2.2505
R37253 PAD.n8085 PAD.n7911 2.2505
R37254 PAD.n8087 PAD.n8086 2.2505
R37255 PAD.n8088 PAD.n7910 2.2505
R37256 PAD.n8093 PAD.n8092 2.2505
R37257 PAD.n8094 PAD.n7906 2.2505
R37258 PAD.n8096 PAD.n8095 2.2505
R37259 PAD.n8097 PAD.n7905 2.2505
R37260 PAD.n8102 PAD.n8101 2.2505
R37261 PAD.n8103 PAD.n7901 2.2505
R37262 PAD.n8105 PAD.n8104 2.2505
R37263 PAD.n8106 PAD.n7900 2.2505
R37264 PAD.n8111 PAD.n8110 2.2505
R37265 PAD.n8112 PAD.n7896 2.2505
R37266 PAD.n8114 PAD.n8113 2.2505
R37267 PAD.n8115 PAD.n7895 2.2505
R37268 PAD.n8120 PAD.n8119 2.2505
R37269 PAD.n8121 PAD.n7891 2.2505
R37270 PAD.n8123 PAD.n8122 2.2505
R37271 PAD.n8124 PAD.n7890 2.2505
R37272 PAD.n8129 PAD.n8128 2.2505
R37273 PAD.n8130 PAD.n7886 2.2505
R37274 PAD.n8132 PAD.n8131 2.2505
R37275 PAD.n8133 PAD.n7885 2.2505
R37276 PAD.n8138 PAD.n8137 2.2505
R37277 PAD.n8139 PAD.n7881 2.2505
R37278 PAD.n8141 PAD.n8140 2.2505
R37279 PAD.n8142 PAD.n7880 2.2505
R37280 PAD.n8147 PAD.n8146 2.2505
R37281 PAD.n8148 PAD.n7876 2.2505
R37282 PAD.n8150 PAD.n8149 2.2505
R37283 PAD.n8151 PAD.n7875 2.2505
R37284 PAD.n8156 PAD.n8155 2.2505
R37285 PAD.n8157 PAD.n7874 2.2505
R37286 PAD.n8159 PAD.n8158 2.2505
R37287 PAD.n8160 PAD.n5193 2.2505
R37288 PAD.n5542 PAD.n5211 2.2505
R37289 PAD.n5541 PAD.n5540 2.2505
R37290 PAD.n5538 PAD.n5212 2.2505
R37291 PAD.n5536 PAD.n5535 2.2505
R37292 PAD.n5528 PAD.n5215 2.2505
R37293 PAD.n5531 PAD.n5530 2.2505
R37294 PAD.n5526 PAD.n5218 2.2505
R37295 PAD.n5524 PAD.n5523 2.2505
R37296 PAD.n5516 PAD.n5220 2.2505
R37297 PAD.n5519 PAD.n5518 2.2505
R37298 PAD.n5514 PAD.n5222 2.2505
R37299 PAD.n5512 PAD.n5511 2.2505
R37300 PAD.n5504 PAD.n5224 2.2505
R37301 PAD.n5507 PAD.n5506 2.2505
R37302 PAD.n5502 PAD.n5226 2.2505
R37303 PAD.n5500 PAD.n5499 2.2505
R37304 PAD.n5492 PAD.n5228 2.2505
R37305 PAD.n5495 PAD.n5494 2.2505
R37306 PAD.n5490 PAD.n5230 2.2505
R37307 PAD.n5488 PAD.n5487 2.2505
R37308 PAD.n5480 PAD.n5232 2.2505
R37309 PAD.n5483 PAD.n5482 2.2505
R37310 PAD.n5478 PAD.n5234 2.2505
R37311 PAD.n5476 PAD.n5475 2.2505
R37312 PAD.n5468 PAD.n5236 2.2505
R37313 PAD.n5471 PAD.n5470 2.2505
R37314 PAD.n5466 PAD.n5238 2.2505
R37315 PAD.n5464 PAD.n5463 2.2505
R37316 PAD.n5456 PAD.n5240 2.2505
R37317 PAD.n5459 PAD.n5458 2.2505
R37318 PAD.n5454 PAD.n5242 2.2505
R37319 PAD.n5452 PAD.n5451 2.2505
R37320 PAD.n5444 PAD.n5244 2.2505
R37321 PAD.n5447 PAD.n5446 2.2505
R37322 PAD.n5442 PAD.n5246 2.2505
R37323 PAD.n5440 PAD.n5439 2.2505
R37324 PAD.n5432 PAD.n5248 2.2505
R37325 PAD.n5435 PAD.n5434 2.2505
R37326 PAD.n5430 PAD.n5250 2.2505
R37327 PAD.n5428 PAD.n5427 2.2505
R37328 PAD.n5420 PAD.n5252 2.2505
R37329 PAD.n5423 PAD.n5422 2.2505
R37330 PAD.n5418 PAD.n5254 2.2505
R37331 PAD.n5416 PAD.n5415 2.2505
R37332 PAD.n5408 PAD.n5256 2.2505
R37333 PAD.n5411 PAD.n5410 2.2505
R37334 PAD.n5406 PAD.n5258 2.2505
R37335 PAD.n5404 PAD.n5403 2.2505
R37336 PAD.n5396 PAD.n5260 2.2505
R37337 PAD.n5399 PAD.n5398 2.2505
R37338 PAD.n5394 PAD.n5262 2.2505
R37339 PAD.n5392 PAD.n5391 2.2505
R37340 PAD.n5384 PAD.n5264 2.2505
R37341 PAD.n5387 PAD.n5386 2.2505
R37342 PAD.n5382 PAD.n5266 2.2505
R37343 PAD.n5380 PAD.n5379 2.2505
R37344 PAD.n5372 PAD.n5268 2.2505
R37345 PAD.n5375 PAD.n5374 2.2505
R37346 PAD.n5370 PAD.n5270 2.2505
R37347 PAD.n5368 PAD.n5367 2.2505
R37348 PAD.n5360 PAD.n5272 2.2505
R37349 PAD.n5363 PAD.n5362 2.2505
R37350 PAD.n5358 PAD.n5274 2.2505
R37351 PAD.n5356 PAD.n5355 2.2505
R37352 PAD.n5348 PAD.n5276 2.2505
R37353 PAD.n5351 PAD.n5350 2.2505
R37354 PAD.n5346 PAD.n5278 2.2505
R37355 PAD.n5344 PAD.n5343 2.2505
R37356 PAD.n5336 PAD.n5280 2.2505
R37357 PAD.n5339 PAD.n5338 2.2505
R37358 PAD.n5334 PAD.n5282 2.2505
R37359 PAD.n5332 PAD.n5331 2.2505
R37360 PAD.n5324 PAD.n5284 2.2505
R37361 PAD.n5327 PAD.n5326 2.2505
R37362 PAD.n5322 PAD.n5286 2.2505
R37363 PAD.n5320 PAD.n5319 2.2505
R37364 PAD.n5312 PAD.n5288 2.2505
R37365 PAD.n5315 PAD.n5314 2.2505
R37366 PAD.n5310 PAD.n5290 2.2505
R37367 PAD.n5308 PAD.n5307 2.2505
R37368 PAD.n5300 PAD.n5292 2.2505
R37369 PAD.n5303 PAD.n5302 2.2505
R37370 PAD.n5298 PAD.n5294 2.2505
R37371 PAD.n5296 PAD.n5295 2.2505
R37372 PAD.n5295 PAD.n5200 2.2505
R37373 PAD.n5294 PAD.n5293 2.2505
R37374 PAD.n5304 PAD.n5303 2.2505
R37375 PAD.n5305 PAD.n5292 2.2505
R37376 PAD.n5307 PAD.n5306 2.2505
R37377 PAD.n5290 PAD.n5289 2.2505
R37378 PAD.n5316 PAD.n5315 2.2505
R37379 PAD.n5317 PAD.n5288 2.2505
R37380 PAD.n5319 PAD.n5318 2.2505
R37381 PAD.n5286 PAD.n5285 2.2505
R37382 PAD.n5328 PAD.n5327 2.2505
R37383 PAD.n5329 PAD.n5284 2.2505
R37384 PAD.n5331 PAD.n5330 2.2505
R37385 PAD.n5282 PAD.n5281 2.2505
R37386 PAD.n5340 PAD.n5339 2.2505
R37387 PAD.n5341 PAD.n5280 2.2505
R37388 PAD.n5343 PAD.n5342 2.2505
R37389 PAD.n5278 PAD.n5277 2.2505
R37390 PAD.n5352 PAD.n5351 2.2505
R37391 PAD.n5353 PAD.n5276 2.2505
R37392 PAD.n5355 PAD.n5354 2.2505
R37393 PAD.n5274 PAD.n5273 2.2505
R37394 PAD.n5364 PAD.n5363 2.2505
R37395 PAD.n5365 PAD.n5272 2.2505
R37396 PAD.n5367 PAD.n5366 2.2505
R37397 PAD.n5270 PAD.n5269 2.2505
R37398 PAD.n5376 PAD.n5375 2.2505
R37399 PAD.n5377 PAD.n5268 2.2505
R37400 PAD.n5379 PAD.n5378 2.2505
R37401 PAD.n5266 PAD.n5265 2.2505
R37402 PAD.n5388 PAD.n5387 2.2505
R37403 PAD.n5389 PAD.n5264 2.2505
R37404 PAD.n5391 PAD.n5390 2.2505
R37405 PAD.n5262 PAD.n5261 2.2505
R37406 PAD.n5400 PAD.n5399 2.2505
R37407 PAD.n5401 PAD.n5260 2.2505
R37408 PAD.n5403 PAD.n5402 2.2505
R37409 PAD.n5258 PAD.n5257 2.2505
R37410 PAD.n5412 PAD.n5411 2.2505
R37411 PAD.n5413 PAD.n5256 2.2505
R37412 PAD.n5415 PAD.n5414 2.2505
R37413 PAD.n5254 PAD.n5253 2.2505
R37414 PAD.n5424 PAD.n5423 2.2505
R37415 PAD.n5425 PAD.n5252 2.2505
R37416 PAD.n5427 PAD.n5426 2.2505
R37417 PAD.n5250 PAD.n5249 2.2505
R37418 PAD.n5436 PAD.n5435 2.2505
R37419 PAD.n5437 PAD.n5248 2.2505
R37420 PAD.n5439 PAD.n5438 2.2505
R37421 PAD.n5246 PAD.n5245 2.2505
R37422 PAD.n5448 PAD.n5447 2.2505
R37423 PAD.n5449 PAD.n5244 2.2505
R37424 PAD.n5451 PAD.n5450 2.2505
R37425 PAD.n5242 PAD.n5241 2.2505
R37426 PAD.n5460 PAD.n5459 2.2505
R37427 PAD.n5461 PAD.n5240 2.2505
R37428 PAD.n5463 PAD.n5462 2.2505
R37429 PAD.n5238 PAD.n5237 2.2505
R37430 PAD.n5472 PAD.n5471 2.2505
R37431 PAD.n5473 PAD.n5236 2.2505
R37432 PAD.n5475 PAD.n5474 2.2505
R37433 PAD.n5234 PAD.n5233 2.2505
R37434 PAD.n5484 PAD.n5483 2.2505
R37435 PAD.n5485 PAD.n5232 2.2505
R37436 PAD.n5487 PAD.n5486 2.2505
R37437 PAD.n5230 PAD.n5229 2.2505
R37438 PAD.n5496 PAD.n5495 2.2505
R37439 PAD.n5497 PAD.n5228 2.2505
R37440 PAD.n5499 PAD.n5498 2.2505
R37441 PAD.n5226 PAD.n5225 2.2505
R37442 PAD.n5508 PAD.n5507 2.2505
R37443 PAD.n5509 PAD.n5224 2.2505
R37444 PAD.n5511 PAD.n5510 2.2505
R37445 PAD.n5222 PAD.n5221 2.2505
R37446 PAD.n5520 PAD.n5519 2.2505
R37447 PAD.n5521 PAD.n5220 2.2505
R37448 PAD.n5523 PAD.n5522 2.2505
R37449 PAD.n5218 PAD.n5217 2.2505
R37450 PAD.n5532 PAD.n5531 2.2505
R37451 PAD.n5533 PAD.n5215 2.2505
R37452 PAD.n5535 PAD.n5534 2.2505
R37453 PAD.n5216 PAD.n5212 2.2505
R37454 PAD.n5541 PAD.n5210 2.2505
R37455 PAD.n5543 PAD.n5542 2.2505
R37456 PAD.n7780 PAD.n7779 2.2505
R37457 PAD.n7106 PAD.n7104 2.2505
R37458 PAD.n7775 PAD.n7774 2.2505
R37459 PAD.n7772 PAD.n7771 2.2505
R37460 PAD.n7769 PAD.n7768 2.2505
R37461 PAD.n7761 PAD.n7108 2.2505
R37462 PAD.n7764 PAD.n7763 2.2505
R37463 PAD.n7760 PAD.n7759 2.2505
R37464 PAD.n7757 PAD.n7756 2.2505
R37465 PAD.n7749 PAD.n7110 2.2505
R37466 PAD.n7752 PAD.n7751 2.2505
R37467 PAD.n7748 PAD.n7747 2.2505
R37468 PAD.n7745 PAD.n7744 2.2505
R37469 PAD.n7737 PAD.n7112 2.2505
R37470 PAD.n7740 PAD.n7739 2.2505
R37471 PAD.n7736 PAD.n7735 2.2505
R37472 PAD.n7733 PAD.n7732 2.2505
R37473 PAD.n7725 PAD.n7114 2.2505
R37474 PAD.n7728 PAD.n7727 2.2505
R37475 PAD.n7724 PAD.n7723 2.2505
R37476 PAD.n7721 PAD.n7720 2.2505
R37477 PAD.n7713 PAD.n7116 2.2505
R37478 PAD.n7716 PAD.n7715 2.2505
R37479 PAD.n7712 PAD.n7711 2.2505
R37480 PAD.n7709 PAD.n7708 2.2505
R37481 PAD.n7701 PAD.n7118 2.2505
R37482 PAD.n7704 PAD.n7703 2.2505
R37483 PAD.n7700 PAD.n7699 2.2505
R37484 PAD.n7697 PAD.n7696 2.2505
R37485 PAD.n7689 PAD.n7120 2.2505
R37486 PAD.n7692 PAD.n7691 2.2505
R37487 PAD.n7688 PAD.n7687 2.2505
R37488 PAD.n7685 PAD.n7684 2.2505
R37489 PAD.n7677 PAD.n7122 2.2505
R37490 PAD.n7680 PAD.n7679 2.2505
R37491 PAD.n7676 PAD.n7675 2.2505
R37492 PAD.n7673 PAD.n7672 2.2505
R37493 PAD.n7665 PAD.n7124 2.2505
R37494 PAD.n7668 PAD.n7667 2.2505
R37495 PAD.n7664 PAD.n7663 2.2505
R37496 PAD.n7661 PAD.n7660 2.2505
R37497 PAD.n7653 PAD.n7126 2.2505
R37498 PAD.n7656 PAD.n7655 2.2505
R37499 PAD.n7652 PAD.n7651 2.2505
R37500 PAD.n7649 PAD.n7648 2.2505
R37501 PAD.n7641 PAD.n7128 2.2505
R37502 PAD.n7644 PAD.n7643 2.2505
R37503 PAD.n7640 PAD.n7639 2.2505
R37504 PAD.n7637 PAD.n7636 2.2505
R37505 PAD.n7629 PAD.n7130 2.2505
R37506 PAD.n7632 PAD.n7631 2.2505
R37507 PAD.n7628 PAD.n7627 2.2505
R37508 PAD.n7625 PAD.n7624 2.2505
R37509 PAD.n7617 PAD.n7132 2.2505
R37510 PAD.n7620 PAD.n7619 2.2505
R37511 PAD.n7616 PAD.n7615 2.2505
R37512 PAD.n7613 PAD.n7612 2.2505
R37513 PAD.n7605 PAD.n7134 2.2505
R37514 PAD.n7608 PAD.n7607 2.2505
R37515 PAD.n7604 PAD.n7603 2.2505
R37516 PAD.n7601 PAD.n7600 2.2505
R37517 PAD.n7593 PAD.n7136 2.2505
R37518 PAD.n7596 PAD.n7595 2.2505
R37519 PAD.n7592 PAD.n7591 2.2505
R37520 PAD.n7589 PAD.n7588 2.2505
R37521 PAD.n7581 PAD.n7138 2.2505
R37522 PAD.n7584 PAD.n7583 2.2505
R37523 PAD.n7580 PAD.n7579 2.2505
R37524 PAD.n7577 PAD.n7576 2.2505
R37525 PAD.n7569 PAD.n7140 2.2505
R37526 PAD.n7572 PAD.n7571 2.2505
R37527 PAD.n7568 PAD.n7567 2.2505
R37528 PAD.n7565 PAD.n7564 2.2505
R37529 PAD.n7557 PAD.n7142 2.2505
R37530 PAD.n7560 PAD.n7559 2.2505
R37531 PAD.n7556 PAD.n7555 2.2505
R37532 PAD.n7553 PAD.n7552 2.2505
R37533 PAD.n7545 PAD.n7144 2.2505
R37534 PAD.n7548 PAD.n7547 2.2505
R37535 PAD.n7544 PAD.n7543 2.2505
R37536 PAD.n7541 PAD.n7540 2.2505
R37537 PAD.n7533 PAD.n7146 2.2505
R37538 PAD.n7536 PAD.n7535 2.2505
R37539 PAD.n7532 PAD.n7531 2.2505
R37540 PAD.n7532 PAD.n7147 2.2505
R37541 PAD.n7537 PAD.n7536 2.2505
R37542 PAD.n7538 PAD.n7146 2.2505
R37543 PAD.n7540 PAD.n7539 2.2505
R37544 PAD.n7544 PAD.n7145 2.2505
R37545 PAD.n7549 PAD.n7548 2.2505
R37546 PAD.n7550 PAD.n7144 2.2505
R37547 PAD.n7552 PAD.n7551 2.2505
R37548 PAD.n7556 PAD.n7143 2.2505
R37549 PAD.n7561 PAD.n7560 2.2505
R37550 PAD.n7562 PAD.n7142 2.2505
R37551 PAD.n7564 PAD.n7563 2.2505
R37552 PAD.n7568 PAD.n7141 2.2505
R37553 PAD.n7573 PAD.n7572 2.2505
R37554 PAD.n7574 PAD.n7140 2.2505
R37555 PAD.n7576 PAD.n7575 2.2505
R37556 PAD.n7580 PAD.n7139 2.2505
R37557 PAD.n7585 PAD.n7584 2.2505
R37558 PAD.n7586 PAD.n7138 2.2505
R37559 PAD.n7588 PAD.n7587 2.2505
R37560 PAD.n7592 PAD.n7137 2.2505
R37561 PAD.n7597 PAD.n7596 2.2505
R37562 PAD.n7598 PAD.n7136 2.2505
R37563 PAD.n7600 PAD.n7599 2.2505
R37564 PAD.n7604 PAD.n7135 2.2505
R37565 PAD.n7609 PAD.n7608 2.2505
R37566 PAD.n7610 PAD.n7134 2.2505
R37567 PAD.n7612 PAD.n7611 2.2505
R37568 PAD.n7616 PAD.n7133 2.2505
R37569 PAD.n7621 PAD.n7620 2.2505
R37570 PAD.n7622 PAD.n7132 2.2505
R37571 PAD.n7624 PAD.n7623 2.2505
R37572 PAD.n7628 PAD.n7131 2.2505
R37573 PAD.n7633 PAD.n7632 2.2505
R37574 PAD.n7634 PAD.n7130 2.2505
R37575 PAD.n7636 PAD.n7635 2.2505
R37576 PAD.n7640 PAD.n7129 2.2505
R37577 PAD.n7645 PAD.n7644 2.2505
R37578 PAD.n7646 PAD.n7128 2.2505
R37579 PAD.n7648 PAD.n7647 2.2505
R37580 PAD.n7652 PAD.n7127 2.2505
R37581 PAD.n7657 PAD.n7656 2.2505
R37582 PAD.n7658 PAD.n7126 2.2505
R37583 PAD.n7660 PAD.n7659 2.2505
R37584 PAD.n7664 PAD.n7125 2.2505
R37585 PAD.n7669 PAD.n7668 2.2505
R37586 PAD.n7670 PAD.n7124 2.2505
R37587 PAD.n7672 PAD.n7671 2.2505
R37588 PAD.n7676 PAD.n7123 2.2505
R37589 PAD.n7681 PAD.n7680 2.2505
R37590 PAD.n7682 PAD.n7122 2.2505
R37591 PAD.n7684 PAD.n7683 2.2505
R37592 PAD.n7688 PAD.n7121 2.2505
R37593 PAD.n7693 PAD.n7692 2.2505
R37594 PAD.n7694 PAD.n7120 2.2505
R37595 PAD.n7696 PAD.n7695 2.2505
R37596 PAD.n7700 PAD.n7119 2.2505
R37597 PAD.n7705 PAD.n7704 2.2505
R37598 PAD.n7706 PAD.n7118 2.2505
R37599 PAD.n7708 PAD.n7707 2.2505
R37600 PAD.n7712 PAD.n7117 2.2505
R37601 PAD.n7717 PAD.n7716 2.2505
R37602 PAD.n7718 PAD.n7116 2.2505
R37603 PAD.n7720 PAD.n7719 2.2505
R37604 PAD.n7724 PAD.n7115 2.2505
R37605 PAD.n7729 PAD.n7728 2.2505
R37606 PAD.n7730 PAD.n7114 2.2505
R37607 PAD.n7732 PAD.n7731 2.2505
R37608 PAD.n7736 PAD.n7113 2.2505
R37609 PAD.n7741 PAD.n7740 2.2505
R37610 PAD.n7742 PAD.n7112 2.2505
R37611 PAD.n7744 PAD.n7743 2.2505
R37612 PAD.n7748 PAD.n7111 2.2505
R37613 PAD.n7753 PAD.n7752 2.2505
R37614 PAD.n7754 PAD.n7110 2.2505
R37615 PAD.n7756 PAD.n7755 2.2505
R37616 PAD.n7760 PAD.n7109 2.2505
R37617 PAD.n7765 PAD.n7764 2.2505
R37618 PAD.n7766 PAD.n7108 2.2505
R37619 PAD.n7768 PAD.n7767 2.2505
R37620 PAD.n7772 PAD.n7107 2.2505
R37621 PAD.n7776 PAD.n7775 2.2505
R37622 PAD.n7777 PAD.n7106 2.2505
R37623 PAD.n7779 PAD.n7778 2.2505
R37624 PAD.n7050 PAD.n6719 2.2505
R37625 PAD.n7049 PAD.n7048 2.2505
R37626 PAD.n7046 PAD.n6720 2.2505
R37627 PAD.n7044 PAD.n7043 2.2505
R37628 PAD.n7036 PAD.n6723 2.2505
R37629 PAD.n7039 PAD.n7038 2.2505
R37630 PAD.n7034 PAD.n6726 2.2505
R37631 PAD.n7032 PAD.n7031 2.2505
R37632 PAD.n7024 PAD.n6728 2.2505
R37633 PAD.n7027 PAD.n7026 2.2505
R37634 PAD.n7022 PAD.n6730 2.2505
R37635 PAD.n7020 PAD.n7019 2.2505
R37636 PAD.n7012 PAD.n6732 2.2505
R37637 PAD.n7015 PAD.n7014 2.2505
R37638 PAD.n7010 PAD.n6734 2.2505
R37639 PAD.n7008 PAD.n7007 2.2505
R37640 PAD.n7000 PAD.n6736 2.2505
R37641 PAD.n7003 PAD.n7002 2.2505
R37642 PAD.n6998 PAD.n6738 2.2505
R37643 PAD.n6996 PAD.n6995 2.2505
R37644 PAD.n6988 PAD.n6740 2.2505
R37645 PAD.n6991 PAD.n6990 2.2505
R37646 PAD.n6986 PAD.n6742 2.2505
R37647 PAD.n6984 PAD.n6983 2.2505
R37648 PAD.n6976 PAD.n6744 2.2505
R37649 PAD.n6979 PAD.n6978 2.2505
R37650 PAD.n6974 PAD.n6746 2.2505
R37651 PAD.n6972 PAD.n6971 2.2505
R37652 PAD.n6964 PAD.n6748 2.2505
R37653 PAD.n6967 PAD.n6966 2.2505
R37654 PAD.n6962 PAD.n6750 2.2505
R37655 PAD.n6960 PAD.n6959 2.2505
R37656 PAD.n6952 PAD.n6752 2.2505
R37657 PAD.n6955 PAD.n6954 2.2505
R37658 PAD.n6950 PAD.n6754 2.2505
R37659 PAD.n6948 PAD.n6947 2.2505
R37660 PAD.n6940 PAD.n6756 2.2505
R37661 PAD.n6943 PAD.n6942 2.2505
R37662 PAD.n6938 PAD.n6758 2.2505
R37663 PAD.n6936 PAD.n6935 2.2505
R37664 PAD.n6928 PAD.n6760 2.2505
R37665 PAD.n6931 PAD.n6930 2.2505
R37666 PAD.n6926 PAD.n6762 2.2505
R37667 PAD.n6924 PAD.n6923 2.2505
R37668 PAD.n6916 PAD.n6764 2.2505
R37669 PAD.n6919 PAD.n6918 2.2505
R37670 PAD.n6914 PAD.n6766 2.2505
R37671 PAD.n6912 PAD.n6911 2.2505
R37672 PAD.n6904 PAD.n6768 2.2505
R37673 PAD.n6907 PAD.n6906 2.2505
R37674 PAD.n6902 PAD.n6770 2.2505
R37675 PAD.n6900 PAD.n6899 2.2505
R37676 PAD.n6892 PAD.n6772 2.2505
R37677 PAD.n6895 PAD.n6894 2.2505
R37678 PAD.n6890 PAD.n6774 2.2505
R37679 PAD.n6888 PAD.n6887 2.2505
R37680 PAD.n6880 PAD.n6776 2.2505
R37681 PAD.n6883 PAD.n6882 2.2505
R37682 PAD.n6878 PAD.n6778 2.2505
R37683 PAD.n6876 PAD.n6875 2.2505
R37684 PAD.n6868 PAD.n6780 2.2505
R37685 PAD.n6871 PAD.n6870 2.2505
R37686 PAD.n6866 PAD.n6782 2.2505
R37687 PAD.n6864 PAD.n6863 2.2505
R37688 PAD.n6856 PAD.n6784 2.2505
R37689 PAD.n6859 PAD.n6858 2.2505
R37690 PAD.n6854 PAD.n6786 2.2505
R37691 PAD.n6852 PAD.n6851 2.2505
R37692 PAD.n6844 PAD.n6788 2.2505
R37693 PAD.n6847 PAD.n6846 2.2505
R37694 PAD.n6842 PAD.n6790 2.2505
R37695 PAD.n6840 PAD.n6839 2.2505
R37696 PAD.n6832 PAD.n6792 2.2505
R37697 PAD.n6835 PAD.n6834 2.2505
R37698 PAD.n6830 PAD.n6794 2.2505
R37699 PAD.n6828 PAD.n6827 2.2505
R37700 PAD.n6820 PAD.n6796 2.2505
R37701 PAD.n6823 PAD.n6822 2.2505
R37702 PAD.n6818 PAD.n6798 2.2505
R37703 PAD.n6816 PAD.n6815 2.2505
R37704 PAD.n6808 PAD.n6800 2.2505
R37705 PAD.n6811 PAD.n6810 2.2505
R37706 PAD.n6806 PAD.n6802 2.2505
R37707 PAD.n6804 PAD.n6803 2.2505
R37708 PAD.n6803 PAD.n6705 2.2505
R37709 PAD.n6802 PAD.n6801 2.2505
R37710 PAD.n6812 PAD.n6811 2.2505
R37711 PAD.n6813 PAD.n6800 2.2505
R37712 PAD.n6815 PAD.n6814 2.2505
R37713 PAD.n6798 PAD.n6797 2.2505
R37714 PAD.n6824 PAD.n6823 2.2505
R37715 PAD.n6825 PAD.n6796 2.2505
R37716 PAD.n6827 PAD.n6826 2.2505
R37717 PAD.n6794 PAD.n6793 2.2505
R37718 PAD.n6836 PAD.n6835 2.2505
R37719 PAD.n6837 PAD.n6792 2.2505
R37720 PAD.n6839 PAD.n6838 2.2505
R37721 PAD.n6790 PAD.n6789 2.2505
R37722 PAD.n6848 PAD.n6847 2.2505
R37723 PAD.n6849 PAD.n6788 2.2505
R37724 PAD.n6851 PAD.n6850 2.2505
R37725 PAD.n6786 PAD.n6785 2.2505
R37726 PAD.n6860 PAD.n6859 2.2505
R37727 PAD.n6861 PAD.n6784 2.2505
R37728 PAD.n6863 PAD.n6862 2.2505
R37729 PAD.n6782 PAD.n6781 2.2505
R37730 PAD.n6872 PAD.n6871 2.2505
R37731 PAD.n6873 PAD.n6780 2.2505
R37732 PAD.n6875 PAD.n6874 2.2505
R37733 PAD.n6778 PAD.n6777 2.2505
R37734 PAD.n6884 PAD.n6883 2.2505
R37735 PAD.n6885 PAD.n6776 2.2505
R37736 PAD.n6887 PAD.n6886 2.2505
R37737 PAD.n6774 PAD.n6773 2.2505
R37738 PAD.n6896 PAD.n6895 2.2505
R37739 PAD.n6897 PAD.n6772 2.2505
R37740 PAD.n6899 PAD.n6898 2.2505
R37741 PAD.n6770 PAD.n6769 2.2505
R37742 PAD.n6908 PAD.n6907 2.2505
R37743 PAD.n6909 PAD.n6768 2.2505
R37744 PAD.n6911 PAD.n6910 2.2505
R37745 PAD.n6766 PAD.n6765 2.2505
R37746 PAD.n6920 PAD.n6919 2.2505
R37747 PAD.n6921 PAD.n6764 2.2505
R37748 PAD.n6923 PAD.n6922 2.2505
R37749 PAD.n6762 PAD.n6761 2.2505
R37750 PAD.n6932 PAD.n6931 2.2505
R37751 PAD.n6933 PAD.n6760 2.2505
R37752 PAD.n6935 PAD.n6934 2.2505
R37753 PAD.n6758 PAD.n6757 2.2505
R37754 PAD.n6944 PAD.n6943 2.2505
R37755 PAD.n6945 PAD.n6756 2.2505
R37756 PAD.n6947 PAD.n6946 2.2505
R37757 PAD.n6754 PAD.n6753 2.2505
R37758 PAD.n6956 PAD.n6955 2.2505
R37759 PAD.n6957 PAD.n6752 2.2505
R37760 PAD.n6959 PAD.n6958 2.2505
R37761 PAD.n6750 PAD.n6749 2.2505
R37762 PAD.n6968 PAD.n6967 2.2505
R37763 PAD.n6969 PAD.n6748 2.2505
R37764 PAD.n6971 PAD.n6970 2.2505
R37765 PAD.n6746 PAD.n6745 2.2505
R37766 PAD.n6980 PAD.n6979 2.2505
R37767 PAD.n6981 PAD.n6744 2.2505
R37768 PAD.n6983 PAD.n6982 2.2505
R37769 PAD.n6742 PAD.n6741 2.2505
R37770 PAD.n6992 PAD.n6991 2.2505
R37771 PAD.n6993 PAD.n6740 2.2505
R37772 PAD.n6995 PAD.n6994 2.2505
R37773 PAD.n6738 PAD.n6737 2.2505
R37774 PAD.n7004 PAD.n7003 2.2505
R37775 PAD.n7005 PAD.n6736 2.2505
R37776 PAD.n7007 PAD.n7006 2.2505
R37777 PAD.n6734 PAD.n6733 2.2505
R37778 PAD.n7016 PAD.n7015 2.2505
R37779 PAD.n7017 PAD.n6732 2.2505
R37780 PAD.n7019 PAD.n7018 2.2505
R37781 PAD.n6730 PAD.n6729 2.2505
R37782 PAD.n7028 PAD.n7027 2.2505
R37783 PAD.n7029 PAD.n6728 2.2505
R37784 PAD.n7031 PAD.n7030 2.2505
R37785 PAD.n6726 PAD.n6725 2.2505
R37786 PAD.n7040 PAD.n7039 2.2505
R37787 PAD.n7041 PAD.n6723 2.2505
R37788 PAD.n7043 PAD.n7042 2.2505
R37789 PAD.n6724 PAD.n6720 2.2505
R37790 PAD.n7049 PAD.n6718 2.2505
R37791 PAD.n7051 PAD.n7050 2.2505
R37792 PAD.n5892 PAD.n5891 2.2505
R37793 PAD.n5890 PAD.n5602 2.2505
R37794 PAD.n5605 PAD.n5604 2.2505
R37795 PAD.n5886 PAD.n5885 2.2505
R37796 PAD.n5883 PAD.n5882 2.2505
R37797 PAD.n5881 PAD.n5610 2.2505
R37798 PAD.n5608 PAD.n5607 2.2505
R37799 PAD.n5877 PAD.n5876 2.2505
R37800 PAD.n5874 PAD.n5873 2.2505
R37801 PAD.n5872 PAD.n5615 2.2505
R37802 PAD.n5613 PAD.n5612 2.2505
R37803 PAD.n5868 PAD.n5867 2.2505
R37804 PAD.n5865 PAD.n5864 2.2505
R37805 PAD.n5863 PAD.n5620 2.2505
R37806 PAD.n5618 PAD.n5617 2.2505
R37807 PAD.n5859 PAD.n5858 2.2505
R37808 PAD.n5856 PAD.n5855 2.2505
R37809 PAD.n5854 PAD.n5625 2.2505
R37810 PAD.n5623 PAD.n5622 2.2505
R37811 PAD.n5850 PAD.n5849 2.2505
R37812 PAD.n5847 PAD.n5846 2.2505
R37813 PAD.n5845 PAD.n5630 2.2505
R37814 PAD.n5628 PAD.n5627 2.2505
R37815 PAD.n5841 PAD.n5840 2.2505
R37816 PAD.n5838 PAD.n5837 2.2505
R37817 PAD.n5836 PAD.n5635 2.2505
R37818 PAD.n5633 PAD.n5632 2.2505
R37819 PAD.n5832 PAD.n5831 2.2505
R37820 PAD.n5829 PAD.n5828 2.2505
R37821 PAD.n5827 PAD.n5640 2.2505
R37822 PAD.n5638 PAD.n5637 2.2505
R37823 PAD.n5823 PAD.n5822 2.2505
R37824 PAD.n5820 PAD.n5819 2.2505
R37825 PAD.n5818 PAD.n5645 2.2505
R37826 PAD.n5643 PAD.n5642 2.2505
R37827 PAD.n5814 PAD.n5813 2.2505
R37828 PAD.n5811 PAD.n5810 2.2505
R37829 PAD.n5809 PAD.n5650 2.2505
R37830 PAD.n5648 PAD.n5647 2.2505
R37831 PAD.n5805 PAD.n5804 2.2505
R37832 PAD.n5802 PAD.n5801 2.2505
R37833 PAD.n5800 PAD.n5655 2.2505
R37834 PAD.n5653 PAD.n5652 2.2505
R37835 PAD.n5796 PAD.n5795 2.2505
R37836 PAD.n5793 PAD.n5792 2.2505
R37837 PAD.n5791 PAD.n5660 2.2505
R37838 PAD.n5658 PAD.n5657 2.2505
R37839 PAD.n5787 PAD.n5786 2.2505
R37840 PAD.n5784 PAD.n5783 2.2505
R37841 PAD.n5782 PAD.n5665 2.2505
R37842 PAD.n5663 PAD.n5662 2.2505
R37843 PAD.n5778 PAD.n5777 2.2505
R37844 PAD.n5775 PAD.n5774 2.2505
R37845 PAD.n5773 PAD.n5670 2.2505
R37846 PAD.n5668 PAD.n5667 2.2505
R37847 PAD.n5769 PAD.n5768 2.2505
R37848 PAD.n5766 PAD.n5765 2.2505
R37849 PAD.n5764 PAD.n5675 2.2505
R37850 PAD.n5673 PAD.n5672 2.2505
R37851 PAD.n5760 PAD.n5759 2.2505
R37852 PAD.n5757 PAD.n5756 2.2505
R37853 PAD.n5755 PAD.n5680 2.2505
R37854 PAD.n5678 PAD.n5677 2.2505
R37855 PAD.n5751 PAD.n5750 2.2505
R37856 PAD.n5748 PAD.n5747 2.2505
R37857 PAD.n5746 PAD.n5685 2.2505
R37858 PAD.n5683 PAD.n5682 2.2505
R37859 PAD.n5742 PAD.n5741 2.2505
R37860 PAD.n5739 PAD.n5738 2.2505
R37861 PAD.n5737 PAD.n5690 2.2505
R37862 PAD.n5688 PAD.n5687 2.2505
R37863 PAD.n5733 PAD.n5732 2.2505
R37864 PAD.n5730 PAD.n5729 2.2505
R37865 PAD.n5728 PAD.n5695 2.2505
R37866 PAD.n5693 PAD.n5692 2.2505
R37867 PAD.n5724 PAD.n5723 2.2505
R37868 PAD.n5721 PAD.n5720 2.2505
R37869 PAD.n5719 PAD.n5700 2.2505
R37870 PAD.n5698 PAD.n5697 2.2505
R37871 PAD.n5715 PAD.n5714 2.2505
R37872 PAD.n5712 PAD.n5711 2.2505
R37873 PAD.n5710 PAD.n5707 2.2505
R37874 PAD.n5705 PAD.n5704 2.2505
R37875 PAD.n5703 PAD.n5702 2.2505
R37876 PAD.n5703 PAD.n5557 2.2505
R37877 PAD.n5708 PAD.n5704 2.2505
R37878 PAD.n5710 PAD.n5709 2.2505
R37879 PAD.n5711 PAD.n5701 2.2505
R37880 PAD.n5716 PAD.n5715 2.2505
R37881 PAD.n5717 PAD.n5697 2.2505
R37882 PAD.n5719 PAD.n5718 2.2505
R37883 PAD.n5720 PAD.n5696 2.2505
R37884 PAD.n5725 PAD.n5724 2.2505
R37885 PAD.n5726 PAD.n5692 2.2505
R37886 PAD.n5728 PAD.n5727 2.2505
R37887 PAD.n5729 PAD.n5691 2.2505
R37888 PAD.n5734 PAD.n5733 2.2505
R37889 PAD.n5735 PAD.n5687 2.2505
R37890 PAD.n5737 PAD.n5736 2.2505
R37891 PAD.n5738 PAD.n5686 2.2505
R37892 PAD.n5743 PAD.n5742 2.2505
R37893 PAD.n5744 PAD.n5682 2.2505
R37894 PAD.n5746 PAD.n5745 2.2505
R37895 PAD.n5747 PAD.n5681 2.2505
R37896 PAD.n5752 PAD.n5751 2.2505
R37897 PAD.n5753 PAD.n5677 2.2505
R37898 PAD.n5755 PAD.n5754 2.2505
R37899 PAD.n5756 PAD.n5676 2.2505
R37900 PAD.n5761 PAD.n5760 2.2505
R37901 PAD.n5762 PAD.n5672 2.2505
R37902 PAD.n5764 PAD.n5763 2.2505
R37903 PAD.n5765 PAD.n5671 2.2505
R37904 PAD.n5770 PAD.n5769 2.2505
R37905 PAD.n5771 PAD.n5667 2.2505
R37906 PAD.n5773 PAD.n5772 2.2505
R37907 PAD.n5774 PAD.n5666 2.2505
R37908 PAD.n5779 PAD.n5778 2.2505
R37909 PAD.n5780 PAD.n5662 2.2505
R37910 PAD.n5782 PAD.n5781 2.2505
R37911 PAD.n5783 PAD.n5661 2.2505
R37912 PAD.n5788 PAD.n5787 2.2505
R37913 PAD.n5789 PAD.n5657 2.2505
R37914 PAD.n5791 PAD.n5790 2.2505
R37915 PAD.n5792 PAD.n5656 2.2505
R37916 PAD.n5797 PAD.n5796 2.2505
R37917 PAD.n5798 PAD.n5652 2.2505
R37918 PAD.n5800 PAD.n5799 2.2505
R37919 PAD.n5801 PAD.n5651 2.2505
R37920 PAD.n5806 PAD.n5805 2.2505
R37921 PAD.n5807 PAD.n5647 2.2505
R37922 PAD.n5809 PAD.n5808 2.2505
R37923 PAD.n5810 PAD.n5646 2.2505
R37924 PAD.n5815 PAD.n5814 2.2505
R37925 PAD.n5816 PAD.n5642 2.2505
R37926 PAD.n5818 PAD.n5817 2.2505
R37927 PAD.n5819 PAD.n5641 2.2505
R37928 PAD.n5824 PAD.n5823 2.2505
R37929 PAD.n5825 PAD.n5637 2.2505
R37930 PAD.n5827 PAD.n5826 2.2505
R37931 PAD.n5828 PAD.n5636 2.2505
R37932 PAD.n5833 PAD.n5832 2.2505
R37933 PAD.n5834 PAD.n5632 2.2505
R37934 PAD.n5836 PAD.n5835 2.2505
R37935 PAD.n5837 PAD.n5631 2.2505
R37936 PAD.n5842 PAD.n5841 2.2505
R37937 PAD.n5843 PAD.n5627 2.2505
R37938 PAD.n5845 PAD.n5844 2.2505
R37939 PAD.n5846 PAD.n5626 2.2505
R37940 PAD.n5851 PAD.n5850 2.2505
R37941 PAD.n5852 PAD.n5622 2.2505
R37942 PAD.n5854 PAD.n5853 2.2505
R37943 PAD.n5855 PAD.n5621 2.2505
R37944 PAD.n5860 PAD.n5859 2.2505
R37945 PAD.n5861 PAD.n5617 2.2505
R37946 PAD.n5863 PAD.n5862 2.2505
R37947 PAD.n5864 PAD.n5616 2.2505
R37948 PAD.n5869 PAD.n5868 2.2505
R37949 PAD.n5870 PAD.n5612 2.2505
R37950 PAD.n5872 PAD.n5871 2.2505
R37951 PAD.n5873 PAD.n5611 2.2505
R37952 PAD.n5878 PAD.n5877 2.2505
R37953 PAD.n5879 PAD.n5607 2.2505
R37954 PAD.n5881 PAD.n5880 2.2505
R37955 PAD.n5882 PAD.n5606 2.2505
R37956 PAD.n5887 PAD.n5886 2.2505
R37957 PAD.n5888 PAD.n5605 2.2505
R37958 PAD.n5890 PAD.n5889 2.2505
R37959 PAD.n5891 PAD.n5545 2.2505
R37960 PAD.n6687 PAD.n5951 2.2505
R37961 PAD.n6672 PAD.n5950 2.2505
R37962 PAD.n6673 PAD.n6439 2.2505
R37963 PAD.n6675 PAD.n6674 2.2505
R37964 PAD.n6671 PAD.n6438 2.2505
R37965 PAD.n6670 PAD.n6669 2.2505
R37966 PAD.n6667 PAD.n6440 2.2505
R37967 PAD.n6665 PAD.n6663 2.2505
R37968 PAD.n6662 PAD.n6442 2.2505
R37969 PAD.n6661 PAD.n6660 2.2505
R37970 PAD.n6658 PAD.n6443 2.2505
R37971 PAD.n6656 PAD.n6654 2.2505
R37972 PAD.n6653 PAD.n6445 2.2505
R37973 PAD.n6652 PAD.n6651 2.2505
R37974 PAD.n6649 PAD.n6446 2.2505
R37975 PAD.n6647 PAD.n6645 2.2505
R37976 PAD.n6644 PAD.n6448 2.2505
R37977 PAD.n6643 PAD.n6642 2.2505
R37978 PAD.n6640 PAD.n6449 2.2505
R37979 PAD.n6638 PAD.n6636 2.2505
R37980 PAD.n6635 PAD.n6451 2.2505
R37981 PAD.n6634 PAD.n6633 2.2505
R37982 PAD.n6631 PAD.n6452 2.2505
R37983 PAD.n6629 PAD.n6627 2.2505
R37984 PAD.n6626 PAD.n6454 2.2505
R37985 PAD.n6625 PAD.n6624 2.2505
R37986 PAD.n6622 PAD.n6455 2.2505
R37987 PAD.n6620 PAD.n6618 2.2505
R37988 PAD.n6617 PAD.n6457 2.2505
R37989 PAD.n6616 PAD.n6615 2.2505
R37990 PAD.n6613 PAD.n6458 2.2505
R37991 PAD.n6611 PAD.n6609 2.2505
R37992 PAD.n6608 PAD.n6460 2.2505
R37993 PAD.n6607 PAD.n6606 2.2505
R37994 PAD.n6604 PAD.n6461 2.2505
R37995 PAD.n6602 PAD.n6600 2.2505
R37996 PAD.n6599 PAD.n6463 2.2505
R37997 PAD.n6598 PAD.n6597 2.2505
R37998 PAD.n6595 PAD.n6464 2.2505
R37999 PAD.n6593 PAD.n6591 2.2505
R38000 PAD.n6590 PAD.n6466 2.2505
R38001 PAD.n6589 PAD.n6588 2.2505
R38002 PAD.n6586 PAD.n6467 2.2505
R38003 PAD.n6584 PAD.n6582 2.2505
R38004 PAD.n6581 PAD.n6469 2.2505
R38005 PAD.n6580 PAD.n6579 2.2505
R38006 PAD.n6577 PAD.n6470 2.2505
R38007 PAD.n6575 PAD.n6573 2.2505
R38008 PAD.n6572 PAD.n6472 2.2505
R38009 PAD.n6571 PAD.n6570 2.2505
R38010 PAD.n6568 PAD.n6473 2.2505
R38011 PAD.n6566 PAD.n6564 2.2505
R38012 PAD.n6563 PAD.n6475 2.2505
R38013 PAD.n6562 PAD.n6561 2.2505
R38014 PAD.n6559 PAD.n6476 2.2505
R38015 PAD.n6557 PAD.n6555 2.2505
R38016 PAD.n6554 PAD.n6478 2.2505
R38017 PAD.n6553 PAD.n6552 2.2505
R38018 PAD.n6550 PAD.n6479 2.2505
R38019 PAD.n6548 PAD.n6546 2.2505
R38020 PAD.n6545 PAD.n6481 2.2505
R38021 PAD.n6544 PAD.n6543 2.2505
R38022 PAD.n6541 PAD.n6482 2.2505
R38023 PAD.n6539 PAD.n6537 2.2505
R38024 PAD.n6536 PAD.n6484 2.2505
R38025 PAD.n6535 PAD.n6534 2.2505
R38026 PAD.n6532 PAD.n6485 2.2505
R38027 PAD.n6530 PAD.n6528 2.2505
R38028 PAD.n6527 PAD.n6487 2.2505
R38029 PAD.n6526 PAD.n6525 2.2505
R38030 PAD.n6523 PAD.n6488 2.2505
R38031 PAD.n6521 PAD.n6519 2.2505
R38032 PAD.n6518 PAD.n6490 2.2505
R38033 PAD.n6517 PAD.n6516 2.2505
R38034 PAD.n6514 PAD.n6491 2.2505
R38035 PAD.n6512 PAD.n6510 2.2505
R38036 PAD.n6509 PAD.n6493 2.2505
R38037 PAD.n6508 PAD.n6507 2.2505
R38038 PAD.n6505 PAD.n6494 2.2505
R38039 PAD.n6503 PAD.n6501 2.2505
R38040 PAD.n6500 PAD.n6496 2.2505
R38041 PAD.n6499 PAD.n6498 2.2505
R38042 PAD.n5900 PAD.n5898 2.2505
R38043 PAD.n6692 PAD.n6691 2.2505
R38044 PAD.n75 PAD.n26 2.2505
R38045 PAD.n363 PAD.n362 2.2505
R38046 PAD.n361 PAD.n76 2.2505
R38047 PAD.n360 PAD.n359 2.2505
R38048 PAD.n355 PAD.n77 2.2505
R38049 PAD.n351 PAD.n350 2.2505
R38050 PAD.n349 PAD.n78 2.2505
R38051 PAD.n348 PAD.n347 2.2505
R38052 PAD.n343 PAD.n79 2.2505
R38053 PAD.n339 PAD.n338 2.2505
R38054 PAD.n337 PAD.n80 2.2505
R38055 PAD.n336 PAD.n335 2.2505
R38056 PAD.n331 PAD.n81 2.2505
R38057 PAD.n327 PAD.n326 2.2505
R38058 PAD.n325 PAD.n82 2.2505
R38059 PAD.n324 PAD.n323 2.2505
R38060 PAD.n319 PAD.n83 2.2505
R38061 PAD.n315 PAD.n314 2.2505
R38062 PAD.n313 PAD.n84 2.2505
R38063 PAD.n312 PAD.n311 2.2505
R38064 PAD.n307 PAD.n85 2.2505
R38065 PAD.n303 PAD.n302 2.2505
R38066 PAD.n301 PAD.n86 2.2505
R38067 PAD.n300 PAD.n299 2.2505
R38068 PAD.n295 PAD.n87 2.2505
R38069 PAD.n291 PAD.n290 2.2505
R38070 PAD.n289 PAD.n88 2.2505
R38071 PAD.n288 PAD.n287 2.2505
R38072 PAD.n283 PAD.n89 2.2505
R38073 PAD.n279 PAD.n278 2.2505
R38074 PAD.n277 PAD.n90 2.2505
R38075 PAD.n276 PAD.n275 2.2505
R38076 PAD.n271 PAD.n91 2.2505
R38077 PAD.n267 PAD.n266 2.2505
R38078 PAD.n265 PAD.n92 2.2505
R38079 PAD.n264 PAD.n263 2.2505
R38080 PAD.n259 PAD.n93 2.2505
R38081 PAD.n255 PAD.n254 2.2505
R38082 PAD.n253 PAD.n94 2.2505
R38083 PAD.n252 PAD.n251 2.2505
R38084 PAD.n247 PAD.n95 2.2505
R38085 PAD.n243 PAD.n242 2.2505
R38086 PAD.n241 PAD.n96 2.2505
R38087 PAD.n240 PAD.n239 2.2505
R38088 PAD.n235 PAD.n97 2.2505
R38089 PAD.n231 PAD.n230 2.2505
R38090 PAD.n229 PAD.n98 2.2505
R38091 PAD.n228 PAD.n227 2.2505
R38092 PAD.n223 PAD.n99 2.2505
R38093 PAD.n219 PAD.n218 2.2505
R38094 PAD.n217 PAD.n100 2.2505
R38095 PAD.n216 PAD.n215 2.2505
R38096 PAD.n211 PAD.n101 2.2505
R38097 PAD.n207 PAD.n206 2.2505
R38098 PAD.n205 PAD.n102 2.2505
R38099 PAD.n204 PAD.n203 2.2505
R38100 PAD.n199 PAD.n103 2.2505
R38101 PAD.n195 PAD.n194 2.2505
R38102 PAD.n193 PAD.n104 2.2505
R38103 PAD.n192 PAD.n191 2.2505
R38104 PAD.n187 PAD.n105 2.2505
R38105 PAD.n183 PAD.n182 2.2505
R38106 PAD.n181 PAD.n106 2.2505
R38107 PAD.n180 PAD.n179 2.2505
R38108 PAD.n175 PAD.n107 2.2505
R38109 PAD.n171 PAD.n170 2.2505
R38110 PAD.n169 PAD.n108 2.2505
R38111 PAD.n168 PAD.n167 2.2505
R38112 PAD.n163 PAD.n109 2.2505
R38113 PAD.n159 PAD.n158 2.2505
R38114 PAD.n157 PAD.n110 2.2505
R38115 PAD.n156 PAD.n155 2.2505
R38116 PAD.n151 PAD.n111 2.2505
R38117 PAD.n147 PAD.n146 2.2505
R38118 PAD.n145 PAD.n112 2.2505
R38119 PAD.n144 PAD.n143 2.2505
R38120 PAD.n139 PAD.n113 2.2505
R38121 PAD.n135 PAD.n134 2.2505
R38122 PAD.n133 PAD.n114 2.2505
R38123 PAD.n132 PAD.n131 2.2505
R38124 PAD.n127 PAD.n115 2.2505
R38125 PAD.n123 PAD.n122 2.2505
R38126 PAD.n121 PAD.n118 2.2505
R38127 PAD.n120 PAD.n119 2.2505
R38128 PAD.n119 PAD.n74 2.2505
R38129 PAD.n118 PAD.n117 2.2505
R38130 PAD.n124 PAD.n123 2.2505
R38131 PAD.n127 PAD.n126 2.2505
R38132 PAD.n131 PAD.n130 2.2505
R38133 PAD.n128 PAD.n114 2.2505
R38134 PAD.n136 PAD.n135 2.2505
R38135 PAD.n139 PAD.n138 2.2505
R38136 PAD.n143 PAD.n142 2.2505
R38137 PAD.n140 PAD.n112 2.2505
R38138 PAD.n148 PAD.n147 2.2505
R38139 PAD.n151 PAD.n150 2.2505
R38140 PAD.n155 PAD.n154 2.2505
R38141 PAD.n152 PAD.n110 2.2505
R38142 PAD.n160 PAD.n159 2.2505
R38143 PAD.n163 PAD.n162 2.2505
R38144 PAD.n167 PAD.n166 2.2505
R38145 PAD.n164 PAD.n108 2.2505
R38146 PAD.n172 PAD.n171 2.2505
R38147 PAD.n175 PAD.n174 2.2505
R38148 PAD.n179 PAD.n178 2.2505
R38149 PAD.n176 PAD.n106 2.2505
R38150 PAD.n184 PAD.n183 2.2505
R38151 PAD.n187 PAD.n186 2.2505
R38152 PAD.n191 PAD.n190 2.2505
R38153 PAD.n188 PAD.n104 2.2505
R38154 PAD.n196 PAD.n195 2.2505
R38155 PAD.n199 PAD.n198 2.2505
R38156 PAD.n203 PAD.n202 2.2505
R38157 PAD.n200 PAD.n102 2.2505
R38158 PAD.n208 PAD.n207 2.2505
R38159 PAD.n211 PAD.n210 2.2505
R38160 PAD.n215 PAD.n214 2.2505
R38161 PAD.n212 PAD.n100 2.2505
R38162 PAD.n220 PAD.n219 2.2505
R38163 PAD.n223 PAD.n222 2.2505
R38164 PAD.n227 PAD.n226 2.2505
R38165 PAD.n224 PAD.n98 2.2505
R38166 PAD.n232 PAD.n231 2.2505
R38167 PAD.n235 PAD.n234 2.2505
R38168 PAD.n239 PAD.n238 2.2505
R38169 PAD.n236 PAD.n96 2.2505
R38170 PAD.n244 PAD.n243 2.2505
R38171 PAD.n247 PAD.n246 2.2505
R38172 PAD.n251 PAD.n250 2.2505
R38173 PAD.n248 PAD.n94 2.2505
R38174 PAD.n256 PAD.n255 2.2505
R38175 PAD.n259 PAD.n258 2.2505
R38176 PAD.n263 PAD.n262 2.2505
R38177 PAD.n260 PAD.n92 2.2505
R38178 PAD.n268 PAD.n267 2.2505
R38179 PAD.n271 PAD.n270 2.2505
R38180 PAD.n275 PAD.n274 2.2505
R38181 PAD.n272 PAD.n90 2.2505
R38182 PAD.n280 PAD.n279 2.2505
R38183 PAD.n283 PAD.n282 2.2505
R38184 PAD.n287 PAD.n286 2.2505
R38185 PAD.n284 PAD.n88 2.2505
R38186 PAD.n292 PAD.n291 2.2505
R38187 PAD.n295 PAD.n294 2.2505
R38188 PAD.n299 PAD.n298 2.2505
R38189 PAD.n296 PAD.n86 2.2505
R38190 PAD.n304 PAD.n303 2.2505
R38191 PAD.n307 PAD.n306 2.2505
R38192 PAD.n311 PAD.n310 2.2505
R38193 PAD.n308 PAD.n84 2.2505
R38194 PAD.n316 PAD.n315 2.2505
R38195 PAD.n319 PAD.n318 2.2505
R38196 PAD.n323 PAD.n322 2.2505
R38197 PAD.n320 PAD.n82 2.2505
R38198 PAD.n328 PAD.n327 2.2505
R38199 PAD.n331 PAD.n330 2.2505
R38200 PAD.n335 PAD.n334 2.2505
R38201 PAD.n332 PAD.n80 2.2505
R38202 PAD.n340 PAD.n339 2.2505
R38203 PAD.n343 PAD.n342 2.2505
R38204 PAD.n347 PAD.n346 2.2505
R38205 PAD.n344 PAD.n78 2.2505
R38206 PAD.n352 PAD.n351 2.2505
R38207 PAD.n355 PAD.n354 2.2505
R38208 PAD.n359 PAD.n358 2.2505
R38209 PAD.n356 PAD.n76 2.2505
R38210 PAD.n364 PAD.n363 2.2505
R38211 PAD.n366 PAD.n75 2.2505
R38212 PAD.n6381 PAD.n6380 2.2505
R38213 PAD.n6379 PAD.n5977 2.2505
R38214 PAD.n6378 PAD.n5952 2.2505
R38215 PAD.n6685 PAD.n5953 2.2505
R38216 PAD.n5559 PAD.n5558 2.2505
R38217 PAD.n6703 PAD.n6702 2.2505
R38218 PAD.n7799 PAD.n7798 2.2505
R38219 PAD.n7797 PAD.n5556 2.2505
R38220 PAD.n7795 PAD.n7794 2.2505
R38221 PAD.n6708 PAD.n6706 2.2505
R38222 PAD.n7153 PAD.n7152 2.2505
R38223 PAD.n7527 PAD.n7526 2.2505
R38224 PAD.n7525 PAD.n7151 2.2505
R38225 PAD.n7524 PAD.n7523 2.2505
R38226 PAD.n7204 PAD.n7203 2.2505
R38227 PAD.n5202 PAD.n5201 2.2505
R38228 PAD.n7823 PAD.n7822 2.2505
R38229 PAD.n7826 PAD.n7825 2.2505
R38230 PAD.n5188 PAD.n5187 2.2505
R38231 PAD.n8178 PAD.n8177 2.2505
R38232 PAD.n8181 PAD.n8180 2.2505
R38233 PAD.n4837 PAD.n4836 2.2505
R38234 PAD.n8198 PAD.n8197 2.2505
R38235 PAD.n8201 PAD.n8200 2.2505
R38236 PAD.n8202 PAD.n4830 2.2505
R38237 PAD.n8208 PAD.n8207 2.2505
R38238 PAD.n4671 PAD.n4670 2.2505
R38239 PAD.n8413 PAD.n8412 2.2505
R38240 PAD.n8417 PAD.n8416 2.2505
R38241 PAD.n8415 PAD.n4317 2.2505
R38242 PAD.n8433 PAD.n4315 2.2505
R38243 PAD.n8436 PAD.n8435 2.2505
R38244 PAD.n4316 PAD.n3975 2.2505
R38245 PAD.n8457 PAD.n3974 2.2505
R38246 PAD.n8460 PAD.n8459 2.2505
R38247 PAD.n3630 PAD.n3629 2.2505
R38248 PAD.n8483 PAD.n8482 2.2505
R38249 PAD.n8484 PAD.n3285 2.2505
R38250 PAD.n8505 PAD.n3284 2.2505
R38251 PAD.n8509 PAD.n8508 2.2505
R38252 PAD.n2900 PAD.n2899 2.2505
R38253 PAD.n8825 PAD.n8824 2.2505
R38254 PAD.n8827 PAD.n2896 2.2505
R38255 PAD.n8829 PAD.n8828 2.2505
R38256 PAD.n2897 PAD.n2882 2.2505
R38257 PAD.n9132 PAD.n9131 2.2505
R38258 PAD.n2492 PAD.n2491 2.2505
R38259 PAD.n9155 PAD.n9154 2.2505
R38260 PAD.n9158 PAD.n9157 2.2505
R38261 PAD.n2144 PAD.n2143 2.2505
R38262 PAD.n9179 PAD.n9178 2.2505
R38263 PAD.n9182 PAD.n9181 2.2505
R38264 PAD.n2042 PAD.n2041 2.2505
R38265 PAD.n9449 PAD.n9448 2.2505
R38266 PAD.n9451 PAD.n2039 2.2505
R38267 PAD.n9453 PAD.n9452 2.2505
R38268 PAD.n9716 PAD.n9715 2.2505
R38269 PAD.n9717 PAD.n1938 2.2505
R38270 PAD.n9719 PAD.n9718 2.2505
R38271 PAD.n9736 PAD.n9735 2.2505
R38272 PAD.n9737 PAD.n1588 2.2505
R38273 PAD.n9739 PAD.n9738 2.2505
R38274 PAD.n10002 PAD.n10001 2.2505
R38275 PAD.n10003 PAD.n1485 2.2505
R38276 PAD.n10005 PAD.n10004 2.2505
R38277 PAD.n10020 PAD.n10019 2.2505
R38278 PAD.n10021 PAD.n1135 2.2505
R38279 PAD.n10359 PAD.n10358 2.2505
R38280 PAD.n10356 PAD.n1116 2.2505
R38281 PAD.n10376 PAD.n1115 2.2505
R38282 PAD.n10380 PAD.n10379 2.2505
R38283 PAD.n774 PAD.n773 2.2505
R38284 PAD.n10401 PAD.n10400 2.2505
R38285 PAD.n10405 PAD.n10404 2.2505
R38286 PAD.n10403 PAD.n423 2.2505
R38287 PAD.n10704 PAD.n422 2.2505
R38288 PAD.n10708 PAD.n10707 2.2505
R38289 PAD.n28 PAD.n27 2.2505
R38290 PAD.n10731 PAD.n10730 2.2505
R38291 PAD.n10733 PAD.n24 2.2505
R38292 PAD.n11530 PAD.n11529 2.2505
R38293 PAD.n11528 PAD.n25 2.2505
R38294 PAD.n11526 PAD.n11525 2.2505
R38295 PAD.n10737 PAD.n10735 2.2505
R38296 PAD.n11504 PAD.n11503 2.2505
R38297 PAD.n10838 PAD.n10734 2.2505
R38298 PAD.n10840 PAD.n10839 2.2505
R38299 PAD.n10835 PAD.n10834 2.2505
R38300 PAD.n10849 PAD.n10848 2.2505
R38301 PAD.n10850 PAD.n10833 2.2505
R38302 PAD.n10852 PAD.n10851 2.2505
R38303 PAD.n10831 PAD.n10830 2.2505
R38304 PAD.n10861 PAD.n10860 2.2505
R38305 PAD.n10862 PAD.n10829 2.2505
R38306 PAD.n10864 PAD.n10863 2.2505
R38307 PAD.n10827 PAD.n10826 2.2505
R38308 PAD.n10873 PAD.n10872 2.2505
R38309 PAD.n10874 PAD.n10825 2.2505
R38310 PAD.n10876 PAD.n10875 2.2505
R38311 PAD.n10823 PAD.n10822 2.2505
R38312 PAD.n10885 PAD.n10884 2.2505
R38313 PAD.n10886 PAD.n10821 2.2505
R38314 PAD.n10888 PAD.n10887 2.2505
R38315 PAD.n10819 PAD.n10818 2.2505
R38316 PAD.n10897 PAD.n10896 2.2505
R38317 PAD.n10898 PAD.n10817 2.2505
R38318 PAD.n10900 PAD.n10899 2.2505
R38319 PAD.n10815 PAD.n10814 2.2505
R38320 PAD.n10909 PAD.n10908 2.2505
R38321 PAD.n10910 PAD.n10813 2.2505
R38322 PAD.n10912 PAD.n10911 2.2505
R38323 PAD.n10811 PAD.n10810 2.2505
R38324 PAD.n10921 PAD.n10920 2.2505
R38325 PAD.n10922 PAD.n10809 2.2505
R38326 PAD.n10924 PAD.n10923 2.2505
R38327 PAD.n10807 PAD.n10806 2.2505
R38328 PAD.n10933 PAD.n10932 2.2505
R38329 PAD.n10934 PAD.n10805 2.2505
R38330 PAD.n10936 PAD.n10935 2.2505
R38331 PAD.n10803 PAD.n10802 2.2505
R38332 PAD.n10945 PAD.n10944 2.2505
R38333 PAD.n10946 PAD.n10801 2.2505
R38334 PAD.n10948 PAD.n10947 2.2505
R38335 PAD.n10799 PAD.n10798 2.2505
R38336 PAD.n10957 PAD.n10956 2.2505
R38337 PAD.n10958 PAD.n10797 2.2505
R38338 PAD.n10960 PAD.n10959 2.2505
R38339 PAD.n10795 PAD.n10794 2.2505
R38340 PAD.n10969 PAD.n10968 2.2505
R38341 PAD.n10970 PAD.n10793 2.2505
R38342 PAD.n10972 PAD.n10971 2.2505
R38343 PAD.n10791 PAD.n10790 2.2505
R38344 PAD.n10981 PAD.n10980 2.2505
R38345 PAD.n10982 PAD.n10789 2.2505
R38346 PAD.n10984 PAD.n10983 2.2505
R38347 PAD.n10787 PAD.n10786 2.2505
R38348 PAD.n10993 PAD.n10992 2.2505
R38349 PAD.n10994 PAD.n10785 2.2505
R38350 PAD.n10996 PAD.n10995 2.2505
R38351 PAD.n10783 PAD.n10782 2.2505
R38352 PAD.n11005 PAD.n11004 2.2505
R38353 PAD.n11006 PAD.n10781 2.2505
R38354 PAD.n11008 PAD.n11007 2.2505
R38355 PAD.n10779 PAD.n10778 2.2505
R38356 PAD.n11017 PAD.n11016 2.2505
R38357 PAD.n11018 PAD.n10777 2.2505
R38358 PAD.n11020 PAD.n11019 2.2505
R38359 PAD.n10775 PAD.n10774 2.2505
R38360 PAD.n11029 PAD.n11028 2.2505
R38361 PAD.n11030 PAD.n10773 2.2505
R38362 PAD.n11032 PAD.n11031 2.2505
R38363 PAD.n10771 PAD.n10770 2.2505
R38364 PAD.n11041 PAD.n11040 2.2505
R38365 PAD.n11042 PAD.n10769 2.2505
R38366 PAD.n11044 PAD.n11043 2.2505
R38367 PAD.n10767 PAD.n10766 2.2505
R38368 PAD.n11053 PAD.n11052 2.2505
R38369 PAD.n11054 PAD.n10765 2.2505
R38370 PAD.n11056 PAD.n11055 2.2505
R38371 PAD.n10763 PAD.n10762 2.2505
R38372 PAD.n11065 PAD.n11064 2.2505
R38373 PAD.n11066 PAD.n10761 2.2505
R38374 PAD.n11068 PAD.n11067 2.2505
R38375 PAD.n10759 PAD.n10758 2.2505
R38376 PAD.n11077 PAD.n11076 2.2505
R38377 PAD.n11078 PAD.n10757 2.2505
R38378 PAD.n11080 PAD.n11079 2.2505
R38379 PAD.n10749 PAD.n10747 2.2505
R38380 PAD.n11087 PAD.n11086 2.2505
R38381 PAD.n11086 PAD.n11085 2.2505
R38382 PAD.n11083 PAD.n10749 2.2505
R38383 PAD.n11081 PAD.n11080 2.2505
R38384 PAD.n11073 PAD.n10757 2.2505
R38385 PAD.n11076 PAD.n11075 2.2505
R38386 PAD.n11071 PAD.n10759 2.2505
R38387 PAD.n11069 PAD.n11068 2.2505
R38388 PAD.n11061 PAD.n10761 2.2505
R38389 PAD.n11064 PAD.n11063 2.2505
R38390 PAD.n11059 PAD.n10763 2.2505
R38391 PAD.n11057 PAD.n11056 2.2505
R38392 PAD.n11049 PAD.n10765 2.2505
R38393 PAD.n11052 PAD.n11051 2.2505
R38394 PAD.n11047 PAD.n10767 2.2505
R38395 PAD.n11045 PAD.n11044 2.2505
R38396 PAD.n11037 PAD.n10769 2.2505
R38397 PAD.n11040 PAD.n11039 2.2505
R38398 PAD.n11035 PAD.n10771 2.2505
R38399 PAD.n11033 PAD.n11032 2.2505
R38400 PAD.n11025 PAD.n10773 2.2505
R38401 PAD.n11028 PAD.n11027 2.2505
R38402 PAD.n11023 PAD.n10775 2.2505
R38403 PAD.n11021 PAD.n11020 2.2505
R38404 PAD.n11013 PAD.n10777 2.2505
R38405 PAD.n11016 PAD.n11015 2.2505
R38406 PAD.n11011 PAD.n10779 2.2505
R38407 PAD.n11009 PAD.n11008 2.2505
R38408 PAD.n11001 PAD.n10781 2.2505
R38409 PAD.n11004 PAD.n11003 2.2505
R38410 PAD.n10999 PAD.n10783 2.2505
R38411 PAD.n10997 PAD.n10996 2.2505
R38412 PAD.n10989 PAD.n10785 2.2505
R38413 PAD.n10992 PAD.n10991 2.2505
R38414 PAD.n10987 PAD.n10787 2.2505
R38415 PAD.n10985 PAD.n10984 2.2505
R38416 PAD.n10977 PAD.n10789 2.2505
R38417 PAD.n10980 PAD.n10979 2.2505
R38418 PAD.n10975 PAD.n10791 2.2505
R38419 PAD.n10973 PAD.n10972 2.2505
R38420 PAD.n10965 PAD.n10793 2.2505
R38421 PAD.n10968 PAD.n10967 2.2505
R38422 PAD.n10963 PAD.n10795 2.2505
R38423 PAD.n10961 PAD.n10960 2.2505
R38424 PAD.n10953 PAD.n10797 2.2505
R38425 PAD.n10956 PAD.n10955 2.2505
R38426 PAD.n10951 PAD.n10799 2.2505
R38427 PAD.n10949 PAD.n10948 2.2505
R38428 PAD.n10941 PAD.n10801 2.2505
R38429 PAD.n10944 PAD.n10943 2.2505
R38430 PAD.n10939 PAD.n10803 2.2505
R38431 PAD.n10937 PAD.n10936 2.2505
R38432 PAD.n10929 PAD.n10805 2.2505
R38433 PAD.n10932 PAD.n10931 2.2505
R38434 PAD.n10927 PAD.n10807 2.2505
R38435 PAD.n10925 PAD.n10924 2.2505
R38436 PAD.n10917 PAD.n10809 2.2505
R38437 PAD.n10920 PAD.n10919 2.2505
R38438 PAD.n10915 PAD.n10811 2.2505
R38439 PAD.n10913 PAD.n10912 2.2505
R38440 PAD.n10905 PAD.n10813 2.2505
R38441 PAD.n10908 PAD.n10907 2.2505
R38442 PAD.n10903 PAD.n10815 2.2505
R38443 PAD.n10901 PAD.n10900 2.2505
R38444 PAD.n10893 PAD.n10817 2.2505
R38445 PAD.n10896 PAD.n10895 2.2505
R38446 PAD.n10891 PAD.n10819 2.2505
R38447 PAD.n10889 PAD.n10888 2.2505
R38448 PAD.n10881 PAD.n10821 2.2505
R38449 PAD.n10884 PAD.n10883 2.2505
R38450 PAD.n10879 PAD.n10823 2.2505
R38451 PAD.n10877 PAD.n10876 2.2505
R38452 PAD.n10869 PAD.n10825 2.2505
R38453 PAD.n10872 PAD.n10871 2.2505
R38454 PAD.n10867 PAD.n10827 2.2505
R38455 PAD.n10865 PAD.n10864 2.2505
R38456 PAD.n10857 PAD.n10829 2.2505
R38457 PAD.n10860 PAD.n10859 2.2505
R38458 PAD.n10855 PAD.n10831 2.2505
R38459 PAD.n10853 PAD.n10852 2.2505
R38460 PAD.n10845 PAD.n10833 2.2505
R38461 PAD.n10848 PAD.n10847 2.2505
R38462 PAD.n10843 PAD.n10835 2.2505
R38463 PAD.n10841 PAD.n10840 2.2505
R38464 PAD.n10838 PAD.n10837 2.2505
R38465 PAD.n6382 PAD.n6381 2.2505
R38466 PAD.n5977 PAD.n5975 2.2505
R38467 PAD.n5973 PAD.n5952 2.2505
R38468 PAD.n6685 PAD.n6684 2.2505
R38469 PAD.n5560 PAD.n5559 2.2505
R38470 PAD.n6702 PAD.n6701 2.2505
R38471 PAD.n7800 PAD.n7799 2.2505
R38472 PAD.n5556 PAD.n5554 2.2505
R38473 PAD.n7794 PAD.n7793 2.2505
R38474 PAD.n6710 PAD.n6708 2.2505
R38475 PAD.n7152 PAD.n7149 2.2505
R38476 PAD.n7529 PAD.n7527 2.2505
R38477 PAD.n7151 PAD.n7150 2.2505
R38478 PAD.n7523 PAD.n7522 2.2505
R38479 PAD.n7205 PAD.n7204 2.2505
R38480 PAD.n5203 PAD.n5202 2.2505
R38481 PAD.n7822 PAD.n7821 2.2505
R38482 PAD.n7827 PAD.n7826 2.2505
R38483 PAD.n5189 PAD.n5188 2.2505
R38484 PAD.n8177 PAD.n8176 2.2505
R38485 PAD.n8182 PAD.n8181 2.2505
R38486 PAD.n4838 PAD.n4837 2.2505
R38487 PAD.n8197 PAD.n8196 2.2505
R38488 PAD.n8201 PAD.n4833 2.2505
R38489 PAD.n8203 PAD.n8202 2.2505
R38490 PAD.n8207 PAD.n8206 2.2505
R38491 PAD.n4672 PAD.n4671 2.2505
R38492 PAD.n8412 PAD.n8411 2.2505
R38493 PAD.n8418 PAD.n8417 2.2505
R38494 PAD.n4318 PAD.n4317 2.2505
R38495 PAD.n8433 PAD.n8432 2.2505
R38496 PAD.n8435 PAD.n3976 2.2505
R38497 PAD.n8455 PAD.n3975 2.2505
R38498 PAD.n8457 PAD.n8456 2.2505
R38499 PAD.n8459 PAD.n3632 2.2505
R38500 PAD.n8480 PAD.n3630 2.2505
R38501 PAD.n8482 PAD.n8481 2.2505
R38502 PAD.n3286 PAD.n3285 2.2505
R38503 PAD.n8505 PAD.n8504 2.2505
R38504 PAD.n8508 PAD.n8507 2.2505
R38505 PAD.n2902 PAD.n2900 2.2505
R38506 PAD.n8824 PAD.n8823 2.2505
R38507 PAD.n2896 PAD.n2893 2.2505
R38508 PAD.n8830 PAD.n8829 2.2505
R38509 PAD.n2897 PAD.n2895 2.2505
R38510 PAD.n9131 PAD.n9130 2.2505
R38511 PAD.n2493 PAD.n2492 2.2505
R38512 PAD.n9154 PAD.n9153 2.2505
R38513 PAD.n9159 PAD.n9158 2.2505
R38514 PAD.n2145 PAD.n2144 2.2505
R38515 PAD.n9178 PAD.n9177 2.2505
R38516 PAD.n9183 PAD.n9182 2.2505
R38517 PAD.n2044 PAD.n2042 2.2505
R38518 PAD.n9448 PAD.n9447 2.2505
R38519 PAD.n2039 PAD.n2038 2.2505
R38520 PAD.n9454 PAD.n9453 2.2505
R38521 PAD.n9715 PAD.n9714 2.2505
R38522 PAD.n1938 PAD.n1937 2.2505
R38523 PAD.n9720 PAD.n9719 2.2505
R38524 PAD.n9735 PAD.n9734 2.2505
R38525 PAD.n1588 PAD.n1587 2.2505
R38526 PAD.n9740 PAD.n9739 2.2505
R38527 PAD.n10001 PAD.n10000 2.2505
R38528 PAD.n1485 PAD.n1484 2.2505
R38529 PAD.n10006 PAD.n10005 2.2505
R38530 PAD.n10019 PAD.n10018 2.2505
R38531 PAD.n1135 PAD.n1133 2.2505
R38532 PAD.n10360 PAD.n10359 2.2505
R38533 PAD.n1117 PAD.n1116 2.2505
R38534 PAD.n10376 PAD.n10375 2.2505
R38535 PAD.n10379 PAD.n10378 2.2505
R38536 PAD.n775 PAD.n774 2.2505
R38537 PAD.n10400 PAD.n10399 2.2505
R38538 PAD.n10406 PAD.n10405 2.2505
R38539 PAD.n424 PAD.n423 2.2505
R38540 PAD.n10704 PAD.n10703 2.2505
R38541 PAD.n10707 PAD.n10706 2.2505
R38542 PAD.n30 PAD.n28 2.2505
R38543 PAD.n10730 PAD.n10729 2.2505
R38544 PAD.n24 PAD.n22 2.2505
R38545 PAD.n11531 PAD.n11530 2.2505
R38546 PAD.n25 PAD.n23 2.2505
R38547 PAD.n11525 PAD.n11524 2.2505
R38548 PAD.n10739 PAD.n10737 2.2505
R38549 PAD.n11503 PAD.n11502 2.2505
R38550 PAD.n6691 PAD.n6690 2.2505
R38551 PAD.n5905 PAD.n5900 2.2505
R38552 PAD.n6498 PAD.n6497 2.2505
R38553 PAD.n6496 PAD.n6495 2.2505
R38554 PAD.n6503 PAD.n6502 2.2505
R38555 PAD.n6505 PAD.n6504 2.2505
R38556 PAD.n6507 PAD.n6506 2.2505
R38557 PAD.n6493 PAD.n6492 2.2505
R38558 PAD.n6512 PAD.n6511 2.2505
R38559 PAD.n6514 PAD.n6513 2.2505
R38560 PAD.n6516 PAD.n6515 2.2505
R38561 PAD.n6490 PAD.n6489 2.2505
R38562 PAD.n6521 PAD.n6520 2.2505
R38563 PAD.n6523 PAD.n6522 2.2505
R38564 PAD.n6525 PAD.n6524 2.2505
R38565 PAD.n6487 PAD.n6486 2.2505
R38566 PAD.n6530 PAD.n6529 2.2505
R38567 PAD.n6532 PAD.n6531 2.2505
R38568 PAD.n6534 PAD.n6533 2.2505
R38569 PAD.n6484 PAD.n6483 2.2505
R38570 PAD.n6539 PAD.n6538 2.2505
R38571 PAD.n6541 PAD.n6540 2.2505
R38572 PAD.n6543 PAD.n6542 2.2505
R38573 PAD.n6481 PAD.n6480 2.2505
R38574 PAD.n6548 PAD.n6547 2.2505
R38575 PAD.n6550 PAD.n6549 2.2505
R38576 PAD.n6552 PAD.n6551 2.2505
R38577 PAD.n6478 PAD.n6477 2.2505
R38578 PAD.n6557 PAD.n6556 2.2505
R38579 PAD.n6559 PAD.n6558 2.2505
R38580 PAD.n6561 PAD.n6560 2.2505
R38581 PAD.n6475 PAD.n6474 2.2505
R38582 PAD.n6566 PAD.n6565 2.2505
R38583 PAD.n6568 PAD.n6567 2.2505
R38584 PAD.n6570 PAD.n6569 2.2505
R38585 PAD.n6472 PAD.n6471 2.2505
R38586 PAD.n6575 PAD.n6574 2.2505
R38587 PAD.n6577 PAD.n6576 2.2505
R38588 PAD.n6579 PAD.n6578 2.2505
R38589 PAD.n6469 PAD.n6468 2.2505
R38590 PAD.n6584 PAD.n6583 2.2505
R38591 PAD.n6586 PAD.n6585 2.2505
R38592 PAD.n6588 PAD.n6587 2.2505
R38593 PAD.n6466 PAD.n6465 2.2505
R38594 PAD.n6593 PAD.n6592 2.2505
R38595 PAD.n6595 PAD.n6594 2.2505
R38596 PAD.n6597 PAD.n6596 2.2505
R38597 PAD.n6463 PAD.n6462 2.2505
R38598 PAD.n6602 PAD.n6601 2.2505
R38599 PAD.n6604 PAD.n6603 2.2505
R38600 PAD.n6606 PAD.n6605 2.2505
R38601 PAD.n6460 PAD.n6459 2.2505
R38602 PAD.n6611 PAD.n6610 2.2505
R38603 PAD.n6613 PAD.n6612 2.2505
R38604 PAD.n6615 PAD.n6614 2.2505
R38605 PAD.n6457 PAD.n6456 2.2505
R38606 PAD.n6620 PAD.n6619 2.2505
R38607 PAD.n6622 PAD.n6621 2.2505
R38608 PAD.n6624 PAD.n6623 2.2505
R38609 PAD.n6454 PAD.n6453 2.2505
R38610 PAD.n6629 PAD.n6628 2.2505
R38611 PAD.n6631 PAD.n6630 2.2505
R38612 PAD.n6633 PAD.n6632 2.2505
R38613 PAD.n6451 PAD.n6450 2.2505
R38614 PAD.n6638 PAD.n6637 2.2505
R38615 PAD.n6640 PAD.n6639 2.2505
R38616 PAD.n6642 PAD.n6641 2.2505
R38617 PAD.n6448 PAD.n6447 2.2505
R38618 PAD.n6647 PAD.n6646 2.2505
R38619 PAD.n6649 PAD.n6648 2.2505
R38620 PAD.n6651 PAD.n6650 2.2505
R38621 PAD.n6445 PAD.n6444 2.2505
R38622 PAD.n6656 PAD.n6655 2.2505
R38623 PAD.n6658 PAD.n6657 2.2505
R38624 PAD.n6660 PAD.n6659 2.2505
R38625 PAD.n6442 PAD.n6441 2.2505
R38626 PAD.n6665 PAD.n6664 2.2505
R38627 PAD.n6667 PAD.n6666 2.2505
R38628 PAD.n6669 PAD.n6668 2.2505
R38629 PAD.n6438 PAD.n6437 2.2505
R38630 PAD.n6676 PAD.n6675 2.2505
R38631 PAD.n6439 PAD.n6436 2.2505
R38632 PAD.n5950 PAD.n5949 2.2505
R38633 PAD.n6688 PAD.n6687 2.2505
R38634 PAD.n6383 PAD.n6382 2.2505
R38635 PAD.n5975 PAD.n5974 2.2505
R38636 PAD.n5973 PAD.n5904 2.2505
R38637 PAD.n6684 PAD.n6683 2.2505
R38638 PAD.n6680 PAD.n5560 2.2505
R38639 PAD.n6701 PAD.n6700 2.2505
R38640 PAD.n7801 PAD.n7800 2.2505
R38641 PAD.n6711 PAD.n5554 2.2505
R38642 PAD.n7793 PAD.n7792 2.2505
R38643 PAD.n7059 PAD.n6710 2.2505
R38644 PAD.n7149 PAD.n7061 2.2505
R38645 PAD.n7529 PAD.n7528 2.2505
R38646 PAD.n7215 PAD.n7150 2.2505
R38647 PAD.n7522 PAD.n7521 2.2505
R38648 PAD.n7206 PAD.n7205 2.2505
R38649 PAD.n7222 PAD.n5203 2.2505
R38650 PAD.n7821 PAD.n7820 2.2505
R38651 PAD.n7828 PAD.n7827 2.2505
R38652 PAD.n8164 PAD.n5189 2.2505
R38653 PAD.n8176 PAD.n8175 2.2505
R38654 PAD.n8183 PAD.n8182 2.2505
R38655 PAD.n8185 PAD.n4838 2.2505
R38656 PAD.n8196 PAD.n8195 2.2505
R38657 PAD.n4842 PAD.n4833 2.2505
R38658 PAD.n8203 PAD.n4682 2.2505
R38659 PAD.n8206 PAD.n8205 2.2505
R38660 PAD.n8408 PAD.n4672 2.2505
R38661 PAD.n8411 PAD.n8410 2.2505
R38662 PAD.n8419 PAD.n8418 2.2505
R38663 PAD.n4319 PAD.n4318 2.2505
R38664 PAD.n8432 PAD.n8431 2.2505
R38665 PAD.n3983 PAD.n3976 2.2505
R38666 PAD.n8455 PAD.n8454 2.2505
R38667 PAD.n8456 PAD.n3641 2.2505
R38668 PAD.n3684 PAD.n3632 2.2505
R38669 PAD.n8480 PAD.n8479 2.2505
R38670 PAD.n8481 PAD.n3296 2.2505
R38671 PAD.n3339 PAD.n3286 2.2505
R38672 PAD.n8504 PAD.n8503 2.2505
R38673 PAD.n8507 PAD.n2952 2.2505
R38674 PAD.n8518 PAD.n2902 2.2505
R38675 PAD.n8823 PAD.n8822 2.2505
R38676 PAD.n2946 PAD.n2893 2.2505
R38677 PAD.n8831 PAD.n8830 2.2505
R38678 PAD.n2895 PAD.n2894 2.2505
R38679 PAD.n9130 PAD.n9129 2.2505
R38680 PAD.n9142 PAD.n2493 2.2505
R38681 PAD.n9153 PAD.n9152 2.2505
R38682 PAD.n9160 PAD.n9159 2.2505
R38683 PAD.n9162 PAD.n2145 2.2505
R38684 PAD.n9177 PAD.n9176 2.2505
R38685 PAD.n9184 PAD.n9183 2.2505
R38686 PAD.n9186 PAD.n2044 2.2505
R38687 PAD.n9447 PAD.n9446 2.2505
R38688 PAD.n2038 PAD.n2037 2.2505
R38689 PAD.n9455 PAD.n9454 2.2505
R38690 PAD.n9714 PAD.n9713 2.2505
R38691 PAD.n1985 PAD.n1937 2.2505
R38692 PAD.n9721 PAD.n9720 2.2505
R38693 PAD.n9734 PAD.n9733 2.2505
R38694 PAD.n1587 PAD.n1586 2.2505
R38695 PAD.n9741 PAD.n9740 2.2505
R38696 PAD.n10000 PAD.n9999 2.2505
R38697 PAD.n1533 PAD.n1484 2.2505
R38698 PAD.n10007 PAD.n10006 2.2505
R38699 PAD.n10018 PAD.n10017 2.2505
R38700 PAD.n1142 PAD.n1133 2.2505
R38701 PAD.n10361 PAD.n10360 2.2505
R38702 PAD.n1118 PAD.n1117 2.2505
R38703 PAD.n10375 PAD.n10374 2.2505
R38704 PAD.n10378 PAD.n782 2.2505
R38705 PAD.n825 PAD.n775 2.2505
R38706 PAD.n10399 PAD.n10398 2.2505
R38707 PAD.n10407 PAD.n10406 2.2505
R38708 PAD.n425 PAD.n424 2.2505
R38709 PAD.n10703 PAD.n10702 2.2505
R38710 PAD.n10706 PAD.n373 2.2505
R38711 PAD.n10718 PAD.n30 2.2505
R38712 PAD.n10729 PAD.n10728 2.2505
R38713 PAD.n22 PAD.n20 2.2505
R38714 PAD.n11532 PAD.n11531 2.2505
R38715 PAD.n10754 PAD.n23 2.2505
R38716 PAD.n11524 PAD.n11523 2.2505
R38717 PAD.n10741 PAD.n10739 2.2505
R38718 PAD.n11502 PAD.n11501 2.2505
R38719 PAD.n11155 PAD.n11105 2.24752
R38720 PAD.n6031 PAD.n5980 2.24752
R38721 PAD.n11157 PAD.n11100 2.24752
R38722 PAD.n11302 PAD.n11254 2.24752
R38723 PAD.n11159 PAD.n11100 2.24752
R38724 PAD.n11302 PAD.n11255 2.24752
R38725 PAD.n11161 PAD.n11100 2.24752
R38726 PAD.n11302 PAD.n11256 2.24752
R38727 PAD.n11163 PAD.n11100 2.24752
R38728 PAD.n11302 PAD.n11257 2.24752
R38729 PAD.n11165 PAD.n11100 2.24752
R38730 PAD.n11302 PAD.n11258 2.24752
R38731 PAD.n11167 PAD.n11100 2.24752
R38732 PAD.n11302 PAD.n11259 2.24752
R38733 PAD.n11169 PAD.n11100 2.24752
R38734 PAD.n11302 PAD.n11260 2.24752
R38735 PAD.n11171 PAD.n11100 2.24752
R38736 PAD.n11302 PAD.n11261 2.24752
R38737 PAD.n11173 PAD.n11100 2.24752
R38738 PAD.n11302 PAD.n11262 2.24752
R38739 PAD.n11175 PAD.n11100 2.24752
R38740 PAD.n11302 PAD.n11263 2.24752
R38741 PAD.n11177 PAD.n11100 2.24752
R38742 PAD.n11302 PAD.n11264 2.24752
R38743 PAD.n11179 PAD.n11100 2.24752
R38744 PAD.n11302 PAD.n11265 2.24752
R38745 PAD.n11181 PAD.n11100 2.24752
R38746 PAD.n11302 PAD.n11266 2.24752
R38747 PAD.n11183 PAD.n11100 2.24752
R38748 PAD.n11302 PAD.n11267 2.24752
R38749 PAD.n11185 PAD.n11100 2.24752
R38750 PAD.n11302 PAD.n11268 2.24752
R38751 PAD.n11187 PAD.n11100 2.24752
R38752 PAD.n11302 PAD.n11269 2.24752
R38753 PAD.n11189 PAD.n11100 2.24752
R38754 PAD.n11302 PAD.n11270 2.24752
R38755 PAD.n11191 PAD.n11100 2.24752
R38756 PAD.n11302 PAD.n11271 2.24752
R38757 PAD.n11193 PAD.n11100 2.24752
R38758 PAD.n11302 PAD.n11272 2.24752
R38759 PAD.n11195 PAD.n11100 2.24752
R38760 PAD.n11302 PAD.n11273 2.24752
R38761 PAD.n11197 PAD.n11100 2.24752
R38762 PAD.n11302 PAD.n11274 2.24752
R38763 PAD.n11199 PAD.n11100 2.24752
R38764 PAD.n11302 PAD.n11275 2.24752
R38765 PAD.n11201 PAD.n11100 2.24752
R38766 PAD.n11302 PAD.n11276 2.24752
R38767 PAD.n11203 PAD.n11100 2.24752
R38768 PAD.n11302 PAD.n11277 2.24752
R38769 PAD.n11205 PAD.n11100 2.24752
R38770 PAD.n11302 PAD.n11278 2.24752
R38771 PAD.n11207 PAD.n11100 2.24752
R38772 PAD.n11302 PAD.n11279 2.24752
R38773 PAD.n11209 PAD.n11100 2.24752
R38774 PAD.n11302 PAD.n11280 2.24752
R38775 PAD.n11211 PAD.n11100 2.24752
R38776 PAD.n11302 PAD.n11281 2.24752
R38777 PAD.n11213 PAD.n11100 2.24752
R38778 PAD.n11302 PAD.n11282 2.24752
R38779 PAD.n11215 PAD.n11100 2.24752
R38780 PAD.n11302 PAD.n11283 2.24752
R38781 PAD.n11217 PAD.n11100 2.24752
R38782 PAD.n11302 PAD.n11284 2.24752
R38783 PAD.n11219 PAD.n11100 2.24752
R38784 PAD.n11302 PAD.n11285 2.24752
R38785 PAD.n11221 PAD.n11100 2.24752
R38786 PAD.n11302 PAD.n11286 2.24752
R38787 PAD.n11223 PAD.n11100 2.24752
R38788 PAD.n11302 PAD.n11287 2.24752
R38789 PAD.n11225 PAD.n11100 2.24752
R38790 PAD.n11302 PAD.n11288 2.24752
R38791 PAD.n11227 PAD.n11100 2.24752
R38792 PAD.n11302 PAD.n11289 2.24752
R38793 PAD.n11229 PAD.n11100 2.24752
R38794 PAD.n11302 PAD.n11290 2.24752
R38795 PAD.n11231 PAD.n11100 2.24752
R38796 PAD.n11302 PAD.n11291 2.24752
R38797 PAD.n11233 PAD.n11100 2.24752
R38798 PAD.n11302 PAD.n11292 2.24752
R38799 PAD.n11235 PAD.n11100 2.24752
R38800 PAD.n11302 PAD.n11293 2.24752
R38801 PAD.n11237 PAD.n11100 2.24752
R38802 PAD.n11302 PAD.n11294 2.24752
R38803 PAD.n11239 PAD.n11100 2.24752
R38804 PAD.n11302 PAD.n11295 2.24752
R38805 PAD.n11241 PAD.n11100 2.24752
R38806 PAD.n11302 PAD.n11296 2.24752
R38807 PAD.n11243 PAD.n11100 2.24752
R38808 PAD.n11302 PAD.n11297 2.24752
R38809 PAD.n11245 PAD.n11100 2.24752
R38810 PAD.n11302 PAD.n11298 2.24752
R38811 PAD.n11247 PAD.n11100 2.24752
R38812 PAD.n11302 PAD.n11299 2.24752
R38813 PAD.n11249 PAD.n11100 2.24752
R38814 PAD.n11302 PAD.n11300 2.24752
R38815 PAD.n11251 PAD.n11100 2.24752
R38816 PAD.n11302 PAD.n11301 2.24752
R38817 PAD.n5966 PAD.n5961 2.24752
R38818 PAD.n11510 PAD.n11095 2.24752
R38819 PAD.n6384 PAD.n5966 2.24752
R38820 PAD.n11511 PAD.n11510 2.24752
R38821 PAD.n6033 PAD.n5982 2.24752
R38822 PAD.n6035 PAD.n5980 2.24752
R38823 PAD.n6036 PAD.n5982 2.24752
R38824 PAD.n6038 PAD.n5980 2.24752
R38825 PAD.n6039 PAD.n5982 2.24752
R38826 PAD.n6041 PAD.n5980 2.24752
R38827 PAD.n6042 PAD.n5982 2.24752
R38828 PAD.n6044 PAD.n5980 2.24752
R38829 PAD.n6045 PAD.n5982 2.24752
R38830 PAD.n6047 PAD.n5980 2.24752
R38831 PAD.n6048 PAD.n5982 2.24752
R38832 PAD.n6050 PAD.n5980 2.24752
R38833 PAD.n6051 PAD.n5982 2.24752
R38834 PAD.n6053 PAD.n5980 2.24752
R38835 PAD.n6054 PAD.n5982 2.24752
R38836 PAD.n6056 PAD.n5980 2.24752
R38837 PAD.n6057 PAD.n5982 2.24752
R38838 PAD.n6059 PAD.n5980 2.24752
R38839 PAD.n6060 PAD.n5982 2.24752
R38840 PAD.n6062 PAD.n5980 2.24752
R38841 PAD.n6063 PAD.n5982 2.24752
R38842 PAD.n6065 PAD.n5980 2.24752
R38843 PAD.n6066 PAD.n5982 2.24752
R38844 PAD.n6068 PAD.n5980 2.24752
R38845 PAD.n6069 PAD.n5982 2.24752
R38846 PAD.n6071 PAD.n5980 2.24752
R38847 PAD.n6072 PAD.n5982 2.24752
R38848 PAD.n6074 PAD.n5980 2.24752
R38849 PAD.n6075 PAD.n5982 2.24752
R38850 PAD.n6077 PAD.n5980 2.24752
R38851 PAD.n6078 PAD.n5982 2.24752
R38852 PAD.n6080 PAD.n5980 2.24752
R38853 PAD.n6081 PAD.n5982 2.24752
R38854 PAD.n6083 PAD.n5980 2.24752
R38855 PAD.n6084 PAD.n5982 2.24752
R38856 PAD.n6086 PAD.n5980 2.24752
R38857 PAD.n6087 PAD.n5982 2.24752
R38858 PAD.n6089 PAD.n5980 2.24752
R38859 PAD.n6090 PAD.n5982 2.24752
R38860 PAD.n6092 PAD.n5980 2.24752
R38861 PAD.n6093 PAD.n5982 2.24752
R38862 PAD.n6095 PAD.n5980 2.24752
R38863 PAD.n6096 PAD.n5982 2.24752
R38864 PAD.n6098 PAD.n5980 2.24752
R38865 PAD.n6099 PAD.n5982 2.24752
R38866 PAD.n6101 PAD.n5980 2.24752
R38867 PAD.n6102 PAD.n5982 2.24752
R38868 PAD.n6104 PAD.n5980 2.24752
R38869 PAD.n6105 PAD.n5982 2.24752
R38870 PAD.n6107 PAD.n5980 2.24752
R38871 PAD.n6108 PAD.n5982 2.24752
R38872 PAD.n6110 PAD.n5980 2.24752
R38873 PAD.n6111 PAD.n5982 2.24752
R38874 PAD.n6113 PAD.n5980 2.24752
R38875 PAD.n6114 PAD.n5982 2.24752
R38876 PAD.n6116 PAD.n5980 2.24752
R38877 PAD.n6117 PAD.n5982 2.24752
R38878 PAD.n6119 PAD.n5980 2.24752
R38879 PAD.n6120 PAD.n5982 2.24752
R38880 PAD.n6122 PAD.n5980 2.24752
R38881 PAD.n6123 PAD.n5982 2.24752
R38882 PAD.n6125 PAD.n5980 2.24752
R38883 PAD.n6126 PAD.n5982 2.24752
R38884 PAD.n6128 PAD.n5980 2.24752
R38885 PAD.n6129 PAD.n5982 2.24752
R38886 PAD.n6131 PAD.n5980 2.24752
R38887 PAD.n6132 PAD.n5982 2.24752
R38888 PAD.n6134 PAD.n5980 2.24752
R38889 PAD.n6135 PAD.n5982 2.24752
R38890 PAD.n6137 PAD.n5980 2.24752
R38891 PAD.n6138 PAD.n5982 2.24752
R38892 PAD.n6140 PAD.n5980 2.24752
R38893 PAD.n6141 PAD.n5982 2.24752
R38894 PAD.n6143 PAD.n5980 2.24752
R38895 PAD.n6144 PAD.n5982 2.24752
R38896 PAD.n6146 PAD.n5980 2.24752
R38897 PAD.n6147 PAD.n5982 2.24752
R38898 PAD.n6149 PAD.n5980 2.24752
R38899 PAD.n6150 PAD.n5982 2.24752
R38900 PAD.n6152 PAD.n5980 2.24752
R38901 PAD.n6153 PAD.n5982 2.24752
R38902 PAD.n6155 PAD.n5980 2.24752
R38903 PAD.n6156 PAD.n5982 2.24752
R38904 PAD.n6158 PAD.n5980 2.24752
R38905 PAD.n6159 PAD.n5982 2.24752
R38906 PAD.n6161 PAD.n5980 2.24752
R38907 PAD.n6162 PAD.n5982 2.24752
R38908 PAD.n6164 PAD.n5980 2.24752
R38909 PAD.n6165 PAD.n5982 2.24752
R38910 PAD.n6167 PAD.n5980 2.24752
R38911 PAD.n6168 PAD.n5982 2.24752
R38912 PAD.n6170 PAD.n5980 2.24752
R38913 PAD.n6171 PAD.n5982 2.24752
R38914 PAD.n6173 PAD.n5980 2.24752
R38915 PAD.n6174 PAD.n5982 2.24752
R38916 PAD.n6176 PAD.n5982 2.24752
R38917 PAD.n11084 PAD.n10755 2.24164
R38918 PAD.n11082 PAD.n21 2.24164
R38919 PAD.n10756 PAD.n10755 2.24164
R38920 PAD.n11074 PAD.n21 2.24164
R38921 PAD.n11072 PAD.n10755 2.24164
R38922 PAD.n11070 PAD.n21 2.24164
R38923 PAD.n10760 PAD.n10755 2.24164
R38924 PAD.n11062 PAD.n21 2.24164
R38925 PAD.n11060 PAD.n10755 2.24164
R38926 PAD.n11058 PAD.n21 2.24164
R38927 PAD.n10764 PAD.n10755 2.24164
R38928 PAD.n11050 PAD.n21 2.24164
R38929 PAD.n11048 PAD.n10755 2.24164
R38930 PAD.n11046 PAD.n21 2.24164
R38931 PAD.n10768 PAD.n10755 2.24164
R38932 PAD.n11038 PAD.n21 2.24164
R38933 PAD.n11036 PAD.n10755 2.24164
R38934 PAD.n11034 PAD.n21 2.24164
R38935 PAD.n10772 PAD.n10755 2.24164
R38936 PAD.n11026 PAD.n21 2.24164
R38937 PAD.n11024 PAD.n10755 2.24164
R38938 PAD.n11022 PAD.n21 2.24164
R38939 PAD.n10776 PAD.n10755 2.24164
R38940 PAD.n11014 PAD.n21 2.24164
R38941 PAD.n11012 PAD.n10755 2.24164
R38942 PAD.n11010 PAD.n21 2.24164
R38943 PAD.n10780 PAD.n10755 2.24164
R38944 PAD.n11002 PAD.n21 2.24164
R38945 PAD.n11000 PAD.n10755 2.24164
R38946 PAD.n10998 PAD.n21 2.24164
R38947 PAD.n10784 PAD.n10755 2.24164
R38948 PAD.n10990 PAD.n21 2.24164
R38949 PAD.n10988 PAD.n10755 2.24164
R38950 PAD.n10986 PAD.n21 2.24164
R38951 PAD.n10788 PAD.n10755 2.24164
R38952 PAD.n10978 PAD.n21 2.24164
R38953 PAD.n10976 PAD.n10755 2.24164
R38954 PAD.n10974 PAD.n21 2.24164
R38955 PAD.n10792 PAD.n10755 2.24164
R38956 PAD.n10966 PAD.n21 2.24164
R38957 PAD.n10964 PAD.n10755 2.24164
R38958 PAD.n10962 PAD.n21 2.24164
R38959 PAD.n10796 PAD.n10755 2.24164
R38960 PAD.n10954 PAD.n21 2.24164
R38961 PAD.n10952 PAD.n10755 2.24164
R38962 PAD.n10950 PAD.n21 2.24164
R38963 PAD.n10800 PAD.n10755 2.24164
R38964 PAD.n10942 PAD.n21 2.24164
R38965 PAD.n10940 PAD.n10755 2.24164
R38966 PAD.n10938 PAD.n21 2.24164
R38967 PAD.n10804 PAD.n10755 2.24164
R38968 PAD.n10930 PAD.n21 2.24164
R38969 PAD.n10928 PAD.n10755 2.24164
R38970 PAD.n10926 PAD.n21 2.24164
R38971 PAD.n10808 PAD.n10755 2.24164
R38972 PAD.n10918 PAD.n21 2.24164
R38973 PAD.n10916 PAD.n10755 2.24164
R38974 PAD.n10914 PAD.n21 2.24164
R38975 PAD.n10812 PAD.n10755 2.24164
R38976 PAD.n10906 PAD.n21 2.24164
R38977 PAD.n10904 PAD.n10755 2.24164
R38978 PAD.n10902 PAD.n21 2.24164
R38979 PAD.n10816 PAD.n10755 2.24164
R38980 PAD.n10894 PAD.n21 2.24164
R38981 PAD.n10892 PAD.n10755 2.24164
R38982 PAD.n10890 PAD.n21 2.24164
R38983 PAD.n10820 PAD.n10755 2.24164
R38984 PAD.n10882 PAD.n21 2.24164
R38985 PAD.n10880 PAD.n10755 2.24164
R38986 PAD.n10878 PAD.n21 2.24164
R38987 PAD.n10824 PAD.n10755 2.24164
R38988 PAD.n10870 PAD.n21 2.24164
R38989 PAD.n10868 PAD.n10755 2.24164
R38990 PAD.n10866 PAD.n21 2.24164
R38991 PAD.n10828 PAD.n10755 2.24164
R38992 PAD.n10858 PAD.n21 2.24164
R38993 PAD.n10856 PAD.n10755 2.24164
R38994 PAD.n10854 PAD.n21 2.24164
R38995 PAD.n10832 PAD.n10755 2.24164
R38996 PAD.n10846 PAD.n21 2.24164
R38997 PAD.n10844 PAD.n10755 2.24164
R38998 PAD.n10842 PAD.n21 2.24164
R38999 PAD.n10836 PAD.n10755 2.24164
R39000 PAD.n116 PAD.n32 2.24164
R39001 PAD.n367 PAD.n73 2.24164
R39002 PAD.n125 PAD.n32 2.24164
R39003 PAD.n367 PAD.n72 2.24164
R39004 PAD.n129 PAD.n32 2.24164
R39005 PAD.n367 PAD.n71 2.24164
R39006 PAD.n137 PAD.n32 2.24164
R39007 PAD.n367 PAD.n70 2.24164
R39008 PAD.n141 PAD.n32 2.24164
R39009 PAD.n367 PAD.n69 2.24164
R39010 PAD.n149 PAD.n32 2.24164
R39011 PAD.n367 PAD.n68 2.24164
R39012 PAD.n153 PAD.n32 2.24164
R39013 PAD.n367 PAD.n67 2.24164
R39014 PAD.n161 PAD.n32 2.24164
R39015 PAD.n367 PAD.n66 2.24164
R39016 PAD.n165 PAD.n32 2.24164
R39017 PAD.n367 PAD.n65 2.24164
R39018 PAD.n173 PAD.n32 2.24164
R39019 PAD.n367 PAD.n64 2.24164
R39020 PAD.n177 PAD.n32 2.24164
R39021 PAD.n367 PAD.n63 2.24164
R39022 PAD.n185 PAD.n32 2.24164
R39023 PAD.n367 PAD.n62 2.24164
R39024 PAD.n189 PAD.n32 2.24164
R39025 PAD.n367 PAD.n61 2.24164
R39026 PAD.n197 PAD.n32 2.24164
R39027 PAD.n367 PAD.n60 2.24164
R39028 PAD.n201 PAD.n32 2.24164
R39029 PAD.n367 PAD.n59 2.24164
R39030 PAD.n209 PAD.n32 2.24164
R39031 PAD.n367 PAD.n58 2.24164
R39032 PAD.n213 PAD.n32 2.24164
R39033 PAD.n367 PAD.n57 2.24164
R39034 PAD.n221 PAD.n32 2.24164
R39035 PAD.n367 PAD.n56 2.24164
R39036 PAD.n225 PAD.n32 2.24164
R39037 PAD.n367 PAD.n55 2.24164
R39038 PAD.n233 PAD.n32 2.24164
R39039 PAD.n367 PAD.n54 2.24164
R39040 PAD.n237 PAD.n32 2.24164
R39041 PAD.n367 PAD.n53 2.24164
R39042 PAD.n245 PAD.n32 2.24164
R39043 PAD.n367 PAD.n52 2.24164
R39044 PAD.n249 PAD.n32 2.24164
R39045 PAD.n367 PAD.n51 2.24164
R39046 PAD.n257 PAD.n32 2.24164
R39047 PAD.n367 PAD.n50 2.24164
R39048 PAD.n261 PAD.n32 2.24164
R39049 PAD.n367 PAD.n49 2.24164
R39050 PAD.n269 PAD.n32 2.24164
R39051 PAD.n367 PAD.n48 2.24164
R39052 PAD.n273 PAD.n32 2.24164
R39053 PAD.n367 PAD.n47 2.24164
R39054 PAD.n281 PAD.n32 2.24164
R39055 PAD.n367 PAD.n46 2.24164
R39056 PAD.n285 PAD.n32 2.24164
R39057 PAD.n367 PAD.n45 2.24164
R39058 PAD.n293 PAD.n32 2.24164
R39059 PAD.n367 PAD.n44 2.24164
R39060 PAD.n297 PAD.n32 2.24164
R39061 PAD.n367 PAD.n43 2.24164
R39062 PAD.n305 PAD.n32 2.24164
R39063 PAD.n367 PAD.n42 2.24164
R39064 PAD.n309 PAD.n32 2.24164
R39065 PAD.n367 PAD.n41 2.24164
R39066 PAD.n317 PAD.n32 2.24164
R39067 PAD.n367 PAD.n40 2.24164
R39068 PAD.n321 PAD.n32 2.24164
R39069 PAD.n367 PAD.n39 2.24164
R39070 PAD.n329 PAD.n32 2.24164
R39071 PAD.n367 PAD.n38 2.24164
R39072 PAD.n333 PAD.n32 2.24164
R39073 PAD.n367 PAD.n37 2.24164
R39074 PAD.n341 PAD.n32 2.24164
R39075 PAD.n367 PAD.n36 2.24164
R39076 PAD.n345 PAD.n32 2.24164
R39077 PAD.n367 PAD.n35 2.24164
R39078 PAD.n353 PAD.n32 2.24164
R39079 PAD.n367 PAD.n34 2.24164
R39080 PAD.n357 PAD.n32 2.24164
R39081 PAD.n367 PAD.n33 2.24164
R39082 PAD.n365 PAD.n32 2.24164
R39083 PAD.n10692 PAD.n419 2.24164
R39084 PAD.n10716 PAD.n414 2.24164
R39085 PAD.n10416 PAD.n419 2.24164
R39086 PAD.n10716 PAD.n413 2.24164
R39087 PAD.n10685 PAD.n419 2.24164
R39088 PAD.n10716 PAD.n412 2.24164
R39089 PAD.n10421 PAD.n419 2.24164
R39090 PAD.n10716 PAD.n411 2.24164
R39091 PAD.n10676 PAD.n419 2.24164
R39092 PAD.n10716 PAD.n410 2.24164
R39093 PAD.n10426 PAD.n419 2.24164
R39094 PAD.n10716 PAD.n409 2.24164
R39095 PAD.n10667 PAD.n419 2.24164
R39096 PAD.n10716 PAD.n408 2.24164
R39097 PAD.n10431 PAD.n419 2.24164
R39098 PAD.n10716 PAD.n407 2.24164
R39099 PAD.n10658 PAD.n419 2.24164
R39100 PAD.n10716 PAD.n406 2.24164
R39101 PAD.n10436 PAD.n419 2.24164
R39102 PAD.n10716 PAD.n405 2.24164
R39103 PAD.n10649 PAD.n419 2.24164
R39104 PAD.n10716 PAD.n404 2.24164
R39105 PAD.n10441 PAD.n419 2.24164
R39106 PAD.n10716 PAD.n403 2.24164
R39107 PAD.n10640 PAD.n419 2.24164
R39108 PAD.n10716 PAD.n402 2.24164
R39109 PAD.n10446 PAD.n419 2.24164
R39110 PAD.n10716 PAD.n401 2.24164
R39111 PAD.n10631 PAD.n419 2.24164
R39112 PAD.n10716 PAD.n400 2.24164
R39113 PAD.n10451 PAD.n419 2.24164
R39114 PAD.n10716 PAD.n399 2.24164
R39115 PAD.n10622 PAD.n419 2.24164
R39116 PAD.n10716 PAD.n398 2.24164
R39117 PAD.n10456 PAD.n419 2.24164
R39118 PAD.n10716 PAD.n397 2.24164
R39119 PAD.n10613 PAD.n419 2.24164
R39120 PAD.n10716 PAD.n396 2.24164
R39121 PAD.n10461 PAD.n419 2.24164
R39122 PAD.n10716 PAD.n395 2.24164
R39123 PAD.n10604 PAD.n419 2.24164
R39124 PAD.n10716 PAD.n394 2.24164
R39125 PAD.n10466 PAD.n419 2.24164
R39126 PAD.n10716 PAD.n393 2.24164
R39127 PAD.n10595 PAD.n419 2.24164
R39128 PAD.n10716 PAD.n392 2.24164
R39129 PAD.n10471 PAD.n419 2.24164
R39130 PAD.n10716 PAD.n391 2.24164
R39131 PAD.n10586 PAD.n419 2.24164
R39132 PAD.n10716 PAD.n390 2.24164
R39133 PAD.n10476 PAD.n419 2.24164
R39134 PAD.n10716 PAD.n389 2.24164
R39135 PAD.n10577 PAD.n419 2.24164
R39136 PAD.n10716 PAD.n388 2.24164
R39137 PAD.n10481 PAD.n419 2.24164
R39138 PAD.n10716 PAD.n387 2.24164
R39139 PAD.n10568 PAD.n419 2.24164
R39140 PAD.n10716 PAD.n386 2.24164
R39141 PAD.n10486 PAD.n419 2.24164
R39142 PAD.n10716 PAD.n385 2.24164
R39143 PAD.n10559 PAD.n419 2.24164
R39144 PAD.n10716 PAD.n384 2.24164
R39145 PAD.n10491 PAD.n419 2.24164
R39146 PAD.n10716 PAD.n383 2.24164
R39147 PAD.n10550 PAD.n419 2.24164
R39148 PAD.n10716 PAD.n382 2.24164
R39149 PAD.n10496 PAD.n419 2.24164
R39150 PAD.n10716 PAD.n381 2.24164
R39151 PAD.n10541 PAD.n419 2.24164
R39152 PAD.n10716 PAD.n380 2.24164
R39153 PAD.n10501 PAD.n419 2.24164
R39154 PAD.n10716 PAD.n379 2.24164
R39155 PAD.n10532 PAD.n419 2.24164
R39156 PAD.n10716 PAD.n378 2.24164
R39157 PAD.n10506 PAD.n419 2.24164
R39158 PAD.n10716 PAD.n377 2.24164
R39159 PAD.n10523 PAD.n419 2.24164
R39160 PAD.n10716 PAD.n376 2.24164
R39161 PAD.n10511 PAD.n419 2.24164
R39162 PAD.n10716 PAD.n375 2.24164
R39163 PAD.n10514 PAD.n419 2.24164
R39164 PAD.n10716 PAD.n374 2.24164
R39165 PAD.n10714 PAD.n419 2.24164
R39166 PAD.n524 PAD.n433 2.24164
R39167 PAD.n526 PAD.n435 2.24164
R39168 PAD.n528 PAD.n433 2.24164
R39169 PAD.n517 PAD.n435 2.24164
R39170 PAD.n536 PAD.n433 2.24164
R39171 PAD.n538 PAD.n435 2.24164
R39172 PAD.n540 PAD.n433 2.24164
R39173 PAD.n513 PAD.n435 2.24164
R39174 PAD.n548 PAD.n433 2.24164
R39175 PAD.n550 PAD.n435 2.24164
R39176 PAD.n552 PAD.n433 2.24164
R39177 PAD.n509 PAD.n435 2.24164
R39178 PAD.n560 PAD.n433 2.24164
R39179 PAD.n562 PAD.n435 2.24164
R39180 PAD.n564 PAD.n433 2.24164
R39181 PAD.n505 PAD.n435 2.24164
R39182 PAD.n572 PAD.n433 2.24164
R39183 PAD.n574 PAD.n435 2.24164
R39184 PAD.n576 PAD.n433 2.24164
R39185 PAD.n501 PAD.n435 2.24164
R39186 PAD.n584 PAD.n433 2.24164
R39187 PAD.n586 PAD.n435 2.24164
R39188 PAD.n588 PAD.n433 2.24164
R39189 PAD.n497 PAD.n435 2.24164
R39190 PAD.n596 PAD.n433 2.24164
R39191 PAD.n598 PAD.n435 2.24164
R39192 PAD.n600 PAD.n433 2.24164
R39193 PAD.n493 PAD.n435 2.24164
R39194 PAD.n608 PAD.n433 2.24164
R39195 PAD.n610 PAD.n435 2.24164
R39196 PAD.n612 PAD.n433 2.24164
R39197 PAD.n489 PAD.n435 2.24164
R39198 PAD.n620 PAD.n433 2.24164
R39199 PAD.n622 PAD.n435 2.24164
R39200 PAD.n624 PAD.n433 2.24164
R39201 PAD.n485 PAD.n435 2.24164
R39202 PAD.n632 PAD.n433 2.24164
R39203 PAD.n634 PAD.n435 2.24164
R39204 PAD.n636 PAD.n433 2.24164
R39205 PAD.n481 PAD.n435 2.24164
R39206 PAD.n644 PAD.n433 2.24164
R39207 PAD.n646 PAD.n435 2.24164
R39208 PAD.n648 PAD.n433 2.24164
R39209 PAD.n477 PAD.n435 2.24164
R39210 PAD.n656 PAD.n433 2.24164
R39211 PAD.n658 PAD.n435 2.24164
R39212 PAD.n660 PAD.n433 2.24164
R39213 PAD.n473 PAD.n435 2.24164
R39214 PAD.n668 PAD.n433 2.24164
R39215 PAD.n670 PAD.n435 2.24164
R39216 PAD.n672 PAD.n433 2.24164
R39217 PAD.n469 PAD.n435 2.24164
R39218 PAD.n680 PAD.n433 2.24164
R39219 PAD.n682 PAD.n435 2.24164
R39220 PAD.n684 PAD.n433 2.24164
R39221 PAD.n465 PAD.n435 2.24164
R39222 PAD.n692 PAD.n433 2.24164
R39223 PAD.n694 PAD.n435 2.24164
R39224 PAD.n696 PAD.n433 2.24164
R39225 PAD.n461 PAD.n435 2.24164
R39226 PAD.n704 PAD.n433 2.24164
R39227 PAD.n706 PAD.n435 2.24164
R39228 PAD.n708 PAD.n433 2.24164
R39229 PAD.n457 PAD.n435 2.24164
R39230 PAD.n716 PAD.n433 2.24164
R39231 PAD.n718 PAD.n435 2.24164
R39232 PAD.n720 PAD.n433 2.24164
R39233 PAD.n453 PAD.n435 2.24164
R39234 PAD.n728 PAD.n433 2.24164
R39235 PAD.n730 PAD.n435 2.24164
R39236 PAD.n732 PAD.n433 2.24164
R39237 PAD.n449 PAD.n435 2.24164
R39238 PAD.n740 PAD.n433 2.24164
R39239 PAD.n742 PAD.n435 2.24164
R39240 PAD.n744 PAD.n433 2.24164
R39241 PAD.n445 PAD.n435 2.24164
R39242 PAD.n752 PAD.n433 2.24164
R39243 PAD.n754 PAD.n435 2.24164
R39244 PAD.n756 PAD.n433 2.24164
R39245 PAD.n441 PAD.n435 2.24164
R39246 PAD.n765 PAD.n433 2.24164
R39247 PAD.n767 PAD.n435 2.24164
R39248 PAD.n769 PAD.n433 2.24164
R39249 PAD.n869 PAD.n828 2.24164
R39250 PAD.n10388 PAD.n823 2.24164
R39251 PAD.n878 PAD.n828 2.24164
R39252 PAD.n10388 PAD.n822 2.24164
R39253 PAD.n882 PAD.n828 2.24164
R39254 PAD.n10388 PAD.n821 2.24164
R39255 PAD.n890 PAD.n828 2.24164
R39256 PAD.n10388 PAD.n820 2.24164
R39257 PAD.n894 PAD.n828 2.24164
R39258 PAD.n10388 PAD.n819 2.24164
R39259 PAD.n902 PAD.n828 2.24164
R39260 PAD.n10388 PAD.n818 2.24164
R39261 PAD.n906 PAD.n828 2.24164
R39262 PAD.n10388 PAD.n817 2.24164
R39263 PAD.n914 PAD.n828 2.24164
R39264 PAD.n10388 PAD.n816 2.24164
R39265 PAD.n918 PAD.n828 2.24164
R39266 PAD.n10388 PAD.n815 2.24164
R39267 PAD.n926 PAD.n828 2.24164
R39268 PAD.n10388 PAD.n814 2.24164
R39269 PAD.n930 PAD.n828 2.24164
R39270 PAD.n10388 PAD.n813 2.24164
R39271 PAD.n938 PAD.n828 2.24164
R39272 PAD.n10388 PAD.n812 2.24164
R39273 PAD.n942 PAD.n828 2.24164
R39274 PAD.n10388 PAD.n811 2.24164
R39275 PAD.n950 PAD.n828 2.24164
R39276 PAD.n10388 PAD.n810 2.24164
R39277 PAD.n954 PAD.n828 2.24164
R39278 PAD.n10388 PAD.n809 2.24164
R39279 PAD.n962 PAD.n828 2.24164
R39280 PAD.n10388 PAD.n808 2.24164
R39281 PAD.n966 PAD.n828 2.24164
R39282 PAD.n10388 PAD.n807 2.24164
R39283 PAD.n974 PAD.n828 2.24164
R39284 PAD.n10388 PAD.n806 2.24164
R39285 PAD.n978 PAD.n828 2.24164
R39286 PAD.n10388 PAD.n805 2.24164
R39287 PAD.n986 PAD.n828 2.24164
R39288 PAD.n10388 PAD.n804 2.24164
R39289 PAD.n990 PAD.n828 2.24164
R39290 PAD.n10388 PAD.n803 2.24164
R39291 PAD.n998 PAD.n828 2.24164
R39292 PAD.n10388 PAD.n802 2.24164
R39293 PAD.n1002 PAD.n828 2.24164
R39294 PAD.n10388 PAD.n801 2.24164
R39295 PAD.n1010 PAD.n828 2.24164
R39296 PAD.n10388 PAD.n800 2.24164
R39297 PAD.n1014 PAD.n828 2.24164
R39298 PAD.n10388 PAD.n799 2.24164
R39299 PAD.n1022 PAD.n828 2.24164
R39300 PAD.n10388 PAD.n798 2.24164
R39301 PAD.n1026 PAD.n828 2.24164
R39302 PAD.n10388 PAD.n797 2.24164
R39303 PAD.n1034 PAD.n828 2.24164
R39304 PAD.n10388 PAD.n796 2.24164
R39305 PAD.n1038 PAD.n828 2.24164
R39306 PAD.n10388 PAD.n795 2.24164
R39307 PAD.n1046 PAD.n828 2.24164
R39308 PAD.n10388 PAD.n794 2.24164
R39309 PAD.n1050 PAD.n828 2.24164
R39310 PAD.n10388 PAD.n793 2.24164
R39311 PAD.n1058 PAD.n828 2.24164
R39312 PAD.n10388 PAD.n792 2.24164
R39313 PAD.n1062 PAD.n828 2.24164
R39314 PAD.n10388 PAD.n791 2.24164
R39315 PAD.n1070 PAD.n828 2.24164
R39316 PAD.n10388 PAD.n790 2.24164
R39317 PAD.n1074 PAD.n828 2.24164
R39318 PAD.n10388 PAD.n789 2.24164
R39319 PAD.n1082 PAD.n828 2.24164
R39320 PAD.n10388 PAD.n788 2.24164
R39321 PAD.n1086 PAD.n828 2.24164
R39322 PAD.n10388 PAD.n787 2.24164
R39323 PAD.n1094 PAD.n828 2.24164
R39324 PAD.n10388 PAD.n786 2.24164
R39325 PAD.n1098 PAD.n828 2.24164
R39326 PAD.n10388 PAD.n785 2.24164
R39327 PAD.n1106 PAD.n828 2.24164
R39328 PAD.n10388 PAD.n784 2.24164
R39329 PAD.n1110 PAD.n828 2.24164
R39330 PAD.n10388 PAD.n783 2.24164
R39331 PAD.n10386 PAD.n828 2.24164
R39332 PAD.n10107 PAD.n1130 2.24164
R39333 PAD.n10109 PAD.n1132 2.24164
R39334 PAD.n10111 PAD.n1130 2.24164
R39335 PAD.n10101 PAD.n1132 2.24164
R39336 PAD.n10119 PAD.n1130 2.24164
R39337 PAD.n10121 PAD.n1132 2.24164
R39338 PAD.n10123 PAD.n1130 2.24164
R39339 PAD.n10097 PAD.n1132 2.24164
R39340 PAD.n10131 PAD.n1130 2.24164
R39341 PAD.n10133 PAD.n1132 2.24164
R39342 PAD.n10135 PAD.n1130 2.24164
R39343 PAD.n10093 PAD.n1132 2.24164
R39344 PAD.n10143 PAD.n1130 2.24164
R39345 PAD.n10145 PAD.n1132 2.24164
R39346 PAD.n10147 PAD.n1130 2.24164
R39347 PAD.n10089 PAD.n1132 2.24164
R39348 PAD.n10155 PAD.n1130 2.24164
R39349 PAD.n10157 PAD.n1132 2.24164
R39350 PAD.n10159 PAD.n1130 2.24164
R39351 PAD.n10085 PAD.n1132 2.24164
R39352 PAD.n10167 PAD.n1130 2.24164
R39353 PAD.n10169 PAD.n1132 2.24164
R39354 PAD.n10171 PAD.n1130 2.24164
R39355 PAD.n10081 PAD.n1132 2.24164
R39356 PAD.n10179 PAD.n1130 2.24164
R39357 PAD.n10181 PAD.n1132 2.24164
R39358 PAD.n10183 PAD.n1130 2.24164
R39359 PAD.n10077 PAD.n1132 2.24164
R39360 PAD.n10191 PAD.n1130 2.24164
R39361 PAD.n10193 PAD.n1132 2.24164
R39362 PAD.n10195 PAD.n1130 2.24164
R39363 PAD.n10073 PAD.n1132 2.24164
R39364 PAD.n10203 PAD.n1130 2.24164
R39365 PAD.n10205 PAD.n1132 2.24164
R39366 PAD.n10207 PAD.n1130 2.24164
R39367 PAD.n10069 PAD.n1132 2.24164
R39368 PAD.n10215 PAD.n1130 2.24164
R39369 PAD.n10217 PAD.n1132 2.24164
R39370 PAD.n10219 PAD.n1130 2.24164
R39371 PAD.n10065 PAD.n1132 2.24164
R39372 PAD.n10227 PAD.n1130 2.24164
R39373 PAD.n10229 PAD.n1132 2.24164
R39374 PAD.n10231 PAD.n1130 2.24164
R39375 PAD.n10061 PAD.n1132 2.24164
R39376 PAD.n10239 PAD.n1130 2.24164
R39377 PAD.n10241 PAD.n1132 2.24164
R39378 PAD.n10243 PAD.n1130 2.24164
R39379 PAD.n10057 PAD.n1132 2.24164
R39380 PAD.n10251 PAD.n1130 2.24164
R39381 PAD.n10253 PAD.n1132 2.24164
R39382 PAD.n10255 PAD.n1130 2.24164
R39383 PAD.n10053 PAD.n1132 2.24164
R39384 PAD.n10263 PAD.n1130 2.24164
R39385 PAD.n10265 PAD.n1132 2.24164
R39386 PAD.n10267 PAD.n1130 2.24164
R39387 PAD.n10049 PAD.n1132 2.24164
R39388 PAD.n10275 PAD.n1130 2.24164
R39389 PAD.n10277 PAD.n1132 2.24164
R39390 PAD.n10279 PAD.n1130 2.24164
R39391 PAD.n10045 PAD.n1132 2.24164
R39392 PAD.n10287 PAD.n1130 2.24164
R39393 PAD.n10289 PAD.n1132 2.24164
R39394 PAD.n10291 PAD.n1130 2.24164
R39395 PAD.n10041 PAD.n1132 2.24164
R39396 PAD.n10299 PAD.n1130 2.24164
R39397 PAD.n10301 PAD.n1132 2.24164
R39398 PAD.n10303 PAD.n1130 2.24164
R39399 PAD.n10037 PAD.n1132 2.24164
R39400 PAD.n10311 PAD.n1130 2.24164
R39401 PAD.n10313 PAD.n1132 2.24164
R39402 PAD.n10315 PAD.n1130 2.24164
R39403 PAD.n10033 PAD.n1132 2.24164
R39404 PAD.n10323 PAD.n1130 2.24164
R39405 PAD.n10325 PAD.n1132 2.24164
R39406 PAD.n10327 PAD.n1130 2.24164
R39407 PAD.n10029 PAD.n1132 2.24164
R39408 PAD.n10335 PAD.n1130 2.24164
R39409 PAD.n10337 PAD.n1132 2.24164
R39410 PAD.n10339 PAD.n1130 2.24164
R39411 PAD.n10025 PAD.n1132 2.24164
R39412 PAD.n10348 PAD.n1130 2.24164
R39413 PAD.n10350 PAD.n1132 2.24164
R39414 PAD.n10352 PAD.n1130 2.24164
R39415 PAD.n1483 PAD.n1482 2.24164
R39416 PAD.n1191 PAD.n1140 2.24164
R39417 PAD.n1483 PAD.n1189 2.24164
R39418 PAD.n1473 PAD.n1140 2.24164
R39419 PAD.n1483 PAD.n1188 2.24164
R39420 PAD.n1197 PAD.n1140 2.24164
R39421 PAD.n1483 PAD.n1187 2.24164
R39422 PAD.n1464 PAD.n1140 2.24164
R39423 PAD.n1483 PAD.n1186 2.24164
R39424 PAD.n1202 PAD.n1140 2.24164
R39425 PAD.n1483 PAD.n1185 2.24164
R39426 PAD.n1455 PAD.n1140 2.24164
R39427 PAD.n1483 PAD.n1184 2.24164
R39428 PAD.n1207 PAD.n1140 2.24164
R39429 PAD.n1483 PAD.n1183 2.24164
R39430 PAD.n1446 PAD.n1140 2.24164
R39431 PAD.n1483 PAD.n1182 2.24164
R39432 PAD.n1212 PAD.n1140 2.24164
R39433 PAD.n1483 PAD.n1181 2.24164
R39434 PAD.n1437 PAD.n1140 2.24164
R39435 PAD.n1483 PAD.n1180 2.24164
R39436 PAD.n1217 PAD.n1140 2.24164
R39437 PAD.n1483 PAD.n1179 2.24164
R39438 PAD.n1428 PAD.n1140 2.24164
R39439 PAD.n1483 PAD.n1178 2.24164
R39440 PAD.n1222 PAD.n1140 2.24164
R39441 PAD.n1483 PAD.n1177 2.24164
R39442 PAD.n1419 PAD.n1140 2.24164
R39443 PAD.n1483 PAD.n1176 2.24164
R39444 PAD.n1227 PAD.n1140 2.24164
R39445 PAD.n1483 PAD.n1175 2.24164
R39446 PAD.n1410 PAD.n1140 2.24164
R39447 PAD.n1483 PAD.n1174 2.24164
R39448 PAD.n1232 PAD.n1140 2.24164
R39449 PAD.n1483 PAD.n1173 2.24164
R39450 PAD.n1401 PAD.n1140 2.24164
R39451 PAD.n1483 PAD.n1172 2.24164
R39452 PAD.n1237 PAD.n1140 2.24164
R39453 PAD.n1483 PAD.n1171 2.24164
R39454 PAD.n1392 PAD.n1140 2.24164
R39455 PAD.n1483 PAD.n1170 2.24164
R39456 PAD.n1242 PAD.n1140 2.24164
R39457 PAD.n1483 PAD.n1169 2.24164
R39458 PAD.n1383 PAD.n1140 2.24164
R39459 PAD.n1483 PAD.n1168 2.24164
R39460 PAD.n1247 PAD.n1140 2.24164
R39461 PAD.n1483 PAD.n1167 2.24164
R39462 PAD.n1374 PAD.n1140 2.24164
R39463 PAD.n1483 PAD.n1166 2.24164
R39464 PAD.n1252 PAD.n1140 2.24164
R39465 PAD.n1483 PAD.n1165 2.24164
R39466 PAD.n1365 PAD.n1140 2.24164
R39467 PAD.n1483 PAD.n1164 2.24164
R39468 PAD.n1257 PAD.n1140 2.24164
R39469 PAD.n1483 PAD.n1163 2.24164
R39470 PAD.n1356 PAD.n1140 2.24164
R39471 PAD.n1483 PAD.n1162 2.24164
R39472 PAD.n1262 PAD.n1140 2.24164
R39473 PAD.n1483 PAD.n1161 2.24164
R39474 PAD.n1347 PAD.n1140 2.24164
R39475 PAD.n1483 PAD.n1160 2.24164
R39476 PAD.n1267 PAD.n1140 2.24164
R39477 PAD.n1483 PAD.n1159 2.24164
R39478 PAD.n1338 PAD.n1140 2.24164
R39479 PAD.n1483 PAD.n1158 2.24164
R39480 PAD.n1272 PAD.n1140 2.24164
R39481 PAD.n1483 PAD.n1157 2.24164
R39482 PAD.n1329 PAD.n1140 2.24164
R39483 PAD.n1483 PAD.n1156 2.24164
R39484 PAD.n1277 PAD.n1140 2.24164
R39485 PAD.n1483 PAD.n1155 2.24164
R39486 PAD.n1320 PAD.n1140 2.24164
R39487 PAD.n1483 PAD.n1154 2.24164
R39488 PAD.n1282 PAD.n1140 2.24164
R39489 PAD.n1483 PAD.n1153 2.24164
R39490 PAD.n1311 PAD.n1140 2.24164
R39491 PAD.n1483 PAD.n1152 2.24164
R39492 PAD.n1287 PAD.n1140 2.24164
R39493 PAD.n1483 PAD.n1151 2.24164
R39494 PAD.n1302 PAD.n1140 2.24164
R39495 PAD.n1483 PAD.n1150 2.24164
R39496 PAD.n1292 PAD.n1140 2.24164
R39497 PAD.n1483 PAD.n1149 2.24164
R39498 PAD.n1577 PAD.n1536 2.24164
R39499 PAD.n9998 PAD.n1530 2.24164
R39500 PAD.n9755 PAD.n1536 2.24164
R39501 PAD.n9998 PAD.n1529 2.24164
R39502 PAD.n9759 PAD.n1536 2.24164
R39503 PAD.n9998 PAD.n1528 2.24164
R39504 PAD.n9767 PAD.n1536 2.24164
R39505 PAD.n9998 PAD.n1527 2.24164
R39506 PAD.n9771 PAD.n1536 2.24164
R39507 PAD.n9998 PAD.n1526 2.24164
R39508 PAD.n9779 PAD.n1536 2.24164
R39509 PAD.n9998 PAD.n1525 2.24164
R39510 PAD.n9783 PAD.n1536 2.24164
R39511 PAD.n9998 PAD.n1524 2.24164
R39512 PAD.n9791 PAD.n1536 2.24164
R39513 PAD.n9998 PAD.n1523 2.24164
R39514 PAD.n9795 PAD.n1536 2.24164
R39515 PAD.n9998 PAD.n1522 2.24164
R39516 PAD.n9803 PAD.n1536 2.24164
R39517 PAD.n9998 PAD.n1521 2.24164
R39518 PAD.n9807 PAD.n1536 2.24164
R39519 PAD.n9998 PAD.n1520 2.24164
R39520 PAD.n9815 PAD.n1536 2.24164
R39521 PAD.n9998 PAD.n1519 2.24164
R39522 PAD.n9819 PAD.n1536 2.24164
R39523 PAD.n9998 PAD.n1518 2.24164
R39524 PAD.n9827 PAD.n1536 2.24164
R39525 PAD.n9998 PAD.n1517 2.24164
R39526 PAD.n9831 PAD.n1536 2.24164
R39527 PAD.n9998 PAD.n1516 2.24164
R39528 PAD.n9839 PAD.n1536 2.24164
R39529 PAD.n9998 PAD.n1515 2.24164
R39530 PAD.n9843 PAD.n1536 2.24164
R39531 PAD.n9998 PAD.n1514 2.24164
R39532 PAD.n9851 PAD.n1536 2.24164
R39533 PAD.n9998 PAD.n1513 2.24164
R39534 PAD.n9855 PAD.n1536 2.24164
R39535 PAD.n9998 PAD.n1512 2.24164
R39536 PAD.n9863 PAD.n1536 2.24164
R39537 PAD.n9998 PAD.n1511 2.24164
R39538 PAD.n9867 PAD.n1536 2.24164
R39539 PAD.n9998 PAD.n1510 2.24164
R39540 PAD.n9875 PAD.n1536 2.24164
R39541 PAD.n9998 PAD.n1509 2.24164
R39542 PAD.n9879 PAD.n1536 2.24164
R39543 PAD.n9998 PAD.n1508 2.24164
R39544 PAD.n9887 PAD.n1536 2.24164
R39545 PAD.n9998 PAD.n1507 2.24164
R39546 PAD.n9891 PAD.n1536 2.24164
R39547 PAD.n9998 PAD.n1506 2.24164
R39548 PAD.n9899 PAD.n1536 2.24164
R39549 PAD.n9998 PAD.n1505 2.24164
R39550 PAD.n9903 PAD.n1536 2.24164
R39551 PAD.n9998 PAD.n1504 2.24164
R39552 PAD.n9911 PAD.n1536 2.24164
R39553 PAD.n9998 PAD.n1503 2.24164
R39554 PAD.n9915 PAD.n1536 2.24164
R39555 PAD.n9998 PAD.n1502 2.24164
R39556 PAD.n9923 PAD.n1536 2.24164
R39557 PAD.n9998 PAD.n1501 2.24164
R39558 PAD.n9927 PAD.n1536 2.24164
R39559 PAD.n9998 PAD.n1500 2.24164
R39560 PAD.n9935 PAD.n1536 2.24164
R39561 PAD.n9998 PAD.n1499 2.24164
R39562 PAD.n9939 PAD.n1536 2.24164
R39563 PAD.n9998 PAD.n1498 2.24164
R39564 PAD.n9947 PAD.n1536 2.24164
R39565 PAD.n9998 PAD.n1497 2.24164
R39566 PAD.n9951 PAD.n1536 2.24164
R39567 PAD.n9998 PAD.n1496 2.24164
R39568 PAD.n9959 PAD.n1536 2.24164
R39569 PAD.n9998 PAD.n1495 2.24164
R39570 PAD.n9963 PAD.n1536 2.24164
R39571 PAD.n9998 PAD.n1494 2.24164
R39572 PAD.n9971 PAD.n1536 2.24164
R39573 PAD.n9998 PAD.n1493 2.24164
R39574 PAD.n9975 PAD.n1536 2.24164
R39575 PAD.n9998 PAD.n1492 2.24164
R39576 PAD.n9983 PAD.n1536 2.24164
R39577 PAD.n9998 PAD.n1491 2.24164
R39578 PAD.n9987 PAD.n1536 2.24164
R39579 PAD.n9998 PAD.n1490 2.24164
R39580 PAD.n9996 PAD.n1536 2.24164
R39581 PAD.n1601 PAD.n1592 2.24164
R39582 PAD.n1928 PAD.n1594 2.24164
R39583 PAD.n1926 PAD.n1592 2.24164
R39584 PAD.n1602 PAD.n1594 2.24164
R39585 PAD.n1918 PAD.n1592 2.24164
R39586 PAD.n1916 PAD.n1594 2.24164
R39587 PAD.n1914 PAD.n1592 2.24164
R39588 PAD.n1607 PAD.n1594 2.24164
R39589 PAD.n1906 PAD.n1592 2.24164
R39590 PAD.n1904 PAD.n1594 2.24164
R39591 PAD.n1902 PAD.n1592 2.24164
R39592 PAD.n1611 PAD.n1594 2.24164
R39593 PAD.n1894 PAD.n1592 2.24164
R39594 PAD.n1892 PAD.n1594 2.24164
R39595 PAD.n1890 PAD.n1592 2.24164
R39596 PAD.n1615 PAD.n1594 2.24164
R39597 PAD.n1882 PAD.n1592 2.24164
R39598 PAD.n1880 PAD.n1594 2.24164
R39599 PAD.n1878 PAD.n1592 2.24164
R39600 PAD.n1619 PAD.n1594 2.24164
R39601 PAD.n1870 PAD.n1592 2.24164
R39602 PAD.n1868 PAD.n1594 2.24164
R39603 PAD.n1866 PAD.n1592 2.24164
R39604 PAD.n1623 PAD.n1594 2.24164
R39605 PAD.n1858 PAD.n1592 2.24164
R39606 PAD.n1856 PAD.n1594 2.24164
R39607 PAD.n1854 PAD.n1592 2.24164
R39608 PAD.n1627 PAD.n1594 2.24164
R39609 PAD.n1846 PAD.n1592 2.24164
R39610 PAD.n1844 PAD.n1594 2.24164
R39611 PAD.n1842 PAD.n1592 2.24164
R39612 PAD.n1631 PAD.n1594 2.24164
R39613 PAD.n1834 PAD.n1592 2.24164
R39614 PAD.n1832 PAD.n1594 2.24164
R39615 PAD.n1830 PAD.n1592 2.24164
R39616 PAD.n1635 PAD.n1594 2.24164
R39617 PAD.n1822 PAD.n1592 2.24164
R39618 PAD.n1820 PAD.n1594 2.24164
R39619 PAD.n1818 PAD.n1592 2.24164
R39620 PAD.n1639 PAD.n1594 2.24164
R39621 PAD.n1810 PAD.n1592 2.24164
R39622 PAD.n1808 PAD.n1594 2.24164
R39623 PAD.n1806 PAD.n1592 2.24164
R39624 PAD.n1643 PAD.n1594 2.24164
R39625 PAD.n1798 PAD.n1592 2.24164
R39626 PAD.n1796 PAD.n1594 2.24164
R39627 PAD.n1794 PAD.n1592 2.24164
R39628 PAD.n1647 PAD.n1594 2.24164
R39629 PAD.n1786 PAD.n1592 2.24164
R39630 PAD.n1784 PAD.n1594 2.24164
R39631 PAD.n1782 PAD.n1592 2.24164
R39632 PAD.n1651 PAD.n1594 2.24164
R39633 PAD.n1774 PAD.n1592 2.24164
R39634 PAD.n1772 PAD.n1594 2.24164
R39635 PAD.n1770 PAD.n1592 2.24164
R39636 PAD.n1655 PAD.n1594 2.24164
R39637 PAD.n1762 PAD.n1592 2.24164
R39638 PAD.n1760 PAD.n1594 2.24164
R39639 PAD.n1758 PAD.n1592 2.24164
R39640 PAD.n1659 PAD.n1594 2.24164
R39641 PAD.n1750 PAD.n1592 2.24164
R39642 PAD.n1748 PAD.n1594 2.24164
R39643 PAD.n1746 PAD.n1592 2.24164
R39644 PAD.n1663 PAD.n1594 2.24164
R39645 PAD.n1738 PAD.n1592 2.24164
R39646 PAD.n1736 PAD.n1594 2.24164
R39647 PAD.n1734 PAD.n1592 2.24164
R39648 PAD.n1667 PAD.n1594 2.24164
R39649 PAD.n1726 PAD.n1592 2.24164
R39650 PAD.n1724 PAD.n1594 2.24164
R39651 PAD.n1722 PAD.n1592 2.24164
R39652 PAD.n1671 PAD.n1594 2.24164
R39653 PAD.n1714 PAD.n1592 2.24164
R39654 PAD.n1712 PAD.n1594 2.24164
R39655 PAD.n1710 PAD.n1592 2.24164
R39656 PAD.n1675 PAD.n1594 2.24164
R39657 PAD.n1702 PAD.n1592 2.24164
R39658 PAD.n1700 PAD.n1594 2.24164
R39659 PAD.n1698 PAD.n1592 2.24164
R39660 PAD.n1679 PAD.n1594 2.24164
R39661 PAD.n1690 PAD.n1592 2.24164
R39662 PAD.n1688 PAD.n1594 2.24164
R39663 PAD.n1686 PAD.n1592 2.24164
R39664 PAD.n2029 PAD.n1988 2.24164
R39665 PAD.n9712 PAD.n1983 2.24164
R39666 PAD.n9469 PAD.n1988 2.24164
R39667 PAD.n9712 PAD.n1982 2.24164
R39668 PAD.n9473 PAD.n1988 2.24164
R39669 PAD.n9712 PAD.n1981 2.24164
R39670 PAD.n9481 PAD.n1988 2.24164
R39671 PAD.n9712 PAD.n1980 2.24164
R39672 PAD.n9485 PAD.n1988 2.24164
R39673 PAD.n9712 PAD.n1979 2.24164
R39674 PAD.n9493 PAD.n1988 2.24164
R39675 PAD.n9712 PAD.n1978 2.24164
R39676 PAD.n9497 PAD.n1988 2.24164
R39677 PAD.n9712 PAD.n1977 2.24164
R39678 PAD.n9505 PAD.n1988 2.24164
R39679 PAD.n9712 PAD.n1976 2.24164
R39680 PAD.n9509 PAD.n1988 2.24164
R39681 PAD.n9712 PAD.n1975 2.24164
R39682 PAD.n9517 PAD.n1988 2.24164
R39683 PAD.n9712 PAD.n1974 2.24164
R39684 PAD.n9521 PAD.n1988 2.24164
R39685 PAD.n9712 PAD.n1973 2.24164
R39686 PAD.n9529 PAD.n1988 2.24164
R39687 PAD.n9712 PAD.n1972 2.24164
R39688 PAD.n9533 PAD.n1988 2.24164
R39689 PAD.n9712 PAD.n1971 2.24164
R39690 PAD.n9541 PAD.n1988 2.24164
R39691 PAD.n9712 PAD.n1970 2.24164
R39692 PAD.n9545 PAD.n1988 2.24164
R39693 PAD.n9712 PAD.n1969 2.24164
R39694 PAD.n9553 PAD.n1988 2.24164
R39695 PAD.n9712 PAD.n1968 2.24164
R39696 PAD.n9557 PAD.n1988 2.24164
R39697 PAD.n9712 PAD.n1967 2.24164
R39698 PAD.n9565 PAD.n1988 2.24164
R39699 PAD.n9712 PAD.n1966 2.24164
R39700 PAD.n9569 PAD.n1988 2.24164
R39701 PAD.n9712 PAD.n1965 2.24164
R39702 PAD.n9577 PAD.n1988 2.24164
R39703 PAD.n9712 PAD.n1964 2.24164
R39704 PAD.n9581 PAD.n1988 2.24164
R39705 PAD.n9712 PAD.n1963 2.24164
R39706 PAD.n9589 PAD.n1988 2.24164
R39707 PAD.n9712 PAD.n1962 2.24164
R39708 PAD.n9593 PAD.n1988 2.24164
R39709 PAD.n9712 PAD.n1961 2.24164
R39710 PAD.n9601 PAD.n1988 2.24164
R39711 PAD.n9712 PAD.n1960 2.24164
R39712 PAD.n9605 PAD.n1988 2.24164
R39713 PAD.n9712 PAD.n1959 2.24164
R39714 PAD.n9613 PAD.n1988 2.24164
R39715 PAD.n9712 PAD.n1958 2.24164
R39716 PAD.n9617 PAD.n1988 2.24164
R39717 PAD.n9712 PAD.n1957 2.24164
R39718 PAD.n9625 PAD.n1988 2.24164
R39719 PAD.n9712 PAD.n1956 2.24164
R39720 PAD.n9629 PAD.n1988 2.24164
R39721 PAD.n9712 PAD.n1955 2.24164
R39722 PAD.n9637 PAD.n1988 2.24164
R39723 PAD.n9712 PAD.n1954 2.24164
R39724 PAD.n9641 PAD.n1988 2.24164
R39725 PAD.n9712 PAD.n1953 2.24164
R39726 PAD.n9649 PAD.n1988 2.24164
R39727 PAD.n9712 PAD.n1952 2.24164
R39728 PAD.n9653 PAD.n1988 2.24164
R39729 PAD.n9712 PAD.n1951 2.24164
R39730 PAD.n9661 PAD.n1988 2.24164
R39731 PAD.n9712 PAD.n1950 2.24164
R39732 PAD.n9665 PAD.n1988 2.24164
R39733 PAD.n9712 PAD.n1949 2.24164
R39734 PAD.n9673 PAD.n1988 2.24164
R39735 PAD.n9712 PAD.n1948 2.24164
R39736 PAD.n9677 PAD.n1988 2.24164
R39737 PAD.n9712 PAD.n1947 2.24164
R39738 PAD.n9685 PAD.n1988 2.24164
R39739 PAD.n9712 PAD.n1946 2.24164
R39740 PAD.n9689 PAD.n1988 2.24164
R39741 PAD.n9712 PAD.n1945 2.24164
R39742 PAD.n9697 PAD.n1988 2.24164
R39743 PAD.n9712 PAD.n1944 2.24164
R39744 PAD.n9701 PAD.n1988 2.24164
R39745 PAD.n9712 PAD.n1943 2.24164
R39746 PAD.n9710 PAD.n1988 2.24164
R39747 PAD.n2132 PAD.n2091 2.24164
R39748 PAD.n9445 PAD.n2087 2.24164
R39749 PAD.n9203 PAD.n2091 2.24164
R39750 PAD.n9445 PAD.n2086 2.24164
R39751 PAD.n9207 PAD.n2091 2.24164
R39752 PAD.n9445 PAD.n2085 2.24164
R39753 PAD.n9215 PAD.n2091 2.24164
R39754 PAD.n9445 PAD.n2084 2.24164
R39755 PAD.n9219 PAD.n2091 2.24164
R39756 PAD.n9445 PAD.n2083 2.24164
R39757 PAD.n9227 PAD.n2091 2.24164
R39758 PAD.n9445 PAD.n2082 2.24164
R39759 PAD.n9231 PAD.n2091 2.24164
R39760 PAD.n9445 PAD.n2081 2.24164
R39761 PAD.n9239 PAD.n2091 2.24164
R39762 PAD.n9445 PAD.n2080 2.24164
R39763 PAD.n9243 PAD.n2091 2.24164
R39764 PAD.n9445 PAD.n2079 2.24164
R39765 PAD.n9251 PAD.n2091 2.24164
R39766 PAD.n9445 PAD.n2078 2.24164
R39767 PAD.n9255 PAD.n2091 2.24164
R39768 PAD.n9445 PAD.n2077 2.24164
R39769 PAD.n9263 PAD.n2091 2.24164
R39770 PAD.n9445 PAD.n2076 2.24164
R39771 PAD.n9267 PAD.n2091 2.24164
R39772 PAD.n9445 PAD.n2075 2.24164
R39773 PAD.n9275 PAD.n2091 2.24164
R39774 PAD.n9445 PAD.n2074 2.24164
R39775 PAD.n9279 PAD.n2091 2.24164
R39776 PAD.n9445 PAD.n2073 2.24164
R39777 PAD.n9287 PAD.n2091 2.24164
R39778 PAD.n9445 PAD.n2072 2.24164
R39779 PAD.n9291 PAD.n2091 2.24164
R39780 PAD.n9445 PAD.n2071 2.24164
R39781 PAD.n9299 PAD.n2091 2.24164
R39782 PAD.n9445 PAD.n2070 2.24164
R39783 PAD.n9303 PAD.n2091 2.24164
R39784 PAD.n9445 PAD.n2069 2.24164
R39785 PAD.n9311 PAD.n2091 2.24164
R39786 PAD.n9445 PAD.n2068 2.24164
R39787 PAD.n9315 PAD.n2091 2.24164
R39788 PAD.n9445 PAD.n2067 2.24164
R39789 PAD.n9323 PAD.n2091 2.24164
R39790 PAD.n9445 PAD.n2066 2.24164
R39791 PAD.n9327 PAD.n2091 2.24164
R39792 PAD.n9445 PAD.n2065 2.24164
R39793 PAD.n9335 PAD.n2091 2.24164
R39794 PAD.n9445 PAD.n2064 2.24164
R39795 PAD.n9339 PAD.n2091 2.24164
R39796 PAD.n9445 PAD.n2063 2.24164
R39797 PAD.n9347 PAD.n2091 2.24164
R39798 PAD.n9445 PAD.n2062 2.24164
R39799 PAD.n9351 PAD.n2091 2.24164
R39800 PAD.n9445 PAD.n2061 2.24164
R39801 PAD.n9359 PAD.n2091 2.24164
R39802 PAD.n9445 PAD.n2060 2.24164
R39803 PAD.n9363 PAD.n2091 2.24164
R39804 PAD.n9445 PAD.n2059 2.24164
R39805 PAD.n9371 PAD.n2091 2.24164
R39806 PAD.n9445 PAD.n2058 2.24164
R39807 PAD.n9375 PAD.n2091 2.24164
R39808 PAD.n9445 PAD.n2057 2.24164
R39809 PAD.n9383 PAD.n2091 2.24164
R39810 PAD.n9445 PAD.n2056 2.24164
R39811 PAD.n9387 PAD.n2091 2.24164
R39812 PAD.n9445 PAD.n2055 2.24164
R39813 PAD.n9395 PAD.n2091 2.24164
R39814 PAD.n9445 PAD.n2054 2.24164
R39815 PAD.n9399 PAD.n2091 2.24164
R39816 PAD.n9445 PAD.n2053 2.24164
R39817 PAD.n9407 PAD.n2091 2.24164
R39818 PAD.n9445 PAD.n2052 2.24164
R39819 PAD.n9411 PAD.n2091 2.24164
R39820 PAD.n9445 PAD.n2051 2.24164
R39821 PAD.n9419 PAD.n2091 2.24164
R39822 PAD.n9445 PAD.n2050 2.24164
R39823 PAD.n9423 PAD.n2091 2.24164
R39824 PAD.n9445 PAD.n2049 2.24164
R39825 PAD.n9431 PAD.n2091 2.24164
R39826 PAD.n9445 PAD.n2048 2.24164
R39827 PAD.n9435 PAD.n2091 2.24164
R39828 PAD.n9445 PAD.n2047 2.24164
R39829 PAD.n9443 PAD.n2091 2.24164
R39830 PAD.n2153 PAD.n2146 2.24164
R39831 PAD.n2479 PAD.n2139 2.24164
R39832 PAD.n2477 PAD.n2146 2.24164
R39833 PAD.n2154 PAD.n2139 2.24164
R39834 PAD.n2469 PAD.n2146 2.24164
R39835 PAD.n2467 PAD.n2139 2.24164
R39836 PAD.n2465 PAD.n2146 2.24164
R39837 PAD.n2159 PAD.n2139 2.24164
R39838 PAD.n2457 PAD.n2146 2.24164
R39839 PAD.n2455 PAD.n2139 2.24164
R39840 PAD.n2453 PAD.n2146 2.24164
R39841 PAD.n2163 PAD.n2139 2.24164
R39842 PAD.n2445 PAD.n2146 2.24164
R39843 PAD.n2443 PAD.n2139 2.24164
R39844 PAD.n2441 PAD.n2146 2.24164
R39845 PAD.n2167 PAD.n2139 2.24164
R39846 PAD.n2433 PAD.n2146 2.24164
R39847 PAD.n2431 PAD.n2139 2.24164
R39848 PAD.n2429 PAD.n2146 2.24164
R39849 PAD.n2171 PAD.n2139 2.24164
R39850 PAD.n2421 PAD.n2146 2.24164
R39851 PAD.n2419 PAD.n2139 2.24164
R39852 PAD.n2417 PAD.n2146 2.24164
R39853 PAD.n2175 PAD.n2139 2.24164
R39854 PAD.n2409 PAD.n2146 2.24164
R39855 PAD.n2407 PAD.n2139 2.24164
R39856 PAD.n2405 PAD.n2146 2.24164
R39857 PAD.n2179 PAD.n2139 2.24164
R39858 PAD.n2397 PAD.n2146 2.24164
R39859 PAD.n2395 PAD.n2139 2.24164
R39860 PAD.n2393 PAD.n2146 2.24164
R39861 PAD.n2183 PAD.n2139 2.24164
R39862 PAD.n2385 PAD.n2146 2.24164
R39863 PAD.n2383 PAD.n2139 2.24164
R39864 PAD.n2381 PAD.n2146 2.24164
R39865 PAD.n2187 PAD.n2139 2.24164
R39866 PAD.n2373 PAD.n2146 2.24164
R39867 PAD.n2371 PAD.n2139 2.24164
R39868 PAD.n2369 PAD.n2146 2.24164
R39869 PAD.n2191 PAD.n2139 2.24164
R39870 PAD.n2361 PAD.n2146 2.24164
R39871 PAD.n2359 PAD.n2139 2.24164
R39872 PAD.n2357 PAD.n2146 2.24164
R39873 PAD.n2195 PAD.n2139 2.24164
R39874 PAD.n2349 PAD.n2146 2.24164
R39875 PAD.n2347 PAD.n2139 2.24164
R39876 PAD.n2345 PAD.n2146 2.24164
R39877 PAD.n2199 PAD.n2139 2.24164
R39878 PAD.n2337 PAD.n2146 2.24164
R39879 PAD.n2335 PAD.n2139 2.24164
R39880 PAD.n2333 PAD.n2146 2.24164
R39881 PAD.n2203 PAD.n2139 2.24164
R39882 PAD.n2325 PAD.n2146 2.24164
R39883 PAD.n2323 PAD.n2139 2.24164
R39884 PAD.n2321 PAD.n2146 2.24164
R39885 PAD.n2207 PAD.n2139 2.24164
R39886 PAD.n2313 PAD.n2146 2.24164
R39887 PAD.n2311 PAD.n2139 2.24164
R39888 PAD.n2309 PAD.n2146 2.24164
R39889 PAD.n2211 PAD.n2139 2.24164
R39890 PAD.n2301 PAD.n2146 2.24164
R39891 PAD.n2299 PAD.n2139 2.24164
R39892 PAD.n2297 PAD.n2146 2.24164
R39893 PAD.n2215 PAD.n2139 2.24164
R39894 PAD.n2289 PAD.n2146 2.24164
R39895 PAD.n2287 PAD.n2139 2.24164
R39896 PAD.n2285 PAD.n2146 2.24164
R39897 PAD.n2219 PAD.n2139 2.24164
R39898 PAD.n2277 PAD.n2146 2.24164
R39899 PAD.n2275 PAD.n2139 2.24164
R39900 PAD.n2273 PAD.n2146 2.24164
R39901 PAD.n2223 PAD.n2139 2.24164
R39902 PAD.n2265 PAD.n2146 2.24164
R39903 PAD.n2263 PAD.n2139 2.24164
R39904 PAD.n2261 PAD.n2146 2.24164
R39905 PAD.n2227 PAD.n2139 2.24164
R39906 PAD.n2253 PAD.n2146 2.24164
R39907 PAD.n2251 PAD.n2139 2.24164
R39908 PAD.n2249 PAD.n2146 2.24164
R39909 PAD.n2231 PAD.n2139 2.24164
R39910 PAD.n2241 PAD.n2146 2.24164
R39911 PAD.n2239 PAD.n2139 2.24164
R39912 PAD.n2237 PAD.n2146 2.24164
R39913 PAD.n2500 PAD.n2494 2.24164
R39914 PAD.n2826 PAD.n2487 2.24164
R39915 PAD.n2824 PAD.n2494 2.24164
R39916 PAD.n2501 PAD.n2487 2.24164
R39917 PAD.n2816 PAD.n2494 2.24164
R39918 PAD.n2814 PAD.n2487 2.24164
R39919 PAD.n2812 PAD.n2494 2.24164
R39920 PAD.n2506 PAD.n2487 2.24164
R39921 PAD.n2804 PAD.n2494 2.24164
R39922 PAD.n2802 PAD.n2487 2.24164
R39923 PAD.n2800 PAD.n2494 2.24164
R39924 PAD.n2510 PAD.n2487 2.24164
R39925 PAD.n2792 PAD.n2494 2.24164
R39926 PAD.n2790 PAD.n2487 2.24164
R39927 PAD.n2788 PAD.n2494 2.24164
R39928 PAD.n2514 PAD.n2487 2.24164
R39929 PAD.n2780 PAD.n2494 2.24164
R39930 PAD.n2778 PAD.n2487 2.24164
R39931 PAD.n2776 PAD.n2494 2.24164
R39932 PAD.n2518 PAD.n2487 2.24164
R39933 PAD.n2768 PAD.n2494 2.24164
R39934 PAD.n2766 PAD.n2487 2.24164
R39935 PAD.n2764 PAD.n2494 2.24164
R39936 PAD.n2522 PAD.n2487 2.24164
R39937 PAD.n2756 PAD.n2494 2.24164
R39938 PAD.n2754 PAD.n2487 2.24164
R39939 PAD.n2752 PAD.n2494 2.24164
R39940 PAD.n2526 PAD.n2487 2.24164
R39941 PAD.n2744 PAD.n2494 2.24164
R39942 PAD.n2742 PAD.n2487 2.24164
R39943 PAD.n2740 PAD.n2494 2.24164
R39944 PAD.n2530 PAD.n2487 2.24164
R39945 PAD.n2732 PAD.n2494 2.24164
R39946 PAD.n2730 PAD.n2487 2.24164
R39947 PAD.n2728 PAD.n2494 2.24164
R39948 PAD.n2534 PAD.n2487 2.24164
R39949 PAD.n2720 PAD.n2494 2.24164
R39950 PAD.n2718 PAD.n2487 2.24164
R39951 PAD.n2716 PAD.n2494 2.24164
R39952 PAD.n2538 PAD.n2487 2.24164
R39953 PAD.n2708 PAD.n2494 2.24164
R39954 PAD.n2706 PAD.n2487 2.24164
R39955 PAD.n2704 PAD.n2494 2.24164
R39956 PAD.n2542 PAD.n2487 2.24164
R39957 PAD.n2696 PAD.n2494 2.24164
R39958 PAD.n2694 PAD.n2487 2.24164
R39959 PAD.n2692 PAD.n2494 2.24164
R39960 PAD.n2546 PAD.n2487 2.24164
R39961 PAD.n2684 PAD.n2494 2.24164
R39962 PAD.n2682 PAD.n2487 2.24164
R39963 PAD.n2680 PAD.n2494 2.24164
R39964 PAD.n2550 PAD.n2487 2.24164
R39965 PAD.n2672 PAD.n2494 2.24164
R39966 PAD.n2670 PAD.n2487 2.24164
R39967 PAD.n2668 PAD.n2494 2.24164
R39968 PAD.n2554 PAD.n2487 2.24164
R39969 PAD.n2660 PAD.n2494 2.24164
R39970 PAD.n2658 PAD.n2487 2.24164
R39971 PAD.n2656 PAD.n2494 2.24164
R39972 PAD.n2558 PAD.n2487 2.24164
R39973 PAD.n2648 PAD.n2494 2.24164
R39974 PAD.n2646 PAD.n2487 2.24164
R39975 PAD.n2644 PAD.n2494 2.24164
R39976 PAD.n2562 PAD.n2487 2.24164
R39977 PAD.n2636 PAD.n2494 2.24164
R39978 PAD.n2634 PAD.n2487 2.24164
R39979 PAD.n2632 PAD.n2494 2.24164
R39980 PAD.n2566 PAD.n2487 2.24164
R39981 PAD.n2624 PAD.n2494 2.24164
R39982 PAD.n2622 PAD.n2487 2.24164
R39983 PAD.n2620 PAD.n2494 2.24164
R39984 PAD.n2570 PAD.n2487 2.24164
R39985 PAD.n2612 PAD.n2494 2.24164
R39986 PAD.n2610 PAD.n2487 2.24164
R39987 PAD.n2608 PAD.n2494 2.24164
R39988 PAD.n2574 PAD.n2487 2.24164
R39989 PAD.n2600 PAD.n2494 2.24164
R39990 PAD.n2598 PAD.n2487 2.24164
R39991 PAD.n2596 PAD.n2494 2.24164
R39992 PAD.n2578 PAD.n2487 2.24164
R39993 PAD.n2588 PAD.n2494 2.24164
R39994 PAD.n2586 PAD.n2487 2.24164
R39995 PAD.n2584 PAD.n2494 2.24164
R39996 PAD.n9116 PAD.n2879 2.24164
R39997 PAD.n9140 PAD.n2875 2.24164
R39998 PAD.n8840 PAD.n2879 2.24164
R39999 PAD.n9140 PAD.n2874 2.24164
R40000 PAD.n9109 PAD.n2879 2.24164
R40001 PAD.n9140 PAD.n2873 2.24164
R40002 PAD.n8845 PAD.n2879 2.24164
R40003 PAD.n9140 PAD.n2872 2.24164
R40004 PAD.n9100 PAD.n2879 2.24164
R40005 PAD.n9140 PAD.n2871 2.24164
R40006 PAD.n8850 PAD.n2879 2.24164
R40007 PAD.n9140 PAD.n2870 2.24164
R40008 PAD.n9091 PAD.n2879 2.24164
R40009 PAD.n9140 PAD.n2869 2.24164
R40010 PAD.n8855 PAD.n2879 2.24164
R40011 PAD.n9140 PAD.n2868 2.24164
R40012 PAD.n9082 PAD.n2879 2.24164
R40013 PAD.n9140 PAD.n2867 2.24164
R40014 PAD.n8860 PAD.n2879 2.24164
R40015 PAD.n9140 PAD.n2866 2.24164
R40016 PAD.n9073 PAD.n2879 2.24164
R40017 PAD.n9140 PAD.n2865 2.24164
R40018 PAD.n8865 PAD.n2879 2.24164
R40019 PAD.n9140 PAD.n2864 2.24164
R40020 PAD.n9064 PAD.n2879 2.24164
R40021 PAD.n9140 PAD.n2863 2.24164
R40022 PAD.n8870 PAD.n2879 2.24164
R40023 PAD.n9140 PAD.n2862 2.24164
R40024 PAD.n9055 PAD.n2879 2.24164
R40025 PAD.n9140 PAD.n2861 2.24164
R40026 PAD.n8875 PAD.n2879 2.24164
R40027 PAD.n9140 PAD.n2860 2.24164
R40028 PAD.n9046 PAD.n2879 2.24164
R40029 PAD.n9140 PAD.n2859 2.24164
R40030 PAD.n8880 PAD.n2879 2.24164
R40031 PAD.n9140 PAD.n2858 2.24164
R40032 PAD.n9037 PAD.n2879 2.24164
R40033 PAD.n9140 PAD.n2857 2.24164
R40034 PAD.n8885 PAD.n2879 2.24164
R40035 PAD.n9140 PAD.n2856 2.24164
R40036 PAD.n9028 PAD.n2879 2.24164
R40037 PAD.n9140 PAD.n2855 2.24164
R40038 PAD.n8890 PAD.n2879 2.24164
R40039 PAD.n9140 PAD.n2854 2.24164
R40040 PAD.n9019 PAD.n2879 2.24164
R40041 PAD.n9140 PAD.n2853 2.24164
R40042 PAD.n8895 PAD.n2879 2.24164
R40043 PAD.n9140 PAD.n2852 2.24164
R40044 PAD.n9010 PAD.n2879 2.24164
R40045 PAD.n9140 PAD.n2851 2.24164
R40046 PAD.n8900 PAD.n2879 2.24164
R40047 PAD.n9140 PAD.n2850 2.24164
R40048 PAD.n9001 PAD.n2879 2.24164
R40049 PAD.n9140 PAD.n2849 2.24164
R40050 PAD.n8905 PAD.n2879 2.24164
R40051 PAD.n9140 PAD.n2848 2.24164
R40052 PAD.n8992 PAD.n2879 2.24164
R40053 PAD.n9140 PAD.n2847 2.24164
R40054 PAD.n8910 PAD.n2879 2.24164
R40055 PAD.n9140 PAD.n2846 2.24164
R40056 PAD.n8983 PAD.n2879 2.24164
R40057 PAD.n9140 PAD.n2845 2.24164
R40058 PAD.n8915 PAD.n2879 2.24164
R40059 PAD.n9140 PAD.n2844 2.24164
R40060 PAD.n8974 PAD.n2879 2.24164
R40061 PAD.n9140 PAD.n2843 2.24164
R40062 PAD.n8920 PAD.n2879 2.24164
R40063 PAD.n9140 PAD.n2842 2.24164
R40064 PAD.n8965 PAD.n2879 2.24164
R40065 PAD.n9140 PAD.n2841 2.24164
R40066 PAD.n8925 PAD.n2879 2.24164
R40067 PAD.n9140 PAD.n2840 2.24164
R40068 PAD.n8956 PAD.n2879 2.24164
R40069 PAD.n9140 PAD.n2839 2.24164
R40070 PAD.n8930 PAD.n2879 2.24164
R40071 PAD.n9140 PAD.n2838 2.24164
R40072 PAD.n8947 PAD.n2879 2.24164
R40073 PAD.n9140 PAD.n2837 2.24164
R40074 PAD.n8935 PAD.n2879 2.24164
R40075 PAD.n9140 PAD.n2836 2.24164
R40076 PAD.n8938 PAD.n2879 2.24164
R40077 PAD.n9140 PAD.n2835 2.24164
R40078 PAD.n9138 PAD.n2879 2.24164
R40079 PAD.n8821 PAD.n8820 2.24164
R40080 PAD.n8812 PAD.n2891 2.24164
R40081 PAD.n8821 PAD.n2945 2.24164
R40082 PAD.n8809 PAD.n2891 2.24164
R40083 PAD.n8821 PAD.n2944 2.24164
R40084 PAD.n8801 PAD.n2891 2.24164
R40085 PAD.n8821 PAD.n2943 2.24164
R40086 PAD.n8797 PAD.n2891 2.24164
R40087 PAD.n8821 PAD.n2942 2.24164
R40088 PAD.n8789 PAD.n2891 2.24164
R40089 PAD.n8821 PAD.n2941 2.24164
R40090 PAD.n8785 PAD.n2891 2.24164
R40091 PAD.n8821 PAD.n2940 2.24164
R40092 PAD.n8777 PAD.n2891 2.24164
R40093 PAD.n8821 PAD.n2939 2.24164
R40094 PAD.n8773 PAD.n2891 2.24164
R40095 PAD.n8821 PAD.n2938 2.24164
R40096 PAD.n8765 PAD.n2891 2.24164
R40097 PAD.n8821 PAD.n2937 2.24164
R40098 PAD.n8761 PAD.n2891 2.24164
R40099 PAD.n8821 PAD.n2936 2.24164
R40100 PAD.n8753 PAD.n2891 2.24164
R40101 PAD.n8821 PAD.n2935 2.24164
R40102 PAD.n8749 PAD.n2891 2.24164
R40103 PAD.n8821 PAD.n2934 2.24164
R40104 PAD.n8741 PAD.n2891 2.24164
R40105 PAD.n8821 PAD.n2933 2.24164
R40106 PAD.n8737 PAD.n2891 2.24164
R40107 PAD.n8821 PAD.n2932 2.24164
R40108 PAD.n8729 PAD.n2891 2.24164
R40109 PAD.n8821 PAD.n2931 2.24164
R40110 PAD.n8725 PAD.n2891 2.24164
R40111 PAD.n8821 PAD.n2930 2.24164
R40112 PAD.n8717 PAD.n2891 2.24164
R40113 PAD.n8821 PAD.n2929 2.24164
R40114 PAD.n8713 PAD.n2891 2.24164
R40115 PAD.n8821 PAD.n2928 2.24164
R40116 PAD.n8705 PAD.n2891 2.24164
R40117 PAD.n8821 PAD.n2927 2.24164
R40118 PAD.n8701 PAD.n2891 2.24164
R40119 PAD.n8821 PAD.n2926 2.24164
R40120 PAD.n8693 PAD.n2891 2.24164
R40121 PAD.n8821 PAD.n2925 2.24164
R40122 PAD.n8689 PAD.n2891 2.24164
R40123 PAD.n8821 PAD.n2924 2.24164
R40124 PAD.n8681 PAD.n2891 2.24164
R40125 PAD.n8821 PAD.n2923 2.24164
R40126 PAD.n8677 PAD.n2891 2.24164
R40127 PAD.n8821 PAD.n2922 2.24164
R40128 PAD.n8669 PAD.n2891 2.24164
R40129 PAD.n8821 PAD.n2921 2.24164
R40130 PAD.n8665 PAD.n2891 2.24164
R40131 PAD.n8821 PAD.n2920 2.24164
R40132 PAD.n8657 PAD.n2891 2.24164
R40133 PAD.n8821 PAD.n2919 2.24164
R40134 PAD.n8653 PAD.n2891 2.24164
R40135 PAD.n8821 PAD.n2918 2.24164
R40136 PAD.n8645 PAD.n2891 2.24164
R40137 PAD.n8821 PAD.n2917 2.24164
R40138 PAD.n8641 PAD.n2891 2.24164
R40139 PAD.n8821 PAD.n2916 2.24164
R40140 PAD.n8633 PAD.n2891 2.24164
R40141 PAD.n8821 PAD.n2915 2.24164
R40142 PAD.n8629 PAD.n2891 2.24164
R40143 PAD.n8821 PAD.n2914 2.24164
R40144 PAD.n8621 PAD.n2891 2.24164
R40145 PAD.n8821 PAD.n2913 2.24164
R40146 PAD.n8617 PAD.n2891 2.24164
R40147 PAD.n8821 PAD.n2912 2.24164
R40148 PAD.n8609 PAD.n2891 2.24164
R40149 PAD.n8821 PAD.n2911 2.24164
R40150 PAD.n8605 PAD.n2891 2.24164
R40151 PAD.n8821 PAD.n2910 2.24164
R40152 PAD.n8597 PAD.n2891 2.24164
R40153 PAD.n8821 PAD.n2909 2.24164
R40154 PAD.n8593 PAD.n2891 2.24164
R40155 PAD.n8821 PAD.n2908 2.24164
R40156 PAD.n8585 PAD.n2891 2.24164
R40157 PAD.n8821 PAD.n2907 2.24164
R40158 PAD.n8581 PAD.n2891 2.24164
R40159 PAD.n8821 PAD.n2906 2.24164
R40160 PAD.n8573 PAD.n2891 2.24164
R40161 PAD.n8821 PAD.n2905 2.24164
R40162 PAD.n3038 PAD.n2997 2.24164
R40163 PAD.n8517 PAD.n2993 2.24164
R40164 PAD.n3047 PAD.n2997 2.24164
R40165 PAD.n8517 PAD.n2992 2.24164
R40166 PAD.n3051 PAD.n2997 2.24164
R40167 PAD.n8517 PAD.n2991 2.24164
R40168 PAD.n3059 PAD.n2997 2.24164
R40169 PAD.n8517 PAD.n2990 2.24164
R40170 PAD.n3063 PAD.n2997 2.24164
R40171 PAD.n8517 PAD.n2989 2.24164
R40172 PAD.n3071 PAD.n2997 2.24164
R40173 PAD.n8517 PAD.n2988 2.24164
R40174 PAD.n3075 PAD.n2997 2.24164
R40175 PAD.n8517 PAD.n2987 2.24164
R40176 PAD.n3083 PAD.n2997 2.24164
R40177 PAD.n8517 PAD.n2986 2.24164
R40178 PAD.n3087 PAD.n2997 2.24164
R40179 PAD.n8517 PAD.n2985 2.24164
R40180 PAD.n3095 PAD.n2997 2.24164
R40181 PAD.n8517 PAD.n2984 2.24164
R40182 PAD.n3099 PAD.n2997 2.24164
R40183 PAD.n8517 PAD.n2983 2.24164
R40184 PAD.n3107 PAD.n2997 2.24164
R40185 PAD.n8517 PAD.n2982 2.24164
R40186 PAD.n3111 PAD.n2997 2.24164
R40187 PAD.n8517 PAD.n2981 2.24164
R40188 PAD.n3119 PAD.n2997 2.24164
R40189 PAD.n8517 PAD.n2980 2.24164
R40190 PAD.n3123 PAD.n2997 2.24164
R40191 PAD.n8517 PAD.n2979 2.24164
R40192 PAD.n3131 PAD.n2997 2.24164
R40193 PAD.n8517 PAD.n2978 2.24164
R40194 PAD.n3135 PAD.n2997 2.24164
R40195 PAD.n8517 PAD.n2977 2.24164
R40196 PAD.n3143 PAD.n2997 2.24164
R40197 PAD.n8517 PAD.n2976 2.24164
R40198 PAD.n3147 PAD.n2997 2.24164
R40199 PAD.n8517 PAD.n2975 2.24164
R40200 PAD.n3155 PAD.n2997 2.24164
R40201 PAD.n8517 PAD.n2974 2.24164
R40202 PAD.n3159 PAD.n2997 2.24164
R40203 PAD.n8517 PAD.n2973 2.24164
R40204 PAD.n3167 PAD.n2997 2.24164
R40205 PAD.n8517 PAD.n2972 2.24164
R40206 PAD.n3171 PAD.n2997 2.24164
R40207 PAD.n8517 PAD.n2971 2.24164
R40208 PAD.n3179 PAD.n2997 2.24164
R40209 PAD.n8517 PAD.n2970 2.24164
R40210 PAD.n3183 PAD.n2997 2.24164
R40211 PAD.n8517 PAD.n2969 2.24164
R40212 PAD.n3191 PAD.n2997 2.24164
R40213 PAD.n8517 PAD.n2968 2.24164
R40214 PAD.n3195 PAD.n2997 2.24164
R40215 PAD.n8517 PAD.n2967 2.24164
R40216 PAD.n3203 PAD.n2997 2.24164
R40217 PAD.n8517 PAD.n2966 2.24164
R40218 PAD.n3207 PAD.n2997 2.24164
R40219 PAD.n8517 PAD.n2965 2.24164
R40220 PAD.n3215 PAD.n2997 2.24164
R40221 PAD.n8517 PAD.n2964 2.24164
R40222 PAD.n3219 PAD.n2997 2.24164
R40223 PAD.n8517 PAD.n2963 2.24164
R40224 PAD.n3227 PAD.n2997 2.24164
R40225 PAD.n8517 PAD.n2962 2.24164
R40226 PAD.n3231 PAD.n2997 2.24164
R40227 PAD.n8517 PAD.n2961 2.24164
R40228 PAD.n3239 PAD.n2997 2.24164
R40229 PAD.n8517 PAD.n2960 2.24164
R40230 PAD.n3243 PAD.n2997 2.24164
R40231 PAD.n8517 PAD.n2959 2.24164
R40232 PAD.n3251 PAD.n2997 2.24164
R40233 PAD.n8517 PAD.n2958 2.24164
R40234 PAD.n3255 PAD.n2997 2.24164
R40235 PAD.n8517 PAD.n2957 2.24164
R40236 PAD.n3263 PAD.n2997 2.24164
R40237 PAD.n8517 PAD.n2956 2.24164
R40238 PAD.n3267 PAD.n2997 2.24164
R40239 PAD.n8517 PAD.n2955 2.24164
R40240 PAD.n3275 PAD.n2997 2.24164
R40241 PAD.n8517 PAD.n2954 2.24164
R40242 PAD.n3279 PAD.n2997 2.24164
R40243 PAD.n8517 PAD.n2953 2.24164
R40244 PAD.n8515 PAD.n2997 2.24164
R40245 PAD.n3383 PAD.n3342 2.24164
R40246 PAD.n8492 PAD.n3337 2.24164
R40247 PAD.n3392 PAD.n3342 2.24164
R40248 PAD.n8492 PAD.n3336 2.24164
R40249 PAD.n3396 PAD.n3342 2.24164
R40250 PAD.n8492 PAD.n3335 2.24164
R40251 PAD.n3404 PAD.n3342 2.24164
R40252 PAD.n8492 PAD.n3334 2.24164
R40253 PAD.n3408 PAD.n3342 2.24164
R40254 PAD.n8492 PAD.n3333 2.24164
R40255 PAD.n3416 PAD.n3342 2.24164
R40256 PAD.n8492 PAD.n3332 2.24164
R40257 PAD.n3420 PAD.n3342 2.24164
R40258 PAD.n8492 PAD.n3331 2.24164
R40259 PAD.n3428 PAD.n3342 2.24164
R40260 PAD.n8492 PAD.n3330 2.24164
R40261 PAD.n3432 PAD.n3342 2.24164
R40262 PAD.n8492 PAD.n3329 2.24164
R40263 PAD.n3440 PAD.n3342 2.24164
R40264 PAD.n8492 PAD.n3328 2.24164
R40265 PAD.n3444 PAD.n3342 2.24164
R40266 PAD.n8492 PAD.n3327 2.24164
R40267 PAD.n3452 PAD.n3342 2.24164
R40268 PAD.n8492 PAD.n3326 2.24164
R40269 PAD.n3456 PAD.n3342 2.24164
R40270 PAD.n8492 PAD.n3325 2.24164
R40271 PAD.n3464 PAD.n3342 2.24164
R40272 PAD.n8492 PAD.n3324 2.24164
R40273 PAD.n3468 PAD.n3342 2.24164
R40274 PAD.n8492 PAD.n3323 2.24164
R40275 PAD.n3476 PAD.n3342 2.24164
R40276 PAD.n8492 PAD.n3322 2.24164
R40277 PAD.n3480 PAD.n3342 2.24164
R40278 PAD.n8492 PAD.n3321 2.24164
R40279 PAD.n3488 PAD.n3342 2.24164
R40280 PAD.n8492 PAD.n3320 2.24164
R40281 PAD.n3492 PAD.n3342 2.24164
R40282 PAD.n8492 PAD.n3319 2.24164
R40283 PAD.n3500 PAD.n3342 2.24164
R40284 PAD.n8492 PAD.n3318 2.24164
R40285 PAD.n3504 PAD.n3342 2.24164
R40286 PAD.n8492 PAD.n3317 2.24164
R40287 PAD.n3512 PAD.n3342 2.24164
R40288 PAD.n8492 PAD.n3316 2.24164
R40289 PAD.n3516 PAD.n3342 2.24164
R40290 PAD.n8492 PAD.n3315 2.24164
R40291 PAD.n3524 PAD.n3342 2.24164
R40292 PAD.n8492 PAD.n3314 2.24164
R40293 PAD.n3528 PAD.n3342 2.24164
R40294 PAD.n8492 PAD.n3313 2.24164
R40295 PAD.n3536 PAD.n3342 2.24164
R40296 PAD.n8492 PAD.n3312 2.24164
R40297 PAD.n3540 PAD.n3342 2.24164
R40298 PAD.n8492 PAD.n3311 2.24164
R40299 PAD.n3548 PAD.n3342 2.24164
R40300 PAD.n8492 PAD.n3310 2.24164
R40301 PAD.n3552 PAD.n3342 2.24164
R40302 PAD.n8492 PAD.n3309 2.24164
R40303 PAD.n3560 PAD.n3342 2.24164
R40304 PAD.n8492 PAD.n3308 2.24164
R40305 PAD.n3564 PAD.n3342 2.24164
R40306 PAD.n8492 PAD.n3307 2.24164
R40307 PAD.n3572 PAD.n3342 2.24164
R40308 PAD.n8492 PAD.n3306 2.24164
R40309 PAD.n3576 PAD.n3342 2.24164
R40310 PAD.n8492 PAD.n3305 2.24164
R40311 PAD.n3584 PAD.n3342 2.24164
R40312 PAD.n8492 PAD.n3304 2.24164
R40313 PAD.n3588 PAD.n3342 2.24164
R40314 PAD.n8492 PAD.n3303 2.24164
R40315 PAD.n3596 PAD.n3342 2.24164
R40316 PAD.n8492 PAD.n3302 2.24164
R40317 PAD.n3600 PAD.n3342 2.24164
R40318 PAD.n8492 PAD.n3301 2.24164
R40319 PAD.n3608 PAD.n3342 2.24164
R40320 PAD.n8492 PAD.n3300 2.24164
R40321 PAD.n3612 PAD.n3342 2.24164
R40322 PAD.n8492 PAD.n3299 2.24164
R40323 PAD.n3620 PAD.n3342 2.24164
R40324 PAD.n8492 PAD.n3298 2.24164
R40325 PAD.n3624 PAD.n3342 2.24164
R40326 PAD.n8492 PAD.n3297 2.24164
R40327 PAD.n8490 PAD.n3342 2.24164
R40328 PAD.n3728 PAD.n3687 2.24164
R40329 PAD.n8468 PAD.n3682 2.24164
R40330 PAD.n3737 PAD.n3687 2.24164
R40331 PAD.n8468 PAD.n3681 2.24164
R40332 PAD.n3741 PAD.n3687 2.24164
R40333 PAD.n8468 PAD.n3680 2.24164
R40334 PAD.n3749 PAD.n3687 2.24164
R40335 PAD.n8468 PAD.n3679 2.24164
R40336 PAD.n3753 PAD.n3687 2.24164
R40337 PAD.n8468 PAD.n3678 2.24164
R40338 PAD.n3761 PAD.n3687 2.24164
R40339 PAD.n8468 PAD.n3677 2.24164
R40340 PAD.n3765 PAD.n3687 2.24164
R40341 PAD.n8468 PAD.n3676 2.24164
R40342 PAD.n3773 PAD.n3687 2.24164
R40343 PAD.n8468 PAD.n3675 2.24164
R40344 PAD.n3777 PAD.n3687 2.24164
R40345 PAD.n8468 PAD.n3674 2.24164
R40346 PAD.n3785 PAD.n3687 2.24164
R40347 PAD.n8468 PAD.n3673 2.24164
R40348 PAD.n3789 PAD.n3687 2.24164
R40349 PAD.n8468 PAD.n3672 2.24164
R40350 PAD.n3797 PAD.n3687 2.24164
R40351 PAD.n8468 PAD.n3671 2.24164
R40352 PAD.n3801 PAD.n3687 2.24164
R40353 PAD.n8468 PAD.n3670 2.24164
R40354 PAD.n3809 PAD.n3687 2.24164
R40355 PAD.n8468 PAD.n3669 2.24164
R40356 PAD.n3813 PAD.n3687 2.24164
R40357 PAD.n8468 PAD.n3668 2.24164
R40358 PAD.n3821 PAD.n3687 2.24164
R40359 PAD.n8468 PAD.n3667 2.24164
R40360 PAD.n3825 PAD.n3687 2.24164
R40361 PAD.n8468 PAD.n3666 2.24164
R40362 PAD.n3833 PAD.n3687 2.24164
R40363 PAD.n8468 PAD.n3665 2.24164
R40364 PAD.n3837 PAD.n3687 2.24164
R40365 PAD.n8468 PAD.n3664 2.24164
R40366 PAD.n3845 PAD.n3687 2.24164
R40367 PAD.n8468 PAD.n3663 2.24164
R40368 PAD.n3849 PAD.n3687 2.24164
R40369 PAD.n8468 PAD.n3662 2.24164
R40370 PAD.n3857 PAD.n3687 2.24164
R40371 PAD.n8468 PAD.n3661 2.24164
R40372 PAD.n3861 PAD.n3687 2.24164
R40373 PAD.n8468 PAD.n3660 2.24164
R40374 PAD.n3869 PAD.n3687 2.24164
R40375 PAD.n8468 PAD.n3659 2.24164
R40376 PAD.n3873 PAD.n3687 2.24164
R40377 PAD.n8468 PAD.n3658 2.24164
R40378 PAD.n3881 PAD.n3687 2.24164
R40379 PAD.n8468 PAD.n3657 2.24164
R40380 PAD.n3885 PAD.n3687 2.24164
R40381 PAD.n8468 PAD.n3656 2.24164
R40382 PAD.n3893 PAD.n3687 2.24164
R40383 PAD.n8468 PAD.n3655 2.24164
R40384 PAD.n3897 PAD.n3687 2.24164
R40385 PAD.n8468 PAD.n3654 2.24164
R40386 PAD.n3905 PAD.n3687 2.24164
R40387 PAD.n8468 PAD.n3653 2.24164
R40388 PAD.n3909 PAD.n3687 2.24164
R40389 PAD.n8468 PAD.n3652 2.24164
R40390 PAD.n3917 PAD.n3687 2.24164
R40391 PAD.n8468 PAD.n3651 2.24164
R40392 PAD.n3921 PAD.n3687 2.24164
R40393 PAD.n8468 PAD.n3650 2.24164
R40394 PAD.n3929 PAD.n3687 2.24164
R40395 PAD.n8468 PAD.n3649 2.24164
R40396 PAD.n3933 PAD.n3687 2.24164
R40397 PAD.n8468 PAD.n3648 2.24164
R40398 PAD.n3941 PAD.n3687 2.24164
R40399 PAD.n8468 PAD.n3647 2.24164
R40400 PAD.n3945 PAD.n3687 2.24164
R40401 PAD.n8468 PAD.n3646 2.24164
R40402 PAD.n3953 PAD.n3687 2.24164
R40403 PAD.n8468 PAD.n3645 2.24164
R40404 PAD.n3957 PAD.n3687 2.24164
R40405 PAD.n8468 PAD.n3644 2.24164
R40406 PAD.n3965 PAD.n3687 2.24164
R40407 PAD.n8468 PAD.n3643 2.24164
R40408 PAD.n3969 PAD.n3687 2.24164
R40409 PAD.n8468 PAD.n3642 2.24164
R40410 PAD.n8466 PAD.n3687 2.24164
R40411 PAD.n4069 PAD.n4028 2.24164
R40412 PAD.n8444 PAD.n4024 2.24164
R40413 PAD.n4078 PAD.n4028 2.24164
R40414 PAD.n8444 PAD.n4023 2.24164
R40415 PAD.n4082 PAD.n4028 2.24164
R40416 PAD.n8444 PAD.n4022 2.24164
R40417 PAD.n4090 PAD.n4028 2.24164
R40418 PAD.n8444 PAD.n4021 2.24164
R40419 PAD.n4094 PAD.n4028 2.24164
R40420 PAD.n8444 PAD.n4020 2.24164
R40421 PAD.n4102 PAD.n4028 2.24164
R40422 PAD.n8444 PAD.n4019 2.24164
R40423 PAD.n4106 PAD.n4028 2.24164
R40424 PAD.n8444 PAD.n4018 2.24164
R40425 PAD.n4114 PAD.n4028 2.24164
R40426 PAD.n8444 PAD.n4017 2.24164
R40427 PAD.n4118 PAD.n4028 2.24164
R40428 PAD.n8444 PAD.n4016 2.24164
R40429 PAD.n4126 PAD.n4028 2.24164
R40430 PAD.n8444 PAD.n4015 2.24164
R40431 PAD.n4130 PAD.n4028 2.24164
R40432 PAD.n8444 PAD.n4014 2.24164
R40433 PAD.n4138 PAD.n4028 2.24164
R40434 PAD.n8444 PAD.n4013 2.24164
R40435 PAD.n4142 PAD.n4028 2.24164
R40436 PAD.n8444 PAD.n4012 2.24164
R40437 PAD.n4150 PAD.n4028 2.24164
R40438 PAD.n8444 PAD.n4011 2.24164
R40439 PAD.n4154 PAD.n4028 2.24164
R40440 PAD.n8444 PAD.n4010 2.24164
R40441 PAD.n4162 PAD.n4028 2.24164
R40442 PAD.n8444 PAD.n4009 2.24164
R40443 PAD.n4166 PAD.n4028 2.24164
R40444 PAD.n8444 PAD.n4008 2.24164
R40445 PAD.n4174 PAD.n4028 2.24164
R40446 PAD.n8444 PAD.n4007 2.24164
R40447 PAD.n4178 PAD.n4028 2.24164
R40448 PAD.n8444 PAD.n4006 2.24164
R40449 PAD.n4186 PAD.n4028 2.24164
R40450 PAD.n8444 PAD.n4005 2.24164
R40451 PAD.n4190 PAD.n4028 2.24164
R40452 PAD.n8444 PAD.n4004 2.24164
R40453 PAD.n4198 PAD.n4028 2.24164
R40454 PAD.n8444 PAD.n4003 2.24164
R40455 PAD.n4202 PAD.n4028 2.24164
R40456 PAD.n8444 PAD.n4002 2.24164
R40457 PAD.n4210 PAD.n4028 2.24164
R40458 PAD.n8444 PAD.n4001 2.24164
R40459 PAD.n4214 PAD.n4028 2.24164
R40460 PAD.n8444 PAD.n4000 2.24164
R40461 PAD.n4222 PAD.n4028 2.24164
R40462 PAD.n8444 PAD.n3999 2.24164
R40463 PAD.n4226 PAD.n4028 2.24164
R40464 PAD.n8444 PAD.n3998 2.24164
R40465 PAD.n4234 PAD.n4028 2.24164
R40466 PAD.n8444 PAD.n3997 2.24164
R40467 PAD.n4238 PAD.n4028 2.24164
R40468 PAD.n8444 PAD.n3996 2.24164
R40469 PAD.n4246 PAD.n4028 2.24164
R40470 PAD.n8444 PAD.n3995 2.24164
R40471 PAD.n4250 PAD.n4028 2.24164
R40472 PAD.n8444 PAD.n3994 2.24164
R40473 PAD.n4258 PAD.n4028 2.24164
R40474 PAD.n8444 PAD.n3993 2.24164
R40475 PAD.n4262 PAD.n4028 2.24164
R40476 PAD.n8444 PAD.n3992 2.24164
R40477 PAD.n4270 PAD.n4028 2.24164
R40478 PAD.n8444 PAD.n3991 2.24164
R40479 PAD.n4274 PAD.n4028 2.24164
R40480 PAD.n8444 PAD.n3990 2.24164
R40481 PAD.n4282 PAD.n4028 2.24164
R40482 PAD.n8444 PAD.n3989 2.24164
R40483 PAD.n4286 PAD.n4028 2.24164
R40484 PAD.n8444 PAD.n3988 2.24164
R40485 PAD.n4294 PAD.n4028 2.24164
R40486 PAD.n8444 PAD.n3987 2.24164
R40487 PAD.n4298 PAD.n4028 2.24164
R40488 PAD.n8444 PAD.n3986 2.24164
R40489 PAD.n4306 PAD.n4028 2.24164
R40490 PAD.n8444 PAD.n3985 2.24164
R40491 PAD.n4310 PAD.n4028 2.24164
R40492 PAD.n8444 PAD.n3984 2.24164
R40493 PAD.n8442 PAD.n4028 2.24164
R40494 PAD.n4421 PAD.n4331 2.24164
R40495 PAD.n4423 PAD.n4333 2.24164
R40496 PAD.n4425 PAD.n4331 2.24164
R40497 PAD.n4415 PAD.n4333 2.24164
R40498 PAD.n4433 PAD.n4331 2.24164
R40499 PAD.n4435 PAD.n4333 2.24164
R40500 PAD.n4437 PAD.n4331 2.24164
R40501 PAD.n4411 PAD.n4333 2.24164
R40502 PAD.n4445 PAD.n4331 2.24164
R40503 PAD.n4447 PAD.n4333 2.24164
R40504 PAD.n4449 PAD.n4331 2.24164
R40505 PAD.n4407 PAD.n4333 2.24164
R40506 PAD.n4457 PAD.n4331 2.24164
R40507 PAD.n4459 PAD.n4333 2.24164
R40508 PAD.n4461 PAD.n4331 2.24164
R40509 PAD.n4403 PAD.n4333 2.24164
R40510 PAD.n4469 PAD.n4331 2.24164
R40511 PAD.n4471 PAD.n4333 2.24164
R40512 PAD.n4473 PAD.n4331 2.24164
R40513 PAD.n4399 PAD.n4333 2.24164
R40514 PAD.n4481 PAD.n4331 2.24164
R40515 PAD.n4483 PAD.n4333 2.24164
R40516 PAD.n4485 PAD.n4331 2.24164
R40517 PAD.n4395 PAD.n4333 2.24164
R40518 PAD.n4493 PAD.n4331 2.24164
R40519 PAD.n4495 PAD.n4333 2.24164
R40520 PAD.n4497 PAD.n4331 2.24164
R40521 PAD.n4391 PAD.n4333 2.24164
R40522 PAD.n4505 PAD.n4331 2.24164
R40523 PAD.n4507 PAD.n4333 2.24164
R40524 PAD.n4509 PAD.n4331 2.24164
R40525 PAD.n4387 PAD.n4333 2.24164
R40526 PAD.n4517 PAD.n4331 2.24164
R40527 PAD.n4519 PAD.n4333 2.24164
R40528 PAD.n4521 PAD.n4331 2.24164
R40529 PAD.n4383 PAD.n4333 2.24164
R40530 PAD.n4529 PAD.n4331 2.24164
R40531 PAD.n4531 PAD.n4333 2.24164
R40532 PAD.n4533 PAD.n4331 2.24164
R40533 PAD.n4379 PAD.n4333 2.24164
R40534 PAD.n4541 PAD.n4331 2.24164
R40535 PAD.n4543 PAD.n4333 2.24164
R40536 PAD.n4545 PAD.n4331 2.24164
R40537 PAD.n4375 PAD.n4333 2.24164
R40538 PAD.n4553 PAD.n4331 2.24164
R40539 PAD.n4555 PAD.n4333 2.24164
R40540 PAD.n4557 PAD.n4331 2.24164
R40541 PAD.n4371 PAD.n4333 2.24164
R40542 PAD.n4565 PAD.n4331 2.24164
R40543 PAD.n4567 PAD.n4333 2.24164
R40544 PAD.n4569 PAD.n4331 2.24164
R40545 PAD.n4367 PAD.n4333 2.24164
R40546 PAD.n4577 PAD.n4331 2.24164
R40547 PAD.n4579 PAD.n4333 2.24164
R40548 PAD.n4581 PAD.n4331 2.24164
R40549 PAD.n4363 PAD.n4333 2.24164
R40550 PAD.n4589 PAD.n4331 2.24164
R40551 PAD.n4591 PAD.n4333 2.24164
R40552 PAD.n4593 PAD.n4331 2.24164
R40553 PAD.n4359 PAD.n4333 2.24164
R40554 PAD.n4601 PAD.n4331 2.24164
R40555 PAD.n4603 PAD.n4333 2.24164
R40556 PAD.n4605 PAD.n4331 2.24164
R40557 PAD.n4355 PAD.n4333 2.24164
R40558 PAD.n4613 PAD.n4331 2.24164
R40559 PAD.n4615 PAD.n4333 2.24164
R40560 PAD.n4617 PAD.n4331 2.24164
R40561 PAD.n4351 PAD.n4333 2.24164
R40562 PAD.n4625 PAD.n4331 2.24164
R40563 PAD.n4627 PAD.n4333 2.24164
R40564 PAD.n4629 PAD.n4331 2.24164
R40565 PAD.n4347 PAD.n4333 2.24164
R40566 PAD.n4637 PAD.n4331 2.24164
R40567 PAD.n4639 PAD.n4333 2.24164
R40568 PAD.n4641 PAD.n4331 2.24164
R40569 PAD.n4343 PAD.n4333 2.24164
R40570 PAD.n4649 PAD.n4331 2.24164
R40571 PAD.n4651 PAD.n4333 2.24164
R40572 PAD.n4653 PAD.n4331 2.24164
R40573 PAD.n4339 PAD.n4333 2.24164
R40574 PAD.n4662 PAD.n4331 2.24164
R40575 PAD.n4664 PAD.n4333 2.24164
R40576 PAD.n4666 PAD.n4331 2.24164
R40577 PAD.n8397 PAD.n8396 2.24164
R40578 PAD.n4726 PAD.n4673 2.24164
R40579 PAD.n8397 PAD.n4723 2.24164
R40580 PAD.n8387 PAD.n4673 2.24164
R40581 PAD.n8397 PAD.n4722 2.24164
R40582 PAD.n4732 PAD.n4673 2.24164
R40583 PAD.n8397 PAD.n4721 2.24164
R40584 PAD.n8378 PAD.n4673 2.24164
R40585 PAD.n8397 PAD.n4720 2.24164
R40586 PAD.n4737 PAD.n4673 2.24164
R40587 PAD.n8397 PAD.n4719 2.24164
R40588 PAD.n8369 PAD.n4673 2.24164
R40589 PAD.n8397 PAD.n4718 2.24164
R40590 PAD.n4742 PAD.n4673 2.24164
R40591 PAD.n8397 PAD.n4717 2.24164
R40592 PAD.n8360 PAD.n4673 2.24164
R40593 PAD.n8397 PAD.n4716 2.24164
R40594 PAD.n4747 PAD.n4673 2.24164
R40595 PAD.n8397 PAD.n4715 2.24164
R40596 PAD.n8351 PAD.n4673 2.24164
R40597 PAD.n8397 PAD.n4714 2.24164
R40598 PAD.n4752 PAD.n4673 2.24164
R40599 PAD.n8397 PAD.n4713 2.24164
R40600 PAD.n8342 PAD.n4673 2.24164
R40601 PAD.n8397 PAD.n4712 2.24164
R40602 PAD.n4757 PAD.n4673 2.24164
R40603 PAD.n8397 PAD.n4711 2.24164
R40604 PAD.n8333 PAD.n4673 2.24164
R40605 PAD.n8397 PAD.n4710 2.24164
R40606 PAD.n4762 PAD.n4673 2.24164
R40607 PAD.n8397 PAD.n4709 2.24164
R40608 PAD.n8324 PAD.n4673 2.24164
R40609 PAD.n8397 PAD.n4708 2.24164
R40610 PAD.n4767 PAD.n4673 2.24164
R40611 PAD.n8397 PAD.n4707 2.24164
R40612 PAD.n8315 PAD.n4673 2.24164
R40613 PAD.n8397 PAD.n4706 2.24164
R40614 PAD.n4772 PAD.n4673 2.24164
R40615 PAD.n8397 PAD.n4705 2.24164
R40616 PAD.n8306 PAD.n4673 2.24164
R40617 PAD.n8397 PAD.n4704 2.24164
R40618 PAD.n4777 PAD.n4673 2.24164
R40619 PAD.n8397 PAD.n4703 2.24164
R40620 PAD.n8297 PAD.n4673 2.24164
R40621 PAD.n8397 PAD.n4702 2.24164
R40622 PAD.n4782 PAD.n4673 2.24164
R40623 PAD.n8397 PAD.n4701 2.24164
R40624 PAD.n8288 PAD.n4673 2.24164
R40625 PAD.n8397 PAD.n4700 2.24164
R40626 PAD.n4787 PAD.n4673 2.24164
R40627 PAD.n8397 PAD.n4699 2.24164
R40628 PAD.n8279 PAD.n4673 2.24164
R40629 PAD.n8397 PAD.n4698 2.24164
R40630 PAD.n4792 PAD.n4673 2.24164
R40631 PAD.n8397 PAD.n4697 2.24164
R40632 PAD.n8270 PAD.n4673 2.24164
R40633 PAD.n8397 PAD.n4696 2.24164
R40634 PAD.n4797 PAD.n4673 2.24164
R40635 PAD.n8397 PAD.n4695 2.24164
R40636 PAD.n8261 PAD.n4673 2.24164
R40637 PAD.n8397 PAD.n4694 2.24164
R40638 PAD.n4802 PAD.n4673 2.24164
R40639 PAD.n8397 PAD.n4693 2.24164
R40640 PAD.n8252 PAD.n4673 2.24164
R40641 PAD.n8397 PAD.n4692 2.24164
R40642 PAD.n4807 PAD.n4673 2.24164
R40643 PAD.n8397 PAD.n4691 2.24164
R40644 PAD.n8243 PAD.n4673 2.24164
R40645 PAD.n8397 PAD.n4690 2.24164
R40646 PAD.n4812 PAD.n4673 2.24164
R40647 PAD.n8397 PAD.n4689 2.24164
R40648 PAD.n8234 PAD.n4673 2.24164
R40649 PAD.n8397 PAD.n4688 2.24164
R40650 PAD.n4817 PAD.n4673 2.24164
R40651 PAD.n8397 PAD.n4687 2.24164
R40652 PAD.n8225 PAD.n4673 2.24164
R40653 PAD.n8397 PAD.n4686 2.24164
R40654 PAD.n4822 PAD.n4673 2.24164
R40655 PAD.n8397 PAD.n4685 2.24164
R40656 PAD.n8216 PAD.n4673 2.24164
R40657 PAD.n8397 PAD.n4684 2.24164
R40658 PAD.n4827 PAD.n4673 2.24164
R40659 PAD.n8397 PAD.n4683 2.24164
R40660 PAD.n4849 PAD.n4840 2.24164
R40661 PAD.n5175 PAD.n4843 2.24164
R40662 PAD.n5173 PAD.n4840 2.24164
R40663 PAD.n4850 PAD.n4843 2.24164
R40664 PAD.n5165 PAD.n4840 2.24164
R40665 PAD.n5163 PAD.n4843 2.24164
R40666 PAD.n5161 PAD.n4840 2.24164
R40667 PAD.n4855 PAD.n4843 2.24164
R40668 PAD.n5153 PAD.n4840 2.24164
R40669 PAD.n5151 PAD.n4843 2.24164
R40670 PAD.n5149 PAD.n4840 2.24164
R40671 PAD.n4859 PAD.n4843 2.24164
R40672 PAD.n5141 PAD.n4840 2.24164
R40673 PAD.n5139 PAD.n4843 2.24164
R40674 PAD.n5137 PAD.n4840 2.24164
R40675 PAD.n4863 PAD.n4843 2.24164
R40676 PAD.n5129 PAD.n4840 2.24164
R40677 PAD.n5127 PAD.n4843 2.24164
R40678 PAD.n5125 PAD.n4840 2.24164
R40679 PAD.n4867 PAD.n4843 2.24164
R40680 PAD.n5117 PAD.n4840 2.24164
R40681 PAD.n5115 PAD.n4843 2.24164
R40682 PAD.n5113 PAD.n4840 2.24164
R40683 PAD.n4871 PAD.n4843 2.24164
R40684 PAD.n5105 PAD.n4840 2.24164
R40685 PAD.n5103 PAD.n4843 2.24164
R40686 PAD.n5101 PAD.n4840 2.24164
R40687 PAD.n4875 PAD.n4843 2.24164
R40688 PAD.n5093 PAD.n4840 2.24164
R40689 PAD.n5091 PAD.n4843 2.24164
R40690 PAD.n5089 PAD.n4840 2.24164
R40691 PAD.n4879 PAD.n4843 2.24164
R40692 PAD.n5081 PAD.n4840 2.24164
R40693 PAD.n5079 PAD.n4843 2.24164
R40694 PAD.n5077 PAD.n4840 2.24164
R40695 PAD.n4883 PAD.n4843 2.24164
R40696 PAD.n5069 PAD.n4840 2.24164
R40697 PAD.n5067 PAD.n4843 2.24164
R40698 PAD.n5065 PAD.n4840 2.24164
R40699 PAD.n4887 PAD.n4843 2.24164
R40700 PAD.n5057 PAD.n4840 2.24164
R40701 PAD.n5055 PAD.n4843 2.24164
R40702 PAD.n5053 PAD.n4840 2.24164
R40703 PAD.n4891 PAD.n4843 2.24164
R40704 PAD.n5045 PAD.n4840 2.24164
R40705 PAD.n5043 PAD.n4843 2.24164
R40706 PAD.n5041 PAD.n4840 2.24164
R40707 PAD.n4895 PAD.n4843 2.24164
R40708 PAD.n5033 PAD.n4840 2.24164
R40709 PAD.n5031 PAD.n4843 2.24164
R40710 PAD.n5029 PAD.n4840 2.24164
R40711 PAD.n4899 PAD.n4843 2.24164
R40712 PAD.n5021 PAD.n4840 2.24164
R40713 PAD.n5019 PAD.n4843 2.24164
R40714 PAD.n5017 PAD.n4840 2.24164
R40715 PAD.n4903 PAD.n4843 2.24164
R40716 PAD.n5009 PAD.n4840 2.24164
R40717 PAD.n5007 PAD.n4843 2.24164
R40718 PAD.n5005 PAD.n4840 2.24164
R40719 PAD.n4907 PAD.n4843 2.24164
R40720 PAD.n4997 PAD.n4840 2.24164
R40721 PAD.n4995 PAD.n4843 2.24164
R40722 PAD.n4993 PAD.n4840 2.24164
R40723 PAD.n4911 PAD.n4843 2.24164
R40724 PAD.n4985 PAD.n4840 2.24164
R40725 PAD.n4983 PAD.n4843 2.24164
R40726 PAD.n4981 PAD.n4840 2.24164
R40727 PAD.n4915 PAD.n4843 2.24164
R40728 PAD.n4973 PAD.n4840 2.24164
R40729 PAD.n4971 PAD.n4843 2.24164
R40730 PAD.n4969 PAD.n4840 2.24164
R40731 PAD.n4919 PAD.n4843 2.24164
R40732 PAD.n4961 PAD.n4840 2.24164
R40733 PAD.n4959 PAD.n4843 2.24164
R40734 PAD.n4957 PAD.n4840 2.24164
R40735 PAD.n4923 PAD.n4843 2.24164
R40736 PAD.n4949 PAD.n4840 2.24164
R40737 PAD.n4947 PAD.n4843 2.24164
R40738 PAD.n4945 PAD.n4840 2.24164
R40739 PAD.n4927 PAD.n4843 2.24164
R40740 PAD.n4937 PAD.n4840 2.24164
R40741 PAD.n4935 PAD.n4843 2.24164
R40742 PAD.n4933 PAD.n4840 2.24164
R40743 PAD.n8163 PAD.n8162 2.24164
R40744 PAD.n7872 PAD.n5183 2.24164
R40745 PAD.n8163 PAD.n7870 2.24164
R40746 PAD.n8153 PAD.n5183 2.24164
R40747 PAD.n8163 PAD.n7869 2.24164
R40748 PAD.n7878 PAD.n5183 2.24164
R40749 PAD.n8163 PAD.n7868 2.24164
R40750 PAD.n8144 PAD.n5183 2.24164
R40751 PAD.n8163 PAD.n7867 2.24164
R40752 PAD.n7883 PAD.n5183 2.24164
R40753 PAD.n8163 PAD.n7866 2.24164
R40754 PAD.n8135 PAD.n5183 2.24164
R40755 PAD.n8163 PAD.n7865 2.24164
R40756 PAD.n7888 PAD.n5183 2.24164
R40757 PAD.n8163 PAD.n7864 2.24164
R40758 PAD.n8126 PAD.n5183 2.24164
R40759 PAD.n8163 PAD.n7863 2.24164
R40760 PAD.n7893 PAD.n5183 2.24164
R40761 PAD.n8163 PAD.n7862 2.24164
R40762 PAD.n8117 PAD.n5183 2.24164
R40763 PAD.n8163 PAD.n7861 2.24164
R40764 PAD.n7898 PAD.n5183 2.24164
R40765 PAD.n8163 PAD.n7860 2.24164
R40766 PAD.n8108 PAD.n5183 2.24164
R40767 PAD.n8163 PAD.n7859 2.24164
R40768 PAD.n7903 PAD.n5183 2.24164
R40769 PAD.n8163 PAD.n7858 2.24164
R40770 PAD.n8099 PAD.n5183 2.24164
R40771 PAD.n8163 PAD.n7857 2.24164
R40772 PAD.n7908 PAD.n5183 2.24164
R40773 PAD.n8163 PAD.n7856 2.24164
R40774 PAD.n8090 PAD.n5183 2.24164
R40775 PAD.n8163 PAD.n7855 2.24164
R40776 PAD.n7913 PAD.n5183 2.24164
R40777 PAD.n8163 PAD.n7854 2.24164
R40778 PAD.n8081 PAD.n5183 2.24164
R40779 PAD.n8163 PAD.n7853 2.24164
R40780 PAD.n7918 PAD.n5183 2.24164
R40781 PAD.n8163 PAD.n7852 2.24164
R40782 PAD.n8072 PAD.n5183 2.24164
R40783 PAD.n8163 PAD.n7851 2.24164
R40784 PAD.n7923 PAD.n5183 2.24164
R40785 PAD.n8163 PAD.n7850 2.24164
R40786 PAD.n8063 PAD.n5183 2.24164
R40787 PAD.n8163 PAD.n7849 2.24164
R40788 PAD.n7928 PAD.n5183 2.24164
R40789 PAD.n8163 PAD.n7848 2.24164
R40790 PAD.n8054 PAD.n5183 2.24164
R40791 PAD.n8163 PAD.n7847 2.24164
R40792 PAD.n7933 PAD.n5183 2.24164
R40793 PAD.n8163 PAD.n7846 2.24164
R40794 PAD.n8045 PAD.n5183 2.24164
R40795 PAD.n8163 PAD.n7845 2.24164
R40796 PAD.n7938 PAD.n5183 2.24164
R40797 PAD.n8163 PAD.n7844 2.24164
R40798 PAD.n8036 PAD.n5183 2.24164
R40799 PAD.n8163 PAD.n7843 2.24164
R40800 PAD.n7943 PAD.n5183 2.24164
R40801 PAD.n8163 PAD.n7842 2.24164
R40802 PAD.n8027 PAD.n5183 2.24164
R40803 PAD.n8163 PAD.n7841 2.24164
R40804 PAD.n7948 PAD.n5183 2.24164
R40805 PAD.n8163 PAD.n7840 2.24164
R40806 PAD.n8018 PAD.n5183 2.24164
R40807 PAD.n8163 PAD.n7839 2.24164
R40808 PAD.n7953 PAD.n5183 2.24164
R40809 PAD.n8163 PAD.n7838 2.24164
R40810 PAD.n8009 PAD.n5183 2.24164
R40811 PAD.n8163 PAD.n7837 2.24164
R40812 PAD.n7958 PAD.n5183 2.24164
R40813 PAD.n8163 PAD.n7836 2.24164
R40814 PAD.n8000 PAD.n5183 2.24164
R40815 PAD.n8163 PAD.n7835 2.24164
R40816 PAD.n7963 PAD.n5183 2.24164
R40817 PAD.n8163 PAD.n7834 2.24164
R40818 PAD.n7991 PAD.n5183 2.24164
R40819 PAD.n8163 PAD.n7833 2.24164
R40820 PAD.n7968 PAD.n5183 2.24164
R40821 PAD.n8163 PAD.n7832 2.24164
R40822 PAD.n7982 PAD.n5183 2.24164
R40823 PAD.n8163 PAD.n7831 2.24164
R40824 PAD.n7975 PAD.n5183 2.24164
R40825 PAD.n8163 PAD.n7830 2.24164
R40826 PAD.n5213 PAD.n5204 2.24164
R40827 PAD.n5539 PAD.n5197 2.24164
R40828 PAD.n5537 PAD.n5204 2.24164
R40829 PAD.n5214 PAD.n5197 2.24164
R40830 PAD.n5529 PAD.n5204 2.24164
R40831 PAD.n5527 PAD.n5197 2.24164
R40832 PAD.n5525 PAD.n5204 2.24164
R40833 PAD.n5219 PAD.n5197 2.24164
R40834 PAD.n5517 PAD.n5204 2.24164
R40835 PAD.n5515 PAD.n5197 2.24164
R40836 PAD.n5513 PAD.n5204 2.24164
R40837 PAD.n5223 PAD.n5197 2.24164
R40838 PAD.n5505 PAD.n5204 2.24164
R40839 PAD.n5503 PAD.n5197 2.24164
R40840 PAD.n5501 PAD.n5204 2.24164
R40841 PAD.n5227 PAD.n5197 2.24164
R40842 PAD.n5493 PAD.n5204 2.24164
R40843 PAD.n5491 PAD.n5197 2.24164
R40844 PAD.n5489 PAD.n5204 2.24164
R40845 PAD.n5231 PAD.n5197 2.24164
R40846 PAD.n5481 PAD.n5204 2.24164
R40847 PAD.n5479 PAD.n5197 2.24164
R40848 PAD.n5477 PAD.n5204 2.24164
R40849 PAD.n5235 PAD.n5197 2.24164
R40850 PAD.n5469 PAD.n5204 2.24164
R40851 PAD.n5467 PAD.n5197 2.24164
R40852 PAD.n5465 PAD.n5204 2.24164
R40853 PAD.n5239 PAD.n5197 2.24164
R40854 PAD.n5457 PAD.n5204 2.24164
R40855 PAD.n5455 PAD.n5197 2.24164
R40856 PAD.n5453 PAD.n5204 2.24164
R40857 PAD.n5243 PAD.n5197 2.24164
R40858 PAD.n5445 PAD.n5204 2.24164
R40859 PAD.n5443 PAD.n5197 2.24164
R40860 PAD.n5441 PAD.n5204 2.24164
R40861 PAD.n5247 PAD.n5197 2.24164
R40862 PAD.n5433 PAD.n5204 2.24164
R40863 PAD.n5431 PAD.n5197 2.24164
R40864 PAD.n5429 PAD.n5204 2.24164
R40865 PAD.n5251 PAD.n5197 2.24164
R40866 PAD.n5421 PAD.n5204 2.24164
R40867 PAD.n5419 PAD.n5197 2.24164
R40868 PAD.n5417 PAD.n5204 2.24164
R40869 PAD.n5255 PAD.n5197 2.24164
R40870 PAD.n5409 PAD.n5204 2.24164
R40871 PAD.n5407 PAD.n5197 2.24164
R40872 PAD.n5405 PAD.n5204 2.24164
R40873 PAD.n5259 PAD.n5197 2.24164
R40874 PAD.n5397 PAD.n5204 2.24164
R40875 PAD.n5395 PAD.n5197 2.24164
R40876 PAD.n5393 PAD.n5204 2.24164
R40877 PAD.n5263 PAD.n5197 2.24164
R40878 PAD.n5385 PAD.n5204 2.24164
R40879 PAD.n5383 PAD.n5197 2.24164
R40880 PAD.n5381 PAD.n5204 2.24164
R40881 PAD.n5267 PAD.n5197 2.24164
R40882 PAD.n5373 PAD.n5204 2.24164
R40883 PAD.n5371 PAD.n5197 2.24164
R40884 PAD.n5369 PAD.n5204 2.24164
R40885 PAD.n5271 PAD.n5197 2.24164
R40886 PAD.n5361 PAD.n5204 2.24164
R40887 PAD.n5359 PAD.n5197 2.24164
R40888 PAD.n5357 PAD.n5204 2.24164
R40889 PAD.n5275 PAD.n5197 2.24164
R40890 PAD.n5349 PAD.n5204 2.24164
R40891 PAD.n5347 PAD.n5197 2.24164
R40892 PAD.n5345 PAD.n5204 2.24164
R40893 PAD.n5279 PAD.n5197 2.24164
R40894 PAD.n5337 PAD.n5204 2.24164
R40895 PAD.n5335 PAD.n5197 2.24164
R40896 PAD.n5333 PAD.n5204 2.24164
R40897 PAD.n5283 PAD.n5197 2.24164
R40898 PAD.n5325 PAD.n5204 2.24164
R40899 PAD.n5323 PAD.n5197 2.24164
R40900 PAD.n5321 PAD.n5204 2.24164
R40901 PAD.n5287 PAD.n5197 2.24164
R40902 PAD.n5313 PAD.n5204 2.24164
R40903 PAD.n5311 PAD.n5197 2.24164
R40904 PAD.n5309 PAD.n5204 2.24164
R40905 PAD.n5291 PAD.n5197 2.24164
R40906 PAD.n5301 PAD.n5204 2.24164
R40907 PAD.n5299 PAD.n5197 2.24164
R40908 PAD.n5297 PAD.n5204 2.24164
R40909 PAD.n7520 PAD.n7519 2.24164
R40910 PAD.n7511 PAD.n7207 2.24164
R40911 PAD.n7520 PAD.n7199 2.24164
R40912 PAD.n7508 PAD.n7207 2.24164
R40913 PAD.n7520 PAD.n7198 2.24164
R40914 PAD.n7500 PAD.n7207 2.24164
R40915 PAD.n7520 PAD.n7197 2.24164
R40916 PAD.n7496 PAD.n7207 2.24164
R40917 PAD.n7520 PAD.n7196 2.24164
R40918 PAD.n7488 PAD.n7207 2.24164
R40919 PAD.n7520 PAD.n7195 2.24164
R40920 PAD.n7484 PAD.n7207 2.24164
R40921 PAD.n7520 PAD.n7194 2.24164
R40922 PAD.n7476 PAD.n7207 2.24164
R40923 PAD.n7520 PAD.n7193 2.24164
R40924 PAD.n7472 PAD.n7207 2.24164
R40925 PAD.n7520 PAD.n7192 2.24164
R40926 PAD.n7464 PAD.n7207 2.24164
R40927 PAD.n7520 PAD.n7191 2.24164
R40928 PAD.n7460 PAD.n7207 2.24164
R40929 PAD.n7520 PAD.n7190 2.24164
R40930 PAD.n7452 PAD.n7207 2.24164
R40931 PAD.n7520 PAD.n7189 2.24164
R40932 PAD.n7448 PAD.n7207 2.24164
R40933 PAD.n7520 PAD.n7188 2.24164
R40934 PAD.n7440 PAD.n7207 2.24164
R40935 PAD.n7520 PAD.n7187 2.24164
R40936 PAD.n7436 PAD.n7207 2.24164
R40937 PAD.n7520 PAD.n7186 2.24164
R40938 PAD.n7428 PAD.n7207 2.24164
R40939 PAD.n7520 PAD.n7185 2.24164
R40940 PAD.n7424 PAD.n7207 2.24164
R40941 PAD.n7520 PAD.n7184 2.24164
R40942 PAD.n7416 PAD.n7207 2.24164
R40943 PAD.n7520 PAD.n7183 2.24164
R40944 PAD.n7412 PAD.n7207 2.24164
R40945 PAD.n7520 PAD.n7182 2.24164
R40946 PAD.n7404 PAD.n7207 2.24164
R40947 PAD.n7520 PAD.n7181 2.24164
R40948 PAD.n7400 PAD.n7207 2.24164
R40949 PAD.n7520 PAD.n7180 2.24164
R40950 PAD.n7392 PAD.n7207 2.24164
R40951 PAD.n7520 PAD.n7179 2.24164
R40952 PAD.n7388 PAD.n7207 2.24164
R40953 PAD.n7520 PAD.n7178 2.24164
R40954 PAD.n7380 PAD.n7207 2.24164
R40955 PAD.n7520 PAD.n7177 2.24164
R40956 PAD.n7376 PAD.n7207 2.24164
R40957 PAD.n7520 PAD.n7176 2.24164
R40958 PAD.n7368 PAD.n7207 2.24164
R40959 PAD.n7520 PAD.n7175 2.24164
R40960 PAD.n7364 PAD.n7207 2.24164
R40961 PAD.n7520 PAD.n7174 2.24164
R40962 PAD.n7356 PAD.n7207 2.24164
R40963 PAD.n7520 PAD.n7173 2.24164
R40964 PAD.n7352 PAD.n7207 2.24164
R40965 PAD.n7520 PAD.n7172 2.24164
R40966 PAD.n7344 PAD.n7207 2.24164
R40967 PAD.n7520 PAD.n7171 2.24164
R40968 PAD.n7340 PAD.n7207 2.24164
R40969 PAD.n7520 PAD.n7170 2.24164
R40970 PAD.n7332 PAD.n7207 2.24164
R40971 PAD.n7520 PAD.n7169 2.24164
R40972 PAD.n7328 PAD.n7207 2.24164
R40973 PAD.n7520 PAD.n7168 2.24164
R40974 PAD.n7320 PAD.n7207 2.24164
R40975 PAD.n7520 PAD.n7167 2.24164
R40976 PAD.n7316 PAD.n7207 2.24164
R40977 PAD.n7520 PAD.n7166 2.24164
R40978 PAD.n7308 PAD.n7207 2.24164
R40979 PAD.n7520 PAD.n7165 2.24164
R40980 PAD.n7304 PAD.n7207 2.24164
R40981 PAD.n7520 PAD.n7164 2.24164
R40982 PAD.n7296 PAD.n7207 2.24164
R40983 PAD.n7520 PAD.n7163 2.24164
R40984 PAD.n7292 PAD.n7207 2.24164
R40985 PAD.n7520 PAD.n7162 2.24164
R40986 PAD.n7284 PAD.n7207 2.24164
R40987 PAD.n7520 PAD.n7161 2.24164
R40988 PAD.n7280 PAD.n7207 2.24164
R40989 PAD.n7520 PAD.n7160 2.24164
R40990 PAD.n7272 PAD.n7207 2.24164
R40991 PAD.n7520 PAD.n7159 2.24164
R40992 PAD.n7782 PAD.n7781 2.24164
R40993 PAD.n7773 PAD.n7105 2.24164
R40994 PAD.n7782 PAD.n7102 2.24164
R40995 PAD.n7770 PAD.n7105 2.24164
R40996 PAD.n7782 PAD.n7101 2.24164
R40997 PAD.n7762 PAD.n7105 2.24164
R40998 PAD.n7782 PAD.n7100 2.24164
R40999 PAD.n7758 PAD.n7105 2.24164
R41000 PAD.n7782 PAD.n7099 2.24164
R41001 PAD.n7750 PAD.n7105 2.24164
R41002 PAD.n7782 PAD.n7098 2.24164
R41003 PAD.n7746 PAD.n7105 2.24164
R41004 PAD.n7782 PAD.n7097 2.24164
R41005 PAD.n7738 PAD.n7105 2.24164
R41006 PAD.n7782 PAD.n7096 2.24164
R41007 PAD.n7734 PAD.n7105 2.24164
R41008 PAD.n7782 PAD.n7095 2.24164
R41009 PAD.n7726 PAD.n7105 2.24164
R41010 PAD.n7782 PAD.n7094 2.24164
R41011 PAD.n7722 PAD.n7105 2.24164
R41012 PAD.n7782 PAD.n7093 2.24164
R41013 PAD.n7714 PAD.n7105 2.24164
R41014 PAD.n7782 PAD.n7092 2.24164
R41015 PAD.n7710 PAD.n7105 2.24164
R41016 PAD.n7782 PAD.n7091 2.24164
R41017 PAD.n7702 PAD.n7105 2.24164
R41018 PAD.n7782 PAD.n7090 2.24164
R41019 PAD.n7698 PAD.n7105 2.24164
R41020 PAD.n7782 PAD.n7089 2.24164
R41021 PAD.n7690 PAD.n7105 2.24164
R41022 PAD.n7782 PAD.n7088 2.24164
R41023 PAD.n7686 PAD.n7105 2.24164
R41024 PAD.n7782 PAD.n7087 2.24164
R41025 PAD.n7678 PAD.n7105 2.24164
R41026 PAD.n7782 PAD.n7086 2.24164
R41027 PAD.n7674 PAD.n7105 2.24164
R41028 PAD.n7782 PAD.n7085 2.24164
R41029 PAD.n7666 PAD.n7105 2.24164
R41030 PAD.n7782 PAD.n7084 2.24164
R41031 PAD.n7662 PAD.n7105 2.24164
R41032 PAD.n7782 PAD.n7083 2.24164
R41033 PAD.n7654 PAD.n7105 2.24164
R41034 PAD.n7782 PAD.n7082 2.24164
R41035 PAD.n7650 PAD.n7105 2.24164
R41036 PAD.n7782 PAD.n7081 2.24164
R41037 PAD.n7642 PAD.n7105 2.24164
R41038 PAD.n7782 PAD.n7080 2.24164
R41039 PAD.n7638 PAD.n7105 2.24164
R41040 PAD.n7782 PAD.n7079 2.24164
R41041 PAD.n7630 PAD.n7105 2.24164
R41042 PAD.n7782 PAD.n7078 2.24164
R41043 PAD.n7626 PAD.n7105 2.24164
R41044 PAD.n7782 PAD.n7077 2.24164
R41045 PAD.n7618 PAD.n7105 2.24164
R41046 PAD.n7782 PAD.n7076 2.24164
R41047 PAD.n7614 PAD.n7105 2.24164
R41048 PAD.n7782 PAD.n7075 2.24164
R41049 PAD.n7606 PAD.n7105 2.24164
R41050 PAD.n7782 PAD.n7074 2.24164
R41051 PAD.n7602 PAD.n7105 2.24164
R41052 PAD.n7782 PAD.n7073 2.24164
R41053 PAD.n7594 PAD.n7105 2.24164
R41054 PAD.n7782 PAD.n7072 2.24164
R41055 PAD.n7590 PAD.n7105 2.24164
R41056 PAD.n7782 PAD.n7071 2.24164
R41057 PAD.n7582 PAD.n7105 2.24164
R41058 PAD.n7782 PAD.n7070 2.24164
R41059 PAD.n7578 PAD.n7105 2.24164
R41060 PAD.n7782 PAD.n7069 2.24164
R41061 PAD.n7570 PAD.n7105 2.24164
R41062 PAD.n7782 PAD.n7068 2.24164
R41063 PAD.n7566 PAD.n7105 2.24164
R41064 PAD.n7782 PAD.n7067 2.24164
R41065 PAD.n7558 PAD.n7105 2.24164
R41066 PAD.n7782 PAD.n7066 2.24164
R41067 PAD.n7554 PAD.n7105 2.24164
R41068 PAD.n7782 PAD.n7065 2.24164
R41069 PAD.n7546 PAD.n7105 2.24164
R41070 PAD.n7782 PAD.n7064 2.24164
R41071 PAD.n7542 PAD.n7105 2.24164
R41072 PAD.n7782 PAD.n7063 2.24164
R41073 PAD.n7534 PAD.n7105 2.24164
R41074 PAD.n7782 PAD.n7062 2.24164
R41075 PAD.n6721 PAD.n6712 2.24164
R41076 PAD.n7047 PAD.n6713 2.24164
R41077 PAD.n7045 PAD.n6712 2.24164
R41078 PAD.n6722 PAD.n6713 2.24164
R41079 PAD.n7037 PAD.n6712 2.24164
R41080 PAD.n7035 PAD.n6713 2.24164
R41081 PAD.n7033 PAD.n6712 2.24164
R41082 PAD.n6727 PAD.n6713 2.24164
R41083 PAD.n7025 PAD.n6712 2.24164
R41084 PAD.n7023 PAD.n6713 2.24164
R41085 PAD.n7021 PAD.n6712 2.24164
R41086 PAD.n6731 PAD.n6713 2.24164
R41087 PAD.n7013 PAD.n6712 2.24164
R41088 PAD.n7011 PAD.n6713 2.24164
R41089 PAD.n7009 PAD.n6712 2.24164
R41090 PAD.n6735 PAD.n6713 2.24164
R41091 PAD.n7001 PAD.n6712 2.24164
R41092 PAD.n6999 PAD.n6713 2.24164
R41093 PAD.n6997 PAD.n6712 2.24164
R41094 PAD.n6739 PAD.n6713 2.24164
R41095 PAD.n6989 PAD.n6712 2.24164
R41096 PAD.n6987 PAD.n6713 2.24164
R41097 PAD.n6985 PAD.n6712 2.24164
R41098 PAD.n6743 PAD.n6713 2.24164
R41099 PAD.n6977 PAD.n6712 2.24164
R41100 PAD.n6975 PAD.n6713 2.24164
R41101 PAD.n6973 PAD.n6712 2.24164
R41102 PAD.n6747 PAD.n6713 2.24164
R41103 PAD.n6965 PAD.n6712 2.24164
R41104 PAD.n6963 PAD.n6713 2.24164
R41105 PAD.n6961 PAD.n6712 2.24164
R41106 PAD.n6751 PAD.n6713 2.24164
R41107 PAD.n6953 PAD.n6712 2.24164
R41108 PAD.n6951 PAD.n6713 2.24164
R41109 PAD.n6949 PAD.n6712 2.24164
R41110 PAD.n6755 PAD.n6713 2.24164
R41111 PAD.n6941 PAD.n6712 2.24164
R41112 PAD.n6939 PAD.n6713 2.24164
R41113 PAD.n6937 PAD.n6712 2.24164
R41114 PAD.n6759 PAD.n6713 2.24164
R41115 PAD.n6929 PAD.n6712 2.24164
R41116 PAD.n6927 PAD.n6713 2.24164
R41117 PAD.n6925 PAD.n6712 2.24164
R41118 PAD.n6763 PAD.n6713 2.24164
R41119 PAD.n6917 PAD.n6712 2.24164
R41120 PAD.n6915 PAD.n6713 2.24164
R41121 PAD.n6913 PAD.n6712 2.24164
R41122 PAD.n6767 PAD.n6713 2.24164
R41123 PAD.n6905 PAD.n6712 2.24164
R41124 PAD.n6903 PAD.n6713 2.24164
R41125 PAD.n6901 PAD.n6712 2.24164
R41126 PAD.n6771 PAD.n6713 2.24164
R41127 PAD.n6893 PAD.n6712 2.24164
R41128 PAD.n6891 PAD.n6713 2.24164
R41129 PAD.n6889 PAD.n6712 2.24164
R41130 PAD.n6775 PAD.n6713 2.24164
R41131 PAD.n6881 PAD.n6712 2.24164
R41132 PAD.n6879 PAD.n6713 2.24164
R41133 PAD.n6877 PAD.n6712 2.24164
R41134 PAD.n6779 PAD.n6713 2.24164
R41135 PAD.n6869 PAD.n6712 2.24164
R41136 PAD.n6867 PAD.n6713 2.24164
R41137 PAD.n6865 PAD.n6712 2.24164
R41138 PAD.n6783 PAD.n6713 2.24164
R41139 PAD.n6857 PAD.n6712 2.24164
R41140 PAD.n6855 PAD.n6713 2.24164
R41141 PAD.n6853 PAD.n6712 2.24164
R41142 PAD.n6787 PAD.n6713 2.24164
R41143 PAD.n6845 PAD.n6712 2.24164
R41144 PAD.n6843 PAD.n6713 2.24164
R41145 PAD.n6841 PAD.n6712 2.24164
R41146 PAD.n6791 PAD.n6713 2.24164
R41147 PAD.n6833 PAD.n6712 2.24164
R41148 PAD.n6831 PAD.n6713 2.24164
R41149 PAD.n6829 PAD.n6712 2.24164
R41150 PAD.n6795 PAD.n6713 2.24164
R41151 PAD.n6821 PAD.n6712 2.24164
R41152 PAD.n6819 PAD.n6713 2.24164
R41153 PAD.n6817 PAD.n6712 2.24164
R41154 PAD.n6799 PAD.n6713 2.24164
R41155 PAD.n6809 PAD.n6712 2.24164
R41156 PAD.n6807 PAD.n6713 2.24164
R41157 PAD.n6805 PAD.n6712 2.24164
R41158 PAD.n5894 PAD.n5893 2.24164
R41159 PAD.n5603 PAD.n5551 2.24164
R41160 PAD.n5894 PAD.n5601 2.24164
R41161 PAD.n5884 PAD.n5551 2.24164
R41162 PAD.n5894 PAD.n5600 2.24164
R41163 PAD.n5609 PAD.n5551 2.24164
R41164 PAD.n5894 PAD.n5599 2.24164
R41165 PAD.n5875 PAD.n5551 2.24164
R41166 PAD.n5894 PAD.n5598 2.24164
R41167 PAD.n5614 PAD.n5551 2.24164
R41168 PAD.n5894 PAD.n5597 2.24164
R41169 PAD.n5866 PAD.n5551 2.24164
R41170 PAD.n5894 PAD.n5596 2.24164
R41171 PAD.n5619 PAD.n5551 2.24164
R41172 PAD.n5894 PAD.n5595 2.24164
R41173 PAD.n5857 PAD.n5551 2.24164
R41174 PAD.n5894 PAD.n5594 2.24164
R41175 PAD.n5624 PAD.n5551 2.24164
R41176 PAD.n5894 PAD.n5593 2.24164
R41177 PAD.n5848 PAD.n5551 2.24164
R41178 PAD.n5894 PAD.n5592 2.24164
R41179 PAD.n5629 PAD.n5551 2.24164
R41180 PAD.n5894 PAD.n5591 2.24164
R41181 PAD.n5839 PAD.n5551 2.24164
R41182 PAD.n5894 PAD.n5590 2.24164
R41183 PAD.n5634 PAD.n5551 2.24164
R41184 PAD.n5894 PAD.n5589 2.24164
R41185 PAD.n5830 PAD.n5551 2.24164
R41186 PAD.n5894 PAD.n5588 2.24164
R41187 PAD.n5639 PAD.n5551 2.24164
R41188 PAD.n5894 PAD.n5587 2.24164
R41189 PAD.n5821 PAD.n5551 2.24164
R41190 PAD.n5894 PAD.n5586 2.24164
R41191 PAD.n5644 PAD.n5551 2.24164
R41192 PAD.n5894 PAD.n5585 2.24164
R41193 PAD.n5812 PAD.n5551 2.24164
R41194 PAD.n5894 PAD.n5584 2.24164
R41195 PAD.n5649 PAD.n5551 2.24164
R41196 PAD.n5894 PAD.n5583 2.24164
R41197 PAD.n5803 PAD.n5551 2.24164
R41198 PAD.n5894 PAD.n5582 2.24164
R41199 PAD.n5654 PAD.n5551 2.24164
R41200 PAD.n5894 PAD.n5581 2.24164
R41201 PAD.n5794 PAD.n5551 2.24164
R41202 PAD.n5894 PAD.n5580 2.24164
R41203 PAD.n5659 PAD.n5551 2.24164
R41204 PAD.n5894 PAD.n5579 2.24164
R41205 PAD.n5785 PAD.n5551 2.24164
R41206 PAD.n5894 PAD.n5578 2.24164
R41207 PAD.n5664 PAD.n5551 2.24164
R41208 PAD.n5894 PAD.n5577 2.24164
R41209 PAD.n5776 PAD.n5551 2.24164
R41210 PAD.n5894 PAD.n5576 2.24164
R41211 PAD.n5669 PAD.n5551 2.24164
R41212 PAD.n5894 PAD.n5575 2.24164
R41213 PAD.n5767 PAD.n5551 2.24164
R41214 PAD.n5894 PAD.n5574 2.24164
R41215 PAD.n5674 PAD.n5551 2.24164
R41216 PAD.n5894 PAD.n5573 2.24164
R41217 PAD.n5758 PAD.n5551 2.24164
R41218 PAD.n5894 PAD.n5572 2.24164
R41219 PAD.n5679 PAD.n5551 2.24164
R41220 PAD.n5894 PAD.n5571 2.24164
R41221 PAD.n5749 PAD.n5551 2.24164
R41222 PAD.n5894 PAD.n5570 2.24164
R41223 PAD.n5684 PAD.n5551 2.24164
R41224 PAD.n5894 PAD.n5569 2.24164
R41225 PAD.n5740 PAD.n5551 2.24164
R41226 PAD.n5894 PAD.n5568 2.24164
R41227 PAD.n5689 PAD.n5551 2.24164
R41228 PAD.n5894 PAD.n5567 2.24164
R41229 PAD.n5731 PAD.n5551 2.24164
R41230 PAD.n5894 PAD.n5566 2.24164
R41231 PAD.n5694 PAD.n5551 2.24164
R41232 PAD.n5894 PAD.n5565 2.24164
R41233 PAD.n5722 PAD.n5551 2.24164
R41234 PAD.n5894 PAD.n5564 2.24164
R41235 PAD.n5699 PAD.n5551 2.24164
R41236 PAD.n5894 PAD.n5563 2.24164
R41237 PAD.n5713 PAD.n5551 2.24164
R41238 PAD.n5894 PAD.n5562 2.24164
R41239 PAD.n5706 PAD.n5551 2.24164
R41240 PAD.n5894 PAD.n5561 2.24164
R41241 PAD.n6678 PAD.n5902 2.24164
R41242 PAD.n6689 PAD.n5906 2.24164
R41243 PAD.n6678 PAD.n6397 2.24164
R41244 PAD.n6689 PAD.n5907 2.24164
R41245 PAD.n6678 PAD.n6398 2.24164
R41246 PAD.n6689 PAD.n5908 2.24164
R41247 PAD.n6678 PAD.n6399 2.24164
R41248 PAD.n6689 PAD.n5909 2.24164
R41249 PAD.n6678 PAD.n6400 2.24164
R41250 PAD.n6689 PAD.n5910 2.24164
R41251 PAD.n6678 PAD.n6401 2.24164
R41252 PAD.n6689 PAD.n5911 2.24164
R41253 PAD.n6678 PAD.n6402 2.24164
R41254 PAD.n6689 PAD.n5912 2.24164
R41255 PAD.n6678 PAD.n6403 2.24164
R41256 PAD.n6689 PAD.n5913 2.24164
R41257 PAD.n6678 PAD.n6404 2.24164
R41258 PAD.n6689 PAD.n5914 2.24164
R41259 PAD.n6678 PAD.n6405 2.24164
R41260 PAD.n6689 PAD.n5915 2.24164
R41261 PAD.n6678 PAD.n6406 2.24164
R41262 PAD.n6689 PAD.n5916 2.24164
R41263 PAD.n6678 PAD.n6407 2.24164
R41264 PAD.n6689 PAD.n5917 2.24164
R41265 PAD.n6678 PAD.n6408 2.24164
R41266 PAD.n6689 PAD.n5918 2.24164
R41267 PAD.n6678 PAD.n6409 2.24164
R41268 PAD.n6689 PAD.n5919 2.24164
R41269 PAD.n6678 PAD.n6410 2.24164
R41270 PAD.n6689 PAD.n5920 2.24164
R41271 PAD.n6678 PAD.n6411 2.24164
R41272 PAD.n6689 PAD.n5921 2.24164
R41273 PAD.n6678 PAD.n6412 2.24164
R41274 PAD.n6689 PAD.n5922 2.24164
R41275 PAD.n6678 PAD.n6413 2.24164
R41276 PAD.n6689 PAD.n5923 2.24164
R41277 PAD.n6678 PAD.n6414 2.24164
R41278 PAD.n6689 PAD.n5924 2.24164
R41279 PAD.n6678 PAD.n6415 2.24164
R41280 PAD.n6689 PAD.n5925 2.24164
R41281 PAD.n6678 PAD.n6416 2.24164
R41282 PAD.n6689 PAD.n5926 2.24164
R41283 PAD.n6678 PAD.n6417 2.24164
R41284 PAD.n6689 PAD.n5927 2.24164
R41285 PAD.n6678 PAD.n6418 2.24164
R41286 PAD.n6689 PAD.n5928 2.24164
R41287 PAD.n6678 PAD.n6419 2.24164
R41288 PAD.n6689 PAD.n5929 2.24164
R41289 PAD.n6678 PAD.n6420 2.24164
R41290 PAD.n6689 PAD.n5930 2.24164
R41291 PAD.n6678 PAD.n6421 2.24164
R41292 PAD.n6689 PAD.n5931 2.24164
R41293 PAD.n6678 PAD.n6422 2.24164
R41294 PAD.n6689 PAD.n5932 2.24164
R41295 PAD.n6678 PAD.n6423 2.24164
R41296 PAD.n6689 PAD.n5933 2.24164
R41297 PAD.n6678 PAD.n6424 2.24164
R41298 PAD.n6689 PAD.n5934 2.24164
R41299 PAD.n6678 PAD.n6425 2.24164
R41300 PAD.n6689 PAD.n5935 2.24164
R41301 PAD.n6678 PAD.n6426 2.24164
R41302 PAD.n6689 PAD.n5936 2.24164
R41303 PAD.n6678 PAD.n6427 2.24164
R41304 PAD.n6689 PAD.n5937 2.24164
R41305 PAD.n6678 PAD.n6428 2.24164
R41306 PAD.n6689 PAD.n5938 2.24164
R41307 PAD.n6678 PAD.n6429 2.24164
R41308 PAD.n6689 PAD.n5939 2.24164
R41309 PAD.n6678 PAD.n6430 2.24164
R41310 PAD.n6689 PAD.n5940 2.24164
R41311 PAD.n6678 PAD.n6431 2.24164
R41312 PAD.n6689 PAD.n5941 2.24164
R41313 PAD.n6678 PAD.n6432 2.24164
R41314 PAD.n6689 PAD.n5942 2.24164
R41315 PAD.n6678 PAD.n6433 2.24164
R41316 PAD.n6689 PAD.n5943 2.24164
R41317 PAD.n6678 PAD.n6434 2.24164
R41318 PAD.n6689 PAD.n5944 2.24164
R41319 PAD.n6678 PAD.n6435 2.24164
R41320 PAD.n6689 PAD.n5945 2.24164
R41321 PAD.n6678 PAD.n6677 2.24164
R41322 PAD.n6689 PAD.n5946 2.24164
R41323 PAD.n6678 PAD.n5947 2.24164
R41324 PAD.n11518 PAD.n10745 1.1255
R41325 PAD.n11520 PAD.n11519 1.1255
R41326 PAD.n11089 PAD.n10744 1.1255
R41327 PAD.n10751 PAD.n10746 1.1255
R41328 PAD.n17 PAD.n15 1.1255
R41329 PAD.n11537 PAD.n11536 1.1255
R41330 PAD.n10725 PAD.n10724 1.1255
R41331 PAD.n10723 PAD.n369 1.1255
R41332 PAD.n10722 PAD.n10721 1.1255
R41333 PAD.n371 PAD.n370 1.1255
R41334 PAD.n10699 PAD.n10698 1.1255
R41335 PAD.n10412 PAD.n428 1.1255
R41336 PAD.n10411 PAD.n10410 1.1255
R41337 PAD.n10395 PAD.n10394 1.1255
R41338 PAD.n10393 PAD.n778 1.1255
R41339 PAD.n10392 PAD.n10391 1.1255
R41340 PAD.n10369 PAD.n1123 1.1255
R41341 PAD.n10371 PAD.n10370 1.1255
R41342 PAD.n10368 PAD.n1122 1.1255
R41343 PAD.n10365 PAD.n10364 1.1255
R41344 PAD.n1126 PAD.n1125 1.1255
R41345 PAD.n10014 PAD.n10013 1.1255
R41346 PAD.n10011 PAD.n10010 1.1255
R41347 PAD.n1147 PAD.n1146 1.1255
R41348 PAD.n1583 PAD.n1582 1.1255
R41349 PAD.n9747 PAD.n1584 1.1255
R41350 PAD.n9727 PAD.n1581 1.1255
R41351 PAD.n9728 PAD.n1597 1.1255
R41352 PAD.n9730 PAD.n9729 1.1255
R41353 PAD.n9725 PAD.n9724 1.1255
R41354 PAD.n1934 PAD.n1933 1.1255
R41355 PAD.n9461 PAD.n2034 1.1255
R41356 PAD.n9192 PAD.n2033 1.1255
R41357 PAD.n9193 PAD.n2036 1.1255
R41358 PAD.n9195 PAD.n9194 1.1255
R41359 PAD.n9191 PAD.n2137 1.1255
R41360 PAD.n9169 PAD.n2136 1.1255
R41361 PAD.n9170 PAD.n2149 1.1255
R41362 PAD.n9173 PAD.n9172 1.1255
R41363 PAD.n9166 PAD.n9165 1.1255
R41364 PAD.n2485 PAD.n2484 1.1255
R41365 PAD.n9149 PAD.n9148 1.1255
R41366 PAD.n9146 PAD.n9145 1.1255
R41367 PAD.n2832 PAD.n2831 1.1255
R41368 PAD.n9123 PAD.n9122 1.1255
R41369 PAD.n9126 PAD.n9125 1.1255
R41370 PAD.n8836 PAD.n2886 1.1255
R41371 PAD.n8835 PAD.n8834 1.1255
R41372 PAD.n8525 PAD.n8524 1.1255
R41373 PAD.n8523 PAD.n2948 1.1255
R41374 PAD.n8522 PAD.n8521 1.1255
R41375 PAD.n8498 PAD.n3292 1.1255
R41376 PAD.n8500 PAD.n8499 1.1255
R41377 PAD.n8497 PAD.n3291 1.1255
R41378 PAD.n8496 PAD.n8495 1.1255
R41379 PAD.n8476 PAD.n8475 1.1255
R41380 PAD.n8474 PAD.n3635 1.1255
R41381 PAD.n8472 PAD.n8471 1.1255
R41382 PAD.n8451 PAD.n8450 1.1255
R41383 PAD.n8449 PAD.n3979 1.1255
R41384 PAD.n8448 PAD.n8447 1.1255
R41385 PAD.n8426 PAD.n4324 1.1255
R41386 PAD.n8428 PAD.n8427 1.1255
R41387 PAD.n8425 PAD.n4323 1.1255
R41388 PAD.n8423 PAD.n8422 1.1255
R41389 PAD.n4327 PAD.n4326 1.1255
R41390 PAD.n8405 PAD.n8404 1.1255
R41391 PAD.n8403 PAD.n4675 1.1255
R41392 PAD.n8401 PAD.n8400 1.1255
R41393 PAD.n4678 PAD.n4677 1.1255
R41394 PAD.n8192 PAD.n8191 1.1255
R41395 PAD.n8189 PAD.n8188 1.1255
R41396 PAD.n5181 PAD.n5180 1.1255
R41397 PAD.n8172 PAD.n8171 1.1255
R41398 PAD.n8169 PAD.n8168 1.1255
R41399 PAD.n5195 PAD.n5194 1.1255
R41400 PAD.n7814 PAD.n7813 1.1255
R41401 PAD.n7817 PAD.n7816 1.1255
R41402 PAD.n5209 PAD.n5207 1.1255
R41403 PAD.n7226 PAD.n7225 1.1255
R41404 PAD.n7227 PAD.n7208 1.1255
R41405 PAD.n7220 PAD.n7219 1.1255
R41406 PAD.n7211 PAD.n7210 1.1255
R41407 PAD.n7213 PAD.n7212 1.1255
R41408 PAD.n7786 PAD.n7785 1.1255
R41409 PAD.n7787 PAD.n6717 1.1255
R41410 PAD.n7789 PAD.n7788 1.1255
R41411 PAD.n7054 PAD.n7053 1.1255
R41412 PAD.n5548 PAD.n5546 1.1255
R41413 PAD.n7805 PAD.n7804 1.1255
R41414 PAD.n6697 PAD.n5544 1.1255
R41415 PAD.n6696 PAD.n6695 1.1255
R41416 PAD.n6694 PAD.n5896 1.1255
R41417 PAD.n6394 PAD.n5897 1.1255
R41418 PAD.n6393 PAD.n6392 1.1255
R41419 PAD.n6391 PAD.n5955 1.1255
R41420 PAD.n5970 PAD.n5955 1.1255
R41421 PAD.n6393 PAD.n5954 1.1255
R41422 PAD.n6395 PAD.n6394 1.1255
R41423 PAD.n6681 PAD.n5896 1.1255
R41424 PAD.n6696 PAD.n5895 1.1255
R41425 PAD.n6698 PAD.n6697 1.1255
R41426 PAD.n7804 PAD.n7803 1.1255
R41427 PAD.n5550 PAD.n5548 1.1255
R41428 PAD.n7053 PAD.n7052 1.1255
R41429 PAD.n7790 PAD.n7789 1.1255
R41430 PAD.n6717 PAD.n6715 1.1255
R41431 PAD.n7785 PAD.n7784 1.1255
R41432 PAD.n7214 PAD.n7213 1.1255
R41433 PAD.n7217 PAD.n7211 1.1255
R41434 PAD.n7219 PAD.n7218 1.1255
R41435 PAD.n7208 PAD.n7202 1.1255
R41436 PAD.n7225 PAD.n7224 1.1255
R41437 PAD.n5207 PAD.n5205 1.1255
R41438 PAD.n7818 PAD.n7817 1.1255
R41439 PAD.n7813 PAD.n5196 1.1255
R41440 PAD.n8166 PAD.n5195 1.1255
R41441 PAD.n8168 PAD.n8167 1.1255
R41442 PAD.n8173 PAD.n8172 1.1255
R41443 PAD.n5182 PAD.n5181 1.1255
R41444 PAD.n8188 PAD.n8187 1.1255
R41445 PAD.n8193 PAD.n8192 1.1255
R41446 PAD.n4680 PAD.n4678 1.1255
R41447 PAD.n8400 PAD.n8399 1.1255
R41448 PAD.n4675 PAD.n4674 1.1255
R41449 PAD.n8406 PAD.n8405 1.1255
R41450 PAD.n4329 PAD.n4327 1.1255
R41451 PAD.n8422 PAD.n8421 1.1255
R41452 PAD.n4323 PAD.n4320 1.1255
R41453 PAD.n8429 PAD.n8428 1.1255
R41454 PAD.n4324 PAD.n4322 1.1255
R41455 PAD.n8447 PAD.n8446 1.1255
R41456 PAD.n3979 PAD.n3978 1.1255
R41457 PAD.n8452 PAD.n8451 1.1255
R41458 PAD.n8471 PAD.n8470 1.1255
R41459 PAD.n3635 PAD.n3634 1.1255
R41460 PAD.n8477 PAD.n8476 1.1255
R41461 PAD.n8495 PAD.n8494 1.1255
R41462 PAD.n3291 PAD.n3288 1.1255
R41463 PAD.n8501 PAD.n8500 1.1255
R41464 PAD.n3292 PAD.n3290 1.1255
R41465 PAD.n8521 PAD.n8520 1.1255
R41466 PAD.n2948 PAD.n2947 1.1255
R41467 PAD.n8526 PAD.n8525 1.1255
R41468 PAD.n8834 PAD.n8833 1.1255
R41469 PAD.n2886 PAD.n2884 1.1255
R41470 PAD.n9127 PAD.n9126 1.1255
R41471 PAD.n9122 PAD.n9121 1.1255
R41472 PAD.n2833 PAD.n2832 1.1255
R41473 PAD.n9145 PAD.n9144 1.1255
R41474 PAD.n9150 PAD.n9149 1.1255
R41475 PAD.n2486 PAD.n2485 1.1255
R41476 PAD.n9165 PAD.n9164 1.1255
R41477 PAD.n9174 PAD.n9173 1.1255
R41478 PAD.n2149 PAD.n2138 1.1255
R41479 PAD.n9188 PAD.n2136 1.1255
R41480 PAD.n9191 PAD.n9190 1.1255
R41481 PAD.n9195 PAD.n2035 1.1255
R41482 PAD.n9457 PAD.n2036 1.1255
R41483 PAD.n9458 PAD.n2033 1.1255
R41484 PAD.n9461 PAD.n9460 1.1255
R41485 PAD.n1935 PAD.n1934 1.1255
R41486 PAD.n9724 PAD.n9723 1.1255
R41487 PAD.n9731 PAD.n9730 1.1255
R41488 PAD.n1597 PAD.n1585 1.1255
R41489 PAD.n9743 PAD.n1581 1.1255
R41490 PAD.n9747 PAD.n9746 1.1255
R41491 PAD.n9745 PAD.n1582 1.1255
R41492 PAD.n1148 PAD.n1147 1.1255
R41493 PAD.n10010 PAD.n10009 1.1255
R41494 PAD.n10015 PAD.n10014 1.1255
R41495 PAD.n1128 PAD.n1126 1.1255
R41496 PAD.n10364 PAD.n10363 1.1255
R41497 PAD.n1122 PAD.n1119 1.1255
R41498 PAD.n10372 PAD.n10371 1.1255
R41499 PAD.n1123 PAD.n1121 1.1255
R41500 PAD.n10391 PAD.n10390 1.1255
R41501 PAD.n778 PAD.n777 1.1255
R41502 PAD.n10396 PAD.n10395 1.1255
R41503 PAD.n10410 PAD.n10409 1.1255
R41504 PAD.n428 PAD.n426 1.1255
R41505 PAD.n10700 PAD.n10699 1.1255
R41506 PAD.n372 PAD.n371 1.1255
R41507 PAD.n10721 PAD.n10720 1.1255
R41508 PAD.n369 PAD.n368 1.1255
R41509 PAD.n10726 PAD.n10725 1.1255
R41510 PAD.n11536 PAD.n11535 1.1255
R41511 PAD.n19 PAD.n17 1.1255
R41512 PAD.n10752 PAD.n10751 1.1255
R41513 PAD.n10744 PAD.n10742 1.1255
R41514 PAD.n11521 PAD.n11520 1.1255
R41515 PAD.n10745 PAD.n10743 1.1255
R41516 PAD.n5971 PAD.n5970 1.1255
R41517 PAD.n5954 PAD.n5903 1.1255
R41518 PAD.n6396 PAD.n6395 1.1255
R41519 PAD.n6682 PAD.n6681 1.1255
R41520 PAD.n6679 PAD.n5895 1.1255
R41521 PAD.n6699 PAD.n6698 1.1255
R41522 PAD.n7803 PAD.n7802 1.1255
R41523 PAD.n5552 PAD.n5550 1.1255
R41524 PAD.n7052 PAD.n6712 1.1255
R41525 PAD.n7791 PAD.n7790 1.1255
R41526 PAD.n7060 PAD.n6715 1.1255
R41527 PAD.n7784 PAD.n7783 1.1255
R41528 PAD.n7214 PAD.n7103 1.1255
R41529 PAD.n7217 PAD.n7216 1.1255
R41530 PAD.n7218 PAD.n7158 1.1255
R41531 PAD.n7202 PAD.n7200 1.1255
R41532 PAD.n7224 PAD.n7223 1.1255
R41533 PAD.n7221 PAD.n5205 1.1255
R41534 PAD.n7819 PAD.n7818 1.1255
R41535 PAD.n7829 PAD.n5196 1.1255
R41536 PAD.n8166 PAD.n8165 1.1255
R41537 PAD.n8167 PAD.n5190 1.1255
R41538 PAD.n8174 PAD.n8173 1.1255
R41539 PAD.n8184 PAD.n5182 1.1255
R41540 PAD.n8187 PAD.n8186 1.1255
R41541 PAD.n8194 PAD.n8193 1.1255
R41542 PAD.n4841 PAD.n4680 1.1255
R41543 PAD.n8399 PAD.n8398 1.1255
R41544 PAD.n4724 PAD.n4674 1.1255
R41545 PAD.n8407 PAD.n8406 1.1255
R41546 PAD.n8409 PAD.n4329 1.1255
R41547 PAD.n8421 PAD.n8420 1.1255
R41548 PAD.n4332 PAD.n4320 1.1255
R41549 PAD.n8430 PAD.n8429 1.1255
R41550 PAD.n4322 PAD.n4321 1.1255
R41551 PAD.n8446 PAD.n8445 1.1255
R41552 PAD.n3978 PAD.n3977 1.1255
R41553 PAD.n8453 PAD.n8452 1.1255
R41554 PAD.n8470 PAD.n8469 1.1255
R41555 PAD.n3634 PAD.n3633 1.1255
R41556 PAD.n8478 PAD.n8477 1.1255
R41557 PAD.n8494 PAD.n8493 1.1255
R41558 PAD.n3288 PAD.n3287 1.1255
R41559 PAD.n8502 PAD.n8501 1.1255
R41560 PAD.n3290 PAD.n3289 1.1255
R41561 PAD.n8520 PAD.n8519 1.1255
R41562 PAD.n2947 PAD.n2904 1.1255
R41563 PAD.n8527 PAD.n8526 1.1255
R41564 PAD.n8833 PAD.n8832 1.1255
R41565 PAD.n2892 PAD.n2884 1.1255
R41566 PAD.n9128 PAD.n9127 1.1255
R41567 PAD.n9121 PAD.n2834 1.1255
R41568 PAD.n9141 PAD.n2833 1.1255
R41569 PAD.n9144 PAD.n9143 1.1255
R41570 PAD.n9151 PAD.n9150 1.1255
R41571 PAD.n9161 PAD.n2486 1.1255
R41572 PAD.n9164 PAD.n9163 1.1255
R41573 PAD.n9175 PAD.n9174 1.1255
R41574 PAD.n9185 PAD.n2138 1.1255
R41575 PAD.n9188 PAD.n9187 1.1255
R41576 PAD.n9190 PAD.n2046 1.1255
R41577 PAD.n2089 PAD.n2035 1.1255
R41578 PAD.n9457 PAD.n9456 1.1255
R41579 PAD.n9458 PAD.n1942 1.1255
R41580 PAD.n9460 PAD.n1986 1.1255
R41581 PAD.n1936 PAD.n1935 1.1255
R41582 PAD.n9723 PAD.n9722 1.1255
R41583 PAD.n9732 PAD.n9731 1.1255
R41584 PAD.n1593 PAD.n1585 1.1255
R41585 PAD.n9743 PAD.n9742 1.1255
R41586 PAD.n9746 PAD.n1489 1.1255
R41587 PAD.n9745 PAD.n1534 1.1255
R41588 PAD.n1532 PAD.n1148 1.1255
R41589 PAD.n10009 PAD.n10008 1.1255
R41590 PAD.n10016 PAD.n10015 1.1255
R41591 PAD.n1141 PAD.n1128 1.1255
R41592 PAD.n10363 PAD.n10362 1.1255
R41593 PAD.n1131 PAD.n1119 1.1255
R41594 PAD.n10373 PAD.n10372 1.1255
R41595 PAD.n1121 PAD.n1120 1.1255
R41596 PAD.n10390 PAD.n10389 1.1255
R41597 PAD.n777 PAD.n776 1.1255
R41598 PAD.n10397 PAD.n10396 1.1255
R41599 PAD.n10409 PAD.n10408 1.1255
R41600 PAD.n434 PAD.n426 1.1255
R41601 PAD.n10701 PAD.n10700 1.1255
R41602 PAD.n418 PAD.n372 1.1255
R41603 PAD.n10720 PAD.n10719 1.1255
R41604 PAD.n10717 PAD.n368 1.1255
R41605 PAD.n10727 PAD.n10726 1.1255
R41606 PAD.n11535 PAD.n11534 1.1255
R41607 PAD.n11533 PAD.n19 1.1255
R41608 PAD.n10753 PAD.n10752 1.1255
R41609 PAD.n10742 PAD.n10740 1.1255
R41610 PAD.n11522 PAD.n11521 1.1255
R41611 PAD.n11500 PAD.n10743 1.1255
R41612 PAD.n4 PAD.t15 0.9641
R41613 PAD.n7 PAD.t6 0.9641
R41614 PAD.n2 PAD.t4 0.9641
R41615 PAD.n11506 PAD.n11505 0.902975
R41616 PAD.n6376 PAD.n6375 0.902975
R41617 PAD.n11498 PAD.n11156 0.9005
R41618 PAD.n11497 PAD.n11154 0.9005
R41619 PAD.n11496 PAD.n11158 0.9005
R41620 PAD.n11305 PAD.n11153 0.9005
R41621 PAD.n11492 PAD.n11160 0.9005
R41622 PAD.n11491 PAD.n11152 0.9005
R41623 PAD.n11490 PAD.n11162 0.9005
R41624 PAD.n11307 PAD.n11151 0.9005
R41625 PAD.n11486 PAD.n11164 0.9005
R41626 PAD.n11485 PAD.n11150 0.9005
R41627 PAD.n11484 PAD.n11166 0.9005
R41628 PAD.n11309 PAD.n11149 0.9005
R41629 PAD.n11480 PAD.n11168 0.9005
R41630 PAD.n11479 PAD.n11148 0.9005
R41631 PAD.n11478 PAD.n11170 0.9005
R41632 PAD.n11311 PAD.n11147 0.9005
R41633 PAD.n11474 PAD.n11172 0.9005
R41634 PAD.n11473 PAD.n11146 0.9005
R41635 PAD.n11472 PAD.n11174 0.9005
R41636 PAD.n11313 PAD.n11145 0.9005
R41637 PAD.n11468 PAD.n11176 0.9005
R41638 PAD.n11467 PAD.n11144 0.9005
R41639 PAD.n11466 PAD.n11178 0.9005
R41640 PAD.n11315 PAD.n11143 0.9005
R41641 PAD.n11462 PAD.n11180 0.9005
R41642 PAD.n11461 PAD.n11142 0.9005
R41643 PAD.n11460 PAD.n11182 0.9005
R41644 PAD.n11317 PAD.n11141 0.9005
R41645 PAD.n11456 PAD.n11184 0.9005
R41646 PAD.n11455 PAD.n11140 0.9005
R41647 PAD.n11454 PAD.n11186 0.9005
R41648 PAD.n11319 PAD.n11139 0.9005
R41649 PAD.n11450 PAD.n11188 0.9005
R41650 PAD.n11449 PAD.n11138 0.9005
R41651 PAD.n11448 PAD.n11190 0.9005
R41652 PAD.n11321 PAD.n11137 0.9005
R41653 PAD.n11444 PAD.n11192 0.9005
R41654 PAD.n11443 PAD.n11136 0.9005
R41655 PAD.n11442 PAD.n11194 0.9005
R41656 PAD.n11323 PAD.n11135 0.9005
R41657 PAD.n11438 PAD.n11196 0.9005
R41658 PAD.n11437 PAD.n11134 0.9005
R41659 PAD.n11436 PAD.n11198 0.9005
R41660 PAD.n11325 PAD.n11133 0.9005
R41661 PAD.n11432 PAD.n11200 0.9005
R41662 PAD.n11431 PAD.n11132 0.9005
R41663 PAD.n11430 PAD.n11202 0.9005
R41664 PAD.n11327 PAD.n11131 0.9005
R41665 PAD.n11426 PAD.n11204 0.9005
R41666 PAD.n11425 PAD.n11130 0.9005
R41667 PAD.n11424 PAD.n11206 0.9005
R41668 PAD.n11329 PAD.n11129 0.9005
R41669 PAD.n11420 PAD.n11208 0.9005
R41670 PAD.n11419 PAD.n11128 0.9005
R41671 PAD.n11418 PAD.n11210 0.9005
R41672 PAD.n11331 PAD.n11127 0.9005
R41673 PAD.n11414 PAD.n11212 0.9005
R41674 PAD.n11413 PAD.n11126 0.9005
R41675 PAD.n11412 PAD.n11214 0.9005
R41676 PAD.n11333 PAD.n11125 0.9005
R41677 PAD.n11408 PAD.n11216 0.9005
R41678 PAD.n11407 PAD.n11124 0.9005
R41679 PAD.n11406 PAD.n11218 0.9005
R41680 PAD.n11335 PAD.n11123 0.9005
R41681 PAD.n11402 PAD.n11220 0.9005
R41682 PAD.n11401 PAD.n11122 0.9005
R41683 PAD.n11400 PAD.n11222 0.9005
R41684 PAD.n11337 PAD.n11121 0.9005
R41685 PAD.n11396 PAD.n11224 0.9005
R41686 PAD.n11395 PAD.n11120 0.9005
R41687 PAD.n11394 PAD.n11226 0.9005
R41688 PAD.n11339 PAD.n11119 0.9005
R41689 PAD.n11390 PAD.n11228 0.9005
R41690 PAD.n11389 PAD.n11118 0.9005
R41691 PAD.n11388 PAD.n11230 0.9005
R41692 PAD.n11341 PAD.n11117 0.9005
R41693 PAD.n11384 PAD.n11232 0.9005
R41694 PAD.n11383 PAD.n11116 0.9005
R41695 PAD.n11382 PAD.n11234 0.9005
R41696 PAD.n11343 PAD.n11115 0.9005
R41697 PAD.n11378 PAD.n11236 0.9005
R41698 PAD.n11377 PAD.n11114 0.9005
R41699 PAD.n11376 PAD.n11238 0.9005
R41700 PAD.n11345 PAD.n11113 0.9005
R41701 PAD.n11372 PAD.n11240 0.9005
R41702 PAD.n11371 PAD.n11112 0.9005
R41703 PAD.n11370 PAD.n11242 0.9005
R41704 PAD.n11347 PAD.n11111 0.9005
R41705 PAD.n11366 PAD.n11244 0.9005
R41706 PAD.n11365 PAD.n11110 0.9005
R41707 PAD.n11364 PAD.n11246 0.9005
R41708 PAD.n11349 PAD.n11109 0.9005
R41709 PAD.n11360 PAD.n11248 0.9005
R41710 PAD.n11359 PAD.n11108 0.9005
R41711 PAD.n11358 PAD.n11250 0.9005
R41712 PAD.n11351 PAD.n11107 0.9005
R41713 PAD.n11354 PAD.n11252 0.9005
R41714 PAD.n11353 PAD.n11106 0.9005
R41715 PAD.n11508 PAD.n11506 0.9005
R41716 PAD.n11497 PAD.n11304 0.9005
R41717 PAD.n11496 PAD.n11495 0.9005
R41718 PAD.n11494 PAD.n11305 0.9005
R41719 PAD.n11493 PAD.n11492 0.9005
R41720 PAD.n11491 PAD.n11306 0.9005
R41721 PAD.n11490 PAD.n11489 0.9005
R41722 PAD.n11488 PAD.n11307 0.9005
R41723 PAD.n11487 PAD.n11486 0.9005
R41724 PAD.n11485 PAD.n11308 0.9005
R41725 PAD.n11484 PAD.n11483 0.9005
R41726 PAD.n11482 PAD.n11309 0.9005
R41727 PAD.n11481 PAD.n11480 0.9005
R41728 PAD.n11479 PAD.n11310 0.9005
R41729 PAD.n11478 PAD.n11477 0.9005
R41730 PAD.n11476 PAD.n11311 0.9005
R41731 PAD.n11475 PAD.n11474 0.9005
R41732 PAD.n11473 PAD.n11312 0.9005
R41733 PAD.n11472 PAD.n11471 0.9005
R41734 PAD.n11470 PAD.n11313 0.9005
R41735 PAD.n11469 PAD.n11468 0.9005
R41736 PAD.n11467 PAD.n11314 0.9005
R41737 PAD.n11466 PAD.n11465 0.9005
R41738 PAD.n11464 PAD.n11315 0.9005
R41739 PAD.n11463 PAD.n11462 0.9005
R41740 PAD.n11461 PAD.n11316 0.9005
R41741 PAD.n11460 PAD.n11459 0.9005
R41742 PAD.n11458 PAD.n11317 0.9005
R41743 PAD.n11457 PAD.n11456 0.9005
R41744 PAD.n11455 PAD.n11318 0.9005
R41745 PAD.n11454 PAD.n11453 0.9005
R41746 PAD.n11452 PAD.n11319 0.9005
R41747 PAD.n11451 PAD.n11450 0.9005
R41748 PAD.n11449 PAD.n11320 0.9005
R41749 PAD.n11448 PAD.n11447 0.9005
R41750 PAD.n11446 PAD.n11321 0.9005
R41751 PAD.n11445 PAD.n11444 0.9005
R41752 PAD.n11443 PAD.n11322 0.9005
R41753 PAD.n11442 PAD.n11441 0.9005
R41754 PAD.n11440 PAD.n11323 0.9005
R41755 PAD.n11439 PAD.n11438 0.9005
R41756 PAD.n11437 PAD.n11324 0.9005
R41757 PAD.n11436 PAD.n11435 0.9005
R41758 PAD.n11434 PAD.n11325 0.9005
R41759 PAD.n11433 PAD.n11432 0.9005
R41760 PAD.n11431 PAD.n11326 0.9005
R41761 PAD.n11430 PAD.n11429 0.9005
R41762 PAD.n11428 PAD.n11327 0.9005
R41763 PAD.n11427 PAD.n11426 0.9005
R41764 PAD.n11425 PAD.n11328 0.9005
R41765 PAD.n11424 PAD.n11423 0.9005
R41766 PAD.n11422 PAD.n11329 0.9005
R41767 PAD.n11421 PAD.n11420 0.9005
R41768 PAD.n11419 PAD.n11330 0.9005
R41769 PAD.n11418 PAD.n11417 0.9005
R41770 PAD.n11416 PAD.n11331 0.9005
R41771 PAD.n11415 PAD.n11414 0.9005
R41772 PAD.n11413 PAD.n11332 0.9005
R41773 PAD.n11412 PAD.n11411 0.9005
R41774 PAD.n11410 PAD.n11333 0.9005
R41775 PAD.n11409 PAD.n11408 0.9005
R41776 PAD.n11407 PAD.n11334 0.9005
R41777 PAD.n11406 PAD.n11405 0.9005
R41778 PAD.n11404 PAD.n11335 0.9005
R41779 PAD.n11403 PAD.n11402 0.9005
R41780 PAD.n11401 PAD.n11336 0.9005
R41781 PAD.n11400 PAD.n11399 0.9005
R41782 PAD.n11398 PAD.n11337 0.9005
R41783 PAD.n11397 PAD.n11396 0.9005
R41784 PAD.n11395 PAD.n11338 0.9005
R41785 PAD.n11394 PAD.n11393 0.9005
R41786 PAD.n11392 PAD.n11339 0.9005
R41787 PAD.n11391 PAD.n11390 0.9005
R41788 PAD.n11389 PAD.n11340 0.9005
R41789 PAD.n11388 PAD.n11387 0.9005
R41790 PAD.n11386 PAD.n11341 0.9005
R41791 PAD.n11385 PAD.n11384 0.9005
R41792 PAD.n11383 PAD.n11342 0.9005
R41793 PAD.n11382 PAD.n11381 0.9005
R41794 PAD.n11380 PAD.n11343 0.9005
R41795 PAD.n11379 PAD.n11378 0.9005
R41796 PAD.n11377 PAD.n11344 0.9005
R41797 PAD.n11376 PAD.n11375 0.9005
R41798 PAD.n11374 PAD.n11345 0.9005
R41799 PAD.n11373 PAD.n11372 0.9005
R41800 PAD.n11371 PAD.n11346 0.9005
R41801 PAD.n11370 PAD.n11369 0.9005
R41802 PAD.n11368 PAD.n11347 0.9005
R41803 PAD.n11367 PAD.n11366 0.9005
R41804 PAD.n11365 PAD.n11348 0.9005
R41805 PAD.n11364 PAD.n11363 0.9005
R41806 PAD.n11362 PAD.n11349 0.9005
R41807 PAD.n11361 PAD.n11360 0.9005
R41808 PAD.n11359 PAD.n11350 0.9005
R41809 PAD.n11358 PAD.n11357 0.9005
R41810 PAD.n11356 PAD.n11351 0.9005
R41811 PAD.n11355 PAD.n11354 0.9005
R41812 PAD.n11353 PAD.n11352 0.9005
R41813 PAD.n11499 PAD.n11498 0.9005
R41814 PAD.n6226 PAD.n6225 0.9005
R41815 PAD.n6227 PAD.n6224 0.9005
R41816 PAD.n6229 PAD.n6228 0.9005
R41817 PAD.n6230 PAD.n6223 0.9005
R41818 PAD.n6232 PAD.n6231 0.9005
R41819 PAD.n6233 PAD.n6222 0.9005
R41820 PAD.n6235 PAD.n6234 0.9005
R41821 PAD.n6236 PAD.n6221 0.9005
R41822 PAD.n6238 PAD.n6237 0.9005
R41823 PAD.n6239 PAD.n6220 0.9005
R41824 PAD.n6241 PAD.n6240 0.9005
R41825 PAD.n6242 PAD.n6219 0.9005
R41826 PAD.n6244 PAD.n6243 0.9005
R41827 PAD.n6245 PAD.n6218 0.9005
R41828 PAD.n6247 PAD.n6246 0.9005
R41829 PAD.n6248 PAD.n6217 0.9005
R41830 PAD.n6250 PAD.n6249 0.9005
R41831 PAD.n6251 PAD.n6216 0.9005
R41832 PAD.n6253 PAD.n6252 0.9005
R41833 PAD.n6254 PAD.n6215 0.9005
R41834 PAD.n6256 PAD.n6255 0.9005
R41835 PAD.n6257 PAD.n6214 0.9005
R41836 PAD.n6259 PAD.n6258 0.9005
R41837 PAD.n6260 PAD.n6213 0.9005
R41838 PAD.n6262 PAD.n6261 0.9005
R41839 PAD.n6263 PAD.n6212 0.9005
R41840 PAD.n6265 PAD.n6264 0.9005
R41841 PAD.n6266 PAD.n6211 0.9005
R41842 PAD.n6268 PAD.n6267 0.9005
R41843 PAD.n6269 PAD.n6210 0.9005
R41844 PAD.n6271 PAD.n6270 0.9005
R41845 PAD.n6272 PAD.n6209 0.9005
R41846 PAD.n6274 PAD.n6273 0.9005
R41847 PAD.n6275 PAD.n6208 0.9005
R41848 PAD.n6277 PAD.n6276 0.9005
R41849 PAD.n6278 PAD.n6207 0.9005
R41850 PAD.n6280 PAD.n6279 0.9005
R41851 PAD.n6281 PAD.n6206 0.9005
R41852 PAD.n6283 PAD.n6282 0.9005
R41853 PAD.n6284 PAD.n6205 0.9005
R41854 PAD.n6286 PAD.n6285 0.9005
R41855 PAD.n6287 PAD.n6204 0.9005
R41856 PAD.n6289 PAD.n6288 0.9005
R41857 PAD.n6290 PAD.n6203 0.9005
R41858 PAD.n6292 PAD.n6291 0.9005
R41859 PAD.n6293 PAD.n6202 0.9005
R41860 PAD.n6295 PAD.n6294 0.9005
R41861 PAD.n6296 PAD.n6201 0.9005
R41862 PAD.n6298 PAD.n6297 0.9005
R41863 PAD.n6299 PAD.n6200 0.9005
R41864 PAD.n6301 PAD.n6300 0.9005
R41865 PAD.n6302 PAD.n6199 0.9005
R41866 PAD.n6304 PAD.n6303 0.9005
R41867 PAD.n6305 PAD.n6198 0.9005
R41868 PAD.n6307 PAD.n6306 0.9005
R41869 PAD.n6308 PAD.n6197 0.9005
R41870 PAD.n6310 PAD.n6309 0.9005
R41871 PAD.n6311 PAD.n6196 0.9005
R41872 PAD.n6313 PAD.n6312 0.9005
R41873 PAD.n6314 PAD.n6195 0.9005
R41874 PAD.n6316 PAD.n6315 0.9005
R41875 PAD.n6317 PAD.n6194 0.9005
R41876 PAD.n6319 PAD.n6318 0.9005
R41877 PAD.n6320 PAD.n6193 0.9005
R41878 PAD.n6322 PAD.n6321 0.9005
R41879 PAD.n6323 PAD.n6192 0.9005
R41880 PAD.n6325 PAD.n6324 0.9005
R41881 PAD.n6326 PAD.n6191 0.9005
R41882 PAD.n6328 PAD.n6327 0.9005
R41883 PAD.n6329 PAD.n6190 0.9005
R41884 PAD.n6331 PAD.n6330 0.9005
R41885 PAD.n6332 PAD.n6189 0.9005
R41886 PAD.n6334 PAD.n6333 0.9005
R41887 PAD.n6335 PAD.n6188 0.9005
R41888 PAD.n6337 PAD.n6336 0.9005
R41889 PAD.n6338 PAD.n6187 0.9005
R41890 PAD.n6340 PAD.n6339 0.9005
R41891 PAD.n6341 PAD.n6186 0.9005
R41892 PAD.n6343 PAD.n6342 0.9005
R41893 PAD.n6344 PAD.n6185 0.9005
R41894 PAD.n6346 PAD.n6345 0.9005
R41895 PAD.n6347 PAD.n6184 0.9005
R41896 PAD.n6349 PAD.n6348 0.9005
R41897 PAD.n6350 PAD.n6183 0.9005
R41898 PAD.n6352 PAD.n6351 0.9005
R41899 PAD.n6353 PAD.n6182 0.9005
R41900 PAD.n6355 PAD.n6354 0.9005
R41901 PAD.n6356 PAD.n6181 0.9005
R41902 PAD.n6358 PAD.n6357 0.9005
R41903 PAD.n6359 PAD.n6180 0.9005
R41904 PAD.n6361 PAD.n6360 0.9005
R41905 PAD.n6362 PAD.n6179 0.9005
R41906 PAD.n6364 PAD.n6363 0.9005
R41907 PAD.n6365 PAD.n6178 0.9005
R41908 PAD.n6367 PAD.n6366 0.9005
R41909 PAD.n6368 PAD.n6177 0.9005
R41910 PAD.n6370 PAD.n6369 0.9005
R41911 PAD.n6371 PAD.n5978 0.9005
R41912 PAD.n6370 PAD.n6032 0.9005
R41913 PAD.n6226 PAD.n6034 0.9005
R41914 PAD.n6227 PAD.n6030 0.9005
R41915 PAD.n6228 PAD.n6037 0.9005
R41916 PAD.n6223 PAD.n6029 0.9005
R41917 PAD.n6232 PAD.n6040 0.9005
R41918 PAD.n6233 PAD.n6028 0.9005
R41919 PAD.n6234 PAD.n6043 0.9005
R41920 PAD.n6221 PAD.n6027 0.9005
R41921 PAD.n6238 PAD.n6046 0.9005
R41922 PAD.n6239 PAD.n6026 0.9005
R41923 PAD.n6240 PAD.n6049 0.9005
R41924 PAD.n6219 PAD.n6025 0.9005
R41925 PAD.n6244 PAD.n6052 0.9005
R41926 PAD.n6245 PAD.n6024 0.9005
R41927 PAD.n6246 PAD.n6055 0.9005
R41928 PAD.n6217 PAD.n6023 0.9005
R41929 PAD.n6250 PAD.n6058 0.9005
R41930 PAD.n6251 PAD.n6022 0.9005
R41931 PAD.n6252 PAD.n6061 0.9005
R41932 PAD.n6215 PAD.n6021 0.9005
R41933 PAD.n6256 PAD.n6064 0.9005
R41934 PAD.n6257 PAD.n6020 0.9005
R41935 PAD.n6258 PAD.n6067 0.9005
R41936 PAD.n6213 PAD.n6019 0.9005
R41937 PAD.n6262 PAD.n6070 0.9005
R41938 PAD.n6263 PAD.n6018 0.9005
R41939 PAD.n6264 PAD.n6073 0.9005
R41940 PAD.n6211 PAD.n6017 0.9005
R41941 PAD.n6268 PAD.n6076 0.9005
R41942 PAD.n6269 PAD.n6016 0.9005
R41943 PAD.n6270 PAD.n6079 0.9005
R41944 PAD.n6209 PAD.n6015 0.9005
R41945 PAD.n6274 PAD.n6082 0.9005
R41946 PAD.n6275 PAD.n6014 0.9005
R41947 PAD.n6276 PAD.n6085 0.9005
R41948 PAD.n6207 PAD.n6013 0.9005
R41949 PAD.n6280 PAD.n6088 0.9005
R41950 PAD.n6281 PAD.n6012 0.9005
R41951 PAD.n6282 PAD.n6091 0.9005
R41952 PAD.n6205 PAD.n6011 0.9005
R41953 PAD.n6286 PAD.n6094 0.9005
R41954 PAD.n6287 PAD.n6010 0.9005
R41955 PAD.n6288 PAD.n6097 0.9005
R41956 PAD.n6203 PAD.n6009 0.9005
R41957 PAD.n6292 PAD.n6100 0.9005
R41958 PAD.n6293 PAD.n6008 0.9005
R41959 PAD.n6294 PAD.n6103 0.9005
R41960 PAD.n6201 PAD.n6007 0.9005
R41961 PAD.n6298 PAD.n6106 0.9005
R41962 PAD.n6299 PAD.n6006 0.9005
R41963 PAD.n6300 PAD.n6109 0.9005
R41964 PAD.n6199 PAD.n6005 0.9005
R41965 PAD.n6304 PAD.n6112 0.9005
R41966 PAD.n6305 PAD.n6004 0.9005
R41967 PAD.n6306 PAD.n6115 0.9005
R41968 PAD.n6197 PAD.n6003 0.9005
R41969 PAD.n6310 PAD.n6118 0.9005
R41970 PAD.n6311 PAD.n6002 0.9005
R41971 PAD.n6312 PAD.n6121 0.9005
R41972 PAD.n6195 PAD.n6001 0.9005
R41973 PAD.n6316 PAD.n6124 0.9005
R41974 PAD.n6317 PAD.n6000 0.9005
R41975 PAD.n6318 PAD.n6127 0.9005
R41976 PAD.n6193 PAD.n5999 0.9005
R41977 PAD.n6322 PAD.n6130 0.9005
R41978 PAD.n6323 PAD.n5998 0.9005
R41979 PAD.n6324 PAD.n6133 0.9005
R41980 PAD.n6191 PAD.n5997 0.9005
R41981 PAD.n6328 PAD.n6136 0.9005
R41982 PAD.n6329 PAD.n5996 0.9005
R41983 PAD.n6330 PAD.n6139 0.9005
R41984 PAD.n6189 PAD.n5995 0.9005
R41985 PAD.n6334 PAD.n6142 0.9005
R41986 PAD.n6335 PAD.n5994 0.9005
R41987 PAD.n6336 PAD.n6145 0.9005
R41988 PAD.n6187 PAD.n5993 0.9005
R41989 PAD.n6340 PAD.n6148 0.9005
R41990 PAD.n6341 PAD.n5992 0.9005
R41991 PAD.n6342 PAD.n6151 0.9005
R41992 PAD.n6185 PAD.n5991 0.9005
R41993 PAD.n6346 PAD.n6154 0.9005
R41994 PAD.n6347 PAD.n5990 0.9005
R41995 PAD.n6348 PAD.n6157 0.9005
R41996 PAD.n6183 PAD.n5989 0.9005
R41997 PAD.n6352 PAD.n6160 0.9005
R41998 PAD.n6353 PAD.n5988 0.9005
R41999 PAD.n6354 PAD.n6163 0.9005
R42000 PAD.n6181 PAD.n5987 0.9005
R42001 PAD.n6358 PAD.n6166 0.9005
R42002 PAD.n6359 PAD.n5986 0.9005
R42003 PAD.n6360 PAD.n6169 0.9005
R42004 PAD.n6179 PAD.n5985 0.9005
R42005 PAD.n6364 PAD.n6172 0.9005
R42006 PAD.n6365 PAD.n5984 0.9005
R42007 PAD.n6366 PAD.n6175 0.9005
R42008 PAD.n6177 PAD.n5983 0.9005
R42009 PAD.n6372 PAD.n6371 0.9005
R42010 PAD.n6375 PAD.n6374 0.9005
R42011 PAD.n7809 PAD.n7808 0.87242
R42012 PAD.n11540 PAD.n11539 0.87242
R42013 PAD.n7810 PAD.n7809 0.79382
R42014 PAD.n3636 PAD.n10 0.79382
R42015 PAD.n11541 PAD.n11 0.79382
R42016 PAD.n11540 PAD.n12 0.79382
R42017 PAD.n11512 PAD.n11090 0.761105
R42018 PAD.n6385 PAD.n5956 0.758684
R42019 PAD.n11104 PAD.n11093 0.7505
R42020 PAD.n11515 PAD.n11514 0.7505
R42021 PAD.n11102 PAD.n11101 0.7505
R42022 PAD.n11516 PAD.n11515 0.7505
R42023 PAD.n11093 PAD.n11091 0.7505
R42024 PAD.n6389 PAD.n6388 0.7505
R42025 PAD.n5959 PAD.n5957 0.7505
R42026 PAD.n5969 PAD.n5959 0.7505
R42027 PAD.n6388 PAD.n6387 0.7505
R42028 PAD.n5968 PAD.n5967 0.7505
R42029 PAD.n10366 PAD.n13 0.407313
R42030 PAD.n9171 PAD.n9168 0.407313
R42031 PAD.n7812 PAD.n7811 0.407313
R42032 PAD.n8473 PAD.n3637 0.407223
R42033 PAD.n11517 PAD.n11090 0.384314
R42034 PAD.n6390 PAD.n5956 0.38336
R42035 PAD.n6 PAD.n5 0.204443
R42036 PAD.n1 PAD.n0 0.199354
R42037 PAD.n9 PAD.n3 0.102972
R42038 PAD PAD.n9 0.0996761
R42039 PAD PAD.n11542 0.09545
R42040 PAD.n1 PAD 0.0811609
R42041 PAD.n8 PAD 0.0811609
R42042 PAD.n7809 PAD.n10 0.0791
R42043 PAD.n11541 PAD.n11540 0.0791
R42044 PAD.n9 PAD.n8 0.0751609
R42045 PAD.n3 PAD 0.0548109
R42046 PAD.n6 PAD 0.0548109
R42047 PAD.n5 PAD 0.0548109
R42048 PAD.n3636 PAD.n11 0.0433318
R42049 PAD.n11542 PAD.n10 0.03995
R42050 PAD.n11542 PAD.n11541 0.03965
R42051 PAD.n7517 PAD.n7209 0.0380882
R42052 PAD.n7513 PAD.n7209 0.0380882
R42053 PAD.n7513 PAD.n7510 0.0380882
R42054 PAD.n7510 PAD.n7506 0.0380882
R42055 PAD.n7506 PAD.n7229 0.0380882
R42056 PAD.n7502 PAD.n7229 0.0380882
R42057 PAD.n7502 PAD.n7498 0.0380882
R42058 PAD.n7498 PAD.n7494 0.0380882
R42059 PAD.n7494 PAD.n7231 0.0380882
R42060 PAD.n7490 PAD.n7231 0.0380882
R42061 PAD.n7490 PAD.n7486 0.0380882
R42062 PAD.n7486 PAD.n7482 0.0380882
R42063 PAD.n7482 PAD.n7233 0.0380882
R42064 PAD.n7478 PAD.n7233 0.0380882
R42065 PAD.n7478 PAD.n7474 0.0380882
R42066 PAD.n7474 PAD.n7470 0.0380882
R42067 PAD.n7470 PAD.n7235 0.0380882
R42068 PAD.n7466 PAD.n7235 0.0380882
R42069 PAD.n7466 PAD.n7462 0.0380882
R42070 PAD.n7462 PAD.n7458 0.0380882
R42071 PAD.n7458 PAD.n7237 0.0380882
R42072 PAD.n7454 PAD.n7237 0.0380882
R42073 PAD.n7454 PAD.n7450 0.0380882
R42074 PAD.n7450 PAD.n7446 0.0380882
R42075 PAD.n7446 PAD.n7239 0.0380882
R42076 PAD.n7442 PAD.n7239 0.0380882
R42077 PAD.n7442 PAD.n7438 0.0380882
R42078 PAD.n7438 PAD.n7434 0.0380882
R42079 PAD.n7434 PAD.n7241 0.0380882
R42080 PAD.n7430 PAD.n7241 0.0380882
R42081 PAD.n7430 PAD.n7426 0.0380882
R42082 PAD.n7426 PAD.n7422 0.0380882
R42083 PAD.n7422 PAD.n7243 0.0380882
R42084 PAD.n7418 PAD.n7243 0.0380882
R42085 PAD.n7418 PAD.n7414 0.0380882
R42086 PAD.n7414 PAD.n7410 0.0380882
R42087 PAD.n7410 PAD.n7245 0.0380882
R42088 PAD.n7406 PAD.n7245 0.0380882
R42089 PAD.n7406 PAD.n7402 0.0380882
R42090 PAD.n7402 PAD.n7398 0.0380882
R42091 PAD.n7398 PAD.n7247 0.0380882
R42092 PAD.n7394 PAD.n7247 0.0380882
R42093 PAD.n7394 PAD.n7390 0.0380882
R42094 PAD.n7390 PAD.n7386 0.0380882
R42095 PAD.n7386 PAD.n7249 0.0380882
R42096 PAD.n7382 PAD.n7249 0.0380882
R42097 PAD.n7382 PAD.n7378 0.0380882
R42098 PAD.n7378 PAD.n7374 0.0380882
R42099 PAD.n7374 PAD.n7251 0.0380882
R42100 PAD.n7370 PAD.n7251 0.0380882
R42101 PAD.n7370 PAD.n7366 0.0380882
R42102 PAD.n7366 PAD.n7362 0.0380882
R42103 PAD.n7362 PAD.n7253 0.0380882
R42104 PAD.n7358 PAD.n7253 0.0380882
R42105 PAD.n7358 PAD.n7354 0.0380882
R42106 PAD.n7354 PAD.n7350 0.0380882
R42107 PAD.n7350 PAD.n7255 0.0380882
R42108 PAD.n7346 PAD.n7255 0.0380882
R42109 PAD.n7346 PAD.n7342 0.0380882
R42110 PAD.n7342 PAD.n7338 0.0380882
R42111 PAD.n7338 PAD.n7257 0.0380882
R42112 PAD.n7334 PAD.n7257 0.0380882
R42113 PAD.n7334 PAD.n7330 0.0380882
R42114 PAD.n7330 PAD.n7326 0.0380882
R42115 PAD.n7326 PAD.n7259 0.0380882
R42116 PAD.n7322 PAD.n7259 0.0380882
R42117 PAD.n7322 PAD.n7318 0.0380882
R42118 PAD.n7318 PAD.n7314 0.0380882
R42119 PAD.n7314 PAD.n7261 0.0380882
R42120 PAD.n7310 PAD.n7261 0.0380882
R42121 PAD.n7310 PAD.n7306 0.0380882
R42122 PAD.n7306 PAD.n7302 0.0380882
R42123 PAD.n7302 PAD.n7263 0.0380882
R42124 PAD.n7298 PAD.n7263 0.0380882
R42125 PAD.n7298 PAD.n7294 0.0380882
R42126 PAD.n7294 PAD.n7290 0.0380882
R42127 PAD.n7290 PAD.n7265 0.0380882
R42128 PAD.n7286 PAD.n7265 0.0380882
R42129 PAD.n7286 PAD.n7282 0.0380882
R42130 PAD.n7282 PAD.n7278 0.0380882
R42131 PAD.n7278 PAD.n7267 0.0380882
R42132 PAD.n7274 PAD.n7267 0.0380882
R42133 PAD.n7274 PAD.n7270 0.0380882
R42134 PAD.n7516 PAD.n7515 0.0380882
R42135 PAD.n7515 PAD.n7514 0.0380882
R42136 PAD.n7514 PAD.n7228 0.0380882
R42137 PAD.n7505 PAD.n7228 0.0380882
R42138 PAD.n7505 PAD.n7504 0.0380882
R42139 PAD.n7504 PAD.n7503 0.0380882
R42140 PAD.n7503 PAD.n7230 0.0380882
R42141 PAD.n7493 PAD.n7230 0.0380882
R42142 PAD.n7493 PAD.n7492 0.0380882
R42143 PAD.n7492 PAD.n7491 0.0380882
R42144 PAD.n7491 PAD.n7232 0.0380882
R42145 PAD.n7481 PAD.n7232 0.0380882
R42146 PAD.n7481 PAD.n7480 0.0380882
R42147 PAD.n7480 PAD.n7479 0.0380882
R42148 PAD.n7479 PAD.n7234 0.0380882
R42149 PAD.n7469 PAD.n7234 0.0380882
R42150 PAD.n7469 PAD.n7468 0.0380882
R42151 PAD.n7468 PAD.n7467 0.0380882
R42152 PAD.n7467 PAD.n7236 0.0380882
R42153 PAD.n7457 PAD.n7236 0.0380882
R42154 PAD.n7457 PAD.n7456 0.0380882
R42155 PAD.n7456 PAD.n7455 0.0380882
R42156 PAD.n7455 PAD.n7238 0.0380882
R42157 PAD.n7445 PAD.n7238 0.0380882
R42158 PAD.n7445 PAD.n7444 0.0380882
R42159 PAD.n7444 PAD.n7443 0.0380882
R42160 PAD.n7443 PAD.n7240 0.0380882
R42161 PAD.n7433 PAD.n7240 0.0380882
R42162 PAD.n7433 PAD.n7432 0.0380882
R42163 PAD.n7432 PAD.n7431 0.0380882
R42164 PAD.n7431 PAD.n7242 0.0380882
R42165 PAD.n7421 PAD.n7242 0.0380882
R42166 PAD.n7421 PAD.n7420 0.0380882
R42167 PAD.n7420 PAD.n7419 0.0380882
R42168 PAD.n7419 PAD.n7244 0.0380882
R42169 PAD.n7409 PAD.n7244 0.0380882
R42170 PAD.n7409 PAD.n7408 0.0380882
R42171 PAD.n7408 PAD.n7407 0.0380882
R42172 PAD.n7407 PAD.n7246 0.0380882
R42173 PAD.n7397 PAD.n7246 0.0380882
R42174 PAD.n7397 PAD.n7396 0.0380882
R42175 PAD.n7396 PAD.n7395 0.0380882
R42176 PAD.n7395 PAD.n7248 0.0380882
R42177 PAD.n7385 PAD.n7248 0.0380882
R42178 PAD.n7385 PAD.n7384 0.0380882
R42179 PAD.n7384 PAD.n7383 0.0380882
R42180 PAD.n7383 PAD.n7250 0.0380882
R42181 PAD.n7373 PAD.n7250 0.0380882
R42182 PAD.n7373 PAD.n7372 0.0380882
R42183 PAD.n7372 PAD.n7371 0.0380882
R42184 PAD.n7371 PAD.n7252 0.0380882
R42185 PAD.n7361 PAD.n7252 0.0380882
R42186 PAD.n7361 PAD.n7360 0.0380882
R42187 PAD.n7360 PAD.n7359 0.0380882
R42188 PAD.n7359 PAD.n7254 0.0380882
R42189 PAD.n7349 PAD.n7254 0.0380882
R42190 PAD.n7349 PAD.n7348 0.0380882
R42191 PAD.n7348 PAD.n7347 0.0380882
R42192 PAD.n7347 PAD.n7256 0.0380882
R42193 PAD.n7337 PAD.n7256 0.0380882
R42194 PAD.n7337 PAD.n7336 0.0380882
R42195 PAD.n7336 PAD.n7335 0.0380882
R42196 PAD.n7335 PAD.n7258 0.0380882
R42197 PAD.n7325 PAD.n7258 0.0380882
R42198 PAD.n7325 PAD.n7324 0.0380882
R42199 PAD.n7324 PAD.n7323 0.0380882
R42200 PAD.n7323 PAD.n7260 0.0380882
R42201 PAD.n7313 PAD.n7260 0.0380882
R42202 PAD.n7313 PAD.n7312 0.0380882
R42203 PAD.n7312 PAD.n7311 0.0380882
R42204 PAD.n7311 PAD.n7262 0.0380882
R42205 PAD.n7301 PAD.n7262 0.0380882
R42206 PAD.n7301 PAD.n7300 0.0380882
R42207 PAD.n7300 PAD.n7299 0.0380882
R42208 PAD.n7299 PAD.n7264 0.0380882
R42209 PAD.n7289 PAD.n7264 0.0380882
R42210 PAD.n7289 PAD.n7288 0.0380882
R42211 PAD.n7288 PAD.n7287 0.0380882
R42212 PAD.n7287 PAD.n7266 0.0380882
R42213 PAD.n7277 PAD.n7266 0.0380882
R42214 PAD.n7277 PAD.n7276 0.0380882
R42215 PAD.n7276 PAD.n7275 0.0380882
R42216 PAD.n7275 PAD.n7268 0.0380882
R42217 PAD.n121 PAD.n120 0.0380882
R42218 PAD.n122 PAD.n121 0.0380882
R42219 PAD.n122 PAD.n115 0.0380882
R42220 PAD.n132 PAD.n115 0.0380882
R42221 PAD.n133 PAD.n132 0.0380882
R42222 PAD.n134 PAD.n133 0.0380882
R42223 PAD.n134 PAD.n113 0.0380882
R42224 PAD.n144 PAD.n113 0.0380882
R42225 PAD.n145 PAD.n144 0.0380882
R42226 PAD.n146 PAD.n145 0.0380882
R42227 PAD.n146 PAD.n111 0.0380882
R42228 PAD.n156 PAD.n111 0.0380882
R42229 PAD.n157 PAD.n156 0.0380882
R42230 PAD.n158 PAD.n157 0.0380882
R42231 PAD.n158 PAD.n109 0.0380882
R42232 PAD.n168 PAD.n109 0.0380882
R42233 PAD.n169 PAD.n168 0.0380882
R42234 PAD.n170 PAD.n169 0.0380882
R42235 PAD.n170 PAD.n107 0.0380882
R42236 PAD.n180 PAD.n107 0.0380882
R42237 PAD.n181 PAD.n180 0.0380882
R42238 PAD.n182 PAD.n181 0.0380882
R42239 PAD.n182 PAD.n105 0.0380882
R42240 PAD.n192 PAD.n105 0.0380882
R42241 PAD.n193 PAD.n192 0.0380882
R42242 PAD.n194 PAD.n193 0.0380882
R42243 PAD.n194 PAD.n103 0.0380882
R42244 PAD.n204 PAD.n103 0.0380882
R42245 PAD.n205 PAD.n204 0.0380882
R42246 PAD.n206 PAD.n205 0.0380882
R42247 PAD.n206 PAD.n101 0.0380882
R42248 PAD.n216 PAD.n101 0.0380882
R42249 PAD.n217 PAD.n216 0.0380882
R42250 PAD.n218 PAD.n217 0.0380882
R42251 PAD.n218 PAD.n99 0.0380882
R42252 PAD.n228 PAD.n99 0.0380882
R42253 PAD.n229 PAD.n228 0.0380882
R42254 PAD.n230 PAD.n229 0.0380882
R42255 PAD.n230 PAD.n97 0.0380882
R42256 PAD.n240 PAD.n97 0.0380882
R42257 PAD.n241 PAD.n240 0.0380882
R42258 PAD.n242 PAD.n241 0.0380882
R42259 PAD.n242 PAD.n95 0.0380882
R42260 PAD.n252 PAD.n95 0.0380882
R42261 PAD.n253 PAD.n252 0.0380882
R42262 PAD.n254 PAD.n253 0.0380882
R42263 PAD.n254 PAD.n93 0.0380882
R42264 PAD.n264 PAD.n93 0.0380882
R42265 PAD.n265 PAD.n264 0.0380882
R42266 PAD.n266 PAD.n265 0.0380882
R42267 PAD.n266 PAD.n91 0.0380882
R42268 PAD.n276 PAD.n91 0.0380882
R42269 PAD.n277 PAD.n276 0.0380882
R42270 PAD.n278 PAD.n277 0.0380882
R42271 PAD.n278 PAD.n89 0.0380882
R42272 PAD.n288 PAD.n89 0.0380882
R42273 PAD.n289 PAD.n288 0.0380882
R42274 PAD.n290 PAD.n289 0.0380882
R42275 PAD.n290 PAD.n87 0.0380882
R42276 PAD.n300 PAD.n87 0.0380882
R42277 PAD.n301 PAD.n300 0.0380882
R42278 PAD.n302 PAD.n301 0.0380882
R42279 PAD.n302 PAD.n85 0.0380882
R42280 PAD.n312 PAD.n85 0.0380882
R42281 PAD.n313 PAD.n312 0.0380882
R42282 PAD.n314 PAD.n313 0.0380882
R42283 PAD.n314 PAD.n83 0.0380882
R42284 PAD.n324 PAD.n83 0.0380882
R42285 PAD.n325 PAD.n324 0.0380882
R42286 PAD.n326 PAD.n325 0.0380882
R42287 PAD.n326 PAD.n81 0.0380882
R42288 PAD.n336 PAD.n81 0.0380882
R42289 PAD.n337 PAD.n336 0.0380882
R42290 PAD.n338 PAD.n337 0.0380882
R42291 PAD.n338 PAD.n79 0.0380882
R42292 PAD.n348 PAD.n79 0.0380882
R42293 PAD.n349 PAD.n348 0.0380882
R42294 PAD.n350 PAD.n349 0.0380882
R42295 PAD.n350 PAD.n77 0.0380882
R42296 PAD.n360 PAD.n77 0.0380882
R42297 PAD.n361 PAD.n360 0.0380882
R42298 PAD.n362 PAD.n361 0.0380882
R42299 PAD.n362 PAD.n26 0.0380882
R42300 PAD.n10695 PAD.n10694 0.0380882
R42301 PAD.n10694 PAD.n10691 0.0380882
R42302 PAD.n10691 PAD.n10414 0.0380882
R42303 PAD.n10687 PAD.n10414 0.0380882
R42304 PAD.n10687 PAD.n10683 0.0380882
R42305 PAD.n10683 PAD.n10682 0.0380882
R42306 PAD.n10682 PAD.n10419 0.0380882
R42307 PAD.n10678 PAD.n10419 0.0380882
R42308 PAD.n10678 PAD.n10674 0.0380882
R42309 PAD.n10674 PAD.n10673 0.0380882
R42310 PAD.n10673 PAD.n10424 0.0380882
R42311 PAD.n10669 PAD.n10424 0.0380882
R42312 PAD.n10669 PAD.n10665 0.0380882
R42313 PAD.n10665 PAD.n10664 0.0380882
R42314 PAD.n10664 PAD.n10429 0.0380882
R42315 PAD.n10660 PAD.n10429 0.0380882
R42316 PAD.n10660 PAD.n10656 0.0380882
R42317 PAD.n10656 PAD.n10655 0.0380882
R42318 PAD.n10655 PAD.n10434 0.0380882
R42319 PAD.n10651 PAD.n10434 0.0380882
R42320 PAD.n10651 PAD.n10647 0.0380882
R42321 PAD.n10647 PAD.n10646 0.0380882
R42322 PAD.n10646 PAD.n10439 0.0380882
R42323 PAD.n10642 PAD.n10439 0.0380882
R42324 PAD.n10642 PAD.n10638 0.0380882
R42325 PAD.n10638 PAD.n10637 0.0380882
R42326 PAD.n10637 PAD.n10444 0.0380882
R42327 PAD.n10633 PAD.n10444 0.0380882
R42328 PAD.n10633 PAD.n10629 0.0380882
R42329 PAD.n10629 PAD.n10628 0.0380882
R42330 PAD.n10628 PAD.n10449 0.0380882
R42331 PAD.n10624 PAD.n10449 0.0380882
R42332 PAD.n10624 PAD.n10620 0.0380882
R42333 PAD.n10620 PAD.n10619 0.0380882
R42334 PAD.n10619 PAD.n10454 0.0380882
R42335 PAD.n10615 PAD.n10454 0.0380882
R42336 PAD.n10615 PAD.n10611 0.0380882
R42337 PAD.n10611 PAD.n10610 0.0380882
R42338 PAD.n10610 PAD.n10459 0.0380882
R42339 PAD.n10606 PAD.n10459 0.0380882
R42340 PAD.n10606 PAD.n10602 0.0380882
R42341 PAD.n10602 PAD.n10601 0.0380882
R42342 PAD.n10601 PAD.n10464 0.0380882
R42343 PAD.n10597 PAD.n10464 0.0380882
R42344 PAD.n10597 PAD.n10593 0.0380882
R42345 PAD.n10593 PAD.n10592 0.0380882
R42346 PAD.n10592 PAD.n10469 0.0380882
R42347 PAD.n10588 PAD.n10469 0.0380882
R42348 PAD.n10588 PAD.n10584 0.0380882
R42349 PAD.n10584 PAD.n10583 0.0380882
R42350 PAD.n10583 PAD.n10474 0.0380882
R42351 PAD.n10579 PAD.n10474 0.0380882
R42352 PAD.n10579 PAD.n10575 0.0380882
R42353 PAD.n10575 PAD.n10574 0.0380882
R42354 PAD.n10574 PAD.n10479 0.0380882
R42355 PAD.n10570 PAD.n10479 0.0380882
R42356 PAD.n10570 PAD.n10566 0.0380882
R42357 PAD.n10566 PAD.n10565 0.0380882
R42358 PAD.n10565 PAD.n10484 0.0380882
R42359 PAD.n10561 PAD.n10484 0.0380882
R42360 PAD.n10561 PAD.n10557 0.0380882
R42361 PAD.n10557 PAD.n10556 0.0380882
R42362 PAD.n10556 PAD.n10489 0.0380882
R42363 PAD.n10552 PAD.n10489 0.0380882
R42364 PAD.n10552 PAD.n10548 0.0380882
R42365 PAD.n10548 PAD.n10547 0.0380882
R42366 PAD.n10547 PAD.n10494 0.0380882
R42367 PAD.n10543 PAD.n10494 0.0380882
R42368 PAD.n10543 PAD.n10539 0.0380882
R42369 PAD.n10539 PAD.n10538 0.0380882
R42370 PAD.n10538 PAD.n10499 0.0380882
R42371 PAD.n10534 PAD.n10499 0.0380882
R42372 PAD.n10534 PAD.n10530 0.0380882
R42373 PAD.n10530 PAD.n10529 0.0380882
R42374 PAD.n10529 PAD.n10504 0.0380882
R42375 PAD.n10525 PAD.n10504 0.0380882
R42376 PAD.n10525 PAD.n10521 0.0380882
R42377 PAD.n10521 PAD.n10520 0.0380882
R42378 PAD.n10520 PAD.n10509 0.0380882
R42379 PAD.n10516 PAD.n10509 0.0380882
R42380 PAD.n10516 PAD.n420 0.0380882
R42381 PAD.n10712 PAD.n420 0.0380882
R42382 PAD.n10712 PAD.n416 0.0380882
R42383 PAD.n10696 PAD.n10413 0.0380882
R42384 PAD.n10690 PAD.n10413 0.0380882
R42385 PAD.n10690 PAD.n10689 0.0380882
R42386 PAD.n10689 PAD.n10688 0.0380882
R42387 PAD.n10688 PAD.n10418 0.0380882
R42388 PAD.n10681 PAD.n10418 0.0380882
R42389 PAD.n10681 PAD.n10680 0.0380882
R42390 PAD.n10680 PAD.n10679 0.0380882
R42391 PAD.n10679 PAD.n10423 0.0380882
R42392 PAD.n10672 PAD.n10423 0.0380882
R42393 PAD.n10672 PAD.n10671 0.0380882
R42394 PAD.n10671 PAD.n10670 0.0380882
R42395 PAD.n10670 PAD.n10428 0.0380882
R42396 PAD.n10663 PAD.n10428 0.0380882
R42397 PAD.n10663 PAD.n10662 0.0380882
R42398 PAD.n10662 PAD.n10661 0.0380882
R42399 PAD.n10661 PAD.n10433 0.0380882
R42400 PAD.n10654 PAD.n10433 0.0380882
R42401 PAD.n10654 PAD.n10653 0.0380882
R42402 PAD.n10653 PAD.n10652 0.0380882
R42403 PAD.n10652 PAD.n10438 0.0380882
R42404 PAD.n10645 PAD.n10438 0.0380882
R42405 PAD.n10645 PAD.n10644 0.0380882
R42406 PAD.n10644 PAD.n10643 0.0380882
R42407 PAD.n10643 PAD.n10443 0.0380882
R42408 PAD.n10636 PAD.n10443 0.0380882
R42409 PAD.n10636 PAD.n10635 0.0380882
R42410 PAD.n10635 PAD.n10634 0.0380882
R42411 PAD.n10634 PAD.n10448 0.0380882
R42412 PAD.n10627 PAD.n10448 0.0380882
R42413 PAD.n10627 PAD.n10626 0.0380882
R42414 PAD.n10626 PAD.n10625 0.0380882
R42415 PAD.n10625 PAD.n10453 0.0380882
R42416 PAD.n10618 PAD.n10453 0.0380882
R42417 PAD.n10618 PAD.n10617 0.0380882
R42418 PAD.n10617 PAD.n10616 0.0380882
R42419 PAD.n10616 PAD.n10458 0.0380882
R42420 PAD.n10609 PAD.n10458 0.0380882
R42421 PAD.n10609 PAD.n10608 0.0380882
R42422 PAD.n10608 PAD.n10607 0.0380882
R42423 PAD.n10607 PAD.n10463 0.0380882
R42424 PAD.n10600 PAD.n10463 0.0380882
R42425 PAD.n10600 PAD.n10599 0.0380882
R42426 PAD.n10599 PAD.n10598 0.0380882
R42427 PAD.n10598 PAD.n10468 0.0380882
R42428 PAD.n10591 PAD.n10468 0.0380882
R42429 PAD.n10591 PAD.n10590 0.0380882
R42430 PAD.n10590 PAD.n10589 0.0380882
R42431 PAD.n10589 PAD.n10473 0.0380882
R42432 PAD.n10582 PAD.n10473 0.0380882
R42433 PAD.n10582 PAD.n10581 0.0380882
R42434 PAD.n10581 PAD.n10580 0.0380882
R42435 PAD.n10580 PAD.n10478 0.0380882
R42436 PAD.n10573 PAD.n10478 0.0380882
R42437 PAD.n10573 PAD.n10572 0.0380882
R42438 PAD.n10572 PAD.n10571 0.0380882
R42439 PAD.n10571 PAD.n10483 0.0380882
R42440 PAD.n10564 PAD.n10483 0.0380882
R42441 PAD.n10564 PAD.n10563 0.0380882
R42442 PAD.n10563 PAD.n10562 0.0380882
R42443 PAD.n10562 PAD.n10488 0.0380882
R42444 PAD.n10555 PAD.n10488 0.0380882
R42445 PAD.n10555 PAD.n10554 0.0380882
R42446 PAD.n10554 PAD.n10553 0.0380882
R42447 PAD.n10553 PAD.n10493 0.0380882
R42448 PAD.n10546 PAD.n10493 0.0380882
R42449 PAD.n10546 PAD.n10545 0.0380882
R42450 PAD.n10545 PAD.n10544 0.0380882
R42451 PAD.n10544 PAD.n10498 0.0380882
R42452 PAD.n10537 PAD.n10498 0.0380882
R42453 PAD.n10537 PAD.n10536 0.0380882
R42454 PAD.n10536 PAD.n10535 0.0380882
R42455 PAD.n10535 PAD.n10503 0.0380882
R42456 PAD.n10528 PAD.n10503 0.0380882
R42457 PAD.n10528 PAD.n10527 0.0380882
R42458 PAD.n10527 PAD.n10526 0.0380882
R42459 PAD.n10526 PAD.n10508 0.0380882
R42460 PAD.n10519 PAD.n10508 0.0380882
R42461 PAD.n10519 PAD.n10518 0.0380882
R42462 PAD.n10518 PAD.n10517 0.0380882
R42463 PAD.n10517 PAD.n421 0.0380882
R42464 PAD.n10711 PAD.n421 0.0380882
R42465 PAD.n10711 PAD.n10710 0.0380882
R42466 PAD.n522 PAD.n520 0.0380882
R42467 PAD.n530 PAD.n520 0.0380882
R42468 PAD.n530 PAD.n518 0.0380882
R42469 PAD.n534 PAD.n518 0.0380882
R42470 PAD.n534 PAD.n516 0.0380882
R42471 PAD.n542 PAD.n516 0.0380882
R42472 PAD.n542 PAD.n514 0.0380882
R42473 PAD.n546 PAD.n514 0.0380882
R42474 PAD.n546 PAD.n512 0.0380882
R42475 PAD.n554 PAD.n512 0.0380882
R42476 PAD.n554 PAD.n510 0.0380882
R42477 PAD.n558 PAD.n510 0.0380882
R42478 PAD.n558 PAD.n508 0.0380882
R42479 PAD.n566 PAD.n508 0.0380882
R42480 PAD.n566 PAD.n506 0.0380882
R42481 PAD.n570 PAD.n506 0.0380882
R42482 PAD.n570 PAD.n504 0.0380882
R42483 PAD.n578 PAD.n504 0.0380882
R42484 PAD.n578 PAD.n502 0.0380882
R42485 PAD.n582 PAD.n502 0.0380882
R42486 PAD.n582 PAD.n500 0.0380882
R42487 PAD.n590 PAD.n500 0.0380882
R42488 PAD.n590 PAD.n498 0.0380882
R42489 PAD.n594 PAD.n498 0.0380882
R42490 PAD.n594 PAD.n496 0.0380882
R42491 PAD.n602 PAD.n496 0.0380882
R42492 PAD.n602 PAD.n494 0.0380882
R42493 PAD.n606 PAD.n494 0.0380882
R42494 PAD.n606 PAD.n492 0.0380882
R42495 PAD.n614 PAD.n492 0.0380882
R42496 PAD.n614 PAD.n490 0.0380882
R42497 PAD.n618 PAD.n490 0.0380882
R42498 PAD.n618 PAD.n488 0.0380882
R42499 PAD.n626 PAD.n488 0.0380882
R42500 PAD.n626 PAD.n486 0.0380882
R42501 PAD.n630 PAD.n486 0.0380882
R42502 PAD.n630 PAD.n484 0.0380882
R42503 PAD.n638 PAD.n484 0.0380882
R42504 PAD.n638 PAD.n482 0.0380882
R42505 PAD.n642 PAD.n482 0.0380882
R42506 PAD.n642 PAD.n480 0.0380882
R42507 PAD.n650 PAD.n480 0.0380882
R42508 PAD.n650 PAD.n478 0.0380882
R42509 PAD.n654 PAD.n478 0.0380882
R42510 PAD.n654 PAD.n476 0.0380882
R42511 PAD.n662 PAD.n476 0.0380882
R42512 PAD.n662 PAD.n474 0.0380882
R42513 PAD.n666 PAD.n474 0.0380882
R42514 PAD.n666 PAD.n472 0.0380882
R42515 PAD.n674 PAD.n472 0.0380882
R42516 PAD.n674 PAD.n470 0.0380882
R42517 PAD.n678 PAD.n470 0.0380882
R42518 PAD.n678 PAD.n468 0.0380882
R42519 PAD.n686 PAD.n468 0.0380882
R42520 PAD.n686 PAD.n466 0.0380882
R42521 PAD.n690 PAD.n466 0.0380882
R42522 PAD.n690 PAD.n464 0.0380882
R42523 PAD.n698 PAD.n464 0.0380882
R42524 PAD.n698 PAD.n462 0.0380882
R42525 PAD.n702 PAD.n462 0.0380882
R42526 PAD.n702 PAD.n460 0.0380882
R42527 PAD.n710 PAD.n460 0.0380882
R42528 PAD.n710 PAD.n458 0.0380882
R42529 PAD.n714 PAD.n458 0.0380882
R42530 PAD.n714 PAD.n456 0.0380882
R42531 PAD.n722 PAD.n456 0.0380882
R42532 PAD.n722 PAD.n454 0.0380882
R42533 PAD.n726 PAD.n454 0.0380882
R42534 PAD.n726 PAD.n452 0.0380882
R42535 PAD.n734 PAD.n452 0.0380882
R42536 PAD.n734 PAD.n450 0.0380882
R42537 PAD.n738 PAD.n450 0.0380882
R42538 PAD.n738 PAD.n448 0.0380882
R42539 PAD.n746 PAD.n448 0.0380882
R42540 PAD.n746 PAD.n446 0.0380882
R42541 PAD.n750 PAD.n446 0.0380882
R42542 PAD.n750 PAD.n444 0.0380882
R42543 PAD.n758 PAD.n444 0.0380882
R42544 PAD.n758 PAD.n442 0.0380882
R42545 PAD.n763 PAD.n442 0.0380882
R42546 PAD.n763 PAD.n440 0.0380882
R42547 PAD.n440 PAD.n439 0.0380882
R42548 PAD.n771 PAD.n439 0.0380882
R42549 PAD.n521 PAD.n519 0.0380882
R42550 PAD.n531 PAD.n519 0.0380882
R42551 PAD.n532 PAD.n531 0.0380882
R42552 PAD.n533 PAD.n532 0.0380882
R42553 PAD.n533 PAD.n515 0.0380882
R42554 PAD.n543 PAD.n515 0.0380882
R42555 PAD.n544 PAD.n543 0.0380882
R42556 PAD.n545 PAD.n544 0.0380882
R42557 PAD.n545 PAD.n511 0.0380882
R42558 PAD.n555 PAD.n511 0.0380882
R42559 PAD.n556 PAD.n555 0.0380882
R42560 PAD.n557 PAD.n556 0.0380882
R42561 PAD.n557 PAD.n507 0.0380882
R42562 PAD.n567 PAD.n507 0.0380882
R42563 PAD.n568 PAD.n567 0.0380882
R42564 PAD.n569 PAD.n568 0.0380882
R42565 PAD.n569 PAD.n503 0.0380882
R42566 PAD.n579 PAD.n503 0.0380882
R42567 PAD.n580 PAD.n579 0.0380882
R42568 PAD.n581 PAD.n580 0.0380882
R42569 PAD.n581 PAD.n499 0.0380882
R42570 PAD.n591 PAD.n499 0.0380882
R42571 PAD.n592 PAD.n591 0.0380882
R42572 PAD.n593 PAD.n592 0.0380882
R42573 PAD.n593 PAD.n495 0.0380882
R42574 PAD.n603 PAD.n495 0.0380882
R42575 PAD.n604 PAD.n603 0.0380882
R42576 PAD.n605 PAD.n604 0.0380882
R42577 PAD.n605 PAD.n491 0.0380882
R42578 PAD.n615 PAD.n491 0.0380882
R42579 PAD.n616 PAD.n615 0.0380882
R42580 PAD.n617 PAD.n616 0.0380882
R42581 PAD.n617 PAD.n487 0.0380882
R42582 PAD.n627 PAD.n487 0.0380882
R42583 PAD.n628 PAD.n627 0.0380882
R42584 PAD.n629 PAD.n628 0.0380882
R42585 PAD.n629 PAD.n483 0.0380882
R42586 PAD.n639 PAD.n483 0.0380882
R42587 PAD.n640 PAD.n639 0.0380882
R42588 PAD.n641 PAD.n640 0.0380882
R42589 PAD.n641 PAD.n479 0.0380882
R42590 PAD.n651 PAD.n479 0.0380882
R42591 PAD.n652 PAD.n651 0.0380882
R42592 PAD.n653 PAD.n652 0.0380882
R42593 PAD.n653 PAD.n475 0.0380882
R42594 PAD.n663 PAD.n475 0.0380882
R42595 PAD.n664 PAD.n663 0.0380882
R42596 PAD.n665 PAD.n664 0.0380882
R42597 PAD.n665 PAD.n471 0.0380882
R42598 PAD.n675 PAD.n471 0.0380882
R42599 PAD.n676 PAD.n675 0.0380882
R42600 PAD.n677 PAD.n676 0.0380882
R42601 PAD.n677 PAD.n467 0.0380882
R42602 PAD.n687 PAD.n467 0.0380882
R42603 PAD.n688 PAD.n687 0.0380882
R42604 PAD.n689 PAD.n688 0.0380882
R42605 PAD.n689 PAD.n463 0.0380882
R42606 PAD.n699 PAD.n463 0.0380882
R42607 PAD.n700 PAD.n699 0.0380882
R42608 PAD.n701 PAD.n700 0.0380882
R42609 PAD.n701 PAD.n459 0.0380882
R42610 PAD.n711 PAD.n459 0.0380882
R42611 PAD.n712 PAD.n711 0.0380882
R42612 PAD.n713 PAD.n712 0.0380882
R42613 PAD.n713 PAD.n455 0.0380882
R42614 PAD.n723 PAD.n455 0.0380882
R42615 PAD.n724 PAD.n723 0.0380882
R42616 PAD.n725 PAD.n724 0.0380882
R42617 PAD.n725 PAD.n451 0.0380882
R42618 PAD.n735 PAD.n451 0.0380882
R42619 PAD.n736 PAD.n735 0.0380882
R42620 PAD.n737 PAD.n736 0.0380882
R42621 PAD.n737 PAD.n447 0.0380882
R42622 PAD.n747 PAD.n447 0.0380882
R42623 PAD.n748 PAD.n747 0.0380882
R42624 PAD.n749 PAD.n748 0.0380882
R42625 PAD.n749 PAD.n443 0.0380882
R42626 PAD.n759 PAD.n443 0.0380882
R42627 PAD.n760 PAD.n759 0.0380882
R42628 PAD.n762 PAD.n760 0.0380882
R42629 PAD.n762 PAD.n761 0.0380882
R42630 PAD.n761 PAD.n438 0.0380882
R42631 PAD.n772 PAD.n438 0.0380882
R42632 PAD.n872 PAD.n871 0.0380882
R42633 PAD.n876 PAD.n871 0.0380882
R42634 PAD.n880 PAD.n876 0.0380882
R42635 PAD.n884 PAD.n880 0.0380882
R42636 PAD.n884 PAD.n867 0.0380882
R42637 PAD.n888 PAD.n867 0.0380882
R42638 PAD.n892 PAD.n888 0.0380882
R42639 PAD.n896 PAD.n892 0.0380882
R42640 PAD.n896 PAD.n865 0.0380882
R42641 PAD.n900 PAD.n865 0.0380882
R42642 PAD.n904 PAD.n900 0.0380882
R42643 PAD.n908 PAD.n904 0.0380882
R42644 PAD.n908 PAD.n863 0.0380882
R42645 PAD.n912 PAD.n863 0.0380882
R42646 PAD.n916 PAD.n912 0.0380882
R42647 PAD.n920 PAD.n916 0.0380882
R42648 PAD.n920 PAD.n861 0.0380882
R42649 PAD.n924 PAD.n861 0.0380882
R42650 PAD.n928 PAD.n924 0.0380882
R42651 PAD.n932 PAD.n928 0.0380882
R42652 PAD.n932 PAD.n859 0.0380882
R42653 PAD.n936 PAD.n859 0.0380882
R42654 PAD.n940 PAD.n936 0.0380882
R42655 PAD.n944 PAD.n940 0.0380882
R42656 PAD.n944 PAD.n857 0.0380882
R42657 PAD.n948 PAD.n857 0.0380882
R42658 PAD.n952 PAD.n948 0.0380882
R42659 PAD.n956 PAD.n952 0.0380882
R42660 PAD.n956 PAD.n855 0.0380882
R42661 PAD.n960 PAD.n855 0.0380882
R42662 PAD.n964 PAD.n960 0.0380882
R42663 PAD.n968 PAD.n964 0.0380882
R42664 PAD.n968 PAD.n853 0.0380882
R42665 PAD.n972 PAD.n853 0.0380882
R42666 PAD.n976 PAD.n972 0.0380882
R42667 PAD.n980 PAD.n976 0.0380882
R42668 PAD.n980 PAD.n851 0.0380882
R42669 PAD.n984 PAD.n851 0.0380882
R42670 PAD.n988 PAD.n984 0.0380882
R42671 PAD.n992 PAD.n988 0.0380882
R42672 PAD.n992 PAD.n849 0.0380882
R42673 PAD.n996 PAD.n849 0.0380882
R42674 PAD.n1000 PAD.n996 0.0380882
R42675 PAD.n1004 PAD.n1000 0.0380882
R42676 PAD.n1004 PAD.n847 0.0380882
R42677 PAD.n1008 PAD.n847 0.0380882
R42678 PAD.n1012 PAD.n1008 0.0380882
R42679 PAD.n1016 PAD.n1012 0.0380882
R42680 PAD.n1016 PAD.n845 0.0380882
R42681 PAD.n1020 PAD.n845 0.0380882
R42682 PAD.n1024 PAD.n1020 0.0380882
R42683 PAD.n1028 PAD.n1024 0.0380882
R42684 PAD.n1028 PAD.n843 0.0380882
R42685 PAD.n1032 PAD.n843 0.0380882
R42686 PAD.n1036 PAD.n1032 0.0380882
R42687 PAD.n1040 PAD.n1036 0.0380882
R42688 PAD.n1040 PAD.n841 0.0380882
R42689 PAD.n1044 PAD.n841 0.0380882
R42690 PAD.n1048 PAD.n1044 0.0380882
R42691 PAD.n1052 PAD.n1048 0.0380882
R42692 PAD.n1052 PAD.n839 0.0380882
R42693 PAD.n1056 PAD.n839 0.0380882
R42694 PAD.n1060 PAD.n1056 0.0380882
R42695 PAD.n1064 PAD.n1060 0.0380882
R42696 PAD.n1064 PAD.n837 0.0380882
R42697 PAD.n1068 PAD.n837 0.0380882
R42698 PAD.n1072 PAD.n1068 0.0380882
R42699 PAD.n1076 PAD.n1072 0.0380882
R42700 PAD.n1076 PAD.n835 0.0380882
R42701 PAD.n1080 PAD.n835 0.0380882
R42702 PAD.n1084 PAD.n1080 0.0380882
R42703 PAD.n1088 PAD.n1084 0.0380882
R42704 PAD.n1088 PAD.n833 0.0380882
R42705 PAD.n1092 PAD.n833 0.0380882
R42706 PAD.n1096 PAD.n1092 0.0380882
R42707 PAD.n1100 PAD.n1096 0.0380882
R42708 PAD.n1100 PAD.n831 0.0380882
R42709 PAD.n1104 PAD.n831 0.0380882
R42710 PAD.n1108 PAD.n1104 0.0380882
R42711 PAD.n1112 PAD.n1108 0.0380882
R42712 PAD.n1112 PAD.n829 0.0380882
R42713 PAD.n10384 PAD.n829 0.0380882
R42714 PAD.n10384 PAD.n826 0.0380882
R42715 PAD.n874 PAD.n873 0.0380882
R42716 PAD.n875 PAD.n874 0.0380882
R42717 PAD.n875 PAD.n868 0.0380882
R42718 PAD.n885 PAD.n868 0.0380882
R42719 PAD.n886 PAD.n885 0.0380882
R42720 PAD.n887 PAD.n886 0.0380882
R42721 PAD.n887 PAD.n866 0.0380882
R42722 PAD.n897 PAD.n866 0.0380882
R42723 PAD.n898 PAD.n897 0.0380882
R42724 PAD.n899 PAD.n898 0.0380882
R42725 PAD.n899 PAD.n864 0.0380882
R42726 PAD.n909 PAD.n864 0.0380882
R42727 PAD.n910 PAD.n909 0.0380882
R42728 PAD.n911 PAD.n910 0.0380882
R42729 PAD.n911 PAD.n862 0.0380882
R42730 PAD.n921 PAD.n862 0.0380882
R42731 PAD.n922 PAD.n921 0.0380882
R42732 PAD.n923 PAD.n922 0.0380882
R42733 PAD.n923 PAD.n860 0.0380882
R42734 PAD.n933 PAD.n860 0.0380882
R42735 PAD.n934 PAD.n933 0.0380882
R42736 PAD.n935 PAD.n934 0.0380882
R42737 PAD.n935 PAD.n858 0.0380882
R42738 PAD.n945 PAD.n858 0.0380882
R42739 PAD.n946 PAD.n945 0.0380882
R42740 PAD.n947 PAD.n946 0.0380882
R42741 PAD.n947 PAD.n856 0.0380882
R42742 PAD.n957 PAD.n856 0.0380882
R42743 PAD.n958 PAD.n957 0.0380882
R42744 PAD.n959 PAD.n958 0.0380882
R42745 PAD.n959 PAD.n854 0.0380882
R42746 PAD.n969 PAD.n854 0.0380882
R42747 PAD.n970 PAD.n969 0.0380882
R42748 PAD.n971 PAD.n970 0.0380882
R42749 PAD.n971 PAD.n852 0.0380882
R42750 PAD.n981 PAD.n852 0.0380882
R42751 PAD.n982 PAD.n981 0.0380882
R42752 PAD.n983 PAD.n982 0.0380882
R42753 PAD.n983 PAD.n850 0.0380882
R42754 PAD.n993 PAD.n850 0.0380882
R42755 PAD.n994 PAD.n993 0.0380882
R42756 PAD.n995 PAD.n994 0.0380882
R42757 PAD.n995 PAD.n848 0.0380882
R42758 PAD.n1005 PAD.n848 0.0380882
R42759 PAD.n1006 PAD.n1005 0.0380882
R42760 PAD.n1007 PAD.n1006 0.0380882
R42761 PAD.n1007 PAD.n846 0.0380882
R42762 PAD.n1017 PAD.n846 0.0380882
R42763 PAD.n1018 PAD.n1017 0.0380882
R42764 PAD.n1019 PAD.n1018 0.0380882
R42765 PAD.n1019 PAD.n844 0.0380882
R42766 PAD.n1029 PAD.n844 0.0380882
R42767 PAD.n1030 PAD.n1029 0.0380882
R42768 PAD.n1031 PAD.n1030 0.0380882
R42769 PAD.n1031 PAD.n842 0.0380882
R42770 PAD.n1041 PAD.n842 0.0380882
R42771 PAD.n1042 PAD.n1041 0.0380882
R42772 PAD.n1043 PAD.n1042 0.0380882
R42773 PAD.n1043 PAD.n840 0.0380882
R42774 PAD.n1053 PAD.n840 0.0380882
R42775 PAD.n1054 PAD.n1053 0.0380882
R42776 PAD.n1055 PAD.n1054 0.0380882
R42777 PAD.n1055 PAD.n838 0.0380882
R42778 PAD.n1065 PAD.n838 0.0380882
R42779 PAD.n1066 PAD.n1065 0.0380882
R42780 PAD.n1067 PAD.n1066 0.0380882
R42781 PAD.n1067 PAD.n836 0.0380882
R42782 PAD.n1077 PAD.n836 0.0380882
R42783 PAD.n1078 PAD.n1077 0.0380882
R42784 PAD.n1079 PAD.n1078 0.0380882
R42785 PAD.n1079 PAD.n834 0.0380882
R42786 PAD.n1089 PAD.n834 0.0380882
R42787 PAD.n1090 PAD.n1089 0.0380882
R42788 PAD.n1091 PAD.n1090 0.0380882
R42789 PAD.n1091 PAD.n832 0.0380882
R42790 PAD.n1101 PAD.n832 0.0380882
R42791 PAD.n1102 PAD.n1101 0.0380882
R42792 PAD.n1103 PAD.n1102 0.0380882
R42793 PAD.n1103 PAD.n830 0.0380882
R42794 PAD.n1113 PAD.n830 0.0380882
R42795 PAD.n1114 PAD.n1113 0.0380882
R42796 PAD.n10383 PAD.n1114 0.0380882
R42797 PAD.n10383 PAD.n10382 0.0380882
R42798 PAD.n10105 PAD.n10104 0.0380882
R42799 PAD.n10113 PAD.n10104 0.0380882
R42800 PAD.n10113 PAD.n10102 0.0380882
R42801 PAD.n10117 PAD.n10102 0.0380882
R42802 PAD.n10117 PAD.n10100 0.0380882
R42803 PAD.n10125 PAD.n10100 0.0380882
R42804 PAD.n10125 PAD.n10098 0.0380882
R42805 PAD.n10129 PAD.n10098 0.0380882
R42806 PAD.n10129 PAD.n10096 0.0380882
R42807 PAD.n10137 PAD.n10096 0.0380882
R42808 PAD.n10137 PAD.n10094 0.0380882
R42809 PAD.n10141 PAD.n10094 0.0380882
R42810 PAD.n10141 PAD.n10092 0.0380882
R42811 PAD.n10149 PAD.n10092 0.0380882
R42812 PAD.n10149 PAD.n10090 0.0380882
R42813 PAD.n10153 PAD.n10090 0.0380882
R42814 PAD.n10153 PAD.n10088 0.0380882
R42815 PAD.n10161 PAD.n10088 0.0380882
R42816 PAD.n10161 PAD.n10086 0.0380882
R42817 PAD.n10165 PAD.n10086 0.0380882
R42818 PAD.n10165 PAD.n10084 0.0380882
R42819 PAD.n10173 PAD.n10084 0.0380882
R42820 PAD.n10173 PAD.n10082 0.0380882
R42821 PAD.n10177 PAD.n10082 0.0380882
R42822 PAD.n10177 PAD.n10080 0.0380882
R42823 PAD.n10185 PAD.n10080 0.0380882
R42824 PAD.n10185 PAD.n10078 0.0380882
R42825 PAD.n10189 PAD.n10078 0.0380882
R42826 PAD.n10189 PAD.n10076 0.0380882
R42827 PAD.n10197 PAD.n10076 0.0380882
R42828 PAD.n10197 PAD.n10074 0.0380882
R42829 PAD.n10201 PAD.n10074 0.0380882
R42830 PAD.n10201 PAD.n10072 0.0380882
R42831 PAD.n10209 PAD.n10072 0.0380882
R42832 PAD.n10209 PAD.n10070 0.0380882
R42833 PAD.n10213 PAD.n10070 0.0380882
R42834 PAD.n10213 PAD.n10068 0.0380882
R42835 PAD.n10221 PAD.n10068 0.0380882
R42836 PAD.n10221 PAD.n10066 0.0380882
R42837 PAD.n10225 PAD.n10066 0.0380882
R42838 PAD.n10225 PAD.n10064 0.0380882
R42839 PAD.n10233 PAD.n10064 0.0380882
R42840 PAD.n10233 PAD.n10062 0.0380882
R42841 PAD.n10237 PAD.n10062 0.0380882
R42842 PAD.n10237 PAD.n10060 0.0380882
R42843 PAD.n10245 PAD.n10060 0.0380882
R42844 PAD.n10245 PAD.n10058 0.0380882
R42845 PAD.n10249 PAD.n10058 0.0380882
R42846 PAD.n10249 PAD.n10056 0.0380882
R42847 PAD.n10257 PAD.n10056 0.0380882
R42848 PAD.n10257 PAD.n10054 0.0380882
R42849 PAD.n10261 PAD.n10054 0.0380882
R42850 PAD.n10261 PAD.n10052 0.0380882
R42851 PAD.n10269 PAD.n10052 0.0380882
R42852 PAD.n10269 PAD.n10050 0.0380882
R42853 PAD.n10273 PAD.n10050 0.0380882
R42854 PAD.n10273 PAD.n10048 0.0380882
R42855 PAD.n10281 PAD.n10048 0.0380882
R42856 PAD.n10281 PAD.n10046 0.0380882
R42857 PAD.n10285 PAD.n10046 0.0380882
R42858 PAD.n10285 PAD.n10044 0.0380882
R42859 PAD.n10293 PAD.n10044 0.0380882
R42860 PAD.n10293 PAD.n10042 0.0380882
R42861 PAD.n10297 PAD.n10042 0.0380882
R42862 PAD.n10297 PAD.n10040 0.0380882
R42863 PAD.n10305 PAD.n10040 0.0380882
R42864 PAD.n10305 PAD.n10038 0.0380882
R42865 PAD.n10309 PAD.n10038 0.0380882
R42866 PAD.n10309 PAD.n10036 0.0380882
R42867 PAD.n10317 PAD.n10036 0.0380882
R42868 PAD.n10317 PAD.n10034 0.0380882
R42869 PAD.n10321 PAD.n10034 0.0380882
R42870 PAD.n10321 PAD.n10032 0.0380882
R42871 PAD.n10329 PAD.n10032 0.0380882
R42872 PAD.n10329 PAD.n10030 0.0380882
R42873 PAD.n10333 PAD.n10030 0.0380882
R42874 PAD.n10333 PAD.n10028 0.0380882
R42875 PAD.n10341 PAD.n10028 0.0380882
R42876 PAD.n10341 PAD.n10026 0.0380882
R42877 PAD.n10346 PAD.n10026 0.0380882
R42878 PAD.n10346 PAD.n10024 0.0380882
R42879 PAD.n10024 PAD.n10023 0.0380882
R42880 PAD.n10354 PAD.n10023 0.0380882
R42881 PAD.n10103 PAD.n1124 0.0380882
R42882 PAD.n10114 PAD.n10103 0.0380882
R42883 PAD.n10115 PAD.n10114 0.0380882
R42884 PAD.n10116 PAD.n10115 0.0380882
R42885 PAD.n10116 PAD.n10099 0.0380882
R42886 PAD.n10126 PAD.n10099 0.0380882
R42887 PAD.n10127 PAD.n10126 0.0380882
R42888 PAD.n10128 PAD.n10127 0.0380882
R42889 PAD.n10128 PAD.n10095 0.0380882
R42890 PAD.n10138 PAD.n10095 0.0380882
R42891 PAD.n10139 PAD.n10138 0.0380882
R42892 PAD.n10140 PAD.n10139 0.0380882
R42893 PAD.n10140 PAD.n10091 0.0380882
R42894 PAD.n10150 PAD.n10091 0.0380882
R42895 PAD.n10151 PAD.n10150 0.0380882
R42896 PAD.n10152 PAD.n10151 0.0380882
R42897 PAD.n10152 PAD.n10087 0.0380882
R42898 PAD.n10162 PAD.n10087 0.0380882
R42899 PAD.n10163 PAD.n10162 0.0380882
R42900 PAD.n10164 PAD.n10163 0.0380882
R42901 PAD.n10164 PAD.n10083 0.0380882
R42902 PAD.n10174 PAD.n10083 0.0380882
R42903 PAD.n10175 PAD.n10174 0.0380882
R42904 PAD.n10176 PAD.n10175 0.0380882
R42905 PAD.n10176 PAD.n10079 0.0380882
R42906 PAD.n10186 PAD.n10079 0.0380882
R42907 PAD.n10187 PAD.n10186 0.0380882
R42908 PAD.n10188 PAD.n10187 0.0380882
R42909 PAD.n10188 PAD.n10075 0.0380882
R42910 PAD.n10198 PAD.n10075 0.0380882
R42911 PAD.n10199 PAD.n10198 0.0380882
R42912 PAD.n10200 PAD.n10199 0.0380882
R42913 PAD.n10200 PAD.n10071 0.0380882
R42914 PAD.n10210 PAD.n10071 0.0380882
R42915 PAD.n10211 PAD.n10210 0.0380882
R42916 PAD.n10212 PAD.n10211 0.0380882
R42917 PAD.n10212 PAD.n10067 0.0380882
R42918 PAD.n10222 PAD.n10067 0.0380882
R42919 PAD.n10223 PAD.n10222 0.0380882
R42920 PAD.n10224 PAD.n10223 0.0380882
R42921 PAD.n10224 PAD.n10063 0.0380882
R42922 PAD.n10234 PAD.n10063 0.0380882
R42923 PAD.n10235 PAD.n10234 0.0380882
R42924 PAD.n10236 PAD.n10235 0.0380882
R42925 PAD.n10236 PAD.n10059 0.0380882
R42926 PAD.n10246 PAD.n10059 0.0380882
R42927 PAD.n10247 PAD.n10246 0.0380882
R42928 PAD.n10248 PAD.n10247 0.0380882
R42929 PAD.n10248 PAD.n10055 0.0380882
R42930 PAD.n10258 PAD.n10055 0.0380882
R42931 PAD.n10259 PAD.n10258 0.0380882
R42932 PAD.n10260 PAD.n10259 0.0380882
R42933 PAD.n10260 PAD.n10051 0.0380882
R42934 PAD.n10270 PAD.n10051 0.0380882
R42935 PAD.n10271 PAD.n10270 0.0380882
R42936 PAD.n10272 PAD.n10271 0.0380882
R42937 PAD.n10272 PAD.n10047 0.0380882
R42938 PAD.n10282 PAD.n10047 0.0380882
R42939 PAD.n10283 PAD.n10282 0.0380882
R42940 PAD.n10284 PAD.n10283 0.0380882
R42941 PAD.n10284 PAD.n10043 0.0380882
R42942 PAD.n10294 PAD.n10043 0.0380882
R42943 PAD.n10295 PAD.n10294 0.0380882
R42944 PAD.n10296 PAD.n10295 0.0380882
R42945 PAD.n10296 PAD.n10039 0.0380882
R42946 PAD.n10306 PAD.n10039 0.0380882
R42947 PAD.n10307 PAD.n10306 0.0380882
R42948 PAD.n10308 PAD.n10307 0.0380882
R42949 PAD.n10308 PAD.n10035 0.0380882
R42950 PAD.n10318 PAD.n10035 0.0380882
R42951 PAD.n10319 PAD.n10318 0.0380882
R42952 PAD.n10320 PAD.n10319 0.0380882
R42953 PAD.n10320 PAD.n10031 0.0380882
R42954 PAD.n10330 PAD.n10031 0.0380882
R42955 PAD.n10331 PAD.n10330 0.0380882
R42956 PAD.n10332 PAD.n10331 0.0380882
R42957 PAD.n10332 PAD.n10027 0.0380882
R42958 PAD.n10342 PAD.n10027 0.0380882
R42959 PAD.n10343 PAD.n10342 0.0380882
R42960 PAD.n10345 PAD.n10343 0.0380882
R42961 PAD.n10345 PAD.n10344 0.0380882
R42962 PAD.n10344 PAD.n10022 0.0380882
R42963 PAD.n10355 PAD.n10022 0.0380882
R42964 PAD.n1480 PAD.n1479 0.0380882
R42965 PAD.n1479 PAD.n1193 0.0380882
R42966 PAD.n1475 PAD.n1193 0.0380882
R42967 PAD.n1475 PAD.n1471 0.0380882
R42968 PAD.n1471 PAD.n1470 0.0380882
R42969 PAD.n1470 PAD.n1195 0.0380882
R42970 PAD.n1466 PAD.n1195 0.0380882
R42971 PAD.n1466 PAD.n1462 0.0380882
R42972 PAD.n1462 PAD.n1461 0.0380882
R42973 PAD.n1461 PAD.n1200 0.0380882
R42974 PAD.n1457 PAD.n1200 0.0380882
R42975 PAD.n1457 PAD.n1453 0.0380882
R42976 PAD.n1453 PAD.n1452 0.0380882
R42977 PAD.n1452 PAD.n1205 0.0380882
R42978 PAD.n1448 PAD.n1205 0.0380882
R42979 PAD.n1448 PAD.n1444 0.0380882
R42980 PAD.n1444 PAD.n1443 0.0380882
R42981 PAD.n1443 PAD.n1210 0.0380882
R42982 PAD.n1439 PAD.n1210 0.0380882
R42983 PAD.n1439 PAD.n1435 0.0380882
R42984 PAD.n1435 PAD.n1434 0.0380882
R42985 PAD.n1434 PAD.n1215 0.0380882
R42986 PAD.n1430 PAD.n1215 0.0380882
R42987 PAD.n1430 PAD.n1426 0.0380882
R42988 PAD.n1426 PAD.n1425 0.0380882
R42989 PAD.n1425 PAD.n1220 0.0380882
R42990 PAD.n1421 PAD.n1220 0.0380882
R42991 PAD.n1421 PAD.n1417 0.0380882
R42992 PAD.n1417 PAD.n1416 0.0380882
R42993 PAD.n1416 PAD.n1225 0.0380882
R42994 PAD.n1412 PAD.n1225 0.0380882
R42995 PAD.n1412 PAD.n1408 0.0380882
R42996 PAD.n1408 PAD.n1407 0.0380882
R42997 PAD.n1407 PAD.n1230 0.0380882
R42998 PAD.n1403 PAD.n1230 0.0380882
R42999 PAD.n1403 PAD.n1399 0.0380882
R43000 PAD.n1399 PAD.n1398 0.0380882
R43001 PAD.n1398 PAD.n1235 0.0380882
R43002 PAD.n1394 PAD.n1235 0.0380882
R43003 PAD.n1394 PAD.n1390 0.0380882
R43004 PAD.n1390 PAD.n1389 0.0380882
R43005 PAD.n1389 PAD.n1240 0.0380882
R43006 PAD.n1385 PAD.n1240 0.0380882
R43007 PAD.n1385 PAD.n1381 0.0380882
R43008 PAD.n1381 PAD.n1380 0.0380882
R43009 PAD.n1380 PAD.n1245 0.0380882
R43010 PAD.n1376 PAD.n1245 0.0380882
R43011 PAD.n1376 PAD.n1372 0.0380882
R43012 PAD.n1372 PAD.n1371 0.0380882
R43013 PAD.n1371 PAD.n1250 0.0380882
R43014 PAD.n1367 PAD.n1250 0.0380882
R43015 PAD.n1367 PAD.n1363 0.0380882
R43016 PAD.n1363 PAD.n1362 0.0380882
R43017 PAD.n1362 PAD.n1255 0.0380882
R43018 PAD.n1358 PAD.n1255 0.0380882
R43019 PAD.n1358 PAD.n1354 0.0380882
R43020 PAD.n1354 PAD.n1353 0.0380882
R43021 PAD.n1353 PAD.n1260 0.0380882
R43022 PAD.n1349 PAD.n1260 0.0380882
R43023 PAD.n1349 PAD.n1345 0.0380882
R43024 PAD.n1345 PAD.n1344 0.0380882
R43025 PAD.n1344 PAD.n1265 0.0380882
R43026 PAD.n1340 PAD.n1265 0.0380882
R43027 PAD.n1340 PAD.n1336 0.0380882
R43028 PAD.n1336 PAD.n1335 0.0380882
R43029 PAD.n1335 PAD.n1270 0.0380882
R43030 PAD.n1331 PAD.n1270 0.0380882
R43031 PAD.n1331 PAD.n1327 0.0380882
R43032 PAD.n1327 PAD.n1326 0.0380882
R43033 PAD.n1326 PAD.n1275 0.0380882
R43034 PAD.n1322 PAD.n1275 0.0380882
R43035 PAD.n1322 PAD.n1318 0.0380882
R43036 PAD.n1318 PAD.n1317 0.0380882
R43037 PAD.n1317 PAD.n1280 0.0380882
R43038 PAD.n1313 PAD.n1280 0.0380882
R43039 PAD.n1313 PAD.n1309 0.0380882
R43040 PAD.n1309 PAD.n1308 0.0380882
R43041 PAD.n1308 PAD.n1285 0.0380882
R43042 PAD.n1304 PAD.n1285 0.0380882
R43043 PAD.n1304 PAD.n1300 0.0380882
R43044 PAD.n1300 PAD.n1299 0.0380882
R43045 PAD.n1299 PAD.n1290 0.0380882
R43046 PAD.n1295 PAD.n1290 0.0380882
R43047 PAD.n1478 PAD.n1145 0.0380882
R43048 PAD.n1478 PAD.n1477 0.0380882
R43049 PAD.n1477 PAD.n1476 0.0380882
R43050 PAD.n1476 PAD.n1194 0.0380882
R43051 PAD.n1469 PAD.n1194 0.0380882
R43052 PAD.n1469 PAD.n1468 0.0380882
R43053 PAD.n1468 PAD.n1467 0.0380882
R43054 PAD.n1467 PAD.n1199 0.0380882
R43055 PAD.n1460 PAD.n1199 0.0380882
R43056 PAD.n1460 PAD.n1459 0.0380882
R43057 PAD.n1459 PAD.n1458 0.0380882
R43058 PAD.n1458 PAD.n1204 0.0380882
R43059 PAD.n1451 PAD.n1204 0.0380882
R43060 PAD.n1451 PAD.n1450 0.0380882
R43061 PAD.n1450 PAD.n1449 0.0380882
R43062 PAD.n1449 PAD.n1209 0.0380882
R43063 PAD.n1442 PAD.n1209 0.0380882
R43064 PAD.n1442 PAD.n1441 0.0380882
R43065 PAD.n1441 PAD.n1440 0.0380882
R43066 PAD.n1440 PAD.n1214 0.0380882
R43067 PAD.n1433 PAD.n1214 0.0380882
R43068 PAD.n1433 PAD.n1432 0.0380882
R43069 PAD.n1432 PAD.n1431 0.0380882
R43070 PAD.n1431 PAD.n1219 0.0380882
R43071 PAD.n1424 PAD.n1219 0.0380882
R43072 PAD.n1424 PAD.n1423 0.0380882
R43073 PAD.n1423 PAD.n1422 0.0380882
R43074 PAD.n1422 PAD.n1224 0.0380882
R43075 PAD.n1415 PAD.n1224 0.0380882
R43076 PAD.n1415 PAD.n1414 0.0380882
R43077 PAD.n1414 PAD.n1413 0.0380882
R43078 PAD.n1413 PAD.n1229 0.0380882
R43079 PAD.n1406 PAD.n1229 0.0380882
R43080 PAD.n1406 PAD.n1405 0.0380882
R43081 PAD.n1405 PAD.n1404 0.0380882
R43082 PAD.n1404 PAD.n1234 0.0380882
R43083 PAD.n1397 PAD.n1234 0.0380882
R43084 PAD.n1397 PAD.n1396 0.0380882
R43085 PAD.n1396 PAD.n1395 0.0380882
R43086 PAD.n1395 PAD.n1239 0.0380882
R43087 PAD.n1388 PAD.n1239 0.0380882
R43088 PAD.n1388 PAD.n1387 0.0380882
R43089 PAD.n1387 PAD.n1386 0.0380882
R43090 PAD.n1386 PAD.n1244 0.0380882
R43091 PAD.n1379 PAD.n1244 0.0380882
R43092 PAD.n1379 PAD.n1378 0.0380882
R43093 PAD.n1378 PAD.n1377 0.0380882
R43094 PAD.n1377 PAD.n1249 0.0380882
R43095 PAD.n1370 PAD.n1249 0.0380882
R43096 PAD.n1370 PAD.n1369 0.0380882
R43097 PAD.n1369 PAD.n1368 0.0380882
R43098 PAD.n1368 PAD.n1254 0.0380882
R43099 PAD.n1361 PAD.n1254 0.0380882
R43100 PAD.n1361 PAD.n1360 0.0380882
R43101 PAD.n1360 PAD.n1359 0.0380882
R43102 PAD.n1359 PAD.n1259 0.0380882
R43103 PAD.n1352 PAD.n1259 0.0380882
R43104 PAD.n1352 PAD.n1351 0.0380882
R43105 PAD.n1351 PAD.n1350 0.0380882
R43106 PAD.n1350 PAD.n1264 0.0380882
R43107 PAD.n1343 PAD.n1264 0.0380882
R43108 PAD.n1343 PAD.n1342 0.0380882
R43109 PAD.n1342 PAD.n1341 0.0380882
R43110 PAD.n1341 PAD.n1269 0.0380882
R43111 PAD.n1334 PAD.n1269 0.0380882
R43112 PAD.n1334 PAD.n1333 0.0380882
R43113 PAD.n1333 PAD.n1332 0.0380882
R43114 PAD.n1332 PAD.n1274 0.0380882
R43115 PAD.n1325 PAD.n1274 0.0380882
R43116 PAD.n1325 PAD.n1324 0.0380882
R43117 PAD.n1324 PAD.n1323 0.0380882
R43118 PAD.n1323 PAD.n1279 0.0380882
R43119 PAD.n1316 PAD.n1279 0.0380882
R43120 PAD.n1316 PAD.n1315 0.0380882
R43121 PAD.n1315 PAD.n1314 0.0380882
R43122 PAD.n1314 PAD.n1284 0.0380882
R43123 PAD.n1307 PAD.n1284 0.0380882
R43124 PAD.n1307 PAD.n1306 0.0380882
R43125 PAD.n1306 PAD.n1305 0.0380882
R43126 PAD.n1305 PAD.n1289 0.0380882
R43127 PAD.n1298 PAD.n1289 0.0380882
R43128 PAD.n1298 PAD.n1297 0.0380882
R43129 PAD.n1297 PAD.n1296 0.0380882
R43130 PAD.n9749 PAD.n1579 0.0380882
R43131 PAD.n9753 PAD.n1579 0.0380882
R43132 PAD.n9757 PAD.n9753 0.0380882
R43133 PAD.n9761 PAD.n9757 0.0380882
R43134 PAD.n9761 PAD.n1575 0.0380882
R43135 PAD.n9765 PAD.n1575 0.0380882
R43136 PAD.n9769 PAD.n9765 0.0380882
R43137 PAD.n9773 PAD.n9769 0.0380882
R43138 PAD.n9773 PAD.n1573 0.0380882
R43139 PAD.n9777 PAD.n1573 0.0380882
R43140 PAD.n9781 PAD.n9777 0.0380882
R43141 PAD.n9785 PAD.n9781 0.0380882
R43142 PAD.n9785 PAD.n1571 0.0380882
R43143 PAD.n9789 PAD.n1571 0.0380882
R43144 PAD.n9793 PAD.n9789 0.0380882
R43145 PAD.n9797 PAD.n9793 0.0380882
R43146 PAD.n9797 PAD.n1569 0.0380882
R43147 PAD.n9801 PAD.n1569 0.0380882
R43148 PAD.n9805 PAD.n9801 0.0380882
R43149 PAD.n9809 PAD.n9805 0.0380882
R43150 PAD.n9809 PAD.n1567 0.0380882
R43151 PAD.n9813 PAD.n1567 0.0380882
R43152 PAD.n9817 PAD.n9813 0.0380882
R43153 PAD.n9821 PAD.n9817 0.0380882
R43154 PAD.n9821 PAD.n1565 0.0380882
R43155 PAD.n9825 PAD.n1565 0.0380882
R43156 PAD.n9829 PAD.n9825 0.0380882
R43157 PAD.n9833 PAD.n9829 0.0380882
R43158 PAD.n9833 PAD.n1563 0.0380882
R43159 PAD.n9837 PAD.n1563 0.0380882
R43160 PAD.n9841 PAD.n9837 0.0380882
R43161 PAD.n9845 PAD.n9841 0.0380882
R43162 PAD.n9845 PAD.n1561 0.0380882
R43163 PAD.n9849 PAD.n1561 0.0380882
R43164 PAD.n9853 PAD.n9849 0.0380882
R43165 PAD.n9857 PAD.n9853 0.0380882
R43166 PAD.n9857 PAD.n1559 0.0380882
R43167 PAD.n9861 PAD.n1559 0.0380882
R43168 PAD.n9865 PAD.n9861 0.0380882
R43169 PAD.n9869 PAD.n9865 0.0380882
R43170 PAD.n9869 PAD.n1557 0.0380882
R43171 PAD.n9873 PAD.n1557 0.0380882
R43172 PAD.n9877 PAD.n9873 0.0380882
R43173 PAD.n9881 PAD.n9877 0.0380882
R43174 PAD.n9881 PAD.n1555 0.0380882
R43175 PAD.n9885 PAD.n1555 0.0380882
R43176 PAD.n9889 PAD.n9885 0.0380882
R43177 PAD.n9893 PAD.n9889 0.0380882
R43178 PAD.n9893 PAD.n1553 0.0380882
R43179 PAD.n9897 PAD.n1553 0.0380882
R43180 PAD.n9901 PAD.n9897 0.0380882
R43181 PAD.n9905 PAD.n9901 0.0380882
R43182 PAD.n9905 PAD.n1551 0.0380882
R43183 PAD.n9909 PAD.n1551 0.0380882
R43184 PAD.n9913 PAD.n9909 0.0380882
R43185 PAD.n9917 PAD.n9913 0.0380882
R43186 PAD.n9917 PAD.n1549 0.0380882
R43187 PAD.n9921 PAD.n1549 0.0380882
R43188 PAD.n9925 PAD.n9921 0.0380882
R43189 PAD.n9929 PAD.n9925 0.0380882
R43190 PAD.n9929 PAD.n1547 0.0380882
R43191 PAD.n9933 PAD.n1547 0.0380882
R43192 PAD.n9937 PAD.n9933 0.0380882
R43193 PAD.n9941 PAD.n9937 0.0380882
R43194 PAD.n9941 PAD.n1545 0.0380882
R43195 PAD.n9945 PAD.n1545 0.0380882
R43196 PAD.n9949 PAD.n9945 0.0380882
R43197 PAD.n9953 PAD.n9949 0.0380882
R43198 PAD.n9953 PAD.n1543 0.0380882
R43199 PAD.n9957 PAD.n1543 0.0380882
R43200 PAD.n9961 PAD.n9957 0.0380882
R43201 PAD.n9965 PAD.n9961 0.0380882
R43202 PAD.n9965 PAD.n1541 0.0380882
R43203 PAD.n9969 PAD.n1541 0.0380882
R43204 PAD.n9973 PAD.n9969 0.0380882
R43205 PAD.n9977 PAD.n9973 0.0380882
R43206 PAD.n9977 PAD.n1539 0.0380882
R43207 PAD.n9981 PAD.n1539 0.0380882
R43208 PAD.n9985 PAD.n9981 0.0380882
R43209 PAD.n9989 PAD.n9985 0.0380882
R43210 PAD.n9989 PAD.n1537 0.0380882
R43211 PAD.n9994 PAD.n1537 0.0380882
R43212 PAD.n9994 PAD.n1535 0.0380882
R43213 PAD.n9751 PAD.n9750 0.0380882
R43214 PAD.n9752 PAD.n9751 0.0380882
R43215 PAD.n9752 PAD.n1576 0.0380882
R43216 PAD.n9762 PAD.n1576 0.0380882
R43217 PAD.n9763 PAD.n9762 0.0380882
R43218 PAD.n9764 PAD.n9763 0.0380882
R43219 PAD.n9764 PAD.n1574 0.0380882
R43220 PAD.n9774 PAD.n1574 0.0380882
R43221 PAD.n9775 PAD.n9774 0.0380882
R43222 PAD.n9776 PAD.n9775 0.0380882
R43223 PAD.n9776 PAD.n1572 0.0380882
R43224 PAD.n9786 PAD.n1572 0.0380882
R43225 PAD.n9787 PAD.n9786 0.0380882
R43226 PAD.n9788 PAD.n9787 0.0380882
R43227 PAD.n9788 PAD.n1570 0.0380882
R43228 PAD.n9798 PAD.n1570 0.0380882
R43229 PAD.n9799 PAD.n9798 0.0380882
R43230 PAD.n9800 PAD.n9799 0.0380882
R43231 PAD.n9800 PAD.n1568 0.0380882
R43232 PAD.n9810 PAD.n1568 0.0380882
R43233 PAD.n9811 PAD.n9810 0.0380882
R43234 PAD.n9812 PAD.n9811 0.0380882
R43235 PAD.n9812 PAD.n1566 0.0380882
R43236 PAD.n9822 PAD.n1566 0.0380882
R43237 PAD.n9823 PAD.n9822 0.0380882
R43238 PAD.n9824 PAD.n9823 0.0380882
R43239 PAD.n9824 PAD.n1564 0.0380882
R43240 PAD.n9834 PAD.n1564 0.0380882
R43241 PAD.n9835 PAD.n9834 0.0380882
R43242 PAD.n9836 PAD.n9835 0.0380882
R43243 PAD.n9836 PAD.n1562 0.0380882
R43244 PAD.n9846 PAD.n1562 0.0380882
R43245 PAD.n9847 PAD.n9846 0.0380882
R43246 PAD.n9848 PAD.n9847 0.0380882
R43247 PAD.n9848 PAD.n1560 0.0380882
R43248 PAD.n9858 PAD.n1560 0.0380882
R43249 PAD.n9859 PAD.n9858 0.0380882
R43250 PAD.n9860 PAD.n9859 0.0380882
R43251 PAD.n9860 PAD.n1558 0.0380882
R43252 PAD.n9870 PAD.n1558 0.0380882
R43253 PAD.n9871 PAD.n9870 0.0380882
R43254 PAD.n9872 PAD.n9871 0.0380882
R43255 PAD.n9872 PAD.n1556 0.0380882
R43256 PAD.n9882 PAD.n1556 0.0380882
R43257 PAD.n9883 PAD.n9882 0.0380882
R43258 PAD.n9884 PAD.n9883 0.0380882
R43259 PAD.n9884 PAD.n1554 0.0380882
R43260 PAD.n9894 PAD.n1554 0.0380882
R43261 PAD.n9895 PAD.n9894 0.0380882
R43262 PAD.n9896 PAD.n9895 0.0380882
R43263 PAD.n9896 PAD.n1552 0.0380882
R43264 PAD.n9906 PAD.n1552 0.0380882
R43265 PAD.n9907 PAD.n9906 0.0380882
R43266 PAD.n9908 PAD.n9907 0.0380882
R43267 PAD.n9908 PAD.n1550 0.0380882
R43268 PAD.n9918 PAD.n1550 0.0380882
R43269 PAD.n9919 PAD.n9918 0.0380882
R43270 PAD.n9920 PAD.n9919 0.0380882
R43271 PAD.n9920 PAD.n1548 0.0380882
R43272 PAD.n9930 PAD.n1548 0.0380882
R43273 PAD.n9931 PAD.n9930 0.0380882
R43274 PAD.n9932 PAD.n9931 0.0380882
R43275 PAD.n9932 PAD.n1546 0.0380882
R43276 PAD.n9942 PAD.n1546 0.0380882
R43277 PAD.n9943 PAD.n9942 0.0380882
R43278 PAD.n9944 PAD.n9943 0.0380882
R43279 PAD.n9944 PAD.n1544 0.0380882
R43280 PAD.n9954 PAD.n1544 0.0380882
R43281 PAD.n9955 PAD.n9954 0.0380882
R43282 PAD.n9956 PAD.n9955 0.0380882
R43283 PAD.n9956 PAD.n1542 0.0380882
R43284 PAD.n9966 PAD.n1542 0.0380882
R43285 PAD.n9967 PAD.n9966 0.0380882
R43286 PAD.n9968 PAD.n9967 0.0380882
R43287 PAD.n9968 PAD.n1540 0.0380882
R43288 PAD.n9978 PAD.n1540 0.0380882
R43289 PAD.n9979 PAD.n9978 0.0380882
R43290 PAD.n9980 PAD.n9979 0.0380882
R43291 PAD.n9980 PAD.n1538 0.0380882
R43292 PAD.n9990 PAD.n1538 0.0380882
R43293 PAD.n9991 PAD.n9990 0.0380882
R43294 PAD.n9993 PAD.n9991 0.0380882
R43295 PAD.n9993 PAD.n9992 0.0380882
R43296 PAD.n1931 PAD.n1930 0.0380882
R43297 PAD.n1930 PAD.n1600 0.0380882
R43298 PAD.n1924 PAD.n1600 0.0380882
R43299 PAD.n1924 PAD.n1603 0.0380882
R43300 PAD.n1920 PAD.n1603 0.0380882
R43301 PAD.n1920 PAD.n1606 0.0380882
R43302 PAD.n1912 PAD.n1606 0.0380882
R43303 PAD.n1912 PAD.n1608 0.0380882
R43304 PAD.n1908 PAD.n1608 0.0380882
R43305 PAD.n1908 PAD.n1610 0.0380882
R43306 PAD.n1900 PAD.n1610 0.0380882
R43307 PAD.n1900 PAD.n1612 0.0380882
R43308 PAD.n1896 PAD.n1612 0.0380882
R43309 PAD.n1896 PAD.n1614 0.0380882
R43310 PAD.n1888 PAD.n1614 0.0380882
R43311 PAD.n1888 PAD.n1616 0.0380882
R43312 PAD.n1884 PAD.n1616 0.0380882
R43313 PAD.n1884 PAD.n1618 0.0380882
R43314 PAD.n1876 PAD.n1618 0.0380882
R43315 PAD.n1876 PAD.n1620 0.0380882
R43316 PAD.n1872 PAD.n1620 0.0380882
R43317 PAD.n1872 PAD.n1622 0.0380882
R43318 PAD.n1864 PAD.n1622 0.0380882
R43319 PAD.n1864 PAD.n1624 0.0380882
R43320 PAD.n1860 PAD.n1624 0.0380882
R43321 PAD.n1860 PAD.n1626 0.0380882
R43322 PAD.n1852 PAD.n1626 0.0380882
R43323 PAD.n1852 PAD.n1628 0.0380882
R43324 PAD.n1848 PAD.n1628 0.0380882
R43325 PAD.n1848 PAD.n1630 0.0380882
R43326 PAD.n1840 PAD.n1630 0.0380882
R43327 PAD.n1840 PAD.n1632 0.0380882
R43328 PAD.n1836 PAD.n1632 0.0380882
R43329 PAD.n1836 PAD.n1634 0.0380882
R43330 PAD.n1828 PAD.n1634 0.0380882
R43331 PAD.n1828 PAD.n1636 0.0380882
R43332 PAD.n1824 PAD.n1636 0.0380882
R43333 PAD.n1824 PAD.n1638 0.0380882
R43334 PAD.n1816 PAD.n1638 0.0380882
R43335 PAD.n1816 PAD.n1640 0.0380882
R43336 PAD.n1812 PAD.n1640 0.0380882
R43337 PAD.n1812 PAD.n1642 0.0380882
R43338 PAD.n1804 PAD.n1642 0.0380882
R43339 PAD.n1804 PAD.n1644 0.0380882
R43340 PAD.n1800 PAD.n1644 0.0380882
R43341 PAD.n1800 PAD.n1646 0.0380882
R43342 PAD.n1792 PAD.n1646 0.0380882
R43343 PAD.n1792 PAD.n1648 0.0380882
R43344 PAD.n1788 PAD.n1648 0.0380882
R43345 PAD.n1788 PAD.n1650 0.0380882
R43346 PAD.n1780 PAD.n1650 0.0380882
R43347 PAD.n1780 PAD.n1652 0.0380882
R43348 PAD.n1776 PAD.n1652 0.0380882
R43349 PAD.n1776 PAD.n1654 0.0380882
R43350 PAD.n1768 PAD.n1654 0.0380882
R43351 PAD.n1768 PAD.n1656 0.0380882
R43352 PAD.n1764 PAD.n1656 0.0380882
R43353 PAD.n1764 PAD.n1658 0.0380882
R43354 PAD.n1756 PAD.n1658 0.0380882
R43355 PAD.n1756 PAD.n1660 0.0380882
R43356 PAD.n1752 PAD.n1660 0.0380882
R43357 PAD.n1752 PAD.n1662 0.0380882
R43358 PAD.n1744 PAD.n1662 0.0380882
R43359 PAD.n1744 PAD.n1664 0.0380882
R43360 PAD.n1740 PAD.n1664 0.0380882
R43361 PAD.n1740 PAD.n1666 0.0380882
R43362 PAD.n1732 PAD.n1666 0.0380882
R43363 PAD.n1732 PAD.n1668 0.0380882
R43364 PAD.n1728 PAD.n1668 0.0380882
R43365 PAD.n1728 PAD.n1670 0.0380882
R43366 PAD.n1720 PAD.n1670 0.0380882
R43367 PAD.n1720 PAD.n1672 0.0380882
R43368 PAD.n1716 PAD.n1672 0.0380882
R43369 PAD.n1716 PAD.n1674 0.0380882
R43370 PAD.n1708 PAD.n1674 0.0380882
R43371 PAD.n1708 PAD.n1676 0.0380882
R43372 PAD.n1704 PAD.n1676 0.0380882
R43373 PAD.n1704 PAD.n1678 0.0380882
R43374 PAD.n1696 PAD.n1678 0.0380882
R43375 PAD.n1696 PAD.n1680 0.0380882
R43376 PAD.n1692 PAD.n1680 0.0380882
R43377 PAD.n1692 PAD.n1682 0.0380882
R43378 PAD.n1684 PAD.n1682 0.0380882
R43379 PAD.n1932 PAD.n1598 0.0380882
R43380 PAD.n1604 PAD.n1598 0.0380882
R43381 PAD.n1923 PAD.n1604 0.0380882
R43382 PAD.n1923 PAD.n1922 0.0380882
R43383 PAD.n1922 PAD.n1921 0.0380882
R43384 PAD.n1921 PAD.n1605 0.0380882
R43385 PAD.n1911 PAD.n1605 0.0380882
R43386 PAD.n1911 PAD.n1910 0.0380882
R43387 PAD.n1910 PAD.n1909 0.0380882
R43388 PAD.n1909 PAD.n1609 0.0380882
R43389 PAD.n1899 PAD.n1609 0.0380882
R43390 PAD.n1899 PAD.n1898 0.0380882
R43391 PAD.n1898 PAD.n1897 0.0380882
R43392 PAD.n1897 PAD.n1613 0.0380882
R43393 PAD.n1887 PAD.n1613 0.0380882
R43394 PAD.n1887 PAD.n1886 0.0380882
R43395 PAD.n1886 PAD.n1885 0.0380882
R43396 PAD.n1885 PAD.n1617 0.0380882
R43397 PAD.n1875 PAD.n1617 0.0380882
R43398 PAD.n1875 PAD.n1874 0.0380882
R43399 PAD.n1874 PAD.n1873 0.0380882
R43400 PAD.n1873 PAD.n1621 0.0380882
R43401 PAD.n1863 PAD.n1621 0.0380882
R43402 PAD.n1863 PAD.n1862 0.0380882
R43403 PAD.n1862 PAD.n1861 0.0380882
R43404 PAD.n1861 PAD.n1625 0.0380882
R43405 PAD.n1851 PAD.n1625 0.0380882
R43406 PAD.n1851 PAD.n1850 0.0380882
R43407 PAD.n1850 PAD.n1849 0.0380882
R43408 PAD.n1849 PAD.n1629 0.0380882
R43409 PAD.n1839 PAD.n1629 0.0380882
R43410 PAD.n1839 PAD.n1838 0.0380882
R43411 PAD.n1838 PAD.n1837 0.0380882
R43412 PAD.n1837 PAD.n1633 0.0380882
R43413 PAD.n1827 PAD.n1633 0.0380882
R43414 PAD.n1827 PAD.n1826 0.0380882
R43415 PAD.n1826 PAD.n1825 0.0380882
R43416 PAD.n1825 PAD.n1637 0.0380882
R43417 PAD.n1815 PAD.n1637 0.0380882
R43418 PAD.n1815 PAD.n1814 0.0380882
R43419 PAD.n1814 PAD.n1813 0.0380882
R43420 PAD.n1813 PAD.n1641 0.0380882
R43421 PAD.n1803 PAD.n1641 0.0380882
R43422 PAD.n1803 PAD.n1802 0.0380882
R43423 PAD.n1802 PAD.n1801 0.0380882
R43424 PAD.n1801 PAD.n1645 0.0380882
R43425 PAD.n1791 PAD.n1645 0.0380882
R43426 PAD.n1791 PAD.n1790 0.0380882
R43427 PAD.n1790 PAD.n1789 0.0380882
R43428 PAD.n1789 PAD.n1649 0.0380882
R43429 PAD.n1779 PAD.n1649 0.0380882
R43430 PAD.n1779 PAD.n1778 0.0380882
R43431 PAD.n1778 PAD.n1777 0.0380882
R43432 PAD.n1777 PAD.n1653 0.0380882
R43433 PAD.n1767 PAD.n1653 0.0380882
R43434 PAD.n1767 PAD.n1766 0.0380882
R43435 PAD.n1766 PAD.n1765 0.0380882
R43436 PAD.n1765 PAD.n1657 0.0380882
R43437 PAD.n1755 PAD.n1657 0.0380882
R43438 PAD.n1755 PAD.n1754 0.0380882
R43439 PAD.n1754 PAD.n1753 0.0380882
R43440 PAD.n1753 PAD.n1661 0.0380882
R43441 PAD.n1743 PAD.n1661 0.0380882
R43442 PAD.n1743 PAD.n1742 0.0380882
R43443 PAD.n1742 PAD.n1741 0.0380882
R43444 PAD.n1741 PAD.n1665 0.0380882
R43445 PAD.n1731 PAD.n1665 0.0380882
R43446 PAD.n1731 PAD.n1730 0.0380882
R43447 PAD.n1730 PAD.n1729 0.0380882
R43448 PAD.n1729 PAD.n1669 0.0380882
R43449 PAD.n1719 PAD.n1669 0.0380882
R43450 PAD.n1719 PAD.n1718 0.0380882
R43451 PAD.n1718 PAD.n1717 0.0380882
R43452 PAD.n1717 PAD.n1673 0.0380882
R43453 PAD.n1707 PAD.n1673 0.0380882
R43454 PAD.n1707 PAD.n1706 0.0380882
R43455 PAD.n1706 PAD.n1705 0.0380882
R43456 PAD.n1705 PAD.n1677 0.0380882
R43457 PAD.n1695 PAD.n1677 0.0380882
R43458 PAD.n1695 PAD.n1694 0.0380882
R43459 PAD.n1694 PAD.n1693 0.0380882
R43460 PAD.n1693 PAD.n1681 0.0380882
R43461 PAD.n1683 PAD.n1681 0.0380882
R43462 PAD.n9463 PAD.n2031 0.0380882
R43463 PAD.n9467 PAD.n2031 0.0380882
R43464 PAD.n9471 PAD.n9467 0.0380882
R43465 PAD.n9475 PAD.n9471 0.0380882
R43466 PAD.n9475 PAD.n2027 0.0380882
R43467 PAD.n9479 PAD.n2027 0.0380882
R43468 PAD.n9483 PAD.n9479 0.0380882
R43469 PAD.n9487 PAD.n9483 0.0380882
R43470 PAD.n9487 PAD.n2025 0.0380882
R43471 PAD.n9491 PAD.n2025 0.0380882
R43472 PAD.n9495 PAD.n9491 0.0380882
R43473 PAD.n9499 PAD.n9495 0.0380882
R43474 PAD.n9499 PAD.n2023 0.0380882
R43475 PAD.n9503 PAD.n2023 0.0380882
R43476 PAD.n9507 PAD.n9503 0.0380882
R43477 PAD.n9511 PAD.n9507 0.0380882
R43478 PAD.n9511 PAD.n2021 0.0380882
R43479 PAD.n9515 PAD.n2021 0.0380882
R43480 PAD.n9519 PAD.n9515 0.0380882
R43481 PAD.n9523 PAD.n9519 0.0380882
R43482 PAD.n9523 PAD.n2019 0.0380882
R43483 PAD.n9527 PAD.n2019 0.0380882
R43484 PAD.n9531 PAD.n9527 0.0380882
R43485 PAD.n9535 PAD.n9531 0.0380882
R43486 PAD.n9535 PAD.n2017 0.0380882
R43487 PAD.n9539 PAD.n2017 0.0380882
R43488 PAD.n9543 PAD.n9539 0.0380882
R43489 PAD.n9547 PAD.n9543 0.0380882
R43490 PAD.n9547 PAD.n2015 0.0380882
R43491 PAD.n9551 PAD.n2015 0.0380882
R43492 PAD.n9555 PAD.n9551 0.0380882
R43493 PAD.n9559 PAD.n9555 0.0380882
R43494 PAD.n9559 PAD.n2013 0.0380882
R43495 PAD.n9563 PAD.n2013 0.0380882
R43496 PAD.n9567 PAD.n9563 0.0380882
R43497 PAD.n9571 PAD.n9567 0.0380882
R43498 PAD.n9571 PAD.n2011 0.0380882
R43499 PAD.n9575 PAD.n2011 0.0380882
R43500 PAD.n9579 PAD.n9575 0.0380882
R43501 PAD.n9583 PAD.n9579 0.0380882
R43502 PAD.n9583 PAD.n2009 0.0380882
R43503 PAD.n9587 PAD.n2009 0.0380882
R43504 PAD.n9591 PAD.n9587 0.0380882
R43505 PAD.n9595 PAD.n9591 0.0380882
R43506 PAD.n9595 PAD.n2007 0.0380882
R43507 PAD.n9599 PAD.n2007 0.0380882
R43508 PAD.n9603 PAD.n9599 0.0380882
R43509 PAD.n9607 PAD.n9603 0.0380882
R43510 PAD.n9607 PAD.n2005 0.0380882
R43511 PAD.n9611 PAD.n2005 0.0380882
R43512 PAD.n9615 PAD.n9611 0.0380882
R43513 PAD.n9619 PAD.n9615 0.0380882
R43514 PAD.n9619 PAD.n2003 0.0380882
R43515 PAD.n9623 PAD.n2003 0.0380882
R43516 PAD.n9627 PAD.n9623 0.0380882
R43517 PAD.n9631 PAD.n9627 0.0380882
R43518 PAD.n9631 PAD.n2001 0.0380882
R43519 PAD.n9635 PAD.n2001 0.0380882
R43520 PAD.n9639 PAD.n9635 0.0380882
R43521 PAD.n9643 PAD.n9639 0.0380882
R43522 PAD.n9643 PAD.n1999 0.0380882
R43523 PAD.n9647 PAD.n1999 0.0380882
R43524 PAD.n9651 PAD.n9647 0.0380882
R43525 PAD.n9655 PAD.n9651 0.0380882
R43526 PAD.n9655 PAD.n1997 0.0380882
R43527 PAD.n9659 PAD.n1997 0.0380882
R43528 PAD.n9663 PAD.n9659 0.0380882
R43529 PAD.n9667 PAD.n9663 0.0380882
R43530 PAD.n9667 PAD.n1995 0.0380882
R43531 PAD.n9671 PAD.n1995 0.0380882
R43532 PAD.n9675 PAD.n9671 0.0380882
R43533 PAD.n9679 PAD.n9675 0.0380882
R43534 PAD.n9679 PAD.n1993 0.0380882
R43535 PAD.n9683 PAD.n1993 0.0380882
R43536 PAD.n9687 PAD.n9683 0.0380882
R43537 PAD.n9691 PAD.n9687 0.0380882
R43538 PAD.n9691 PAD.n1991 0.0380882
R43539 PAD.n9695 PAD.n1991 0.0380882
R43540 PAD.n9699 PAD.n9695 0.0380882
R43541 PAD.n9703 PAD.n9699 0.0380882
R43542 PAD.n9703 PAD.n1989 0.0380882
R43543 PAD.n9708 PAD.n1989 0.0380882
R43544 PAD.n9708 PAD.n1987 0.0380882
R43545 PAD.n9465 PAD.n9464 0.0380882
R43546 PAD.n9466 PAD.n9465 0.0380882
R43547 PAD.n9466 PAD.n2028 0.0380882
R43548 PAD.n9476 PAD.n2028 0.0380882
R43549 PAD.n9477 PAD.n9476 0.0380882
R43550 PAD.n9478 PAD.n9477 0.0380882
R43551 PAD.n9478 PAD.n2026 0.0380882
R43552 PAD.n9488 PAD.n2026 0.0380882
R43553 PAD.n9489 PAD.n9488 0.0380882
R43554 PAD.n9490 PAD.n9489 0.0380882
R43555 PAD.n9490 PAD.n2024 0.0380882
R43556 PAD.n9500 PAD.n2024 0.0380882
R43557 PAD.n9501 PAD.n9500 0.0380882
R43558 PAD.n9502 PAD.n9501 0.0380882
R43559 PAD.n9502 PAD.n2022 0.0380882
R43560 PAD.n9512 PAD.n2022 0.0380882
R43561 PAD.n9513 PAD.n9512 0.0380882
R43562 PAD.n9514 PAD.n9513 0.0380882
R43563 PAD.n9514 PAD.n2020 0.0380882
R43564 PAD.n9524 PAD.n2020 0.0380882
R43565 PAD.n9525 PAD.n9524 0.0380882
R43566 PAD.n9526 PAD.n9525 0.0380882
R43567 PAD.n9526 PAD.n2018 0.0380882
R43568 PAD.n9536 PAD.n2018 0.0380882
R43569 PAD.n9537 PAD.n9536 0.0380882
R43570 PAD.n9538 PAD.n9537 0.0380882
R43571 PAD.n9538 PAD.n2016 0.0380882
R43572 PAD.n9548 PAD.n2016 0.0380882
R43573 PAD.n9549 PAD.n9548 0.0380882
R43574 PAD.n9550 PAD.n9549 0.0380882
R43575 PAD.n9550 PAD.n2014 0.0380882
R43576 PAD.n9560 PAD.n2014 0.0380882
R43577 PAD.n9561 PAD.n9560 0.0380882
R43578 PAD.n9562 PAD.n9561 0.0380882
R43579 PAD.n9562 PAD.n2012 0.0380882
R43580 PAD.n9572 PAD.n2012 0.0380882
R43581 PAD.n9573 PAD.n9572 0.0380882
R43582 PAD.n9574 PAD.n9573 0.0380882
R43583 PAD.n9574 PAD.n2010 0.0380882
R43584 PAD.n9584 PAD.n2010 0.0380882
R43585 PAD.n9585 PAD.n9584 0.0380882
R43586 PAD.n9586 PAD.n9585 0.0380882
R43587 PAD.n9586 PAD.n2008 0.0380882
R43588 PAD.n9596 PAD.n2008 0.0380882
R43589 PAD.n9597 PAD.n9596 0.0380882
R43590 PAD.n9598 PAD.n9597 0.0380882
R43591 PAD.n9598 PAD.n2006 0.0380882
R43592 PAD.n9608 PAD.n2006 0.0380882
R43593 PAD.n9609 PAD.n9608 0.0380882
R43594 PAD.n9610 PAD.n9609 0.0380882
R43595 PAD.n9610 PAD.n2004 0.0380882
R43596 PAD.n9620 PAD.n2004 0.0380882
R43597 PAD.n9621 PAD.n9620 0.0380882
R43598 PAD.n9622 PAD.n9621 0.0380882
R43599 PAD.n9622 PAD.n2002 0.0380882
R43600 PAD.n9632 PAD.n2002 0.0380882
R43601 PAD.n9633 PAD.n9632 0.0380882
R43602 PAD.n9634 PAD.n9633 0.0380882
R43603 PAD.n9634 PAD.n2000 0.0380882
R43604 PAD.n9644 PAD.n2000 0.0380882
R43605 PAD.n9645 PAD.n9644 0.0380882
R43606 PAD.n9646 PAD.n9645 0.0380882
R43607 PAD.n9646 PAD.n1998 0.0380882
R43608 PAD.n9656 PAD.n1998 0.0380882
R43609 PAD.n9657 PAD.n9656 0.0380882
R43610 PAD.n9658 PAD.n9657 0.0380882
R43611 PAD.n9658 PAD.n1996 0.0380882
R43612 PAD.n9668 PAD.n1996 0.0380882
R43613 PAD.n9669 PAD.n9668 0.0380882
R43614 PAD.n9670 PAD.n9669 0.0380882
R43615 PAD.n9670 PAD.n1994 0.0380882
R43616 PAD.n9680 PAD.n1994 0.0380882
R43617 PAD.n9681 PAD.n9680 0.0380882
R43618 PAD.n9682 PAD.n9681 0.0380882
R43619 PAD.n9682 PAD.n1992 0.0380882
R43620 PAD.n9692 PAD.n1992 0.0380882
R43621 PAD.n9693 PAD.n9692 0.0380882
R43622 PAD.n9694 PAD.n9693 0.0380882
R43623 PAD.n9694 PAD.n1990 0.0380882
R43624 PAD.n9704 PAD.n1990 0.0380882
R43625 PAD.n9705 PAD.n9704 0.0380882
R43626 PAD.n9707 PAD.n9705 0.0380882
R43627 PAD.n9707 PAD.n9706 0.0380882
R43628 PAD.n9197 PAD.n2134 0.0380882
R43629 PAD.n9201 PAD.n2134 0.0380882
R43630 PAD.n9205 PAD.n9201 0.0380882
R43631 PAD.n9209 PAD.n9205 0.0380882
R43632 PAD.n9209 PAD.n2130 0.0380882
R43633 PAD.n9213 PAD.n2130 0.0380882
R43634 PAD.n9217 PAD.n9213 0.0380882
R43635 PAD.n9221 PAD.n9217 0.0380882
R43636 PAD.n9221 PAD.n2128 0.0380882
R43637 PAD.n9225 PAD.n2128 0.0380882
R43638 PAD.n9229 PAD.n9225 0.0380882
R43639 PAD.n9233 PAD.n9229 0.0380882
R43640 PAD.n9233 PAD.n2126 0.0380882
R43641 PAD.n9237 PAD.n2126 0.0380882
R43642 PAD.n9241 PAD.n9237 0.0380882
R43643 PAD.n9245 PAD.n9241 0.0380882
R43644 PAD.n9245 PAD.n2124 0.0380882
R43645 PAD.n9249 PAD.n2124 0.0380882
R43646 PAD.n9253 PAD.n9249 0.0380882
R43647 PAD.n9257 PAD.n9253 0.0380882
R43648 PAD.n9257 PAD.n2122 0.0380882
R43649 PAD.n9261 PAD.n2122 0.0380882
R43650 PAD.n9265 PAD.n9261 0.0380882
R43651 PAD.n9269 PAD.n9265 0.0380882
R43652 PAD.n9269 PAD.n2120 0.0380882
R43653 PAD.n9273 PAD.n2120 0.0380882
R43654 PAD.n9277 PAD.n9273 0.0380882
R43655 PAD.n9281 PAD.n9277 0.0380882
R43656 PAD.n9281 PAD.n2118 0.0380882
R43657 PAD.n9285 PAD.n2118 0.0380882
R43658 PAD.n9289 PAD.n9285 0.0380882
R43659 PAD.n9293 PAD.n9289 0.0380882
R43660 PAD.n9293 PAD.n2116 0.0380882
R43661 PAD.n9297 PAD.n2116 0.0380882
R43662 PAD.n9301 PAD.n9297 0.0380882
R43663 PAD.n9305 PAD.n9301 0.0380882
R43664 PAD.n9305 PAD.n2114 0.0380882
R43665 PAD.n9309 PAD.n2114 0.0380882
R43666 PAD.n9313 PAD.n9309 0.0380882
R43667 PAD.n9317 PAD.n9313 0.0380882
R43668 PAD.n9317 PAD.n2112 0.0380882
R43669 PAD.n9321 PAD.n2112 0.0380882
R43670 PAD.n9325 PAD.n9321 0.0380882
R43671 PAD.n9329 PAD.n9325 0.0380882
R43672 PAD.n9329 PAD.n2110 0.0380882
R43673 PAD.n9333 PAD.n2110 0.0380882
R43674 PAD.n9337 PAD.n9333 0.0380882
R43675 PAD.n9341 PAD.n9337 0.0380882
R43676 PAD.n9341 PAD.n2108 0.0380882
R43677 PAD.n9345 PAD.n2108 0.0380882
R43678 PAD.n9349 PAD.n9345 0.0380882
R43679 PAD.n9353 PAD.n9349 0.0380882
R43680 PAD.n9353 PAD.n2106 0.0380882
R43681 PAD.n9357 PAD.n2106 0.0380882
R43682 PAD.n9361 PAD.n9357 0.0380882
R43683 PAD.n9365 PAD.n9361 0.0380882
R43684 PAD.n9365 PAD.n2104 0.0380882
R43685 PAD.n9369 PAD.n2104 0.0380882
R43686 PAD.n9373 PAD.n9369 0.0380882
R43687 PAD.n9377 PAD.n9373 0.0380882
R43688 PAD.n9377 PAD.n2102 0.0380882
R43689 PAD.n9381 PAD.n2102 0.0380882
R43690 PAD.n9385 PAD.n9381 0.0380882
R43691 PAD.n9389 PAD.n9385 0.0380882
R43692 PAD.n9389 PAD.n2100 0.0380882
R43693 PAD.n9393 PAD.n2100 0.0380882
R43694 PAD.n9397 PAD.n9393 0.0380882
R43695 PAD.n9401 PAD.n9397 0.0380882
R43696 PAD.n9401 PAD.n2098 0.0380882
R43697 PAD.n9405 PAD.n2098 0.0380882
R43698 PAD.n9409 PAD.n9405 0.0380882
R43699 PAD.n9413 PAD.n9409 0.0380882
R43700 PAD.n9413 PAD.n2096 0.0380882
R43701 PAD.n9417 PAD.n2096 0.0380882
R43702 PAD.n9421 PAD.n9417 0.0380882
R43703 PAD.n9425 PAD.n9421 0.0380882
R43704 PAD.n9425 PAD.n2094 0.0380882
R43705 PAD.n9429 PAD.n2094 0.0380882
R43706 PAD.n9433 PAD.n9429 0.0380882
R43707 PAD.n9437 PAD.n9433 0.0380882
R43708 PAD.n9437 PAD.n2092 0.0380882
R43709 PAD.n9441 PAD.n2092 0.0380882
R43710 PAD.n9441 PAD.n2090 0.0380882
R43711 PAD.n9199 PAD.n9198 0.0380882
R43712 PAD.n9200 PAD.n9199 0.0380882
R43713 PAD.n9200 PAD.n2131 0.0380882
R43714 PAD.n9210 PAD.n2131 0.0380882
R43715 PAD.n9211 PAD.n9210 0.0380882
R43716 PAD.n9212 PAD.n9211 0.0380882
R43717 PAD.n9212 PAD.n2129 0.0380882
R43718 PAD.n9222 PAD.n2129 0.0380882
R43719 PAD.n9223 PAD.n9222 0.0380882
R43720 PAD.n9224 PAD.n9223 0.0380882
R43721 PAD.n9224 PAD.n2127 0.0380882
R43722 PAD.n9234 PAD.n2127 0.0380882
R43723 PAD.n9235 PAD.n9234 0.0380882
R43724 PAD.n9236 PAD.n9235 0.0380882
R43725 PAD.n9236 PAD.n2125 0.0380882
R43726 PAD.n9246 PAD.n2125 0.0380882
R43727 PAD.n9247 PAD.n9246 0.0380882
R43728 PAD.n9248 PAD.n9247 0.0380882
R43729 PAD.n9248 PAD.n2123 0.0380882
R43730 PAD.n9258 PAD.n2123 0.0380882
R43731 PAD.n9259 PAD.n9258 0.0380882
R43732 PAD.n9260 PAD.n9259 0.0380882
R43733 PAD.n9260 PAD.n2121 0.0380882
R43734 PAD.n9270 PAD.n2121 0.0380882
R43735 PAD.n9271 PAD.n9270 0.0380882
R43736 PAD.n9272 PAD.n9271 0.0380882
R43737 PAD.n9272 PAD.n2119 0.0380882
R43738 PAD.n9282 PAD.n2119 0.0380882
R43739 PAD.n9283 PAD.n9282 0.0380882
R43740 PAD.n9284 PAD.n9283 0.0380882
R43741 PAD.n9284 PAD.n2117 0.0380882
R43742 PAD.n9294 PAD.n2117 0.0380882
R43743 PAD.n9295 PAD.n9294 0.0380882
R43744 PAD.n9296 PAD.n9295 0.0380882
R43745 PAD.n9296 PAD.n2115 0.0380882
R43746 PAD.n9306 PAD.n2115 0.0380882
R43747 PAD.n9307 PAD.n9306 0.0380882
R43748 PAD.n9308 PAD.n9307 0.0380882
R43749 PAD.n9308 PAD.n2113 0.0380882
R43750 PAD.n9318 PAD.n2113 0.0380882
R43751 PAD.n9319 PAD.n9318 0.0380882
R43752 PAD.n9320 PAD.n9319 0.0380882
R43753 PAD.n9320 PAD.n2111 0.0380882
R43754 PAD.n9330 PAD.n2111 0.0380882
R43755 PAD.n9331 PAD.n9330 0.0380882
R43756 PAD.n9332 PAD.n9331 0.0380882
R43757 PAD.n9332 PAD.n2109 0.0380882
R43758 PAD.n9342 PAD.n2109 0.0380882
R43759 PAD.n9343 PAD.n9342 0.0380882
R43760 PAD.n9344 PAD.n9343 0.0380882
R43761 PAD.n9344 PAD.n2107 0.0380882
R43762 PAD.n9354 PAD.n2107 0.0380882
R43763 PAD.n9355 PAD.n9354 0.0380882
R43764 PAD.n9356 PAD.n9355 0.0380882
R43765 PAD.n9356 PAD.n2105 0.0380882
R43766 PAD.n9366 PAD.n2105 0.0380882
R43767 PAD.n9367 PAD.n9366 0.0380882
R43768 PAD.n9368 PAD.n9367 0.0380882
R43769 PAD.n9368 PAD.n2103 0.0380882
R43770 PAD.n9378 PAD.n2103 0.0380882
R43771 PAD.n9379 PAD.n9378 0.0380882
R43772 PAD.n9380 PAD.n9379 0.0380882
R43773 PAD.n9380 PAD.n2101 0.0380882
R43774 PAD.n9390 PAD.n2101 0.0380882
R43775 PAD.n9391 PAD.n9390 0.0380882
R43776 PAD.n9392 PAD.n9391 0.0380882
R43777 PAD.n9392 PAD.n2099 0.0380882
R43778 PAD.n9402 PAD.n2099 0.0380882
R43779 PAD.n9403 PAD.n9402 0.0380882
R43780 PAD.n9404 PAD.n9403 0.0380882
R43781 PAD.n9404 PAD.n2097 0.0380882
R43782 PAD.n9414 PAD.n2097 0.0380882
R43783 PAD.n9415 PAD.n9414 0.0380882
R43784 PAD.n9416 PAD.n9415 0.0380882
R43785 PAD.n9416 PAD.n2095 0.0380882
R43786 PAD.n9426 PAD.n2095 0.0380882
R43787 PAD.n9427 PAD.n9426 0.0380882
R43788 PAD.n9428 PAD.n9427 0.0380882
R43789 PAD.n9428 PAD.n2093 0.0380882
R43790 PAD.n9438 PAD.n2093 0.0380882
R43791 PAD.n9439 PAD.n9438 0.0380882
R43792 PAD.n9440 PAD.n9439 0.0380882
R43793 PAD.n9440 PAD.n2040 0.0380882
R43794 PAD.n2482 PAD.n2481 0.0380882
R43795 PAD.n2481 PAD.n2152 0.0380882
R43796 PAD.n2475 PAD.n2152 0.0380882
R43797 PAD.n2475 PAD.n2155 0.0380882
R43798 PAD.n2471 PAD.n2155 0.0380882
R43799 PAD.n2471 PAD.n2158 0.0380882
R43800 PAD.n2463 PAD.n2158 0.0380882
R43801 PAD.n2463 PAD.n2160 0.0380882
R43802 PAD.n2459 PAD.n2160 0.0380882
R43803 PAD.n2459 PAD.n2162 0.0380882
R43804 PAD.n2451 PAD.n2162 0.0380882
R43805 PAD.n2451 PAD.n2164 0.0380882
R43806 PAD.n2447 PAD.n2164 0.0380882
R43807 PAD.n2447 PAD.n2166 0.0380882
R43808 PAD.n2439 PAD.n2166 0.0380882
R43809 PAD.n2439 PAD.n2168 0.0380882
R43810 PAD.n2435 PAD.n2168 0.0380882
R43811 PAD.n2435 PAD.n2170 0.0380882
R43812 PAD.n2427 PAD.n2170 0.0380882
R43813 PAD.n2427 PAD.n2172 0.0380882
R43814 PAD.n2423 PAD.n2172 0.0380882
R43815 PAD.n2423 PAD.n2174 0.0380882
R43816 PAD.n2415 PAD.n2174 0.0380882
R43817 PAD.n2415 PAD.n2176 0.0380882
R43818 PAD.n2411 PAD.n2176 0.0380882
R43819 PAD.n2411 PAD.n2178 0.0380882
R43820 PAD.n2403 PAD.n2178 0.0380882
R43821 PAD.n2403 PAD.n2180 0.0380882
R43822 PAD.n2399 PAD.n2180 0.0380882
R43823 PAD.n2399 PAD.n2182 0.0380882
R43824 PAD.n2391 PAD.n2182 0.0380882
R43825 PAD.n2391 PAD.n2184 0.0380882
R43826 PAD.n2387 PAD.n2184 0.0380882
R43827 PAD.n2387 PAD.n2186 0.0380882
R43828 PAD.n2379 PAD.n2186 0.0380882
R43829 PAD.n2379 PAD.n2188 0.0380882
R43830 PAD.n2375 PAD.n2188 0.0380882
R43831 PAD.n2375 PAD.n2190 0.0380882
R43832 PAD.n2367 PAD.n2190 0.0380882
R43833 PAD.n2367 PAD.n2192 0.0380882
R43834 PAD.n2363 PAD.n2192 0.0380882
R43835 PAD.n2363 PAD.n2194 0.0380882
R43836 PAD.n2355 PAD.n2194 0.0380882
R43837 PAD.n2355 PAD.n2196 0.0380882
R43838 PAD.n2351 PAD.n2196 0.0380882
R43839 PAD.n2351 PAD.n2198 0.0380882
R43840 PAD.n2343 PAD.n2198 0.0380882
R43841 PAD.n2343 PAD.n2200 0.0380882
R43842 PAD.n2339 PAD.n2200 0.0380882
R43843 PAD.n2339 PAD.n2202 0.0380882
R43844 PAD.n2331 PAD.n2202 0.0380882
R43845 PAD.n2331 PAD.n2204 0.0380882
R43846 PAD.n2327 PAD.n2204 0.0380882
R43847 PAD.n2327 PAD.n2206 0.0380882
R43848 PAD.n2319 PAD.n2206 0.0380882
R43849 PAD.n2319 PAD.n2208 0.0380882
R43850 PAD.n2315 PAD.n2208 0.0380882
R43851 PAD.n2315 PAD.n2210 0.0380882
R43852 PAD.n2307 PAD.n2210 0.0380882
R43853 PAD.n2307 PAD.n2212 0.0380882
R43854 PAD.n2303 PAD.n2212 0.0380882
R43855 PAD.n2303 PAD.n2214 0.0380882
R43856 PAD.n2295 PAD.n2214 0.0380882
R43857 PAD.n2295 PAD.n2216 0.0380882
R43858 PAD.n2291 PAD.n2216 0.0380882
R43859 PAD.n2291 PAD.n2218 0.0380882
R43860 PAD.n2283 PAD.n2218 0.0380882
R43861 PAD.n2283 PAD.n2220 0.0380882
R43862 PAD.n2279 PAD.n2220 0.0380882
R43863 PAD.n2279 PAD.n2222 0.0380882
R43864 PAD.n2271 PAD.n2222 0.0380882
R43865 PAD.n2271 PAD.n2224 0.0380882
R43866 PAD.n2267 PAD.n2224 0.0380882
R43867 PAD.n2267 PAD.n2226 0.0380882
R43868 PAD.n2259 PAD.n2226 0.0380882
R43869 PAD.n2259 PAD.n2228 0.0380882
R43870 PAD.n2255 PAD.n2228 0.0380882
R43871 PAD.n2255 PAD.n2230 0.0380882
R43872 PAD.n2247 PAD.n2230 0.0380882
R43873 PAD.n2247 PAD.n2232 0.0380882
R43874 PAD.n2243 PAD.n2232 0.0380882
R43875 PAD.n2243 PAD.n2234 0.0380882
R43876 PAD.n2235 PAD.n2234 0.0380882
R43877 PAD.n2483 PAD.n2150 0.0380882
R43878 PAD.n2156 PAD.n2150 0.0380882
R43879 PAD.n2474 PAD.n2156 0.0380882
R43880 PAD.n2474 PAD.n2473 0.0380882
R43881 PAD.n2473 PAD.n2472 0.0380882
R43882 PAD.n2472 PAD.n2157 0.0380882
R43883 PAD.n2462 PAD.n2157 0.0380882
R43884 PAD.n2462 PAD.n2461 0.0380882
R43885 PAD.n2461 PAD.n2460 0.0380882
R43886 PAD.n2460 PAD.n2161 0.0380882
R43887 PAD.n2450 PAD.n2161 0.0380882
R43888 PAD.n2450 PAD.n2449 0.0380882
R43889 PAD.n2449 PAD.n2448 0.0380882
R43890 PAD.n2448 PAD.n2165 0.0380882
R43891 PAD.n2438 PAD.n2165 0.0380882
R43892 PAD.n2438 PAD.n2437 0.0380882
R43893 PAD.n2437 PAD.n2436 0.0380882
R43894 PAD.n2436 PAD.n2169 0.0380882
R43895 PAD.n2426 PAD.n2169 0.0380882
R43896 PAD.n2426 PAD.n2425 0.0380882
R43897 PAD.n2425 PAD.n2424 0.0380882
R43898 PAD.n2424 PAD.n2173 0.0380882
R43899 PAD.n2414 PAD.n2173 0.0380882
R43900 PAD.n2414 PAD.n2413 0.0380882
R43901 PAD.n2413 PAD.n2412 0.0380882
R43902 PAD.n2412 PAD.n2177 0.0380882
R43903 PAD.n2402 PAD.n2177 0.0380882
R43904 PAD.n2402 PAD.n2401 0.0380882
R43905 PAD.n2401 PAD.n2400 0.0380882
R43906 PAD.n2400 PAD.n2181 0.0380882
R43907 PAD.n2390 PAD.n2181 0.0380882
R43908 PAD.n2390 PAD.n2389 0.0380882
R43909 PAD.n2389 PAD.n2388 0.0380882
R43910 PAD.n2388 PAD.n2185 0.0380882
R43911 PAD.n2378 PAD.n2185 0.0380882
R43912 PAD.n2378 PAD.n2377 0.0380882
R43913 PAD.n2377 PAD.n2376 0.0380882
R43914 PAD.n2376 PAD.n2189 0.0380882
R43915 PAD.n2366 PAD.n2189 0.0380882
R43916 PAD.n2366 PAD.n2365 0.0380882
R43917 PAD.n2365 PAD.n2364 0.0380882
R43918 PAD.n2364 PAD.n2193 0.0380882
R43919 PAD.n2354 PAD.n2193 0.0380882
R43920 PAD.n2354 PAD.n2353 0.0380882
R43921 PAD.n2353 PAD.n2352 0.0380882
R43922 PAD.n2352 PAD.n2197 0.0380882
R43923 PAD.n2342 PAD.n2197 0.0380882
R43924 PAD.n2342 PAD.n2341 0.0380882
R43925 PAD.n2341 PAD.n2340 0.0380882
R43926 PAD.n2340 PAD.n2201 0.0380882
R43927 PAD.n2330 PAD.n2201 0.0380882
R43928 PAD.n2330 PAD.n2329 0.0380882
R43929 PAD.n2329 PAD.n2328 0.0380882
R43930 PAD.n2328 PAD.n2205 0.0380882
R43931 PAD.n2318 PAD.n2205 0.0380882
R43932 PAD.n2318 PAD.n2317 0.0380882
R43933 PAD.n2317 PAD.n2316 0.0380882
R43934 PAD.n2316 PAD.n2209 0.0380882
R43935 PAD.n2306 PAD.n2209 0.0380882
R43936 PAD.n2306 PAD.n2305 0.0380882
R43937 PAD.n2305 PAD.n2304 0.0380882
R43938 PAD.n2304 PAD.n2213 0.0380882
R43939 PAD.n2294 PAD.n2213 0.0380882
R43940 PAD.n2294 PAD.n2293 0.0380882
R43941 PAD.n2293 PAD.n2292 0.0380882
R43942 PAD.n2292 PAD.n2217 0.0380882
R43943 PAD.n2282 PAD.n2217 0.0380882
R43944 PAD.n2282 PAD.n2281 0.0380882
R43945 PAD.n2281 PAD.n2280 0.0380882
R43946 PAD.n2280 PAD.n2221 0.0380882
R43947 PAD.n2270 PAD.n2221 0.0380882
R43948 PAD.n2270 PAD.n2269 0.0380882
R43949 PAD.n2269 PAD.n2268 0.0380882
R43950 PAD.n2268 PAD.n2225 0.0380882
R43951 PAD.n2258 PAD.n2225 0.0380882
R43952 PAD.n2258 PAD.n2257 0.0380882
R43953 PAD.n2257 PAD.n2256 0.0380882
R43954 PAD.n2256 PAD.n2229 0.0380882
R43955 PAD.n2246 PAD.n2229 0.0380882
R43956 PAD.n2246 PAD.n2245 0.0380882
R43957 PAD.n2245 PAD.n2244 0.0380882
R43958 PAD.n2244 PAD.n2233 0.0380882
R43959 PAD.n2233 PAD.n2142 0.0380882
R43960 PAD.n2829 PAD.n2828 0.0380882
R43961 PAD.n2828 PAD.n2499 0.0380882
R43962 PAD.n2822 PAD.n2499 0.0380882
R43963 PAD.n2822 PAD.n2502 0.0380882
R43964 PAD.n2818 PAD.n2502 0.0380882
R43965 PAD.n2818 PAD.n2505 0.0380882
R43966 PAD.n2810 PAD.n2505 0.0380882
R43967 PAD.n2810 PAD.n2507 0.0380882
R43968 PAD.n2806 PAD.n2507 0.0380882
R43969 PAD.n2806 PAD.n2509 0.0380882
R43970 PAD.n2798 PAD.n2509 0.0380882
R43971 PAD.n2798 PAD.n2511 0.0380882
R43972 PAD.n2794 PAD.n2511 0.0380882
R43973 PAD.n2794 PAD.n2513 0.0380882
R43974 PAD.n2786 PAD.n2513 0.0380882
R43975 PAD.n2786 PAD.n2515 0.0380882
R43976 PAD.n2782 PAD.n2515 0.0380882
R43977 PAD.n2782 PAD.n2517 0.0380882
R43978 PAD.n2774 PAD.n2517 0.0380882
R43979 PAD.n2774 PAD.n2519 0.0380882
R43980 PAD.n2770 PAD.n2519 0.0380882
R43981 PAD.n2770 PAD.n2521 0.0380882
R43982 PAD.n2762 PAD.n2521 0.0380882
R43983 PAD.n2762 PAD.n2523 0.0380882
R43984 PAD.n2758 PAD.n2523 0.0380882
R43985 PAD.n2758 PAD.n2525 0.0380882
R43986 PAD.n2750 PAD.n2525 0.0380882
R43987 PAD.n2750 PAD.n2527 0.0380882
R43988 PAD.n2746 PAD.n2527 0.0380882
R43989 PAD.n2746 PAD.n2529 0.0380882
R43990 PAD.n2738 PAD.n2529 0.0380882
R43991 PAD.n2738 PAD.n2531 0.0380882
R43992 PAD.n2734 PAD.n2531 0.0380882
R43993 PAD.n2734 PAD.n2533 0.0380882
R43994 PAD.n2726 PAD.n2533 0.0380882
R43995 PAD.n2726 PAD.n2535 0.0380882
R43996 PAD.n2722 PAD.n2535 0.0380882
R43997 PAD.n2722 PAD.n2537 0.0380882
R43998 PAD.n2714 PAD.n2537 0.0380882
R43999 PAD.n2714 PAD.n2539 0.0380882
R44000 PAD.n2710 PAD.n2539 0.0380882
R44001 PAD.n2710 PAD.n2541 0.0380882
R44002 PAD.n2702 PAD.n2541 0.0380882
R44003 PAD.n2702 PAD.n2543 0.0380882
R44004 PAD.n2698 PAD.n2543 0.0380882
R44005 PAD.n2698 PAD.n2545 0.0380882
R44006 PAD.n2690 PAD.n2545 0.0380882
R44007 PAD.n2690 PAD.n2547 0.0380882
R44008 PAD.n2686 PAD.n2547 0.0380882
R44009 PAD.n2686 PAD.n2549 0.0380882
R44010 PAD.n2678 PAD.n2549 0.0380882
R44011 PAD.n2678 PAD.n2551 0.0380882
R44012 PAD.n2674 PAD.n2551 0.0380882
R44013 PAD.n2674 PAD.n2553 0.0380882
R44014 PAD.n2666 PAD.n2553 0.0380882
R44015 PAD.n2666 PAD.n2555 0.0380882
R44016 PAD.n2662 PAD.n2555 0.0380882
R44017 PAD.n2662 PAD.n2557 0.0380882
R44018 PAD.n2654 PAD.n2557 0.0380882
R44019 PAD.n2654 PAD.n2559 0.0380882
R44020 PAD.n2650 PAD.n2559 0.0380882
R44021 PAD.n2650 PAD.n2561 0.0380882
R44022 PAD.n2642 PAD.n2561 0.0380882
R44023 PAD.n2642 PAD.n2563 0.0380882
R44024 PAD.n2638 PAD.n2563 0.0380882
R44025 PAD.n2638 PAD.n2565 0.0380882
R44026 PAD.n2630 PAD.n2565 0.0380882
R44027 PAD.n2630 PAD.n2567 0.0380882
R44028 PAD.n2626 PAD.n2567 0.0380882
R44029 PAD.n2626 PAD.n2569 0.0380882
R44030 PAD.n2618 PAD.n2569 0.0380882
R44031 PAD.n2618 PAD.n2571 0.0380882
R44032 PAD.n2614 PAD.n2571 0.0380882
R44033 PAD.n2614 PAD.n2573 0.0380882
R44034 PAD.n2606 PAD.n2573 0.0380882
R44035 PAD.n2606 PAD.n2575 0.0380882
R44036 PAD.n2602 PAD.n2575 0.0380882
R44037 PAD.n2602 PAD.n2577 0.0380882
R44038 PAD.n2594 PAD.n2577 0.0380882
R44039 PAD.n2594 PAD.n2579 0.0380882
R44040 PAD.n2590 PAD.n2579 0.0380882
R44041 PAD.n2590 PAD.n2581 0.0380882
R44042 PAD.n2582 PAD.n2581 0.0380882
R44043 PAD.n2830 PAD.n2497 0.0380882
R44044 PAD.n2503 PAD.n2497 0.0380882
R44045 PAD.n2821 PAD.n2503 0.0380882
R44046 PAD.n2821 PAD.n2820 0.0380882
R44047 PAD.n2820 PAD.n2819 0.0380882
R44048 PAD.n2819 PAD.n2504 0.0380882
R44049 PAD.n2809 PAD.n2504 0.0380882
R44050 PAD.n2809 PAD.n2808 0.0380882
R44051 PAD.n2808 PAD.n2807 0.0380882
R44052 PAD.n2807 PAD.n2508 0.0380882
R44053 PAD.n2797 PAD.n2508 0.0380882
R44054 PAD.n2797 PAD.n2796 0.0380882
R44055 PAD.n2796 PAD.n2795 0.0380882
R44056 PAD.n2795 PAD.n2512 0.0380882
R44057 PAD.n2785 PAD.n2512 0.0380882
R44058 PAD.n2785 PAD.n2784 0.0380882
R44059 PAD.n2784 PAD.n2783 0.0380882
R44060 PAD.n2783 PAD.n2516 0.0380882
R44061 PAD.n2773 PAD.n2516 0.0380882
R44062 PAD.n2773 PAD.n2772 0.0380882
R44063 PAD.n2772 PAD.n2771 0.0380882
R44064 PAD.n2771 PAD.n2520 0.0380882
R44065 PAD.n2761 PAD.n2520 0.0380882
R44066 PAD.n2761 PAD.n2760 0.0380882
R44067 PAD.n2760 PAD.n2759 0.0380882
R44068 PAD.n2759 PAD.n2524 0.0380882
R44069 PAD.n2749 PAD.n2524 0.0380882
R44070 PAD.n2749 PAD.n2748 0.0380882
R44071 PAD.n2748 PAD.n2747 0.0380882
R44072 PAD.n2747 PAD.n2528 0.0380882
R44073 PAD.n2737 PAD.n2528 0.0380882
R44074 PAD.n2737 PAD.n2736 0.0380882
R44075 PAD.n2736 PAD.n2735 0.0380882
R44076 PAD.n2735 PAD.n2532 0.0380882
R44077 PAD.n2725 PAD.n2532 0.0380882
R44078 PAD.n2725 PAD.n2724 0.0380882
R44079 PAD.n2724 PAD.n2723 0.0380882
R44080 PAD.n2723 PAD.n2536 0.0380882
R44081 PAD.n2713 PAD.n2536 0.0380882
R44082 PAD.n2713 PAD.n2712 0.0380882
R44083 PAD.n2712 PAD.n2711 0.0380882
R44084 PAD.n2711 PAD.n2540 0.0380882
R44085 PAD.n2701 PAD.n2540 0.0380882
R44086 PAD.n2701 PAD.n2700 0.0380882
R44087 PAD.n2700 PAD.n2699 0.0380882
R44088 PAD.n2699 PAD.n2544 0.0380882
R44089 PAD.n2689 PAD.n2544 0.0380882
R44090 PAD.n2689 PAD.n2688 0.0380882
R44091 PAD.n2688 PAD.n2687 0.0380882
R44092 PAD.n2687 PAD.n2548 0.0380882
R44093 PAD.n2677 PAD.n2548 0.0380882
R44094 PAD.n2677 PAD.n2676 0.0380882
R44095 PAD.n2676 PAD.n2675 0.0380882
R44096 PAD.n2675 PAD.n2552 0.0380882
R44097 PAD.n2665 PAD.n2552 0.0380882
R44098 PAD.n2665 PAD.n2664 0.0380882
R44099 PAD.n2664 PAD.n2663 0.0380882
R44100 PAD.n2663 PAD.n2556 0.0380882
R44101 PAD.n2653 PAD.n2556 0.0380882
R44102 PAD.n2653 PAD.n2652 0.0380882
R44103 PAD.n2652 PAD.n2651 0.0380882
R44104 PAD.n2651 PAD.n2560 0.0380882
R44105 PAD.n2641 PAD.n2560 0.0380882
R44106 PAD.n2641 PAD.n2640 0.0380882
R44107 PAD.n2640 PAD.n2639 0.0380882
R44108 PAD.n2639 PAD.n2564 0.0380882
R44109 PAD.n2629 PAD.n2564 0.0380882
R44110 PAD.n2629 PAD.n2628 0.0380882
R44111 PAD.n2628 PAD.n2627 0.0380882
R44112 PAD.n2627 PAD.n2568 0.0380882
R44113 PAD.n2617 PAD.n2568 0.0380882
R44114 PAD.n2617 PAD.n2616 0.0380882
R44115 PAD.n2616 PAD.n2615 0.0380882
R44116 PAD.n2615 PAD.n2572 0.0380882
R44117 PAD.n2605 PAD.n2572 0.0380882
R44118 PAD.n2605 PAD.n2604 0.0380882
R44119 PAD.n2604 PAD.n2603 0.0380882
R44120 PAD.n2603 PAD.n2576 0.0380882
R44121 PAD.n2593 PAD.n2576 0.0380882
R44122 PAD.n2593 PAD.n2592 0.0380882
R44123 PAD.n2592 PAD.n2591 0.0380882
R44124 PAD.n2591 PAD.n2580 0.0380882
R44125 PAD.n2580 PAD.n2490 0.0380882
R44126 PAD.n9119 PAD.n9118 0.0380882
R44127 PAD.n9118 PAD.n9115 0.0380882
R44128 PAD.n9115 PAD.n8838 0.0380882
R44129 PAD.n9111 PAD.n8838 0.0380882
R44130 PAD.n9111 PAD.n9107 0.0380882
R44131 PAD.n9107 PAD.n9106 0.0380882
R44132 PAD.n9106 PAD.n8843 0.0380882
R44133 PAD.n9102 PAD.n8843 0.0380882
R44134 PAD.n9102 PAD.n9098 0.0380882
R44135 PAD.n9098 PAD.n9097 0.0380882
R44136 PAD.n9097 PAD.n8848 0.0380882
R44137 PAD.n9093 PAD.n8848 0.0380882
R44138 PAD.n9093 PAD.n9089 0.0380882
R44139 PAD.n9089 PAD.n9088 0.0380882
R44140 PAD.n9088 PAD.n8853 0.0380882
R44141 PAD.n9084 PAD.n8853 0.0380882
R44142 PAD.n9084 PAD.n9080 0.0380882
R44143 PAD.n9080 PAD.n9079 0.0380882
R44144 PAD.n9079 PAD.n8858 0.0380882
R44145 PAD.n9075 PAD.n8858 0.0380882
R44146 PAD.n9075 PAD.n9071 0.0380882
R44147 PAD.n9071 PAD.n9070 0.0380882
R44148 PAD.n9070 PAD.n8863 0.0380882
R44149 PAD.n9066 PAD.n8863 0.0380882
R44150 PAD.n9066 PAD.n9062 0.0380882
R44151 PAD.n9062 PAD.n9061 0.0380882
R44152 PAD.n9061 PAD.n8868 0.0380882
R44153 PAD.n9057 PAD.n8868 0.0380882
R44154 PAD.n9057 PAD.n9053 0.0380882
R44155 PAD.n9053 PAD.n9052 0.0380882
R44156 PAD.n9052 PAD.n8873 0.0380882
R44157 PAD.n9048 PAD.n8873 0.0380882
R44158 PAD.n9048 PAD.n9044 0.0380882
R44159 PAD.n9044 PAD.n9043 0.0380882
R44160 PAD.n9043 PAD.n8878 0.0380882
R44161 PAD.n9039 PAD.n8878 0.0380882
R44162 PAD.n9039 PAD.n9035 0.0380882
R44163 PAD.n9035 PAD.n9034 0.0380882
R44164 PAD.n9034 PAD.n8883 0.0380882
R44165 PAD.n9030 PAD.n8883 0.0380882
R44166 PAD.n9030 PAD.n9026 0.0380882
R44167 PAD.n9026 PAD.n9025 0.0380882
R44168 PAD.n9025 PAD.n8888 0.0380882
R44169 PAD.n9021 PAD.n8888 0.0380882
R44170 PAD.n9021 PAD.n9017 0.0380882
R44171 PAD.n9017 PAD.n9016 0.0380882
R44172 PAD.n9016 PAD.n8893 0.0380882
R44173 PAD.n9012 PAD.n8893 0.0380882
R44174 PAD.n9012 PAD.n9008 0.0380882
R44175 PAD.n9008 PAD.n9007 0.0380882
R44176 PAD.n9007 PAD.n8898 0.0380882
R44177 PAD.n9003 PAD.n8898 0.0380882
R44178 PAD.n9003 PAD.n8999 0.0380882
R44179 PAD.n8999 PAD.n8998 0.0380882
R44180 PAD.n8998 PAD.n8903 0.0380882
R44181 PAD.n8994 PAD.n8903 0.0380882
R44182 PAD.n8994 PAD.n8990 0.0380882
R44183 PAD.n8990 PAD.n8989 0.0380882
R44184 PAD.n8989 PAD.n8908 0.0380882
R44185 PAD.n8985 PAD.n8908 0.0380882
R44186 PAD.n8985 PAD.n8981 0.0380882
R44187 PAD.n8981 PAD.n8980 0.0380882
R44188 PAD.n8980 PAD.n8913 0.0380882
R44189 PAD.n8976 PAD.n8913 0.0380882
R44190 PAD.n8976 PAD.n8972 0.0380882
R44191 PAD.n8972 PAD.n8971 0.0380882
R44192 PAD.n8971 PAD.n8918 0.0380882
R44193 PAD.n8967 PAD.n8918 0.0380882
R44194 PAD.n8967 PAD.n8963 0.0380882
R44195 PAD.n8963 PAD.n8962 0.0380882
R44196 PAD.n8962 PAD.n8923 0.0380882
R44197 PAD.n8958 PAD.n8923 0.0380882
R44198 PAD.n8958 PAD.n8954 0.0380882
R44199 PAD.n8954 PAD.n8953 0.0380882
R44200 PAD.n8953 PAD.n8928 0.0380882
R44201 PAD.n8949 PAD.n8928 0.0380882
R44202 PAD.n8949 PAD.n8945 0.0380882
R44203 PAD.n8945 PAD.n8944 0.0380882
R44204 PAD.n8944 PAD.n8933 0.0380882
R44205 PAD.n8940 PAD.n8933 0.0380882
R44206 PAD.n8940 PAD.n2880 0.0380882
R44207 PAD.n9136 PAD.n2880 0.0380882
R44208 PAD.n9136 PAD.n2877 0.0380882
R44209 PAD.n9120 PAD.n8837 0.0380882
R44210 PAD.n9114 PAD.n8837 0.0380882
R44211 PAD.n9114 PAD.n9113 0.0380882
R44212 PAD.n9113 PAD.n9112 0.0380882
R44213 PAD.n9112 PAD.n8842 0.0380882
R44214 PAD.n9105 PAD.n8842 0.0380882
R44215 PAD.n9105 PAD.n9104 0.0380882
R44216 PAD.n9104 PAD.n9103 0.0380882
R44217 PAD.n9103 PAD.n8847 0.0380882
R44218 PAD.n9096 PAD.n8847 0.0380882
R44219 PAD.n9096 PAD.n9095 0.0380882
R44220 PAD.n9095 PAD.n9094 0.0380882
R44221 PAD.n9094 PAD.n8852 0.0380882
R44222 PAD.n9087 PAD.n8852 0.0380882
R44223 PAD.n9087 PAD.n9086 0.0380882
R44224 PAD.n9086 PAD.n9085 0.0380882
R44225 PAD.n9085 PAD.n8857 0.0380882
R44226 PAD.n9078 PAD.n8857 0.0380882
R44227 PAD.n9078 PAD.n9077 0.0380882
R44228 PAD.n9077 PAD.n9076 0.0380882
R44229 PAD.n9076 PAD.n8862 0.0380882
R44230 PAD.n9069 PAD.n8862 0.0380882
R44231 PAD.n9069 PAD.n9068 0.0380882
R44232 PAD.n9068 PAD.n9067 0.0380882
R44233 PAD.n9067 PAD.n8867 0.0380882
R44234 PAD.n9060 PAD.n8867 0.0380882
R44235 PAD.n9060 PAD.n9059 0.0380882
R44236 PAD.n9059 PAD.n9058 0.0380882
R44237 PAD.n9058 PAD.n8872 0.0380882
R44238 PAD.n9051 PAD.n8872 0.0380882
R44239 PAD.n9051 PAD.n9050 0.0380882
R44240 PAD.n9050 PAD.n9049 0.0380882
R44241 PAD.n9049 PAD.n8877 0.0380882
R44242 PAD.n9042 PAD.n8877 0.0380882
R44243 PAD.n9042 PAD.n9041 0.0380882
R44244 PAD.n9041 PAD.n9040 0.0380882
R44245 PAD.n9040 PAD.n8882 0.0380882
R44246 PAD.n9033 PAD.n8882 0.0380882
R44247 PAD.n9033 PAD.n9032 0.0380882
R44248 PAD.n9032 PAD.n9031 0.0380882
R44249 PAD.n9031 PAD.n8887 0.0380882
R44250 PAD.n9024 PAD.n8887 0.0380882
R44251 PAD.n9024 PAD.n9023 0.0380882
R44252 PAD.n9023 PAD.n9022 0.0380882
R44253 PAD.n9022 PAD.n8892 0.0380882
R44254 PAD.n9015 PAD.n8892 0.0380882
R44255 PAD.n9015 PAD.n9014 0.0380882
R44256 PAD.n9014 PAD.n9013 0.0380882
R44257 PAD.n9013 PAD.n8897 0.0380882
R44258 PAD.n9006 PAD.n8897 0.0380882
R44259 PAD.n9006 PAD.n9005 0.0380882
R44260 PAD.n9005 PAD.n9004 0.0380882
R44261 PAD.n9004 PAD.n8902 0.0380882
R44262 PAD.n8997 PAD.n8902 0.0380882
R44263 PAD.n8997 PAD.n8996 0.0380882
R44264 PAD.n8996 PAD.n8995 0.0380882
R44265 PAD.n8995 PAD.n8907 0.0380882
R44266 PAD.n8988 PAD.n8907 0.0380882
R44267 PAD.n8988 PAD.n8987 0.0380882
R44268 PAD.n8987 PAD.n8986 0.0380882
R44269 PAD.n8986 PAD.n8912 0.0380882
R44270 PAD.n8979 PAD.n8912 0.0380882
R44271 PAD.n8979 PAD.n8978 0.0380882
R44272 PAD.n8978 PAD.n8977 0.0380882
R44273 PAD.n8977 PAD.n8917 0.0380882
R44274 PAD.n8970 PAD.n8917 0.0380882
R44275 PAD.n8970 PAD.n8969 0.0380882
R44276 PAD.n8969 PAD.n8968 0.0380882
R44277 PAD.n8968 PAD.n8922 0.0380882
R44278 PAD.n8961 PAD.n8922 0.0380882
R44279 PAD.n8961 PAD.n8960 0.0380882
R44280 PAD.n8960 PAD.n8959 0.0380882
R44281 PAD.n8959 PAD.n8927 0.0380882
R44282 PAD.n8952 PAD.n8927 0.0380882
R44283 PAD.n8952 PAD.n8951 0.0380882
R44284 PAD.n8951 PAD.n8950 0.0380882
R44285 PAD.n8950 PAD.n8932 0.0380882
R44286 PAD.n8943 PAD.n8932 0.0380882
R44287 PAD.n8943 PAD.n8942 0.0380882
R44288 PAD.n8942 PAD.n8941 0.0380882
R44289 PAD.n8941 PAD.n2881 0.0380882
R44290 PAD.n9135 PAD.n2881 0.0380882
R44291 PAD.n9135 PAD.n9134 0.0380882
R44292 PAD.n8818 PAD.n8529 0.0380882
R44293 PAD.n8814 PAD.n8529 0.0380882
R44294 PAD.n8814 PAD.n8811 0.0380882
R44295 PAD.n8811 PAD.n8807 0.0380882
R44296 PAD.n8807 PAD.n8531 0.0380882
R44297 PAD.n8803 PAD.n8531 0.0380882
R44298 PAD.n8803 PAD.n8799 0.0380882
R44299 PAD.n8799 PAD.n8795 0.0380882
R44300 PAD.n8795 PAD.n8533 0.0380882
R44301 PAD.n8791 PAD.n8533 0.0380882
R44302 PAD.n8791 PAD.n8787 0.0380882
R44303 PAD.n8787 PAD.n8783 0.0380882
R44304 PAD.n8783 PAD.n8535 0.0380882
R44305 PAD.n8779 PAD.n8535 0.0380882
R44306 PAD.n8779 PAD.n8775 0.0380882
R44307 PAD.n8775 PAD.n8771 0.0380882
R44308 PAD.n8771 PAD.n8537 0.0380882
R44309 PAD.n8767 PAD.n8537 0.0380882
R44310 PAD.n8767 PAD.n8763 0.0380882
R44311 PAD.n8763 PAD.n8759 0.0380882
R44312 PAD.n8759 PAD.n8539 0.0380882
R44313 PAD.n8755 PAD.n8539 0.0380882
R44314 PAD.n8755 PAD.n8751 0.0380882
R44315 PAD.n8751 PAD.n8747 0.0380882
R44316 PAD.n8747 PAD.n8541 0.0380882
R44317 PAD.n8743 PAD.n8541 0.0380882
R44318 PAD.n8743 PAD.n8739 0.0380882
R44319 PAD.n8739 PAD.n8735 0.0380882
R44320 PAD.n8735 PAD.n8543 0.0380882
R44321 PAD.n8731 PAD.n8543 0.0380882
R44322 PAD.n8731 PAD.n8727 0.0380882
R44323 PAD.n8727 PAD.n8723 0.0380882
R44324 PAD.n8723 PAD.n8545 0.0380882
R44325 PAD.n8719 PAD.n8545 0.0380882
R44326 PAD.n8719 PAD.n8715 0.0380882
R44327 PAD.n8715 PAD.n8711 0.0380882
R44328 PAD.n8711 PAD.n8547 0.0380882
R44329 PAD.n8707 PAD.n8547 0.0380882
R44330 PAD.n8707 PAD.n8703 0.0380882
R44331 PAD.n8703 PAD.n8699 0.0380882
R44332 PAD.n8699 PAD.n8549 0.0380882
R44333 PAD.n8695 PAD.n8549 0.0380882
R44334 PAD.n8695 PAD.n8691 0.0380882
R44335 PAD.n8691 PAD.n8687 0.0380882
R44336 PAD.n8687 PAD.n8551 0.0380882
R44337 PAD.n8683 PAD.n8551 0.0380882
R44338 PAD.n8683 PAD.n8679 0.0380882
R44339 PAD.n8679 PAD.n8675 0.0380882
R44340 PAD.n8675 PAD.n8553 0.0380882
R44341 PAD.n8671 PAD.n8553 0.0380882
R44342 PAD.n8671 PAD.n8667 0.0380882
R44343 PAD.n8667 PAD.n8663 0.0380882
R44344 PAD.n8663 PAD.n8555 0.0380882
R44345 PAD.n8659 PAD.n8555 0.0380882
R44346 PAD.n8659 PAD.n8655 0.0380882
R44347 PAD.n8655 PAD.n8651 0.0380882
R44348 PAD.n8651 PAD.n8557 0.0380882
R44349 PAD.n8647 PAD.n8557 0.0380882
R44350 PAD.n8647 PAD.n8643 0.0380882
R44351 PAD.n8643 PAD.n8639 0.0380882
R44352 PAD.n8639 PAD.n8559 0.0380882
R44353 PAD.n8635 PAD.n8559 0.0380882
R44354 PAD.n8635 PAD.n8631 0.0380882
R44355 PAD.n8631 PAD.n8627 0.0380882
R44356 PAD.n8627 PAD.n8561 0.0380882
R44357 PAD.n8623 PAD.n8561 0.0380882
R44358 PAD.n8623 PAD.n8619 0.0380882
R44359 PAD.n8619 PAD.n8615 0.0380882
R44360 PAD.n8615 PAD.n8563 0.0380882
R44361 PAD.n8611 PAD.n8563 0.0380882
R44362 PAD.n8611 PAD.n8607 0.0380882
R44363 PAD.n8607 PAD.n8603 0.0380882
R44364 PAD.n8603 PAD.n8565 0.0380882
R44365 PAD.n8599 PAD.n8565 0.0380882
R44366 PAD.n8599 PAD.n8595 0.0380882
R44367 PAD.n8595 PAD.n8591 0.0380882
R44368 PAD.n8591 PAD.n8567 0.0380882
R44369 PAD.n8587 PAD.n8567 0.0380882
R44370 PAD.n8587 PAD.n8583 0.0380882
R44371 PAD.n8583 PAD.n8579 0.0380882
R44372 PAD.n8579 PAD.n8569 0.0380882
R44373 PAD.n8575 PAD.n8569 0.0380882
R44374 PAD.n8575 PAD.n8571 0.0380882
R44375 PAD.n8817 PAD.n8816 0.0380882
R44376 PAD.n8816 PAD.n8815 0.0380882
R44377 PAD.n8815 PAD.n8530 0.0380882
R44378 PAD.n8806 PAD.n8530 0.0380882
R44379 PAD.n8806 PAD.n8805 0.0380882
R44380 PAD.n8805 PAD.n8804 0.0380882
R44381 PAD.n8804 PAD.n8532 0.0380882
R44382 PAD.n8794 PAD.n8532 0.0380882
R44383 PAD.n8794 PAD.n8793 0.0380882
R44384 PAD.n8793 PAD.n8792 0.0380882
R44385 PAD.n8792 PAD.n8534 0.0380882
R44386 PAD.n8782 PAD.n8534 0.0380882
R44387 PAD.n8782 PAD.n8781 0.0380882
R44388 PAD.n8781 PAD.n8780 0.0380882
R44389 PAD.n8780 PAD.n8536 0.0380882
R44390 PAD.n8770 PAD.n8536 0.0380882
R44391 PAD.n8770 PAD.n8769 0.0380882
R44392 PAD.n8769 PAD.n8768 0.0380882
R44393 PAD.n8768 PAD.n8538 0.0380882
R44394 PAD.n8758 PAD.n8538 0.0380882
R44395 PAD.n8758 PAD.n8757 0.0380882
R44396 PAD.n8757 PAD.n8756 0.0380882
R44397 PAD.n8756 PAD.n8540 0.0380882
R44398 PAD.n8746 PAD.n8540 0.0380882
R44399 PAD.n8746 PAD.n8745 0.0380882
R44400 PAD.n8745 PAD.n8744 0.0380882
R44401 PAD.n8744 PAD.n8542 0.0380882
R44402 PAD.n8734 PAD.n8542 0.0380882
R44403 PAD.n8734 PAD.n8733 0.0380882
R44404 PAD.n8733 PAD.n8732 0.0380882
R44405 PAD.n8732 PAD.n8544 0.0380882
R44406 PAD.n8722 PAD.n8544 0.0380882
R44407 PAD.n8722 PAD.n8721 0.0380882
R44408 PAD.n8721 PAD.n8720 0.0380882
R44409 PAD.n8720 PAD.n8546 0.0380882
R44410 PAD.n8710 PAD.n8546 0.0380882
R44411 PAD.n8710 PAD.n8709 0.0380882
R44412 PAD.n8709 PAD.n8708 0.0380882
R44413 PAD.n8708 PAD.n8548 0.0380882
R44414 PAD.n8698 PAD.n8548 0.0380882
R44415 PAD.n8698 PAD.n8697 0.0380882
R44416 PAD.n8697 PAD.n8696 0.0380882
R44417 PAD.n8696 PAD.n8550 0.0380882
R44418 PAD.n8686 PAD.n8550 0.0380882
R44419 PAD.n8686 PAD.n8685 0.0380882
R44420 PAD.n8685 PAD.n8684 0.0380882
R44421 PAD.n8684 PAD.n8552 0.0380882
R44422 PAD.n8674 PAD.n8552 0.0380882
R44423 PAD.n8674 PAD.n8673 0.0380882
R44424 PAD.n8673 PAD.n8672 0.0380882
R44425 PAD.n8672 PAD.n8554 0.0380882
R44426 PAD.n8662 PAD.n8554 0.0380882
R44427 PAD.n8662 PAD.n8661 0.0380882
R44428 PAD.n8661 PAD.n8660 0.0380882
R44429 PAD.n8660 PAD.n8556 0.0380882
R44430 PAD.n8650 PAD.n8556 0.0380882
R44431 PAD.n8650 PAD.n8649 0.0380882
R44432 PAD.n8649 PAD.n8648 0.0380882
R44433 PAD.n8648 PAD.n8558 0.0380882
R44434 PAD.n8638 PAD.n8558 0.0380882
R44435 PAD.n8638 PAD.n8637 0.0380882
R44436 PAD.n8637 PAD.n8636 0.0380882
R44437 PAD.n8636 PAD.n8560 0.0380882
R44438 PAD.n8626 PAD.n8560 0.0380882
R44439 PAD.n8626 PAD.n8625 0.0380882
R44440 PAD.n8625 PAD.n8624 0.0380882
R44441 PAD.n8624 PAD.n8562 0.0380882
R44442 PAD.n8614 PAD.n8562 0.0380882
R44443 PAD.n8614 PAD.n8613 0.0380882
R44444 PAD.n8613 PAD.n8612 0.0380882
R44445 PAD.n8612 PAD.n8564 0.0380882
R44446 PAD.n8602 PAD.n8564 0.0380882
R44447 PAD.n8602 PAD.n8601 0.0380882
R44448 PAD.n8601 PAD.n8600 0.0380882
R44449 PAD.n8600 PAD.n8566 0.0380882
R44450 PAD.n8590 PAD.n8566 0.0380882
R44451 PAD.n8590 PAD.n8589 0.0380882
R44452 PAD.n8589 PAD.n8588 0.0380882
R44453 PAD.n8588 PAD.n8568 0.0380882
R44454 PAD.n8578 PAD.n8568 0.0380882
R44455 PAD.n8578 PAD.n8577 0.0380882
R44456 PAD.n8577 PAD.n8576 0.0380882
R44457 PAD.n8576 PAD.n2898 0.0380882
R44458 PAD.n3041 PAD.n3040 0.0380882
R44459 PAD.n3045 PAD.n3040 0.0380882
R44460 PAD.n3049 PAD.n3045 0.0380882
R44461 PAD.n3053 PAD.n3049 0.0380882
R44462 PAD.n3053 PAD.n3036 0.0380882
R44463 PAD.n3057 PAD.n3036 0.0380882
R44464 PAD.n3061 PAD.n3057 0.0380882
R44465 PAD.n3065 PAD.n3061 0.0380882
R44466 PAD.n3065 PAD.n3034 0.0380882
R44467 PAD.n3069 PAD.n3034 0.0380882
R44468 PAD.n3073 PAD.n3069 0.0380882
R44469 PAD.n3077 PAD.n3073 0.0380882
R44470 PAD.n3077 PAD.n3032 0.0380882
R44471 PAD.n3081 PAD.n3032 0.0380882
R44472 PAD.n3085 PAD.n3081 0.0380882
R44473 PAD.n3089 PAD.n3085 0.0380882
R44474 PAD.n3089 PAD.n3030 0.0380882
R44475 PAD.n3093 PAD.n3030 0.0380882
R44476 PAD.n3097 PAD.n3093 0.0380882
R44477 PAD.n3101 PAD.n3097 0.0380882
R44478 PAD.n3101 PAD.n3028 0.0380882
R44479 PAD.n3105 PAD.n3028 0.0380882
R44480 PAD.n3109 PAD.n3105 0.0380882
R44481 PAD.n3113 PAD.n3109 0.0380882
R44482 PAD.n3113 PAD.n3026 0.0380882
R44483 PAD.n3117 PAD.n3026 0.0380882
R44484 PAD.n3121 PAD.n3117 0.0380882
R44485 PAD.n3125 PAD.n3121 0.0380882
R44486 PAD.n3125 PAD.n3024 0.0380882
R44487 PAD.n3129 PAD.n3024 0.0380882
R44488 PAD.n3133 PAD.n3129 0.0380882
R44489 PAD.n3137 PAD.n3133 0.0380882
R44490 PAD.n3137 PAD.n3022 0.0380882
R44491 PAD.n3141 PAD.n3022 0.0380882
R44492 PAD.n3145 PAD.n3141 0.0380882
R44493 PAD.n3149 PAD.n3145 0.0380882
R44494 PAD.n3149 PAD.n3020 0.0380882
R44495 PAD.n3153 PAD.n3020 0.0380882
R44496 PAD.n3157 PAD.n3153 0.0380882
R44497 PAD.n3161 PAD.n3157 0.0380882
R44498 PAD.n3161 PAD.n3018 0.0380882
R44499 PAD.n3165 PAD.n3018 0.0380882
R44500 PAD.n3169 PAD.n3165 0.0380882
R44501 PAD.n3173 PAD.n3169 0.0380882
R44502 PAD.n3173 PAD.n3016 0.0380882
R44503 PAD.n3177 PAD.n3016 0.0380882
R44504 PAD.n3181 PAD.n3177 0.0380882
R44505 PAD.n3185 PAD.n3181 0.0380882
R44506 PAD.n3185 PAD.n3014 0.0380882
R44507 PAD.n3189 PAD.n3014 0.0380882
R44508 PAD.n3193 PAD.n3189 0.0380882
R44509 PAD.n3197 PAD.n3193 0.0380882
R44510 PAD.n3197 PAD.n3012 0.0380882
R44511 PAD.n3201 PAD.n3012 0.0380882
R44512 PAD.n3205 PAD.n3201 0.0380882
R44513 PAD.n3209 PAD.n3205 0.0380882
R44514 PAD.n3209 PAD.n3010 0.0380882
R44515 PAD.n3213 PAD.n3010 0.0380882
R44516 PAD.n3217 PAD.n3213 0.0380882
R44517 PAD.n3221 PAD.n3217 0.0380882
R44518 PAD.n3221 PAD.n3008 0.0380882
R44519 PAD.n3225 PAD.n3008 0.0380882
R44520 PAD.n3229 PAD.n3225 0.0380882
R44521 PAD.n3233 PAD.n3229 0.0380882
R44522 PAD.n3233 PAD.n3006 0.0380882
R44523 PAD.n3237 PAD.n3006 0.0380882
R44524 PAD.n3241 PAD.n3237 0.0380882
R44525 PAD.n3245 PAD.n3241 0.0380882
R44526 PAD.n3245 PAD.n3004 0.0380882
R44527 PAD.n3249 PAD.n3004 0.0380882
R44528 PAD.n3253 PAD.n3249 0.0380882
R44529 PAD.n3257 PAD.n3253 0.0380882
R44530 PAD.n3257 PAD.n3002 0.0380882
R44531 PAD.n3261 PAD.n3002 0.0380882
R44532 PAD.n3265 PAD.n3261 0.0380882
R44533 PAD.n3269 PAD.n3265 0.0380882
R44534 PAD.n3269 PAD.n3000 0.0380882
R44535 PAD.n3273 PAD.n3000 0.0380882
R44536 PAD.n3277 PAD.n3273 0.0380882
R44537 PAD.n3281 PAD.n3277 0.0380882
R44538 PAD.n3281 PAD.n2998 0.0380882
R44539 PAD.n8513 PAD.n2998 0.0380882
R44540 PAD.n8513 PAD.n2995 0.0380882
R44541 PAD.n3043 PAD.n3042 0.0380882
R44542 PAD.n3044 PAD.n3043 0.0380882
R44543 PAD.n3044 PAD.n3037 0.0380882
R44544 PAD.n3054 PAD.n3037 0.0380882
R44545 PAD.n3055 PAD.n3054 0.0380882
R44546 PAD.n3056 PAD.n3055 0.0380882
R44547 PAD.n3056 PAD.n3035 0.0380882
R44548 PAD.n3066 PAD.n3035 0.0380882
R44549 PAD.n3067 PAD.n3066 0.0380882
R44550 PAD.n3068 PAD.n3067 0.0380882
R44551 PAD.n3068 PAD.n3033 0.0380882
R44552 PAD.n3078 PAD.n3033 0.0380882
R44553 PAD.n3079 PAD.n3078 0.0380882
R44554 PAD.n3080 PAD.n3079 0.0380882
R44555 PAD.n3080 PAD.n3031 0.0380882
R44556 PAD.n3090 PAD.n3031 0.0380882
R44557 PAD.n3091 PAD.n3090 0.0380882
R44558 PAD.n3092 PAD.n3091 0.0380882
R44559 PAD.n3092 PAD.n3029 0.0380882
R44560 PAD.n3102 PAD.n3029 0.0380882
R44561 PAD.n3103 PAD.n3102 0.0380882
R44562 PAD.n3104 PAD.n3103 0.0380882
R44563 PAD.n3104 PAD.n3027 0.0380882
R44564 PAD.n3114 PAD.n3027 0.0380882
R44565 PAD.n3115 PAD.n3114 0.0380882
R44566 PAD.n3116 PAD.n3115 0.0380882
R44567 PAD.n3116 PAD.n3025 0.0380882
R44568 PAD.n3126 PAD.n3025 0.0380882
R44569 PAD.n3127 PAD.n3126 0.0380882
R44570 PAD.n3128 PAD.n3127 0.0380882
R44571 PAD.n3128 PAD.n3023 0.0380882
R44572 PAD.n3138 PAD.n3023 0.0380882
R44573 PAD.n3139 PAD.n3138 0.0380882
R44574 PAD.n3140 PAD.n3139 0.0380882
R44575 PAD.n3140 PAD.n3021 0.0380882
R44576 PAD.n3150 PAD.n3021 0.0380882
R44577 PAD.n3151 PAD.n3150 0.0380882
R44578 PAD.n3152 PAD.n3151 0.0380882
R44579 PAD.n3152 PAD.n3019 0.0380882
R44580 PAD.n3162 PAD.n3019 0.0380882
R44581 PAD.n3163 PAD.n3162 0.0380882
R44582 PAD.n3164 PAD.n3163 0.0380882
R44583 PAD.n3164 PAD.n3017 0.0380882
R44584 PAD.n3174 PAD.n3017 0.0380882
R44585 PAD.n3175 PAD.n3174 0.0380882
R44586 PAD.n3176 PAD.n3175 0.0380882
R44587 PAD.n3176 PAD.n3015 0.0380882
R44588 PAD.n3186 PAD.n3015 0.0380882
R44589 PAD.n3187 PAD.n3186 0.0380882
R44590 PAD.n3188 PAD.n3187 0.0380882
R44591 PAD.n3188 PAD.n3013 0.0380882
R44592 PAD.n3198 PAD.n3013 0.0380882
R44593 PAD.n3199 PAD.n3198 0.0380882
R44594 PAD.n3200 PAD.n3199 0.0380882
R44595 PAD.n3200 PAD.n3011 0.0380882
R44596 PAD.n3210 PAD.n3011 0.0380882
R44597 PAD.n3211 PAD.n3210 0.0380882
R44598 PAD.n3212 PAD.n3211 0.0380882
R44599 PAD.n3212 PAD.n3009 0.0380882
R44600 PAD.n3222 PAD.n3009 0.0380882
R44601 PAD.n3223 PAD.n3222 0.0380882
R44602 PAD.n3224 PAD.n3223 0.0380882
R44603 PAD.n3224 PAD.n3007 0.0380882
R44604 PAD.n3234 PAD.n3007 0.0380882
R44605 PAD.n3235 PAD.n3234 0.0380882
R44606 PAD.n3236 PAD.n3235 0.0380882
R44607 PAD.n3236 PAD.n3005 0.0380882
R44608 PAD.n3246 PAD.n3005 0.0380882
R44609 PAD.n3247 PAD.n3246 0.0380882
R44610 PAD.n3248 PAD.n3247 0.0380882
R44611 PAD.n3248 PAD.n3003 0.0380882
R44612 PAD.n3258 PAD.n3003 0.0380882
R44613 PAD.n3259 PAD.n3258 0.0380882
R44614 PAD.n3260 PAD.n3259 0.0380882
R44615 PAD.n3260 PAD.n3001 0.0380882
R44616 PAD.n3270 PAD.n3001 0.0380882
R44617 PAD.n3271 PAD.n3270 0.0380882
R44618 PAD.n3272 PAD.n3271 0.0380882
R44619 PAD.n3272 PAD.n2999 0.0380882
R44620 PAD.n3282 PAD.n2999 0.0380882
R44621 PAD.n3283 PAD.n3282 0.0380882
R44622 PAD.n8512 PAD.n3283 0.0380882
R44623 PAD.n8512 PAD.n8511 0.0380882
R44624 PAD.n3386 PAD.n3385 0.0380882
R44625 PAD.n3390 PAD.n3385 0.0380882
R44626 PAD.n3394 PAD.n3390 0.0380882
R44627 PAD.n3398 PAD.n3394 0.0380882
R44628 PAD.n3398 PAD.n3381 0.0380882
R44629 PAD.n3402 PAD.n3381 0.0380882
R44630 PAD.n3406 PAD.n3402 0.0380882
R44631 PAD.n3410 PAD.n3406 0.0380882
R44632 PAD.n3410 PAD.n3379 0.0380882
R44633 PAD.n3414 PAD.n3379 0.0380882
R44634 PAD.n3418 PAD.n3414 0.0380882
R44635 PAD.n3422 PAD.n3418 0.0380882
R44636 PAD.n3422 PAD.n3377 0.0380882
R44637 PAD.n3426 PAD.n3377 0.0380882
R44638 PAD.n3430 PAD.n3426 0.0380882
R44639 PAD.n3434 PAD.n3430 0.0380882
R44640 PAD.n3434 PAD.n3375 0.0380882
R44641 PAD.n3438 PAD.n3375 0.0380882
R44642 PAD.n3442 PAD.n3438 0.0380882
R44643 PAD.n3446 PAD.n3442 0.0380882
R44644 PAD.n3446 PAD.n3373 0.0380882
R44645 PAD.n3450 PAD.n3373 0.0380882
R44646 PAD.n3454 PAD.n3450 0.0380882
R44647 PAD.n3458 PAD.n3454 0.0380882
R44648 PAD.n3458 PAD.n3371 0.0380882
R44649 PAD.n3462 PAD.n3371 0.0380882
R44650 PAD.n3466 PAD.n3462 0.0380882
R44651 PAD.n3470 PAD.n3466 0.0380882
R44652 PAD.n3470 PAD.n3369 0.0380882
R44653 PAD.n3474 PAD.n3369 0.0380882
R44654 PAD.n3478 PAD.n3474 0.0380882
R44655 PAD.n3482 PAD.n3478 0.0380882
R44656 PAD.n3482 PAD.n3367 0.0380882
R44657 PAD.n3486 PAD.n3367 0.0380882
R44658 PAD.n3490 PAD.n3486 0.0380882
R44659 PAD.n3494 PAD.n3490 0.0380882
R44660 PAD.n3494 PAD.n3365 0.0380882
R44661 PAD.n3498 PAD.n3365 0.0380882
R44662 PAD.n3502 PAD.n3498 0.0380882
R44663 PAD.n3506 PAD.n3502 0.0380882
R44664 PAD.n3506 PAD.n3363 0.0380882
R44665 PAD.n3510 PAD.n3363 0.0380882
R44666 PAD.n3514 PAD.n3510 0.0380882
R44667 PAD.n3518 PAD.n3514 0.0380882
R44668 PAD.n3518 PAD.n3361 0.0380882
R44669 PAD.n3522 PAD.n3361 0.0380882
R44670 PAD.n3526 PAD.n3522 0.0380882
R44671 PAD.n3530 PAD.n3526 0.0380882
R44672 PAD.n3530 PAD.n3359 0.0380882
R44673 PAD.n3534 PAD.n3359 0.0380882
R44674 PAD.n3538 PAD.n3534 0.0380882
R44675 PAD.n3542 PAD.n3538 0.0380882
R44676 PAD.n3542 PAD.n3357 0.0380882
R44677 PAD.n3546 PAD.n3357 0.0380882
R44678 PAD.n3550 PAD.n3546 0.0380882
R44679 PAD.n3554 PAD.n3550 0.0380882
R44680 PAD.n3554 PAD.n3355 0.0380882
R44681 PAD.n3558 PAD.n3355 0.0380882
R44682 PAD.n3562 PAD.n3558 0.0380882
R44683 PAD.n3566 PAD.n3562 0.0380882
R44684 PAD.n3566 PAD.n3353 0.0380882
R44685 PAD.n3570 PAD.n3353 0.0380882
R44686 PAD.n3574 PAD.n3570 0.0380882
R44687 PAD.n3578 PAD.n3574 0.0380882
R44688 PAD.n3578 PAD.n3351 0.0380882
R44689 PAD.n3582 PAD.n3351 0.0380882
R44690 PAD.n3586 PAD.n3582 0.0380882
R44691 PAD.n3590 PAD.n3586 0.0380882
R44692 PAD.n3590 PAD.n3349 0.0380882
R44693 PAD.n3594 PAD.n3349 0.0380882
R44694 PAD.n3598 PAD.n3594 0.0380882
R44695 PAD.n3602 PAD.n3598 0.0380882
R44696 PAD.n3602 PAD.n3347 0.0380882
R44697 PAD.n3606 PAD.n3347 0.0380882
R44698 PAD.n3610 PAD.n3606 0.0380882
R44699 PAD.n3614 PAD.n3610 0.0380882
R44700 PAD.n3614 PAD.n3345 0.0380882
R44701 PAD.n3618 PAD.n3345 0.0380882
R44702 PAD.n3622 PAD.n3618 0.0380882
R44703 PAD.n3626 PAD.n3622 0.0380882
R44704 PAD.n3626 PAD.n3343 0.0380882
R44705 PAD.n8488 PAD.n3343 0.0380882
R44706 PAD.n8488 PAD.n3340 0.0380882
R44707 PAD.n3388 PAD.n3387 0.0380882
R44708 PAD.n3389 PAD.n3388 0.0380882
R44709 PAD.n3389 PAD.n3382 0.0380882
R44710 PAD.n3399 PAD.n3382 0.0380882
R44711 PAD.n3400 PAD.n3399 0.0380882
R44712 PAD.n3401 PAD.n3400 0.0380882
R44713 PAD.n3401 PAD.n3380 0.0380882
R44714 PAD.n3411 PAD.n3380 0.0380882
R44715 PAD.n3412 PAD.n3411 0.0380882
R44716 PAD.n3413 PAD.n3412 0.0380882
R44717 PAD.n3413 PAD.n3378 0.0380882
R44718 PAD.n3423 PAD.n3378 0.0380882
R44719 PAD.n3424 PAD.n3423 0.0380882
R44720 PAD.n3425 PAD.n3424 0.0380882
R44721 PAD.n3425 PAD.n3376 0.0380882
R44722 PAD.n3435 PAD.n3376 0.0380882
R44723 PAD.n3436 PAD.n3435 0.0380882
R44724 PAD.n3437 PAD.n3436 0.0380882
R44725 PAD.n3437 PAD.n3374 0.0380882
R44726 PAD.n3447 PAD.n3374 0.0380882
R44727 PAD.n3448 PAD.n3447 0.0380882
R44728 PAD.n3449 PAD.n3448 0.0380882
R44729 PAD.n3449 PAD.n3372 0.0380882
R44730 PAD.n3459 PAD.n3372 0.0380882
R44731 PAD.n3460 PAD.n3459 0.0380882
R44732 PAD.n3461 PAD.n3460 0.0380882
R44733 PAD.n3461 PAD.n3370 0.0380882
R44734 PAD.n3471 PAD.n3370 0.0380882
R44735 PAD.n3472 PAD.n3471 0.0380882
R44736 PAD.n3473 PAD.n3472 0.0380882
R44737 PAD.n3473 PAD.n3368 0.0380882
R44738 PAD.n3483 PAD.n3368 0.0380882
R44739 PAD.n3484 PAD.n3483 0.0380882
R44740 PAD.n3485 PAD.n3484 0.0380882
R44741 PAD.n3485 PAD.n3366 0.0380882
R44742 PAD.n3495 PAD.n3366 0.0380882
R44743 PAD.n3496 PAD.n3495 0.0380882
R44744 PAD.n3497 PAD.n3496 0.0380882
R44745 PAD.n3497 PAD.n3364 0.0380882
R44746 PAD.n3507 PAD.n3364 0.0380882
R44747 PAD.n3508 PAD.n3507 0.0380882
R44748 PAD.n3509 PAD.n3508 0.0380882
R44749 PAD.n3509 PAD.n3362 0.0380882
R44750 PAD.n3519 PAD.n3362 0.0380882
R44751 PAD.n3520 PAD.n3519 0.0380882
R44752 PAD.n3521 PAD.n3520 0.0380882
R44753 PAD.n3521 PAD.n3360 0.0380882
R44754 PAD.n3531 PAD.n3360 0.0380882
R44755 PAD.n3532 PAD.n3531 0.0380882
R44756 PAD.n3533 PAD.n3532 0.0380882
R44757 PAD.n3533 PAD.n3358 0.0380882
R44758 PAD.n3543 PAD.n3358 0.0380882
R44759 PAD.n3544 PAD.n3543 0.0380882
R44760 PAD.n3545 PAD.n3544 0.0380882
R44761 PAD.n3545 PAD.n3356 0.0380882
R44762 PAD.n3555 PAD.n3356 0.0380882
R44763 PAD.n3556 PAD.n3555 0.0380882
R44764 PAD.n3557 PAD.n3556 0.0380882
R44765 PAD.n3557 PAD.n3354 0.0380882
R44766 PAD.n3567 PAD.n3354 0.0380882
R44767 PAD.n3568 PAD.n3567 0.0380882
R44768 PAD.n3569 PAD.n3568 0.0380882
R44769 PAD.n3569 PAD.n3352 0.0380882
R44770 PAD.n3579 PAD.n3352 0.0380882
R44771 PAD.n3580 PAD.n3579 0.0380882
R44772 PAD.n3581 PAD.n3580 0.0380882
R44773 PAD.n3581 PAD.n3350 0.0380882
R44774 PAD.n3591 PAD.n3350 0.0380882
R44775 PAD.n3592 PAD.n3591 0.0380882
R44776 PAD.n3593 PAD.n3592 0.0380882
R44777 PAD.n3593 PAD.n3348 0.0380882
R44778 PAD.n3603 PAD.n3348 0.0380882
R44779 PAD.n3604 PAD.n3603 0.0380882
R44780 PAD.n3605 PAD.n3604 0.0380882
R44781 PAD.n3605 PAD.n3346 0.0380882
R44782 PAD.n3615 PAD.n3346 0.0380882
R44783 PAD.n3616 PAD.n3615 0.0380882
R44784 PAD.n3617 PAD.n3616 0.0380882
R44785 PAD.n3617 PAD.n3344 0.0380882
R44786 PAD.n3627 PAD.n3344 0.0380882
R44787 PAD.n3628 PAD.n3627 0.0380882
R44788 PAD.n8487 PAD.n3628 0.0380882
R44789 PAD.n8487 PAD.n8486 0.0380882
R44790 PAD.n3731 PAD.n3730 0.0380882
R44791 PAD.n3735 PAD.n3730 0.0380882
R44792 PAD.n3739 PAD.n3735 0.0380882
R44793 PAD.n3743 PAD.n3739 0.0380882
R44794 PAD.n3743 PAD.n3726 0.0380882
R44795 PAD.n3747 PAD.n3726 0.0380882
R44796 PAD.n3751 PAD.n3747 0.0380882
R44797 PAD.n3755 PAD.n3751 0.0380882
R44798 PAD.n3755 PAD.n3724 0.0380882
R44799 PAD.n3759 PAD.n3724 0.0380882
R44800 PAD.n3763 PAD.n3759 0.0380882
R44801 PAD.n3767 PAD.n3763 0.0380882
R44802 PAD.n3767 PAD.n3722 0.0380882
R44803 PAD.n3771 PAD.n3722 0.0380882
R44804 PAD.n3775 PAD.n3771 0.0380882
R44805 PAD.n3779 PAD.n3775 0.0380882
R44806 PAD.n3779 PAD.n3720 0.0380882
R44807 PAD.n3783 PAD.n3720 0.0380882
R44808 PAD.n3787 PAD.n3783 0.0380882
R44809 PAD.n3791 PAD.n3787 0.0380882
R44810 PAD.n3791 PAD.n3718 0.0380882
R44811 PAD.n3795 PAD.n3718 0.0380882
R44812 PAD.n3799 PAD.n3795 0.0380882
R44813 PAD.n3803 PAD.n3799 0.0380882
R44814 PAD.n3803 PAD.n3716 0.0380882
R44815 PAD.n3807 PAD.n3716 0.0380882
R44816 PAD.n3811 PAD.n3807 0.0380882
R44817 PAD.n3815 PAD.n3811 0.0380882
R44818 PAD.n3815 PAD.n3714 0.0380882
R44819 PAD.n3819 PAD.n3714 0.0380882
R44820 PAD.n3823 PAD.n3819 0.0380882
R44821 PAD.n3827 PAD.n3823 0.0380882
R44822 PAD.n3827 PAD.n3712 0.0380882
R44823 PAD.n3831 PAD.n3712 0.0380882
R44824 PAD.n3835 PAD.n3831 0.0380882
R44825 PAD.n3839 PAD.n3835 0.0380882
R44826 PAD.n3839 PAD.n3710 0.0380882
R44827 PAD.n3843 PAD.n3710 0.0380882
R44828 PAD.n3847 PAD.n3843 0.0380882
R44829 PAD.n3851 PAD.n3847 0.0380882
R44830 PAD.n3851 PAD.n3708 0.0380882
R44831 PAD.n3855 PAD.n3708 0.0380882
R44832 PAD.n3859 PAD.n3855 0.0380882
R44833 PAD.n3863 PAD.n3859 0.0380882
R44834 PAD.n3863 PAD.n3706 0.0380882
R44835 PAD.n3867 PAD.n3706 0.0380882
R44836 PAD.n3871 PAD.n3867 0.0380882
R44837 PAD.n3875 PAD.n3871 0.0380882
R44838 PAD.n3875 PAD.n3704 0.0380882
R44839 PAD.n3879 PAD.n3704 0.0380882
R44840 PAD.n3883 PAD.n3879 0.0380882
R44841 PAD.n3887 PAD.n3883 0.0380882
R44842 PAD.n3887 PAD.n3702 0.0380882
R44843 PAD.n3891 PAD.n3702 0.0380882
R44844 PAD.n3895 PAD.n3891 0.0380882
R44845 PAD.n3899 PAD.n3895 0.0380882
R44846 PAD.n3899 PAD.n3700 0.0380882
R44847 PAD.n3903 PAD.n3700 0.0380882
R44848 PAD.n3907 PAD.n3903 0.0380882
R44849 PAD.n3911 PAD.n3907 0.0380882
R44850 PAD.n3911 PAD.n3698 0.0380882
R44851 PAD.n3915 PAD.n3698 0.0380882
R44852 PAD.n3919 PAD.n3915 0.0380882
R44853 PAD.n3923 PAD.n3919 0.0380882
R44854 PAD.n3923 PAD.n3696 0.0380882
R44855 PAD.n3927 PAD.n3696 0.0380882
R44856 PAD.n3931 PAD.n3927 0.0380882
R44857 PAD.n3935 PAD.n3931 0.0380882
R44858 PAD.n3935 PAD.n3694 0.0380882
R44859 PAD.n3939 PAD.n3694 0.0380882
R44860 PAD.n3943 PAD.n3939 0.0380882
R44861 PAD.n3947 PAD.n3943 0.0380882
R44862 PAD.n3947 PAD.n3692 0.0380882
R44863 PAD.n3951 PAD.n3692 0.0380882
R44864 PAD.n3955 PAD.n3951 0.0380882
R44865 PAD.n3959 PAD.n3955 0.0380882
R44866 PAD.n3959 PAD.n3690 0.0380882
R44867 PAD.n3963 PAD.n3690 0.0380882
R44868 PAD.n3967 PAD.n3963 0.0380882
R44869 PAD.n3971 PAD.n3967 0.0380882
R44870 PAD.n3971 PAD.n3688 0.0380882
R44871 PAD.n8464 PAD.n3688 0.0380882
R44872 PAD.n8464 PAD.n3685 0.0380882
R44873 PAD.n3733 PAD.n3732 0.0380882
R44874 PAD.n3734 PAD.n3733 0.0380882
R44875 PAD.n3734 PAD.n3727 0.0380882
R44876 PAD.n3744 PAD.n3727 0.0380882
R44877 PAD.n3745 PAD.n3744 0.0380882
R44878 PAD.n3746 PAD.n3745 0.0380882
R44879 PAD.n3746 PAD.n3725 0.0380882
R44880 PAD.n3756 PAD.n3725 0.0380882
R44881 PAD.n3757 PAD.n3756 0.0380882
R44882 PAD.n3758 PAD.n3757 0.0380882
R44883 PAD.n3758 PAD.n3723 0.0380882
R44884 PAD.n3768 PAD.n3723 0.0380882
R44885 PAD.n3769 PAD.n3768 0.0380882
R44886 PAD.n3770 PAD.n3769 0.0380882
R44887 PAD.n3770 PAD.n3721 0.0380882
R44888 PAD.n3780 PAD.n3721 0.0380882
R44889 PAD.n3781 PAD.n3780 0.0380882
R44890 PAD.n3782 PAD.n3781 0.0380882
R44891 PAD.n3782 PAD.n3719 0.0380882
R44892 PAD.n3792 PAD.n3719 0.0380882
R44893 PAD.n3793 PAD.n3792 0.0380882
R44894 PAD.n3794 PAD.n3793 0.0380882
R44895 PAD.n3794 PAD.n3717 0.0380882
R44896 PAD.n3804 PAD.n3717 0.0380882
R44897 PAD.n3805 PAD.n3804 0.0380882
R44898 PAD.n3806 PAD.n3805 0.0380882
R44899 PAD.n3806 PAD.n3715 0.0380882
R44900 PAD.n3816 PAD.n3715 0.0380882
R44901 PAD.n3817 PAD.n3816 0.0380882
R44902 PAD.n3818 PAD.n3817 0.0380882
R44903 PAD.n3818 PAD.n3713 0.0380882
R44904 PAD.n3828 PAD.n3713 0.0380882
R44905 PAD.n3829 PAD.n3828 0.0380882
R44906 PAD.n3830 PAD.n3829 0.0380882
R44907 PAD.n3830 PAD.n3711 0.0380882
R44908 PAD.n3840 PAD.n3711 0.0380882
R44909 PAD.n3841 PAD.n3840 0.0380882
R44910 PAD.n3842 PAD.n3841 0.0380882
R44911 PAD.n3842 PAD.n3709 0.0380882
R44912 PAD.n3852 PAD.n3709 0.0380882
R44913 PAD.n3853 PAD.n3852 0.0380882
R44914 PAD.n3854 PAD.n3853 0.0380882
R44915 PAD.n3854 PAD.n3707 0.0380882
R44916 PAD.n3864 PAD.n3707 0.0380882
R44917 PAD.n3865 PAD.n3864 0.0380882
R44918 PAD.n3866 PAD.n3865 0.0380882
R44919 PAD.n3866 PAD.n3705 0.0380882
R44920 PAD.n3876 PAD.n3705 0.0380882
R44921 PAD.n3877 PAD.n3876 0.0380882
R44922 PAD.n3878 PAD.n3877 0.0380882
R44923 PAD.n3878 PAD.n3703 0.0380882
R44924 PAD.n3888 PAD.n3703 0.0380882
R44925 PAD.n3889 PAD.n3888 0.0380882
R44926 PAD.n3890 PAD.n3889 0.0380882
R44927 PAD.n3890 PAD.n3701 0.0380882
R44928 PAD.n3900 PAD.n3701 0.0380882
R44929 PAD.n3901 PAD.n3900 0.0380882
R44930 PAD.n3902 PAD.n3901 0.0380882
R44931 PAD.n3902 PAD.n3699 0.0380882
R44932 PAD.n3912 PAD.n3699 0.0380882
R44933 PAD.n3913 PAD.n3912 0.0380882
R44934 PAD.n3914 PAD.n3913 0.0380882
R44935 PAD.n3914 PAD.n3697 0.0380882
R44936 PAD.n3924 PAD.n3697 0.0380882
R44937 PAD.n3925 PAD.n3924 0.0380882
R44938 PAD.n3926 PAD.n3925 0.0380882
R44939 PAD.n3926 PAD.n3695 0.0380882
R44940 PAD.n3936 PAD.n3695 0.0380882
R44941 PAD.n3937 PAD.n3936 0.0380882
R44942 PAD.n3938 PAD.n3937 0.0380882
R44943 PAD.n3938 PAD.n3693 0.0380882
R44944 PAD.n3948 PAD.n3693 0.0380882
R44945 PAD.n3949 PAD.n3948 0.0380882
R44946 PAD.n3950 PAD.n3949 0.0380882
R44947 PAD.n3950 PAD.n3691 0.0380882
R44948 PAD.n3960 PAD.n3691 0.0380882
R44949 PAD.n3961 PAD.n3960 0.0380882
R44950 PAD.n3962 PAD.n3961 0.0380882
R44951 PAD.n3962 PAD.n3689 0.0380882
R44952 PAD.n3972 PAD.n3689 0.0380882
R44953 PAD.n3973 PAD.n3972 0.0380882
R44954 PAD.n8463 PAD.n3973 0.0380882
R44955 PAD.n8463 PAD.n8462 0.0380882
R44956 PAD.n4072 PAD.n4071 0.0380882
R44957 PAD.n4076 PAD.n4071 0.0380882
R44958 PAD.n4080 PAD.n4076 0.0380882
R44959 PAD.n4084 PAD.n4080 0.0380882
R44960 PAD.n4084 PAD.n4067 0.0380882
R44961 PAD.n4088 PAD.n4067 0.0380882
R44962 PAD.n4092 PAD.n4088 0.0380882
R44963 PAD.n4096 PAD.n4092 0.0380882
R44964 PAD.n4096 PAD.n4065 0.0380882
R44965 PAD.n4100 PAD.n4065 0.0380882
R44966 PAD.n4104 PAD.n4100 0.0380882
R44967 PAD.n4108 PAD.n4104 0.0380882
R44968 PAD.n4108 PAD.n4063 0.0380882
R44969 PAD.n4112 PAD.n4063 0.0380882
R44970 PAD.n4116 PAD.n4112 0.0380882
R44971 PAD.n4120 PAD.n4116 0.0380882
R44972 PAD.n4120 PAD.n4061 0.0380882
R44973 PAD.n4124 PAD.n4061 0.0380882
R44974 PAD.n4128 PAD.n4124 0.0380882
R44975 PAD.n4132 PAD.n4128 0.0380882
R44976 PAD.n4132 PAD.n4059 0.0380882
R44977 PAD.n4136 PAD.n4059 0.0380882
R44978 PAD.n4140 PAD.n4136 0.0380882
R44979 PAD.n4144 PAD.n4140 0.0380882
R44980 PAD.n4144 PAD.n4057 0.0380882
R44981 PAD.n4148 PAD.n4057 0.0380882
R44982 PAD.n4152 PAD.n4148 0.0380882
R44983 PAD.n4156 PAD.n4152 0.0380882
R44984 PAD.n4156 PAD.n4055 0.0380882
R44985 PAD.n4160 PAD.n4055 0.0380882
R44986 PAD.n4164 PAD.n4160 0.0380882
R44987 PAD.n4168 PAD.n4164 0.0380882
R44988 PAD.n4168 PAD.n4053 0.0380882
R44989 PAD.n4172 PAD.n4053 0.0380882
R44990 PAD.n4176 PAD.n4172 0.0380882
R44991 PAD.n4180 PAD.n4176 0.0380882
R44992 PAD.n4180 PAD.n4051 0.0380882
R44993 PAD.n4184 PAD.n4051 0.0380882
R44994 PAD.n4188 PAD.n4184 0.0380882
R44995 PAD.n4192 PAD.n4188 0.0380882
R44996 PAD.n4192 PAD.n4049 0.0380882
R44997 PAD.n4196 PAD.n4049 0.0380882
R44998 PAD.n4200 PAD.n4196 0.0380882
R44999 PAD.n4204 PAD.n4200 0.0380882
R45000 PAD.n4204 PAD.n4047 0.0380882
R45001 PAD.n4208 PAD.n4047 0.0380882
R45002 PAD.n4212 PAD.n4208 0.0380882
R45003 PAD.n4216 PAD.n4212 0.0380882
R45004 PAD.n4216 PAD.n4045 0.0380882
R45005 PAD.n4220 PAD.n4045 0.0380882
R45006 PAD.n4224 PAD.n4220 0.0380882
R45007 PAD.n4228 PAD.n4224 0.0380882
R45008 PAD.n4228 PAD.n4043 0.0380882
R45009 PAD.n4232 PAD.n4043 0.0380882
R45010 PAD.n4236 PAD.n4232 0.0380882
R45011 PAD.n4240 PAD.n4236 0.0380882
R45012 PAD.n4240 PAD.n4041 0.0380882
R45013 PAD.n4244 PAD.n4041 0.0380882
R45014 PAD.n4248 PAD.n4244 0.0380882
R45015 PAD.n4252 PAD.n4248 0.0380882
R45016 PAD.n4252 PAD.n4039 0.0380882
R45017 PAD.n4256 PAD.n4039 0.0380882
R45018 PAD.n4260 PAD.n4256 0.0380882
R45019 PAD.n4264 PAD.n4260 0.0380882
R45020 PAD.n4264 PAD.n4037 0.0380882
R45021 PAD.n4268 PAD.n4037 0.0380882
R45022 PAD.n4272 PAD.n4268 0.0380882
R45023 PAD.n4276 PAD.n4272 0.0380882
R45024 PAD.n4276 PAD.n4035 0.0380882
R45025 PAD.n4280 PAD.n4035 0.0380882
R45026 PAD.n4284 PAD.n4280 0.0380882
R45027 PAD.n4288 PAD.n4284 0.0380882
R45028 PAD.n4288 PAD.n4033 0.0380882
R45029 PAD.n4292 PAD.n4033 0.0380882
R45030 PAD.n4296 PAD.n4292 0.0380882
R45031 PAD.n4300 PAD.n4296 0.0380882
R45032 PAD.n4300 PAD.n4031 0.0380882
R45033 PAD.n4304 PAD.n4031 0.0380882
R45034 PAD.n4308 PAD.n4304 0.0380882
R45035 PAD.n4312 PAD.n4308 0.0380882
R45036 PAD.n4312 PAD.n4029 0.0380882
R45037 PAD.n8440 PAD.n4029 0.0380882
R45038 PAD.n8440 PAD.n4026 0.0380882
R45039 PAD.n4074 PAD.n4073 0.0380882
R45040 PAD.n4075 PAD.n4074 0.0380882
R45041 PAD.n4075 PAD.n4068 0.0380882
R45042 PAD.n4085 PAD.n4068 0.0380882
R45043 PAD.n4086 PAD.n4085 0.0380882
R45044 PAD.n4087 PAD.n4086 0.0380882
R45045 PAD.n4087 PAD.n4066 0.0380882
R45046 PAD.n4097 PAD.n4066 0.0380882
R45047 PAD.n4098 PAD.n4097 0.0380882
R45048 PAD.n4099 PAD.n4098 0.0380882
R45049 PAD.n4099 PAD.n4064 0.0380882
R45050 PAD.n4109 PAD.n4064 0.0380882
R45051 PAD.n4110 PAD.n4109 0.0380882
R45052 PAD.n4111 PAD.n4110 0.0380882
R45053 PAD.n4111 PAD.n4062 0.0380882
R45054 PAD.n4121 PAD.n4062 0.0380882
R45055 PAD.n4122 PAD.n4121 0.0380882
R45056 PAD.n4123 PAD.n4122 0.0380882
R45057 PAD.n4123 PAD.n4060 0.0380882
R45058 PAD.n4133 PAD.n4060 0.0380882
R45059 PAD.n4134 PAD.n4133 0.0380882
R45060 PAD.n4135 PAD.n4134 0.0380882
R45061 PAD.n4135 PAD.n4058 0.0380882
R45062 PAD.n4145 PAD.n4058 0.0380882
R45063 PAD.n4146 PAD.n4145 0.0380882
R45064 PAD.n4147 PAD.n4146 0.0380882
R45065 PAD.n4147 PAD.n4056 0.0380882
R45066 PAD.n4157 PAD.n4056 0.0380882
R45067 PAD.n4158 PAD.n4157 0.0380882
R45068 PAD.n4159 PAD.n4158 0.0380882
R45069 PAD.n4159 PAD.n4054 0.0380882
R45070 PAD.n4169 PAD.n4054 0.0380882
R45071 PAD.n4170 PAD.n4169 0.0380882
R45072 PAD.n4171 PAD.n4170 0.0380882
R45073 PAD.n4171 PAD.n4052 0.0380882
R45074 PAD.n4181 PAD.n4052 0.0380882
R45075 PAD.n4182 PAD.n4181 0.0380882
R45076 PAD.n4183 PAD.n4182 0.0380882
R45077 PAD.n4183 PAD.n4050 0.0380882
R45078 PAD.n4193 PAD.n4050 0.0380882
R45079 PAD.n4194 PAD.n4193 0.0380882
R45080 PAD.n4195 PAD.n4194 0.0380882
R45081 PAD.n4195 PAD.n4048 0.0380882
R45082 PAD.n4205 PAD.n4048 0.0380882
R45083 PAD.n4206 PAD.n4205 0.0380882
R45084 PAD.n4207 PAD.n4206 0.0380882
R45085 PAD.n4207 PAD.n4046 0.0380882
R45086 PAD.n4217 PAD.n4046 0.0380882
R45087 PAD.n4218 PAD.n4217 0.0380882
R45088 PAD.n4219 PAD.n4218 0.0380882
R45089 PAD.n4219 PAD.n4044 0.0380882
R45090 PAD.n4229 PAD.n4044 0.0380882
R45091 PAD.n4230 PAD.n4229 0.0380882
R45092 PAD.n4231 PAD.n4230 0.0380882
R45093 PAD.n4231 PAD.n4042 0.0380882
R45094 PAD.n4241 PAD.n4042 0.0380882
R45095 PAD.n4242 PAD.n4241 0.0380882
R45096 PAD.n4243 PAD.n4242 0.0380882
R45097 PAD.n4243 PAD.n4040 0.0380882
R45098 PAD.n4253 PAD.n4040 0.0380882
R45099 PAD.n4254 PAD.n4253 0.0380882
R45100 PAD.n4255 PAD.n4254 0.0380882
R45101 PAD.n4255 PAD.n4038 0.0380882
R45102 PAD.n4265 PAD.n4038 0.0380882
R45103 PAD.n4266 PAD.n4265 0.0380882
R45104 PAD.n4267 PAD.n4266 0.0380882
R45105 PAD.n4267 PAD.n4036 0.0380882
R45106 PAD.n4277 PAD.n4036 0.0380882
R45107 PAD.n4278 PAD.n4277 0.0380882
R45108 PAD.n4279 PAD.n4278 0.0380882
R45109 PAD.n4279 PAD.n4034 0.0380882
R45110 PAD.n4289 PAD.n4034 0.0380882
R45111 PAD.n4290 PAD.n4289 0.0380882
R45112 PAD.n4291 PAD.n4290 0.0380882
R45113 PAD.n4291 PAD.n4032 0.0380882
R45114 PAD.n4301 PAD.n4032 0.0380882
R45115 PAD.n4302 PAD.n4301 0.0380882
R45116 PAD.n4303 PAD.n4302 0.0380882
R45117 PAD.n4303 PAD.n4030 0.0380882
R45118 PAD.n4313 PAD.n4030 0.0380882
R45119 PAD.n4314 PAD.n4313 0.0380882
R45120 PAD.n8439 PAD.n4314 0.0380882
R45121 PAD.n8439 PAD.n8438 0.0380882
R45122 PAD.n4419 PAD.n4418 0.0380882
R45123 PAD.n4427 PAD.n4418 0.0380882
R45124 PAD.n4427 PAD.n4416 0.0380882
R45125 PAD.n4431 PAD.n4416 0.0380882
R45126 PAD.n4431 PAD.n4414 0.0380882
R45127 PAD.n4439 PAD.n4414 0.0380882
R45128 PAD.n4439 PAD.n4412 0.0380882
R45129 PAD.n4443 PAD.n4412 0.0380882
R45130 PAD.n4443 PAD.n4410 0.0380882
R45131 PAD.n4451 PAD.n4410 0.0380882
R45132 PAD.n4451 PAD.n4408 0.0380882
R45133 PAD.n4455 PAD.n4408 0.0380882
R45134 PAD.n4455 PAD.n4406 0.0380882
R45135 PAD.n4463 PAD.n4406 0.0380882
R45136 PAD.n4463 PAD.n4404 0.0380882
R45137 PAD.n4467 PAD.n4404 0.0380882
R45138 PAD.n4467 PAD.n4402 0.0380882
R45139 PAD.n4475 PAD.n4402 0.0380882
R45140 PAD.n4475 PAD.n4400 0.0380882
R45141 PAD.n4479 PAD.n4400 0.0380882
R45142 PAD.n4479 PAD.n4398 0.0380882
R45143 PAD.n4487 PAD.n4398 0.0380882
R45144 PAD.n4487 PAD.n4396 0.0380882
R45145 PAD.n4491 PAD.n4396 0.0380882
R45146 PAD.n4491 PAD.n4394 0.0380882
R45147 PAD.n4499 PAD.n4394 0.0380882
R45148 PAD.n4499 PAD.n4392 0.0380882
R45149 PAD.n4503 PAD.n4392 0.0380882
R45150 PAD.n4503 PAD.n4390 0.0380882
R45151 PAD.n4511 PAD.n4390 0.0380882
R45152 PAD.n4511 PAD.n4388 0.0380882
R45153 PAD.n4515 PAD.n4388 0.0380882
R45154 PAD.n4515 PAD.n4386 0.0380882
R45155 PAD.n4523 PAD.n4386 0.0380882
R45156 PAD.n4523 PAD.n4384 0.0380882
R45157 PAD.n4527 PAD.n4384 0.0380882
R45158 PAD.n4527 PAD.n4382 0.0380882
R45159 PAD.n4535 PAD.n4382 0.0380882
R45160 PAD.n4535 PAD.n4380 0.0380882
R45161 PAD.n4539 PAD.n4380 0.0380882
R45162 PAD.n4539 PAD.n4378 0.0380882
R45163 PAD.n4547 PAD.n4378 0.0380882
R45164 PAD.n4547 PAD.n4376 0.0380882
R45165 PAD.n4551 PAD.n4376 0.0380882
R45166 PAD.n4551 PAD.n4374 0.0380882
R45167 PAD.n4559 PAD.n4374 0.0380882
R45168 PAD.n4559 PAD.n4372 0.0380882
R45169 PAD.n4563 PAD.n4372 0.0380882
R45170 PAD.n4563 PAD.n4370 0.0380882
R45171 PAD.n4571 PAD.n4370 0.0380882
R45172 PAD.n4571 PAD.n4368 0.0380882
R45173 PAD.n4575 PAD.n4368 0.0380882
R45174 PAD.n4575 PAD.n4366 0.0380882
R45175 PAD.n4583 PAD.n4366 0.0380882
R45176 PAD.n4583 PAD.n4364 0.0380882
R45177 PAD.n4587 PAD.n4364 0.0380882
R45178 PAD.n4587 PAD.n4362 0.0380882
R45179 PAD.n4595 PAD.n4362 0.0380882
R45180 PAD.n4595 PAD.n4360 0.0380882
R45181 PAD.n4599 PAD.n4360 0.0380882
R45182 PAD.n4599 PAD.n4358 0.0380882
R45183 PAD.n4607 PAD.n4358 0.0380882
R45184 PAD.n4607 PAD.n4356 0.0380882
R45185 PAD.n4611 PAD.n4356 0.0380882
R45186 PAD.n4611 PAD.n4354 0.0380882
R45187 PAD.n4619 PAD.n4354 0.0380882
R45188 PAD.n4619 PAD.n4352 0.0380882
R45189 PAD.n4623 PAD.n4352 0.0380882
R45190 PAD.n4623 PAD.n4350 0.0380882
R45191 PAD.n4631 PAD.n4350 0.0380882
R45192 PAD.n4631 PAD.n4348 0.0380882
R45193 PAD.n4635 PAD.n4348 0.0380882
R45194 PAD.n4635 PAD.n4346 0.0380882
R45195 PAD.n4643 PAD.n4346 0.0380882
R45196 PAD.n4643 PAD.n4344 0.0380882
R45197 PAD.n4647 PAD.n4344 0.0380882
R45198 PAD.n4647 PAD.n4342 0.0380882
R45199 PAD.n4655 PAD.n4342 0.0380882
R45200 PAD.n4655 PAD.n4340 0.0380882
R45201 PAD.n4660 PAD.n4340 0.0380882
R45202 PAD.n4660 PAD.n4338 0.0380882
R45203 PAD.n4338 PAD.n4337 0.0380882
R45204 PAD.n4668 PAD.n4337 0.0380882
R45205 PAD.n4417 PAD.n4325 0.0380882
R45206 PAD.n4428 PAD.n4417 0.0380882
R45207 PAD.n4429 PAD.n4428 0.0380882
R45208 PAD.n4430 PAD.n4429 0.0380882
R45209 PAD.n4430 PAD.n4413 0.0380882
R45210 PAD.n4440 PAD.n4413 0.0380882
R45211 PAD.n4441 PAD.n4440 0.0380882
R45212 PAD.n4442 PAD.n4441 0.0380882
R45213 PAD.n4442 PAD.n4409 0.0380882
R45214 PAD.n4452 PAD.n4409 0.0380882
R45215 PAD.n4453 PAD.n4452 0.0380882
R45216 PAD.n4454 PAD.n4453 0.0380882
R45217 PAD.n4454 PAD.n4405 0.0380882
R45218 PAD.n4464 PAD.n4405 0.0380882
R45219 PAD.n4465 PAD.n4464 0.0380882
R45220 PAD.n4466 PAD.n4465 0.0380882
R45221 PAD.n4466 PAD.n4401 0.0380882
R45222 PAD.n4476 PAD.n4401 0.0380882
R45223 PAD.n4477 PAD.n4476 0.0380882
R45224 PAD.n4478 PAD.n4477 0.0380882
R45225 PAD.n4478 PAD.n4397 0.0380882
R45226 PAD.n4488 PAD.n4397 0.0380882
R45227 PAD.n4489 PAD.n4488 0.0380882
R45228 PAD.n4490 PAD.n4489 0.0380882
R45229 PAD.n4490 PAD.n4393 0.0380882
R45230 PAD.n4500 PAD.n4393 0.0380882
R45231 PAD.n4501 PAD.n4500 0.0380882
R45232 PAD.n4502 PAD.n4501 0.0380882
R45233 PAD.n4502 PAD.n4389 0.0380882
R45234 PAD.n4512 PAD.n4389 0.0380882
R45235 PAD.n4513 PAD.n4512 0.0380882
R45236 PAD.n4514 PAD.n4513 0.0380882
R45237 PAD.n4514 PAD.n4385 0.0380882
R45238 PAD.n4524 PAD.n4385 0.0380882
R45239 PAD.n4525 PAD.n4524 0.0380882
R45240 PAD.n4526 PAD.n4525 0.0380882
R45241 PAD.n4526 PAD.n4381 0.0380882
R45242 PAD.n4536 PAD.n4381 0.0380882
R45243 PAD.n4537 PAD.n4536 0.0380882
R45244 PAD.n4538 PAD.n4537 0.0380882
R45245 PAD.n4538 PAD.n4377 0.0380882
R45246 PAD.n4548 PAD.n4377 0.0380882
R45247 PAD.n4549 PAD.n4548 0.0380882
R45248 PAD.n4550 PAD.n4549 0.0380882
R45249 PAD.n4550 PAD.n4373 0.0380882
R45250 PAD.n4560 PAD.n4373 0.0380882
R45251 PAD.n4561 PAD.n4560 0.0380882
R45252 PAD.n4562 PAD.n4561 0.0380882
R45253 PAD.n4562 PAD.n4369 0.0380882
R45254 PAD.n4572 PAD.n4369 0.0380882
R45255 PAD.n4573 PAD.n4572 0.0380882
R45256 PAD.n4574 PAD.n4573 0.0380882
R45257 PAD.n4574 PAD.n4365 0.0380882
R45258 PAD.n4584 PAD.n4365 0.0380882
R45259 PAD.n4585 PAD.n4584 0.0380882
R45260 PAD.n4586 PAD.n4585 0.0380882
R45261 PAD.n4586 PAD.n4361 0.0380882
R45262 PAD.n4596 PAD.n4361 0.0380882
R45263 PAD.n4597 PAD.n4596 0.0380882
R45264 PAD.n4598 PAD.n4597 0.0380882
R45265 PAD.n4598 PAD.n4357 0.0380882
R45266 PAD.n4608 PAD.n4357 0.0380882
R45267 PAD.n4609 PAD.n4608 0.0380882
R45268 PAD.n4610 PAD.n4609 0.0380882
R45269 PAD.n4610 PAD.n4353 0.0380882
R45270 PAD.n4620 PAD.n4353 0.0380882
R45271 PAD.n4621 PAD.n4620 0.0380882
R45272 PAD.n4622 PAD.n4621 0.0380882
R45273 PAD.n4622 PAD.n4349 0.0380882
R45274 PAD.n4632 PAD.n4349 0.0380882
R45275 PAD.n4633 PAD.n4632 0.0380882
R45276 PAD.n4634 PAD.n4633 0.0380882
R45277 PAD.n4634 PAD.n4345 0.0380882
R45278 PAD.n4644 PAD.n4345 0.0380882
R45279 PAD.n4645 PAD.n4644 0.0380882
R45280 PAD.n4646 PAD.n4645 0.0380882
R45281 PAD.n4646 PAD.n4341 0.0380882
R45282 PAD.n4656 PAD.n4341 0.0380882
R45283 PAD.n4657 PAD.n4656 0.0380882
R45284 PAD.n4659 PAD.n4657 0.0380882
R45285 PAD.n4659 PAD.n4658 0.0380882
R45286 PAD.n4658 PAD.n4336 0.0380882
R45287 PAD.n4669 PAD.n4336 0.0380882
R45288 PAD.n8394 PAD.n8393 0.0380882
R45289 PAD.n8393 PAD.n4728 0.0380882
R45290 PAD.n8389 PAD.n4728 0.0380882
R45291 PAD.n8389 PAD.n8385 0.0380882
R45292 PAD.n8385 PAD.n8384 0.0380882
R45293 PAD.n8384 PAD.n4730 0.0380882
R45294 PAD.n8380 PAD.n4730 0.0380882
R45295 PAD.n8380 PAD.n8376 0.0380882
R45296 PAD.n8376 PAD.n8375 0.0380882
R45297 PAD.n8375 PAD.n4735 0.0380882
R45298 PAD.n8371 PAD.n4735 0.0380882
R45299 PAD.n8371 PAD.n8367 0.0380882
R45300 PAD.n8367 PAD.n8366 0.0380882
R45301 PAD.n8366 PAD.n4740 0.0380882
R45302 PAD.n8362 PAD.n4740 0.0380882
R45303 PAD.n8362 PAD.n8358 0.0380882
R45304 PAD.n8358 PAD.n8357 0.0380882
R45305 PAD.n8357 PAD.n4745 0.0380882
R45306 PAD.n8353 PAD.n4745 0.0380882
R45307 PAD.n8353 PAD.n8349 0.0380882
R45308 PAD.n8349 PAD.n8348 0.0380882
R45309 PAD.n8348 PAD.n4750 0.0380882
R45310 PAD.n8344 PAD.n4750 0.0380882
R45311 PAD.n8344 PAD.n8340 0.0380882
R45312 PAD.n8340 PAD.n8339 0.0380882
R45313 PAD.n8339 PAD.n4755 0.0380882
R45314 PAD.n8335 PAD.n4755 0.0380882
R45315 PAD.n8335 PAD.n8331 0.0380882
R45316 PAD.n8331 PAD.n8330 0.0380882
R45317 PAD.n8330 PAD.n4760 0.0380882
R45318 PAD.n8326 PAD.n4760 0.0380882
R45319 PAD.n8326 PAD.n8322 0.0380882
R45320 PAD.n8322 PAD.n8321 0.0380882
R45321 PAD.n8321 PAD.n4765 0.0380882
R45322 PAD.n8317 PAD.n4765 0.0380882
R45323 PAD.n8317 PAD.n8313 0.0380882
R45324 PAD.n8313 PAD.n8312 0.0380882
R45325 PAD.n8312 PAD.n4770 0.0380882
R45326 PAD.n8308 PAD.n4770 0.0380882
R45327 PAD.n8308 PAD.n8304 0.0380882
R45328 PAD.n8304 PAD.n8303 0.0380882
R45329 PAD.n8303 PAD.n4775 0.0380882
R45330 PAD.n8299 PAD.n4775 0.0380882
R45331 PAD.n8299 PAD.n8295 0.0380882
R45332 PAD.n8295 PAD.n8294 0.0380882
R45333 PAD.n8294 PAD.n4780 0.0380882
R45334 PAD.n8290 PAD.n4780 0.0380882
R45335 PAD.n8290 PAD.n8286 0.0380882
R45336 PAD.n8286 PAD.n8285 0.0380882
R45337 PAD.n8285 PAD.n4785 0.0380882
R45338 PAD.n8281 PAD.n4785 0.0380882
R45339 PAD.n8281 PAD.n8277 0.0380882
R45340 PAD.n8277 PAD.n8276 0.0380882
R45341 PAD.n8276 PAD.n4790 0.0380882
R45342 PAD.n8272 PAD.n4790 0.0380882
R45343 PAD.n8272 PAD.n8268 0.0380882
R45344 PAD.n8268 PAD.n8267 0.0380882
R45345 PAD.n8267 PAD.n4795 0.0380882
R45346 PAD.n8263 PAD.n4795 0.0380882
R45347 PAD.n8263 PAD.n8259 0.0380882
R45348 PAD.n8259 PAD.n8258 0.0380882
R45349 PAD.n8258 PAD.n4800 0.0380882
R45350 PAD.n8254 PAD.n4800 0.0380882
R45351 PAD.n8254 PAD.n8250 0.0380882
R45352 PAD.n8250 PAD.n8249 0.0380882
R45353 PAD.n8249 PAD.n4805 0.0380882
R45354 PAD.n8245 PAD.n4805 0.0380882
R45355 PAD.n8245 PAD.n8241 0.0380882
R45356 PAD.n8241 PAD.n8240 0.0380882
R45357 PAD.n8240 PAD.n4810 0.0380882
R45358 PAD.n8236 PAD.n4810 0.0380882
R45359 PAD.n8236 PAD.n8232 0.0380882
R45360 PAD.n8232 PAD.n8231 0.0380882
R45361 PAD.n8231 PAD.n4815 0.0380882
R45362 PAD.n8227 PAD.n4815 0.0380882
R45363 PAD.n8227 PAD.n8223 0.0380882
R45364 PAD.n8223 PAD.n8222 0.0380882
R45365 PAD.n8222 PAD.n4820 0.0380882
R45366 PAD.n8218 PAD.n4820 0.0380882
R45367 PAD.n8218 PAD.n8214 0.0380882
R45368 PAD.n8214 PAD.n8213 0.0380882
R45369 PAD.n8213 PAD.n4825 0.0380882
R45370 PAD.n4829 PAD.n4825 0.0380882
R45371 PAD.n8392 PAD.n4676 0.0380882
R45372 PAD.n8392 PAD.n8391 0.0380882
R45373 PAD.n8391 PAD.n8390 0.0380882
R45374 PAD.n8390 PAD.n4729 0.0380882
R45375 PAD.n8383 PAD.n4729 0.0380882
R45376 PAD.n8383 PAD.n8382 0.0380882
R45377 PAD.n8382 PAD.n8381 0.0380882
R45378 PAD.n8381 PAD.n4734 0.0380882
R45379 PAD.n8374 PAD.n4734 0.0380882
R45380 PAD.n8374 PAD.n8373 0.0380882
R45381 PAD.n8373 PAD.n8372 0.0380882
R45382 PAD.n8372 PAD.n4739 0.0380882
R45383 PAD.n8365 PAD.n4739 0.0380882
R45384 PAD.n8365 PAD.n8364 0.0380882
R45385 PAD.n8364 PAD.n8363 0.0380882
R45386 PAD.n8363 PAD.n4744 0.0380882
R45387 PAD.n8356 PAD.n4744 0.0380882
R45388 PAD.n8356 PAD.n8355 0.0380882
R45389 PAD.n8355 PAD.n8354 0.0380882
R45390 PAD.n8354 PAD.n4749 0.0380882
R45391 PAD.n8347 PAD.n4749 0.0380882
R45392 PAD.n8347 PAD.n8346 0.0380882
R45393 PAD.n8346 PAD.n8345 0.0380882
R45394 PAD.n8345 PAD.n4754 0.0380882
R45395 PAD.n8338 PAD.n4754 0.0380882
R45396 PAD.n8338 PAD.n8337 0.0380882
R45397 PAD.n8337 PAD.n8336 0.0380882
R45398 PAD.n8336 PAD.n4759 0.0380882
R45399 PAD.n8329 PAD.n4759 0.0380882
R45400 PAD.n8329 PAD.n8328 0.0380882
R45401 PAD.n8328 PAD.n8327 0.0380882
R45402 PAD.n8327 PAD.n4764 0.0380882
R45403 PAD.n8320 PAD.n4764 0.0380882
R45404 PAD.n8320 PAD.n8319 0.0380882
R45405 PAD.n8319 PAD.n8318 0.0380882
R45406 PAD.n8318 PAD.n4769 0.0380882
R45407 PAD.n8311 PAD.n4769 0.0380882
R45408 PAD.n8311 PAD.n8310 0.0380882
R45409 PAD.n8310 PAD.n8309 0.0380882
R45410 PAD.n8309 PAD.n4774 0.0380882
R45411 PAD.n8302 PAD.n4774 0.0380882
R45412 PAD.n8302 PAD.n8301 0.0380882
R45413 PAD.n8301 PAD.n8300 0.0380882
R45414 PAD.n8300 PAD.n4779 0.0380882
R45415 PAD.n8293 PAD.n4779 0.0380882
R45416 PAD.n8293 PAD.n8292 0.0380882
R45417 PAD.n8292 PAD.n8291 0.0380882
R45418 PAD.n8291 PAD.n4784 0.0380882
R45419 PAD.n8284 PAD.n4784 0.0380882
R45420 PAD.n8284 PAD.n8283 0.0380882
R45421 PAD.n8283 PAD.n8282 0.0380882
R45422 PAD.n8282 PAD.n4789 0.0380882
R45423 PAD.n8275 PAD.n4789 0.0380882
R45424 PAD.n8275 PAD.n8274 0.0380882
R45425 PAD.n8274 PAD.n8273 0.0380882
R45426 PAD.n8273 PAD.n4794 0.0380882
R45427 PAD.n8266 PAD.n4794 0.0380882
R45428 PAD.n8266 PAD.n8265 0.0380882
R45429 PAD.n8265 PAD.n8264 0.0380882
R45430 PAD.n8264 PAD.n4799 0.0380882
R45431 PAD.n8257 PAD.n4799 0.0380882
R45432 PAD.n8257 PAD.n8256 0.0380882
R45433 PAD.n8256 PAD.n8255 0.0380882
R45434 PAD.n8255 PAD.n4804 0.0380882
R45435 PAD.n8248 PAD.n4804 0.0380882
R45436 PAD.n8248 PAD.n8247 0.0380882
R45437 PAD.n8247 PAD.n8246 0.0380882
R45438 PAD.n8246 PAD.n4809 0.0380882
R45439 PAD.n8239 PAD.n4809 0.0380882
R45440 PAD.n8239 PAD.n8238 0.0380882
R45441 PAD.n8238 PAD.n8237 0.0380882
R45442 PAD.n8237 PAD.n4814 0.0380882
R45443 PAD.n8230 PAD.n4814 0.0380882
R45444 PAD.n8230 PAD.n8229 0.0380882
R45445 PAD.n8229 PAD.n8228 0.0380882
R45446 PAD.n8228 PAD.n4819 0.0380882
R45447 PAD.n8221 PAD.n4819 0.0380882
R45448 PAD.n8221 PAD.n8220 0.0380882
R45449 PAD.n8220 PAD.n8219 0.0380882
R45450 PAD.n8219 PAD.n4824 0.0380882
R45451 PAD.n8212 PAD.n4824 0.0380882
R45452 PAD.n8212 PAD.n8211 0.0380882
R45453 PAD.n8211 PAD.n8210 0.0380882
R45454 PAD.n5178 PAD.n5177 0.0380882
R45455 PAD.n5177 PAD.n4848 0.0380882
R45456 PAD.n5171 PAD.n4848 0.0380882
R45457 PAD.n5171 PAD.n4851 0.0380882
R45458 PAD.n5167 PAD.n4851 0.0380882
R45459 PAD.n5167 PAD.n4854 0.0380882
R45460 PAD.n5159 PAD.n4854 0.0380882
R45461 PAD.n5159 PAD.n4856 0.0380882
R45462 PAD.n5155 PAD.n4856 0.0380882
R45463 PAD.n5155 PAD.n4858 0.0380882
R45464 PAD.n5147 PAD.n4858 0.0380882
R45465 PAD.n5147 PAD.n4860 0.0380882
R45466 PAD.n5143 PAD.n4860 0.0380882
R45467 PAD.n5143 PAD.n4862 0.0380882
R45468 PAD.n5135 PAD.n4862 0.0380882
R45469 PAD.n5135 PAD.n4864 0.0380882
R45470 PAD.n5131 PAD.n4864 0.0380882
R45471 PAD.n5131 PAD.n4866 0.0380882
R45472 PAD.n5123 PAD.n4866 0.0380882
R45473 PAD.n5123 PAD.n4868 0.0380882
R45474 PAD.n5119 PAD.n4868 0.0380882
R45475 PAD.n5119 PAD.n4870 0.0380882
R45476 PAD.n5111 PAD.n4870 0.0380882
R45477 PAD.n5111 PAD.n4872 0.0380882
R45478 PAD.n5107 PAD.n4872 0.0380882
R45479 PAD.n5107 PAD.n4874 0.0380882
R45480 PAD.n5099 PAD.n4874 0.0380882
R45481 PAD.n5099 PAD.n4876 0.0380882
R45482 PAD.n5095 PAD.n4876 0.0380882
R45483 PAD.n5095 PAD.n4878 0.0380882
R45484 PAD.n5087 PAD.n4878 0.0380882
R45485 PAD.n5087 PAD.n4880 0.0380882
R45486 PAD.n5083 PAD.n4880 0.0380882
R45487 PAD.n5083 PAD.n4882 0.0380882
R45488 PAD.n5075 PAD.n4882 0.0380882
R45489 PAD.n5075 PAD.n4884 0.0380882
R45490 PAD.n5071 PAD.n4884 0.0380882
R45491 PAD.n5071 PAD.n4886 0.0380882
R45492 PAD.n5063 PAD.n4886 0.0380882
R45493 PAD.n5063 PAD.n4888 0.0380882
R45494 PAD.n5059 PAD.n4888 0.0380882
R45495 PAD.n5059 PAD.n4890 0.0380882
R45496 PAD.n5051 PAD.n4890 0.0380882
R45497 PAD.n5051 PAD.n4892 0.0380882
R45498 PAD.n5047 PAD.n4892 0.0380882
R45499 PAD.n5047 PAD.n4894 0.0380882
R45500 PAD.n5039 PAD.n4894 0.0380882
R45501 PAD.n5039 PAD.n4896 0.0380882
R45502 PAD.n5035 PAD.n4896 0.0380882
R45503 PAD.n5035 PAD.n4898 0.0380882
R45504 PAD.n5027 PAD.n4898 0.0380882
R45505 PAD.n5027 PAD.n4900 0.0380882
R45506 PAD.n5023 PAD.n4900 0.0380882
R45507 PAD.n5023 PAD.n4902 0.0380882
R45508 PAD.n5015 PAD.n4902 0.0380882
R45509 PAD.n5015 PAD.n4904 0.0380882
R45510 PAD.n5011 PAD.n4904 0.0380882
R45511 PAD.n5011 PAD.n4906 0.0380882
R45512 PAD.n5003 PAD.n4906 0.0380882
R45513 PAD.n5003 PAD.n4908 0.0380882
R45514 PAD.n4999 PAD.n4908 0.0380882
R45515 PAD.n4999 PAD.n4910 0.0380882
R45516 PAD.n4991 PAD.n4910 0.0380882
R45517 PAD.n4991 PAD.n4912 0.0380882
R45518 PAD.n4987 PAD.n4912 0.0380882
R45519 PAD.n4987 PAD.n4914 0.0380882
R45520 PAD.n4979 PAD.n4914 0.0380882
R45521 PAD.n4979 PAD.n4916 0.0380882
R45522 PAD.n4975 PAD.n4916 0.0380882
R45523 PAD.n4975 PAD.n4918 0.0380882
R45524 PAD.n4967 PAD.n4918 0.0380882
R45525 PAD.n4967 PAD.n4920 0.0380882
R45526 PAD.n4963 PAD.n4920 0.0380882
R45527 PAD.n4963 PAD.n4922 0.0380882
R45528 PAD.n4955 PAD.n4922 0.0380882
R45529 PAD.n4955 PAD.n4924 0.0380882
R45530 PAD.n4951 PAD.n4924 0.0380882
R45531 PAD.n4951 PAD.n4926 0.0380882
R45532 PAD.n4943 PAD.n4926 0.0380882
R45533 PAD.n4943 PAD.n4928 0.0380882
R45534 PAD.n4939 PAD.n4928 0.0380882
R45535 PAD.n4939 PAD.n4930 0.0380882
R45536 PAD.n4931 PAD.n4930 0.0380882
R45537 PAD.n5179 PAD.n4846 0.0380882
R45538 PAD.n4852 PAD.n4846 0.0380882
R45539 PAD.n5170 PAD.n4852 0.0380882
R45540 PAD.n5170 PAD.n5169 0.0380882
R45541 PAD.n5169 PAD.n5168 0.0380882
R45542 PAD.n5168 PAD.n4853 0.0380882
R45543 PAD.n5158 PAD.n4853 0.0380882
R45544 PAD.n5158 PAD.n5157 0.0380882
R45545 PAD.n5157 PAD.n5156 0.0380882
R45546 PAD.n5156 PAD.n4857 0.0380882
R45547 PAD.n5146 PAD.n4857 0.0380882
R45548 PAD.n5146 PAD.n5145 0.0380882
R45549 PAD.n5145 PAD.n5144 0.0380882
R45550 PAD.n5144 PAD.n4861 0.0380882
R45551 PAD.n5134 PAD.n4861 0.0380882
R45552 PAD.n5134 PAD.n5133 0.0380882
R45553 PAD.n5133 PAD.n5132 0.0380882
R45554 PAD.n5132 PAD.n4865 0.0380882
R45555 PAD.n5122 PAD.n4865 0.0380882
R45556 PAD.n5122 PAD.n5121 0.0380882
R45557 PAD.n5121 PAD.n5120 0.0380882
R45558 PAD.n5120 PAD.n4869 0.0380882
R45559 PAD.n5110 PAD.n4869 0.0380882
R45560 PAD.n5110 PAD.n5109 0.0380882
R45561 PAD.n5109 PAD.n5108 0.0380882
R45562 PAD.n5108 PAD.n4873 0.0380882
R45563 PAD.n5098 PAD.n4873 0.0380882
R45564 PAD.n5098 PAD.n5097 0.0380882
R45565 PAD.n5097 PAD.n5096 0.0380882
R45566 PAD.n5096 PAD.n4877 0.0380882
R45567 PAD.n5086 PAD.n4877 0.0380882
R45568 PAD.n5086 PAD.n5085 0.0380882
R45569 PAD.n5085 PAD.n5084 0.0380882
R45570 PAD.n5084 PAD.n4881 0.0380882
R45571 PAD.n5074 PAD.n4881 0.0380882
R45572 PAD.n5074 PAD.n5073 0.0380882
R45573 PAD.n5073 PAD.n5072 0.0380882
R45574 PAD.n5072 PAD.n4885 0.0380882
R45575 PAD.n5062 PAD.n4885 0.0380882
R45576 PAD.n5062 PAD.n5061 0.0380882
R45577 PAD.n5061 PAD.n5060 0.0380882
R45578 PAD.n5060 PAD.n4889 0.0380882
R45579 PAD.n5050 PAD.n4889 0.0380882
R45580 PAD.n5050 PAD.n5049 0.0380882
R45581 PAD.n5049 PAD.n5048 0.0380882
R45582 PAD.n5048 PAD.n4893 0.0380882
R45583 PAD.n5038 PAD.n4893 0.0380882
R45584 PAD.n5038 PAD.n5037 0.0380882
R45585 PAD.n5037 PAD.n5036 0.0380882
R45586 PAD.n5036 PAD.n4897 0.0380882
R45587 PAD.n5026 PAD.n4897 0.0380882
R45588 PAD.n5026 PAD.n5025 0.0380882
R45589 PAD.n5025 PAD.n5024 0.0380882
R45590 PAD.n5024 PAD.n4901 0.0380882
R45591 PAD.n5014 PAD.n4901 0.0380882
R45592 PAD.n5014 PAD.n5013 0.0380882
R45593 PAD.n5013 PAD.n5012 0.0380882
R45594 PAD.n5012 PAD.n4905 0.0380882
R45595 PAD.n5002 PAD.n4905 0.0380882
R45596 PAD.n5002 PAD.n5001 0.0380882
R45597 PAD.n5001 PAD.n5000 0.0380882
R45598 PAD.n5000 PAD.n4909 0.0380882
R45599 PAD.n4990 PAD.n4909 0.0380882
R45600 PAD.n4990 PAD.n4989 0.0380882
R45601 PAD.n4989 PAD.n4988 0.0380882
R45602 PAD.n4988 PAD.n4913 0.0380882
R45603 PAD.n4978 PAD.n4913 0.0380882
R45604 PAD.n4978 PAD.n4977 0.0380882
R45605 PAD.n4977 PAD.n4976 0.0380882
R45606 PAD.n4976 PAD.n4917 0.0380882
R45607 PAD.n4966 PAD.n4917 0.0380882
R45608 PAD.n4966 PAD.n4965 0.0380882
R45609 PAD.n4965 PAD.n4964 0.0380882
R45610 PAD.n4964 PAD.n4921 0.0380882
R45611 PAD.n4954 PAD.n4921 0.0380882
R45612 PAD.n4954 PAD.n4953 0.0380882
R45613 PAD.n4953 PAD.n4952 0.0380882
R45614 PAD.n4952 PAD.n4925 0.0380882
R45615 PAD.n4942 PAD.n4925 0.0380882
R45616 PAD.n4942 PAD.n4941 0.0380882
R45617 PAD.n4941 PAD.n4940 0.0380882
R45618 PAD.n4940 PAD.n4929 0.0380882
R45619 PAD.n4929 PAD.n4835 0.0380882
R45620 PAD.n8160 PAD.n8159 0.0380882
R45621 PAD.n8159 PAD.n7874 0.0380882
R45622 PAD.n8155 PAD.n7874 0.0380882
R45623 PAD.n8155 PAD.n8151 0.0380882
R45624 PAD.n8151 PAD.n8150 0.0380882
R45625 PAD.n8150 PAD.n7876 0.0380882
R45626 PAD.n8146 PAD.n7876 0.0380882
R45627 PAD.n8146 PAD.n8142 0.0380882
R45628 PAD.n8142 PAD.n8141 0.0380882
R45629 PAD.n8141 PAD.n7881 0.0380882
R45630 PAD.n8137 PAD.n7881 0.0380882
R45631 PAD.n8137 PAD.n8133 0.0380882
R45632 PAD.n8133 PAD.n8132 0.0380882
R45633 PAD.n8132 PAD.n7886 0.0380882
R45634 PAD.n8128 PAD.n7886 0.0380882
R45635 PAD.n8128 PAD.n8124 0.0380882
R45636 PAD.n8124 PAD.n8123 0.0380882
R45637 PAD.n8123 PAD.n7891 0.0380882
R45638 PAD.n8119 PAD.n7891 0.0380882
R45639 PAD.n8119 PAD.n8115 0.0380882
R45640 PAD.n8115 PAD.n8114 0.0380882
R45641 PAD.n8114 PAD.n7896 0.0380882
R45642 PAD.n8110 PAD.n7896 0.0380882
R45643 PAD.n8110 PAD.n8106 0.0380882
R45644 PAD.n8106 PAD.n8105 0.0380882
R45645 PAD.n8105 PAD.n7901 0.0380882
R45646 PAD.n8101 PAD.n7901 0.0380882
R45647 PAD.n8101 PAD.n8097 0.0380882
R45648 PAD.n8097 PAD.n8096 0.0380882
R45649 PAD.n8096 PAD.n7906 0.0380882
R45650 PAD.n8092 PAD.n7906 0.0380882
R45651 PAD.n8092 PAD.n8088 0.0380882
R45652 PAD.n8088 PAD.n8087 0.0380882
R45653 PAD.n8087 PAD.n7911 0.0380882
R45654 PAD.n8083 PAD.n7911 0.0380882
R45655 PAD.n8083 PAD.n8079 0.0380882
R45656 PAD.n8079 PAD.n8078 0.0380882
R45657 PAD.n8078 PAD.n7916 0.0380882
R45658 PAD.n8074 PAD.n7916 0.0380882
R45659 PAD.n8074 PAD.n8070 0.0380882
R45660 PAD.n8070 PAD.n8069 0.0380882
R45661 PAD.n8069 PAD.n7921 0.0380882
R45662 PAD.n8065 PAD.n7921 0.0380882
R45663 PAD.n8065 PAD.n8061 0.0380882
R45664 PAD.n8061 PAD.n8060 0.0380882
R45665 PAD.n8060 PAD.n7926 0.0380882
R45666 PAD.n8056 PAD.n7926 0.0380882
R45667 PAD.n8056 PAD.n8052 0.0380882
R45668 PAD.n8052 PAD.n8051 0.0380882
R45669 PAD.n8051 PAD.n7931 0.0380882
R45670 PAD.n8047 PAD.n7931 0.0380882
R45671 PAD.n8047 PAD.n8043 0.0380882
R45672 PAD.n8043 PAD.n8042 0.0380882
R45673 PAD.n8042 PAD.n7936 0.0380882
R45674 PAD.n8038 PAD.n7936 0.0380882
R45675 PAD.n8038 PAD.n8034 0.0380882
R45676 PAD.n8034 PAD.n8033 0.0380882
R45677 PAD.n8033 PAD.n7941 0.0380882
R45678 PAD.n8029 PAD.n7941 0.0380882
R45679 PAD.n8029 PAD.n8025 0.0380882
R45680 PAD.n8025 PAD.n8024 0.0380882
R45681 PAD.n8024 PAD.n7946 0.0380882
R45682 PAD.n8020 PAD.n7946 0.0380882
R45683 PAD.n8020 PAD.n8016 0.0380882
R45684 PAD.n8016 PAD.n8015 0.0380882
R45685 PAD.n8015 PAD.n7951 0.0380882
R45686 PAD.n8011 PAD.n7951 0.0380882
R45687 PAD.n8011 PAD.n8007 0.0380882
R45688 PAD.n8007 PAD.n8006 0.0380882
R45689 PAD.n8006 PAD.n7956 0.0380882
R45690 PAD.n8002 PAD.n7956 0.0380882
R45691 PAD.n8002 PAD.n7998 0.0380882
R45692 PAD.n7998 PAD.n7997 0.0380882
R45693 PAD.n7997 PAD.n7961 0.0380882
R45694 PAD.n7993 PAD.n7961 0.0380882
R45695 PAD.n7993 PAD.n7989 0.0380882
R45696 PAD.n7989 PAD.n7988 0.0380882
R45697 PAD.n7988 PAD.n7966 0.0380882
R45698 PAD.n7984 PAD.n7966 0.0380882
R45699 PAD.n7984 PAD.n7980 0.0380882
R45700 PAD.n7980 PAD.n7979 0.0380882
R45701 PAD.n7979 PAD.n7973 0.0380882
R45702 PAD.n7973 PAD.n7972 0.0380882
R45703 PAD.n8158 PAD.n5193 0.0380882
R45704 PAD.n8158 PAD.n8157 0.0380882
R45705 PAD.n8157 PAD.n8156 0.0380882
R45706 PAD.n8156 PAD.n7875 0.0380882
R45707 PAD.n8149 PAD.n7875 0.0380882
R45708 PAD.n8149 PAD.n8148 0.0380882
R45709 PAD.n8148 PAD.n8147 0.0380882
R45710 PAD.n8147 PAD.n7880 0.0380882
R45711 PAD.n8140 PAD.n7880 0.0380882
R45712 PAD.n8140 PAD.n8139 0.0380882
R45713 PAD.n8139 PAD.n8138 0.0380882
R45714 PAD.n8138 PAD.n7885 0.0380882
R45715 PAD.n8131 PAD.n7885 0.0380882
R45716 PAD.n8131 PAD.n8130 0.0380882
R45717 PAD.n8130 PAD.n8129 0.0380882
R45718 PAD.n8129 PAD.n7890 0.0380882
R45719 PAD.n8122 PAD.n7890 0.0380882
R45720 PAD.n8122 PAD.n8121 0.0380882
R45721 PAD.n8121 PAD.n8120 0.0380882
R45722 PAD.n8120 PAD.n7895 0.0380882
R45723 PAD.n8113 PAD.n7895 0.0380882
R45724 PAD.n8113 PAD.n8112 0.0380882
R45725 PAD.n8112 PAD.n8111 0.0380882
R45726 PAD.n8111 PAD.n7900 0.0380882
R45727 PAD.n8104 PAD.n7900 0.0380882
R45728 PAD.n8104 PAD.n8103 0.0380882
R45729 PAD.n8103 PAD.n8102 0.0380882
R45730 PAD.n8102 PAD.n7905 0.0380882
R45731 PAD.n8095 PAD.n7905 0.0380882
R45732 PAD.n8095 PAD.n8094 0.0380882
R45733 PAD.n8094 PAD.n8093 0.0380882
R45734 PAD.n8093 PAD.n7910 0.0380882
R45735 PAD.n8086 PAD.n7910 0.0380882
R45736 PAD.n8086 PAD.n8085 0.0380882
R45737 PAD.n8085 PAD.n8084 0.0380882
R45738 PAD.n8084 PAD.n7915 0.0380882
R45739 PAD.n8077 PAD.n7915 0.0380882
R45740 PAD.n8077 PAD.n8076 0.0380882
R45741 PAD.n8076 PAD.n8075 0.0380882
R45742 PAD.n8075 PAD.n7920 0.0380882
R45743 PAD.n8068 PAD.n7920 0.0380882
R45744 PAD.n8068 PAD.n8067 0.0380882
R45745 PAD.n8067 PAD.n8066 0.0380882
R45746 PAD.n8066 PAD.n7925 0.0380882
R45747 PAD.n8059 PAD.n7925 0.0380882
R45748 PAD.n8059 PAD.n8058 0.0380882
R45749 PAD.n8058 PAD.n8057 0.0380882
R45750 PAD.n8057 PAD.n7930 0.0380882
R45751 PAD.n8050 PAD.n7930 0.0380882
R45752 PAD.n8050 PAD.n8049 0.0380882
R45753 PAD.n8049 PAD.n8048 0.0380882
R45754 PAD.n8048 PAD.n7935 0.0380882
R45755 PAD.n8041 PAD.n7935 0.0380882
R45756 PAD.n8041 PAD.n8040 0.0380882
R45757 PAD.n8040 PAD.n8039 0.0380882
R45758 PAD.n8039 PAD.n7940 0.0380882
R45759 PAD.n8032 PAD.n7940 0.0380882
R45760 PAD.n8032 PAD.n8031 0.0380882
R45761 PAD.n8031 PAD.n8030 0.0380882
R45762 PAD.n8030 PAD.n7945 0.0380882
R45763 PAD.n8023 PAD.n7945 0.0380882
R45764 PAD.n8023 PAD.n8022 0.0380882
R45765 PAD.n8022 PAD.n8021 0.0380882
R45766 PAD.n8021 PAD.n7950 0.0380882
R45767 PAD.n8014 PAD.n7950 0.0380882
R45768 PAD.n8014 PAD.n8013 0.0380882
R45769 PAD.n8013 PAD.n8012 0.0380882
R45770 PAD.n8012 PAD.n7955 0.0380882
R45771 PAD.n8005 PAD.n7955 0.0380882
R45772 PAD.n8005 PAD.n8004 0.0380882
R45773 PAD.n8004 PAD.n8003 0.0380882
R45774 PAD.n8003 PAD.n7960 0.0380882
R45775 PAD.n7996 PAD.n7960 0.0380882
R45776 PAD.n7996 PAD.n7995 0.0380882
R45777 PAD.n7995 PAD.n7994 0.0380882
R45778 PAD.n7994 PAD.n7965 0.0380882
R45779 PAD.n7987 PAD.n7965 0.0380882
R45780 PAD.n7987 PAD.n7986 0.0380882
R45781 PAD.n7986 PAD.n7985 0.0380882
R45782 PAD.n7985 PAD.n7970 0.0380882
R45783 PAD.n7978 PAD.n7970 0.0380882
R45784 PAD.n7978 PAD.n7977 0.0380882
R45785 PAD.n7977 PAD.n5186 0.0380882
R45786 PAD.n5542 PAD.n5541 0.0380882
R45787 PAD.n5541 PAD.n5212 0.0380882
R45788 PAD.n5535 PAD.n5212 0.0380882
R45789 PAD.n5535 PAD.n5215 0.0380882
R45790 PAD.n5531 PAD.n5215 0.0380882
R45791 PAD.n5531 PAD.n5218 0.0380882
R45792 PAD.n5523 PAD.n5218 0.0380882
R45793 PAD.n5523 PAD.n5220 0.0380882
R45794 PAD.n5519 PAD.n5220 0.0380882
R45795 PAD.n5519 PAD.n5222 0.0380882
R45796 PAD.n5511 PAD.n5222 0.0380882
R45797 PAD.n5511 PAD.n5224 0.0380882
R45798 PAD.n5507 PAD.n5224 0.0380882
R45799 PAD.n5507 PAD.n5226 0.0380882
R45800 PAD.n5499 PAD.n5226 0.0380882
R45801 PAD.n5499 PAD.n5228 0.0380882
R45802 PAD.n5495 PAD.n5228 0.0380882
R45803 PAD.n5495 PAD.n5230 0.0380882
R45804 PAD.n5487 PAD.n5230 0.0380882
R45805 PAD.n5487 PAD.n5232 0.0380882
R45806 PAD.n5483 PAD.n5232 0.0380882
R45807 PAD.n5483 PAD.n5234 0.0380882
R45808 PAD.n5475 PAD.n5234 0.0380882
R45809 PAD.n5475 PAD.n5236 0.0380882
R45810 PAD.n5471 PAD.n5236 0.0380882
R45811 PAD.n5471 PAD.n5238 0.0380882
R45812 PAD.n5463 PAD.n5238 0.0380882
R45813 PAD.n5463 PAD.n5240 0.0380882
R45814 PAD.n5459 PAD.n5240 0.0380882
R45815 PAD.n5459 PAD.n5242 0.0380882
R45816 PAD.n5451 PAD.n5242 0.0380882
R45817 PAD.n5451 PAD.n5244 0.0380882
R45818 PAD.n5447 PAD.n5244 0.0380882
R45819 PAD.n5447 PAD.n5246 0.0380882
R45820 PAD.n5439 PAD.n5246 0.0380882
R45821 PAD.n5439 PAD.n5248 0.0380882
R45822 PAD.n5435 PAD.n5248 0.0380882
R45823 PAD.n5435 PAD.n5250 0.0380882
R45824 PAD.n5427 PAD.n5250 0.0380882
R45825 PAD.n5427 PAD.n5252 0.0380882
R45826 PAD.n5423 PAD.n5252 0.0380882
R45827 PAD.n5423 PAD.n5254 0.0380882
R45828 PAD.n5415 PAD.n5254 0.0380882
R45829 PAD.n5415 PAD.n5256 0.0380882
R45830 PAD.n5411 PAD.n5256 0.0380882
R45831 PAD.n5411 PAD.n5258 0.0380882
R45832 PAD.n5403 PAD.n5258 0.0380882
R45833 PAD.n5403 PAD.n5260 0.0380882
R45834 PAD.n5399 PAD.n5260 0.0380882
R45835 PAD.n5399 PAD.n5262 0.0380882
R45836 PAD.n5391 PAD.n5262 0.0380882
R45837 PAD.n5391 PAD.n5264 0.0380882
R45838 PAD.n5387 PAD.n5264 0.0380882
R45839 PAD.n5387 PAD.n5266 0.0380882
R45840 PAD.n5379 PAD.n5266 0.0380882
R45841 PAD.n5379 PAD.n5268 0.0380882
R45842 PAD.n5375 PAD.n5268 0.0380882
R45843 PAD.n5375 PAD.n5270 0.0380882
R45844 PAD.n5367 PAD.n5270 0.0380882
R45845 PAD.n5367 PAD.n5272 0.0380882
R45846 PAD.n5363 PAD.n5272 0.0380882
R45847 PAD.n5363 PAD.n5274 0.0380882
R45848 PAD.n5355 PAD.n5274 0.0380882
R45849 PAD.n5355 PAD.n5276 0.0380882
R45850 PAD.n5351 PAD.n5276 0.0380882
R45851 PAD.n5351 PAD.n5278 0.0380882
R45852 PAD.n5343 PAD.n5278 0.0380882
R45853 PAD.n5343 PAD.n5280 0.0380882
R45854 PAD.n5339 PAD.n5280 0.0380882
R45855 PAD.n5339 PAD.n5282 0.0380882
R45856 PAD.n5331 PAD.n5282 0.0380882
R45857 PAD.n5331 PAD.n5284 0.0380882
R45858 PAD.n5327 PAD.n5284 0.0380882
R45859 PAD.n5327 PAD.n5286 0.0380882
R45860 PAD.n5319 PAD.n5286 0.0380882
R45861 PAD.n5319 PAD.n5288 0.0380882
R45862 PAD.n5315 PAD.n5288 0.0380882
R45863 PAD.n5315 PAD.n5290 0.0380882
R45864 PAD.n5307 PAD.n5290 0.0380882
R45865 PAD.n5307 PAD.n5292 0.0380882
R45866 PAD.n5303 PAD.n5292 0.0380882
R45867 PAD.n5303 PAD.n5294 0.0380882
R45868 PAD.n5295 PAD.n5294 0.0380882
R45869 PAD.n5543 PAD.n5210 0.0380882
R45870 PAD.n5216 PAD.n5210 0.0380882
R45871 PAD.n5534 PAD.n5216 0.0380882
R45872 PAD.n5534 PAD.n5533 0.0380882
R45873 PAD.n5533 PAD.n5532 0.0380882
R45874 PAD.n5532 PAD.n5217 0.0380882
R45875 PAD.n5522 PAD.n5217 0.0380882
R45876 PAD.n5522 PAD.n5521 0.0380882
R45877 PAD.n5521 PAD.n5520 0.0380882
R45878 PAD.n5520 PAD.n5221 0.0380882
R45879 PAD.n5510 PAD.n5221 0.0380882
R45880 PAD.n5510 PAD.n5509 0.0380882
R45881 PAD.n5509 PAD.n5508 0.0380882
R45882 PAD.n5508 PAD.n5225 0.0380882
R45883 PAD.n5498 PAD.n5225 0.0380882
R45884 PAD.n5498 PAD.n5497 0.0380882
R45885 PAD.n5497 PAD.n5496 0.0380882
R45886 PAD.n5496 PAD.n5229 0.0380882
R45887 PAD.n5486 PAD.n5229 0.0380882
R45888 PAD.n5486 PAD.n5485 0.0380882
R45889 PAD.n5485 PAD.n5484 0.0380882
R45890 PAD.n5484 PAD.n5233 0.0380882
R45891 PAD.n5474 PAD.n5233 0.0380882
R45892 PAD.n5474 PAD.n5473 0.0380882
R45893 PAD.n5473 PAD.n5472 0.0380882
R45894 PAD.n5472 PAD.n5237 0.0380882
R45895 PAD.n5462 PAD.n5237 0.0380882
R45896 PAD.n5462 PAD.n5461 0.0380882
R45897 PAD.n5461 PAD.n5460 0.0380882
R45898 PAD.n5460 PAD.n5241 0.0380882
R45899 PAD.n5450 PAD.n5241 0.0380882
R45900 PAD.n5450 PAD.n5449 0.0380882
R45901 PAD.n5449 PAD.n5448 0.0380882
R45902 PAD.n5448 PAD.n5245 0.0380882
R45903 PAD.n5438 PAD.n5245 0.0380882
R45904 PAD.n5438 PAD.n5437 0.0380882
R45905 PAD.n5437 PAD.n5436 0.0380882
R45906 PAD.n5436 PAD.n5249 0.0380882
R45907 PAD.n5426 PAD.n5249 0.0380882
R45908 PAD.n5426 PAD.n5425 0.0380882
R45909 PAD.n5425 PAD.n5424 0.0380882
R45910 PAD.n5424 PAD.n5253 0.0380882
R45911 PAD.n5414 PAD.n5253 0.0380882
R45912 PAD.n5414 PAD.n5413 0.0380882
R45913 PAD.n5413 PAD.n5412 0.0380882
R45914 PAD.n5412 PAD.n5257 0.0380882
R45915 PAD.n5402 PAD.n5257 0.0380882
R45916 PAD.n5402 PAD.n5401 0.0380882
R45917 PAD.n5401 PAD.n5400 0.0380882
R45918 PAD.n5400 PAD.n5261 0.0380882
R45919 PAD.n5390 PAD.n5261 0.0380882
R45920 PAD.n5390 PAD.n5389 0.0380882
R45921 PAD.n5389 PAD.n5388 0.0380882
R45922 PAD.n5388 PAD.n5265 0.0380882
R45923 PAD.n5378 PAD.n5265 0.0380882
R45924 PAD.n5378 PAD.n5377 0.0380882
R45925 PAD.n5377 PAD.n5376 0.0380882
R45926 PAD.n5376 PAD.n5269 0.0380882
R45927 PAD.n5366 PAD.n5269 0.0380882
R45928 PAD.n5366 PAD.n5365 0.0380882
R45929 PAD.n5365 PAD.n5364 0.0380882
R45930 PAD.n5364 PAD.n5273 0.0380882
R45931 PAD.n5354 PAD.n5273 0.0380882
R45932 PAD.n5354 PAD.n5353 0.0380882
R45933 PAD.n5353 PAD.n5352 0.0380882
R45934 PAD.n5352 PAD.n5277 0.0380882
R45935 PAD.n5342 PAD.n5277 0.0380882
R45936 PAD.n5342 PAD.n5341 0.0380882
R45937 PAD.n5341 PAD.n5340 0.0380882
R45938 PAD.n5340 PAD.n5281 0.0380882
R45939 PAD.n5330 PAD.n5281 0.0380882
R45940 PAD.n5330 PAD.n5329 0.0380882
R45941 PAD.n5329 PAD.n5328 0.0380882
R45942 PAD.n5328 PAD.n5285 0.0380882
R45943 PAD.n5318 PAD.n5285 0.0380882
R45944 PAD.n5318 PAD.n5317 0.0380882
R45945 PAD.n5317 PAD.n5316 0.0380882
R45946 PAD.n5316 PAD.n5289 0.0380882
R45947 PAD.n5306 PAD.n5289 0.0380882
R45948 PAD.n5306 PAD.n5305 0.0380882
R45949 PAD.n5305 PAD.n5304 0.0380882
R45950 PAD.n5304 PAD.n5293 0.0380882
R45951 PAD.n5293 PAD.n5200 0.0380882
R45952 PAD.n7779 PAD.n7106 0.0380882
R45953 PAD.n7775 PAD.n7106 0.0380882
R45954 PAD.n7775 PAD.n7772 0.0380882
R45955 PAD.n7772 PAD.n7768 0.0380882
R45956 PAD.n7768 PAD.n7108 0.0380882
R45957 PAD.n7764 PAD.n7108 0.0380882
R45958 PAD.n7764 PAD.n7760 0.0380882
R45959 PAD.n7760 PAD.n7756 0.0380882
R45960 PAD.n7756 PAD.n7110 0.0380882
R45961 PAD.n7752 PAD.n7110 0.0380882
R45962 PAD.n7752 PAD.n7748 0.0380882
R45963 PAD.n7748 PAD.n7744 0.0380882
R45964 PAD.n7744 PAD.n7112 0.0380882
R45965 PAD.n7740 PAD.n7112 0.0380882
R45966 PAD.n7740 PAD.n7736 0.0380882
R45967 PAD.n7736 PAD.n7732 0.0380882
R45968 PAD.n7732 PAD.n7114 0.0380882
R45969 PAD.n7728 PAD.n7114 0.0380882
R45970 PAD.n7728 PAD.n7724 0.0380882
R45971 PAD.n7724 PAD.n7720 0.0380882
R45972 PAD.n7720 PAD.n7116 0.0380882
R45973 PAD.n7716 PAD.n7116 0.0380882
R45974 PAD.n7716 PAD.n7712 0.0380882
R45975 PAD.n7712 PAD.n7708 0.0380882
R45976 PAD.n7708 PAD.n7118 0.0380882
R45977 PAD.n7704 PAD.n7118 0.0380882
R45978 PAD.n7704 PAD.n7700 0.0380882
R45979 PAD.n7700 PAD.n7696 0.0380882
R45980 PAD.n7696 PAD.n7120 0.0380882
R45981 PAD.n7692 PAD.n7120 0.0380882
R45982 PAD.n7692 PAD.n7688 0.0380882
R45983 PAD.n7688 PAD.n7684 0.0380882
R45984 PAD.n7684 PAD.n7122 0.0380882
R45985 PAD.n7680 PAD.n7122 0.0380882
R45986 PAD.n7680 PAD.n7676 0.0380882
R45987 PAD.n7676 PAD.n7672 0.0380882
R45988 PAD.n7672 PAD.n7124 0.0380882
R45989 PAD.n7668 PAD.n7124 0.0380882
R45990 PAD.n7668 PAD.n7664 0.0380882
R45991 PAD.n7664 PAD.n7660 0.0380882
R45992 PAD.n7660 PAD.n7126 0.0380882
R45993 PAD.n7656 PAD.n7126 0.0380882
R45994 PAD.n7656 PAD.n7652 0.0380882
R45995 PAD.n7652 PAD.n7648 0.0380882
R45996 PAD.n7648 PAD.n7128 0.0380882
R45997 PAD.n7644 PAD.n7128 0.0380882
R45998 PAD.n7644 PAD.n7640 0.0380882
R45999 PAD.n7640 PAD.n7636 0.0380882
R46000 PAD.n7636 PAD.n7130 0.0380882
R46001 PAD.n7632 PAD.n7130 0.0380882
R46002 PAD.n7632 PAD.n7628 0.0380882
R46003 PAD.n7628 PAD.n7624 0.0380882
R46004 PAD.n7624 PAD.n7132 0.0380882
R46005 PAD.n7620 PAD.n7132 0.0380882
R46006 PAD.n7620 PAD.n7616 0.0380882
R46007 PAD.n7616 PAD.n7612 0.0380882
R46008 PAD.n7612 PAD.n7134 0.0380882
R46009 PAD.n7608 PAD.n7134 0.0380882
R46010 PAD.n7608 PAD.n7604 0.0380882
R46011 PAD.n7604 PAD.n7600 0.0380882
R46012 PAD.n7600 PAD.n7136 0.0380882
R46013 PAD.n7596 PAD.n7136 0.0380882
R46014 PAD.n7596 PAD.n7592 0.0380882
R46015 PAD.n7592 PAD.n7588 0.0380882
R46016 PAD.n7588 PAD.n7138 0.0380882
R46017 PAD.n7584 PAD.n7138 0.0380882
R46018 PAD.n7584 PAD.n7580 0.0380882
R46019 PAD.n7580 PAD.n7576 0.0380882
R46020 PAD.n7576 PAD.n7140 0.0380882
R46021 PAD.n7572 PAD.n7140 0.0380882
R46022 PAD.n7572 PAD.n7568 0.0380882
R46023 PAD.n7568 PAD.n7564 0.0380882
R46024 PAD.n7564 PAD.n7142 0.0380882
R46025 PAD.n7560 PAD.n7142 0.0380882
R46026 PAD.n7560 PAD.n7556 0.0380882
R46027 PAD.n7556 PAD.n7552 0.0380882
R46028 PAD.n7552 PAD.n7144 0.0380882
R46029 PAD.n7548 PAD.n7144 0.0380882
R46030 PAD.n7548 PAD.n7544 0.0380882
R46031 PAD.n7544 PAD.n7540 0.0380882
R46032 PAD.n7540 PAD.n7146 0.0380882
R46033 PAD.n7536 PAD.n7146 0.0380882
R46034 PAD.n7536 PAD.n7532 0.0380882
R46035 PAD.n7778 PAD.n7777 0.0380882
R46036 PAD.n7777 PAD.n7776 0.0380882
R46037 PAD.n7776 PAD.n7107 0.0380882
R46038 PAD.n7767 PAD.n7107 0.0380882
R46039 PAD.n7767 PAD.n7766 0.0380882
R46040 PAD.n7766 PAD.n7765 0.0380882
R46041 PAD.n7765 PAD.n7109 0.0380882
R46042 PAD.n7755 PAD.n7109 0.0380882
R46043 PAD.n7755 PAD.n7754 0.0380882
R46044 PAD.n7754 PAD.n7753 0.0380882
R46045 PAD.n7753 PAD.n7111 0.0380882
R46046 PAD.n7743 PAD.n7111 0.0380882
R46047 PAD.n7743 PAD.n7742 0.0380882
R46048 PAD.n7742 PAD.n7741 0.0380882
R46049 PAD.n7741 PAD.n7113 0.0380882
R46050 PAD.n7731 PAD.n7113 0.0380882
R46051 PAD.n7731 PAD.n7730 0.0380882
R46052 PAD.n7730 PAD.n7729 0.0380882
R46053 PAD.n7729 PAD.n7115 0.0380882
R46054 PAD.n7719 PAD.n7115 0.0380882
R46055 PAD.n7719 PAD.n7718 0.0380882
R46056 PAD.n7718 PAD.n7717 0.0380882
R46057 PAD.n7717 PAD.n7117 0.0380882
R46058 PAD.n7707 PAD.n7117 0.0380882
R46059 PAD.n7707 PAD.n7706 0.0380882
R46060 PAD.n7706 PAD.n7705 0.0380882
R46061 PAD.n7705 PAD.n7119 0.0380882
R46062 PAD.n7695 PAD.n7119 0.0380882
R46063 PAD.n7695 PAD.n7694 0.0380882
R46064 PAD.n7694 PAD.n7693 0.0380882
R46065 PAD.n7693 PAD.n7121 0.0380882
R46066 PAD.n7683 PAD.n7121 0.0380882
R46067 PAD.n7683 PAD.n7682 0.0380882
R46068 PAD.n7682 PAD.n7681 0.0380882
R46069 PAD.n7681 PAD.n7123 0.0380882
R46070 PAD.n7671 PAD.n7123 0.0380882
R46071 PAD.n7671 PAD.n7670 0.0380882
R46072 PAD.n7670 PAD.n7669 0.0380882
R46073 PAD.n7669 PAD.n7125 0.0380882
R46074 PAD.n7659 PAD.n7125 0.0380882
R46075 PAD.n7659 PAD.n7658 0.0380882
R46076 PAD.n7658 PAD.n7657 0.0380882
R46077 PAD.n7657 PAD.n7127 0.0380882
R46078 PAD.n7647 PAD.n7127 0.0380882
R46079 PAD.n7647 PAD.n7646 0.0380882
R46080 PAD.n7646 PAD.n7645 0.0380882
R46081 PAD.n7645 PAD.n7129 0.0380882
R46082 PAD.n7635 PAD.n7129 0.0380882
R46083 PAD.n7635 PAD.n7634 0.0380882
R46084 PAD.n7634 PAD.n7633 0.0380882
R46085 PAD.n7633 PAD.n7131 0.0380882
R46086 PAD.n7623 PAD.n7131 0.0380882
R46087 PAD.n7623 PAD.n7622 0.0380882
R46088 PAD.n7622 PAD.n7621 0.0380882
R46089 PAD.n7621 PAD.n7133 0.0380882
R46090 PAD.n7611 PAD.n7133 0.0380882
R46091 PAD.n7611 PAD.n7610 0.0380882
R46092 PAD.n7610 PAD.n7609 0.0380882
R46093 PAD.n7609 PAD.n7135 0.0380882
R46094 PAD.n7599 PAD.n7135 0.0380882
R46095 PAD.n7599 PAD.n7598 0.0380882
R46096 PAD.n7598 PAD.n7597 0.0380882
R46097 PAD.n7597 PAD.n7137 0.0380882
R46098 PAD.n7587 PAD.n7137 0.0380882
R46099 PAD.n7587 PAD.n7586 0.0380882
R46100 PAD.n7586 PAD.n7585 0.0380882
R46101 PAD.n7585 PAD.n7139 0.0380882
R46102 PAD.n7575 PAD.n7139 0.0380882
R46103 PAD.n7575 PAD.n7574 0.0380882
R46104 PAD.n7574 PAD.n7573 0.0380882
R46105 PAD.n7573 PAD.n7141 0.0380882
R46106 PAD.n7563 PAD.n7141 0.0380882
R46107 PAD.n7563 PAD.n7562 0.0380882
R46108 PAD.n7562 PAD.n7561 0.0380882
R46109 PAD.n7561 PAD.n7143 0.0380882
R46110 PAD.n7551 PAD.n7143 0.0380882
R46111 PAD.n7551 PAD.n7550 0.0380882
R46112 PAD.n7550 PAD.n7549 0.0380882
R46113 PAD.n7549 PAD.n7145 0.0380882
R46114 PAD.n7539 PAD.n7145 0.0380882
R46115 PAD.n7539 PAD.n7538 0.0380882
R46116 PAD.n7538 PAD.n7537 0.0380882
R46117 PAD.n7537 PAD.n7147 0.0380882
R46118 PAD.n7050 PAD.n7049 0.0380882
R46119 PAD.n7049 PAD.n6720 0.0380882
R46120 PAD.n7043 PAD.n6720 0.0380882
R46121 PAD.n7043 PAD.n6723 0.0380882
R46122 PAD.n7039 PAD.n6723 0.0380882
R46123 PAD.n7039 PAD.n6726 0.0380882
R46124 PAD.n7031 PAD.n6726 0.0380882
R46125 PAD.n7031 PAD.n6728 0.0380882
R46126 PAD.n7027 PAD.n6728 0.0380882
R46127 PAD.n7027 PAD.n6730 0.0380882
R46128 PAD.n7019 PAD.n6730 0.0380882
R46129 PAD.n7019 PAD.n6732 0.0380882
R46130 PAD.n7015 PAD.n6732 0.0380882
R46131 PAD.n7015 PAD.n6734 0.0380882
R46132 PAD.n7007 PAD.n6734 0.0380882
R46133 PAD.n7007 PAD.n6736 0.0380882
R46134 PAD.n7003 PAD.n6736 0.0380882
R46135 PAD.n7003 PAD.n6738 0.0380882
R46136 PAD.n6995 PAD.n6738 0.0380882
R46137 PAD.n6995 PAD.n6740 0.0380882
R46138 PAD.n6991 PAD.n6740 0.0380882
R46139 PAD.n6991 PAD.n6742 0.0380882
R46140 PAD.n6983 PAD.n6742 0.0380882
R46141 PAD.n6983 PAD.n6744 0.0380882
R46142 PAD.n6979 PAD.n6744 0.0380882
R46143 PAD.n6979 PAD.n6746 0.0380882
R46144 PAD.n6971 PAD.n6746 0.0380882
R46145 PAD.n6971 PAD.n6748 0.0380882
R46146 PAD.n6967 PAD.n6748 0.0380882
R46147 PAD.n6967 PAD.n6750 0.0380882
R46148 PAD.n6959 PAD.n6750 0.0380882
R46149 PAD.n6959 PAD.n6752 0.0380882
R46150 PAD.n6955 PAD.n6752 0.0380882
R46151 PAD.n6955 PAD.n6754 0.0380882
R46152 PAD.n6947 PAD.n6754 0.0380882
R46153 PAD.n6947 PAD.n6756 0.0380882
R46154 PAD.n6943 PAD.n6756 0.0380882
R46155 PAD.n6943 PAD.n6758 0.0380882
R46156 PAD.n6935 PAD.n6758 0.0380882
R46157 PAD.n6935 PAD.n6760 0.0380882
R46158 PAD.n6931 PAD.n6760 0.0380882
R46159 PAD.n6931 PAD.n6762 0.0380882
R46160 PAD.n6923 PAD.n6762 0.0380882
R46161 PAD.n6923 PAD.n6764 0.0380882
R46162 PAD.n6919 PAD.n6764 0.0380882
R46163 PAD.n6919 PAD.n6766 0.0380882
R46164 PAD.n6911 PAD.n6766 0.0380882
R46165 PAD.n6911 PAD.n6768 0.0380882
R46166 PAD.n6907 PAD.n6768 0.0380882
R46167 PAD.n6907 PAD.n6770 0.0380882
R46168 PAD.n6899 PAD.n6770 0.0380882
R46169 PAD.n6899 PAD.n6772 0.0380882
R46170 PAD.n6895 PAD.n6772 0.0380882
R46171 PAD.n6895 PAD.n6774 0.0380882
R46172 PAD.n6887 PAD.n6774 0.0380882
R46173 PAD.n6887 PAD.n6776 0.0380882
R46174 PAD.n6883 PAD.n6776 0.0380882
R46175 PAD.n6883 PAD.n6778 0.0380882
R46176 PAD.n6875 PAD.n6778 0.0380882
R46177 PAD.n6875 PAD.n6780 0.0380882
R46178 PAD.n6871 PAD.n6780 0.0380882
R46179 PAD.n6871 PAD.n6782 0.0380882
R46180 PAD.n6863 PAD.n6782 0.0380882
R46181 PAD.n6863 PAD.n6784 0.0380882
R46182 PAD.n6859 PAD.n6784 0.0380882
R46183 PAD.n6859 PAD.n6786 0.0380882
R46184 PAD.n6851 PAD.n6786 0.0380882
R46185 PAD.n6851 PAD.n6788 0.0380882
R46186 PAD.n6847 PAD.n6788 0.0380882
R46187 PAD.n6847 PAD.n6790 0.0380882
R46188 PAD.n6839 PAD.n6790 0.0380882
R46189 PAD.n6839 PAD.n6792 0.0380882
R46190 PAD.n6835 PAD.n6792 0.0380882
R46191 PAD.n6835 PAD.n6794 0.0380882
R46192 PAD.n6827 PAD.n6794 0.0380882
R46193 PAD.n6827 PAD.n6796 0.0380882
R46194 PAD.n6823 PAD.n6796 0.0380882
R46195 PAD.n6823 PAD.n6798 0.0380882
R46196 PAD.n6815 PAD.n6798 0.0380882
R46197 PAD.n6815 PAD.n6800 0.0380882
R46198 PAD.n6811 PAD.n6800 0.0380882
R46199 PAD.n6811 PAD.n6802 0.0380882
R46200 PAD.n6803 PAD.n6802 0.0380882
R46201 PAD.n7051 PAD.n6718 0.0380882
R46202 PAD.n6724 PAD.n6718 0.0380882
R46203 PAD.n7042 PAD.n6724 0.0380882
R46204 PAD.n7042 PAD.n7041 0.0380882
R46205 PAD.n7041 PAD.n7040 0.0380882
R46206 PAD.n7040 PAD.n6725 0.0380882
R46207 PAD.n7030 PAD.n6725 0.0380882
R46208 PAD.n7030 PAD.n7029 0.0380882
R46209 PAD.n7029 PAD.n7028 0.0380882
R46210 PAD.n7028 PAD.n6729 0.0380882
R46211 PAD.n7018 PAD.n6729 0.0380882
R46212 PAD.n7018 PAD.n7017 0.0380882
R46213 PAD.n7017 PAD.n7016 0.0380882
R46214 PAD.n7016 PAD.n6733 0.0380882
R46215 PAD.n7006 PAD.n6733 0.0380882
R46216 PAD.n7006 PAD.n7005 0.0380882
R46217 PAD.n7005 PAD.n7004 0.0380882
R46218 PAD.n7004 PAD.n6737 0.0380882
R46219 PAD.n6994 PAD.n6737 0.0380882
R46220 PAD.n6994 PAD.n6993 0.0380882
R46221 PAD.n6993 PAD.n6992 0.0380882
R46222 PAD.n6992 PAD.n6741 0.0380882
R46223 PAD.n6982 PAD.n6741 0.0380882
R46224 PAD.n6982 PAD.n6981 0.0380882
R46225 PAD.n6981 PAD.n6980 0.0380882
R46226 PAD.n6980 PAD.n6745 0.0380882
R46227 PAD.n6970 PAD.n6745 0.0380882
R46228 PAD.n6970 PAD.n6969 0.0380882
R46229 PAD.n6969 PAD.n6968 0.0380882
R46230 PAD.n6968 PAD.n6749 0.0380882
R46231 PAD.n6958 PAD.n6749 0.0380882
R46232 PAD.n6958 PAD.n6957 0.0380882
R46233 PAD.n6957 PAD.n6956 0.0380882
R46234 PAD.n6956 PAD.n6753 0.0380882
R46235 PAD.n6946 PAD.n6753 0.0380882
R46236 PAD.n6946 PAD.n6945 0.0380882
R46237 PAD.n6945 PAD.n6944 0.0380882
R46238 PAD.n6944 PAD.n6757 0.0380882
R46239 PAD.n6934 PAD.n6757 0.0380882
R46240 PAD.n6934 PAD.n6933 0.0380882
R46241 PAD.n6933 PAD.n6932 0.0380882
R46242 PAD.n6932 PAD.n6761 0.0380882
R46243 PAD.n6922 PAD.n6761 0.0380882
R46244 PAD.n6922 PAD.n6921 0.0380882
R46245 PAD.n6921 PAD.n6920 0.0380882
R46246 PAD.n6920 PAD.n6765 0.0380882
R46247 PAD.n6910 PAD.n6765 0.0380882
R46248 PAD.n6910 PAD.n6909 0.0380882
R46249 PAD.n6909 PAD.n6908 0.0380882
R46250 PAD.n6908 PAD.n6769 0.0380882
R46251 PAD.n6898 PAD.n6769 0.0380882
R46252 PAD.n6898 PAD.n6897 0.0380882
R46253 PAD.n6897 PAD.n6896 0.0380882
R46254 PAD.n6896 PAD.n6773 0.0380882
R46255 PAD.n6886 PAD.n6773 0.0380882
R46256 PAD.n6886 PAD.n6885 0.0380882
R46257 PAD.n6885 PAD.n6884 0.0380882
R46258 PAD.n6884 PAD.n6777 0.0380882
R46259 PAD.n6874 PAD.n6777 0.0380882
R46260 PAD.n6874 PAD.n6873 0.0380882
R46261 PAD.n6873 PAD.n6872 0.0380882
R46262 PAD.n6872 PAD.n6781 0.0380882
R46263 PAD.n6862 PAD.n6781 0.0380882
R46264 PAD.n6862 PAD.n6861 0.0380882
R46265 PAD.n6861 PAD.n6860 0.0380882
R46266 PAD.n6860 PAD.n6785 0.0380882
R46267 PAD.n6850 PAD.n6785 0.0380882
R46268 PAD.n6850 PAD.n6849 0.0380882
R46269 PAD.n6849 PAD.n6848 0.0380882
R46270 PAD.n6848 PAD.n6789 0.0380882
R46271 PAD.n6838 PAD.n6789 0.0380882
R46272 PAD.n6838 PAD.n6837 0.0380882
R46273 PAD.n6837 PAD.n6836 0.0380882
R46274 PAD.n6836 PAD.n6793 0.0380882
R46275 PAD.n6826 PAD.n6793 0.0380882
R46276 PAD.n6826 PAD.n6825 0.0380882
R46277 PAD.n6825 PAD.n6824 0.0380882
R46278 PAD.n6824 PAD.n6797 0.0380882
R46279 PAD.n6814 PAD.n6797 0.0380882
R46280 PAD.n6814 PAD.n6813 0.0380882
R46281 PAD.n6813 PAD.n6812 0.0380882
R46282 PAD.n6812 PAD.n6801 0.0380882
R46283 PAD.n6801 PAD.n6705 0.0380882
R46284 PAD.n5891 PAD.n5890 0.0380882
R46285 PAD.n5890 PAD.n5605 0.0380882
R46286 PAD.n5886 PAD.n5605 0.0380882
R46287 PAD.n5886 PAD.n5882 0.0380882
R46288 PAD.n5882 PAD.n5881 0.0380882
R46289 PAD.n5881 PAD.n5607 0.0380882
R46290 PAD.n5877 PAD.n5607 0.0380882
R46291 PAD.n5877 PAD.n5873 0.0380882
R46292 PAD.n5873 PAD.n5872 0.0380882
R46293 PAD.n5872 PAD.n5612 0.0380882
R46294 PAD.n5868 PAD.n5612 0.0380882
R46295 PAD.n5868 PAD.n5864 0.0380882
R46296 PAD.n5864 PAD.n5863 0.0380882
R46297 PAD.n5863 PAD.n5617 0.0380882
R46298 PAD.n5859 PAD.n5617 0.0380882
R46299 PAD.n5859 PAD.n5855 0.0380882
R46300 PAD.n5855 PAD.n5854 0.0380882
R46301 PAD.n5854 PAD.n5622 0.0380882
R46302 PAD.n5850 PAD.n5622 0.0380882
R46303 PAD.n5850 PAD.n5846 0.0380882
R46304 PAD.n5846 PAD.n5845 0.0380882
R46305 PAD.n5845 PAD.n5627 0.0380882
R46306 PAD.n5841 PAD.n5627 0.0380882
R46307 PAD.n5841 PAD.n5837 0.0380882
R46308 PAD.n5837 PAD.n5836 0.0380882
R46309 PAD.n5836 PAD.n5632 0.0380882
R46310 PAD.n5832 PAD.n5632 0.0380882
R46311 PAD.n5832 PAD.n5828 0.0380882
R46312 PAD.n5828 PAD.n5827 0.0380882
R46313 PAD.n5827 PAD.n5637 0.0380882
R46314 PAD.n5823 PAD.n5637 0.0380882
R46315 PAD.n5823 PAD.n5819 0.0380882
R46316 PAD.n5819 PAD.n5818 0.0380882
R46317 PAD.n5818 PAD.n5642 0.0380882
R46318 PAD.n5814 PAD.n5642 0.0380882
R46319 PAD.n5814 PAD.n5810 0.0380882
R46320 PAD.n5810 PAD.n5809 0.0380882
R46321 PAD.n5809 PAD.n5647 0.0380882
R46322 PAD.n5805 PAD.n5647 0.0380882
R46323 PAD.n5805 PAD.n5801 0.0380882
R46324 PAD.n5801 PAD.n5800 0.0380882
R46325 PAD.n5800 PAD.n5652 0.0380882
R46326 PAD.n5796 PAD.n5652 0.0380882
R46327 PAD.n5796 PAD.n5792 0.0380882
R46328 PAD.n5792 PAD.n5791 0.0380882
R46329 PAD.n5791 PAD.n5657 0.0380882
R46330 PAD.n5787 PAD.n5657 0.0380882
R46331 PAD.n5787 PAD.n5783 0.0380882
R46332 PAD.n5783 PAD.n5782 0.0380882
R46333 PAD.n5782 PAD.n5662 0.0380882
R46334 PAD.n5778 PAD.n5662 0.0380882
R46335 PAD.n5778 PAD.n5774 0.0380882
R46336 PAD.n5774 PAD.n5773 0.0380882
R46337 PAD.n5773 PAD.n5667 0.0380882
R46338 PAD.n5769 PAD.n5667 0.0380882
R46339 PAD.n5769 PAD.n5765 0.0380882
R46340 PAD.n5765 PAD.n5764 0.0380882
R46341 PAD.n5764 PAD.n5672 0.0380882
R46342 PAD.n5760 PAD.n5672 0.0380882
R46343 PAD.n5760 PAD.n5756 0.0380882
R46344 PAD.n5756 PAD.n5755 0.0380882
R46345 PAD.n5755 PAD.n5677 0.0380882
R46346 PAD.n5751 PAD.n5677 0.0380882
R46347 PAD.n5751 PAD.n5747 0.0380882
R46348 PAD.n5747 PAD.n5746 0.0380882
R46349 PAD.n5746 PAD.n5682 0.0380882
R46350 PAD.n5742 PAD.n5682 0.0380882
R46351 PAD.n5742 PAD.n5738 0.0380882
R46352 PAD.n5738 PAD.n5737 0.0380882
R46353 PAD.n5737 PAD.n5687 0.0380882
R46354 PAD.n5733 PAD.n5687 0.0380882
R46355 PAD.n5733 PAD.n5729 0.0380882
R46356 PAD.n5729 PAD.n5728 0.0380882
R46357 PAD.n5728 PAD.n5692 0.0380882
R46358 PAD.n5724 PAD.n5692 0.0380882
R46359 PAD.n5724 PAD.n5720 0.0380882
R46360 PAD.n5720 PAD.n5719 0.0380882
R46361 PAD.n5719 PAD.n5697 0.0380882
R46362 PAD.n5715 PAD.n5697 0.0380882
R46363 PAD.n5715 PAD.n5711 0.0380882
R46364 PAD.n5711 PAD.n5710 0.0380882
R46365 PAD.n5710 PAD.n5704 0.0380882
R46366 PAD.n5704 PAD.n5703 0.0380882
R46367 PAD.n5889 PAD.n5545 0.0380882
R46368 PAD.n5889 PAD.n5888 0.0380882
R46369 PAD.n5888 PAD.n5887 0.0380882
R46370 PAD.n5887 PAD.n5606 0.0380882
R46371 PAD.n5880 PAD.n5606 0.0380882
R46372 PAD.n5880 PAD.n5879 0.0380882
R46373 PAD.n5879 PAD.n5878 0.0380882
R46374 PAD.n5878 PAD.n5611 0.0380882
R46375 PAD.n5871 PAD.n5611 0.0380882
R46376 PAD.n5871 PAD.n5870 0.0380882
R46377 PAD.n5870 PAD.n5869 0.0380882
R46378 PAD.n5869 PAD.n5616 0.0380882
R46379 PAD.n5862 PAD.n5616 0.0380882
R46380 PAD.n5862 PAD.n5861 0.0380882
R46381 PAD.n5861 PAD.n5860 0.0380882
R46382 PAD.n5860 PAD.n5621 0.0380882
R46383 PAD.n5853 PAD.n5621 0.0380882
R46384 PAD.n5853 PAD.n5852 0.0380882
R46385 PAD.n5852 PAD.n5851 0.0380882
R46386 PAD.n5851 PAD.n5626 0.0380882
R46387 PAD.n5844 PAD.n5626 0.0380882
R46388 PAD.n5844 PAD.n5843 0.0380882
R46389 PAD.n5843 PAD.n5842 0.0380882
R46390 PAD.n5842 PAD.n5631 0.0380882
R46391 PAD.n5835 PAD.n5631 0.0380882
R46392 PAD.n5835 PAD.n5834 0.0380882
R46393 PAD.n5834 PAD.n5833 0.0380882
R46394 PAD.n5833 PAD.n5636 0.0380882
R46395 PAD.n5826 PAD.n5636 0.0380882
R46396 PAD.n5826 PAD.n5825 0.0380882
R46397 PAD.n5825 PAD.n5824 0.0380882
R46398 PAD.n5824 PAD.n5641 0.0380882
R46399 PAD.n5817 PAD.n5641 0.0380882
R46400 PAD.n5817 PAD.n5816 0.0380882
R46401 PAD.n5816 PAD.n5815 0.0380882
R46402 PAD.n5815 PAD.n5646 0.0380882
R46403 PAD.n5808 PAD.n5646 0.0380882
R46404 PAD.n5808 PAD.n5807 0.0380882
R46405 PAD.n5807 PAD.n5806 0.0380882
R46406 PAD.n5806 PAD.n5651 0.0380882
R46407 PAD.n5799 PAD.n5651 0.0380882
R46408 PAD.n5799 PAD.n5798 0.0380882
R46409 PAD.n5798 PAD.n5797 0.0380882
R46410 PAD.n5797 PAD.n5656 0.0380882
R46411 PAD.n5790 PAD.n5656 0.0380882
R46412 PAD.n5790 PAD.n5789 0.0380882
R46413 PAD.n5789 PAD.n5788 0.0380882
R46414 PAD.n5788 PAD.n5661 0.0380882
R46415 PAD.n5781 PAD.n5661 0.0380882
R46416 PAD.n5781 PAD.n5780 0.0380882
R46417 PAD.n5780 PAD.n5779 0.0380882
R46418 PAD.n5779 PAD.n5666 0.0380882
R46419 PAD.n5772 PAD.n5666 0.0380882
R46420 PAD.n5772 PAD.n5771 0.0380882
R46421 PAD.n5771 PAD.n5770 0.0380882
R46422 PAD.n5770 PAD.n5671 0.0380882
R46423 PAD.n5763 PAD.n5671 0.0380882
R46424 PAD.n5763 PAD.n5762 0.0380882
R46425 PAD.n5762 PAD.n5761 0.0380882
R46426 PAD.n5761 PAD.n5676 0.0380882
R46427 PAD.n5754 PAD.n5676 0.0380882
R46428 PAD.n5754 PAD.n5753 0.0380882
R46429 PAD.n5753 PAD.n5752 0.0380882
R46430 PAD.n5752 PAD.n5681 0.0380882
R46431 PAD.n5745 PAD.n5681 0.0380882
R46432 PAD.n5745 PAD.n5744 0.0380882
R46433 PAD.n5744 PAD.n5743 0.0380882
R46434 PAD.n5743 PAD.n5686 0.0380882
R46435 PAD.n5736 PAD.n5686 0.0380882
R46436 PAD.n5736 PAD.n5735 0.0380882
R46437 PAD.n5735 PAD.n5734 0.0380882
R46438 PAD.n5734 PAD.n5691 0.0380882
R46439 PAD.n5727 PAD.n5691 0.0380882
R46440 PAD.n5727 PAD.n5726 0.0380882
R46441 PAD.n5726 PAD.n5725 0.0380882
R46442 PAD.n5725 PAD.n5696 0.0380882
R46443 PAD.n5718 PAD.n5696 0.0380882
R46444 PAD.n5718 PAD.n5717 0.0380882
R46445 PAD.n5717 PAD.n5716 0.0380882
R46446 PAD.n5716 PAD.n5701 0.0380882
R46447 PAD.n5709 PAD.n5701 0.0380882
R46448 PAD.n5709 PAD.n5708 0.0380882
R46449 PAD.n5708 PAD.n5557 0.0380882
R46450 PAD.n11087 PAD.n10747 0.0380882
R46451 PAD.n11079 PAD.n10747 0.0380882
R46452 PAD.n11079 PAD.n11078 0.0380882
R46453 PAD.n11078 PAD.n11077 0.0380882
R46454 PAD.n11077 PAD.n10758 0.0380882
R46455 PAD.n11067 PAD.n10758 0.0380882
R46456 PAD.n11067 PAD.n11066 0.0380882
R46457 PAD.n11066 PAD.n11065 0.0380882
R46458 PAD.n11065 PAD.n10762 0.0380882
R46459 PAD.n11055 PAD.n10762 0.0380882
R46460 PAD.n11055 PAD.n11054 0.0380882
R46461 PAD.n11054 PAD.n11053 0.0380882
R46462 PAD.n11053 PAD.n10766 0.0380882
R46463 PAD.n11043 PAD.n10766 0.0380882
R46464 PAD.n11043 PAD.n11042 0.0380882
R46465 PAD.n11042 PAD.n11041 0.0380882
R46466 PAD.n11041 PAD.n10770 0.0380882
R46467 PAD.n11031 PAD.n10770 0.0380882
R46468 PAD.n11031 PAD.n11030 0.0380882
R46469 PAD.n11030 PAD.n11029 0.0380882
R46470 PAD.n11029 PAD.n10774 0.0380882
R46471 PAD.n11019 PAD.n10774 0.0380882
R46472 PAD.n11019 PAD.n11018 0.0380882
R46473 PAD.n11018 PAD.n11017 0.0380882
R46474 PAD.n11017 PAD.n10778 0.0380882
R46475 PAD.n11007 PAD.n10778 0.0380882
R46476 PAD.n11007 PAD.n11006 0.0380882
R46477 PAD.n11006 PAD.n11005 0.0380882
R46478 PAD.n11005 PAD.n10782 0.0380882
R46479 PAD.n10995 PAD.n10782 0.0380882
R46480 PAD.n10995 PAD.n10994 0.0380882
R46481 PAD.n10994 PAD.n10993 0.0380882
R46482 PAD.n10993 PAD.n10786 0.0380882
R46483 PAD.n10983 PAD.n10786 0.0380882
R46484 PAD.n10983 PAD.n10982 0.0380882
R46485 PAD.n10982 PAD.n10981 0.0380882
R46486 PAD.n10981 PAD.n10790 0.0380882
R46487 PAD.n10971 PAD.n10790 0.0380882
R46488 PAD.n10971 PAD.n10970 0.0380882
R46489 PAD.n10970 PAD.n10969 0.0380882
R46490 PAD.n10969 PAD.n10794 0.0380882
R46491 PAD.n10959 PAD.n10794 0.0380882
R46492 PAD.n10959 PAD.n10958 0.0380882
R46493 PAD.n10958 PAD.n10957 0.0380882
R46494 PAD.n10957 PAD.n10798 0.0380882
R46495 PAD.n10947 PAD.n10798 0.0380882
R46496 PAD.n10947 PAD.n10946 0.0380882
R46497 PAD.n10946 PAD.n10945 0.0380882
R46498 PAD.n10945 PAD.n10802 0.0380882
R46499 PAD.n10935 PAD.n10802 0.0380882
R46500 PAD.n10935 PAD.n10934 0.0380882
R46501 PAD.n10934 PAD.n10933 0.0380882
R46502 PAD.n10933 PAD.n10806 0.0380882
R46503 PAD.n10923 PAD.n10806 0.0380882
R46504 PAD.n10923 PAD.n10922 0.0380882
R46505 PAD.n10922 PAD.n10921 0.0380882
R46506 PAD.n10921 PAD.n10810 0.0380882
R46507 PAD.n10911 PAD.n10810 0.0380882
R46508 PAD.n10911 PAD.n10910 0.0380882
R46509 PAD.n10910 PAD.n10909 0.0380882
R46510 PAD.n10909 PAD.n10814 0.0380882
R46511 PAD.n10899 PAD.n10814 0.0380882
R46512 PAD.n10899 PAD.n10898 0.0380882
R46513 PAD.n10898 PAD.n10897 0.0380882
R46514 PAD.n10897 PAD.n10818 0.0380882
R46515 PAD.n10887 PAD.n10818 0.0380882
R46516 PAD.n10887 PAD.n10886 0.0380882
R46517 PAD.n10886 PAD.n10885 0.0380882
R46518 PAD.n10885 PAD.n10822 0.0380882
R46519 PAD.n10875 PAD.n10822 0.0380882
R46520 PAD.n10875 PAD.n10874 0.0380882
R46521 PAD.n10874 PAD.n10873 0.0380882
R46522 PAD.n10873 PAD.n10826 0.0380882
R46523 PAD.n10863 PAD.n10826 0.0380882
R46524 PAD.n10863 PAD.n10862 0.0380882
R46525 PAD.n10862 PAD.n10861 0.0380882
R46526 PAD.n10861 PAD.n10830 0.0380882
R46527 PAD.n10851 PAD.n10830 0.0380882
R46528 PAD.n10851 PAD.n10850 0.0380882
R46529 PAD.n10850 PAD.n10849 0.0380882
R46530 PAD.n10849 PAD.n10834 0.0380882
R46531 PAD.n10839 PAD.n10834 0.0380882
R46532 PAD.n10839 PAD.n10734 0.0380882
R46533 PAD.n6692 PAD.n5898 0.0380882
R46534 PAD.n6499 PAD.n5898 0.0380882
R46535 PAD.n6500 PAD.n6499 0.0380882
R46536 PAD.n6501 PAD.n6500 0.0380882
R46537 PAD.n6501 PAD.n6494 0.0380882
R46538 PAD.n6508 PAD.n6494 0.0380882
R46539 PAD.n6509 PAD.n6508 0.0380882
R46540 PAD.n6510 PAD.n6509 0.0380882
R46541 PAD.n6510 PAD.n6491 0.0380882
R46542 PAD.n6517 PAD.n6491 0.0380882
R46543 PAD.n6518 PAD.n6517 0.0380882
R46544 PAD.n6519 PAD.n6518 0.0380882
R46545 PAD.n6519 PAD.n6488 0.0380882
R46546 PAD.n6526 PAD.n6488 0.0380882
R46547 PAD.n6527 PAD.n6526 0.0380882
R46548 PAD.n6528 PAD.n6527 0.0380882
R46549 PAD.n6528 PAD.n6485 0.0380882
R46550 PAD.n6535 PAD.n6485 0.0380882
R46551 PAD.n6536 PAD.n6535 0.0380882
R46552 PAD.n6537 PAD.n6536 0.0380882
R46553 PAD.n6537 PAD.n6482 0.0380882
R46554 PAD.n6544 PAD.n6482 0.0380882
R46555 PAD.n6545 PAD.n6544 0.0380882
R46556 PAD.n6546 PAD.n6545 0.0380882
R46557 PAD.n6546 PAD.n6479 0.0380882
R46558 PAD.n6553 PAD.n6479 0.0380882
R46559 PAD.n6554 PAD.n6553 0.0380882
R46560 PAD.n6555 PAD.n6554 0.0380882
R46561 PAD.n6555 PAD.n6476 0.0380882
R46562 PAD.n6562 PAD.n6476 0.0380882
R46563 PAD.n6563 PAD.n6562 0.0380882
R46564 PAD.n6564 PAD.n6563 0.0380882
R46565 PAD.n6564 PAD.n6473 0.0380882
R46566 PAD.n6571 PAD.n6473 0.0380882
R46567 PAD.n6572 PAD.n6571 0.0380882
R46568 PAD.n6573 PAD.n6572 0.0380882
R46569 PAD.n6573 PAD.n6470 0.0380882
R46570 PAD.n6580 PAD.n6470 0.0380882
R46571 PAD.n6581 PAD.n6580 0.0380882
R46572 PAD.n6582 PAD.n6581 0.0380882
R46573 PAD.n6582 PAD.n6467 0.0380882
R46574 PAD.n6589 PAD.n6467 0.0380882
R46575 PAD.n6590 PAD.n6589 0.0380882
R46576 PAD.n6591 PAD.n6590 0.0380882
R46577 PAD.n6591 PAD.n6464 0.0380882
R46578 PAD.n6598 PAD.n6464 0.0380882
R46579 PAD.n6599 PAD.n6598 0.0380882
R46580 PAD.n6600 PAD.n6599 0.0380882
R46581 PAD.n6600 PAD.n6461 0.0380882
R46582 PAD.n6607 PAD.n6461 0.0380882
R46583 PAD.n6608 PAD.n6607 0.0380882
R46584 PAD.n6609 PAD.n6608 0.0380882
R46585 PAD.n6609 PAD.n6458 0.0380882
R46586 PAD.n6616 PAD.n6458 0.0380882
R46587 PAD.n6617 PAD.n6616 0.0380882
R46588 PAD.n6618 PAD.n6617 0.0380882
R46589 PAD.n6618 PAD.n6455 0.0380882
R46590 PAD.n6625 PAD.n6455 0.0380882
R46591 PAD.n6626 PAD.n6625 0.0380882
R46592 PAD.n6627 PAD.n6626 0.0380882
R46593 PAD.n6627 PAD.n6452 0.0380882
R46594 PAD.n6634 PAD.n6452 0.0380882
R46595 PAD.n6635 PAD.n6634 0.0380882
R46596 PAD.n6636 PAD.n6635 0.0380882
R46597 PAD.n6636 PAD.n6449 0.0380882
R46598 PAD.n6643 PAD.n6449 0.0380882
R46599 PAD.n6644 PAD.n6643 0.0380882
R46600 PAD.n6645 PAD.n6644 0.0380882
R46601 PAD.n6645 PAD.n6446 0.0380882
R46602 PAD.n6652 PAD.n6446 0.0380882
R46603 PAD.n6653 PAD.n6652 0.0380882
R46604 PAD.n6654 PAD.n6653 0.0380882
R46605 PAD.n6654 PAD.n6443 0.0380882
R46606 PAD.n6661 PAD.n6443 0.0380882
R46607 PAD.n6662 PAD.n6661 0.0380882
R46608 PAD.n6663 PAD.n6662 0.0380882
R46609 PAD.n6663 PAD.n6440 0.0380882
R46610 PAD.n6670 PAD.n6440 0.0380882
R46611 PAD.n6671 PAD.n6670 0.0380882
R46612 PAD.n6674 PAD.n6671 0.0380882
R46613 PAD.n6674 PAD.n6673 0.0380882
R46614 PAD.n6673 PAD.n6672 0.0380882
R46615 PAD.n6672 PAD.n5951 0.0380882
R46616 PAD.n6691 PAD.n5900 0.0380882
R46617 PAD.n6498 PAD.n5900 0.0380882
R46618 PAD.n6498 PAD.n6496 0.0380882
R46619 PAD.n6503 PAD.n6496 0.0380882
R46620 PAD.n6505 PAD.n6503 0.0380882
R46621 PAD.n6507 PAD.n6505 0.0380882
R46622 PAD.n6507 PAD.n6493 0.0380882
R46623 PAD.n6512 PAD.n6493 0.0380882
R46624 PAD.n6514 PAD.n6512 0.0380882
R46625 PAD.n6516 PAD.n6514 0.0380882
R46626 PAD.n6516 PAD.n6490 0.0380882
R46627 PAD.n6521 PAD.n6490 0.0380882
R46628 PAD.n6523 PAD.n6521 0.0380882
R46629 PAD.n6525 PAD.n6523 0.0380882
R46630 PAD.n6525 PAD.n6487 0.0380882
R46631 PAD.n6530 PAD.n6487 0.0380882
R46632 PAD.n6532 PAD.n6530 0.0380882
R46633 PAD.n6534 PAD.n6532 0.0380882
R46634 PAD.n6534 PAD.n6484 0.0380882
R46635 PAD.n6539 PAD.n6484 0.0380882
R46636 PAD.n6541 PAD.n6539 0.0380882
R46637 PAD.n6543 PAD.n6541 0.0380882
R46638 PAD.n6543 PAD.n6481 0.0380882
R46639 PAD.n6548 PAD.n6481 0.0380882
R46640 PAD.n6550 PAD.n6548 0.0380882
R46641 PAD.n6552 PAD.n6550 0.0380882
R46642 PAD.n6552 PAD.n6478 0.0380882
R46643 PAD.n6557 PAD.n6478 0.0380882
R46644 PAD.n6559 PAD.n6557 0.0380882
R46645 PAD.n6561 PAD.n6559 0.0380882
R46646 PAD.n6561 PAD.n6475 0.0380882
R46647 PAD.n6566 PAD.n6475 0.0380882
R46648 PAD.n6568 PAD.n6566 0.0380882
R46649 PAD.n6570 PAD.n6568 0.0380882
R46650 PAD.n6570 PAD.n6472 0.0380882
R46651 PAD.n6575 PAD.n6472 0.0380882
R46652 PAD.n6577 PAD.n6575 0.0380882
R46653 PAD.n6579 PAD.n6577 0.0380882
R46654 PAD.n6579 PAD.n6469 0.0380882
R46655 PAD.n6584 PAD.n6469 0.0380882
R46656 PAD.n6586 PAD.n6584 0.0380882
R46657 PAD.n6588 PAD.n6586 0.0380882
R46658 PAD.n6588 PAD.n6466 0.0380882
R46659 PAD.n6593 PAD.n6466 0.0380882
R46660 PAD.n6595 PAD.n6593 0.0380882
R46661 PAD.n6597 PAD.n6595 0.0380882
R46662 PAD.n6597 PAD.n6463 0.0380882
R46663 PAD.n6602 PAD.n6463 0.0380882
R46664 PAD.n6604 PAD.n6602 0.0380882
R46665 PAD.n6606 PAD.n6604 0.0380882
R46666 PAD.n6606 PAD.n6460 0.0380882
R46667 PAD.n6611 PAD.n6460 0.0380882
R46668 PAD.n6613 PAD.n6611 0.0380882
R46669 PAD.n6615 PAD.n6613 0.0380882
R46670 PAD.n6615 PAD.n6457 0.0380882
R46671 PAD.n6620 PAD.n6457 0.0380882
R46672 PAD.n6622 PAD.n6620 0.0380882
R46673 PAD.n6624 PAD.n6622 0.0380882
R46674 PAD.n6624 PAD.n6454 0.0380882
R46675 PAD.n6629 PAD.n6454 0.0380882
R46676 PAD.n6631 PAD.n6629 0.0380882
R46677 PAD.n6633 PAD.n6631 0.0380882
R46678 PAD.n6633 PAD.n6451 0.0380882
R46679 PAD.n6638 PAD.n6451 0.0380882
R46680 PAD.n6640 PAD.n6638 0.0380882
R46681 PAD.n6642 PAD.n6640 0.0380882
R46682 PAD.n6642 PAD.n6448 0.0380882
R46683 PAD.n6647 PAD.n6448 0.0380882
R46684 PAD.n6649 PAD.n6647 0.0380882
R46685 PAD.n6651 PAD.n6649 0.0380882
R46686 PAD.n6651 PAD.n6445 0.0380882
R46687 PAD.n6656 PAD.n6445 0.0380882
R46688 PAD.n6658 PAD.n6656 0.0380882
R46689 PAD.n6660 PAD.n6658 0.0380882
R46690 PAD.n6660 PAD.n6442 0.0380882
R46691 PAD.n6665 PAD.n6442 0.0380882
R46692 PAD.n6667 PAD.n6665 0.0380882
R46693 PAD.n6669 PAD.n6667 0.0380882
R46694 PAD.n6669 PAD.n6438 0.0380882
R46695 PAD.n6675 PAD.n6438 0.0380882
R46696 PAD.n6675 PAD.n6439 0.0380882
R46697 PAD.n6439 PAD.n5950 0.0380882
R46698 PAD.n6687 PAD.n5950 0.0380882
R46699 PAD.n119 PAD.n118 0.0380882
R46700 PAD.n123 PAD.n118 0.0380882
R46701 PAD.n127 PAD.n123 0.0380882
R46702 PAD.n131 PAD.n127 0.0380882
R46703 PAD.n131 PAD.n114 0.0380882
R46704 PAD.n135 PAD.n114 0.0380882
R46705 PAD.n139 PAD.n135 0.0380882
R46706 PAD.n143 PAD.n139 0.0380882
R46707 PAD.n143 PAD.n112 0.0380882
R46708 PAD.n147 PAD.n112 0.0380882
R46709 PAD.n151 PAD.n147 0.0380882
R46710 PAD.n155 PAD.n151 0.0380882
R46711 PAD.n155 PAD.n110 0.0380882
R46712 PAD.n159 PAD.n110 0.0380882
R46713 PAD.n163 PAD.n159 0.0380882
R46714 PAD.n167 PAD.n163 0.0380882
R46715 PAD.n167 PAD.n108 0.0380882
R46716 PAD.n171 PAD.n108 0.0380882
R46717 PAD.n175 PAD.n171 0.0380882
R46718 PAD.n179 PAD.n175 0.0380882
R46719 PAD.n179 PAD.n106 0.0380882
R46720 PAD.n183 PAD.n106 0.0380882
R46721 PAD.n187 PAD.n183 0.0380882
R46722 PAD.n191 PAD.n187 0.0380882
R46723 PAD.n191 PAD.n104 0.0380882
R46724 PAD.n195 PAD.n104 0.0380882
R46725 PAD.n199 PAD.n195 0.0380882
R46726 PAD.n203 PAD.n199 0.0380882
R46727 PAD.n203 PAD.n102 0.0380882
R46728 PAD.n207 PAD.n102 0.0380882
R46729 PAD.n211 PAD.n207 0.0380882
R46730 PAD.n215 PAD.n211 0.0380882
R46731 PAD.n215 PAD.n100 0.0380882
R46732 PAD.n219 PAD.n100 0.0380882
R46733 PAD.n223 PAD.n219 0.0380882
R46734 PAD.n227 PAD.n223 0.0380882
R46735 PAD.n227 PAD.n98 0.0380882
R46736 PAD.n231 PAD.n98 0.0380882
R46737 PAD.n235 PAD.n231 0.0380882
R46738 PAD.n239 PAD.n235 0.0380882
R46739 PAD.n239 PAD.n96 0.0380882
R46740 PAD.n243 PAD.n96 0.0380882
R46741 PAD.n247 PAD.n243 0.0380882
R46742 PAD.n251 PAD.n247 0.0380882
R46743 PAD.n251 PAD.n94 0.0380882
R46744 PAD.n255 PAD.n94 0.0380882
R46745 PAD.n259 PAD.n255 0.0380882
R46746 PAD.n263 PAD.n259 0.0380882
R46747 PAD.n263 PAD.n92 0.0380882
R46748 PAD.n267 PAD.n92 0.0380882
R46749 PAD.n271 PAD.n267 0.0380882
R46750 PAD.n275 PAD.n271 0.0380882
R46751 PAD.n275 PAD.n90 0.0380882
R46752 PAD.n279 PAD.n90 0.0380882
R46753 PAD.n283 PAD.n279 0.0380882
R46754 PAD.n287 PAD.n283 0.0380882
R46755 PAD.n287 PAD.n88 0.0380882
R46756 PAD.n291 PAD.n88 0.0380882
R46757 PAD.n295 PAD.n291 0.0380882
R46758 PAD.n299 PAD.n295 0.0380882
R46759 PAD.n299 PAD.n86 0.0380882
R46760 PAD.n303 PAD.n86 0.0380882
R46761 PAD.n307 PAD.n303 0.0380882
R46762 PAD.n311 PAD.n307 0.0380882
R46763 PAD.n311 PAD.n84 0.0380882
R46764 PAD.n315 PAD.n84 0.0380882
R46765 PAD.n319 PAD.n315 0.0380882
R46766 PAD.n323 PAD.n319 0.0380882
R46767 PAD.n323 PAD.n82 0.0380882
R46768 PAD.n327 PAD.n82 0.0380882
R46769 PAD.n331 PAD.n327 0.0380882
R46770 PAD.n335 PAD.n331 0.0380882
R46771 PAD.n335 PAD.n80 0.0380882
R46772 PAD.n339 PAD.n80 0.0380882
R46773 PAD.n343 PAD.n339 0.0380882
R46774 PAD.n347 PAD.n343 0.0380882
R46775 PAD.n347 PAD.n78 0.0380882
R46776 PAD.n351 PAD.n78 0.0380882
R46777 PAD.n355 PAD.n351 0.0380882
R46778 PAD.n359 PAD.n355 0.0380882
R46779 PAD.n359 PAD.n76 0.0380882
R46780 PAD.n363 PAD.n76 0.0380882
R46781 PAD.n363 PAD.n75 0.0380882
R46782 PAD.n11086 PAD.n10749 0.0380882
R46783 PAD.n11080 PAD.n10749 0.0380882
R46784 PAD.n11080 PAD.n10757 0.0380882
R46785 PAD.n11076 PAD.n10757 0.0380882
R46786 PAD.n11076 PAD.n10759 0.0380882
R46787 PAD.n11068 PAD.n10759 0.0380882
R46788 PAD.n11068 PAD.n10761 0.0380882
R46789 PAD.n11064 PAD.n10761 0.0380882
R46790 PAD.n11064 PAD.n10763 0.0380882
R46791 PAD.n11056 PAD.n10763 0.0380882
R46792 PAD.n11056 PAD.n10765 0.0380882
R46793 PAD.n11052 PAD.n10765 0.0380882
R46794 PAD.n11052 PAD.n10767 0.0380882
R46795 PAD.n11044 PAD.n10767 0.0380882
R46796 PAD.n11044 PAD.n10769 0.0380882
R46797 PAD.n11040 PAD.n10769 0.0380882
R46798 PAD.n11040 PAD.n10771 0.0380882
R46799 PAD.n11032 PAD.n10771 0.0380882
R46800 PAD.n11032 PAD.n10773 0.0380882
R46801 PAD.n11028 PAD.n10773 0.0380882
R46802 PAD.n11028 PAD.n10775 0.0380882
R46803 PAD.n11020 PAD.n10775 0.0380882
R46804 PAD.n11020 PAD.n10777 0.0380882
R46805 PAD.n11016 PAD.n10777 0.0380882
R46806 PAD.n11016 PAD.n10779 0.0380882
R46807 PAD.n11008 PAD.n10779 0.0380882
R46808 PAD.n11008 PAD.n10781 0.0380882
R46809 PAD.n11004 PAD.n10781 0.0380882
R46810 PAD.n11004 PAD.n10783 0.0380882
R46811 PAD.n10996 PAD.n10783 0.0380882
R46812 PAD.n10996 PAD.n10785 0.0380882
R46813 PAD.n10992 PAD.n10785 0.0380882
R46814 PAD.n10992 PAD.n10787 0.0380882
R46815 PAD.n10984 PAD.n10787 0.0380882
R46816 PAD.n10984 PAD.n10789 0.0380882
R46817 PAD.n10980 PAD.n10789 0.0380882
R46818 PAD.n10980 PAD.n10791 0.0380882
R46819 PAD.n10972 PAD.n10791 0.0380882
R46820 PAD.n10972 PAD.n10793 0.0380882
R46821 PAD.n10968 PAD.n10793 0.0380882
R46822 PAD.n10968 PAD.n10795 0.0380882
R46823 PAD.n10960 PAD.n10795 0.0380882
R46824 PAD.n10960 PAD.n10797 0.0380882
R46825 PAD.n10956 PAD.n10797 0.0380882
R46826 PAD.n10956 PAD.n10799 0.0380882
R46827 PAD.n10948 PAD.n10799 0.0380882
R46828 PAD.n10948 PAD.n10801 0.0380882
R46829 PAD.n10944 PAD.n10801 0.0380882
R46830 PAD.n10944 PAD.n10803 0.0380882
R46831 PAD.n10936 PAD.n10803 0.0380882
R46832 PAD.n10936 PAD.n10805 0.0380882
R46833 PAD.n10932 PAD.n10805 0.0380882
R46834 PAD.n10932 PAD.n10807 0.0380882
R46835 PAD.n10924 PAD.n10807 0.0380882
R46836 PAD.n10924 PAD.n10809 0.0380882
R46837 PAD.n10920 PAD.n10809 0.0380882
R46838 PAD.n10920 PAD.n10811 0.0380882
R46839 PAD.n10912 PAD.n10811 0.0380882
R46840 PAD.n10912 PAD.n10813 0.0380882
R46841 PAD.n10908 PAD.n10813 0.0380882
R46842 PAD.n10908 PAD.n10815 0.0380882
R46843 PAD.n10900 PAD.n10815 0.0380882
R46844 PAD.n10900 PAD.n10817 0.0380882
R46845 PAD.n10896 PAD.n10817 0.0380882
R46846 PAD.n10896 PAD.n10819 0.0380882
R46847 PAD.n10888 PAD.n10819 0.0380882
R46848 PAD.n10888 PAD.n10821 0.0380882
R46849 PAD.n10884 PAD.n10821 0.0380882
R46850 PAD.n10884 PAD.n10823 0.0380882
R46851 PAD.n10876 PAD.n10823 0.0380882
R46852 PAD.n10876 PAD.n10825 0.0380882
R46853 PAD.n10872 PAD.n10825 0.0380882
R46854 PAD.n10872 PAD.n10827 0.0380882
R46855 PAD.n10864 PAD.n10827 0.0380882
R46856 PAD.n10864 PAD.n10829 0.0380882
R46857 PAD.n10860 PAD.n10829 0.0380882
R46858 PAD.n10860 PAD.n10831 0.0380882
R46859 PAD.n10852 PAD.n10831 0.0380882
R46860 PAD.n10852 PAD.n10833 0.0380882
R46861 PAD.n10848 PAD.n10833 0.0380882
R46862 PAD.n10848 PAD.n10835 0.0380882
R46863 PAD.n10840 PAD.n10835 0.0380882
R46864 PAD.n10840 PAD.n10838 0.0380882
R46865 PAD.n7810 PAD.n3637 0.0368392
R46866 PAD.n9168 PAD.n12 0.035749
R46867 PAD.n0 PAD 0.0336535
R46868 PAD.n6380 PAD.n6379 0.03245
R46869 PAD.n6379 PAD.n6378 0.03245
R46870 PAD.n5953 PAD.n5558 0.03245
R46871 PAD.n6703 PAD.n5558 0.03245
R46872 PAD.n7798 PAD.n7797 0.03245
R46873 PAD.n7795 PAD.n6706 0.03245
R46874 PAD.n7153 PAD.n6706 0.03245
R46875 PAD.n7526 PAD.n7525 0.03245
R46876 PAD.n7525 PAD.n7524 0.03245
R46877 PAD.n7203 PAD.n5201 0.03245
R46878 PAD.n7823 PAD.n5201 0.03245
R46879 PAD.n7825 PAD.n5187 0.03245
R46880 PAD.n8178 PAD.n5187 0.03245
R46881 PAD.n8180 PAD.n4836 0.03245
R46882 PAD.n8198 PAD.n4836 0.03245
R46883 PAD.n8200 PAD.n4830 0.03245
R46884 PAD.n8208 PAD.n4670 0.03245
R46885 PAD.n8413 PAD.n4670 0.03245
R46886 PAD.n8416 PAD.n8415 0.03245
R46887 PAD.n8415 PAD.n4315 0.03245
R46888 PAD.n8436 PAD.n4316 0.03245
R46889 PAD.n4316 PAD.n3974 0.03245
R46890 PAD.n8460 PAD.n3629 0.03245
R46891 PAD.n8483 PAD.n3629 0.03245
R46892 PAD.n8484 PAD.n3284 0.03245
R46893 PAD.n8509 PAD.n2899 0.03245
R46894 PAD.n8825 PAD.n2899 0.03245
R46895 PAD.n8828 PAD.n8827 0.03245
R46896 PAD.n8828 PAD.n2882 0.03245
R46897 PAD.n9132 PAD.n2491 0.03245
R46898 PAD.n9155 PAD.n2491 0.03245
R46899 PAD.n9157 PAD.n2143 0.03245
R46900 PAD.n9179 PAD.n2143 0.03245
R46901 PAD.n9181 PAD.n2041 0.03245
R46902 PAD.n9449 PAD.n2041 0.03245
R46903 PAD.n9452 PAD.n9451 0.03245
R46904 PAD.n9717 PAD.n9716 0.03245
R46905 PAD.n9718 PAD.n9717 0.03245
R46906 PAD.n9737 PAD.n9736 0.03245
R46907 PAD.n9738 PAD.n9737 0.03245
R46908 PAD.n10003 PAD.n10002 0.03245
R46909 PAD.n10004 PAD.n10003 0.03245
R46910 PAD.n10021 PAD.n10020 0.03245
R46911 PAD.n10358 PAD.n10021 0.03245
R46912 PAD.n10356 PAD.n1115 0.03245
R46913 PAD.n10380 PAD.n773 0.03245
R46914 PAD.n10401 PAD.n773 0.03245
R46915 PAD.n10404 PAD.n10403 0.03245
R46916 PAD.n10403 PAD.n422 0.03245
R46917 PAD.n10708 PAD.n27 0.03245
R46918 PAD.n10731 PAD.n27 0.03245
R46919 PAD.n11529 PAD.n10733 0.03245
R46920 PAD.n11529 PAD.n11528 0.03245
R46921 PAD.n11526 PAD.n10735 0.03245
R46922 PAD.n11504 PAD.n10735 0.03245
R46923 PAD.n7797 PAD.n7796 0.031775
R46924 PAD.n7516 PAD.n7227 0.0317353
R46925 PAD.n120 PAD.n14 0.0317353
R46926 PAD.n10697 PAD.n10696 0.0317353
R46927 PAD.n521 PAD.n430 0.0317353
R46928 PAD.n873 PAD.n779 0.0317353
R46929 PAD.n10367 PAD.n1124 0.0317353
R46930 PAD.n10012 PAD.n1145 0.0317353
R46931 PAD.n9750 PAD.n1580 0.0317353
R46932 PAD.n9726 PAD.n1932 0.0317353
R46933 PAD.n9464 PAD.n2032 0.0317353
R46934 PAD.n9198 PAD.n2135 0.0317353
R46935 PAD.n9167 PAD.n2483 0.0317353
R46936 PAD.n9147 PAD.n2830 0.0317353
R46937 PAD.n9124 PAD.n9120 0.0317353
R46938 PAD.n8817 PAD.n2888 0.0317353
R46939 PAD.n3042 PAD.n2949 0.0317353
R46940 PAD.n3387 PAD.n3293 0.0317353
R46941 PAD.n3732 PAD.n3638 0.0317353
R46942 PAD.n4073 PAD.n3980 0.0317353
R46943 PAD.n8424 PAD.n4325 0.0317353
R46944 PAD.n8402 PAD.n4676 0.0317353
R46945 PAD.n8190 PAD.n5179 0.0317353
R46946 PAD.n8170 PAD.n5193 0.0317353
R46947 PAD.n7815 PAD.n5543 0.0317353
R46948 PAD.n7778 PAD.n7056 0.0317353
R46949 PAD.n7055 PAD.n7051 0.0317353
R46950 PAD.n7806 PAD.n5545 0.0317353
R46951 PAD.n11088 PAD.n11087 0.0317353
R46952 PAD.n6693 PAD.n6692 0.0317353
R46953 PAD.n8510 PAD.n3284 0.031325
R46954 PAD.n9451 PAD.n9450 0.030875
R46955 PAD.n10381 PAD.n1115 0.030875
R46956 PAD.n8200 PAD.n8199 0.030425
R46957 PAD.n8209 PAD.n4830 0.028625
R46958 PAD.n6381 PAD.n5977 0.0284039
R46959 PAD.n5977 PAD.n5952 0.0284039
R46960 PAD.n6685 PAD.n5559 0.0284039
R46961 PAD.n6702 PAD.n5559 0.0284039
R46962 PAD.n7799 PAD.n5556 0.0284039
R46963 PAD.n7794 PAD.n6708 0.0284039
R46964 PAD.n7152 PAD.n6708 0.0284039
R46965 PAD.n7527 PAD.n7151 0.0284039
R46966 PAD.n7523 PAD.n7151 0.0284039
R46967 PAD.n7204 PAD.n5202 0.0284039
R46968 PAD.n7822 PAD.n5202 0.0284039
R46969 PAD.n7826 PAD.n5188 0.0284039
R46970 PAD.n8177 PAD.n5188 0.0284039
R46971 PAD.n8181 PAD.n4837 0.0284039
R46972 PAD.n8197 PAD.n4837 0.0284039
R46973 PAD.n8202 PAD.n8201 0.0284039
R46974 PAD.n8207 PAD.n4671 0.0284039
R46975 PAD.n8412 PAD.n4671 0.0284039
R46976 PAD.n8417 PAD.n4317 0.0284039
R46977 PAD.n8433 PAD.n4317 0.0284039
R46978 PAD.n8435 PAD.n3975 0.0284039
R46979 PAD.n8457 PAD.n3975 0.0284039
R46980 PAD.n8459 PAD.n3630 0.0284039
R46981 PAD.n8482 PAD.n3630 0.0284039
R46982 PAD.n8505 PAD.n3285 0.0284039
R46983 PAD.n8508 PAD.n2900 0.0284039
R46984 PAD.n8824 PAD.n2900 0.0284039
R46985 PAD.n8829 PAD.n2896 0.0284039
R46986 PAD.n8829 PAD.n2897 0.0284039
R46987 PAD.n9131 PAD.n2492 0.0284039
R46988 PAD.n9154 PAD.n2492 0.0284039
R46989 PAD.n9158 PAD.n2144 0.0284039
R46990 PAD.n9178 PAD.n2144 0.0284039
R46991 PAD.n9182 PAD.n2042 0.0284039
R46992 PAD.n9448 PAD.n2042 0.0284039
R46993 PAD.n9453 PAD.n2039 0.0284039
R46994 PAD.n9715 PAD.n1938 0.0284039
R46995 PAD.n9719 PAD.n1938 0.0284039
R46996 PAD.n9735 PAD.n1588 0.0284039
R46997 PAD.n9739 PAD.n1588 0.0284039
R46998 PAD.n10001 PAD.n1485 0.0284039
R46999 PAD.n10005 PAD.n1485 0.0284039
R47000 PAD.n10019 PAD.n1135 0.0284039
R47001 PAD.n10359 PAD.n1135 0.0284039
R47002 PAD.n10376 PAD.n1116 0.0284039
R47003 PAD.n10379 PAD.n774 0.0284039
R47004 PAD.n10400 PAD.n774 0.0284039
R47005 PAD.n10405 PAD.n423 0.0284039
R47006 PAD.n10704 PAD.n423 0.0284039
R47007 PAD.n10707 PAD.n28 0.0284039
R47008 PAD.n10730 PAD.n28 0.0284039
R47009 PAD.n11530 PAD.n24 0.0284039
R47010 PAD.n11530 PAD.n25 0.0284039
R47011 PAD.n11525 PAD.n10737 0.0284039
R47012 PAD.n11503 PAD.n10737 0.0284039
R47013 PAD.n6382 PAD.n5975 0.0284039
R47014 PAD.n5975 PAD.n5973 0.0284039
R47015 PAD.n6684 PAD.n5560 0.0284039
R47016 PAD.n6701 PAD.n5560 0.0284039
R47017 PAD.n7800 PAD.n5554 0.0284039
R47018 PAD.n7793 PAD.n6710 0.0284039
R47019 PAD.n7149 PAD.n6710 0.0284039
R47020 PAD.n7529 PAD.n7150 0.0284039
R47021 PAD.n7522 PAD.n7150 0.0284039
R47022 PAD.n7205 PAD.n5203 0.0284039
R47023 PAD.n7821 PAD.n5203 0.0284039
R47024 PAD.n7827 PAD.n5189 0.0284039
R47025 PAD.n8176 PAD.n5189 0.0284039
R47026 PAD.n8182 PAD.n4838 0.0284039
R47027 PAD.n8196 PAD.n4838 0.0284039
R47028 PAD.n8203 PAD.n4833 0.0284039
R47029 PAD.n8206 PAD.n4672 0.0284039
R47030 PAD.n8411 PAD.n4672 0.0284039
R47031 PAD.n8418 PAD.n4318 0.0284039
R47032 PAD.n8432 PAD.n4318 0.0284039
R47033 PAD.n8455 PAD.n3976 0.0284039
R47034 PAD.n8456 PAD.n8455 0.0284039
R47035 PAD.n8480 PAD.n3632 0.0284039
R47036 PAD.n8481 PAD.n8480 0.0284039
R47037 PAD.n8504 PAD.n3286 0.0284039
R47038 PAD.n8507 PAD.n2902 0.0284039
R47039 PAD.n8823 PAD.n2902 0.0284039
R47040 PAD.n8830 PAD.n2893 0.0284039
R47041 PAD.n8830 PAD.n2895 0.0284039
R47042 PAD.n9130 PAD.n2493 0.0284039
R47043 PAD.n9153 PAD.n2493 0.0284039
R47044 PAD.n9159 PAD.n2145 0.0284039
R47045 PAD.n9177 PAD.n2145 0.0284039
R47046 PAD.n9183 PAD.n2044 0.0284039
R47047 PAD.n9447 PAD.n2044 0.0284039
R47048 PAD.n9454 PAD.n2038 0.0284039
R47049 PAD.n9714 PAD.n1937 0.0284039
R47050 PAD.n9720 PAD.n1937 0.0284039
R47051 PAD.n9734 PAD.n1587 0.0284039
R47052 PAD.n9740 PAD.n1587 0.0284039
R47053 PAD.n10000 PAD.n1484 0.0284039
R47054 PAD.n10006 PAD.n1484 0.0284039
R47055 PAD.n10018 PAD.n1133 0.0284039
R47056 PAD.n10360 PAD.n1133 0.0284039
R47057 PAD.n10375 PAD.n1117 0.0284039
R47058 PAD.n10378 PAD.n775 0.0284039
R47059 PAD.n10399 PAD.n775 0.0284039
R47060 PAD.n10406 PAD.n424 0.0284039
R47061 PAD.n10703 PAD.n424 0.0284039
R47062 PAD.n10706 PAD.n30 0.0284039
R47063 PAD.n10729 PAD.n30 0.0284039
R47064 PAD.n11531 PAD.n22 0.0284039
R47065 PAD.n11531 PAD.n23 0.0284039
R47066 PAD.n11524 PAD.n10739 0.0284039
R47067 PAD.n11502 PAD.n10739 0.0284039
R47068 PAD.n9452 PAD.n1939 0.028175
R47069 PAD.n10357 PAD.n10356 0.028175
R47070 PAD.n6707 PAD.n5556 0.0278144
R47071 PAD.n6709 PAD.n5554 0.0278144
R47072 PAD.n8485 PAD.n8484 0.027725
R47073 PAD.n8506 PAD.n8505 0.0274214
R47074 PAD.n8504 PAD.n2996 0.0274214
R47075 PAD.n7798 PAD.n6704 0.027275
R47076 PAD.n2043 PAD.n2039 0.0270284
R47077 PAD.n10377 PAD.n10376 0.0270284
R47078 PAD.n2045 PAD.n2038 0.0270284
R47079 PAD.n10375 PAD.n827 0.0270284
R47080 PAD.n8201 PAD.n4834 0.0266354
R47081 PAD.n4839 PAD.n4833 0.0266354
R47082 PAD.n7154 PAD.n7153 0.025925
R47083 PAD.n7268 PAD.n7155 0.0259118
R47084 PAD.n10732 PAD.n26 0.0259118
R47085 PAD.n10710 PAD.n10709 0.0259118
R47086 PAD.n10402 PAD.n772 0.0259118
R47087 PAD.n10382 PAD.n10381 0.0259118
R47088 PAD.n10357 PAD.n10355 0.0259118
R47089 PAD.n1296 PAD.n1137 0.0259118
R47090 PAD.n9992 PAD.n1486 0.0259118
R47091 PAD.n1683 PAD.n1589 0.0259118
R47092 PAD.n9706 PAD.n1939 0.0259118
R47093 PAD.n9450 PAD.n2040 0.0259118
R47094 PAD.n9180 PAD.n2142 0.0259118
R47095 PAD.n9156 PAD.n2490 0.0259118
R47096 PAD.n9134 PAD.n9133 0.0259118
R47097 PAD.n8826 PAD.n2898 0.0259118
R47098 PAD.n8511 PAD.n8510 0.0259118
R47099 PAD.n8486 PAD.n8485 0.0259118
R47100 PAD.n8462 PAD.n8461 0.0259118
R47101 PAD.n8438 PAD.n8437 0.0259118
R47102 PAD.n8414 PAD.n4669 0.0259118
R47103 PAD.n8210 PAD.n8209 0.0259118
R47104 PAD.n8199 PAD.n4835 0.0259118
R47105 PAD.n8179 PAD.n5186 0.0259118
R47106 PAD.n7824 PAD.n5200 0.0259118
R47107 PAD.n7154 PAD.n7147 0.0259118
R47108 PAD.n7796 PAD.n6705 0.0259118
R47109 PAD.n6704 PAD.n5557 0.0259118
R47110 PAD.n11527 PAD.n10734 0.0259118
R47111 PAD.n6377 PAD.n5951 0.0259118
R47112 PAD.n8826 PAD.n8825 0.025475
R47113 PAD.n11527 PAD.n11526 0.025475
R47114 PAD.n11106 PAD.n11104 0.0251375
R47115 PAD.n11353 PAD.n11093 0.0251375
R47116 PAD.n11352 PAD.n11091 0.0251375
R47117 PAD.n6226 PAD.n5959 0.0251375
R47118 PAD.n6225 PAD.n5957 0.0251375
R47119 PAD.n6034 PAD.n5969 0.0251375
R47120 PAD.n8202 PAD.n4831 0.0250633
R47121 PAD.n8204 PAD.n8203 0.0250633
R47122 PAD.n9181 PAD.n9180 0.025025
R47123 PAD.n10402 PAD.n10401 0.025025
R47124 PAD.n9453 PAD.n1940 0.0246703
R47125 PAD.n1136 PAD.n1116 0.0246703
R47126 PAD.n9454 PAD.n1941 0.0246703
R47127 PAD.n1134 PAD.n1117 0.0246703
R47128 PAD.n8180 PAD.n8179 0.024575
R47129 PAD.n3631 PAD.n3285 0.0242773
R47130 PAD.n3341 PAD.n3286 0.0242773
R47131 PAD.n7799 PAD.n5555 0.0238843
R47132 PAD.n7800 PAD.n5553 0.0238843
R47133 PAD.n7811 PAD.n7808 0.0228122
R47134 PAD.n8414 PAD.n8413 0.022775
R47135 PAD.n7152 PAD.n7148 0.0227052
R47136 PAD.n7530 PAD.n7149 0.0227052
R47137 PAD.n9718 PAD.n1589 0.022325
R47138 PAD.n10020 PAD.n1137 0.022325
R47139 PAD.n8824 PAD.n2901 0.0223122
R47140 PAD.n11525 PAD.n10736 0.0223122
R47141 PAD.n8823 PAD.n2903 0.0223122
R47142 PAD.n11524 PAD.n10738 0.0223122
R47143 PAD.n13 PAD.n12 0.0221339
R47144 PAD.n9182 PAD.n2141 0.0219192
R47145 PAD.n10400 PAD.n437 0.0219192
R47146 PAD.n9183 PAD.n2140 0.0219192
R47147 PAD.n10399 PAD.n436 0.0219192
R47148 PAD.n8461 PAD.n8460 0.021875
R47149 PAD.n11539 PAD.n13 0.0216978
R47150 PAD.n8181 PAD.n5185 0.0215262
R47151 PAD.n8182 PAD.n5184 0.0215262
R47152 PAD.n6377 PAD.n5953 0.021425
R47153 PAD.n7811 PAD.n7810 0.0210195
R47154 PAD.n7524 PAD.n7155 0.020075
R47155 PAD.n8412 PAD.n4335 0.0199541
R47156 PAD.n8411 PAD.n4334 0.0199541
R47157 PAD.n117 PAD.n116 0.019716
R47158 PAD.n124 PAD.n73 0.019716
R47159 PAD.n125 PAD.n124 0.019716
R47160 PAD.n130 PAD.n72 0.019716
R47161 PAD.n130 PAD.n129 0.019716
R47162 PAD.n136 PAD.n71 0.019716
R47163 PAD.n137 PAD.n136 0.019716
R47164 PAD.n142 PAD.n70 0.019716
R47165 PAD.n142 PAD.n141 0.019716
R47166 PAD.n148 PAD.n69 0.019716
R47167 PAD.n149 PAD.n148 0.019716
R47168 PAD.n154 PAD.n68 0.019716
R47169 PAD.n154 PAD.n153 0.019716
R47170 PAD.n160 PAD.n67 0.019716
R47171 PAD.n161 PAD.n160 0.019716
R47172 PAD.n166 PAD.n66 0.019716
R47173 PAD.n166 PAD.n165 0.019716
R47174 PAD.n172 PAD.n65 0.019716
R47175 PAD.n173 PAD.n172 0.019716
R47176 PAD.n178 PAD.n64 0.019716
R47177 PAD.n178 PAD.n177 0.019716
R47178 PAD.n184 PAD.n63 0.019716
R47179 PAD.n185 PAD.n184 0.019716
R47180 PAD.n190 PAD.n62 0.019716
R47181 PAD.n190 PAD.n189 0.019716
R47182 PAD.n196 PAD.n61 0.019716
R47183 PAD.n197 PAD.n196 0.019716
R47184 PAD.n202 PAD.n60 0.019716
R47185 PAD.n202 PAD.n201 0.019716
R47186 PAD.n208 PAD.n59 0.019716
R47187 PAD.n209 PAD.n208 0.019716
R47188 PAD.n214 PAD.n58 0.019716
R47189 PAD.n214 PAD.n213 0.019716
R47190 PAD.n220 PAD.n57 0.019716
R47191 PAD.n221 PAD.n220 0.019716
R47192 PAD.n226 PAD.n56 0.019716
R47193 PAD.n226 PAD.n225 0.019716
R47194 PAD.n232 PAD.n55 0.019716
R47195 PAD.n233 PAD.n232 0.019716
R47196 PAD.n238 PAD.n54 0.019716
R47197 PAD.n238 PAD.n237 0.019716
R47198 PAD.n244 PAD.n53 0.019716
R47199 PAD.n245 PAD.n244 0.019716
R47200 PAD.n250 PAD.n52 0.019716
R47201 PAD.n250 PAD.n249 0.019716
R47202 PAD.n256 PAD.n51 0.019716
R47203 PAD.n257 PAD.n256 0.019716
R47204 PAD.n262 PAD.n50 0.019716
R47205 PAD.n262 PAD.n261 0.019716
R47206 PAD.n268 PAD.n49 0.019716
R47207 PAD.n269 PAD.n268 0.019716
R47208 PAD.n274 PAD.n48 0.019716
R47209 PAD.n274 PAD.n273 0.019716
R47210 PAD.n280 PAD.n47 0.019716
R47211 PAD.n281 PAD.n280 0.019716
R47212 PAD.n286 PAD.n46 0.019716
R47213 PAD.n286 PAD.n285 0.019716
R47214 PAD.n292 PAD.n45 0.019716
R47215 PAD.n293 PAD.n292 0.019716
R47216 PAD.n298 PAD.n44 0.019716
R47217 PAD.n298 PAD.n297 0.019716
R47218 PAD.n304 PAD.n43 0.019716
R47219 PAD.n305 PAD.n304 0.019716
R47220 PAD.n310 PAD.n42 0.019716
R47221 PAD.n310 PAD.n309 0.019716
R47222 PAD.n316 PAD.n41 0.019716
R47223 PAD.n317 PAD.n316 0.019716
R47224 PAD.n322 PAD.n40 0.019716
R47225 PAD.n322 PAD.n321 0.019716
R47226 PAD.n328 PAD.n39 0.019716
R47227 PAD.n329 PAD.n328 0.019716
R47228 PAD.n334 PAD.n38 0.019716
R47229 PAD.n334 PAD.n333 0.019716
R47230 PAD.n340 PAD.n37 0.019716
R47231 PAD.n341 PAD.n340 0.019716
R47232 PAD.n346 PAD.n36 0.019716
R47233 PAD.n346 PAD.n345 0.019716
R47234 PAD.n352 PAD.n35 0.019716
R47235 PAD.n353 PAD.n352 0.019716
R47236 PAD.n358 PAD.n34 0.019716
R47237 PAD.n358 PAD.n357 0.019716
R47238 PAD.n364 PAD.n33 0.019716
R47239 PAD.n365 PAD.n364 0.019716
R47240 PAD.n7519 PAD.n7201 0.019716
R47241 PAD.n7512 PAD.n7511 0.019716
R47242 PAD.n7512 PAD.n7199 0.019716
R47243 PAD.n7508 PAD.n7507 0.019716
R47244 PAD.n7507 PAD.n7198 0.019716
R47245 PAD.n7501 PAD.n7500 0.019716
R47246 PAD.n7501 PAD.n7197 0.019716
R47247 PAD.n7496 PAD.n7495 0.019716
R47248 PAD.n7495 PAD.n7196 0.019716
R47249 PAD.n7489 PAD.n7488 0.019716
R47250 PAD.n7489 PAD.n7195 0.019716
R47251 PAD.n7484 PAD.n7483 0.019716
R47252 PAD.n7483 PAD.n7194 0.019716
R47253 PAD.n7477 PAD.n7476 0.019716
R47254 PAD.n7477 PAD.n7193 0.019716
R47255 PAD.n7472 PAD.n7471 0.019716
R47256 PAD.n7471 PAD.n7192 0.019716
R47257 PAD.n7465 PAD.n7464 0.019716
R47258 PAD.n7465 PAD.n7191 0.019716
R47259 PAD.n7460 PAD.n7459 0.019716
R47260 PAD.n7459 PAD.n7190 0.019716
R47261 PAD.n7453 PAD.n7452 0.019716
R47262 PAD.n7453 PAD.n7189 0.019716
R47263 PAD.n7448 PAD.n7447 0.019716
R47264 PAD.n7447 PAD.n7188 0.019716
R47265 PAD.n7441 PAD.n7440 0.019716
R47266 PAD.n7441 PAD.n7187 0.019716
R47267 PAD.n7436 PAD.n7435 0.019716
R47268 PAD.n7435 PAD.n7186 0.019716
R47269 PAD.n7429 PAD.n7428 0.019716
R47270 PAD.n7429 PAD.n7185 0.019716
R47271 PAD.n7424 PAD.n7423 0.019716
R47272 PAD.n7423 PAD.n7184 0.019716
R47273 PAD.n7417 PAD.n7416 0.019716
R47274 PAD.n7417 PAD.n7183 0.019716
R47275 PAD.n7412 PAD.n7411 0.019716
R47276 PAD.n7411 PAD.n7182 0.019716
R47277 PAD.n7405 PAD.n7404 0.019716
R47278 PAD.n7405 PAD.n7181 0.019716
R47279 PAD.n7400 PAD.n7399 0.019716
R47280 PAD.n7399 PAD.n7180 0.019716
R47281 PAD.n7393 PAD.n7392 0.019716
R47282 PAD.n7393 PAD.n7179 0.019716
R47283 PAD.n7388 PAD.n7387 0.019716
R47284 PAD.n7387 PAD.n7178 0.019716
R47285 PAD.n7381 PAD.n7380 0.019716
R47286 PAD.n7381 PAD.n7177 0.019716
R47287 PAD.n7376 PAD.n7375 0.019716
R47288 PAD.n7375 PAD.n7176 0.019716
R47289 PAD.n7369 PAD.n7368 0.019716
R47290 PAD.n7369 PAD.n7175 0.019716
R47291 PAD.n7364 PAD.n7363 0.019716
R47292 PAD.n7363 PAD.n7174 0.019716
R47293 PAD.n7357 PAD.n7356 0.019716
R47294 PAD.n7357 PAD.n7173 0.019716
R47295 PAD.n7352 PAD.n7351 0.019716
R47296 PAD.n7351 PAD.n7172 0.019716
R47297 PAD.n7345 PAD.n7344 0.019716
R47298 PAD.n7345 PAD.n7171 0.019716
R47299 PAD.n7340 PAD.n7339 0.019716
R47300 PAD.n7339 PAD.n7170 0.019716
R47301 PAD.n7333 PAD.n7332 0.019716
R47302 PAD.n7333 PAD.n7169 0.019716
R47303 PAD.n7328 PAD.n7327 0.019716
R47304 PAD.n7327 PAD.n7168 0.019716
R47305 PAD.n7321 PAD.n7320 0.019716
R47306 PAD.n7321 PAD.n7167 0.019716
R47307 PAD.n7316 PAD.n7315 0.019716
R47308 PAD.n7315 PAD.n7166 0.019716
R47309 PAD.n7309 PAD.n7308 0.019716
R47310 PAD.n7309 PAD.n7165 0.019716
R47311 PAD.n7304 PAD.n7303 0.019716
R47312 PAD.n7303 PAD.n7164 0.019716
R47313 PAD.n7297 PAD.n7296 0.019716
R47314 PAD.n7297 PAD.n7163 0.019716
R47315 PAD.n7292 PAD.n7291 0.019716
R47316 PAD.n7291 PAD.n7162 0.019716
R47317 PAD.n7285 PAD.n7284 0.019716
R47318 PAD.n7285 PAD.n7161 0.019716
R47319 PAD.n7280 PAD.n7279 0.019716
R47320 PAD.n7279 PAD.n7160 0.019716
R47321 PAD.n7273 PAD.n7272 0.019716
R47322 PAD.n7273 PAD.n7159 0.019716
R47323 PAD.n10693 PAD.n10692 0.019716
R47324 PAD.n10417 PAD.n414 0.019716
R47325 PAD.n10417 PAD.n10416 0.019716
R47326 PAD.n10686 PAD.n413 0.019716
R47327 PAD.n10686 PAD.n10685 0.019716
R47328 PAD.n10422 PAD.n412 0.019716
R47329 PAD.n10422 PAD.n10421 0.019716
R47330 PAD.n10677 PAD.n411 0.019716
R47331 PAD.n10677 PAD.n10676 0.019716
R47332 PAD.n10427 PAD.n410 0.019716
R47333 PAD.n10427 PAD.n10426 0.019716
R47334 PAD.n10668 PAD.n409 0.019716
R47335 PAD.n10668 PAD.n10667 0.019716
R47336 PAD.n10432 PAD.n408 0.019716
R47337 PAD.n10432 PAD.n10431 0.019716
R47338 PAD.n10659 PAD.n407 0.019716
R47339 PAD.n10659 PAD.n10658 0.019716
R47340 PAD.n10437 PAD.n406 0.019716
R47341 PAD.n10437 PAD.n10436 0.019716
R47342 PAD.n10650 PAD.n405 0.019716
R47343 PAD.n10650 PAD.n10649 0.019716
R47344 PAD.n10442 PAD.n404 0.019716
R47345 PAD.n10442 PAD.n10441 0.019716
R47346 PAD.n10641 PAD.n403 0.019716
R47347 PAD.n10641 PAD.n10640 0.019716
R47348 PAD.n10447 PAD.n402 0.019716
R47349 PAD.n10447 PAD.n10446 0.019716
R47350 PAD.n10632 PAD.n401 0.019716
R47351 PAD.n10632 PAD.n10631 0.019716
R47352 PAD.n10452 PAD.n400 0.019716
R47353 PAD.n10452 PAD.n10451 0.019716
R47354 PAD.n10623 PAD.n399 0.019716
R47355 PAD.n10623 PAD.n10622 0.019716
R47356 PAD.n10457 PAD.n398 0.019716
R47357 PAD.n10457 PAD.n10456 0.019716
R47358 PAD.n10614 PAD.n397 0.019716
R47359 PAD.n10614 PAD.n10613 0.019716
R47360 PAD.n10462 PAD.n396 0.019716
R47361 PAD.n10462 PAD.n10461 0.019716
R47362 PAD.n10605 PAD.n395 0.019716
R47363 PAD.n10605 PAD.n10604 0.019716
R47364 PAD.n10467 PAD.n394 0.019716
R47365 PAD.n10467 PAD.n10466 0.019716
R47366 PAD.n10596 PAD.n393 0.019716
R47367 PAD.n10596 PAD.n10595 0.019716
R47368 PAD.n10472 PAD.n392 0.019716
R47369 PAD.n10472 PAD.n10471 0.019716
R47370 PAD.n10587 PAD.n391 0.019716
R47371 PAD.n10587 PAD.n10586 0.019716
R47372 PAD.n10477 PAD.n390 0.019716
R47373 PAD.n10477 PAD.n10476 0.019716
R47374 PAD.n10578 PAD.n389 0.019716
R47375 PAD.n10578 PAD.n10577 0.019716
R47376 PAD.n10482 PAD.n388 0.019716
R47377 PAD.n10482 PAD.n10481 0.019716
R47378 PAD.n10569 PAD.n387 0.019716
R47379 PAD.n10569 PAD.n10568 0.019716
R47380 PAD.n10487 PAD.n386 0.019716
R47381 PAD.n10487 PAD.n10486 0.019716
R47382 PAD.n10560 PAD.n385 0.019716
R47383 PAD.n10560 PAD.n10559 0.019716
R47384 PAD.n10492 PAD.n384 0.019716
R47385 PAD.n10492 PAD.n10491 0.019716
R47386 PAD.n10551 PAD.n383 0.019716
R47387 PAD.n10551 PAD.n10550 0.019716
R47388 PAD.n10497 PAD.n382 0.019716
R47389 PAD.n10497 PAD.n10496 0.019716
R47390 PAD.n10542 PAD.n381 0.019716
R47391 PAD.n10542 PAD.n10541 0.019716
R47392 PAD.n10502 PAD.n380 0.019716
R47393 PAD.n10502 PAD.n10501 0.019716
R47394 PAD.n10533 PAD.n379 0.019716
R47395 PAD.n10533 PAD.n10532 0.019716
R47396 PAD.n10507 PAD.n378 0.019716
R47397 PAD.n10507 PAD.n10506 0.019716
R47398 PAD.n10524 PAD.n377 0.019716
R47399 PAD.n10524 PAD.n10523 0.019716
R47400 PAD.n10512 PAD.n376 0.019716
R47401 PAD.n10512 PAD.n10511 0.019716
R47402 PAD.n10515 PAD.n375 0.019716
R47403 PAD.n10515 PAD.n10514 0.019716
R47404 PAD.n10713 PAD.n374 0.019716
R47405 PAD.n10714 PAD.n10713 0.019716
R47406 PAD.n525 PAD.n524 0.019716
R47407 PAD.n529 PAD.n526 0.019716
R47408 PAD.n529 PAD.n528 0.019716
R47409 PAD.n535 PAD.n517 0.019716
R47410 PAD.n536 PAD.n535 0.019716
R47411 PAD.n541 PAD.n538 0.019716
R47412 PAD.n541 PAD.n540 0.019716
R47413 PAD.n547 PAD.n513 0.019716
R47414 PAD.n548 PAD.n547 0.019716
R47415 PAD.n553 PAD.n550 0.019716
R47416 PAD.n553 PAD.n552 0.019716
R47417 PAD.n559 PAD.n509 0.019716
R47418 PAD.n560 PAD.n559 0.019716
R47419 PAD.n565 PAD.n562 0.019716
R47420 PAD.n565 PAD.n564 0.019716
R47421 PAD.n571 PAD.n505 0.019716
R47422 PAD.n572 PAD.n571 0.019716
R47423 PAD.n577 PAD.n574 0.019716
R47424 PAD.n577 PAD.n576 0.019716
R47425 PAD.n583 PAD.n501 0.019716
R47426 PAD.n584 PAD.n583 0.019716
R47427 PAD.n589 PAD.n586 0.019716
R47428 PAD.n589 PAD.n588 0.019716
R47429 PAD.n595 PAD.n497 0.019716
R47430 PAD.n596 PAD.n595 0.019716
R47431 PAD.n601 PAD.n598 0.019716
R47432 PAD.n601 PAD.n600 0.019716
R47433 PAD.n607 PAD.n493 0.019716
R47434 PAD.n608 PAD.n607 0.019716
R47435 PAD.n613 PAD.n610 0.019716
R47436 PAD.n613 PAD.n612 0.019716
R47437 PAD.n619 PAD.n489 0.019716
R47438 PAD.n620 PAD.n619 0.019716
R47439 PAD.n625 PAD.n622 0.019716
R47440 PAD.n625 PAD.n624 0.019716
R47441 PAD.n631 PAD.n485 0.019716
R47442 PAD.n632 PAD.n631 0.019716
R47443 PAD.n637 PAD.n634 0.019716
R47444 PAD.n637 PAD.n636 0.019716
R47445 PAD.n643 PAD.n481 0.019716
R47446 PAD.n644 PAD.n643 0.019716
R47447 PAD.n649 PAD.n646 0.019716
R47448 PAD.n649 PAD.n648 0.019716
R47449 PAD.n655 PAD.n477 0.019716
R47450 PAD.n656 PAD.n655 0.019716
R47451 PAD.n661 PAD.n658 0.019716
R47452 PAD.n661 PAD.n660 0.019716
R47453 PAD.n667 PAD.n473 0.019716
R47454 PAD.n668 PAD.n667 0.019716
R47455 PAD.n673 PAD.n670 0.019716
R47456 PAD.n673 PAD.n672 0.019716
R47457 PAD.n679 PAD.n469 0.019716
R47458 PAD.n680 PAD.n679 0.019716
R47459 PAD.n685 PAD.n682 0.019716
R47460 PAD.n685 PAD.n684 0.019716
R47461 PAD.n691 PAD.n465 0.019716
R47462 PAD.n692 PAD.n691 0.019716
R47463 PAD.n697 PAD.n694 0.019716
R47464 PAD.n697 PAD.n696 0.019716
R47465 PAD.n703 PAD.n461 0.019716
R47466 PAD.n704 PAD.n703 0.019716
R47467 PAD.n709 PAD.n706 0.019716
R47468 PAD.n709 PAD.n708 0.019716
R47469 PAD.n715 PAD.n457 0.019716
R47470 PAD.n716 PAD.n715 0.019716
R47471 PAD.n721 PAD.n718 0.019716
R47472 PAD.n721 PAD.n720 0.019716
R47473 PAD.n727 PAD.n453 0.019716
R47474 PAD.n728 PAD.n727 0.019716
R47475 PAD.n733 PAD.n730 0.019716
R47476 PAD.n733 PAD.n732 0.019716
R47477 PAD.n739 PAD.n449 0.019716
R47478 PAD.n740 PAD.n739 0.019716
R47479 PAD.n745 PAD.n742 0.019716
R47480 PAD.n745 PAD.n744 0.019716
R47481 PAD.n751 PAD.n445 0.019716
R47482 PAD.n752 PAD.n751 0.019716
R47483 PAD.n757 PAD.n754 0.019716
R47484 PAD.n757 PAD.n756 0.019716
R47485 PAD.n764 PAD.n441 0.019716
R47486 PAD.n765 PAD.n764 0.019716
R47487 PAD.n768 PAD.n767 0.019716
R47488 PAD.n769 PAD.n768 0.019716
R47489 PAD.n870 PAD.n869 0.019716
R47490 PAD.n877 PAD.n823 0.019716
R47491 PAD.n878 PAD.n877 0.019716
R47492 PAD.n883 PAD.n822 0.019716
R47493 PAD.n883 PAD.n882 0.019716
R47494 PAD.n889 PAD.n821 0.019716
R47495 PAD.n890 PAD.n889 0.019716
R47496 PAD.n895 PAD.n820 0.019716
R47497 PAD.n895 PAD.n894 0.019716
R47498 PAD.n901 PAD.n819 0.019716
R47499 PAD.n902 PAD.n901 0.019716
R47500 PAD.n907 PAD.n818 0.019716
R47501 PAD.n907 PAD.n906 0.019716
R47502 PAD.n913 PAD.n817 0.019716
R47503 PAD.n914 PAD.n913 0.019716
R47504 PAD.n919 PAD.n816 0.019716
R47505 PAD.n919 PAD.n918 0.019716
R47506 PAD.n925 PAD.n815 0.019716
R47507 PAD.n926 PAD.n925 0.019716
R47508 PAD.n931 PAD.n814 0.019716
R47509 PAD.n931 PAD.n930 0.019716
R47510 PAD.n937 PAD.n813 0.019716
R47511 PAD.n938 PAD.n937 0.019716
R47512 PAD.n943 PAD.n812 0.019716
R47513 PAD.n943 PAD.n942 0.019716
R47514 PAD.n949 PAD.n811 0.019716
R47515 PAD.n950 PAD.n949 0.019716
R47516 PAD.n955 PAD.n810 0.019716
R47517 PAD.n955 PAD.n954 0.019716
R47518 PAD.n961 PAD.n809 0.019716
R47519 PAD.n962 PAD.n961 0.019716
R47520 PAD.n967 PAD.n808 0.019716
R47521 PAD.n967 PAD.n966 0.019716
R47522 PAD.n973 PAD.n807 0.019716
R47523 PAD.n974 PAD.n973 0.019716
R47524 PAD.n979 PAD.n806 0.019716
R47525 PAD.n979 PAD.n978 0.019716
R47526 PAD.n985 PAD.n805 0.019716
R47527 PAD.n986 PAD.n985 0.019716
R47528 PAD.n991 PAD.n804 0.019716
R47529 PAD.n991 PAD.n990 0.019716
R47530 PAD.n997 PAD.n803 0.019716
R47531 PAD.n998 PAD.n997 0.019716
R47532 PAD.n1003 PAD.n802 0.019716
R47533 PAD.n1003 PAD.n1002 0.019716
R47534 PAD.n1009 PAD.n801 0.019716
R47535 PAD.n1010 PAD.n1009 0.019716
R47536 PAD.n1015 PAD.n800 0.019716
R47537 PAD.n1015 PAD.n1014 0.019716
R47538 PAD.n1021 PAD.n799 0.019716
R47539 PAD.n1022 PAD.n1021 0.019716
R47540 PAD.n1027 PAD.n798 0.019716
R47541 PAD.n1027 PAD.n1026 0.019716
R47542 PAD.n1033 PAD.n797 0.019716
R47543 PAD.n1034 PAD.n1033 0.019716
R47544 PAD.n1039 PAD.n796 0.019716
R47545 PAD.n1039 PAD.n1038 0.019716
R47546 PAD.n1045 PAD.n795 0.019716
R47547 PAD.n1046 PAD.n1045 0.019716
R47548 PAD.n1051 PAD.n794 0.019716
R47549 PAD.n1051 PAD.n1050 0.019716
R47550 PAD.n1057 PAD.n793 0.019716
R47551 PAD.n1058 PAD.n1057 0.019716
R47552 PAD.n1063 PAD.n792 0.019716
R47553 PAD.n1063 PAD.n1062 0.019716
R47554 PAD.n1069 PAD.n791 0.019716
R47555 PAD.n1070 PAD.n1069 0.019716
R47556 PAD.n1075 PAD.n790 0.019716
R47557 PAD.n1075 PAD.n1074 0.019716
R47558 PAD.n1081 PAD.n789 0.019716
R47559 PAD.n1082 PAD.n1081 0.019716
R47560 PAD.n1087 PAD.n788 0.019716
R47561 PAD.n1087 PAD.n1086 0.019716
R47562 PAD.n1093 PAD.n787 0.019716
R47563 PAD.n1094 PAD.n1093 0.019716
R47564 PAD.n1099 PAD.n786 0.019716
R47565 PAD.n1099 PAD.n1098 0.019716
R47566 PAD.n1105 PAD.n785 0.019716
R47567 PAD.n1106 PAD.n1105 0.019716
R47568 PAD.n1111 PAD.n784 0.019716
R47569 PAD.n1111 PAD.n1110 0.019716
R47570 PAD.n10385 PAD.n783 0.019716
R47571 PAD.n10386 PAD.n10385 0.019716
R47572 PAD.n10108 PAD.n10107 0.019716
R47573 PAD.n10112 PAD.n10109 0.019716
R47574 PAD.n10112 PAD.n10111 0.019716
R47575 PAD.n10118 PAD.n10101 0.019716
R47576 PAD.n10119 PAD.n10118 0.019716
R47577 PAD.n10124 PAD.n10121 0.019716
R47578 PAD.n10124 PAD.n10123 0.019716
R47579 PAD.n10130 PAD.n10097 0.019716
R47580 PAD.n10131 PAD.n10130 0.019716
R47581 PAD.n10136 PAD.n10133 0.019716
R47582 PAD.n10136 PAD.n10135 0.019716
R47583 PAD.n10142 PAD.n10093 0.019716
R47584 PAD.n10143 PAD.n10142 0.019716
R47585 PAD.n10148 PAD.n10145 0.019716
R47586 PAD.n10148 PAD.n10147 0.019716
R47587 PAD.n10154 PAD.n10089 0.019716
R47588 PAD.n10155 PAD.n10154 0.019716
R47589 PAD.n10160 PAD.n10157 0.019716
R47590 PAD.n10160 PAD.n10159 0.019716
R47591 PAD.n10166 PAD.n10085 0.019716
R47592 PAD.n10167 PAD.n10166 0.019716
R47593 PAD.n10172 PAD.n10169 0.019716
R47594 PAD.n10172 PAD.n10171 0.019716
R47595 PAD.n10178 PAD.n10081 0.019716
R47596 PAD.n10179 PAD.n10178 0.019716
R47597 PAD.n10184 PAD.n10181 0.019716
R47598 PAD.n10184 PAD.n10183 0.019716
R47599 PAD.n10190 PAD.n10077 0.019716
R47600 PAD.n10191 PAD.n10190 0.019716
R47601 PAD.n10196 PAD.n10193 0.019716
R47602 PAD.n10196 PAD.n10195 0.019716
R47603 PAD.n10202 PAD.n10073 0.019716
R47604 PAD.n10203 PAD.n10202 0.019716
R47605 PAD.n10208 PAD.n10205 0.019716
R47606 PAD.n10208 PAD.n10207 0.019716
R47607 PAD.n10214 PAD.n10069 0.019716
R47608 PAD.n10215 PAD.n10214 0.019716
R47609 PAD.n10220 PAD.n10217 0.019716
R47610 PAD.n10220 PAD.n10219 0.019716
R47611 PAD.n10226 PAD.n10065 0.019716
R47612 PAD.n10227 PAD.n10226 0.019716
R47613 PAD.n10232 PAD.n10229 0.019716
R47614 PAD.n10232 PAD.n10231 0.019716
R47615 PAD.n10238 PAD.n10061 0.019716
R47616 PAD.n10239 PAD.n10238 0.019716
R47617 PAD.n10244 PAD.n10241 0.019716
R47618 PAD.n10244 PAD.n10243 0.019716
R47619 PAD.n10250 PAD.n10057 0.019716
R47620 PAD.n10251 PAD.n10250 0.019716
R47621 PAD.n10256 PAD.n10253 0.019716
R47622 PAD.n10256 PAD.n10255 0.019716
R47623 PAD.n10262 PAD.n10053 0.019716
R47624 PAD.n10263 PAD.n10262 0.019716
R47625 PAD.n10268 PAD.n10265 0.019716
R47626 PAD.n10268 PAD.n10267 0.019716
R47627 PAD.n10274 PAD.n10049 0.019716
R47628 PAD.n10275 PAD.n10274 0.019716
R47629 PAD.n10280 PAD.n10277 0.019716
R47630 PAD.n10280 PAD.n10279 0.019716
R47631 PAD.n10286 PAD.n10045 0.019716
R47632 PAD.n10287 PAD.n10286 0.019716
R47633 PAD.n10292 PAD.n10289 0.019716
R47634 PAD.n10292 PAD.n10291 0.019716
R47635 PAD.n10298 PAD.n10041 0.019716
R47636 PAD.n10299 PAD.n10298 0.019716
R47637 PAD.n10304 PAD.n10301 0.019716
R47638 PAD.n10304 PAD.n10303 0.019716
R47639 PAD.n10310 PAD.n10037 0.019716
R47640 PAD.n10311 PAD.n10310 0.019716
R47641 PAD.n10316 PAD.n10313 0.019716
R47642 PAD.n10316 PAD.n10315 0.019716
R47643 PAD.n10322 PAD.n10033 0.019716
R47644 PAD.n10323 PAD.n10322 0.019716
R47645 PAD.n10328 PAD.n10325 0.019716
R47646 PAD.n10328 PAD.n10327 0.019716
R47647 PAD.n10334 PAD.n10029 0.019716
R47648 PAD.n10335 PAD.n10334 0.019716
R47649 PAD.n10340 PAD.n10337 0.019716
R47650 PAD.n10340 PAD.n10339 0.019716
R47651 PAD.n10347 PAD.n10025 0.019716
R47652 PAD.n10348 PAD.n10347 0.019716
R47653 PAD.n10351 PAD.n10350 0.019716
R47654 PAD.n10352 PAD.n10351 0.019716
R47655 PAD.n1482 PAD.n1190 0.019716
R47656 PAD.n1192 PAD.n1191 0.019716
R47657 PAD.n1192 PAD.n1189 0.019716
R47658 PAD.n1473 PAD.n1472 0.019716
R47659 PAD.n1472 PAD.n1188 0.019716
R47660 PAD.n1197 PAD.n1196 0.019716
R47661 PAD.n1196 PAD.n1187 0.019716
R47662 PAD.n1464 PAD.n1463 0.019716
R47663 PAD.n1463 PAD.n1186 0.019716
R47664 PAD.n1202 PAD.n1201 0.019716
R47665 PAD.n1201 PAD.n1185 0.019716
R47666 PAD.n1455 PAD.n1454 0.019716
R47667 PAD.n1454 PAD.n1184 0.019716
R47668 PAD.n1207 PAD.n1206 0.019716
R47669 PAD.n1206 PAD.n1183 0.019716
R47670 PAD.n1446 PAD.n1445 0.019716
R47671 PAD.n1445 PAD.n1182 0.019716
R47672 PAD.n1212 PAD.n1211 0.019716
R47673 PAD.n1211 PAD.n1181 0.019716
R47674 PAD.n1437 PAD.n1436 0.019716
R47675 PAD.n1436 PAD.n1180 0.019716
R47676 PAD.n1217 PAD.n1216 0.019716
R47677 PAD.n1216 PAD.n1179 0.019716
R47678 PAD.n1428 PAD.n1427 0.019716
R47679 PAD.n1427 PAD.n1178 0.019716
R47680 PAD.n1222 PAD.n1221 0.019716
R47681 PAD.n1221 PAD.n1177 0.019716
R47682 PAD.n1419 PAD.n1418 0.019716
R47683 PAD.n1418 PAD.n1176 0.019716
R47684 PAD.n1227 PAD.n1226 0.019716
R47685 PAD.n1226 PAD.n1175 0.019716
R47686 PAD.n1410 PAD.n1409 0.019716
R47687 PAD.n1409 PAD.n1174 0.019716
R47688 PAD.n1232 PAD.n1231 0.019716
R47689 PAD.n1231 PAD.n1173 0.019716
R47690 PAD.n1401 PAD.n1400 0.019716
R47691 PAD.n1400 PAD.n1172 0.019716
R47692 PAD.n1237 PAD.n1236 0.019716
R47693 PAD.n1236 PAD.n1171 0.019716
R47694 PAD.n1392 PAD.n1391 0.019716
R47695 PAD.n1391 PAD.n1170 0.019716
R47696 PAD.n1242 PAD.n1241 0.019716
R47697 PAD.n1241 PAD.n1169 0.019716
R47698 PAD.n1383 PAD.n1382 0.019716
R47699 PAD.n1382 PAD.n1168 0.019716
R47700 PAD.n1247 PAD.n1246 0.019716
R47701 PAD.n1246 PAD.n1167 0.019716
R47702 PAD.n1374 PAD.n1373 0.019716
R47703 PAD.n1373 PAD.n1166 0.019716
R47704 PAD.n1252 PAD.n1251 0.019716
R47705 PAD.n1251 PAD.n1165 0.019716
R47706 PAD.n1365 PAD.n1364 0.019716
R47707 PAD.n1364 PAD.n1164 0.019716
R47708 PAD.n1257 PAD.n1256 0.019716
R47709 PAD.n1256 PAD.n1163 0.019716
R47710 PAD.n1356 PAD.n1355 0.019716
R47711 PAD.n1355 PAD.n1162 0.019716
R47712 PAD.n1262 PAD.n1261 0.019716
R47713 PAD.n1261 PAD.n1161 0.019716
R47714 PAD.n1347 PAD.n1346 0.019716
R47715 PAD.n1346 PAD.n1160 0.019716
R47716 PAD.n1267 PAD.n1266 0.019716
R47717 PAD.n1266 PAD.n1159 0.019716
R47718 PAD.n1338 PAD.n1337 0.019716
R47719 PAD.n1337 PAD.n1158 0.019716
R47720 PAD.n1272 PAD.n1271 0.019716
R47721 PAD.n1271 PAD.n1157 0.019716
R47722 PAD.n1329 PAD.n1328 0.019716
R47723 PAD.n1328 PAD.n1156 0.019716
R47724 PAD.n1277 PAD.n1276 0.019716
R47725 PAD.n1276 PAD.n1155 0.019716
R47726 PAD.n1320 PAD.n1319 0.019716
R47727 PAD.n1319 PAD.n1154 0.019716
R47728 PAD.n1282 PAD.n1281 0.019716
R47729 PAD.n1281 PAD.n1153 0.019716
R47730 PAD.n1311 PAD.n1310 0.019716
R47731 PAD.n1310 PAD.n1152 0.019716
R47732 PAD.n1287 PAD.n1286 0.019716
R47733 PAD.n1286 PAD.n1151 0.019716
R47734 PAD.n1302 PAD.n1301 0.019716
R47735 PAD.n1301 PAD.n1150 0.019716
R47736 PAD.n1292 PAD.n1291 0.019716
R47737 PAD.n1291 PAD.n1149 0.019716
R47738 PAD.n1578 PAD.n1577 0.019716
R47739 PAD.n9754 PAD.n1530 0.019716
R47740 PAD.n9755 PAD.n9754 0.019716
R47741 PAD.n9760 PAD.n1529 0.019716
R47742 PAD.n9760 PAD.n9759 0.019716
R47743 PAD.n9766 PAD.n1528 0.019716
R47744 PAD.n9767 PAD.n9766 0.019716
R47745 PAD.n9772 PAD.n1527 0.019716
R47746 PAD.n9772 PAD.n9771 0.019716
R47747 PAD.n9778 PAD.n1526 0.019716
R47748 PAD.n9779 PAD.n9778 0.019716
R47749 PAD.n9784 PAD.n1525 0.019716
R47750 PAD.n9784 PAD.n9783 0.019716
R47751 PAD.n9790 PAD.n1524 0.019716
R47752 PAD.n9791 PAD.n9790 0.019716
R47753 PAD.n9796 PAD.n1523 0.019716
R47754 PAD.n9796 PAD.n9795 0.019716
R47755 PAD.n9802 PAD.n1522 0.019716
R47756 PAD.n9803 PAD.n9802 0.019716
R47757 PAD.n9808 PAD.n1521 0.019716
R47758 PAD.n9808 PAD.n9807 0.019716
R47759 PAD.n9814 PAD.n1520 0.019716
R47760 PAD.n9815 PAD.n9814 0.019716
R47761 PAD.n9820 PAD.n1519 0.019716
R47762 PAD.n9820 PAD.n9819 0.019716
R47763 PAD.n9826 PAD.n1518 0.019716
R47764 PAD.n9827 PAD.n9826 0.019716
R47765 PAD.n9832 PAD.n1517 0.019716
R47766 PAD.n9832 PAD.n9831 0.019716
R47767 PAD.n9838 PAD.n1516 0.019716
R47768 PAD.n9839 PAD.n9838 0.019716
R47769 PAD.n9844 PAD.n1515 0.019716
R47770 PAD.n9844 PAD.n9843 0.019716
R47771 PAD.n9850 PAD.n1514 0.019716
R47772 PAD.n9851 PAD.n9850 0.019716
R47773 PAD.n9856 PAD.n1513 0.019716
R47774 PAD.n9856 PAD.n9855 0.019716
R47775 PAD.n9862 PAD.n1512 0.019716
R47776 PAD.n9863 PAD.n9862 0.019716
R47777 PAD.n9868 PAD.n1511 0.019716
R47778 PAD.n9868 PAD.n9867 0.019716
R47779 PAD.n9874 PAD.n1510 0.019716
R47780 PAD.n9875 PAD.n9874 0.019716
R47781 PAD.n9880 PAD.n1509 0.019716
R47782 PAD.n9880 PAD.n9879 0.019716
R47783 PAD.n9886 PAD.n1508 0.019716
R47784 PAD.n9887 PAD.n9886 0.019716
R47785 PAD.n9892 PAD.n1507 0.019716
R47786 PAD.n9892 PAD.n9891 0.019716
R47787 PAD.n9898 PAD.n1506 0.019716
R47788 PAD.n9899 PAD.n9898 0.019716
R47789 PAD.n9904 PAD.n1505 0.019716
R47790 PAD.n9904 PAD.n9903 0.019716
R47791 PAD.n9910 PAD.n1504 0.019716
R47792 PAD.n9911 PAD.n9910 0.019716
R47793 PAD.n9916 PAD.n1503 0.019716
R47794 PAD.n9916 PAD.n9915 0.019716
R47795 PAD.n9922 PAD.n1502 0.019716
R47796 PAD.n9923 PAD.n9922 0.019716
R47797 PAD.n9928 PAD.n1501 0.019716
R47798 PAD.n9928 PAD.n9927 0.019716
R47799 PAD.n9934 PAD.n1500 0.019716
R47800 PAD.n9935 PAD.n9934 0.019716
R47801 PAD.n9940 PAD.n1499 0.019716
R47802 PAD.n9940 PAD.n9939 0.019716
R47803 PAD.n9946 PAD.n1498 0.019716
R47804 PAD.n9947 PAD.n9946 0.019716
R47805 PAD.n9952 PAD.n1497 0.019716
R47806 PAD.n9952 PAD.n9951 0.019716
R47807 PAD.n9958 PAD.n1496 0.019716
R47808 PAD.n9959 PAD.n9958 0.019716
R47809 PAD.n9964 PAD.n1495 0.019716
R47810 PAD.n9964 PAD.n9963 0.019716
R47811 PAD.n9970 PAD.n1494 0.019716
R47812 PAD.n9971 PAD.n9970 0.019716
R47813 PAD.n9976 PAD.n1493 0.019716
R47814 PAD.n9976 PAD.n9975 0.019716
R47815 PAD.n9982 PAD.n1492 0.019716
R47816 PAD.n9983 PAD.n9982 0.019716
R47817 PAD.n9988 PAD.n1491 0.019716
R47818 PAD.n9988 PAD.n9987 0.019716
R47819 PAD.n9995 PAD.n1490 0.019716
R47820 PAD.n9996 PAD.n9995 0.019716
R47821 PAD.n1929 PAD.n1601 0.019716
R47822 PAD.n1928 PAD.n1927 0.019716
R47823 PAD.n1927 PAD.n1926 0.019716
R47824 PAD.n1917 PAD.n1602 0.019716
R47825 PAD.n1918 PAD.n1917 0.019716
R47826 PAD.n1916 PAD.n1915 0.019716
R47827 PAD.n1915 PAD.n1914 0.019716
R47828 PAD.n1905 PAD.n1607 0.019716
R47829 PAD.n1906 PAD.n1905 0.019716
R47830 PAD.n1904 PAD.n1903 0.019716
R47831 PAD.n1903 PAD.n1902 0.019716
R47832 PAD.n1893 PAD.n1611 0.019716
R47833 PAD.n1894 PAD.n1893 0.019716
R47834 PAD.n1892 PAD.n1891 0.019716
R47835 PAD.n1891 PAD.n1890 0.019716
R47836 PAD.n1881 PAD.n1615 0.019716
R47837 PAD.n1882 PAD.n1881 0.019716
R47838 PAD.n1880 PAD.n1879 0.019716
R47839 PAD.n1879 PAD.n1878 0.019716
R47840 PAD.n1869 PAD.n1619 0.019716
R47841 PAD.n1870 PAD.n1869 0.019716
R47842 PAD.n1868 PAD.n1867 0.019716
R47843 PAD.n1867 PAD.n1866 0.019716
R47844 PAD.n1857 PAD.n1623 0.019716
R47845 PAD.n1858 PAD.n1857 0.019716
R47846 PAD.n1856 PAD.n1855 0.019716
R47847 PAD.n1855 PAD.n1854 0.019716
R47848 PAD.n1845 PAD.n1627 0.019716
R47849 PAD.n1846 PAD.n1845 0.019716
R47850 PAD.n1844 PAD.n1843 0.019716
R47851 PAD.n1843 PAD.n1842 0.019716
R47852 PAD.n1833 PAD.n1631 0.019716
R47853 PAD.n1834 PAD.n1833 0.019716
R47854 PAD.n1832 PAD.n1831 0.019716
R47855 PAD.n1831 PAD.n1830 0.019716
R47856 PAD.n1821 PAD.n1635 0.019716
R47857 PAD.n1822 PAD.n1821 0.019716
R47858 PAD.n1820 PAD.n1819 0.019716
R47859 PAD.n1819 PAD.n1818 0.019716
R47860 PAD.n1809 PAD.n1639 0.019716
R47861 PAD.n1810 PAD.n1809 0.019716
R47862 PAD.n1808 PAD.n1807 0.019716
R47863 PAD.n1807 PAD.n1806 0.019716
R47864 PAD.n1797 PAD.n1643 0.019716
R47865 PAD.n1798 PAD.n1797 0.019716
R47866 PAD.n1796 PAD.n1795 0.019716
R47867 PAD.n1795 PAD.n1794 0.019716
R47868 PAD.n1785 PAD.n1647 0.019716
R47869 PAD.n1786 PAD.n1785 0.019716
R47870 PAD.n1784 PAD.n1783 0.019716
R47871 PAD.n1783 PAD.n1782 0.019716
R47872 PAD.n1773 PAD.n1651 0.019716
R47873 PAD.n1774 PAD.n1773 0.019716
R47874 PAD.n1772 PAD.n1771 0.019716
R47875 PAD.n1771 PAD.n1770 0.019716
R47876 PAD.n1761 PAD.n1655 0.019716
R47877 PAD.n1762 PAD.n1761 0.019716
R47878 PAD.n1760 PAD.n1759 0.019716
R47879 PAD.n1759 PAD.n1758 0.019716
R47880 PAD.n1749 PAD.n1659 0.019716
R47881 PAD.n1750 PAD.n1749 0.019716
R47882 PAD.n1748 PAD.n1747 0.019716
R47883 PAD.n1747 PAD.n1746 0.019716
R47884 PAD.n1737 PAD.n1663 0.019716
R47885 PAD.n1738 PAD.n1737 0.019716
R47886 PAD.n1736 PAD.n1735 0.019716
R47887 PAD.n1735 PAD.n1734 0.019716
R47888 PAD.n1725 PAD.n1667 0.019716
R47889 PAD.n1726 PAD.n1725 0.019716
R47890 PAD.n1724 PAD.n1723 0.019716
R47891 PAD.n1723 PAD.n1722 0.019716
R47892 PAD.n1713 PAD.n1671 0.019716
R47893 PAD.n1714 PAD.n1713 0.019716
R47894 PAD.n1712 PAD.n1711 0.019716
R47895 PAD.n1711 PAD.n1710 0.019716
R47896 PAD.n1701 PAD.n1675 0.019716
R47897 PAD.n1702 PAD.n1701 0.019716
R47898 PAD.n1700 PAD.n1699 0.019716
R47899 PAD.n1699 PAD.n1698 0.019716
R47900 PAD.n1689 PAD.n1679 0.019716
R47901 PAD.n1690 PAD.n1689 0.019716
R47902 PAD.n1688 PAD.n1687 0.019716
R47903 PAD.n1687 PAD.n1686 0.019716
R47904 PAD.n2030 PAD.n2029 0.019716
R47905 PAD.n9468 PAD.n1983 0.019716
R47906 PAD.n9469 PAD.n9468 0.019716
R47907 PAD.n9474 PAD.n1982 0.019716
R47908 PAD.n9474 PAD.n9473 0.019716
R47909 PAD.n9480 PAD.n1981 0.019716
R47910 PAD.n9481 PAD.n9480 0.019716
R47911 PAD.n9486 PAD.n1980 0.019716
R47912 PAD.n9486 PAD.n9485 0.019716
R47913 PAD.n9492 PAD.n1979 0.019716
R47914 PAD.n9493 PAD.n9492 0.019716
R47915 PAD.n9498 PAD.n1978 0.019716
R47916 PAD.n9498 PAD.n9497 0.019716
R47917 PAD.n9504 PAD.n1977 0.019716
R47918 PAD.n9505 PAD.n9504 0.019716
R47919 PAD.n9510 PAD.n1976 0.019716
R47920 PAD.n9510 PAD.n9509 0.019716
R47921 PAD.n9516 PAD.n1975 0.019716
R47922 PAD.n9517 PAD.n9516 0.019716
R47923 PAD.n9522 PAD.n1974 0.019716
R47924 PAD.n9522 PAD.n9521 0.019716
R47925 PAD.n9528 PAD.n1973 0.019716
R47926 PAD.n9529 PAD.n9528 0.019716
R47927 PAD.n9534 PAD.n1972 0.019716
R47928 PAD.n9534 PAD.n9533 0.019716
R47929 PAD.n9540 PAD.n1971 0.019716
R47930 PAD.n9541 PAD.n9540 0.019716
R47931 PAD.n9546 PAD.n1970 0.019716
R47932 PAD.n9546 PAD.n9545 0.019716
R47933 PAD.n9552 PAD.n1969 0.019716
R47934 PAD.n9553 PAD.n9552 0.019716
R47935 PAD.n9558 PAD.n1968 0.019716
R47936 PAD.n9558 PAD.n9557 0.019716
R47937 PAD.n9564 PAD.n1967 0.019716
R47938 PAD.n9565 PAD.n9564 0.019716
R47939 PAD.n9570 PAD.n1966 0.019716
R47940 PAD.n9570 PAD.n9569 0.019716
R47941 PAD.n9576 PAD.n1965 0.019716
R47942 PAD.n9577 PAD.n9576 0.019716
R47943 PAD.n9582 PAD.n1964 0.019716
R47944 PAD.n9582 PAD.n9581 0.019716
R47945 PAD.n9588 PAD.n1963 0.019716
R47946 PAD.n9589 PAD.n9588 0.019716
R47947 PAD.n9594 PAD.n1962 0.019716
R47948 PAD.n9594 PAD.n9593 0.019716
R47949 PAD.n9600 PAD.n1961 0.019716
R47950 PAD.n9601 PAD.n9600 0.019716
R47951 PAD.n9606 PAD.n1960 0.019716
R47952 PAD.n9606 PAD.n9605 0.019716
R47953 PAD.n9612 PAD.n1959 0.019716
R47954 PAD.n9613 PAD.n9612 0.019716
R47955 PAD.n9618 PAD.n1958 0.019716
R47956 PAD.n9618 PAD.n9617 0.019716
R47957 PAD.n9624 PAD.n1957 0.019716
R47958 PAD.n9625 PAD.n9624 0.019716
R47959 PAD.n9630 PAD.n1956 0.019716
R47960 PAD.n9630 PAD.n9629 0.019716
R47961 PAD.n9636 PAD.n1955 0.019716
R47962 PAD.n9637 PAD.n9636 0.019716
R47963 PAD.n9642 PAD.n1954 0.019716
R47964 PAD.n9642 PAD.n9641 0.019716
R47965 PAD.n9648 PAD.n1953 0.019716
R47966 PAD.n9649 PAD.n9648 0.019716
R47967 PAD.n9654 PAD.n1952 0.019716
R47968 PAD.n9654 PAD.n9653 0.019716
R47969 PAD.n9660 PAD.n1951 0.019716
R47970 PAD.n9661 PAD.n9660 0.019716
R47971 PAD.n9666 PAD.n1950 0.019716
R47972 PAD.n9666 PAD.n9665 0.019716
R47973 PAD.n9672 PAD.n1949 0.019716
R47974 PAD.n9673 PAD.n9672 0.019716
R47975 PAD.n9678 PAD.n1948 0.019716
R47976 PAD.n9678 PAD.n9677 0.019716
R47977 PAD.n9684 PAD.n1947 0.019716
R47978 PAD.n9685 PAD.n9684 0.019716
R47979 PAD.n9690 PAD.n1946 0.019716
R47980 PAD.n9690 PAD.n9689 0.019716
R47981 PAD.n9696 PAD.n1945 0.019716
R47982 PAD.n9697 PAD.n9696 0.019716
R47983 PAD.n9702 PAD.n1944 0.019716
R47984 PAD.n9702 PAD.n9701 0.019716
R47985 PAD.n9709 PAD.n1943 0.019716
R47986 PAD.n9710 PAD.n9709 0.019716
R47987 PAD.n2133 PAD.n2132 0.019716
R47988 PAD.n9202 PAD.n2087 0.019716
R47989 PAD.n9203 PAD.n9202 0.019716
R47990 PAD.n9208 PAD.n2086 0.019716
R47991 PAD.n9208 PAD.n9207 0.019716
R47992 PAD.n9214 PAD.n2085 0.019716
R47993 PAD.n9215 PAD.n9214 0.019716
R47994 PAD.n9220 PAD.n2084 0.019716
R47995 PAD.n9220 PAD.n9219 0.019716
R47996 PAD.n9226 PAD.n2083 0.019716
R47997 PAD.n9227 PAD.n9226 0.019716
R47998 PAD.n9232 PAD.n2082 0.019716
R47999 PAD.n9232 PAD.n9231 0.019716
R48000 PAD.n9238 PAD.n2081 0.019716
R48001 PAD.n9239 PAD.n9238 0.019716
R48002 PAD.n9244 PAD.n2080 0.019716
R48003 PAD.n9244 PAD.n9243 0.019716
R48004 PAD.n9250 PAD.n2079 0.019716
R48005 PAD.n9251 PAD.n9250 0.019716
R48006 PAD.n9256 PAD.n2078 0.019716
R48007 PAD.n9256 PAD.n9255 0.019716
R48008 PAD.n9262 PAD.n2077 0.019716
R48009 PAD.n9263 PAD.n9262 0.019716
R48010 PAD.n9268 PAD.n2076 0.019716
R48011 PAD.n9268 PAD.n9267 0.019716
R48012 PAD.n9274 PAD.n2075 0.019716
R48013 PAD.n9275 PAD.n9274 0.019716
R48014 PAD.n9280 PAD.n2074 0.019716
R48015 PAD.n9280 PAD.n9279 0.019716
R48016 PAD.n9286 PAD.n2073 0.019716
R48017 PAD.n9287 PAD.n9286 0.019716
R48018 PAD.n9292 PAD.n2072 0.019716
R48019 PAD.n9292 PAD.n9291 0.019716
R48020 PAD.n9298 PAD.n2071 0.019716
R48021 PAD.n9299 PAD.n9298 0.019716
R48022 PAD.n9304 PAD.n2070 0.019716
R48023 PAD.n9304 PAD.n9303 0.019716
R48024 PAD.n9310 PAD.n2069 0.019716
R48025 PAD.n9311 PAD.n9310 0.019716
R48026 PAD.n9316 PAD.n2068 0.019716
R48027 PAD.n9316 PAD.n9315 0.019716
R48028 PAD.n9322 PAD.n2067 0.019716
R48029 PAD.n9323 PAD.n9322 0.019716
R48030 PAD.n9328 PAD.n2066 0.019716
R48031 PAD.n9328 PAD.n9327 0.019716
R48032 PAD.n9334 PAD.n2065 0.019716
R48033 PAD.n9335 PAD.n9334 0.019716
R48034 PAD.n9340 PAD.n2064 0.019716
R48035 PAD.n9340 PAD.n9339 0.019716
R48036 PAD.n9346 PAD.n2063 0.019716
R48037 PAD.n9347 PAD.n9346 0.019716
R48038 PAD.n9352 PAD.n2062 0.019716
R48039 PAD.n9352 PAD.n9351 0.019716
R48040 PAD.n9358 PAD.n2061 0.019716
R48041 PAD.n9359 PAD.n9358 0.019716
R48042 PAD.n9364 PAD.n2060 0.019716
R48043 PAD.n9364 PAD.n9363 0.019716
R48044 PAD.n9370 PAD.n2059 0.019716
R48045 PAD.n9371 PAD.n9370 0.019716
R48046 PAD.n9376 PAD.n2058 0.019716
R48047 PAD.n9376 PAD.n9375 0.019716
R48048 PAD.n9382 PAD.n2057 0.019716
R48049 PAD.n9383 PAD.n9382 0.019716
R48050 PAD.n9388 PAD.n2056 0.019716
R48051 PAD.n9388 PAD.n9387 0.019716
R48052 PAD.n9394 PAD.n2055 0.019716
R48053 PAD.n9395 PAD.n9394 0.019716
R48054 PAD.n9400 PAD.n2054 0.019716
R48055 PAD.n9400 PAD.n9399 0.019716
R48056 PAD.n9406 PAD.n2053 0.019716
R48057 PAD.n9407 PAD.n9406 0.019716
R48058 PAD.n9412 PAD.n2052 0.019716
R48059 PAD.n9412 PAD.n9411 0.019716
R48060 PAD.n9418 PAD.n2051 0.019716
R48061 PAD.n9419 PAD.n9418 0.019716
R48062 PAD.n9424 PAD.n2050 0.019716
R48063 PAD.n9424 PAD.n9423 0.019716
R48064 PAD.n9430 PAD.n2049 0.019716
R48065 PAD.n9431 PAD.n9430 0.019716
R48066 PAD.n9436 PAD.n2048 0.019716
R48067 PAD.n9436 PAD.n9435 0.019716
R48068 PAD.n9442 PAD.n2047 0.019716
R48069 PAD.n9443 PAD.n9442 0.019716
R48070 PAD.n2480 PAD.n2153 0.019716
R48071 PAD.n2479 PAD.n2478 0.019716
R48072 PAD.n2478 PAD.n2477 0.019716
R48073 PAD.n2468 PAD.n2154 0.019716
R48074 PAD.n2469 PAD.n2468 0.019716
R48075 PAD.n2467 PAD.n2466 0.019716
R48076 PAD.n2466 PAD.n2465 0.019716
R48077 PAD.n2456 PAD.n2159 0.019716
R48078 PAD.n2457 PAD.n2456 0.019716
R48079 PAD.n2455 PAD.n2454 0.019716
R48080 PAD.n2454 PAD.n2453 0.019716
R48081 PAD.n2444 PAD.n2163 0.019716
R48082 PAD.n2445 PAD.n2444 0.019716
R48083 PAD.n2443 PAD.n2442 0.019716
R48084 PAD.n2442 PAD.n2441 0.019716
R48085 PAD.n2432 PAD.n2167 0.019716
R48086 PAD.n2433 PAD.n2432 0.019716
R48087 PAD.n2431 PAD.n2430 0.019716
R48088 PAD.n2430 PAD.n2429 0.019716
R48089 PAD.n2420 PAD.n2171 0.019716
R48090 PAD.n2421 PAD.n2420 0.019716
R48091 PAD.n2419 PAD.n2418 0.019716
R48092 PAD.n2418 PAD.n2417 0.019716
R48093 PAD.n2408 PAD.n2175 0.019716
R48094 PAD.n2409 PAD.n2408 0.019716
R48095 PAD.n2407 PAD.n2406 0.019716
R48096 PAD.n2406 PAD.n2405 0.019716
R48097 PAD.n2396 PAD.n2179 0.019716
R48098 PAD.n2397 PAD.n2396 0.019716
R48099 PAD.n2395 PAD.n2394 0.019716
R48100 PAD.n2394 PAD.n2393 0.019716
R48101 PAD.n2384 PAD.n2183 0.019716
R48102 PAD.n2385 PAD.n2384 0.019716
R48103 PAD.n2383 PAD.n2382 0.019716
R48104 PAD.n2382 PAD.n2381 0.019716
R48105 PAD.n2372 PAD.n2187 0.019716
R48106 PAD.n2373 PAD.n2372 0.019716
R48107 PAD.n2371 PAD.n2370 0.019716
R48108 PAD.n2370 PAD.n2369 0.019716
R48109 PAD.n2360 PAD.n2191 0.019716
R48110 PAD.n2361 PAD.n2360 0.019716
R48111 PAD.n2359 PAD.n2358 0.019716
R48112 PAD.n2358 PAD.n2357 0.019716
R48113 PAD.n2348 PAD.n2195 0.019716
R48114 PAD.n2349 PAD.n2348 0.019716
R48115 PAD.n2347 PAD.n2346 0.019716
R48116 PAD.n2346 PAD.n2345 0.019716
R48117 PAD.n2336 PAD.n2199 0.019716
R48118 PAD.n2337 PAD.n2336 0.019716
R48119 PAD.n2335 PAD.n2334 0.019716
R48120 PAD.n2334 PAD.n2333 0.019716
R48121 PAD.n2324 PAD.n2203 0.019716
R48122 PAD.n2325 PAD.n2324 0.019716
R48123 PAD.n2323 PAD.n2322 0.019716
R48124 PAD.n2322 PAD.n2321 0.019716
R48125 PAD.n2312 PAD.n2207 0.019716
R48126 PAD.n2313 PAD.n2312 0.019716
R48127 PAD.n2311 PAD.n2310 0.019716
R48128 PAD.n2310 PAD.n2309 0.019716
R48129 PAD.n2300 PAD.n2211 0.019716
R48130 PAD.n2301 PAD.n2300 0.019716
R48131 PAD.n2299 PAD.n2298 0.019716
R48132 PAD.n2298 PAD.n2297 0.019716
R48133 PAD.n2288 PAD.n2215 0.019716
R48134 PAD.n2289 PAD.n2288 0.019716
R48135 PAD.n2287 PAD.n2286 0.019716
R48136 PAD.n2286 PAD.n2285 0.019716
R48137 PAD.n2276 PAD.n2219 0.019716
R48138 PAD.n2277 PAD.n2276 0.019716
R48139 PAD.n2275 PAD.n2274 0.019716
R48140 PAD.n2274 PAD.n2273 0.019716
R48141 PAD.n2264 PAD.n2223 0.019716
R48142 PAD.n2265 PAD.n2264 0.019716
R48143 PAD.n2263 PAD.n2262 0.019716
R48144 PAD.n2262 PAD.n2261 0.019716
R48145 PAD.n2252 PAD.n2227 0.019716
R48146 PAD.n2253 PAD.n2252 0.019716
R48147 PAD.n2251 PAD.n2250 0.019716
R48148 PAD.n2250 PAD.n2249 0.019716
R48149 PAD.n2240 PAD.n2231 0.019716
R48150 PAD.n2241 PAD.n2240 0.019716
R48151 PAD.n2239 PAD.n2238 0.019716
R48152 PAD.n2238 PAD.n2237 0.019716
R48153 PAD.n2827 PAD.n2500 0.019716
R48154 PAD.n2826 PAD.n2825 0.019716
R48155 PAD.n2825 PAD.n2824 0.019716
R48156 PAD.n2815 PAD.n2501 0.019716
R48157 PAD.n2816 PAD.n2815 0.019716
R48158 PAD.n2814 PAD.n2813 0.019716
R48159 PAD.n2813 PAD.n2812 0.019716
R48160 PAD.n2803 PAD.n2506 0.019716
R48161 PAD.n2804 PAD.n2803 0.019716
R48162 PAD.n2802 PAD.n2801 0.019716
R48163 PAD.n2801 PAD.n2800 0.019716
R48164 PAD.n2791 PAD.n2510 0.019716
R48165 PAD.n2792 PAD.n2791 0.019716
R48166 PAD.n2790 PAD.n2789 0.019716
R48167 PAD.n2789 PAD.n2788 0.019716
R48168 PAD.n2779 PAD.n2514 0.019716
R48169 PAD.n2780 PAD.n2779 0.019716
R48170 PAD.n2778 PAD.n2777 0.019716
R48171 PAD.n2777 PAD.n2776 0.019716
R48172 PAD.n2767 PAD.n2518 0.019716
R48173 PAD.n2768 PAD.n2767 0.019716
R48174 PAD.n2766 PAD.n2765 0.019716
R48175 PAD.n2765 PAD.n2764 0.019716
R48176 PAD.n2755 PAD.n2522 0.019716
R48177 PAD.n2756 PAD.n2755 0.019716
R48178 PAD.n2754 PAD.n2753 0.019716
R48179 PAD.n2753 PAD.n2752 0.019716
R48180 PAD.n2743 PAD.n2526 0.019716
R48181 PAD.n2744 PAD.n2743 0.019716
R48182 PAD.n2742 PAD.n2741 0.019716
R48183 PAD.n2741 PAD.n2740 0.019716
R48184 PAD.n2731 PAD.n2530 0.019716
R48185 PAD.n2732 PAD.n2731 0.019716
R48186 PAD.n2730 PAD.n2729 0.019716
R48187 PAD.n2729 PAD.n2728 0.019716
R48188 PAD.n2719 PAD.n2534 0.019716
R48189 PAD.n2720 PAD.n2719 0.019716
R48190 PAD.n2718 PAD.n2717 0.019716
R48191 PAD.n2717 PAD.n2716 0.019716
R48192 PAD.n2707 PAD.n2538 0.019716
R48193 PAD.n2708 PAD.n2707 0.019716
R48194 PAD.n2706 PAD.n2705 0.019716
R48195 PAD.n2705 PAD.n2704 0.019716
R48196 PAD.n2695 PAD.n2542 0.019716
R48197 PAD.n2696 PAD.n2695 0.019716
R48198 PAD.n2694 PAD.n2693 0.019716
R48199 PAD.n2693 PAD.n2692 0.019716
R48200 PAD.n2683 PAD.n2546 0.019716
R48201 PAD.n2684 PAD.n2683 0.019716
R48202 PAD.n2682 PAD.n2681 0.019716
R48203 PAD.n2681 PAD.n2680 0.019716
R48204 PAD.n2671 PAD.n2550 0.019716
R48205 PAD.n2672 PAD.n2671 0.019716
R48206 PAD.n2670 PAD.n2669 0.019716
R48207 PAD.n2669 PAD.n2668 0.019716
R48208 PAD.n2659 PAD.n2554 0.019716
R48209 PAD.n2660 PAD.n2659 0.019716
R48210 PAD.n2658 PAD.n2657 0.019716
R48211 PAD.n2657 PAD.n2656 0.019716
R48212 PAD.n2647 PAD.n2558 0.019716
R48213 PAD.n2648 PAD.n2647 0.019716
R48214 PAD.n2646 PAD.n2645 0.019716
R48215 PAD.n2645 PAD.n2644 0.019716
R48216 PAD.n2635 PAD.n2562 0.019716
R48217 PAD.n2636 PAD.n2635 0.019716
R48218 PAD.n2634 PAD.n2633 0.019716
R48219 PAD.n2633 PAD.n2632 0.019716
R48220 PAD.n2623 PAD.n2566 0.019716
R48221 PAD.n2624 PAD.n2623 0.019716
R48222 PAD.n2622 PAD.n2621 0.019716
R48223 PAD.n2621 PAD.n2620 0.019716
R48224 PAD.n2611 PAD.n2570 0.019716
R48225 PAD.n2612 PAD.n2611 0.019716
R48226 PAD.n2610 PAD.n2609 0.019716
R48227 PAD.n2609 PAD.n2608 0.019716
R48228 PAD.n2599 PAD.n2574 0.019716
R48229 PAD.n2600 PAD.n2599 0.019716
R48230 PAD.n2598 PAD.n2597 0.019716
R48231 PAD.n2597 PAD.n2596 0.019716
R48232 PAD.n2587 PAD.n2578 0.019716
R48233 PAD.n2588 PAD.n2587 0.019716
R48234 PAD.n2586 PAD.n2585 0.019716
R48235 PAD.n2585 PAD.n2584 0.019716
R48236 PAD.n9117 PAD.n9116 0.019716
R48237 PAD.n8841 PAD.n2875 0.019716
R48238 PAD.n8841 PAD.n8840 0.019716
R48239 PAD.n9110 PAD.n2874 0.019716
R48240 PAD.n9110 PAD.n9109 0.019716
R48241 PAD.n8846 PAD.n2873 0.019716
R48242 PAD.n8846 PAD.n8845 0.019716
R48243 PAD.n9101 PAD.n2872 0.019716
R48244 PAD.n9101 PAD.n9100 0.019716
R48245 PAD.n8851 PAD.n2871 0.019716
R48246 PAD.n8851 PAD.n8850 0.019716
R48247 PAD.n9092 PAD.n2870 0.019716
R48248 PAD.n9092 PAD.n9091 0.019716
R48249 PAD.n8856 PAD.n2869 0.019716
R48250 PAD.n8856 PAD.n8855 0.019716
R48251 PAD.n9083 PAD.n2868 0.019716
R48252 PAD.n9083 PAD.n9082 0.019716
R48253 PAD.n8861 PAD.n2867 0.019716
R48254 PAD.n8861 PAD.n8860 0.019716
R48255 PAD.n9074 PAD.n2866 0.019716
R48256 PAD.n9074 PAD.n9073 0.019716
R48257 PAD.n8866 PAD.n2865 0.019716
R48258 PAD.n8866 PAD.n8865 0.019716
R48259 PAD.n9065 PAD.n2864 0.019716
R48260 PAD.n9065 PAD.n9064 0.019716
R48261 PAD.n8871 PAD.n2863 0.019716
R48262 PAD.n8871 PAD.n8870 0.019716
R48263 PAD.n9056 PAD.n2862 0.019716
R48264 PAD.n9056 PAD.n9055 0.019716
R48265 PAD.n8876 PAD.n2861 0.019716
R48266 PAD.n8876 PAD.n8875 0.019716
R48267 PAD.n9047 PAD.n2860 0.019716
R48268 PAD.n9047 PAD.n9046 0.019716
R48269 PAD.n8881 PAD.n2859 0.019716
R48270 PAD.n8881 PAD.n8880 0.019716
R48271 PAD.n9038 PAD.n2858 0.019716
R48272 PAD.n9038 PAD.n9037 0.019716
R48273 PAD.n8886 PAD.n2857 0.019716
R48274 PAD.n8886 PAD.n8885 0.019716
R48275 PAD.n9029 PAD.n2856 0.019716
R48276 PAD.n9029 PAD.n9028 0.019716
R48277 PAD.n8891 PAD.n2855 0.019716
R48278 PAD.n8891 PAD.n8890 0.019716
R48279 PAD.n9020 PAD.n2854 0.019716
R48280 PAD.n9020 PAD.n9019 0.019716
R48281 PAD.n8896 PAD.n2853 0.019716
R48282 PAD.n8896 PAD.n8895 0.019716
R48283 PAD.n9011 PAD.n2852 0.019716
R48284 PAD.n9011 PAD.n9010 0.019716
R48285 PAD.n8901 PAD.n2851 0.019716
R48286 PAD.n8901 PAD.n8900 0.019716
R48287 PAD.n9002 PAD.n2850 0.019716
R48288 PAD.n9002 PAD.n9001 0.019716
R48289 PAD.n8906 PAD.n2849 0.019716
R48290 PAD.n8906 PAD.n8905 0.019716
R48291 PAD.n8993 PAD.n2848 0.019716
R48292 PAD.n8993 PAD.n8992 0.019716
R48293 PAD.n8911 PAD.n2847 0.019716
R48294 PAD.n8911 PAD.n8910 0.019716
R48295 PAD.n8984 PAD.n2846 0.019716
R48296 PAD.n8984 PAD.n8983 0.019716
R48297 PAD.n8916 PAD.n2845 0.019716
R48298 PAD.n8916 PAD.n8915 0.019716
R48299 PAD.n8975 PAD.n2844 0.019716
R48300 PAD.n8975 PAD.n8974 0.019716
R48301 PAD.n8921 PAD.n2843 0.019716
R48302 PAD.n8921 PAD.n8920 0.019716
R48303 PAD.n8966 PAD.n2842 0.019716
R48304 PAD.n8966 PAD.n8965 0.019716
R48305 PAD.n8926 PAD.n2841 0.019716
R48306 PAD.n8926 PAD.n8925 0.019716
R48307 PAD.n8957 PAD.n2840 0.019716
R48308 PAD.n8957 PAD.n8956 0.019716
R48309 PAD.n8931 PAD.n2839 0.019716
R48310 PAD.n8931 PAD.n8930 0.019716
R48311 PAD.n8948 PAD.n2838 0.019716
R48312 PAD.n8948 PAD.n8947 0.019716
R48313 PAD.n8936 PAD.n2837 0.019716
R48314 PAD.n8936 PAD.n8935 0.019716
R48315 PAD.n8939 PAD.n2836 0.019716
R48316 PAD.n8939 PAD.n8938 0.019716
R48317 PAD.n9137 PAD.n2835 0.019716
R48318 PAD.n9138 PAD.n9137 0.019716
R48319 PAD.n8820 PAD.n8528 0.019716
R48320 PAD.n8813 PAD.n8812 0.019716
R48321 PAD.n8813 PAD.n2945 0.019716
R48322 PAD.n8809 PAD.n8808 0.019716
R48323 PAD.n8808 PAD.n2944 0.019716
R48324 PAD.n8802 PAD.n8801 0.019716
R48325 PAD.n8802 PAD.n2943 0.019716
R48326 PAD.n8797 PAD.n8796 0.019716
R48327 PAD.n8796 PAD.n2942 0.019716
R48328 PAD.n8790 PAD.n8789 0.019716
R48329 PAD.n8790 PAD.n2941 0.019716
R48330 PAD.n8785 PAD.n8784 0.019716
R48331 PAD.n8784 PAD.n2940 0.019716
R48332 PAD.n8778 PAD.n8777 0.019716
R48333 PAD.n8778 PAD.n2939 0.019716
R48334 PAD.n8773 PAD.n8772 0.019716
R48335 PAD.n8772 PAD.n2938 0.019716
R48336 PAD.n8766 PAD.n8765 0.019716
R48337 PAD.n8766 PAD.n2937 0.019716
R48338 PAD.n8761 PAD.n8760 0.019716
R48339 PAD.n8760 PAD.n2936 0.019716
R48340 PAD.n8754 PAD.n8753 0.019716
R48341 PAD.n8754 PAD.n2935 0.019716
R48342 PAD.n8749 PAD.n8748 0.019716
R48343 PAD.n8748 PAD.n2934 0.019716
R48344 PAD.n8742 PAD.n8741 0.019716
R48345 PAD.n8742 PAD.n2933 0.019716
R48346 PAD.n8737 PAD.n8736 0.019716
R48347 PAD.n8736 PAD.n2932 0.019716
R48348 PAD.n8730 PAD.n8729 0.019716
R48349 PAD.n8730 PAD.n2931 0.019716
R48350 PAD.n8725 PAD.n8724 0.019716
R48351 PAD.n8724 PAD.n2930 0.019716
R48352 PAD.n8718 PAD.n8717 0.019716
R48353 PAD.n8718 PAD.n2929 0.019716
R48354 PAD.n8713 PAD.n8712 0.019716
R48355 PAD.n8712 PAD.n2928 0.019716
R48356 PAD.n8706 PAD.n8705 0.019716
R48357 PAD.n8706 PAD.n2927 0.019716
R48358 PAD.n8701 PAD.n8700 0.019716
R48359 PAD.n8700 PAD.n2926 0.019716
R48360 PAD.n8694 PAD.n8693 0.019716
R48361 PAD.n8694 PAD.n2925 0.019716
R48362 PAD.n8689 PAD.n8688 0.019716
R48363 PAD.n8688 PAD.n2924 0.019716
R48364 PAD.n8682 PAD.n8681 0.019716
R48365 PAD.n8682 PAD.n2923 0.019716
R48366 PAD.n8677 PAD.n8676 0.019716
R48367 PAD.n8676 PAD.n2922 0.019716
R48368 PAD.n8670 PAD.n8669 0.019716
R48369 PAD.n8670 PAD.n2921 0.019716
R48370 PAD.n8665 PAD.n8664 0.019716
R48371 PAD.n8664 PAD.n2920 0.019716
R48372 PAD.n8658 PAD.n8657 0.019716
R48373 PAD.n8658 PAD.n2919 0.019716
R48374 PAD.n8653 PAD.n8652 0.019716
R48375 PAD.n8652 PAD.n2918 0.019716
R48376 PAD.n8646 PAD.n8645 0.019716
R48377 PAD.n8646 PAD.n2917 0.019716
R48378 PAD.n8641 PAD.n8640 0.019716
R48379 PAD.n8640 PAD.n2916 0.019716
R48380 PAD.n8634 PAD.n8633 0.019716
R48381 PAD.n8634 PAD.n2915 0.019716
R48382 PAD.n8629 PAD.n8628 0.019716
R48383 PAD.n8628 PAD.n2914 0.019716
R48384 PAD.n8622 PAD.n8621 0.019716
R48385 PAD.n8622 PAD.n2913 0.019716
R48386 PAD.n8617 PAD.n8616 0.019716
R48387 PAD.n8616 PAD.n2912 0.019716
R48388 PAD.n8610 PAD.n8609 0.019716
R48389 PAD.n8610 PAD.n2911 0.019716
R48390 PAD.n8605 PAD.n8604 0.019716
R48391 PAD.n8604 PAD.n2910 0.019716
R48392 PAD.n8598 PAD.n8597 0.019716
R48393 PAD.n8598 PAD.n2909 0.019716
R48394 PAD.n8593 PAD.n8592 0.019716
R48395 PAD.n8592 PAD.n2908 0.019716
R48396 PAD.n8586 PAD.n8585 0.019716
R48397 PAD.n8586 PAD.n2907 0.019716
R48398 PAD.n8581 PAD.n8580 0.019716
R48399 PAD.n8580 PAD.n2906 0.019716
R48400 PAD.n8574 PAD.n8573 0.019716
R48401 PAD.n8574 PAD.n2905 0.019716
R48402 PAD.n3039 PAD.n3038 0.019716
R48403 PAD.n3046 PAD.n2993 0.019716
R48404 PAD.n3047 PAD.n3046 0.019716
R48405 PAD.n3052 PAD.n2992 0.019716
R48406 PAD.n3052 PAD.n3051 0.019716
R48407 PAD.n3058 PAD.n2991 0.019716
R48408 PAD.n3059 PAD.n3058 0.019716
R48409 PAD.n3064 PAD.n2990 0.019716
R48410 PAD.n3064 PAD.n3063 0.019716
R48411 PAD.n3070 PAD.n2989 0.019716
R48412 PAD.n3071 PAD.n3070 0.019716
R48413 PAD.n3076 PAD.n2988 0.019716
R48414 PAD.n3076 PAD.n3075 0.019716
R48415 PAD.n3082 PAD.n2987 0.019716
R48416 PAD.n3083 PAD.n3082 0.019716
R48417 PAD.n3088 PAD.n2986 0.019716
R48418 PAD.n3088 PAD.n3087 0.019716
R48419 PAD.n3094 PAD.n2985 0.019716
R48420 PAD.n3095 PAD.n3094 0.019716
R48421 PAD.n3100 PAD.n2984 0.019716
R48422 PAD.n3100 PAD.n3099 0.019716
R48423 PAD.n3106 PAD.n2983 0.019716
R48424 PAD.n3107 PAD.n3106 0.019716
R48425 PAD.n3112 PAD.n2982 0.019716
R48426 PAD.n3112 PAD.n3111 0.019716
R48427 PAD.n3118 PAD.n2981 0.019716
R48428 PAD.n3119 PAD.n3118 0.019716
R48429 PAD.n3124 PAD.n2980 0.019716
R48430 PAD.n3124 PAD.n3123 0.019716
R48431 PAD.n3130 PAD.n2979 0.019716
R48432 PAD.n3131 PAD.n3130 0.019716
R48433 PAD.n3136 PAD.n2978 0.019716
R48434 PAD.n3136 PAD.n3135 0.019716
R48435 PAD.n3142 PAD.n2977 0.019716
R48436 PAD.n3143 PAD.n3142 0.019716
R48437 PAD.n3148 PAD.n2976 0.019716
R48438 PAD.n3148 PAD.n3147 0.019716
R48439 PAD.n3154 PAD.n2975 0.019716
R48440 PAD.n3155 PAD.n3154 0.019716
R48441 PAD.n3160 PAD.n2974 0.019716
R48442 PAD.n3160 PAD.n3159 0.019716
R48443 PAD.n3166 PAD.n2973 0.019716
R48444 PAD.n3167 PAD.n3166 0.019716
R48445 PAD.n3172 PAD.n2972 0.019716
R48446 PAD.n3172 PAD.n3171 0.019716
R48447 PAD.n3178 PAD.n2971 0.019716
R48448 PAD.n3179 PAD.n3178 0.019716
R48449 PAD.n3184 PAD.n2970 0.019716
R48450 PAD.n3184 PAD.n3183 0.019716
R48451 PAD.n3190 PAD.n2969 0.019716
R48452 PAD.n3191 PAD.n3190 0.019716
R48453 PAD.n3196 PAD.n2968 0.019716
R48454 PAD.n3196 PAD.n3195 0.019716
R48455 PAD.n3202 PAD.n2967 0.019716
R48456 PAD.n3203 PAD.n3202 0.019716
R48457 PAD.n3208 PAD.n2966 0.019716
R48458 PAD.n3208 PAD.n3207 0.019716
R48459 PAD.n3214 PAD.n2965 0.019716
R48460 PAD.n3215 PAD.n3214 0.019716
R48461 PAD.n3220 PAD.n2964 0.019716
R48462 PAD.n3220 PAD.n3219 0.019716
R48463 PAD.n3226 PAD.n2963 0.019716
R48464 PAD.n3227 PAD.n3226 0.019716
R48465 PAD.n3232 PAD.n2962 0.019716
R48466 PAD.n3232 PAD.n3231 0.019716
R48467 PAD.n3238 PAD.n2961 0.019716
R48468 PAD.n3239 PAD.n3238 0.019716
R48469 PAD.n3244 PAD.n2960 0.019716
R48470 PAD.n3244 PAD.n3243 0.019716
R48471 PAD.n3250 PAD.n2959 0.019716
R48472 PAD.n3251 PAD.n3250 0.019716
R48473 PAD.n3256 PAD.n2958 0.019716
R48474 PAD.n3256 PAD.n3255 0.019716
R48475 PAD.n3262 PAD.n2957 0.019716
R48476 PAD.n3263 PAD.n3262 0.019716
R48477 PAD.n3268 PAD.n2956 0.019716
R48478 PAD.n3268 PAD.n3267 0.019716
R48479 PAD.n3274 PAD.n2955 0.019716
R48480 PAD.n3275 PAD.n3274 0.019716
R48481 PAD.n3280 PAD.n2954 0.019716
R48482 PAD.n3280 PAD.n3279 0.019716
R48483 PAD.n8514 PAD.n2953 0.019716
R48484 PAD.n8515 PAD.n8514 0.019716
R48485 PAD.n3384 PAD.n3383 0.019716
R48486 PAD.n3391 PAD.n3337 0.019716
R48487 PAD.n3392 PAD.n3391 0.019716
R48488 PAD.n3397 PAD.n3336 0.019716
R48489 PAD.n3397 PAD.n3396 0.019716
R48490 PAD.n3403 PAD.n3335 0.019716
R48491 PAD.n3404 PAD.n3403 0.019716
R48492 PAD.n3409 PAD.n3334 0.019716
R48493 PAD.n3409 PAD.n3408 0.019716
R48494 PAD.n3415 PAD.n3333 0.019716
R48495 PAD.n3416 PAD.n3415 0.019716
R48496 PAD.n3421 PAD.n3332 0.019716
R48497 PAD.n3421 PAD.n3420 0.019716
R48498 PAD.n3427 PAD.n3331 0.019716
R48499 PAD.n3428 PAD.n3427 0.019716
R48500 PAD.n3433 PAD.n3330 0.019716
R48501 PAD.n3433 PAD.n3432 0.019716
R48502 PAD.n3439 PAD.n3329 0.019716
R48503 PAD.n3440 PAD.n3439 0.019716
R48504 PAD.n3445 PAD.n3328 0.019716
R48505 PAD.n3445 PAD.n3444 0.019716
R48506 PAD.n3451 PAD.n3327 0.019716
R48507 PAD.n3452 PAD.n3451 0.019716
R48508 PAD.n3457 PAD.n3326 0.019716
R48509 PAD.n3457 PAD.n3456 0.019716
R48510 PAD.n3463 PAD.n3325 0.019716
R48511 PAD.n3464 PAD.n3463 0.019716
R48512 PAD.n3469 PAD.n3324 0.019716
R48513 PAD.n3469 PAD.n3468 0.019716
R48514 PAD.n3475 PAD.n3323 0.019716
R48515 PAD.n3476 PAD.n3475 0.019716
R48516 PAD.n3481 PAD.n3322 0.019716
R48517 PAD.n3481 PAD.n3480 0.019716
R48518 PAD.n3487 PAD.n3321 0.019716
R48519 PAD.n3488 PAD.n3487 0.019716
R48520 PAD.n3493 PAD.n3320 0.019716
R48521 PAD.n3493 PAD.n3492 0.019716
R48522 PAD.n3499 PAD.n3319 0.019716
R48523 PAD.n3500 PAD.n3499 0.019716
R48524 PAD.n3505 PAD.n3318 0.019716
R48525 PAD.n3505 PAD.n3504 0.019716
R48526 PAD.n3511 PAD.n3317 0.019716
R48527 PAD.n3512 PAD.n3511 0.019716
R48528 PAD.n3517 PAD.n3316 0.019716
R48529 PAD.n3517 PAD.n3516 0.019716
R48530 PAD.n3523 PAD.n3315 0.019716
R48531 PAD.n3524 PAD.n3523 0.019716
R48532 PAD.n3529 PAD.n3314 0.019716
R48533 PAD.n3529 PAD.n3528 0.019716
R48534 PAD.n3535 PAD.n3313 0.019716
R48535 PAD.n3536 PAD.n3535 0.019716
R48536 PAD.n3541 PAD.n3312 0.019716
R48537 PAD.n3541 PAD.n3540 0.019716
R48538 PAD.n3547 PAD.n3311 0.019716
R48539 PAD.n3548 PAD.n3547 0.019716
R48540 PAD.n3553 PAD.n3310 0.019716
R48541 PAD.n3553 PAD.n3552 0.019716
R48542 PAD.n3559 PAD.n3309 0.019716
R48543 PAD.n3560 PAD.n3559 0.019716
R48544 PAD.n3565 PAD.n3308 0.019716
R48545 PAD.n3565 PAD.n3564 0.019716
R48546 PAD.n3571 PAD.n3307 0.019716
R48547 PAD.n3572 PAD.n3571 0.019716
R48548 PAD.n3577 PAD.n3306 0.019716
R48549 PAD.n3577 PAD.n3576 0.019716
R48550 PAD.n3583 PAD.n3305 0.019716
R48551 PAD.n3584 PAD.n3583 0.019716
R48552 PAD.n3589 PAD.n3304 0.019716
R48553 PAD.n3589 PAD.n3588 0.019716
R48554 PAD.n3595 PAD.n3303 0.019716
R48555 PAD.n3596 PAD.n3595 0.019716
R48556 PAD.n3601 PAD.n3302 0.019716
R48557 PAD.n3601 PAD.n3600 0.019716
R48558 PAD.n3607 PAD.n3301 0.019716
R48559 PAD.n3608 PAD.n3607 0.019716
R48560 PAD.n3613 PAD.n3300 0.019716
R48561 PAD.n3613 PAD.n3612 0.019716
R48562 PAD.n3619 PAD.n3299 0.019716
R48563 PAD.n3620 PAD.n3619 0.019716
R48564 PAD.n3625 PAD.n3298 0.019716
R48565 PAD.n3625 PAD.n3624 0.019716
R48566 PAD.n8489 PAD.n3297 0.019716
R48567 PAD.n8490 PAD.n8489 0.019716
R48568 PAD.n3729 PAD.n3728 0.019716
R48569 PAD.n3736 PAD.n3682 0.019716
R48570 PAD.n3737 PAD.n3736 0.019716
R48571 PAD.n3742 PAD.n3681 0.019716
R48572 PAD.n3742 PAD.n3741 0.019716
R48573 PAD.n3748 PAD.n3680 0.019716
R48574 PAD.n3749 PAD.n3748 0.019716
R48575 PAD.n3754 PAD.n3679 0.019716
R48576 PAD.n3754 PAD.n3753 0.019716
R48577 PAD.n3760 PAD.n3678 0.019716
R48578 PAD.n3761 PAD.n3760 0.019716
R48579 PAD.n3766 PAD.n3677 0.019716
R48580 PAD.n3766 PAD.n3765 0.019716
R48581 PAD.n3772 PAD.n3676 0.019716
R48582 PAD.n3773 PAD.n3772 0.019716
R48583 PAD.n3778 PAD.n3675 0.019716
R48584 PAD.n3778 PAD.n3777 0.019716
R48585 PAD.n3784 PAD.n3674 0.019716
R48586 PAD.n3785 PAD.n3784 0.019716
R48587 PAD.n3790 PAD.n3673 0.019716
R48588 PAD.n3790 PAD.n3789 0.019716
R48589 PAD.n3796 PAD.n3672 0.019716
R48590 PAD.n3797 PAD.n3796 0.019716
R48591 PAD.n3802 PAD.n3671 0.019716
R48592 PAD.n3802 PAD.n3801 0.019716
R48593 PAD.n3808 PAD.n3670 0.019716
R48594 PAD.n3809 PAD.n3808 0.019716
R48595 PAD.n3814 PAD.n3669 0.019716
R48596 PAD.n3814 PAD.n3813 0.019716
R48597 PAD.n3820 PAD.n3668 0.019716
R48598 PAD.n3821 PAD.n3820 0.019716
R48599 PAD.n3826 PAD.n3667 0.019716
R48600 PAD.n3826 PAD.n3825 0.019716
R48601 PAD.n3832 PAD.n3666 0.019716
R48602 PAD.n3833 PAD.n3832 0.019716
R48603 PAD.n3838 PAD.n3665 0.019716
R48604 PAD.n3838 PAD.n3837 0.019716
R48605 PAD.n3844 PAD.n3664 0.019716
R48606 PAD.n3845 PAD.n3844 0.019716
R48607 PAD.n3850 PAD.n3663 0.019716
R48608 PAD.n3850 PAD.n3849 0.019716
R48609 PAD.n3856 PAD.n3662 0.019716
R48610 PAD.n3857 PAD.n3856 0.019716
R48611 PAD.n3862 PAD.n3661 0.019716
R48612 PAD.n3862 PAD.n3861 0.019716
R48613 PAD.n3868 PAD.n3660 0.019716
R48614 PAD.n3869 PAD.n3868 0.019716
R48615 PAD.n3874 PAD.n3659 0.019716
R48616 PAD.n3874 PAD.n3873 0.019716
R48617 PAD.n3880 PAD.n3658 0.019716
R48618 PAD.n3881 PAD.n3880 0.019716
R48619 PAD.n3886 PAD.n3657 0.019716
R48620 PAD.n3886 PAD.n3885 0.019716
R48621 PAD.n3892 PAD.n3656 0.019716
R48622 PAD.n3893 PAD.n3892 0.019716
R48623 PAD.n3898 PAD.n3655 0.019716
R48624 PAD.n3898 PAD.n3897 0.019716
R48625 PAD.n3904 PAD.n3654 0.019716
R48626 PAD.n3905 PAD.n3904 0.019716
R48627 PAD.n3910 PAD.n3653 0.019716
R48628 PAD.n3910 PAD.n3909 0.019716
R48629 PAD.n3916 PAD.n3652 0.019716
R48630 PAD.n3917 PAD.n3916 0.019716
R48631 PAD.n3922 PAD.n3651 0.019716
R48632 PAD.n3922 PAD.n3921 0.019716
R48633 PAD.n3928 PAD.n3650 0.019716
R48634 PAD.n3929 PAD.n3928 0.019716
R48635 PAD.n3934 PAD.n3649 0.019716
R48636 PAD.n3934 PAD.n3933 0.019716
R48637 PAD.n3940 PAD.n3648 0.019716
R48638 PAD.n3941 PAD.n3940 0.019716
R48639 PAD.n3946 PAD.n3647 0.019716
R48640 PAD.n3946 PAD.n3945 0.019716
R48641 PAD.n3952 PAD.n3646 0.019716
R48642 PAD.n3953 PAD.n3952 0.019716
R48643 PAD.n3958 PAD.n3645 0.019716
R48644 PAD.n3958 PAD.n3957 0.019716
R48645 PAD.n3964 PAD.n3644 0.019716
R48646 PAD.n3965 PAD.n3964 0.019716
R48647 PAD.n3970 PAD.n3643 0.019716
R48648 PAD.n3970 PAD.n3969 0.019716
R48649 PAD.n8465 PAD.n3642 0.019716
R48650 PAD.n8466 PAD.n8465 0.019716
R48651 PAD.n4070 PAD.n4069 0.019716
R48652 PAD.n4077 PAD.n4024 0.019716
R48653 PAD.n4078 PAD.n4077 0.019716
R48654 PAD.n4083 PAD.n4023 0.019716
R48655 PAD.n4083 PAD.n4082 0.019716
R48656 PAD.n4089 PAD.n4022 0.019716
R48657 PAD.n4090 PAD.n4089 0.019716
R48658 PAD.n4095 PAD.n4021 0.019716
R48659 PAD.n4095 PAD.n4094 0.019716
R48660 PAD.n4101 PAD.n4020 0.019716
R48661 PAD.n4102 PAD.n4101 0.019716
R48662 PAD.n4107 PAD.n4019 0.019716
R48663 PAD.n4107 PAD.n4106 0.019716
R48664 PAD.n4113 PAD.n4018 0.019716
R48665 PAD.n4114 PAD.n4113 0.019716
R48666 PAD.n4119 PAD.n4017 0.019716
R48667 PAD.n4119 PAD.n4118 0.019716
R48668 PAD.n4125 PAD.n4016 0.019716
R48669 PAD.n4126 PAD.n4125 0.019716
R48670 PAD.n4131 PAD.n4015 0.019716
R48671 PAD.n4131 PAD.n4130 0.019716
R48672 PAD.n4137 PAD.n4014 0.019716
R48673 PAD.n4138 PAD.n4137 0.019716
R48674 PAD.n4143 PAD.n4013 0.019716
R48675 PAD.n4143 PAD.n4142 0.019716
R48676 PAD.n4149 PAD.n4012 0.019716
R48677 PAD.n4150 PAD.n4149 0.019716
R48678 PAD.n4155 PAD.n4011 0.019716
R48679 PAD.n4155 PAD.n4154 0.019716
R48680 PAD.n4161 PAD.n4010 0.019716
R48681 PAD.n4162 PAD.n4161 0.019716
R48682 PAD.n4167 PAD.n4009 0.019716
R48683 PAD.n4167 PAD.n4166 0.019716
R48684 PAD.n4173 PAD.n4008 0.019716
R48685 PAD.n4174 PAD.n4173 0.019716
R48686 PAD.n4179 PAD.n4007 0.019716
R48687 PAD.n4179 PAD.n4178 0.019716
R48688 PAD.n4185 PAD.n4006 0.019716
R48689 PAD.n4186 PAD.n4185 0.019716
R48690 PAD.n4191 PAD.n4005 0.019716
R48691 PAD.n4191 PAD.n4190 0.019716
R48692 PAD.n4197 PAD.n4004 0.019716
R48693 PAD.n4198 PAD.n4197 0.019716
R48694 PAD.n4203 PAD.n4003 0.019716
R48695 PAD.n4203 PAD.n4202 0.019716
R48696 PAD.n4209 PAD.n4002 0.019716
R48697 PAD.n4210 PAD.n4209 0.019716
R48698 PAD.n4215 PAD.n4001 0.019716
R48699 PAD.n4215 PAD.n4214 0.019716
R48700 PAD.n4221 PAD.n4000 0.019716
R48701 PAD.n4222 PAD.n4221 0.019716
R48702 PAD.n4227 PAD.n3999 0.019716
R48703 PAD.n4227 PAD.n4226 0.019716
R48704 PAD.n4233 PAD.n3998 0.019716
R48705 PAD.n4234 PAD.n4233 0.019716
R48706 PAD.n4239 PAD.n3997 0.019716
R48707 PAD.n4239 PAD.n4238 0.019716
R48708 PAD.n4245 PAD.n3996 0.019716
R48709 PAD.n4246 PAD.n4245 0.019716
R48710 PAD.n4251 PAD.n3995 0.019716
R48711 PAD.n4251 PAD.n4250 0.019716
R48712 PAD.n4257 PAD.n3994 0.019716
R48713 PAD.n4258 PAD.n4257 0.019716
R48714 PAD.n4263 PAD.n3993 0.019716
R48715 PAD.n4263 PAD.n4262 0.019716
R48716 PAD.n4269 PAD.n3992 0.019716
R48717 PAD.n4270 PAD.n4269 0.019716
R48718 PAD.n4275 PAD.n3991 0.019716
R48719 PAD.n4275 PAD.n4274 0.019716
R48720 PAD.n4281 PAD.n3990 0.019716
R48721 PAD.n4282 PAD.n4281 0.019716
R48722 PAD.n4287 PAD.n3989 0.019716
R48723 PAD.n4287 PAD.n4286 0.019716
R48724 PAD.n4293 PAD.n3988 0.019716
R48725 PAD.n4294 PAD.n4293 0.019716
R48726 PAD.n4299 PAD.n3987 0.019716
R48727 PAD.n4299 PAD.n4298 0.019716
R48728 PAD.n4305 PAD.n3986 0.019716
R48729 PAD.n4306 PAD.n4305 0.019716
R48730 PAD.n4311 PAD.n3985 0.019716
R48731 PAD.n4311 PAD.n4310 0.019716
R48732 PAD.n8441 PAD.n3984 0.019716
R48733 PAD.n8442 PAD.n8441 0.019716
R48734 PAD.n4422 PAD.n4421 0.019716
R48735 PAD.n4426 PAD.n4423 0.019716
R48736 PAD.n4426 PAD.n4425 0.019716
R48737 PAD.n4432 PAD.n4415 0.019716
R48738 PAD.n4433 PAD.n4432 0.019716
R48739 PAD.n4438 PAD.n4435 0.019716
R48740 PAD.n4438 PAD.n4437 0.019716
R48741 PAD.n4444 PAD.n4411 0.019716
R48742 PAD.n4445 PAD.n4444 0.019716
R48743 PAD.n4450 PAD.n4447 0.019716
R48744 PAD.n4450 PAD.n4449 0.019716
R48745 PAD.n4456 PAD.n4407 0.019716
R48746 PAD.n4457 PAD.n4456 0.019716
R48747 PAD.n4462 PAD.n4459 0.019716
R48748 PAD.n4462 PAD.n4461 0.019716
R48749 PAD.n4468 PAD.n4403 0.019716
R48750 PAD.n4469 PAD.n4468 0.019716
R48751 PAD.n4474 PAD.n4471 0.019716
R48752 PAD.n4474 PAD.n4473 0.019716
R48753 PAD.n4480 PAD.n4399 0.019716
R48754 PAD.n4481 PAD.n4480 0.019716
R48755 PAD.n4486 PAD.n4483 0.019716
R48756 PAD.n4486 PAD.n4485 0.019716
R48757 PAD.n4492 PAD.n4395 0.019716
R48758 PAD.n4493 PAD.n4492 0.019716
R48759 PAD.n4498 PAD.n4495 0.019716
R48760 PAD.n4498 PAD.n4497 0.019716
R48761 PAD.n4504 PAD.n4391 0.019716
R48762 PAD.n4505 PAD.n4504 0.019716
R48763 PAD.n4510 PAD.n4507 0.019716
R48764 PAD.n4510 PAD.n4509 0.019716
R48765 PAD.n4516 PAD.n4387 0.019716
R48766 PAD.n4517 PAD.n4516 0.019716
R48767 PAD.n4522 PAD.n4519 0.019716
R48768 PAD.n4522 PAD.n4521 0.019716
R48769 PAD.n4528 PAD.n4383 0.019716
R48770 PAD.n4529 PAD.n4528 0.019716
R48771 PAD.n4534 PAD.n4531 0.019716
R48772 PAD.n4534 PAD.n4533 0.019716
R48773 PAD.n4540 PAD.n4379 0.019716
R48774 PAD.n4541 PAD.n4540 0.019716
R48775 PAD.n4546 PAD.n4543 0.019716
R48776 PAD.n4546 PAD.n4545 0.019716
R48777 PAD.n4552 PAD.n4375 0.019716
R48778 PAD.n4553 PAD.n4552 0.019716
R48779 PAD.n4558 PAD.n4555 0.019716
R48780 PAD.n4558 PAD.n4557 0.019716
R48781 PAD.n4564 PAD.n4371 0.019716
R48782 PAD.n4565 PAD.n4564 0.019716
R48783 PAD.n4570 PAD.n4567 0.019716
R48784 PAD.n4570 PAD.n4569 0.019716
R48785 PAD.n4576 PAD.n4367 0.019716
R48786 PAD.n4577 PAD.n4576 0.019716
R48787 PAD.n4582 PAD.n4579 0.019716
R48788 PAD.n4582 PAD.n4581 0.019716
R48789 PAD.n4588 PAD.n4363 0.019716
R48790 PAD.n4589 PAD.n4588 0.019716
R48791 PAD.n4594 PAD.n4591 0.019716
R48792 PAD.n4594 PAD.n4593 0.019716
R48793 PAD.n4600 PAD.n4359 0.019716
R48794 PAD.n4601 PAD.n4600 0.019716
R48795 PAD.n4606 PAD.n4603 0.019716
R48796 PAD.n4606 PAD.n4605 0.019716
R48797 PAD.n4612 PAD.n4355 0.019716
R48798 PAD.n4613 PAD.n4612 0.019716
R48799 PAD.n4618 PAD.n4615 0.019716
R48800 PAD.n4618 PAD.n4617 0.019716
R48801 PAD.n4624 PAD.n4351 0.019716
R48802 PAD.n4625 PAD.n4624 0.019716
R48803 PAD.n4630 PAD.n4627 0.019716
R48804 PAD.n4630 PAD.n4629 0.019716
R48805 PAD.n4636 PAD.n4347 0.019716
R48806 PAD.n4637 PAD.n4636 0.019716
R48807 PAD.n4642 PAD.n4639 0.019716
R48808 PAD.n4642 PAD.n4641 0.019716
R48809 PAD.n4648 PAD.n4343 0.019716
R48810 PAD.n4649 PAD.n4648 0.019716
R48811 PAD.n4654 PAD.n4651 0.019716
R48812 PAD.n4654 PAD.n4653 0.019716
R48813 PAD.n4661 PAD.n4339 0.019716
R48814 PAD.n4662 PAD.n4661 0.019716
R48815 PAD.n4665 PAD.n4664 0.019716
R48816 PAD.n4666 PAD.n4665 0.019716
R48817 PAD.n8396 PAD.n4725 0.019716
R48818 PAD.n4727 PAD.n4726 0.019716
R48819 PAD.n4727 PAD.n4723 0.019716
R48820 PAD.n8387 PAD.n8386 0.019716
R48821 PAD.n8386 PAD.n4722 0.019716
R48822 PAD.n4732 PAD.n4731 0.019716
R48823 PAD.n4731 PAD.n4721 0.019716
R48824 PAD.n8378 PAD.n8377 0.019716
R48825 PAD.n8377 PAD.n4720 0.019716
R48826 PAD.n4737 PAD.n4736 0.019716
R48827 PAD.n4736 PAD.n4719 0.019716
R48828 PAD.n8369 PAD.n8368 0.019716
R48829 PAD.n8368 PAD.n4718 0.019716
R48830 PAD.n4742 PAD.n4741 0.019716
R48831 PAD.n4741 PAD.n4717 0.019716
R48832 PAD.n8360 PAD.n8359 0.019716
R48833 PAD.n8359 PAD.n4716 0.019716
R48834 PAD.n4747 PAD.n4746 0.019716
R48835 PAD.n4746 PAD.n4715 0.019716
R48836 PAD.n8351 PAD.n8350 0.019716
R48837 PAD.n8350 PAD.n4714 0.019716
R48838 PAD.n4752 PAD.n4751 0.019716
R48839 PAD.n4751 PAD.n4713 0.019716
R48840 PAD.n8342 PAD.n8341 0.019716
R48841 PAD.n8341 PAD.n4712 0.019716
R48842 PAD.n4757 PAD.n4756 0.019716
R48843 PAD.n4756 PAD.n4711 0.019716
R48844 PAD.n8333 PAD.n8332 0.019716
R48845 PAD.n8332 PAD.n4710 0.019716
R48846 PAD.n4762 PAD.n4761 0.019716
R48847 PAD.n4761 PAD.n4709 0.019716
R48848 PAD.n8324 PAD.n8323 0.019716
R48849 PAD.n8323 PAD.n4708 0.019716
R48850 PAD.n4767 PAD.n4766 0.019716
R48851 PAD.n4766 PAD.n4707 0.019716
R48852 PAD.n8315 PAD.n8314 0.019716
R48853 PAD.n8314 PAD.n4706 0.019716
R48854 PAD.n4772 PAD.n4771 0.019716
R48855 PAD.n4771 PAD.n4705 0.019716
R48856 PAD.n8306 PAD.n8305 0.019716
R48857 PAD.n8305 PAD.n4704 0.019716
R48858 PAD.n4777 PAD.n4776 0.019716
R48859 PAD.n4776 PAD.n4703 0.019716
R48860 PAD.n8297 PAD.n8296 0.019716
R48861 PAD.n8296 PAD.n4702 0.019716
R48862 PAD.n4782 PAD.n4781 0.019716
R48863 PAD.n4781 PAD.n4701 0.019716
R48864 PAD.n8288 PAD.n8287 0.019716
R48865 PAD.n8287 PAD.n4700 0.019716
R48866 PAD.n4787 PAD.n4786 0.019716
R48867 PAD.n4786 PAD.n4699 0.019716
R48868 PAD.n8279 PAD.n8278 0.019716
R48869 PAD.n8278 PAD.n4698 0.019716
R48870 PAD.n4792 PAD.n4791 0.019716
R48871 PAD.n4791 PAD.n4697 0.019716
R48872 PAD.n8270 PAD.n8269 0.019716
R48873 PAD.n8269 PAD.n4696 0.019716
R48874 PAD.n4797 PAD.n4796 0.019716
R48875 PAD.n4796 PAD.n4695 0.019716
R48876 PAD.n8261 PAD.n8260 0.019716
R48877 PAD.n8260 PAD.n4694 0.019716
R48878 PAD.n4802 PAD.n4801 0.019716
R48879 PAD.n4801 PAD.n4693 0.019716
R48880 PAD.n8252 PAD.n8251 0.019716
R48881 PAD.n8251 PAD.n4692 0.019716
R48882 PAD.n4807 PAD.n4806 0.019716
R48883 PAD.n4806 PAD.n4691 0.019716
R48884 PAD.n8243 PAD.n8242 0.019716
R48885 PAD.n8242 PAD.n4690 0.019716
R48886 PAD.n4812 PAD.n4811 0.019716
R48887 PAD.n4811 PAD.n4689 0.019716
R48888 PAD.n8234 PAD.n8233 0.019716
R48889 PAD.n8233 PAD.n4688 0.019716
R48890 PAD.n4817 PAD.n4816 0.019716
R48891 PAD.n4816 PAD.n4687 0.019716
R48892 PAD.n8225 PAD.n8224 0.019716
R48893 PAD.n8224 PAD.n4686 0.019716
R48894 PAD.n4822 PAD.n4821 0.019716
R48895 PAD.n4821 PAD.n4685 0.019716
R48896 PAD.n8216 PAD.n8215 0.019716
R48897 PAD.n8215 PAD.n4684 0.019716
R48898 PAD.n4827 PAD.n4826 0.019716
R48899 PAD.n4826 PAD.n4683 0.019716
R48900 PAD.n5176 PAD.n4849 0.019716
R48901 PAD.n5175 PAD.n5174 0.019716
R48902 PAD.n5174 PAD.n5173 0.019716
R48903 PAD.n5164 PAD.n4850 0.019716
R48904 PAD.n5165 PAD.n5164 0.019716
R48905 PAD.n5163 PAD.n5162 0.019716
R48906 PAD.n5162 PAD.n5161 0.019716
R48907 PAD.n5152 PAD.n4855 0.019716
R48908 PAD.n5153 PAD.n5152 0.019716
R48909 PAD.n5151 PAD.n5150 0.019716
R48910 PAD.n5150 PAD.n5149 0.019716
R48911 PAD.n5140 PAD.n4859 0.019716
R48912 PAD.n5141 PAD.n5140 0.019716
R48913 PAD.n5139 PAD.n5138 0.019716
R48914 PAD.n5138 PAD.n5137 0.019716
R48915 PAD.n5128 PAD.n4863 0.019716
R48916 PAD.n5129 PAD.n5128 0.019716
R48917 PAD.n5127 PAD.n5126 0.019716
R48918 PAD.n5126 PAD.n5125 0.019716
R48919 PAD.n5116 PAD.n4867 0.019716
R48920 PAD.n5117 PAD.n5116 0.019716
R48921 PAD.n5115 PAD.n5114 0.019716
R48922 PAD.n5114 PAD.n5113 0.019716
R48923 PAD.n5104 PAD.n4871 0.019716
R48924 PAD.n5105 PAD.n5104 0.019716
R48925 PAD.n5103 PAD.n5102 0.019716
R48926 PAD.n5102 PAD.n5101 0.019716
R48927 PAD.n5092 PAD.n4875 0.019716
R48928 PAD.n5093 PAD.n5092 0.019716
R48929 PAD.n5091 PAD.n5090 0.019716
R48930 PAD.n5090 PAD.n5089 0.019716
R48931 PAD.n5080 PAD.n4879 0.019716
R48932 PAD.n5081 PAD.n5080 0.019716
R48933 PAD.n5079 PAD.n5078 0.019716
R48934 PAD.n5078 PAD.n5077 0.019716
R48935 PAD.n5068 PAD.n4883 0.019716
R48936 PAD.n5069 PAD.n5068 0.019716
R48937 PAD.n5067 PAD.n5066 0.019716
R48938 PAD.n5066 PAD.n5065 0.019716
R48939 PAD.n5056 PAD.n4887 0.019716
R48940 PAD.n5057 PAD.n5056 0.019716
R48941 PAD.n5055 PAD.n5054 0.019716
R48942 PAD.n5054 PAD.n5053 0.019716
R48943 PAD.n5044 PAD.n4891 0.019716
R48944 PAD.n5045 PAD.n5044 0.019716
R48945 PAD.n5043 PAD.n5042 0.019716
R48946 PAD.n5042 PAD.n5041 0.019716
R48947 PAD.n5032 PAD.n4895 0.019716
R48948 PAD.n5033 PAD.n5032 0.019716
R48949 PAD.n5031 PAD.n5030 0.019716
R48950 PAD.n5030 PAD.n5029 0.019716
R48951 PAD.n5020 PAD.n4899 0.019716
R48952 PAD.n5021 PAD.n5020 0.019716
R48953 PAD.n5019 PAD.n5018 0.019716
R48954 PAD.n5018 PAD.n5017 0.019716
R48955 PAD.n5008 PAD.n4903 0.019716
R48956 PAD.n5009 PAD.n5008 0.019716
R48957 PAD.n5007 PAD.n5006 0.019716
R48958 PAD.n5006 PAD.n5005 0.019716
R48959 PAD.n4996 PAD.n4907 0.019716
R48960 PAD.n4997 PAD.n4996 0.019716
R48961 PAD.n4995 PAD.n4994 0.019716
R48962 PAD.n4994 PAD.n4993 0.019716
R48963 PAD.n4984 PAD.n4911 0.019716
R48964 PAD.n4985 PAD.n4984 0.019716
R48965 PAD.n4983 PAD.n4982 0.019716
R48966 PAD.n4982 PAD.n4981 0.019716
R48967 PAD.n4972 PAD.n4915 0.019716
R48968 PAD.n4973 PAD.n4972 0.019716
R48969 PAD.n4971 PAD.n4970 0.019716
R48970 PAD.n4970 PAD.n4969 0.019716
R48971 PAD.n4960 PAD.n4919 0.019716
R48972 PAD.n4961 PAD.n4960 0.019716
R48973 PAD.n4959 PAD.n4958 0.019716
R48974 PAD.n4958 PAD.n4957 0.019716
R48975 PAD.n4948 PAD.n4923 0.019716
R48976 PAD.n4949 PAD.n4948 0.019716
R48977 PAD.n4947 PAD.n4946 0.019716
R48978 PAD.n4946 PAD.n4945 0.019716
R48979 PAD.n4936 PAD.n4927 0.019716
R48980 PAD.n4937 PAD.n4936 0.019716
R48981 PAD.n4935 PAD.n4934 0.019716
R48982 PAD.n4934 PAD.n4933 0.019716
R48983 PAD.n8162 PAD.n7871 0.019716
R48984 PAD.n7873 PAD.n7872 0.019716
R48985 PAD.n7873 PAD.n7870 0.019716
R48986 PAD.n8153 PAD.n8152 0.019716
R48987 PAD.n8152 PAD.n7869 0.019716
R48988 PAD.n7878 PAD.n7877 0.019716
R48989 PAD.n7877 PAD.n7868 0.019716
R48990 PAD.n8144 PAD.n8143 0.019716
R48991 PAD.n8143 PAD.n7867 0.019716
R48992 PAD.n7883 PAD.n7882 0.019716
R48993 PAD.n7882 PAD.n7866 0.019716
R48994 PAD.n8135 PAD.n8134 0.019716
R48995 PAD.n8134 PAD.n7865 0.019716
R48996 PAD.n7888 PAD.n7887 0.019716
R48997 PAD.n7887 PAD.n7864 0.019716
R48998 PAD.n8126 PAD.n8125 0.019716
R48999 PAD.n8125 PAD.n7863 0.019716
R49000 PAD.n7893 PAD.n7892 0.019716
R49001 PAD.n7892 PAD.n7862 0.019716
R49002 PAD.n8117 PAD.n8116 0.019716
R49003 PAD.n8116 PAD.n7861 0.019716
R49004 PAD.n7898 PAD.n7897 0.019716
R49005 PAD.n7897 PAD.n7860 0.019716
R49006 PAD.n8108 PAD.n8107 0.019716
R49007 PAD.n8107 PAD.n7859 0.019716
R49008 PAD.n7903 PAD.n7902 0.019716
R49009 PAD.n7902 PAD.n7858 0.019716
R49010 PAD.n8099 PAD.n8098 0.019716
R49011 PAD.n8098 PAD.n7857 0.019716
R49012 PAD.n7908 PAD.n7907 0.019716
R49013 PAD.n7907 PAD.n7856 0.019716
R49014 PAD.n8090 PAD.n8089 0.019716
R49015 PAD.n8089 PAD.n7855 0.019716
R49016 PAD.n7913 PAD.n7912 0.019716
R49017 PAD.n7912 PAD.n7854 0.019716
R49018 PAD.n8081 PAD.n8080 0.019716
R49019 PAD.n8080 PAD.n7853 0.019716
R49020 PAD.n7918 PAD.n7917 0.019716
R49021 PAD.n7917 PAD.n7852 0.019716
R49022 PAD.n8072 PAD.n8071 0.019716
R49023 PAD.n8071 PAD.n7851 0.019716
R49024 PAD.n7923 PAD.n7922 0.019716
R49025 PAD.n7922 PAD.n7850 0.019716
R49026 PAD.n8063 PAD.n8062 0.019716
R49027 PAD.n8062 PAD.n7849 0.019716
R49028 PAD.n7928 PAD.n7927 0.019716
R49029 PAD.n7927 PAD.n7848 0.019716
R49030 PAD.n8054 PAD.n8053 0.019716
R49031 PAD.n8053 PAD.n7847 0.019716
R49032 PAD.n7933 PAD.n7932 0.019716
R49033 PAD.n7932 PAD.n7846 0.019716
R49034 PAD.n8045 PAD.n8044 0.019716
R49035 PAD.n8044 PAD.n7845 0.019716
R49036 PAD.n7938 PAD.n7937 0.019716
R49037 PAD.n7937 PAD.n7844 0.019716
R49038 PAD.n8036 PAD.n8035 0.019716
R49039 PAD.n8035 PAD.n7843 0.019716
R49040 PAD.n7943 PAD.n7942 0.019716
R49041 PAD.n7942 PAD.n7842 0.019716
R49042 PAD.n8027 PAD.n8026 0.019716
R49043 PAD.n8026 PAD.n7841 0.019716
R49044 PAD.n7948 PAD.n7947 0.019716
R49045 PAD.n7947 PAD.n7840 0.019716
R49046 PAD.n8018 PAD.n8017 0.019716
R49047 PAD.n8017 PAD.n7839 0.019716
R49048 PAD.n7953 PAD.n7952 0.019716
R49049 PAD.n7952 PAD.n7838 0.019716
R49050 PAD.n8009 PAD.n8008 0.019716
R49051 PAD.n8008 PAD.n7837 0.019716
R49052 PAD.n7958 PAD.n7957 0.019716
R49053 PAD.n7957 PAD.n7836 0.019716
R49054 PAD.n8000 PAD.n7999 0.019716
R49055 PAD.n7999 PAD.n7835 0.019716
R49056 PAD.n7963 PAD.n7962 0.019716
R49057 PAD.n7962 PAD.n7834 0.019716
R49058 PAD.n7991 PAD.n7990 0.019716
R49059 PAD.n7990 PAD.n7833 0.019716
R49060 PAD.n7968 PAD.n7967 0.019716
R49061 PAD.n7967 PAD.n7832 0.019716
R49062 PAD.n7982 PAD.n7981 0.019716
R49063 PAD.n7981 PAD.n7831 0.019716
R49064 PAD.n7975 PAD.n7974 0.019716
R49065 PAD.n7974 PAD.n7830 0.019716
R49066 PAD.n5540 PAD.n5213 0.019716
R49067 PAD.n5539 PAD.n5538 0.019716
R49068 PAD.n5538 PAD.n5537 0.019716
R49069 PAD.n5528 PAD.n5214 0.019716
R49070 PAD.n5529 PAD.n5528 0.019716
R49071 PAD.n5527 PAD.n5526 0.019716
R49072 PAD.n5526 PAD.n5525 0.019716
R49073 PAD.n5516 PAD.n5219 0.019716
R49074 PAD.n5517 PAD.n5516 0.019716
R49075 PAD.n5515 PAD.n5514 0.019716
R49076 PAD.n5514 PAD.n5513 0.019716
R49077 PAD.n5504 PAD.n5223 0.019716
R49078 PAD.n5505 PAD.n5504 0.019716
R49079 PAD.n5503 PAD.n5502 0.019716
R49080 PAD.n5502 PAD.n5501 0.019716
R49081 PAD.n5492 PAD.n5227 0.019716
R49082 PAD.n5493 PAD.n5492 0.019716
R49083 PAD.n5491 PAD.n5490 0.019716
R49084 PAD.n5490 PAD.n5489 0.019716
R49085 PAD.n5480 PAD.n5231 0.019716
R49086 PAD.n5481 PAD.n5480 0.019716
R49087 PAD.n5479 PAD.n5478 0.019716
R49088 PAD.n5478 PAD.n5477 0.019716
R49089 PAD.n5468 PAD.n5235 0.019716
R49090 PAD.n5469 PAD.n5468 0.019716
R49091 PAD.n5467 PAD.n5466 0.019716
R49092 PAD.n5466 PAD.n5465 0.019716
R49093 PAD.n5456 PAD.n5239 0.019716
R49094 PAD.n5457 PAD.n5456 0.019716
R49095 PAD.n5455 PAD.n5454 0.019716
R49096 PAD.n5454 PAD.n5453 0.019716
R49097 PAD.n5444 PAD.n5243 0.019716
R49098 PAD.n5445 PAD.n5444 0.019716
R49099 PAD.n5443 PAD.n5442 0.019716
R49100 PAD.n5442 PAD.n5441 0.019716
R49101 PAD.n5432 PAD.n5247 0.019716
R49102 PAD.n5433 PAD.n5432 0.019716
R49103 PAD.n5431 PAD.n5430 0.019716
R49104 PAD.n5430 PAD.n5429 0.019716
R49105 PAD.n5420 PAD.n5251 0.019716
R49106 PAD.n5421 PAD.n5420 0.019716
R49107 PAD.n5419 PAD.n5418 0.019716
R49108 PAD.n5418 PAD.n5417 0.019716
R49109 PAD.n5408 PAD.n5255 0.019716
R49110 PAD.n5409 PAD.n5408 0.019716
R49111 PAD.n5407 PAD.n5406 0.019716
R49112 PAD.n5406 PAD.n5405 0.019716
R49113 PAD.n5396 PAD.n5259 0.019716
R49114 PAD.n5397 PAD.n5396 0.019716
R49115 PAD.n5395 PAD.n5394 0.019716
R49116 PAD.n5394 PAD.n5393 0.019716
R49117 PAD.n5384 PAD.n5263 0.019716
R49118 PAD.n5385 PAD.n5384 0.019716
R49119 PAD.n5383 PAD.n5382 0.019716
R49120 PAD.n5382 PAD.n5381 0.019716
R49121 PAD.n5372 PAD.n5267 0.019716
R49122 PAD.n5373 PAD.n5372 0.019716
R49123 PAD.n5371 PAD.n5370 0.019716
R49124 PAD.n5370 PAD.n5369 0.019716
R49125 PAD.n5360 PAD.n5271 0.019716
R49126 PAD.n5361 PAD.n5360 0.019716
R49127 PAD.n5359 PAD.n5358 0.019716
R49128 PAD.n5358 PAD.n5357 0.019716
R49129 PAD.n5348 PAD.n5275 0.019716
R49130 PAD.n5349 PAD.n5348 0.019716
R49131 PAD.n5347 PAD.n5346 0.019716
R49132 PAD.n5346 PAD.n5345 0.019716
R49133 PAD.n5336 PAD.n5279 0.019716
R49134 PAD.n5337 PAD.n5336 0.019716
R49135 PAD.n5335 PAD.n5334 0.019716
R49136 PAD.n5334 PAD.n5333 0.019716
R49137 PAD.n5324 PAD.n5283 0.019716
R49138 PAD.n5325 PAD.n5324 0.019716
R49139 PAD.n5323 PAD.n5322 0.019716
R49140 PAD.n5322 PAD.n5321 0.019716
R49141 PAD.n5312 PAD.n5287 0.019716
R49142 PAD.n5313 PAD.n5312 0.019716
R49143 PAD.n5311 PAD.n5310 0.019716
R49144 PAD.n5310 PAD.n5309 0.019716
R49145 PAD.n5300 PAD.n5291 0.019716
R49146 PAD.n5301 PAD.n5300 0.019716
R49147 PAD.n5299 PAD.n5298 0.019716
R49148 PAD.n5298 PAD.n5297 0.019716
R49149 PAD.n7781 PAD.n7104 0.019716
R49150 PAD.n7774 PAD.n7773 0.019716
R49151 PAD.n7774 PAD.n7102 0.019716
R49152 PAD.n7770 PAD.n7769 0.019716
R49153 PAD.n7769 PAD.n7101 0.019716
R49154 PAD.n7763 PAD.n7762 0.019716
R49155 PAD.n7763 PAD.n7100 0.019716
R49156 PAD.n7758 PAD.n7757 0.019716
R49157 PAD.n7757 PAD.n7099 0.019716
R49158 PAD.n7751 PAD.n7750 0.019716
R49159 PAD.n7751 PAD.n7098 0.019716
R49160 PAD.n7746 PAD.n7745 0.019716
R49161 PAD.n7745 PAD.n7097 0.019716
R49162 PAD.n7739 PAD.n7738 0.019716
R49163 PAD.n7739 PAD.n7096 0.019716
R49164 PAD.n7734 PAD.n7733 0.019716
R49165 PAD.n7733 PAD.n7095 0.019716
R49166 PAD.n7727 PAD.n7726 0.019716
R49167 PAD.n7727 PAD.n7094 0.019716
R49168 PAD.n7722 PAD.n7721 0.019716
R49169 PAD.n7721 PAD.n7093 0.019716
R49170 PAD.n7715 PAD.n7714 0.019716
R49171 PAD.n7715 PAD.n7092 0.019716
R49172 PAD.n7710 PAD.n7709 0.019716
R49173 PAD.n7709 PAD.n7091 0.019716
R49174 PAD.n7703 PAD.n7702 0.019716
R49175 PAD.n7703 PAD.n7090 0.019716
R49176 PAD.n7698 PAD.n7697 0.019716
R49177 PAD.n7697 PAD.n7089 0.019716
R49178 PAD.n7691 PAD.n7690 0.019716
R49179 PAD.n7691 PAD.n7088 0.019716
R49180 PAD.n7686 PAD.n7685 0.019716
R49181 PAD.n7685 PAD.n7087 0.019716
R49182 PAD.n7679 PAD.n7678 0.019716
R49183 PAD.n7679 PAD.n7086 0.019716
R49184 PAD.n7674 PAD.n7673 0.019716
R49185 PAD.n7673 PAD.n7085 0.019716
R49186 PAD.n7667 PAD.n7666 0.019716
R49187 PAD.n7667 PAD.n7084 0.019716
R49188 PAD.n7662 PAD.n7661 0.019716
R49189 PAD.n7661 PAD.n7083 0.019716
R49190 PAD.n7655 PAD.n7654 0.019716
R49191 PAD.n7655 PAD.n7082 0.019716
R49192 PAD.n7650 PAD.n7649 0.019716
R49193 PAD.n7649 PAD.n7081 0.019716
R49194 PAD.n7643 PAD.n7642 0.019716
R49195 PAD.n7643 PAD.n7080 0.019716
R49196 PAD.n7638 PAD.n7637 0.019716
R49197 PAD.n7637 PAD.n7079 0.019716
R49198 PAD.n7631 PAD.n7630 0.019716
R49199 PAD.n7631 PAD.n7078 0.019716
R49200 PAD.n7626 PAD.n7625 0.019716
R49201 PAD.n7625 PAD.n7077 0.019716
R49202 PAD.n7619 PAD.n7618 0.019716
R49203 PAD.n7619 PAD.n7076 0.019716
R49204 PAD.n7614 PAD.n7613 0.019716
R49205 PAD.n7613 PAD.n7075 0.019716
R49206 PAD.n7607 PAD.n7606 0.019716
R49207 PAD.n7607 PAD.n7074 0.019716
R49208 PAD.n7602 PAD.n7601 0.019716
R49209 PAD.n7601 PAD.n7073 0.019716
R49210 PAD.n7595 PAD.n7594 0.019716
R49211 PAD.n7595 PAD.n7072 0.019716
R49212 PAD.n7590 PAD.n7589 0.019716
R49213 PAD.n7589 PAD.n7071 0.019716
R49214 PAD.n7583 PAD.n7582 0.019716
R49215 PAD.n7583 PAD.n7070 0.019716
R49216 PAD.n7578 PAD.n7577 0.019716
R49217 PAD.n7577 PAD.n7069 0.019716
R49218 PAD.n7571 PAD.n7570 0.019716
R49219 PAD.n7571 PAD.n7068 0.019716
R49220 PAD.n7566 PAD.n7565 0.019716
R49221 PAD.n7565 PAD.n7067 0.019716
R49222 PAD.n7559 PAD.n7558 0.019716
R49223 PAD.n7559 PAD.n7066 0.019716
R49224 PAD.n7554 PAD.n7553 0.019716
R49225 PAD.n7553 PAD.n7065 0.019716
R49226 PAD.n7547 PAD.n7546 0.019716
R49227 PAD.n7547 PAD.n7064 0.019716
R49228 PAD.n7542 PAD.n7541 0.019716
R49229 PAD.n7541 PAD.n7063 0.019716
R49230 PAD.n7535 PAD.n7534 0.019716
R49231 PAD.n7535 PAD.n7062 0.019716
R49232 PAD.n7048 PAD.n6721 0.019716
R49233 PAD.n7047 PAD.n7046 0.019716
R49234 PAD.n7046 PAD.n7045 0.019716
R49235 PAD.n7036 PAD.n6722 0.019716
R49236 PAD.n7037 PAD.n7036 0.019716
R49237 PAD.n7035 PAD.n7034 0.019716
R49238 PAD.n7034 PAD.n7033 0.019716
R49239 PAD.n7024 PAD.n6727 0.019716
R49240 PAD.n7025 PAD.n7024 0.019716
R49241 PAD.n7023 PAD.n7022 0.019716
R49242 PAD.n7022 PAD.n7021 0.019716
R49243 PAD.n7012 PAD.n6731 0.019716
R49244 PAD.n7013 PAD.n7012 0.019716
R49245 PAD.n7011 PAD.n7010 0.019716
R49246 PAD.n7010 PAD.n7009 0.019716
R49247 PAD.n7000 PAD.n6735 0.019716
R49248 PAD.n7001 PAD.n7000 0.019716
R49249 PAD.n6999 PAD.n6998 0.019716
R49250 PAD.n6998 PAD.n6997 0.019716
R49251 PAD.n6988 PAD.n6739 0.019716
R49252 PAD.n6989 PAD.n6988 0.019716
R49253 PAD.n6987 PAD.n6986 0.019716
R49254 PAD.n6986 PAD.n6985 0.019716
R49255 PAD.n6976 PAD.n6743 0.019716
R49256 PAD.n6977 PAD.n6976 0.019716
R49257 PAD.n6975 PAD.n6974 0.019716
R49258 PAD.n6974 PAD.n6973 0.019716
R49259 PAD.n6964 PAD.n6747 0.019716
R49260 PAD.n6965 PAD.n6964 0.019716
R49261 PAD.n6963 PAD.n6962 0.019716
R49262 PAD.n6962 PAD.n6961 0.019716
R49263 PAD.n6952 PAD.n6751 0.019716
R49264 PAD.n6953 PAD.n6952 0.019716
R49265 PAD.n6951 PAD.n6950 0.019716
R49266 PAD.n6950 PAD.n6949 0.019716
R49267 PAD.n6940 PAD.n6755 0.019716
R49268 PAD.n6941 PAD.n6940 0.019716
R49269 PAD.n6939 PAD.n6938 0.019716
R49270 PAD.n6938 PAD.n6937 0.019716
R49271 PAD.n6928 PAD.n6759 0.019716
R49272 PAD.n6929 PAD.n6928 0.019716
R49273 PAD.n6927 PAD.n6926 0.019716
R49274 PAD.n6926 PAD.n6925 0.019716
R49275 PAD.n6916 PAD.n6763 0.019716
R49276 PAD.n6917 PAD.n6916 0.019716
R49277 PAD.n6915 PAD.n6914 0.019716
R49278 PAD.n6914 PAD.n6913 0.019716
R49279 PAD.n6904 PAD.n6767 0.019716
R49280 PAD.n6905 PAD.n6904 0.019716
R49281 PAD.n6903 PAD.n6902 0.019716
R49282 PAD.n6902 PAD.n6901 0.019716
R49283 PAD.n6892 PAD.n6771 0.019716
R49284 PAD.n6893 PAD.n6892 0.019716
R49285 PAD.n6891 PAD.n6890 0.019716
R49286 PAD.n6890 PAD.n6889 0.019716
R49287 PAD.n6880 PAD.n6775 0.019716
R49288 PAD.n6881 PAD.n6880 0.019716
R49289 PAD.n6879 PAD.n6878 0.019716
R49290 PAD.n6878 PAD.n6877 0.019716
R49291 PAD.n6868 PAD.n6779 0.019716
R49292 PAD.n6869 PAD.n6868 0.019716
R49293 PAD.n6867 PAD.n6866 0.019716
R49294 PAD.n6866 PAD.n6865 0.019716
R49295 PAD.n6856 PAD.n6783 0.019716
R49296 PAD.n6857 PAD.n6856 0.019716
R49297 PAD.n6855 PAD.n6854 0.019716
R49298 PAD.n6854 PAD.n6853 0.019716
R49299 PAD.n6844 PAD.n6787 0.019716
R49300 PAD.n6845 PAD.n6844 0.019716
R49301 PAD.n6843 PAD.n6842 0.019716
R49302 PAD.n6842 PAD.n6841 0.019716
R49303 PAD.n6832 PAD.n6791 0.019716
R49304 PAD.n6833 PAD.n6832 0.019716
R49305 PAD.n6831 PAD.n6830 0.019716
R49306 PAD.n6830 PAD.n6829 0.019716
R49307 PAD.n6820 PAD.n6795 0.019716
R49308 PAD.n6821 PAD.n6820 0.019716
R49309 PAD.n6819 PAD.n6818 0.019716
R49310 PAD.n6818 PAD.n6817 0.019716
R49311 PAD.n6808 PAD.n6799 0.019716
R49312 PAD.n6809 PAD.n6808 0.019716
R49313 PAD.n6807 PAD.n6806 0.019716
R49314 PAD.n6806 PAD.n6805 0.019716
R49315 PAD.n5893 PAD.n5602 0.019716
R49316 PAD.n5604 PAD.n5603 0.019716
R49317 PAD.n5604 PAD.n5601 0.019716
R49318 PAD.n5884 PAD.n5883 0.019716
R49319 PAD.n5883 PAD.n5600 0.019716
R49320 PAD.n5609 PAD.n5608 0.019716
R49321 PAD.n5608 PAD.n5599 0.019716
R49322 PAD.n5875 PAD.n5874 0.019716
R49323 PAD.n5874 PAD.n5598 0.019716
R49324 PAD.n5614 PAD.n5613 0.019716
R49325 PAD.n5613 PAD.n5597 0.019716
R49326 PAD.n5866 PAD.n5865 0.019716
R49327 PAD.n5865 PAD.n5596 0.019716
R49328 PAD.n5619 PAD.n5618 0.019716
R49329 PAD.n5618 PAD.n5595 0.019716
R49330 PAD.n5857 PAD.n5856 0.019716
R49331 PAD.n5856 PAD.n5594 0.019716
R49332 PAD.n5624 PAD.n5623 0.019716
R49333 PAD.n5623 PAD.n5593 0.019716
R49334 PAD.n5848 PAD.n5847 0.019716
R49335 PAD.n5847 PAD.n5592 0.019716
R49336 PAD.n5629 PAD.n5628 0.019716
R49337 PAD.n5628 PAD.n5591 0.019716
R49338 PAD.n5839 PAD.n5838 0.019716
R49339 PAD.n5838 PAD.n5590 0.019716
R49340 PAD.n5634 PAD.n5633 0.019716
R49341 PAD.n5633 PAD.n5589 0.019716
R49342 PAD.n5830 PAD.n5829 0.019716
R49343 PAD.n5829 PAD.n5588 0.019716
R49344 PAD.n5639 PAD.n5638 0.019716
R49345 PAD.n5638 PAD.n5587 0.019716
R49346 PAD.n5821 PAD.n5820 0.019716
R49347 PAD.n5820 PAD.n5586 0.019716
R49348 PAD.n5644 PAD.n5643 0.019716
R49349 PAD.n5643 PAD.n5585 0.019716
R49350 PAD.n5812 PAD.n5811 0.019716
R49351 PAD.n5811 PAD.n5584 0.019716
R49352 PAD.n5649 PAD.n5648 0.019716
R49353 PAD.n5648 PAD.n5583 0.019716
R49354 PAD.n5803 PAD.n5802 0.019716
R49355 PAD.n5802 PAD.n5582 0.019716
R49356 PAD.n5654 PAD.n5653 0.019716
R49357 PAD.n5653 PAD.n5581 0.019716
R49358 PAD.n5794 PAD.n5793 0.019716
R49359 PAD.n5793 PAD.n5580 0.019716
R49360 PAD.n5659 PAD.n5658 0.019716
R49361 PAD.n5658 PAD.n5579 0.019716
R49362 PAD.n5785 PAD.n5784 0.019716
R49363 PAD.n5784 PAD.n5578 0.019716
R49364 PAD.n5664 PAD.n5663 0.019716
R49365 PAD.n5663 PAD.n5577 0.019716
R49366 PAD.n5776 PAD.n5775 0.019716
R49367 PAD.n5775 PAD.n5576 0.019716
R49368 PAD.n5669 PAD.n5668 0.019716
R49369 PAD.n5668 PAD.n5575 0.019716
R49370 PAD.n5767 PAD.n5766 0.019716
R49371 PAD.n5766 PAD.n5574 0.019716
R49372 PAD.n5674 PAD.n5673 0.019716
R49373 PAD.n5673 PAD.n5573 0.019716
R49374 PAD.n5758 PAD.n5757 0.019716
R49375 PAD.n5757 PAD.n5572 0.019716
R49376 PAD.n5679 PAD.n5678 0.019716
R49377 PAD.n5678 PAD.n5571 0.019716
R49378 PAD.n5749 PAD.n5748 0.019716
R49379 PAD.n5748 PAD.n5570 0.019716
R49380 PAD.n5684 PAD.n5683 0.019716
R49381 PAD.n5683 PAD.n5569 0.019716
R49382 PAD.n5740 PAD.n5739 0.019716
R49383 PAD.n5739 PAD.n5568 0.019716
R49384 PAD.n5689 PAD.n5688 0.019716
R49385 PAD.n5688 PAD.n5567 0.019716
R49386 PAD.n5731 PAD.n5730 0.019716
R49387 PAD.n5730 PAD.n5566 0.019716
R49388 PAD.n5694 PAD.n5693 0.019716
R49389 PAD.n5693 PAD.n5565 0.019716
R49390 PAD.n5722 PAD.n5721 0.019716
R49391 PAD.n5721 PAD.n5564 0.019716
R49392 PAD.n5699 PAD.n5698 0.019716
R49393 PAD.n5698 PAD.n5563 0.019716
R49394 PAD.n5713 PAD.n5712 0.019716
R49395 PAD.n5712 PAD.n5562 0.019716
R49396 PAD.n5706 PAD.n5705 0.019716
R49397 PAD.n5705 PAD.n5561 0.019716
R49398 PAD.n11084 PAD.n11083 0.019716
R49399 PAD.n11083 PAD.n11082 0.019716
R49400 PAD.n11073 PAD.n10756 0.019716
R49401 PAD.n11074 PAD.n11073 0.019716
R49402 PAD.n11072 PAD.n11071 0.019716
R49403 PAD.n11071 PAD.n11070 0.019716
R49404 PAD.n11061 PAD.n10760 0.019716
R49405 PAD.n11062 PAD.n11061 0.019716
R49406 PAD.n11060 PAD.n11059 0.019716
R49407 PAD.n11059 PAD.n11058 0.019716
R49408 PAD.n11049 PAD.n10764 0.019716
R49409 PAD.n11050 PAD.n11049 0.019716
R49410 PAD.n11048 PAD.n11047 0.019716
R49411 PAD.n11047 PAD.n11046 0.019716
R49412 PAD.n11037 PAD.n10768 0.019716
R49413 PAD.n11038 PAD.n11037 0.019716
R49414 PAD.n11036 PAD.n11035 0.019716
R49415 PAD.n11035 PAD.n11034 0.019716
R49416 PAD.n11025 PAD.n10772 0.019716
R49417 PAD.n11026 PAD.n11025 0.019716
R49418 PAD.n11024 PAD.n11023 0.019716
R49419 PAD.n11023 PAD.n11022 0.019716
R49420 PAD.n11013 PAD.n10776 0.019716
R49421 PAD.n11014 PAD.n11013 0.019716
R49422 PAD.n11012 PAD.n11011 0.019716
R49423 PAD.n11011 PAD.n11010 0.019716
R49424 PAD.n11001 PAD.n10780 0.019716
R49425 PAD.n11002 PAD.n11001 0.019716
R49426 PAD.n11000 PAD.n10999 0.019716
R49427 PAD.n10999 PAD.n10998 0.019716
R49428 PAD.n10989 PAD.n10784 0.019716
R49429 PAD.n10990 PAD.n10989 0.019716
R49430 PAD.n10988 PAD.n10987 0.019716
R49431 PAD.n10987 PAD.n10986 0.019716
R49432 PAD.n10977 PAD.n10788 0.019716
R49433 PAD.n10978 PAD.n10977 0.019716
R49434 PAD.n10976 PAD.n10975 0.019716
R49435 PAD.n10975 PAD.n10974 0.019716
R49436 PAD.n10965 PAD.n10792 0.019716
R49437 PAD.n10966 PAD.n10965 0.019716
R49438 PAD.n10964 PAD.n10963 0.019716
R49439 PAD.n10963 PAD.n10962 0.019716
R49440 PAD.n10953 PAD.n10796 0.019716
R49441 PAD.n10954 PAD.n10953 0.019716
R49442 PAD.n10952 PAD.n10951 0.019716
R49443 PAD.n10951 PAD.n10950 0.019716
R49444 PAD.n10941 PAD.n10800 0.019716
R49445 PAD.n10942 PAD.n10941 0.019716
R49446 PAD.n10940 PAD.n10939 0.019716
R49447 PAD.n10939 PAD.n10938 0.019716
R49448 PAD.n10929 PAD.n10804 0.019716
R49449 PAD.n10930 PAD.n10929 0.019716
R49450 PAD.n10928 PAD.n10927 0.019716
R49451 PAD.n10927 PAD.n10926 0.019716
R49452 PAD.n10917 PAD.n10808 0.019716
R49453 PAD.n10918 PAD.n10917 0.019716
R49454 PAD.n10916 PAD.n10915 0.019716
R49455 PAD.n10915 PAD.n10914 0.019716
R49456 PAD.n10905 PAD.n10812 0.019716
R49457 PAD.n10906 PAD.n10905 0.019716
R49458 PAD.n10904 PAD.n10903 0.019716
R49459 PAD.n10903 PAD.n10902 0.019716
R49460 PAD.n10893 PAD.n10816 0.019716
R49461 PAD.n10894 PAD.n10893 0.019716
R49462 PAD.n10892 PAD.n10891 0.019716
R49463 PAD.n10891 PAD.n10890 0.019716
R49464 PAD.n10881 PAD.n10820 0.019716
R49465 PAD.n10882 PAD.n10881 0.019716
R49466 PAD.n10880 PAD.n10879 0.019716
R49467 PAD.n10879 PAD.n10878 0.019716
R49468 PAD.n10869 PAD.n10824 0.019716
R49469 PAD.n10870 PAD.n10869 0.019716
R49470 PAD.n10868 PAD.n10867 0.019716
R49471 PAD.n10867 PAD.n10866 0.019716
R49472 PAD.n10857 PAD.n10828 0.019716
R49473 PAD.n10858 PAD.n10857 0.019716
R49474 PAD.n10856 PAD.n10855 0.019716
R49475 PAD.n10855 PAD.n10854 0.019716
R49476 PAD.n10845 PAD.n10832 0.019716
R49477 PAD.n10846 PAD.n10845 0.019716
R49478 PAD.n10844 PAD.n10843 0.019716
R49479 PAD.n10843 PAD.n10842 0.019716
R49480 PAD.n10837 PAD.n10836 0.019716
R49481 PAD.n5905 PAD.n5902 0.019716
R49482 PAD.n5906 PAD.n5905 0.019716
R49483 PAD.n6495 PAD.n6397 0.019716
R49484 PAD.n6495 PAD.n5907 0.019716
R49485 PAD.n6504 PAD.n6398 0.019716
R49486 PAD.n6504 PAD.n5908 0.019716
R49487 PAD.n6492 PAD.n6399 0.019716
R49488 PAD.n6492 PAD.n5909 0.019716
R49489 PAD.n6513 PAD.n6400 0.019716
R49490 PAD.n6513 PAD.n5910 0.019716
R49491 PAD.n6489 PAD.n6401 0.019716
R49492 PAD.n6489 PAD.n5911 0.019716
R49493 PAD.n6522 PAD.n6402 0.019716
R49494 PAD.n6522 PAD.n5912 0.019716
R49495 PAD.n6486 PAD.n6403 0.019716
R49496 PAD.n6486 PAD.n5913 0.019716
R49497 PAD.n6531 PAD.n6404 0.019716
R49498 PAD.n6531 PAD.n5914 0.019716
R49499 PAD.n6483 PAD.n6405 0.019716
R49500 PAD.n6483 PAD.n5915 0.019716
R49501 PAD.n6540 PAD.n6406 0.019716
R49502 PAD.n6540 PAD.n5916 0.019716
R49503 PAD.n6480 PAD.n6407 0.019716
R49504 PAD.n6480 PAD.n5917 0.019716
R49505 PAD.n6549 PAD.n6408 0.019716
R49506 PAD.n6549 PAD.n5918 0.019716
R49507 PAD.n6477 PAD.n6409 0.019716
R49508 PAD.n6477 PAD.n5919 0.019716
R49509 PAD.n6558 PAD.n6410 0.019716
R49510 PAD.n6558 PAD.n5920 0.019716
R49511 PAD.n6474 PAD.n6411 0.019716
R49512 PAD.n6474 PAD.n5921 0.019716
R49513 PAD.n6567 PAD.n6412 0.019716
R49514 PAD.n6567 PAD.n5922 0.019716
R49515 PAD.n6471 PAD.n6413 0.019716
R49516 PAD.n6471 PAD.n5923 0.019716
R49517 PAD.n6576 PAD.n6414 0.019716
R49518 PAD.n6576 PAD.n5924 0.019716
R49519 PAD.n6468 PAD.n6415 0.019716
R49520 PAD.n6468 PAD.n5925 0.019716
R49521 PAD.n6585 PAD.n6416 0.019716
R49522 PAD.n6585 PAD.n5926 0.019716
R49523 PAD.n6465 PAD.n6417 0.019716
R49524 PAD.n6465 PAD.n5927 0.019716
R49525 PAD.n6594 PAD.n6418 0.019716
R49526 PAD.n6594 PAD.n5928 0.019716
R49527 PAD.n6462 PAD.n6419 0.019716
R49528 PAD.n6462 PAD.n5929 0.019716
R49529 PAD.n6603 PAD.n6420 0.019716
R49530 PAD.n6603 PAD.n5930 0.019716
R49531 PAD.n6459 PAD.n6421 0.019716
R49532 PAD.n6459 PAD.n5931 0.019716
R49533 PAD.n6612 PAD.n6422 0.019716
R49534 PAD.n6612 PAD.n5932 0.019716
R49535 PAD.n6456 PAD.n6423 0.019716
R49536 PAD.n6456 PAD.n5933 0.019716
R49537 PAD.n6621 PAD.n6424 0.019716
R49538 PAD.n6621 PAD.n5934 0.019716
R49539 PAD.n6453 PAD.n6425 0.019716
R49540 PAD.n6453 PAD.n5935 0.019716
R49541 PAD.n6630 PAD.n6426 0.019716
R49542 PAD.n6630 PAD.n5936 0.019716
R49543 PAD.n6450 PAD.n6427 0.019716
R49544 PAD.n6450 PAD.n5937 0.019716
R49545 PAD.n6639 PAD.n6428 0.019716
R49546 PAD.n6639 PAD.n5938 0.019716
R49547 PAD.n6447 PAD.n6429 0.019716
R49548 PAD.n6447 PAD.n5939 0.019716
R49549 PAD.n6648 PAD.n6430 0.019716
R49550 PAD.n6648 PAD.n5940 0.019716
R49551 PAD.n6444 PAD.n6431 0.019716
R49552 PAD.n6444 PAD.n5941 0.019716
R49553 PAD.n6657 PAD.n6432 0.019716
R49554 PAD.n6657 PAD.n5942 0.019716
R49555 PAD.n6441 PAD.n6433 0.019716
R49556 PAD.n6441 PAD.n5943 0.019716
R49557 PAD.n6666 PAD.n6434 0.019716
R49558 PAD.n6666 PAD.n5944 0.019716
R49559 PAD.n6437 PAD.n6435 0.019716
R49560 PAD.n6437 PAD.n5945 0.019716
R49561 PAD.n6677 PAD.n6436 0.019716
R49562 PAD.n6436 PAD.n5946 0.019716
R49563 PAD.n6688 PAD.n5947 0.019716
R49564 PAD.n11085 PAD.n11084 0.019716
R49565 PAD.n11081 PAD.n10756 0.019716
R49566 PAD.n11082 PAD.n11081 0.019716
R49567 PAD.n11075 PAD.n11072 0.019716
R49568 PAD.n11075 PAD.n11074 0.019716
R49569 PAD.n11069 PAD.n10760 0.019716
R49570 PAD.n11070 PAD.n11069 0.019716
R49571 PAD.n11063 PAD.n11060 0.019716
R49572 PAD.n11063 PAD.n11062 0.019716
R49573 PAD.n11057 PAD.n10764 0.019716
R49574 PAD.n11058 PAD.n11057 0.019716
R49575 PAD.n11051 PAD.n11048 0.019716
R49576 PAD.n11051 PAD.n11050 0.019716
R49577 PAD.n11045 PAD.n10768 0.019716
R49578 PAD.n11046 PAD.n11045 0.019716
R49579 PAD.n11039 PAD.n11036 0.019716
R49580 PAD.n11039 PAD.n11038 0.019716
R49581 PAD.n11033 PAD.n10772 0.019716
R49582 PAD.n11034 PAD.n11033 0.019716
R49583 PAD.n11027 PAD.n11024 0.019716
R49584 PAD.n11027 PAD.n11026 0.019716
R49585 PAD.n11021 PAD.n10776 0.019716
R49586 PAD.n11022 PAD.n11021 0.019716
R49587 PAD.n11015 PAD.n11012 0.019716
R49588 PAD.n11015 PAD.n11014 0.019716
R49589 PAD.n11009 PAD.n10780 0.019716
R49590 PAD.n11010 PAD.n11009 0.019716
R49591 PAD.n11003 PAD.n11000 0.019716
R49592 PAD.n11003 PAD.n11002 0.019716
R49593 PAD.n10997 PAD.n10784 0.019716
R49594 PAD.n10998 PAD.n10997 0.019716
R49595 PAD.n10991 PAD.n10988 0.019716
R49596 PAD.n10991 PAD.n10990 0.019716
R49597 PAD.n10985 PAD.n10788 0.019716
R49598 PAD.n10986 PAD.n10985 0.019716
R49599 PAD.n10979 PAD.n10976 0.019716
R49600 PAD.n10979 PAD.n10978 0.019716
R49601 PAD.n10973 PAD.n10792 0.019716
R49602 PAD.n10974 PAD.n10973 0.019716
R49603 PAD.n10967 PAD.n10964 0.019716
R49604 PAD.n10967 PAD.n10966 0.019716
R49605 PAD.n10961 PAD.n10796 0.019716
R49606 PAD.n10962 PAD.n10961 0.019716
R49607 PAD.n10955 PAD.n10952 0.019716
R49608 PAD.n10955 PAD.n10954 0.019716
R49609 PAD.n10949 PAD.n10800 0.019716
R49610 PAD.n10950 PAD.n10949 0.019716
R49611 PAD.n10943 PAD.n10940 0.019716
R49612 PAD.n10943 PAD.n10942 0.019716
R49613 PAD.n10937 PAD.n10804 0.019716
R49614 PAD.n10938 PAD.n10937 0.019716
R49615 PAD.n10931 PAD.n10928 0.019716
R49616 PAD.n10931 PAD.n10930 0.019716
R49617 PAD.n10925 PAD.n10808 0.019716
R49618 PAD.n10926 PAD.n10925 0.019716
R49619 PAD.n10919 PAD.n10916 0.019716
R49620 PAD.n10919 PAD.n10918 0.019716
R49621 PAD.n10913 PAD.n10812 0.019716
R49622 PAD.n10914 PAD.n10913 0.019716
R49623 PAD.n10907 PAD.n10904 0.019716
R49624 PAD.n10907 PAD.n10906 0.019716
R49625 PAD.n10901 PAD.n10816 0.019716
R49626 PAD.n10902 PAD.n10901 0.019716
R49627 PAD.n10895 PAD.n10892 0.019716
R49628 PAD.n10895 PAD.n10894 0.019716
R49629 PAD.n10889 PAD.n10820 0.019716
R49630 PAD.n10890 PAD.n10889 0.019716
R49631 PAD.n10883 PAD.n10880 0.019716
R49632 PAD.n10883 PAD.n10882 0.019716
R49633 PAD.n10877 PAD.n10824 0.019716
R49634 PAD.n10878 PAD.n10877 0.019716
R49635 PAD.n10871 PAD.n10868 0.019716
R49636 PAD.n10871 PAD.n10870 0.019716
R49637 PAD.n10865 PAD.n10828 0.019716
R49638 PAD.n10866 PAD.n10865 0.019716
R49639 PAD.n10859 PAD.n10856 0.019716
R49640 PAD.n10859 PAD.n10858 0.019716
R49641 PAD.n10853 PAD.n10832 0.019716
R49642 PAD.n10854 PAD.n10853 0.019716
R49643 PAD.n10847 PAD.n10844 0.019716
R49644 PAD.n10847 PAD.n10846 0.019716
R49645 PAD.n10841 PAD.n10836 0.019716
R49646 PAD.n10842 PAD.n10841 0.019716
R49647 PAD.n116 PAD.n74 0.019716
R49648 PAD.n117 PAD.n73 0.019716
R49649 PAD.n126 PAD.n72 0.019716
R49650 PAD.n126 PAD.n125 0.019716
R49651 PAD.n128 PAD.n71 0.019716
R49652 PAD.n129 PAD.n128 0.019716
R49653 PAD.n138 PAD.n70 0.019716
R49654 PAD.n138 PAD.n137 0.019716
R49655 PAD.n140 PAD.n69 0.019716
R49656 PAD.n141 PAD.n140 0.019716
R49657 PAD.n150 PAD.n68 0.019716
R49658 PAD.n150 PAD.n149 0.019716
R49659 PAD.n152 PAD.n67 0.019716
R49660 PAD.n153 PAD.n152 0.019716
R49661 PAD.n162 PAD.n66 0.019716
R49662 PAD.n162 PAD.n161 0.019716
R49663 PAD.n164 PAD.n65 0.019716
R49664 PAD.n165 PAD.n164 0.019716
R49665 PAD.n174 PAD.n64 0.019716
R49666 PAD.n174 PAD.n173 0.019716
R49667 PAD.n176 PAD.n63 0.019716
R49668 PAD.n177 PAD.n176 0.019716
R49669 PAD.n186 PAD.n62 0.019716
R49670 PAD.n186 PAD.n185 0.019716
R49671 PAD.n188 PAD.n61 0.019716
R49672 PAD.n189 PAD.n188 0.019716
R49673 PAD.n198 PAD.n60 0.019716
R49674 PAD.n198 PAD.n197 0.019716
R49675 PAD.n200 PAD.n59 0.019716
R49676 PAD.n201 PAD.n200 0.019716
R49677 PAD.n210 PAD.n58 0.019716
R49678 PAD.n210 PAD.n209 0.019716
R49679 PAD.n212 PAD.n57 0.019716
R49680 PAD.n213 PAD.n212 0.019716
R49681 PAD.n222 PAD.n56 0.019716
R49682 PAD.n222 PAD.n221 0.019716
R49683 PAD.n224 PAD.n55 0.019716
R49684 PAD.n225 PAD.n224 0.019716
R49685 PAD.n234 PAD.n54 0.019716
R49686 PAD.n234 PAD.n233 0.019716
R49687 PAD.n236 PAD.n53 0.019716
R49688 PAD.n237 PAD.n236 0.019716
R49689 PAD.n246 PAD.n52 0.019716
R49690 PAD.n246 PAD.n245 0.019716
R49691 PAD.n248 PAD.n51 0.019716
R49692 PAD.n249 PAD.n248 0.019716
R49693 PAD.n258 PAD.n50 0.019716
R49694 PAD.n258 PAD.n257 0.019716
R49695 PAD.n260 PAD.n49 0.019716
R49696 PAD.n261 PAD.n260 0.019716
R49697 PAD.n270 PAD.n48 0.019716
R49698 PAD.n270 PAD.n269 0.019716
R49699 PAD.n272 PAD.n47 0.019716
R49700 PAD.n273 PAD.n272 0.019716
R49701 PAD.n282 PAD.n46 0.019716
R49702 PAD.n282 PAD.n281 0.019716
R49703 PAD.n284 PAD.n45 0.019716
R49704 PAD.n285 PAD.n284 0.019716
R49705 PAD.n294 PAD.n44 0.019716
R49706 PAD.n294 PAD.n293 0.019716
R49707 PAD.n296 PAD.n43 0.019716
R49708 PAD.n297 PAD.n296 0.019716
R49709 PAD.n306 PAD.n42 0.019716
R49710 PAD.n306 PAD.n305 0.019716
R49711 PAD.n308 PAD.n41 0.019716
R49712 PAD.n309 PAD.n308 0.019716
R49713 PAD.n318 PAD.n40 0.019716
R49714 PAD.n318 PAD.n317 0.019716
R49715 PAD.n320 PAD.n39 0.019716
R49716 PAD.n321 PAD.n320 0.019716
R49717 PAD.n330 PAD.n38 0.019716
R49718 PAD.n330 PAD.n329 0.019716
R49719 PAD.n332 PAD.n37 0.019716
R49720 PAD.n333 PAD.n332 0.019716
R49721 PAD.n342 PAD.n36 0.019716
R49722 PAD.n342 PAD.n341 0.019716
R49723 PAD.n344 PAD.n35 0.019716
R49724 PAD.n345 PAD.n344 0.019716
R49725 PAD.n354 PAD.n34 0.019716
R49726 PAD.n354 PAD.n353 0.019716
R49727 PAD.n356 PAD.n33 0.019716
R49728 PAD.n357 PAD.n356 0.019716
R49729 PAD.n366 PAD.n365 0.019716
R49730 PAD.n10692 PAD.n415 0.019716
R49731 PAD.n10693 PAD.n414 0.019716
R49732 PAD.n10415 PAD.n413 0.019716
R49733 PAD.n10416 PAD.n10415 0.019716
R49734 PAD.n10684 PAD.n412 0.019716
R49735 PAD.n10685 PAD.n10684 0.019716
R49736 PAD.n10420 PAD.n411 0.019716
R49737 PAD.n10421 PAD.n10420 0.019716
R49738 PAD.n10675 PAD.n410 0.019716
R49739 PAD.n10676 PAD.n10675 0.019716
R49740 PAD.n10425 PAD.n409 0.019716
R49741 PAD.n10426 PAD.n10425 0.019716
R49742 PAD.n10666 PAD.n408 0.019716
R49743 PAD.n10667 PAD.n10666 0.019716
R49744 PAD.n10430 PAD.n407 0.019716
R49745 PAD.n10431 PAD.n10430 0.019716
R49746 PAD.n10657 PAD.n406 0.019716
R49747 PAD.n10658 PAD.n10657 0.019716
R49748 PAD.n10435 PAD.n405 0.019716
R49749 PAD.n10436 PAD.n10435 0.019716
R49750 PAD.n10648 PAD.n404 0.019716
R49751 PAD.n10649 PAD.n10648 0.019716
R49752 PAD.n10440 PAD.n403 0.019716
R49753 PAD.n10441 PAD.n10440 0.019716
R49754 PAD.n10639 PAD.n402 0.019716
R49755 PAD.n10640 PAD.n10639 0.019716
R49756 PAD.n10445 PAD.n401 0.019716
R49757 PAD.n10446 PAD.n10445 0.019716
R49758 PAD.n10630 PAD.n400 0.019716
R49759 PAD.n10631 PAD.n10630 0.019716
R49760 PAD.n10450 PAD.n399 0.019716
R49761 PAD.n10451 PAD.n10450 0.019716
R49762 PAD.n10621 PAD.n398 0.019716
R49763 PAD.n10622 PAD.n10621 0.019716
R49764 PAD.n10455 PAD.n397 0.019716
R49765 PAD.n10456 PAD.n10455 0.019716
R49766 PAD.n10612 PAD.n396 0.019716
R49767 PAD.n10613 PAD.n10612 0.019716
R49768 PAD.n10460 PAD.n395 0.019716
R49769 PAD.n10461 PAD.n10460 0.019716
R49770 PAD.n10603 PAD.n394 0.019716
R49771 PAD.n10604 PAD.n10603 0.019716
R49772 PAD.n10465 PAD.n393 0.019716
R49773 PAD.n10466 PAD.n10465 0.019716
R49774 PAD.n10594 PAD.n392 0.019716
R49775 PAD.n10595 PAD.n10594 0.019716
R49776 PAD.n10470 PAD.n391 0.019716
R49777 PAD.n10471 PAD.n10470 0.019716
R49778 PAD.n10585 PAD.n390 0.019716
R49779 PAD.n10586 PAD.n10585 0.019716
R49780 PAD.n10475 PAD.n389 0.019716
R49781 PAD.n10476 PAD.n10475 0.019716
R49782 PAD.n10576 PAD.n388 0.019716
R49783 PAD.n10577 PAD.n10576 0.019716
R49784 PAD.n10480 PAD.n387 0.019716
R49785 PAD.n10481 PAD.n10480 0.019716
R49786 PAD.n10567 PAD.n386 0.019716
R49787 PAD.n10568 PAD.n10567 0.019716
R49788 PAD.n10485 PAD.n385 0.019716
R49789 PAD.n10486 PAD.n10485 0.019716
R49790 PAD.n10558 PAD.n384 0.019716
R49791 PAD.n10559 PAD.n10558 0.019716
R49792 PAD.n10490 PAD.n383 0.019716
R49793 PAD.n10491 PAD.n10490 0.019716
R49794 PAD.n10549 PAD.n382 0.019716
R49795 PAD.n10550 PAD.n10549 0.019716
R49796 PAD.n10495 PAD.n381 0.019716
R49797 PAD.n10496 PAD.n10495 0.019716
R49798 PAD.n10540 PAD.n380 0.019716
R49799 PAD.n10541 PAD.n10540 0.019716
R49800 PAD.n10500 PAD.n379 0.019716
R49801 PAD.n10501 PAD.n10500 0.019716
R49802 PAD.n10531 PAD.n378 0.019716
R49803 PAD.n10532 PAD.n10531 0.019716
R49804 PAD.n10505 PAD.n377 0.019716
R49805 PAD.n10506 PAD.n10505 0.019716
R49806 PAD.n10522 PAD.n376 0.019716
R49807 PAD.n10523 PAD.n10522 0.019716
R49808 PAD.n10510 PAD.n375 0.019716
R49809 PAD.n10511 PAD.n10510 0.019716
R49810 PAD.n10513 PAD.n374 0.019716
R49811 PAD.n10514 PAD.n10513 0.019716
R49812 PAD.n10715 PAD.n10714 0.019716
R49813 PAD.n524 PAD.n523 0.019716
R49814 PAD.n526 PAD.n525 0.019716
R49815 PAD.n527 PAD.n517 0.019716
R49816 PAD.n528 PAD.n527 0.019716
R49817 PAD.n538 PAD.n537 0.019716
R49818 PAD.n537 PAD.n536 0.019716
R49819 PAD.n539 PAD.n513 0.019716
R49820 PAD.n540 PAD.n539 0.019716
R49821 PAD.n550 PAD.n549 0.019716
R49822 PAD.n549 PAD.n548 0.019716
R49823 PAD.n551 PAD.n509 0.019716
R49824 PAD.n552 PAD.n551 0.019716
R49825 PAD.n562 PAD.n561 0.019716
R49826 PAD.n561 PAD.n560 0.019716
R49827 PAD.n563 PAD.n505 0.019716
R49828 PAD.n564 PAD.n563 0.019716
R49829 PAD.n574 PAD.n573 0.019716
R49830 PAD.n573 PAD.n572 0.019716
R49831 PAD.n575 PAD.n501 0.019716
R49832 PAD.n576 PAD.n575 0.019716
R49833 PAD.n586 PAD.n585 0.019716
R49834 PAD.n585 PAD.n584 0.019716
R49835 PAD.n587 PAD.n497 0.019716
R49836 PAD.n588 PAD.n587 0.019716
R49837 PAD.n598 PAD.n597 0.019716
R49838 PAD.n597 PAD.n596 0.019716
R49839 PAD.n599 PAD.n493 0.019716
R49840 PAD.n600 PAD.n599 0.019716
R49841 PAD.n610 PAD.n609 0.019716
R49842 PAD.n609 PAD.n608 0.019716
R49843 PAD.n611 PAD.n489 0.019716
R49844 PAD.n612 PAD.n611 0.019716
R49845 PAD.n622 PAD.n621 0.019716
R49846 PAD.n621 PAD.n620 0.019716
R49847 PAD.n623 PAD.n485 0.019716
R49848 PAD.n624 PAD.n623 0.019716
R49849 PAD.n634 PAD.n633 0.019716
R49850 PAD.n633 PAD.n632 0.019716
R49851 PAD.n635 PAD.n481 0.019716
R49852 PAD.n636 PAD.n635 0.019716
R49853 PAD.n646 PAD.n645 0.019716
R49854 PAD.n645 PAD.n644 0.019716
R49855 PAD.n647 PAD.n477 0.019716
R49856 PAD.n648 PAD.n647 0.019716
R49857 PAD.n658 PAD.n657 0.019716
R49858 PAD.n657 PAD.n656 0.019716
R49859 PAD.n659 PAD.n473 0.019716
R49860 PAD.n660 PAD.n659 0.019716
R49861 PAD.n670 PAD.n669 0.019716
R49862 PAD.n669 PAD.n668 0.019716
R49863 PAD.n671 PAD.n469 0.019716
R49864 PAD.n672 PAD.n671 0.019716
R49865 PAD.n682 PAD.n681 0.019716
R49866 PAD.n681 PAD.n680 0.019716
R49867 PAD.n683 PAD.n465 0.019716
R49868 PAD.n684 PAD.n683 0.019716
R49869 PAD.n694 PAD.n693 0.019716
R49870 PAD.n693 PAD.n692 0.019716
R49871 PAD.n695 PAD.n461 0.019716
R49872 PAD.n696 PAD.n695 0.019716
R49873 PAD.n706 PAD.n705 0.019716
R49874 PAD.n705 PAD.n704 0.019716
R49875 PAD.n707 PAD.n457 0.019716
R49876 PAD.n708 PAD.n707 0.019716
R49877 PAD.n718 PAD.n717 0.019716
R49878 PAD.n717 PAD.n716 0.019716
R49879 PAD.n719 PAD.n453 0.019716
R49880 PAD.n720 PAD.n719 0.019716
R49881 PAD.n730 PAD.n729 0.019716
R49882 PAD.n729 PAD.n728 0.019716
R49883 PAD.n731 PAD.n449 0.019716
R49884 PAD.n732 PAD.n731 0.019716
R49885 PAD.n742 PAD.n741 0.019716
R49886 PAD.n741 PAD.n740 0.019716
R49887 PAD.n743 PAD.n445 0.019716
R49888 PAD.n744 PAD.n743 0.019716
R49889 PAD.n754 PAD.n753 0.019716
R49890 PAD.n753 PAD.n752 0.019716
R49891 PAD.n755 PAD.n441 0.019716
R49892 PAD.n756 PAD.n755 0.019716
R49893 PAD.n767 PAD.n766 0.019716
R49894 PAD.n766 PAD.n765 0.019716
R49895 PAD.n770 PAD.n769 0.019716
R49896 PAD.n869 PAD.n824 0.019716
R49897 PAD.n870 PAD.n823 0.019716
R49898 PAD.n879 PAD.n822 0.019716
R49899 PAD.n879 PAD.n878 0.019716
R49900 PAD.n881 PAD.n821 0.019716
R49901 PAD.n882 PAD.n881 0.019716
R49902 PAD.n891 PAD.n820 0.019716
R49903 PAD.n891 PAD.n890 0.019716
R49904 PAD.n893 PAD.n819 0.019716
R49905 PAD.n894 PAD.n893 0.019716
R49906 PAD.n903 PAD.n818 0.019716
R49907 PAD.n903 PAD.n902 0.019716
R49908 PAD.n905 PAD.n817 0.019716
R49909 PAD.n906 PAD.n905 0.019716
R49910 PAD.n915 PAD.n816 0.019716
R49911 PAD.n915 PAD.n914 0.019716
R49912 PAD.n917 PAD.n815 0.019716
R49913 PAD.n918 PAD.n917 0.019716
R49914 PAD.n927 PAD.n814 0.019716
R49915 PAD.n927 PAD.n926 0.019716
R49916 PAD.n929 PAD.n813 0.019716
R49917 PAD.n930 PAD.n929 0.019716
R49918 PAD.n939 PAD.n812 0.019716
R49919 PAD.n939 PAD.n938 0.019716
R49920 PAD.n941 PAD.n811 0.019716
R49921 PAD.n942 PAD.n941 0.019716
R49922 PAD.n951 PAD.n810 0.019716
R49923 PAD.n951 PAD.n950 0.019716
R49924 PAD.n953 PAD.n809 0.019716
R49925 PAD.n954 PAD.n953 0.019716
R49926 PAD.n963 PAD.n808 0.019716
R49927 PAD.n963 PAD.n962 0.019716
R49928 PAD.n965 PAD.n807 0.019716
R49929 PAD.n966 PAD.n965 0.019716
R49930 PAD.n975 PAD.n806 0.019716
R49931 PAD.n975 PAD.n974 0.019716
R49932 PAD.n977 PAD.n805 0.019716
R49933 PAD.n978 PAD.n977 0.019716
R49934 PAD.n987 PAD.n804 0.019716
R49935 PAD.n987 PAD.n986 0.019716
R49936 PAD.n989 PAD.n803 0.019716
R49937 PAD.n990 PAD.n989 0.019716
R49938 PAD.n999 PAD.n802 0.019716
R49939 PAD.n999 PAD.n998 0.019716
R49940 PAD.n1001 PAD.n801 0.019716
R49941 PAD.n1002 PAD.n1001 0.019716
R49942 PAD.n1011 PAD.n800 0.019716
R49943 PAD.n1011 PAD.n1010 0.019716
R49944 PAD.n1013 PAD.n799 0.019716
R49945 PAD.n1014 PAD.n1013 0.019716
R49946 PAD.n1023 PAD.n798 0.019716
R49947 PAD.n1023 PAD.n1022 0.019716
R49948 PAD.n1025 PAD.n797 0.019716
R49949 PAD.n1026 PAD.n1025 0.019716
R49950 PAD.n1035 PAD.n796 0.019716
R49951 PAD.n1035 PAD.n1034 0.019716
R49952 PAD.n1037 PAD.n795 0.019716
R49953 PAD.n1038 PAD.n1037 0.019716
R49954 PAD.n1047 PAD.n794 0.019716
R49955 PAD.n1047 PAD.n1046 0.019716
R49956 PAD.n1049 PAD.n793 0.019716
R49957 PAD.n1050 PAD.n1049 0.019716
R49958 PAD.n1059 PAD.n792 0.019716
R49959 PAD.n1059 PAD.n1058 0.019716
R49960 PAD.n1061 PAD.n791 0.019716
R49961 PAD.n1062 PAD.n1061 0.019716
R49962 PAD.n1071 PAD.n790 0.019716
R49963 PAD.n1071 PAD.n1070 0.019716
R49964 PAD.n1073 PAD.n789 0.019716
R49965 PAD.n1074 PAD.n1073 0.019716
R49966 PAD.n1083 PAD.n788 0.019716
R49967 PAD.n1083 PAD.n1082 0.019716
R49968 PAD.n1085 PAD.n787 0.019716
R49969 PAD.n1086 PAD.n1085 0.019716
R49970 PAD.n1095 PAD.n786 0.019716
R49971 PAD.n1095 PAD.n1094 0.019716
R49972 PAD.n1097 PAD.n785 0.019716
R49973 PAD.n1098 PAD.n1097 0.019716
R49974 PAD.n1107 PAD.n784 0.019716
R49975 PAD.n1107 PAD.n1106 0.019716
R49976 PAD.n1109 PAD.n783 0.019716
R49977 PAD.n1110 PAD.n1109 0.019716
R49978 PAD.n10387 PAD.n10386 0.019716
R49979 PAD.n10107 PAD.n10106 0.019716
R49980 PAD.n10109 PAD.n10108 0.019716
R49981 PAD.n10110 PAD.n10101 0.019716
R49982 PAD.n10111 PAD.n10110 0.019716
R49983 PAD.n10121 PAD.n10120 0.019716
R49984 PAD.n10120 PAD.n10119 0.019716
R49985 PAD.n10122 PAD.n10097 0.019716
R49986 PAD.n10123 PAD.n10122 0.019716
R49987 PAD.n10133 PAD.n10132 0.019716
R49988 PAD.n10132 PAD.n10131 0.019716
R49989 PAD.n10134 PAD.n10093 0.019716
R49990 PAD.n10135 PAD.n10134 0.019716
R49991 PAD.n10145 PAD.n10144 0.019716
R49992 PAD.n10144 PAD.n10143 0.019716
R49993 PAD.n10146 PAD.n10089 0.019716
R49994 PAD.n10147 PAD.n10146 0.019716
R49995 PAD.n10157 PAD.n10156 0.019716
R49996 PAD.n10156 PAD.n10155 0.019716
R49997 PAD.n10158 PAD.n10085 0.019716
R49998 PAD.n10159 PAD.n10158 0.019716
R49999 PAD.n10169 PAD.n10168 0.019716
R50000 PAD.n10168 PAD.n10167 0.019716
R50001 PAD.n10170 PAD.n10081 0.019716
R50002 PAD.n10171 PAD.n10170 0.019716
R50003 PAD.n10181 PAD.n10180 0.019716
R50004 PAD.n10180 PAD.n10179 0.019716
R50005 PAD.n10182 PAD.n10077 0.019716
R50006 PAD.n10183 PAD.n10182 0.019716
R50007 PAD.n10193 PAD.n10192 0.019716
R50008 PAD.n10192 PAD.n10191 0.019716
R50009 PAD.n10194 PAD.n10073 0.019716
R50010 PAD.n10195 PAD.n10194 0.019716
R50011 PAD.n10205 PAD.n10204 0.019716
R50012 PAD.n10204 PAD.n10203 0.019716
R50013 PAD.n10206 PAD.n10069 0.019716
R50014 PAD.n10207 PAD.n10206 0.019716
R50015 PAD.n10217 PAD.n10216 0.019716
R50016 PAD.n10216 PAD.n10215 0.019716
R50017 PAD.n10218 PAD.n10065 0.019716
R50018 PAD.n10219 PAD.n10218 0.019716
R50019 PAD.n10229 PAD.n10228 0.019716
R50020 PAD.n10228 PAD.n10227 0.019716
R50021 PAD.n10230 PAD.n10061 0.019716
R50022 PAD.n10231 PAD.n10230 0.019716
R50023 PAD.n10241 PAD.n10240 0.019716
R50024 PAD.n10240 PAD.n10239 0.019716
R50025 PAD.n10242 PAD.n10057 0.019716
R50026 PAD.n10243 PAD.n10242 0.019716
R50027 PAD.n10253 PAD.n10252 0.019716
R50028 PAD.n10252 PAD.n10251 0.019716
R50029 PAD.n10254 PAD.n10053 0.019716
R50030 PAD.n10255 PAD.n10254 0.019716
R50031 PAD.n10265 PAD.n10264 0.019716
R50032 PAD.n10264 PAD.n10263 0.019716
R50033 PAD.n10266 PAD.n10049 0.019716
R50034 PAD.n10267 PAD.n10266 0.019716
R50035 PAD.n10277 PAD.n10276 0.019716
R50036 PAD.n10276 PAD.n10275 0.019716
R50037 PAD.n10278 PAD.n10045 0.019716
R50038 PAD.n10279 PAD.n10278 0.019716
R50039 PAD.n10289 PAD.n10288 0.019716
R50040 PAD.n10288 PAD.n10287 0.019716
R50041 PAD.n10290 PAD.n10041 0.019716
R50042 PAD.n10291 PAD.n10290 0.019716
R50043 PAD.n10301 PAD.n10300 0.019716
R50044 PAD.n10300 PAD.n10299 0.019716
R50045 PAD.n10302 PAD.n10037 0.019716
R50046 PAD.n10303 PAD.n10302 0.019716
R50047 PAD.n10313 PAD.n10312 0.019716
R50048 PAD.n10312 PAD.n10311 0.019716
R50049 PAD.n10314 PAD.n10033 0.019716
R50050 PAD.n10315 PAD.n10314 0.019716
R50051 PAD.n10325 PAD.n10324 0.019716
R50052 PAD.n10324 PAD.n10323 0.019716
R50053 PAD.n10326 PAD.n10029 0.019716
R50054 PAD.n10327 PAD.n10326 0.019716
R50055 PAD.n10337 PAD.n10336 0.019716
R50056 PAD.n10336 PAD.n10335 0.019716
R50057 PAD.n10338 PAD.n10025 0.019716
R50058 PAD.n10339 PAD.n10338 0.019716
R50059 PAD.n10350 PAD.n10349 0.019716
R50060 PAD.n10349 PAD.n10348 0.019716
R50061 PAD.n10353 PAD.n10352 0.019716
R50062 PAD.n1482 PAD.n1481 0.019716
R50063 PAD.n1191 PAD.n1190 0.019716
R50064 PAD.n1474 PAD.n1473 0.019716
R50065 PAD.n1474 PAD.n1189 0.019716
R50066 PAD.n1198 PAD.n1197 0.019716
R50067 PAD.n1198 PAD.n1188 0.019716
R50068 PAD.n1465 PAD.n1464 0.019716
R50069 PAD.n1465 PAD.n1187 0.019716
R50070 PAD.n1203 PAD.n1202 0.019716
R50071 PAD.n1203 PAD.n1186 0.019716
R50072 PAD.n1456 PAD.n1455 0.019716
R50073 PAD.n1456 PAD.n1185 0.019716
R50074 PAD.n1208 PAD.n1207 0.019716
R50075 PAD.n1208 PAD.n1184 0.019716
R50076 PAD.n1447 PAD.n1446 0.019716
R50077 PAD.n1447 PAD.n1183 0.019716
R50078 PAD.n1213 PAD.n1212 0.019716
R50079 PAD.n1213 PAD.n1182 0.019716
R50080 PAD.n1438 PAD.n1437 0.019716
R50081 PAD.n1438 PAD.n1181 0.019716
R50082 PAD.n1218 PAD.n1217 0.019716
R50083 PAD.n1218 PAD.n1180 0.019716
R50084 PAD.n1429 PAD.n1428 0.019716
R50085 PAD.n1429 PAD.n1179 0.019716
R50086 PAD.n1223 PAD.n1222 0.019716
R50087 PAD.n1223 PAD.n1178 0.019716
R50088 PAD.n1420 PAD.n1419 0.019716
R50089 PAD.n1420 PAD.n1177 0.019716
R50090 PAD.n1228 PAD.n1227 0.019716
R50091 PAD.n1228 PAD.n1176 0.019716
R50092 PAD.n1411 PAD.n1410 0.019716
R50093 PAD.n1411 PAD.n1175 0.019716
R50094 PAD.n1233 PAD.n1232 0.019716
R50095 PAD.n1233 PAD.n1174 0.019716
R50096 PAD.n1402 PAD.n1401 0.019716
R50097 PAD.n1402 PAD.n1173 0.019716
R50098 PAD.n1238 PAD.n1237 0.019716
R50099 PAD.n1238 PAD.n1172 0.019716
R50100 PAD.n1393 PAD.n1392 0.019716
R50101 PAD.n1393 PAD.n1171 0.019716
R50102 PAD.n1243 PAD.n1242 0.019716
R50103 PAD.n1243 PAD.n1170 0.019716
R50104 PAD.n1384 PAD.n1383 0.019716
R50105 PAD.n1384 PAD.n1169 0.019716
R50106 PAD.n1248 PAD.n1247 0.019716
R50107 PAD.n1248 PAD.n1168 0.019716
R50108 PAD.n1375 PAD.n1374 0.019716
R50109 PAD.n1375 PAD.n1167 0.019716
R50110 PAD.n1253 PAD.n1252 0.019716
R50111 PAD.n1253 PAD.n1166 0.019716
R50112 PAD.n1366 PAD.n1365 0.019716
R50113 PAD.n1366 PAD.n1165 0.019716
R50114 PAD.n1258 PAD.n1257 0.019716
R50115 PAD.n1258 PAD.n1164 0.019716
R50116 PAD.n1357 PAD.n1356 0.019716
R50117 PAD.n1357 PAD.n1163 0.019716
R50118 PAD.n1263 PAD.n1262 0.019716
R50119 PAD.n1263 PAD.n1162 0.019716
R50120 PAD.n1348 PAD.n1347 0.019716
R50121 PAD.n1348 PAD.n1161 0.019716
R50122 PAD.n1268 PAD.n1267 0.019716
R50123 PAD.n1268 PAD.n1160 0.019716
R50124 PAD.n1339 PAD.n1338 0.019716
R50125 PAD.n1339 PAD.n1159 0.019716
R50126 PAD.n1273 PAD.n1272 0.019716
R50127 PAD.n1273 PAD.n1158 0.019716
R50128 PAD.n1330 PAD.n1329 0.019716
R50129 PAD.n1330 PAD.n1157 0.019716
R50130 PAD.n1278 PAD.n1277 0.019716
R50131 PAD.n1278 PAD.n1156 0.019716
R50132 PAD.n1321 PAD.n1320 0.019716
R50133 PAD.n1321 PAD.n1155 0.019716
R50134 PAD.n1283 PAD.n1282 0.019716
R50135 PAD.n1283 PAD.n1154 0.019716
R50136 PAD.n1312 PAD.n1311 0.019716
R50137 PAD.n1312 PAD.n1153 0.019716
R50138 PAD.n1288 PAD.n1287 0.019716
R50139 PAD.n1288 PAD.n1152 0.019716
R50140 PAD.n1303 PAD.n1302 0.019716
R50141 PAD.n1303 PAD.n1151 0.019716
R50142 PAD.n1293 PAD.n1292 0.019716
R50143 PAD.n1293 PAD.n1150 0.019716
R50144 PAD.n1294 PAD.n1149 0.019716
R50145 PAD.n1577 PAD.n1531 0.019716
R50146 PAD.n1578 PAD.n1530 0.019716
R50147 PAD.n9756 PAD.n1529 0.019716
R50148 PAD.n9756 PAD.n9755 0.019716
R50149 PAD.n9758 PAD.n1528 0.019716
R50150 PAD.n9759 PAD.n9758 0.019716
R50151 PAD.n9768 PAD.n1527 0.019716
R50152 PAD.n9768 PAD.n9767 0.019716
R50153 PAD.n9770 PAD.n1526 0.019716
R50154 PAD.n9771 PAD.n9770 0.019716
R50155 PAD.n9780 PAD.n1525 0.019716
R50156 PAD.n9780 PAD.n9779 0.019716
R50157 PAD.n9782 PAD.n1524 0.019716
R50158 PAD.n9783 PAD.n9782 0.019716
R50159 PAD.n9792 PAD.n1523 0.019716
R50160 PAD.n9792 PAD.n9791 0.019716
R50161 PAD.n9794 PAD.n1522 0.019716
R50162 PAD.n9795 PAD.n9794 0.019716
R50163 PAD.n9804 PAD.n1521 0.019716
R50164 PAD.n9804 PAD.n9803 0.019716
R50165 PAD.n9806 PAD.n1520 0.019716
R50166 PAD.n9807 PAD.n9806 0.019716
R50167 PAD.n9816 PAD.n1519 0.019716
R50168 PAD.n9816 PAD.n9815 0.019716
R50169 PAD.n9818 PAD.n1518 0.019716
R50170 PAD.n9819 PAD.n9818 0.019716
R50171 PAD.n9828 PAD.n1517 0.019716
R50172 PAD.n9828 PAD.n9827 0.019716
R50173 PAD.n9830 PAD.n1516 0.019716
R50174 PAD.n9831 PAD.n9830 0.019716
R50175 PAD.n9840 PAD.n1515 0.019716
R50176 PAD.n9840 PAD.n9839 0.019716
R50177 PAD.n9842 PAD.n1514 0.019716
R50178 PAD.n9843 PAD.n9842 0.019716
R50179 PAD.n9852 PAD.n1513 0.019716
R50180 PAD.n9852 PAD.n9851 0.019716
R50181 PAD.n9854 PAD.n1512 0.019716
R50182 PAD.n9855 PAD.n9854 0.019716
R50183 PAD.n9864 PAD.n1511 0.019716
R50184 PAD.n9864 PAD.n9863 0.019716
R50185 PAD.n9866 PAD.n1510 0.019716
R50186 PAD.n9867 PAD.n9866 0.019716
R50187 PAD.n9876 PAD.n1509 0.019716
R50188 PAD.n9876 PAD.n9875 0.019716
R50189 PAD.n9878 PAD.n1508 0.019716
R50190 PAD.n9879 PAD.n9878 0.019716
R50191 PAD.n9888 PAD.n1507 0.019716
R50192 PAD.n9888 PAD.n9887 0.019716
R50193 PAD.n9890 PAD.n1506 0.019716
R50194 PAD.n9891 PAD.n9890 0.019716
R50195 PAD.n9900 PAD.n1505 0.019716
R50196 PAD.n9900 PAD.n9899 0.019716
R50197 PAD.n9902 PAD.n1504 0.019716
R50198 PAD.n9903 PAD.n9902 0.019716
R50199 PAD.n9912 PAD.n1503 0.019716
R50200 PAD.n9912 PAD.n9911 0.019716
R50201 PAD.n9914 PAD.n1502 0.019716
R50202 PAD.n9915 PAD.n9914 0.019716
R50203 PAD.n9924 PAD.n1501 0.019716
R50204 PAD.n9924 PAD.n9923 0.019716
R50205 PAD.n9926 PAD.n1500 0.019716
R50206 PAD.n9927 PAD.n9926 0.019716
R50207 PAD.n9936 PAD.n1499 0.019716
R50208 PAD.n9936 PAD.n9935 0.019716
R50209 PAD.n9938 PAD.n1498 0.019716
R50210 PAD.n9939 PAD.n9938 0.019716
R50211 PAD.n9948 PAD.n1497 0.019716
R50212 PAD.n9948 PAD.n9947 0.019716
R50213 PAD.n9950 PAD.n1496 0.019716
R50214 PAD.n9951 PAD.n9950 0.019716
R50215 PAD.n9960 PAD.n1495 0.019716
R50216 PAD.n9960 PAD.n9959 0.019716
R50217 PAD.n9962 PAD.n1494 0.019716
R50218 PAD.n9963 PAD.n9962 0.019716
R50219 PAD.n9972 PAD.n1493 0.019716
R50220 PAD.n9972 PAD.n9971 0.019716
R50221 PAD.n9974 PAD.n1492 0.019716
R50222 PAD.n9975 PAD.n9974 0.019716
R50223 PAD.n9984 PAD.n1491 0.019716
R50224 PAD.n9984 PAD.n9983 0.019716
R50225 PAD.n9986 PAD.n1490 0.019716
R50226 PAD.n9987 PAD.n9986 0.019716
R50227 PAD.n9997 PAD.n9996 0.019716
R50228 PAD.n1601 PAD.n1599 0.019716
R50229 PAD.n1929 PAD.n1928 0.019716
R50230 PAD.n1925 PAD.n1602 0.019716
R50231 PAD.n1926 PAD.n1925 0.019716
R50232 PAD.n1919 PAD.n1916 0.019716
R50233 PAD.n1919 PAD.n1918 0.019716
R50234 PAD.n1913 PAD.n1607 0.019716
R50235 PAD.n1914 PAD.n1913 0.019716
R50236 PAD.n1907 PAD.n1904 0.019716
R50237 PAD.n1907 PAD.n1906 0.019716
R50238 PAD.n1901 PAD.n1611 0.019716
R50239 PAD.n1902 PAD.n1901 0.019716
R50240 PAD.n1895 PAD.n1892 0.019716
R50241 PAD.n1895 PAD.n1894 0.019716
R50242 PAD.n1889 PAD.n1615 0.019716
R50243 PAD.n1890 PAD.n1889 0.019716
R50244 PAD.n1883 PAD.n1880 0.019716
R50245 PAD.n1883 PAD.n1882 0.019716
R50246 PAD.n1877 PAD.n1619 0.019716
R50247 PAD.n1878 PAD.n1877 0.019716
R50248 PAD.n1871 PAD.n1868 0.019716
R50249 PAD.n1871 PAD.n1870 0.019716
R50250 PAD.n1865 PAD.n1623 0.019716
R50251 PAD.n1866 PAD.n1865 0.019716
R50252 PAD.n1859 PAD.n1856 0.019716
R50253 PAD.n1859 PAD.n1858 0.019716
R50254 PAD.n1853 PAD.n1627 0.019716
R50255 PAD.n1854 PAD.n1853 0.019716
R50256 PAD.n1847 PAD.n1844 0.019716
R50257 PAD.n1847 PAD.n1846 0.019716
R50258 PAD.n1841 PAD.n1631 0.019716
R50259 PAD.n1842 PAD.n1841 0.019716
R50260 PAD.n1835 PAD.n1832 0.019716
R50261 PAD.n1835 PAD.n1834 0.019716
R50262 PAD.n1829 PAD.n1635 0.019716
R50263 PAD.n1830 PAD.n1829 0.019716
R50264 PAD.n1823 PAD.n1820 0.019716
R50265 PAD.n1823 PAD.n1822 0.019716
R50266 PAD.n1817 PAD.n1639 0.019716
R50267 PAD.n1818 PAD.n1817 0.019716
R50268 PAD.n1811 PAD.n1808 0.019716
R50269 PAD.n1811 PAD.n1810 0.019716
R50270 PAD.n1805 PAD.n1643 0.019716
R50271 PAD.n1806 PAD.n1805 0.019716
R50272 PAD.n1799 PAD.n1796 0.019716
R50273 PAD.n1799 PAD.n1798 0.019716
R50274 PAD.n1793 PAD.n1647 0.019716
R50275 PAD.n1794 PAD.n1793 0.019716
R50276 PAD.n1787 PAD.n1784 0.019716
R50277 PAD.n1787 PAD.n1786 0.019716
R50278 PAD.n1781 PAD.n1651 0.019716
R50279 PAD.n1782 PAD.n1781 0.019716
R50280 PAD.n1775 PAD.n1772 0.019716
R50281 PAD.n1775 PAD.n1774 0.019716
R50282 PAD.n1769 PAD.n1655 0.019716
R50283 PAD.n1770 PAD.n1769 0.019716
R50284 PAD.n1763 PAD.n1760 0.019716
R50285 PAD.n1763 PAD.n1762 0.019716
R50286 PAD.n1757 PAD.n1659 0.019716
R50287 PAD.n1758 PAD.n1757 0.019716
R50288 PAD.n1751 PAD.n1748 0.019716
R50289 PAD.n1751 PAD.n1750 0.019716
R50290 PAD.n1745 PAD.n1663 0.019716
R50291 PAD.n1746 PAD.n1745 0.019716
R50292 PAD.n1739 PAD.n1736 0.019716
R50293 PAD.n1739 PAD.n1738 0.019716
R50294 PAD.n1733 PAD.n1667 0.019716
R50295 PAD.n1734 PAD.n1733 0.019716
R50296 PAD.n1727 PAD.n1724 0.019716
R50297 PAD.n1727 PAD.n1726 0.019716
R50298 PAD.n1721 PAD.n1671 0.019716
R50299 PAD.n1722 PAD.n1721 0.019716
R50300 PAD.n1715 PAD.n1712 0.019716
R50301 PAD.n1715 PAD.n1714 0.019716
R50302 PAD.n1709 PAD.n1675 0.019716
R50303 PAD.n1710 PAD.n1709 0.019716
R50304 PAD.n1703 PAD.n1700 0.019716
R50305 PAD.n1703 PAD.n1702 0.019716
R50306 PAD.n1697 PAD.n1679 0.019716
R50307 PAD.n1698 PAD.n1697 0.019716
R50308 PAD.n1691 PAD.n1688 0.019716
R50309 PAD.n1691 PAD.n1690 0.019716
R50310 PAD.n1686 PAD.n1685 0.019716
R50311 PAD.n2029 PAD.n1984 0.019716
R50312 PAD.n2030 PAD.n1983 0.019716
R50313 PAD.n9470 PAD.n1982 0.019716
R50314 PAD.n9470 PAD.n9469 0.019716
R50315 PAD.n9472 PAD.n1981 0.019716
R50316 PAD.n9473 PAD.n9472 0.019716
R50317 PAD.n9482 PAD.n1980 0.019716
R50318 PAD.n9482 PAD.n9481 0.019716
R50319 PAD.n9484 PAD.n1979 0.019716
R50320 PAD.n9485 PAD.n9484 0.019716
R50321 PAD.n9494 PAD.n1978 0.019716
R50322 PAD.n9494 PAD.n9493 0.019716
R50323 PAD.n9496 PAD.n1977 0.019716
R50324 PAD.n9497 PAD.n9496 0.019716
R50325 PAD.n9506 PAD.n1976 0.019716
R50326 PAD.n9506 PAD.n9505 0.019716
R50327 PAD.n9508 PAD.n1975 0.019716
R50328 PAD.n9509 PAD.n9508 0.019716
R50329 PAD.n9518 PAD.n1974 0.019716
R50330 PAD.n9518 PAD.n9517 0.019716
R50331 PAD.n9520 PAD.n1973 0.019716
R50332 PAD.n9521 PAD.n9520 0.019716
R50333 PAD.n9530 PAD.n1972 0.019716
R50334 PAD.n9530 PAD.n9529 0.019716
R50335 PAD.n9532 PAD.n1971 0.019716
R50336 PAD.n9533 PAD.n9532 0.019716
R50337 PAD.n9542 PAD.n1970 0.019716
R50338 PAD.n9542 PAD.n9541 0.019716
R50339 PAD.n9544 PAD.n1969 0.019716
R50340 PAD.n9545 PAD.n9544 0.019716
R50341 PAD.n9554 PAD.n1968 0.019716
R50342 PAD.n9554 PAD.n9553 0.019716
R50343 PAD.n9556 PAD.n1967 0.019716
R50344 PAD.n9557 PAD.n9556 0.019716
R50345 PAD.n9566 PAD.n1966 0.019716
R50346 PAD.n9566 PAD.n9565 0.019716
R50347 PAD.n9568 PAD.n1965 0.019716
R50348 PAD.n9569 PAD.n9568 0.019716
R50349 PAD.n9578 PAD.n1964 0.019716
R50350 PAD.n9578 PAD.n9577 0.019716
R50351 PAD.n9580 PAD.n1963 0.019716
R50352 PAD.n9581 PAD.n9580 0.019716
R50353 PAD.n9590 PAD.n1962 0.019716
R50354 PAD.n9590 PAD.n9589 0.019716
R50355 PAD.n9592 PAD.n1961 0.019716
R50356 PAD.n9593 PAD.n9592 0.019716
R50357 PAD.n9602 PAD.n1960 0.019716
R50358 PAD.n9602 PAD.n9601 0.019716
R50359 PAD.n9604 PAD.n1959 0.019716
R50360 PAD.n9605 PAD.n9604 0.019716
R50361 PAD.n9614 PAD.n1958 0.019716
R50362 PAD.n9614 PAD.n9613 0.019716
R50363 PAD.n9616 PAD.n1957 0.019716
R50364 PAD.n9617 PAD.n9616 0.019716
R50365 PAD.n9626 PAD.n1956 0.019716
R50366 PAD.n9626 PAD.n9625 0.019716
R50367 PAD.n9628 PAD.n1955 0.019716
R50368 PAD.n9629 PAD.n9628 0.019716
R50369 PAD.n9638 PAD.n1954 0.019716
R50370 PAD.n9638 PAD.n9637 0.019716
R50371 PAD.n9640 PAD.n1953 0.019716
R50372 PAD.n9641 PAD.n9640 0.019716
R50373 PAD.n9650 PAD.n1952 0.019716
R50374 PAD.n9650 PAD.n9649 0.019716
R50375 PAD.n9652 PAD.n1951 0.019716
R50376 PAD.n9653 PAD.n9652 0.019716
R50377 PAD.n9662 PAD.n1950 0.019716
R50378 PAD.n9662 PAD.n9661 0.019716
R50379 PAD.n9664 PAD.n1949 0.019716
R50380 PAD.n9665 PAD.n9664 0.019716
R50381 PAD.n9674 PAD.n1948 0.019716
R50382 PAD.n9674 PAD.n9673 0.019716
R50383 PAD.n9676 PAD.n1947 0.019716
R50384 PAD.n9677 PAD.n9676 0.019716
R50385 PAD.n9686 PAD.n1946 0.019716
R50386 PAD.n9686 PAD.n9685 0.019716
R50387 PAD.n9688 PAD.n1945 0.019716
R50388 PAD.n9689 PAD.n9688 0.019716
R50389 PAD.n9698 PAD.n1944 0.019716
R50390 PAD.n9698 PAD.n9697 0.019716
R50391 PAD.n9700 PAD.n1943 0.019716
R50392 PAD.n9701 PAD.n9700 0.019716
R50393 PAD.n9711 PAD.n9710 0.019716
R50394 PAD.n2132 PAD.n2088 0.019716
R50395 PAD.n2133 PAD.n2087 0.019716
R50396 PAD.n9204 PAD.n2086 0.019716
R50397 PAD.n9204 PAD.n9203 0.019716
R50398 PAD.n9206 PAD.n2085 0.019716
R50399 PAD.n9207 PAD.n9206 0.019716
R50400 PAD.n9216 PAD.n2084 0.019716
R50401 PAD.n9216 PAD.n9215 0.019716
R50402 PAD.n9218 PAD.n2083 0.019716
R50403 PAD.n9219 PAD.n9218 0.019716
R50404 PAD.n9228 PAD.n2082 0.019716
R50405 PAD.n9228 PAD.n9227 0.019716
R50406 PAD.n9230 PAD.n2081 0.019716
R50407 PAD.n9231 PAD.n9230 0.019716
R50408 PAD.n9240 PAD.n2080 0.019716
R50409 PAD.n9240 PAD.n9239 0.019716
R50410 PAD.n9242 PAD.n2079 0.019716
R50411 PAD.n9243 PAD.n9242 0.019716
R50412 PAD.n9252 PAD.n2078 0.019716
R50413 PAD.n9252 PAD.n9251 0.019716
R50414 PAD.n9254 PAD.n2077 0.019716
R50415 PAD.n9255 PAD.n9254 0.019716
R50416 PAD.n9264 PAD.n2076 0.019716
R50417 PAD.n9264 PAD.n9263 0.019716
R50418 PAD.n9266 PAD.n2075 0.019716
R50419 PAD.n9267 PAD.n9266 0.019716
R50420 PAD.n9276 PAD.n2074 0.019716
R50421 PAD.n9276 PAD.n9275 0.019716
R50422 PAD.n9278 PAD.n2073 0.019716
R50423 PAD.n9279 PAD.n9278 0.019716
R50424 PAD.n9288 PAD.n2072 0.019716
R50425 PAD.n9288 PAD.n9287 0.019716
R50426 PAD.n9290 PAD.n2071 0.019716
R50427 PAD.n9291 PAD.n9290 0.019716
R50428 PAD.n9300 PAD.n2070 0.019716
R50429 PAD.n9300 PAD.n9299 0.019716
R50430 PAD.n9302 PAD.n2069 0.019716
R50431 PAD.n9303 PAD.n9302 0.019716
R50432 PAD.n9312 PAD.n2068 0.019716
R50433 PAD.n9312 PAD.n9311 0.019716
R50434 PAD.n9314 PAD.n2067 0.019716
R50435 PAD.n9315 PAD.n9314 0.019716
R50436 PAD.n9324 PAD.n2066 0.019716
R50437 PAD.n9324 PAD.n9323 0.019716
R50438 PAD.n9326 PAD.n2065 0.019716
R50439 PAD.n9327 PAD.n9326 0.019716
R50440 PAD.n9336 PAD.n2064 0.019716
R50441 PAD.n9336 PAD.n9335 0.019716
R50442 PAD.n9338 PAD.n2063 0.019716
R50443 PAD.n9339 PAD.n9338 0.019716
R50444 PAD.n9348 PAD.n2062 0.019716
R50445 PAD.n9348 PAD.n9347 0.019716
R50446 PAD.n9350 PAD.n2061 0.019716
R50447 PAD.n9351 PAD.n9350 0.019716
R50448 PAD.n9360 PAD.n2060 0.019716
R50449 PAD.n9360 PAD.n9359 0.019716
R50450 PAD.n9362 PAD.n2059 0.019716
R50451 PAD.n9363 PAD.n9362 0.019716
R50452 PAD.n9372 PAD.n2058 0.019716
R50453 PAD.n9372 PAD.n9371 0.019716
R50454 PAD.n9374 PAD.n2057 0.019716
R50455 PAD.n9375 PAD.n9374 0.019716
R50456 PAD.n9384 PAD.n2056 0.019716
R50457 PAD.n9384 PAD.n9383 0.019716
R50458 PAD.n9386 PAD.n2055 0.019716
R50459 PAD.n9387 PAD.n9386 0.019716
R50460 PAD.n9396 PAD.n2054 0.019716
R50461 PAD.n9396 PAD.n9395 0.019716
R50462 PAD.n9398 PAD.n2053 0.019716
R50463 PAD.n9399 PAD.n9398 0.019716
R50464 PAD.n9408 PAD.n2052 0.019716
R50465 PAD.n9408 PAD.n9407 0.019716
R50466 PAD.n9410 PAD.n2051 0.019716
R50467 PAD.n9411 PAD.n9410 0.019716
R50468 PAD.n9420 PAD.n2050 0.019716
R50469 PAD.n9420 PAD.n9419 0.019716
R50470 PAD.n9422 PAD.n2049 0.019716
R50471 PAD.n9423 PAD.n9422 0.019716
R50472 PAD.n9432 PAD.n2048 0.019716
R50473 PAD.n9432 PAD.n9431 0.019716
R50474 PAD.n9434 PAD.n2047 0.019716
R50475 PAD.n9435 PAD.n9434 0.019716
R50476 PAD.n9444 PAD.n9443 0.019716
R50477 PAD.n2153 PAD.n2151 0.019716
R50478 PAD.n2480 PAD.n2479 0.019716
R50479 PAD.n2476 PAD.n2154 0.019716
R50480 PAD.n2477 PAD.n2476 0.019716
R50481 PAD.n2470 PAD.n2467 0.019716
R50482 PAD.n2470 PAD.n2469 0.019716
R50483 PAD.n2464 PAD.n2159 0.019716
R50484 PAD.n2465 PAD.n2464 0.019716
R50485 PAD.n2458 PAD.n2455 0.019716
R50486 PAD.n2458 PAD.n2457 0.019716
R50487 PAD.n2452 PAD.n2163 0.019716
R50488 PAD.n2453 PAD.n2452 0.019716
R50489 PAD.n2446 PAD.n2443 0.019716
R50490 PAD.n2446 PAD.n2445 0.019716
R50491 PAD.n2440 PAD.n2167 0.019716
R50492 PAD.n2441 PAD.n2440 0.019716
R50493 PAD.n2434 PAD.n2431 0.019716
R50494 PAD.n2434 PAD.n2433 0.019716
R50495 PAD.n2428 PAD.n2171 0.019716
R50496 PAD.n2429 PAD.n2428 0.019716
R50497 PAD.n2422 PAD.n2419 0.019716
R50498 PAD.n2422 PAD.n2421 0.019716
R50499 PAD.n2416 PAD.n2175 0.019716
R50500 PAD.n2417 PAD.n2416 0.019716
R50501 PAD.n2410 PAD.n2407 0.019716
R50502 PAD.n2410 PAD.n2409 0.019716
R50503 PAD.n2404 PAD.n2179 0.019716
R50504 PAD.n2405 PAD.n2404 0.019716
R50505 PAD.n2398 PAD.n2395 0.019716
R50506 PAD.n2398 PAD.n2397 0.019716
R50507 PAD.n2392 PAD.n2183 0.019716
R50508 PAD.n2393 PAD.n2392 0.019716
R50509 PAD.n2386 PAD.n2383 0.019716
R50510 PAD.n2386 PAD.n2385 0.019716
R50511 PAD.n2380 PAD.n2187 0.019716
R50512 PAD.n2381 PAD.n2380 0.019716
R50513 PAD.n2374 PAD.n2371 0.019716
R50514 PAD.n2374 PAD.n2373 0.019716
R50515 PAD.n2368 PAD.n2191 0.019716
R50516 PAD.n2369 PAD.n2368 0.019716
R50517 PAD.n2362 PAD.n2359 0.019716
R50518 PAD.n2362 PAD.n2361 0.019716
R50519 PAD.n2356 PAD.n2195 0.019716
R50520 PAD.n2357 PAD.n2356 0.019716
R50521 PAD.n2350 PAD.n2347 0.019716
R50522 PAD.n2350 PAD.n2349 0.019716
R50523 PAD.n2344 PAD.n2199 0.019716
R50524 PAD.n2345 PAD.n2344 0.019716
R50525 PAD.n2338 PAD.n2335 0.019716
R50526 PAD.n2338 PAD.n2337 0.019716
R50527 PAD.n2332 PAD.n2203 0.019716
R50528 PAD.n2333 PAD.n2332 0.019716
R50529 PAD.n2326 PAD.n2323 0.019716
R50530 PAD.n2326 PAD.n2325 0.019716
R50531 PAD.n2320 PAD.n2207 0.019716
R50532 PAD.n2321 PAD.n2320 0.019716
R50533 PAD.n2314 PAD.n2311 0.019716
R50534 PAD.n2314 PAD.n2313 0.019716
R50535 PAD.n2308 PAD.n2211 0.019716
R50536 PAD.n2309 PAD.n2308 0.019716
R50537 PAD.n2302 PAD.n2299 0.019716
R50538 PAD.n2302 PAD.n2301 0.019716
R50539 PAD.n2296 PAD.n2215 0.019716
R50540 PAD.n2297 PAD.n2296 0.019716
R50541 PAD.n2290 PAD.n2287 0.019716
R50542 PAD.n2290 PAD.n2289 0.019716
R50543 PAD.n2284 PAD.n2219 0.019716
R50544 PAD.n2285 PAD.n2284 0.019716
R50545 PAD.n2278 PAD.n2275 0.019716
R50546 PAD.n2278 PAD.n2277 0.019716
R50547 PAD.n2272 PAD.n2223 0.019716
R50548 PAD.n2273 PAD.n2272 0.019716
R50549 PAD.n2266 PAD.n2263 0.019716
R50550 PAD.n2266 PAD.n2265 0.019716
R50551 PAD.n2260 PAD.n2227 0.019716
R50552 PAD.n2261 PAD.n2260 0.019716
R50553 PAD.n2254 PAD.n2251 0.019716
R50554 PAD.n2254 PAD.n2253 0.019716
R50555 PAD.n2248 PAD.n2231 0.019716
R50556 PAD.n2249 PAD.n2248 0.019716
R50557 PAD.n2242 PAD.n2239 0.019716
R50558 PAD.n2242 PAD.n2241 0.019716
R50559 PAD.n2237 PAD.n2236 0.019716
R50560 PAD.n2500 PAD.n2498 0.019716
R50561 PAD.n2827 PAD.n2826 0.019716
R50562 PAD.n2823 PAD.n2501 0.019716
R50563 PAD.n2824 PAD.n2823 0.019716
R50564 PAD.n2817 PAD.n2814 0.019716
R50565 PAD.n2817 PAD.n2816 0.019716
R50566 PAD.n2811 PAD.n2506 0.019716
R50567 PAD.n2812 PAD.n2811 0.019716
R50568 PAD.n2805 PAD.n2802 0.019716
R50569 PAD.n2805 PAD.n2804 0.019716
R50570 PAD.n2799 PAD.n2510 0.019716
R50571 PAD.n2800 PAD.n2799 0.019716
R50572 PAD.n2793 PAD.n2790 0.019716
R50573 PAD.n2793 PAD.n2792 0.019716
R50574 PAD.n2787 PAD.n2514 0.019716
R50575 PAD.n2788 PAD.n2787 0.019716
R50576 PAD.n2781 PAD.n2778 0.019716
R50577 PAD.n2781 PAD.n2780 0.019716
R50578 PAD.n2775 PAD.n2518 0.019716
R50579 PAD.n2776 PAD.n2775 0.019716
R50580 PAD.n2769 PAD.n2766 0.019716
R50581 PAD.n2769 PAD.n2768 0.019716
R50582 PAD.n2763 PAD.n2522 0.019716
R50583 PAD.n2764 PAD.n2763 0.019716
R50584 PAD.n2757 PAD.n2754 0.019716
R50585 PAD.n2757 PAD.n2756 0.019716
R50586 PAD.n2751 PAD.n2526 0.019716
R50587 PAD.n2752 PAD.n2751 0.019716
R50588 PAD.n2745 PAD.n2742 0.019716
R50589 PAD.n2745 PAD.n2744 0.019716
R50590 PAD.n2739 PAD.n2530 0.019716
R50591 PAD.n2740 PAD.n2739 0.019716
R50592 PAD.n2733 PAD.n2730 0.019716
R50593 PAD.n2733 PAD.n2732 0.019716
R50594 PAD.n2727 PAD.n2534 0.019716
R50595 PAD.n2728 PAD.n2727 0.019716
R50596 PAD.n2721 PAD.n2718 0.019716
R50597 PAD.n2721 PAD.n2720 0.019716
R50598 PAD.n2715 PAD.n2538 0.019716
R50599 PAD.n2716 PAD.n2715 0.019716
R50600 PAD.n2709 PAD.n2706 0.019716
R50601 PAD.n2709 PAD.n2708 0.019716
R50602 PAD.n2703 PAD.n2542 0.019716
R50603 PAD.n2704 PAD.n2703 0.019716
R50604 PAD.n2697 PAD.n2694 0.019716
R50605 PAD.n2697 PAD.n2696 0.019716
R50606 PAD.n2691 PAD.n2546 0.019716
R50607 PAD.n2692 PAD.n2691 0.019716
R50608 PAD.n2685 PAD.n2682 0.019716
R50609 PAD.n2685 PAD.n2684 0.019716
R50610 PAD.n2679 PAD.n2550 0.019716
R50611 PAD.n2680 PAD.n2679 0.019716
R50612 PAD.n2673 PAD.n2670 0.019716
R50613 PAD.n2673 PAD.n2672 0.019716
R50614 PAD.n2667 PAD.n2554 0.019716
R50615 PAD.n2668 PAD.n2667 0.019716
R50616 PAD.n2661 PAD.n2658 0.019716
R50617 PAD.n2661 PAD.n2660 0.019716
R50618 PAD.n2655 PAD.n2558 0.019716
R50619 PAD.n2656 PAD.n2655 0.019716
R50620 PAD.n2649 PAD.n2646 0.019716
R50621 PAD.n2649 PAD.n2648 0.019716
R50622 PAD.n2643 PAD.n2562 0.019716
R50623 PAD.n2644 PAD.n2643 0.019716
R50624 PAD.n2637 PAD.n2634 0.019716
R50625 PAD.n2637 PAD.n2636 0.019716
R50626 PAD.n2631 PAD.n2566 0.019716
R50627 PAD.n2632 PAD.n2631 0.019716
R50628 PAD.n2625 PAD.n2622 0.019716
R50629 PAD.n2625 PAD.n2624 0.019716
R50630 PAD.n2619 PAD.n2570 0.019716
R50631 PAD.n2620 PAD.n2619 0.019716
R50632 PAD.n2613 PAD.n2610 0.019716
R50633 PAD.n2613 PAD.n2612 0.019716
R50634 PAD.n2607 PAD.n2574 0.019716
R50635 PAD.n2608 PAD.n2607 0.019716
R50636 PAD.n2601 PAD.n2598 0.019716
R50637 PAD.n2601 PAD.n2600 0.019716
R50638 PAD.n2595 PAD.n2578 0.019716
R50639 PAD.n2596 PAD.n2595 0.019716
R50640 PAD.n2589 PAD.n2586 0.019716
R50641 PAD.n2589 PAD.n2588 0.019716
R50642 PAD.n2584 PAD.n2583 0.019716
R50643 PAD.n9116 PAD.n2876 0.019716
R50644 PAD.n9117 PAD.n2875 0.019716
R50645 PAD.n8839 PAD.n2874 0.019716
R50646 PAD.n8840 PAD.n8839 0.019716
R50647 PAD.n9108 PAD.n2873 0.019716
R50648 PAD.n9109 PAD.n9108 0.019716
R50649 PAD.n8844 PAD.n2872 0.019716
R50650 PAD.n8845 PAD.n8844 0.019716
R50651 PAD.n9099 PAD.n2871 0.019716
R50652 PAD.n9100 PAD.n9099 0.019716
R50653 PAD.n8849 PAD.n2870 0.019716
R50654 PAD.n8850 PAD.n8849 0.019716
R50655 PAD.n9090 PAD.n2869 0.019716
R50656 PAD.n9091 PAD.n9090 0.019716
R50657 PAD.n8854 PAD.n2868 0.019716
R50658 PAD.n8855 PAD.n8854 0.019716
R50659 PAD.n9081 PAD.n2867 0.019716
R50660 PAD.n9082 PAD.n9081 0.019716
R50661 PAD.n8859 PAD.n2866 0.019716
R50662 PAD.n8860 PAD.n8859 0.019716
R50663 PAD.n9072 PAD.n2865 0.019716
R50664 PAD.n9073 PAD.n9072 0.019716
R50665 PAD.n8864 PAD.n2864 0.019716
R50666 PAD.n8865 PAD.n8864 0.019716
R50667 PAD.n9063 PAD.n2863 0.019716
R50668 PAD.n9064 PAD.n9063 0.019716
R50669 PAD.n8869 PAD.n2862 0.019716
R50670 PAD.n8870 PAD.n8869 0.019716
R50671 PAD.n9054 PAD.n2861 0.019716
R50672 PAD.n9055 PAD.n9054 0.019716
R50673 PAD.n8874 PAD.n2860 0.019716
R50674 PAD.n8875 PAD.n8874 0.019716
R50675 PAD.n9045 PAD.n2859 0.019716
R50676 PAD.n9046 PAD.n9045 0.019716
R50677 PAD.n8879 PAD.n2858 0.019716
R50678 PAD.n8880 PAD.n8879 0.019716
R50679 PAD.n9036 PAD.n2857 0.019716
R50680 PAD.n9037 PAD.n9036 0.019716
R50681 PAD.n8884 PAD.n2856 0.019716
R50682 PAD.n8885 PAD.n8884 0.019716
R50683 PAD.n9027 PAD.n2855 0.019716
R50684 PAD.n9028 PAD.n9027 0.019716
R50685 PAD.n8889 PAD.n2854 0.019716
R50686 PAD.n8890 PAD.n8889 0.019716
R50687 PAD.n9018 PAD.n2853 0.019716
R50688 PAD.n9019 PAD.n9018 0.019716
R50689 PAD.n8894 PAD.n2852 0.019716
R50690 PAD.n8895 PAD.n8894 0.019716
R50691 PAD.n9009 PAD.n2851 0.019716
R50692 PAD.n9010 PAD.n9009 0.019716
R50693 PAD.n8899 PAD.n2850 0.019716
R50694 PAD.n8900 PAD.n8899 0.019716
R50695 PAD.n9000 PAD.n2849 0.019716
R50696 PAD.n9001 PAD.n9000 0.019716
R50697 PAD.n8904 PAD.n2848 0.019716
R50698 PAD.n8905 PAD.n8904 0.019716
R50699 PAD.n8991 PAD.n2847 0.019716
R50700 PAD.n8992 PAD.n8991 0.019716
R50701 PAD.n8909 PAD.n2846 0.019716
R50702 PAD.n8910 PAD.n8909 0.019716
R50703 PAD.n8982 PAD.n2845 0.019716
R50704 PAD.n8983 PAD.n8982 0.019716
R50705 PAD.n8914 PAD.n2844 0.019716
R50706 PAD.n8915 PAD.n8914 0.019716
R50707 PAD.n8973 PAD.n2843 0.019716
R50708 PAD.n8974 PAD.n8973 0.019716
R50709 PAD.n8919 PAD.n2842 0.019716
R50710 PAD.n8920 PAD.n8919 0.019716
R50711 PAD.n8964 PAD.n2841 0.019716
R50712 PAD.n8965 PAD.n8964 0.019716
R50713 PAD.n8924 PAD.n2840 0.019716
R50714 PAD.n8925 PAD.n8924 0.019716
R50715 PAD.n8955 PAD.n2839 0.019716
R50716 PAD.n8956 PAD.n8955 0.019716
R50717 PAD.n8929 PAD.n2838 0.019716
R50718 PAD.n8930 PAD.n8929 0.019716
R50719 PAD.n8946 PAD.n2837 0.019716
R50720 PAD.n8947 PAD.n8946 0.019716
R50721 PAD.n8934 PAD.n2836 0.019716
R50722 PAD.n8935 PAD.n8934 0.019716
R50723 PAD.n8937 PAD.n2835 0.019716
R50724 PAD.n8938 PAD.n8937 0.019716
R50725 PAD.n9139 PAD.n9138 0.019716
R50726 PAD.n8820 PAD.n8819 0.019716
R50727 PAD.n8812 PAD.n8528 0.019716
R50728 PAD.n8810 PAD.n8809 0.019716
R50729 PAD.n8810 PAD.n2945 0.019716
R50730 PAD.n8801 PAD.n8800 0.019716
R50731 PAD.n8800 PAD.n2944 0.019716
R50732 PAD.n8798 PAD.n8797 0.019716
R50733 PAD.n8798 PAD.n2943 0.019716
R50734 PAD.n8789 PAD.n8788 0.019716
R50735 PAD.n8788 PAD.n2942 0.019716
R50736 PAD.n8786 PAD.n8785 0.019716
R50737 PAD.n8786 PAD.n2941 0.019716
R50738 PAD.n8777 PAD.n8776 0.019716
R50739 PAD.n8776 PAD.n2940 0.019716
R50740 PAD.n8774 PAD.n8773 0.019716
R50741 PAD.n8774 PAD.n2939 0.019716
R50742 PAD.n8765 PAD.n8764 0.019716
R50743 PAD.n8764 PAD.n2938 0.019716
R50744 PAD.n8762 PAD.n8761 0.019716
R50745 PAD.n8762 PAD.n2937 0.019716
R50746 PAD.n8753 PAD.n8752 0.019716
R50747 PAD.n8752 PAD.n2936 0.019716
R50748 PAD.n8750 PAD.n8749 0.019716
R50749 PAD.n8750 PAD.n2935 0.019716
R50750 PAD.n8741 PAD.n8740 0.019716
R50751 PAD.n8740 PAD.n2934 0.019716
R50752 PAD.n8738 PAD.n8737 0.019716
R50753 PAD.n8738 PAD.n2933 0.019716
R50754 PAD.n8729 PAD.n8728 0.019716
R50755 PAD.n8728 PAD.n2932 0.019716
R50756 PAD.n8726 PAD.n8725 0.019716
R50757 PAD.n8726 PAD.n2931 0.019716
R50758 PAD.n8717 PAD.n8716 0.019716
R50759 PAD.n8716 PAD.n2930 0.019716
R50760 PAD.n8714 PAD.n8713 0.019716
R50761 PAD.n8714 PAD.n2929 0.019716
R50762 PAD.n8705 PAD.n8704 0.019716
R50763 PAD.n8704 PAD.n2928 0.019716
R50764 PAD.n8702 PAD.n8701 0.019716
R50765 PAD.n8702 PAD.n2927 0.019716
R50766 PAD.n8693 PAD.n8692 0.019716
R50767 PAD.n8692 PAD.n2926 0.019716
R50768 PAD.n8690 PAD.n8689 0.019716
R50769 PAD.n8690 PAD.n2925 0.019716
R50770 PAD.n8681 PAD.n8680 0.019716
R50771 PAD.n8680 PAD.n2924 0.019716
R50772 PAD.n8678 PAD.n8677 0.019716
R50773 PAD.n8678 PAD.n2923 0.019716
R50774 PAD.n8669 PAD.n8668 0.019716
R50775 PAD.n8668 PAD.n2922 0.019716
R50776 PAD.n8666 PAD.n8665 0.019716
R50777 PAD.n8666 PAD.n2921 0.019716
R50778 PAD.n8657 PAD.n8656 0.019716
R50779 PAD.n8656 PAD.n2920 0.019716
R50780 PAD.n8654 PAD.n8653 0.019716
R50781 PAD.n8654 PAD.n2919 0.019716
R50782 PAD.n8645 PAD.n8644 0.019716
R50783 PAD.n8644 PAD.n2918 0.019716
R50784 PAD.n8642 PAD.n8641 0.019716
R50785 PAD.n8642 PAD.n2917 0.019716
R50786 PAD.n8633 PAD.n8632 0.019716
R50787 PAD.n8632 PAD.n2916 0.019716
R50788 PAD.n8630 PAD.n8629 0.019716
R50789 PAD.n8630 PAD.n2915 0.019716
R50790 PAD.n8621 PAD.n8620 0.019716
R50791 PAD.n8620 PAD.n2914 0.019716
R50792 PAD.n8618 PAD.n8617 0.019716
R50793 PAD.n8618 PAD.n2913 0.019716
R50794 PAD.n8609 PAD.n8608 0.019716
R50795 PAD.n8608 PAD.n2912 0.019716
R50796 PAD.n8606 PAD.n8605 0.019716
R50797 PAD.n8606 PAD.n2911 0.019716
R50798 PAD.n8597 PAD.n8596 0.019716
R50799 PAD.n8596 PAD.n2910 0.019716
R50800 PAD.n8594 PAD.n8593 0.019716
R50801 PAD.n8594 PAD.n2909 0.019716
R50802 PAD.n8585 PAD.n8584 0.019716
R50803 PAD.n8584 PAD.n2908 0.019716
R50804 PAD.n8582 PAD.n8581 0.019716
R50805 PAD.n8582 PAD.n2907 0.019716
R50806 PAD.n8573 PAD.n8572 0.019716
R50807 PAD.n8572 PAD.n2906 0.019716
R50808 PAD.n8570 PAD.n2905 0.019716
R50809 PAD.n3038 PAD.n2994 0.019716
R50810 PAD.n3039 PAD.n2993 0.019716
R50811 PAD.n3048 PAD.n2992 0.019716
R50812 PAD.n3048 PAD.n3047 0.019716
R50813 PAD.n3050 PAD.n2991 0.019716
R50814 PAD.n3051 PAD.n3050 0.019716
R50815 PAD.n3060 PAD.n2990 0.019716
R50816 PAD.n3060 PAD.n3059 0.019716
R50817 PAD.n3062 PAD.n2989 0.019716
R50818 PAD.n3063 PAD.n3062 0.019716
R50819 PAD.n3072 PAD.n2988 0.019716
R50820 PAD.n3072 PAD.n3071 0.019716
R50821 PAD.n3074 PAD.n2987 0.019716
R50822 PAD.n3075 PAD.n3074 0.019716
R50823 PAD.n3084 PAD.n2986 0.019716
R50824 PAD.n3084 PAD.n3083 0.019716
R50825 PAD.n3086 PAD.n2985 0.019716
R50826 PAD.n3087 PAD.n3086 0.019716
R50827 PAD.n3096 PAD.n2984 0.019716
R50828 PAD.n3096 PAD.n3095 0.019716
R50829 PAD.n3098 PAD.n2983 0.019716
R50830 PAD.n3099 PAD.n3098 0.019716
R50831 PAD.n3108 PAD.n2982 0.019716
R50832 PAD.n3108 PAD.n3107 0.019716
R50833 PAD.n3110 PAD.n2981 0.019716
R50834 PAD.n3111 PAD.n3110 0.019716
R50835 PAD.n3120 PAD.n2980 0.019716
R50836 PAD.n3120 PAD.n3119 0.019716
R50837 PAD.n3122 PAD.n2979 0.019716
R50838 PAD.n3123 PAD.n3122 0.019716
R50839 PAD.n3132 PAD.n2978 0.019716
R50840 PAD.n3132 PAD.n3131 0.019716
R50841 PAD.n3134 PAD.n2977 0.019716
R50842 PAD.n3135 PAD.n3134 0.019716
R50843 PAD.n3144 PAD.n2976 0.019716
R50844 PAD.n3144 PAD.n3143 0.019716
R50845 PAD.n3146 PAD.n2975 0.019716
R50846 PAD.n3147 PAD.n3146 0.019716
R50847 PAD.n3156 PAD.n2974 0.019716
R50848 PAD.n3156 PAD.n3155 0.019716
R50849 PAD.n3158 PAD.n2973 0.019716
R50850 PAD.n3159 PAD.n3158 0.019716
R50851 PAD.n3168 PAD.n2972 0.019716
R50852 PAD.n3168 PAD.n3167 0.019716
R50853 PAD.n3170 PAD.n2971 0.019716
R50854 PAD.n3171 PAD.n3170 0.019716
R50855 PAD.n3180 PAD.n2970 0.019716
R50856 PAD.n3180 PAD.n3179 0.019716
R50857 PAD.n3182 PAD.n2969 0.019716
R50858 PAD.n3183 PAD.n3182 0.019716
R50859 PAD.n3192 PAD.n2968 0.019716
R50860 PAD.n3192 PAD.n3191 0.019716
R50861 PAD.n3194 PAD.n2967 0.019716
R50862 PAD.n3195 PAD.n3194 0.019716
R50863 PAD.n3204 PAD.n2966 0.019716
R50864 PAD.n3204 PAD.n3203 0.019716
R50865 PAD.n3206 PAD.n2965 0.019716
R50866 PAD.n3207 PAD.n3206 0.019716
R50867 PAD.n3216 PAD.n2964 0.019716
R50868 PAD.n3216 PAD.n3215 0.019716
R50869 PAD.n3218 PAD.n2963 0.019716
R50870 PAD.n3219 PAD.n3218 0.019716
R50871 PAD.n3228 PAD.n2962 0.019716
R50872 PAD.n3228 PAD.n3227 0.019716
R50873 PAD.n3230 PAD.n2961 0.019716
R50874 PAD.n3231 PAD.n3230 0.019716
R50875 PAD.n3240 PAD.n2960 0.019716
R50876 PAD.n3240 PAD.n3239 0.019716
R50877 PAD.n3242 PAD.n2959 0.019716
R50878 PAD.n3243 PAD.n3242 0.019716
R50879 PAD.n3252 PAD.n2958 0.019716
R50880 PAD.n3252 PAD.n3251 0.019716
R50881 PAD.n3254 PAD.n2957 0.019716
R50882 PAD.n3255 PAD.n3254 0.019716
R50883 PAD.n3264 PAD.n2956 0.019716
R50884 PAD.n3264 PAD.n3263 0.019716
R50885 PAD.n3266 PAD.n2955 0.019716
R50886 PAD.n3267 PAD.n3266 0.019716
R50887 PAD.n3276 PAD.n2954 0.019716
R50888 PAD.n3276 PAD.n3275 0.019716
R50889 PAD.n3278 PAD.n2953 0.019716
R50890 PAD.n3279 PAD.n3278 0.019716
R50891 PAD.n8516 PAD.n8515 0.019716
R50892 PAD.n3383 PAD.n3338 0.019716
R50893 PAD.n3384 PAD.n3337 0.019716
R50894 PAD.n3393 PAD.n3336 0.019716
R50895 PAD.n3393 PAD.n3392 0.019716
R50896 PAD.n3395 PAD.n3335 0.019716
R50897 PAD.n3396 PAD.n3395 0.019716
R50898 PAD.n3405 PAD.n3334 0.019716
R50899 PAD.n3405 PAD.n3404 0.019716
R50900 PAD.n3407 PAD.n3333 0.019716
R50901 PAD.n3408 PAD.n3407 0.019716
R50902 PAD.n3417 PAD.n3332 0.019716
R50903 PAD.n3417 PAD.n3416 0.019716
R50904 PAD.n3419 PAD.n3331 0.019716
R50905 PAD.n3420 PAD.n3419 0.019716
R50906 PAD.n3429 PAD.n3330 0.019716
R50907 PAD.n3429 PAD.n3428 0.019716
R50908 PAD.n3431 PAD.n3329 0.019716
R50909 PAD.n3432 PAD.n3431 0.019716
R50910 PAD.n3441 PAD.n3328 0.019716
R50911 PAD.n3441 PAD.n3440 0.019716
R50912 PAD.n3443 PAD.n3327 0.019716
R50913 PAD.n3444 PAD.n3443 0.019716
R50914 PAD.n3453 PAD.n3326 0.019716
R50915 PAD.n3453 PAD.n3452 0.019716
R50916 PAD.n3455 PAD.n3325 0.019716
R50917 PAD.n3456 PAD.n3455 0.019716
R50918 PAD.n3465 PAD.n3324 0.019716
R50919 PAD.n3465 PAD.n3464 0.019716
R50920 PAD.n3467 PAD.n3323 0.019716
R50921 PAD.n3468 PAD.n3467 0.019716
R50922 PAD.n3477 PAD.n3322 0.019716
R50923 PAD.n3477 PAD.n3476 0.019716
R50924 PAD.n3479 PAD.n3321 0.019716
R50925 PAD.n3480 PAD.n3479 0.019716
R50926 PAD.n3489 PAD.n3320 0.019716
R50927 PAD.n3489 PAD.n3488 0.019716
R50928 PAD.n3491 PAD.n3319 0.019716
R50929 PAD.n3492 PAD.n3491 0.019716
R50930 PAD.n3501 PAD.n3318 0.019716
R50931 PAD.n3501 PAD.n3500 0.019716
R50932 PAD.n3503 PAD.n3317 0.019716
R50933 PAD.n3504 PAD.n3503 0.019716
R50934 PAD.n3513 PAD.n3316 0.019716
R50935 PAD.n3513 PAD.n3512 0.019716
R50936 PAD.n3515 PAD.n3315 0.019716
R50937 PAD.n3516 PAD.n3515 0.019716
R50938 PAD.n3525 PAD.n3314 0.019716
R50939 PAD.n3525 PAD.n3524 0.019716
R50940 PAD.n3527 PAD.n3313 0.019716
R50941 PAD.n3528 PAD.n3527 0.019716
R50942 PAD.n3537 PAD.n3312 0.019716
R50943 PAD.n3537 PAD.n3536 0.019716
R50944 PAD.n3539 PAD.n3311 0.019716
R50945 PAD.n3540 PAD.n3539 0.019716
R50946 PAD.n3549 PAD.n3310 0.019716
R50947 PAD.n3549 PAD.n3548 0.019716
R50948 PAD.n3551 PAD.n3309 0.019716
R50949 PAD.n3552 PAD.n3551 0.019716
R50950 PAD.n3561 PAD.n3308 0.019716
R50951 PAD.n3561 PAD.n3560 0.019716
R50952 PAD.n3563 PAD.n3307 0.019716
R50953 PAD.n3564 PAD.n3563 0.019716
R50954 PAD.n3573 PAD.n3306 0.019716
R50955 PAD.n3573 PAD.n3572 0.019716
R50956 PAD.n3575 PAD.n3305 0.019716
R50957 PAD.n3576 PAD.n3575 0.019716
R50958 PAD.n3585 PAD.n3304 0.019716
R50959 PAD.n3585 PAD.n3584 0.019716
R50960 PAD.n3587 PAD.n3303 0.019716
R50961 PAD.n3588 PAD.n3587 0.019716
R50962 PAD.n3597 PAD.n3302 0.019716
R50963 PAD.n3597 PAD.n3596 0.019716
R50964 PAD.n3599 PAD.n3301 0.019716
R50965 PAD.n3600 PAD.n3599 0.019716
R50966 PAD.n3609 PAD.n3300 0.019716
R50967 PAD.n3609 PAD.n3608 0.019716
R50968 PAD.n3611 PAD.n3299 0.019716
R50969 PAD.n3612 PAD.n3611 0.019716
R50970 PAD.n3621 PAD.n3298 0.019716
R50971 PAD.n3621 PAD.n3620 0.019716
R50972 PAD.n3623 PAD.n3297 0.019716
R50973 PAD.n3624 PAD.n3623 0.019716
R50974 PAD.n8491 PAD.n8490 0.019716
R50975 PAD.n3728 PAD.n3683 0.019716
R50976 PAD.n3729 PAD.n3682 0.019716
R50977 PAD.n3738 PAD.n3681 0.019716
R50978 PAD.n3738 PAD.n3737 0.019716
R50979 PAD.n3740 PAD.n3680 0.019716
R50980 PAD.n3741 PAD.n3740 0.019716
R50981 PAD.n3750 PAD.n3679 0.019716
R50982 PAD.n3750 PAD.n3749 0.019716
R50983 PAD.n3752 PAD.n3678 0.019716
R50984 PAD.n3753 PAD.n3752 0.019716
R50985 PAD.n3762 PAD.n3677 0.019716
R50986 PAD.n3762 PAD.n3761 0.019716
R50987 PAD.n3764 PAD.n3676 0.019716
R50988 PAD.n3765 PAD.n3764 0.019716
R50989 PAD.n3774 PAD.n3675 0.019716
R50990 PAD.n3774 PAD.n3773 0.019716
R50991 PAD.n3776 PAD.n3674 0.019716
R50992 PAD.n3777 PAD.n3776 0.019716
R50993 PAD.n3786 PAD.n3673 0.019716
R50994 PAD.n3786 PAD.n3785 0.019716
R50995 PAD.n3788 PAD.n3672 0.019716
R50996 PAD.n3789 PAD.n3788 0.019716
R50997 PAD.n3798 PAD.n3671 0.019716
R50998 PAD.n3798 PAD.n3797 0.019716
R50999 PAD.n3800 PAD.n3670 0.019716
R51000 PAD.n3801 PAD.n3800 0.019716
R51001 PAD.n3810 PAD.n3669 0.019716
R51002 PAD.n3810 PAD.n3809 0.019716
R51003 PAD.n3812 PAD.n3668 0.019716
R51004 PAD.n3813 PAD.n3812 0.019716
R51005 PAD.n3822 PAD.n3667 0.019716
R51006 PAD.n3822 PAD.n3821 0.019716
R51007 PAD.n3824 PAD.n3666 0.019716
R51008 PAD.n3825 PAD.n3824 0.019716
R51009 PAD.n3834 PAD.n3665 0.019716
R51010 PAD.n3834 PAD.n3833 0.019716
R51011 PAD.n3836 PAD.n3664 0.019716
R51012 PAD.n3837 PAD.n3836 0.019716
R51013 PAD.n3846 PAD.n3663 0.019716
R51014 PAD.n3846 PAD.n3845 0.019716
R51015 PAD.n3848 PAD.n3662 0.019716
R51016 PAD.n3849 PAD.n3848 0.019716
R51017 PAD.n3858 PAD.n3661 0.019716
R51018 PAD.n3858 PAD.n3857 0.019716
R51019 PAD.n3860 PAD.n3660 0.019716
R51020 PAD.n3861 PAD.n3860 0.019716
R51021 PAD.n3870 PAD.n3659 0.019716
R51022 PAD.n3870 PAD.n3869 0.019716
R51023 PAD.n3872 PAD.n3658 0.019716
R51024 PAD.n3873 PAD.n3872 0.019716
R51025 PAD.n3882 PAD.n3657 0.019716
R51026 PAD.n3882 PAD.n3881 0.019716
R51027 PAD.n3884 PAD.n3656 0.019716
R51028 PAD.n3885 PAD.n3884 0.019716
R51029 PAD.n3894 PAD.n3655 0.019716
R51030 PAD.n3894 PAD.n3893 0.019716
R51031 PAD.n3896 PAD.n3654 0.019716
R51032 PAD.n3897 PAD.n3896 0.019716
R51033 PAD.n3906 PAD.n3653 0.019716
R51034 PAD.n3906 PAD.n3905 0.019716
R51035 PAD.n3908 PAD.n3652 0.019716
R51036 PAD.n3909 PAD.n3908 0.019716
R51037 PAD.n3918 PAD.n3651 0.019716
R51038 PAD.n3918 PAD.n3917 0.019716
R51039 PAD.n3920 PAD.n3650 0.019716
R51040 PAD.n3921 PAD.n3920 0.019716
R51041 PAD.n3930 PAD.n3649 0.019716
R51042 PAD.n3930 PAD.n3929 0.019716
R51043 PAD.n3932 PAD.n3648 0.019716
R51044 PAD.n3933 PAD.n3932 0.019716
R51045 PAD.n3942 PAD.n3647 0.019716
R51046 PAD.n3942 PAD.n3941 0.019716
R51047 PAD.n3944 PAD.n3646 0.019716
R51048 PAD.n3945 PAD.n3944 0.019716
R51049 PAD.n3954 PAD.n3645 0.019716
R51050 PAD.n3954 PAD.n3953 0.019716
R51051 PAD.n3956 PAD.n3644 0.019716
R51052 PAD.n3957 PAD.n3956 0.019716
R51053 PAD.n3966 PAD.n3643 0.019716
R51054 PAD.n3966 PAD.n3965 0.019716
R51055 PAD.n3968 PAD.n3642 0.019716
R51056 PAD.n3969 PAD.n3968 0.019716
R51057 PAD.n8467 PAD.n8466 0.019716
R51058 PAD.n4069 PAD.n4025 0.019716
R51059 PAD.n4070 PAD.n4024 0.019716
R51060 PAD.n4079 PAD.n4023 0.019716
R51061 PAD.n4079 PAD.n4078 0.019716
R51062 PAD.n4081 PAD.n4022 0.019716
R51063 PAD.n4082 PAD.n4081 0.019716
R51064 PAD.n4091 PAD.n4021 0.019716
R51065 PAD.n4091 PAD.n4090 0.019716
R51066 PAD.n4093 PAD.n4020 0.019716
R51067 PAD.n4094 PAD.n4093 0.019716
R51068 PAD.n4103 PAD.n4019 0.019716
R51069 PAD.n4103 PAD.n4102 0.019716
R51070 PAD.n4105 PAD.n4018 0.019716
R51071 PAD.n4106 PAD.n4105 0.019716
R51072 PAD.n4115 PAD.n4017 0.019716
R51073 PAD.n4115 PAD.n4114 0.019716
R51074 PAD.n4117 PAD.n4016 0.019716
R51075 PAD.n4118 PAD.n4117 0.019716
R51076 PAD.n4127 PAD.n4015 0.019716
R51077 PAD.n4127 PAD.n4126 0.019716
R51078 PAD.n4129 PAD.n4014 0.019716
R51079 PAD.n4130 PAD.n4129 0.019716
R51080 PAD.n4139 PAD.n4013 0.019716
R51081 PAD.n4139 PAD.n4138 0.019716
R51082 PAD.n4141 PAD.n4012 0.019716
R51083 PAD.n4142 PAD.n4141 0.019716
R51084 PAD.n4151 PAD.n4011 0.019716
R51085 PAD.n4151 PAD.n4150 0.019716
R51086 PAD.n4153 PAD.n4010 0.019716
R51087 PAD.n4154 PAD.n4153 0.019716
R51088 PAD.n4163 PAD.n4009 0.019716
R51089 PAD.n4163 PAD.n4162 0.019716
R51090 PAD.n4165 PAD.n4008 0.019716
R51091 PAD.n4166 PAD.n4165 0.019716
R51092 PAD.n4175 PAD.n4007 0.019716
R51093 PAD.n4175 PAD.n4174 0.019716
R51094 PAD.n4177 PAD.n4006 0.019716
R51095 PAD.n4178 PAD.n4177 0.019716
R51096 PAD.n4187 PAD.n4005 0.019716
R51097 PAD.n4187 PAD.n4186 0.019716
R51098 PAD.n4189 PAD.n4004 0.019716
R51099 PAD.n4190 PAD.n4189 0.019716
R51100 PAD.n4199 PAD.n4003 0.019716
R51101 PAD.n4199 PAD.n4198 0.019716
R51102 PAD.n4201 PAD.n4002 0.019716
R51103 PAD.n4202 PAD.n4201 0.019716
R51104 PAD.n4211 PAD.n4001 0.019716
R51105 PAD.n4211 PAD.n4210 0.019716
R51106 PAD.n4213 PAD.n4000 0.019716
R51107 PAD.n4214 PAD.n4213 0.019716
R51108 PAD.n4223 PAD.n3999 0.019716
R51109 PAD.n4223 PAD.n4222 0.019716
R51110 PAD.n4225 PAD.n3998 0.019716
R51111 PAD.n4226 PAD.n4225 0.019716
R51112 PAD.n4235 PAD.n3997 0.019716
R51113 PAD.n4235 PAD.n4234 0.019716
R51114 PAD.n4237 PAD.n3996 0.019716
R51115 PAD.n4238 PAD.n4237 0.019716
R51116 PAD.n4247 PAD.n3995 0.019716
R51117 PAD.n4247 PAD.n4246 0.019716
R51118 PAD.n4249 PAD.n3994 0.019716
R51119 PAD.n4250 PAD.n4249 0.019716
R51120 PAD.n4259 PAD.n3993 0.019716
R51121 PAD.n4259 PAD.n4258 0.019716
R51122 PAD.n4261 PAD.n3992 0.019716
R51123 PAD.n4262 PAD.n4261 0.019716
R51124 PAD.n4271 PAD.n3991 0.019716
R51125 PAD.n4271 PAD.n4270 0.019716
R51126 PAD.n4273 PAD.n3990 0.019716
R51127 PAD.n4274 PAD.n4273 0.019716
R51128 PAD.n4283 PAD.n3989 0.019716
R51129 PAD.n4283 PAD.n4282 0.019716
R51130 PAD.n4285 PAD.n3988 0.019716
R51131 PAD.n4286 PAD.n4285 0.019716
R51132 PAD.n4295 PAD.n3987 0.019716
R51133 PAD.n4295 PAD.n4294 0.019716
R51134 PAD.n4297 PAD.n3986 0.019716
R51135 PAD.n4298 PAD.n4297 0.019716
R51136 PAD.n4307 PAD.n3985 0.019716
R51137 PAD.n4307 PAD.n4306 0.019716
R51138 PAD.n4309 PAD.n3984 0.019716
R51139 PAD.n4310 PAD.n4309 0.019716
R51140 PAD.n8443 PAD.n8442 0.019716
R51141 PAD.n4421 PAD.n4420 0.019716
R51142 PAD.n4423 PAD.n4422 0.019716
R51143 PAD.n4424 PAD.n4415 0.019716
R51144 PAD.n4425 PAD.n4424 0.019716
R51145 PAD.n4435 PAD.n4434 0.019716
R51146 PAD.n4434 PAD.n4433 0.019716
R51147 PAD.n4436 PAD.n4411 0.019716
R51148 PAD.n4437 PAD.n4436 0.019716
R51149 PAD.n4447 PAD.n4446 0.019716
R51150 PAD.n4446 PAD.n4445 0.019716
R51151 PAD.n4448 PAD.n4407 0.019716
R51152 PAD.n4449 PAD.n4448 0.019716
R51153 PAD.n4459 PAD.n4458 0.019716
R51154 PAD.n4458 PAD.n4457 0.019716
R51155 PAD.n4460 PAD.n4403 0.019716
R51156 PAD.n4461 PAD.n4460 0.019716
R51157 PAD.n4471 PAD.n4470 0.019716
R51158 PAD.n4470 PAD.n4469 0.019716
R51159 PAD.n4472 PAD.n4399 0.019716
R51160 PAD.n4473 PAD.n4472 0.019716
R51161 PAD.n4483 PAD.n4482 0.019716
R51162 PAD.n4482 PAD.n4481 0.019716
R51163 PAD.n4484 PAD.n4395 0.019716
R51164 PAD.n4485 PAD.n4484 0.019716
R51165 PAD.n4495 PAD.n4494 0.019716
R51166 PAD.n4494 PAD.n4493 0.019716
R51167 PAD.n4496 PAD.n4391 0.019716
R51168 PAD.n4497 PAD.n4496 0.019716
R51169 PAD.n4507 PAD.n4506 0.019716
R51170 PAD.n4506 PAD.n4505 0.019716
R51171 PAD.n4508 PAD.n4387 0.019716
R51172 PAD.n4509 PAD.n4508 0.019716
R51173 PAD.n4519 PAD.n4518 0.019716
R51174 PAD.n4518 PAD.n4517 0.019716
R51175 PAD.n4520 PAD.n4383 0.019716
R51176 PAD.n4521 PAD.n4520 0.019716
R51177 PAD.n4531 PAD.n4530 0.019716
R51178 PAD.n4530 PAD.n4529 0.019716
R51179 PAD.n4532 PAD.n4379 0.019716
R51180 PAD.n4533 PAD.n4532 0.019716
R51181 PAD.n4543 PAD.n4542 0.019716
R51182 PAD.n4542 PAD.n4541 0.019716
R51183 PAD.n4544 PAD.n4375 0.019716
R51184 PAD.n4545 PAD.n4544 0.019716
R51185 PAD.n4555 PAD.n4554 0.019716
R51186 PAD.n4554 PAD.n4553 0.019716
R51187 PAD.n4556 PAD.n4371 0.019716
R51188 PAD.n4557 PAD.n4556 0.019716
R51189 PAD.n4567 PAD.n4566 0.019716
R51190 PAD.n4566 PAD.n4565 0.019716
R51191 PAD.n4568 PAD.n4367 0.019716
R51192 PAD.n4569 PAD.n4568 0.019716
R51193 PAD.n4579 PAD.n4578 0.019716
R51194 PAD.n4578 PAD.n4577 0.019716
R51195 PAD.n4580 PAD.n4363 0.019716
R51196 PAD.n4581 PAD.n4580 0.019716
R51197 PAD.n4591 PAD.n4590 0.019716
R51198 PAD.n4590 PAD.n4589 0.019716
R51199 PAD.n4592 PAD.n4359 0.019716
R51200 PAD.n4593 PAD.n4592 0.019716
R51201 PAD.n4603 PAD.n4602 0.019716
R51202 PAD.n4602 PAD.n4601 0.019716
R51203 PAD.n4604 PAD.n4355 0.019716
R51204 PAD.n4605 PAD.n4604 0.019716
R51205 PAD.n4615 PAD.n4614 0.019716
R51206 PAD.n4614 PAD.n4613 0.019716
R51207 PAD.n4616 PAD.n4351 0.019716
R51208 PAD.n4617 PAD.n4616 0.019716
R51209 PAD.n4627 PAD.n4626 0.019716
R51210 PAD.n4626 PAD.n4625 0.019716
R51211 PAD.n4628 PAD.n4347 0.019716
R51212 PAD.n4629 PAD.n4628 0.019716
R51213 PAD.n4639 PAD.n4638 0.019716
R51214 PAD.n4638 PAD.n4637 0.019716
R51215 PAD.n4640 PAD.n4343 0.019716
R51216 PAD.n4641 PAD.n4640 0.019716
R51217 PAD.n4651 PAD.n4650 0.019716
R51218 PAD.n4650 PAD.n4649 0.019716
R51219 PAD.n4652 PAD.n4339 0.019716
R51220 PAD.n4653 PAD.n4652 0.019716
R51221 PAD.n4664 PAD.n4663 0.019716
R51222 PAD.n4663 PAD.n4662 0.019716
R51223 PAD.n4667 PAD.n4666 0.019716
R51224 PAD.n8396 PAD.n8395 0.019716
R51225 PAD.n4726 PAD.n4725 0.019716
R51226 PAD.n8388 PAD.n8387 0.019716
R51227 PAD.n8388 PAD.n4723 0.019716
R51228 PAD.n4733 PAD.n4732 0.019716
R51229 PAD.n4733 PAD.n4722 0.019716
R51230 PAD.n8379 PAD.n8378 0.019716
R51231 PAD.n8379 PAD.n4721 0.019716
R51232 PAD.n4738 PAD.n4737 0.019716
R51233 PAD.n4738 PAD.n4720 0.019716
R51234 PAD.n8370 PAD.n8369 0.019716
R51235 PAD.n8370 PAD.n4719 0.019716
R51236 PAD.n4743 PAD.n4742 0.019716
R51237 PAD.n4743 PAD.n4718 0.019716
R51238 PAD.n8361 PAD.n8360 0.019716
R51239 PAD.n8361 PAD.n4717 0.019716
R51240 PAD.n4748 PAD.n4747 0.019716
R51241 PAD.n4748 PAD.n4716 0.019716
R51242 PAD.n8352 PAD.n8351 0.019716
R51243 PAD.n8352 PAD.n4715 0.019716
R51244 PAD.n4753 PAD.n4752 0.019716
R51245 PAD.n4753 PAD.n4714 0.019716
R51246 PAD.n8343 PAD.n8342 0.019716
R51247 PAD.n8343 PAD.n4713 0.019716
R51248 PAD.n4758 PAD.n4757 0.019716
R51249 PAD.n4758 PAD.n4712 0.019716
R51250 PAD.n8334 PAD.n8333 0.019716
R51251 PAD.n8334 PAD.n4711 0.019716
R51252 PAD.n4763 PAD.n4762 0.019716
R51253 PAD.n4763 PAD.n4710 0.019716
R51254 PAD.n8325 PAD.n8324 0.019716
R51255 PAD.n8325 PAD.n4709 0.019716
R51256 PAD.n4768 PAD.n4767 0.019716
R51257 PAD.n4768 PAD.n4708 0.019716
R51258 PAD.n8316 PAD.n8315 0.019716
R51259 PAD.n8316 PAD.n4707 0.019716
R51260 PAD.n4773 PAD.n4772 0.019716
R51261 PAD.n4773 PAD.n4706 0.019716
R51262 PAD.n8307 PAD.n8306 0.019716
R51263 PAD.n8307 PAD.n4705 0.019716
R51264 PAD.n4778 PAD.n4777 0.019716
R51265 PAD.n4778 PAD.n4704 0.019716
R51266 PAD.n8298 PAD.n8297 0.019716
R51267 PAD.n8298 PAD.n4703 0.019716
R51268 PAD.n4783 PAD.n4782 0.019716
R51269 PAD.n4783 PAD.n4702 0.019716
R51270 PAD.n8289 PAD.n8288 0.019716
R51271 PAD.n8289 PAD.n4701 0.019716
R51272 PAD.n4788 PAD.n4787 0.019716
R51273 PAD.n4788 PAD.n4700 0.019716
R51274 PAD.n8280 PAD.n8279 0.019716
R51275 PAD.n8280 PAD.n4699 0.019716
R51276 PAD.n4793 PAD.n4792 0.019716
R51277 PAD.n4793 PAD.n4698 0.019716
R51278 PAD.n8271 PAD.n8270 0.019716
R51279 PAD.n8271 PAD.n4697 0.019716
R51280 PAD.n4798 PAD.n4797 0.019716
R51281 PAD.n4798 PAD.n4696 0.019716
R51282 PAD.n8262 PAD.n8261 0.019716
R51283 PAD.n8262 PAD.n4695 0.019716
R51284 PAD.n4803 PAD.n4802 0.019716
R51285 PAD.n4803 PAD.n4694 0.019716
R51286 PAD.n8253 PAD.n8252 0.019716
R51287 PAD.n8253 PAD.n4693 0.019716
R51288 PAD.n4808 PAD.n4807 0.019716
R51289 PAD.n4808 PAD.n4692 0.019716
R51290 PAD.n8244 PAD.n8243 0.019716
R51291 PAD.n8244 PAD.n4691 0.019716
R51292 PAD.n4813 PAD.n4812 0.019716
R51293 PAD.n4813 PAD.n4690 0.019716
R51294 PAD.n8235 PAD.n8234 0.019716
R51295 PAD.n8235 PAD.n4689 0.019716
R51296 PAD.n4818 PAD.n4817 0.019716
R51297 PAD.n4818 PAD.n4688 0.019716
R51298 PAD.n8226 PAD.n8225 0.019716
R51299 PAD.n8226 PAD.n4687 0.019716
R51300 PAD.n4823 PAD.n4822 0.019716
R51301 PAD.n4823 PAD.n4686 0.019716
R51302 PAD.n8217 PAD.n8216 0.019716
R51303 PAD.n8217 PAD.n4685 0.019716
R51304 PAD.n4828 PAD.n4827 0.019716
R51305 PAD.n4828 PAD.n4684 0.019716
R51306 PAD.n4832 PAD.n4683 0.019716
R51307 PAD.n4849 PAD.n4847 0.019716
R51308 PAD.n5176 PAD.n5175 0.019716
R51309 PAD.n5172 PAD.n4850 0.019716
R51310 PAD.n5173 PAD.n5172 0.019716
R51311 PAD.n5166 PAD.n5163 0.019716
R51312 PAD.n5166 PAD.n5165 0.019716
R51313 PAD.n5160 PAD.n4855 0.019716
R51314 PAD.n5161 PAD.n5160 0.019716
R51315 PAD.n5154 PAD.n5151 0.019716
R51316 PAD.n5154 PAD.n5153 0.019716
R51317 PAD.n5148 PAD.n4859 0.019716
R51318 PAD.n5149 PAD.n5148 0.019716
R51319 PAD.n5142 PAD.n5139 0.019716
R51320 PAD.n5142 PAD.n5141 0.019716
R51321 PAD.n5136 PAD.n4863 0.019716
R51322 PAD.n5137 PAD.n5136 0.019716
R51323 PAD.n5130 PAD.n5127 0.019716
R51324 PAD.n5130 PAD.n5129 0.019716
R51325 PAD.n5124 PAD.n4867 0.019716
R51326 PAD.n5125 PAD.n5124 0.019716
R51327 PAD.n5118 PAD.n5115 0.019716
R51328 PAD.n5118 PAD.n5117 0.019716
R51329 PAD.n5112 PAD.n4871 0.019716
R51330 PAD.n5113 PAD.n5112 0.019716
R51331 PAD.n5106 PAD.n5103 0.019716
R51332 PAD.n5106 PAD.n5105 0.019716
R51333 PAD.n5100 PAD.n4875 0.019716
R51334 PAD.n5101 PAD.n5100 0.019716
R51335 PAD.n5094 PAD.n5091 0.019716
R51336 PAD.n5094 PAD.n5093 0.019716
R51337 PAD.n5088 PAD.n4879 0.019716
R51338 PAD.n5089 PAD.n5088 0.019716
R51339 PAD.n5082 PAD.n5079 0.019716
R51340 PAD.n5082 PAD.n5081 0.019716
R51341 PAD.n5076 PAD.n4883 0.019716
R51342 PAD.n5077 PAD.n5076 0.019716
R51343 PAD.n5070 PAD.n5067 0.019716
R51344 PAD.n5070 PAD.n5069 0.019716
R51345 PAD.n5064 PAD.n4887 0.019716
R51346 PAD.n5065 PAD.n5064 0.019716
R51347 PAD.n5058 PAD.n5055 0.019716
R51348 PAD.n5058 PAD.n5057 0.019716
R51349 PAD.n5052 PAD.n4891 0.019716
R51350 PAD.n5053 PAD.n5052 0.019716
R51351 PAD.n5046 PAD.n5043 0.019716
R51352 PAD.n5046 PAD.n5045 0.019716
R51353 PAD.n5040 PAD.n4895 0.019716
R51354 PAD.n5041 PAD.n5040 0.019716
R51355 PAD.n5034 PAD.n5031 0.019716
R51356 PAD.n5034 PAD.n5033 0.019716
R51357 PAD.n5028 PAD.n4899 0.019716
R51358 PAD.n5029 PAD.n5028 0.019716
R51359 PAD.n5022 PAD.n5019 0.019716
R51360 PAD.n5022 PAD.n5021 0.019716
R51361 PAD.n5016 PAD.n4903 0.019716
R51362 PAD.n5017 PAD.n5016 0.019716
R51363 PAD.n5010 PAD.n5007 0.019716
R51364 PAD.n5010 PAD.n5009 0.019716
R51365 PAD.n5004 PAD.n4907 0.019716
R51366 PAD.n5005 PAD.n5004 0.019716
R51367 PAD.n4998 PAD.n4995 0.019716
R51368 PAD.n4998 PAD.n4997 0.019716
R51369 PAD.n4992 PAD.n4911 0.019716
R51370 PAD.n4993 PAD.n4992 0.019716
R51371 PAD.n4986 PAD.n4983 0.019716
R51372 PAD.n4986 PAD.n4985 0.019716
R51373 PAD.n4980 PAD.n4915 0.019716
R51374 PAD.n4981 PAD.n4980 0.019716
R51375 PAD.n4974 PAD.n4971 0.019716
R51376 PAD.n4974 PAD.n4973 0.019716
R51377 PAD.n4968 PAD.n4919 0.019716
R51378 PAD.n4969 PAD.n4968 0.019716
R51379 PAD.n4962 PAD.n4959 0.019716
R51380 PAD.n4962 PAD.n4961 0.019716
R51381 PAD.n4956 PAD.n4923 0.019716
R51382 PAD.n4957 PAD.n4956 0.019716
R51383 PAD.n4950 PAD.n4947 0.019716
R51384 PAD.n4950 PAD.n4949 0.019716
R51385 PAD.n4944 PAD.n4927 0.019716
R51386 PAD.n4945 PAD.n4944 0.019716
R51387 PAD.n4938 PAD.n4935 0.019716
R51388 PAD.n4938 PAD.n4937 0.019716
R51389 PAD.n4933 PAD.n4932 0.019716
R51390 PAD.n8162 PAD.n8161 0.019716
R51391 PAD.n7872 PAD.n7871 0.019716
R51392 PAD.n8154 PAD.n8153 0.019716
R51393 PAD.n8154 PAD.n7870 0.019716
R51394 PAD.n7879 PAD.n7878 0.019716
R51395 PAD.n7879 PAD.n7869 0.019716
R51396 PAD.n8145 PAD.n8144 0.019716
R51397 PAD.n8145 PAD.n7868 0.019716
R51398 PAD.n7884 PAD.n7883 0.019716
R51399 PAD.n7884 PAD.n7867 0.019716
R51400 PAD.n8136 PAD.n8135 0.019716
R51401 PAD.n8136 PAD.n7866 0.019716
R51402 PAD.n7889 PAD.n7888 0.019716
R51403 PAD.n7889 PAD.n7865 0.019716
R51404 PAD.n8127 PAD.n8126 0.019716
R51405 PAD.n8127 PAD.n7864 0.019716
R51406 PAD.n7894 PAD.n7893 0.019716
R51407 PAD.n7894 PAD.n7863 0.019716
R51408 PAD.n8118 PAD.n8117 0.019716
R51409 PAD.n8118 PAD.n7862 0.019716
R51410 PAD.n7899 PAD.n7898 0.019716
R51411 PAD.n7899 PAD.n7861 0.019716
R51412 PAD.n8109 PAD.n8108 0.019716
R51413 PAD.n8109 PAD.n7860 0.019716
R51414 PAD.n7904 PAD.n7903 0.019716
R51415 PAD.n7904 PAD.n7859 0.019716
R51416 PAD.n8100 PAD.n8099 0.019716
R51417 PAD.n8100 PAD.n7858 0.019716
R51418 PAD.n7909 PAD.n7908 0.019716
R51419 PAD.n7909 PAD.n7857 0.019716
R51420 PAD.n8091 PAD.n8090 0.019716
R51421 PAD.n8091 PAD.n7856 0.019716
R51422 PAD.n7914 PAD.n7913 0.019716
R51423 PAD.n7914 PAD.n7855 0.019716
R51424 PAD.n8082 PAD.n8081 0.019716
R51425 PAD.n8082 PAD.n7854 0.019716
R51426 PAD.n7919 PAD.n7918 0.019716
R51427 PAD.n7919 PAD.n7853 0.019716
R51428 PAD.n8073 PAD.n8072 0.019716
R51429 PAD.n8073 PAD.n7852 0.019716
R51430 PAD.n7924 PAD.n7923 0.019716
R51431 PAD.n7924 PAD.n7851 0.019716
R51432 PAD.n8064 PAD.n8063 0.019716
R51433 PAD.n8064 PAD.n7850 0.019716
R51434 PAD.n7929 PAD.n7928 0.019716
R51435 PAD.n7929 PAD.n7849 0.019716
R51436 PAD.n8055 PAD.n8054 0.019716
R51437 PAD.n8055 PAD.n7848 0.019716
R51438 PAD.n7934 PAD.n7933 0.019716
R51439 PAD.n7934 PAD.n7847 0.019716
R51440 PAD.n8046 PAD.n8045 0.019716
R51441 PAD.n8046 PAD.n7846 0.019716
R51442 PAD.n7939 PAD.n7938 0.019716
R51443 PAD.n7939 PAD.n7845 0.019716
R51444 PAD.n8037 PAD.n8036 0.019716
R51445 PAD.n8037 PAD.n7844 0.019716
R51446 PAD.n7944 PAD.n7943 0.019716
R51447 PAD.n7944 PAD.n7843 0.019716
R51448 PAD.n8028 PAD.n8027 0.019716
R51449 PAD.n8028 PAD.n7842 0.019716
R51450 PAD.n7949 PAD.n7948 0.019716
R51451 PAD.n7949 PAD.n7841 0.019716
R51452 PAD.n8019 PAD.n8018 0.019716
R51453 PAD.n8019 PAD.n7840 0.019716
R51454 PAD.n7954 PAD.n7953 0.019716
R51455 PAD.n7954 PAD.n7839 0.019716
R51456 PAD.n8010 PAD.n8009 0.019716
R51457 PAD.n8010 PAD.n7838 0.019716
R51458 PAD.n7959 PAD.n7958 0.019716
R51459 PAD.n7959 PAD.n7837 0.019716
R51460 PAD.n8001 PAD.n8000 0.019716
R51461 PAD.n8001 PAD.n7836 0.019716
R51462 PAD.n7964 PAD.n7963 0.019716
R51463 PAD.n7964 PAD.n7835 0.019716
R51464 PAD.n7992 PAD.n7991 0.019716
R51465 PAD.n7992 PAD.n7834 0.019716
R51466 PAD.n7969 PAD.n7968 0.019716
R51467 PAD.n7969 PAD.n7833 0.019716
R51468 PAD.n7983 PAD.n7982 0.019716
R51469 PAD.n7983 PAD.n7832 0.019716
R51470 PAD.n7976 PAD.n7975 0.019716
R51471 PAD.n7976 PAD.n7831 0.019716
R51472 PAD.n7971 PAD.n7830 0.019716
R51473 PAD.n5213 PAD.n5211 0.019716
R51474 PAD.n5540 PAD.n5539 0.019716
R51475 PAD.n5536 PAD.n5214 0.019716
R51476 PAD.n5537 PAD.n5536 0.019716
R51477 PAD.n5530 PAD.n5527 0.019716
R51478 PAD.n5530 PAD.n5529 0.019716
R51479 PAD.n5524 PAD.n5219 0.019716
R51480 PAD.n5525 PAD.n5524 0.019716
R51481 PAD.n5518 PAD.n5515 0.019716
R51482 PAD.n5518 PAD.n5517 0.019716
R51483 PAD.n5512 PAD.n5223 0.019716
R51484 PAD.n5513 PAD.n5512 0.019716
R51485 PAD.n5506 PAD.n5503 0.019716
R51486 PAD.n5506 PAD.n5505 0.019716
R51487 PAD.n5500 PAD.n5227 0.019716
R51488 PAD.n5501 PAD.n5500 0.019716
R51489 PAD.n5494 PAD.n5491 0.019716
R51490 PAD.n5494 PAD.n5493 0.019716
R51491 PAD.n5488 PAD.n5231 0.019716
R51492 PAD.n5489 PAD.n5488 0.019716
R51493 PAD.n5482 PAD.n5479 0.019716
R51494 PAD.n5482 PAD.n5481 0.019716
R51495 PAD.n5476 PAD.n5235 0.019716
R51496 PAD.n5477 PAD.n5476 0.019716
R51497 PAD.n5470 PAD.n5467 0.019716
R51498 PAD.n5470 PAD.n5469 0.019716
R51499 PAD.n5464 PAD.n5239 0.019716
R51500 PAD.n5465 PAD.n5464 0.019716
R51501 PAD.n5458 PAD.n5455 0.019716
R51502 PAD.n5458 PAD.n5457 0.019716
R51503 PAD.n5452 PAD.n5243 0.019716
R51504 PAD.n5453 PAD.n5452 0.019716
R51505 PAD.n5446 PAD.n5443 0.019716
R51506 PAD.n5446 PAD.n5445 0.019716
R51507 PAD.n5440 PAD.n5247 0.019716
R51508 PAD.n5441 PAD.n5440 0.019716
R51509 PAD.n5434 PAD.n5431 0.019716
R51510 PAD.n5434 PAD.n5433 0.019716
R51511 PAD.n5428 PAD.n5251 0.019716
R51512 PAD.n5429 PAD.n5428 0.019716
R51513 PAD.n5422 PAD.n5419 0.019716
R51514 PAD.n5422 PAD.n5421 0.019716
R51515 PAD.n5416 PAD.n5255 0.019716
R51516 PAD.n5417 PAD.n5416 0.019716
R51517 PAD.n5410 PAD.n5407 0.019716
R51518 PAD.n5410 PAD.n5409 0.019716
R51519 PAD.n5404 PAD.n5259 0.019716
R51520 PAD.n5405 PAD.n5404 0.019716
R51521 PAD.n5398 PAD.n5395 0.019716
R51522 PAD.n5398 PAD.n5397 0.019716
R51523 PAD.n5392 PAD.n5263 0.019716
R51524 PAD.n5393 PAD.n5392 0.019716
R51525 PAD.n5386 PAD.n5383 0.019716
R51526 PAD.n5386 PAD.n5385 0.019716
R51527 PAD.n5380 PAD.n5267 0.019716
R51528 PAD.n5381 PAD.n5380 0.019716
R51529 PAD.n5374 PAD.n5371 0.019716
R51530 PAD.n5374 PAD.n5373 0.019716
R51531 PAD.n5368 PAD.n5271 0.019716
R51532 PAD.n5369 PAD.n5368 0.019716
R51533 PAD.n5362 PAD.n5359 0.019716
R51534 PAD.n5362 PAD.n5361 0.019716
R51535 PAD.n5356 PAD.n5275 0.019716
R51536 PAD.n5357 PAD.n5356 0.019716
R51537 PAD.n5350 PAD.n5347 0.019716
R51538 PAD.n5350 PAD.n5349 0.019716
R51539 PAD.n5344 PAD.n5279 0.019716
R51540 PAD.n5345 PAD.n5344 0.019716
R51541 PAD.n5338 PAD.n5335 0.019716
R51542 PAD.n5338 PAD.n5337 0.019716
R51543 PAD.n5332 PAD.n5283 0.019716
R51544 PAD.n5333 PAD.n5332 0.019716
R51545 PAD.n5326 PAD.n5323 0.019716
R51546 PAD.n5326 PAD.n5325 0.019716
R51547 PAD.n5320 PAD.n5287 0.019716
R51548 PAD.n5321 PAD.n5320 0.019716
R51549 PAD.n5314 PAD.n5311 0.019716
R51550 PAD.n5314 PAD.n5313 0.019716
R51551 PAD.n5308 PAD.n5291 0.019716
R51552 PAD.n5309 PAD.n5308 0.019716
R51553 PAD.n5302 PAD.n5299 0.019716
R51554 PAD.n5302 PAD.n5301 0.019716
R51555 PAD.n5297 PAD.n5296 0.019716
R51556 PAD.n7519 PAD.n7518 0.019716
R51557 PAD.n7511 PAD.n7201 0.019716
R51558 PAD.n7509 PAD.n7508 0.019716
R51559 PAD.n7509 PAD.n7199 0.019716
R51560 PAD.n7500 PAD.n7499 0.019716
R51561 PAD.n7499 PAD.n7198 0.019716
R51562 PAD.n7497 PAD.n7496 0.019716
R51563 PAD.n7497 PAD.n7197 0.019716
R51564 PAD.n7488 PAD.n7487 0.019716
R51565 PAD.n7487 PAD.n7196 0.019716
R51566 PAD.n7485 PAD.n7484 0.019716
R51567 PAD.n7485 PAD.n7195 0.019716
R51568 PAD.n7476 PAD.n7475 0.019716
R51569 PAD.n7475 PAD.n7194 0.019716
R51570 PAD.n7473 PAD.n7472 0.019716
R51571 PAD.n7473 PAD.n7193 0.019716
R51572 PAD.n7464 PAD.n7463 0.019716
R51573 PAD.n7463 PAD.n7192 0.019716
R51574 PAD.n7461 PAD.n7460 0.019716
R51575 PAD.n7461 PAD.n7191 0.019716
R51576 PAD.n7452 PAD.n7451 0.019716
R51577 PAD.n7451 PAD.n7190 0.019716
R51578 PAD.n7449 PAD.n7448 0.019716
R51579 PAD.n7449 PAD.n7189 0.019716
R51580 PAD.n7440 PAD.n7439 0.019716
R51581 PAD.n7439 PAD.n7188 0.019716
R51582 PAD.n7437 PAD.n7436 0.019716
R51583 PAD.n7437 PAD.n7187 0.019716
R51584 PAD.n7428 PAD.n7427 0.019716
R51585 PAD.n7427 PAD.n7186 0.019716
R51586 PAD.n7425 PAD.n7424 0.019716
R51587 PAD.n7425 PAD.n7185 0.019716
R51588 PAD.n7416 PAD.n7415 0.019716
R51589 PAD.n7415 PAD.n7184 0.019716
R51590 PAD.n7413 PAD.n7412 0.019716
R51591 PAD.n7413 PAD.n7183 0.019716
R51592 PAD.n7404 PAD.n7403 0.019716
R51593 PAD.n7403 PAD.n7182 0.019716
R51594 PAD.n7401 PAD.n7400 0.019716
R51595 PAD.n7401 PAD.n7181 0.019716
R51596 PAD.n7392 PAD.n7391 0.019716
R51597 PAD.n7391 PAD.n7180 0.019716
R51598 PAD.n7389 PAD.n7388 0.019716
R51599 PAD.n7389 PAD.n7179 0.019716
R51600 PAD.n7380 PAD.n7379 0.019716
R51601 PAD.n7379 PAD.n7178 0.019716
R51602 PAD.n7377 PAD.n7376 0.019716
R51603 PAD.n7377 PAD.n7177 0.019716
R51604 PAD.n7368 PAD.n7367 0.019716
R51605 PAD.n7367 PAD.n7176 0.019716
R51606 PAD.n7365 PAD.n7364 0.019716
R51607 PAD.n7365 PAD.n7175 0.019716
R51608 PAD.n7356 PAD.n7355 0.019716
R51609 PAD.n7355 PAD.n7174 0.019716
R51610 PAD.n7353 PAD.n7352 0.019716
R51611 PAD.n7353 PAD.n7173 0.019716
R51612 PAD.n7344 PAD.n7343 0.019716
R51613 PAD.n7343 PAD.n7172 0.019716
R51614 PAD.n7341 PAD.n7340 0.019716
R51615 PAD.n7341 PAD.n7171 0.019716
R51616 PAD.n7332 PAD.n7331 0.019716
R51617 PAD.n7331 PAD.n7170 0.019716
R51618 PAD.n7329 PAD.n7328 0.019716
R51619 PAD.n7329 PAD.n7169 0.019716
R51620 PAD.n7320 PAD.n7319 0.019716
R51621 PAD.n7319 PAD.n7168 0.019716
R51622 PAD.n7317 PAD.n7316 0.019716
R51623 PAD.n7317 PAD.n7167 0.019716
R51624 PAD.n7308 PAD.n7307 0.019716
R51625 PAD.n7307 PAD.n7166 0.019716
R51626 PAD.n7305 PAD.n7304 0.019716
R51627 PAD.n7305 PAD.n7165 0.019716
R51628 PAD.n7296 PAD.n7295 0.019716
R51629 PAD.n7295 PAD.n7164 0.019716
R51630 PAD.n7293 PAD.n7292 0.019716
R51631 PAD.n7293 PAD.n7163 0.019716
R51632 PAD.n7284 PAD.n7283 0.019716
R51633 PAD.n7283 PAD.n7162 0.019716
R51634 PAD.n7281 PAD.n7280 0.019716
R51635 PAD.n7281 PAD.n7161 0.019716
R51636 PAD.n7272 PAD.n7271 0.019716
R51637 PAD.n7271 PAD.n7160 0.019716
R51638 PAD.n7269 PAD.n7159 0.019716
R51639 PAD.n7781 PAD.n7780 0.019716
R51640 PAD.n7773 PAD.n7104 0.019716
R51641 PAD.n7771 PAD.n7770 0.019716
R51642 PAD.n7771 PAD.n7102 0.019716
R51643 PAD.n7762 PAD.n7761 0.019716
R51644 PAD.n7761 PAD.n7101 0.019716
R51645 PAD.n7759 PAD.n7758 0.019716
R51646 PAD.n7759 PAD.n7100 0.019716
R51647 PAD.n7750 PAD.n7749 0.019716
R51648 PAD.n7749 PAD.n7099 0.019716
R51649 PAD.n7747 PAD.n7746 0.019716
R51650 PAD.n7747 PAD.n7098 0.019716
R51651 PAD.n7738 PAD.n7737 0.019716
R51652 PAD.n7737 PAD.n7097 0.019716
R51653 PAD.n7735 PAD.n7734 0.019716
R51654 PAD.n7735 PAD.n7096 0.019716
R51655 PAD.n7726 PAD.n7725 0.019716
R51656 PAD.n7725 PAD.n7095 0.019716
R51657 PAD.n7723 PAD.n7722 0.019716
R51658 PAD.n7723 PAD.n7094 0.019716
R51659 PAD.n7714 PAD.n7713 0.019716
R51660 PAD.n7713 PAD.n7093 0.019716
R51661 PAD.n7711 PAD.n7710 0.019716
R51662 PAD.n7711 PAD.n7092 0.019716
R51663 PAD.n7702 PAD.n7701 0.019716
R51664 PAD.n7701 PAD.n7091 0.019716
R51665 PAD.n7699 PAD.n7698 0.019716
R51666 PAD.n7699 PAD.n7090 0.019716
R51667 PAD.n7690 PAD.n7689 0.019716
R51668 PAD.n7689 PAD.n7089 0.019716
R51669 PAD.n7687 PAD.n7686 0.019716
R51670 PAD.n7687 PAD.n7088 0.019716
R51671 PAD.n7678 PAD.n7677 0.019716
R51672 PAD.n7677 PAD.n7087 0.019716
R51673 PAD.n7675 PAD.n7674 0.019716
R51674 PAD.n7675 PAD.n7086 0.019716
R51675 PAD.n7666 PAD.n7665 0.019716
R51676 PAD.n7665 PAD.n7085 0.019716
R51677 PAD.n7663 PAD.n7662 0.019716
R51678 PAD.n7663 PAD.n7084 0.019716
R51679 PAD.n7654 PAD.n7653 0.019716
R51680 PAD.n7653 PAD.n7083 0.019716
R51681 PAD.n7651 PAD.n7650 0.019716
R51682 PAD.n7651 PAD.n7082 0.019716
R51683 PAD.n7642 PAD.n7641 0.019716
R51684 PAD.n7641 PAD.n7081 0.019716
R51685 PAD.n7639 PAD.n7638 0.019716
R51686 PAD.n7639 PAD.n7080 0.019716
R51687 PAD.n7630 PAD.n7629 0.019716
R51688 PAD.n7629 PAD.n7079 0.019716
R51689 PAD.n7627 PAD.n7626 0.019716
R51690 PAD.n7627 PAD.n7078 0.019716
R51691 PAD.n7618 PAD.n7617 0.019716
R51692 PAD.n7617 PAD.n7077 0.019716
R51693 PAD.n7615 PAD.n7614 0.019716
R51694 PAD.n7615 PAD.n7076 0.019716
R51695 PAD.n7606 PAD.n7605 0.019716
R51696 PAD.n7605 PAD.n7075 0.019716
R51697 PAD.n7603 PAD.n7602 0.019716
R51698 PAD.n7603 PAD.n7074 0.019716
R51699 PAD.n7594 PAD.n7593 0.019716
R51700 PAD.n7593 PAD.n7073 0.019716
R51701 PAD.n7591 PAD.n7590 0.019716
R51702 PAD.n7591 PAD.n7072 0.019716
R51703 PAD.n7582 PAD.n7581 0.019716
R51704 PAD.n7581 PAD.n7071 0.019716
R51705 PAD.n7579 PAD.n7578 0.019716
R51706 PAD.n7579 PAD.n7070 0.019716
R51707 PAD.n7570 PAD.n7569 0.019716
R51708 PAD.n7569 PAD.n7069 0.019716
R51709 PAD.n7567 PAD.n7566 0.019716
R51710 PAD.n7567 PAD.n7068 0.019716
R51711 PAD.n7558 PAD.n7557 0.019716
R51712 PAD.n7557 PAD.n7067 0.019716
R51713 PAD.n7555 PAD.n7554 0.019716
R51714 PAD.n7555 PAD.n7066 0.019716
R51715 PAD.n7546 PAD.n7545 0.019716
R51716 PAD.n7545 PAD.n7065 0.019716
R51717 PAD.n7543 PAD.n7542 0.019716
R51718 PAD.n7543 PAD.n7064 0.019716
R51719 PAD.n7534 PAD.n7533 0.019716
R51720 PAD.n7533 PAD.n7063 0.019716
R51721 PAD.n7531 PAD.n7062 0.019716
R51722 PAD.n6721 PAD.n6719 0.019716
R51723 PAD.n7048 PAD.n7047 0.019716
R51724 PAD.n7044 PAD.n6722 0.019716
R51725 PAD.n7045 PAD.n7044 0.019716
R51726 PAD.n7038 PAD.n7035 0.019716
R51727 PAD.n7038 PAD.n7037 0.019716
R51728 PAD.n7032 PAD.n6727 0.019716
R51729 PAD.n7033 PAD.n7032 0.019716
R51730 PAD.n7026 PAD.n7023 0.019716
R51731 PAD.n7026 PAD.n7025 0.019716
R51732 PAD.n7020 PAD.n6731 0.019716
R51733 PAD.n7021 PAD.n7020 0.019716
R51734 PAD.n7014 PAD.n7011 0.019716
R51735 PAD.n7014 PAD.n7013 0.019716
R51736 PAD.n7008 PAD.n6735 0.019716
R51737 PAD.n7009 PAD.n7008 0.019716
R51738 PAD.n7002 PAD.n6999 0.019716
R51739 PAD.n7002 PAD.n7001 0.019716
R51740 PAD.n6996 PAD.n6739 0.019716
R51741 PAD.n6997 PAD.n6996 0.019716
R51742 PAD.n6990 PAD.n6987 0.019716
R51743 PAD.n6990 PAD.n6989 0.019716
R51744 PAD.n6984 PAD.n6743 0.019716
R51745 PAD.n6985 PAD.n6984 0.019716
R51746 PAD.n6978 PAD.n6975 0.019716
R51747 PAD.n6978 PAD.n6977 0.019716
R51748 PAD.n6972 PAD.n6747 0.019716
R51749 PAD.n6973 PAD.n6972 0.019716
R51750 PAD.n6966 PAD.n6963 0.019716
R51751 PAD.n6966 PAD.n6965 0.019716
R51752 PAD.n6960 PAD.n6751 0.019716
R51753 PAD.n6961 PAD.n6960 0.019716
R51754 PAD.n6954 PAD.n6951 0.019716
R51755 PAD.n6954 PAD.n6953 0.019716
R51756 PAD.n6948 PAD.n6755 0.019716
R51757 PAD.n6949 PAD.n6948 0.019716
R51758 PAD.n6942 PAD.n6939 0.019716
R51759 PAD.n6942 PAD.n6941 0.019716
R51760 PAD.n6936 PAD.n6759 0.019716
R51761 PAD.n6937 PAD.n6936 0.019716
R51762 PAD.n6930 PAD.n6927 0.019716
R51763 PAD.n6930 PAD.n6929 0.019716
R51764 PAD.n6924 PAD.n6763 0.019716
R51765 PAD.n6925 PAD.n6924 0.019716
R51766 PAD.n6918 PAD.n6915 0.019716
R51767 PAD.n6918 PAD.n6917 0.019716
R51768 PAD.n6912 PAD.n6767 0.019716
R51769 PAD.n6913 PAD.n6912 0.019716
R51770 PAD.n6906 PAD.n6903 0.019716
R51771 PAD.n6906 PAD.n6905 0.019716
R51772 PAD.n6900 PAD.n6771 0.019716
R51773 PAD.n6901 PAD.n6900 0.019716
R51774 PAD.n6894 PAD.n6891 0.019716
R51775 PAD.n6894 PAD.n6893 0.019716
R51776 PAD.n6888 PAD.n6775 0.019716
R51777 PAD.n6889 PAD.n6888 0.019716
R51778 PAD.n6882 PAD.n6879 0.019716
R51779 PAD.n6882 PAD.n6881 0.019716
R51780 PAD.n6876 PAD.n6779 0.019716
R51781 PAD.n6877 PAD.n6876 0.019716
R51782 PAD.n6870 PAD.n6867 0.019716
R51783 PAD.n6870 PAD.n6869 0.019716
R51784 PAD.n6864 PAD.n6783 0.019716
R51785 PAD.n6865 PAD.n6864 0.019716
R51786 PAD.n6858 PAD.n6855 0.019716
R51787 PAD.n6858 PAD.n6857 0.019716
R51788 PAD.n6852 PAD.n6787 0.019716
R51789 PAD.n6853 PAD.n6852 0.019716
R51790 PAD.n6846 PAD.n6843 0.019716
R51791 PAD.n6846 PAD.n6845 0.019716
R51792 PAD.n6840 PAD.n6791 0.019716
R51793 PAD.n6841 PAD.n6840 0.019716
R51794 PAD.n6834 PAD.n6831 0.019716
R51795 PAD.n6834 PAD.n6833 0.019716
R51796 PAD.n6828 PAD.n6795 0.019716
R51797 PAD.n6829 PAD.n6828 0.019716
R51798 PAD.n6822 PAD.n6819 0.019716
R51799 PAD.n6822 PAD.n6821 0.019716
R51800 PAD.n6816 PAD.n6799 0.019716
R51801 PAD.n6817 PAD.n6816 0.019716
R51802 PAD.n6810 PAD.n6807 0.019716
R51803 PAD.n6810 PAD.n6809 0.019716
R51804 PAD.n6805 PAD.n6804 0.019716
R51805 PAD.n5893 PAD.n5892 0.019716
R51806 PAD.n5603 PAD.n5602 0.019716
R51807 PAD.n5885 PAD.n5884 0.019716
R51808 PAD.n5885 PAD.n5601 0.019716
R51809 PAD.n5610 PAD.n5609 0.019716
R51810 PAD.n5610 PAD.n5600 0.019716
R51811 PAD.n5876 PAD.n5875 0.019716
R51812 PAD.n5876 PAD.n5599 0.019716
R51813 PAD.n5615 PAD.n5614 0.019716
R51814 PAD.n5615 PAD.n5598 0.019716
R51815 PAD.n5867 PAD.n5866 0.019716
R51816 PAD.n5867 PAD.n5597 0.019716
R51817 PAD.n5620 PAD.n5619 0.019716
R51818 PAD.n5620 PAD.n5596 0.019716
R51819 PAD.n5858 PAD.n5857 0.019716
R51820 PAD.n5858 PAD.n5595 0.019716
R51821 PAD.n5625 PAD.n5624 0.019716
R51822 PAD.n5625 PAD.n5594 0.019716
R51823 PAD.n5849 PAD.n5848 0.019716
R51824 PAD.n5849 PAD.n5593 0.019716
R51825 PAD.n5630 PAD.n5629 0.019716
R51826 PAD.n5630 PAD.n5592 0.019716
R51827 PAD.n5840 PAD.n5839 0.019716
R51828 PAD.n5840 PAD.n5591 0.019716
R51829 PAD.n5635 PAD.n5634 0.019716
R51830 PAD.n5635 PAD.n5590 0.019716
R51831 PAD.n5831 PAD.n5830 0.019716
R51832 PAD.n5831 PAD.n5589 0.019716
R51833 PAD.n5640 PAD.n5639 0.019716
R51834 PAD.n5640 PAD.n5588 0.019716
R51835 PAD.n5822 PAD.n5821 0.019716
R51836 PAD.n5822 PAD.n5587 0.019716
R51837 PAD.n5645 PAD.n5644 0.019716
R51838 PAD.n5645 PAD.n5586 0.019716
R51839 PAD.n5813 PAD.n5812 0.019716
R51840 PAD.n5813 PAD.n5585 0.019716
R51841 PAD.n5650 PAD.n5649 0.019716
R51842 PAD.n5650 PAD.n5584 0.019716
R51843 PAD.n5804 PAD.n5803 0.019716
R51844 PAD.n5804 PAD.n5583 0.019716
R51845 PAD.n5655 PAD.n5654 0.019716
R51846 PAD.n5655 PAD.n5582 0.019716
R51847 PAD.n5795 PAD.n5794 0.019716
R51848 PAD.n5795 PAD.n5581 0.019716
R51849 PAD.n5660 PAD.n5659 0.019716
R51850 PAD.n5660 PAD.n5580 0.019716
R51851 PAD.n5786 PAD.n5785 0.019716
R51852 PAD.n5786 PAD.n5579 0.019716
R51853 PAD.n5665 PAD.n5664 0.019716
R51854 PAD.n5665 PAD.n5578 0.019716
R51855 PAD.n5777 PAD.n5776 0.019716
R51856 PAD.n5777 PAD.n5577 0.019716
R51857 PAD.n5670 PAD.n5669 0.019716
R51858 PAD.n5670 PAD.n5576 0.019716
R51859 PAD.n5768 PAD.n5767 0.019716
R51860 PAD.n5768 PAD.n5575 0.019716
R51861 PAD.n5675 PAD.n5674 0.019716
R51862 PAD.n5675 PAD.n5574 0.019716
R51863 PAD.n5759 PAD.n5758 0.019716
R51864 PAD.n5759 PAD.n5573 0.019716
R51865 PAD.n5680 PAD.n5679 0.019716
R51866 PAD.n5680 PAD.n5572 0.019716
R51867 PAD.n5750 PAD.n5749 0.019716
R51868 PAD.n5750 PAD.n5571 0.019716
R51869 PAD.n5685 PAD.n5684 0.019716
R51870 PAD.n5685 PAD.n5570 0.019716
R51871 PAD.n5741 PAD.n5740 0.019716
R51872 PAD.n5741 PAD.n5569 0.019716
R51873 PAD.n5690 PAD.n5689 0.019716
R51874 PAD.n5690 PAD.n5568 0.019716
R51875 PAD.n5732 PAD.n5731 0.019716
R51876 PAD.n5732 PAD.n5567 0.019716
R51877 PAD.n5695 PAD.n5694 0.019716
R51878 PAD.n5695 PAD.n5566 0.019716
R51879 PAD.n5723 PAD.n5722 0.019716
R51880 PAD.n5723 PAD.n5565 0.019716
R51881 PAD.n5700 PAD.n5699 0.019716
R51882 PAD.n5700 PAD.n5564 0.019716
R51883 PAD.n5714 PAD.n5713 0.019716
R51884 PAD.n5714 PAD.n5563 0.019716
R51885 PAD.n5707 PAD.n5706 0.019716
R51886 PAD.n5707 PAD.n5562 0.019716
R51887 PAD.n5702 PAD.n5561 0.019716
R51888 PAD.n6690 PAD.n5902 0.019716
R51889 PAD.n6497 PAD.n6397 0.019716
R51890 PAD.n6497 PAD.n5906 0.019716
R51891 PAD.n6502 PAD.n6398 0.019716
R51892 PAD.n6502 PAD.n5907 0.019716
R51893 PAD.n6506 PAD.n6399 0.019716
R51894 PAD.n6506 PAD.n5908 0.019716
R51895 PAD.n6511 PAD.n6400 0.019716
R51896 PAD.n6511 PAD.n5909 0.019716
R51897 PAD.n6515 PAD.n6401 0.019716
R51898 PAD.n6515 PAD.n5910 0.019716
R51899 PAD.n6520 PAD.n6402 0.019716
R51900 PAD.n6520 PAD.n5911 0.019716
R51901 PAD.n6524 PAD.n6403 0.019716
R51902 PAD.n6524 PAD.n5912 0.019716
R51903 PAD.n6529 PAD.n6404 0.019716
R51904 PAD.n6529 PAD.n5913 0.019716
R51905 PAD.n6533 PAD.n6405 0.019716
R51906 PAD.n6533 PAD.n5914 0.019716
R51907 PAD.n6538 PAD.n6406 0.019716
R51908 PAD.n6538 PAD.n5915 0.019716
R51909 PAD.n6542 PAD.n6407 0.019716
R51910 PAD.n6542 PAD.n5916 0.019716
R51911 PAD.n6547 PAD.n6408 0.019716
R51912 PAD.n6547 PAD.n5917 0.019716
R51913 PAD.n6551 PAD.n6409 0.019716
R51914 PAD.n6551 PAD.n5918 0.019716
R51915 PAD.n6556 PAD.n6410 0.019716
R51916 PAD.n6556 PAD.n5919 0.019716
R51917 PAD.n6560 PAD.n6411 0.019716
R51918 PAD.n6560 PAD.n5920 0.019716
R51919 PAD.n6565 PAD.n6412 0.019716
R51920 PAD.n6565 PAD.n5921 0.019716
R51921 PAD.n6569 PAD.n6413 0.019716
R51922 PAD.n6569 PAD.n5922 0.019716
R51923 PAD.n6574 PAD.n6414 0.019716
R51924 PAD.n6574 PAD.n5923 0.019716
R51925 PAD.n6578 PAD.n6415 0.019716
R51926 PAD.n6578 PAD.n5924 0.019716
R51927 PAD.n6583 PAD.n6416 0.019716
R51928 PAD.n6583 PAD.n5925 0.019716
R51929 PAD.n6587 PAD.n6417 0.019716
R51930 PAD.n6587 PAD.n5926 0.019716
R51931 PAD.n6592 PAD.n6418 0.019716
R51932 PAD.n6592 PAD.n5927 0.019716
R51933 PAD.n6596 PAD.n6419 0.019716
R51934 PAD.n6596 PAD.n5928 0.019716
R51935 PAD.n6601 PAD.n6420 0.019716
R51936 PAD.n6601 PAD.n5929 0.019716
R51937 PAD.n6605 PAD.n6421 0.019716
R51938 PAD.n6605 PAD.n5930 0.019716
R51939 PAD.n6610 PAD.n6422 0.019716
R51940 PAD.n6610 PAD.n5931 0.019716
R51941 PAD.n6614 PAD.n6423 0.019716
R51942 PAD.n6614 PAD.n5932 0.019716
R51943 PAD.n6619 PAD.n6424 0.019716
R51944 PAD.n6619 PAD.n5933 0.019716
R51945 PAD.n6623 PAD.n6425 0.019716
R51946 PAD.n6623 PAD.n5934 0.019716
R51947 PAD.n6628 PAD.n6426 0.019716
R51948 PAD.n6628 PAD.n5935 0.019716
R51949 PAD.n6632 PAD.n6427 0.019716
R51950 PAD.n6632 PAD.n5936 0.019716
R51951 PAD.n6637 PAD.n6428 0.019716
R51952 PAD.n6637 PAD.n5937 0.019716
R51953 PAD.n6641 PAD.n6429 0.019716
R51954 PAD.n6641 PAD.n5938 0.019716
R51955 PAD.n6646 PAD.n6430 0.019716
R51956 PAD.n6646 PAD.n5939 0.019716
R51957 PAD.n6650 PAD.n6431 0.019716
R51958 PAD.n6650 PAD.n5940 0.019716
R51959 PAD.n6655 PAD.n6432 0.019716
R51960 PAD.n6655 PAD.n5941 0.019716
R51961 PAD.n6659 PAD.n6433 0.019716
R51962 PAD.n6659 PAD.n5942 0.019716
R51963 PAD.n6664 PAD.n6434 0.019716
R51964 PAD.n6664 PAD.n5943 0.019716
R51965 PAD.n6668 PAD.n6435 0.019716
R51966 PAD.n6668 PAD.n5944 0.019716
R51967 PAD.n6677 PAD.n6676 0.019716
R51968 PAD.n6676 PAD.n5945 0.019716
R51969 PAD.n5949 PAD.n5947 0.019716
R51970 PAD.n5949 PAD.n5946 0.019716
R51971 PAD.n9133 PAD.n2882 0.019625
R51972 PAD.n10733 PAD.n10732 0.019625
R51973 PAD.n9719 PAD.n1590 0.0195611
R51974 PAD.n10019 PAD.n1138 0.0195611
R51975 PAD.n9720 PAD.n1591 0.0195611
R51976 PAD.n10018 PAD.n1139 0.0195611
R51977 PAD.n9157 PAD.n9156 0.019175
R51978 PAD.n10709 PAD.n422 0.019175
R51979 PAD.n8459 PAD.n8458 0.0191681
R51980 PAD.n3686 PAD.n3632 0.0191681
R51981 PAD.n6686 PAD.n6685 0.0187751
R51982 PAD.n6684 PAD.n5948 0.0187751
R51983 PAD.n7825 PAD.n7824 0.018725
R51984 PAD.n7523 PAD.n7156 0.0175961
R51985 PAD.n7522 PAD.n7157 0.0175961
R51986 PAD.n6392 PAD.n6391 0.017282
R51987 PAD.n6392 PAD.n5897 0.017282
R51988 PAD.n6695 PAD.n6694 0.017282
R51989 PAD.n6695 PAD.n5544 0.017282
R51990 PAD.n7805 PAD.n5546 0.017282
R51991 PAD.n7054 PAD.n5546 0.017282
R51992 PAD.n7788 PAD.n7787 0.017282
R51993 PAD.n7787 PAD.n7786 0.017282
R51994 PAD.n7212 PAD.n7210 0.017282
R51995 PAD.n7220 PAD.n7210 0.017282
R51996 PAD.n7227 PAD.n7220 0.017282
R51997 PAD.n7227 PAD.n7226 0.017282
R51998 PAD.n7226 PAD.n5209 0.017282
R51999 PAD.n7816 PAD.n5209 0.017282
R52000 PAD.n8169 PAD.n5194 0.017282
R52001 PAD.n8171 PAD.n5180 0.017282
R52002 PAD.n8189 PAD.n5180 0.017282
R52003 PAD.n8191 PAD.n4677 0.017282
R52004 PAD.n8401 PAD.n4677 0.017282
R52005 PAD.n8404 PAD.n8403 0.017282
R52006 PAD.n8404 PAD.n4326 0.017282
R52007 PAD.n8423 PAD.n4326 0.017282
R52008 PAD.n8427 PAD.n8425 0.017282
R52009 PAD.n8427 PAD.n8426 0.017282
R52010 PAD.n8449 PAD.n8448 0.017282
R52011 PAD.n8450 PAD.n8449 0.017282
R52012 PAD.n8475 PAD.n8474 0.017282
R52013 PAD.n8497 PAD.n8496 0.017282
R52014 PAD.n8499 PAD.n8497 0.017282
R52015 PAD.n8499 PAD.n8498 0.017282
R52016 PAD.n8523 PAD.n8522 0.017282
R52017 PAD.n8524 PAD.n8523 0.017282
R52018 PAD.n8836 PAD.n8835 0.017282
R52019 PAD.n9125 PAD.n8836 0.017282
R52020 PAD.n9123 PAD.n2831 0.017282
R52021 PAD.n9146 PAD.n2831 0.017282
R52022 PAD.n9148 PAD.n2484 0.017282
R52023 PAD.n9166 PAD.n2484 0.017282
R52024 PAD.n9170 PAD.n9169 0.017282
R52025 PAD.n9169 PAD.n2137 0.017282
R52026 PAD.n9194 PAD.n9193 0.017282
R52027 PAD.n9193 PAD.n9192 0.017282
R52028 PAD.n2034 PAD.n1933 0.017282
R52029 PAD.n9725 PAD.n1933 0.017282
R52030 PAD.n9729 PAD.n9728 0.017282
R52031 PAD.n9728 PAD.n9727 0.017282
R52032 PAD.n1584 PAD.n1583 0.017282
R52033 PAD.n1583 PAD.n1146 0.017282
R52034 PAD.n10011 PAD.n1146 0.017282
R52035 PAD.n10013 PAD.n1125 0.017282
R52036 PAD.n10365 PAD.n1125 0.017282
R52037 PAD.n10370 PAD.n10368 0.017282
R52038 PAD.n10370 PAD.n10369 0.017282
R52039 PAD.n10393 PAD.n10392 0.017282
R52040 PAD.n10394 PAD.n10393 0.017282
R52041 PAD.n10412 PAD.n10411 0.017282
R52042 PAD.n10698 PAD.n10412 0.017282
R52043 PAD.n10722 PAD.n370 0.017282
R52044 PAD.n10723 PAD.n10722 0.017282
R52045 PAD.n10724 PAD.n10723 0.017282
R52046 PAD.n11537 PAD.n15 0.017282
R52047 PAD.n10746 PAD.n15 0.017282
R52048 PAD.n11519 PAD.n11089 0.017282
R52049 PAD.n11519 PAD.n11518 0.017282
R52050 PAD.n2897 PAD.n2883 0.0172031
R52051 PAD.n29 PAD.n24 0.0172031
R52052 PAD.n2895 PAD.n2878 0.0172031
R52053 PAD.n31 PAD.n22 0.0172031
R52054 PAD.n8437 PAD.n4315 0.016925
R52055 PAD.n9158 PAD.n2489 0.01681
R52056 PAD.n10705 PAD.n10704 0.01681
R52057 PAD.n9159 PAD.n2488 0.01681
R52058 PAD.n10703 PAD.n417 0.01681
R52059 PAD.n8522 PAD.n2949 0.0167406
R52060 PAD.n10698 PAD.n10697 0.0167406
R52061 PAD.n9738 PAD.n1486 0.016475
R52062 PAD.n10002 PAD.n1486 0.016475
R52063 PAD.n11518 PAD.n11517 0.0164699
R52064 PAD.n7826 PAD.n5199 0.016417
R52065 PAD.n7827 PAD.n5198 0.016417
R52066 PAD.n9167 PAD.n9166 0.0161992
R52067 PAD.n10013 PAD.n10012 0.0161992
R52068 PAD.n8437 PAD.n8436 0.016025
R52069 PAD.n6694 PAD.n6693 0.0156579
R52070 PAD.n8402 PAD.n8401 0.0156579
R52071 PAD.n6393 PAD.n5955 0.0154799
R52072 PAD.n6394 PAD.n6393 0.0154799
R52073 PAD.n6696 PAD.n5896 0.0154799
R52074 PAD.n6697 PAD.n6696 0.0154799
R52075 PAD.n7804 PAD.n5548 0.0154799
R52076 PAD.n7053 PAD.n5548 0.0154799
R52077 PAD.n7789 PAD.n6717 0.0154799
R52078 PAD.n7785 PAD.n6717 0.0154799
R52079 PAD.n7213 PAD.n7211 0.0154799
R52080 PAD.n7219 PAD.n7211 0.0154799
R52081 PAD.n7219 PAD.n7208 0.0154799
R52082 PAD.n7225 PAD.n7208 0.0154799
R52083 PAD.n7225 PAD.n5207 0.0154799
R52084 PAD.n7817 PAD.n5207 0.0154799
R52085 PAD.n7813 PAD.n5195 0.0154799
R52086 PAD.n8168 PAD.n5195 0.0154799
R52087 PAD.n8172 PAD.n5181 0.0154799
R52088 PAD.n8188 PAD.n5181 0.0154799
R52089 PAD.n8192 PAD.n4678 0.0154799
R52090 PAD.n8400 PAD.n4678 0.0154799
R52091 PAD.n8405 PAD.n4675 0.0154799
R52092 PAD.n8405 PAD.n4327 0.0154799
R52093 PAD.n8422 PAD.n4327 0.0154799
R52094 PAD.n8428 PAD.n4323 0.0154799
R52095 PAD.n8428 PAD.n4324 0.0154799
R52096 PAD.n8447 PAD.n3979 0.0154799
R52097 PAD.n8451 PAD.n3979 0.0154799
R52098 PAD.n8471 PAD.n3635 0.0154799
R52099 PAD.n8476 PAD.n3635 0.0154799
R52100 PAD.n8495 PAD.n3291 0.0154799
R52101 PAD.n8500 PAD.n3291 0.0154799
R52102 PAD.n8500 PAD.n3292 0.0154799
R52103 PAD.n8521 PAD.n2948 0.0154799
R52104 PAD.n8525 PAD.n2948 0.0154799
R52105 PAD.n8834 PAD.n2886 0.0154799
R52106 PAD.n9126 PAD.n2886 0.0154799
R52107 PAD.n9122 PAD.n2832 0.0154799
R52108 PAD.n9145 PAD.n2832 0.0154799
R52109 PAD.n9149 PAD.n2485 0.0154799
R52110 PAD.n9165 PAD.n2485 0.0154799
R52111 PAD.n9173 PAD.n2149 0.0154799
R52112 PAD.n2149 PAD.n2136 0.0154799
R52113 PAD.n9191 PAD.n2136 0.0154799
R52114 PAD.n9195 PAD.n2036 0.0154799
R52115 PAD.n2036 PAD.n2033 0.0154799
R52116 PAD.n9461 PAD.n1934 0.0154799
R52117 PAD.n9724 PAD.n1934 0.0154799
R52118 PAD.n9730 PAD.n1597 0.0154799
R52119 PAD.n1597 PAD.n1581 0.0154799
R52120 PAD.n9747 PAD.n1582 0.0154799
R52121 PAD.n1582 PAD.n1147 0.0154799
R52122 PAD.n10010 PAD.n1147 0.0154799
R52123 PAD.n10014 PAD.n1126 0.0154799
R52124 PAD.n10364 PAD.n1126 0.0154799
R52125 PAD.n10371 PAD.n1122 0.0154799
R52126 PAD.n10371 PAD.n1123 0.0154799
R52127 PAD.n10391 PAD.n778 0.0154799
R52128 PAD.n10395 PAD.n778 0.0154799
R52129 PAD.n10410 PAD.n428 0.0154799
R52130 PAD.n10699 PAD.n428 0.0154799
R52131 PAD.n10721 PAD.n371 0.0154799
R52132 PAD.n10721 PAD.n369 0.0154799
R52133 PAD.n10725 PAD.n369 0.0154799
R52134 PAD.n11536 PAD.n17 0.0154799
R52135 PAD.n10751 PAD.n17 0.0154799
R52136 PAD.n11520 PAD.n10744 0.0154799
R52137 PAD.n11520 PAD.n10745 0.0154799
R52138 PAD.n5970 PAD.n5954 0.0154799
R52139 PAD.n6395 PAD.n5954 0.0154799
R52140 PAD.n6681 PAD.n5895 0.0154799
R52141 PAD.n6698 PAD.n5895 0.0154799
R52142 PAD.n7803 PAD.n5550 0.0154799
R52143 PAD.n7052 PAD.n5550 0.0154799
R52144 PAD.n7790 PAD.n6715 0.0154799
R52145 PAD.n7784 PAD.n6715 0.0154799
R52146 PAD.n7217 PAD.n7214 0.0154799
R52147 PAD.n7218 PAD.n7217 0.0154799
R52148 PAD.n7218 PAD.n7202 0.0154799
R52149 PAD.n7224 PAD.n7202 0.0154799
R52150 PAD.n7224 PAD.n5205 0.0154799
R52151 PAD.n7818 PAD.n5205 0.0154799
R52152 PAD.n8166 PAD.n5196 0.0154799
R52153 PAD.n8167 PAD.n8166 0.0154799
R52154 PAD.n8173 PAD.n5182 0.0154799
R52155 PAD.n8187 PAD.n5182 0.0154799
R52156 PAD.n8193 PAD.n4680 0.0154799
R52157 PAD.n8399 PAD.n4680 0.0154799
R52158 PAD.n8406 PAD.n4674 0.0154799
R52159 PAD.n8406 PAD.n4329 0.0154799
R52160 PAD.n8421 PAD.n4329 0.0154799
R52161 PAD.n8429 PAD.n4320 0.0154799
R52162 PAD.n8429 PAD.n4322 0.0154799
R52163 PAD.n8446 PAD.n3978 0.0154799
R52164 PAD.n8452 PAD.n3978 0.0154799
R52165 PAD.n8470 PAD.n3634 0.0154799
R52166 PAD.n8477 PAD.n3634 0.0154799
R52167 PAD.n8494 PAD.n3288 0.0154799
R52168 PAD.n8501 PAD.n3288 0.0154799
R52169 PAD.n8501 PAD.n3290 0.0154799
R52170 PAD.n8520 PAD.n2947 0.0154799
R52171 PAD.n8526 PAD.n2947 0.0154799
R52172 PAD.n8833 PAD.n2884 0.0154799
R52173 PAD.n9127 PAD.n2884 0.0154799
R52174 PAD.n9121 PAD.n2833 0.0154799
R52175 PAD.n9144 PAD.n2833 0.0154799
R52176 PAD.n9150 PAD.n2486 0.0154799
R52177 PAD.n9164 PAD.n2486 0.0154799
R52178 PAD.n9174 PAD.n2138 0.0154799
R52179 PAD.n9188 PAD.n2138 0.0154799
R52180 PAD.n9190 PAD.n9188 0.0154799
R52181 PAD.n9457 PAD.n2035 0.0154799
R52182 PAD.n9458 PAD.n9457 0.0154799
R52183 PAD.n9460 PAD.n1935 0.0154799
R52184 PAD.n9723 PAD.n1935 0.0154799
R52185 PAD.n9731 PAD.n1585 0.0154799
R52186 PAD.n9743 PAD.n1585 0.0154799
R52187 PAD.n9746 PAD.n9745 0.0154799
R52188 PAD.n9745 PAD.n1148 0.0154799
R52189 PAD.n10009 PAD.n1148 0.0154799
R52190 PAD.n10015 PAD.n1128 0.0154799
R52191 PAD.n10363 PAD.n1128 0.0154799
R52192 PAD.n10372 PAD.n1119 0.0154799
R52193 PAD.n10372 PAD.n1121 0.0154799
R52194 PAD.n10390 PAD.n777 0.0154799
R52195 PAD.n10396 PAD.n777 0.0154799
R52196 PAD.n10409 PAD.n426 0.0154799
R52197 PAD.n10700 PAD.n426 0.0154799
R52198 PAD.n10720 PAD.n372 0.0154799
R52199 PAD.n10720 PAD.n368 0.0154799
R52200 PAD.n10726 PAD.n368 0.0154799
R52201 PAD.n11535 PAD.n19 0.0154799
R52202 PAD.n10752 PAD.n19 0.0154799
R52203 PAD.n11521 PAD.n10742 0.0154799
R52204 PAD.n11521 PAD.n10743 0.0154799
R52205 PAD.n8425 PAD.n8424 0.0151165
R52206 PAD.n8521 PAD.n2950 0.0149966
R52207 PAD.n10699 PAD.n429 0.0149966
R52208 PAD.n8520 PAD.n2951 0.0149966
R52209 PAD.n10700 PAD.n427 0.0149966
R52210 PAD.n8434 PAD.n8433 0.014845
R52211 PAD.n8432 PAD.n4027 0.014845
R52212 PAD.n11092 PAD.n10745 0.014755
R52213 PAD.n11094 PAD.n10743 0.014755
R52214 PAD.n9194 PAD.n2135 0.0145752
R52215 PAD.n9727 PAD.n1580 0.0145752
R52216 PAD.n9165 PAD.n2148 0.0145134
R52217 PAD.n10014 PAD.n1144 0.0145134
R52218 PAD.n9164 PAD.n2147 0.0145134
R52219 PAD.n10015 PAD.n1143 0.0145134
R52220 PAD.n9739 PAD.n1487 0.014452
R52221 PAD.n10001 PAD.n1487 0.014452
R52222 PAD.n9740 PAD.n1488 0.014452
R52223 PAD.n10000 PAD.n1488 0.014452
R52224 PAD.n11515 PAD.n11093 0.01445
R52225 PAD.n11354 PAD.n11353 0.01445
R52226 PAD.n11354 PAD.n11351 0.01445
R52227 PAD.n11358 PAD.n11351 0.01445
R52228 PAD.n11359 PAD.n11358 0.01445
R52229 PAD.n11360 PAD.n11359 0.01445
R52230 PAD.n11360 PAD.n11349 0.01445
R52231 PAD.n11364 PAD.n11349 0.01445
R52232 PAD.n11365 PAD.n11364 0.01445
R52233 PAD.n11366 PAD.n11365 0.01445
R52234 PAD.n11366 PAD.n11347 0.01445
R52235 PAD.n11370 PAD.n11347 0.01445
R52236 PAD.n11371 PAD.n11370 0.01445
R52237 PAD.n11372 PAD.n11371 0.01445
R52238 PAD.n11372 PAD.n11345 0.01445
R52239 PAD.n11376 PAD.n11345 0.01445
R52240 PAD.n11377 PAD.n11376 0.01445
R52241 PAD.n11378 PAD.n11377 0.01445
R52242 PAD.n11378 PAD.n11343 0.01445
R52243 PAD.n11382 PAD.n11343 0.01445
R52244 PAD.n11383 PAD.n11382 0.01445
R52245 PAD.n11384 PAD.n11383 0.01445
R52246 PAD.n11384 PAD.n11341 0.01445
R52247 PAD.n11388 PAD.n11341 0.01445
R52248 PAD.n11389 PAD.n11388 0.01445
R52249 PAD.n11390 PAD.n11389 0.01445
R52250 PAD.n11390 PAD.n11339 0.01445
R52251 PAD.n11394 PAD.n11339 0.01445
R52252 PAD.n11395 PAD.n11394 0.01445
R52253 PAD.n11396 PAD.n11395 0.01445
R52254 PAD.n11396 PAD.n11337 0.01445
R52255 PAD.n11400 PAD.n11337 0.01445
R52256 PAD.n11401 PAD.n11400 0.01445
R52257 PAD.n11402 PAD.n11401 0.01445
R52258 PAD.n11402 PAD.n11335 0.01445
R52259 PAD.n11406 PAD.n11335 0.01445
R52260 PAD.n11407 PAD.n11406 0.01445
R52261 PAD.n11408 PAD.n11407 0.01445
R52262 PAD.n11408 PAD.n11333 0.01445
R52263 PAD.n11412 PAD.n11333 0.01445
R52264 PAD.n11413 PAD.n11412 0.01445
R52265 PAD.n11414 PAD.n11413 0.01445
R52266 PAD.n11414 PAD.n11331 0.01445
R52267 PAD.n11418 PAD.n11331 0.01445
R52268 PAD.n11419 PAD.n11418 0.01445
R52269 PAD.n11420 PAD.n11419 0.01445
R52270 PAD.n11420 PAD.n11329 0.01445
R52271 PAD.n11424 PAD.n11329 0.01445
R52272 PAD.n11425 PAD.n11424 0.01445
R52273 PAD.n11426 PAD.n11425 0.01445
R52274 PAD.n11426 PAD.n11327 0.01445
R52275 PAD.n11430 PAD.n11327 0.01445
R52276 PAD.n11431 PAD.n11430 0.01445
R52277 PAD.n11432 PAD.n11431 0.01445
R52278 PAD.n11432 PAD.n11325 0.01445
R52279 PAD.n11436 PAD.n11325 0.01445
R52280 PAD.n11437 PAD.n11436 0.01445
R52281 PAD.n11438 PAD.n11437 0.01445
R52282 PAD.n11438 PAD.n11323 0.01445
R52283 PAD.n11442 PAD.n11323 0.01445
R52284 PAD.n11443 PAD.n11442 0.01445
R52285 PAD.n11444 PAD.n11443 0.01445
R52286 PAD.n11444 PAD.n11321 0.01445
R52287 PAD.n11448 PAD.n11321 0.01445
R52288 PAD.n11449 PAD.n11448 0.01445
R52289 PAD.n11450 PAD.n11449 0.01445
R52290 PAD.n11450 PAD.n11319 0.01445
R52291 PAD.n11454 PAD.n11319 0.01445
R52292 PAD.n11455 PAD.n11454 0.01445
R52293 PAD.n11456 PAD.n11455 0.01445
R52294 PAD.n11456 PAD.n11317 0.01445
R52295 PAD.n11460 PAD.n11317 0.01445
R52296 PAD.n11461 PAD.n11460 0.01445
R52297 PAD.n11462 PAD.n11461 0.01445
R52298 PAD.n11462 PAD.n11315 0.01445
R52299 PAD.n11466 PAD.n11315 0.01445
R52300 PAD.n11467 PAD.n11466 0.01445
R52301 PAD.n11468 PAD.n11467 0.01445
R52302 PAD.n11468 PAD.n11313 0.01445
R52303 PAD.n11472 PAD.n11313 0.01445
R52304 PAD.n11473 PAD.n11472 0.01445
R52305 PAD.n11474 PAD.n11473 0.01445
R52306 PAD.n11474 PAD.n11311 0.01445
R52307 PAD.n11478 PAD.n11311 0.01445
R52308 PAD.n11479 PAD.n11478 0.01445
R52309 PAD.n11480 PAD.n11479 0.01445
R52310 PAD.n11480 PAD.n11309 0.01445
R52311 PAD.n11484 PAD.n11309 0.01445
R52312 PAD.n11485 PAD.n11484 0.01445
R52313 PAD.n11486 PAD.n11485 0.01445
R52314 PAD.n11486 PAD.n11307 0.01445
R52315 PAD.n11490 PAD.n11307 0.01445
R52316 PAD.n11491 PAD.n11490 0.01445
R52317 PAD.n11492 PAD.n11491 0.01445
R52318 PAD.n11492 PAD.n11305 0.01445
R52319 PAD.n11496 PAD.n11305 0.01445
R52320 PAD.n11497 PAD.n11496 0.01445
R52321 PAD.n11498 PAD.n11497 0.01445
R52322 PAD.n11516 PAD.n11091 0.01445
R52323 PAD.n11355 PAD.n11352 0.01445
R52324 PAD.n11356 PAD.n11355 0.01445
R52325 PAD.n11357 PAD.n11356 0.01445
R52326 PAD.n11357 PAD.n11350 0.01445
R52327 PAD.n11361 PAD.n11350 0.01445
R52328 PAD.n11362 PAD.n11361 0.01445
R52329 PAD.n11363 PAD.n11362 0.01445
R52330 PAD.n11363 PAD.n11348 0.01445
R52331 PAD.n11367 PAD.n11348 0.01445
R52332 PAD.n11368 PAD.n11367 0.01445
R52333 PAD.n11369 PAD.n11368 0.01445
R52334 PAD.n11369 PAD.n11346 0.01445
R52335 PAD.n11373 PAD.n11346 0.01445
R52336 PAD.n11374 PAD.n11373 0.01445
R52337 PAD.n11375 PAD.n11374 0.01445
R52338 PAD.n11375 PAD.n11344 0.01445
R52339 PAD.n11379 PAD.n11344 0.01445
R52340 PAD.n11380 PAD.n11379 0.01445
R52341 PAD.n11381 PAD.n11380 0.01445
R52342 PAD.n11381 PAD.n11342 0.01445
R52343 PAD.n11385 PAD.n11342 0.01445
R52344 PAD.n11386 PAD.n11385 0.01445
R52345 PAD.n11387 PAD.n11386 0.01445
R52346 PAD.n11387 PAD.n11340 0.01445
R52347 PAD.n11391 PAD.n11340 0.01445
R52348 PAD.n11392 PAD.n11391 0.01445
R52349 PAD.n11393 PAD.n11392 0.01445
R52350 PAD.n11393 PAD.n11338 0.01445
R52351 PAD.n11397 PAD.n11338 0.01445
R52352 PAD.n11398 PAD.n11397 0.01445
R52353 PAD.n11399 PAD.n11398 0.01445
R52354 PAD.n11399 PAD.n11336 0.01445
R52355 PAD.n11403 PAD.n11336 0.01445
R52356 PAD.n11404 PAD.n11403 0.01445
R52357 PAD.n11405 PAD.n11404 0.01445
R52358 PAD.n11405 PAD.n11334 0.01445
R52359 PAD.n11409 PAD.n11334 0.01445
R52360 PAD.n11410 PAD.n11409 0.01445
R52361 PAD.n11411 PAD.n11410 0.01445
R52362 PAD.n11411 PAD.n11332 0.01445
R52363 PAD.n11415 PAD.n11332 0.01445
R52364 PAD.n11416 PAD.n11415 0.01445
R52365 PAD.n11417 PAD.n11416 0.01445
R52366 PAD.n11417 PAD.n11330 0.01445
R52367 PAD.n11421 PAD.n11330 0.01445
R52368 PAD.n11422 PAD.n11421 0.01445
R52369 PAD.n11423 PAD.n11422 0.01445
R52370 PAD.n11423 PAD.n11328 0.01445
R52371 PAD.n11427 PAD.n11328 0.01445
R52372 PAD.n11428 PAD.n11427 0.01445
R52373 PAD.n11429 PAD.n11428 0.01445
R52374 PAD.n11429 PAD.n11326 0.01445
R52375 PAD.n11433 PAD.n11326 0.01445
R52376 PAD.n11434 PAD.n11433 0.01445
R52377 PAD.n11435 PAD.n11434 0.01445
R52378 PAD.n11435 PAD.n11324 0.01445
R52379 PAD.n11439 PAD.n11324 0.01445
R52380 PAD.n11440 PAD.n11439 0.01445
R52381 PAD.n11441 PAD.n11440 0.01445
R52382 PAD.n11441 PAD.n11322 0.01445
R52383 PAD.n11445 PAD.n11322 0.01445
R52384 PAD.n11446 PAD.n11445 0.01445
R52385 PAD.n11447 PAD.n11446 0.01445
R52386 PAD.n11447 PAD.n11320 0.01445
R52387 PAD.n11451 PAD.n11320 0.01445
R52388 PAD.n11452 PAD.n11451 0.01445
R52389 PAD.n11453 PAD.n11452 0.01445
R52390 PAD.n11453 PAD.n11318 0.01445
R52391 PAD.n11457 PAD.n11318 0.01445
R52392 PAD.n11458 PAD.n11457 0.01445
R52393 PAD.n11459 PAD.n11458 0.01445
R52394 PAD.n11459 PAD.n11316 0.01445
R52395 PAD.n11463 PAD.n11316 0.01445
R52396 PAD.n11464 PAD.n11463 0.01445
R52397 PAD.n11465 PAD.n11464 0.01445
R52398 PAD.n11465 PAD.n11314 0.01445
R52399 PAD.n11469 PAD.n11314 0.01445
R52400 PAD.n11470 PAD.n11469 0.01445
R52401 PAD.n11471 PAD.n11470 0.01445
R52402 PAD.n11471 PAD.n11312 0.01445
R52403 PAD.n11475 PAD.n11312 0.01445
R52404 PAD.n11476 PAD.n11475 0.01445
R52405 PAD.n11477 PAD.n11476 0.01445
R52406 PAD.n11477 PAD.n11310 0.01445
R52407 PAD.n11481 PAD.n11310 0.01445
R52408 PAD.n11482 PAD.n11481 0.01445
R52409 PAD.n11483 PAD.n11482 0.01445
R52410 PAD.n11483 PAD.n11308 0.01445
R52411 PAD.n11487 PAD.n11308 0.01445
R52412 PAD.n11488 PAD.n11487 0.01445
R52413 PAD.n11489 PAD.n11488 0.01445
R52414 PAD.n11489 PAD.n11306 0.01445
R52415 PAD.n11493 PAD.n11306 0.01445
R52416 PAD.n11494 PAD.n11493 0.01445
R52417 PAD.n11495 PAD.n11494 0.01445
R52418 PAD.n11495 PAD.n11304 0.01445
R52419 PAD.n11499 PAD.n11304 0.01445
R52420 PAD.n6388 PAD.n5959 0.01445
R52421 PAD.n6227 PAD.n6226 0.01445
R52422 PAD.n6228 PAD.n6227 0.01445
R52423 PAD.n6228 PAD.n6223 0.01445
R52424 PAD.n6232 PAD.n6223 0.01445
R52425 PAD.n6233 PAD.n6232 0.01445
R52426 PAD.n6234 PAD.n6233 0.01445
R52427 PAD.n6234 PAD.n6221 0.01445
R52428 PAD.n6238 PAD.n6221 0.01445
R52429 PAD.n6239 PAD.n6238 0.01445
R52430 PAD.n6240 PAD.n6239 0.01445
R52431 PAD.n6240 PAD.n6219 0.01445
R52432 PAD.n6244 PAD.n6219 0.01445
R52433 PAD.n6245 PAD.n6244 0.01445
R52434 PAD.n6246 PAD.n6245 0.01445
R52435 PAD.n6246 PAD.n6217 0.01445
R52436 PAD.n6250 PAD.n6217 0.01445
R52437 PAD.n6251 PAD.n6250 0.01445
R52438 PAD.n6252 PAD.n6251 0.01445
R52439 PAD.n6252 PAD.n6215 0.01445
R52440 PAD.n6256 PAD.n6215 0.01445
R52441 PAD.n6257 PAD.n6256 0.01445
R52442 PAD.n6258 PAD.n6257 0.01445
R52443 PAD.n6258 PAD.n6213 0.01445
R52444 PAD.n6262 PAD.n6213 0.01445
R52445 PAD.n6263 PAD.n6262 0.01445
R52446 PAD.n6264 PAD.n6263 0.01445
R52447 PAD.n6264 PAD.n6211 0.01445
R52448 PAD.n6268 PAD.n6211 0.01445
R52449 PAD.n6269 PAD.n6268 0.01445
R52450 PAD.n6270 PAD.n6269 0.01445
R52451 PAD.n6270 PAD.n6209 0.01445
R52452 PAD.n6274 PAD.n6209 0.01445
R52453 PAD.n6275 PAD.n6274 0.01445
R52454 PAD.n6276 PAD.n6275 0.01445
R52455 PAD.n6276 PAD.n6207 0.01445
R52456 PAD.n6280 PAD.n6207 0.01445
R52457 PAD.n6281 PAD.n6280 0.01445
R52458 PAD.n6282 PAD.n6281 0.01445
R52459 PAD.n6282 PAD.n6205 0.01445
R52460 PAD.n6286 PAD.n6205 0.01445
R52461 PAD.n6287 PAD.n6286 0.01445
R52462 PAD.n6288 PAD.n6287 0.01445
R52463 PAD.n6288 PAD.n6203 0.01445
R52464 PAD.n6292 PAD.n6203 0.01445
R52465 PAD.n6293 PAD.n6292 0.01445
R52466 PAD.n6294 PAD.n6293 0.01445
R52467 PAD.n6294 PAD.n6201 0.01445
R52468 PAD.n6298 PAD.n6201 0.01445
R52469 PAD.n6299 PAD.n6298 0.01445
R52470 PAD.n6300 PAD.n6299 0.01445
R52471 PAD.n6300 PAD.n6199 0.01445
R52472 PAD.n6304 PAD.n6199 0.01445
R52473 PAD.n6305 PAD.n6304 0.01445
R52474 PAD.n6306 PAD.n6305 0.01445
R52475 PAD.n6306 PAD.n6197 0.01445
R52476 PAD.n6310 PAD.n6197 0.01445
R52477 PAD.n6311 PAD.n6310 0.01445
R52478 PAD.n6312 PAD.n6311 0.01445
R52479 PAD.n6312 PAD.n6195 0.01445
R52480 PAD.n6316 PAD.n6195 0.01445
R52481 PAD.n6317 PAD.n6316 0.01445
R52482 PAD.n6318 PAD.n6317 0.01445
R52483 PAD.n6318 PAD.n6193 0.01445
R52484 PAD.n6322 PAD.n6193 0.01445
R52485 PAD.n6323 PAD.n6322 0.01445
R52486 PAD.n6324 PAD.n6323 0.01445
R52487 PAD.n6324 PAD.n6191 0.01445
R52488 PAD.n6328 PAD.n6191 0.01445
R52489 PAD.n6329 PAD.n6328 0.01445
R52490 PAD.n6330 PAD.n6329 0.01445
R52491 PAD.n6330 PAD.n6189 0.01445
R52492 PAD.n6334 PAD.n6189 0.01445
R52493 PAD.n6335 PAD.n6334 0.01445
R52494 PAD.n6336 PAD.n6335 0.01445
R52495 PAD.n6336 PAD.n6187 0.01445
R52496 PAD.n6340 PAD.n6187 0.01445
R52497 PAD.n6341 PAD.n6340 0.01445
R52498 PAD.n6342 PAD.n6341 0.01445
R52499 PAD.n6342 PAD.n6185 0.01445
R52500 PAD.n6346 PAD.n6185 0.01445
R52501 PAD.n6347 PAD.n6346 0.01445
R52502 PAD.n6348 PAD.n6347 0.01445
R52503 PAD.n6348 PAD.n6183 0.01445
R52504 PAD.n6352 PAD.n6183 0.01445
R52505 PAD.n6353 PAD.n6352 0.01445
R52506 PAD.n6354 PAD.n6353 0.01445
R52507 PAD.n6354 PAD.n6181 0.01445
R52508 PAD.n6358 PAD.n6181 0.01445
R52509 PAD.n6359 PAD.n6358 0.01445
R52510 PAD.n6360 PAD.n6359 0.01445
R52511 PAD.n6360 PAD.n6179 0.01445
R52512 PAD.n6364 PAD.n6179 0.01445
R52513 PAD.n6365 PAD.n6364 0.01445
R52514 PAD.n6366 PAD.n6365 0.01445
R52515 PAD.n6366 PAD.n6177 0.01445
R52516 PAD.n6370 PAD.n6177 0.01445
R52517 PAD.n6371 PAD.n6370 0.01445
R52518 PAD.n6389 PAD.n5957 0.01445
R52519 PAD.n6225 PAD.n6224 0.01445
R52520 PAD.n6229 PAD.n6224 0.01445
R52521 PAD.n6230 PAD.n6229 0.01445
R52522 PAD.n6231 PAD.n6230 0.01445
R52523 PAD.n6231 PAD.n6222 0.01445
R52524 PAD.n6235 PAD.n6222 0.01445
R52525 PAD.n6236 PAD.n6235 0.01445
R52526 PAD.n6237 PAD.n6236 0.01445
R52527 PAD.n6237 PAD.n6220 0.01445
R52528 PAD.n6241 PAD.n6220 0.01445
R52529 PAD.n6242 PAD.n6241 0.01445
R52530 PAD.n6243 PAD.n6242 0.01445
R52531 PAD.n6243 PAD.n6218 0.01445
R52532 PAD.n6247 PAD.n6218 0.01445
R52533 PAD.n6248 PAD.n6247 0.01445
R52534 PAD.n6249 PAD.n6248 0.01445
R52535 PAD.n6249 PAD.n6216 0.01445
R52536 PAD.n6253 PAD.n6216 0.01445
R52537 PAD.n6254 PAD.n6253 0.01445
R52538 PAD.n6255 PAD.n6254 0.01445
R52539 PAD.n6255 PAD.n6214 0.01445
R52540 PAD.n6259 PAD.n6214 0.01445
R52541 PAD.n6260 PAD.n6259 0.01445
R52542 PAD.n6261 PAD.n6260 0.01445
R52543 PAD.n6261 PAD.n6212 0.01445
R52544 PAD.n6265 PAD.n6212 0.01445
R52545 PAD.n6266 PAD.n6265 0.01445
R52546 PAD.n6267 PAD.n6266 0.01445
R52547 PAD.n6267 PAD.n6210 0.01445
R52548 PAD.n6271 PAD.n6210 0.01445
R52549 PAD.n6272 PAD.n6271 0.01445
R52550 PAD.n6273 PAD.n6272 0.01445
R52551 PAD.n6273 PAD.n6208 0.01445
R52552 PAD.n6277 PAD.n6208 0.01445
R52553 PAD.n6278 PAD.n6277 0.01445
R52554 PAD.n6279 PAD.n6278 0.01445
R52555 PAD.n6279 PAD.n6206 0.01445
R52556 PAD.n6283 PAD.n6206 0.01445
R52557 PAD.n6284 PAD.n6283 0.01445
R52558 PAD.n6285 PAD.n6284 0.01445
R52559 PAD.n6285 PAD.n6204 0.01445
R52560 PAD.n6289 PAD.n6204 0.01445
R52561 PAD.n6290 PAD.n6289 0.01445
R52562 PAD.n6291 PAD.n6290 0.01445
R52563 PAD.n6291 PAD.n6202 0.01445
R52564 PAD.n6295 PAD.n6202 0.01445
R52565 PAD.n6296 PAD.n6295 0.01445
R52566 PAD.n6297 PAD.n6296 0.01445
R52567 PAD.n6297 PAD.n6200 0.01445
R52568 PAD.n6301 PAD.n6200 0.01445
R52569 PAD.n6302 PAD.n6301 0.01445
R52570 PAD.n6303 PAD.n6302 0.01445
R52571 PAD.n6303 PAD.n6198 0.01445
R52572 PAD.n6307 PAD.n6198 0.01445
R52573 PAD.n6308 PAD.n6307 0.01445
R52574 PAD.n6309 PAD.n6308 0.01445
R52575 PAD.n6309 PAD.n6196 0.01445
R52576 PAD.n6313 PAD.n6196 0.01445
R52577 PAD.n6314 PAD.n6313 0.01445
R52578 PAD.n6315 PAD.n6314 0.01445
R52579 PAD.n6315 PAD.n6194 0.01445
R52580 PAD.n6319 PAD.n6194 0.01445
R52581 PAD.n6320 PAD.n6319 0.01445
R52582 PAD.n6321 PAD.n6320 0.01445
R52583 PAD.n6321 PAD.n6192 0.01445
R52584 PAD.n6325 PAD.n6192 0.01445
R52585 PAD.n6326 PAD.n6325 0.01445
R52586 PAD.n6327 PAD.n6326 0.01445
R52587 PAD.n6327 PAD.n6190 0.01445
R52588 PAD.n6331 PAD.n6190 0.01445
R52589 PAD.n6332 PAD.n6331 0.01445
R52590 PAD.n6333 PAD.n6332 0.01445
R52591 PAD.n6333 PAD.n6188 0.01445
R52592 PAD.n6337 PAD.n6188 0.01445
R52593 PAD.n6338 PAD.n6337 0.01445
R52594 PAD.n6339 PAD.n6338 0.01445
R52595 PAD.n6339 PAD.n6186 0.01445
R52596 PAD.n6343 PAD.n6186 0.01445
R52597 PAD.n6344 PAD.n6343 0.01445
R52598 PAD.n6345 PAD.n6344 0.01445
R52599 PAD.n6345 PAD.n6184 0.01445
R52600 PAD.n6349 PAD.n6184 0.01445
R52601 PAD.n6350 PAD.n6349 0.01445
R52602 PAD.n6351 PAD.n6350 0.01445
R52603 PAD.n6351 PAD.n6182 0.01445
R52604 PAD.n6355 PAD.n6182 0.01445
R52605 PAD.n6356 PAD.n6355 0.01445
R52606 PAD.n6357 PAD.n6356 0.01445
R52607 PAD.n6357 PAD.n6180 0.01445
R52608 PAD.n6361 PAD.n6180 0.01445
R52609 PAD.n6362 PAD.n6361 0.01445
R52610 PAD.n6363 PAD.n6362 0.01445
R52611 PAD.n6363 PAD.n6178 0.01445
R52612 PAD.n6367 PAD.n6178 0.01445
R52613 PAD.n6368 PAD.n6367 0.01445
R52614 PAD.n6369 PAD.n6368 0.01445
R52615 PAD.n6369 PAD.n5978 0.01445
R52616 PAD.n6391 PAD.n6390 0.0143045
R52617 PAD.n7824 PAD.n7823 0.014225
R52618 PAD.n8435 PAD.n8434 0.014059
R52619 PAD.n4027 PAD.n3976 0.014059
R52620 PAD.n8475 PAD.n3293 0.0140338
R52621 PAD.n5899 PAD.n5896 0.0140302
R52622 PAD.n8400 PAD.n4679 0.0140302
R52623 PAD.n6681 PAD.n5901 0.0140302
R52624 PAD.n8399 PAD.n4681 0.0140302
R52625 PAD.n9156 PAD.n9155 0.013775
R52626 PAD.n10709 PAD.n10708 0.013775
R52627 PAD.n9171 PAD.n9170 0.0137632
R52628 PAD.n4328 PAD.n4323 0.013547
R52629 PAD.n4330 PAD.n4320 0.013547
R52630 PAD.n7786 PAD.n7056 0.0134925
R52631 PAD.n7815 PAD.n7814 0.0134925
R52632 PAD.n9133 PAD.n9132 0.013325
R52633 PAD.n10732 PAD.n10731 0.013325
R52634 PAD.n9196 PAD.n9195 0.0130638
R52635 PAD.n9748 PAD.n1581 0.0130638
R52636 PAD.n9189 PAD.n2035 0.0130638
R52637 PAD.n9744 PAD.n9743 0.0130638
R52638 PAD.n8835 PAD.n2888 0.0129511
R52639 PAD.n10394 PAD.n430 0.0129511
R52640 PAD.n7203 PAD.n7155 0.012875
R52641 PAD.n5958 PAD.n5955 0.0128221
R52642 PAD.n5970 PAD.n5960 0.0128221
R52643 PAD.n8474 PAD.n8473 0.0128158
R52644 PAD.n8476 PAD.n3294 0.0125805
R52645 PAD.n11536 PAD.n16 0.0125805
R52646 PAD.n8477 PAD.n3295 0.0125805
R52647 PAD.n11535 PAD.n18 0.0125805
R52648 PAD.n7822 PAD.n5199 0.0124869
R52649 PAD.n7821 PAD.n5198 0.0124869
R52650 PAD.n9147 PAD.n9146 0.0124098
R52651 PAD.n10368 PAD.n10367 0.0124098
R52652 PAD.n11538 PAD.n14 0.0124098
R52653 PAD.n11102 PAD.n11094 0.0123125
R52654 PAD.n11101 PAD.n11092 0.0123125
R52655 PAD.n5967 PAD.n5958 0.0123125
R52656 PAD.n5968 PAD.n5960 0.0123125
R52657 PAD.n7785 PAD.n7057 0.0120973
R52658 PAD.n7813 PAD.n5208 0.0120973
R52659 PAD.n7784 PAD.n7058 0.0120973
R52660 PAD.n5206 PAD.n5196 0.0120973
R52661 PAD.n9154 PAD.n2489 0.0120939
R52662 PAD.n10707 PAD.n10705 0.0120939
R52663 PAD.n9153 PAD.n2488 0.0120939
R52664 PAD.n10706 PAD.n417 0.0120939
R52665 PAD.n11505 PAD.n11499 0.011975
R52666 PAD.n6376 PAD.n5978 0.011975
R52667 PAD.n7806 PAD.n7805 0.0118684
R52668 PAD.n8190 PAD.n8189 0.0118684
R52669 PAD.n9131 PAD.n2883 0.0117009
R52670 PAD.n10730 PAD.n29 0.0117009
R52671 PAD.n9130 PAD.n2878 0.0117009
R52672 PAD.n10729 PAD.n31 0.0117009
R52673 PAD.n8834 PAD.n2889 0.0116141
R52674 PAD.n10395 PAD.n431 0.0116141
R52675 PAD.n8833 PAD.n2890 0.0116141
R52676 PAD.n10396 PAD.n432 0.0116141
R52677 PAD.n7812 PAD.n5194 0.0115977
R52678 PAD.n6378 PAD.n6377 0.011525
R52679 PAD.n8448 PAD.n3980 0.0113271
R52680 PAD.n7204 PAD.n7156 0.0113079
R52681 PAD.n7205 PAD.n7157 0.0113079
R52682 PAD.n9145 PAD.n2496 0.0111309
R52683 PAD.n1127 PAD.n1122 0.0111309
R52684 PAD.n9144 PAD.n2495 0.0111309
R52685 PAD.n1129 PAD.n1119 0.0111309
R52686 PAD.n8461 PAD.n3974 0.011075
R52687 PAD.n2034 PAD.n2032 0.0107857
R52688 PAD.n9726 PAD.n9725 0.0107857
R52689 PAD.n7804 PAD.n5547 0.0106477
R52690 PAD.n8188 PAD.n4845 0.0106477
R52691 PAD.n7803 PAD.n5549 0.0106477
R52692 PAD.n8187 PAD.n4844 0.0106477
R52693 PAD.n9736 PAD.n1589 0.010625
R52694 PAD.n10004 PAD.n1137 0.010625
R52695 PAD.n74 PAD.n18 0.0105588
R52696 PAD.n366 PAD.n31 0.0105588
R52697 PAD.n7518 PAD.n7202 0.0105588
R52698 PAD.n7269 PAD.n7157 0.0105588
R52699 PAD.n7517 PAD.n7208 0.0105588
R52700 PAD.n7270 PAD.n7156 0.0105588
R52701 PAD.n427 PAD.n415 0.0105588
R52702 PAD.n10715 PAD.n417 0.0105588
R52703 PAD.n10695 PAD.n429 0.0105588
R52704 PAD.n10705 PAD.n416 0.0105588
R52705 PAD.n523 PAD.n432 0.0105588
R52706 PAD.n770 PAD.n436 0.0105588
R52707 PAD.n522 PAD.n431 0.0105588
R52708 PAD.n771 PAD.n437 0.0105588
R52709 PAD.n824 PAD.n781 0.0105588
R52710 PAD.n10387 PAD.n827 0.0105588
R52711 PAD.n872 PAD.n780 0.0105588
R52712 PAD.n10377 PAD.n826 0.0105588
R52713 PAD.n10106 PAD.n1129 0.0105588
R52714 PAD.n10353 PAD.n1134 0.0105588
R52715 PAD.n10105 PAD.n1127 0.0105588
R52716 PAD.n10354 PAD.n1136 0.0105588
R52717 PAD.n1481 PAD.n1143 0.0105588
R52718 PAD.n1294 PAD.n1139 0.0105588
R52719 PAD.n1480 PAD.n1144 0.0105588
R52720 PAD.n1295 PAD.n1138 0.0105588
R52721 PAD.n9744 PAD.n1531 0.0105588
R52722 PAD.n9997 PAD.n1488 0.0105588
R52723 PAD.n9749 PAD.n9748 0.0105588
R52724 PAD.n1535 PAD.n1487 0.0105588
R52725 PAD.n1599 PAD.n1595 0.0105588
R52726 PAD.n1685 PAD.n1591 0.0105588
R52727 PAD.n1931 PAD.n1596 0.0105588
R52728 PAD.n1684 PAD.n1590 0.0105588
R52729 PAD.n9459 PAD.n1984 0.0105588
R52730 PAD.n9711 PAD.n1941 0.0105588
R52731 PAD.n9463 PAD.n9462 0.0105588
R52732 PAD.n1987 PAD.n1940 0.0105588
R52733 PAD.n9189 PAD.n2088 0.0105588
R52734 PAD.n9444 PAD.n2045 0.0105588
R52735 PAD.n9197 PAD.n9196 0.0105588
R52736 PAD.n2090 PAD.n2043 0.0105588
R52737 PAD.n2151 PAD.n2147 0.0105588
R52738 PAD.n2236 PAD.n2140 0.0105588
R52739 PAD.n2482 PAD.n2148 0.0105588
R52740 PAD.n2235 PAD.n2141 0.0105588
R52741 PAD.n2498 PAD.n2495 0.0105588
R52742 PAD.n2583 PAD.n2488 0.0105588
R52743 PAD.n2829 PAD.n2496 0.0105588
R52744 PAD.n2582 PAD.n2489 0.0105588
R52745 PAD.n2885 PAD.n2876 0.0105588
R52746 PAD.n9139 PAD.n2878 0.0105588
R52747 PAD.n9119 PAD.n2887 0.0105588
R52748 PAD.n2883 PAD.n2877 0.0105588
R52749 PAD.n8819 PAD.n2890 0.0105588
R52750 PAD.n8570 PAD.n2903 0.0105588
R52751 PAD.n8818 PAD.n2889 0.0105588
R52752 PAD.n8571 PAD.n2901 0.0105588
R52753 PAD.n2994 PAD.n2951 0.0105588
R52754 PAD.n8516 PAD.n2996 0.0105588
R52755 PAD.n3041 PAD.n2950 0.0105588
R52756 PAD.n8506 PAD.n2995 0.0105588
R52757 PAD.n3338 PAD.n3295 0.0105588
R52758 PAD.n8491 PAD.n3341 0.0105588
R52759 PAD.n3386 PAD.n3294 0.0105588
R52760 PAD.n3631 PAD.n3340 0.0105588
R52761 PAD.n3683 PAD.n3640 0.0105588
R52762 PAD.n8467 PAD.n3686 0.0105588
R52763 PAD.n3731 PAD.n3639 0.0105588
R52764 PAD.n8458 PAD.n3685 0.0105588
R52765 PAD.n4025 PAD.n3982 0.0105588
R52766 PAD.n8443 PAD.n4027 0.0105588
R52767 PAD.n4072 PAD.n3981 0.0105588
R52768 PAD.n8434 PAD.n4026 0.0105588
R52769 PAD.n4420 PAD.n4330 0.0105588
R52770 PAD.n4667 PAD.n4334 0.0105588
R52771 PAD.n4419 PAD.n4328 0.0105588
R52772 PAD.n4668 PAD.n4335 0.0105588
R52773 PAD.n8395 PAD.n4681 0.0105588
R52774 PAD.n8204 PAD.n4832 0.0105588
R52775 PAD.n8394 PAD.n4679 0.0105588
R52776 PAD.n4831 PAD.n4829 0.0105588
R52777 PAD.n4847 PAD.n4844 0.0105588
R52778 PAD.n4932 PAD.n4839 0.0105588
R52779 PAD.n5178 PAD.n4845 0.0105588
R52780 PAD.n4931 PAD.n4834 0.0105588
R52781 PAD.n8161 PAD.n5191 0.0105588
R52782 PAD.n7971 PAD.n5184 0.0105588
R52783 PAD.n8160 PAD.n5192 0.0105588
R52784 PAD.n7972 PAD.n5185 0.0105588
R52785 PAD.n5211 PAD.n5206 0.0105588
R52786 PAD.n5296 PAD.n5198 0.0105588
R52787 PAD.n5542 PAD.n5208 0.0105588
R52788 PAD.n5295 PAD.n5199 0.0105588
R52789 PAD.n7780 PAD.n7058 0.0105588
R52790 PAD.n7531 PAD.n7530 0.0105588
R52791 PAD.n7779 PAD.n7057 0.0105588
R52792 PAD.n7532 PAD.n7148 0.0105588
R52793 PAD.n6719 PAD.n6714 0.0105588
R52794 PAD.n6804 PAD.n6709 0.0105588
R52795 PAD.n7050 PAD.n6716 0.0105588
R52796 PAD.n6803 PAD.n6707 0.0105588
R52797 PAD.n5892 PAD.n5549 0.0105588
R52798 PAD.n5702 PAD.n5553 0.0105588
R52799 PAD.n5891 PAD.n5547 0.0105588
R52800 PAD.n5703 PAD.n5555 0.0105588
R52801 PAD.n6691 PAD.n5899 0.0105588
R52802 PAD.n6687 PAD.n6686 0.0105588
R52803 PAD.n119 PAD.n16 0.0105588
R52804 PAD.n75 PAD.n29 0.0105588
R52805 PAD.n11086 PAD.n10748 0.0105588
R52806 PAD.n10838 PAD.n10736 0.0105588
R52807 PAD.n11085 PAD.n10750 0.0105588
R52808 PAD.n10837 PAD.n10738 0.0105588
R52809 PAD.n6690 PAD.n5901 0.0105588
R52810 PAD.n6688 PAD.n5948 0.0105588
R52811 PAD.n8450 PAD.n3638 0.0102444
R52812 PAD.n11089 PAD.n11088 0.0102444
R52813 PAD.n8416 PAD.n8414 0.010175
R52814 PAD.n11505 PAD.n11504 0.010175
R52815 PAD.n8447 PAD.n3981 0.0101644
R52816 PAD.n8446 PAD.n3982 0.0101644
R52817 PAD.n6686 PAD.n5952 0.0101288
R52818 PAD.n5973 PAD.n5948 0.0101288
R52819 PAD.n8458 PAD.n8457 0.00973581
R52820 PAD.n8456 PAD.n3686 0.00973581
R52821 PAD.n7055 PAD.n7054 0.00970301
R52822 PAD.n8171 PAD.n8170 0.00970301
R52823 PAD.n11101 PAD.n11090 0.00969267
R52824 PAD.n9462 PAD.n9461 0.00968121
R52825 PAD.n9724 PAD.n1596 0.00968121
R52826 PAD.n9460 PAD.n9459 0.00968121
R52827 PAD.n9723 PAD.n1595 0.00968121
R52828 PAD.n9735 PAD.n1590 0.00934279
R52829 PAD.n10005 PAD.n1138 0.00934279
R52830 PAD.n9734 PAD.n1591 0.00934279
R52831 PAD.n10006 PAD.n1139 0.00934279
R52832 PAD.n8451 PAD.n3639 0.00919799
R52833 PAD.n10748 PAD.n10744 0.00919799
R52834 PAD.n8452 PAD.n3640 0.00919799
R52835 PAD.n10750 PAD.n10742 0.00919799
R52836 PAD.n9124 PAD.n9123 0.00916165
R52837 PAD.n10369 PAD.n779 0.00916165
R52838 PAD.n8417 PAD.n4335 0.00894978
R52839 PAD.n11503 PAD.n11303 0.00894978
R52840 PAD.n8418 PAD.n4334 0.00894978
R52841 PAD.n11502 PAD.n11253 0.00894978
R52842 PAD.n7053 PAD.n6716 0.00871477
R52843 PAD.n8172 PAD.n5192 0.00871477
R52844 PAD.n7052 PAD.n6714 0.00871477
R52845 PAD.n8173 PAD.n5191 0.00871477
R52846 PAD.n11253 PAD.n11156 0.0087125
R52847 PAD.n11498 PAD.n11303 0.0087125
R52848 PAD.n6371 PAD.n5976 0.0087125
R52849 PAD.n6372 PAD.n5972 0.0087125
R52850 PAD.n9125 PAD.n9124 0.0086203
R52851 PAD.n10392 PAD.n779 0.0086203
R52852 PAD.n8179 PAD.n8178 0.008375
R52853 PAD.n9122 PAD.n2887 0.00823154
R52854 PAD.n1123 PAD.n780 0.00823154
R52855 PAD.n9121 PAD.n2885 0.00823154
R52856 PAD.n1121 PAD.n781 0.00823154
R52857 PAD.n5967 PAD.n5956 0.00813094
R52858 PAD.n9168 PAD.n11 0.00808277
R52859 PAD.n7788 PAD.n7055 0.00807895
R52860 PAD.n8170 PAD.n8169 0.00807895
R52861 PAD.n11511 PAD.n11102 0.00796421
R52862 PAD.n11104 PAD.n11095 0.00796421
R52863 PAD.n11301 PAD.n11252 0.00796421
R52864 PAD.n11251 PAD.n11107 0.00796421
R52865 PAD.n11300 PAD.n11250 0.00796421
R52866 PAD.n11249 PAD.n11108 0.00796421
R52867 PAD.n11299 PAD.n11248 0.00796421
R52868 PAD.n11247 PAD.n11109 0.00796421
R52869 PAD.n11298 PAD.n11246 0.00796421
R52870 PAD.n11245 PAD.n11110 0.00796421
R52871 PAD.n11297 PAD.n11244 0.00796421
R52872 PAD.n11243 PAD.n11111 0.00796421
R52873 PAD.n11296 PAD.n11242 0.00796421
R52874 PAD.n11241 PAD.n11112 0.00796421
R52875 PAD.n11295 PAD.n11240 0.00796421
R52876 PAD.n11239 PAD.n11113 0.00796421
R52877 PAD.n11294 PAD.n11238 0.00796421
R52878 PAD.n11237 PAD.n11114 0.00796421
R52879 PAD.n11293 PAD.n11236 0.00796421
R52880 PAD.n11235 PAD.n11115 0.00796421
R52881 PAD.n11292 PAD.n11234 0.00796421
R52882 PAD.n11233 PAD.n11116 0.00796421
R52883 PAD.n11291 PAD.n11232 0.00796421
R52884 PAD.n11231 PAD.n11117 0.00796421
R52885 PAD.n11290 PAD.n11230 0.00796421
R52886 PAD.n11229 PAD.n11118 0.00796421
R52887 PAD.n11289 PAD.n11228 0.00796421
R52888 PAD.n11227 PAD.n11119 0.00796421
R52889 PAD.n11288 PAD.n11226 0.00796421
R52890 PAD.n11225 PAD.n11120 0.00796421
R52891 PAD.n11287 PAD.n11224 0.00796421
R52892 PAD.n11223 PAD.n11121 0.00796421
R52893 PAD.n11286 PAD.n11222 0.00796421
R52894 PAD.n11221 PAD.n11122 0.00796421
R52895 PAD.n11285 PAD.n11220 0.00796421
R52896 PAD.n11219 PAD.n11123 0.00796421
R52897 PAD.n11284 PAD.n11218 0.00796421
R52898 PAD.n11217 PAD.n11124 0.00796421
R52899 PAD.n11283 PAD.n11216 0.00796421
R52900 PAD.n11215 PAD.n11125 0.00796421
R52901 PAD.n11282 PAD.n11214 0.00796421
R52902 PAD.n11213 PAD.n11126 0.00796421
R52903 PAD.n11281 PAD.n11212 0.00796421
R52904 PAD.n11211 PAD.n11127 0.00796421
R52905 PAD.n11280 PAD.n11210 0.00796421
R52906 PAD.n11209 PAD.n11128 0.00796421
R52907 PAD.n11279 PAD.n11208 0.00796421
R52908 PAD.n11207 PAD.n11129 0.00796421
R52909 PAD.n11278 PAD.n11206 0.00796421
R52910 PAD.n11205 PAD.n11130 0.00796421
R52911 PAD.n11277 PAD.n11204 0.00796421
R52912 PAD.n11203 PAD.n11131 0.00796421
R52913 PAD.n11276 PAD.n11202 0.00796421
R52914 PAD.n11201 PAD.n11132 0.00796421
R52915 PAD.n11275 PAD.n11200 0.00796421
R52916 PAD.n11199 PAD.n11133 0.00796421
R52917 PAD.n11274 PAD.n11198 0.00796421
R52918 PAD.n11197 PAD.n11134 0.00796421
R52919 PAD.n11273 PAD.n11196 0.00796421
R52920 PAD.n11195 PAD.n11135 0.00796421
R52921 PAD.n11272 PAD.n11194 0.00796421
R52922 PAD.n11193 PAD.n11136 0.00796421
R52923 PAD.n11271 PAD.n11192 0.00796421
R52924 PAD.n11191 PAD.n11137 0.00796421
R52925 PAD.n11270 PAD.n11190 0.00796421
R52926 PAD.n11189 PAD.n11138 0.00796421
R52927 PAD.n11269 PAD.n11188 0.00796421
R52928 PAD.n11187 PAD.n11139 0.00796421
R52929 PAD.n11268 PAD.n11186 0.00796421
R52930 PAD.n11185 PAD.n11140 0.00796421
R52931 PAD.n11267 PAD.n11184 0.00796421
R52932 PAD.n11183 PAD.n11141 0.00796421
R52933 PAD.n11266 PAD.n11182 0.00796421
R52934 PAD.n11181 PAD.n11142 0.00796421
R52935 PAD.n11265 PAD.n11180 0.00796421
R52936 PAD.n11179 PAD.n11143 0.00796421
R52937 PAD.n11264 PAD.n11178 0.00796421
R52938 PAD.n11177 PAD.n11144 0.00796421
R52939 PAD.n11263 PAD.n11176 0.00796421
R52940 PAD.n11175 PAD.n11145 0.00796421
R52941 PAD.n11262 PAD.n11174 0.00796421
R52942 PAD.n11173 PAD.n11146 0.00796421
R52943 PAD.n11261 PAD.n11172 0.00796421
R52944 PAD.n11171 PAD.n11147 0.00796421
R52945 PAD.n11260 PAD.n11170 0.00796421
R52946 PAD.n11169 PAD.n11148 0.00796421
R52947 PAD.n11259 PAD.n11168 0.00796421
R52948 PAD.n11167 PAD.n11149 0.00796421
R52949 PAD.n11258 PAD.n11166 0.00796421
R52950 PAD.n11165 PAD.n11150 0.00796421
R52951 PAD.n11257 PAD.n11164 0.00796421
R52952 PAD.n11163 PAD.n11151 0.00796421
R52953 PAD.n11256 PAD.n11162 0.00796421
R52954 PAD.n11161 PAD.n11152 0.00796421
R52955 PAD.n11255 PAD.n11160 0.00796421
R52956 PAD.n11159 PAD.n11153 0.00796421
R52957 PAD.n11254 PAD.n11158 0.00796421
R52958 PAD.n11157 PAD.n11154 0.00796421
R52959 PAD.n11156 PAD.n11155 0.00796421
R52960 PAD.n6384 PAD.n5968 0.00796421
R52961 PAD.n5969 PAD.n5961 0.00796421
R52962 PAD.n6033 PAD.n6030 0.00796421
R52963 PAD.n6037 PAD.n6035 0.00796421
R52964 PAD.n6036 PAD.n6029 0.00796421
R52965 PAD.n6040 PAD.n6038 0.00796421
R52966 PAD.n6039 PAD.n6028 0.00796421
R52967 PAD.n6043 PAD.n6041 0.00796421
R52968 PAD.n6042 PAD.n6027 0.00796421
R52969 PAD.n6046 PAD.n6044 0.00796421
R52970 PAD.n6045 PAD.n6026 0.00796421
R52971 PAD.n6049 PAD.n6047 0.00796421
R52972 PAD.n6048 PAD.n6025 0.00796421
R52973 PAD.n6052 PAD.n6050 0.00796421
R52974 PAD.n6051 PAD.n6024 0.00796421
R52975 PAD.n6055 PAD.n6053 0.00796421
R52976 PAD.n6054 PAD.n6023 0.00796421
R52977 PAD.n6058 PAD.n6056 0.00796421
R52978 PAD.n6057 PAD.n6022 0.00796421
R52979 PAD.n6061 PAD.n6059 0.00796421
R52980 PAD.n6060 PAD.n6021 0.00796421
R52981 PAD.n6064 PAD.n6062 0.00796421
R52982 PAD.n6063 PAD.n6020 0.00796421
R52983 PAD.n6067 PAD.n6065 0.00796421
R52984 PAD.n6066 PAD.n6019 0.00796421
R52985 PAD.n6070 PAD.n6068 0.00796421
R52986 PAD.n6069 PAD.n6018 0.00796421
R52987 PAD.n6073 PAD.n6071 0.00796421
R52988 PAD.n6072 PAD.n6017 0.00796421
R52989 PAD.n6076 PAD.n6074 0.00796421
R52990 PAD.n6075 PAD.n6016 0.00796421
R52991 PAD.n6079 PAD.n6077 0.00796421
R52992 PAD.n6078 PAD.n6015 0.00796421
R52993 PAD.n6082 PAD.n6080 0.00796421
R52994 PAD.n6081 PAD.n6014 0.00796421
R52995 PAD.n6085 PAD.n6083 0.00796421
R52996 PAD.n6084 PAD.n6013 0.00796421
R52997 PAD.n6088 PAD.n6086 0.00796421
R52998 PAD.n6087 PAD.n6012 0.00796421
R52999 PAD.n6091 PAD.n6089 0.00796421
R53000 PAD.n6090 PAD.n6011 0.00796421
R53001 PAD.n6094 PAD.n6092 0.00796421
R53002 PAD.n6093 PAD.n6010 0.00796421
R53003 PAD.n6097 PAD.n6095 0.00796421
R53004 PAD.n6096 PAD.n6009 0.00796421
R53005 PAD.n6100 PAD.n6098 0.00796421
R53006 PAD.n6099 PAD.n6008 0.00796421
R53007 PAD.n6103 PAD.n6101 0.00796421
R53008 PAD.n6102 PAD.n6007 0.00796421
R53009 PAD.n6106 PAD.n6104 0.00796421
R53010 PAD.n6105 PAD.n6006 0.00796421
R53011 PAD.n6109 PAD.n6107 0.00796421
R53012 PAD.n6108 PAD.n6005 0.00796421
R53013 PAD.n6112 PAD.n6110 0.00796421
R53014 PAD.n6111 PAD.n6004 0.00796421
R53015 PAD.n6115 PAD.n6113 0.00796421
R53016 PAD.n6114 PAD.n6003 0.00796421
R53017 PAD.n6118 PAD.n6116 0.00796421
R53018 PAD.n6117 PAD.n6002 0.00796421
R53019 PAD.n6121 PAD.n6119 0.00796421
R53020 PAD.n6120 PAD.n6001 0.00796421
R53021 PAD.n6124 PAD.n6122 0.00796421
R53022 PAD.n6123 PAD.n6000 0.00796421
R53023 PAD.n6127 PAD.n6125 0.00796421
R53024 PAD.n6126 PAD.n5999 0.00796421
R53025 PAD.n6130 PAD.n6128 0.00796421
R53026 PAD.n6129 PAD.n5998 0.00796421
R53027 PAD.n6133 PAD.n6131 0.00796421
R53028 PAD.n6132 PAD.n5997 0.00796421
R53029 PAD.n6136 PAD.n6134 0.00796421
R53030 PAD.n6135 PAD.n5996 0.00796421
R53031 PAD.n6139 PAD.n6137 0.00796421
R53032 PAD.n6138 PAD.n5995 0.00796421
R53033 PAD.n6142 PAD.n6140 0.00796421
R53034 PAD.n6141 PAD.n5994 0.00796421
R53035 PAD.n6145 PAD.n6143 0.00796421
R53036 PAD.n6144 PAD.n5993 0.00796421
R53037 PAD.n6148 PAD.n6146 0.00796421
R53038 PAD.n6147 PAD.n5992 0.00796421
R53039 PAD.n6151 PAD.n6149 0.00796421
R53040 PAD.n6150 PAD.n5991 0.00796421
R53041 PAD.n6154 PAD.n6152 0.00796421
R53042 PAD.n6153 PAD.n5990 0.00796421
R53043 PAD.n6157 PAD.n6155 0.00796421
R53044 PAD.n6156 PAD.n5989 0.00796421
R53045 PAD.n6160 PAD.n6158 0.00796421
R53046 PAD.n6159 PAD.n5988 0.00796421
R53047 PAD.n6163 PAD.n6161 0.00796421
R53048 PAD.n6162 PAD.n5987 0.00796421
R53049 PAD.n6166 PAD.n6164 0.00796421
R53050 PAD.n6165 PAD.n5986 0.00796421
R53051 PAD.n6169 PAD.n6167 0.00796421
R53052 PAD.n6168 PAD.n5985 0.00796421
R53053 PAD.n6172 PAD.n6170 0.00796421
R53054 PAD.n6171 PAD.n5984 0.00796421
R53055 PAD.n6175 PAD.n6173 0.00796421
R53056 PAD.n6174 PAD.n5983 0.00796421
R53057 PAD.n6032 PAD.n6031 0.00796421
R53058 PAD.n6372 PAD.n6176 0.00796421
R53059 PAD.n6176 PAD.n6032 0.00796421
R53060 PAD.n11155 PAD.n11154 0.00796421
R53061 PAD.n11158 PAD.n11157 0.00796421
R53062 PAD.n11254 PAD.n11153 0.00796421
R53063 PAD.n11160 PAD.n11159 0.00796421
R53064 PAD.n11255 PAD.n11152 0.00796421
R53065 PAD.n11162 PAD.n11161 0.00796421
R53066 PAD.n11256 PAD.n11151 0.00796421
R53067 PAD.n11164 PAD.n11163 0.00796421
R53068 PAD.n11257 PAD.n11150 0.00796421
R53069 PAD.n11166 PAD.n11165 0.00796421
R53070 PAD.n11258 PAD.n11149 0.00796421
R53071 PAD.n11168 PAD.n11167 0.00796421
R53072 PAD.n11259 PAD.n11148 0.00796421
R53073 PAD.n11170 PAD.n11169 0.00796421
R53074 PAD.n11260 PAD.n11147 0.00796421
R53075 PAD.n11172 PAD.n11171 0.00796421
R53076 PAD.n11261 PAD.n11146 0.00796421
R53077 PAD.n11174 PAD.n11173 0.00796421
R53078 PAD.n11262 PAD.n11145 0.00796421
R53079 PAD.n11176 PAD.n11175 0.00796421
R53080 PAD.n11263 PAD.n11144 0.00796421
R53081 PAD.n11178 PAD.n11177 0.00796421
R53082 PAD.n11264 PAD.n11143 0.00796421
R53083 PAD.n11180 PAD.n11179 0.00796421
R53084 PAD.n11265 PAD.n11142 0.00796421
R53085 PAD.n11182 PAD.n11181 0.00796421
R53086 PAD.n11266 PAD.n11141 0.00796421
R53087 PAD.n11184 PAD.n11183 0.00796421
R53088 PAD.n11267 PAD.n11140 0.00796421
R53089 PAD.n11186 PAD.n11185 0.00796421
R53090 PAD.n11268 PAD.n11139 0.00796421
R53091 PAD.n11188 PAD.n11187 0.00796421
R53092 PAD.n11269 PAD.n11138 0.00796421
R53093 PAD.n11190 PAD.n11189 0.00796421
R53094 PAD.n11270 PAD.n11137 0.00796421
R53095 PAD.n11192 PAD.n11191 0.00796421
R53096 PAD.n11271 PAD.n11136 0.00796421
R53097 PAD.n11194 PAD.n11193 0.00796421
R53098 PAD.n11272 PAD.n11135 0.00796421
R53099 PAD.n11196 PAD.n11195 0.00796421
R53100 PAD.n11273 PAD.n11134 0.00796421
R53101 PAD.n11198 PAD.n11197 0.00796421
R53102 PAD.n11274 PAD.n11133 0.00796421
R53103 PAD.n11200 PAD.n11199 0.00796421
R53104 PAD.n11275 PAD.n11132 0.00796421
R53105 PAD.n11202 PAD.n11201 0.00796421
R53106 PAD.n11276 PAD.n11131 0.00796421
R53107 PAD.n11204 PAD.n11203 0.00796421
R53108 PAD.n11277 PAD.n11130 0.00796421
R53109 PAD.n11206 PAD.n11205 0.00796421
R53110 PAD.n11278 PAD.n11129 0.00796421
R53111 PAD.n11208 PAD.n11207 0.00796421
R53112 PAD.n11279 PAD.n11128 0.00796421
R53113 PAD.n11210 PAD.n11209 0.00796421
R53114 PAD.n11280 PAD.n11127 0.00796421
R53115 PAD.n11212 PAD.n11211 0.00796421
R53116 PAD.n11281 PAD.n11126 0.00796421
R53117 PAD.n11214 PAD.n11213 0.00796421
R53118 PAD.n11282 PAD.n11125 0.00796421
R53119 PAD.n11216 PAD.n11215 0.00796421
R53120 PAD.n11283 PAD.n11124 0.00796421
R53121 PAD.n11218 PAD.n11217 0.00796421
R53122 PAD.n11284 PAD.n11123 0.00796421
R53123 PAD.n11220 PAD.n11219 0.00796421
R53124 PAD.n11285 PAD.n11122 0.00796421
R53125 PAD.n11222 PAD.n11221 0.00796421
R53126 PAD.n11286 PAD.n11121 0.00796421
R53127 PAD.n11224 PAD.n11223 0.00796421
R53128 PAD.n11287 PAD.n11120 0.00796421
R53129 PAD.n11226 PAD.n11225 0.00796421
R53130 PAD.n11288 PAD.n11119 0.00796421
R53131 PAD.n11228 PAD.n11227 0.00796421
R53132 PAD.n11289 PAD.n11118 0.00796421
R53133 PAD.n11230 PAD.n11229 0.00796421
R53134 PAD.n11290 PAD.n11117 0.00796421
R53135 PAD.n11232 PAD.n11231 0.00796421
R53136 PAD.n11291 PAD.n11116 0.00796421
R53137 PAD.n11234 PAD.n11233 0.00796421
R53138 PAD.n11292 PAD.n11115 0.00796421
R53139 PAD.n11236 PAD.n11235 0.00796421
R53140 PAD.n11293 PAD.n11114 0.00796421
R53141 PAD.n11238 PAD.n11237 0.00796421
R53142 PAD.n11294 PAD.n11113 0.00796421
R53143 PAD.n11240 PAD.n11239 0.00796421
R53144 PAD.n11295 PAD.n11112 0.00796421
R53145 PAD.n11242 PAD.n11241 0.00796421
R53146 PAD.n11296 PAD.n11111 0.00796421
R53147 PAD.n11244 PAD.n11243 0.00796421
R53148 PAD.n11297 PAD.n11110 0.00796421
R53149 PAD.n11246 PAD.n11245 0.00796421
R53150 PAD.n11298 PAD.n11109 0.00796421
R53151 PAD.n11248 PAD.n11247 0.00796421
R53152 PAD.n11299 PAD.n11108 0.00796421
R53153 PAD.n11250 PAD.n11249 0.00796421
R53154 PAD.n11300 PAD.n11107 0.00796421
R53155 PAD.n11252 PAD.n11251 0.00796421
R53156 PAD.n11301 PAD.n11106 0.00796421
R53157 PAD.n6387 PAD.n5961 0.00796421
R53158 PAD.n11514 PAD.n11095 0.00796421
R53159 PAD.n6385 PAD.n6384 0.00796421
R53160 PAD.n11512 PAD.n11511 0.00796421
R53161 PAD.n6034 PAD.n6033 0.00796421
R53162 PAD.n6035 PAD.n6030 0.00796421
R53163 PAD.n6037 PAD.n6036 0.00796421
R53164 PAD.n6038 PAD.n6029 0.00796421
R53165 PAD.n6040 PAD.n6039 0.00796421
R53166 PAD.n6041 PAD.n6028 0.00796421
R53167 PAD.n6043 PAD.n6042 0.00796421
R53168 PAD.n6044 PAD.n6027 0.00796421
R53169 PAD.n6046 PAD.n6045 0.00796421
R53170 PAD.n6047 PAD.n6026 0.00796421
R53171 PAD.n6049 PAD.n6048 0.00796421
R53172 PAD.n6050 PAD.n6025 0.00796421
R53173 PAD.n6052 PAD.n6051 0.00796421
R53174 PAD.n6053 PAD.n6024 0.00796421
R53175 PAD.n6055 PAD.n6054 0.00796421
R53176 PAD.n6056 PAD.n6023 0.00796421
R53177 PAD.n6058 PAD.n6057 0.00796421
R53178 PAD.n6059 PAD.n6022 0.00796421
R53179 PAD.n6061 PAD.n6060 0.00796421
R53180 PAD.n6062 PAD.n6021 0.00796421
R53181 PAD.n6064 PAD.n6063 0.00796421
R53182 PAD.n6065 PAD.n6020 0.00796421
R53183 PAD.n6067 PAD.n6066 0.00796421
R53184 PAD.n6068 PAD.n6019 0.00796421
R53185 PAD.n6070 PAD.n6069 0.00796421
R53186 PAD.n6071 PAD.n6018 0.00796421
R53187 PAD.n6073 PAD.n6072 0.00796421
R53188 PAD.n6074 PAD.n6017 0.00796421
R53189 PAD.n6076 PAD.n6075 0.00796421
R53190 PAD.n6077 PAD.n6016 0.00796421
R53191 PAD.n6079 PAD.n6078 0.00796421
R53192 PAD.n6080 PAD.n6015 0.00796421
R53193 PAD.n6082 PAD.n6081 0.00796421
R53194 PAD.n6083 PAD.n6014 0.00796421
R53195 PAD.n6085 PAD.n6084 0.00796421
R53196 PAD.n6086 PAD.n6013 0.00796421
R53197 PAD.n6088 PAD.n6087 0.00796421
R53198 PAD.n6089 PAD.n6012 0.00796421
R53199 PAD.n6091 PAD.n6090 0.00796421
R53200 PAD.n6092 PAD.n6011 0.00796421
R53201 PAD.n6094 PAD.n6093 0.00796421
R53202 PAD.n6095 PAD.n6010 0.00796421
R53203 PAD.n6097 PAD.n6096 0.00796421
R53204 PAD.n6098 PAD.n6009 0.00796421
R53205 PAD.n6100 PAD.n6099 0.00796421
R53206 PAD.n6101 PAD.n6008 0.00796421
R53207 PAD.n6103 PAD.n6102 0.00796421
R53208 PAD.n6104 PAD.n6007 0.00796421
R53209 PAD.n6106 PAD.n6105 0.00796421
R53210 PAD.n6107 PAD.n6006 0.00796421
R53211 PAD.n6109 PAD.n6108 0.00796421
R53212 PAD.n6110 PAD.n6005 0.00796421
R53213 PAD.n6112 PAD.n6111 0.00796421
R53214 PAD.n6113 PAD.n6004 0.00796421
R53215 PAD.n6115 PAD.n6114 0.00796421
R53216 PAD.n6116 PAD.n6003 0.00796421
R53217 PAD.n6118 PAD.n6117 0.00796421
R53218 PAD.n6119 PAD.n6002 0.00796421
R53219 PAD.n6121 PAD.n6120 0.00796421
R53220 PAD.n6122 PAD.n6001 0.00796421
R53221 PAD.n6124 PAD.n6123 0.00796421
R53222 PAD.n6125 PAD.n6000 0.00796421
R53223 PAD.n6127 PAD.n6126 0.00796421
R53224 PAD.n6128 PAD.n5999 0.00796421
R53225 PAD.n6130 PAD.n6129 0.00796421
R53226 PAD.n6131 PAD.n5998 0.00796421
R53227 PAD.n6133 PAD.n6132 0.00796421
R53228 PAD.n6134 PAD.n5997 0.00796421
R53229 PAD.n6136 PAD.n6135 0.00796421
R53230 PAD.n6137 PAD.n5996 0.00796421
R53231 PAD.n6139 PAD.n6138 0.00796421
R53232 PAD.n6140 PAD.n5995 0.00796421
R53233 PAD.n6142 PAD.n6141 0.00796421
R53234 PAD.n6143 PAD.n5994 0.00796421
R53235 PAD.n6145 PAD.n6144 0.00796421
R53236 PAD.n6146 PAD.n5993 0.00796421
R53237 PAD.n6148 PAD.n6147 0.00796421
R53238 PAD.n6149 PAD.n5992 0.00796421
R53239 PAD.n6151 PAD.n6150 0.00796421
R53240 PAD.n6152 PAD.n5991 0.00796421
R53241 PAD.n6154 PAD.n6153 0.00796421
R53242 PAD.n6155 PAD.n5990 0.00796421
R53243 PAD.n6157 PAD.n6156 0.00796421
R53244 PAD.n6158 PAD.n5989 0.00796421
R53245 PAD.n6160 PAD.n6159 0.00796421
R53246 PAD.n6161 PAD.n5988 0.00796421
R53247 PAD.n6163 PAD.n6162 0.00796421
R53248 PAD.n6164 PAD.n5987 0.00796421
R53249 PAD.n6166 PAD.n6165 0.00796421
R53250 PAD.n6167 PAD.n5986 0.00796421
R53251 PAD.n6169 PAD.n6168 0.00796421
R53252 PAD.n6170 PAD.n5985 0.00796421
R53253 PAD.n6172 PAD.n6171 0.00796421
R53254 PAD.n6173 PAD.n5984 0.00796421
R53255 PAD.n6175 PAD.n6174 0.00796421
R53256 PAD.n6031 PAD.n5983 0.00796421
R53257 PAD.n9180 PAD.n9179 0.007925
R53258 PAD.n10404 PAD.n10402 0.007925
R53259 PAD.n9126 PAD.n2887 0.00774832
R53260 PAD.n10391 PAD.n780 0.00774832
R53261 PAD.n9127 PAD.n2885 0.00774832
R53262 PAD.n10390 PAD.n781 0.00774832
R53263 PAD.n8472 PAD.n3638 0.00753759
R53264 PAD.n11088 PAD.n10746 0.00753759
R53265 PAD.n8827 PAD.n8826 0.007475
R53266 PAD.n11528 PAD.n11527 0.007475
R53267 PAD.n8177 PAD.n5185 0.00737773
R53268 PAD.n8176 PAD.n5184 0.00737773
R53269 PAD.n7789 PAD.n6716 0.0072651
R53270 PAD.n8168 PAD.n5192 0.0072651
R53271 PAD.n7790 PAD.n6714 0.0072651
R53272 PAD.n8167 PAD.n5191 0.0072651
R53273 PAD.n11517 PAD.n11516 0.0071375
R53274 PAD.n6390 PAD.n6389 0.0071375
R53275 PAD.n6380 PAD.n6376 0.007025
R53276 PAD.n7526 PAD.n7154 0.007025
R53277 PAD.n9192 PAD.n2032 0.00699624
R53278 PAD.n9729 PAD.n9726 0.00699624
R53279 PAD.n3637 PAD.n3636 0.0069926
R53280 PAD.n9178 PAD.n2141 0.00698472
R53281 PAD.n10405 PAD.n437 0.00698472
R53282 PAD.n9177 PAD.n2140 0.00698472
R53283 PAD.n10406 PAD.n436 0.00698472
R53284 PAD.n8471 PAD.n3639 0.00678188
R53285 PAD.n10751 PAD.n10748 0.00678188
R53286 PAD.n8470 PAD.n3640 0.00678188
R53287 PAD.n10752 PAD.n10750 0.00678188
R53288 PAD.n2901 PAD.n2896 0.0065917
R53289 PAD.n10736 PAD.n25 0.0065917
R53290 PAD.n2903 PAD.n2893 0.0065917
R53291 PAD.n10738 PAD.n23 0.0065917
R53292 PAD.n8426 PAD.n3980 0.00645489
R53293 PAD.n9462 PAD.n2033 0.00629866
R53294 PAD.n9730 PAD.n1596 0.00629866
R53295 PAD.n9459 PAD.n9458 0.00629866
R53296 PAD.n9731 PAD.n1595 0.00629866
R53297 PAD.n11508 PAD.n11253 0.0062375
R53298 PAD.n11506 PAD.n11303 0.0062375
R53299 PAD.n6375 PAD.n5976 0.0062375
R53300 PAD.n6374 PAD.n5972 0.0062375
R53301 PAD.n6381 PAD.n5976 0.00619869
R53302 PAD.n7527 PAD.n7148 0.00619869
R53303 PAD.n6382 PAD.n5972 0.00619869
R53304 PAD.n7530 PAD.n7529 0.00619869
R53305 PAD.n7814 PAD.n7812 0.00618421
R53306 PAD.n8191 PAD.n8190 0.00591353
R53307 PAD.n4324 PAD.n3981 0.00581544
R53308 PAD.n4322 PAD.n3982 0.00581544
R53309 PAD.n6704 PAD.n6703 0.005675
R53310 PAD.n9148 PAD.n9147 0.00537218
R53311 PAD.n6697 PAD.n5547 0.00533221
R53312 PAD.n8192 PAD.n4845 0.00533221
R53313 PAD.n6698 PAD.n5549 0.00533221
R53314 PAD.n8193 PAD.n4844 0.00533221
R53315 PAD.n8485 PAD.n8483 0.005225
R53316 PAD.n6702 PAD.n5555 0.00501965
R53317 PAD.n6701 PAD.n5553 0.00501965
R53318 PAD.n8473 PAD.n8472 0.00496617
R53319 PAD.n9149 PAD.n2496 0.00484899
R53320 PAD.n10364 PAD.n1127 0.00484899
R53321 PAD.n9150 PAD.n2495 0.00484899
R53322 PAD.n10363 PAD.n1129 0.00484899
R53323 PAD.n8524 PAD.n2888 0.00483083
R53324 PAD.n10411 PAD.n430 0.00483083
R53325 PAD.n9716 PAD.n1939 0.004775
R53326 PAD.n10358 PAD.n10357 0.004775
R53327 PAD.n8482 PAD.n3631 0.00462664
R53328 PAD.n8481 PAD.n3341 0.00462664
R53329 PAD.n8525 PAD.n2889 0.00436577
R53330 PAD.n10410 PAD.n431 0.00436577
R53331 PAD.n8526 PAD.n2890 0.00436577
R53332 PAD.n10409 PAD.n432 0.00436577
R53333 PAD.n8209 PAD.n8208 0.004325
R53334 PAD.n7212 PAD.n7056 0.00428947
R53335 PAD.n7816 PAD.n7815 0.00428947
R53336 PAD.n9715 PAD.n1940 0.00423362
R53337 PAD.n10359 PAD.n1136 0.00423362
R53338 PAD.n9714 PAD.n1941 0.00423362
R53339 PAD.n10360 PAD.n1134 0.00423362
R53340 PAD.n9172 PAD.n9171 0.0040188
R53341 PAD.n7213 PAD.n7057 0.00388255
R53342 PAD.n7817 PAD.n5208 0.00388255
R53343 PAD.n7214 PAD.n7058 0.00388255
R53344 PAD.n7818 PAD.n5206 0.00388255
R53345 PAD.n8207 PAD.n4831 0.00384061
R53346 PAD.n8206 PAD.n8204 0.00384061
R53347 PAD.n8496 PAD.n3293 0.00374812
R53348 PAD.n10724 PAD.n14 0.00374812
R53349 PAD.n7807 PAD.n7806 0.00347744
R53350 PAD.n8495 PAD.n3294 0.00339933
R53351 PAD.n10725 PAD.n16 0.00339933
R53352 PAD.n8494 PAD.n3295 0.00339933
R53353 PAD.n10726 PAD.n18 0.00339933
R53354 PAD.n2137 PAD.n2135 0.00320677
R53355 PAD.n1584 PAD.n1580 0.00320677
R53356 PAD.n7807 PAD.n5544 0.00293609
R53357 PAD.n10366 PAD.n10365 0.00293609
R53358 PAD.n10367 PAD.n10366 0.00293609
R53359 PAD.n9196 PAD.n9191 0.00291611
R53360 PAD.n9748 PAD.n9747 0.00291611
R53361 PAD.n9190 PAD.n9189 0.00291611
R53362 PAD.n9746 PAD.n9744 0.00291611
R53363 PAD.n8424 PAD.n8423 0.00266541
R53364 PAD.n11514 PAD.n11094 0.0026375
R53365 PAD.n11515 PAD.n11092 0.0026375
R53366 PAD.n6388 PAD.n5958 0.0026375
R53367 PAD.n6387 PAD.n5960 0.0026375
R53368 PAD.n8199 PAD.n8198 0.002525
R53369 PAD.n8422 PAD.n4328 0.00243289
R53370 PAD.n8421 PAD.n4330 0.00243289
R53371 PAD.n8197 PAD.n4834 0.00226856
R53372 PAD.n8196 PAD.n4839 0.00226856
R53373 PAD.n6693 PAD.n5897 0.00212406
R53374 PAD.n8403 PAD.n8402 0.00212406
R53375 PAD.n11538 PAD.n11537 0.00212406
R53376 PAD.n9450 PAD.n9449 0.002075
R53377 PAD.n10381 PAD.n10380 0.002075
R53378 PAD.n6394 PAD.n5899 0.00194966
R53379 PAD.n4679 PAD.n4675 0.00194966
R53380 PAD.n6395 PAD.n5901 0.00194966
R53381 PAD.n4681 PAD.n4674 0.00194966
R53382 PAD.n9448 PAD.n2043 0.00187555
R53383 PAD.n10379 PAD.n10377 0.00187555
R53384 PAD.n9447 PAD.n2045 0.00187555
R53385 PAD.n10378 PAD.n827 0.00187555
R53386 PAD.n8510 PAD.n8509 0.001625
R53387 PAD.n9172 PAD.n9167 0.00158271
R53388 PAD.n10012 PAD.n10011 0.00158271
R53389 PAD.n8508 PAD.n8506 0.00148253
R53390 PAD.n8507 PAD.n2996 0.00148253
R53391 PAD.n9173 PAD.n2148 0.00146644
R53392 PAD.n10010 PAD.n1144 0.00146644
R53393 PAD.n9174 PAD.n2147 0.00146644
R53394 PAD.n10009 PAD.n1143 0.00146644
R53395 PAD.n11103 PAD.n11097 0.00128471
R53396 PAD.n11103 PAD.n11098 0.00128471
R53397 PAD.n7796 PAD.n7795 0.001175
R53398 PAD.n7794 PAD.n6707 0.00108952
R53399 PAD.n7793 PAD.n6709 0.00108952
R53400 PAD.n6386 PAD.n5966 0.00106946
R53401 PAD.n8165 PAD.n7829 0.00106946
R53402 PAD.n8445 PAD.n3977 0.00106946
R53403 PAD.n11534 PAD.n11533 0.00106946
R53404 PAD.n6682 PAD.n6680 0.00106487
R53405 PAD.n10016 PAD.n1142 0.00106487
R53406 PAD.n9186 PAD.n9185 0.0010465
R53407 PAD.n8498 PAD.n2949 0.00104135
R53408 PAD.n10697 PAD.n370 0.00104135
R53409 PAD.n8454 PAD.n8453 0.00103731
R53410 PAD.n9129 PAD.n9128 0.00103731
R53411 PAD.n5982 PAD.n5963 0.00103272
R53412 PAD.n5981 PAD.n5964 0.00103272
R53413 PAD.n5980 PAD.n5962 0.00103272
R53414 PAD.n5979 PAD.n5965 0.00103272
R53415 PAD.n8503 PAD.n3287 0.00102813
R53416 PAD.n9141 PAD.n9140 0.00102813
R53417 PAD.n4321 PAD.n3983 0.00101894
R53418 PAD.n9143 PAD.n9142 0.00101894
R53419 PAD.n4841 PAD.n4682 0.00100976
R53420 PAD.n9733 PAD.n1592 0.00100517
R53421 PAD.n9742 PAD.n1586 0.00100057
R53422 PAD.n7061 PAD.n7060 0.000991389
R53423 PAD.n8164 PAD.n8163 0.000991389
R53424 PAD.n10398 PAD.n776 0.000991389
R53425 PAD.n3292 PAD.n2950 0.000983221
R53426 PAD.n429 PAD.n371 0.000983221
R53427 PAD.n3290 PAD.n2951 0.000983221
R53428 PAD.n427 PAD.n372 0.000983221
R53429 PAD.n7215 PAD.n7158 0.000982204
R53430 PAD.n10701 PAD.n425 0.000982204
R53431 PAD.n7819 PAD.n5197 0.000977612
R53432 PAD.n8175 PAD.n8174 0.00097302
R53433 PAD.n9721 PAD.n1936 0.00097302
R53434 PAD.n10408 PAD.n433 0.00097302
R53435 PAD.n8409 PAD.n8408 0.000963835
R53436 PAD.n11532 PAD.n21 0.000959242
R53437 PAD.n10755 PAD.n10754 0.000959242
R53438 PAD.n8469 PAD.n3641 0.00095465
R53439 PAD.n2894 PAD.n2892 0.00095465
R53440 PAD.n6700 PAD.n5551 0.000945465
R53441 PAD.n8518 PAD.n2904 0.000945465
R53442 PAD.n6679 PAD.n5894 0.000940873
R53443 PAD.n8431 PAD.n8430 0.00093628
R53444 PAD.n9152 PAD.n9151 0.00093628
R53445 PAD.n1594 PAD.n1593 0.00093628
R53446 PAD.n9456 PAD.n2037 0.000927095
R53447 PAD.n10727 PAD.n367 0.000922503
R53448 PAD.n11507 PAD.n11096 0.000922503
R53449 PAD.n11302 PAD.n11099 0.000922503
R53450 PAD.n11510 PAD.n11509 0.000922503
R53451 PAD.n11513 PAD.n11100 0.000922503
R53452 PAD.n7782 PAD.n7103 0.00091791
R53453 PAD.n7801 PAD.n5552 0.000908726
R53454 PAD.n10361 PAD.n1132 0.000908726
R53455 PAD.n10373 PAD.n1118 0.000908726
R53456 PAD.n1536 PAD.n1489 0.000904133
R53457 PAD.n1141 PAD.n1130 0.000904133
R53458 PAD.n7221 PAD.n5204 0.000894948
R53459 PAD.n8184 PAD.n8183 0.000890356
R53460 PAD.n1986 PAD.n1985 0.000890356
R53461 PAD.n435 PAD.n434 0.000890356
R53462 PAD.n11523 PAD.n11522 0.000890356
R53463 PAD.n10008 PAD.n1140 0.000876579
R53464 PAD.n6678 PAD.n6396 0.000871986
R53465 PAD.n8397 PAD.n4724 0.000871986
R53466 PAD.n3684 PAD.n3633 0.000871986
R53467 PAD.n8832 PAD.n8831 0.000871986
R53468 PAD.n9446 PAD.n9445 0.000862801
R53469 PAD.n419 PAD.n418 0.000858209
R53470 PAD.n4332 PAD.n4319 0.000853617
R53471 PAD.n9161 PAD.n9160 0.000853617
R53472 PAD.n10388 PAD.n825 0.000844432
R53473 PAD.n11501 PAD.n11500 0.000844432
R53474 PAD.n9187 PAD.n2091 0.000839839
R53475 PAD.n10717 PAD.n32 0.000839839
R53476 PAD.n6383 PAD.n5971 0.000835247
R53477 PAD.n7216 PAD.n7105 0.000835247
R53478 PAD.n7223 PAD.n7222 0.000835247
R53479 PAD.n10719 PAD.n10718 0.000835247
R53480 PAD.n6712 PAD.n6711 0.000826062
R53481 PAD.n7792 PAD.n6712 0.000826062
R53482 PAD.n7059 PAD.n6713 0.000826062
R53483 PAD.n1120 PAD.n782 0.000826062
R53484 PAD.n3289 PAD.n2997 0.00082147
R53485 PAD.n9998 PAD.n1534 0.00082147
R53486 PAD.n5974 PAD.n5971 0.000816877
R53487 PAD.n1534 PAD.n1533 0.000816877
R53488 PAD.n8186 PAD.n8185 0.000807692
R53489 PAD.n9713 PAD.n1942 0.000807692
R53490 PAD.n10374 PAD.n828 0.000807692
R53491 PAD.n11500 PAD.n10741 0.000807692
R53492 PAD.n7520 PAD.n7200 0.0008031
R53493 PAD.n9162 PAD.n9161 0.000798507
R53494 PAD.n1532 PAD.n1483 0.000793915
R53495 PAD.n6689 PAD.n5903 0.000789323
R53496 PAD.n8407 PAD.n4673 0.000789323
R53497 PAD.n8479 PAD.n8478 0.000789323
R53498 PAD.n8517 PAD.n2952 0.000789323
R53499 PAD PAD.n2946 0.00078473
R53500 PAD.n8479 PAD.n3633 0.000780138
R53501 PAD.n10719 PAD.n10716 0.000775545
R53502 PAD.n8420 PAD.n8419 0.000770953
R53503 PAD.n9163 PAD.n9162 0.000770953
R53504 PAD.n9175 PAD.n2139 0.000770953
R53505 PAD.n8185 PAD.n8184 0.000761768
R53506 PAD.n8195 PAD.n4840 0.000761768
R53507 PAD.n4843 PAD.n4842 0.000761768
R53508 PAD.n11522 PAD.n10741 0.000761768
R53509 PAD.n8205 PAD.n4673 0.000757176
R53510 PAD.n8420 PAD.n4331 0.000757176
R53511 PAD.n3342 PAD.n3296 0.000757176
R53512 PAD.n8492 PAD.n3339 0.000757176
R53513 PAD.n5974 PAD.n5903 0.000752583
R53514 PAD.n7206 PAD.n7200 0.000752583
R53515 PAD.n1533 PAD.n1532 0.000752583
R53516 PAD.n418 PAD.n373 0.000752583
R53517 PAD.n8502 PAD.n2997 0.000747991
R53518 PAD.n6711 PAD.n5552 0.000743398
R53519 PAD.n7792 PAD.n7791 0.000743398
R53520 PAD.n9455 PAD.n1988 0.000743398
R53521 PAD.n9713 PAD.n9712 0.000743398
R53522 PAD.n10374 PAD.n10373 0.000743398
R53523 PAD.n10389 PAD.n782 0.000743398
R53524 PAD.n8519 PAD.n8517 0.000738806
R53525 PAD.n6386 PAD.n6383 0.000734214
R53526 PAD.n7222 PAD.n7221 0.000734214
R53527 PAD.n9999 PAD.n1489 0.000734214
R53528 PAD.n10718 PAD.n10717 0.000734214
R53529 PAD.n7528 PAD.n7105 0.000729621
R53530 PAD.n2091 PAD.n2046 0.000729621
R53531 PAD.n8195 PAD.n8194 0.000725029
R53532 PAD.n9456 PAD.n9455 0.000725029
R53533 PAD.n11501 PAD.n11097 0.000725029
R53534 PAD.n7223 PAD.n7207 0.000720436
R53535 PAD.n8430 PAD.n4319 0.000715844
R53536 PAD.n8493 PAD.n3296 0.000706659
R53537 PAD.n8822 PAD.n2904 0.000706659
R53538 PAD.n8398 PAD.n8397 0.000697474
R53539 PAD.n8831 PAD.n2892 0.000697474
R53540 PAD.n9176 PAD.n2146 0.000692882
R53541 PAD.n9184 PAD.n2139 0.000692882
R53542 PAD.n8410 PAD.n8409 0.000688289
R53543 PAD.n8493 PAD.n8492 0.000688289
R53544 PAD.n9163 PAD.n2146 0.000688289
R53545 PAD.n9176 PAD.n9175 0.000688289
R53546 PAD.n8821 PAD.n8527 0.000683697
R53547 PAD.n8822 PAD.n8821 0.000679104
R53548 PAD.n2946 PAD.n2891 0.000679104
R53549 PAD.n1985 PAD.n1936 0.000679104
R53550 PAD.n11523 PAD.n10740 0.000679104
R53551 PAD.n4333 PAD.n4332 0.000674512
R53552 PAD.n10407 PAD.n435 0.000674512
R53553 PAD.n6396 PAD.n5904 0.00066992
R53554 PAD.n7521 PAD.n7158 0.00066992
R53555 PAD.n10008 PAD.n10007 0.00066992
R53556 PAD.n10702 PAD.n10701 0.00066992
R53557 PAD.n8194 PAD.n4843 0.000665327
R53558 PAD.n10362 PAD.n1130 0.000665327
R53559 PAD.n7802 PAD.n7801 0.000660735
R53560 PAD.n7060 PAD.n7059 0.000660735
R53561 PAD.n8183 PAD.n5183 0.000660735
R53562 PAD.n1131 PAD.n1118 0.000660735
R53563 PAD.n825 PAD.n776 0.000660735
R53564 PAD.n9151 PAD.n2487 0.000656142
R53565 PAD.n7783 PAD.n7782 0.00065155
R53566 PAD.n7820 PAD.n7819 0.00065155
R53567 PAD.n9742 PAD.n9741 0.00065155
R53568 PAD.n10728 PAD.n10727 0.00065155
R53569 PAD.n9445 PAD.n2089 0.000646958
R53570 PAD.n11507 PAD.n11098 0.000646958
R53571 PAD.n11302 PAD.n11096 0.000646958
R53572 PAD.n11509 PAD.n11099 0.000646958
R53573 PAD.n11510 PAD.n11100 0.000646958
R53574 PAD.n11513 PAD.n11105 0.000646958
R53575 PAD.n4842 PAD.n4841 0.000642365
R53576 PAD.n2089 PAD.n2037 0.000642365
R53577 PAD.n9732 PAD.n1594 0.00063318
R53578 PAD.n6699 PAD.n5894 0.000628588
R53579 PAD.n4321 PAD.n4028 0.000628588
R53580 PAD.n8410 PAD.n4331 0.000623995
R53581 PAD.n8419 PAD.n4333 0.000623995
R53582 PAD.n3339 PAD.n3287 0.000623995
R53583 PAD.n8519 PAD.n8518 0.000623995
R53584 PAD.n6689 PAD.n5904 0.000610218
R53585 PAD.n6683 PAD.n6678 0.000610218
R53586 PAD.n3687 PAD.n3641 0.000610218
R53587 PAD.n8468 PAD.n3684 0.000610218
R53588 PAD.n8408 PAD.n8407 0.000605626
R53589 PAD.n8478 PAD.n3342 0.000605626
R53590 PAD.n9185 PAD.n9184 0.000605626
R53591 PAD.n10007 PAD.n1483 0.000605626
R53592 PAD.n10017 PAD.n1140 0.000605626
R53593 PAD.n8832 PAD.n2891 0.000601033
R53594 PAD.n1988 PAD.n1942 0.000601033
R53595 PAD.n7521 PAD.n7520 0.000596441
R53596 PAD.n7207 PAD.n7206 0.000596441
R53597 PAD.n8175 PAD.n5190 0.000596441
R53598 PAD.n9722 PAD.n9721 0.000596441
R53599 PAD.n10397 PAD.n433 0.000596441
R53600 PAD.n10753 PAD.n21 0.000596441
R53601 PAD.n10754 PAD.n10753 0.000596441
R53602 PAD.n6683 PAD.n6682 0.000587256
R53603 PAD.n7216 PAD.n7215 0.000587256
R53604 PAD.n8469 PAD.n8468 0.000587256
R53605 PAD.n10017 PAD.n10016 0.000587256
R53606 PAD.n434 PAD.n425 0.000587256
R53607 PAD.n7791 PAD.n6713 0.000582664
R53608 PAD.n8186 PAD.n4840 0.000582664
R53609 PAD.n1132 PAD.n1131 0.000582664
R53610 PAD.n6700 PAD.n6699 0.000578071
R53611 PAD.n7783 PAD.n7061 0.000578071
R53612 PAD.n10362 PAD.n10361 0.000578071
R53613 PAD.n10398 PAD.n10397 0.000578071
R53614 PAD.n10728 PAD.n32 0.000578071
R53615 PAD.n367 PAD.n20 0.000578071
R53616 PAD.n2894 PAD.n2879 0.000573479
R53617 PAD.n9143 PAD.n2494 0.000573479
R53618 PAD.n7829 PAD.n7828 0.000568886
R53619 PAD.n1593 PAD.n1586 0.000568886
R53620 PAD.n11534 PAD.n20 0.000568886
R53621 PAD.n8163 PAD.n5190 0.000564294
R53622 PAD.n10389 PAD.n10388 0.000564294
R53623 PAD.n8398 PAD.n4682 0.000559702
R53624 PAD.n9152 PAD.n2494 0.000559702
R53625 PAD.n9160 PAD.n2487 0.000559702
R53626 PAD.n9446 PAD.n2046 0.000559702
R53627 PAD.n9142 PAD.n9141 0.000550517
R53628 PAD.n9722 PAD.n1592 0.000550517
R53629 PAD.n7802 PAD.n5551 0.000545924
R53630 PAD.n8445 PAD.n8444 0.000545924
R53631 PAD.n8503 PAD.n8502 0.000541332
R53632 PAD.n3289 PAD.n2952 0.000541332
R53633 PAD.n9128 PAD.n2879 0.000541332
R53634 PAD.n9140 PAD.n2834 0.000541332
R53635 PAD.n10702 PAD.n419 0.000541332
R53636 PAD.n10716 PAD.n373 0.000541332
R53637 PAD.n6373 PAD.n5963 0.000536739
R53638 PAD.n5982 PAD.n5964 0.000536739
R53639 PAD.n5981 PAD.n5962 0.000536739
R53640 PAD.n5980 PAD.n5965 0.000536739
R53641 PAD.n5979 PAD.n5966 0.000536739
R53642 PAD.n8454 PAD.n3977 0.000532147
R53643 PAD.n9129 PAD.n2834 0.000532147
R53644 PAD.n7820 PAD.n5204 0.000522962
R53645 PAD.n7828 PAD.n5197 0.000522962
R53646 PAD.n8205 PAD.n4724 0.000522962
R53647 PAD.n9187 PAD.n9186 0.000522962
R53648 PAD.n8174 PAD.n5183 0.00051837
R53649 PAD.n9712 PAD.n1986 0.00051837
R53650 PAD.n1120 PAD.n828 0.00051837
R53651 PAD.n8165 PAD.n8164 0.000513777
R53652 PAD.n9733 PAD.n9732 0.000513777
R53653 PAD.n9741 PAD.n1536 0.000513777
R53654 PAD.n9999 PAD.n9998 0.000513777
R53655 PAD.n11533 PAD.n11532 0.000513777
R53656 PAD.n10755 PAD.n10740 0.000513777
R53657 PAD.n6680 PAD.n6679 0.000504592
R53658 PAD.n7528 PAD.n7103 0.000504592
R53659 PAD.n8431 PAD.n4028 0.000504592
R53660 PAD.n8444 PAD.n3983 0.000504592
R53661 PAD.n8453 PAD.n3687 0.000504592
R53662 PAD.n8527 PAD 0.000504592
R53663 PAD.n1142 PAD.n1141 0.000504592
R53664 PAD.n10408 PAD.n10407 0.000504592
R53665 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_1.nmos_6p0_CDNS_4066195314530_0.D.n0 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_1.nmos_6p0_CDNS_4066195314530_0.D.t4 37.5434
R53666 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_1.nmos_6p0_CDNS_4066195314530_0.D.n1 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_1.nmos_6p0_CDNS_4066195314530_0.D.t5 37.5434
R53667 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_1.nmos_6p0_CDNS_4066195314530_0.D.n0 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_1.nmos_6p0_CDNS_4066195314530_0.D.t2 25.3941
R53668 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_1.nmos_6p0_CDNS_4066195314530_0.D.n1 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_1.nmos_6p0_CDNS_4066195314530_0.D.t3 25.3941
R53669 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_1.nmos_6p0_CDNS_4066195314530_0.D.n1 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_1.nmos_6p0_CDNS_4066195314530_0.D.n0 8.44221
R53670 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_1.nmos_6p0_CDNS_4066195314530_0.D.t1 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_1.nmos_6p0_CDNS_4066195314530_0.D.n1 4.90922
R53671 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_1.nmos_6p0_CDNS_4066195314530_0.D.t1 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_1.nmos_6p0_CDNS_4066195314530_0.D.t0 2.6373
R53672 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_1.Z.n2 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_1.Z.t4 37.5434
R53673 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_1.Z.n3 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_1.Z.t5 37.5434
R53674 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_1.Z.n0 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_1.Z.t7 29.034
R53675 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_1.Z.n0 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_1.Z.t12 28.9248
R53676 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_1.Z.n0 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_1.Z.t11 28.9248
R53677 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_1.Z.n0 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_1.Z.t3 28.9248
R53678 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_1.Z.n0 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_1.Z.t2 28.9248
R53679 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_1.Z.n2 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_1.Z.t9 25.3941
R53680 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_1.Z.n3 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_1.Z.t10 25.3941
R53681 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_1.Z.n1 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_1.Z.t13 24.9104
R53682 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_1.Z.n1 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_1.Z.t6 24.8782
R53683 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_1.Z.n1 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_1.Z.t8 24.5969
R53684 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_1.Z GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_1.Z.n0 10.2118
R53685 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_1.Z.n3 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_1.Z.n2 8.44221
R53686 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_1.Z GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_1.Z.n3 4.40816
R53687 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_1.Z.n0 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_1.Z 3.54046
R53688 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_1.Z GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_1.Z.n1 2.40605
R53689 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_1.Z GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_1.Z.t1 2.2999
R53690 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_1.Z GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_1.Z.t0 2.0632
R53691 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_drv_0.Z.n2 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_drv_0.Z.t5 40.4112
R53692 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_drv_0.Z.n3 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_drv_0.Z.t4 40.4112
R53693 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_drv_0.Z.n4 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_drv_0.Z.t11 40.4112
R53694 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_drv_0.Z.n5 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_drv_0.Z.t7 40.4112
R53695 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_drv_0.Z.n1 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_drv_0.Z.t1 40.4112
R53696 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_drv_0.Z.n0 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_drv_0.Z.t9 40.4112
R53697 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_drv_0.Z.n2 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_drv_0.Z.t3 35.3012
R53698 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_drv_0.Z.n3 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_drv_0.Z.t2 35.3012
R53699 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_drv_0.Z.n4 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_drv_0.Z.t10 35.3012
R53700 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_drv_0.Z.n5 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_drv_0.Z.t6 35.3012
R53701 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_drv_0.Z.n1 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_drv_0.Z.t12 35.3012
R53702 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_drv_0.Z.n0 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_drv_0.Z.t8 35.3012
R53703 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_drv_0.Z.t0 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_drv_0.nmos_6p0_CDNS_4066195314550_0.D 6.07134
R53704 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_drv_0.nmos_6p0_CDNS_4066195314550_0.D GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_drv_0.Z.n0 4.13606
R53705 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_drv_0.nmos_6p0_CDNS_4066195314550_0.D GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_drv_0.Z.n1 4.0005
R53706 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_drv_0.nmos_6p0_CDNS_4066195314550_0.D GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_drv_0.Z.n5 4.0005
R53707 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_drv_0.nmos_6p0_CDNS_4066195314550_0.D GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_drv_0.Z.n4 4.0005
R53708 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_drv_0.nmos_6p0_CDNS_4066195314550_0.D GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_drv_0.Z.n3 4.0005
R53709 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_drv_0.nmos_6p0_CDNS_4066195314550_0.D GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_drv_0.Z.n2 4.0005
R53710 Y Y.n13 9.7577
R53711 Y.n5 Y.n4 6.3005
R53712 Y.n4 Y 3.18489
R53713 Y.n1 Y.n0 2.08611
R53714 Y.n3 Y.n2 2.08611
R53715 Y.n11 Y.n10 1.67295
R53716 Y.n11 Y.n9 1.09506
R53717 Y.n12 Y.n8 1.09506
R53718 Y.n0 Y.t1 1.0925
R53719 Y.n0 Y.t5 1.0925
R53720 Y.n2 Y.t2 1.0925
R53721 Y.n2 Y.t0 1.0925
R53722 Y.n4 Y.t4 1.0925
R53723 Y.n4 Y.t3 1.0925
R53724 Y.n6 Y.n5 0.825895
R53725 Y.n13 Y.n7 0.770237
R53726 Y.n12 Y.n11 0.578395
R53727 Y.n7 Y.n6 0.578395
R53728 Y.n10 Y.t11 0.5205
R53729 Y.n10 Y.t10 0.5205
R53730 Y.n9 Y.t9 0.5205
R53731 Y.n9 Y.t7 0.5205
R53732 Y.n8 Y.t8 0.5205
R53733 Y.n8 Y.t6 0.5205
R53734 Y.n13 Y.n12 0.457605
R53735 Y.n7 Y.n1 0.336924
R53736 Y.n6 Y.n3 0.336924
R53737 Y.n5 Y 0.1355
R53738 Y.n1 Y 0.0456808
R53739 Y.n3 Y 0.0456808
R53740 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.nmos_6p0_CDNS_4066195314511_1.S.n0 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.nmos_6p0_CDNS_4066195314511_1.S.t3 38.8469
R53741 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.nmos_6p0_CDNS_4066195314511_1.S.n0 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.nmos_6p0_CDNS_4066195314511_1.S.t2 22.5262
R53742 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.nmos_6p0_CDNS_4066195314511_1.S GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.nmos_6p0_CDNS_4066195314511_1.S.n0 12.9666
R53743 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.nmos_6p0_CDNS_4066195314511_1.S GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.nmos_6p0_CDNS_4066195314511_1.S.t0 2.19095
R53744 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.nmos_6p0_CDNS_4066195314511_1.S GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.nmos_6p0_CDNS_4066195314511_1.S.t1 1.9977
R53745 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_1.nmos_6p0_CDNS_4066195314511_1.S.n0 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_1.nmos_6p0_CDNS_4066195314511_1.S.t3 38.8469
R53746 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_1.nmos_6p0_CDNS_4066195314511_1.S.n0 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_1.nmos_6p0_CDNS_4066195314511_1.S.t2 22.5262
R53747 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_1.nmos_6p0_CDNS_4066195314511_1.S GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_1.nmos_6p0_CDNS_4066195314511_1.S.n0 12.9666
R53748 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_1.nmos_6p0_CDNS_4066195314511_1.S GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_1.nmos_6p0_CDNS_4066195314511_1.S.t1 2.19095
R53749 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_1.nmos_6p0_CDNS_4066195314511_1.S GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_1.nmos_6p0_CDNS_4066195314511_1.S.t0 1.9977
R53750 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_a_0.nmos_6p0_CDNS_4066195314511_2.D GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_a_0.nmos_6p0_CDNS_4066195314511_1.S.n0 1.15854
R53751 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_a_0.nmos_6p0_CDNS_4066195314511_1.S.n0 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_a_0.nmos_6p0_CDNS_4066195314511_1.S.t1 0.5465
R53752 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_a_0.nmos_6p0_CDNS_4066195314511_1.S.n0 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_a_0.nmos_6p0_CDNS_4066195314511_1.S.t0 0.5465
R53753 GF_NI_IN_C_BASE_0.comp018green_out_predrv_3.nmos_6p0_CDNS_4066195314519_2.S.n1 GF_NI_IN_C_BASE_0.comp018green_out_predrv_3.nmos_6p0_CDNS_4066195314519_2.S.t2 79.0838
R53754 GF_NI_IN_C_BASE_0.comp018green_out_predrv_3.nmos_6p0_CDNS_4066195314519_2.S.n1 GF_NI_IN_C_BASE_0.comp018green_out_predrv_3.nmos_6p0_CDNS_4066195314519_2.S.t5 78.041
R53755 GF_NI_IN_C_BASE_0.comp018green_out_predrv_3.nmos_6p0_CDNS_4066195314519_2.S.n5 GF_NI_IN_C_BASE_0.comp018green_out_predrv_3.nmos_6p0_CDNS_4066195314519_2.S.t4 34.4148
R53756 GF_NI_IN_C_BASE_0.comp018green_out_predrv_3.nmos_6p0_CDNS_4066195314519_2.S.n2 GF_NI_IN_C_BASE_0.comp018green_out_predrv_3.nmos_6p0_CDNS_4066195314519_2.S.t3 34.4148
R53757 GF_NI_IN_C_BASE_0.comp018green_out_predrv_3.nmos_6p0_CDNS_4066195314519_2.S.n3 GF_NI_IN_C_BASE_0.comp018green_out_predrv_3.nmos_6p0_CDNS_4066195314519_2.S.t6 34.4148
R53758 GF_NI_IN_C_BASE_0.comp018green_out_predrv_3.nmos_6p0_CDNS_4066195314519_2.S.n4 GF_NI_IN_C_BASE_0.comp018green_out_predrv_3.nmos_6p0_CDNS_4066195314519_2.S.t7 34.4148
R53759 GF_NI_IN_C_BASE_0.comp018green_out_predrv_3.nmos_6p0_CDNS_4066195314519_2.S.n3 GF_NI_IN_C_BASE_0.comp018green_out_predrv_3.nmos_6p0_CDNS_4066195314519_2.S.n2 10.9956
R53760 GF_NI_IN_C_BASE_0.comp018green_out_predrv_3.nmos_6p0_CDNS_4066195314519_2.S.n4 GF_NI_IN_C_BASE_0.comp018green_out_predrv_3.nmos_6p0_CDNS_4066195314519_2.S.n3 10.9956
R53761 GF_NI_IN_C_BASE_0.comp018green_out_predrv_3.nmos_6p0_CDNS_4066195314519_2.S.n5 GF_NI_IN_C_BASE_0.comp018green_out_predrv_3.nmos_6p0_CDNS_4066195314519_2.S.n4 10.9956
R53762 GF_NI_IN_C_BASE_0.comp018green_out_predrv_3.nmos_6p0_CDNS_4066195314519_2.S.n6 GF_NI_IN_C_BASE_0.comp018green_out_predrv_3.nmos_6p0_CDNS_4066195314519_2.S.n5 9.95826
R53763 GF_NI_IN_C_BASE_0.comp018green_out_predrv_3.nmos_6p0_CDNS_4066195314519_2.S.n2 GF_NI_IN_C_BASE_0.comp018green_out_predrv_3.nmos_6p0_CDNS_4066195314519_2.S.n1 8.49628
R53764 GF_NI_IN_C_BASE_0.comp018green_out_predrv_3.nmos_6p0_CDNS_4066195314519_2.S.n0 GF_NI_IN_C_BASE_0.comp018green_out_predrv_3.nmos_6p0_CDNS_4066195314519_2.S.t1 2.12938
R53765 GF_NI_IN_C_BASE_0.comp018green_out_predrv_3.nmos_6p0_CDNS_4066195314519_2.S.n0 GF_NI_IN_C_BASE_0.comp018green_out_predrv_3.nmos_6p0_CDNS_4066195314519_2.S.t0 1.97771
R53766 GF_NI_IN_C_BASE_0.comp018green_out_predrv_3.nmos_6p0_CDNS_4066195314519_2.S.n6 GF_NI_IN_C_BASE_0.comp018green_out_predrv_3.nmos_6p0_CDNS_4066195314519_2.S.n0 1.32326
R53767 GF_NI_IN_C_BASE_0.comp018green_out_predrv_3.nmos_6p0_CDNS_4066195314519_2.S GF_NI_IN_C_BASE_0.comp018green_out_predrv_3.nmos_6p0_CDNS_4066195314519_2.S.n6 1.25751
R53768 GF_NI_IN_C_BASE_0.ndrive_Y_<1> GF_NI_IN_C_BASE_0.ndrive_Y_<1>.t5 90.7338
R53769 GF_NI_IN_C_BASE_0.ndrive_Y_<1>.n0 GF_NI_IN_C_BASE_0.ndrive_Y_<1>.t1 5.90425
R53770 GF_NI_IN_C_BASE_0.ndrive_Y_<1>.n2 GF_NI_IN_C_BASE_0.ndrive_Y_<1>.t4 2.41832
R53771 GF_NI_IN_C_BASE_0.ndrive_Y_<1>.n1 GF_NI_IN_C_BASE_0.ndrive_Y_<1>.t2 1.84043
R53772 GF_NI_IN_C_BASE_0.ndrive_Y_<1>.n0 GF_NI_IN_C_BASE_0.ndrive_Y_<1> 1.5749
R53773 GF_NI_IN_C_BASE_0.ndrive_Y_<1>.n3 GF_NI_IN_C_BASE_0.ndrive_Y_<1>.n2 1.48076
R53774 GF_NI_IN_C_BASE_0.ndrive_Y_<1>.n1 GF_NI_IN_C_BASE_0.ndrive_Y_<1>.n0 1.09118
R53775 GF_NI_IN_C_BASE_0.ndrive_Y_<1> GF_NI_IN_C_BASE_0.ndrive_Y_<1>.n3 0.9455
R53776 GF_NI_IN_C_BASE_0.ndrive_Y_<1>.n2 GF_NI_IN_C_BASE_0.ndrive_Y_<1>.n1 0.578395
R53777 GF_NI_IN_C_BASE_0.ndrive_Y_<1> GF_NI_IN_C_BASE_0.ndrive_Y_<1>.t3 0.500893
R53778 GF_NI_IN_C_BASE_0.ndrive_Y_<1>.n3 GF_NI_IN_C_BASE_0.ndrive_Y_<1>.t0 0.360167
R53779 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_drv_0.nmos_6p0_CDNS_4066195314547_0.S.n3 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_drv_0.nmos_6p0_CDNS_4066195314547_0.S.t8 41.7148
R53780 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_drv_0.nmos_6p0_CDNS_4066195314547_0.S.n2 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_drv_0.nmos_6p0_CDNS_4066195314547_0.S.t7 41.7148
R53781 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_drv_0.nmos_6p0_CDNS_4066195314547_0.S.n1 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_drv_0.nmos_6p0_CDNS_4066195314547_0.S.t4 34.2225
R53782 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_drv_0.nmos_6p0_CDNS_4066195314547_0.S.n1 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_drv_0.nmos_6p0_CDNS_4066195314547_0.S.t3 34.0869
R53783 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_drv_0.nmos_6p0_CDNS_4066195314547_0.S.n3 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_drv_0.nmos_6p0_CDNS_4066195314547_0.S.t6 30.0869
R53784 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_drv_0.nmos_6p0_CDNS_4066195314547_0.S.n2 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_drv_0.nmos_6p0_CDNS_4066195314547_0.S.t5 30.0869
R53785 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_drv_0.nmos_6p0_CDNS_4066195314547_0.S.n0 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_drv_0.nmos_6p0_CDNS_4066195314547_0.S.t2 4.67357
R53786 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_drv_0.nmos_6p0_CDNS_4066195314547_0.S.n1 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_drv_0.nmos_6p0_CDNS_4066195314547_0.S.n2 4.0005
R53787 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_drv_0.nmos_6p0_CDNS_4066195314547_0.S.n1 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_drv_0.nmos_6p0_CDNS_4066195314547_0.S.n3 4.0005
R53788 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_drv_0.nmos_6p0_CDNS_4066195314547_0.S.n0 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_drv_0.nmos_6p0_CDNS_4066195314547_0.S 2.87207
R53789 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_drv_0.nmos_6p0_CDNS_4066195314547_0.S.n0 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_drv_0.nmos_6p0_CDNS_4066195314547_0.S.t1 1.81789
R53790 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_drv_0.nmos_6p0_CDNS_4066195314547_0.S GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_drv_0.nmos_6p0_CDNS_4066195314547_0.S.t0 1.22475
R53791 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_drv_0.nmos_6p0_CDNS_4066195314547_0.S.n1 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_drv_0.nmos_6p0_CDNS_4066195314547_0.S.n0 1.14881
R53792 GF_NI_IN_C_BASE_0.comp018green_out_predrv_2.nmos_6p0_CDNS_4066195314519_2.S.n1 GF_NI_IN_C_BASE_0.comp018green_out_predrv_2.nmos_6p0_CDNS_4066195314519_2.S.t6 79.0838
R53793 GF_NI_IN_C_BASE_0.comp018green_out_predrv_2.nmos_6p0_CDNS_4066195314519_2.S.n1 GF_NI_IN_C_BASE_0.comp018green_out_predrv_2.nmos_6p0_CDNS_4066195314519_2.S.t5 78.041
R53794 GF_NI_IN_C_BASE_0.comp018green_out_predrv_2.nmos_6p0_CDNS_4066195314519_2.S.n5 GF_NI_IN_C_BASE_0.comp018green_out_predrv_2.nmos_6p0_CDNS_4066195314519_2.S.t3 34.4148
R53795 GF_NI_IN_C_BASE_0.comp018green_out_predrv_2.nmos_6p0_CDNS_4066195314519_2.S.n2 GF_NI_IN_C_BASE_0.comp018green_out_predrv_2.nmos_6p0_CDNS_4066195314519_2.S.t2 34.4148
R53796 GF_NI_IN_C_BASE_0.comp018green_out_predrv_2.nmos_6p0_CDNS_4066195314519_2.S.n4 GF_NI_IN_C_BASE_0.comp018green_out_predrv_2.nmos_6p0_CDNS_4066195314519_2.S.t4 34.4148
R53797 GF_NI_IN_C_BASE_0.comp018green_out_predrv_2.nmos_6p0_CDNS_4066195314519_2.S.n3 GF_NI_IN_C_BASE_0.comp018green_out_predrv_2.nmos_6p0_CDNS_4066195314519_2.S.t7 34.4148
R53798 GF_NI_IN_C_BASE_0.comp018green_out_predrv_2.nmos_6p0_CDNS_4066195314519_2.S.n5 GF_NI_IN_C_BASE_0.comp018green_out_predrv_2.nmos_6p0_CDNS_4066195314519_2.S.n4 10.9956
R53799 GF_NI_IN_C_BASE_0.comp018green_out_predrv_2.nmos_6p0_CDNS_4066195314519_2.S.n4 GF_NI_IN_C_BASE_0.comp018green_out_predrv_2.nmos_6p0_CDNS_4066195314519_2.S.n3 10.9956
R53800 GF_NI_IN_C_BASE_0.comp018green_out_predrv_2.nmos_6p0_CDNS_4066195314519_2.S.n3 GF_NI_IN_C_BASE_0.comp018green_out_predrv_2.nmos_6p0_CDNS_4066195314519_2.S.n2 10.9956
R53801 GF_NI_IN_C_BASE_0.comp018green_out_predrv_2.nmos_6p0_CDNS_4066195314519_2.S.n6 GF_NI_IN_C_BASE_0.comp018green_out_predrv_2.nmos_6p0_CDNS_4066195314519_2.S.n5 9.95826
R53802 GF_NI_IN_C_BASE_0.comp018green_out_predrv_2.nmos_6p0_CDNS_4066195314519_2.S.n2 GF_NI_IN_C_BASE_0.comp018green_out_predrv_2.nmos_6p0_CDNS_4066195314519_2.S.n1 8.49628
R53803 GF_NI_IN_C_BASE_0.comp018green_out_predrv_2.nmos_6p0_CDNS_4066195314519_2.S.n0 GF_NI_IN_C_BASE_0.comp018green_out_predrv_2.nmos_6p0_CDNS_4066195314519_2.S.t1 2.12938
R53804 GF_NI_IN_C_BASE_0.comp018green_out_predrv_2.nmos_6p0_CDNS_4066195314519_2.S.n0 GF_NI_IN_C_BASE_0.comp018green_out_predrv_2.nmos_6p0_CDNS_4066195314519_2.S.t0 1.97771
R53805 GF_NI_IN_C_BASE_0.comp018green_out_predrv_2.nmos_6p0_CDNS_4066195314519_2.S.n6 GF_NI_IN_C_BASE_0.comp018green_out_predrv_2.nmos_6p0_CDNS_4066195314519_2.S.n0 1.32326
R53806 GF_NI_IN_C_BASE_0.comp018green_out_predrv_2.nmos_6p0_CDNS_4066195314519_2.S GF_NI_IN_C_BASE_0.comp018green_out_predrv_2.nmos_6p0_CDNS_4066195314519_2.S.n6 1.25751
R53807 GF_NI_IN_C_BASE_0.ndrive_x_<2> GF_NI_IN_C_BASE_0.ndrive_x_<2>.t3 90.7537
R53808 GF_NI_IN_C_BASE_0.ndrive_x_<2>.t0 GF_NI_IN_C_BASE_0.ndrive_x_<2>.n0 7.28458
R53809 GF_NI_IN_C_BASE_0.ndrive_x_<2>.n0 GF_NI_IN_C_BASE_0.ndrive_x_<2>.t1 6.03391
R53810 GF_NI_IN_C_BASE_0.ndrive_x_<2>.n0 GF_NI_IN_C_BASE_0.ndrive_x_<2> 1.45646
R53811 GF_NI_IN_C_BASE_0.ndrive_x_<2> GF_NI_IN_C_BASE_0.ndrive_x_<2>.t0 0.951421
R53812 GF_NI_IN_C_BASE_0.ndrive_x_<2>.t2 GF_NI_IN_C_BASE_0.ndrive_x_<2> 0.773893
R53813 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_a_0.nmos_6p0_CDNS_4066195314511_1.D.n0 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_a_0.nmos_6p0_CDNS_4066195314511_1.D.t3 38.8469
R53814 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_a_0.nmos_6p0_CDNS_4066195314511_1.D.n0 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_a_0.nmos_6p0_CDNS_4066195314511_1.D.t2 22.5262
R53815 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_a_0.nmos_6p0_CDNS_4066195314511_1.D GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_a_0.nmos_6p0_CDNS_4066195314511_1.D.n0 12.9564
R53816 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_a_0.nmos_6p0_CDNS_4066195314511_1.D GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_a_0.nmos_6p0_CDNS_4066195314511_1.D.t1 2.19095
R53817 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_a_0.nmos_6p0_CDNS_4066195314511_1.D GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_a_0.nmos_6p0_CDNS_4066195314511_1.D.t0 1.9977
R53818 GF_NI_IN_C_BASE_0.ndrive_x_<0> GF_NI_IN_C_BASE_0.ndrive_x_<0>.t3 89.2634
R53819 GF_NI_IN_C_BASE_0.ndrive_x_<0>.t0 GF_NI_IN_C_BASE_0.ndrive_x_<0>.n0 7.28458
R53820 GF_NI_IN_C_BASE_0.ndrive_x_<0>.n0 GF_NI_IN_C_BASE_0.ndrive_x_<0>.t1 6.03391
R53821 GF_NI_IN_C_BASE_0.ndrive_x_<0>.n0 GF_NI_IN_C_BASE_0.ndrive_x_<0> 1.45646
R53822 GF_NI_IN_C_BASE_0.ndrive_x_<0> GF_NI_IN_C_BASE_0.ndrive_x_<0>.t0 0.951421
R53823 GF_NI_IN_C_BASE_0.ndrive_x_<0>.t2 GF_NI_IN_C_BASE_0.ndrive_x_<0> 0.773893
R53824 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_1.EN GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_1.EN.t2 82.1164
R53825 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_1.EN GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_1.EN.t3 82.1164
R53826 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_1.EN.n1 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_1.EN.t5 44.3219
R53827 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_1.EN GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_1.EN.t6 42.2319
R53828 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_1.EN GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_1.EN.t7 42.2319
R53829 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_1.EN.n1 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_1.EN.t4 28.0534
R53830 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_1.EN.n0 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_1.EN 11.0504
R53831 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_1.EN GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_1.EN.n0 7.90454
R53832 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_1.EN.n0 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_1.EN 7.30826
R53833 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_1.EN GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_1.EN.n1 4.09808
R53834 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_1.EN GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_1.EN.t0 1.53534
R53835 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_1.EN GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_1.EN.t1 1.33388
R53836 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_logic_pupd_0.PDB_OUT.n0 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_logic_pupd_0.PDB_OUT.t1 35.9269
R53837 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_logic_pupd_0.PDB_OUT.n0 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_logic_pupd_0.PDB_OUT.t2 30.9212
R53838 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_logic_pupd_0.PDB_OUT.t0 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_0.A 25.1335
R53839 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_0.A GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_logic_pupd_0.PDB_OUT.n0 4.0005
R53840 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_0.nmos_6p0_CDNS_4066195314530_0.D.n0 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_0.nmos_6p0_CDNS_4066195314530_0.D.t3 37.5434
R53841 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_0.nmos_6p0_CDNS_4066195314530_0.D.n1 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_0.nmos_6p0_CDNS_4066195314530_0.D.t4 37.5434
R53842 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_0.nmos_6p0_CDNS_4066195314530_0.D.n0 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_0.nmos_6p0_CDNS_4066195314530_0.D.t5 25.3941
R53843 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_0.nmos_6p0_CDNS_4066195314530_0.D.n1 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_0.nmos_6p0_CDNS_4066195314530_0.D.t2 25.3941
R53844 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_0.nmos_6p0_CDNS_4066195314530_0.D.n1 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_0.nmos_6p0_CDNS_4066195314530_0.D.n0 8.44221
R53845 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_0.nmos_6p0_CDNS_4066195314530_0.D.t1 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_0.nmos_6p0_CDNS_4066195314530_0.D.n1 4.90922
R53846 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_0.nmos_6p0_CDNS_4066195314530_0.D.t1 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_0.nmos_6p0_CDNS_4066195314530_0.D.t0 2.6373
R53847 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_pupd_0.ppolyf_u_CDNS_4066195314533_0.PLUS.t0 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_pupd_0.ppolyf_u_CDNS_4066195314533_0.PLUS 11.0117
R53848 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_pupd_0.ppolyf_u_CDNS_4066195314533_0.PLUS GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_pupd_0.ppolyf_u_CDNS_4066195314533_0.PLUS.t1 11.0117
R53849 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_pupd_0.ppolyf_u_CDNS_4066195314533_0.MINUS.t0 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_pupd_0.ppolyf_u_CDNS_4066195314533_0.MINUS.t1 22.3936
R53850 GF_NI_IN_C_BASE_0.comp018green_out_predrv_0.SL.n6 GF_NI_IN_C_BASE_0.comp018green_out_predrv_0.SL.t7 79.2576
R53851 GF_NI_IN_C_BASE_0.comp018green_out_predrv_0.SL.n5 GF_NI_IN_C_BASE_0.comp018green_out_predrv_0.SL.t11 79.2576
R53852 GF_NI_IN_C_BASE_0.comp018green_out_predrv_0.SL.n4 GF_NI_IN_C_BASE_0.comp018green_out_predrv_0.SL.t13 79.2576
R53853 GF_NI_IN_C_BASE_0.comp018green_out_predrv_0.SL.n3 GF_NI_IN_C_BASE_0.comp018green_out_predrv_0.SL.t3 79.2576
R53854 GF_NI_IN_C_BASE_0.comp018green_out_predrv_0.SL.n6 GF_NI_IN_C_BASE_0.comp018green_out_predrv_0.SL.t4 77.8672
R53855 GF_NI_IN_C_BASE_0.comp018green_out_predrv_0.SL.n5 GF_NI_IN_C_BASE_0.comp018green_out_predrv_0.SL.t5 77.8672
R53856 GF_NI_IN_C_BASE_0.comp018green_out_predrv_0.SL.n4 GF_NI_IN_C_BASE_0.comp018green_out_predrv_0.SL.t12 77.8672
R53857 GF_NI_IN_C_BASE_0.comp018green_out_predrv_0.SL.n3 GF_NI_IN_C_BASE_0.comp018green_out_predrv_0.SL.t10 77.8672
R53858 GF_NI_IN_C_BASE_0.comp018green_out_predrv_0.SL.n1 GF_NI_IN_C_BASE_0.comp018green_out_predrv_0.SL.t8 37.5434
R53859 GF_NI_IN_C_BASE_0.comp018green_out_predrv_0.SL.n2 GF_NI_IN_C_BASE_0.comp018green_out_predrv_0.SL.t2 37.5434
R53860 GF_NI_IN_C_BASE_0.comp018green_out_predrv_0.SL.n1 GF_NI_IN_C_BASE_0.comp018green_out_predrv_0.SL.t6 25.3941
R53861 GF_NI_IN_C_BASE_0.comp018green_out_predrv_0.SL.n2 GF_NI_IN_C_BASE_0.comp018green_out_predrv_0.SL.t9 25.3941
R53862 GF_NI_IN_C_BASE_0.comp018green_out_predrv_0.SL.n0 GF_NI_IN_C_BASE_0.comp018green_out_predrv_0.SL 12.2973
R53863 GF_NI_IN_C_BASE_0.comp018green_out_predrv_0.SL.n7 GF_NI_IN_C_BASE_0.comp018green_out_predrv_0.SL.n0 8.47471
R53864 GF_NI_IN_C_BASE_0.comp018green_out_predrv_0.SL.n2 GF_NI_IN_C_BASE_0.comp018green_out_predrv_0.SL.n1 8.44221
R53865 GF_NI_IN_C_BASE_0.comp018green_out_predrv_0.SL.n0 GF_NI_IN_C_BASE_0.comp018green_out_predrv_0.SL 8.14787
R53866 GF_NI_IN_C_BASE_0.comp018green_out_predrv_0.SL.n0 GF_NI_IN_C_BASE_0.comp018green_out_predrv_0.SL 6.07313
R53867 GF_NI_IN_C_BASE_0.comp018green_out_predrv_0.SL GF_NI_IN_C_BASE_0.comp018green_out_predrv_0.SL.n7 5.15345
R53868 GF_NI_IN_C_BASE_0.comp018green_out_predrv_0.SL GF_NI_IN_C_BASE_0.comp018green_out_predrv_0.SL.n3 5.13701
R53869 GF_NI_IN_C_BASE_0.comp018green_out_predrv_0.SL GF_NI_IN_C_BASE_0.comp018green_out_predrv_0.SL.n4 5.13701
R53870 GF_NI_IN_C_BASE_0.comp018green_out_predrv_0.SL GF_NI_IN_C_BASE_0.comp018green_out_predrv_0.SL.n5 5.13701
R53871 GF_NI_IN_C_BASE_0.comp018green_out_predrv_0.SL GF_NI_IN_C_BASE_0.comp018green_out_predrv_0.SL.n6 5.13701
R53872 GF_NI_IN_C_BASE_0.comp018green_out_predrv_0.SL GF_NI_IN_C_BASE_0.comp018green_out_predrv_0.SL.n2 4.34849
R53873 GF_NI_IN_C_BASE_0.comp018green_out_predrv_0.SL.n7 GF_NI_IN_C_BASE_0.comp018green_out_predrv_0.SL 3.78055
R53874 GF_NI_IN_C_BASE_0.comp018green_out_predrv_0.SL.t0 GF_NI_IN_C_BASE_0.comp018green_out_predrv_0.SL 3.17854
R53875 GF_NI_IN_C_BASE_0.comp018green_out_predrv_0.SL GF_NI_IN_C_BASE_0.comp018green_out_predrv_0.SL.t1 2.94253
R53876 GF_NI_IN_C_BASE_0.pdrive_x_<2>.n2 GF_NI_IN_C_BASE_0.pdrive_x_<2>.t5 113.415
R53877 GF_NI_IN_C_BASE_0.pdrive_x_<2>.n2 GF_NI_IN_C_BASE_0.pdrive_x_<2>.t4 112.603
R53878 GF_NI_IN_C_BASE_0.pdrive_x_<2>.t2 GF_NI_IN_C_BASE_0.pdrive_x_<2>.n1 6.12025
R53879 GF_NI_IN_C_BASE_0.pdrive_x_<2> GF_NI_IN_C_BASE_0.pdrive_x_<2>.n2 2.40448
R53880 GF_NI_IN_C_BASE_0.pdrive_x_<2>.t3 GF_NI_IN_C_BASE_0.pdrive_x_<2>.n1 2.26404
R53881 GF_NI_IN_C_BASE_0.pdrive_x_<2> GF_NI_IN_C_BASE_0.pdrive_x_<2>.n0 1.4357
R53882 GF_NI_IN_C_BASE_0.pdrive_x_<2>.n1 GF_NI_IN_C_BASE_0.pdrive_x_<2>.n0 1.03582
R53883 GF_NI_IN_C_BASE_0.pdrive_x_<2> GF_NI_IN_C_BASE_0.pdrive_x_<2>.t0 0.779294
R53884 GF_NI_IN_C_BASE_0.pdrive_x_<2> GF_NI_IN_C_BASE_0.pdrive_x_<2>.t3 0.7439
R53885 GF_NI_IN_C_BASE_0.pdrive_x_<2>.n0 GF_NI_IN_C_BASE_0.pdrive_x_<2>.t1 0.66992
R53886 GF_NI_IN_C_BASE_0.ppolyf_u_CDNS_4066195314551_0.MINUS.t0 GF_NI_IN_C_BASE_0.ppolyf_u_CDNS_4066195314551_0.MINUS.t1 60.8949
R53887 GF_NI_IN_C_BASE_0.comp018green_out_predrv_0.nmos_6p0_CDNS_4066195314519_2.S.n1 GF_NI_IN_C_BASE_0.comp018green_out_predrv_0.nmos_6p0_CDNS_4066195314519_2.S.t6 79.0838
R53888 GF_NI_IN_C_BASE_0.comp018green_out_predrv_0.nmos_6p0_CDNS_4066195314519_2.S.n1 GF_NI_IN_C_BASE_0.comp018green_out_predrv_0.nmos_6p0_CDNS_4066195314519_2.S.t4 78.041
R53889 GF_NI_IN_C_BASE_0.comp018green_out_predrv_0.nmos_6p0_CDNS_4066195314519_2.S.n5 GF_NI_IN_C_BASE_0.comp018green_out_predrv_0.nmos_6p0_CDNS_4066195314519_2.S.t2 34.4148
R53890 GF_NI_IN_C_BASE_0.comp018green_out_predrv_0.nmos_6p0_CDNS_4066195314519_2.S.n2 GF_NI_IN_C_BASE_0.comp018green_out_predrv_0.nmos_6p0_CDNS_4066195314519_2.S.t7 34.4148
R53891 GF_NI_IN_C_BASE_0.comp018green_out_predrv_0.nmos_6p0_CDNS_4066195314519_2.S.n4 GF_NI_IN_C_BASE_0.comp018green_out_predrv_0.nmos_6p0_CDNS_4066195314519_2.S.t3 34.4148
R53892 GF_NI_IN_C_BASE_0.comp018green_out_predrv_0.nmos_6p0_CDNS_4066195314519_2.S.n3 GF_NI_IN_C_BASE_0.comp018green_out_predrv_0.nmos_6p0_CDNS_4066195314519_2.S.t5 34.4148
R53893 GF_NI_IN_C_BASE_0.comp018green_out_predrv_0.nmos_6p0_CDNS_4066195314519_2.S.n5 GF_NI_IN_C_BASE_0.comp018green_out_predrv_0.nmos_6p0_CDNS_4066195314519_2.S.n4 10.9956
R53894 GF_NI_IN_C_BASE_0.comp018green_out_predrv_0.nmos_6p0_CDNS_4066195314519_2.S.n4 GF_NI_IN_C_BASE_0.comp018green_out_predrv_0.nmos_6p0_CDNS_4066195314519_2.S.n3 10.9956
R53895 GF_NI_IN_C_BASE_0.comp018green_out_predrv_0.nmos_6p0_CDNS_4066195314519_2.S.n3 GF_NI_IN_C_BASE_0.comp018green_out_predrv_0.nmos_6p0_CDNS_4066195314519_2.S.n2 10.9956
R53896 GF_NI_IN_C_BASE_0.comp018green_out_predrv_0.nmos_6p0_CDNS_4066195314519_2.S.n6 GF_NI_IN_C_BASE_0.comp018green_out_predrv_0.nmos_6p0_CDNS_4066195314519_2.S.n5 9.95826
R53897 GF_NI_IN_C_BASE_0.comp018green_out_predrv_0.nmos_6p0_CDNS_4066195314519_2.S.n2 GF_NI_IN_C_BASE_0.comp018green_out_predrv_0.nmos_6p0_CDNS_4066195314519_2.S.n1 8.49628
R53898 GF_NI_IN_C_BASE_0.comp018green_out_predrv_0.nmos_6p0_CDNS_4066195314519_2.S.n0 GF_NI_IN_C_BASE_0.comp018green_out_predrv_0.nmos_6p0_CDNS_4066195314519_2.S.t0 2.12938
R53899 GF_NI_IN_C_BASE_0.comp018green_out_predrv_0.nmos_6p0_CDNS_4066195314519_2.S.n0 GF_NI_IN_C_BASE_0.comp018green_out_predrv_0.nmos_6p0_CDNS_4066195314519_2.S.t1 1.97771
R53900 GF_NI_IN_C_BASE_0.comp018green_out_predrv_0.nmos_6p0_CDNS_4066195314519_2.S.n6 GF_NI_IN_C_BASE_0.comp018green_out_predrv_0.nmos_6p0_CDNS_4066195314519_2.S.n0 1.32326
R53901 GF_NI_IN_C_BASE_0.comp018green_out_predrv_0.nmos_6p0_CDNS_4066195314519_2.S GF_NI_IN_C_BASE_0.comp018green_out_predrv_0.nmos_6p0_CDNS_4066195314519_2.S.n6 1.25751
R53902 GF_NI_IN_C_BASE_0.ndrive_y_<0> GF_NI_IN_C_BASE_0.ndrive_y_<0>.t5 90.6729
R53903 GF_NI_IN_C_BASE_0.ndrive_y_<0>.n1 GF_NI_IN_C_BASE_0.ndrive_y_<0>.t3 5.90425
R53904 GF_NI_IN_C_BASE_0.ndrive_y_<0>.n2 GF_NI_IN_C_BASE_0.ndrive_y_<0> 3.52102
R53905 GF_NI_IN_C_BASE_0.ndrive_y_<0>.n4 GF_NI_IN_C_BASE_0.ndrive_y_<0>.t1 2.41832
R53906 GF_NI_IN_C_BASE_0.ndrive_y_<0>.n1 GF_NI_IN_C_BASE_0.ndrive_y_<0> 1.5749
R53907 GF_NI_IN_C_BASE_0.ndrive_y_<0>.n3 GF_NI_IN_C_BASE_0.ndrive_y_<0>.n2 1.48076
R53908 GF_NI_IN_C_BASE_0.ndrive_y_<0>.n0 GF_NI_IN_C_BASE_0.ndrive_y_<0>.n4 1.48076
R53909 GF_NI_IN_C_BASE_0.ndrive_y_<0>.n3 GF_NI_IN_C_BASE_0.ndrive_y_<0>.n1 1.09118
R53910 GF_NI_IN_C_BASE_0.ndrive_y_<0> GF_NI_IN_C_BASE_0.ndrive_y_<0>.n0 0.9455
R53911 GF_NI_IN_C_BASE_0.ndrive_y_<0>.n4 GF_NI_IN_C_BASE_0.ndrive_y_<0>.n3 0.578395
R53912 GF_NI_IN_C_BASE_0.ndrive_y_<0> GF_NI_IN_C_BASE_0.ndrive_y_<0>.t0 0.500893
R53913 GF_NI_IN_C_BASE_0.ndrive_y_<0>.n2 GF_NI_IN_C_BASE_0.ndrive_y_<0>.t4 0.360167
R53914 GF_NI_IN_C_BASE_0.ndrive_y_<0>.n0 GF_NI_IN_C_BASE_0.ndrive_y_<0>.t2 0.360167
R53915 GF_NI_IN_C_BASE_0.pdrive_x_<0>.n2 GF_NI_IN_C_BASE_0.pdrive_x_<0>.t4 113.251
R53916 GF_NI_IN_C_BASE_0.pdrive_x_<0>.n2 GF_NI_IN_C_BASE_0.pdrive_x_<0>.t5 112.769
R53917 GF_NI_IN_C_BASE_0.pdrive_x_<0>.t2 GF_NI_IN_C_BASE_0.pdrive_x_<0>.n1 6.12025
R53918 GF_NI_IN_C_BASE_0.pdrive_x_<0> GF_NI_IN_C_BASE_0.pdrive_x_<0>.n2 2.39
R53919 GF_NI_IN_C_BASE_0.pdrive_x_<0>.t3 GF_NI_IN_C_BASE_0.pdrive_x_<0>.n1 2.26404
R53920 GF_NI_IN_C_BASE_0.pdrive_x_<0> GF_NI_IN_C_BASE_0.pdrive_x_<0>.n0 1.4357
R53921 GF_NI_IN_C_BASE_0.pdrive_x_<0>.n1 GF_NI_IN_C_BASE_0.pdrive_x_<0>.n0 1.03582
R53922 GF_NI_IN_C_BASE_0.pdrive_x_<0> GF_NI_IN_C_BASE_0.pdrive_x_<0>.t0 0.779294
R53923 GF_NI_IN_C_BASE_0.pdrive_x_<0> GF_NI_IN_C_BASE_0.pdrive_x_<0>.t3 0.7466
R53924 GF_NI_IN_C_BASE_0.pdrive_x_<0>.n0 GF_NI_IN_C_BASE_0.pdrive_x_<0>.t1 0.66992
R53925 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_2.nmos_6p0_CDNS_4066195314530_0.D.n1 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_2.nmos_6p0_CDNS_4066195314530_0.D.t4 37.5434
R53926 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_2.nmos_6p0_CDNS_4066195314530_0.D.n0 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_2.nmos_6p0_CDNS_4066195314530_0.D.t5 37.5434
R53927 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_2.nmos_6p0_CDNS_4066195314530_0.D.n1 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_2.nmos_6p0_CDNS_4066195314530_0.D.t2 25.3941
R53928 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_2.nmos_6p0_CDNS_4066195314530_0.D.n0 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_2.nmos_6p0_CDNS_4066195314530_0.D.t3 25.3941
R53929 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_2.nmos_6p0_CDNS_4066195314530_0.D.n1 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_2.nmos_6p0_CDNS_4066195314530_0.D.n0 8.44221
R53930 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_2.nmos_6p0_CDNS_4066195314530_0.D.t1 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_2.nmos_6p0_CDNS_4066195314530_0.D.n1 4.90922
R53931 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_2.nmos_6p0_CDNS_4066195314530_0.D.t1 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_2.nmos_6p0_CDNS_4066195314530_0.D.t0 2.6373
R53932 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_pupd_0.PU_B.n1 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_pupd_0.PU_B.t3 37.5434
R53933 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_pupd_0.PU_B.n0 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_pupd_0.PU_B.t4 37.5434
R53934 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_pupd_0.PU_B GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_pupd_0.PU_B.t2 26.1617
R53935 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_pupd_0.PU_B.n1 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_pupd_0.PU_B.t5 25.3941
R53936 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_pupd_0.PU_B.n0 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_pupd_0.PU_B.t6 25.3941
R53937 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_pupd_0.PU_B.n1 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_pupd_0.PU_B.n0 8.44221
R53938 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_pupd_0.PU_B GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_pupd_0.PU_B.n1 4.40816
R53939 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_pupd_0.PU_B GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_pupd_0.PU_B.t1 2.2999
R53940 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_pupd_0.PU_B GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_pupd_0.PU_B.t0 2.0632
R53941 GF_NI_IN_C_BASE_0.comp018green_out_predrv_0.nmos_6p0_CDNS_4066195314519_0.D.n1 GF_NI_IN_C_BASE_0.comp018green_out_predrv_0.nmos_6p0_CDNS_4066195314519_0.D.t4 80.4772
R53942 GF_NI_IN_C_BASE_0.comp018green_out_predrv_0.nmos_6p0_CDNS_4066195314519_0.D.n0 GF_NI_IN_C_BASE_0.comp018green_out_predrv_0.nmos_6p0_CDNS_4066195314519_0.D.t3 80.4772
R53943 GF_NI_IN_C_BASE_0.comp018green_out_predrv_0.nmos_6p0_CDNS_4066195314519_0.D.n1 GF_NI_IN_C_BASE_0.comp018green_out_predrv_0.nmos_6p0_CDNS_4066195314519_0.D.t8 62.5719
R53944 GF_NI_IN_C_BASE_0.comp018green_out_predrv_0.nmos_6p0_CDNS_4066195314519_0.D.n0 GF_NI_IN_C_BASE_0.comp018green_out_predrv_0.nmos_6p0_CDNS_4066195314519_0.D.t7 62.5719
R53945 GF_NI_IN_C_BASE_0.comp018green_out_predrv_0.nmos_6p0_CDNS_4066195314519_0.D.n4 GF_NI_IN_C_BASE_0.comp018green_out_predrv_0.nmos_6p0_CDNS_4066195314519_0.D.t5 45.4098
R53946 GF_NI_IN_C_BASE_0.comp018green_out_predrv_0.nmos_6p0_CDNS_4066195314519_0.D.n4 GF_NI_IN_C_BASE_0.comp018green_out_predrv_0.nmos_6p0_CDNS_4066195314519_0.D.t6 34.4148
R53947 GF_NI_IN_C_BASE_0.comp018green_out_predrv_0.nmos_6p0_CDNS_4066195314519_0.D.n2 GF_NI_IN_C_BASE_0.comp018green_out_predrv_0.nmos_6p0_CDNS_4066195314519_0.D.n1 8.06816
R53948 GF_NI_IN_C_BASE_0.comp018green_out_predrv_0.nmos_6p0_CDNS_4066195314519_0.D.n2 GF_NI_IN_C_BASE_0.comp018green_out_predrv_0.nmos_6p0_CDNS_4066195314519_0.D.n0 8.06816
R53949 GF_NI_IN_C_BASE_0.comp018green_out_predrv_0.nmos_6p0_CDNS_4066195314519_0.D.n3 GF_NI_IN_C_BASE_0.comp018green_out_predrv_0.nmos_6p0_CDNS_4066195314519_0.D.n2 6.31953
R53950 GF_NI_IN_C_BASE_0.comp018green_out_predrv_0.nmos_6p0_CDNS_4066195314519_0.D.t0 GF_NI_IN_C_BASE_0.comp018green_out_predrv_0.nmos_6p0_CDNS_4066195314519_0.D.n4 6.08116
R53951 GF_NI_IN_C_BASE_0.comp018green_out_predrv_0.nmos_6p0_CDNS_4066195314519_0.D.t2 GF_NI_IN_C_BASE_0.comp018green_out_predrv_0.nmos_6p0_CDNS_4066195314519_0.D.n3 4.80357
R53952 GF_NI_IN_C_BASE_0.comp018green_out_predrv_0.nmos_6p0_CDNS_4066195314519_0.D.n3 GF_NI_IN_C_BASE_0.comp018green_out_predrv_0.nmos_6p0_CDNS_4066195314519_0.D.t1 4.54043
R53953 GF_NI_IN_C_BASE_0.comp018green_out_predrv_0.nmos_6p0_CDNS_4066195314519_0.D.t2 GF_NI_IN_C_BASE_0.comp018green_out_predrv_0.nmos_6p0_CDNS_4066195314519_0.D.t0 1.1409
R53954 GF_NI_IN_C_BASE_0.comp018green_out_predrv_0.nmos_6p0_CDNS_4066195314519_0.D.t0 GF_NI_IN_C_BASE_0.comp018green_out_predrv_0.nmos_6p0_CDNS_4066195314519_0.D 0.702585
R53955 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_0.Z.n0 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_0.Z.t4 37.5434
R53956 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_0.Z.n1 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_0.Z.t3 37.5434
R53957 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_0.Z.n0 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_0.Z.t2 25.3941
R53958 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_0.Z.n1 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_0.Z.t5 25.3941
R53959 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_0.Z.n1 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_0.Z.n0 8.44221
R53960 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_0.nmos_6p0_CDNS_4066195314531_1.D GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_0.Z.n1 4.40816
R53961 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_0.nmos_6p0_CDNS_4066195314531_1.D GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_0.Z.t1 2.2762
R53962 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_0.Z.t0 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_0.nmos_6p0_CDNS_4066195314531_1.D 2.08654
R53963 GF_NI_IN_C_BASE_0.comp018green_out_predrv_2.nmos_6p0_CDNS_4066195314519_0.D.n1 GF_NI_IN_C_BASE_0.comp018green_out_predrv_2.nmos_6p0_CDNS_4066195314519_0.D.t4 80.4772
R53964 GF_NI_IN_C_BASE_0.comp018green_out_predrv_2.nmos_6p0_CDNS_4066195314519_0.D.n0 GF_NI_IN_C_BASE_0.comp018green_out_predrv_2.nmos_6p0_CDNS_4066195314519_0.D.t5 80.4772
R53965 GF_NI_IN_C_BASE_0.comp018green_out_predrv_2.nmos_6p0_CDNS_4066195314519_0.D.n1 GF_NI_IN_C_BASE_0.comp018green_out_predrv_2.nmos_6p0_CDNS_4066195314519_0.D.t3 62.5719
R53966 GF_NI_IN_C_BASE_0.comp018green_out_predrv_2.nmos_6p0_CDNS_4066195314519_0.D.n0 GF_NI_IN_C_BASE_0.comp018green_out_predrv_2.nmos_6p0_CDNS_4066195314519_0.D.t8 62.5719
R53967 GF_NI_IN_C_BASE_0.comp018green_out_predrv_2.nmos_6p0_CDNS_4066195314519_0.D.n4 GF_NI_IN_C_BASE_0.comp018green_out_predrv_2.nmos_6p0_CDNS_4066195314519_0.D.t6 45.4098
R53968 GF_NI_IN_C_BASE_0.comp018green_out_predrv_2.nmos_6p0_CDNS_4066195314519_0.D.n4 GF_NI_IN_C_BASE_0.comp018green_out_predrv_2.nmos_6p0_CDNS_4066195314519_0.D.t7 34.4148
R53969 GF_NI_IN_C_BASE_0.comp018green_out_predrv_2.nmos_6p0_CDNS_4066195314519_0.D.n2 GF_NI_IN_C_BASE_0.comp018green_out_predrv_2.nmos_6p0_CDNS_4066195314519_0.D.n1 8.06816
R53970 GF_NI_IN_C_BASE_0.comp018green_out_predrv_2.nmos_6p0_CDNS_4066195314519_0.D.n2 GF_NI_IN_C_BASE_0.comp018green_out_predrv_2.nmos_6p0_CDNS_4066195314519_0.D.n0 8.06816
R53971 GF_NI_IN_C_BASE_0.comp018green_out_predrv_2.nmos_6p0_CDNS_4066195314519_0.D.n3 GF_NI_IN_C_BASE_0.comp018green_out_predrv_2.nmos_6p0_CDNS_4066195314519_0.D.n2 6.31953
R53972 GF_NI_IN_C_BASE_0.comp018green_out_predrv_2.nmos_6p0_CDNS_4066195314519_0.D.t2 GF_NI_IN_C_BASE_0.comp018green_out_predrv_2.nmos_6p0_CDNS_4066195314519_0.D.n4 6.08116
R53973 GF_NI_IN_C_BASE_0.comp018green_out_predrv_2.nmos_6p0_CDNS_4066195314519_0.D.t1 GF_NI_IN_C_BASE_0.comp018green_out_predrv_2.nmos_6p0_CDNS_4066195314519_0.D.n3 4.80357
R53974 GF_NI_IN_C_BASE_0.comp018green_out_predrv_2.nmos_6p0_CDNS_4066195314519_0.D.n3 GF_NI_IN_C_BASE_0.comp018green_out_predrv_2.nmos_6p0_CDNS_4066195314519_0.D.t0 4.54043
R53975 GF_NI_IN_C_BASE_0.comp018green_out_predrv_2.nmos_6p0_CDNS_4066195314519_0.D.t1 GF_NI_IN_C_BASE_0.comp018green_out_predrv_2.nmos_6p0_CDNS_4066195314519_0.D.t2 1.1409
R53976 GF_NI_IN_C_BASE_0.comp018green_out_predrv_2.nmos_6p0_CDNS_4066195314519_0.D.t2 GF_NI_IN_C_BASE_0.comp018green_out_predrv_2.nmos_6p0_CDNS_4066195314519_0.D 0.702585
R53977 GF_NI_IN_C_BASE_0.pdrive_y_<2> GF_NI_IN_C_BASE_0.pdrive_y_<2>.t4 115.388
R53978 GF_NI_IN_C_BASE_0.pdrive_y_<2>.t1 GF_NI_IN_C_BASE_0.pdrive_y_<2>.n1 6.10848
R53979 GF_NI_IN_C_BASE_0.pdrive_y_<2>.n0 GF_NI_IN_C_BASE_0.pdrive_y_<2>.n1 2.68197
R53980 GF_NI_IN_C_BASE_0.pdrive_y_<2>.n2 GF_NI_IN_C_BASE_0.pdrive_y_<2> 1.59856
R53981 GF_NI_IN_C_BASE_0.pdrive_y_<2>.n2 GF_NI_IN_C_BASE_0.pdrive_y_<2> 0.780424
R53982 GF_NI_IN_C_BASE_0.pdrive_y_<2> GF_NI_IN_C_BASE_0.pdrive_y_<2>.n0 0.7304
R53983 GF_NI_IN_C_BASE_0.pdrive_y_<2>.t2 GF_NI_IN_C_BASE_0.pdrive_y_<2> 0.500893
R53984 GF_NI_IN_C_BASE_0.pdrive_y_<2> GF_NI_IN_C_BASE_0.pdrive_y_<2>.t0 0.494197
R53985 GF_NI_IN_C_BASE_0.pdrive_y_<2>.n0 GF_NI_IN_C_BASE_0.pdrive_y_<2>.t3 0.360167
R53986 GF_NI_IN_C_BASE_0.pdrive_y_<2>.n1 GF_NI_IN_C_BASE_0.pdrive_y_<2>.n2 0.336519
R53987 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_cms_smt_0.nmos_6p0_CDNS_4066195314537_0.D.t1 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_cms_smt_0.nmos_6p0_CDNS_4066195314537_0.D.n2 4.05318
R53988 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_cms_smt_0.nmos_6p0_CDNS_4066195314537_0.D GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_cms_smt_0.nmos_6p0_CDNS_4066195314537_0.D.n1 1.23426
R53989 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_cms_smt_0.nmos_6p0_CDNS_4066195314537_0.D GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_cms_smt_0.nmos_6p0_CDNS_4066195314537_0.D.n0 1.23426
R53990 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_cms_smt_0.nmos_6p0_CDNS_4066195314537_0.D GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_cms_smt_0.nmos_6p0_CDNS_4066195314537_0.D.n2 1.10335
R53991 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_cms_smt_0.nmos_6p0_CDNS_4066195314537_0.D GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_cms_smt_0.nmos_6p0_CDNS_4066195314537_0.D.t0 1.02238
R53992 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_cms_smt_0.nmos_6p0_CDNS_4066195314537_0.D GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_cms_smt_0.nmos_6p0_CDNS_4066195314537_0.D.t2 1.02224
R53993 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_cms_smt_0.nmos_6p0_CDNS_4066195314537_0.D.n2 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_cms_smt_0.nmos_6p0_CDNS_4066195314537_0.D 0.943559
R53994 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_cms_smt_0.nmos_6p0_CDNS_4066195314537_0.D.n1 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_cms_smt_0.nmos_6p0_CDNS_4066195314537_0.D.t6 0.618613
R53995 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_cms_smt_0.nmos_6p0_CDNS_4066195314537_0.D.n1 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_cms_smt_0.nmos_6p0_CDNS_4066195314537_0.D.t4 0.618613
R53996 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_cms_smt_0.nmos_6p0_CDNS_4066195314537_0.D.n0 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_cms_smt_0.nmos_6p0_CDNS_4066195314537_0.D.t3 0.618613
R53997 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_cms_smt_0.nmos_6p0_CDNS_4066195314537_0.D.n0 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_cms_smt_0.nmos_6p0_CDNS_4066195314537_0.D.t5 0.618613
R53998 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_3.Z.n3 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_3.Z.t7 40.5676
R53999 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_3.Z.n2 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_3.Z.t11 40.5676
R54000 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_3.Z.n5 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_3.Z.t3 37.5434
R54001 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_3.Z.n4 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_3.Z.t12 37.5434
R54002 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_3.Z.n5 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_3.Z.t9 25.3941
R54003 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_3.Z.n4 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_3.Z.t4 25.3941
R54004 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_3.Z.n3 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_3.Z.t6 24.8726
R54005 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_3.Z.n2 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_3.Z.t10 24.8726
R54006 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_3.Z.n0 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_3.Z.t5 22.3127
R54007 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_3.Z.n0 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_3.Z.t1 21.9898
R54008 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_3.Z.n1 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_3.Z.t8 20.6262
R54009 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_3.Z.n1 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_3.Z.t2 20.1126
R54010 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_3.Z.n5 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_3.Z.n4 8.44221
R54011 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_3.Z.n0 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_3.Z.n1 6.88071
R54012 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_3.Z GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_3.Z.n0 6.22439
R54013 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_3.Z GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_3.Z.n5 4.40816
R54014 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_3.Z GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_3.Z.n3 4.09994
R54015 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_3.Z GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_3.Z.n2 4.03661
R54016 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_3.Z GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_3.Z.t0 2.75597
R54017 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_cms_smt_0.nmos_6p0_CDNS_4066195314536_1.S.n0 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_cms_smt_0.nmos_6p0_CDNS_4066195314536_1.S.t4 14.2306
R54018 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_cms_smt_0.nmos_6p0_CDNS_4066195314536_1.S.n0 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_cms_smt_0.nmos_6p0_CDNS_4066195314536_1.S.t3 13.9076
R54019 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_cms_smt_0.nmos_6p0_CDNS_4066195314536_1.S.n1 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_cms_smt_0.nmos_6p0_CDNS_4066195314536_1.S.t2 11.6919
R54020 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_cms_smt_0.nmos_6p0_CDNS_4066195314536_1.S.n1 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_cms_smt_0.nmos_6p0_CDNS_4066195314536_1.S.t1 4.40522
R54021 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_cms_smt_0.nmos_6p0_CDNS_4066195314536_1.S.n0 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_cms_smt_0.nmos_6p0_CDNS_4066195314536_1.S.t0 4.13853
R54022 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_cms_smt_0.nmos_6p0_CDNS_4066195314536_1.S.n1 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_cms_smt_0.nmos_6p0_CDNS_4066195314536_1.S.n0 4.13772
R54023 GF_NI_IN_C_BASE_0.comp018green_out_predrv_1.nmos_6p0_CDNS_4066195314519_2.S.n1 GF_NI_IN_C_BASE_0.comp018green_out_predrv_1.nmos_6p0_CDNS_4066195314519_2.S.t5 79.0838
R54024 GF_NI_IN_C_BASE_0.comp018green_out_predrv_1.nmos_6p0_CDNS_4066195314519_2.S.n1 GF_NI_IN_C_BASE_0.comp018green_out_predrv_1.nmos_6p0_CDNS_4066195314519_2.S.t2 78.041
R54025 GF_NI_IN_C_BASE_0.comp018green_out_predrv_1.nmos_6p0_CDNS_4066195314519_2.S.n5 GF_NI_IN_C_BASE_0.comp018green_out_predrv_1.nmos_6p0_CDNS_4066195314519_2.S.t7 34.4148
R54026 GF_NI_IN_C_BASE_0.comp018green_out_predrv_1.nmos_6p0_CDNS_4066195314519_2.S.n2 GF_NI_IN_C_BASE_0.comp018green_out_predrv_1.nmos_6p0_CDNS_4066195314519_2.S.t6 34.4148
R54027 GF_NI_IN_C_BASE_0.comp018green_out_predrv_1.nmos_6p0_CDNS_4066195314519_2.S.n3 GF_NI_IN_C_BASE_0.comp018green_out_predrv_1.nmos_6p0_CDNS_4066195314519_2.S.t3 34.4148
R54028 GF_NI_IN_C_BASE_0.comp018green_out_predrv_1.nmos_6p0_CDNS_4066195314519_2.S.n4 GF_NI_IN_C_BASE_0.comp018green_out_predrv_1.nmos_6p0_CDNS_4066195314519_2.S.t4 34.4148
R54029 GF_NI_IN_C_BASE_0.comp018green_out_predrv_1.nmos_6p0_CDNS_4066195314519_2.S.n3 GF_NI_IN_C_BASE_0.comp018green_out_predrv_1.nmos_6p0_CDNS_4066195314519_2.S.n2 10.9956
R54030 GF_NI_IN_C_BASE_0.comp018green_out_predrv_1.nmos_6p0_CDNS_4066195314519_2.S.n4 GF_NI_IN_C_BASE_0.comp018green_out_predrv_1.nmos_6p0_CDNS_4066195314519_2.S.n3 10.9956
R54031 GF_NI_IN_C_BASE_0.comp018green_out_predrv_1.nmos_6p0_CDNS_4066195314519_2.S.n5 GF_NI_IN_C_BASE_0.comp018green_out_predrv_1.nmos_6p0_CDNS_4066195314519_2.S.n4 10.9956
R54032 GF_NI_IN_C_BASE_0.comp018green_out_predrv_1.nmos_6p0_CDNS_4066195314519_2.S.n6 GF_NI_IN_C_BASE_0.comp018green_out_predrv_1.nmos_6p0_CDNS_4066195314519_2.S.n5 9.95826
R54033 GF_NI_IN_C_BASE_0.comp018green_out_predrv_1.nmos_6p0_CDNS_4066195314519_2.S.n2 GF_NI_IN_C_BASE_0.comp018green_out_predrv_1.nmos_6p0_CDNS_4066195314519_2.S.n1 8.49628
R54034 GF_NI_IN_C_BASE_0.comp018green_out_predrv_1.nmos_6p0_CDNS_4066195314519_2.S.n0 GF_NI_IN_C_BASE_0.comp018green_out_predrv_1.nmos_6p0_CDNS_4066195314519_2.S.t0 2.12938
R54035 GF_NI_IN_C_BASE_0.comp018green_out_predrv_1.nmos_6p0_CDNS_4066195314519_2.S.n0 GF_NI_IN_C_BASE_0.comp018green_out_predrv_1.nmos_6p0_CDNS_4066195314519_2.S.t1 1.97771
R54036 GF_NI_IN_C_BASE_0.comp018green_out_predrv_1.nmos_6p0_CDNS_4066195314519_2.S.n6 GF_NI_IN_C_BASE_0.comp018green_out_predrv_1.nmos_6p0_CDNS_4066195314519_2.S.n0 1.32326
R54037 GF_NI_IN_C_BASE_0.comp018green_out_predrv_1.nmos_6p0_CDNS_4066195314519_2.S GF_NI_IN_C_BASE_0.comp018green_out_predrv_1.nmos_6p0_CDNS_4066195314519_2.S.n6 1.25751
R54038 GF_NI_IN_C_BASE_0.ndrive_Y_<3> GF_NI_IN_C_BASE_0.ndrive_Y_<3>.t5 89.3064
R54039 GF_NI_IN_C_BASE_0.ndrive_Y_<3>.n1 GF_NI_IN_C_BASE_0.ndrive_Y_<3>.t3 5.90425
R54040 GF_NI_IN_C_BASE_0.ndrive_Y_<3>.n3 GF_NI_IN_C_BASE_0.ndrive_Y_<3>.t1 2.41832
R54041 GF_NI_IN_C_BASE_0.ndrive_Y_<3>.n2 GF_NI_IN_C_BASE_0.ndrive_Y_<3>.t4 1.84043
R54042 GF_NI_IN_C_BASE_0.ndrive_Y_<3>.n1 GF_NI_IN_C_BASE_0.ndrive_Y_<3> 1.5749
R54043 GF_NI_IN_C_BASE_0.ndrive_Y_<3>.n0 GF_NI_IN_C_BASE_0.ndrive_Y_<3>.n3 1.48076
R54044 GF_NI_IN_C_BASE_0.ndrive_Y_<3>.n2 GF_NI_IN_C_BASE_0.ndrive_Y_<3>.n1 1.09118
R54045 GF_NI_IN_C_BASE_0.ndrive_Y_<3> GF_NI_IN_C_BASE_0.ndrive_Y_<3>.n0 0.9455
R54046 GF_NI_IN_C_BASE_0.ndrive_Y_<3>.n3 GF_NI_IN_C_BASE_0.ndrive_Y_<3>.n2 0.578395
R54047 GF_NI_IN_C_BASE_0.ndrive_Y_<3> GF_NI_IN_C_BASE_0.ndrive_Y_<3>.t0 0.500893
R54048 GF_NI_IN_C_BASE_0.ndrive_Y_<3>.n0 GF_NI_IN_C_BASE_0.ndrive_Y_<3>.t2 0.360167
R54049 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_pupd_0.ppolyf_u_CDNS_4066195314533_1.PLUS.t0 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_pupd_0.ppolyf_u_CDNS_4066195314533_1.PLUS 11.0117
R54050 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_pupd_0.ppolyf_u_CDNS_4066195314533_1.PLUS GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_pupd_0.ppolyf_u_CDNS_4066195314533_1.PLUS.t1 11.0117
R54051 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_pupd_0.ppolyf_u_CDNS_4066195314533_1.MINUS.t0 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_pupd_0.ppolyf_u_CDNS_4066195314533_1.MINUS.t1 22.3936
R54052 GF_NI_IN_C_BASE_0.comp018green_out_predrv_3.nmos_6p0_CDNS_4066195314519_0.D.n1 GF_NI_IN_C_BASE_0.comp018green_out_predrv_3.nmos_6p0_CDNS_4066195314519_0.D.t8 80.4772
R54053 GF_NI_IN_C_BASE_0.comp018green_out_predrv_3.nmos_6p0_CDNS_4066195314519_0.D.n0 GF_NI_IN_C_BASE_0.comp018green_out_predrv_3.nmos_6p0_CDNS_4066195314519_0.D.t3 80.4772
R54054 GF_NI_IN_C_BASE_0.comp018green_out_predrv_3.nmos_6p0_CDNS_4066195314519_0.D.n1 GF_NI_IN_C_BASE_0.comp018green_out_predrv_3.nmos_6p0_CDNS_4066195314519_0.D.t6 62.5719
R54055 GF_NI_IN_C_BASE_0.comp018green_out_predrv_3.nmos_6p0_CDNS_4066195314519_0.D.n0 GF_NI_IN_C_BASE_0.comp018green_out_predrv_3.nmos_6p0_CDNS_4066195314519_0.D.t4 62.5719
R54056 GF_NI_IN_C_BASE_0.comp018green_out_predrv_3.nmos_6p0_CDNS_4066195314519_0.D.n4 GF_NI_IN_C_BASE_0.comp018green_out_predrv_3.nmos_6p0_CDNS_4066195314519_0.D.t5 45.4098
R54057 GF_NI_IN_C_BASE_0.comp018green_out_predrv_3.nmos_6p0_CDNS_4066195314519_0.D.n4 GF_NI_IN_C_BASE_0.comp018green_out_predrv_3.nmos_6p0_CDNS_4066195314519_0.D.t7 34.4148
R54058 GF_NI_IN_C_BASE_0.comp018green_out_predrv_3.nmos_6p0_CDNS_4066195314519_0.D.n2 GF_NI_IN_C_BASE_0.comp018green_out_predrv_3.nmos_6p0_CDNS_4066195314519_0.D.n1 8.06816
R54059 GF_NI_IN_C_BASE_0.comp018green_out_predrv_3.nmos_6p0_CDNS_4066195314519_0.D.n2 GF_NI_IN_C_BASE_0.comp018green_out_predrv_3.nmos_6p0_CDNS_4066195314519_0.D.n0 8.06816
R54060 GF_NI_IN_C_BASE_0.comp018green_out_predrv_3.nmos_6p0_CDNS_4066195314519_0.D.n3 GF_NI_IN_C_BASE_0.comp018green_out_predrv_3.nmos_6p0_CDNS_4066195314519_0.D.n2 6.31953
R54061 GF_NI_IN_C_BASE_0.comp018green_out_predrv_3.nmos_6p0_CDNS_4066195314519_0.D.t2 GF_NI_IN_C_BASE_0.comp018green_out_predrv_3.nmos_6p0_CDNS_4066195314519_0.D.n4 6.08116
R54062 GF_NI_IN_C_BASE_0.comp018green_out_predrv_3.nmos_6p0_CDNS_4066195314519_0.D.t0 GF_NI_IN_C_BASE_0.comp018green_out_predrv_3.nmos_6p0_CDNS_4066195314519_0.D.n3 4.80357
R54063 GF_NI_IN_C_BASE_0.comp018green_out_predrv_3.nmos_6p0_CDNS_4066195314519_0.D.n3 GF_NI_IN_C_BASE_0.comp018green_out_predrv_3.nmos_6p0_CDNS_4066195314519_0.D.t1 4.54043
R54064 GF_NI_IN_C_BASE_0.comp018green_out_predrv_3.nmos_6p0_CDNS_4066195314519_0.D.t0 GF_NI_IN_C_BASE_0.comp018green_out_predrv_3.nmos_6p0_CDNS_4066195314519_0.D.t2 1.1409
R54065 GF_NI_IN_C_BASE_0.comp018green_out_predrv_3.nmos_6p0_CDNS_4066195314519_0.D.t2 GF_NI_IN_C_BASE_0.comp018green_out_predrv_3.nmos_6p0_CDNS_4066195314519_0.D 0.702557
R54066 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_3.nmos_6p0_CDNS_4066195314530_0.D.n1 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_3.nmos_6p0_CDNS_4066195314530_0.D.t5 37.5434
R54067 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_3.nmos_6p0_CDNS_4066195314530_0.D.n0 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_3.nmos_6p0_CDNS_4066195314530_0.D.t3 37.5434
R54068 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_3.nmos_6p0_CDNS_4066195314530_0.D.n1 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_3.nmos_6p0_CDNS_4066195314530_0.D.t2 25.3941
R54069 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_3.nmos_6p0_CDNS_4066195314530_0.D.n0 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_3.nmos_6p0_CDNS_4066195314530_0.D.t4 25.3941
R54070 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_3.nmos_6p0_CDNS_4066195314530_0.D.n1 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_3.nmos_6p0_CDNS_4066195314530_0.D.n0 8.44221
R54071 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_3.nmos_6p0_CDNS_4066195314530_0.D.t1 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_3.nmos_6p0_CDNS_4066195314530_0.D.n1 4.90922
R54072 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_3.nmos_6p0_CDNS_4066195314530_0.D.t1 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_3.nmos_6p0_CDNS_4066195314530_0.D.t0 2.6373
R54073 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_pupd_0.PD GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_pupd_0.PD.t2 24.9619
R54074 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_pupd_0.PD GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_pupd_0.PD.t1 2.39238
R54075 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_pupd_0.PD GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_pupd_0.PD.t0 2.0632
R54076 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_cms_smt_0.nmos_6p0_CDNS_4066195314530_0.D GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_cms_smt_0.nmos_6p0_CDNS_4066195314530_0.D.t2 19.4535
R54077 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_cms_smt_0.nmos_6p0_CDNS_4066195314530_0.D GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_cms_smt_0.nmos_6p0_CDNS_4066195314530_0.D.t1 13.1326
R54078 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_cms_smt_0.nmos_6p0_CDNS_4066195314530_0.D.n0 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_cms_smt_0.nmos_6p0_CDNS_4066195314530_0.D.t0 8.30501
R54079 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_cms_smt_0.nmos_6p0_CDNS_4066195314530_0.D.n0 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_cms_smt_0.nmos_6p0_CDNS_4066195314530_0.D.t0 8.14999
R54080 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_cms_smt_0.nmos_6p0_CDNS_4066195314530_0.D GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_cms_smt_0.nmos_6p0_CDNS_4066195314530_0.D.n0 5.61641
R54081 GF_NI_IN_C_BASE_0.ndrive_x_<3> GF_NI_IN_C_BASE_0.ndrive_x_<3>.t3 90.7152
R54082 GF_NI_IN_C_BASE_0.ndrive_x_<3>.n0 GF_NI_IN_C_BASE_0.ndrive_x_<3>.n1 7.28458
R54083 GF_NI_IN_C_BASE_0.ndrive_x_<3>.n1 GF_NI_IN_C_BASE_0.ndrive_x_<3>.t1 6.03391
R54084 GF_NI_IN_C_BASE_0.ndrive_x_<3>.n1 GF_NI_IN_C_BASE_0.ndrive_x_<3> 1.45646
R54085 GF_NI_IN_C_BASE_0.ndrive_x_<3> GF_NI_IN_C_BASE_0.ndrive_x_<3>.n0 0.951421
R54086 GF_NI_IN_C_BASE_0.ndrive_x_<3>.t0 GF_NI_IN_C_BASE_0.ndrive_x_<3> 0.500893
R54087 GF_NI_IN_C_BASE_0.ndrive_x_<3>.n0 GF_NI_IN_C_BASE_0.ndrive_x_<3>.t2 0.360167
R54088 GF_NI_IN_C_BASE_0.ndrive_y_<2> GF_NI_IN_C_BASE_0.ndrive_y_<2>.t5 90.9292
R54089 GF_NI_IN_C_BASE_0.ndrive_y_<2>.n1 GF_NI_IN_C_BASE_0.ndrive_y_<2> 12.0008
R54090 GF_NI_IN_C_BASE_0.ndrive_y_<2>.n0 GF_NI_IN_C_BASE_0.ndrive_y_<2>.t0 5.90425
R54091 GF_NI_IN_C_BASE_0.ndrive_y_<2>.n3 GF_NI_IN_C_BASE_0.ndrive_y_<2>.t4 2.41832
R54092 GF_NI_IN_C_BASE_0.ndrive_y_<2>.n0 GF_NI_IN_C_BASE_0.ndrive_y_<2> 1.5749
R54093 GF_NI_IN_C_BASE_0.ndrive_y_<2>.n4 GF_NI_IN_C_BASE_0.ndrive_y_<2>.n3 1.48076
R54094 GF_NI_IN_C_BASE_0.ndrive_y_<2>.n2 GF_NI_IN_C_BASE_0.ndrive_y_<2>.n1 1.48076
R54095 GF_NI_IN_C_BASE_0.ndrive_y_<2>.n2 GF_NI_IN_C_BASE_0.ndrive_y_<2>.n0 1.09118
R54096 GF_NI_IN_C_BASE_0.ndrive_y_<2> GF_NI_IN_C_BASE_0.ndrive_y_<2>.n4 0.9455
R54097 GF_NI_IN_C_BASE_0.ndrive_y_<2>.n3 GF_NI_IN_C_BASE_0.ndrive_y_<2>.n2 0.578395
R54098 GF_NI_IN_C_BASE_0.ndrive_y_<2> GF_NI_IN_C_BASE_0.ndrive_y_<2>.t3 0.500893
R54099 GF_NI_IN_C_BASE_0.ndrive_y_<2>.n4 GF_NI_IN_C_BASE_0.ndrive_y_<2>.t1 0.360167
R54100 GF_NI_IN_C_BASE_0.ndrive_y_<2>.n1 GF_NI_IN_C_BASE_0.ndrive_y_<2>.t2 0.360167
R54101 GF_NI_IN_C_BASE_0.ndrive_x_<1> GF_NI_IN_C_BASE_0.ndrive_x_<1>.t3 90.8824
R54102 GF_NI_IN_C_BASE_0.ndrive_x_<1>.n0 GF_NI_IN_C_BASE_0.ndrive_x_<1>.n1 7.28458
R54103 GF_NI_IN_C_BASE_0.ndrive_x_<1>.n1 GF_NI_IN_C_BASE_0.ndrive_x_<1>.t0 6.03391
R54104 GF_NI_IN_C_BASE_0.ndrive_x_<1>.n1 GF_NI_IN_C_BASE_0.ndrive_x_<1> 1.45646
R54105 GF_NI_IN_C_BASE_0.ndrive_x_<1> GF_NI_IN_C_BASE_0.ndrive_x_<1>.n0 0.951421
R54106 GF_NI_IN_C_BASE_0.ndrive_x_<1>.t1 GF_NI_IN_C_BASE_0.ndrive_x_<1> 0.500893
R54107 GF_NI_IN_C_BASE_0.ndrive_x_<1>.n0 GF_NI_IN_C_BASE_0.ndrive_x_<1>.t2 0.360167
R54108 GF_NI_IN_C_BASE_0.pdrive_y_<0> GF_NI_IN_C_BASE_0.pdrive_y_<0>.t4 115.13
R54109 GF_NI_IN_C_BASE_0.pdrive_y_<0>.t1 GF_NI_IN_C_BASE_0.pdrive_y_<0>.n1 6.10848
R54110 GF_NI_IN_C_BASE_0.pdrive_y_<0>.n0 GF_NI_IN_C_BASE_0.pdrive_y_<0>.n1 2.68197
R54111 GF_NI_IN_C_BASE_0.pdrive_y_<0>.n2 GF_NI_IN_C_BASE_0.pdrive_y_<0> 1.59856
R54112 GF_NI_IN_C_BASE_0.pdrive_y_<0>.n2 GF_NI_IN_C_BASE_0.pdrive_y_<0> 0.780424
R54113 GF_NI_IN_C_BASE_0.pdrive_y_<0> GF_NI_IN_C_BASE_0.pdrive_y_<0>.n0 0.7304
R54114 GF_NI_IN_C_BASE_0.pdrive_y_<0>.t2 GF_NI_IN_C_BASE_0.pdrive_y_<0> 0.500893
R54115 GF_NI_IN_C_BASE_0.pdrive_y_<0> GF_NI_IN_C_BASE_0.pdrive_y_<0>.t0 0.494197
R54116 GF_NI_IN_C_BASE_0.pdrive_y_<0>.n0 GF_NI_IN_C_BASE_0.pdrive_y_<0>.t3 0.360167
R54117 GF_NI_IN_C_BASE_0.pdrive_y_<0>.n1 GF_NI_IN_C_BASE_0.pdrive_y_<0>.n2 0.336519
R54118 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_1.nmos_6p0_CDNS_4066195314531_0.D GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_1.ZB.t1 2.36868
R54119 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_1.nmos_6p0_CDNS_4066195314531_0.D GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_1.ZB.t0 2.08654
R54120 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_logic_pupd_0.comp018green_std_nand2_1.nmos_6p0_CDNS_4066195314511_1.S GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_logic_pupd_0.comp018green_std_nand2_1.nmos_6p0_CDNS_4066195314511_0.D.n0 1.15854
R54121 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_logic_pupd_0.comp018green_std_nand2_1.nmos_6p0_CDNS_4066195314511_0.D.n0 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_logic_pupd_0.comp018green_std_nand2_1.nmos_6p0_CDNS_4066195314511_0.D.t1 0.5465
R54122 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_logic_pupd_0.comp018green_std_nand2_1.nmos_6p0_CDNS_4066195314511_0.D.n0 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_logic_pupd_0.comp018green_std_nand2_1.nmos_6p0_CDNS_4066195314511_0.D.t0 0.5465
R54123 a_5575_62984.t0 a_5575_62984.n2 4.28715
R54124 a_5575_62984.n3 a_5575_62984.t5 5.32188
R54125 a_5575_62984.t1 a_5575_62984.n0 4.29256
R54126 a_5575_62984.n3 a_5575_62984.n1 2.84024
R54127 a_5575_62984.t4 a_5575_62984.n0 1.30198
R54128 a_5575_62984.n1 a_5575_62984.n2 0.00322045
R54129 a_5575_62984.n1 a_5575_62984.t3 2.34839
R54130 a_5575_62984.n0 a_5575_62984.n3 2.28727
R54131 a_5575_62984.n2 a_5575_62984.t2 8.1298
R54132 GF_NI_IN_C_BASE_0.comp018green_sigbuf_1_0.nmos_6p0_CDNS_4066195314530_0.D.n0 GF_NI_IN_C_BASE_0.comp018green_sigbuf_1_0.nmos_6p0_CDNS_4066195314530_0.D.t4 37.5434
R54133 GF_NI_IN_C_BASE_0.comp018green_sigbuf_1_0.nmos_6p0_CDNS_4066195314530_0.D.n1 GF_NI_IN_C_BASE_0.comp018green_sigbuf_1_0.nmos_6p0_CDNS_4066195314530_0.D.t5 37.5434
R54134 GF_NI_IN_C_BASE_0.comp018green_sigbuf_1_0.nmos_6p0_CDNS_4066195314530_0.D.n0 GF_NI_IN_C_BASE_0.comp018green_sigbuf_1_0.nmos_6p0_CDNS_4066195314530_0.D.t2 25.3941
R54135 GF_NI_IN_C_BASE_0.comp018green_sigbuf_1_0.nmos_6p0_CDNS_4066195314530_0.D.n1 GF_NI_IN_C_BASE_0.comp018green_sigbuf_1_0.nmos_6p0_CDNS_4066195314530_0.D.t3 25.3941
R54136 GF_NI_IN_C_BASE_0.comp018green_sigbuf_1_0.nmos_6p0_CDNS_4066195314530_0.D.n1 GF_NI_IN_C_BASE_0.comp018green_sigbuf_1_0.nmos_6p0_CDNS_4066195314530_0.D.n0 8.44221
R54137 GF_NI_IN_C_BASE_0.comp018green_sigbuf_1_0.nmos_6p0_CDNS_4066195314530_0.D.t1 GF_NI_IN_C_BASE_0.comp018green_sigbuf_1_0.nmos_6p0_CDNS_4066195314530_0.D.n1 4.93097
R54138 GF_NI_IN_C_BASE_0.comp018green_sigbuf_1_0.nmos_6p0_CDNS_4066195314530_0.D.t1 GF_NI_IN_C_BASE_0.comp018green_sigbuf_1_0.nmos_6p0_CDNS_4066195314530_0.D.t0 2.6373
R54139 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_logic_pupd_0.PUB_OUT.n0 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_logic_pupd_0.PUB_OUT.t3 35.9269
R54140 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_logic_pupd_0.PUB_OUT.n0 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_logic_pupd_0.PUB_OUT.t2 30.9212
R54141 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_logic_pupd_0.PUB_OUT.t0 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_2.A 23.5268
R54142 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_2.A GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_logic_pupd_0.PUB_OUT.n0 4.0005
R54143 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_logic_pupd_0.PUB_OUT.t0 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_logic_pupd_0.PUB_OUT.t1 3.23447
R54144 GF_NI_IN_C_BASE_0.pdrive_x_<3>.n3 GF_NI_IN_C_BASE_0.pdrive_x_<3>.t5 113.317
R54145 GF_NI_IN_C_BASE_0.pdrive_x_<3>.n3 GF_NI_IN_C_BASE_0.pdrive_x_<3>.t4 112.746
R54146 GF_NI_IN_C_BASE_0.pdrive_x_<3>.t2 GF_NI_IN_C_BASE_0.pdrive_x_<3>.n1 6.12025
R54147 GF_NI_IN_C_BASE_0.pdrive_x_<3> GF_NI_IN_C_BASE_0.pdrive_x_<3>.n3 2.39
R54148 GF_NI_IN_C_BASE_0.pdrive_x_<3>.n0 GF_NI_IN_C_BASE_0.pdrive_x_<3>.n1 2.26404
R54149 GF_NI_IN_C_BASE_0.pdrive_x_<3>.n2 GF_NI_IN_C_BASE_0.pdrive_x_<3> 1.43572
R54150 GF_NI_IN_C_BASE_0.pdrive_x_<3>.n1 GF_NI_IN_C_BASE_0.pdrive_x_<3>.n2 1.0357
R54151 GF_NI_IN_C_BASE_0.pdrive_x_<3> GF_NI_IN_C_BASE_0.pdrive_x_<3>.t1 0.779435
R54152 GF_NI_IN_C_BASE_0.pdrive_x_<3> GF_NI_IN_C_BASE_0.pdrive_x_<3>.n0 0.7466
R54153 GF_NI_IN_C_BASE_0.pdrive_x_<3>.t0 GF_NI_IN_C_BASE_0.pdrive_x_<3>.n2 0.396936
R54154 GF_NI_IN_C_BASE_0.pdrive_x_<3>.n0 GF_NI_IN_C_BASE_0.pdrive_x_<3>.t3 0.360167
R54155 GF_NI_IN_C_BASE_0.pdrive_y_<3> GF_NI_IN_C_BASE_0.pdrive_y_<3>.t4 115.088
R54156 GF_NI_IN_C_BASE_0.pdrive_y_<3>.t1 GF_NI_IN_C_BASE_0.pdrive_y_<3>.n1 6.10848
R54157 GF_NI_IN_C_BASE_0.pdrive_y_<3>.n0 GF_NI_IN_C_BASE_0.pdrive_y_<3>.n1 2.68197
R54158 GF_NI_IN_C_BASE_0.pdrive_y_<3>.n2 GF_NI_IN_C_BASE_0.pdrive_y_<3> 1.59857
R54159 GF_NI_IN_C_BASE_0.pdrive_y_<3>.n2 GF_NI_IN_C_BASE_0.pdrive_y_<3> 0.781133
R54160 GF_NI_IN_C_BASE_0.pdrive_y_<3> GF_NI_IN_C_BASE_0.pdrive_y_<3>.n0 0.7304
R54161 GF_NI_IN_C_BASE_0.pdrive_y_<3> GF_NI_IN_C_BASE_0.pdrive_y_<3>.t2 0.500875
R54162 GF_NI_IN_C_BASE_0.pdrive_y_<3> GF_NI_IN_C_BASE_0.pdrive_y_<3>.t0 0.493858
R54163 GF_NI_IN_C_BASE_0.pdrive_y_<3>.n0 GF_NI_IN_C_BASE_0.pdrive_y_<3>.t3 0.360167
R54164 GF_NI_IN_C_BASE_0.pdrive_y_<3>.n1 GF_NI_IN_C_BASE_0.pdrive_y_<3>.n2 0.336519
R54165 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_3.nmos_6p0_CDNS_4066195314531_0.D GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_3.ZB.t1 2.36868
R54166 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_3.nmos_6p0_CDNS_4066195314531_0.D GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_3.ZB.t0 2.08654
R54167 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.ENB GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.ENB.t2 82.1164
R54168 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.ENB GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.ENB.t3 42.2319
R54169 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.ENB GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.ENB.t0 2.04837
R54170 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.ENB GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.ENB.t1 1.49421
R54171 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_cms_smt_0.nmos_6p0_CDNS_4066195314535_0.D.n1 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_cms_smt_0.nmos_6p0_CDNS_4066195314535_0.D.t2 22.8162
R54172 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_cms_smt_0.nmos_6p0_CDNS_4066195314535_0.D.n1 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_cms_smt_0.nmos_6p0_CDNS_4066195314535_0.D.t4 22.3026
R54173 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_cms_smt_0.nmos_6p0_CDNS_4066195314535_0.D.n0 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_cms_smt_0.nmos_6p0_CDNS_4066195314535_0.D.t3 20.1892
R54174 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_cms_smt_0.nmos_6p0_CDNS_4066195314535_0.D.n0 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_cms_smt_0.nmos_6p0_CDNS_4066195314535_0.D.n1 11.9677
R54175 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_cms_smt_0.nmos_6p0_CDNS_4066195314535_0.D GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_cms_smt_0.nmos_6p0_CDNS_4066195314535_0.D.t0 1.55917
R54176 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_cms_smt_0.nmos_6p0_CDNS_4066195314535_0.D.n0 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_cms_smt_0.nmos_6p0_CDNS_4066195314535_0.D.t1 1.45173
R54177 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_cms_smt_0.nmos_6p0_CDNS_4066195314535_0.D GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_cms_smt_0.nmos_6p0_CDNS_4066195314535_0.D.n0 1.38831
R54178 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_pupd_0.ppolyf_u_CDNS_4066195314533_2.PLUS.t1 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_pupd_0.ppolyf_u_CDNS_4066195314533_2.PLUS.t0 22.3936
R54179 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_pupd_0.ppolyf_u_CDNS_4066195314533_5.MINUS.n0 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_pupd_0.ppolyf_u_CDNS_4066195314533_5.MINUS.n1 3.11956
R54180 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_pupd_0.ppolyf_u_CDNS_4066195314533_5.MINUS.t0 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_pupd_0.ppolyf_u_CDNS_4066195314533_5.MINUS.n0 2.91689
R54181 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_pupd_0.ppolyf_u_CDNS_4066195314533_5.MINUS GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_pupd_0.ppolyf_u_CDNS_4066195314533_5.MINUS.n0 0.0638785
R54182 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_pupd_0.ppolyf_u_CDNS_4066195314533_5.MINUS GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_pupd_0.ppolyf_u_CDNS_4066195314533_5.MINUS.n2 0.055602
R54183 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_pupd_0.ppolyf_u_CDNS_4066195314533_5.MINUS.n2 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_pupd_0.ppolyf_u_CDNS_4066195314533_5.MINUS.n1 6.35009
R54184 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_pupd_0.ppolyf_u_CDNS_4066195314533_5.MINUS GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_pupd_0.ppolyf_u_CDNS_4066195314533_5.MINUS.n2 11.9543
R54185 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_pupd_0.ppolyf_u_CDNS_4066195314533_5.MINUS.t2 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_pupd_0.ppolyf_u_CDNS_4066195314533_5.MINUS 11.0117
R54186 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_pupd_0.ppolyf_u_CDNS_4066195314533_5.MINUS.n1 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_pupd_0.ppolyf_u_CDNS_4066195314533_5.MINUS.t1 1.0925
R54187 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_a_0.nmos_6p0_CDNS_4066195314511_3.S.n0 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_a_0.nmos_6p0_CDNS_4066195314511_3.S.t3 44.3219
R54188 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_a_0.nmos_6p0_CDNS_4066195314511_3.S.n0 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_a_0.nmos_6p0_CDNS_4066195314511_3.S.t2 28.0534
R54189 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_a_0.nmos_6p0_CDNS_4066195314511_3.S GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_a_0.nmos_6p0_CDNS_4066195314511_3.S.n0 4.18151
R54190 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_a_0.nmos_6p0_CDNS_4066195314511_3.S GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_a_0.nmos_6p0_CDNS_4066195314511_3.S.t1 1.76195
R54191 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_a_0.nmos_6p0_CDNS_4066195314511_3.S GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_a_0.nmos_6p0_CDNS_4066195314511_3.S.t0 1.56963
R54192 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_2.nmos_6p0_CDNS_4066195314531_0.D GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_2.ZB.t1 2.36868
R54193 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_2.nmos_6p0_CDNS_4066195314531_0.D GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_2.ZB.t0 2.08654
R54194 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.EN GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.EN.t5 82.1164
R54195 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.EN.n0 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.EN.t4 44.3219
R54196 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.EN GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.EN.t2 42.2319
R54197 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.EN.n0 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.EN.t3 28.0534
R54198 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.EN GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.EN.n0 4.09808
R54199 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.EN GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.EN.t0 1.53534
R54200 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.EN GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.EN.t1 1.33388
R54201 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_2.nmos_6p0_CDNS_4066195314511_1.D GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_2.nmos_6p0_CDNS_4066195314511_0.S.n0 1.15854
R54202 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_2.nmos_6p0_CDNS_4066195314511_0.S.n0 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_2.nmos_6p0_CDNS_4066195314511_0.S.t1 0.5465
R54203 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_2.nmos_6p0_CDNS_4066195314511_0.S.n0 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_2.nmos_6p0_CDNS_4066195314511_0.S.t0 0.5465
R54204 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_2.nmos_6p0_CDNS_4066195314511_1.S.n0 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_2.nmos_6p0_CDNS_4066195314511_1.S.t3 38.8469
R54205 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_2.nmos_6p0_CDNS_4066195314511_1.S.n0 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_2.nmos_6p0_CDNS_4066195314511_1.S.t2 22.5262
R54206 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_2.nmos_6p0_CDNS_4066195314511_1.S.t0 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_2.nmos_6p0_CDNS_4066195314511_1.S.n0 12.9666
R54207 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_2.nmos_6p0_CDNS_4066195314511_1.S.t0 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_2.nmos_6p0_CDNS_4066195314511_1.S.t1 2.79762
R54208 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_1.ENB GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_1.ENB.t3 82.1164
R54209 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_1.ENB GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_1.ENB.t4 82.1164
R54210 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_1.ENB GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_1.ENB.t5 42.2319
R54211 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_1.ENB GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_1.ENB.t2 42.2319
R54212 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_1.ENB.n0 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_1.ENB 10.4346
R54213 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_1.ENB.n0 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_1.ENB 9.25386
R54214 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_1.ENB GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_1.ENB.n0 7.14721
R54215 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_1.ENB GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_1.ENB.t1 2.04837
R54216 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_1.ENB GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_1.ENB.t0 1.49421
R54217 PD.n5 PD.t3 35.5619
R54218 PD PD.t2 35.4693
R54219 PD.n5 PD.t4 34.9362
R54220 PD.n2 PD.t1 33.3819
R54221 PD.n3 PD.t0 28.9398
R54222 PD PD.n7 23.3129
R54223 PD.n2 PD.t5 16.3212
R54224 PD.n3 PD.n2 12.3062
R54225 PD.n1 PD 4.88182
R54226 PD.n7 PD.n4 4.73379
R54227 PD.n7 PD.n6 4.00668
R54228 PD PD.n3 4.00168
R54229 PD.n6 PD.n5 4.0005
R54230 PD.n4 PD 2.3055
R54231 PD.n1 PD.n0 2.25122
R54232 PD.n0 PD.t6 1.31518
R54233 PD PD.n1 0.4505
R54234 PD.n6 PD 0.00642105
R54235 PD.n4 PD 0.00405263
R54236 PD.n0 PD 0.001225
R54237 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.nmos_6p0_CDNS_4066195314511_1.D GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.nmos_6p0_CDNS_4066195314511_0.S.n0 1.15854
R54238 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.nmos_6p0_CDNS_4066195314511_0.S.t0 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.nmos_6p0_CDNS_4066195314511_0.S.n0 0.5465
R54239 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.nmos_6p0_CDNS_4066195314511_0.S.n0 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.nmos_6p0_CDNS_4066195314511_0.S.t1 0.5465
R54240 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_pupd_0.ppolyf_u_CDNS_4066195314533_4.PLUS.t0 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_pupd_0.ppolyf_u_CDNS_4066195314533_4.PLUS.t1 22.3936
R54241 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_logic_pupd_0.comp018green_std_nand2_0.nmos_6p0_CDNS_4066195314511_1.S GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_logic_pupd_0.comp018green_std_nand2_0.nmos_6p0_CDNS_4066195314511_0.D.n0 1.15854
R54242 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_logic_pupd_0.comp018green_std_nand2_0.nmos_6p0_CDNS_4066195314511_0.D.n0 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_logic_pupd_0.comp018green_std_nand2_0.nmos_6p0_CDNS_4066195314511_0.D.t1 0.5465
R54243 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_logic_pupd_0.comp018green_std_nand2_0.nmos_6p0_CDNS_4066195314511_0.D.n0 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_logic_pupd_0.comp018green_std_nand2_0.nmos_6p0_CDNS_4066195314511_0.D.t0 0.5465
R54244 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_pupd_0.ppolyf_u_CDNS_4066195314533_3.MINUS.t0 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_pupd_0.ppolyf_u_CDNS_4066195314533_3.MINUS 11.0117
R54245 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_pupd_0.ppolyf_u_CDNS_4066195314533_3.MINUS GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_pupd_0.ppolyf_u_CDNS_4066195314533_3.MINUS.t1 11.0117
C0 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_1.EN 0.31341f
C1 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_1.EN GF_NI_IN_C_BASE_0.pdrive_x_<2> 0.055041f
C2 GF_NI_IN_C_BASE_0.pdrive_y_<0> DVSS 2.40128f
C3 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE VDD 26.6474f
C4 GF_NI_IN_C_BASE_0.comp018green_out_predrv_0.SL GF_NI_IN_C_BASE_0.ndrive_x_<3> 0.864692f
C5 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_cms_smt_0.nmos_6p0_CDNS_4066195314537_0.D DVDD 6.16e-19
C6 GF_NI_IN_C_BASE_0.comp018green_out_predrv_1.EN GF_NI_IN_C_BASE_0.comp018green_out_predrv_1.nmos_6p0_CDNS_4066195314519_0.D 2.21816f
C7 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_cms_smt_0.nmos_6p0_CDNS_4066195314535_0.D PU 2.31e-19
C8 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.ENB GF_NI_IN_C_BASE_0.comp018green_out_predrv_0.SL 0.407297f
C9 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_pupd_0.PD VDD 0.595879f
C10 GF_NI_IN_C_BASE_0.comp018green_out_predrv_1.ENB GF_NI_IN_C_BASE_0.pdrive_x_<3> 6.39e-19
C11 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE GF_NI_IN_C_BASE_0.comp018green_out_predrv_1.ENB 0.024125f
C12 GF_NI_IN_C_BASE_0.pdrive_y_<1> DVDD 16.7876f
C13 GF_NI_IN_C_BASE_0.ndrive_y_<2> GF_NI_IN_C_BASE_0.pdrive_y_<2> 0.06919f
C14 GF_NI_IN_C_BASE_0.comp018green_out_predrv_3.nmos_6p0_CDNS_4066195314519_0.D DVDD 3.94638f
C15 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_cms_smt_0.nmos_6p0_CDNS_4066195314537_0.D GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_cms_smt_0.nmos_6p0_CDNS_4066195314540_0.S 1.03718f
C16 w_4468_53312# VDD 0.007089f
C17 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_1.EN GF_NI_IN_C_BASE_0.ndrive_x_<2> 0.003319f
C18 PU Y 0.228424f
C19 GF_NI_IN_C_BASE_0.comp018green_out_predrv_1.EN GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_a_0.nmos_6p0_CDNS_4066195314511_3.S 0.014957f
C20 DVDD PAD 0.31019p
C21 GF_NI_IN_C_BASE_0.comp018green_out_predrv_1.EN GF_NI_IN_C_BASE_0.comp018green_out_predrv_2.nmos_6p0_CDNS_4066195314519_2.S 6.5e-19
C22 GF_NI_IN_C_BASE_0.comp018green_out_predrv_1.ENB GF_NI_IN_C_BASE_0.ndrive_x_<2> 3.42e-19
C23 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.EN GF_NI_IN_C_BASE_0.pdrive_x_<0> 9.2e-19
C24 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_drv_0.nmos_6p0_CDNS_4066195314547_0.S VDD 1.49069f
C25 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_cms_smt_0.nmos_6p0_CDNS_4066195314530_0.D DVDD 0.09529f
C26 GF_NI_IN_C_BASE_0.comp018green_out_predrv_0.nmos_6p0_CDNS_4066195314519_2.S DVDD 5.46753f
C27 GF_NI_IN_C_BASE_0.comp018green_out_predrv_1.nmos_6p0_CDNS_4066195314519_2.S DVDD 5.6228f
C28 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_1.EN GF_NI_IN_C_BASE_0.pdrive_x_<1> 0.05515f
C29 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_cms_smt_0.nmos_6p0_CDNS_4066195314535_0.D PD 1.33e-19
C30 GF_NI_IN_C_BASE_0.pdrive_y_<3> PAD 10.1904f
C31 GF_NI_IN_C_BASE_0.comp018green_out_predrv_0.SL GF_NI_IN_C_BASE_0.ndrive_x_<1> 0.858187f
C32 DVDD DVSS 0.353198p
C33 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.EN GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_1.ENB 0.001515f
C34 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_cms_smt_0.nmos_6p0_CDNS_4066195314530_0.D GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_cms_smt_0.nmos_6p0_CDNS_4066195314540_0.S 0.395973f
C35 PD Y 1.13e-19
C36 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.EN GF_NI_IN_C_BASE_0.ndrive_x_<0> 0.002977f
C37 GF_NI_IN_C_BASE_0.comp018green_out_predrv_1.EN PAD 0.227696f
C38 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.ENB GF_NI_IN_C_BASE_0.comp018green_out_predrv_0.SLB 4.24e-20
C39 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_1.ENB VDD 0.136356f
C40 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_1.EN GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_1.ENB 5.44729f
C41 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_1.Z DVDD 3.50468f
C42 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_1.nmos_6p0_CDNS_4066195314511_1.S 0.991052f
C43 GF_NI_IN_C_BASE_0.comp018green_out_predrv_0.A GF_NI_IN_C_BASE_0.ndrive_Y_<1> 6.85e-19
C44 GF_NI_IN_C_BASE_0.comp018green_out_predrv_1.nmos_6p0_CDNS_4066195314519_0.D GF_NI_IN_C_BASE_0.comp018green_out_predrv_1.nmos_6p0_CDNS_4066195314519_2.S 1.90189f
C45 GF_NI_IN_C_BASE_0.comp018green_out_predrv_1.nmos_6p0_CDNS_4066195314519_2.S GF_NI_IN_C_BASE_0.pdrive_y_<3> 0.020536f
C46 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_a_0.nmos_6p0_CDNS_4066195314511_3.S PAD 0.005824f
C47 GF_NI_IN_C_BASE_0.comp018green_out_predrv_2.nmos_6p0_CDNS_4066195314519_2.S PAD 0.289643f
C48 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_cms_smt_0.nmos_6p0_CDNS_4066195314540_0.S DVSS 0.758941f
C49 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_pupd_0.PU_B GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_drv_0.A 0.001819f
C50 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_pupd_0.ppolyf_u_CDNS_4066195314533_0.PLUS 0.003198f
C51 GF_NI_IN_C_BASE_0.pdrive_y_<3> DVSS 2.51388f
C52 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_1.ENB GF_NI_IN_C_BASE_0.comp018green_out_predrv_1.ENB 0.002247f
C53 GF_NI_IN_C_BASE_0.comp018green_out_predrv_1.nmos_6p0_CDNS_4066195314519_0.D DVSS 4.61993f
C54 GF_NI_IN_C_BASE_0.comp018green_out_predrv_1.EN GF_NI_IN_C_BASE_0.comp018green_out_predrv_1.nmos_6p0_CDNS_4066195314519_2.S 2.30331f
C55 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_pupd_0.ppolyf_u_CDNS_4066195314533_5.MINUS PD 0.106114f
C56 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_1.Z GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_cms_smt_0.nmos_6p0_CDNS_4066195314540_0.S 0.001012f
C57 GF_NI_IN_C_BASE_0.comp018green_out_predrv_3.nmos_6p0_CDNS_4066195314519_0.D GF_NI_IN_C_BASE_0.pdrive_y_<1> 2.80754f
C58 GF_NI_IN_C_BASE_0.comp018green_out_predrv_3.nmos_6p0_CDNS_4066195314519_2.S DVDD 5.24558f
C59 GF_NI_IN_C_BASE_0.comp018green_out_predrv_1.EN DVSS 2.69014f
C60 GF_NI_IN_C_BASE_0.pdrive_y_<1> PAD 10.1967f
C61 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_cms_smt_0.nmos_6p0_CDNS_4066195314530_0.D GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_cms_smt_0.nmos_6p0_CDNS_4066195314537_0.D 0.178647f
C62 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_a_0.nmos_6p0_CDNS_4066195314511_3.S DVSS 0.733838f
C63 GF_NI_IN_C_BASE_0.comp018green_out_predrv_0.SL GF_NI_IN_C_BASE_0.comp018green_out_predrv_2.nmos_6p0_CDNS_4066195314519_0.D 0.01198f
C64 GF_NI_IN_C_BASE_0.comp018green_out_predrv_2.nmos_6p0_CDNS_4066195314519_2.S DVSS 2.81189f
C65 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.nmos_6p0_CDNS_4066195314511_1.S GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.ENB 0.013931f
C66 GF_NI_IN_C_BASE_0.ndrive_y_<0> GF_NI_IN_C_BASE_0.pdrive_y_<0> 2.38e-19
C67 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_cms_smt_0.nmos_6p0_CDNS_4066195314537_0.D DVSS 1.72154f
C68 GF_NI_IN_C_BASE_0.ndrive_y_<2> DVDD 11.7314f
C69 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_pupd_0.PD GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_drv_0.A 9.98e-19
C70 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_1.Z GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_cms_smt_0.nmos_6p0_CDNS_4066195314537_0.D 0.575641f
C71 DVDD PU 2.82121f
C72 GF_NI_IN_C_BASE_0.comp018green_out_predrv_3.nmos_6p0_CDNS_4066195314519_0.D DVSS 4.60391f
C73 GF_NI_IN_C_BASE_0.pdrive_y_<1> DVSS 2.57275f
C74 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_1.nmos_6p0_CDNS_4066195314511_1.S GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_1.ENB 0.013931f
C75 PAD DVSS 0.238705p
C76 GF_NI_IN_C_BASE_0.comp018green_out_predrv_3.nmos_6p0_CDNS_4066195314519_2.S GF_NI_IN_C_BASE_0.comp018green_out_predrv_2.nmos_6p0_CDNS_4066195314519_2.S 0.032032f
C77 GF_NI_IN_C_BASE_0.comp018green_out_predrv_1.ENB GF_NI_IN_C_BASE_0.ndrive_Y_<3> 0.360444f
C78 GF_NI_IN_C_BASE_0.ndrive_y_<2> GF_NI_IN_C_BASE_0.pdrive_y_<3> 0.069955f
C79 GF_NI_IN_C_BASE_0.ndrive_y_<2> GF_NI_IN_C_BASE_0.comp018green_out_predrv_1.nmos_6p0_CDNS_4066195314519_0.D 0.00245f
C80 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.EN GF_NI_IN_C_BASE_0.comp018green_out_predrv_0.A 0.328973f
C81 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_drv_0.A GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_drv_0.nmos_6p0_CDNS_4066195314547_0.S 0.520068f
C82 GF_NI_IN_C_BASE_0.comp018green_out_predrv_0.nmos_6p0_CDNS_4066195314519_2.S DVSS 2.84499f
C83 GF_NI_IN_C_BASE_0.comp018green_out_predrv_0.SL GF_NI_IN_C_BASE_0.comp018green_out_predrv_0.nmos_6p0_CDNS_4066195314519_0.D 0.01198f
C84 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_cms_smt_0.nmos_6p0_CDNS_4066195314530_0.D DVSS 2.02847f
C85 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_1.EN GF_NI_IN_C_BASE_0.comp018green_out_predrv_0.A 0.80907f
C86 GF_NI_IN_C_BASE_0.comp018green_out_predrv_0.A VDD 0.154321f
C87 GF_NI_IN_C_BASE_0.comp018green_out_predrv_1.nmos_6p0_CDNS_4066195314519_2.S DVSS 2.74665f
C88 GF_NI_IN_C_BASE_0.comp018green_out_predrv_0.SLB GF_NI_IN_C_BASE_0.comp018green_out_predrv_2.nmos_6p0_CDNS_4066195314519_0.D 0.026278f
C89 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE GF_NI_IN_C_BASE_0.comp018green_out_predrv_0.SL 0.027335f
C90 GF_NI_IN_C_BASE_0.comp018green_out_predrv_0.SL GF_NI_IN_C_BASE_0.pdrive_x_<2> 0.005985f
C91 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_a_0.nmos_6p0_CDNS_4066195314511_1.D 0.845232f
C92 GF_NI_IN_C_BASE_0.comp018green_out_predrv_1.EN GF_NI_IN_C_BASE_0.ndrive_y_<2> 6.12e-19
C93 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_1.Z GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_cms_smt_0.nmos_6p0_CDNS_4066195314530_0.D 0.316661f
C94 GF_NI_IN_C_BASE_0.comp018green_out_predrv_3.nmos_6p0_CDNS_4066195314519_2.S GF_NI_IN_C_BASE_0.pdrive_y_<1> 0.026792f
C95 DVDD PD 2.8238f
C96 GF_NI_IN_C_BASE_0.comp018green_out_predrv_3.nmos_6p0_CDNS_4066195314519_0.D GF_NI_IN_C_BASE_0.comp018green_out_predrv_3.nmos_6p0_CDNS_4066195314519_2.S 1.90189f
C97 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_logic_pupd_0.comp018green_std_xor2_0.nmos_6p0_CDNS_4066195314530_2.D VDD 0.74012f
C98 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.EN GF_NI_IN_C_BASE_0.ndrive_Y_<1> 3.42e-19
C99 GF_NI_IN_C_BASE_0.comp018green_out_predrv_1.ENB GF_NI_IN_C_BASE_0.comp018green_out_predrv_0.A 0.091634f
C100 GF_NI_IN_C_BASE_0.comp018green_out_predrv_2.nmos_6p0_CDNS_4066195314519_2.S GF_NI_IN_C_BASE_0.ndrive_y_<2> 1.8828f
C101 GF_NI_IN_C_BASE_0.ndrive_y_<0> DVDD 8.5375f
C102 GF_NI_IN_C_BASE_0.comp018green_out_predrv_3.nmos_6p0_CDNS_4066195314519_2.S PAD 0.289643f
C103 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_1.EN GF_NI_IN_C_BASE_0.ndrive_Y_<1> 3.42e-19
C104 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_1.Z DVSS 5.63042f
C105 GF_NI_IN_C_BASE_0.comp018green_out_predrv_0.SL GF_NI_IN_C_BASE_0.ndrive_x_<2> 0.861977f
C106 w_4468_53312# GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_a_0.nmos_6p0_CDNS_4066195314511_1.D 0.001239f
C107 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_3.Z 0.093529f
C108 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_pupd_0.ppolyf_u_CDNS_4066195314533_3.MINUS 0.065372f
C109 GF_NI_IN_C_BASE_0.comp018green_out_predrv_3.nmos_6p0_CDNS_4066195314519_2.S DVSS 2.74619f
C110 GF_NI_IN_C_BASE_0.ndrive_y_<2> PAD 6.37203f
C111 GF_NI_IN_C_BASE_0.comp018green_out_predrv_0.SL GF_NI_IN_C_BASE_0.pdrive_x_<1> 0.013839f
C112 GF_NI_IN_C_BASE_0.comp018green_out_predrv_0.SLB GF_NI_IN_C_BASE_0.comp018green_out_predrv_0.nmos_6p0_CDNS_4066195314519_0.D 0.024516f
C113 GF_NI_IN_C_BASE_0.comp018green_out_predrv_0.SLB GF_NI_IN_C_BASE_0.pdrive_x_<3> 0.544964f
C114 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE GF_NI_IN_C_BASE_0.comp018green_out_predrv_0.SLB 0.001199f
C115 GF_NI_IN_C_BASE_0.comp018green_out_predrv_0.SLB GF_NI_IN_C_BASE_0.pdrive_x_<2> 0.544964f
C116 GF_NI_IN_C_BASE_0.pdrive_y_<0> GF_NI_IN_C_BASE_0.ndrive_x_<1> 0.069442f
C117 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_pupd_0.ppolyf_u_CDNS_4066195314533_1.PLUS VDD 0.001237f
C118 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_cms_smt_0.nmos_6p0_CDNS_4066195314530_0.D PU 0.029892f
C119 GF_NI_IN_C_BASE_0.comp018green_out_predrv_2.nmos_6p0_CDNS_4066195314519_0.D GF_NI_IN_C_BASE_0.pdrive_y_<2> 2.80754f
C120 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_1.nmos_6p0_CDNS_4066195314511_1.S GF_NI_IN_C_BASE_0.comp018green_out_predrv_0.A 5.93e-20
C121 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_1.ENB GF_NI_IN_C_BASE_0.comp018green_out_predrv_0.SL 0.34223f
C122 GF_NI_IN_C_BASE_0.ndrive_x_<3> DVDD 5.84068f
C123 GF_NI_IN_C_BASE_0.comp018green_out_predrv_0.SL GF_NI_IN_C_BASE_0.ndrive_x_<0> 0.869906f
C124 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_3.Z GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_drv_0.nmos_6p0_CDNS_4066195314547_0.S 6.92e-19
C125 GF_NI_IN_C_BASE_0.ndrive_y_<2> DVSS 9.637599f
C126 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.ENB DVDD 1.30292f
C127 DVSS PU 6.57534f
C128 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_1.Z PU 0.05345f
C129 GF_NI_IN_C_BASE_0.comp018green_out_predrv_1.nmos_6p0_CDNS_4066195314519_0.D GF_NI_IN_C_BASE_0.ndrive_x_<3> 0.039995f
C130 GF_NI_IN_C_BASE_0.pdrive_y_<3> GF_NI_IN_C_BASE_0.ndrive_x_<3> 3.33e-19
C131 GF_NI_IN_C_BASE_0.ndrive_y_<0> PAD 5.88153f
C132 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.EN VDD 0.289021f
C133 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.EN GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_1.EN 0.011456f
C134 GF_NI_IN_C_BASE_0.comp018green_out_predrv_0.SLB GF_NI_IN_C_BASE_0.pdrive_x_<1> 0.544964f
C135 GF_NI_IN_C_BASE_0.comp018green_out_predrv_0.SLB GF_NI_IN_C_BASE_0.pdrive_x_<0> 0.544964f
C136 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.nmos_6p0_CDNS_4066195314511_1.S 0.991848f
C137 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_cms_smt_0.nmos_6p0_CDNS_4066195314530_0.D PD 0.011323f
C138 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_cms_smt_0.nmos_6p0_CDNS_4066195314535_0.D 0.003102f
C139 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_1.EN VDD 0.363481f
C140 GF_NI_IN_C_BASE_0.comp018green_out_predrv_1.EN GF_NI_IN_C_BASE_0.ndrive_x_<3> 0.007481f
C141 GF_NI_IN_C_BASE_0.comp018green_out_predrv_0.nmos_6p0_CDNS_4066195314519_2.S GF_NI_IN_C_BASE_0.ndrive_y_<0> 1.8897f
C142 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_pupd_0.PU_B GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_pupd_0.ppolyf_u_CDNS_4066195314533_5.MINUS 0.426986f
C143 GF_NI_IN_C_BASE_0.comp018green_out_predrv_3.nmos_6p0_CDNS_4066195314519_2.S GF_NI_IN_C_BASE_0.ndrive_y_<2> 3.7e-19
C144 GF_NI_IN_C_BASE_0.ndrive_x_<1> DVDD 9.37134f
C145 GF_NI_IN_C_BASE_0.pdrive_y_<2> GF_NI_IN_C_BASE_0.pdrive_x_<2> 2.31053f
C146 DVSS PD 6.40624f
C147 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_1.ENB GF_NI_IN_C_BASE_0.comp018green_out_predrv_0.SLB 0.077321f
C148 GF_NI_IN_C_BASE_0.comp018green_out_predrv_1.ENB VDD 0.136026f
C149 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_1.EN GF_NI_IN_C_BASE_0.comp018green_out_predrv_1.ENB 0.005324f
C150 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE Y 2.57356f
C151 GF_NI_IN_C_BASE_0.ndrive_y_<0> DVSS 12.1872f
C152 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_1.Z PD 0.046863f
C153 GF_NI_IN_C_BASE_0.comp018green_out_predrv_0.SL GF_NI_IN_C_BASE_0.ndrive_Y_<3> 1.11322f
C154 GF_NI_IN_C_BASE_0.ndrive_x_<2> GF_NI_IN_C_BASE_0.pdrive_y_<2> 0.465424f
C155 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_pupd_0.ppolyf_u_CDNS_4066195314533_5.MINUS 0.287174f
C156 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_pupd_0.ppolyf_u_CDNS_4066195314533_0.PLUS GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_pupd_0.ppolyf_u_CDNS_4066195314533_1.PLUS 0.034604f
C157 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_cms_smt_0.nmos_6p0_CDNS_4066195314535_0.D GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_drv_0.nmos_6p0_CDNS_4066195314547_0.S 7.55e-19
C158 GF_NI_IN_C_BASE_0.ndrive_x_<3> PAD 6.09734f
C159 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_pupd_0.PD GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_pupd_0.ppolyf_u_CDNS_4066195314533_5.MINUS 1.10297f
C160 GF_NI_IN_C_BASE_0.comp018green_out_predrv_0.A GF_NI_IN_C_BASE_0.comp018green_out_predrv_0.SL 8.486509f
C161 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_a_0.nmos_6p0_CDNS_4066195314511_1.D GF_NI_IN_C_BASE_0.comp018green_out_predrv_0.A 0.045759f
C162 GF_NI_IN_C_BASE_0.comp018green_out_predrv_0.nmos_6p0_CDNS_4066195314519_0.D GF_NI_IN_C_BASE_0.pdrive_y_<0> 2.92427f
C163 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_drv_0.nmos_6p0_CDNS_4066195314547_0.S Y 0.002641f
C164 GF_NI_IN_C_BASE_0.comp018green_out_predrv_1.nmos_6p0_CDNS_4066195314519_2.S GF_NI_IN_C_BASE_0.ndrive_x_<3> 1.76852f
C165 GF_NI_IN_C_BASE_0.comp018green_out_predrv_2.nmos_6p0_CDNS_4066195314519_0.D DVDD 3.94147f
C166 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.ENB GF_NI_IN_C_BASE_0.comp018green_out_predrv_0.nmos_6p0_CDNS_4066195314519_2.S 0.561221f
C167 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_1.nmos_6p0_CDNS_4066195314511_1.S VDD 1.20038f
C168 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_1.EN GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_1.nmos_6p0_CDNS_4066195314511_1.S 0.594367f
C169 GF_NI_IN_C_BASE_0.comp018green_out_predrv_0.SL GF_NI_IN_C_BASE_0.ndrive_Y_<1> 1.11846f
C170 GF_NI_IN_C_BASE_0.ndrive_x_<3> DVSS 12.0448f
C171 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_drv_0.nmos_6p0_CDNS_4066195314547_0.S GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_pupd_0.ppolyf_u_CDNS_4066195314533_5.MINUS 0.016985f
C172 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_pupd_0.ppolyf_u_CDNS_4066195314533_0.PLUS VDD 0.001144f
C173 PU PD 0.788434f
C174 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.ENB DVSS 2.66771f
C175 GF_NI_IN_C_BASE_0.pdrive_y_<1> GF_NI_IN_C_BASE_0.ndrive_x_<1> 0.069353f
C176 GF_NI_IN_C_BASE_0.comp018green_out_predrv_3.nmos_6p0_CDNS_4066195314519_0.D GF_NI_IN_C_BASE_0.ndrive_x_<1> 0.041607f
C177 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_pupd_0.PU_B DVDD 2.29092f
C178 GF_NI_IN_C_BASE_0.comp018green_out_predrv_2.nmos_6p0_CDNS_4066195314519_0.D GF_NI_IN_C_BASE_0.comp018green_out_predrv_1.nmos_6p0_CDNS_4066195314519_0.D 0.00366f
C179 GF_NI_IN_C_BASE_0.comp018green_out_predrv_2.nmos_6p0_CDNS_4066195314519_0.D GF_NI_IN_C_BASE_0.pdrive_y_<3> 0.02501f
C180 GF_NI_IN_C_BASE_0.ndrive_x_<1> PAD 5.87598f
C181 GF_NI_IN_C_BASE_0.comp018green_out_predrv_1.EN GF_NI_IN_C_BASE_0.comp018green_out_predrv_2.nmos_6p0_CDNS_4066195314519_0.D 2.31e-19
C182 GF_NI_IN_C_BASE_0.comp018green_out_predrv_0.A GF_NI_IN_C_BASE_0.comp018green_out_predrv_0.SLB 0.215003f
C183 GF_NI_IN_C_BASE_0.pdrive_y_<0> GF_NI_IN_C_BASE_0.pdrive_x_<0> 2.34844f
C184 GF_NI_IN_C_BASE_0.pdrive_y_<0> GF_NI_IN_C_BASE_0.pdrive_x_<1> 0.071453f
C185 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_drv_0.A VDD 0.655203f
C186 GF_NI_IN_C_BASE_0.comp018green_out_predrv_0.nmos_6p0_CDNS_4066195314519_0.D DVDD 4.0074f
C187 GF_NI_IN_C_BASE_0.comp018green_out_predrv_2.nmos_6p0_CDNS_4066195314519_2.S GF_NI_IN_C_BASE_0.comp018green_out_predrv_2.nmos_6p0_CDNS_4066195314519_0.D 1.90189f
C188 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE DVDD 24.3242f
C189 GF_NI_IN_C_BASE_0.pdrive_x_<2> DVDD 30.1606f
C190 GF_NI_IN_C_BASE_0.pdrive_x_<3> DVDD 29.843401f
C191 GF_NI_IN_C_BASE_0.ndrive_x_<1> DVSS 9.78923f
C192 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_pupd_0.PD DVDD 0.603095f
C193 GF_NI_IN_C_BASE_0.ndrive_x_<0> GF_NI_IN_C_BASE_0.pdrive_y_<0> 1.64e-19
C194 GF_NI_IN_C_BASE_0.comp018green_out_predrv_1.nmos_6p0_CDNS_4066195314519_0.D GF_NI_IN_C_BASE_0.pdrive_x_<3> 0.718047f
C195 GF_NI_IN_C_BASE_0.pdrive_x_<3> GF_NI_IN_C_BASE_0.pdrive_y_<3> 2.34446f
C196 GF_NI_IN_C_BASE_0.ndrive_y_<2> GF_NI_IN_C_BASE_0.ndrive_x_<3> 9.95829f
C197 GF_NI_IN_C_BASE_0.pdrive_x_<2> GF_NI_IN_C_BASE_0.pdrive_y_<3> 0.071453f
C198 GF_NI_IN_C_BASE_0.ndrive_x_<2> DVDD 15.290899f
C199 w_4468_53312# DVDD 3.90127f
C200 GF_NI_IN_C_BASE_0.pdrive_x_<2> GF_NI_IN_C_BASE_0.comp018green_out_predrv_1.nmos_6p0_CDNS_4066195314519_0.D 5.58e-20
C201 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.nmos_6p0_CDNS_4066195314511_1.S GF_NI_IN_C_BASE_0.comp018green_out_predrv_0.A 5.93e-20
C202 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.EN GF_NI_IN_C_BASE_0.comp018green_out_predrv_0.SL 0.051023f
C203 GF_NI_IN_C_BASE_0.comp018green_out_predrv_1.EN GF_NI_IN_C_BASE_0.pdrive_x_<3> 9.56e-19
C204 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE GF_NI_IN_C_BASE_0.comp018green_out_predrv_1.EN 0.032326f
C205 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_drv_0.nmos_6p0_CDNS_4066195314547_0.S DVDD 0.415966f
C206 GF_NI_IN_C_BASE_0.comp018green_out_predrv_0.SL VDD 0.646847f
C207 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_1.EN GF_NI_IN_C_BASE_0.comp018green_out_predrv_0.SL 0.08661f
C208 GF_NI_IN_C_BASE_0.comp018green_out_predrv_3.nmos_6p0_CDNS_4066195314519_2.S GF_NI_IN_C_BASE_0.ndrive_x_<1> 1.76505f
C209 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_a_0.nmos_6p0_CDNS_4066195314511_1.D VDD 1.29558f
C210 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_a_0.nmos_6p0_CDNS_4066195314511_3.S 0.001798f
C211 GF_NI_IN_C_BASE_0.ndrive_x_<2> GF_NI_IN_C_BASE_0.pdrive_y_<3> 0.158648f
C212 GF_NI_IN_C_BASE_0.ndrive_x_<2> GF_NI_IN_C_BASE_0.comp018green_out_predrv_1.nmos_6p0_CDNS_4066195314519_0.D 0.001369f
C213 GF_NI_IN_C_BASE_0.pdrive_x_<1> DVDD 30.2148f
C214 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE GF_NI_IN_C_BASE_0.comp018green_out_predrv_2.nmos_6p0_CDNS_4066195314519_2.S 0.001031f
C215 GF_NI_IN_C_BASE_0.comp018green_out_predrv_2.nmos_6p0_CDNS_4066195314519_2.S GF_NI_IN_C_BASE_0.pdrive_x_<2> 0.184422f
C216 GF_NI_IN_C_BASE_0.pdrive_x_<0> DVDD 29.688799f
C217 GF_NI_IN_C_BASE_0.comp018green_out_predrv_0.A GF_NI_IN_C_BASE_0.pdrive_y_<2> 0.06401f
C218 GF_NI_IN_C_BASE_0.comp018green_out_predrv_1.ENB GF_NI_IN_C_BASE_0.comp018green_out_predrv_0.SL 0.247434f
C219 GF_NI_IN_C_BASE_0.comp018green_out_predrv_1.ENB GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_a_0.nmos_6p0_CDNS_4066195314511_1.D 1.6e-19
C220 GF_NI_IN_C_BASE_0.comp018green_out_predrv_2.nmos_6p0_CDNS_4066195314519_0.D DVSS 4.60296f
C221 GF_NI_IN_C_BASE_0.comp018green_out_predrv_1.EN GF_NI_IN_C_BASE_0.ndrive_x_<2> 3.42e-19
C222 w_4468_53312# GF_NI_IN_C_BASE_0.comp018green_out_predrv_1.EN 0.001159f
C223 w_4468_53312# GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_a_0.nmos_6p0_CDNS_4066195314511_3.S 0.001239f
C224 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_1.ENB DVDD 1.73896f
C225 GF_NI_IN_C_BASE_0.comp018green_out_predrv_0.nmos_6p0_CDNS_4066195314519_0.D GF_NI_IN_C_BASE_0.comp018green_out_predrv_3.nmos_6p0_CDNS_4066195314519_0.D 0.00366f
C226 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE GF_NI_IN_C_BASE_0.comp018green_out_predrv_3.nmos_6p0_CDNS_4066195314519_0.D 0.001902f
C227 GF_NI_IN_C_BASE_0.comp018green_out_predrv_2.nmos_6p0_CDNS_4066195314519_2.S GF_NI_IN_C_BASE_0.ndrive_x_<2> 1.77749f
C228 GF_NI_IN_C_BASE_0.ndrive_x_<0> DVDD 7.912839f
C229 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_3.Z VDD 0.186935f
C230 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_pupd_0.PU_B DVSS 4.79611f
C231 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.ENB GF_NI_IN_C_BASE_0.ndrive_y_<0> 0.371612f
C232 GF_NI_IN_C_BASE_0.pdrive_x_<3> PAD 20.2053f
C233 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE PAD 1.52682f
C234 GF_NI_IN_C_BASE_0.pdrive_x_<2> PAD 20.8838f
C235 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_pupd_0.ppolyf_u_CDNS_4066195314533_3.MINUS VDD 8.14e-19
C236 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.EN GF_NI_IN_C_BASE_0.comp018green_out_predrv_0.SLB 5.97e-20
C237 GF_NI_IN_C_BASE_0.comp018green_out_predrv_0.nmos_6p0_CDNS_4066195314519_2.S GF_NI_IN_C_BASE_0.comp018green_out_predrv_0.nmos_6p0_CDNS_4066195314519_0.D 1.90189f
C238 GF_NI_IN_C_BASE_0.comp018green_out_predrv_0.SLB VDD 0.131856f
C239 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_1.EN GF_NI_IN_C_BASE_0.comp018green_out_predrv_0.SLB 0.088175f
C240 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE GF_NI_IN_C_BASE_0.comp018green_out_predrv_0.nmos_6p0_CDNS_4066195314519_2.S 0.0011f
C241 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_cms_smt_0.nmos_6p0_CDNS_4066195314530_0.D 0.016805f
C242 GF_NI_IN_C_BASE_0.comp018green_out_predrv_1.nmos_6p0_CDNS_4066195314519_2.S GF_NI_IN_C_BASE_0.pdrive_x_<3> 8.77e-19
C243 GF_NI_IN_C_BASE_0.comp018green_out_predrv_0.A GF_NI_IN_C_BASE_0.pdrive_y_<0> 0.055976f
C244 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_1.ENB GF_NI_IN_C_BASE_0.comp018green_out_predrv_1.EN 0.007733f
C245 w_4468_53312# PAD 1.7719f
C246 GF_NI_IN_C_BASE_0.ndrive_x_<2> PAD 7.42368f
C247 GF_NI_IN_C_BASE_0.comp018green_out_predrv_0.nmos_6p0_CDNS_4066195314519_0.D DVSS 4.60007f
C248 GF_NI_IN_C_BASE_0.comp018green_out_predrv_1.ENB GF_NI_IN_C_BASE_0.comp018green_out_predrv_0.SLB 0.211601f
C249 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_1.nmos_6p0_CDNS_4066195314511_1.S GF_NI_IN_C_BASE_0.comp018green_out_predrv_0.SL 4.94e-20
C250 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_1.ENB GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_a_0.nmos_6p0_CDNS_4066195314511_3.S 1.29e-20
C251 GF_NI_IN_C_BASE_0.pdrive_x_<3> DVSS 5.56609f
C252 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE DVSS 30.9421f
C253 GF_NI_IN_C_BASE_0.pdrive_x_<2> DVSS 4.80365f
C254 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_1.ENB GF_NI_IN_C_BASE_0.comp018green_out_predrv_2.nmos_6p0_CDNS_4066195314519_2.S 0.519126f
C255 GF_NI_IN_C_BASE_0.comp018green_out_predrv_3.nmos_6p0_CDNS_4066195314519_0.D GF_NI_IN_C_BASE_0.pdrive_x_<1> 0.86434f
C256 GF_NI_IN_C_BASE_0.pdrive_y_<0> GF_NI_IN_C_BASE_0.ndrive_Y_<1> 0.158279f
C257 GF_NI_IN_C_BASE_0.pdrive_x_<1> GF_NI_IN_C_BASE_0.pdrive_y_<1> 2.29406f
C258 GF_NI_IN_C_BASE_0.ndrive_y_<0> GF_NI_IN_C_BASE_0.ndrive_x_<1> 10.0071f
C259 GF_NI_IN_C_BASE_0.pdrive_x_<0> GF_NI_IN_C_BASE_0.comp018green_out_predrv_3.nmos_6p0_CDNS_4066195314519_0.D 5.58e-20
C260 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_1.Z 0.05398f
C261 GF_NI_IN_C_BASE_0.comp018green_out_predrv_2.nmos_6p0_CDNS_4066195314519_0.D GF_NI_IN_C_BASE_0.ndrive_y_<2> 1.2931f
C262 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_pupd_0.PD DVSS 2.0042f
C263 GF_NI_IN_C_BASE_0.ndrive_Y_<3> DVDD 12.3616f
C264 GF_NI_IN_C_BASE_0.pdrive_x_<0> PAD 20.2173f
C265 GF_NI_IN_C_BASE_0.pdrive_x_<1> PAD 20.890501f
C266 w_4468_53312# DVSS 0.22053f
C267 GF_NI_IN_C_BASE_0.ndrive_x_<2> DVSS 11.0547f
C268 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.nmos_6p0_CDNS_4066195314511_1.S GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.EN 0.594367f
C269 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_cms_smt_0.nmos_6p0_CDNS_4066195314530_0.D GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_drv_0.nmos_6p0_CDNS_4066195314547_0.S 6.63e-20
C270 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_1.ENB GF_NI_IN_C_BASE_0.comp018green_out_predrv_3.nmos_6p0_CDNS_4066195314519_0.D 2.42579f
C271 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_pupd_0.ppolyf_u_CDNS_4066195314533_5.MINUS GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_pupd_0.ppolyf_u_CDNS_4066195314533_1.PLUS 4.05e-19
C272 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.nmos_6p0_CDNS_4066195314511_1.S VDD 1.18218f
C273 GF_NI_IN_C_BASE_0.comp018green_out_predrv_0.nmos_6p0_CDNS_4066195314519_2.S GF_NI_IN_C_BASE_0.pdrive_x_<0> 8.77e-19
C274 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_pupd_0.PU_B PU 0.200243f
C275 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_cms_smt_0.nmos_6p0_CDNS_4066195314535_0.D VDD 0.227715f
C276 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_1.ENB PAD 0.1164f
C277 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_drv_0.nmos_6p0_CDNS_4066195314547_0.S DVSS 1.23422f
C278 GF_NI_IN_C_BASE_0.comp018green_out_predrv_1.nmos_6p0_CDNS_4066195314519_0.D GF_NI_IN_C_BASE_0.ndrive_Y_<3> 1.27008f
C279 GF_NI_IN_C_BASE_0.ndrive_x_<0> PAD 5.05035f
C280 GF_NI_IN_C_BASE_0.comp018green_out_predrv_0.A DVDD 3.82271f
C281 GF_NI_IN_C_BASE_0.pdrive_x_<1> DVSS 4.80778f
C282 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_1.EN GF_NI_IN_C_BASE_0.pdrive_y_<2> 0.004504f
C283 GF_NI_IN_C_BASE_0.pdrive_x_<0> DVSS 5.52502f
C284 VDD Y 1.79605f
C285 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_pupd_0.ppolyf_u_CDNS_4066195314533_3.MINUS GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_pupd_0.ppolyf_u_CDNS_4066195314533_0.PLUS 0.034604f
C286 GF_NI_IN_C_BASE_0.comp018green_out_predrv_0.nmos_6p0_CDNS_4066195314519_2.S GF_NI_IN_C_BASE_0.ndrive_x_<0> 1.79768f
C287 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_logic_pupd_0.comp018green_std_xor2_0.nmos_6p0_CDNS_4066195314530_2.D DVDD 0.171184f
C288 GF_NI_IN_C_BASE_0.ndrive_y_<2> GF_NI_IN_C_BASE_0.pdrive_x_<3> 0.074402f
C289 GF_NI_IN_C_BASE_0.ndrive_Y_<1> DVDD 17.769402f
C290 GF_NI_IN_C_BASE_0.ndrive_y_<2> GF_NI_IN_C_BASE_0.pdrive_x_<2> 0.217482f
C291 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_1.ENB DVSS 4.90648f
C292 GF_NI_IN_C_BASE_0.comp018green_out_predrv_0.A GF_NI_IN_C_BASE_0.comp018green_out_predrv_1.nmos_6p0_CDNS_4066195314519_0.D 0.491713f
C293 GF_NI_IN_C_BASE_0.comp018green_out_predrv_0.A GF_NI_IN_C_BASE_0.pdrive_y_<3> 0.055976f
C294 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE PU 5.05097f
C295 GF_NI_IN_C_BASE_0.ndrive_x_<0> DVSS 17.7576f
C296 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.ENB GF_NI_IN_C_BASE_0.ndrive_x_<1> 6.12e-19
C297 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_pupd_0.ppolyf_u_CDNS_4066195314533_5.MINUS VDD 1.53792f
C298 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_3.Z GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_drv_0.A 3.36825f
C299 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_pupd_0.PU_B PD 1.53932f
C300 GF_NI_IN_C_BASE_0.comp018green_out_predrv_1.EN GF_NI_IN_C_BASE_0.comp018green_out_predrv_0.A 0.835267f
C301 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_pupd_0.PD PU 0.052014f
C302 GF_NI_IN_C_BASE_0.comp018green_out_predrv_3.nmos_6p0_CDNS_4066195314519_2.S GF_NI_IN_C_BASE_0.pdrive_x_<1> 0.184422f
C303 GF_NI_IN_C_BASE_0.ndrive_x_<2> GF_NI_IN_C_BASE_0.ndrive_y_<2> 14.653599f
C304 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_a_0.nmos_6p0_CDNS_4066195314511_3.S GF_NI_IN_C_BASE_0.comp018green_out_predrv_0.A 0.5167f
C305 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_a_0.nmos_6p0_CDNS_4066195314511_1.D GF_NI_IN_C_BASE_0.comp018green_out_predrv_0.SL 4.94e-20
C306 GF_NI_IN_C_BASE_0.comp018green_out_predrv_0.A GF_NI_IN_C_BASE_0.comp018green_out_predrv_2.nmos_6p0_CDNS_4066195314519_2.S 1.67859f
C307 GF_NI_IN_C_BASE_0.ndrive_Y_<3> PAD 5.0955f
C308 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_1.ENB GF_NI_IN_C_BASE_0.comp018green_out_predrv_3.nmos_6p0_CDNS_4066195314519_2.S 0.562071f
C309 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE PD 4.86189f
C310 GF_NI_IN_C_BASE_0.comp018green_out_predrv_0.nmos_6p0_CDNS_4066195314519_0.D GF_NI_IN_C_BASE_0.ndrive_y_<0> 1.29246f
C311 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_pupd_0.ppolyf_u_CDNS_4066195314533_1.PLUS DVDD 0.373802f
C312 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_drv_0.nmos_6p0_CDNS_4066195314547_0.S PU 0.021163f
C313 GF_NI_IN_C_BASE_0.ndrive_Y_<1> GF_NI_IN_C_BASE_0.comp018green_out_predrv_2.nmos_6p0_CDNS_4066195314519_2.S 3.7e-19
C314 GF_NI_IN_C_BASE_0.comp018green_out_predrv_1.nmos_6p0_CDNS_4066195314519_2.S GF_NI_IN_C_BASE_0.ndrive_Y_<3> 1.92044f
C315 GF_NI_IN_C_BASE_0.comp018green_out_predrv_0.A GF_NI_IN_C_BASE_0.pdrive_y_<1> 0.064015f
C316 GF_NI_IN_C_BASE_0.comp018green_out_predrv_0.A GF_NI_IN_C_BASE_0.comp018green_out_predrv_3.nmos_6p0_CDNS_4066195314519_0.D 0.505117f
C317 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_pupd_0.PD PD 0.013731f
C318 GF_NI_IN_C_BASE_0.comp018green_out_predrv_0.A PAD 0.107351f
C319 GF_NI_IN_C_BASE_0.ndrive_Y_<3> DVSS 16.0763f
C320 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_1.ENB GF_NI_IN_C_BASE_0.ndrive_y_<2> 0.34647f
C321 GF_NI_IN_C_BASE_0.pdrive_y_<1> GF_NI_IN_C_BASE_0.ndrive_Y_<1> 0.463637f
C322 GF_NI_IN_C_BASE_0.comp018green_out_predrv_3.nmos_6p0_CDNS_4066195314519_0.D GF_NI_IN_C_BASE_0.ndrive_Y_<1> 1.27145f
C323 GF_NI_IN_C_BASE_0.comp018green_out_predrv_0.SL GF_NI_IN_C_BASE_0.comp018green_out_predrv_0.SLB 9.573371f
C324 GF_NI_IN_C_BASE_0.comp018green_out_predrv_0.A GF_NI_IN_C_BASE_0.comp018green_out_predrv_0.nmos_6p0_CDNS_4066195314519_2.S 1.67734f
C325 GF_NI_IN_C_BASE_0.comp018green_out_predrv_0.A GF_NI_IN_C_BASE_0.comp018green_out_predrv_1.nmos_6p0_CDNS_4066195314519_2.S 1.67734f
C326 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.EN DVDD 1.75575f
C327 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_cms_smt_0.nmos_6p0_CDNS_4066195314535_0.D GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_drv_0.A 3.40047f
C328 GF_NI_IN_C_BASE_0.ndrive_Y_<1> PAD 7.99617f
C329 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_drv_0.nmos_6p0_CDNS_4066195314547_0.S PD 0.223029f
C330 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_pupd_0.ppolyf_u_CDNS_4066195314533_5.MINUS GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_pupd_0.ppolyf_u_CDNS_4066195314533_0.PLUS 4.22e-19
C331 DVDD VDD 48.8373f
C332 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_1.EN DVDD 2.35753f
C333 GF_NI_IN_C_BASE_0.comp018green_out_predrv_0.A DVSS 11.039001f
C334 GF_NI_IN_C_BASE_0.ndrive_y_<0> GF_NI_IN_C_BASE_0.pdrive_x_<0> 7.63e-19
C335 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_logic_pupd_0.comp018green_std_xor2_0.nmos_6p0_CDNS_4066195314530_2.D DVSS 0.369885f
C336 GF_NI_IN_C_BASE_0.comp018green_out_predrv_1.ENB DVDD 1.3057f
C337 GF_NI_IN_C_BASE_0.pdrive_x_<3> GF_NI_IN_C_BASE_0.ndrive_x_<3> 7.34e-19
C338 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.ENB GF_NI_IN_C_BASE_0.comp018green_out_predrv_0.nmos_6p0_CDNS_4066195314519_0.D 2.42579f
C339 GF_NI_IN_C_BASE_0.ndrive_Y_<1> DVSS 10.7603f
C340 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.ENB 0.047579f
C341 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_drv_0.A GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_pupd_0.ppolyf_u_CDNS_4066195314533_5.MINUS 0.001033f
C342 GF_NI_IN_C_BASE_0.ndrive_x_<0> GF_NI_IN_C_BASE_0.ndrive_y_<0> 10.427401f
C343 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.nmos_6p0_CDNS_4066195314511_1.S GF_NI_IN_C_BASE_0.comp018green_out_predrv_0.SL 4.94e-20
C344 GF_NI_IN_C_BASE_0.comp018green_out_predrv_1.EN VDD 0.402841f
C345 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_1.EN GF_NI_IN_C_BASE_0.comp018green_out_predrv_1.EN 0.712898f
C346 GF_NI_IN_C_BASE_0.comp018green_out_predrv_1.ENB GF_NI_IN_C_BASE_0.comp018green_out_predrv_1.nmos_6p0_CDNS_4066195314519_0.D 2.42388f
C347 GF_NI_IN_C_BASE_0.comp018green_out_predrv_0.A GF_NI_IN_C_BASE_0.comp018green_out_predrv_3.nmos_6p0_CDNS_4066195314519_2.S 1.67859f
C348 GF_NI_IN_C_BASE_0.ndrive_y_<2> GF_NI_IN_C_BASE_0.ndrive_Y_<3> 0.003823f
C349 GF_NI_IN_C_BASE_0.ndrive_x_<2> GF_NI_IN_C_BASE_0.ndrive_x_<3> 0.003209f
C350 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_a_0.nmos_6p0_CDNS_4066195314511_3.S VDD 0.28821f
C351 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_1.EN GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_a_0.nmos_6p0_CDNS_4066195314511_3.S 4.38e-19
C352 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_1.EN GF_NI_IN_C_BASE_0.comp018green_out_predrv_2.nmos_6p0_CDNS_4066195314519_2.S 2.30393f
C353 GF_NI_IN_C_BASE_0.comp018green_out_predrv_1.EN GF_NI_IN_C_BASE_0.comp018green_out_predrv_1.ENB 5.39405f
C354 GF_NI_IN_C_BASE_0.comp018green_out_predrv_0.SL GF_NI_IN_C_BASE_0.pdrive_y_<2> 1.53e-19
C355 GF_NI_IN_C_BASE_0.comp018green_out_predrv_1.ENB GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_a_0.nmos_6p0_CDNS_4066195314511_3.S 0.001643f
C356 GF_NI_IN_C_BASE_0.comp018green_out_predrv_3.nmos_6p0_CDNS_4066195314519_2.S GF_NI_IN_C_BASE_0.ndrive_Y_<1> 1.90029f
C357 GF_NI_IN_C_BASE_0.comp018green_out_predrv_0.nmos_6p0_CDNS_4066195314519_0.D GF_NI_IN_C_BASE_0.ndrive_x_<1> 0.00245f
C358 GF_NI_IN_C_BASE_0.comp018green_out_predrv_1.ENB GF_NI_IN_C_BASE_0.comp018green_out_predrv_2.nmos_6p0_CDNS_4066195314519_2.S 1.28e-19
C359 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_pupd_0.ppolyf_u_CDNS_4066195314533_1.PLUS DVSS 0.073601f
C360 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_1.nmos_6p0_CDNS_4066195314511_1.S DVDD 0.487748f
C361 GF_NI_IN_C_BASE_0.comp018green_out_predrv_0.A GF_NI_IN_C_BASE_0.ndrive_y_<2> 0.001225f
C362 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_1.EN GF_NI_IN_C_BASE_0.pdrive_y_<1> 0.005045f
C363 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_1.EN GF_NI_IN_C_BASE_0.comp018green_out_predrv_3.nmos_6p0_CDNS_4066195314519_0.D 2.2174f
C364 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.ENB GF_NI_IN_C_BASE_0.pdrive_x_<0> 6.39e-19
C365 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_3.Z GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_cms_smt_0.nmos_6p0_CDNS_4066195314535_0.D 1.98091f
C366 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_pupd_0.ppolyf_u_CDNS_4066195314533_0.PLUS DVDD 0.353843f
C367 PAD VDD 1.40846f
C368 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_1.EN PAD 0.109854f
C369 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_logic_pupd_0.comp018green_std_xor2_0.nmos_6p0_CDNS_4066195314530_2.D PU 0.840559f
C370 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.EN GF_NI_IN_C_BASE_0.comp018green_out_predrv_0.nmos_6p0_CDNS_4066195314519_2.S 2.30471f
C371 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.ENB GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_1.ENB 0.042012f
C372 GF_NI_IN_C_BASE_0.comp018green_out_predrv_1.ENB PAD 0.005919f
C373 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.ENB GF_NI_IN_C_BASE_0.ndrive_x_<0> 0.00719f
C374 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_cms_smt_0.nmos_6p0_CDNS_4066195314530_0.D VDD 0.083541f
C375 GF_NI_IN_C_BASE_0.comp018green_out_predrv_0.SL GF_NI_IN_C_BASE_0.pdrive_y_<0> 1.53e-19
C376 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.EN DVSS 2.27601f
C377 GF_NI_IN_C_BASE_0.comp018green_out_predrv_0.SLB GF_NI_IN_C_BASE_0.pdrive_y_<2> 0.737025f
C378 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_3.Z GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_pupd_0.ppolyf_u_CDNS_4066195314533_5.MINUS 0.002397f
C379 DVSS VDD 31.514502f
C380 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_1.EN DVSS 3.81168f
C381 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_drv_0.A DVDD 2.37178f
C382 GF_NI_IN_C_BASE_0.pdrive_x_<1> GF_NI_IN_C_BASE_0.ndrive_x_<1> 0.156934f
C383 GF_NI_IN_C_BASE_0.pdrive_x_<0> GF_NI_IN_C_BASE_0.ndrive_x_<1> 0.074382f
C384 GF_NI_IN_C_BASE_0.comp018green_out_predrv_1.ENB GF_NI_IN_C_BASE_0.comp018green_out_predrv_1.nmos_6p0_CDNS_4066195314519_2.S 0.561221f
C385 GF_NI_IN_C_BASE_0.comp018green_out_predrv_0.A GF_NI_IN_C_BASE_0.ndrive_y_<0> 0.001918f
C386 GF_NI_IN_C_BASE_0.comp018green_out_predrv_2.nmos_6p0_CDNS_4066195314519_0.D GF_NI_IN_C_BASE_0.pdrive_x_<3> 5.58e-20
C387 GF_NI_IN_C_BASE_0.comp018green_out_predrv_2.nmos_6p0_CDNS_4066195314519_0.D GF_NI_IN_C_BASE_0.pdrive_x_<2> 0.86434f
C388 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_logic_pupd_0.comp018green_std_xor2_0.nmos_6p0_CDNS_4066195314530_2.D PD 0.100418f
C389 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_pupd_0.ppolyf_u_CDNS_4066195314533_5.MINUS GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_pupd_0.ppolyf_u_CDNS_4066195314533_3.MINUS 0.035159f
C390 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_1.Z VDD 0.182038f
C391 GF_NI_IN_C_BASE_0.comp018green_out_predrv_1.ENB DVSS 2.5731f
C392 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_1.ENB GF_NI_IN_C_BASE_0.ndrive_x_<1> 0.012707f
C393 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_cms_smt_0.nmos_6p0_CDNS_4066195314540_0.S GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_drv_0.A 0.894376f
C394 GF_NI_IN_C_BASE_0.ndrive_y_<0> GF_NI_IN_C_BASE_0.ndrive_Y_<1> 0.031279f
C395 GF_NI_IN_C_BASE_0.ndrive_x_<0> GF_NI_IN_C_BASE_0.ndrive_x_<1> 0.003886f
C396 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_pupd_0.PU_B 1.71e-19
C397 GF_NI_IN_C_BASE_0.comp018green_out_predrv_2.nmos_6p0_CDNS_4066195314519_0.D GF_NI_IN_C_BASE_0.ndrive_x_<2> 0.035148f
C398 GF_NI_IN_C_BASE_0.ndrive_Y_<3> GF_NI_IN_C_BASE_0.ndrive_x_<3> 10.302f
C399 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_1.EN GF_NI_IN_C_BASE_0.comp018green_out_predrv_3.nmos_6p0_CDNS_4066195314519_2.S 2.30509f
C400 GF_NI_IN_C_BASE_0.comp018green_out_predrv_3.nmos_6p0_CDNS_4066195314519_2.S VDD 0.002554f
C401 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_pupd_0.PD GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_pupd_0.PU_B 2.46651f
C402 GF_NI_IN_C_BASE_0.comp018green_out_predrv_0.SLB GF_NI_IN_C_BASE_0.pdrive_y_<0> 0.737025f
C403 GF_NI_IN_C_BASE_0.comp018green_out_predrv_0.SL DVDD 7.04964f
C404 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_a_0.nmos_6p0_CDNS_4066195314511_1.D DVDD 0.48747f
C405 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE GF_NI_IN_C_BASE_0.comp018green_out_predrv_0.nmos_6p0_CDNS_4066195314519_0.D 9.09e-19
C406 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_cms_smt_0.nmos_6p0_CDNS_4066195314537_0.D GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_drv_0.A 0.007263f
C407 GF_NI_IN_C_BASE_0.pdrive_x_<2> GF_NI_IN_C_BASE_0.pdrive_x_<3> 0.048189f
C408 GF_NI_IN_C_BASE_0.comp018green_out_predrv_0.A GF_NI_IN_C_BASE_0.ndrive_x_<3> 0.001965f
C409 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_1.EN GF_NI_IN_C_BASE_0.ndrive_y_<2> 6.12e-19
C410 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_pupd_0.PU_B GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_drv_0.nmos_6p0_CDNS_4066195314547_0.S 0.060445f
C411 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_1.nmos_6p0_CDNS_4066195314511_1.S DVSS 0.624553f
C412 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.ENB GF_NI_IN_C_BASE_0.comp018green_out_predrv_0.A 0.658049f
C413 VDD PU 3.47633f
C414 GF_NI_IN_C_BASE_0.comp018green_out_predrv_0.SL GF_NI_IN_C_BASE_0.pdrive_y_<3> 1.53e-19
C415 GF_NI_IN_C_BASE_0.comp018green_out_predrv_0.SL GF_NI_IN_C_BASE_0.comp018green_out_predrv_1.nmos_6p0_CDNS_4066195314519_0.D 0.01198f
C416 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_cms_smt_0.nmos_6p0_CDNS_4066195314535_0.D GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_pupd_0.ppolyf_u_CDNS_4066195314533_5.MINUS 0.001011f
C417 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_1.ENB GF_NI_IN_C_BASE_0.comp018green_out_predrv_2.nmos_6p0_CDNS_4066195314519_0.D 2.42536f
C418 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_3.Z DVDD 3.12747f
C419 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_pupd_0.ppolyf_u_CDNS_4066195314533_0.PLUS DVSS 0.069602f
C420 GF_NI_IN_C_BASE_0.comp018green_out_predrv_1.ENB GF_NI_IN_C_BASE_0.ndrive_y_<2> 7.22e-19
C421 GF_NI_IN_C_BASE_0.ndrive_x_<2> GF_NI_IN_C_BASE_0.pdrive_x_<3> 0.981343f
C422 w_4468_53312# GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE 0.161159f
C423 GF_NI_IN_C_BASE_0.ndrive_x_<2> GF_NI_IN_C_BASE_0.pdrive_x_<2> 0.523505f
C424 GF_NI_IN_C_BASE_0.comp018green_out_predrv_1.EN GF_NI_IN_C_BASE_0.comp018green_out_predrv_0.SL 0.09891f
C425 GF_NI_IN_C_BASE_0.comp018green_out_predrv_1.EN GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_a_0.nmos_6p0_CDNS_4066195314511_1.D 0.001593f
C426 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.ENB GF_NI_IN_C_BASE_0.ndrive_Y_<1> 3.42e-19
C427 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_pupd_0.ppolyf_u_CDNS_4066195314533_3.MINUS DVDD 0.352299f
C428 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_a_0.nmos_6p0_CDNS_4066195314511_3.S GF_NI_IN_C_BASE_0.comp018green_out_predrv_0.SL 4.94e-20
C429 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_a_0.nmos_6p0_CDNS_4066195314511_3.S GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_a_0.nmos_6p0_CDNS_4066195314511_1.D 0.589096f
C430 GF_NI_IN_C_BASE_0.comp018green_out_predrv_0.SL GF_NI_IN_C_BASE_0.comp018green_out_predrv_2.nmos_6p0_CDNS_4066195314519_2.S 0.324691f
C431 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_cms_smt_0.nmos_6p0_CDNS_4066195314530_0.D GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_drv_0.A 0.504632f
C432 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_3.Z GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_cms_smt_0.nmos_6p0_CDNS_4066195314540_0.S 0.050642f
C433 GF_NI_IN_C_BASE_0.comp018green_out_predrv_0.SLB DVDD 0.478425f
C434 GF_NI_IN_C_BASE_0.comp018green_out_predrv_0.nmos_6p0_CDNS_4066195314519_0.D GF_NI_IN_C_BASE_0.pdrive_x_<1> 5.58e-20
C435 GF_NI_IN_C_BASE_0.comp018green_out_predrv_0.nmos_6p0_CDNS_4066195314519_0.D GF_NI_IN_C_BASE_0.pdrive_x_<0> 0.718068f
C436 GF_NI_IN_C_BASE_0.pdrive_x_<1> GF_NI_IN_C_BASE_0.pdrive_x_<2> 0.925558f
C437 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.EN GF_NI_IN_C_BASE_0.ndrive_y_<0> 0.00714f
C438 VDD PD 4.66804f
C439 GF_NI_IN_C_BASE_0.comp018green_out_predrv_0.A GF_NI_IN_C_BASE_0.ndrive_x_<1> 0.00192f
C440 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_drv_0.A DVSS 1.44026f
C441 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_pupd_0.PD GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_drv_0.nmos_6p0_CDNS_4066195314547_0.S 0.08422f
C442 GF_NI_IN_C_BASE_0.comp018green_out_predrv_0.SL GF_NI_IN_C_BASE_0.pdrive_y_<1> 1.53e-19
C443 GF_NI_IN_C_BASE_0.comp018green_out_predrv_0.SL GF_NI_IN_C_BASE_0.comp018green_out_predrv_3.nmos_6p0_CDNS_4066195314519_0.D 0.01198f
C444 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_1.Z GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_drv_0.A 0.290394f
C445 GF_NI_IN_C_BASE_0.comp018green_out_predrv_0.SLB GF_NI_IN_C_BASE_0.comp018green_out_predrv_1.nmos_6p0_CDNS_4066195314519_0.D 0.026278f
C446 GF_NI_IN_C_BASE_0.comp018green_out_predrv_0.SLB GF_NI_IN_C_BASE_0.pdrive_y_<3> 0.737025f
C447 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_1.ENB 0.037834f
C448 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_1.ENB GF_NI_IN_C_BASE_0.pdrive_x_<2> 0.035199f
C449 GF_NI_IN_C_BASE_0.comp018green_out_predrv_0.nmos_6p0_CDNS_4066195314519_0.D GF_NI_IN_C_BASE_0.ndrive_x_<0> 0.033783f
C450 GF_NI_IN_C_BASE_0.comp018green_out_predrv_0.SL PAD 0.598535f
C451 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_a_0.nmos_6p0_CDNS_4066195314511_1.D PAD 0.003241f
C452 GF_NI_IN_C_BASE_0.ndrive_Y_<1> GF_NI_IN_C_BASE_0.ndrive_x_<1> 14.8135f
C453 GF_NI_IN_C_BASE_0.comp018green_out_predrv_1.EN GF_NI_IN_C_BASE_0.comp018green_out_predrv_0.SLB 0.039646f
C454 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_3.Z GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_cms_smt_0.nmos_6p0_CDNS_4066195314537_0.D 0.079431f
C455 GF_NI_IN_C_BASE_0.comp018green_out_predrv_0.SL GF_NI_IN_C_BASE_0.comp018green_out_predrv_0.nmos_6p0_CDNS_4066195314519_2.S 0.328757f
C456 GF_NI_IN_C_BASE_0.comp018green_out_predrv_0.SL GF_NI_IN_C_BASE_0.comp018green_out_predrv_1.nmos_6p0_CDNS_4066195314519_2.S 0.329817f
C457 GF_NI_IN_C_BASE_0.comp018green_out_predrv_0.SLB GF_NI_IN_C_BASE_0.comp018green_out_predrv_2.nmos_6p0_CDNS_4066195314519_2.S 0.003533f
C458 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_1.ENB GF_NI_IN_C_BASE_0.ndrive_x_<2> 0.007532f
C459 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.nmos_6p0_CDNS_4066195314511_1.S DVDD 0.488555f
C460 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_cms_smt_0.nmos_6p0_CDNS_4066195314535_0.D DVDD 1.95425f
C461 GF_NI_IN_C_BASE_0.pdrive_x_<0> GF_NI_IN_C_BASE_0.pdrive_x_<1> 0.048189f
C462 GF_NI_IN_C_BASE_0.comp018green_out_predrv_0.SL DVSS 9.61187f
C463 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_a_0.nmos_6p0_CDNS_4066195314511_1.D DVSS 0.627513f
C464 GF_NI_IN_C_BASE_0.comp018green_out_predrv_0.A GF_NI_IN_C_BASE_0.comp018green_out_predrv_2.nmos_6p0_CDNS_4066195314519_0.D 0.505117f
C465 GF_NI_IN_C_BASE_0.pdrive_y_<2> DVDD 16.792099f
C466 DVDD Y 2.10224f
C467 GF_NI_IN_C_BASE_0.comp018green_out_predrv_0.SLB GF_NI_IN_C_BASE_0.pdrive_y_<1> 0.737025f
C468 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.EN GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.ENB 1.47047f
C469 GF_NI_IN_C_BASE_0.comp018green_out_predrv_0.SLB GF_NI_IN_C_BASE_0.comp018green_out_predrv_3.nmos_6p0_CDNS_4066195314519_0.D 0.026278f
C470 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_1.ENB GF_NI_IN_C_BASE_0.pdrive_x_<1> 0.035214f
C471 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_1.ENB GF_NI_IN_C_BASE_0.pdrive_x_<0> 0.003333f
C472 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_3.Z GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_cms_smt_0.nmos_6p0_CDNS_4066195314530_0.D 0.303391f
C473 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.ENB VDD 0.13593f
C474 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.ENB GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_1.EN 0.001515f
C475 GF_NI_IN_C_BASE_0.ndrive_x_<0> GF_NI_IN_C_BASE_0.pdrive_x_<0> 4.33e-19
C476 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_drv_0.A PU 0.001361f
C477 GF_NI_IN_C_BASE_0.comp018green_out_predrv_0.SLB PAD 0.10231f
C478 GF_NI_IN_C_BASE_0.comp018green_out_predrv_1.ENB GF_NI_IN_C_BASE_0.ndrive_x_<3> 0.01433f
C479 GF_NI_IN_C_BASE_0.pdrive_x_<3> GF_NI_IN_C_BASE_0.ndrive_Y_<3> 4.4e-19
C480 GF_NI_IN_C_BASE_0.pdrive_y_<2> GF_NI_IN_C_BASE_0.pdrive_y_<3> 0.124712f
C481 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_pupd_0.ppolyf_u_CDNS_4066195314533_5.MINUS DVDD 5.16836f
C482 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_3.Z DVSS 4.87161f
C483 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_pupd_0.PU_B GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_logic_pupd_0.comp018green_std_xor2_0.nmos_6p0_CDNS_4066195314530_2.D 3.11e-20
C484 GF_NI_IN_C_BASE_0.comp018green_out_predrv_0.SL GF_NI_IN_C_BASE_0.comp018green_out_predrv_3.nmos_6p0_CDNS_4066195314519_2.S 0.329551f
C485 GF_NI_IN_C_BASE_0.comp018green_out_predrv_0.SLB GF_NI_IN_C_BASE_0.comp018green_out_predrv_1.nmos_6p0_CDNS_4066195314519_2.S 0.014194f
C486 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_1.Z GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_3.Z 1.53428f
C487 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_pupd_0.ppolyf_u_CDNS_4066195314533_3.MINUS DVSS 0.053116f
C488 GF_NI_IN_C_BASE_0.ndrive_x_<2> GF_NI_IN_C_BASE_0.ndrive_Y_<3> 0.003293f
C489 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.EN GF_NI_IN_C_BASE_0.ndrive_x_<1> 6.12e-19
C490 GF_NI_IN_C_BASE_0.comp018green_out_predrv_0.SLB DVSS 17.344698f
C491 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_cms_smt_0.nmos_6p0_CDNS_4066195314535_0.D GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_cms_smt_0.nmos_6p0_CDNS_4066195314537_0.D 1.21e-19
C492 GF_NI_IN_C_BASE_0.comp018green_out_predrv_0.A GF_NI_IN_C_BASE_0.comp018green_out_predrv_0.nmos_6p0_CDNS_4066195314519_0.D 0.505117f
C493 GF_NI_IN_C_BASE_0.comp018green_out_predrv_2.nmos_6p0_CDNS_4066195314519_2.S GF_NI_IN_C_BASE_0.pdrive_y_<2> 0.026792f
C494 GF_NI_IN_C_BASE_0.pdrive_y_<0> DVDD 18.050402f
C495 GF_NI_IN_C_BASE_0.comp018green_out_predrv_0.A GF_NI_IN_C_BASE_0.pdrive_x_<3> 0.00224f
C496 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE GF_NI_IN_C_BASE_0.comp018green_out_predrv_0.A 0.011497f
C497 GF_NI_IN_C_BASE_0.comp018green_out_predrv_0.A GF_NI_IN_C_BASE_0.pdrive_x_<2> 0.051146f
C498 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_drv_0.A PD 0.055616f
C499 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_1.EN GF_NI_IN_C_BASE_0.ndrive_x_<1> 0.003589f
C500 GF_NI_IN_C_BASE_0.comp018green_out_predrv_0.SL GF_NI_IN_C_BASE_0.ndrive_y_<2> 1.11498f
C501 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_logic_pupd_0.comp018green_std_xor2_0.nmos_6p0_CDNS_4066195314530_2.D 0.397451f
C502 GF_NI_IN_C_BASE_0.comp018green_out_predrv_0.nmos_6p0_CDNS_4066195314519_0.D GF_NI_IN_C_BASE_0.ndrive_Y_<1> 0.001369f
C503 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_pupd_0.PD GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_logic_pupd_0.comp018green_std_xor2_0.nmos_6p0_CDNS_4066195314530_2.D 3.68e-20
C504 GF_NI_IN_C_BASE_0.comp018green_out_predrv_0.A GF_NI_IN_C_BASE_0.ndrive_x_<2> 0.00138f
C505 GF_NI_IN_C_BASE_0.pdrive_y_<2> PAD 10.1896f
C506 GF_NI_IN_C_BASE_0.comp018green_out_predrv_0.SLB GF_NI_IN_C_BASE_0.comp018green_out_predrv_3.nmos_6p0_CDNS_4066195314519_2.S 0.003533f
C507 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_cms_smt_0.nmos_6p0_CDNS_4066195314535_0.D GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_cms_smt_0.nmos_6p0_CDNS_4066195314530_0.D 0.217321f
C508 GF_NI_IN_C_BASE_0.ndrive_Y_<1> GF_NI_IN_C_BASE_0.ndrive_x_<2> 0.13555f
C509 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.nmos_6p0_CDNS_4066195314511_1.S DVSS 0.624553f
C510 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_3.Z PU 2.62886f
C511 GF_NI_IN_C_BASE_0.comp018green_out_predrv_0.A GF_NI_IN_C_BASE_0.pdrive_x_<1> 0.051146f
C512 GF_NI_IN_C_BASE_0.comp018green_out_predrv_0.A GF_NI_IN_C_BASE_0.pdrive_x_<0> 0.002263f
C513 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_cms_smt_0.nmos_6p0_CDNS_4066195314535_0.D DVSS 0.663933f
C514 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_1.EN GF_NI_IN_C_BASE_0.comp018green_out_predrv_2.nmos_6p0_CDNS_4066195314519_0.D 2.21763f
C515 GF_NI_IN_C_BASE_0.comp018green_out_predrv_0.SL GF_NI_IN_C_BASE_0.ndrive_y_<0> 1.12772f
C516 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_1.Z GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_cms_smt_0.nmos_6p0_CDNS_4066195314535_0.D 0.66544f
C517 GF_NI_IN_C_BASE_0.pdrive_y_<2> DVSS 2.51221f
C518 DVSS Y 0.982246f
C519 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_pupd_0.ppolyf_u_CDNS_4066195314533_1.PLUS 9.81e-19
C520 GF_NI_IN_C_BASE_0.pdrive_x_<1> GF_NI_IN_C_BASE_0.ndrive_Y_<1> 0.668765f
C521 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_1.ENB GF_NI_IN_C_BASE_0.comp018green_out_predrv_0.A 4.43546f
C522 GF_NI_IN_C_BASE_0.pdrive_y_<0> GF_NI_IN_C_BASE_0.pdrive_y_<1> 0.124934f
C523 GF_NI_IN_C_BASE_0.pdrive_x_<0> GF_NI_IN_C_BASE_0.ndrive_Y_<1> 0.981139f
C524 GF_NI_IN_C_BASE_0.pdrive_y_<0> GF_NI_IN_C_BASE_0.comp018green_out_predrv_3.nmos_6p0_CDNS_4066195314519_0.D 0.02501f
C525 GF_NI_IN_C_BASE_0.comp018green_out_predrv_1.ENB GF_NI_IN_C_BASE_0.comp018green_out_predrv_2.nmos_6p0_CDNS_4066195314519_0.D 1.8e-19
C526 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_cms_smt_0.nmos_6p0_CDNS_4066195314530_0.D GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_pupd_0.ppolyf_u_CDNS_4066195314533_5.MINUS 5.42e-20
C527 GF_NI_IN_C_BASE_0.comp018green_out_predrv_0.A GF_NI_IN_C_BASE_0.ndrive_x_<0> 7.02e-19
C528 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_cms_smt_0.nmos_6p0_CDNS_4066195314540_0.S DVDD 0.355101f
C529 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_pupd_0.PU_B VDD 0.516636f
C530 GF_NI_IN_C_BASE_0.pdrive_y_<3> DVDD 17.9215f
C531 GF_NI_IN_C_BASE_0.comp018green_out_predrv_1.nmos_6p0_CDNS_4066195314519_0.D DVDD 4.00784f
C532 GF_NI_IN_C_BASE_0.pdrive_y_<0> PAD 10.1953f
C533 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_3.Z PD 2.63281f
C534 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_pupd_0.ppolyf_u_CDNS_4066195314533_5.MINUS DVSS 1.09337f
C535 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_1.ENB GF_NI_IN_C_BASE_0.ndrive_Y_<1> 0.360786f
C536 GF_NI_IN_C_BASE_0.ndrive_x_<0> GF_NI_IN_C_BASE_0.ndrive_Y_<1> 0.002206f
C537 GF_NI_IN_C_BASE_0.comp018green_out_predrv_1.EN DVDD 1.74689f
C538 GF_NI_IN_C_BASE_0.comp018green_out_predrv_0.nmos_6p0_CDNS_4066195314519_2.S GF_NI_IN_C_BASE_0.pdrive_y_<0> 0.020536f
C539 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_1.Z GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_pupd_0.ppolyf_u_CDNS_4066195314533_5.MINUS 0.002385f
C540 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.EN GF_NI_IN_C_BASE_0.comp018green_out_predrv_0.nmos_6p0_CDNS_4066195314519_0.D 2.21936f
C541 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_a_0.nmos_6p0_CDNS_4066195314511_3.S DVDD 1.05814f
C542 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.EN 0.218225f
C543 GF_NI_IN_C_BASE_0.comp018green_out_predrv_2.nmos_6p0_CDNS_4066195314519_2.S DVDD 5.24568f
C544 GF_NI_IN_C_BASE_0.comp018green_out_predrv_1.nmos_6p0_CDNS_4066195314519_0.D GF_NI_IN_C_BASE_0.pdrive_y_<3> 2.92427f
C545 Y VSS 4.754909f
C546 PD VSS 14.931949f
C547 PU VSS 11.908794f
C548 VDD VSS 0.158878p
C549 DVSS VSS 0.200993p
C550 PAD VSS 96.433205f
C551 DVDD VSS 1.073183p
C552 GF_NI_IN_C_BASE_0.ndrive_x_<3> VSS 26.701586f
C553 GF_NI_IN_C_BASE_0.ndrive_Y_<3> VSS 22.96035f
C554 GF_NI_IN_C_BASE_0.pdrive_y_<3> VSS 21.603668f
C555 GF_NI_IN_C_BASE_0.pdrive_x_<3> VSS 5.376266f
C556 GF_NI_IN_C_BASE_0.comp018green_out_predrv_1.nmos_6p0_CDNS_4066195314519_2.S VSS 1.790432f
C557 GF_NI_IN_C_BASE_0.comp018green_out_predrv_1.nmos_6p0_CDNS_4066195314519_0.D VSS 1.300081f
C558 GF_NI_IN_C_BASE_0.pdrive_x_<2> VSS 7.15483f
C559 GF_NI_IN_C_BASE_0.pdrive_y_<2> VSS 20.644226f
C560 GF_NI_IN_C_BASE_0.ndrive_y_<2> VSS 28.465302f
C561 GF_NI_IN_C_BASE_0.ndrive_x_<2> VSS 32.978447f
C562 GF_NI_IN_C_BASE_0.comp018green_out_predrv_2.nmos_6p0_CDNS_4066195314519_0.D VSS 1.297007f
C563 GF_NI_IN_C_BASE_0.comp018green_out_predrv_2.nmos_6p0_CDNS_4066195314519_2.S VSS 1.730357f
C564 GF_NI_IN_C_BASE_0.ndrive_x_<1> VSS 32.483826f
C565 GF_NI_IN_C_BASE_0.ndrive_Y_<1> VSS 31.33064f
C566 GF_NI_IN_C_BASE_0.pdrive_y_<1> VSS 21.372349f
C567 GF_NI_IN_C_BASE_0.pdrive_x_<1> VSS 7.13999f
C568 GF_NI_IN_C_BASE_0.comp018green_out_predrv_3.nmos_6p0_CDNS_4066195314519_2.S VSS 1.724805f
C569 GF_NI_IN_C_BASE_0.comp018green_out_predrv_3.nmos_6p0_CDNS_4066195314519_0.D VSS 1.297141f
C570 GF_NI_IN_C_BASE_0.pdrive_x_<0> VSS 5.363458f
C571 GF_NI_IN_C_BASE_0.pdrive_y_<0> VSS 21.647776f
C572 GF_NI_IN_C_BASE_0.ndrive_y_<0> VSS 25.177105f
C573 GF_NI_IN_C_BASE_0.ndrive_x_<0> VSS 25.017963f
C574 GF_NI_IN_C_BASE_0.comp018green_out_predrv_0.nmos_6p0_CDNS_4066195314519_0.D VSS 1.300759f
C575 GF_NI_IN_C_BASE_0.comp018green_out_predrv_0.nmos_6p0_CDNS_4066195314519_2.S VSS 1.793422f
C576 GF_NI_IN_C_BASE_0.comp018green_out_predrv_0.SLB VSS 6.851561f
C577 GF_NI_IN_C_BASE_0.comp018green_out_predrv_0.SL VSS 11.020435f
C578 GF_NI_IN_C_BASE_0.comp018green_out_predrv_0.A VSS 15.25784f
C579 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_a_0.nmos_6p0_CDNS_4066195314511_1.D VSS 1.038f
C580 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_a_0.nmos_6p0_CDNS_4066195314511_3.S VSS 0.331655f
C581 GF_NI_IN_C_BASE_0.comp018green_out_predrv_1.ENB VSS 9.62785f
C582 GF_NI_IN_C_BASE_0.comp018green_out_predrv_1.EN VSS 10.112769f
C583 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_1.ENB VSS 10.52142f
C584 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_1.nmos_6p0_CDNS_4066195314511_1.S VSS 0.982221f
C585 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_1.EN VSS 12.747739f
C586 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.ENB VSS 4.6969f
C587 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.EN VSS 5.6328f
C588 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.nmos_6p0_CDNS_4066195314511_1.S VSS 1.01104f
C589 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_logic_pupd_0.comp018green_std_xor2_0.nmos_6p0_CDNS_4066195314530_2.D VSS 0.810347f
C590 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_pupd_0.ppolyf_u_CDNS_4066195314533_1.PLUS VSS 0.15084f
C591 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_pupd_0.ppolyf_u_CDNS_4066195314533_0.PLUS VSS 0.148863f
C592 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_pupd_0.ppolyf_u_CDNS_4066195314533_3.MINUS VSS 0.148863f
C593 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_pupd_0.ppolyf_u_CDNS_4066195314533_5.MINUS VSS 6.718775f
C594 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_drv_0.nmos_6p0_CDNS_4066195314547_0.S VSS 4.00792f
C595 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_drv_0.A VSS 3.577513f
C596 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_cms_smt_0.nmos_6p0_CDNS_4066195314540_0.S VSS 2.347956f
C597 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_cms_smt_0.nmos_6p0_CDNS_4066195314537_0.D VSS 0.632754f
C598 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_cms_smt_0.nmos_6p0_CDNS_4066195314530_0.D VSS 4.30132f
C599 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_cms_smt_0.nmos_6p0_CDNS_4066195314535_0.D VSS 1.270011f
C600 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_pupd_0.PU_B VSS 7.37483f
C601 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_pupd_0.PD VSS 4.77241f
C602 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_3.Z VSS 10.80828f
C603 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_1.Z VSS 4.827301f
C604 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE VSS 57.476803f
C605 w_4468_53312# VSS 39.222f
C606 PD.t6 VSS 0.328461f
C607 PD.n0 VSS 0.160976f
C608 PD.n1 VSS 1.4255f
C609 PD.t5 VSS 0.299567f
C610 PD.t1 VSS 0.597f
C611 PD.n2 VSS 1.00116f
C612 PD.t0 VSS 0.608834f
C613 PD.n3 VSS 0.451354f
C614 PD.t2 VSS 0.697402f
C615 PD.n4 VSS 0.940613f
C616 PD.t4 VSS 0.674453f
C617 PD.t3 VSS 0.6813f
C618 PD.n5 VSS 0.771456f
C619 PD.n6 VSS 0.284198f
C620 PD.n7 VSS 6.72437f
C621 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_1.ENB.t5 VSS 1.00379f
C622 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_1.ENB.t3 VSS 2.03153f
C623 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_1.ENB.t0 VSS 0.291265f
C624 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_1.ENB.t1 VSS 1.00909f
C625 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_1.ENB.n0 VSS 3.98221f
C626 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_1.ENB.t2 VSS 1.00379f
C627 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_1.ENB.t4 VSS 2.03153f
C628 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.EN.t4 VSS 0.536852f
C629 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.EN.t3 VSS 0.287306f
C630 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.EN.n0 VSS 0.382086f
C631 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.EN.t0 VSS 0.206579f
C632 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.EN.t2 VSS 0.528517f
C633 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.EN.t5 VSS 1.06955f
C634 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.EN.t1 VSS 0.505447f
C635 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_pupd_0.ppolyf_u_CDNS_4066195314533_5.MINUS.t0 VSS 0.210383f
C636 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_pupd_0.ppolyf_u_CDNS_4066195314533_5.MINUS.n0 VSS 0.232277f
C637 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_pupd_0.ppolyf_u_CDNS_4066195314533_5.MINUS.n1 VSS 0.046696f
C638 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_pupd_0.ppolyf_u_CDNS_4066195314533_5.MINUS.t1 VSS 0.019531f
C639 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_pupd_0.ppolyf_u_CDNS_4066195314533_5.MINUS.n2 VSS 1.35751f
C640 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_pupd_0.ppolyf_u_CDNS_4066195314533_5.MINUS.t2 VSS 0.033306f
C641 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_cms_smt_0.nmos_6p0_CDNS_4066195314535_0.D.t0 VSS 0.159919f
C642 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_cms_smt_0.nmos_6p0_CDNS_4066195314535_0.D.t1 VSS 0.463729f
C643 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_cms_smt_0.nmos_6p0_CDNS_4066195314535_0.D.n0 VSS 1.04783f
C644 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_cms_smt_0.nmos_6p0_CDNS_4066195314535_0.D.t2 VSS 0.198371f
C645 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_cms_smt_0.nmos_6p0_CDNS_4066195314535_0.D.t4 VSS 0.195341f
C646 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_cms_smt_0.nmos_6p0_CDNS_4066195314535_0.D.n1 VSS 0.973754f
C647 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_cms_smt_0.nmos_6p0_CDNS_4066195314535_0.D.t3 VSS 0.157997f
C648 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.ENB.t1 VSS 0.138169f
C649 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.ENB.t0 VSS 0.478686f
C650 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.ENB.t3 VSS 0.476171f
C651 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.ENB.t2 VSS 0.963705f
C652 GF_NI_IN_C_BASE_0.pdrive_y_<3>.t0 VSS 1.26189f
C653 GF_NI_IN_C_BASE_0.pdrive_y_<3>.t2 VSS 1.25662f
C654 GF_NI_IN_C_BASE_0.pdrive_y_<3>.t3 VSS 1.61254f
C655 GF_NI_IN_C_BASE_0.pdrive_y_<3>.n0 VSS 2.51077f
C656 GF_NI_IN_C_BASE_0.pdrive_y_<3>.n1 VSS 1.27701f
C657 GF_NI_IN_C_BASE_0.pdrive_y_<3>.n2 VSS 0.913487f
C658 GF_NI_IN_C_BASE_0.pdrive_y_<3>.t1 VSS 0.13621f
C659 GF_NI_IN_C_BASE_0.pdrive_y_<3>.t4 VSS 6.32474f
C660 GF_NI_IN_C_BASE_0.pdrive_x_<3>.t3 VSS 1.61065f
C661 GF_NI_IN_C_BASE_0.pdrive_x_<3>.n0 VSS 2.36388f
C662 GF_NI_IN_C_BASE_0.pdrive_x_<3>.n1 VSS 1.88831f
C663 GF_NI_IN_C_BASE_0.pdrive_x_<3>.n2 VSS 1.37203f
C664 GF_NI_IN_C_BASE_0.pdrive_x_<3>.t0 VSS 0.99663f
C665 GF_NI_IN_C_BASE_0.pdrive_x_<3>.t1 VSS 0.803601f
C666 GF_NI_IN_C_BASE_0.pdrive_x_<3>.t2 VSS 0.136052f
C667 GF_NI_IN_C_BASE_0.pdrive_x_<3>.t5 VSS 6.08062f
C668 GF_NI_IN_C_BASE_0.pdrive_x_<3>.t4 VSS 6.00179f
C669 GF_NI_IN_C_BASE_0.pdrive_x_<3>.n3 VSS 33.0065f
C670 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_logic_pupd_0.PUB_OUT.t0 VSS 0.924776f
C671 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_logic_pupd_0.PUB_OUT.t1 VSS 0.146537f
C672 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_2.A VSS 0.561385f
C673 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_logic_pupd_0.PUB_OUT.t3 VSS 0.134163f
C674 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_logic_pupd_0.PUB_OUT.t2 VSS 0.089926f
C675 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_logic_pupd_0.PUB_OUT.n0 VSS 0.143212f
C676 GF_NI_IN_C_BASE_0.pdrive_y_<0>.t0 VSS 1.26541f
C677 GF_NI_IN_C_BASE_0.pdrive_y_<0>.t2 VSS 1.26004f
C678 GF_NI_IN_C_BASE_0.pdrive_y_<0>.t3 VSS 1.61704f
C679 GF_NI_IN_C_BASE_0.pdrive_y_<0>.n0 VSS 2.51778f
C680 GF_NI_IN_C_BASE_0.pdrive_y_<0>.n1 VSS 1.28058f
C681 GF_NI_IN_C_BASE_0.pdrive_y_<0>.n2 VSS 0.915927f
C682 GF_NI_IN_C_BASE_0.pdrive_y_<0>.t1 VSS 0.136591f
C683 GF_NI_IN_C_BASE_0.pdrive_y_<0>.t4 VSS 6.34406f
C684 GF_NI_IN_C_BASE_0.ndrive_x_<1>.t1 VSS 1.08312f
C685 GF_NI_IN_C_BASE_0.ndrive_x_<1>.t2 VSS 1.38999f
C686 GF_NI_IN_C_BASE_0.ndrive_x_<1>.n0 VSS 1.80704f
C687 GF_NI_IN_C_BASE_0.ndrive_x_<1>.t0 VSS 0.114393f
C688 GF_NI_IN_C_BASE_0.ndrive_x_<1>.n1 VSS 1.84967f
C689 GF_NI_IN_C_BASE_0.ndrive_x_<1>.t3 VSS 12.944799f
C690 GF_NI_IN_C_BASE_0.ndrive_y_<2>.t3 VSS 1.01484f
C691 GF_NI_IN_C_BASE_0.ndrive_y_<2>.t0 VSS 0.10226f
C692 GF_NI_IN_C_BASE_0.ndrive_y_<2>.n0 VSS 0.746002f
C693 GF_NI_IN_C_BASE_0.ndrive_y_<2>.t5 VSS 12.126599f
C694 GF_NI_IN_C_BASE_0.ndrive_y_<2>.t2 VSS 1.13289f
C695 GF_NI_IN_C_BASE_0.ndrive_y_<2>.n1 VSS 3.49749f
C696 GF_NI_IN_C_BASE_0.ndrive_y_<2>.n2 VSS 0.805369f
C697 GF_NI_IN_C_BASE_0.ndrive_y_<2>.t4 VSS 2.56725f
C698 GF_NI_IN_C_BASE_0.ndrive_y_<2>.n3 VSS 1.27451f
C699 GF_NI_IN_C_BASE_0.ndrive_y_<2>.t1 VSS 1.30236f
C700 GF_NI_IN_C_BASE_0.ndrive_y_<2>.n4 VSS 1.19632f
C701 GF_NI_IN_C_BASE_0.ndrive_x_<3>.t0 VSS 1.05175f
C702 GF_NI_IN_C_BASE_0.ndrive_x_<3>.t2 VSS 1.34973f
C703 GF_NI_IN_C_BASE_0.ndrive_x_<3>.n0 VSS 1.7547f
C704 GF_NI_IN_C_BASE_0.ndrive_x_<3>.t1 VSS 0.111079f
C705 GF_NI_IN_C_BASE_0.ndrive_x_<3>.n1 VSS 1.79609f
C706 GF_NI_IN_C_BASE_0.ndrive_x_<3>.t3 VSS 12.4708f
C707 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_cms_smt_0.nmos_6p0_CDNS_4066195314530_0.D.n0 VSS 0.131232f
C708 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_cms_smt_0.nmos_6p0_CDNS_4066195314530_0.D.t2 VSS 0.097441f
C709 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_cms_smt_0.nmos_6p0_CDNS_4066195314530_0.D.t1 VSS 0.418367f
C710 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_cms_smt_0.nmos_6p0_CDNS_4066195314530_0.D.t0 VSS 0.035864f
C711 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_pupd_0.PD.t0 VSS 0.162139f
C712 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_pupd_0.PD.t1 VSS 0.477818f
C713 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_pupd_0.PD.t2 VSS 0.256771f
C714 GF_NI_IN_C_BASE_0.comp018green_out_predrv_3.nmos_6p0_CDNS_4066195314519_0.D.t2 VSS 1.55639f
C715 GF_NI_IN_C_BASE_0.comp018green_out_predrv_3.nmos_6p0_CDNS_4066195314519_0.D.t0 VSS 1.49904f
C716 GF_NI_IN_C_BASE_0.comp018green_out_predrv_3.nmos_6p0_CDNS_4066195314519_0.D.t1 VSS 1.87506f
C717 GF_NI_IN_C_BASE_0.comp018green_out_predrv_3.nmos_6p0_CDNS_4066195314519_0.D.t4 VSS 1.23679f
C718 GF_NI_IN_C_BASE_0.comp018green_out_predrv_3.nmos_6p0_CDNS_4066195314519_0.D.t3 VSS 1.35457f
C719 GF_NI_IN_C_BASE_0.comp018green_out_predrv_3.nmos_6p0_CDNS_4066195314519_0.D.n0 VSS 0.969197f
C720 GF_NI_IN_C_BASE_0.comp018green_out_predrv_3.nmos_6p0_CDNS_4066195314519_0.D.t6 VSS 1.23679f
C721 GF_NI_IN_C_BASE_0.comp018green_out_predrv_3.nmos_6p0_CDNS_4066195314519_0.D.t8 VSS 1.35457f
C722 GF_NI_IN_C_BASE_0.comp018green_out_predrv_3.nmos_6p0_CDNS_4066195314519_0.D.n1 VSS 0.969197f
C723 GF_NI_IN_C_BASE_0.comp018green_out_predrv_3.nmos_6p0_CDNS_4066195314519_0.D.n2 VSS 0.255239f
C724 GF_NI_IN_C_BASE_0.comp018green_out_predrv_3.nmos_6p0_CDNS_4066195314519_0.D.n3 VSS 1.17912f
C725 GF_NI_IN_C_BASE_0.comp018green_out_predrv_3.nmos_6p0_CDNS_4066195314519_0.D.t7 VSS 0.624028f
C726 GF_NI_IN_C_BASE_0.comp018green_out_predrv_3.nmos_6p0_CDNS_4066195314519_0.D.t5 VSS 0.718195f
C727 GF_NI_IN_C_BASE_0.comp018green_out_predrv_3.nmos_6p0_CDNS_4066195314519_0.D.n4 VSS 0.810212f
C728 GF_NI_IN_C_BASE_0.ndrive_Y_<3>.t0 VSS 0.94601f
C729 GF_NI_IN_C_BASE_0.ndrive_Y_<3>.t2 VSS 1.21403f
C730 GF_NI_IN_C_BASE_0.ndrive_Y_<3>.n0 VSS 1.11518f
C731 GF_NI_IN_C_BASE_0.ndrive_Y_<3>.t1 VSS 2.39313f
C732 GF_NI_IN_C_BASE_0.ndrive_Y_<3>.t3 VSS 0.095324f
C733 GF_NI_IN_C_BASE_0.ndrive_Y_<3>.n1 VSS 0.695405f
C734 GF_NI_IN_C_BASE_0.ndrive_Y_<3>.t4 VSS 2.20897f
C735 GF_NI_IN_C_BASE_0.ndrive_Y_<3>.n2 VSS 1.03087f
C736 GF_NI_IN_C_BASE_0.ndrive_Y_<3>.n3 VSS 1.18807f
C737 GF_NI_IN_C_BASE_0.ndrive_Y_<3>.t5 VSS 10.826099f
C738 GF_NI_IN_C_BASE_0.comp018green_out_predrv_1.nmos_6p0_CDNS_4066195314519_2.S.t1 VSS 1.33525f
C739 GF_NI_IN_C_BASE_0.comp018green_out_predrv_1.nmos_6p0_CDNS_4066195314519_2.S.t0 VSS 1.13112f
C740 GF_NI_IN_C_BASE_0.comp018green_out_predrv_1.nmos_6p0_CDNS_4066195314519_2.S.n0 VSS 0.741389f
C741 GF_NI_IN_C_BASE_0.comp018green_out_predrv_1.nmos_6p0_CDNS_4066195314519_2.S.t7 VSS 0.433086f
C742 GF_NI_IN_C_BASE_0.comp018green_out_predrv_1.nmos_6p0_CDNS_4066195314519_2.S.t4 VSS 0.433086f
C743 GF_NI_IN_C_BASE_0.comp018green_out_predrv_1.nmos_6p0_CDNS_4066195314519_2.S.t3 VSS 0.433086f
C744 GF_NI_IN_C_BASE_0.comp018green_out_predrv_1.nmos_6p0_CDNS_4066195314519_2.S.t6 VSS 0.433086f
C745 GF_NI_IN_C_BASE_0.comp018green_out_predrv_1.nmos_6p0_CDNS_4066195314519_2.S.t5 VSS 0.93609f
C746 GF_NI_IN_C_BASE_0.comp018green_out_predrv_1.nmos_6p0_CDNS_4066195314519_2.S.t2 VSS 0.931295f
C747 GF_NI_IN_C_BASE_0.comp018green_out_predrv_1.nmos_6p0_CDNS_4066195314519_2.S.n1 VSS 0.993039f
C748 GF_NI_IN_C_BASE_0.comp018green_out_predrv_1.nmos_6p0_CDNS_4066195314519_2.S.n2 VSS 0.464839f
C749 GF_NI_IN_C_BASE_0.comp018green_out_predrv_1.nmos_6p0_CDNS_4066195314519_2.S.n3 VSS 0.299319f
C750 GF_NI_IN_C_BASE_0.comp018green_out_predrv_1.nmos_6p0_CDNS_4066195314519_2.S.n4 VSS 0.299319f
C751 GF_NI_IN_C_BASE_0.comp018green_out_predrv_1.nmos_6p0_CDNS_4066195314519_2.S.n5 VSS 0.442492f
C752 GF_NI_IN_C_BASE_0.comp018green_out_predrv_1.nmos_6p0_CDNS_4066195314519_2.S.n6 VSS 0.576756f
C753 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_3.Z.n0 VSS 1.82434f
C754 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_3.Z.t0 VSS 0.228818f
C755 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_3.Z.t8 VSS 0.308392f
C756 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_3.Z.t2 VSS 0.302472f
C757 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_3.Z.n1 VSS 1.36191f
C758 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_3.Z.t5 VSS 0.325049f
C759 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_3.Z.t1 VSS 0.321259f
C760 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_3.Z.t10 VSS 0.404429f
C761 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_3.Z.t11 VSS 0.76375f
C762 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_3.Z.n2 VSS 0.644041f
C763 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_3.Z.t6 VSS 0.404429f
C764 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_3.Z.t7 VSS 0.76375f
C765 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_3.Z.n3 VSS 0.646847f
C766 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_3.Z.t3 VSS 0.631504f
C767 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_3.Z.t9 VSS 0.358296f
C768 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_3.Z.t12 VSS 0.631504f
C769 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_3.Z.t4 VSS 0.358296f
C770 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_3.Z.n4 VSS 0.915343f
C771 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_3.Z.n5 VSS 0.909193f
C772 GF_NI_IN_C_BASE_0.pdrive_y_<2>.t0 VSS 1.24183f
C773 GF_NI_IN_C_BASE_0.pdrive_y_<2>.t2 VSS 1.23656f
C774 GF_NI_IN_C_BASE_0.pdrive_y_<2>.t3 VSS 1.58691f
C775 GF_NI_IN_C_BASE_0.pdrive_y_<2>.n0 VSS 2.47086f
C776 GF_NI_IN_C_BASE_0.pdrive_y_<2>.n1 VSS 1.25671f
C777 GF_NI_IN_C_BASE_0.pdrive_y_<2>.n2 VSS 0.898858f
C778 GF_NI_IN_C_BASE_0.pdrive_y_<2>.t1 VSS 0.134046f
C779 GF_NI_IN_C_BASE_0.pdrive_y_<2>.t4 VSS 6.27852f
C780 GF_NI_IN_C_BASE_0.comp018green_out_predrv_2.nmos_6p0_CDNS_4066195314519_0.D.t2 VSS 1.55629f
C781 GF_NI_IN_C_BASE_0.comp018green_out_predrv_2.nmos_6p0_CDNS_4066195314519_0.D.t1 VSS 1.49904f
C782 GF_NI_IN_C_BASE_0.comp018green_out_predrv_2.nmos_6p0_CDNS_4066195314519_0.D.t8 VSS 1.23679f
C783 GF_NI_IN_C_BASE_0.comp018green_out_predrv_2.nmos_6p0_CDNS_4066195314519_0.D.t5 VSS 1.35457f
C784 GF_NI_IN_C_BASE_0.comp018green_out_predrv_2.nmos_6p0_CDNS_4066195314519_0.D.n0 VSS 0.969197f
C785 GF_NI_IN_C_BASE_0.comp018green_out_predrv_2.nmos_6p0_CDNS_4066195314519_0.D.t3 VSS 1.23679f
C786 GF_NI_IN_C_BASE_0.comp018green_out_predrv_2.nmos_6p0_CDNS_4066195314519_0.D.t4 VSS 1.35457f
C787 GF_NI_IN_C_BASE_0.comp018green_out_predrv_2.nmos_6p0_CDNS_4066195314519_0.D.n1 VSS 0.969197f
C788 GF_NI_IN_C_BASE_0.comp018green_out_predrv_2.nmos_6p0_CDNS_4066195314519_0.D.n2 VSS 0.255239f
C789 GF_NI_IN_C_BASE_0.comp018green_out_predrv_2.nmos_6p0_CDNS_4066195314519_0.D.t0 VSS 1.87506f
C790 GF_NI_IN_C_BASE_0.comp018green_out_predrv_2.nmos_6p0_CDNS_4066195314519_0.D.n3 VSS 1.17912f
C791 GF_NI_IN_C_BASE_0.comp018green_out_predrv_2.nmos_6p0_CDNS_4066195314519_0.D.t7 VSS 0.624028f
C792 GF_NI_IN_C_BASE_0.comp018green_out_predrv_2.nmos_6p0_CDNS_4066195314519_0.D.t6 VSS 0.718195f
C793 GF_NI_IN_C_BASE_0.comp018green_out_predrv_2.nmos_6p0_CDNS_4066195314519_0.D.n4 VSS 0.810212f
C794 GF_NI_IN_C_BASE_0.comp018green_out_predrv_0.nmos_6p0_CDNS_4066195314519_0.D.t0 VSS 1.57587f
C795 GF_NI_IN_C_BASE_0.comp018green_out_predrv_0.nmos_6p0_CDNS_4066195314519_0.D.t2 VSS 1.51789f
C796 GF_NI_IN_C_BASE_0.comp018green_out_predrv_0.nmos_6p0_CDNS_4066195314519_0.D.t7 VSS 1.25234f
C797 GF_NI_IN_C_BASE_0.comp018green_out_predrv_0.nmos_6p0_CDNS_4066195314519_0.D.t3 VSS 1.37161f
C798 GF_NI_IN_C_BASE_0.comp018green_out_predrv_0.nmos_6p0_CDNS_4066195314519_0.D.n0 VSS 0.981388f
C799 GF_NI_IN_C_BASE_0.comp018green_out_predrv_0.nmos_6p0_CDNS_4066195314519_0.D.t8 VSS 1.25234f
C800 GF_NI_IN_C_BASE_0.comp018green_out_predrv_0.nmos_6p0_CDNS_4066195314519_0.D.t4 VSS 1.37161f
C801 GF_NI_IN_C_BASE_0.comp018green_out_predrv_0.nmos_6p0_CDNS_4066195314519_0.D.n1 VSS 0.981388f
C802 GF_NI_IN_C_BASE_0.comp018green_out_predrv_0.nmos_6p0_CDNS_4066195314519_0.D.n2 VSS 0.25845f
C803 GF_NI_IN_C_BASE_0.comp018green_out_predrv_0.nmos_6p0_CDNS_4066195314519_0.D.t1 VSS 1.89864f
C804 GF_NI_IN_C_BASE_0.comp018green_out_predrv_0.nmos_6p0_CDNS_4066195314519_0.D.n3 VSS 1.19395f
C805 GF_NI_IN_C_BASE_0.comp018green_out_predrv_0.nmos_6p0_CDNS_4066195314519_0.D.t6 VSS 0.631878f
C806 GF_NI_IN_C_BASE_0.comp018green_out_predrv_0.nmos_6p0_CDNS_4066195314519_0.D.t5 VSS 0.727229f
C807 GF_NI_IN_C_BASE_0.comp018green_out_predrv_0.nmos_6p0_CDNS_4066195314519_0.D.n4 VSS 0.820403f
C808 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_pupd_0.PU_B.t1 VSS 0.51572f
C809 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_pupd_0.PU_B.t0 VSS 0.181706f
C810 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_pupd_0.PU_B.t2 VSS 0.418935f
C811 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_pupd_0.PU_B.t3 VSS 0.50148f
C812 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_pupd_0.PU_B.t5 VSS 0.284525f
C813 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_pupd_0.PU_B.t4 VSS 0.50148f
C814 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_pupd_0.PU_B.t6 VSS 0.284525f
C815 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_pupd_0.PU_B.n0 VSS 0.726879f
C816 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_pupd_0.PU_B.n1 VSS 0.721995f
C817 GF_NI_IN_C_BASE_0.pdrive_x_<0>.t3 VSS 3.96081f
C818 GF_NI_IN_C_BASE_0.pdrive_x_<0>.t0 VSS 0.800753f
C819 GF_NI_IN_C_BASE_0.pdrive_x_<0>.t1 VSS 0.70782f
C820 GF_NI_IN_C_BASE_0.pdrive_x_<0>.n0 VSS 1.65277f
C821 GF_NI_IN_C_BASE_0.pdrive_x_<0>.n1 VSS 1.88173f
C822 GF_NI_IN_C_BASE_0.pdrive_x_<0>.t2 VSS 0.135582f
C823 GF_NI_IN_C_BASE_0.pdrive_x_<0>.t5 VSS 5.98219f
C824 GF_NI_IN_C_BASE_0.pdrive_x_<0>.t4 VSS 6.05673f
C825 GF_NI_IN_C_BASE_0.pdrive_x_<0>.n2 VSS 32.894302f
C826 GF_NI_IN_C_BASE_0.ndrive_y_<0>.t0 VSS 0.978804f
C827 GF_NI_IN_C_BASE_0.ndrive_y_<0>.t2 VSS 1.25612f
C828 GF_NI_IN_C_BASE_0.ndrive_y_<0>.n0 VSS 1.15384f
C829 GF_NI_IN_C_BASE_0.ndrive_y_<0>.t3 VSS 0.098628f
C830 GF_NI_IN_C_BASE_0.ndrive_y_<0>.n1 VSS 0.719511f
C831 GF_NI_IN_C_BASE_0.ndrive_y_<0>.t5 VSS 11.609401f
C832 GF_NI_IN_C_BASE_0.ndrive_y_<0>.t4 VSS 1.09267f
C833 GF_NI_IN_C_BASE_0.ndrive_y_<0>.n2 VSS 1.57958f
C834 GF_NI_IN_C_BASE_0.ndrive_y_<0>.n3 VSS 0.77677f
C835 GF_NI_IN_C_BASE_0.ndrive_y_<0>.t1 VSS 2.47609f
C836 GF_NI_IN_C_BASE_0.ndrive_y_<0>.n4 VSS 1.22926f
C837 GF_NI_IN_C_BASE_0.comp018green_out_predrv_0.nmos_6p0_CDNS_4066195314519_2.S.t1 VSS 1.33525f
C838 GF_NI_IN_C_BASE_0.comp018green_out_predrv_0.nmos_6p0_CDNS_4066195314519_2.S.t0 VSS 1.13112f
C839 GF_NI_IN_C_BASE_0.comp018green_out_predrv_0.nmos_6p0_CDNS_4066195314519_2.S.n0 VSS 0.741389f
C840 GF_NI_IN_C_BASE_0.comp018green_out_predrv_0.nmos_6p0_CDNS_4066195314519_2.S.t2 VSS 0.433086f
C841 GF_NI_IN_C_BASE_0.comp018green_out_predrv_0.nmos_6p0_CDNS_4066195314519_2.S.t3 VSS 0.433086f
C842 GF_NI_IN_C_BASE_0.comp018green_out_predrv_0.nmos_6p0_CDNS_4066195314519_2.S.t5 VSS 0.433086f
C843 GF_NI_IN_C_BASE_0.comp018green_out_predrv_0.nmos_6p0_CDNS_4066195314519_2.S.t7 VSS 0.433086f
C844 GF_NI_IN_C_BASE_0.comp018green_out_predrv_0.nmos_6p0_CDNS_4066195314519_2.S.t4 VSS 0.931295f
C845 GF_NI_IN_C_BASE_0.comp018green_out_predrv_0.nmos_6p0_CDNS_4066195314519_2.S.t6 VSS 0.93609f
C846 GF_NI_IN_C_BASE_0.comp018green_out_predrv_0.nmos_6p0_CDNS_4066195314519_2.S.n1 VSS 0.993039f
C847 GF_NI_IN_C_BASE_0.comp018green_out_predrv_0.nmos_6p0_CDNS_4066195314519_2.S.n2 VSS 0.464839f
C848 GF_NI_IN_C_BASE_0.comp018green_out_predrv_0.nmos_6p0_CDNS_4066195314519_2.S.n3 VSS 0.299319f
C849 GF_NI_IN_C_BASE_0.comp018green_out_predrv_0.nmos_6p0_CDNS_4066195314519_2.S.n4 VSS 0.299319f
C850 GF_NI_IN_C_BASE_0.comp018green_out_predrv_0.nmos_6p0_CDNS_4066195314519_2.S.n5 VSS 0.442492f
C851 GF_NI_IN_C_BASE_0.comp018green_out_predrv_0.nmos_6p0_CDNS_4066195314519_2.S.n6 VSS 0.576756f
C852 GF_NI_IN_C_BASE_0.pdrive_x_<2>.t3 VSS 3.87079f
C853 GF_NI_IN_C_BASE_0.pdrive_x_<2>.t0 VSS 0.782832f
C854 GF_NI_IN_C_BASE_0.pdrive_x_<2>.t1 VSS 0.691979f
C855 GF_NI_IN_C_BASE_0.pdrive_x_<2>.n0 VSS 1.61579f
C856 GF_NI_IN_C_BASE_0.pdrive_x_<2>.n1 VSS 1.83962f
C857 GF_NI_IN_C_BASE_0.pdrive_x_<2>.t2 VSS 0.132547f
C858 GF_NI_IN_C_BASE_0.pdrive_x_<2>.t4 VSS 5.82992f
C859 GF_NI_IN_C_BASE_0.pdrive_x_<2>.t5 VSS 5.94087f
C860 GF_NI_IN_C_BASE_0.pdrive_x_<2>.n2 VSS 32.157803f
C861 GF_NI_IN_C_BASE_0.comp018green_out_predrv_0.SL.n0 VSS 5.05896f
C862 GF_NI_IN_C_BASE_0.comp018green_out_predrv_0.SL.t1 VSS 0.387109f
C863 GF_NI_IN_C_BASE_0.comp018green_out_predrv_0.SL.t2 VSS 0.48626f
C864 GF_NI_IN_C_BASE_0.comp018green_out_predrv_0.SL.t9 VSS 0.27589f
C865 GF_NI_IN_C_BASE_0.comp018green_out_predrv_0.SL.t8 VSS 0.48626f
C866 GF_NI_IN_C_BASE_0.comp018green_out_predrv_0.SL.t6 VSS 0.27589f
C867 GF_NI_IN_C_BASE_0.comp018green_out_predrv_0.SL.n1 VSS 0.704818f
C868 GF_NI_IN_C_BASE_0.comp018green_out_predrv_0.SL.n2 VSS 0.698682f
C869 GF_NI_IN_C_BASE_0.comp018green_out_predrv_0.SL.t3 VSS 1.51298f
C870 GF_NI_IN_C_BASE_0.comp018green_out_predrv_0.SL.t10 VSS 1.50265f
C871 GF_NI_IN_C_BASE_0.comp018green_out_predrv_0.SL.n3 VSS 1.24529f
C872 GF_NI_IN_C_BASE_0.comp018green_out_predrv_0.SL.t12 VSS 1.50265f
C873 GF_NI_IN_C_BASE_0.comp018green_out_predrv_0.SL.t13 VSS 1.51298f
C874 GF_NI_IN_C_BASE_0.comp018green_out_predrv_0.SL.n4 VSS 1.24529f
C875 GF_NI_IN_C_BASE_0.comp018green_out_predrv_0.SL.t11 VSS 1.51298f
C876 GF_NI_IN_C_BASE_0.comp018green_out_predrv_0.SL.t5 VSS 1.50265f
C877 GF_NI_IN_C_BASE_0.comp018green_out_predrv_0.SL.n5 VSS 1.24529f
C878 GF_NI_IN_C_BASE_0.comp018green_out_predrv_0.SL.t4 VSS 1.50265f
C879 GF_NI_IN_C_BASE_0.comp018green_out_predrv_0.SL.t7 VSS 1.51298f
C880 GF_NI_IN_C_BASE_0.comp018green_out_predrv_0.SL.n6 VSS 1.24529f
C881 GF_NI_IN_C_BASE_0.comp018green_out_predrv_0.SL.n7 VSS 2.53456f
C882 GF_NI_IN_C_BASE_0.comp018green_out_predrv_0.SL.t0 VSS 0.131137f
C883 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_logic_pupd_0.PDB_OUT.t0 VSS 4.43443f
C884 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_0.A VSS 2.41435f
C885 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_logic_pupd_0.PDB_OUT.t1 VSS 0.457031f
C886 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_logic_pupd_0.PDB_OUT.t2 VSS 0.306336f
C887 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_logic_pupd_0.PDB_OUT.n0 VSS 0.487855f
C888 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_1.EN.t6 VSS 0.923628f
C889 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_1.EN.t2 VSS 1.86913f
C890 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_1.EN.t7 VSS 0.923628f
C891 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_1.EN.t3 VSS 1.86913f
C892 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_1.EN.n0 VSS 3.58291f
C893 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_1.EN.t0 VSS 0.361015f
C894 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_1.EN.t1 VSS 0.88331f
C895 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_1.EN.t5 VSS 0.938193f
C896 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_1.EN.t4 VSS 0.502091f
C897 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_1.EN.n1 VSS 0.667727f
C898 GF_NI_IN_C_BASE_0.ndrive_x_<0>.t0 VSS 2.97732f
C899 GF_NI_IN_C_BASE_0.ndrive_x_<0>.t2 VSS 0.736166f
C900 GF_NI_IN_C_BASE_0.ndrive_x_<0>.t1 VSS 0.106531f
C901 GF_NI_IN_C_BASE_0.ndrive_x_<0>.n0 VSS 1.72255f
C902 GF_NI_IN_C_BASE_0.ndrive_x_<0>.t3 VSS 11.547501f
C903 GF_NI_IN_C_BASE_0.ndrive_x_<2>.t0 VSS 2.93739f
C904 GF_NI_IN_C_BASE_0.ndrive_x_<2>.t2 VSS 0.726293f
C905 GF_NI_IN_C_BASE_0.ndrive_x_<2>.t1 VSS 0.105102f
C906 GF_NI_IN_C_BASE_0.ndrive_x_<2>.n0 VSS 1.69945f
C907 GF_NI_IN_C_BASE_0.ndrive_x_<2>.t3 VSS 12.238501f
C908 GF_NI_IN_C_BASE_0.comp018green_out_predrv_2.nmos_6p0_CDNS_4066195314519_2.S.t0 VSS 1.29746f
C909 GF_NI_IN_C_BASE_0.comp018green_out_predrv_2.nmos_6p0_CDNS_4066195314519_2.S.t1 VSS 1.09911f
C910 GF_NI_IN_C_BASE_0.comp018green_out_predrv_2.nmos_6p0_CDNS_4066195314519_2.S.n0 VSS 0.720406f
C911 GF_NI_IN_C_BASE_0.comp018green_out_predrv_2.nmos_6p0_CDNS_4066195314519_2.S.t3 VSS 0.420829f
C912 GF_NI_IN_C_BASE_0.comp018green_out_predrv_2.nmos_6p0_CDNS_4066195314519_2.S.t4 VSS 0.420829f
C913 GF_NI_IN_C_BASE_0.comp018green_out_predrv_2.nmos_6p0_CDNS_4066195314519_2.S.t7 VSS 0.420829f
C914 GF_NI_IN_C_BASE_0.comp018green_out_predrv_2.nmos_6p0_CDNS_4066195314519_2.S.t2 VSS 0.420829f
C915 GF_NI_IN_C_BASE_0.comp018green_out_predrv_2.nmos_6p0_CDNS_4066195314519_2.S.t5 VSS 0.904937f
C916 GF_NI_IN_C_BASE_0.comp018green_out_predrv_2.nmos_6p0_CDNS_4066195314519_2.S.t6 VSS 0.909597f
C917 GF_NI_IN_C_BASE_0.comp018green_out_predrv_2.nmos_6p0_CDNS_4066195314519_2.S.n1 VSS 0.964934f
C918 GF_NI_IN_C_BASE_0.comp018green_out_predrv_2.nmos_6p0_CDNS_4066195314519_2.S.n2 VSS 0.451683f
C919 GF_NI_IN_C_BASE_0.comp018green_out_predrv_2.nmos_6p0_CDNS_4066195314519_2.S.n3 VSS 0.290848f
C920 GF_NI_IN_C_BASE_0.comp018green_out_predrv_2.nmos_6p0_CDNS_4066195314519_2.S.n4 VSS 0.290848f
C921 GF_NI_IN_C_BASE_0.comp018green_out_predrv_2.nmos_6p0_CDNS_4066195314519_2.S.n5 VSS 0.429969f
C922 GF_NI_IN_C_BASE_0.comp018green_out_predrv_2.nmos_6p0_CDNS_4066195314519_2.S.n6 VSS 0.560433f
C923 GF_NI_IN_C_BASE_0.ndrive_Y_<1>.t3 VSS 0.93914f
C924 GF_NI_IN_C_BASE_0.ndrive_Y_<1>.t4 VSS 2.37575f
C925 GF_NI_IN_C_BASE_0.ndrive_Y_<1>.t1 VSS 0.094632f
C926 GF_NI_IN_C_BASE_0.ndrive_Y_<1>.n0 VSS 0.690355f
C927 GF_NI_IN_C_BASE_0.ndrive_Y_<1>.t2 VSS 2.19293f
C928 GF_NI_IN_C_BASE_0.ndrive_Y_<1>.n1 VSS 1.02339f
C929 GF_NI_IN_C_BASE_0.ndrive_Y_<1>.n2 VSS 1.17944f
C930 GF_NI_IN_C_BASE_0.ndrive_Y_<1>.t0 VSS 1.20522f
C931 GF_NI_IN_C_BASE_0.ndrive_Y_<1>.n3 VSS 1.10708f
C932 GF_NI_IN_C_BASE_0.ndrive_Y_<1>.t5 VSS 11.5531f
C933 GF_NI_IN_C_BASE_0.comp018green_out_predrv_3.nmos_6p0_CDNS_4066195314519_2.S.t0 VSS 1.28486f
C934 GF_NI_IN_C_BASE_0.comp018green_out_predrv_3.nmos_6p0_CDNS_4066195314519_2.S.t1 VSS 1.08844f
C935 GF_NI_IN_C_BASE_0.comp018green_out_predrv_3.nmos_6p0_CDNS_4066195314519_2.S.n0 VSS 0.713412f
C936 GF_NI_IN_C_BASE_0.comp018green_out_predrv_3.nmos_6p0_CDNS_4066195314519_2.S.t4 VSS 0.416743f
C937 GF_NI_IN_C_BASE_0.comp018green_out_predrv_3.nmos_6p0_CDNS_4066195314519_2.S.t7 VSS 0.416743f
C938 GF_NI_IN_C_BASE_0.comp018green_out_predrv_3.nmos_6p0_CDNS_4066195314519_2.S.t6 VSS 0.416743f
C939 GF_NI_IN_C_BASE_0.comp018green_out_predrv_3.nmos_6p0_CDNS_4066195314519_2.S.t3 VSS 0.416743f
C940 GF_NI_IN_C_BASE_0.comp018green_out_predrv_3.nmos_6p0_CDNS_4066195314519_2.S.t2 VSS 0.900766f
C941 GF_NI_IN_C_BASE_0.comp018green_out_predrv_3.nmos_6p0_CDNS_4066195314519_2.S.t5 VSS 0.896151f
C942 GF_NI_IN_C_BASE_0.comp018green_out_predrv_3.nmos_6p0_CDNS_4066195314519_2.S.n1 VSS 0.955566f
C943 GF_NI_IN_C_BASE_0.comp018green_out_predrv_3.nmos_6p0_CDNS_4066195314519_2.S.n2 VSS 0.447298f
C944 GF_NI_IN_C_BASE_0.comp018green_out_predrv_3.nmos_6p0_CDNS_4066195314519_2.S.n3 VSS 0.288024f
C945 GF_NI_IN_C_BASE_0.comp018green_out_predrv_3.nmos_6p0_CDNS_4066195314519_2.S.n4 VSS 0.288024f
C946 GF_NI_IN_C_BASE_0.comp018green_out_predrv_3.nmos_6p0_CDNS_4066195314519_2.S.n5 VSS 0.425794f
C947 GF_NI_IN_C_BASE_0.comp018green_out_predrv_3.nmos_6p0_CDNS_4066195314519_2.S.n6 VSS 0.554992f
C948 Y.t1 VSS 0.040502f
C949 Y.t5 VSS 0.040502f
C950 Y.n0 VSS 0.081775f
C951 Y.n1 VSS 0.046888f
C952 Y.t2 VSS 0.040502f
C953 Y.t0 VSS 0.040502f
C954 Y.n2 VSS 0.081775f
C955 Y.n3 VSS 0.046888f
C956 Y.t4 VSS 0.040502f
C957 Y.t3 VSS 0.040502f
C958 Y.n4 VSS 0.08178f
C959 Y.n5 VSS 0.170526f
C960 Y.n6 VSS 0.296406f
C961 Y.n7 VSS 0.290688f
C962 Y.t8 VSS 0.094506f
C963 Y.t6 VSS 0.094506f
C964 Y.n8 VSS 0.278921f
C965 Y.t9 VSS 0.094506f
C966 Y.t7 VSS 0.094506f
C967 Y.n9 VSS 0.278921f
C968 Y.t11 VSS 0.094506f
C969 Y.t10 VSS 0.094506f
C970 Y.n10 VSS 0.39267f
C971 Y.n11 VSS 0.62594f
C972 Y.n12 VSS 0.393669f
C973 Y.n13 VSS 1.41386f
C974 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_drv_0.nmos_6p0_CDNS_4066195314550_0.D VSS 1.49697f
C975 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_drv_0.Z.t0 VSS 0.063962f
C976 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_drv_0.Z.t9 VSS 0.169311f
C977 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_drv_0.Z.t8 VSS 0.221117f
C978 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_drv_0.Z.n0 VSS 0.251108f
C979 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_drv_0.Z.t1 VSS 0.169311f
C980 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_drv_0.Z.t12 VSS 0.221117f
C981 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_drv_0.Z.n1 VSS 0.249078f
C982 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_drv_0.Z.t5 VSS 0.169311f
C983 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_drv_0.Z.t3 VSS 0.221117f
C984 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_drv_0.Z.n2 VSS 0.249078f
C985 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_drv_0.Z.t4 VSS 0.169311f
C986 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_drv_0.Z.t2 VSS 0.221117f
C987 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_drv_0.Z.n3 VSS 0.249078f
C988 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_drv_0.Z.t11 VSS 0.169311f
C989 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_drv_0.Z.t10 VSS 0.221117f
C990 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_drv_0.Z.n4 VSS 0.249078f
C991 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_drv_0.Z.t7 VSS 0.169311f
C992 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_drv_0.Z.t6 VSS 0.221117f
C993 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_drv_0.Z.n5 VSS 0.249078f
C994 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_1.Z.n0 VSS 1.81515f
C995 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_1.Z.t1 VSS 0.365536f
C996 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_1.Z.n1 VSS 0.505169f
C997 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_1.Z.t5 VSS 0.355443f
C998 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_1.Z.t10 VSS 0.201668f
C999 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_1.Z.t4 VSS 0.355443f
C1000 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_1.Z.t9 VSS 0.201668f
C1001 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_1.Z.n2 VSS 0.515203f
C1002 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_1.Z.n3 VSS 0.511741f
C1003 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_1.Z.t0 VSS 0.128791f
C1004 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_1.Z.t7 VSS 0.31839f
C1005 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_1.Z.t6 VSS 0.2261f
C1006 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_1.Z.t13 VSS 0.226338f
C1007 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_1.Z.t8 VSS 0.22431f
C1008 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_1.Z.t2 VSS 0.317768f
C1009 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_1.Z.t3 VSS 0.317768f
C1010 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_1.Z.t11 VSS 0.317768f
C1011 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_1.Z.t12 VSS 0.317768f
C1012 PAD.t4 VSS 0.012458f
C1013 PAD.t21 VSS 0.028949f
C1014 PAD.n0 VSS 0.032683f
C1015 PAD.n1 VSS 0.037314f
C1016 PAD.n2 VSS 0.026049f
C1017 PAD.n3 VSS 0.013703f
C1018 PAD.t6 VSS 0.012458f
C1019 PAD.t15 VSS 0.012458f
C1020 PAD.n4 VSS 0.02649f
C1021 PAD.n5 VSS 0.030039f
C1022 PAD.n6 VSS 0.030039f
C1023 PAD.n7 VSS 0.026049f
C1024 PAD.n8 VSS 0.018379f
C1025 PAD.n9 VSS 0.024671f
C1026 PAD.n10 VSS 10.1398f
C1027 PAD.n11 VSS 12.7698f
C1028 PAD.n12 VSS 13.1442f
C1029 PAD.n13 VSS 14.504801f
C1030 PAD.n14 VSS 0.043265f
C1031 PAD.n15 VSS 0.062262f
C1032 PAD.n16 VSS 0.039754f
C1033 PAD.n17 VSS 0.069752f
C1034 PAD.n18 VSS 0.039754f
C1035 PAD.n19 VSS 0.069752f
C1036 PAD.n20 VSS 0.157837f
C1037 PAD.n21 VSS 0.596822f
C1038 PAD.n22 VSS 0.03925f
C1039 PAD.n23 VSS 0.029913f
C1040 PAD.n24 VSS 0.03925f
C1041 PAD.n25 VSS 0.029913f
C1042 PAD.n26 VSS 0.03055f
C1043 PAD.n27 VSS 0.042887f
C1044 PAD.n28 VSS 0.049106f
C1045 PAD.n29 VSS 0.029431f
C1046 PAD.n30 VSS 0.049106f
C1047 PAD.n31 VSS 0.029431f
C1048 PAD.n32 VSS 0.44885f
C1049 PAD.n74 VSS 0.023105f
C1050 PAD.n75 VSS 0.023105f
C1051 PAD.n76 VSS 0.036454f
C1052 PAD.n77 VSS 0.036454f
C1053 PAD.n78 VSS 0.036454f
C1054 PAD.n79 VSS 0.036454f
C1055 PAD.n80 VSS 0.036454f
C1056 PAD.n81 VSS 0.036454f
C1057 PAD.n82 VSS 0.036454f
C1058 PAD.n83 VSS 0.036454f
C1059 PAD.n84 VSS 0.036454f
C1060 PAD.n85 VSS 0.036454f
C1061 PAD.n86 VSS 0.036454f
C1062 PAD.n87 VSS 0.036454f
C1063 PAD.n88 VSS 0.036454f
C1064 PAD.n89 VSS 0.036454f
C1065 PAD.n90 VSS 0.036454f
C1066 PAD.n91 VSS 0.036454f
C1067 PAD.n92 VSS 0.036454f
C1068 PAD.n93 VSS 0.036454f
C1069 PAD.n94 VSS 0.036454f
C1070 PAD.n95 VSS 0.036454f
C1071 PAD.n96 VSS 0.036454f
C1072 PAD.n97 VSS 0.036454f
C1073 PAD.n98 VSS 0.036454f
C1074 PAD.n99 VSS 0.036454f
C1075 PAD.n100 VSS 0.036454f
C1076 PAD.n101 VSS 0.036454f
C1077 PAD.n102 VSS 0.036454f
C1078 PAD.n103 VSS 0.036454f
C1079 PAD.n104 VSS 0.036454f
C1080 PAD.n105 VSS 0.036454f
C1081 PAD.n106 VSS 0.036454f
C1082 PAD.n107 VSS 0.036454f
C1083 PAD.n108 VSS 0.036454f
C1084 PAD.n109 VSS 0.036454f
C1085 PAD.n110 VSS 0.036454f
C1086 PAD.n111 VSS 0.036454f
C1087 PAD.n112 VSS 0.036454f
C1088 PAD.n113 VSS 0.036454f
C1089 PAD.n114 VSS 0.036454f
C1090 PAD.n115 VSS 0.036454f
C1091 PAD.n117 VSS 0.036454f
C1092 PAD.n118 VSS 0.036454f
C1093 PAD.n119 VSS 0.023105f
C1094 PAD.n120 VSS 0.033374f
C1095 PAD.n121 VSS 0.036454f
C1096 PAD.n122 VSS 0.036454f
C1097 PAD.n123 VSS 0.036454f
C1098 PAD.n124 VSS 0.036454f
C1099 PAD.n126 VSS 0.036454f
C1100 PAD.n127 VSS 0.036454f
C1101 PAD.n128 VSS 0.036454f
C1102 PAD.n130 VSS 0.036454f
C1103 PAD.n131 VSS 0.036454f
C1104 PAD.n132 VSS 0.036454f
C1105 PAD.n133 VSS 0.036454f
C1106 PAD.n134 VSS 0.036454f
C1107 PAD.n135 VSS 0.036454f
C1108 PAD.n136 VSS 0.036454f
C1109 PAD.n138 VSS 0.036454f
C1110 PAD.n139 VSS 0.036454f
C1111 PAD.n140 VSS 0.036454f
C1112 PAD.n142 VSS 0.036454f
C1113 PAD.n143 VSS 0.036454f
C1114 PAD.n144 VSS 0.036454f
C1115 PAD.n145 VSS 0.036454f
C1116 PAD.n146 VSS 0.036454f
C1117 PAD.n147 VSS 0.036454f
C1118 PAD.n148 VSS 0.036454f
C1119 PAD.n150 VSS 0.036454f
C1120 PAD.n151 VSS 0.036454f
C1121 PAD.n152 VSS 0.036454f
C1122 PAD.n154 VSS 0.036454f
C1123 PAD.n155 VSS 0.036454f
C1124 PAD.n156 VSS 0.036454f
C1125 PAD.n157 VSS 0.036454f
C1126 PAD.n158 VSS 0.036454f
C1127 PAD.n159 VSS 0.036454f
C1128 PAD.n160 VSS 0.036454f
C1129 PAD.n162 VSS 0.036454f
C1130 PAD.n163 VSS 0.036454f
C1131 PAD.n164 VSS 0.036454f
C1132 PAD.n166 VSS 0.036454f
C1133 PAD.n167 VSS 0.036454f
C1134 PAD.n168 VSS 0.036454f
C1135 PAD.n169 VSS 0.036454f
C1136 PAD.n170 VSS 0.036454f
C1137 PAD.n171 VSS 0.036454f
C1138 PAD.n172 VSS 0.036454f
C1139 PAD.n174 VSS 0.036454f
C1140 PAD.n175 VSS 0.036454f
C1141 PAD.n176 VSS 0.036454f
C1142 PAD.n178 VSS 0.036454f
C1143 PAD.n179 VSS 0.036454f
C1144 PAD.n180 VSS 0.036454f
C1145 PAD.n181 VSS 0.036454f
C1146 PAD.n182 VSS 0.036454f
C1147 PAD.n183 VSS 0.036454f
C1148 PAD.n184 VSS 0.036454f
C1149 PAD.n186 VSS 0.036454f
C1150 PAD.n187 VSS 0.036454f
C1151 PAD.n188 VSS 0.036454f
C1152 PAD.n190 VSS 0.036454f
C1153 PAD.n191 VSS 0.036454f
C1154 PAD.n192 VSS 0.036454f
C1155 PAD.n193 VSS 0.036454f
C1156 PAD.n194 VSS 0.036454f
C1157 PAD.n195 VSS 0.036454f
C1158 PAD.n196 VSS 0.036454f
C1159 PAD.n198 VSS 0.036454f
C1160 PAD.n199 VSS 0.036454f
C1161 PAD.n200 VSS 0.036454f
C1162 PAD.n202 VSS 0.036454f
C1163 PAD.n203 VSS 0.036454f
C1164 PAD.n204 VSS 0.036454f
C1165 PAD.n205 VSS 0.036454f
C1166 PAD.n206 VSS 0.036454f
C1167 PAD.n207 VSS 0.036454f
C1168 PAD.n208 VSS 0.036454f
C1169 PAD.n210 VSS 0.036454f
C1170 PAD.n211 VSS 0.036454f
C1171 PAD.n212 VSS 0.036454f
C1172 PAD.n214 VSS 0.036454f
C1173 PAD.n215 VSS 0.036454f
C1174 PAD.n216 VSS 0.036454f
C1175 PAD.n217 VSS 0.036454f
C1176 PAD.n218 VSS 0.036454f
C1177 PAD.n219 VSS 0.036454f
C1178 PAD.n220 VSS 0.036454f
C1179 PAD.n222 VSS 0.036454f
C1180 PAD.n223 VSS 0.036454f
C1181 PAD.n224 VSS 0.036454f
C1182 PAD.n226 VSS 0.036454f
C1183 PAD.n227 VSS 0.036454f
C1184 PAD.n228 VSS 0.036454f
C1185 PAD.n229 VSS 0.036454f
C1186 PAD.n230 VSS 0.036454f
C1187 PAD.n231 VSS 0.036454f
C1188 PAD.n232 VSS 0.036454f
C1189 PAD.n234 VSS 0.036454f
C1190 PAD.n235 VSS 0.036454f
C1191 PAD.n236 VSS 0.036454f
C1192 PAD.n238 VSS 0.036454f
C1193 PAD.n239 VSS 0.036454f
C1194 PAD.n240 VSS 0.036454f
C1195 PAD.n241 VSS 0.036454f
C1196 PAD.n242 VSS 0.036454f
C1197 PAD.n243 VSS 0.036454f
C1198 PAD.n244 VSS 0.036454f
C1199 PAD.n246 VSS 0.036454f
C1200 PAD.n247 VSS 0.036454f
C1201 PAD.n248 VSS 0.036454f
C1202 PAD.n250 VSS 0.036454f
C1203 PAD.n251 VSS 0.036454f
C1204 PAD.n252 VSS 0.036454f
C1205 PAD.n253 VSS 0.036454f
C1206 PAD.n254 VSS 0.036454f
C1207 PAD.n255 VSS 0.036454f
C1208 PAD.n256 VSS 0.036454f
C1209 PAD.n258 VSS 0.036454f
C1210 PAD.n259 VSS 0.036454f
C1211 PAD.n260 VSS 0.036454f
C1212 PAD.n262 VSS 0.036454f
C1213 PAD.n263 VSS 0.036454f
C1214 PAD.n264 VSS 0.036454f
C1215 PAD.n265 VSS 0.036454f
C1216 PAD.n266 VSS 0.036454f
C1217 PAD.n267 VSS 0.036454f
C1218 PAD.n268 VSS 0.036454f
C1219 PAD.n270 VSS 0.036454f
C1220 PAD.n271 VSS 0.036454f
C1221 PAD.n272 VSS 0.036454f
C1222 PAD.n274 VSS 0.036454f
C1223 PAD.n275 VSS 0.036454f
C1224 PAD.n276 VSS 0.036454f
C1225 PAD.n277 VSS 0.036454f
C1226 PAD.n278 VSS 0.036454f
C1227 PAD.n279 VSS 0.036454f
C1228 PAD.n280 VSS 0.036454f
C1229 PAD.n282 VSS 0.036454f
C1230 PAD.n283 VSS 0.036454f
C1231 PAD.n284 VSS 0.036454f
C1232 PAD.n286 VSS 0.036454f
C1233 PAD.n287 VSS 0.036454f
C1234 PAD.n288 VSS 0.036454f
C1235 PAD.n289 VSS 0.036454f
C1236 PAD.n290 VSS 0.036454f
C1237 PAD.n291 VSS 0.036454f
C1238 PAD.n292 VSS 0.036454f
C1239 PAD.n294 VSS 0.036454f
C1240 PAD.n295 VSS 0.036454f
C1241 PAD.n296 VSS 0.036454f
C1242 PAD.n298 VSS 0.036454f
C1243 PAD.n299 VSS 0.036454f
C1244 PAD.n300 VSS 0.036454f
C1245 PAD.n301 VSS 0.036454f
C1246 PAD.n302 VSS 0.036454f
C1247 PAD.n303 VSS 0.036454f
C1248 PAD.n304 VSS 0.036454f
C1249 PAD.n306 VSS 0.036454f
C1250 PAD.n307 VSS 0.036454f
C1251 PAD.n308 VSS 0.036454f
C1252 PAD.n310 VSS 0.036454f
C1253 PAD.n311 VSS 0.036454f
C1254 PAD.n312 VSS 0.036454f
C1255 PAD.n313 VSS 0.036454f
C1256 PAD.n314 VSS 0.036454f
C1257 PAD.n315 VSS 0.036454f
C1258 PAD.n316 VSS 0.036454f
C1259 PAD.n318 VSS 0.036454f
C1260 PAD.n319 VSS 0.036454f
C1261 PAD.n320 VSS 0.036454f
C1262 PAD.n322 VSS 0.036454f
C1263 PAD.n323 VSS 0.036454f
C1264 PAD.n324 VSS 0.036454f
C1265 PAD.n325 VSS 0.036454f
C1266 PAD.n326 VSS 0.036454f
C1267 PAD.n327 VSS 0.036454f
C1268 PAD.n328 VSS 0.036454f
C1269 PAD.n330 VSS 0.036454f
C1270 PAD.n331 VSS 0.036454f
C1271 PAD.n332 VSS 0.036454f
C1272 PAD.n334 VSS 0.036454f
C1273 PAD.n335 VSS 0.036454f
C1274 PAD.n336 VSS 0.036454f
C1275 PAD.n337 VSS 0.036454f
C1276 PAD.n338 VSS 0.036454f
C1277 PAD.n339 VSS 0.036454f
C1278 PAD.n340 VSS 0.036454f
C1279 PAD.n342 VSS 0.036454f
C1280 PAD.n343 VSS 0.036454f
C1281 PAD.n344 VSS 0.036454f
C1282 PAD.n346 VSS 0.036454f
C1283 PAD.n347 VSS 0.036454f
C1284 PAD.n348 VSS 0.036454f
C1285 PAD.n349 VSS 0.036454f
C1286 PAD.n350 VSS 0.036454f
C1287 PAD.n351 VSS 0.036454f
C1288 PAD.n352 VSS 0.036454f
C1289 PAD.n354 VSS 0.036454f
C1290 PAD.n355 VSS 0.036454f
C1291 PAD.n356 VSS 0.036454f
C1292 PAD.n358 VSS 0.036454f
C1293 PAD.n359 VSS 0.036454f
C1294 PAD.n360 VSS 0.036454f
C1295 PAD.n361 VSS 0.036454f
C1296 PAD.n362 VSS 0.036454f
C1297 PAD.n363 VSS 0.036454f
C1298 PAD.n364 VSS 0.036454f
C1299 PAD.n366 VSS 0.023105f
C1300 PAD.n367 VSS 0.537633f
C1301 PAD.n368 VSS 0.069752f
C1302 PAD.n369 VSS 0.069752f
C1303 PAD.n370 VSS 0.032135f
C1304 PAD.n371 VSS 0.036001f
C1305 PAD.n372 VSS 0.036001f
C1306 PAD.n373 VSS 0.315674f
C1307 PAD.n415 VSS 0.023105f
C1308 PAD.n416 VSS 0.023105f
C1309 PAD.n417 VSS 0.029431f
C1310 PAD.n418 VSS 0.656011f
C1311 PAD.n419 VSS 0.42912f
C1312 PAD.n420 VSS 0.036454f
C1313 PAD.n421 VSS 0.036454f
C1314 PAD.n422 VSS 0.033978f
C1315 PAD.n423 VSS 0.049106f
C1316 PAD.n424 VSS 0.049106f
C1317 PAD.n425 VSS 0.611619f
C1318 PAD.n426 VSS 0.069752f
C1319 PAD.n427 VSS 0.039754f
C1320 PAD.n428 VSS 0.069752f
C1321 PAD.n429 VSS 0.039754f
C1322 PAD.n430 VSS 0.046278f
C1323 PAD.n431 VSS 0.039754f
C1324 PAD.n432 VSS 0.039754f
C1325 PAD.n433 VSS 0.611619f
C1326 PAD.n434 VSS 0.512971f
C1327 PAD.n435 VSS 0.606687f
C1328 PAD.n436 VSS 0.029431f
C1329 PAD.n437 VSS 0.029431f
C1330 PAD.n438 VSS 0.036454f
C1331 PAD.n439 VSS 0.036454f
C1332 PAD.n440 VSS 0.036454f
C1333 PAD.n442 VSS 0.036454f
C1334 PAD.n443 VSS 0.036454f
C1335 PAD.n444 VSS 0.036454f
C1336 PAD.n446 VSS 0.036454f
C1337 PAD.n447 VSS 0.036454f
C1338 PAD.n448 VSS 0.036454f
C1339 PAD.n450 VSS 0.036454f
C1340 PAD.n451 VSS 0.036454f
C1341 PAD.n452 VSS 0.036454f
C1342 PAD.n454 VSS 0.036454f
C1343 PAD.n455 VSS 0.036454f
C1344 PAD.n456 VSS 0.036454f
C1345 PAD.n458 VSS 0.036454f
C1346 PAD.n459 VSS 0.036454f
C1347 PAD.n460 VSS 0.036454f
C1348 PAD.n462 VSS 0.036454f
C1349 PAD.n463 VSS 0.036454f
C1350 PAD.n464 VSS 0.036454f
C1351 PAD.n466 VSS 0.036454f
C1352 PAD.n467 VSS 0.036454f
C1353 PAD.n468 VSS 0.036454f
C1354 PAD.n470 VSS 0.036454f
C1355 PAD.n471 VSS 0.036454f
C1356 PAD.n472 VSS 0.036454f
C1357 PAD.n474 VSS 0.036454f
C1358 PAD.n475 VSS 0.036454f
C1359 PAD.n476 VSS 0.036454f
C1360 PAD.n478 VSS 0.036454f
C1361 PAD.n479 VSS 0.036454f
C1362 PAD.n480 VSS 0.036454f
C1363 PAD.n482 VSS 0.036454f
C1364 PAD.n483 VSS 0.036454f
C1365 PAD.n484 VSS 0.036454f
C1366 PAD.n486 VSS 0.036454f
C1367 PAD.n487 VSS 0.036454f
C1368 PAD.n488 VSS 0.036454f
C1369 PAD.n490 VSS 0.036454f
C1370 PAD.n491 VSS 0.036454f
C1371 PAD.n492 VSS 0.036454f
C1372 PAD.n494 VSS 0.036454f
C1373 PAD.n495 VSS 0.036454f
C1374 PAD.n496 VSS 0.036454f
C1375 PAD.n498 VSS 0.036454f
C1376 PAD.n499 VSS 0.036454f
C1377 PAD.n500 VSS 0.036454f
C1378 PAD.n502 VSS 0.036454f
C1379 PAD.n503 VSS 0.036454f
C1380 PAD.n504 VSS 0.036454f
C1381 PAD.n506 VSS 0.036454f
C1382 PAD.n507 VSS 0.036454f
C1383 PAD.n508 VSS 0.036454f
C1384 PAD.n510 VSS 0.036454f
C1385 PAD.n511 VSS 0.036454f
C1386 PAD.n512 VSS 0.036454f
C1387 PAD.n514 VSS 0.036454f
C1388 PAD.n515 VSS 0.036454f
C1389 PAD.n516 VSS 0.036454f
C1390 PAD.n518 VSS 0.036454f
C1391 PAD.n519 VSS 0.036454f
C1392 PAD.n520 VSS 0.036454f
C1393 PAD.n521 VSS 0.033374f
C1394 PAD.n522 VSS 0.023105f
C1395 PAD.n523 VSS 0.023105f
C1396 PAD.n525 VSS 0.036454f
C1397 PAD.n527 VSS 0.036454f
C1398 PAD.n529 VSS 0.036454f
C1399 PAD.n530 VSS 0.036454f
C1400 PAD.n531 VSS 0.036454f
C1401 PAD.n532 VSS 0.036454f
C1402 PAD.n533 VSS 0.036454f
C1403 PAD.n534 VSS 0.036454f
C1404 PAD.n535 VSS 0.036454f
C1405 PAD.n537 VSS 0.036454f
C1406 PAD.n539 VSS 0.036454f
C1407 PAD.n541 VSS 0.036454f
C1408 PAD.n542 VSS 0.036454f
C1409 PAD.n543 VSS 0.036454f
C1410 PAD.n544 VSS 0.036454f
C1411 PAD.n545 VSS 0.036454f
C1412 PAD.n546 VSS 0.036454f
C1413 PAD.n547 VSS 0.036454f
C1414 PAD.n549 VSS 0.036454f
C1415 PAD.n551 VSS 0.036454f
C1416 PAD.n553 VSS 0.036454f
C1417 PAD.n554 VSS 0.036454f
C1418 PAD.n555 VSS 0.036454f
C1419 PAD.n556 VSS 0.036454f
C1420 PAD.n557 VSS 0.036454f
C1421 PAD.n558 VSS 0.036454f
C1422 PAD.n559 VSS 0.036454f
C1423 PAD.n561 VSS 0.036454f
C1424 PAD.n563 VSS 0.036454f
C1425 PAD.n565 VSS 0.036454f
C1426 PAD.n566 VSS 0.036454f
C1427 PAD.n567 VSS 0.036454f
C1428 PAD.n568 VSS 0.036454f
C1429 PAD.n569 VSS 0.036454f
C1430 PAD.n570 VSS 0.036454f
C1431 PAD.n571 VSS 0.036454f
C1432 PAD.n573 VSS 0.036454f
C1433 PAD.n575 VSS 0.036454f
C1434 PAD.n577 VSS 0.036454f
C1435 PAD.n578 VSS 0.036454f
C1436 PAD.n579 VSS 0.036454f
C1437 PAD.n580 VSS 0.036454f
C1438 PAD.n581 VSS 0.036454f
C1439 PAD.n582 VSS 0.036454f
C1440 PAD.n583 VSS 0.036454f
C1441 PAD.n585 VSS 0.036454f
C1442 PAD.n587 VSS 0.036454f
C1443 PAD.n589 VSS 0.036454f
C1444 PAD.n590 VSS 0.036454f
C1445 PAD.n591 VSS 0.036454f
C1446 PAD.n592 VSS 0.036454f
C1447 PAD.n593 VSS 0.036454f
C1448 PAD.n594 VSS 0.036454f
C1449 PAD.n595 VSS 0.036454f
C1450 PAD.n597 VSS 0.036454f
C1451 PAD.n599 VSS 0.036454f
C1452 PAD.n601 VSS 0.036454f
C1453 PAD.n602 VSS 0.036454f
C1454 PAD.n603 VSS 0.036454f
C1455 PAD.n604 VSS 0.036454f
C1456 PAD.n605 VSS 0.036454f
C1457 PAD.n606 VSS 0.036454f
C1458 PAD.n607 VSS 0.036454f
C1459 PAD.n609 VSS 0.036454f
C1460 PAD.n611 VSS 0.036454f
C1461 PAD.n613 VSS 0.036454f
C1462 PAD.n614 VSS 0.036454f
C1463 PAD.n615 VSS 0.036454f
C1464 PAD.n616 VSS 0.036454f
C1465 PAD.n617 VSS 0.036454f
C1466 PAD.n618 VSS 0.036454f
C1467 PAD.n619 VSS 0.036454f
C1468 PAD.n621 VSS 0.036454f
C1469 PAD.n623 VSS 0.036454f
C1470 PAD.n625 VSS 0.036454f
C1471 PAD.n626 VSS 0.036454f
C1472 PAD.n627 VSS 0.036454f
C1473 PAD.n628 VSS 0.036454f
C1474 PAD.n629 VSS 0.036454f
C1475 PAD.n630 VSS 0.036454f
C1476 PAD.n631 VSS 0.036454f
C1477 PAD.n633 VSS 0.036454f
C1478 PAD.n635 VSS 0.036454f
C1479 PAD.n637 VSS 0.036454f
C1480 PAD.n638 VSS 0.036454f
C1481 PAD.n639 VSS 0.036454f
C1482 PAD.n640 VSS 0.036454f
C1483 PAD.n641 VSS 0.036454f
C1484 PAD.n642 VSS 0.036454f
C1485 PAD.n643 VSS 0.036454f
C1486 PAD.n645 VSS 0.036454f
C1487 PAD.n647 VSS 0.036454f
C1488 PAD.n649 VSS 0.036454f
C1489 PAD.n650 VSS 0.036454f
C1490 PAD.n651 VSS 0.036454f
C1491 PAD.n652 VSS 0.036454f
C1492 PAD.n653 VSS 0.036454f
C1493 PAD.n654 VSS 0.036454f
C1494 PAD.n655 VSS 0.036454f
C1495 PAD.n657 VSS 0.036454f
C1496 PAD.n659 VSS 0.036454f
C1497 PAD.n661 VSS 0.036454f
C1498 PAD.n662 VSS 0.036454f
C1499 PAD.n663 VSS 0.036454f
C1500 PAD.n664 VSS 0.036454f
C1501 PAD.n665 VSS 0.036454f
C1502 PAD.n666 VSS 0.036454f
C1503 PAD.n667 VSS 0.036454f
C1504 PAD.n669 VSS 0.036454f
C1505 PAD.n671 VSS 0.036454f
C1506 PAD.n673 VSS 0.036454f
C1507 PAD.n674 VSS 0.036454f
C1508 PAD.n675 VSS 0.036454f
C1509 PAD.n676 VSS 0.036454f
C1510 PAD.n677 VSS 0.036454f
C1511 PAD.n678 VSS 0.036454f
C1512 PAD.n679 VSS 0.036454f
C1513 PAD.n681 VSS 0.036454f
C1514 PAD.n683 VSS 0.036454f
C1515 PAD.n685 VSS 0.036454f
C1516 PAD.n686 VSS 0.036454f
C1517 PAD.n687 VSS 0.036454f
C1518 PAD.n688 VSS 0.036454f
C1519 PAD.n689 VSS 0.036454f
C1520 PAD.n690 VSS 0.036454f
C1521 PAD.n691 VSS 0.036454f
C1522 PAD.n693 VSS 0.036454f
C1523 PAD.n695 VSS 0.036454f
C1524 PAD.n697 VSS 0.036454f
C1525 PAD.n698 VSS 0.036454f
C1526 PAD.n699 VSS 0.036454f
C1527 PAD.n700 VSS 0.036454f
C1528 PAD.n701 VSS 0.036454f
C1529 PAD.n702 VSS 0.036454f
C1530 PAD.n703 VSS 0.036454f
C1531 PAD.n705 VSS 0.036454f
C1532 PAD.n707 VSS 0.036454f
C1533 PAD.n709 VSS 0.036454f
C1534 PAD.n710 VSS 0.036454f
C1535 PAD.n711 VSS 0.036454f
C1536 PAD.n712 VSS 0.036454f
C1537 PAD.n713 VSS 0.036454f
C1538 PAD.n714 VSS 0.036454f
C1539 PAD.n715 VSS 0.036454f
C1540 PAD.n717 VSS 0.036454f
C1541 PAD.n719 VSS 0.036454f
C1542 PAD.n721 VSS 0.036454f
C1543 PAD.n722 VSS 0.036454f
C1544 PAD.n723 VSS 0.036454f
C1545 PAD.n724 VSS 0.036454f
C1546 PAD.n725 VSS 0.036454f
C1547 PAD.n726 VSS 0.036454f
C1548 PAD.n727 VSS 0.036454f
C1549 PAD.n729 VSS 0.036454f
C1550 PAD.n731 VSS 0.036454f
C1551 PAD.n733 VSS 0.036454f
C1552 PAD.n734 VSS 0.036454f
C1553 PAD.n735 VSS 0.036454f
C1554 PAD.n736 VSS 0.036454f
C1555 PAD.n737 VSS 0.036454f
C1556 PAD.n738 VSS 0.036454f
C1557 PAD.n739 VSS 0.036454f
C1558 PAD.n741 VSS 0.036454f
C1559 PAD.n743 VSS 0.036454f
C1560 PAD.n745 VSS 0.036454f
C1561 PAD.n746 VSS 0.036454f
C1562 PAD.n747 VSS 0.036454f
C1563 PAD.n748 VSS 0.036454f
C1564 PAD.n749 VSS 0.036454f
C1565 PAD.n750 VSS 0.036454f
C1566 PAD.n751 VSS 0.036454f
C1567 PAD.n753 VSS 0.036454f
C1568 PAD.n755 VSS 0.036454f
C1569 PAD.n757 VSS 0.036454f
C1570 PAD.n758 VSS 0.036454f
C1571 PAD.n759 VSS 0.036454f
C1572 PAD.n760 VSS 0.036454f
C1573 PAD.n761 VSS 0.036454f
C1574 PAD.n762 VSS 0.036454f
C1575 PAD.n763 VSS 0.036454f
C1576 PAD.n764 VSS 0.036454f
C1577 PAD.n766 VSS 0.036454f
C1578 PAD.n768 VSS 0.036454f
C1579 PAD.n770 VSS 0.023105f
C1580 PAD.n771 VSS 0.023105f
C1581 PAD.n772 VSS 0.03055f
C1582 PAD.n773 VSS 0.042887f
C1583 PAD.n774 VSS 0.049106f
C1584 PAD.n775 VSS 0.049106f
C1585 PAD.n776 VSS 0.700403f
C1586 PAD.n777 VSS 0.069752f
C1587 PAD.n778 VSS 0.069752f
C1588 PAD.n779 VSS 0.046278f
C1589 PAD.n780 VSS 0.039754f
C1590 PAD.n781 VSS 0.039754f
C1591 PAD.n782 VSS 0.611619f
C1592 PAD.n824 VSS 0.023105f
C1593 PAD.n825 VSS 0.542565f
C1594 PAD.n826 VSS 0.023105f
C1595 PAD.n827 VSS 0.029431f
C1596 PAD.n828 VSS 0.350201f
C1597 PAD.n829 VSS 0.036454f
C1598 PAD.n830 VSS 0.036454f
C1599 PAD.n831 VSS 0.036454f
C1600 PAD.n832 VSS 0.036454f
C1601 PAD.n833 VSS 0.036454f
C1602 PAD.n834 VSS 0.036454f
C1603 PAD.n835 VSS 0.036454f
C1604 PAD.n836 VSS 0.036454f
C1605 PAD.n837 VSS 0.036454f
C1606 PAD.n838 VSS 0.036454f
C1607 PAD.n839 VSS 0.036454f
C1608 PAD.n840 VSS 0.036454f
C1609 PAD.n841 VSS 0.036454f
C1610 PAD.n842 VSS 0.036454f
C1611 PAD.n843 VSS 0.036454f
C1612 PAD.n844 VSS 0.036454f
C1613 PAD.n845 VSS 0.036454f
C1614 PAD.n846 VSS 0.036454f
C1615 PAD.n847 VSS 0.036454f
C1616 PAD.n848 VSS 0.036454f
C1617 PAD.n849 VSS 0.036454f
C1618 PAD.n850 VSS 0.036454f
C1619 PAD.n851 VSS 0.036454f
C1620 PAD.n852 VSS 0.036454f
C1621 PAD.n853 VSS 0.036454f
C1622 PAD.n854 VSS 0.036454f
C1623 PAD.n855 VSS 0.036454f
C1624 PAD.n856 VSS 0.036454f
C1625 PAD.n857 VSS 0.036454f
C1626 PAD.n858 VSS 0.036454f
C1627 PAD.n859 VSS 0.036454f
C1628 PAD.n860 VSS 0.036454f
C1629 PAD.n861 VSS 0.036454f
C1630 PAD.n862 VSS 0.036454f
C1631 PAD.n863 VSS 0.036454f
C1632 PAD.n864 VSS 0.036454f
C1633 PAD.n865 VSS 0.036454f
C1634 PAD.n866 VSS 0.036454f
C1635 PAD.n867 VSS 0.036454f
C1636 PAD.n868 VSS 0.036454f
C1637 PAD.n870 VSS 0.036454f
C1638 PAD.n871 VSS 0.036454f
C1639 PAD.n872 VSS 0.023105f
C1640 PAD.n873 VSS 0.033374f
C1641 PAD.n874 VSS 0.036454f
C1642 PAD.n875 VSS 0.036454f
C1643 PAD.n876 VSS 0.036454f
C1644 PAD.n877 VSS 0.036454f
C1645 PAD.n879 VSS 0.036454f
C1646 PAD.n880 VSS 0.036454f
C1647 PAD.n881 VSS 0.036454f
C1648 PAD.n883 VSS 0.036454f
C1649 PAD.n884 VSS 0.036454f
C1650 PAD.n885 VSS 0.036454f
C1651 PAD.n886 VSS 0.036454f
C1652 PAD.n887 VSS 0.036454f
C1653 PAD.n888 VSS 0.036454f
C1654 PAD.n889 VSS 0.036454f
C1655 PAD.n891 VSS 0.036454f
C1656 PAD.n892 VSS 0.036454f
C1657 PAD.n893 VSS 0.036454f
C1658 PAD.n895 VSS 0.036454f
C1659 PAD.n896 VSS 0.036454f
C1660 PAD.n897 VSS 0.036454f
C1661 PAD.n898 VSS 0.036454f
C1662 PAD.n899 VSS 0.036454f
C1663 PAD.n900 VSS 0.036454f
C1664 PAD.n901 VSS 0.036454f
C1665 PAD.n903 VSS 0.036454f
C1666 PAD.n904 VSS 0.036454f
C1667 PAD.n905 VSS 0.036454f
C1668 PAD.n907 VSS 0.036454f
C1669 PAD.n908 VSS 0.036454f
C1670 PAD.n909 VSS 0.036454f
C1671 PAD.n910 VSS 0.036454f
C1672 PAD.n911 VSS 0.036454f
C1673 PAD.n912 VSS 0.036454f
C1674 PAD.n913 VSS 0.036454f
C1675 PAD.n915 VSS 0.036454f
C1676 PAD.n916 VSS 0.036454f
C1677 PAD.n917 VSS 0.036454f
C1678 PAD.n919 VSS 0.036454f
C1679 PAD.n920 VSS 0.036454f
C1680 PAD.n921 VSS 0.036454f
C1681 PAD.n922 VSS 0.036454f
C1682 PAD.n923 VSS 0.036454f
C1683 PAD.n924 VSS 0.036454f
C1684 PAD.n925 VSS 0.036454f
C1685 PAD.n927 VSS 0.036454f
C1686 PAD.n928 VSS 0.036454f
C1687 PAD.n929 VSS 0.036454f
C1688 PAD.n931 VSS 0.036454f
C1689 PAD.n932 VSS 0.036454f
C1690 PAD.n933 VSS 0.036454f
C1691 PAD.n934 VSS 0.036454f
C1692 PAD.n935 VSS 0.036454f
C1693 PAD.n936 VSS 0.036454f
C1694 PAD.n937 VSS 0.036454f
C1695 PAD.n939 VSS 0.036454f
C1696 PAD.n940 VSS 0.036454f
C1697 PAD.n941 VSS 0.036454f
C1698 PAD.n943 VSS 0.036454f
C1699 PAD.n944 VSS 0.036454f
C1700 PAD.n945 VSS 0.036454f
C1701 PAD.n946 VSS 0.036454f
C1702 PAD.n947 VSS 0.036454f
C1703 PAD.n948 VSS 0.036454f
C1704 PAD.n949 VSS 0.036454f
C1705 PAD.n951 VSS 0.036454f
C1706 PAD.n952 VSS 0.036454f
C1707 PAD.n953 VSS 0.036454f
C1708 PAD.n955 VSS 0.036454f
C1709 PAD.n956 VSS 0.036454f
C1710 PAD.n957 VSS 0.036454f
C1711 PAD.n958 VSS 0.036454f
C1712 PAD.n959 VSS 0.036454f
C1713 PAD.n960 VSS 0.036454f
C1714 PAD.n961 VSS 0.036454f
C1715 PAD.n963 VSS 0.036454f
C1716 PAD.n964 VSS 0.036454f
C1717 PAD.n965 VSS 0.036454f
C1718 PAD.n967 VSS 0.036454f
C1719 PAD.n968 VSS 0.036454f
C1720 PAD.n969 VSS 0.036454f
C1721 PAD.n970 VSS 0.036454f
C1722 PAD.n971 VSS 0.036454f
C1723 PAD.n972 VSS 0.036454f
C1724 PAD.n973 VSS 0.036454f
C1725 PAD.n975 VSS 0.036454f
C1726 PAD.n976 VSS 0.036454f
C1727 PAD.n977 VSS 0.036454f
C1728 PAD.n979 VSS 0.036454f
C1729 PAD.n980 VSS 0.036454f
C1730 PAD.n981 VSS 0.036454f
C1731 PAD.n982 VSS 0.036454f
C1732 PAD.n983 VSS 0.036454f
C1733 PAD.n984 VSS 0.036454f
C1734 PAD.n985 VSS 0.036454f
C1735 PAD.n987 VSS 0.036454f
C1736 PAD.n988 VSS 0.036454f
C1737 PAD.n989 VSS 0.036454f
C1738 PAD.n991 VSS 0.036454f
C1739 PAD.n992 VSS 0.036454f
C1740 PAD.n993 VSS 0.036454f
C1741 PAD.n994 VSS 0.036454f
C1742 PAD.n995 VSS 0.036454f
C1743 PAD.n996 VSS 0.036454f
C1744 PAD.n997 VSS 0.036454f
C1745 PAD.n999 VSS 0.036454f
C1746 PAD.n1000 VSS 0.036454f
C1747 PAD.n1001 VSS 0.036454f
C1748 PAD.n1003 VSS 0.036454f
C1749 PAD.n1004 VSS 0.036454f
C1750 PAD.n1005 VSS 0.036454f
C1751 PAD.n1006 VSS 0.036454f
C1752 PAD.n1007 VSS 0.036454f
C1753 PAD.n1008 VSS 0.036454f
C1754 PAD.n1009 VSS 0.036454f
C1755 PAD.n1011 VSS 0.036454f
C1756 PAD.n1012 VSS 0.036454f
C1757 PAD.n1013 VSS 0.036454f
C1758 PAD.n1015 VSS 0.036454f
C1759 PAD.n1016 VSS 0.036454f
C1760 PAD.n1017 VSS 0.036454f
C1761 PAD.n1018 VSS 0.036454f
C1762 PAD.n1019 VSS 0.036454f
C1763 PAD.n1020 VSS 0.036454f
C1764 PAD.n1021 VSS 0.036454f
C1765 PAD.n1023 VSS 0.036454f
C1766 PAD.n1024 VSS 0.036454f
C1767 PAD.n1025 VSS 0.036454f
C1768 PAD.n1027 VSS 0.036454f
C1769 PAD.n1028 VSS 0.036454f
C1770 PAD.n1029 VSS 0.036454f
C1771 PAD.n1030 VSS 0.036454f
C1772 PAD.n1031 VSS 0.036454f
C1773 PAD.n1032 VSS 0.036454f
C1774 PAD.n1033 VSS 0.036454f
C1775 PAD.n1035 VSS 0.036454f
C1776 PAD.n1036 VSS 0.036454f
C1777 PAD.n1037 VSS 0.036454f
C1778 PAD.n1039 VSS 0.036454f
C1779 PAD.n1040 VSS 0.036454f
C1780 PAD.n1041 VSS 0.036454f
C1781 PAD.n1042 VSS 0.036454f
C1782 PAD.n1043 VSS 0.036454f
C1783 PAD.n1044 VSS 0.036454f
C1784 PAD.n1045 VSS 0.036454f
C1785 PAD.n1047 VSS 0.036454f
C1786 PAD.n1048 VSS 0.036454f
C1787 PAD.n1049 VSS 0.036454f
C1788 PAD.n1051 VSS 0.036454f
C1789 PAD.n1052 VSS 0.036454f
C1790 PAD.n1053 VSS 0.036454f
C1791 PAD.n1054 VSS 0.036454f
C1792 PAD.n1055 VSS 0.036454f
C1793 PAD.n1056 VSS 0.036454f
C1794 PAD.n1057 VSS 0.036454f
C1795 PAD.n1059 VSS 0.036454f
C1796 PAD.n1060 VSS 0.036454f
C1797 PAD.n1061 VSS 0.036454f
C1798 PAD.n1063 VSS 0.036454f
C1799 PAD.n1064 VSS 0.036454f
C1800 PAD.n1065 VSS 0.036454f
C1801 PAD.n1066 VSS 0.036454f
C1802 PAD.n1067 VSS 0.036454f
C1803 PAD.n1068 VSS 0.036454f
C1804 PAD.n1069 VSS 0.036454f
C1805 PAD.n1071 VSS 0.036454f
C1806 PAD.n1072 VSS 0.036454f
C1807 PAD.n1073 VSS 0.036454f
C1808 PAD.n1075 VSS 0.036454f
C1809 PAD.n1076 VSS 0.036454f
C1810 PAD.n1077 VSS 0.036454f
C1811 PAD.n1078 VSS 0.036454f
C1812 PAD.n1079 VSS 0.036454f
C1813 PAD.n1080 VSS 0.036454f
C1814 PAD.n1081 VSS 0.036454f
C1815 PAD.n1083 VSS 0.036454f
C1816 PAD.n1084 VSS 0.036454f
C1817 PAD.n1085 VSS 0.036454f
C1818 PAD.n1087 VSS 0.036454f
C1819 PAD.n1088 VSS 0.036454f
C1820 PAD.n1089 VSS 0.036454f
C1821 PAD.n1090 VSS 0.036454f
C1822 PAD.n1091 VSS 0.036454f
C1823 PAD.n1092 VSS 0.036454f
C1824 PAD.n1093 VSS 0.036454f
C1825 PAD.n1095 VSS 0.036454f
C1826 PAD.n1096 VSS 0.036454f
C1827 PAD.n1097 VSS 0.036454f
C1828 PAD.n1099 VSS 0.036454f
C1829 PAD.n1100 VSS 0.036454f
C1830 PAD.n1101 VSS 0.036454f
C1831 PAD.n1102 VSS 0.036454f
C1832 PAD.n1103 VSS 0.036454f
C1833 PAD.n1104 VSS 0.036454f
C1834 PAD.n1105 VSS 0.036454f
C1835 PAD.n1107 VSS 0.036454f
C1836 PAD.n1108 VSS 0.036454f
C1837 PAD.n1109 VSS 0.036454f
C1838 PAD.n1111 VSS 0.036454f
C1839 PAD.n1112 VSS 0.036454f
C1840 PAD.n1113 VSS 0.036454f
C1841 PAD.n1114 VSS 0.036454f
C1842 PAD.n1115 VSS 0.04183f
C1843 PAD.n1116 VSS 0.045821f
C1844 PAD.n1117 VSS 0.045821f
C1845 PAD.n1118 VSS 0.611619f
C1846 PAD.n1119 VSS 0.059627f
C1847 PAD.n1120 VSS 0.369931f
C1848 PAD.n1121 VSS 0.052877f
C1849 PAD.n1122 VSS 0.059627f
C1850 PAD.n1123 VSS 0.052877f
C1851 PAD.n1124 VSS 0.033374f
C1852 PAD.n1125 VSS 0.062262f
C1853 PAD.n1126 VSS 0.069752f
C1854 PAD.n1127 VSS 0.039754f
C1855 PAD.n1128 VSS 0.069752f
C1856 PAD.n1129 VSS 0.039754f
C1857 PAD.n1130 VSS 0.61162f
C1858 PAD.n1131 VSS 0.261418f
C1859 PAD.n1132 VSS 0.527768f
C1860 PAD.n1133 VSS 0.049106f
C1861 PAD.n1134 VSS 0.029431f
C1862 PAD.n1135 VSS 0.049106f
C1863 PAD.n1136 VSS 0.029431f
C1864 PAD.n1137 VSS 0.033766f
C1865 PAD.n1138 VSS 0.029431f
C1866 PAD.n1139 VSS 0.029431f
C1867 PAD.n1140 VSS 0.517904f
C1868 PAD.n1141 VSS 0.438985f
C1869 PAD.n1142 VSS 0.611619f
C1870 PAD.n1143 VSS 0.039754f
C1871 PAD.n1144 VSS 0.039754f
C1872 PAD.n1145 VSS 0.033374f
C1873 PAD.n1146 VSS 0.062262f
C1874 PAD.n1147 VSS 0.069752f
C1875 PAD.n1148 VSS 0.069752f
C1876 PAD.n1190 VSS 0.036454f
C1877 PAD.n1192 VSS 0.036454f
C1878 PAD.n1193 VSS 0.036454f
C1879 PAD.n1194 VSS 0.036454f
C1880 PAD.n1195 VSS 0.036454f
C1881 PAD.n1196 VSS 0.036454f
C1882 PAD.n1198 VSS 0.036454f
C1883 PAD.n1199 VSS 0.036454f
C1884 PAD.n1200 VSS 0.036454f
C1885 PAD.n1201 VSS 0.036454f
C1886 PAD.n1203 VSS 0.036454f
C1887 PAD.n1204 VSS 0.036454f
C1888 PAD.n1205 VSS 0.036454f
C1889 PAD.n1206 VSS 0.036454f
C1890 PAD.n1208 VSS 0.036454f
C1891 PAD.n1209 VSS 0.036454f
C1892 PAD.n1210 VSS 0.036454f
C1893 PAD.n1211 VSS 0.036454f
C1894 PAD.n1213 VSS 0.036454f
C1895 PAD.n1214 VSS 0.036454f
C1896 PAD.n1215 VSS 0.036454f
C1897 PAD.n1216 VSS 0.036454f
C1898 PAD.n1218 VSS 0.036454f
C1899 PAD.n1219 VSS 0.036454f
C1900 PAD.n1220 VSS 0.036454f
C1901 PAD.n1221 VSS 0.036454f
C1902 PAD.n1223 VSS 0.036454f
C1903 PAD.n1224 VSS 0.036454f
C1904 PAD.n1225 VSS 0.036454f
C1905 PAD.n1226 VSS 0.036454f
C1906 PAD.n1228 VSS 0.036454f
C1907 PAD.n1229 VSS 0.036454f
C1908 PAD.n1230 VSS 0.036454f
C1909 PAD.n1231 VSS 0.036454f
C1910 PAD.n1233 VSS 0.036454f
C1911 PAD.n1234 VSS 0.036454f
C1912 PAD.n1235 VSS 0.036454f
C1913 PAD.n1236 VSS 0.036454f
C1914 PAD.n1238 VSS 0.036454f
C1915 PAD.n1239 VSS 0.036454f
C1916 PAD.n1240 VSS 0.036454f
C1917 PAD.n1241 VSS 0.036454f
C1918 PAD.n1243 VSS 0.036454f
C1919 PAD.n1244 VSS 0.036454f
C1920 PAD.n1245 VSS 0.036454f
C1921 PAD.n1246 VSS 0.036454f
C1922 PAD.n1248 VSS 0.036454f
C1923 PAD.n1249 VSS 0.036454f
C1924 PAD.n1250 VSS 0.036454f
C1925 PAD.n1251 VSS 0.036454f
C1926 PAD.n1253 VSS 0.036454f
C1927 PAD.n1254 VSS 0.036454f
C1928 PAD.n1255 VSS 0.036454f
C1929 PAD.n1256 VSS 0.036454f
C1930 PAD.n1258 VSS 0.036454f
C1931 PAD.n1259 VSS 0.036454f
C1932 PAD.n1260 VSS 0.036454f
C1933 PAD.n1261 VSS 0.036454f
C1934 PAD.n1263 VSS 0.036454f
C1935 PAD.n1264 VSS 0.036454f
C1936 PAD.n1265 VSS 0.036454f
C1937 PAD.n1266 VSS 0.036454f
C1938 PAD.n1268 VSS 0.036454f
C1939 PAD.n1269 VSS 0.036454f
C1940 PAD.n1270 VSS 0.036454f
C1941 PAD.n1271 VSS 0.036454f
C1942 PAD.n1273 VSS 0.036454f
C1943 PAD.n1274 VSS 0.036454f
C1944 PAD.n1275 VSS 0.036454f
C1945 PAD.n1276 VSS 0.036454f
C1946 PAD.n1278 VSS 0.036454f
C1947 PAD.n1279 VSS 0.036454f
C1948 PAD.n1280 VSS 0.036454f
C1949 PAD.n1281 VSS 0.036454f
C1950 PAD.n1283 VSS 0.036454f
C1951 PAD.n1284 VSS 0.036454f
C1952 PAD.n1285 VSS 0.036454f
C1953 PAD.n1286 VSS 0.036454f
C1954 PAD.n1288 VSS 0.036454f
C1955 PAD.n1289 VSS 0.036454f
C1956 PAD.n1290 VSS 0.036454f
C1957 PAD.n1291 VSS 0.036454f
C1958 PAD.n1293 VSS 0.036454f
C1959 PAD.n1294 VSS 0.023105f
C1960 PAD.n1295 VSS 0.023105f
C1961 PAD.n1296 VSS 0.03055f
C1962 PAD.n1297 VSS 0.036454f
C1963 PAD.n1298 VSS 0.036454f
C1964 PAD.n1299 VSS 0.036454f
C1965 PAD.n1300 VSS 0.036454f
C1966 PAD.n1301 VSS 0.036454f
C1967 PAD.n1303 VSS 0.036454f
C1968 PAD.n1304 VSS 0.036454f
C1969 PAD.n1305 VSS 0.036454f
C1970 PAD.n1306 VSS 0.036454f
C1971 PAD.n1307 VSS 0.036454f
C1972 PAD.n1308 VSS 0.036454f
C1973 PAD.n1309 VSS 0.036454f
C1974 PAD.n1310 VSS 0.036454f
C1975 PAD.n1312 VSS 0.036454f
C1976 PAD.n1313 VSS 0.036454f
C1977 PAD.n1314 VSS 0.036454f
C1978 PAD.n1315 VSS 0.036454f
C1979 PAD.n1316 VSS 0.036454f
C1980 PAD.n1317 VSS 0.036454f
C1981 PAD.n1318 VSS 0.036454f
C1982 PAD.n1319 VSS 0.036454f
C1983 PAD.n1321 VSS 0.036454f
C1984 PAD.n1322 VSS 0.036454f
C1985 PAD.n1323 VSS 0.036454f
C1986 PAD.n1324 VSS 0.036454f
C1987 PAD.n1325 VSS 0.036454f
C1988 PAD.n1326 VSS 0.036454f
C1989 PAD.n1327 VSS 0.036454f
C1990 PAD.n1328 VSS 0.036454f
C1991 PAD.n1330 VSS 0.036454f
C1992 PAD.n1331 VSS 0.036454f
C1993 PAD.n1332 VSS 0.036454f
C1994 PAD.n1333 VSS 0.036454f
C1995 PAD.n1334 VSS 0.036454f
C1996 PAD.n1335 VSS 0.036454f
C1997 PAD.n1336 VSS 0.036454f
C1998 PAD.n1337 VSS 0.036454f
C1999 PAD.n1339 VSS 0.036454f
C2000 PAD.n1340 VSS 0.036454f
C2001 PAD.n1341 VSS 0.036454f
C2002 PAD.n1342 VSS 0.036454f
C2003 PAD.n1343 VSS 0.036454f
C2004 PAD.n1344 VSS 0.036454f
C2005 PAD.n1345 VSS 0.036454f
C2006 PAD.n1346 VSS 0.036454f
C2007 PAD.n1348 VSS 0.036454f
C2008 PAD.n1349 VSS 0.036454f
C2009 PAD.n1350 VSS 0.036454f
C2010 PAD.n1351 VSS 0.036454f
C2011 PAD.n1352 VSS 0.036454f
C2012 PAD.n1353 VSS 0.036454f
C2013 PAD.n1354 VSS 0.036454f
C2014 PAD.n1355 VSS 0.036454f
C2015 PAD.n1357 VSS 0.036454f
C2016 PAD.n1358 VSS 0.036454f
C2017 PAD.n1359 VSS 0.036454f
C2018 PAD.n1360 VSS 0.036454f
C2019 PAD.n1361 VSS 0.036454f
C2020 PAD.n1362 VSS 0.036454f
C2021 PAD.n1363 VSS 0.036454f
C2022 PAD.n1364 VSS 0.036454f
C2023 PAD.n1366 VSS 0.036454f
C2024 PAD.n1367 VSS 0.036454f
C2025 PAD.n1368 VSS 0.036454f
C2026 PAD.n1369 VSS 0.036454f
C2027 PAD.n1370 VSS 0.036454f
C2028 PAD.n1371 VSS 0.036454f
C2029 PAD.n1372 VSS 0.036454f
C2030 PAD.n1373 VSS 0.036454f
C2031 PAD.n1375 VSS 0.036454f
C2032 PAD.n1376 VSS 0.036454f
C2033 PAD.n1377 VSS 0.036454f
C2034 PAD.n1378 VSS 0.036454f
C2035 PAD.n1379 VSS 0.036454f
C2036 PAD.n1380 VSS 0.036454f
C2037 PAD.n1381 VSS 0.036454f
C2038 PAD.n1382 VSS 0.036454f
C2039 PAD.n1384 VSS 0.036454f
C2040 PAD.n1385 VSS 0.036454f
C2041 PAD.n1386 VSS 0.036454f
C2042 PAD.n1387 VSS 0.036454f
C2043 PAD.n1388 VSS 0.036454f
C2044 PAD.n1389 VSS 0.036454f
C2045 PAD.n1390 VSS 0.036454f
C2046 PAD.n1391 VSS 0.036454f
C2047 PAD.n1393 VSS 0.036454f
C2048 PAD.n1394 VSS 0.036454f
C2049 PAD.n1395 VSS 0.036454f
C2050 PAD.n1396 VSS 0.036454f
C2051 PAD.n1397 VSS 0.036454f
C2052 PAD.n1398 VSS 0.036454f
C2053 PAD.n1399 VSS 0.036454f
C2054 PAD.n1400 VSS 0.036454f
C2055 PAD.n1402 VSS 0.036454f
C2056 PAD.n1403 VSS 0.036454f
C2057 PAD.n1404 VSS 0.036454f
C2058 PAD.n1405 VSS 0.036454f
C2059 PAD.n1406 VSS 0.036454f
C2060 PAD.n1407 VSS 0.036454f
C2061 PAD.n1408 VSS 0.036454f
C2062 PAD.n1409 VSS 0.036454f
C2063 PAD.n1411 VSS 0.036454f
C2064 PAD.n1412 VSS 0.036454f
C2065 PAD.n1413 VSS 0.036454f
C2066 PAD.n1414 VSS 0.036454f
C2067 PAD.n1415 VSS 0.036454f
C2068 PAD.n1416 VSS 0.036454f
C2069 PAD.n1417 VSS 0.036454f
C2070 PAD.n1418 VSS 0.036454f
C2071 PAD.n1420 VSS 0.036454f
C2072 PAD.n1421 VSS 0.036454f
C2073 PAD.n1422 VSS 0.036454f
C2074 PAD.n1423 VSS 0.036454f
C2075 PAD.n1424 VSS 0.036454f
C2076 PAD.n1425 VSS 0.036454f
C2077 PAD.n1426 VSS 0.036454f
C2078 PAD.n1427 VSS 0.036454f
C2079 PAD.n1429 VSS 0.036454f
C2080 PAD.n1430 VSS 0.036454f
C2081 PAD.n1431 VSS 0.036454f
C2082 PAD.n1432 VSS 0.036454f
C2083 PAD.n1433 VSS 0.036454f
C2084 PAD.n1434 VSS 0.036454f
C2085 PAD.n1435 VSS 0.036454f
C2086 PAD.n1436 VSS 0.036454f
C2087 PAD.n1438 VSS 0.036454f
C2088 PAD.n1439 VSS 0.036454f
C2089 PAD.n1440 VSS 0.036454f
C2090 PAD.n1441 VSS 0.036454f
C2091 PAD.n1442 VSS 0.036454f
C2092 PAD.n1443 VSS 0.036454f
C2093 PAD.n1444 VSS 0.036454f
C2094 PAD.n1445 VSS 0.036454f
C2095 PAD.n1447 VSS 0.036454f
C2096 PAD.n1448 VSS 0.036454f
C2097 PAD.n1449 VSS 0.036454f
C2098 PAD.n1450 VSS 0.036454f
C2099 PAD.n1451 VSS 0.036454f
C2100 PAD.n1452 VSS 0.036454f
C2101 PAD.n1453 VSS 0.036454f
C2102 PAD.n1454 VSS 0.036454f
C2103 PAD.n1456 VSS 0.036454f
C2104 PAD.n1457 VSS 0.036454f
C2105 PAD.n1458 VSS 0.036454f
C2106 PAD.n1459 VSS 0.036454f
C2107 PAD.n1460 VSS 0.036454f
C2108 PAD.n1461 VSS 0.036454f
C2109 PAD.n1462 VSS 0.036454f
C2110 PAD.n1463 VSS 0.036454f
C2111 PAD.n1465 VSS 0.036454f
C2112 PAD.n1466 VSS 0.036454f
C2113 PAD.n1467 VSS 0.036454f
C2114 PAD.n1468 VSS 0.036454f
C2115 PAD.n1469 VSS 0.036454f
C2116 PAD.n1470 VSS 0.036454f
C2117 PAD.n1471 VSS 0.036454f
C2118 PAD.n1472 VSS 0.036454f
C2119 PAD.n1474 VSS 0.036454f
C2120 PAD.n1475 VSS 0.036454f
C2121 PAD.n1476 VSS 0.036454f
C2122 PAD.n1477 VSS 0.036454f
C2123 PAD.n1478 VSS 0.036454f
C2124 PAD.n1479 VSS 0.036454f
C2125 PAD.n1480 VSS 0.023105f
C2126 PAD.n1481 VSS 0.023105f
C2127 PAD.n1483 VSS 0.42912f
C2128 PAD.n1484 VSS 0.049106f
C2129 PAD.n1485 VSS 0.049106f
C2130 PAD.n1486 VSS 0.033766f
C2131 PAD.n1487 VSS 0.029431f
C2132 PAD.n1488 VSS 0.029431f
C2133 PAD.n1489 VSS 0.685606f
C2134 PAD.n1531 VSS 0.023105f
C2135 PAD.n1532 VSS 0.586957f
C2136 PAD.n1533 VSS 0.611619f
C2137 PAD.n1534 VSS 0.685606f
C2138 PAD.n1535 VSS 0.023105f
C2139 PAD.n1536 VSS 0.44885f
C2140 PAD.n1537 VSS 0.036454f
C2141 PAD.n1538 VSS 0.036454f
C2142 PAD.n1539 VSS 0.036454f
C2143 PAD.n1540 VSS 0.036454f
C2144 PAD.n1541 VSS 0.036454f
C2145 PAD.n1542 VSS 0.036454f
C2146 PAD.n1543 VSS 0.036454f
C2147 PAD.n1544 VSS 0.036454f
C2148 PAD.n1545 VSS 0.036454f
C2149 PAD.n1546 VSS 0.036454f
C2150 PAD.n1547 VSS 0.036454f
C2151 PAD.n1548 VSS 0.036454f
C2152 PAD.n1549 VSS 0.036454f
C2153 PAD.n1550 VSS 0.036454f
C2154 PAD.n1551 VSS 0.036454f
C2155 PAD.n1552 VSS 0.036454f
C2156 PAD.n1553 VSS 0.036454f
C2157 PAD.n1554 VSS 0.036454f
C2158 PAD.n1555 VSS 0.036454f
C2159 PAD.n1556 VSS 0.036454f
C2160 PAD.n1557 VSS 0.036454f
C2161 PAD.n1558 VSS 0.036454f
C2162 PAD.n1559 VSS 0.036454f
C2163 PAD.n1560 VSS 0.036454f
C2164 PAD.n1561 VSS 0.036454f
C2165 PAD.n1562 VSS 0.036454f
C2166 PAD.n1563 VSS 0.036454f
C2167 PAD.n1564 VSS 0.036454f
C2168 PAD.n1565 VSS 0.036454f
C2169 PAD.n1566 VSS 0.036454f
C2170 PAD.n1567 VSS 0.036454f
C2171 PAD.n1568 VSS 0.036454f
C2172 PAD.n1569 VSS 0.036454f
C2173 PAD.n1570 VSS 0.036454f
C2174 PAD.n1571 VSS 0.036454f
C2175 PAD.n1572 VSS 0.036454f
C2176 PAD.n1573 VSS 0.036454f
C2177 PAD.n1574 VSS 0.036454f
C2178 PAD.n1575 VSS 0.036454f
C2179 PAD.n1576 VSS 0.036454f
C2180 PAD.n1578 VSS 0.036454f
C2181 PAD.n1579 VSS 0.036454f
C2182 PAD.n1580 VSS 0.046278f
C2183 PAD.n1581 VSS 0.064127f
C2184 PAD.n1582 VSS 0.069752f
C2185 PAD.n1583 VSS 0.062262f
C2186 PAD.n1584 VSS 0.036152f
C2187 PAD.n1585 VSS 0.069752f
C2188 PAD.n1586 VSS 0.611619f
C2189 PAD.n1587 VSS 0.049106f
C2190 PAD.n1588 VSS 0.049106f
C2191 PAD.n1589 VSS 0.033766f
C2192 PAD.n1590 VSS 0.029431f
C2193 PAD.n1591 VSS 0.029431f
C2194 PAD.n1592 VSS 0.596822f
C2195 PAD.n1593 VSS 0.542565f
C2196 PAD.n1594 VSS 0.611619f
C2197 PAD.n1595 VSS 0.039754f
C2198 PAD.n1596 VSS 0.039754f
C2199 PAD.n1597 VSS 0.069752f
C2200 PAD.n1598 VSS 0.036454f
C2201 PAD.n1599 VSS 0.023105f
C2202 PAD.n1600 VSS 0.036454f
C2203 PAD.n1603 VSS 0.036454f
C2204 PAD.n1604 VSS 0.036454f
C2205 PAD.n1605 VSS 0.036454f
C2206 PAD.n1606 VSS 0.036454f
C2207 PAD.n1608 VSS 0.036454f
C2208 PAD.n1609 VSS 0.036454f
C2209 PAD.n1610 VSS 0.036454f
C2210 PAD.n1612 VSS 0.036454f
C2211 PAD.n1613 VSS 0.036454f
C2212 PAD.n1614 VSS 0.036454f
C2213 PAD.n1616 VSS 0.036454f
C2214 PAD.n1617 VSS 0.036454f
C2215 PAD.n1618 VSS 0.036454f
C2216 PAD.n1620 VSS 0.036454f
C2217 PAD.n1621 VSS 0.036454f
C2218 PAD.n1622 VSS 0.036454f
C2219 PAD.n1624 VSS 0.036454f
C2220 PAD.n1625 VSS 0.036454f
C2221 PAD.n1626 VSS 0.036454f
C2222 PAD.n1628 VSS 0.036454f
C2223 PAD.n1629 VSS 0.036454f
C2224 PAD.n1630 VSS 0.036454f
C2225 PAD.n1632 VSS 0.036454f
C2226 PAD.n1633 VSS 0.036454f
C2227 PAD.n1634 VSS 0.036454f
C2228 PAD.n1636 VSS 0.036454f
C2229 PAD.n1637 VSS 0.036454f
C2230 PAD.n1638 VSS 0.036454f
C2231 PAD.n1640 VSS 0.036454f
C2232 PAD.n1641 VSS 0.036454f
C2233 PAD.n1642 VSS 0.036454f
C2234 PAD.n1644 VSS 0.036454f
C2235 PAD.n1645 VSS 0.036454f
C2236 PAD.n1646 VSS 0.036454f
C2237 PAD.n1648 VSS 0.036454f
C2238 PAD.n1649 VSS 0.036454f
C2239 PAD.n1650 VSS 0.036454f
C2240 PAD.n1652 VSS 0.036454f
C2241 PAD.n1653 VSS 0.036454f
C2242 PAD.n1654 VSS 0.036454f
C2243 PAD.n1656 VSS 0.036454f
C2244 PAD.n1657 VSS 0.036454f
C2245 PAD.n1658 VSS 0.036454f
C2246 PAD.n1660 VSS 0.036454f
C2247 PAD.n1661 VSS 0.036454f
C2248 PAD.n1662 VSS 0.036454f
C2249 PAD.n1664 VSS 0.036454f
C2250 PAD.n1665 VSS 0.036454f
C2251 PAD.n1666 VSS 0.036454f
C2252 PAD.n1668 VSS 0.036454f
C2253 PAD.n1669 VSS 0.036454f
C2254 PAD.n1670 VSS 0.036454f
C2255 PAD.n1672 VSS 0.036454f
C2256 PAD.n1673 VSS 0.036454f
C2257 PAD.n1674 VSS 0.036454f
C2258 PAD.n1676 VSS 0.036454f
C2259 PAD.n1677 VSS 0.036454f
C2260 PAD.n1678 VSS 0.036454f
C2261 PAD.n1680 VSS 0.036454f
C2262 PAD.n1681 VSS 0.036454f
C2263 PAD.n1682 VSS 0.036454f
C2264 PAD.n1683 VSS 0.03055f
C2265 PAD.n1684 VSS 0.023105f
C2266 PAD.n1685 VSS 0.023105f
C2267 PAD.n1687 VSS 0.036454f
C2268 PAD.n1689 VSS 0.036454f
C2269 PAD.n1691 VSS 0.036454f
C2270 PAD.n1692 VSS 0.036454f
C2271 PAD.n1693 VSS 0.036454f
C2272 PAD.n1694 VSS 0.036454f
C2273 PAD.n1695 VSS 0.036454f
C2274 PAD.n1696 VSS 0.036454f
C2275 PAD.n1697 VSS 0.036454f
C2276 PAD.n1699 VSS 0.036454f
C2277 PAD.n1701 VSS 0.036454f
C2278 PAD.n1703 VSS 0.036454f
C2279 PAD.n1704 VSS 0.036454f
C2280 PAD.n1705 VSS 0.036454f
C2281 PAD.n1706 VSS 0.036454f
C2282 PAD.n1707 VSS 0.036454f
C2283 PAD.n1708 VSS 0.036454f
C2284 PAD.n1709 VSS 0.036454f
C2285 PAD.n1711 VSS 0.036454f
C2286 PAD.n1713 VSS 0.036454f
C2287 PAD.n1715 VSS 0.036454f
C2288 PAD.n1716 VSS 0.036454f
C2289 PAD.n1717 VSS 0.036454f
C2290 PAD.n1718 VSS 0.036454f
C2291 PAD.n1719 VSS 0.036454f
C2292 PAD.n1720 VSS 0.036454f
C2293 PAD.n1721 VSS 0.036454f
C2294 PAD.n1723 VSS 0.036454f
C2295 PAD.n1725 VSS 0.036454f
C2296 PAD.n1727 VSS 0.036454f
C2297 PAD.n1728 VSS 0.036454f
C2298 PAD.n1729 VSS 0.036454f
C2299 PAD.n1730 VSS 0.036454f
C2300 PAD.n1731 VSS 0.036454f
C2301 PAD.n1732 VSS 0.036454f
C2302 PAD.n1733 VSS 0.036454f
C2303 PAD.n1735 VSS 0.036454f
C2304 PAD.n1737 VSS 0.036454f
C2305 PAD.n1739 VSS 0.036454f
C2306 PAD.n1740 VSS 0.036454f
C2307 PAD.n1741 VSS 0.036454f
C2308 PAD.n1742 VSS 0.036454f
C2309 PAD.n1743 VSS 0.036454f
C2310 PAD.n1744 VSS 0.036454f
C2311 PAD.n1745 VSS 0.036454f
C2312 PAD.n1747 VSS 0.036454f
C2313 PAD.n1749 VSS 0.036454f
C2314 PAD.n1751 VSS 0.036454f
C2315 PAD.n1752 VSS 0.036454f
C2316 PAD.n1753 VSS 0.036454f
C2317 PAD.n1754 VSS 0.036454f
C2318 PAD.n1755 VSS 0.036454f
C2319 PAD.n1756 VSS 0.036454f
C2320 PAD.n1757 VSS 0.036454f
C2321 PAD.n1759 VSS 0.036454f
C2322 PAD.n1761 VSS 0.036454f
C2323 PAD.n1763 VSS 0.036454f
C2324 PAD.n1764 VSS 0.036454f
C2325 PAD.n1765 VSS 0.036454f
C2326 PAD.n1766 VSS 0.036454f
C2327 PAD.n1767 VSS 0.036454f
C2328 PAD.n1768 VSS 0.036454f
C2329 PAD.n1769 VSS 0.036454f
C2330 PAD.n1771 VSS 0.036454f
C2331 PAD.n1773 VSS 0.036454f
C2332 PAD.n1775 VSS 0.036454f
C2333 PAD.n1776 VSS 0.036454f
C2334 PAD.n1777 VSS 0.036454f
C2335 PAD.n1778 VSS 0.036454f
C2336 PAD.n1779 VSS 0.036454f
C2337 PAD.n1780 VSS 0.036454f
C2338 PAD.n1781 VSS 0.036454f
C2339 PAD.n1783 VSS 0.036454f
C2340 PAD.n1785 VSS 0.036454f
C2341 PAD.n1787 VSS 0.036454f
C2342 PAD.n1788 VSS 0.036454f
C2343 PAD.n1789 VSS 0.036454f
C2344 PAD.n1790 VSS 0.036454f
C2345 PAD.n1791 VSS 0.036454f
C2346 PAD.n1792 VSS 0.036454f
C2347 PAD.n1793 VSS 0.036454f
C2348 PAD.n1795 VSS 0.036454f
C2349 PAD.n1797 VSS 0.036454f
C2350 PAD.n1799 VSS 0.036454f
C2351 PAD.n1800 VSS 0.036454f
C2352 PAD.n1801 VSS 0.036454f
C2353 PAD.n1802 VSS 0.036454f
C2354 PAD.n1803 VSS 0.036454f
C2355 PAD.n1804 VSS 0.036454f
C2356 PAD.n1805 VSS 0.036454f
C2357 PAD.n1807 VSS 0.036454f
C2358 PAD.n1809 VSS 0.036454f
C2359 PAD.n1811 VSS 0.036454f
C2360 PAD.n1812 VSS 0.036454f
C2361 PAD.n1813 VSS 0.036454f
C2362 PAD.n1814 VSS 0.036454f
C2363 PAD.n1815 VSS 0.036454f
C2364 PAD.n1816 VSS 0.036454f
C2365 PAD.n1817 VSS 0.036454f
C2366 PAD.n1819 VSS 0.036454f
C2367 PAD.n1821 VSS 0.036454f
C2368 PAD.n1823 VSS 0.036454f
C2369 PAD.n1824 VSS 0.036454f
C2370 PAD.n1825 VSS 0.036454f
C2371 PAD.n1826 VSS 0.036454f
C2372 PAD.n1827 VSS 0.036454f
C2373 PAD.n1828 VSS 0.036454f
C2374 PAD.n1829 VSS 0.036454f
C2375 PAD.n1831 VSS 0.036454f
C2376 PAD.n1833 VSS 0.036454f
C2377 PAD.n1835 VSS 0.036454f
C2378 PAD.n1836 VSS 0.036454f
C2379 PAD.n1837 VSS 0.036454f
C2380 PAD.n1838 VSS 0.036454f
C2381 PAD.n1839 VSS 0.036454f
C2382 PAD.n1840 VSS 0.036454f
C2383 PAD.n1841 VSS 0.036454f
C2384 PAD.n1843 VSS 0.036454f
C2385 PAD.n1845 VSS 0.036454f
C2386 PAD.n1847 VSS 0.036454f
C2387 PAD.n1848 VSS 0.036454f
C2388 PAD.n1849 VSS 0.036454f
C2389 PAD.n1850 VSS 0.036454f
C2390 PAD.n1851 VSS 0.036454f
C2391 PAD.n1852 VSS 0.036454f
C2392 PAD.n1853 VSS 0.036454f
C2393 PAD.n1855 VSS 0.036454f
C2394 PAD.n1857 VSS 0.036454f
C2395 PAD.n1859 VSS 0.036454f
C2396 PAD.n1860 VSS 0.036454f
C2397 PAD.n1861 VSS 0.036454f
C2398 PAD.n1862 VSS 0.036454f
C2399 PAD.n1863 VSS 0.036454f
C2400 PAD.n1864 VSS 0.036454f
C2401 PAD.n1865 VSS 0.036454f
C2402 PAD.n1867 VSS 0.036454f
C2403 PAD.n1869 VSS 0.036454f
C2404 PAD.n1871 VSS 0.036454f
C2405 PAD.n1872 VSS 0.036454f
C2406 PAD.n1873 VSS 0.036454f
C2407 PAD.n1874 VSS 0.036454f
C2408 PAD.n1875 VSS 0.036454f
C2409 PAD.n1876 VSS 0.036454f
C2410 PAD.n1877 VSS 0.036454f
C2411 PAD.n1879 VSS 0.036454f
C2412 PAD.n1881 VSS 0.036454f
C2413 PAD.n1883 VSS 0.036454f
C2414 PAD.n1884 VSS 0.036454f
C2415 PAD.n1885 VSS 0.036454f
C2416 PAD.n1886 VSS 0.036454f
C2417 PAD.n1887 VSS 0.036454f
C2418 PAD.n1888 VSS 0.036454f
C2419 PAD.n1889 VSS 0.036454f
C2420 PAD.n1891 VSS 0.036454f
C2421 PAD.n1893 VSS 0.036454f
C2422 PAD.n1895 VSS 0.036454f
C2423 PAD.n1896 VSS 0.036454f
C2424 PAD.n1897 VSS 0.036454f
C2425 PAD.n1898 VSS 0.036454f
C2426 PAD.n1899 VSS 0.036454f
C2427 PAD.n1900 VSS 0.036454f
C2428 PAD.n1901 VSS 0.036454f
C2429 PAD.n1903 VSS 0.036454f
C2430 PAD.n1905 VSS 0.036454f
C2431 PAD.n1907 VSS 0.036454f
C2432 PAD.n1908 VSS 0.036454f
C2433 PAD.n1909 VSS 0.036454f
C2434 PAD.n1910 VSS 0.036454f
C2435 PAD.n1911 VSS 0.036454f
C2436 PAD.n1912 VSS 0.036454f
C2437 PAD.n1913 VSS 0.036454f
C2438 PAD.n1915 VSS 0.036454f
C2439 PAD.n1917 VSS 0.036454f
C2440 PAD.n1919 VSS 0.036454f
C2441 PAD.n1920 VSS 0.036454f
C2442 PAD.n1921 VSS 0.036454f
C2443 PAD.n1922 VSS 0.036454f
C2444 PAD.n1923 VSS 0.036454f
C2445 PAD.n1924 VSS 0.036454f
C2446 PAD.n1925 VSS 0.036454f
C2447 PAD.n1927 VSS 0.036454f
C2448 PAD.n1929 VSS 0.036454f
C2449 PAD.n1930 VSS 0.036454f
C2450 PAD.n1931 VSS 0.023105f
C2451 PAD.n1932 VSS 0.033374f
C2452 PAD.n1933 VSS 0.062262f
C2453 PAD.n1934 VSS 0.069752f
C2454 PAD.n1935 VSS 0.069752f
C2455 PAD.n1936 VSS 0.700403f
C2456 PAD.n1937 VSS 0.049106f
C2457 PAD.n1938 VSS 0.049106f
C2458 PAD.n1939 VSS 0.033766f
C2459 PAD.n1940 VSS 0.029431f
C2460 PAD.n1941 VSS 0.029431f
C2461 PAD.n1942 VSS 0.438985f
C2462 PAD.n1984 VSS 0.023105f
C2463 PAD.n1985 VSS 0.611619f
C2464 PAD.n1986 VSS 0.438985f
C2465 PAD.n1987 VSS 0.023105f
C2466 PAD.n1988 VSS 0.369931f
C2467 PAD.n1989 VSS 0.036454f
C2468 PAD.n1990 VSS 0.036454f
C2469 PAD.n1991 VSS 0.036454f
C2470 PAD.n1992 VSS 0.036454f
C2471 PAD.n1993 VSS 0.036454f
C2472 PAD.n1994 VSS 0.036454f
C2473 PAD.n1995 VSS 0.036454f
C2474 PAD.n1996 VSS 0.036454f
C2475 PAD.n1997 VSS 0.036454f
C2476 PAD.n1998 VSS 0.036454f
C2477 PAD.n1999 VSS 0.036454f
C2478 PAD.n2000 VSS 0.036454f
C2479 PAD.n2001 VSS 0.036454f
C2480 PAD.n2002 VSS 0.036454f
C2481 PAD.n2003 VSS 0.036454f
C2482 PAD.n2004 VSS 0.036454f
C2483 PAD.n2005 VSS 0.036454f
C2484 PAD.n2006 VSS 0.036454f
C2485 PAD.n2007 VSS 0.036454f
C2486 PAD.n2008 VSS 0.036454f
C2487 PAD.n2009 VSS 0.036454f
C2488 PAD.n2010 VSS 0.036454f
C2489 PAD.n2011 VSS 0.036454f
C2490 PAD.n2012 VSS 0.036454f
C2491 PAD.n2013 VSS 0.036454f
C2492 PAD.n2014 VSS 0.036454f
C2493 PAD.n2015 VSS 0.036454f
C2494 PAD.n2016 VSS 0.036454f
C2495 PAD.n2017 VSS 0.036454f
C2496 PAD.n2018 VSS 0.036454f
C2497 PAD.n2019 VSS 0.036454f
C2498 PAD.n2020 VSS 0.036454f
C2499 PAD.n2021 VSS 0.036454f
C2500 PAD.n2022 VSS 0.036454f
C2501 PAD.n2023 VSS 0.036454f
C2502 PAD.n2024 VSS 0.036454f
C2503 PAD.n2025 VSS 0.036454f
C2504 PAD.n2026 VSS 0.036454f
C2505 PAD.n2027 VSS 0.036454f
C2506 PAD.n2028 VSS 0.036454f
C2507 PAD.n2030 VSS 0.036454f
C2508 PAD.n2031 VSS 0.036454f
C2509 PAD.n2032 VSS 0.046278f
C2510 PAD.n2033 VSS 0.048377f
C2511 PAD.n2034 VSS 0.050211f
C2512 PAD.n2035 VSS 0.064127f
C2513 PAD.n2036 VSS 0.069752f
C2514 PAD.n2037 VSS 0.611619f
C2515 PAD.n2038 VSS 0.047896f
C2516 PAD.n2039 VSS 0.047896f
C2517 PAD.n2040 VSS 0.03055f
C2518 PAD.n2041 VSS 0.042887f
C2519 PAD.n2042 VSS 0.049106f
C2520 PAD.n2043 VSS 0.029431f
C2521 PAD.n2044 VSS 0.049106f
C2522 PAD.n2045 VSS 0.029431f
C2523 PAD.n2046 VSS 0.310742f
C2524 PAD.n2088 VSS 0.023105f
C2525 PAD.n2089 VSS 0.310742f
C2526 PAD.n2090 VSS 0.023105f
C2527 PAD.n2091 VSS 0.61162f
C2528 PAD.n2092 VSS 0.036454f
C2529 PAD.n2093 VSS 0.036454f
C2530 PAD.n2094 VSS 0.036454f
C2531 PAD.n2095 VSS 0.036454f
C2532 PAD.n2096 VSS 0.036454f
C2533 PAD.n2097 VSS 0.036454f
C2534 PAD.n2098 VSS 0.036454f
C2535 PAD.n2099 VSS 0.036454f
C2536 PAD.n2100 VSS 0.036454f
C2537 PAD.n2101 VSS 0.036454f
C2538 PAD.n2102 VSS 0.036454f
C2539 PAD.n2103 VSS 0.036454f
C2540 PAD.n2104 VSS 0.036454f
C2541 PAD.n2105 VSS 0.036454f
C2542 PAD.n2106 VSS 0.036454f
C2543 PAD.n2107 VSS 0.036454f
C2544 PAD.n2108 VSS 0.036454f
C2545 PAD.n2109 VSS 0.036454f
C2546 PAD.n2110 VSS 0.036454f
C2547 PAD.n2111 VSS 0.036454f
C2548 PAD.n2112 VSS 0.036454f
C2549 PAD.n2113 VSS 0.036454f
C2550 PAD.n2114 VSS 0.036454f
C2551 PAD.n2115 VSS 0.036454f
C2552 PAD.n2116 VSS 0.036454f
C2553 PAD.n2117 VSS 0.036454f
C2554 PAD.n2118 VSS 0.036454f
C2555 PAD.n2119 VSS 0.036454f
C2556 PAD.n2120 VSS 0.036454f
C2557 PAD.n2121 VSS 0.036454f
C2558 PAD.n2122 VSS 0.036454f
C2559 PAD.n2123 VSS 0.036454f
C2560 PAD.n2124 VSS 0.036454f
C2561 PAD.n2125 VSS 0.036454f
C2562 PAD.n2126 VSS 0.036454f
C2563 PAD.n2127 VSS 0.036454f
C2564 PAD.n2128 VSS 0.036454f
C2565 PAD.n2129 VSS 0.036454f
C2566 PAD.n2130 VSS 0.036454f
C2567 PAD.n2131 VSS 0.036454f
C2568 PAD.n2133 VSS 0.036454f
C2569 PAD.n2134 VSS 0.036454f
C2570 PAD.n2135 VSS 0.046278f
C2571 PAD.n2136 VSS 0.069752f
C2572 PAD.n2137 VSS 0.036152f
C2573 PAD.n2138 VSS 0.069752f
C2574 PAD.n2139 VSS 0.498174f
C2575 PAD.n2140 VSS 0.029431f
C2576 PAD.n2141 VSS 0.029431f
C2577 PAD.n2142 VSS 0.03055f
C2578 PAD.n2143 VSS 0.042887f
C2579 PAD.n2144 VSS 0.049106f
C2580 PAD.n2145 VSS 0.049106f
C2581 PAD.n2146 VSS 0.40939f
C2582 PAD.n2147 VSS 0.039754f
C2583 PAD.n2148 VSS 0.039754f
C2584 PAD.n2149 VSS 0.069752f
C2585 PAD.n2150 VSS 0.036454f
C2586 PAD.n2151 VSS 0.023105f
C2587 PAD.n2152 VSS 0.036454f
C2588 PAD.n2155 VSS 0.036454f
C2589 PAD.n2156 VSS 0.036454f
C2590 PAD.n2157 VSS 0.036454f
C2591 PAD.n2158 VSS 0.036454f
C2592 PAD.n2160 VSS 0.036454f
C2593 PAD.n2161 VSS 0.036454f
C2594 PAD.n2162 VSS 0.036454f
C2595 PAD.n2164 VSS 0.036454f
C2596 PAD.n2165 VSS 0.036454f
C2597 PAD.n2166 VSS 0.036454f
C2598 PAD.n2168 VSS 0.036454f
C2599 PAD.n2169 VSS 0.036454f
C2600 PAD.n2170 VSS 0.036454f
C2601 PAD.n2172 VSS 0.036454f
C2602 PAD.n2173 VSS 0.036454f
C2603 PAD.n2174 VSS 0.036454f
C2604 PAD.n2176 VSS 0.036454f
C2605 PAD.n2177 VSS 0.036454f
C2606 PAD.n2178 VSS 0.036454f
C2607 PAD.n2180 VSS 0.036454f
C2608 PAD.n2181 VSS 0.036454f
C2609 PAD.n2182 VSS 0.036454f
C2610 PAD.n2184 VSS 0.036454f
C2611 PAD.n2185 VSS 0.036454f
C2612 PAD.n2186 VSS 0.036454f
C2613 PAD.n2188 VSS 0.036454f
C2614 PAD.n2189 VSS 0.036454f
C2615 PAD.n2190 VSS 0.036454f
C2616 PAD.n2192 VSS 0.036454f
C2617 PAD.n2193 VSS 0.036454f
C2618 PAD.n2194 VSS 0.036454f
C2619 PAD.n2196 VSS 0.036454f
C2620 PAD.n2197 VSS 0.036454f
C2621 PAD.n2198 VSS 0.036454f
C2622 PAD.n2200 VSS 0.036454f
C2623 PAD.n2201 VSS 0.036454f
C2624 PAD.n2202 VSS 0.036454f
C2625 PAD.n2204 VSS 0.036454f
C2626 PAD.n2205 VSS 0.036454f
C2627 PAD.n2206 VSS 0.036454f
C2628 PAD.n2208 VSS 0.036454f
C2629 PAD.n2209 VSS 0.036454f
C2630 PAD.n2210 VSS 0.036454f
C2631 PAD.n2212 VSS 0.036454f
C2632 PAD.n2213 VSS 0.036454f
C2633 PAD.n2214 VSS 0.036454f
C2634 PAD.n2216 VSS 0.036454f
C2635 PAD.n2217 VSS 0.036454f
C2636 PAD.n2218 VSS 0.036454f
C2637 PAD.n2220 VSS 0.036454f
C2638 PAD.n2221 VSS 0.036454f
C2639 PAD.n2222 VSS 0.036454f
C2640 PAD.n2224 VSS 0.036454f
C2641 PAD.n2225 VSS 0.036454f
C2642 PAD.n2226 VSS 0.036454f
C2643 PAD.n2228 VSS 0.036454f
C2644 PAD.n2229 VSS 0.036454f
C2645 PAD.n2230 VSS 0.036454f
C2646 PAD.n2232 VSS 0.036454f
C2647 PAD.n2233 VSS 0.036454f
C2648 PAD.n2234 VSS 0.036454f
C2649 PAD.n2235 VSS 0.023105f
C2650 PAD.n2236 VSS 0.023105f
C2651 PAD.n2238 VSS 0.036454f
C2652 PAD.n2240 VSS 0.036454f
C2653 PAD.n2242 VSS 0.036454f
C2654 PAD.n2243 VSS 0.036454f
C2655 PAD.n2244 VSS 0.036454f
C2656 PAD.n2245 VSS 0.036454f
C2657 PAD.n2246 VSS 0.036454f
C2658 PAD.n2247 VSS 0.036454f
C2659 PAD.n2248 VSS 0.036454f
C2660 PAD.n2250 VSS 0.036454f
C2661 PAD.n2252 VSS 0.036454f
C2662 PAD.n2254 VSS 0.036454f
C2663 PAD.n2255 VSS 0.036454f
C2664 PAD.n2256 VSS 0.036454f
C2665 PAD.n2257 VSS 0.036454f
C2666 PAD.n2258 VSS 0.036454f
C2667 PAD.n2259 VSS 0.036454f
C2668 PAD.n2260 VSS 0.036454f
C2669 PAD.n2262 VSS 0.036454f
C2670 PAD.n2264 VSS 0.036454f
C2671 PAD.n2266 VSS 0.036454f
C2672 PAD.n2267 VSS 0.036454f
C2673 PAD.n2268 VSS 0.036454f
C2674 PAD.n2269 VSS 0.036454f
C2675 PAD.n2270 VSS 0.036454f
C2676 PAD.n2271 VSS 0.036454f
C2677 PAD.n2272 VSS 0.036454f
C2678 PAD.n2274 VSS 0.036454f
C2679 PAD.n2276 VSS 0.036454f
C2680 PAD.n2278 VSS 0.036454f
C2681 PAD.n2279 VSS 0.036454f
C2682 PAD.n2280 VSS 0.036454f
C2683 PAD.n2281 VSS 0.036454f
C2684 PAD.n2282 VSS 0.036454f
C2685 PAD.n2283 VSS 0.036454f
C2686 PAD.n2284 VSS 0.036454f
C2687 PAD.n2286 VSS 0.036454f
C2688 PAD.n2288 VSS 0.036454f
C2689 PAD.n2290 VSS 0.036454f
C2690 PAD.n2291 VSS 0.036454f
C2691 PAD.n2292 VSS 0.036454f
C2692 PAD.n2293 VSS 0.036454f
C2693 PAD.n2294 VSS 0.036454f
C2694 PAD.n2295 VSS 0.036454f
C2695 PAD.n2296 VSS 0.036454f
C2696 PAD.n2298 VSS 0.036454f
C2697 PAD.n2300 VSS 0.036454f
C2698 PAD.n2302 VSS 0.036454f
C2699 PAD.n2303 VSS 0.036454f
C2700 PAD.n2304 VSS 0.036454f
C2701 PAD.n2305 VSS 0.036454f
C2702 PAD.n2306 VSS 0.036454f
C2703 PAD.n2307 VSS 0.036454f
C2704 PAD.n2308 VSS 0.036454f
C2705 PAD.n2310 VSS 0.036454f
C2706 PAD.n2312 VSS 0.036454f
C2707 PAD.n2314 VSS 0.036454f
C2708 PAD.n2315 VSS 0.036454f
C2709 PAD.n2316 VSS 0.036454f
C2710 PAD.n2317 VSS 0.036454f
C2711 PAD.n2318 VSS 0.036454f
C2712 PAD.n2319 VSS 0.036454f
C2713 PAD.n2320 VSS 0.036454f
C2714 PAD.n2322 VSS 0.036454f
C2715 PAD.n2324 VSS 0.036454f
C2716 PAD.n2326 VSS 0.036454f
C2717 PAD.n2327 VSS 0.036454f
C2718 PAD.n2328 VSS 0.036454f
C2719 PAD.n2329 VSS 0.036454f
C2720 PAD.n2330 VSS 0.036454f
C2721 PAD.n2331 VSS 0.036454f
C2722 PAD.n2332 VSS 0.036454f
C2723 PAD.n2334 VSS 0.036454f
C2724 PAD.n2336 VSS 0.036454f
C2725 PAD.n2338 VSS 0.036454f
C2726 PAD.n2339 VSS 0.036454f
C2727 PAD.n2340 VSS 0.036454f
C2728 PAD.n2341 VSS 0.036454f
C2729 PAD.n2342 VSS 0.036454f
C2730 PAD.n2343 VSS 0.036454f
C2731 PAD.n2344 VSS 0.036454f
C2732 PAD.n2346 VSS 0.036454f
C2733 PAD.n2348 VSS 0.036454f
C2734 PAD.n2350 VSS 0.036454f
C2735 PAD.n2351 VSS 0.036454f
C2736 PAD.n2352 VSS 0.036454f
C2737 PAD.n2353 VSS 0.036454f
C2738 PAD.n2354 VSS 0.036454f
C2739 PAD.n2355 VSS 0.036454f
C2740 PAD.n2356 VSS 0.036454f
C2741 PAD.n2358 VSS 0.036454f
C2742 PAD.n2360 VSS 0.036454f
C2743 PAD.n2362 VSS 0.036454f
C2744 PAD.n2363 VSS 0.036454f
C2745 PAD.n2364 VSS 0.036454f
C2746 PAD.n2365 VSS 0.036454f
C2747 PAD.n2366 VSS 0.036454f
C2748 PAD.n2367 VSS 0.036454f
C2749 PAD.n2368 VSS 0.036454f
C2750 PAD.n2370 VSS 0.036454f
C2751 PAD.n2372 VSS 0.036454f
C2752 PAD.n2374 VSS 0.036454f
C2753 PAD.n2375 VSS 0.036454f
C2754 PAD.n2376 VSS 0.036454f
C2755 PAD.n2377 VSS 0.036454f
C2756 PAD.n2378 VSS 0.036454f
C2757 PAD.n2379 VSS 0.036454f
C2758 PAD.n2380 VSS 0.036454f
C2759 PAD.n2382 VSS 0.036454f
C2760 PAD.n2384 VSS 0.036454f
C2761 PAD.n2386 VSS 0.036454f
C2762 PAD.n2387 VSS 0.036454f
C2763 PAD.n2388 VSS 0.036454f
C2764 PAD.n2389 VSS 0.036454f
C2765 PAD.n2390 VSS 0.036454f
C2766 PAD.n2391 VSS 0.036454f
C2767 PAD.n2392 VSS 0.036454f
C2768 PAD.n2394 VSS 0.036454f
C2769 PAD.n2396 VSS 0.036454f
C2770 PAD.n2398 VSS 0.036454f
C2771 PAD.n2399 VSS 0.036454f
C2772 PAD.n2400 VSS 0.036454f
C2773 PAD.n2401 VSS 0.036454f
C2774 PAD.n2402 VSS 0.036454f
C2775 PAD.n2403 VSS 0.036454f
C2776 PAD.n2404 VSS 0.036454f
C2777 PAD.n2406 VSS 0.036454f
C2778 PAD.n2408 VSS 0.036454f
C2779 PAD.n2410 VSS 0.036454f
C2780 PAD.n2411 VSS 0.036454f
C2781 PAD.n2412 VSS 0.036454f
C2782 PAD.n2413 VSS 0.036454f
C2783 PAD.n2414 VSS 0.036454f
C2784 PAD.n2415 VSS 0.036454f
C2785 PAD.n2416 VSS 0.036454f
C2786 PAD.n2418 VSS 0.036454f
C2787 PAD.n2420 VSS 0.036454f
C2788 PAD.n2422 VSS 0.036454f
C2789 PAD.n2423 VSS 0.036454f
C2790 PAD.n2424 VSS 0.036454f
C2791 PAD.n2425 VSS 0.036454f
C2792 PAD.n2426 VSS 0.036454f
C2793 PAD.n2427 VSS 0.036454f
C2794 PAD.n2428 VSS 0.036454f
C2795 PAD.n2430 VSS 0.036454f
C2796 PAD.n2432 VSS 0.036454f
C2797 PAD.n2434 VSS 0.036454f
C2798 PAD.n2435 VSS 0.036454f
C2799 PAD.n2436 VSS 0.036454f
C2800 PAD.n2437 VSS 0.036454f
C2801 PAD.n2438 VSS 0.036454f
C2802 PAD.n2439 VSS 0.036454f
C2803 PAD.n2440 VSS 0.036454f
C2804 PAD.n2442 VSS 0.036454f
C2805 PAD.n2444 VSS 0.036454f
C2806 PAD.n2446 VSS 0.036454f
C2807 PAD.n2447 VSS 0.036454f
C2808 PAD.n2448 VSS 0.036454f
C2809 PAD.n2449 VSS 0.036454f
C2810 PAD.n2450 VSS 0.036454f
C2811 PAD.n2451 VSS 0.036454f
C2812 PAD.n2452 VSS 0.036454f
C2813 PAD.n2454 VSS 0.036454f
C2814 PAD.n2456 VSS 0.036454f
C2815 PAD.n2458 VSS 0.036454f
C2816 PAD.n2459 VSS 0.036454f
C2817 PAD.n2460 VSS 0.036454f
C2818 PAD.n2461 VSS 0.036454f
C2819 PAD.n2462 VSS 0.036454f
C2820 PAD.n2463 VSS 0.036454f
C2821 PAD.n2464 VSS 0.036454f
C2822 PAD.n2466 VSS 0.036454f
C2823 PAD.n2468 VSS 0.036454f
C2824 PAD.n2470 VSS 0.036454f
C2825 PAD.n2471 VSS 0.036454f
C2826 PAD.n2472 VSS 0.036454f
C2827 PAD.n2473 VSS 0.036454f
C2828 PAD.n2474 VSS 0.036454f
C2829 PAD.n2475 VSS 0.036454f
C2830 PAD.n2476 VSS 0.036454f
C2831 PAD.n2478 VSS 0.036454f
C2832 PAD.n2480 VSS 0.036454f
C2833 PAD.n2481 VSS 0.036454f
C2834 PAD.n2482 VSS 0.023105f
C2835 PAD.n2483 VSS 0.033374f
C2836 PAD.n2484 VSS 0.062262f
C2837 PAD.n2485 VSS 0.069752f
C2838 PAD.n2486 VSS 0.069752f
C2839 PAD.n2487 VSS 0.231823f
C2840 PAD.n2488 VSS 0.029431f
C2841 PAD.n2489 VSS 0.029431f
C2842 PAD.n2490 VSS 0.03055f
C2843 PAD.n2491 VSS 0.042887f
C2844 PAD.n2492 VSS 0.049106f
C2845 PAD.n2493 VSS 0.049106f
C2846 PAD.n2494 VSS 0.14304f
C2847 PAD.n2495 VSS 0.039754f
C2848 PAD.n2496 VSS 0.039754f
C2849 PAD.n2497 VSS 0.036454f
C2850 PAD.n2498 VSS 0.023105f
C2851 PAD.n2499 VSS 0.036454f
C2852 PAD.n2502 VSS 0.036454f
C2853 PAD.n2503 VSS 0.036454f
C2854 PAD.n2504 VSS 0.036454f
C2855 PAD.n2505 VSS 0.036454f
C2856 PAD.n2507 VSS 0.036454f
C2857 PAD.n2508 VSS 0.036454f
C2858 PAD.n2509 VSS 0.036454f
C2859 PAD.n2511 VSS 0.036454f
C2860 PAD.n2512 VSS 0.036454f
C2861 PAD.n2513 VSS 0.036454f
C2862 PAD.n2515 VSS 0.036454f
C2863 PAD.n2516 VSS 0.036454f
C2864 PAD.n2517 VSS 0.036454f
C2865 PAD.n2519 VSS 0.036454f
C2866 PAD.n2520 VSS 0.036454f
C2867 PAD.n2521 VSS 0.036454f
C2868 PAD.n2523 VSS 0.036454f
C2869 PAD.n2524 VSS 0.036454f
C2870 PAD.n2525 VSS 0.036454f
C2871 PAD.n2527 VSS 0.036454f
C2872 PAD.n2528 VSS 0.036454f
C2873 PAD.n2529 VSS 0.036454f
C2874 PAD.n2531 VSS 0.036454f
C2875 PAD.n2532 VSS 0.036454f
C2876 PAD.n2533 VSS 0.036454f
C2877 PAD.n2535 VSS 0.036454f
C2878 PAD.n2536 VSS 0.036454f
C2879 PAD.n2537 VSS 0.036454f
C2880 PAD.n2539 VSS 0.036454f
C2881 PAD.n2540 VSS 0.036454f
C2882 PAD.n2541 VSS 0.036454f
C2883 PAD.n2543 VSS 0.036454f
C2884 PAD.n2544 VSS 0.036454f
C2885 PAD.n2545 VSS 0.036454f
C2886 PAD.n2547 VSS 0.036454f
C2887 PAD.n2548 VSS 0.036454f
C2888 PAD.n2549 VSS 0.036454f
C2889 PAD.n2551 VSS 0.036454f
C2890 PAD.n2552 VSS 0.036454f
C2891 PAD.n2553 VSS 0.036454f
C2892 PAD.n2555 VSS 0.036454f
C2893 PAD.n2556 VSS 0.036454f
C2894 PAD.n2557 VSS 0.036454f
C2895 PAD.n2559 VSS 0.036454f
C2896 PAD.n2560 VSS 0.036454f
C2897 PAD.n2561 VSS 0.036454f
C2898 PAD.n2563 VSS 0.036454f
C2899 PAD.n2564 VSS 0.036454f
C2900 PAD.n2565 VSS 0.036454f
C2901 PAD.n2567 VSS 0.036454f
C2902 PAD.n2568 VSS 0.036454f
C2903 PAD.n2569 VSS 0.036454f
C2904 PAD.n2571 VSS 0.036454f
C2905 PAD.n2572 VSS 0.036454f
C2906 PAD.n2573 VSS 0.036454f
C2907 PAD.n2575 VSS 0.036454f
C2908 PAD.n2576 VSS 0.036454f
C2909 PAD.n2577 VSS 0.036454f
C2910 PAD.n2579 VSS 0.036454f
C2911 PAD.n2580 VSS 0.036454f
C2912 PAD.n2581 VSS 0.036454f
C2913 PAD.n2582 VSS 0.023105f
C2914 PAD.n2583 VSS 0.023105f
C2915 PAD.n2585 VSS 0.036454f
C2916 PAD.n2587 VSS 0.036454f
C2917 PAD.n2589 VSS 0.036454f
C2918 PAD.n2590 VSS 0.036454f
C2919 PAD.n2591 VSS 0.036454f
C2920 PAD.n2592 VSS 0.036454f
C2921 PAD.n2593 VSS 0.036454f
C2922 PAD.n2594 VSS 0.036454f
C2923 PAD.n2595 VSS 0.036454f
C2924 PAD.n2597 VSS 0.036454f
C2925 PAD.n2599 VSS 0.036454f
C2926 PAD.n2601 VSS 0.036454f
C2927 PAD.n2602 VSS 0.036454f
C2928 PAD.n2603 VSS 0.036454f
C2929 PAD.n2604 VSS 0.036454f
C2930 PAD.n2605 VSS 0.036454f
C2931 PAD.n2606 VSS 0.036454f
C2932 PAD.n2607 VSS 0.036454f
C2933 PAD.n2609 VSS 0.036454f
C2934 PAD.n2611 VSS 0.036454f
C2935 PAD.n2613 VSS 0.036454f
C2936 PAD.n2614 VSS 0.036454f
C2937 PAD.n2615 VSS 0.036454f
C2938 PAD.n2616 VSS 0.036454f
C2939 PAD.n2617 VSS 0.036454f
C2940 PAD.n2618 VSS 0.036454f
C2941 PAD.n2619 VSS 0.036454f
C2942 PAD.n2621 VSS 0.036454f
C2943 PAD.n2623 VSS 0.036454f
C2944 PAD.n2625 VSS 0.036454f
C2945 PAD.n2626 VSS 0.036454f
C2946 PAD.n2627 VSS 0.036454f
C2947 PAD.n2628 VSS 0.036454f
C2948 PAD.n2629 VSS 0.036454f
C2949 PAD.n2630 VSS 0.036454f
C2950 PAD.n2631 VSS 0.036454f
C2951 PAD.n2633 VSS 0.036454f
C2952 PAD.n2635 VSS 0.036454f
C2953 PAD.n2637 VSS 0.036454f
C2954 PAD.n2638 VSS 0.036454f
C2955 PAD.n2639 VSS 0.036454f
C2956 PAD.n2640 VSS 0.036454f
C2957 PAD.n2641 VSS 0.036454f
C2958 PAD.n2642 VSS 0.036454f
C2959 PAD.n2643 VSS 0.036454f
C2960 PAD.n2645 VSS 0.036454f
C2961 PAD.n2647 VSS 0.036454f
C2962 PAD.n2649 VSS 0.036454f
C2963 PAD.n2650 VSS 0.036454f
C2964 PAD.n2651 VSS 0.036454f
C2965 PAD.n2652 VSS 0.036454f
C2966 PAD.n2653 VSS 0.036454f
C2967 PAD.n2654 VSS 0.036454f
C2968 PAD.n2655 VSS 0.036454f
C2969 PAD.n2657 VSS 0.036454f
C2970 PAD.n2659 VSS 0.036454f
C2971 PAD.n2661 VSS 0.036454f
C2972 PAD.n2662 VSS 0.036454f
C2973 PAD.n2663 VSS 0.036454f
C2974 PAD.n2664 VSS 0.036454f
C2975 PAD.n2665 VSS 0.036454f
C2976 PAD.n2666 VSS 0.036454f
C2977 PAD.n2667 VSS 0.036454f
C2978 PAD.n2669 VSS 0.036454f
C2979 PAD.n2671 VSS 0.036454f
C2980 PAD.n2673 VSS 0.036454f
C2981 PAD.n2674 VSS 0.036454f
C2982 PAD.n2675 VSS 0.036454f
C2983 PAD.n2676 VSS 0.036454f
C2984 PAD.n2677 VSS 0.036454f
C2985 PAD.n2678 VSS 0.036454f
C2986 PAD.n2679 VSS 0.036454f
C2987 PAD.n2681 VSS 0.036454f
C2988 PAD.n2683 VSS 0.036454f
C2989 PAD.n2685 VSS 0.036454f
C2990 PAD.n2686 VSS 0.036454f
C2991 PAD.n2687 VSS 0.036454f
C2992 PAD.n2688 VSS 0.036454f
C2993 PAD.n2689 VSS 0.036454f
C2994 PAD.n2690 VSS 0.036454f
C2995 PAD.n2691 VSS 0.036454f
C2996 PAD.n2693 VSS 0.036454f
C2997 PAD.n2695 VSS 0.036454f
C2998 PAD.n2697 VSS 0.036454f
C2999 PAD.n2698 VSS 0.036454f
C3000 PAD.n2699 VSS 0.036454f
C3001 PAD.n2700 VSS 0.036454f
C3002 PAD.n2701 VSS 0.036454f
C3003 PAD.n2702 VSS 0.036454f
C3004 PAD.n2703 VSS 0.036454f
C3005 PAD.n2705 VSS 0.036454f
C3006 PAD.n2707 VSS 0.036454f
C3007 PAD.n2709 VSS 0.036454f
C3008 PAD.n2710 VSS 0.036454f
C3009 PAD.n2711 VSS 0.036454f
C3010 PAD.n2712 VSS 0.036454f
C3011 PAD.n2713 VSS 0.036454f
C3012 PAD.n2714 VSS 0.036454f
C3013 PAD.n2715 VSS 0.036454f
C3014 PAD.n2717 VSS 0.036454f
C3015 PAD.n2719 VSS 0.036454f
C3016 PAD.n2721 VSS 0.036454f
C3017 PAD.n2722 VSS 0.036454f
C3018 PAD.n2723 VSS 0.036454f
C3019 PAD.n2724 VSS 0.036454f
C3020 PAD.n2725 VSS 0.036454f
C3021 PAD.n2726 VSS 0.036454f
C3022 PAD.n2727 VSS 0.036454f
C3023 PAD.n2729 VSS 0.036454f
C3024 PAD.n2731 VSS 0.036454f
C3025 PAD.n2733 VSS 0.036454f
C3026 PAD.n2734 VSS 0.036454f
C3027 PAD.n2735 VSS 0.036454f
C3028 PAD.n2736 VSS 0.036454f
C3029 PAD.n2737 VSS 0.036454f
C3030 PAD.n2738 VSS 0.036454f
C3031 PAD.n2739 VSS 0.036454f
C3032 PAD.n2741 VSS 0.036454f
C3033 PAD.n2743 VSS 0.036454f
C3034 PAD.n2745 VSS 0.036454f
C3035 PAD.n2746 VSS 0.036454f
C3036 PAD.n2747 VSS 0.036454f
C3037 PAD.n2748 VSS 0.036454f
C3038 PAD.n2749 VSS 0.036454f
C3039 PAD.n2750 VSS 0.036454f
C3040 PAD.n2751 VSS 0.036454f
C3041 PAD.n2753 VSS 0.036454f
C3042 PAD.n2755 VSS 0.036454f
C3043 PAD.n2757 VSS 0.036454f
C3044 PAD.n2758 VSS 0.036454f
C3045 PAD.n2759 VSS 0.036454f
C3046 PAD.n2760 VSS 0.036454f
C3047 PAD.n2761 VSS 0.036454f
C3048 PAD.n2762 VSS 0.036454f
C3049 PAD.n2763 VSS 0.036454f
C3050 PAD.n2765 VSS 0.036454f
C3051 PAD.n2767 VSS 0.036454f
C3052 PAD.n2769 VSS 0.036454f
C3053 PAD.n2770 VSS 0.036454f
C3054 PAD.n2771 VSS 0.036454f
C3055 PAD.n2772 VSS 0.036454f
C3056 PAD.n2773 VSS 0.036454f
C3057 PAD.n2774 VSS 0.036454f
C3058 PAD.n2775 VSS 0.036454f
C3059 PAD.n2777 VSS 0.036454f
C3060 PAD.n2779 VSS 0.036454f
C3061 PAD.n2781 VSS 0.036454f
C3062 PAD.n2782 VSS 0.036454f
C3063 PAD.n2783 VSS 0.036454f
C3064 PAD.n2784 VSS 0.036454f
C3065 PAD.n2785 VSS 0.036454f
C3066 PAD.n2786 VSS 0.036454f
C3067 PAD.n2787 VSS 0.036454f
C3068 PAD.n2789 VSS 0.036454f
C3069 PAD.n2791 VSS 0.036454f
C3070 PAD.n2793 VSS 0.036454f
C3071 PAD.n2794 VSS 0.036454f
C3072 PAD.n2795 VSS 0.036454f
C3073 PAD.n2796 VSS 0.036454f
C3074 PAD.n2797 VSS 0.036454f
C3075 PAD.n2798 VSS 0.036454f
C3076 PAD.n2799 VSS 0.036454f
C3077 PAD.n2801 VSS 0.036454f
C3078 PAD.n2803 VSS 0.036454f
C3079 PAD.n2805 VSS 0.036454f
C3080 PAD.n2806 VSS 0.036454f
C3081 PAD.n2807 VSS 0.036454f
C3082 PAD.n2808 VSS 0.036454f
C3083 PAD.n2809 VSS 0.036454f
C3084 PAD.n2810 VSS 0.036454f
C3085 PAD.n2811 VSS 0.036454f
C3086 PAD.n2813 VSS 0.036454f
C3087 PAD.n2815 VSS 0.036454f
C3088 PAD.n2817 VSS 0.036454f
C3089 PAD.n2818 VSS 0.036454f
C3090 PAD.n2819 VSS 0.036454f
C3091 PAD.n2820 VSS 0.036454f
C3092 PAD.n2821 VSS 0.036454f
C3093 PAD.n2822 VSS 0.036454f
C3094 PAD.n2823 VSS 0.036454f
C3095 PAD.n2825 VSS 0.036454f
C3096 PAD.n2827 VSS 0.036454f
C3097 PAD.n2828 VSS 0.036454f
C3098 PAD.n2829 VSS 0.023105f
C3099 PAD.n2830 VSS 0.033374f
C3100 PAD.n2831 VSS 0.062262f
C3101 PAD.n2832 VSS 0.069752f
C3102 PAD.n2833 VSS 0.069752f
C3103 PAD.n2834 VSS 0.078918f
C3104 PAD.n2876 VSS 0.023105f
C3105 PAD.n2877 VSS 0.023105f
C3106 PAD.n2878 VSS 0.029431f
C3107 PAD.n2879 VSS 0.12331f
C3108 PAD.n2880 VSS 0.036454f
C3109 PAD.n2881 VSS 0.036454f
C3110 PAD.n2882 VSS 0.03428f
C3111 PAD.n2883 VSS 0.029431f
C3112 PAD.n2884 VSS 0.069752f
C3113 PAD.n2885 VSS 0.039754f
C3114 PAD.n2886 VSS 0.069752f
C3115 PAD.n2887 VSS 0.039754f
C3116 PAD.n2888 VSS 0.046278f
C3117 PAD.n2889 VSS 0.039754f
C3118 PAD.n2890 VSS 0.039754f
C3119 PAD.n2891 VSS 0.300877f
C3120 PAD.n2892 VSS 0.700403f
C3121 PAD.n2893 VSS 0.029913f
C3122 PAD.n2894 VSS 0.567228f
C3123 PAD.n2895 VSS 0.03925f
C3124 PAD.n2896 VSS 0.029913f
C3125 PAD.n2897 VSS 0.03925f
C3126 PAD.n2898 VSS 0.03055f
C3127 PAD.n2899 VSS 0.042887f
C3128 PAD.n2900 VSS 0.049106f
C3129 PAD.n2901 VSS 0.029431f
C3130 PAD.n2902 VSS 0.049106f
C3131 PAD.n2903 VSS 0.029431f
C3132 PAD.n2904 VSS 0.700403f
C3133 PAD.n2946 VSS 0.498174f
C3134 PAD.n2947 VSS 0.069752f
C3135 PAD.n2948 VSS 0.069752f
C3136 PAD.n2949 VSS 0.046278f
C3137 PAD.n2950 VSS 0.039754f
C3138 PAD.n2951 VSS 0.039754f
C3139 PAD.n2952 VSS 0.355133f
C3140 PAD.n2994 VSS 0.023105f
C3141 PAD.n2995 VSS 0.023105f
C3142 PAD.n2996 VSS 0.029431f
C3143 PAD.n2997 VSS 0.61162f
C3144 PAD.n2998 VSS 0.036454f
C3145 PAD.n2999 VSS 0.036454f
C3146 PAD.n3000 VSS 0.036454f
C3147 PAD.n3001 VSS 0.036454f
C3148 PAD.n3002 VSS 0.036454f
C3149 PAD.n3003 VSS 0.036454f
C3150 PAD.n3004 VSS 0.036454f
C3151 PAD.n3005 VSS 0.036454f
C3152 PAD.n3006 VSS 0.036454f
C3153 PAD.n3007 VSS 0.036454f
C3154 PAD.n3008 VSS 0.036454f
C3155 PAD.n3009 VSS 0.036454f
C3156 PAD.n3010 VSS 0.036454f
C3157 PAD.n3011 VSS 0.036454f
C3158 PAD.n3012 VSS 0.036454f
C3159 PAD.n3013 VSS 0.036454f
C3160 PAD.n3014 VSS 0.036454f
C3161 PAD.n3015 VSS 0.036454f
C3162 PAD.n3016 VSS 0.036454f
C3163 PAD.n3017 VSS 0.036454f
C3164 PAD.n3018 VSS 0.036454f
C3165 PAD.n3019 VSS 0.036454f
C3166 PAD.n3020 VSS 0.036454f
C3167 PAD.n3021 VSS 0.036454f
C3168 PAD.n3022 VSS 0.036454f
C3169 PAD.n3023 VSS 0.036454f
C3170 PAD.n3024 VSS 0.036454f
C3171 PAD.n3025 VSS 0.036454f
C3172 PAD.n3026 VSS 0.036454f
C3173 PAD.n3027 VSS 0.036454f
C3174 PAD.n3028 VSS 0.036454f
C3175 PAD.n3029 VSS 0.036454f
C3176 PAD.n3030 VSS 0.036454f
C3177 PAD.n3031 VSS 0.036454f
C3178 PAD.n3032 VSS 0.036454f
C3179 PAD.n3033 VSS 0.036454f
C3180 PAD.n3034 VSS 0.036454f
C3181 PAD.n3035 VSS 0.036454f
C3182 PAD.n3036 VSS 0.036454f
C3183 PAD.n3037 VSS 0.036454f
C3184 PAD.n3039 VSS 0.036454f
C3185 PAD.n3040 VSS 0.036454f
C3186 PAD.n3041 VSS 0.023105f
C3187 PAD.n3042 VSS 0.033374f
C3188 PAD.n3043 VSS 0.036454f
C3189 PAD.n3044 VSS 0.036454f
C3190 PAD.n3045 VSS 0.036454f
C3191 PAD.n3046 VSS 0.036454f
C3192 PAD.n3048 VSS 0.036454f
C3193 PAD.n3049 VSS 0.036454f
C3194 PAD.n3050 VSS 0.036454f
C3195 PAD.n3052 VSS 0.036454f
C3196 PAD.n3053 VSS 0.036454f
C3197 PAD.n3054 VSS 0.036454f
C3198 PAD.n3055 VSS 0.036454f
C3199 PAD.n3056 VSS 0.036454f
C3200 PAD.n3057 VSS 0.036454f
C3201 PAD.n3058 VSS 0.036454f
C3202 PAD.n3060 VSS 0.036454f
C3203 PAD.n3061 VSS 0.036454f
C3204 PAD.n3062 VSS 0.036454f
C3205 PAD.n3064 VSS 0.036454f
C3206 PAD.n3065 VSS 0.036454f
C3207 PAD.n3066 VSS 0.036454f
C3208 PAD.n3067 VSS 0.036454f
C3209 PAD.n3068 VSS 0.036454f
C3210 PAD.n3069 VSS 0.036454f
C3211 PAD.n3070 VSS 0.036454f
C3212 PAD.n3072 VSS 0.036454f
C3213 PAD.n3073 VSS 0.036454f
C3214 PAD.n3074 VSS 0.036454f
C3215 PAD.n3076 VSS 0.036454f
C3216 PAD.n3077 VSS 0.036454f
C3217 PAD.n3078 VSS 0.036454f
C3218 PAD.n3079 VSS 0.036454f
C3219 PAD.n3080 VSS 0.036454f
C3220 PAD.n3081 VSS 0.036454f
C3221 PAD.n3082 VSS 0.036454f
C3222 PAD.n3084 VSS 0.036454f
C3223 PAD.n3085 VSS 0.036454f
C3224 PAD.n3086 VSS 0.036454f
C3225 PAD.n3088 VSS 0.036454f
C3226 PAD.n3089 VSS 0.036454f
C3227 PAD.n3090 VSS 0.036454f
C3228 PAD.n3091 VSS 0.036454f
C3229 PAD.n3092 VSS 0.036454f
C3230 PAD.n3093 VSS 0.036454f
C3231 PAD.n3094 VSS 0.036454f
C3232 PAD.n3096 VSS 0.036454f
C3233 PAD.n3097 VSS 0.036454f
C3234 PAD.n3098 VSS 0.036454f
C3235 PAD.n3100 VSS 0.036454f
C3236 PAD.n3101 VSS 0.036454f
C3237 PAD.n3102 VSS 0.036454f
C3238 PAD.n3103 VSS 0.036454f
C3239 PAD.n3104 VSS 0.036454f
C3240 PAD.n3105 VSS 0.036454f
C3241 PAD.n3106 VSS 0.036454f
C3242 PAD.n3108 VSS 0.036454f
C3243 PAD.n3109 VSS 0.036454f
C3244 PAD.n3110 VSS 0.036454f
C3245 PAD.n3112 VSS 0.036454f
C3246 PAD.n3113 VSS 0.036454f
C3247 PAD.n3114 VSS 0.036454f
C3248 PAD.n3115 VSS 0.036454f
C3249 PAD.n3116 VSS 0.036454f
C3250 PAD.n3117 VSS 0.036454f
C3251 PAD.n3118 VSS 0.036454f
C3252 PAD.n3120 VSS 0.036454f
C3253 PAD.n3121 VSS 0.036454f
C3254 PAD.n3122 VSS 0.036454f
C3255 PAD.n3124 VSS 0.036454f
C3256 PAD.n3125 VSS 0.036454f
C3257 PAD.n3126 VSS 0.036454f
C3258 PAD.n3127 VSS 0.036454f
C3259 PAD.n3128 VSS 0.036454f
C3260 PAD.n3129 VSS 0.036454f
C3261 PAD.n3130 VSS 0.036454f
C3262 PAD.n3132 VSS 0.036454f
C3263 PAD.n3133 VSS 0.036454f
C3264 PAD.n3134 VSS 0.036454f
C3265 PAD.n3136 VSS 0.036454f
C3266 PAD.n3137 VSS 0.036454f
C3267 PAD.n3138 VSS 0.036454f
C3268 PAD.n3139 VSS 0.036454f
C3269 PAD.n3140 VSS 0.036454f
C3270 PAD.n3141 VSS 0.036454f
C3271 PAD.n3142 VSS 0.036454f
C3272 PAD.n3144 VSS 0.036454f
C3273 PAD.n3145 VSS 0.036454f
C3274 PAD.n3146 VSS 0.036454f
C3275 PAD.n3148 VSS 0.036454f
C3276 PAD.n3149 VSS 0.036454f
C3277 PAD.n3150 VSS 0.036454f
C3278 PAD.n3151 VSS 0.036454f
C3279 PAD.n3152 VSS 0.036454f
C3280 PAD.n3153 VSS 0.036454f
C3281 PAD.n3154 VSS 0.036454f
C3282 PAD.n3156 VSS 0.036454f
C3283 PAD.n3157 VSS 0.036454f
C3284 PAD.n3158 VSS 0.036454f
C3285 PAD.n3160 VSS 0.036454f
C3286 PAD.n3161 VSS 0.036454f
C3287 PAD.n3162 VSS 0.036454f
C3288 PAD.n3163 VSS 0.036454f
C3289 PAD.n3164 VSS 0.036454f
C3290 PAD.n3165 VSS 0.036454f
C3291 PAD.n3166 VSS 0.036454f
C3292 PAD.n3168 VSS 0.036454f
C3293 PAD.n3169 VSS 0.036454f
C3294 PAD.n3170 VSS 0.036454f
C3295 PAD.n3172 VSS 0.036454f
C3296 PAD.n3173 VSS 0.036454f
C3297 PAD.n3174 VSS 0.036454f
C3298 PAD.n3175 VSS 0.036454f
C3299 PAD.n3176 VSS 0.036454f
C3300 PAD.n3177 VSS 0.036454f
C3301 PAD.n3178 VSS 0.036454f
C3302 PAD.n3180 VSS 0.036454f
C3303 PAD.n3181 VSS 0.036454f
C3304 PAD.n3182 VSS 0.036454f
C3305 PAD.n3184 VSS 0.036454f
C3306 PAD.n3185 VSS 0.036454f
C3307 PAD.n3186 VSS 0.036454f
C3308 PAD.n3187 VSS 0.036454f
C3309 PAD.n3188 VSS 0.036454f
C3310 PAD.n3189 VSS 0.036454f
C3311 PAD.n3190 VSS 0.036454f
C3312 PAD.n3192 VSS 0.036454f
C3313 PAD.n3193 VSS 0.036454f
C3314 PAD.n3194 VSS 0.036454f
C3315 PAD.n3196 VSS 0.036454f
C3316 PAD.n3197 VSS 0.036454f
C3317 PAD.n3198 VSS 0.036454f
C3318 PAD.n3199 VSS 0.036454f
C3319 PAD.n3200 VSS 0.036454f
C3320 PAD.n3201 VSS 0.036454f
C3321 PAD.n3202 VSS 0.036454f
C3322 PAD.n3204 VSS 0.036454f
C3323 PAD.n3205 VSS 0.036454f
C3324 PAD.n3206 VSS 0.036454f
C3325 PAD.n3208 VSS 0.036454f
C3326 PAD.n3209 VSS 0.036454f
C3327 PAD.n3210 VSS 0.036454f
C3328 PAD.n3211 VSS 0.036454f
C3329 PAD.n3212 VSS 0.036454f
C3330 PAD.n3213 VSS 0.036454f
C3331 PAD.n3214 VSS 0.036454f
C3332 PAD.n3216 VSS 0.036454f
C3333 PAD.n3217 VSS 0.036454f
C3334 PAD.n3218 VSS 0.036454f
C3335 PAD.n3220 VSS 0.036454f
C3336 PAD.n3221 VSS 0.036454f
C3337 PAD.n3222 VSS 0.036454f
C3338 PAD.n3223 VSS 0.036454f
C3339 PAD.n3224 VSS 0.036454f
C3340 PAD.n3225 VSS 0.036454f
C3341 PAD.n3226 VSS 0.036454f
C3342 PAD.n3228 VSS 0.036454f
C3343 PAD.n3229 VSS 0.036454f
C3344 PAD.n3230 VSS 0.036454f
C3345 PAD.n3232 VSS 0.036454f
C3346 PAD.n3233 VSS 0.036454f
C3347 PAD.n3234 VSS 0.036454f
C3348 PAD.n3235 VSS 0.036454f
C3349 PAD.n3236 VSS 0.036454f
C3350 PAD.n3237 VSS 0.036454f
C3351 PAD.n3238 VSS 0.036454f
C3352 PAD.n3240 VSS 0.036454f
C3353 PAD.n3241 VSS 0.036454f
C3354 PAD.n3242 VSS 0.036454f
C3355 PAD.n3244 VSS 0.036454f
C3356 PAD.n3245 VSS 0.036454f
C3357 PAD.n3246 VSS 0.036454f
C3358 PAD.n3247 VSS 0.036454f
C3359 PAD.n3248 VSS 0.036454f
C3360 PAD.n3249 VSS 0.036454f
C3361 PAD.n3250 VSS 0.036454f
C3362 PAD.n3252 VSS 0.036454f
C3363 PAD.n3253 VSS 0.036454f
C3364 PAD.n3254 VSS 0.036454f
C3365 PAD.n3256 VSS 0.036454f
C3366 PAD.n3257 VSS 0.036454f
C3367 PAD.n3258 VSS 0.036454f
C3368 PAD.n3259 VSS 0.036454f
C3369 PAD.n3260 VSS 0.036454f
C3370 PAD.n3261 VSS 0.036454f
C3371 PAD.n3262 VSS 0.036454f
C3372 PAD.n3264 VSS 0.036454f
C3373 PAD.n3265 VSS 0.036454f
C3374 PAD.n3266 VSS 0.036454f
C3375 PAD.n3268 VSS 0.036454f
C3376 PAD.n3269 VSS 0.036454f
C3377 PAD.n3270 VSS 0.036454f
C3378 PAD.n3271 VSS 0.036454f
C3379 PAD.n3272 VSS 0.036454f
C3380 PAD.n3273 VSS 0.036454f
C3381 PAD.n3274 VSS 0.036454f
C3382 PAD.n3276 VSS 0.036454f
C3383 PAD.n3277 VSS 0.036454f
C3384 PAD.n3278 VSS 0.036454f
C3385 PAD.n3280 VSS 0.036454f
C3386 PAD.n3281 VSS 0.036454f
C3387 PAD.n3282 VSS 0.036454f
C3388 PAD.n3283 VSS 0.036454f
C3389 PAD.n3284 VSS 0.042132f
C3390 PAD.n3285 VSS 0.045475f
C3391 PAD.n3286 VSS 0.045475f
C3392 PAD.n3287 VSS 0.700403f
C3393 PAD.n3288 VSS 0.069752f
C3394 PAD.n3289 VSS 0.389661f
C3395 PAD.n3290 VSS 0.036001f
C3396 PAD.n3291 VSS 0.069752f
C3397 PAD.n3292 VSS 0.036001f
C3398 PAD.n3293 VSS 0.046278f
C3399 PAD.n3294 VSS 0.039754f
C3400 PAD.n3295 VSS 0.039754f
C3401 PAD.n3296 VSS 0.498174f
C3402 PAD.n3338 VSS 0.023105f
C3403 PAD.n3339 VSS 0.40939f
C3404 PAD.n3340 VSS 0.023105f
C3405 PAD.n3341 VSS 0.029431f
C3406 PAD.n3342 VSS 0.389661f
C3407 PAD.n3343 VSS 0.036454f
C3408 PAD.n3344 VSS 0.036454f
C3409 PAD.n3345 VSS 0.036454f
C3410 PAD.n3346 VSS 0.036454f
C3411 PAD.n3347 VSS 0.036454f
C3412 PAD.n3348 VSS 0.036454f
C3413 PAD.n3349 VSS 0.036454f
C3414 PAD.n3350 VSS 0.036454f
C3415 PAD.n3351 VSS 0.036454f
C3416 PAD.n3352 VSS 0.036454f
C3417 PAD.n3353 VSS 0.036454f
C3418 PAD.n3354 VSS 0.036454f
C3419 PAD.n3355 VSS 0.036454f
C3420 PAD.n3356 VSS 0.036454f
C3421 PAD.n3357 VSS 0.036454f
C3422 PAD.n3358 VSS 0.036454f
C3423 PAD.n3359 VSS 0.036454f
C3424 PAD.n3360 VSS 0.036454f
C3425 PAD.n3361 VSS 0.036454f
C3426 PAD.n3362 VSS 0.036454f
C3427 PAD.n3363 VSS 0.036454f
C3428 PAD.n3364 VSS 0.036454f
C3429 PAD.n3365 VSS 0.036454f
C3430 PAD.n3366 VSS 0.036454f
C3431 PAD.n3367 VSS 0.036454f
C3432 PAD.n3368 VSS 0.036454f
C3433 PAD.n3369 VSS 0.036454f
C3434 PAD.n3370 VSS 0.036454f
C3435 PAD.n3371 VSS 0.036454f
C3436 PAD.n3372 VSS 0.036454f
C3437 PAD.n3373 VSS 0.036454f
C3438 PAD.n3374 VSS 0.036454f
C3439 PAD.n3375 VSS 0.036454f
C3440 PAD.n3376 VSS 0.036454f
C3441 PAD.n3377 VSS 0.036454f
C3442 PAD.n3378 VSS 0.036454f
C3443 PAD.n3379 VSS 0.036454f
C3444 PAD.n3380 VSS 0.036454f
C3445 PAD.n3381 VSS 0.036454f
C3446 PAD.n3382 VSS 0.036454f
C3447 PAD.n3384 VSS 0.036454f
C3448 PAD.n3385 VSS 0.036454f
C3449 PAD.n3386 VSS 0.023105f
C3450 PAD.n3387 VSS 0.033374f
C3451 PAD.n3388 VSS 0.036454f
C3452 PAD.n3389 VSS 0.036454f
C3453 PAD.n3390 VSS 0.036454f
C3454 PAD.n3391 VSS 0.036454f
C3455 PAD.n3393 VSS 0.036454f
C3456 PAD.n3394 VSS 0.036454f
C3457 PAD.n3395 VSS 0.036454f
C3458 PAD.n3397 VSS 0.036454f
C3459 PAD.n3398 VSS 0.036454f
C3460 PAD.n3399 VSS 0.036454f
C3461 PAD.n3400 VSS 0.036454f
C3462 PAD.n3401 VSS 0.036454f
C3463 PAD.n3402 VSS 0.036454f
C3464 PAD.n3403 VSS 0.036454f
C3465 PAD.n3405 VSS 0.036454f
C3466 PAD.n3406 VSS 0.036454f
C3467 PAD.n3407 VSS 0.036454f
C3468 PAD.n3409 VSS 0.036454f
C3469 PAD.n3410 VSS 0.036454f
C3470 PAD.n3411 VSS 0.036454f
C3471 PAD.n3412 VSS 0.036454f
C3472 PAD.n3413 VSS 0.036454f
C3473 PAD.n3414 VSS 0.036454f
C3474 PAD.n3415 VSS 0.036454f
C3475 PAD.n3417 VSS 0.036454f
C3476 PAD.n3418 VSS 0.036454f
C3477 PAD.n3419 VSS 0.036454f
C3478 PAD.n3421 VSS 0.036454f
C3479 PAD.n3422 VSS 0.036454f
C3480 PAD.n3423 VSS 0.036454f
C3481 PAD.n3424 VSS 0.036454f
C3482 PAD.n3425 VSS 0.036454f
C3483 PAD.n3426 VSS 0.036454f
C3484 PAD.n3427 VSS 0.036454f
C3485 PAD.n3429 VSS 0.036454f
C3486 PAD.n3430 VSS 0.036454f
C3487 PAD.n3431 VSS 0.036454f
C3488 PAD.n3433 VSS 0.036454f
C3489 PAD.n3434 VSS 0.036454f
C3490 PAD.n3435 VSS 0.036454f
C3491 PAD.n3436 VSS 0.036454f
C3492 PAD.n3437 VSS 0.036454f
C3493 PAD.n3438 VSS 0.036454f
C3494 PAD.n3439 VSS 0.036454f
C3495 PAD.n3441 VSS 0.036454f
C3496 PAD.n3442 VSS 0.036454f
C3497 PAD.n3443 VSS 0.036454f
C3498 PAD.n3445 VSS 0.036454f
C3499 PAD.n3446 VSS 0.036454f
C3500 PAD.n3447 VSS 0.036454f
C3501 PAD.n3448 VSS 0.036454f
C3502 PAD.n3449 VSS 0.036454f
C3503 PAD.n3450 VSS 0.036454f
C3504 PAD.n3451 VSS 0.036454f
C3505 PAD.n3453 VSS 0.036454f
C3506 PAD.n3454 VSS 0.036454f
C3507 PAD.n3455 VSS 0.036454f
C3508 PAD.n3457 VSS 0.036454f
C3509 PAD.n3458 VSS 0.036454f
C3510 PAD.n3459 VSS 0.036454f
C3511 PAD.n3460 VSS 0.036454f
C3512 PAD.n3461 VSS 0.036454f
C3513 PAD.n3462 VSS 0.036454f
C3514 PAD.n3463 VSS 0.036454f
C3515 PAD.n3465 VSS 0.036454f
C3516 PAD.n3466 VSS 0.036454f
C3517 PAD.n3467 VSS 0.036454f
C3518 PAD.n3469 VSS 0.036454f
C3519 PAD.n3470 VSS 0.036454f
C3520 PAD.n3471 VSS 0.036454f
C3521 PAD.n3472 VSS 0.036454f
C3522 PAD.n3473 VSS 0.036454f
C3523 PAD.n3474 VSS 0.036454f
C3524 PAD.n3475 VSS 0.036454f
C3525 PAD.n3477 VSS 0.036454f
C3526 PAD.n3478 VSS 0.036454f
C3527 PAD.n3479 VSS 0.036454f
C3528 PAD.n3481 VSS 0.036454f
C3529 PAD.n3482 VSS 0.036454f
C3530 PAD.n3483 VSS 0.036454f
C3531 PAD.n3484 VSS 0.036454f
C3532 PAD.n3485 VSS 0.036454f
C3533 PAD.n3486 VSS 0.036454f
C3534 PAD.n3487 VSS 0.036454f
C3535 PAD.n3489 VSS 0.036454f
C3536 PAD.n3490 VSS 0.036454f
C3537 PAD.n3491 VSS 0.036454f
C3538 PAD.n3493 VSS 0.036454f
C3539 PAD.n3494 VSS 0.036454f
C3540 PAD.n3495 VSS 0.036454f
C3541 PAD.n3496 VSS 0.036454f
C3542 PAD.n3497 VSS 0.036454f
C3543 PAD.n3498 VSS 0.036454f
C3544 PAD.n3499 VSS 0.036454f
C3545 PAD.n3501 VSS 0.036454f
C3546 PAD.n3502 VSS 0.036454f
C3547 PAD.n3503 VSS 0.036454f
C3548 PAD.n3505 VSS 0.036454f
C3549 PAD.n3506 VSS 0.036454f
C3550 PAD.n3507 VSS 0.036454f
C3551 PAD.n3508 VSS 0.036454f
C3552 PAD.n3509 VSS 0.036454f
C3553 PAD.n3510 VSS 0.036454f
C3554 PAD.n3511 VSS 0.036454f
C3555 PAD.n3513 VSS 0.036454f
C3556 PAD.n3514 VSS 0.036454f
C3557 PAD.n3515 VSS 0.036454f
C3558 PAD.n3517 VSS 0.036454f
C3559 PAD.n3518 VSS 0.036454f
C3560 PAD.n3519 VSS 0.036454f
C3561 PAD.n3520 VSS 0.036454f
C3562 PAD.n3521 VSS 0.036454f
C3563 PAD.n3522 VSS 0.036454f
C3564 PAD.n3523 VSS 0.036454f
C3565 PAD.n3525 VSS 0.036454f
C3566 PAD.n3526 VSS 0.036454f
C3567 PAD.n3527 VSS 0.036454f
C3568 PAD.n3529 VSS 0.036454f
C3569 PAD.n3530 VSS 0.036454f
C3570 PAD.n3531 VSS 0.036454f
C3571 PAD.n3532 VSS 0.036454f
C3572 PAD.n3533 VSS 0.036454f
C3573 PAD.n3534 VSS 0.036454f
C3574 PAD.n3535 VSS 0.036454f
C3575 PAD.n3537 VSS 0.036454f
C3576 PAD.n3538 VSS 0.036454f
C3577 PAD.n3539 VSS 0.036454f
C3578 PAD.n3541 VSS 0.036454f
C3579 PAD.n3542 VSS 0.036454f
C3580 PAD.n3543 VSS 0.036454f
C3581 PAD.n3544 VSS 0.036454f
C3582 PAD.n3545 VSS 0.036454f
C3583 PAD.n3546 VSS 0.036454f
C3584 PAD.n3547 VSS 0.036454f
C3585 PAD.n3549 VSS 0.036454f
C3586 PAD.n3550 VSS 0.036454f
C3587 PAD.n3551 VSS 0.036454f
C3588 PAD.n3553 VSS 0.036454f
C3589 PAD.n3554 VSS 0.036454f
C3590 PAD.n3555 VSS 0.036454f
C3591 PAD.n3556 VSS 0.036454f
C3592 PAD.n3557 VSS 0.036454f
C3593 PAD.n3558 VSS 0.036454f
C3594 PAD.n3559 VSS 0.036454f
C3595 PAD.n3561 VSS 0.036454f
C3596 PAD.n3562 VSS 0.036454f
C3597 PAD.n3563 VSS 0.036454f
C3598 PAD.n3565 VSS 0.036454f
C3599 PAD.n3566 VSS 0.036454f
C3600 PAD.n3567 VSS 0.036454f
C3601 PAD.n3568 VSS 0.036454f
C3602 PAD.n3569 VSS 0.036454f
C3603 PAD.n3570 VSS 0.036454f
C3604 PAD.n3571 VSS 0.036454f
C3605 PAD.n3573 VSS 0.036454f
C3606 PAD.n3574 VSS 0.036454f
C3607 PAD.n3575 VSS 0.036454f
C3608 PAD.n3577 VSS 0.036454f
C3609 PAD.n3578 VSS 0.036454f
C3610 PAD.n3579 VSS 0.036454f
C3611 PAD.n3580 VSS 0.036454f
C3612 PAD.n3581 VSS 0.036454f
C3613 PAD.n3582 VSS 0.036454f
C3614 PAD.n3583 VSS 0.036454f
C3615 PAD.n3585 VSS 0.036454f
C3616 PAD.n3586 VSS 0.036454f
C3617 PAD.n3587 VSS 0.036454f
C3618 PAD.n3589 VSS 0.036454f
C3619 PAD.n3590 VSS 0.036454f
C3620 PAD.n3591 VSS 0.036454f
C3621 PAD.n3592 VSS 0.036454f
C3622 PAD.n3593 VSS 0.036454f
C3623 PAD.n3594 VSS 0.036454f
C3624 PAD.n3595 VSS 0.036454f
C3625 PAD.n3597 VSS 0.036454f
C3626 PAD.n3598 VSS 0.036454f
C3627 PAD.n3599 VSS 0.036454f
C3628 PAD.n3601 VSS 0.036454f
C3629 PAD.n3602 VSS 0.036454f
C3630 PAD.n3603 VSS 0.036454f
C3631 PAD.n3604 VSS 0.036454f
C3632 PAD.n3605 VSS 0.036454f
C3633 PAD.n3606 VSS 0.036454f
C3634 PAD.n3607 VSS 0.036454f
C3635 PAD.n3609 VSS 0.036454f
C3636 PAD.n3610 VSS 0.036454f
C3637 PAD.n3611 VSS 0.036454f
C3638 PAD.n3613 VSS 0.036454f
C3639 PAD.n3614 VSS 0.036454f
C3640 PAD.n3615 VSS 0.036454f
C3641 PAD.n3616 VSS 0.036454f
C3642 PAD.n3617 VSS 0.036454f
C3643 PAD.n3618 VSS 0.036454f
C3644 PAD.n3619 VSS 0.036454f
C3645 PAD.n3621 VSS 0.036454f
C3646 PAD.n3622 VSS 0.036454f
C3647 PAD.n3623 VSS 0.036454f
C3648 PAD.n3625 VSS 0.036454f
C3649 PAD.n3626 VSS 0.036454f
C3650 PAD.n3627 VSS 0.036454f
C3651 PAD.n3628 VSS 0.036454f
C3652 PAD.n3629 VSS 0.042887f
C3653 PAD.n3630 VSS 0.049106f
C3654 PAD.n3631 VSS 0.029431f
C3655 PAD.n3632 VSS 0.040979f
C3656 PAD.n3633 VSS 0.700403f
C3657 PAD.n3634 VSS 0.069752f
C3658 PAD.n3635 VSS 0.069752f
C3659 PAD.n3636 VSS 12.7067f
C3660 PAD.n3637 VSS 14.5091f
C3661 PAD.n3638 VSS 0.046278f
C3662 PAD.n3639 VSS 0.039754f
C3663 PAD.n3640 VSS 0.039754f
C3664 PAD.n3641 VSS 0.606687f
C3665 PAD.n3683 VSS 0.023105f
C3666 PAD.n3684 VSS 0.517904f
C3667 PAD.n3685 VSS 0.023105f
C3668 PAD.n3686 VSS 0.029431f
C3669 PAD.n3687 VSS 0.12331f
C3670 PAD.n3688 VSS 0.036454f
C3671 PAD.n3689 VSS 0.036454f
C3672 PAD.n3690 VSS 0.036454f
C3673 PAD.n3691 VSS 0.036454f
C3674 PAD.n3692 VSS 0.036454f
C3675 PAD.n3693 VSS 0.036454f
C3676 PAD.n3694 VSS 0.036454f
C3677 PAD.n3695 VSS 0.036454f
C3678 PAD.n3696 VSS 0.036454f
C3679 PAD.n3697 VSS 0.036454f
C3680 PAD.n3698 VSS 0.036454f
C3681 PAD.n3699 VSS 0.036454f
C3682 PAD.n3700 VSS 0.036454f
C3683 PAD.n3701 VSS 0.036454f
C3684 PAD.n3702 VSS 0.036454f
C3685 PAD.n3703 VSS 0.036454f
C3686 PAD.n3704 VSS 0.036454f
C3687 PAD.n3705 VSS 0.036454f
C3688 PAD.n3706 VSS 0.036454f
C3689 PAD.n3707 VSS 0.036454f
C3690 PAD.n3708 VSS 0.036454f
C3691 PAD.n3709 VSS 0.036454f
C3692 PAD.n3710 VSS 0.036454f
C3693 PAD.n3711 VSS 0.036454f
C3694 PAD.n3712 VSS 0.036454f
C3695 PAD.n3713 VSS 0.036454f
C3696 PAD.n3714 VSS 0.036454f
C3697 PAD.n3715 VSS 0.036454f
C3698 PAD.n3716 VSS 0.036454f
C3699 PAD.n3717 VSS 0.036454f
C3700 PAD.n3718 VSS 0.036454f
C3701 PAD.n3719 VSS 0.036454f
C3702 PAD.n3720 VSS 0.036454f
C3703 PAD.n3721 VSS 0.036454f
C3704 PAD.n3722 VSS 0.036454f
C3705 PAD.n3723 VSS 0.036454f
C3706 PAD.n3724 VSS 0.036454f
C3707 PAD.n3725 VSS 0.036454f
C3708 PAD.n3726 VSS 0.036454f
C3709 PAD.n3727 VSS 0.036454f
C3710 PAD.n3729 VSS 0.036454f
C3711 PAD.n3730 VSS 0.036454f
C3712 PAD.n3731 VSS 0.023105f
C3713 PAD.n3732 VSS 0.033374f
C3714 PAD.n3733 VSS 0.036454f
C3715 PAD.n3734 VSS 0.036454f
C3716 PAD.n3735 VSS 0.036454f
C3717 PAD.n3736 VSS 0.036454f
C3718 PAD.n3738 VSS 0.036454f
C3719 PAD.n3739 VSS 0.036454f
C3720 PAD.n3740 VSS 0.036454f
C3721 PAD.n3742 VSS 0.036454f
C3722 PAD.n3743 VSS 0.036454f
C3723 PAD.n3744 VSS 0.036454f
C3724 PAD.n3745 VSS 0.036454f
C3725 PAD.n3746 VSS 0.036454f
C3726 PAD.n3747 VSS 0.036454f
C3727 PAD.n3748 VSS 0.036454f
C3728 PAD.n3750 VSS 0.036454f
C3729 PAD.n3751 VSS 0.036454f
C3730 PAD.n3752 VSS 0.036454f
C3731 PAD.n3754 VSS 0.036454f
C3732 PAD.n3755 VSS 0.036454f
C3733 PAD.n3756 VSS 0.036454f
C3734 PAD.n3757 VSS 0.036454f
C3735 PAD.n3758 VSS 0.036454f
C3736 PAD.n3759 VSS 0.036454f
C3737 PAD.n3760 VSS 0.036454f
C3738 PAD.n3762 VSS 0.036454f
C3739 PAD.n3763 VSS 0.036454f
C3740 PAD.n3764 VSS 0.036454f
C3741 PAD.n3766 VSS 0.036454f
C3742 PAD.n3767 VSS 0.036454f
C3743 PAD.n3768 VSS 0.036454f
C3744 PAD.n3769 VSS 0.036454f
C3745 PAD.n3770 VSS 0.036454f
C3746 PAD.n3771 VSS 0.036454f
C3747 PAD.n3772 VSS 0.036454f
C3748 PAD.n3774 VSS 0.036454f
C3749 PAD.n3775 VSS 0.036454f
C3750 PAD.n3776 VSS 0.036454f
C3751 PAD.n3778 VSS 0.036454f
C3752 PAD.n3779 VSS 0.036454f
C3753 PAD.n3780 VSS 0.036454f
C3754 PAD.n3781 VSS 0.036454f
C3755 PAD.n3782 VSS 0.036454f
C3756 PAD.n3783 VSS 0.036454f
C3757 PAD.n3784 VSS 0.036454f
C3758 PAD.n3786 VSS 0.036454f
C3759 PAD.n3787 VSS 0.036454f
C3760 PAD.n3788 VSS 0.036454f
C3761 PAD.n3790 VSS 0.036454f
C3762 PAD.n3791 VSS 0.036454f
C3763 PAD.n3792 VSS 0.036454f
C3764 PAD.n3793 VSS 0.036454f
C3765 PAD.n3794 VSS 0.036454f
C3766 PAD.n3795 VSS 0.036454f
C3767 PAD.n3796 VSS 0.036454f
C3768 PAD.n3798 VSS 0.036454f
C3769 PAD.n3799 VSS 0.036454f
C3770 PAD.n3800 VSS 0.036454f
C3771 PAD.n3802 VSS 0.036454f
C3772 PAD.n3803 VSS 0.036454f
C3773 PAD.n3804 VSS 0.036454f
C3774 PAD.n3805 VSS 0.036454f
C3775 PAD.n3806 VSS 0.036454f
C3776 PAD.n3807 VSS 0.036454f
C3777 PAD.n3808 VSS 0.036454f
C3778 PAD.n3810 VSS 0.036454f
C3779 PAD.n3811 VSS 0.036454f
C3780 PAD.n3812 VSS 0.036454f
C3781 PAD.n3814 VSS 0.036454f
C3782 PAD.n3815 VSS 0.036454f
C3783 PAD.n3816 VSS 0.036454f
C3784 PAD.n3817 VSS 0.036454f
C3785 PAD.n3818 VSS 0.036454f
C3786 PAD.n3819 VSS 0.036454f
C3787 PAD.n3820 VSS 0.036454f
C3788 PAD.n3822 VSS 0.036454f
C3789 PAD.n3823 VSS 0.036454f
C3790 PAD.n3824 VSS 0.036454f
C3791 PAD.n3826 VSS 0.036454f
C3792 PAD.n3827 VSS 0.036454f
C3793 PAD.n3828 VSS 0.036454f
C3794 PAD.n3829 VSS 0.036454f
C3795 PAD.n3830 VSS 0.036454f
C3796 PAD.n3831 VSS 0.036454f
C3797 PAD.n3832 VSS 0.036454f
C3798 PAD.n3834 VSS 0.036454f
C3799 PAD.n3835 VSS 0.036454f
C3800 PAD.n3836 VSS 0.036454f
C3801 PAD.n3838 VSS 0.036454f
C3802 PAD.n3839 VSS 0.036454f
C3803 PAD.n3840 VSS 0.036454f
C3804 PAD.n3841 VSS 0.036454f
C3805 PAD.n3842 VSS 0.036454f
C3806 PAD.n3843 VSS 0.036454f
C3807 PAD.n3844 VSS 0.036454f
C3808 PAD.n3846 VSS 0.036454f
C3809 PAD.n3847 VSS 0.036454f
C3810 PAD.n3848 VSS 0.036454f
C3811 PAD.n3850 VSS 0.036454f
C3812 PAD.n3851 VSS 0.036454f
C3813 PAD.n3852 VSS 0.036454f
C3814 PAD.n3853 VSS 0.036454f
C3815 PAD.n3854 VSS 0.036454f
C3816 PAD.n3855 VSS 0.036454f
C3817 PAD.n3856 VSS 0.036454f
C3818 PAD.n3858 VSS 0.036454f
C3819 PAD.n3859 VSS 0.036454f
C3820 PAD.n3860 VSS 0.036454f
C3821 PAD.n3862 VSS 0.036454f
C3822 PAD.n3863 VSS 0.036454f
C3823 PAD.n3864 VSS 0.036454f
C3824 PAD.n3865 VSS 0.036454f
C3825 PAD.n3866 VSS 0.036454f
C3826 PAD.n3867 VSS 0.036454f
C3827 PAD.n3868 VSS 0.036454f
C3828 PAD.n3870 VSS 0.036454f
C3829 PAD.n3871 VSS 0.036454f
C3830 PAD.n3872 VSS 0.036454f
C3831 PAD.n3874 VSS 0.036454f
C3832 PAD.n3875 VSS 0.036454f
C3833 PAD.n3876 VSS 0.036454f
C3834 PAD.n3877 VSS 0.036454f
C3835 PAD.n3878 VSS 0.036454f
C3836 PAD.n3879 VSS 0.036454f
C3837 PAD.n3880 VSS 0.036454f
C3838 PAD.n3882 VSS 0.036454f
C3839 PAD.n3883 VSS 0.036454f
C3840 PAD.n3884 VSS 0.036454f
C3841 PAD.n3886 VSS 0.036454f
C3842 PAD.n3887 VSS 0.036454f
C3843 PAD.n3888 VSS 0.036454f
C3844 PAD.n3889 VSS 0.036454f
C3845 PAD.n3890 VSS 0.036454f
C3846 PAD.n3891 VSS 0.036454f
C3847 PAD.n3892 VSS 0.036454f
C3848 PAD.n3894 VSS 0.036454f
C3849 PAD.n3895 VSS 0.036454f
C3850 PAD.n3896 VSS 0.036454f
C3851 PAD.n3898 VSS 0.036454f
C3852 PAD.n3899 VSS 0.036454f
C3853 PAD.n3900 VSS 0.036454f
C3854 PAD.n3901 VSS 0.036454f
C3855 PAD.n3902 VSS 0.036454f
C3856 PAD.n3903 VSS 0.036454f
C3857 PAD.n3904 VSS 0.036454f
C3858 PAD.n3906 VSS 0.036454f
C3859 PAD.n3907 VSS 0.036454f
C3860 PAD.n3908 VSS 0.036454f
C3861 PAD.n3910 VSS 0.036454f
C3862 PAD.n3911 VSS 0.036454f
C3863 PAD.n3912 VSS 0.036454f
C3864 PAD.n3913 VSS 0.036454f
C3865 PAD.n3914 VSS 0.036454f
C3866 PAD.n3915 VSS 0.036454f
C3867 PAD.n3916 VSS 0.036454f
C3868 PAD.n3918 VSS 0.036454f
C3869 PAD.n3919 VSS 0.036454f
C3870 PAD.n3920 VSS 0.036454f
C3871 PAD.n3922 VSS 0.036454f
C3872 PAD.n3923 VSS 0.036454f
C3873 PAD.n3924 VSS 0.036454f
C3874 PAD.n3925 VSS 0.036454f
C3875 PAD.n3926 VSS 0.036454f
C3876 PAD.n3927 VSS 0.036454f
C3877 PAD.n3928 VSS 0.036454f
C3878 PAD.n3930 VSS 0.036454f
C3879 PAD.n3931 VSS 0.036454f
C3880 PAD.n3932 VSS 0.036454f
C3881 PAD.n3934 VSS 0.036454f
C3882 PAD.n3935 VSS 0.036454f
C3883 PAD.n3936 VSS 0.036454f
C3884 PAD.n3937 VSS 0.036454f
C3885 PAD.n3938 VSS 0.036454f
C3886 PAD.n3939 VSS 0.036454f
C3887 PAD.n3940 VSS 0.036454f
C3888 PAD.n3942 VSS 0.036454f
C3889 PAD.n3943 VSS 0.036454f
C3890 PAD.n3944 VSS 0.036454f
C3891 PAD.n3946 VSS 0.036454f
C3892 PAD.n3947 VSS 0.036454f
C3893 PAD.n3948 VSS 0.036454f
C3894 PAD.n3949 VSS 0.036454f
C3895 PAD.n3950 VSS 0.036454f
C3896 PAD.n3951 VSS 0.036454f
C3897 PAD.n3952 VSS 0.036454f
C3898 PAD.n3954 VSS 0.036454f
C3899 PAD.n3955 VSS 0.036454f
C3900 PAD.n3956 VSS 0.036454f
C3901 PAD.n3958 VSS 0.036454f
C3902 PAD.n3959 VSS 0.036454f
C3903 PAD.n3960 VSS 0.036454f
C3904 PAD.n3961 VSS 0.036454f
C3905 PAD.n3962 VSS 0.036454f
C3906 PAD.n3963 VSS 0.036454f
C3907 PAD.n3964 VSS 0.036454f
C3908 PAD.n3966 VSS 0.036454f
C3909 PAD.n3967 VSS 0.036454f
C3910 PAD.n3968 VSS 0.036454f
C3911 PAD.n3970 VSS 0.036454f
C3912 PAD.n3971 VSS 0.036454f
C3913 PAD.n3972 VSS 0.036454f
C3914 PAD.n3973 VSS 0.036454f
C3915 PAD.n3974 VSS 0.028541f
C3916 PAD.n3975 VSS 0.049106f
C3917 PAD.n3976 VSS 0.036484f
C3918 PAD.n3977 VSS 0.646146f
C3919 PAD.n3978 VSS 0.069752f
C3920 PAD.n3979 VSS 0.069752f
C3921 PAD.n3980 VSS 0.046278f
C3922 PAD.n3981 VSS 0.039754f
C3923 PAD.n3982 VSS 0.039754f
C3924 PAD.n3983 VSS 0.562295f
C3925 PAD.n4025 VSS 0.023105f
C3926 PAD.n4026 VSS 0.023105f
C3927 PAD.n4027 VSS 0.029431f
C3928 PAD.n4028 VSS 0.14304f
C3929 PAD.n4029 VSS 0.036454f
C3930 PAD.n4030 VSS 0.036454f
C3931 PAD.n4031 VSS 0.036454f
C3932 PAD.n4032 VSS 0.036454f
C3933 PAD.n4033 VSS 0.036454f
C3934 PAD.n4034 VSS 0.036454f
C3935 PAD.n4035 VSS 0.036454f
C3936 PAD.n4036 VSS 0.036454f
C3937 PAD.n4037 VSS 0.036454f
C3938 PAD.n4038 VSS 0.036454f
C3939 PAD.n4039 VSS 0.036454f
C3940 PAD.n4040 VSS 0.036454f
C3941 PAD.n4041 VSS 0.036454f
C3942 PAD.n4042 VSS 0.036454f
C3943 PAD.n4043 VSS 0.036454f
C3944 PAD.n4044 VSS 0.036454f
C3945 PAD.n4045 VSS 0.036454f
C3946 PAD.n4046 VSS 0.036454f
C3947 PAD.n4047 VSS 0.036454f
C3948 PAD.n4048 VSS 0.036454f
C3949 PAD.n4049 VSS 0.036454f
C3950 PAD.n4050 VSS 0.036454f
C3951 PAD.n4051 VSS 0.036454f
C3952 PAD.n4052 VSS 0.036454f
C3953 PAD.n4053 VSS 0.036454f
C3954 PAD.n4054 VSS 0.036454f
C3955 PAD.n4055 VSS 0.036454f
C3956 PAD.n4056 VSS 0.036454f
C3957 PAD.n4057 VSS 0.036454f
C3958 PAD.n4058 VSS 0.036454f
C3959 PAD.n4059 VSS 0.036454f
C3960 PAD.n4060 VSS 0.036454f
C3961 PAD.n4061 VSS 0.036454f
C3962 PAD.n4062 VSS 0.036454f
C3963 PAD.n4063 VSS 0.036454f
C3964 PAD.n4064 VSS 0.036454f
C3965 PAD.n4065 VSS 0.036454f
C3966 PAD.n4066 VSS 0.036454f
C3967 PAD.n4067 VSS 0.036454f
C3968 PAD.n4068 VSS 0.036454f
C3969 PAD.n4070 VSS 0.036454f
C3970 PAD.n4071 VSS 0.036454f
C3971 PAD.n4072 VSS 0.023105f
C3972 PAD.n4073 VSS 0.033374f
C3973 PAD.n4074 VSS 0.036454f
C3974 PAD.n4075 VSS 0.036454f
C3975 PAD.n4076 VSS 0.036454f
C3976 PAD.n4077 VSS 0.036454f
C3977 PAD.n4079 VSS 0.036454f
C3978 PAD.n4080 VSS 0.036454f
C3979 PAD.n4081 VSS 0.036454f
C3980 PAD.n4083 VSS 0.036454f
C3981 PAD.n4084 VSS 0.036454f
C3982 PAD.n4085 VSS 0.036454f
C3983 PAD.n4086 VSS 0.036454f
C3984 PAD.n4087 VSS 0.036454f
C3985 PAD.n4088 VSS 0.036454f
C3986 PAD.n4089 VSS 0.036454f
C3987 PAD.n4091 VSS 0.036454f
C3988 PAD.n4092 VSS 0.036454f
C3989 PAD.n4093 VSS 0.036454f
C3990 PAD.n4095 VSS 0.036454f
C3991 PAD.n4096 VSS 0.036454f
C3992 PAD.n4097 VSS 0.036454f
C3993 PAD.n4098 VSS 0.036454f
C3994 PAD.n4099 VSS 0.036454f
C3995 PAD.n4100 VSS 0.036454f
C3996 PAD.n4101 VSS 0.036454f
C3997 PAD.n4103 VSS 0.036454f
C3998 PAD.n4104 VSS 0.036454f
C3999 PAD.n4105 VSS 0.036454f
C4000 PAD.n4107 VSS 0.036454f
C4001 PAD.n4108 VSS 0.036454f
C4002 PAD.n4109 VSS 0.036454f
C4003 PAD.n4110 VSS 0.036454f
C4004 PAD.n4111 VSS 0.036454f
C4005 PAD.n4112 VSS 0.036454f
C4006 PAD.n4113 VSS 0.036454f
C4007 PAD.n4115 VSS 0.036454f
C4008 PAD.n4116 VSS 0.036454f
C4009 PAD.n4117 VSS 0.036454f
C4010 PAD.n4119 VSS 0.036454f
C4011 PAD.n4120 VSS 0.036454f
C4012 PAD.n4121 VSS 0.036454f
C4013 PAD.n4122 VSS 0.036454f
C4014 PAD.n4123 VSS 0.036454f
C4015 PAD.n4124 VSS 0.036454f
C4016 PAD.n4125 VSS 0.036454f
C4017 PAD.n4127 VSS 0.036454f
C4018 PAD.n4128 VSS 0.036454f
C4019 PAD.n4129 VSS 0.036454f
C4020 PAD.n4131 VSS 0.036454f
C4021 PAD.n4132 VSS 0.036454f
C4022 PAD.n4133 VSS 0.036454f
C4023 PAD.n4134 VSS 0.036454f
C4024 PAD.n4135 VSS 0.036454f
C4025 PAD.n4136 VSS 0.036454f
C4026 PAD.n4137 VSS 0.036454f
C4027 PAD.n4139 VSS 0.036454f
C4028 PAD.n4140 VSS 0.036454f
C4029 PAD.n4141 VSS 0.036454f
C4030 PAD.n4143 VSS 0.036454f
C4031 PAD.n4144 VSS 0.036454f
C4032 PAD.n4145 VSS 0.036454f
C4033 PAD.n4146 VSS 0.036454f
C4034 PAD.n4147 VSS 0.036454f
C4035 PAD.n4148 VSS 0.036454f
C4036 PAD.n4149 VSS 0.036454f
C4037 PAD.n4151 VSS 0.036454f
C4038 PAD.n4152 VSS 0.036454f
C4039 PAD.n4153 VSS 0.036454f
C4040 PAD.n4155 VSS 0.036454f
C4041 PAD.n4156 VSS 0.036454f
C4042 PAD.n4157 VSS 0.036454f
C4043 PAD.n4158 VSS 0.036454f
C4044 PAD.n4159 VSS 0.036454f
C4045 PAD.n4160 VSS 0.036454f
C4046 PAD.n4161 VSS 0.036454f
C4047 PAD.n4163 VSS 0.036454f
C4048 PAD.n4164 VSS 0.036454f
C4049 PAD.n4165 VSS 0.036454f
C4050 PAD.n4167 VSS 0.036454f
C4051 PAD.n4168 VSS 0.036454f
C4052 PAD.n4169 VSS 0.036454f
C4053 PAD.n4170 VSS 0.036454f
C4054 PAD.n4171 VSS 0.036454f
C4055 PAD.n4172 VSS 0.036454f
C4056 PAD.n4173 VSS 0.036454f
C4057 PAD.n4175 VSS 0.036454f
C4058 PAD.n4176 VSS 0.036454f
C4059 PAD.n4177 VSS 0.036454f
C4060 PAD.n4179 VSS 0.036454f
C4061 PAD.n4180 VSS 0.036454f
C4062 PAD.n4181 VSS 0.036454f
C4063 PAD.n4182 VSS 0.036454f
C4064 PAD.n4183 VSS 0.036454f
C4065 PAD.n4184 VSS 0.036454f
C4066 PAD.n4185 VSS 0.036454f
C4067 PAD.n4187 VSS 0.036454f
C4068 PAD.n4188 VSS 0.036454f
C4069 PAD.n4189 VSS 0.036454f
C4070 PAD.n4191 VSS 0.036454f
C4071 PAD.n4192 VSS 0.036454f
C4072 PAD.n4193 VSS 0.036454f
C4073 PAD.n4194 VSS 0.036454f
C4074 PAD.n4195 VSS 0.036454f
C4075 PAD.n4196 VSS 0.036454f
C4076 PAD.n4197 VSS 0.036454f
C4077 PAD.n4199 VSS 0.036454f
C4078 PAD.n4200 VSS 0.036454f
C4079 PAD.n4201 VSS 0.036454f
C4080 PAD.n4203 VSS 0.036454f
C4081 PAD.n4204 VSS 0.036454f
C4082 PAD.n4205 VSS 0.036454f
C4083 PAD.n4206 VSS 0.036454f
C4084 PAD.n4207 VSS 0.036454f
C4085 PAD.n4208 VSS 0.036454f
C4086 PAD.n4209 VSS 0.036454f
C4087 PAD.n4211 VSS 0.036454f
C4088 PAD.n4212 VSS 0.036454f
C4089 PAD.n4213 VSS 0.036454f
C4090 PAD.n4215 VSS 0.036454f
C4091 PAD.n4216 VSS 0.036454f
C4092 PAD.n4217 VSS 0.036454f
C4093 PAD.n4218 VSS 0.036454f
C4094 PAD.n4219 VSS 0.036454f
C4095 PAD.n4220 VSS 0.036454f
C4096 PAD.n4221 VSS 0.036454f
C4097 PAD.n4223 VSS 0.036454f
C4098 PAD.n4224 VSS 0.036454f
C4099 PAD.n4225 VSS 0.036454f
C4100 PAD.n4227 VSS 0.036454f
C4101 PAD.n4228 VSS 0.036454f
C4102 PAD.n4229 VSS 0.036454f
C4103 PAD.n4230 VSS 0.036454f
C4104 PAD.n4231 VSS 0.036454f
C4105 PAD.n4232 VSS 0.036454f
C4106 PAD.n4233 VSS 0.036454f
C4107 PAD.n4235 VSS 0.036454f
C4108 PAD.n4236 VSS 0.036454f
C4109 PAD.n4237 VSS 0.036454f
C4110 PAD.n4239 VSS 0.036454f
C4111 PAD.n4240 VSS 0.036454f
C4112 PAD.n4241 VSS 0.036454f
C4113 PAD.n4242 VSS 0.036454f
C4114 PAD.n4243 VSS 0.036454f
C4115 PAD.n4244 VSS 0.036454f
C4116 PAD.n4245 VSS 0.036454f
C4117 PAD.n4247 VSS 0.036454f
C4118 PAD.n4248 VSS 0.036454f
C4119 PAD.n4249 VSS 0.036454f
C4120 PAD.n4251 VSS 0.036454f
C4121 PAD.n4252 VSS 0.036454f
C4122 PAD.n4253 VSS 0.036454f
C4123 PAD.n4254 VSS 0.036454f
C4124 PAD.n4255 VSS 0.036454f
C4125 PAD.n4256 VSS 0.036454f
C4126 PAD.n4257 VSS 0.036454f
C4127 PAD.n4259 VSS 0.036454f
C4128 PAD.n4260 VSS 0.036454f
C4129 PAD.n4261 VSS 0.036454f
C4130 PAD.n4263 VSS 0.036454f
C4131 PAD.n4264 VSS 0.036454f
C4132 PAD.n4265 VSS 0.036454f
C4133 PAD.n4266 VSS 0.036454f
C4134 PAD.n4267 VSS 0.036454f
C4135 PAD.n4268 VSS 0.036454f
C4136 PAD.n4269 VSS 0.036454f
C4137 PAD.n4271 VSS 0.036454f
C4138 PAD.n4272 VSS 0.036454f
C4139 PAD.n4273 VSS 0.036454f
C4140 PAD.n4275 VSS 0.036454f
C4141 PAD.n4276 VSS 0.036454f
C4142 PAD.n4277 VSS 0.036454f
C4143 PAD.n4278 VSS 0.036454f
C4144 PAD.n4279 VSS 0.036454f
C4145 PAD.n4280 VSS 0.036454f
C4146 PAD.n4281 VSS 0.036454f
C4147 PAD.n4283 VSS 0.036454f
C4148 PAD.n4284 VSS 0.036454f
C4149 PAD.n4285 VSS 0.036454f
C4150 PAD.n4287 VSS 0.036454f
C4151 PAD.n4288 VSS 0.036454f
C4152 PAD.n4289 VSS 0.036454f
C4153 PAD.n4290 VSS 0.036454f
C4154 PAD.n4291 VSS 0.036454f
C4155 PAD.n4292 VSS 0.036454f
C4156 PAD.n4293 VSS 0.036454f
C4157 PAD.n4295 VSS 0.036454f
C4158 PAD.n4296 VSS 0.036454f
C4159 PAD.n4297 VSS 0.036454f
C4160 PAD.n4299 VSS 0.036454f
C4161 PAD.n4300 VSS 0.036454f
C4162 PAD.n4301 VSS 0.036454f
C4163 PAD.n4302 VSS 0.036454f
C4164 PAD.n4303 VSS 0.036454f
C4165 PAD.n4304 VSS 0.036454f
C4166 PAD.n4305 VSS 0.036454f
C4167 PAD.n4307 VSS 0.036454f
C4168 PAD.n4308 VSS 0.036454f
C4169 PAD.n4309 VSS 0.036454f
C4170 PAD.n4311 VSS 0.036454f
C4171 PAD.n4312 VSS 0.036454f
C4172 PAD.n4313 VSS 0.036454f
C4173 PAD.n4314 VSS 0.036454f
C4174 PAD.n4315 VSS 0.032467f
C4175 PAD.n4316 VSS 0.042887f
C4176 PAD.n4317 VSS 0.049106f
C4177 PAD.n4318 VSS 0.049106f
C4178 PAD.n4319 VSS 0.611619f
C4179 PAD.n4320 VSS 0.065252f
C4180 PAD.n4321 VSS 0.695471f
C4181 PAD.n4322 VSS 0.047251f
C4182 PAD.n4323 VSS 0.065252f
C4183 PAD.n4324 VSS 0.047251f
C4184 PAD.n4325 VSS 0.033374f
C4185 PAD.n4326 VSS 0.062262f
C4186 PAD.n4327 VSS 0.069752f
C4187 PAD.n4328 VSS 0.039754f
C4188 PAD.n4329 VSS 0.069752f
C4189 PAD.n4330 VSS 0.039754f
C4190 PAD.n4331 VSS 0.40939f
C4191 PAD.n4332 VSS 0.567228f
C4192 PAD.n4333 VSS 0.320607f
C4193 PAD.n4334 VSS 0.029431f
C4194 PAD.n4335 VSS 0.029431f
C4195 PAD.n4336 VSS 0.036454f
C4196 PAD.n4337 VSS 0.036454f
C4197 PAD.n4338 VSS 0.036454f
C4198 PAD.n4340 VSS 0.036454f
C4199 PAD.n4341 VSS 0.036454f
C4200 PAD.n4342 VSS 0.036454f
C4201 PAD.n4344 VSS 0.036454f
C4202 PAD.n4345 VSS 0.036454f
C4203 PAD.n4346 VSS 0.036454f
C4204 PAD.n4348 VSS 0.036454f
C4205 PAD.n4349 VSS 0.036454f
C4206 PAD.n4350 VSS 0.036454f
C4207 PAD.n4352 VSS 0.036454f
C4208 PAD.n4353 VSS 0.036454f
C4209 PAD.n4354 VSS 0.036454f
C4210 PAD.n4356 VSS 0.036454f
C4211 PAD.n4357 VSS 0.036454f
C4212 PAD.n4358 VSS 0.036454f
C4213 PAD.n4360 VSS 0.036454f
C4214 PAD.n4361 VSS 0.036454f
C4215 PAD.n4362 VSS 0.036454f
C4216 PAD.n4364 VSS 0.036454f
C4217 PAD.n4365 VSS 0.036454f
C4218 PAD.n4366 VSS 0.036454f
C4219 PAD.n4368 VSS 0.036454f
C4220 PAD.n4369 VSS 0.036454f
C4221 PAD.n4370 VSS 0.036454f
C4222 PAD.n4372 VSS 0.036454f
C4223 PAD.n4373 VSS 0.036454f
C4224 PAD.n4374 VSS 0.036454f
C4225 PAD.n4376 VSS 0.036454f
C4226 PAD.n4377 VSS 0.036454f
C4227 PAD.n4378 VSS 0.036454f
C4228 PAD.n4380 VSS 0.036454f
C4229 PAD.n4381 VSS 0.036454f
C4230 PAD.n4382 VSS 0.036454f
C4231 PAD.n4384 VSS 0.036454f
C4232 PAD.n4385 VSS 0.036454f
C4233 PAD.n4386 VSS 0.036454f
C4234 PAD.n4388 VSS 0.036454f
C4235 PAD.n4389 VSS 0.036454f
C4236 PAD.n4390 VSS 0.036454f
C4237 PAD.n4392 VSS 0.036454f
C4238 PAD.n4393 VSS 0.036454f
C4239 PAD.n4394 VSS 0.036454f
C4240 PAD.n4396 VSS 0.036454f
C4241 PAD.n4397 VSS 0.036454f
C4242 PAD.n4398 VSS 0.036454f
C4243 PAD.n4400 VSS 0.036454f
C4244 PAD.n4401 VSS 0.036454f
C4245 PAD.n4402 VSS 0.036454f
C4246 PAD.n4404 VSS 0.036454f
C4247 PAD.n4405 VSS 0.036454f
C4248 PAD.n4406 VSS 0.036454f
C4249 PAD.n4408 VSS 0.036454f
C4250 PAD.n4409 VSS 0.036454f
C4251 PAD.n4410 VSS 0.036454f
C4252 PAD.n4412 VSS 0.036454f
C4253 PAD.n4413 VSS 0.036454f
C4254 PAD.n4414 VSS 0.036454f
C4255 PAD.n4416 VSS 0.036454f
C4256 PAD.n4417 VSS 0.036454f
C4257 PAD.n4418 VSS 0.036454f
C4258 PAD.n4419 VSS 0.023105f
C4259 PAD.n4420 VSS 0.023105f
C4260 PAD.n4422 VSS 0.036454f
C4261 PAD.n4424 VSS 0.036454f
C4262 PAD.n4426 VSS 0.036454f
C4263 PAD.n4427 VSS 0.036454f
C4264 PAD.n4428 VSS 0.036454f
C4265 PAD.n4429 VSS 0.036454f
C4266 PAD.n4430 VSS 0.036454f
C4267 PAD.n4431 VSS 0.036454f
C4268 PAD.n4432 VSS 0.036454f
C4269 PAD.n4434 VSS 0.036454f
C4270 PAD.n4436 VSS 0.036454f
C4271 PAD.n4438 VSS 0.036454f
C4272 PAD.n4439 VSS 0.036454f
C4273 PAD.n4440 VSS 0.036454f
C4274 PAD.n4441 VSS 0.036454f
C4275 PAD.n4442 VSS 0.036454f
C4276 PAD.n4443 VSS 0.036454f
C4277 PAD.n4444 VSS 0.036454f
C4278 PAD.n4446 VSS 0.036454f
C4279 PAD.n4448 VSS 0.036454f
C4280 PAD.n4450 VSS 0.036454f
C4281 PAD.n4451 VSS 0.036454f
C4282 PAD.n4452 VSS 0.036454f
C4283 PAD.n4453 VSS 0.036454f
C4284 PAD.n4454 VSS 0.036454f
C4285 PAD.n4455 VSS 0.036454f
C4286 PAD.n4456 VSS 0.036454f
C4287 PAD.n4458 VSS 0.036454f
C4288 PAD.n4460 VSS 0.036454f
C4289 PAD.n4462 VSS 0.036454f
C4290 PAD.n4463 VSS 0.036454f
C4291 PAD.n4464 VSS 0.036454f
C4292 PAD.n4465 VSS 0.036454f
C4293 PAD.n4466 VSS 0.036454f
C4294 PAD.n4467 VSS 0.036454f
C4295 PAD.n4468 VSS 0.036454f
C4296 PAD.n4470 VSS 0.036454f
C4297 PAD.n4472 VSS 0.036454f
C4298 PAD.n4474 VSS 0.036454f
C4299 PAD.n4475 VSS 0.036454f
C4300 PAD.n4476 VSS 0.036454f
C4301 PAD.n4477 VSS 0.036454f
C4302 PAD.n4478 VSS 0.036454f
C4303 PAD.n4479 VSS 0.036454f
C4304 PAD.n4480 VSS 0.036454f
C4305 PAD.n4482 VSS 0.036454f
C4306 PAD.n4484 VSS 0.036454f
C4307 PAD.n4486 VSS 0.036454f
C4308 PAD.n4487 VSS 0.036454f
C4309 PAD.n4488 VSS 0.036454f
C4310 PAD.n4489 VSS 0.036454f
C4311 PAD.n4490 VSS 0.036454f
C4312 PAD.n4491 VSS 0.036454f
C4313 PAD.n4492 VSS 0.036454f
C4314 PAD.n4494 VSS 0.036454f
C4315 PAD.n4496 VSS 0.036454f
C4316 PAD.n4498 VSS 0.036454f
C4317 PAD.n4499 VSS 0.036454f
C4318 PAD.n4500 VSS 0.036454f
C4319 PAD.n4501 VSS 0.036454f
C4320 PAD.n4502 VSS 0.036454f
C4321 PAD.n4503 VSS 0.036454f
C4322 PAD.n4504 VSS 0.036454f
C4323 PAD.n4506 VSS 0.036454f
C4324 PAD.n4508 VSS 0.036454f
C4325 PAD.n4510 VSS 0.036454f
C4326 PAD.n4511 VSS 0.036454f
C4327 PAD.n4512 VSS 0.036454f
C4328 PAD.n4513 VSS 0.036454f
C4329 PAD.n4514 VSS 0.036454f
C4330 PAD.n4515 VSS 0.036454f
C4331 PAD.n4516 VSS 0.036454f
C4332 PAD.n4518 VSS 0.036454f
C4333 PAD.n4520 VSS 0.036454f
C4334 PAD.n4522 VSS 0.036454f
C4335 PAD.n4523 VSS 0.036454f
C4336 PAD.n4524 VSS 0.036454f
C4337 PAD.n4525 VSS 0.036454f
C4338 PAD.n4526 VSS 0.036454f
C4339 PAD.n4527 VSS 0.036454f
C4340 PAD.n4528 VSS 0.036454f
C4341 PAD.n4530 VSS 0.036454f
C4342 PAD.n4532 VSS 0.036454f
C4343 PAD.n4534 VSS 0.036454f
C4344 PAD.n4535 VSS 0.036454f
C4345 PAD.n4536 VSS 0.036454f
C4346 PAD.n4537 VSS 0.036454f
C4347 PAD.n4538 VSS 0.036454f
C4348 PAD.n4539 VSS 0.036454f
C4349 PAD.n4540 VSS 0.036454f
C4350 PAD.n4542 VSS 0.036454f
C4351 PAD.n4544 VSS 0.036454f
C4352 PAD.n4546 VSS 0.036454f
C4353 PAD.n4547 VSS 0.036454f
C4354 PAD.n4548 VSS 0.036454f
C4355 PAD.n4549 VSS 0.036454f
C4356 PAD.n4550 VSS 0.036454f
C4357 PAD.n4551 VSS 0.036454f
C4358 PAD.n4552 VSS 0.036454f
C4359 PAD.n4554 VSS 0.036454f
C4360 PAD.n4556 VSS 0.036454f
C4361 PAD.n4558 VSS 0.036454f
C4362 PAD.n4559 VSS 0.036454f
C4363 PAD.n4560 VSS 0.036454f
C4364 PAD.n4561 VSS 0.036454f
C4365 PAD.n4562 VSS 0.036454f
C4366 PAD.n4563 VSS 0.036454f
C4367 PAD.n4564 VSS 0.036454f
C4368 PAD.n4566 VSS 0.036454f
C4369 PAD.n4568 VSS 0.036454f
C4370 PAD.n4570 VSS 0.036454f
C4371 PAD.n4571 VSS 0.036454f
C4372 PAD.n4572 VSS 0.036454f
C4373 PAD.n4573 VSS 0.036454f
C4374 PAD.n4574 VSS 0.036454f
C4375 PAD.n4575 VSS 0.036454f
C4376 PAD.n4576 VSS 0.036454f
C4377 PAD.n4578 VSS 0.036454f
C4378 PAD.n4580 VSS 0.036454f
C4379 PAD.n4582 VSS 0.036454f
C4380 PAD.n4583 VSS 0.036454f
C4381 PAD.n4584 VSS 0.036454f
C4382 PAD.n4585 VSS 0.036454f
C4383 PAD.n4586 VSS 0.036454f
C4384 PAD.n4587 VSS 0.036454f
C4385 PAD.n4588 VSS 0.036454f
C4386 PAD.n4590 VSS 0.036454f
C4387 PAD.n4592 VSS 0.036454f
C4388 PAD.n4594 VSS 0.036454f
C4389 PAD.n4595 VSS 0.036454f
C4390 PAD.n4596 VSS 0.036454f
C4391 PAD.n4597 VSS 0.036454f
C4392 PAD.n4598 VSS 0.036454f
C4393 PAD.n4599 VSS 0.036454f
C4394 PAD.n4600 VSS 0.036454f
C4395 PAD.n4602 VSS 0.036454f
C4396 PAD.n4604 VSS 0.036454f
C4397 PAD.n4606 VSS 0.036454f
C4398 PAD.n4607 VSS 0.036454f
C4399 PAD.n4608 VSS 0.036454f
C4400 PAD.n4609 VSS 0.036454f
C4401 PAD.n4610 VSS 0.036454f
C4402 PAD.n4611 VSS 0.036454f
C4403 PAD.n4612 VSS 0.036454f
C4404 PAD.n4614 VSS 0.036454f
C4405 PAD.n4616 VSS 0.036454f
C4406 PAD.n4618 VSS 0.036454f
C4407 PAD.n4619 VSS 0.036454f
C4408 PAD.n4620 VSS 0.036454f
C4409 PAD.n4621 VSS 0.036454f
C4410 PAD.n4622 VSS 0.036454f
C4411 PAD.n4623 VSS 0.036454f
C4412 PAD.n4624 VSS 0.036454f
C4413 PAD.n4626 VSS 0.036454f
C4414 PAD.n4628 VSS 0.036454f
C4415 PAD.n4630 VSS 0.036454f
C4416 PAD.n4631 VSS 0.036454f
C4417 PAD.n4632 VSS 0.036454f
C4418 PAD.n4633 VSS 0.036454f
C4419 PAD.n4634 VSS 0.036454f
C4420 PAD.n4635 VSS 0.036454f
C4421 PAD.n4636 VSS 0.036454f
C4422 PAD.n4638 VSS 0.036454f
C4423 PAD.n4640 VSS 0.036454f
C4424 PAD.n4642 VSS 0.036454f
C4425 PAD.n4643 VSS 0.036454f
C4426 PAD.n4644 VSS 0.036454f
C4427 PAD.n4645 VSS 0.036454f
C4428 PAD.n4646 VSS 0.036454f
C4429 PAD.n4647 VSS 0.036454f
C4430 PAD.n4648 VSS 0.036454f
C4431 PAD.n4650 VSS 0.036454f
C4432 PAD.n4652 VSS 0.036454f
C4433 PAD.n4654 VSS 0.036454f
C4434 PAD.n4655 VSS 0.036454f
C4435 PAD.n4656 VSS 0.036454f
C4436 PAD.n4657 VSS 0.036454f
C4437 PAD.n4658 VSS 0.036454f
C4438 PAD.n4659 VSS 0.036454f
C4439 PAD.n4660 VSS 0.036454f
C4440 PAD.n4661 VSS 0.036454f
C4441 PAD.n4663 VSS 0.036454f
C4442 PAD.n4665 VSS 0.036454f
C4443 PAD.n4667 VSS 0.023105f
C4444 PAD.n4668 VSS 0.023105f
C4445 PAD.n4669 VSS 0.03055f
C4446 PAD.n4670 VSS 0.042887f
C4447 PAD.n4671 VSS 0.049106f
C4448 PAD.n4672 VSS 0.049106f
C4449 PAD.n4673 VSS 0.586957f
C4450 PAD.n4674 VSS 0.038251f
C4451 PAD.n4675 VSS 0.038251f
C4452 PAD.n4676 VSS 0.033374f
C4453 PAD.n4677 VSS 0.062262f
C4454 PAD.n4678 VSS 0.069752f
C4455 PAD.n4679 VSS 0.039754f
C4456 PAD.n4680 VSS 0.069752f
C4457 PAD.n4681 VSS 0.039754f
C4458 PAD.n4682 VSS 0.611619f
C4459 PAD.n4724 VSS 0.424187f
C4460 PAD.n4725 VSS 0.036454f
C4461 PAD.n4727 VSS 0.036454f
C4462 PAD.n4728 VSS 0.036454f
C4463 PAD.n4729 VSS 0.036454f
C4464 PAD.n4730 VSS 0.036454f
C4465 PAD.n4731 VSS 0.036454f
C4466 PAD.n4733 VSS 0.036454f
C4467 PAD.n4734 VSS 0.036454f
C4468 PAD.n4735 VSS 0.036454f
C4469 PAD.n4736 VSS 0.036454f
C4470 PAD.n4738 VSS 0.036454f
C4471 PAD.n4739 VSS 0.036454f
C4472 PAD.n4740 VSS 0.036454f
C4473 PAD.n4741 VSS 0.036454f
C4474 PAD.n4743 VSS 0.036454f
C4475 PAD.n4744 VSS 0.036454f
C4476 PAD.n4745 VSS 0.036454f
C4477 PAD.n4746 VSS 0.036454f
C4478 PAD.n4748 VSS 0.036454f
C4479 PAD.n4749 VSS 0.036454f
C4480 PAD.n4750 VSS 0.036454f
C4481 PAD.n4751 VSS 0.036454f
C4482 PAD.n4753 VSS 0.036454f
C4483 PAD.n4754 VSS 0.036454f
C4484 PAD.n4755 VSS 0.036454f
C4485 PAD.n4756 VSS 0.036454f
C4486 PAD.n4758 VSS 0.036454f
C4487 PAD.n4759 VSS 0.036454f
C4488 PAD.n4760 VSS 0.036454f
C4489 PAD.n4761 VSS 0.036454f
C4490 PAD.n4763 VSS 0.036454f
C4491 PAD.n4764 VSS 0.036454f
C4492 PAD.n4765 VSS 0.036454f
C4493 PAD.n4766 VSS 0.036454f
C4494 PAD.n4768 VSS 0.036454f
C4495 PAD.n4769 VSS 0.036454f
C4496 PAD.n4770 VSS 0.036454f
C4497 PAD.n4771 VSS 0.036454f
C4498 PAD.n4773 VSS 0.036454f
C4499 PAD.n4774 VSS 0.036454f
C4500 PAD.n4775 VSS 0.036454f
C4501 PAD.n4776 VSS 0.036454f
C4502 PAD.n4778 VSS 0.036454f
C4503 PAD.n4779 VSS 0.036454f
C4504 PAD.n4780 VSS 0.036454f
C4505 PAD.n4781 VSS 0.036454f
C4506 PAD.n4783 VSS 0.036454f
C4507 PAD.n4784 VSS 0.036454f
C4508 PAD.n4785 VSS 0.036454f
C4509 PAD.n4786 VSS 0.036454f
C4510 PAD.n4788 VSS 0.036454f
C4511 PAD.n4789 VSS 0.036454f
C4512 PAD.n4790 VSS 0.036454f
C4513 PAD.n4791 VSS 0.036454f
C4514 PAD.n4793 VSS 0.036454f
C4515 PAD.n4794 VSS 0.036454f
C4516 PAD.n4795 VSS 0.036454f
C4517 PAD.n4796 VSS 0.036454f
C4518 PAD.n4798 VSS 0.036454f
C4519 PAD.n4799 VSS 0.036454f
C4520 PAD.n4800 VSS 0.036454f
C4521 PAD.n4801 VSS 0.036454f
C4522 PAD.n4803 VSS 0.036454f
C4523 PAD.n4804 VSS 0.036454f
C4524 PAD.n4805 VSS 0.036454f
C4525 PAD.n4806 VSS 0.036454f
C4526 PAD.n4808 VSS 0.036454f
C4527 PAD.n4809 VSS 0.036454f
C4528 PAD.n4810 VSS 0.036454f
C4529 PAD.n4811 VSS 0.036454f
C4530 PAD.n4813 VSS 0.036454f
C4531 PAD.n4814 VSS 0.036454f
C4532 PAD.n4815 VSS 0.036454f
C4533 PAD.n4816 VSS 0.036454f
C4534 PAD.n4818 VSS 0.036454f
C4535 PAD.n4819 VSS 0.036454f
C4536 PAD.n4820 VSS 0.036454f
C4537 PAD.n4821 VSS 0.036454f
C4538 PAD.n4823 VSS 0.036454f
C4539 PAD.n4824 VSS 0.036454f
C4540 PAD.n4825 VSS 0.036454f
C4541 PAD.n4826 VSS 0.036454f
C4542 PAD.n4828 VSS 0.036454f
C4543 PAD.n4829 VSS 0.023105f
C4544 PAD.n4830 VSS 0.04032f
C4545 PAD.n4831 VSS 0.029431f
C4546 PAD.n4832 VSS 0.023105f
C4547 PAD.n4833 VSS 0.04755f
C4548 PAD.n4834 VSS 0.029431f
C4549 PAD.n4835 VSS 0.03055f
C4550 PAD.n4836 VSS 0.042887f
C4551 PAD.n4837 VSS 0.049106f
C4552 PAD.n4838 VSS 0.049106f
C4553 PAD.n4839 VSS 0.029431f
C4554 PAD.n4840 VSS 0.369931f
C4555 PAD.n4841 VSS 0.700403f
C4556 PAD.n4842 VSS 0.434052f
C4557 PAD.n4843 VSS 0.458715f
C4558 PAD.n4844 VSS 0.039754f
C4559 PAD.n4845 VSS 0.039754f
C4560 PAD.n4846 VSS 0.036454f
C4561 PAD.n4847 VSS 0.023105f
C4562 PAD.n4848 VSS 0.036454f
C4563 PAD.n4851 VSS 0.036454f
C4564 PAD.n4852 VSS 0.036454f
C4565 PAD.n4853 VSS 0.036454f
C4566 PAD.n4854 VSS 0.036454f
C4567 PAD.n4856 VSS 0.036454f
C4568 PAD.n4857 VSS 0.036454f
C4569 PAD.n4858 VSS 0.036454f
C4570 PAD.n4860 VSS 0.036454f
C4571 PAD.n4861 VSS 0.036454f
C4572 PAD.n4862 VSS 0.036454f
C4573 PAD.n4864 VSS 0.036454f
C4574 PAD.n4865 VSS 0.036454f
C4575 PAD.n4866 VSS 0.036454f
C4576 PAD.n4868 VSS 0.036454f
C4577 PAD.n4869 VSS 0.036454f
C4578 PAD.n4870 VSS 0.036454f
C4579 PAD.n4872 VSS 0.036454f
C4580 PAD.n4873 VSS 0.036454f
C4581 PAD.n4874 VSS 0.036454f
C4582 PAD.n4876 VSS 0.036454f
C4583 PAD.n4877 VSS 0.036454f
C4584 PAD.n4878 VSS 0.036454f
C4585 PAD.n4880 VSS 0.036454f
C4586 PAD.n4881 VSS 0.036454f
C4587 PAD.n4882 VSS 0.036454f
C4588 PAD.n4884 VSS 0.036454f
C4589 PAD.n4885 VSS 0.036454f
C4590 PAD.n4886 VSS 0.036454f
C4591 PAD.n4888 VSS 0.036454f
C4592 PAD.n4889 VSS 0.036454f
C4593 PAD.n4890 VSS 0.036454f
C4594 PAD.n4892 VSS 0.036454f
C4595 PAD.n4893 VSS 0.036454f
C4596 PAD.n4894 VSS 0.036454f
C4597 PAD.n4896 VSS 0.036454f
C4598 PAD.n4897 VSS 0.036454f
C4599 PAD.n4898 VSS 0.036454f
C4600 PAD.n4900 VSS 0.036454f
C4601 PAD.n4901 VSS 0.036454f
C4602 PAD.n4902 VSS 0.036454f
C4603 PAD.n4904 VSS 0.036454f
C4604 PAD.n4905 VSS 0.036454f
C4605 PAD.n4906 VSS 0.036454f
C4606 PAD.n4908 VSS 0.036454f
C4607 PAD.n4909 VSS 0.036454f
C4608 PAD.n4910 VSS 0.036454f
C4609 PAD.n4912 VSS 0.036454f
C4610 PAD.n4913 VSS 0.036454f
C4611 PAD.n4914 VSS 0.036454f
C4612 PAD.n4916 VSS 0.036454f
C4613 PAD.n4917 VSS 0.036454f
C4614 PAD.n4918 VSS 0.036454f
C4615 PAD.n4920 VSS 0.036454f
C4616 PAD.n4921 VSS 0.036454f
C4617 PAD.n4922 VSS 0.036454f
C4618 PAD.n4924 VSS 0.036454f
C4619 PAD.n4925 VSS 0.036454f
C4620 PAD.n4926 VSS 0.036454f
C4621 PAD.n4928 VSS 0.036454f
C4622 PAD.n4929 VSS 0.036454f
C4623 PAD.n4930 VSS 0.036454f
C4624 PAD.n4931 VSS 0.023105f
C4625 PAD.n4932 VSS 0.023105f
C4626 PAD.n4934 VSS 0.036454f
C4627 PAD.n4936 VSS 0.036454f
C4628 PAD.n4938 VSS 0.036454f
C4629 PAD.n4939 VSS 0.036454f
C4630 PAD.n4940 VSS 0.036454f
C4631 PAD.n4941 VSS 0.036454f
C4632 PAD.n4942 VSS 0.036454f
C4633 PAD.n4943 VSS 0.036454f
C4634 PAD.n4944 VSS 0.036454f
C4635 PAD.n4946 VSS 0.036454f
C4636 PAD.n4948 VSS 0.036454f
C4637 PAD.n4950 VSS 0.036454f
C4638 PAD.n4951 VSS 0.036454f
C4639 PAD.n4952 VSS 0.036454f
C4640 PAD.n4953 VSS 0.036454f
C4641 PAD.n4954 VSS 0.036454f
C4642 PAD.n4955 VSS 0.036454f
C4643 PAD.n4956 VSS 0.036454f
C4644 PAD.n4958 VSS 0.036454f
C4645 PAD.n4960 VSS 0.036454f
C4646 PAD.n4962 VSS 0.036454f
C4647 PAD.n4963 VSS 0.036454f
C4648 PAD.n4964 VSS 0.036454f
C4649 PAD.n4965 VSS 0.036454f
C4650 PAD.n4966 VSS 0.036454f
C4651 PAD.n4967 VSS 0.036454f
C4652 PAD.n4968 VSS 0.036454f
C4653 PAD.n4970 VSS 0.036454f
C4654 PAD.n4972 VSS 0.036454f
C4655 PAD.n4974 VSS 0.036454f
C4656 PAD.n4975 VSS 0.036454f
C4657 PAD.n4976 VSS 0.036454f
C4658 PAD.n4977 VSS 0.036454f
C4659 PAD.n4978 VSS 0.036454f
C4660 PAD.n4979 VSS 0.036454f
C4661 PAD.n4980 VSS 0.036454f
C4662 PAD.n4982 VSS 0.036454f
C4663 PAD.n4984 VSS 0.036454f
C4664 PAD.n4986 VSS 0.036454f
C4665 PAD.n4987 VSS 0.036454f
C4666 PAD.n4988 VSS 0.036454f
C4667 PAD.n4989 VSS 0.036454f
C4668 PAD.n4990 VSS 0.036454f
C4669 PAD.n4991 VSS 0.036454f
C4670 PAD.n4992 VSS 0.036454f
C4671 PAD.n4994 VSS 0.036454f
C4672 PAD.n4996 VSS 0.036454f
C4673 PAD.n4998 VSS 0.036454f
C4674 PAD.n4999 VSS 0.036454f
C4675 PAD.n5000 VSS 0.036454f
C4676 PAD.n5001 VSS 0.036454f
C4677 PAD.n5002 VSS 0.036454f
C4678 PAD.n5003 VSS 0.036454f
C4679 PAD.n5004 VSS 0.036454f
C4680 PAD.n5006 VSS 0.036454f
C4681 PAD.n5008 VSS 0.036454f
C4682 PAD.n5010 VSS 0.036454f
C4683 PAD.n5011 VSS 0.036454f
C4684 PAD.n5012 VSS 0.036454f
C4685 PAD.n5013 VSS 0.036454f
C4686 PAD.n5014 VSS 0.036454f
C4687 PAD.n5015 VSS 0.036454f
C4688 PAD.n5016 VSS 0.036454f
C4689 PAD.n5018 VSS 0.036454f
C4690 PAD.n5020 VSS 0.036454f
C4691 PAD.n5022 VSS 0.036454f
C4692 PAD.n5023 VSS 0.036454f
C4693 PAD.n5024 VSS 0.036454f
C4694 PAD.n5025 VSS 0.036454f
C4695 PAD.n5026 VSS 0.036454f
C4696 PAD.n5027 VSS 0.036454f
C4697 PAD.n5028 VSS 0.036454f
C4698 PAD.n5030 VSS 0.036454f
C4699 PAD.n5032 VSS 0.036454f
C4700 PAD.n5034 VSS 0.036454f
C4701 PAD.n5035 VSS 0.036454f
C4702 PAD.n5036 VSS 0.036454f
C4703 PAD.n5037 VSS 0.036454f
C4704 PAD.n5038 VSS 0.036454f
C4705 PAD.n5039 VSS 0.036454f
C4706 PAD.n5040 VSS 0.036454f
C4707 PAD.n5042 VSS 0.036454f
C4708 PAD.n5044 VSS 0.036454f
C4709 PAD.n5046 VSS 0.036454f
C4710 PAD.n5047 VSS 0.036454f
C4711 PAD.n5048 VSS 0.036454f
C4712 PAD.n5049 VSS 0.036454f
C4713 PAD.n5050 VSS 0.036454f
C4714 PAD.n5051 VSS 0.036454f
C4715 PAD.n5052 VSS 0.036454f
C4716 PAD.n5054 VSS 0.036454f
C4717 PAD.n5056 VSS 0.036454f
C4718 PAD.n5058 VSS 0.036454f
C4719 PAD.n5059 VSS 0.036454f
C4720 PAD.n5060 VSS 0.036454f
C4721 PAD.n5061 VSS 0.036454f
C4722 PAD.n5062 VSS 0.036454f
C4723 PAD.n5063 VSS 0.036454f
C4724 PAD.n5064 VSS 0.036454f
C4725 PAD.n5066 VSS 0.036454f
C4726 PAD.n5068 VSS 0.036454f
C4727 PAD.n5070 VSS 0.036454f
C4728 PAD.n5071 VSS 0.036454f
C4729 PAD.n5072 VSS 0.036454f
C4730 PAD.n5073 VSS 0.036454f
C4731 PAD.n5074 VSS 0.036454f
C4732 PAD.n5075 VSS 0.036454f
C4733 PAD.n5076 VSS 0.036454f
C4734 PAD.n5078 VSS 0.036454f
C4735 PAD.n5080 VSS 0.036454f
C4736 PAD.n5082 VSS 0.036454f
C4737 PAD.n5083 VSS 0.036454f
C4738 PAD.n5084 VSS 0.036454f
C4739 PAD.n5085 VSS 0.036454f
C4740 PAD.n5086 VSS 0.036454f
C4741 PAD.n5087 VSS 0.036454f
C4742 PAD.n5088 VSS 0.036454f
C4743 PAD.n5090 VSS 0.036454f
C4744 PAD.n5092 VSS 0.036454f
C4745 PAD.n5094 VSS 0.036454f
C4746 PAD.n5095 VSS 0.036454f
C4747 PAD.n5096 VSS 0.036454f
C4748 PAD.n5097 VSS 0.036454f
C4749 PAD.n5098 VSS 0.036454f
C4750 PAD.n5099 VSS 0.036454f
C4751 PAD.n5100 VSS 0.036454f
C4752 PAD.n5102 VSS 0.036454f
C4753 PAD.n5104 VSS 0.036454f
C4754 PAD.n5106 VSS 0.036454f
C4755 PAD.n5107 VSS 0.036454f
C4756 PAD.n5108 VSS 0.036454f
C4757 PAD.n5109 VSS 0.036454f
C4758 PAD.n5110 VSS 0.036454f
C4759 PAD.n5111 VSS 0.036454f
C4760 PAD.n5112 VSS 0.036454f
C4761 PAD.n5114 VSS 0.036454f
C4762 PAD.n5116 VSS 0.036454f
C4763 PAD.n5118 VSS 0.036454f
C4764 PAD.n5119 VSS 0.036454f
C4765 PAD.n5120 VSS 0.036454f
C4766 PAD.n5121 VSS 0.036454f
C4767 PAD.n5122 VSS 0.036454f
C4768 PAD.n5123 VSS 0.036454f
C4769 PAD.n5124 VSS 0.036454f
C4770 PAD.n5126 VSS 0.036454f
C4771 PAD.n5128 VSS 0.036454f
C4772 PAD.n5130 VSS 0.036454f
C4773 PAD.n5131 VSS 0.036454f
C4774 PAD.n5132 VSS 0.036454f
C4775 PAD.n5133 VSS 0.036454f
C4776 PAD.n5134 VSS 0.036454f
C4777 PAD.n5135 VSS 0.036454f
C4778 PAD.n5136 VSS 0.036454f
C4779 PAD.n5138 VSS 0.036454f
C4780 PAD.n5140 VSS 0.036454f
C4781 PAD.n5142 VSS 0.036454f
C4782 PAD.n5143 VSS 0.036454f
C4783 PAD.n5144 VSS 0.036454f
C4784 PAD.n5145 VSS 0.036454f
C4785 PAD.n5146 VSS 0.036454f
C4786 PAD.n5147 VSS 0.036454f
C4787 PAD.n5148 VSS 0.036454f
C4788 PAD.n5150 VSS 0.036454f
C4789 PAD.n5152 VSS 0.036454f
C4790 PAD.n5154 VSS 0.036454f
C4791 PAD.n5155 VSS 0.036454f
C4792 PAD.n5156 VSS 0.036454f
C4793 PAD.n5157 VSS 0.036454f
C4794 PAD.n5158 VSS 0.036454f
C4795 PAD.n5159 VSS 0.036454f
C4796 PAD.n5160 VSS 0.036454f
C4797 PAD.n5162 VSS 0.036454f
C4798 PAD.n5164 VSS 0.036454f
C4799 PAD.n5166 VSS 0.036454f
C4800 PAD.n5167 VSS 0.036454f
C4801 PAD.n5168 VSS 0.036454f
C4802 PAD.n5169 VSS 0.036454f
C4803 PAD.n5170 VSS 0.036454f
C4804 PAD.n5171 VSS 0.036454f
C4805 PAD.n5172 VSS 0.036454f
C4806 PAD.n5174 VSS 0.036454f
C4807 PAD.n5176 VSS 0.036454f
C4808 PAD.n5177 VSS 0.036454f
C4809 PAD.n5178 VSS 0.023105f
C4810 PAD.n5179 VSS 0.033374f
C4811 PAD.n5180 VSS 0.062262f
C4812 PAD.n5181 VSS 0.069752f
C4813 PAD.n5182 VSS 0.069752f
C4814 PAD.n5183 VSS 0.192364f
C4815 PAD.n5184 VSS 0.029431f
C4816 PAD.n5185 VSS 0.029431f
C4817 PAD.n5186 VSS 0.03055f
C4818 PAD.n5187 VSS 0.042887f
C4819 PAD.n5188 VSS 0.049106f
C4820 PAD.n5189 VSS 0.049106f
C4821 PAD.n5190 VSS 0.172634f
C4822 PAD.n5191 VSS 0.039754f
C4823 PAD.n5192 VSS 0.039754f
C4824 PAD.n5193 VSS 0.033374f
C4825 PAD.n5194 VSS 0.051718f
C4826 PAD.n5195 VSS 0.069752f
C4827 PAD.n5196 VSS 0.061877f
C4828 PAD.n5197 VSS 0.537633f
C4829 PAD.n5198 VSS 0.029431f
C4830 PAD.n5199 VSS 0.029431f
C4831 PAD.n5200 VSS 0.03055f
C4832 PAD.n5201 VSS 0.042887f
C4833 PAD.n5202 VSS 0.049106f
C4834 PAD.n5203 VSS 0.049106f
C4835 PAD.n5204 VSS 0.44885f
C4836 PAD.n5205 VSS 0.069752f
C4837 PAD.n5206 VSS 0.039754f
C4838 PAD.n5207 VSS 0.069752f
C4839 PAD.n5208 VSS 0.039754f
C4840 PAD.n5209 VSS 0.062262f
C4841 PAD.n5210 VSS 0.036454f
C4842 PAD.n5211 VSS 0.023105f
C4843 PAD.n5212 VSS 0.036454f
C4844 PAD.n5215 VSS 0.036454f
C4845 PAD.n5216 VSS 0.036454f
C4846 PAD.n5217 VSS 0.036454f
C4847 PAD.n5218 VSS 0.036454f
C4848 PAD.n5220 VSS 0.036454f
C4849 PAD.n5221 VSS 0.036454f
C4850 PAD.n5222 VSS 0.036454f
C4851 PAD.n5224 VSS 0.036454f
C4852 PAD.n5225 VSS 0.036454f
C4853 PAD.n5226 VSS 0.036454f
C4854 PAD.n5228 VSS 0.036454f
C4855 PAD.n5229 VSS 0.036454f
C4856 PAD.n5230 VSS 0.036454f
C4857 PAD.n5232 VSS 0.036454f
C4858 PAD.n5233 VSS 0.036454f
C4859 PAD.n5234 VSS 0.036454f
C4860 PAD.n5236 VSS 0.036454f
C4861 PAD.n5237 VSS 0.036454f
C4862 PAD.n5238 VSS 0.036454f
C4863 PAD.n5240 VSS 0.036454f
C4864 PAD.n5241 VSS 0.036454f
C4865 PAD.n5242 VSS 0.036454f
C4866 PAD.n5244 VSS 0.036454f
C4867 PAD.n5245 VSS 0.036454f
C4868 PAD.n5246 VSS 0.036454f
C4869 PAD.n5248 VSS 0.036454f
C4870 PAD.n5249 VSS 0.036454f
C4871 PAD.n5250 VSS 0.036454f
C4872 PAD.n5252 VSS 0.036454f
C4873 PAD.n5253 VSS 0.036454f
C4874 PAD.n5254 VSS 0.036454f
C4875 PAD.n5256 VSS 0.036454f
C4876 PAD.n5257 VSS 0.036454f
C4877 PAD.n5258 VSS 0.036454f
C4878 PAD.n5260 VSS 0.036454f
C4879 PAD.n5261 VSS 0.036454f
C4880 PAD.n5262 VSS 0.036454f
C4881 PAD.n5264 VSS 0.036454f
C4882 PAD.n5265 VSS 0.036454f
C4883 PAD.n5266 VSS 0.036454f
C4884 PAD.n5268 VSS 0.036454f
C4885 PAD.n5269 VSS 0.036454f
C4886 PAD.n5270 VSS 0.036454f
C4887 PAD.n5272 VSS 0.036454f
C4888 PAD.n5273 VSS 0.036454f
C4889 PAD.n5274 VSS 0.036454f
C4890 PAD.n5276 VSS 0.036454f
C4891 PAD.n5277 VSS 0.036454f
C4892 PAD.n5278 VSS 0.036454f
C4893 PAD.n5280 VSS 0.036454f
C4894 PAD.n5281 VSS 0.036454f
C4895 PAD.n5282 VSS 0.036454f
C4896 PAD.n5284 VSS 0.036454f
C4897 PAD.n5285 VSS 0.036454f
C4898 PAD.n5286 VSS 0.036454f
C4899 PAD.n5288 VSS 0.036454f
C4900 PAD.n5289 VSS 0.036454f
C4901 PAD.n5290 VSS 0.036454f
C4902 PAD.n5292 VSS 0.036454f
C4903 PAD.n5293 VSS 0.036454f
C4904 PAD.n5294 VSS 0.036454f
C4905 PAD.n5295 VSS 0.023105f
C4906 PAD.n5296 VSS 0.023105f
C4907 PAD.n5298 VSS 0.036454f
C4908 PAD.n5300 VSS 0.036454f
C4909 PAD.n5302 VSS 0.036454f
C4910 PAD.n5303 VSS 0.036454f
C4911 PAD.n5304 VSS 0.036454f
C4912 PAD.n5305 VSS 0.036454f
C4913 PAD.n5306 VSS 0.036454f
C4914 PAD.n5307 VSS 0.036454f
C4915 PAD.n5308 VSS 0.036454f
C4916 PAD.n5310 VSS 0.036454f
C4917 PAD.n5312 VSS 0.036454f
C4918 PAD.n5314 VSS 0.036454f
C4919 PAD.n5315 VSS 0.036454f
C4920 PAD.n5316 VSS 0.036454f
C4921 PAD.n5317 VSS 0.036454f
C4922 PAD.n5318 VSS 0.036454f
C4923 PAD.n5319 VSS 0.036454f
C4924 PAD.n5320 VSS 0.036454f
C4925 PAD.n5322 VSS 0.036454f
C4926 PAD.n5324 VSS 0.036454f
C4927 PAD.n5326 VSS 0.036454f
C4928 PAD.n5327 VSS 0.036454f
C4929 PAD.n5328 VSS 0.036454f
C4930 PAD.n5329 VSS 0.036454f
C4931 PAD.n5330 VSS 0.036454f
C4932 PAD.n5331 VSS 0.036454f
C4933 PAD.n5332 VSS 0.036454f
C4934 PAD.n5334 VSS 0.036454f
C4935 PAD.n5336 VSS 0.036454f
C4936 PAD.n5338 VSS 0.036454f
C4937 PAD.n5339 VSS 0.036454f
C4938 PAD.n5340 VSS 0.036454f
C4939 PAD.n5341 VSS 0.036454f
C4940 PAD.n5342 VSS 0.036454f
C4941 PAD.n5343 VSS 0.036454f
C4942 PAD.n5344 VSS 0.036454f
C4943 PAD.n5346 VSS 0.036454f
C4944 PAD.n5348 VSS 0.036454f
C4945 PAD.n5350 VSS 0.036454f
C4946 PAD.n5351 VSS 0.036454f
C4947 PAD.n5352 VSS 0.036454f
C4948 PAD.n5353 VSS 0.036454f
C4949 PAD.n5354 VSS 0.036454f
C4950 PAD.n5355 VSS 0.036454f
C4951 PAD.n5356 VSS 0.036454f
C4952 PAD.n5358 VSS 0.036454f
C4953 PAD.n5360 VSS 0.036454f
C4954 PAD.n5362 VSS 0.036454f
C4955 PAD.n5363 VSS 0.036454f
C4956 PAD.n5364 VSS 0.036454f
C4957 PAD.n5365 VSS 0.036454f
C4958 PAD.n5366 VSS 0.036454f
C4959 PAD.n5367 VSS 0.036454f
C4960 PAD.n5368 VSS 0.036454f
C4961 PAD.n5370 VSS 0.036454f
C4962 PAD.n5372 VSS 0.036454f
C4963 PAD.n5374 VSS 0.036454f
C4964 PAD.n5375 VSS 0.036454f
C4965 PAD.n5376 VSS 0.036454f
C4966 PAD.n5377 VSS 0.036454f
C4967 PAD.n5378 VSS 0.036454f
C4968 PAD.n5379 VSS 0.036454f
C4969 PAD.n5380 VSS 0.036454f
C4970 PAD.n5382 VSS 0.036454f
C4971 PAD.n5384 VSS 0.036454f
C4972 PAD.n5386 VSS 0.036454f
C4973 PAD.n5387 VSS 0.036454f
C4974 PAD.n5388 VSS 0.036454f
C4975 PAD.n5389 VSS 0.036454f
C4976 PAD.n5390 VSS 0.036454f
C4977 PAD.n5391 VSS 0.036454f
C4978 PAD.n5392 VSS 0.036454f
C4979 PAD.n5394 VSS 0.036454f
C4980 PAD.n5396 VSS 0.036454f
C4981 PAD.n5398 VSS 0.036454f
C4982 PAD.n5399 VSS 0.036454f
C4983 PAD.n5400 VSS 0.036454f
C4984 PAD.n5401 VSS 0.036454f
C4985 PAD.n5402 VSS 0.036454f
C4986 PAD.n5403 VSS 0.036454f
C4987 PAD.n5404 VSS 0.036454f
C4988 PAD.n5406 VSS 0.036454f
C4989 PAD.n5408 VSS 0.036454f
C4990 PAD.n5410 VSS 0.036454f
C4991 PAD.n5411 VSS 0.036454f
C4992 PAD.n5412 VSS 0.036454f
C4993 PAD.n5413 VSS 0.036454f
C4994 PAD.n5414 VSS 0.036454f
C4995 PAD.n5415 VSS 0.036454f
C4996 PAD.n5416 VSS 0.036454f
C4997 PAD.n5418 VSS 0.036454f
C4998 PAD.n5420 VSS 0.036454f
C4999 PAD.n5422 VSS 0.036454f
C5000 PAD.n5423 VSS 0.036454f
C5001 PAD.n5424 VSS 0.036454f
C5002 PAD.n5425 VSS 0.036454f
C5003 PAD.n5426 VSS 0.036454f
C5004 PAD.n5427 VSS 0.036454f
C5005 PAD.n5428 VSS 0.036454f
C5006 PAD.n5430 VSS 0.036454f
C5007 PAD.n5432 VSS 0.036454f
C5008 PAD.n5434 VSS 0.036454f
C5009 PAD.n5435 VSS 0.036454f
C5010 PAD.n5436 VSS 0.036454f
C5011 PAD.n5437 VSS 0.036454f
C5012 PAD.n5438 VSS 0.036454f
C5013 PAD.n5439 VSS 0.036454f
C5014 PAD.n5440 VSS 0.036454f
C5015 PAD.n5442 VSS 0.036454f
C5016 PAD.n5444 VSS 0.036454f
C5017 PAD.n5446 VSS 0.036454f
C5018 PAD.n5447 VSS 0.036454f
C5019 PAD.n5448 VSS 0.036454f
C5020 PAD.n5449 VSS 0.036454f
C5021 PAD.n5450 VSS 0.036454f
C5022 PAD.n5451 VSS 0.036454f
C5023 PAD.n5452 VSS 0.036454f
C5024 PAD.n5454 VSS 0.036454f
C5025 PAD.n5456 VSS 0.036454f
C5026 PAD.n5458 VSS 0.036454f
C5027 PAD.n5459 VSS 0.036454f
C5028 PAD.n5460 VSS 0.036454f
C5029 PAD.n5461 VSS 0.036454f
C5030 PAD.n5462 VSS 0.036454f
C5031 PAD.n5463 VSS 0.036454f
C5032 PAD.n5464 VSS 0.036454f
C5033 PAD.n5466 VSS 0.036454f
C5034 PAD.n5468 VSS 0.036454f
C5035 PAD.n5470 VSS 0.036454f
C5036 PAD.n5471 VSS 0.036454f
C5037 PAD.n5472 VSS 0.036454f
C5038 PAD.n5473 VSS 0.036454f
C5039 PAD.n5474 VSS 0.036454f
C5040 PAD.n5475 VSS 0.036454f
C5041 PAD.n5476 VSS 0.036454f
C5042 PAD.n5478 VSS 0.036454f
C5043 PAD.n5480 VSS 0.036454f
C5044 PAD.n5482 VSS 0.036454f
C5045 PAD.n5483 VSS 0.036454f
C5046 PAD.n5484 VSS 0.036454f
C5047 PAD.n5485 VSS 0.036454f
C5048 PAD.n5486 VSS 0.036454f
C5049 PAD.n5487 VSS 0.036454f
C5050 PAD.n5488 VSS 0.036454f
C5051 PAD.n5490 VSS 0.036454f
C5052 PAD.n5492 VSS 0.036454f
C5053 PAD.n5494 VSS 0.036454f
C5054 PAD.n5495 VSS 0.036454f
C5055 PAD.n5496 VSS 0.036454f
C5056 PAD.n5497 VSS 0.036454f
C5057 PAD.n5498 VSS 0.036454f
C5058 PAD.n5499 VSS 0.036454f
C5059 PAD.n5500 VSS 0.036454f
C5060 PAD.n5502 VSS 0.036454f
C5061 PAD.n5504 VSS 0.036454f
C5062 PAD.n5506 VSS 0.036454f
C5063 PAD.n5507 VSS 0.036454f
C5064 PAD.n5508 VSS 0.036454f
C5065 PAD.n5509 VSS 0.036454f
C5066 PAD.n5510 VSS 0.036454f
C5067 PAD.n5511 VSS 0.036454f
C5068 PAD.n5512 VSS 0.036454f
C5069 PAD.n5514 VSS 0.036454f
C5070 PAD.n5516 VSS 0.036454f
C5071 PAD.n5518 VSS 0.036454f
C5072 PAD.n5519 VSS 0.036454f
C5073 PAD.n5520 VSS 0.036454f
C5074 PAD.n5521 VSS 0.036454f
C5075 PAD.n5522 VSS 0.036454f
C5076 PAD.n5523 VSS 0.036454f
C5077 PAD.n5524 VSS 0.036454f
C5078 PAD.n5526 VSS 0.036454f
C5079 PAD.n5528 VSS 0.036454f
C5080 PAD.n5530 VSS 0.036454f
C5081 PAD.n5531 VSS 0.036454f
C5082 PAD.n5532 VSS 0.036454f
C5083 PAD.n5533 VSS 0.036454f
C5084 PAD.n5534 VSS 0.036454f
C5085 PAD.n5535 VSS 0.036454f
C5086 PAD.n5536 VSS 0.036454f
C5087 PAD.n5538 VSS 0.036454f
C5088 PAD.n5540 VSS 0.036454f
C5089 PAD.n5541 VSS 0.036454f
C5090 PAD.n5542 VSS 0.023105f
C5091 PAD.n5543 VSS 0.033374f
C5092 PAD.n5544 VSS 0.03565f
C5093 PAD.n5545 VSS 0.033374f
C5094 PAD.n5546 VSS 0.062262f
C5095 PAD.n5547 VSS 0.039754f
C5096 PAD.n5548 VSS 0.069752f
C5097 PAD.n5549 VSS 0.039754f
C5098 PAD.n5550 VSS 0.069752f
C5099 PAD.n5551 VSS 0.527768f
C5100 PAD.n5552 VSS 0.700403f
C5101 PAD.n5553 VSS 0.029431f
C5102 PAD.n5554 VSS 0.048587f
C5103 PAD.n5555 VSS 0.029431f
C5104 PAD.n5556 VSS 0.048587f
C5105 PAD.n5557 VSS 0.03055f
C5106 PAD.n5558 VSS 0.042887f
C5107 PAD.n5559 VSS 0.049106f
C5108 PAD.n5560 VSS 0.049106f
C5109 PAD.n5602 VSS 0.036454f
C5110 PAD.n5604 VSS 0.036454f
C5111 PAD.n5605 VSS 0.036454f
C5112 PAD.n5606 VSS 0.036454f
C5113 PAD.n5607 VSS 0.036454f
C5114 PAD.n5608 VSS 0.036454f
C5115 PAD.n5610 VSS 0.036454f
C5116 PAD.n5611 VSS 0.036454f
C5117 PAD.n5612 VSS 0.036454f
C5118 PAD.n5613 VSS 0.036454f
C5119 PAD.n5615 VSS 0.036454f
C5120 PAD.n5616 VSS 0.036454f
C5121 PAD.n5617 VSS 0.036454f
C5122 PAD.n5618 VSS 0.036454f
C5123 PAD.n5620 VSS 0.036454f
C5124 PAD.n5621 VSS 0.036454f
C5125 PAD.n5622 VSS 0.036454f
C5126 PAD.n5623 VSS 0.036454f
C5127 PAD.n5625 VSS 0.036454f
C5128 PAD.n5626 VSS 0.036454f
C5129 PAD.n5627 VSS 0.036454f
C5130 PAD.n5628 VSS 0.036454f
C5131 PAD.n5630 VSS 0.036454f
C5132 PAD.n5631 VSS 0.036454f
C5133 PAD.n5632 VSS 0.036454f
C5134 PAD.n5633 VSS 0.036454f
C5135 PAD.n5635 VSS 0.036454f
C5136 PAD.n5636 VSS 0.036454f
C5137 PAD.n5637 VSS 0.036454f
C5138 PAD.n5638 VSS 0.036454f
C5139 PAD.n5640 VSS 0.036454f
C5140 PAD.n5641 VSS 0.036454f
C5141 PAD.n5642 VSS 0.036454f
C5142 PAD.n5643 VSS 0.036454f
C5143 PAD.n5645 VSS 0.036454f
C5144 PAD.n5646 VSS 0.036454f
C5145 PAD.n5647 VSS 0.036454f
C5146 PAD.n5648 VSS 0.036454f
C5147 PAD.n5650 VSS 0.036454f
C5148 PAD.n5651 VSS 0.036454f
C5149 PAD.n5652 VSS 0.036454f
C5150 PAD.n5653 VSS 0.036454f
C5151 PAD.n5655 VSS 0.036454f
C5152 PAD.n5656 VSS 0.036454f
C5153 PAD.n5657 VSS 0.036454f
C5154 PAD.n5658 VSS 0.036454f
C5155 PAD.n5660 VSS 0.036454f
C5156 PAD.n5661 VSS 0.036454f
C5157 PAD.n5662 VSS 0.036454f
C5158 PAD.n5663 VSS 0.036454f
C5159 PAD.n5665 VSS 0.036454f
C5160 PAD.n5666 VSS 0.036454f
C5161 PAD.n5667 VSS 0.036454f
C5162 PAD.n5668 VSS 0.036454f
C5163 PAD.n5670 VSS 0.036454f
C5164 PAD.n5671 VSS 0.036454f
C5165 PAD.n5672 VSS 0.036454f
C5166 PAD.n5673 VSS 0.036454f
C5167 PAD.n5675 VSS 0.036454f
C5168 PAD.n5676 VSS 0.036454f
C5169 PAD.n5677 VSS 0.036454f
C5170 PAD.n5678 VSS 0.036454f
C5171 PAD.n5680 VSS 0.036454f
C5172 PAD.n5681 VSS 0.036454f
C5173 PAD.n5682 VSS 0.036454f
C5174 PAD.n5683 VSS 0.036454f
C5175 PAD.n5685 VSS 0.036454f
C5176 PAD.n5686 VSS 0.036454f
C5177 PAD.n5687 VSS 0.036454f
C5178 PAD.n5688 VSS 0.036454f
C5179 PAD.n5690 VSS 0.036454f
C5180 PAD.n5691 VSS 0.036454f
C5181 PAD.n5692 VSS 0.036454f
C5182 PAD.n5693 VSS 0.036454f
C5183 PAD.n5695 VSS 0.036454f
C5184 PAD.n5696 VSS 0.036454f
C5185 PAD.n5697 VSS 0.036454f
C5186 PAD.n5698 VSS 0.036454f
C5187 PAD.n5700 VSS 0.036454f
C5188 PAD.n5701 VSS 0.036454f
C5189 PAD.n5702 VSS 0.023105f
C5190 PAD.n5703 VSS 0.023105f
C5191 PAD.n5704 VSS 0.036454f
C5192 PAD.n5705 VSS 0.036454f
C5193 PAD.n5707 VSS 0.036454f
C5194 PAD.n5708 VSS 0.036454f
C5195 PAD.n5709 VSS 0.036454f
C5196 PAD.n5710 VSS 0.036454f
C5197 PAD.n5711 VSS 0.036454f
C5198 PAD.n5712 VSS 0.036454f
C5199 PAD.n5714 VSS 0.036454f
C5200 PAD.n5715 VSS 0.036454f
C5201 PAD.n5716 VSS 0.036454f
C5202 PAD.n5717 VSS 0.036454f
C5203 PAD.n5718 VSS 0.036454f
C5204 PAD.n5719 VSS 0.036454f
C5205 PAD.n5720 VSS 0.036454f
C5206 PAD.n5721 VSS 0.036454f
C5207 PAD.n5723 VSS 0.036454f
C5208 PAD.n5724 VSS 0.036454f
C5209 PAD.n5725 VSS 0.036454f
C5210 PAD.n5726 VSS 0.036454f
C5211 PAD.n5727 VSS 0.036454f
C5212 PAD.n5728 VSS 0.036454f
C5213 PAD.n5729 VSS 0.036454f
C5214 PAD.n5730 VSS 0.036454f
C5215 PAD.n5732 VSS 0.036454f
C5216 PAD.n5733 VSS 0.036454f
C5217 PAD.n5734 VSS 0.036454f
C5218 PAD.n5735 VSS 0.036454f
C5219 PAD.n5736 VSS 0.036454f
C5220 PAD.n5737 VSS 0.036454f
C5221 PAD.n5738 VSS 0.036454f
C5222 PAD.n5739 VSS 0.036454f
C5223 PAD.n5741 VSS 0.036454f
C5224 PAD.n5742 VSS 0.036454f
C5225 PAD.n5743 VSS 0.036454f
C5226 PAD.n5744 VSS 0.036454f
C5227 PAD.n5745 VSS 0.036454f
C5228 PAD.n5746 VSS 0.036454f
C5229 PAD.n5747 VSS 0.036454f
C5230 PAD.n5748 VSS 0.036454f
C5231 PAD.n5750 VSS 0.036454f
C5232 PAD.n5751 VSS 0.036454f
C5233 PAD.n5752 VSS 0.036454f
C5234 PAD.n5753 VSS 0.036454f
C5235 PAD.n5754 VSS 0.036454f
C5236 PAD.n5755 VSS 0.036454f
C5237 PAD.n5756 VSS 0.036454f
C5238 PAD.n5757 VSS 0.036454f
C5239 PAD.n5759 VSS 0.036454f
C5240 PAD.n5760 VSS 0.036454f
C5241 PAD.n5761 VSS 0.036454f
C5242 PAD.n5762 VSS 0.036454f
C5243 PAD.n5763 VSS 0.036454f
C5244 PAD.n5764 VSS 0.036454f
C5245 PAD.n5765 VSS 0.036454f
C5246 PAD.n5766 VSS 0.036454f
C5247 PAD.n5768 VSS 0.036454f
C5248 PAD.n5769 VSS 0.036454f
C5249 PAD.n5770 VSS 0.036454f
C5250 PAD.n5771 VSS 0.036454f
C5251 PAD.n5772 VSS 0.036454f
C5252 PAD.n5773 VSS 0.036454f
C5253 PAD.n5774 VSS 0.036454f
C5254 PAD.n5775 VSS 0.036454f
C5255 PAD.n5777 VSS 0.036454f
C5256 PAD.n5778 VSS 0.036454f
C5257 PAD.n5779 VSS 0.036454f
C5258 PAD.n5780 VSS 0.036454f
C5259 PAD.n5781 VSS 0.036454f
C5260 PAD.n5782 VSS 0.036454f
C5261 PAD.n5783 VSS 0.036454f
C5262 PAD.n5784 VSS 0.036454f
C5263 PAD.n5786 VSS 0.036454f
C5264 PAD.n5787 VSS 0.036454f
C5265 PAD.n5788 VSS 0.036454f
C5266 PAD.n5789 VSS 0.036454f
C5267 PAD.n5790 VSS 0.036454f
C5268 PAD.n5791 VSS 0.036454f
C5269 PAD.n5792 VSS 0.036454f
C5270 PAD.n5793 VSS 0.036454f
C5271 PAD.n5795 VSS 0.036454f
C5272 PAD.n5796 VSS 0.036454f
C5273 PAD.n5797 VSS 0.036454f
C5274 PAD.n5798 VSS 0.036454f
C5275 PAD.n5799 VSS 0.036454f
C5276 PAD.n5800 VSS 0.036454f
C5277 PAD.n5801 VSS 0.036454f
C5278 PAD.n5802 VSS 0.036454f
C5279 PAD.n5804 VSS 0.036454f
C5280 PAD.n5805 VSS 0.036454f
C5281 PAD.n5806 VSS 0.036454f
C5282 PAD.n5807 VSS 0.036454f
C5283 PAD.n5808 VSS 0.036454f
C5284 PAD.n5809 VSS 0.036454f
C5285 PAD.n5810 VSS 0.036454f
C5286 PAD.n5811 VSS 0.036454f
C5287 PAD.n5813 VSS 0.036454f
C5288 PAD.n5814 VSS 0.036454f
C5289 PAD.n5815 VSS 0.036454f
C5290 PAD.n5816 VSS 0.036454f
C5291 PAD.n5817 VSS 0.036454f
C5292 PAD.n5818 VSS 0.036454f
C5293 PAD.n5819 VSS 0.036454f
C5294 PAD.n5820 VSS 0.036454f
C5295 PAD.n5822 VSS 0.036454f
C5296 PAD.n5823 VSS 0.036454f
C5297 PAD.n5824 VSS 0.036454f
C5298 PAD.n5825 VSS 0.036454f
C5299 PAD.n5826 VSS 0.036454f
C5300 PAD.n5827 VSS 0.036454f
C5301 PAD.n5828 VSS 0.036454f
C5302 PAD.n5829 VSS 0.036454f
C5303 PAD.n5831 VSS 0.036454f
C5304 PAD.n5832 VSS 0.036454f
C5305 PAD.n5833 VSS 0.036454f
C5306 PAD.n5834 VSS 0.036454f
C5307 PAD.n5835 VSS 0.036454f
C5308 PAD.n5836 VSS 0.036454f
C5309 PAD.n5837 VSS 0.036454f
C5310 PAD.n5838 VSS 0.036454f
C5311 PAD.n5840 VSS 0.036454f
C5312 PAD.n5841 VSS 0.036454f
C5313 PAD.n5842 VSS 0.036454f
C5314 PAD.n5843 VSS 0.036454f
C5315 PAD.n5844 VSS 0.036454f
C5316 PAD.n5845 VSS 0.036454f
C5317 PAD.n5846 VSS 0.036454f
C5318 PAD.n5847 VSS 0.036454f
C5319 PAD.n5849 VSS 0.036454f
C5320 PAD.n5850 VSS 0.036454f
C5321 PAD.n5851 VSS 0.036454f
C5322 PAD.n5852 VSS 0.036454f
C5323 PAD.n5853 VSS 0.036454f
C5324 PAD.n5854 VSS 0.036454f
C5325 PAD.n5855 VSS 0.036454f
C5326 PAD.n5856 VSS 0.036454f
C5327 PAD.n5858 VSS 0.036454f
C5328 PAD.n5859 VSS 0.036454f
C5329 PAD.n5860 VSS 0.036454f
C5330 PAD.n5861 VSS 0.036454f
C5331 PAD.n5862 VSS 0.036454f
C5332 PAD.n5863 VSS 0.036454f
C5333 PAD.n5864 VSS 0.036454f
C5334 PAD.n5865 VSS 0.036454f
C5335 PAD.n5867 VSS 0.036454f
C5336 PAD.n5868 VSS 0.036454f
C5337 PAD.n5869 VSS 0.036454f
C5338 PAD.n5870 VSS 0.036454f
C5339 PAD.n5871 VSS 0.036454f
C5340 PAD.n5872 VSS 0.036454f
C5341 PAD.n5873 VSS 0.036454f
C5342 PAD.n5874 VSS 0.036454f
C5343 PAD.n5876 VSS 0.036454f
C5344 PAD.n5877 VSS 0.036454f
C5345 PAD.n5878 VSS 0.036454f
C5346 PAD.n5879 VSS 0.036454f
C5347 PAD.n5880 VSS 0.036454f
C5348 PAD.n5881 VSS 0.036454f
C5349 PAD.n5882 VSS 0.036454f
C5350 PAD.n5883 VSS 0.036454f
C5351 PAD.n5885 VSS 0.036454f
C5352 PAD.n5886 VSS 0.036454f
C5353 PAD.n5887 VSS 0.036454f
C5354 PAD.n5888 VSS 0.036454f
C5355 PAD.n5889 VSS 0.036454f
C5356 PAD.n5890 VSS 0.036454f
C5357 PAD.n5891 VSS 0.023105f
C5358 PAD.n5892 VSS 0.023105f
C5359 PAD.n5894 VSS 0.61162f
C5360 PAD.n5895 VSS 0.069752f
C5361 PAD.n5896 VSS 0.066377f
C5362 PAD.n5897 VSS 0.034144f
C5363 PAD.n5898 VSS 0.036454f
C5364 PAD.n5899 VSS 0.039754f
C5365 PAD.n5900 VSS 0.036454f
C5366 PAD.n5901 VSS 0.039754f
C5367 PAD.n5903 VSS 0.582025f
C5368 PAD.n5904 VSS 0.300877f
C5369 PAD.n5905 VSS 0.036454f
C5370 PAD.n5948 VSS 0.029431f
C5371 PAD.n5949 VSS 0.036454f
C5372 PAD.n5950 VSS 0.036454f
C5373 PAD.n5951 VSS 0.03055f
C5374 PAD.n5952 VSS 0.033025f
C5375 PAD.n5953 VSS 0.035488f
C5376 PAD.n5954 VSS 0.069752f
C5377 PAD.n5955 VSS 0.063565f
C5378 PAD.n5956 VSS 0.128762f
C5379 PAD.n5957 VSS 0.103594f
C5380 PAD.n5958 VSS 0.066139f
C5381 PAD.n5959 VSS 0.103594f
C5382 PAD.n5960 VSS 0.066139f
C5383 PAD.n5962 VSS 0.61162f
C5384 PAD.n5963 VSS 0.61162f
C5385 PAD.n5964 VSS 0.61162f
C5386 PAD.n5965 VSS 0.61162f
C5387 PAD.n5966 VSS 0.651079f
C5388 PAD.n5967 VSS 0.069163f
C5389 PAD.n5968 VSS 0.069163f
C5390 PAD.n5969 VSS 0.103594f
C5391 PAD.n5970 VSS 0.063565f
C5392 PAD.n5971 VSS 0.700403f
C5393 PAD.n5972 VSS 0.042465f
C5394 PAD.n5973 VSS 0.033025f
C5395 PAD.n5974 VSS 0.611619f
C5396 PAD.n5975 VSS 0.049106f
C5397 PAD.n5976 VSS 0.042465f
C5398 PAD.n5977 VSS 0.049106f
C5399 PAD.n5978 VSS 0.068257f
C5400 PAD.n5979 VSS 0.61162f
C5401 PAD.n5980 VSS 0.61162f
C5402 PAD.n5981 VSS 0.61162f
C5403 PAD.n5982 VSS 0.61162f
C5404 PAD.n5983 VSS 0.074902f
C5405 PAD.n5984 VSS 0.074902f
C5406 PAD.n5985 VSS 0.074902f
C5407 PAD.n5986 VSS 0.074902f
C5408 PAD.n5987 VSS 0.074902f
C5409 PAD.n5988 VSS 0.074902f
C5410 PAD.n5989 VSS 0.074902f
C5411 PAD.n5990 VSS 0.074902f
C5412 PAD.n5991 VSS 0.074902f
C5413 PAD.n5992 VSS 0.074902f
C5414 PAD.n5993 VSS 0.074902f
C5415 PAD.n5994 VSS 0.074902f
C5416 PAD.n5995 VSS 0.074902f
C5417 PAD.n5996 VSS 0.074902f
C5418 PAD.n5997 VSS 0.074902f
C5419 PAD.n5998 VSS 0.074902f
C5420 PAD.n5999 VSS 0.074902f
C5421 PAD.n6000 VSS 0.074902f
C5422 PAD.n6001 VSS 0.074902f
C5423 PAD.n6002 VSS 0.074902f
C5424 PAD.n6003 VSS 0.074902f
C5425 PAD.n6004 VSS 0.074902f
C5426 PAD.n6005 VSS 0.074902f
C5427 PAD.n6006 VSS 0.074902f
C5428 PAD.n6007 VSS 0.074902f
C5429 PAD.n6008 VSS 0.074902f
C5430 PAD.n6009 VSS 0.074902f
C5431 PAD.n6010 VSS 0.074902f
C5432 PAD.n6011 VSS 0.074902f
C5433 PAD.n6012 VSS 0.074902f
C5434 PAD.n6013 VSS 0.074902f
C5435 PAD.n6014 VSS 0.074902f
C5436 PAD.n6015 VSS 0.074902f
C5437 PAD.n6016 VSS 0.074902f
C5438 PAD.n6017 VSS 0.074902f
C5439 PAD.n6018 VSS 0.074902f
C5440 PAD.n6019 VSS 0.074902f
C5441 PAD.n6020 VSS 0.074902f
C5442 PAD.n6021 VSS 0.074902f
C5443 PAD.n6022 VSS 0.074902f
C5444 PAD.n6023 VSS 0.074902f
C5445 PAD.n6024 VSS 0.074902f
C5446 PAD.n6025 VSS 0.074902f
C5447 PAD.n6026 VSS 0.074902f
C5448 PAD.n6027 VSS 0.074902f
C5449 PAD.n6028 VSS 0.074902f
C5450 PAD.n6029 VSS 0.074902f
C5451 PAD.n6030 VSS 0.074902f
C5452 PAD.n6032 VSS 0.074902f
C5453 PAD.n6034 VSS 0.103594f
C5454 PAD.n6037 VSS 0.074902f
C5455 PAD.n6040 VSS 0.074902f
C5456 PAD.n6043 VSS 0.074902f
C5457 PAD.n6046 VSS 0.074902f
C5458 PAD.n6049 VSS 0.074902f
C5459 PAD.n6052 VSS 0.074902f
C5460 PAD.n6055 VSS 0.074902f
C5461 PAD.n6058 VSS 0.074902f
C5462 PAD.n6061 VSS 0.074902f
C5463 PAD.n6064 VSS 0.074902f
C5464 PAD.n6067 VSS 0.074902f
C5465 PAD.n6070 VSS 0.074902f
C5466 PAD.n6073 VSS 0.074902f
C5467 PAD.n6076 VSS 0.074902f
C5468 PAD.n6079 VSS 0.074902f
C5469 PAD.n6082 VSS 0.074902f
C5470 PAD.n6085 VSS 0.074902f
C5471 PAD.n6088 VSS 0.074902f
C5472 PAD.n6091 VSS 0.074902f
C5473 PAD.n6094 VSS 0.074902f
C5474 PAD.n6097 VSS 0.074902f
C5475 PAD.n6100 VSS 0.074902f
C5476 PAD.n6103 VSS 0.074902f
C5477 PAD.n6106 VSS 0.074902f
C5478 PAD.n6109 VSS 0.074902f
C5479 PAD.n6112 VSS 0.074902f
C5480 PAD.n6115 VSS 0.074902f
C5481 PAD.n6118 VSS 0.074902f
C5482 PAD.n6121 VSS 0.074902f
C5483 PAD.n6124 VSS 0.074902f
C5484 PAD.n6127 VSS 0.074902f
C5485 PAD.n6130 VSS 0.074902f
C5486 PAD.n6133 VSS 0.074902f
C5487 PAD.n6136 VSS 0.074902f
C5488 PAD.n6139 VSS 0.074902f
C5489 PAD.n6142 VSS 0.074902f
C5490 PAD.n6145 VSS 0.074902f
C5491 PAD.n6148 VSS 0.074902f
C5492 PAD.n6151 VSS 0.074902f
C5493 PAD.n6154 VSS 0.074902f
C5494 PAD.n6157 VSS 0.074902f
C5495 PAD.n6160 VSS 0.074902f
C5496 PAD.n6163 VSS 0.074902f
C5497 PAD.n6166 VSS 0.074902f
C5498 PAD.n6169 VSS 0.074902f
C5499 PAD.n6172 VSS 0.074902f
C5500 PAD.n6175 VSS 0.074902f
C5501 PAD.n6177 VSS 0.074902f
C5502 PAD.n6178 VSS 0.074902f
C5503 PAD.n6179 VSS 0.074902f
C5504 PAD.n6180 VSS 0.074902f
C5505 PAD.n6181 VSS 0.074902f
C5506 PAD.n6182 VSS 0.074902f
C5507 PAD.n6183 VSS 0.074902f
C5508 PAD.n6184 VSS 0.074902f
C5509 PAD.n6185 VSS 0.074902f
C5510 PAD.n6186 VSS 0.074902f
C5511 PAD.n6187 VSS 0.074902f
C5512 PAD.n6188 VSS 0.074902f
C5513 PAD.n6189 VSS 0.074902f
C5514 PAD.n6190 VSS 0.074902f
C5515 PAD.n6191 VSS 0.074902f
C5516 PAD.n6192 VSS 0.074902f
C5517 PAD.n6193 VSS 0.074902f
C5518 PAD.n6194 VSS 0.074902f
C5519 PAD.n6195 VSS 0.074902f
C5520 PAD.n6196 VSS 0.074902f
C5521 PAD.n6197 VSS 0.074902f
C5522 PAD.n6198 VSS 0.074902f
C5523 PAD.n6199 VSS 0.074902f
C5524 PAD.n6200 VSS 0.074902f
C5525 PAD.n6201 VSS 0.074902f
C5526 PAD.n6202 VSS 0.074902f
C5527 PAD.n6203 VSS 0.074902f
C5528 PAD.n6204 VSS 0.074902f
C5529 PAD.n6205 VSS 0.074902f
C5530 PAD.n6206 VSS 0.074902f
C5531 PAD.n6207 VSS 0.074902f
C5532 PAD.n6208 VSS 0.074902f
C5533 PAD.n6209 VSS 0.074902f
C5534 PAD.n6210 VSS 0.074902f
C5535 PAD.n6211 VSS 0.074902f
C5536 PAD.n6212 VSS 0.074902f
C5537 PAD.n6213 VSS 0.074902f
C5538 PAD.n6214 VSS 0.074902f
C5539 PAD.n6215 VSS 0.074902f
C5540 PAD.n6216 VSS 0.074902f
C5541 PAD.n6217 VSS 0.074902f
C5542 PAD.n6218 VSS 0.074902f
C5543 PAD.n6219 VSS 0.074902f
C5544 PAD.n6220 VSS 0.074902f
C5545 PAD.n6221 VSS 0.074902f
C5546 PAD.n6222 VSS 0.074902f
C5547 PAD.n6223 VSS 0.074902f
C5548 PAD.n6224 VSS 0.074902f
C5549 PAD.n6225 VSS 0.103594f
C5550 PAD.n6226 VSS 0.103594f
C5551 PAD.n6227 VSS 0.074902f
C5552 PAD.n6228 VSS 0.074902f
C5553 PAD.n6229 VSS 0.074902f
C5554 PAD.n6230 VSS 0.074902f
C5555 PAD.n6231 VSS 0.074902f
C5556 PAD.n6232 VSS 0.074902f
C5557 PAD.n6233 VSS 0.074902f
C5558 PAD.n6234 VSS 0.074902f
C5559 PAD.n6235 VSS 0.074902f
C5560 PAD.n6236 VSS 0.074902f
C5561 PAD.n6237 VSS 0.074902f
C5562 PAD.n6238 VSS 0.074902f
C5563 PAD.n6239 VSS 0.074902f
C5564 PAD.n6240 VSS 0.074902f
C5565 PAD.n6241 VSS 0.074902f
C5566 PAD.n6242 VSS 0.074902f
C5567 PAD.n6243 VSS 0.074902f
C5568 PAD.n6244 VSS 0.074902f
C5569 PAD.n6245 VSS 0.074902f
C5570 PAD.n6246 VSS 0.074902f
C5571 PAD.n6247 VSS 0.074902f
C5572 PAD.n6248 VSS 0.074902f
C5573 PAD.n6249 VSS 0.074902f
C5574 PAD.n6250 VSS 0.074902f
C5575 PAD.n6251 VSS 0.074902f
C5576 PAD.n6252 VSS 0.074902f
C5577 PAD.n6253 VSS 0.074902f
C5578 PAD.n6254 VSS 0.074902f
C5579 PAD.n6255 VSS 0.074902f
C5580 PAD.n6256 VSS 0.074902f
C5581 PAD.n6257 VSS 0.074902f
C5582 PAD.n6258 VSS 0.074902f
C5583 PAD.n6259 VSS 0.074902f
C5584 PAD.n6260 VSS 0.074902f
C5585 PAD.n6261 VSS 0.074902f
C5586 PAD.n6262 VSS 0.074902f
C5587 PAD.n6263 VSS 0.074902f
C5588 PAD.n6264 VSS 0.074902f
C5589 PAD.n6265 VSS 0.074902f
C5590 PAD.n6266 VSS 0.074902f
C5591 PAD.n6267 VSS 0.074902f
C5592 PAD.n6268 VSS 0.074902f
C5593 PAD.n6269 VSS 0.074902f
C5594 PAD.n6270 VSS 0.074902f
C5595 PAD.n6271 VSS 0.074902f
C5596 PAD.n6272 VSS 0.074902f
C5597 PAD.n6273 VSS 0.074902f
C5598 PAD.n6274 VSS 0.074902f
C5599 PAD.n6275 VSS 0.074902f
C5600 PAD.n6276 VSS 0.074902f
C5601 PAD.n6277 VSS 0.074902f
C5602 PAD.n6278 VSS 0.074902f
C5603 PAD.n6279 VSS 0.074902f
C5604 PAD.n6280 VSS 0.074902f
C5605 PAD.n6281 VSS 0.074902f
C5606 PAD.n6282 VSS 0.074902f
C5607 PAD.n6283 VSS 0.074902f
C5608 PAD.n6284 VSS 0.074902f
C5609 PAD.n6285 VSS 0.074902f
C5610 PAD.n6286 VSS 0.074902f
C5611 PAD.n6287 VSS 0.074902f
C5612 PAD.n6288 VSS 0.074902f
C5613 PAD.n6289 VSS 0.074902f
C5614 PAD.n6290 VSS 0.074902f
C5615 PAD.n6291 VSS 0.074902f
C5616 PAD.n6292 VSS 0.074902f
C5617 PAD.n6293 VSS 0.074902f
C5618 PAD.n6294 VSS 0.074902f
C5619 PAD.n6295 VSS 0.074902f
C5620 PAD.n6296 VSS 0.074902f
C5621 PAD.n6297 VSS 0.074902f
C5622 PAD.n6298 VSS 0.074902f
C5623 PAD.n6299 VSS 0.074902f
C5624 PAD.n6300 VSS 0.074902f
C5625 PAD.n6301 VSS 0.074902f
C5626 PAD.n6302 VSS 0.074902f
C5627 PAD.n6303 VSS 0.074902f
C5628 PAD.n6304 VSS 0.074902f
C5629 PAD.n6305 VSS 0.074902f
C5630 PAD.n6306 VSS 0.074902f
C5631 PAD.n6307 VSS 0.074902f
C5632 PAD.n6308 VSS 0.074902f
C5633 PAD.n6309 VSS 0.074902f
C5634 PAD.n6310 VSS 0.074902f
C5635 PAD.n6311 VSS 0.074902f
C5636 PAD.n6312 VSS 0.074902f
C5637 PAD.n6313 VSS 0.074902f
C5638 PAD.n6314 VSS 0.074902f
C5639 PAD.n6315 VSS 0.074902f
C5640 PAD.n6316 VSS 0.074902f
C5641 PAD.n6317 VSS 0.074902f
C5642 PAD.n6318 VSS 0.074902f
C5643 PAD.n6319 VSS 0.074902f
C5644 PAD.n6320 VSS 0.074902f
C5645 PAD.n6321 VSS 0.074902f
C5646 PAD.n6322 VSS 0.074902f
C5647 PAD.n6323 VSS 0.074902f
C5648 PAD.n6324 VSS 0.074902f
C5649 PAD.n6325 VSS 0.074902f
C5650 PAD.n6326 VSS 0.074902f
C5651 PAD.n6327 VSS 0.074902f
C5652 PAD.n6328 VSS 0.074902f
C5653 PAD.n6329 VSS 0.074902f
C5654 PAD.n6330 VSS 0.074902f
C5655 PAD.n6331 VSS 0.074902f
C5656 PAD.n6332 VSS 0.074902f
C5657 PAD.n6333 VSS 0.074902f
C5658 PAD.n6334 VSS 0.074902f
C5659 PAD.n6335 VSS 0.074902f
C5660 PAD.n6336 VSS 0.074902f
C5661 PAD.n6337 VSS 0.074902f
C5662 PAD.n6338 VSS 0.074902f
C5663 PAD.n6339 VSS 0.074902f
C5664 PAD.n6340 VSS 0.074902f
C5665 PAD.n6341 VSS 0.074902f
C5666 PAD.n6342 VSS 0.074902f
C5667 PAD.n6343 VSS 0.074902f
C5668 PAD.n6344 VSS 0.074902f
C5669 PAD.n6345 VSS 0.074902f
C5670 PAD.n6346 VSS 0.074902f
C5671 PAD.n6347 VSS 0.074902f
C5672 PAD.n6348 VSS 0.074902f
C5673 PAD.n6349 VSS 0.074902f
C5674 PAD.n6350 VSS 0.074902f
C5675 PAD.n6351 VSS 0.074902f
C5676 PAD.n6352 VSS 0.074902f
C5677 PAD.n6353 VSS 0.074902f
C5678 PAD.n6354 VSS 0.074902f
C5679 PAD.n6355 VSS 0.074902f
C5680 PAD.n6356 VSS 0.074902f
C5681 PAD.n6357 VSS 0.074902f
C5682 PAD.n6358 VSS 0.074902f
C5683 PAD.n6359 VSS 0.074902f
C5684 PAD.n6360 VSS 0.074902f
C5685 PAD.n6361 VSS 0.074902f
C5686 PAD.n6362 VSS 0.074902f
C5687 PAD.n6363 VSS 0.074902f
C5688 PAD.n6364 VSS 0.074902f
C5689 PAD.n6365 VSS 0.074902f
C5690 PAD.n6366 VSS 0.074902f
C5691 PAD.n6367 VSS 0.074902f
C5692 PAD.n6368 VSS 0.074902f
C5693 PAD.n6369 VSS 0.074902f
C5694 PAD.n6370 VSS 0.074902f
C5695 PAD.n6371 VSS 0.059499f
C5696 PAD.n6372 VSS 0.059499f
C5697 PAD.n6373 VSS 1.51918f
C5698 PAD.n6374 VSS 0.122923f
C5699 PAD.n6375 VSS 0.123237f
C5700 PAD.n6376 VSS 0.155682f
C5701 PAD.n6377 VSS 0.033766f
C5702 PAD.n6378 VSS 0.028843f
C5703 PAD.n6379 VSS 0.042887f
C5704 PAD.n6380 VSS 0.025823f
C5705 PAD.n6381 VSS 0.029567f
C5706 PAD.n6382 VSS 0.029567f
C5707 PAD.n6383 VSS 0.611619f
C5708 PAD.n6385 VSS 0.125801f
C5709 PAD.n6386 VSS 0.863173f
C5710 PAD.n6387 VSS 0.043189f
C5711 PAD.n6388 VSS 0.043189f
C5712 PAD.n6389 VSS 0.05527f
C5713 PAD.n6390 VSS 0.238879f
C5714 PAD.n6391 VSS 0.056739f
C5715 PAD.n6392 VSS 0.062262f
C5716 PAD.n6393 VSS 0.069752f
C5717 PAD.n6394 VSS 0.038251f
C5718 PAD.n6395 VSS 0.038251f
C5719 PAD.n6396 VSS 0.582025f
C5720 PAD.n6436 VSS 0.036454f
C5721 PAD.n6437 VSS 0.036454f
C5722 PAD.n6438 VSS 0.036454f
C5723 PAD.n6439 VSS 0.036454f
C5724 PAD.n6440 VSS 0.036454f
C5725 PAD.n6441 VSS 0.036454f
C5726 PAD.n6442 VSS 0.036454f
C5727 PAD.n6443 VSS 0.036454f
C5728 PAD.n6444 VSS 0.036454f
C5729 PAD.n6445 VSS 0.036454f
C5730 PAD.n6446 VSS 0.036454f
C5731 PAD.n6447 VSS 0.036454f
C5732 PAD.n6448 VSS 0.036454f
C5733 PAD.n6449 VSS 0.036454f
C5734 PAD.n6450 VSS 0.036454f
C5735 PAD.n6451 VSS 0.036454f
C5736 PAD.n6452 VSS 0.036454f
C5737 PAD.n6453 VSS 0.036454f
C5738 PAD.n6454 VSS 0.036454f
C5739 PAD.n6455 VSS 0.036454f
C5740 PAD.n6456 VSS 0.036454f
C5741 PAD.n6457 VSS 0.036454f
C5742 PAD.n6458 VSS 0.036454f
C5743 PAD.n6459 VSS 0.036454f
C5744 PAD.n6460 VSS 0.036454f
C5745 PAD.n6461 VSS 0.036454f
C5746 PAD.n6462 VSS 0.036454f
C5747 PAD.n6463 VSS 0.036454f
C5748 PAD.n6464 VSS 0.036454f
C5749 PAD.n6465 VSS 0.036454f
C5750 PAD.n6466 VSS 0.036454f
C5751 PAD.n6467 VSS 0.036454f
C5752 PAD.n6468 VSS 0.036454f
C5753 PAD.n6469 VSS 0.036454f
C5754 PAD.n6470 VSS 0.036454f
C5755 PAD.n6471 VSS 0.036454f
C5756 PAD.n6472 VSS 0.036454f
C5757 PAD.n6473 VSS 0.036454f
C5758 PAD.n6474 VSS 0.036454f
C5759 PAD.n6475 VSS 0.036454f
C5760 PAD.n6476 VSS 0.036454f
C5761 PAD.n6477 VSS 0.036454f
C5762 PAD.n6478 VSS 0.036454f
C5763 PAD.n6479 VSS 0.036454f
C5764 PAD.n6480 VSS 0.036454f
C5765 PAD.n6481 VSS 0.036454f
C5766 PAD.n6482 VSS 0.036454f
C5767 PAD.n6483 VSS 0.036454f
C5768 PAD.n6484 VSS 0.036454f
C5769 PAD.n6485 VSS 0.036454f
C5770 PAD.n6486 VSS 0.036454f
C5771 PAD.n6487 VSS 0.036454f
C5772 PAD.n6488 VSS 0.036454f
C5773 PAD.n6489 VSS 0.036454f
C5774 PAD.n6490 VSS 0.036454f
C5775 PAD.n6491 VSS 0.036454f
C5776 PAD.n6492 VSS 0.036454f
C5777 PAD.n6493 VSS 0.036454f
C5778 PAD.n6494 VSS 0.036454f
C5779 PAD.n6495 VSS 0.036454f
C5780 PAD.n6496 VSS 0.036454f
C5781 PAD.n6497 VSS 0.036454f
C5782 PAD.n6498 VSS 0.036454f
C5783 PAD.n6499 VSS 0.036454f
C5784 PAD.n6500 VSS 0.036454f
C5785 PAD.n6501 VSS 0.036454f
C5786 PAD.n6502 VSS 0.036454f
C5787 PAD.n6503 VSS 0.036454f
C5788 PAD.n6504 VSS 0.036454f
C5789 PAD.n6505 VSS 0.036454f
C5790 PAD.n6506 VSS 0.036454f
C5791 PAD.n6507 VSS 0.036454f
C5792 PAD.n6508 VSS 0.036454f
C5793 PAD.n6509 VSS 0.036454f
C5794 PAD.n6510 VSS 0.036454f
C5795 PAD.n6511 VSS 0.036454f
C5796 PAD.n6512 VSS 0.036454f
C5797 PAD.n6513 VSS 0.036454f
C5798 PAD.n6514 VSS 0.036454f
C5799 PAD.n6515 VSS 0.036454f
C5800 PAD.n6516 VSS 0.036454f
C5801 PAD.n6517 VSS 0.036454f
C5802 PAD.n6518 VSS 0.036454f
C5803 PAD.n6519 VSS 0.036454f
C5804 PAD.n6520 VSS 0.036454f
C5805 PAD.n6521 VSS 0.036454f
C5806 PAD.n6522 VSS 0.036454f
C5807 PAD.n6523 VSS 0.036454f
C5808 PAD.n6524 VSS 0.036454f
C5809 PAD.n6525 VSS 0.036454f
C5810 PAD.n6526 VSS 0.036454f
C5811 PAD.n6527 VSS 0.036454f
C5812 PAD.n6528 VSS 0.036454f
C5813 PAD.n6529 VSS 0.036454f
C5814 PAD.n6530 VSS 0.036454f
C5815 PAD.n6531 VSS 0.036454f
C5816 PAD.n6532 VSS 0.036454f
C5817 PAD.n6533 VSS 0.036454f
C5818 PAD.n6534 VSS 0.036454f
C5819 PAD.n6535 VSS 0.036454f
C5820 PAD.n6536 VSS 0.036454f
C5821 PAD.n6537 VSS 0.036454f
C5822 PAD.n6538 VSS 0.036454f
C5823 PAD.n6539 VSS 0.036454f
C5824 PAD.n6540 VSS 0.036454f
C5825 PAD.n6541 VSS 0.036454f
C5826 PAD.n6542 VSS 0.036454f
C5827 PAD.n6543 VSS 0.036454f
C5828 PAD.n6544 VSS 0.036454f
C5829 PAD.n6545 VSS 0.036454f
C5830 PAD.n6546 VSS 0.036454f
C5831 PAD.n6547 VSS 0.036454f
C5832 PAD.n6548 VSS 0.036454f
C5833 PAD.n6549 VSS 0.036454f
C5834 PAD.n6550 VSS 0.036454f
C5835 PAD.n6551 VSS 0.036454f
C5836 PAD.n6552 VSS 0.036454f
C5837 PAD.n6553 VSS 0.036454f
C5838 PAD.n6554 VSS 0.036454f
C5839 PAD.n6555 VSS 0.036454f
C5840 PAD.n6556 VSS 0.036454f
C5841 PAD.n6557 VSS 0.036454f
C5842 PAD.n6558 VSS 0.036454f
C5843 PAD.n6559 VSS 0.036454f
C5844 PAD.n6560 VSS 0.036454f
C5845 PAD.n6561 VSS 0.036454f
C5846 PAD.n6562 VSS 0.036454f
C5847 PAD.n6563 VSS 0.036454f
C5848 PAD.n6564 VSS 0.036454f
C5849 PAD.n6565 VSS 0.036454f
C5850 PAD.n6566 VSS 0.036454f
C5851 PAD.n6567 VSS 0.036454f
C5852 PAD.n6568 VSS 0.036454f
C5853 PAD.n6569 VSS 0.036454f
C5854 PAD.n6570 VSS 0.036454f
C5855 PAD.n6571 VSS 0.036454f
C5856 PAD.n6572 VSS 0.036454f
C5857 PAD.n6573 VSS 0.036454f
C5858 PAD.n6574 VSS 0.036454f
C5859 PAD.n6575 VSS 0.036454f
C5860 PAD.n6576 VSS 0.036454f
C5861 PAD.n6577 VSS 0.036454f
C5862 PAD.n6578 VSS 0.036454f
C5863 PAD.n6579 VSS 0.036454f
C5864 PAD.n6580 VSS 0.036454f
C5865 PAD.n6581 VSS 0.036454f
C5866 PAD.n6582 VSS 0.036454f
C5867 PAD.n6583 VSS 0.036454f
C5868 PAD.n6584 VSS 0.036454f
C5869 PAD.n6585 VSS 0.036454f
C5870 PAD.n6586 VSS 0.036454f
C5871 PAD.n6587 VSS 0.036454f
C5872 PAD.n6588 VSS 0.036454f
C5873 PAD.n6589 VSS 0.036454f
C5874 PAD.n6590 VSS 0.036454f
C5875 PAD.n6591 VSS 0.036454f
C5876 PAD.n6592 VSS 0.036454f
C5877 PAD.n6593 VSS 0.036454f
C5878 PAD.n6594 VSS 0.036454f
C5879 PAD.n6595 VSS 0.036454f
C5880 PAD.n6596 VSS 0.036454f
C5881 PAD.n6597 VSS 0.036454f
C5882 PAD.n6598 VSS 0.036454f
C5883 PAD.n6599 VSS 0.036454f
C5884 PAD.n6600 VSS 0.036454f
C5885 PAD.n6601 VSS 0.036454f
C5886 PAD.n6602 VSS 0.036454f
C5887 PAD.n6603 VSS 0.036454f
C5888 PAD.n6604 VSS 0.036454f
C5889 PAD.n6605 VSS 0.036454f
C5890 PAD.n6606 VSS 0.036454f
C5891 PAD.n6607 VSS 0.036454f
C5892 PAD.n6608 VSS 0.036454f
C5893 PAD.n6609 VSS 0.036454f
C5894 PAD.n6610 VSS 0.036454f
C5895 PAD.n6611 VSS 0.036454f
C5896 PAD.n6612 VSS 0.036454f
C5897 PAD.n6613 VSS 0.036454f
C5898 PAD.n6614 VSS 0.036454f
C5899 PAD.n6615 VSS 0.036454f
C5900 PAD.n6616 VSS 0.036454f
C5901 PAD.n6617 VSS 0.036454f
C5902 PAD.n6618 VSS 0.036454f
C5903 PAD.n6619 VSS 0.036454f
C5904 PAD.n6620 VSS 0.036454f
C5905 PAD.n6621 VSS 0.036454f
C5906 PAD.n6622 VSS 0.036454f
C5907 PAD.n6623 VSS 0.036454f
C5908 PAD.n6624 VSS 0.036454f
C5909 PAD.n6625 VSS 0.036454f
C5910 PAD.n6626 VSS 0.036454f
C5911 PAD.n6627 VSS 0.036454f
C5912 PAD.n6628 VSS 0.036454f
C5913 PAD.n6629 VSS 0.036454f
C5914 PAD.n6630 VSS 0.036454f
C5915 PAD.n6631 VSS 0.036454f
C5916 PAD.n6632 VSS 0.036454f
C5917 PAD.n6633 VSS 0.036454f
C5918 PAD.n6634 VSS 0.036454f
C5919 PAD.n6635 VSS 0.036454f
C5920 PAD.n6636 VSS 0.036454f
C5921 PAD.n6637 VSS 0.036454f
C5922 PAD.n6638 VSS 0.036454f
C5923 PAD.n6639 VSS 0.036454f
C5924 PAD.n6640 VSS 0.036454f
C5925 PAD.n6641 VSS 0.036454f
C5926 PAD.n6642 VSS 0.036454f
C5927 PAD.n6643 VSS 0.036454f
C5928 PAD.n6644 VSS 0.036454f
C5929 PAD.n6645 VSS 0.036454f
C5930 PAD.n6646 VSS 0.036454f
C5931 PAD.n6647 VSS 0.036454f
C5932 PAD.n6648 VSS 0.036454f
C5933 PAD.n6649 VSS 0.036454f
C5934 PAD.n6650 VSS 0.036454f
C5935 PAD.n6651 VSS 0.036454f
C5936 PAD.n6652 VSS 0.036454f
C5937 PAD.n6653 VSS 0.036454f
C5938 PAD.n6654 VSS 0.036454f
C5939 PAD.n6655 VSS 0.036454f
C5940 PAD.n6656 VSS 0.036454f
C5941 PAD.n6657 VSS 0.036454f
C5942 PAD.n6658 VSS 0.036454f
C5943 PAD.n6659 VSS 0.036454f
C5944 PAD.n6660 VSS 0.036454f
C5945 PAD.n6661 VSS 0.036454f
C5946 PAD.n6662 VSS 0.036454f
C5947 PAD.n6663 VSS 0.036454f
C5948 PAD.n6664 VSS 0.036454f
C5949 PAD.n6665 VSS 0.036454f
C5950 PAD.n6666 VSS 0.036454f
C5951 PAD.n6667 VSS 0.036454f
C5952 PAD.n6668 VSS 0.036454f
C5953 PAD.n6669 VSS 0.036454f
C5954 PAD.n6670 VSS 0.036454f
C5955 PAD.n6671 VSS 0.036454f
C5956 PAD.n6672 VSS 0.036454f
C5957 PAD.n6673 VSS 0.036454f
C5958 PAD.n6674 VSS 0.036454f
C5959 PAD.n6675 VSS 0.036454f
C5960 PAD.n6676 VSS 0.036454f
C5961 PAD.n6678 VSS 0.517904f
C5962 PAD.n6679 VSS 0.478444f
C5963 PAD.n6680 VSS 0.611619f
C5964 PAD.n6681 VSS 0.066377f
C5965 PAD.n6682 VSS 0.700403f
C5966 PAD.n6683 VSS 0.212094f
C5967 PAD.n6684 VSS 0.040633f
C5968 PAD.n6685 VSS 0.040633f
C5969 PAD.n6686 VSS 0.029431f
C5970 PAD.n6687 VSS 0.023105f
C5971 PAD.n6688 VSS 0.023105f
C5972 PAD.n6689 VSS 0.42912f
C5973 PAD.n6690 VSS 0.023105f
C5974 PAD.n6691 VSS 0.023105f
C5975 PAD.n6692 VSS 0.033374f
C5976 PAD.n6693 VSS 0.046278f
C5977 PAD.n6694 VSS 0.059249f
C5978 PAD.n6695 VSS 0.062262f
C5979 PAD.n6696 VSS 0.069752f
C5980 PAD.n6697 VSS 0.046126f
C5981 PAD.n6698 VSS 0.046126f
C5982 PAD.n6699 VSS 0.221958f
C5983 PAD.n6700 VSS 0.562295f
C5984 PAD.n6701 VSS 0.02853f
C5985 PAD.n6702 VSS 0.02853f
C5986 PAD.n6703 VSS 0.024917f
C5987 PAD.n6704 VSS 0.033766f
C5988 PAD.n6705 VSS 0.03055f
C5989 PAD.n6706 VSS 0.042887f
C5990 PAD.n6707 VSS 0.029431f
C5991 PAD.n6708 VSS 0.049106f
C5992 PAD.n6709 VSS 0.029431f
C5993 PAD.n6710 VSS 0.049106f
C5994 PAD.n6711 VSS 0.611619f
C5995 PAD.n6712 VSS 0.700403f
C5996 PAD.n6713 VSS 0.438985f
C5997 PAD.n6714 VSS 0.039754f
C5998 PAD.n6715 VSS 0.069752f
C5999 PAD.n6716 VSS 0.039754f
C6000 PAD.n6717 VSS 0.069752f
C6001 PAD.n6718 VSS 0.036454f
C6002 PAD.n6719 VSS 0.023105f
C6003 PAD.n6720 VSS 0.036454f
C6004 PAD.n6723 VSS 0.036454f
C6005 PAD.n6724 VSS 0.036454f
C6006 PAD.n6725 VSS 0.036454f
C6007 PAD.n6726 VSS 0.036454f
C6008 PAD.n6728 VSS 0.036454f
C6009 PAD.n6729 VSS 0.036454f
C6010 PAD.n6730 VSS 0.036454f
C6011 PAD.n6732 VSS 0.036454f
C6012 PAD.n6733 VSS 0.036454f
C6013 PAD.n6734 VSS 0.036454f
C6014 PAD.n6736 VSS 0.036454f
C6015 PAD.n6737 VSS 0.036454f
C6016 PAD.n6738 VSS 0.036454f
C6017 PAD.n6740 VSS 0.036454f
C6018 PAD.n6741 VSS 0.036454f
C6019 PAD.n6742 VSS 0.036454f
C6020 PAD.n6744 VSS 0.036454f
C6021 PAD.n6745 VSS 0.036454f
C6022 PAD.n6746 VSS 0.036454f
C6023 PAD.n6748 VSS 0.036454f
C6024 PAD.n6749 VSS 0.036454f
C6025 PAD.n6750 VSS 0.036454f
C6026 PAD.n6752 VSS 0.036454f
C6027 PAD.n6753 VSS 0.036454f
C6028 PAD.n6754 VSS 0.036454f
C6029 PAD.n6756 VSS 0.036454f
C6030 PAD.n6757 VSS 0.036454f
C6031 PAD.n6758 VSS 0.036454f
C6032 PAD.n6760 VSS 0.036454f
C6033 PAD.n6761 VSS 0.036454f
C6034 PAD.n6762 VSS 0.036454f
C6035 PAD.n6764 VSS 0.036454f
C6036 PAD.n6765 VSS 0.036454f
C6037 PAD.n6766 VSS 0.036454f
C6038 PAD.n6768 VSS 0.036454f
C6039 PAD.n6769 VSS 0.036454f
C6040 PAD.n6770 VSS 0.036454f
C6041 PAD.n6772 VSS 0.036454f
C6042 PAD.n6773 VSS 0.036454f
C6043 PAD.n6774 VSS 0.036454f
C6044 PAD.n6776 VSS 0.036454f
C6045 PAD.n6777 VSS 0.036454f
C6046 PAD.n6778 VSS 0.036454f
C6047 PAD.n6780 VSS 0.036454f
C6048 PAD.n6781 VSS 0.036454f
C6049 PAD.n6782 VSS 0.036454f
C6050 PAD.n6784 VSS 0.036454f
C6051 PAD.n6785 VSS 0.036454f
C6052 PAD.n6786 VSS 0.036454f
C6053 PAD.n6788 VSS 0.036454f
C6054 PAD.n6789 VSS 0.036454f
C6055 PAD.n6790 VSS 0.036454f
C6056 PAD.n6792 VSS 0.036454f
C6057 PAD.n6793 VSS 0.036454f
C6058 PAD.n6794 VSS 0.036454f
C6059 PAD.n6796 VSS 0.036454f
C6060 PAD.n6797 VSS 0.036454f
C6061 PAD.n6798 VSS 0.036454f
C6062 PAD.n6800 VSS 0.036454f
C6063 PAD.n6801 VSS 0.036454f
C6064 PAD.n6802 VSS 0.036454f
C6065 PAD.n6803 VSS 0.023105f
C6066 PAD.n6804 VSS 0.023105f
C6067 PAD.n6806 VSS 0.036454f
C6068 PAD.n6808 VSS 0.036454f
C6069 PAD.n6810 VSS 0.036454f
C6070 PAD.n6811 VSS 0.036454f
C6071 PAD.n6812 VSS 0.036454f
C6072 PAD.n6813 VSS 0.036454f
C6073 PAD.n6814 VSS 0.036454f
C6074 PAD.n6815 VSS 0.036454f
C6075 PAD.n6816 VSS 0.036454f
C6076 PAD.n6818 VSS 0.036454f
C6077 PAD.n6820 VSS 0.036454f
C6078 PAD.n6822 VSS 0.036454f
C6079 PAD.n6823 VSS 0.036454f
C6080 PAD.n6824 VSS 0.036454f
C6081 PAD.n6825 VSS 0.036454f
C6082 PAD.n6826 VSS 0.036454f
C6083 PAD.n6827 VSS 0.036454f
C6084 PAD.n6828 VSS 0.036454f
C6085 PAD.n6830 VSS 0.036454f
C6086 PAD.n6832 VSS 0.036454f
C6087 PAD.n6834 VSS 0.036454f
C6088 PAD.n6835 VSS 0.036454f
C6089 PAD.n6836 VSS 0.036454f
C6090 PAD.n6837 VSS 0.036454f
C6091 PAD.n6838 VSS 0.036454f
C6092 PAD.n6839 VSS 0.036454f
C6093 PAD.n6840 VSS 0.036454f
C6094 PAD.n6842 VSS 0.036454f
C6095 PAD.n6844 VSS 0.036454f
C6096 PAD.n6846 VSS 0.036454f
C6097 PAD.n6847 VSS 0.036454f
C6098 PAD.n6848 VSS 0.036454f
C6099 PAD.n6849 VSS 0.036454f
C6100 PAD.n6850 VSS 0.036454f
C6101 PAD.n6851 VSS 0.036454f
C6102 PAD.n6852 VSS 0.036454f
C6103 PAD.n6854 VSS 0.036454f
C6104 PAD.n6856 VSS 0.036454f
C6105 PAD.n6858 VSS 0.036454f
C6106 PAD.n6859 VSS 0.036454f
C6107 PAD.n6860 VSS 0.036454f
C6108 PAD.n6861 VSS 0.036454f
C6109 PAD.n6862 VSS 0.036454f
C6110 PAD.n6863 VSS 0.036454f
C6111 PAD.n6864 VSS 0.036454f
C6112 PAD.n6866 VSS 0.036454f
C6113 PAD.n6868 VSS 0.036454f
C6114 PAD.n6870 VSS 0.036454f
C6115 PAD.n6871 VSS 0.036454f
C6116 PAD.n6872 VSS 0.036454f
C6117 PAD.n6873 VSS 0.036454f
C6118 PAD.n6874 VSS 0.036454f
C6119 PAD.n6875 VSS 0.036454f
C6120 PAD.n6876 VSS 0.036454f
C6121 PAD.n6878 VSS 0.036454f
C6122 PAD.n6880 VSS 0.036454f
C6123 PAD.n6882 VSS 0.036454f
C6124 PAD.n6883 VSS 0.036454f
C6125 PAD.n6884 VSS 0.036454f
C6126 PAD.n6885 VSS 0.036454f
C6127 PAD.n6886 VSS 0.036454f
C6128 PAD.n6887 VSS 0.036454f
C6129 PAD.n6888 VSS 0.036454f
C6130 PAD.n6890 VSS 0.036454f
C6131 PAD.n6892 VSS 0.036454f
C6132 PAD.n6894 VSS 0.036454f
C6133 PAD.n6895 VSS 0.036454f
C6134 PAD.n6896 VSS 0.036454f
C6135 PAD.n6897 VSS 0.036454f
C6136 PAD.n6898 VSS 0.036454f
C6137 PAD.n6899 VSS 0.036454f
C6138 PAD.n6900 VSS 0.036454f
C6139 PAD.n6902 VSS 0.036454f
C6140 PAD.n6904 VSS 0.036454f
C6141 PAD.n6906 VSS 0.036454f
C6142 PAD.n6907 VSS 0.036454f
C6143 PAD.n6908 VSS 0.036454f
C6144 PAD.n6909 VSS 0.036454f
C6145 PAD.n6910 VSS 0.036454f
C6146 PAD.n6911 VSS 0.036454f
C6147 PAD.n6912 VSS 0.036454f
C6148 PAD.n6914 VSS 0.036454f
C6149 PAD.n6916 VSS 0.036454f
C6150 PAD.n6918 VSS 0.036454f
C6151 PAD.n6919 VSS 0.036454f
C6152 PAD.n6920 VSS 0.036454f
C6153 PAD.n6921 VSS 0.036454f
C6154 PAD.n6922 VSS 0.036454f
C6155 PAD.n6923 VSS 0.036454f
C6156 PAD.n6924 VSS 0.036454f
C6157 PAD.n6926 VSS 0.036454f
C6158 PAD.n6928 VSS 0.036454f
C6159 PAD.n6930 VSS 0.036454f
C6160 PAD.n6931 VSS 0.036454f
C6161 PAD.n6932 VSS 0.036454f
C6162 PAD.n6933 VSS 0.036454f
C6163 PAD.n6934 VSS 0.036454f
C6164 PAD.n6935 VSS 0.036454f
C6165 PAD.n6936 VSS 0.036454f
C6166 PAD.n6938 VSS 0.036454f
C6167 PAD.n6940 VSS 0.036454f
C6168 PAD.n6942 VSS 0.036454f
C6169 PAD.n6943 VSS 0.036454f
C6170 PAD.n6944 VSS 0.036454f
C6171 PAD.n6945 VSS 0.036454f
C6172 PAD.n6946 VSS 0.036454f
C6173 PAD.n6947 VSS 0.036454f
C6174 PAD.n6948 VSS 0.036454f
C6175 PAD.n6950 VSS 0.036454f
C6176 PAD.n6952 VSS 0.036454f
C6177 PAD.n6954 VSS 0.036454f
C6178 PAD.n6955 VSS 0.036454f
C6179 PAD.n6956 VSS 0.036454f
C6180 PAD.n6957 VSS 0.036454f
C6181 PAD.n6958 VSS 0.036454f
C6182 PAD.n6959 VSS 0.036454f
C6183 PAD.n6960 VSS 0.036454f
C6184 PAD.n6962 VSS 0.036454f
C6185 PAD.n6964 VSS 0.036454f
C6186 PAD.n6966 VSS 0.036454f
C6187 PAD.n6967 VSS 0.036454f
C6188 PAD.n6968 VSS 0.036454f
C6189 PAD.n6969 VSS 0.036454f
C6190 PAD.n6970 VSS 0.036454f
C6191 PAD.n6971 VSS 0.036454f
C6192 PAD.n6972 VSS 0.036454f
C6193 PAD.n6974 VSS 0.036454f
C6194 PAD.n6976 VSS 0.036454f
C6195 PAD.n6978 VSS 0.036454f
C6196 PAD.n6979 VSS 0.036454f
C6197 PAD.n6980 VSS 0.036454f
C6198 PAD.n6981 VSS 0.036454f
C6199 PAD.n6982 VSS 0.036454f
C6200 PAD.n6983 VSS 0.036454f
C6201 PAD.n6984 VSS 0.036454f
C6202 PAD.n6986 VSS 0.036454f
C6203 PAD.n6988 VSS 0.036454f
C6204 PAD.n6990 VSS 0.036454f
C6205 PAD.n6991 VSS 0.036454f
C6206 PAD.n6992 VSS 0.036454f
C6207 PAD.n6993 VSS 0.036454f
C6208 PAD.n6994 VSS 0.036454f
C6209 PAD.n6995 VSS 0.036454f
C6210 PAD.n6996 VSS 0.036454f
C6211 PAD.n6998 VSS 0.036454f
C6212 PAD.n7000 VSS 0.036454f
C6213 PAD.n7002 VSS 0.036454f
C6214 PAD.n7003 VSS 0.036454f
C6215 PAD.n7004 VSS 0.036454f
C6216 PAD.n7005 VSS 0.036454f
C6217 PAD.n7006 VSS 0.036454f
C6218 PAD.n7007 VSS 0.036454f
C6219 PAD.n7008 VSS 0.036454f
C6220 PAD.n7010 VSS 0.036454f
C6221 PAD.n7012 VSS 0.036454f
C6222 PAD.n7014 VSS 0.036454f
C6223 PAD.n7015 VSS 0.036454f
C6224 PAD.n7016 VSS 0.036454f
C6225 PAD.n7017 VSS 0.036454f
C6226 PAD.n7018 VSS 0.036454f
C6227 PAD.n7019 VSS 0.036454f
C6228 PAD.n7020 VSS 0.036454f
C6229 PAD.n7022 VSS 0.036454f
C6230 PAD.n7024 VSS 0.036454f
C6231 PAD.n7026 VSS 0.036454f
C6232 PAD.n7027 VSS 0.036454f
C6233 PAD.n7028 VSS 0.036454f
C6234 PAD.n7029 VSS 0.036454f
C6235 PAD.n7030 VSS 0.036454f
C6236 PAD.n7031 VSS 0.036454f
C6237 PAD.n7032 VSS 0.036454f
C6238 PAD.n7034 VSS 0.036454f
C6239 PAD.n7036 VSS 0.036454f
C6240 PAD.n7038 VSS 0.036454f
C6241 PAD.n7039 VSS 0.036454f
C6242 PAD.n7040 VSS 0.036454f
C6243 PAD.n7041 VSS 0.036454f
C6244 PAD.n7042 VSS 0.036454f
C6245 PAD.n7043 VSS 0.036454f
C6246 PAD.n7044 VSS 0.036454f
C6247 PAD.n7046 VSS 0.036454f
C6248 PAD.n7048 VSS 0.036454f
C6249 PAD.n7049 VSS 0.036454f
C6250 PAD.n7050 VSS 0.023105f
C6251 PAD.n7051 VSS 0.033374f
C6252 PAD.n7052 VSS 0.054002f
C6253 PAD.n7053 VSS 0.054002f
C6254 PAD.n7054 VSS 0.048203f
C6255 PAD.n7055 VSS 0.046278f
C6256 PAD.n7056 VSS 0.046278f
C6257 PAD.n7057 VSS 0.039754f
C6258 PAD.n7058 VSS 0.039754f
C6259 PAD.n7059 VSS 0.522836f
C6260 PAD.n7060 VSS 0.700403f
C6261 PAD.n7061 VSS 0.611619f
C6262 PAD.n7103 VSS 0.453782f
C6263 PAD.n7104 VSS 0.036454f
C6264 PAD.n7105 VSS 0.606687f
C6265 PAD.n7106 VSS 0.036454f
C6266 PAD.n7107 VSS 0.036454f
C6267 PAD.n7108 VSS 0.036454f
C6268 PAD.n7109 VSS 0.036454f
C6269 PAD.n7110 VSS 0.036454f
C6270 PAD.n7111 VSS 0.036454f
C6271 PAD.n7112 VSS 0.036454f
C6272 PAD.n7113 VSS 0.036454f
C6273 PAD.n7114 VSS 0.036454f
C6274 PAD.n7115 VSS 0.036454f
C6275 PAD.n7116 VSS 0.036454f
C6276 PAD.n7117 VSS 0.036454f
C6277 PAD.n7118 VSS 0.036454f
C6278 PAD.n7119 VSS 0.036454f
C6279 PAD.n7120 VSS 0.036454f
C6280 PAD.n7121 VSS 0.036454f
C6281 PAD.n7122 VSS 0.036454f
C6282 PAD.n7123 VSS 0.036454f
C6283 PAD.n7124 VSS 0.036454f
C6284 PAD.n7125 VSS 0.036454f
C6285 PAD.n7126 VSS 0.036454f
C6286 PAD.n7127 VSS 0.036454f
C6287 PAD.n7128 VSS 0.036454f
C6288 PAD.n7129 VSS 0.036454f
C6289 PAD.n7130 VSS 0.036454f
C6290 PAD.n7131 VSS 0.036454f
C6291 PAD.n7132 VSS 0.036454f
C6292 PAD.n7133 VSS 0.036454f
C6293 PAD.n7134 VSS 0.036454f
C6294 PAD.n7135 VSS 0.036454f
C6295 PAD.n7136 VSS 0.036454f
C6296 PAD.n7137 VSS 0.036454f
C6297 PAD.n7138 VSS 0.036454f
C6298 PAD.n7139 VSS 0.036454f
C6299 PAD.n7140 VSS 0.036454f
C6300 PAD.n7141 VSS 0.036454f
C6301 PAD.n7142 VSS 0.036454f
C6302 PAD.n7143 VSS 0.036454f
C6303 PAD.n7144 VSS 0.036454f
C6304 PAD.n7145 VSS 0.036454f
C6305 PAD.n7146 VSS 0.036454f
C6306 PAD.n7147 VSS 0.03055f
C6307 PAD.n7148 VSS 0.029431f
C6308 PAD.n7149 VSS 0.044092f
C6309 PAD.n7150 VSS 0.049106f
C6310 PAD.n7151 VSS 0.049106f
C6311 PAD.n7152 VSS 0.044092f
C6312 PAD.n7153 VSS 0.038508f
C6313 PAD.n7154 VSS 0.033766f
C6314 PAD.n7155 VSS 0.033766f
C6315 PAD.n7156 VSS 0.029431f
C6316 PAD.n7157 VSS 0.029431f
C6317 PAD.n7158 VSS 0.700403f
C6318 PAD.n7200 VSS 0.596822f
C6319 PAD.n7201 VSS 0.036454f
C6320 PAD.n7202 VSS 0.07463f
C6321 PAD.n7203 VSS 0.029749f
C6322 PAD.n7204 VSS 0.034063f
C6323 PAD.n7205 VSS 0.034063f
C6324 PAD.n7206 VSS 0.374863f
C6325 PAD.n7207 VSS 0.340336f
C6326 PAD.n7208 VSS 0.07463f
C6327 PAD.n7209 VSS 0.036454f
C6328 PAD.n7210 VSS 0.062262f
C6329 PAD.n7211 VSS 0.069752f
C6330 PAD.n7212 VSS 0.038161f
C6331 PAD.n7213 VSS 0.042751f
C6332 PAD.n7214 VSS 0.042751f
C6333 PAD.n7215 VSS 0.611619f
C6334 PAD.n7216 VSS 0.453782f
C6335 PAD.n7217 VSS 0.069752f
C6336 PAD.n7218 VSS 0.069752f
C6337 PAD.n7219 VSS 0.069752f
C6338 PAD.n7220 VSS 0.062262f
C6339 PAD.n7221 VSS 0.675741f
C6340 PAD.n7222 VSS 0.611619f
C6341 PAD.n7223 VSS 0.596822f
C6342 PAD.n7224 VSS 0.069752f
C6343 PAD.n7225 VSS 0.069752f
C6344 PAD.n7226 VSS 0.062262f
C6345 PAD.n7227 VSS 0.077409f
C6346 PAD.n7228 VSS 0.036454f
C6347 PAD.n7229 VSS 0.036454f
C6348 PAD.n7230 VSS 0.036454f
C6349 PAD.n7231 VSS 0.036454f
C6350 PAD.n7232 VSS 0.036454f
C6351 PAD.n7233 VSS 0.036454f
C6352 PAD.n7234 VSS 0.036454f
C6353 PAD.n7235 VSS 0.036454f
C6354 PAD.n7236 VSS 0.036454f
C6355 PAD.n7237 VSS 0.036454f
C6356 PAD.n7238 VSS 0.036454f
C6357 PAD.n7239 VSS 0.036454f
C6358 PAD.n7240 VSS 0.036454f
C6359 PAD.n7241 VSS 0.036454f
C6360 PAD.n7242 VSS 0.036454f
C6361 PAD.n7243 VSS 0.036454f
C6362 PAD.n7244 VSS 0.036454f
C6363 PAD.n7245 VSS 0.036454f
C6364 PAD.n7246 VSS 0.036454f
C6365 PAD.n7247 VSS 0.036454f
C6366 PAD.n7248 VSS 0.036454f
C6367 PAD.n7249 VSS 0.036454f
C6368 PAD.n7250 VSS 0.036454f
C6369 PAD.n7251 VSS 0.036454f
C6370 PAD.n7252 VSS 0.036454f
C6371 PAD.n7253 VSS 0.036454f
C6372 PAD.n7254 VSS 0.036454f
C6373 PAD.n7255 VSS 0.036454f
C6374 PAD.n7256 VSS 0.036454f
C6375 PAD.n7257 VSS 0.036454f
C6376 PAD.n7258 VSS 0.036454f
C6377 PAD.n7259 VSS 0.036454f
C6378 PAD.n7260 VSS 0.036454f
C6379 PAD.n7261 VSS 0.036454f
C6380 PAD.n7262 VSS 0.036454f
C6381 PAD.n7263 VSS 0.036454f
C6382 PAD.n7264 VSS 0.036454f
C6383 PAD.n7265 VSS 0.036454f
C6384 PAD.n7266 VSS 0.036454f
C6385 PAD.n7267 VSS 0.036454f
C6386 PAD.n7268 VSS 0.03055f
C6387 PAD.n7269 VSS 0.023105f
C6388 PAD.n7270 VSS 0.023105f
C6389 PAD.n7271 VSS 0.036454f
C6390 PAD.n7273 VSS 0.036454f
C6391 PAD.n7274 VSS 0.036454f
C6392 PAD.n7275 VSS 0.036454f
C6393 PAD.n7276 VSS 0.036454f
C6394 PAD.n7277 VSS 0.036454f
C6395 PAD.n7278 VSS 0.036454f
C6396 PAD.n7279 VSS 0.036454f
C6397 PAD.n7281 VSS 0.036454f
C6398 PAD.n7282 VSS 0.036454f
C6399 PAD.n7283 VSS 0.036454f
C6400 PAD.n7285 VSS 0.036454f
C6401 PAD.n7286 VSS 0.036454f
C6402 PAD.n7287 VSS 0.036454f
C6403 PAD.n7288 VSS 0.036454f
C6404 PAD.n7289 VSS 0.036454f
C6405 PAD.n7290 VSS 0.036454f
C6406 PAD.n7291 VSS 0.036454f
C6407 PAD.n7293 VSS 0.036454f
C6408 PAD.n7294 VSS 0.036454f
C6409 PAD.n7295 VSS 0.036454f
C6410 PAD.n7297 VSS 0.036454f
C6411 PAD.n7298 VSS 0.036454f
C6412 PAD.n7299 VSS 0.036454f
C6413 PAD.n7300 VSS 0.036454f
C6414 PAD.n7301 VSS 0.036454f
C6415 PAD.n7302 VSS 0.036454f
C6416 PAD.n7303 VSS 0.036454f
C6417 PAD.n7305 VSS 0.036454f
C6418 PAD.n7306 VSS 0.036454f
C6419 PAD.n7307 VSS 0.036454f
C6420 PAD.n7309 VSS 0.036454f
C6421 PAD.n7310 VSS 0.036454f
C6422 PAD.n7311 VSS 0.036454f
C6423 PAD.n7312 VSS 0.036454f
C6424 PAD.n7313 VSS 0.036454f
C6425 PAD.n7314 VSS 0.036454f
C6426 PAD.n7315 VSS 0.036454f
C6427 PAD.n7317 VSS 0.036454f
C6428 PAD.n7318 VSS 0.036454f
C6429 PAD.n7319 VSS 0.036454f
C6430 PAD.n7321 VSS 0.036454f
C6431 PAD.n7322 VSS 0.036454f
C6432 PAD.n7323 VSS 0.036454f
C6433 PAD.n7324 VSS 0.036454f
C6434 PAD.n7325 VSS 0.036454f
C6435 PAD.n7326 VSS 0.036454f
C6436 PAD.n7327 VSS 0.036454f
C6437 PAD.n7329 VSS 0.036454f
C6438 PAD.n7330 VSS 0.036454f
C6439 PAD.n7331 VSS 0.036454f
C6440 PAD.n7333 VSS 0.036454f
C6441 PAD.n7334 VSS 0.036454f
C6442 PAD.n7335 VSS 0.036454f
C6443 PAD.n7336 VSS 0.036454f
C6444 PAD.n7337 VSS 0.036454f
C6445 PAD.n7338 VSS 0.036454f
C6446 PAD.n7339 VSS 0.036454f
C6447 PAD.n7341 VSS 0.036454f
C6448 PAD.n7342 VSS 0.036454f
C6449 PAD.n7343 VSS 0.036454f
C6450 PAD.n7345 VSS 0.036454f
C6451 PAD.n7346 VSS 0.036454f
C6452 PAD.n7347 VSS 0.036454f
C6453 PAD.n7348 VSS 0.036454f
C6454 PAD.n7349 VSS 0.036454f
C6455 PAD.n7350 VSS 0.036454f
C6456 PAD.n7351 VSS 0.036454f
C6457 PAD.n7353 VSS 0.036454f
C6458 PAD.n7354 VSS 0.036454f
C6459 PAD.n7355 VSS 0.036454f
C6460 PAD.n7357 VSS 0.036454f
C6461 PAD.n7358 VSS 0.036454f
C6462 PAD.n7359 VSS 0.036454f
C6463 PAD.n7360 VSS 0.036454f
C6464 PAD.n7361 VSS 0.036454f
C6465 PAD.n7362 VSS 0.036454f
C6466 PAD.n7363 VSS 0.036454f
C6467 PAD.n7365 VSS 0.036454f
C6468 PAD.n7366 VSS 0.036454f
C6469 PAD.n7367 VSS 0.036454f
C6470 PAD.n7369 VSS 0.036454f
C6471 PAD.n7370 VSS 0.036454f
C6472 PAD.n7371 VSS 0.036454f
C6473 PAD.n7372 VSS 0.036454f
C6474 PAD.n7373 VSS 0.036454f
C6475 PAD.n7374 VSS 0.036454f
C6476 PAD.n7375 VSS 0.036454f
C6477 PAD.n7377 VSS 0.036454f
C6478 PAD.n7378 VSS 0.036454f
C6479 PAD.n7379 VSS 0.036454f
C6480 PAD.n7381 VSS 0.036454f
C6481 PAD.n7382 VSS 0.036454f
C6482 PAD.n7383 VSS 0.036454f
C6483 PAD.n7384 VSS 0.036454f
C6484 PAD.n7385 VSS 0.036454f
C6485 PAD.n7386 VSS 0.036454f
C6486 PAD.n7387 VSS 0.036454f
C6487 PAD.n7389 VSS 0.036454f
C6488 PAD.n7390 VSS 0.036454f
C6489 PAD.n7391 VSS 0.036454f
C6490 PAD.n7393 VSS 0.036454f
C6491 PAD.n7394 VSS 0.036454f
C6492 PAD.n7395 VSS 0.036454f
C6493 PAD.n7396 VSS 0.036454f
C6494 PAD.n7397 VSS 0.036454f
C6495 PAD.n7398 VSS 0.036454f
C6496 PAD.n7399 VSS 0.036454f
C6497 PAD.n7401 VSS 0.036454f
C6498 PAD.n7402 VSS 0.036454f
C6499 PAD.n7403 VSS 0.036454f
C6500 PAD.n7405 VSS 0.036454f
C6501 PAD.n7406 VSS 0.036454f
C6502 PAD.n7407 VSS 0.036454f
C6503 PAD.n7408 VSS 0.036454f
C6504 PAD.n7409 VSS 0.036454f
C6505 PAD.n7410 VSS 0.036454f
C6506 PAD.n7411 VSS 0.036454f
C6507 PAD.n7413 VSS 0.036454f
C6508 PAD.n7414 VSS 0.036454f
C6509 PAD.n7415 VSS 0.036454f
C6510 PAD.n7417 VSS 0.036454f
C6511 PAD.n7418 VSS 0.036454f
C6512 PAD.n7419 VSS 0.036454f
C6513 PAD.n7420 VSS 0.036454f
C6514 PAD.n7421 VSS 0.036454f
C6515 PAD.n7422 VSS 0.036454f
C6516 PAD.n7423 VSS 0.036454f
C6517 PAD.n7425 VSS 0.036454f
C6518 PAD.n7426 VSS 0.036454f
C6519 PAD.n7427 VSS 0.036454f
C6520 PAD.n7429 VSS 0.036454f
C6521 PAD.n7430 VSS 0.036454f
C6522 PAD.n7431 VSS 0.036454f
C6523 PAD.n7432 VSS 0.036454f
C6524 PAD.n7433 VSS 0.036454f
C6525 PAD.n7434 VSS 0.036454f
C6526 PAD.n7435 VSS 0.036454f
C6527 PAD.n7437 VSS 0.036454f
C6528 PAD.n7438 VSS 0.036454f
C6529 PAD.n7439 VSS 0.036454f
C6530 PAD.n7441 VSS 0.036454f
C6531 PAD.n7442 VSS 0.036454f
C6532 PAD.n7443 VSS 0.036454f
C6533 PAD.n7444 VSS 0.036454f
C6534 PAD.n7445 VSS 0.036454f
C6535 PAD.n7446 VSS 0.036454f
C6536 PAD.n7447 VSS 0.036454f
C6537 PAD.n7449 VSS 0.036454f
C6538 PAD.n7450 VSS 0.036454f
C6539 PAD.n7451 VSS 0.036454f
C6540 PAD.n7453 VSS 0.036454f
C6541 PAD.n7454 VSS 0.036454f
C6542 PAD.n7455 VSS 0.036454f
C6543 PAD.n7456 VSS 0.036454f
C6544 PAD.n7457 VSS 0.036454f
C6545 PAD.n7458 VSS 0.036454f
C6546 PAD.n7459 VSS 0.036454f
C6547 PAD.n7461 VSS 0.036454f
C6548 PAD.n7462 VSS 0.036454f
C6549 PAD.n7463 VSS 0.036454f
C6550 PAD.n7465 VSS 0.036454f
C6551 PAD.n7466 VSS 0.036454f
C6552 PAD.n7467 VSS 0.036454f
C6553 PAD.n7468 VSS 0.036454f
C6554 PAD.n7469 VSS 0.036454f
C6555 PAD.n7470 VSS 0.036454f
C6556 PAD.n7471 VSS 0.036454f
C6557 PAD.n7473 VSS 0.036454f
C6558 PAD.n7474 VSS 0.036454f
C6559 PAD.n7475 VSS 0.036454f
C6560 PAD.n7477 VSS 0.036454f
C6561 PAD.n7478 VSS 0.036454f
C6562 PAD.n7479 VSS 0.036454f
C6563 PAD.n7480 VSS 0.036454f
C6564 PAD.n7481 VSS 0.036454f
C6565 PAD.n7482 VSS 0.036454f
C6566 PAD.n7483 VSS 0.036454f
C6567 PAD.n7485 VSS 0.036454f
C6568 PAD.n7486 VSS 0.036454f
C6569 PAD.n7487 VSS 0.036454f
C6570 PAD.n7489 VSS 0.036454f
C6571 PAD.n7490 VSS 0.036454f
C6572 PAD.n7491 VSS 0.036454f
C6573 PAD.n7492 VSS 0.036454f
C6574 PAD.n7493 VSS 0.036454f
C6575 PAD.n7494 VSS 0.036454f
C6576 PAD.n7495 VSS 0.036454f
C6577 PAD.n7497 VSS 0.036454f
C6578 PAD.n7498 VSS 0.036454f
C6579 PAD.n7499 VSS 0.036454f
C6580 PAD.n7501 VSS 0.036454f
C6581 PAD.n7502 VSS 0.036454f
C6582 PAD.n7503 VSS 0.036454f
C6583 PAD.n7504 VSS 0.036454f
C6584 PAD.n7505 VSS 0.036454f
C6585 PAD.n7506 VSS 0.036454f
C6586 PAD.n7507 VSS 0.036454f
C6587 PAD.n7509 VSS 0.036454f
C6588 PAD.n7510 VSS 0.036454f
C6589 PAD.n7512 VSS 0.036454f
C6590 PAD.n7513 VSS 0.036454f
C6591 PAD.n7514 VSS 0.036454f
C6592 PAD.n7515 VSS 0.036454f
C6593 PAD.n7516 VSS 0.033374f
C6594 PAD.n7517 VSS 0.023105f
C6595 PAD.n7518 VSS 0.023105f
C6596 PAD.n7520 VSS 0.42912f
C6597 PAD.n7521 VSS 0.286079f
C6598 PAD.n7522 VSS 0.039596f
C6599 PAD.n7523 VSS 0.039596f
C6600 PAD.n7524 VSS 0.034582f
C6601 PAD.n7525 VSS 0.042887f
C6602 PAD.n7526 VSS 0.025823f
C6603 PAD.n7527 VSS 0.029567f
C6604 PAD.n7528 VSS 0.251553f
C6605 PAD.n7529 VSS 0.029567f
C6606 PAD.n7530 VSS 0.029431f
C6607 PAD.n7531 VSS 0.023105f
C6608 PAD.n7532 VSS 0.023105f
C6609 PAD.n7533 VSS 0.036454f
C6610 PAD.n7535 VSS 0.036454f
C6611 PAD.n7536 VSS 0.036454f
C6612 PAD.n7537 VSS 0.036454f
C6613 PAD.n7538 VSS 0.036454f
C6614 PAD.n7539 VSS 0.036454f
C6615 PAD.n7540 VSS 0.036454f
C6616 PAD.n7541 VSS 0.036454f
C6617 PAD.n7543 VSS 0.036454f
C6618 PAD.n7544 VSS 0.036454f
C6619 PAD.n7545 VSS 0.036454f
C6620 PAD.n7547 VSS 0.036454f
C6621 PAD.n7548 VSS 0.036454f
C6622 PAD.n7549 VSS 0.036454f
C6623 PAD.n7550 VSS 0.036454f
C6624 PAD.n7551 VSS 0.036454f
C6625 PAD.n7552 VSS 0.036454f
C6626 PAD.n7553 VSS 0.036454f
C6627 PAD.n7555 VSS 0.036454f
C6628 PAD.n7556 VSS 0.036454f
C6629 PAD.n7557 VSS 0.036454f
C6630 PAD.n7559 VSS 0.036454f
C6631 PAD.n7560 VSS 0.036454f
C6632 PAD.n7561 VSS 0.036454f
C6633 PAD.n7562 VSS 0.036454f
C6634 PAD.n7563 VSS 0.036454f
C6635 PAD.n7564 VSS 0.036454f
C6636 PAD.n7565 VSS 0.036454f
C6637 PAD.n7567 VSS 0.036454f
C6638 PAD.n7568 VSS 0.036454f
C6639 PAD.n7569 VSS 0.036454f
C6640 PAD.n7571 VSS 0.036454f
C6641 PAD.n7572 VSS 0.036454f
C6642 PAD.n7573 VSS 0.036454f
C6643 PAD.n7574 VSS 0.036454f
C6644 PAD.n7575 VSS 0.036454f
C6645 PAD.n7576 VSS 0.036454f
C6646 PAD.n7577 VSS 0.036454f
C6647 PAD.n7579 VSS 0.036454f
C6648 PAD.n7580 VSS 0.036454f
C6649 PAD.n7581 VSS 0.036454f
C6650 PAD.n7583 VSS 0.036454f
C6651 PAD.n7584 VSS 0.036454f
C6652 PAD.n7585 VSS 0.036454f
C6653 PAD.n7586 VSS 0.036454f
C6654 PAD.n7587 VSS 0.036454f
C6655 PAD.n7588 VSS 0.036454f
C6656 PAD.n7589 VSS 0.036454f
C6657 PAD.n7591 VSS 0.036454f
C6658 PAD.n7592 VSS 0.036454f
C6659 PAD.n7593 VSS 0.036454f
C6660 PAD.n7595 VSS 0.036454f
C6661 PAD.n7596 VSS 0.036454f
C6662 PAD.n7597 VSS 0.036454f
C6663 PAD.n7598 VSS 0.036454f
C6664 PAD.n7599 VSS 0.036454f
C6665 PAD.n7600 VSS 0.036454f
C6666 PAD.n7601 VSS 0.036454f
C6667 PAD.n7603 VSS 0.036454f
C6668 PAD.n7604 VSS 0.036454f
C6669 PAD.n7605 VSS 0.036454f
C6670 PAD.n7607 VSS 0.036454f
C6671 PAD.n7608 VSS 0.036454f
C6672 PAD.n7609 VSS 0.036454f
C6673 PAD.n7610 VSS 0.036454f
C6674 PAD.n7611 VSS 0.036454f
C6675 PAD.n7612 VSS 0.036454f
C6676 PAD.n7613 VSS 0.036454f
C6677 PAD.n7615 VSS 0.036454f
C6678 PAD.n7616 VSS 0.036454f
C6679 PAD.n7617 VSS 0.036454f
C6680 PAD.n7619 VSS 0.036454f
C6681 PAD.n7620 VSS 0.036454f
C6682 PAD.n7621 VSS 0.036454f
C6683 PAD.n7622 VSS 0.036454f
C6684 PAD.n7623 VSS 0.036454f
C6685 PAD.n7624 VSS 0.036454f
C6686 PAD.n7625 VSS 0.036454f
C6687 PAD.n7627 VSS 0.036454f
C6688 PAD.n7628 VSS 0.036454f
C6689 PAD.n7629 VSS 0.036454f
C6690 PAD.n7631 VSS 0.036454f
C6691 PAD.n7632 VSS 0.036454f
C6692 PAD.n7633 VSS 0.036454f
C6693 PAD.n7634 VSS 0.036454f
C6694 PAD.n7635 VSS 0.036454f
C6695 PAD.n7636 VSS 0.036454f
C6696 PAD.n7637 VSS 0.036454f
C6697 PAD.n7639 VSS 0.036454f
C6698 PAD.n7640 VSS 0.036454f
C6699 PAD.n7641 VSS 0.036454f
C6700 PAD.n7643 VSS 0.036454f
C6701 PAD.n7644 VSS 0.036454f
C6702 PAD.n7645 VSS 0.036454f
C6703 PAD.n7646 VSS 0.036454f
C6704 PAD.n7647 VSS 0.036454f
C6705 PAD.n7648 VSS 0.036454f
C6706 PAD.n7649 VSS 0.036454f
C6707 PAD.n7651 VSS 0.036454f
C6708 PAD.n7652 VSS 0.036454f
C6709 PAD.n7653 VSS 0.036454f
C6710 PAD.n7655 VSS 0.036454f
C6711 PAD.n7656 VSS 0.036454f
C6712 PAD.n7657 VSS 0.036454f
C6713 PAD.n7658 VSS 0.036454f
C6714 PAD.n7659 VSS 0.036454f
C6715 PAD.n7660 VSS 0.036454f
C6716 PAD.n7661 VSS 0.036454f
C6717 PAD.n7663 VSS 0.036454f
C6718 PAD.n7664 VSS 0.036454f
C6719 PAD.n7665 VSS 0.036454f
C6720 PAD.n7667 VSS 0.036454f
C6721 PAD.n7668 VSS 0.036454f
C6722 PAD.n7669 VSS 0.036454f
C6723 PAD.n7670 VSS 0.036454f
C6724 PAD.n7671 VSS 0.036454f
C6725 PAD.n7672 VSS 0.036454f
C6726 PAD.n7673 VSS 0.036454f
C6727 PAD.n7675 VSS 0.036454f
C6728 PAD.n7676 VSS 0.036454f
C6729 PAD.n7677 VSS 0.036454f
C6730 PAD.n7679 VSS 0.036454f
C6731 PAD.n7680 VSS 0.036454f
C6732 PAD.n7681 VSS 0.036454f
C6733 PAD.n7682 VSS 0.036454f
C6734 PAD.n7683 VSS 0.036454f
C6735 PAD.n7684 VSS 0.036454f
C6736 PAD.n7685 VSS 0.036454f
C6737 PAD.n7687 VSS 0.036454f
C6738 PAD.n7688 VSS 0.036454f
C6739 PAD.n7689 VSS 0.036454f
C6740 PAD.n7691 VSS 0.036454f
C6741 PAD.n7692 VSS 0.036454f
C6742 PAD.n7693 VSS 0.036454f
C6743 PAD.n7694 VSS 0.036454f
C6744 PAD.n7695 VSS 0.036454f
C6745 PAD.n7696 VSS 0.036454f
C6746 PAD.n7697 VSS 0.036454f
C6747 PAD.n7699 VSS 0.036454f
C6748 PAD.n7700 VSS 0.036454f
C6749 PAD.n7701 VSS 0.036454f
C6750 PAD.n7703 VSS 0.036454f
C6751 PAD.n7704 VSS 0.036454f
C6752 PAD.n7705 VSS 0.036454f
C6753 PAD.n7706 VSS 0.036454f
C6754 PAD.n7707 VSS 0.036454f
C6755 PAD.n7708 VSS 0.036454f
C6756 PAD.n7709 VSS 0.036454f
C6757 PAD.n7711 VSS 0.036454f
C6758 PAD.n7712 VSS 0.036454f
C6759 PAD.n7713 VSS 0.036454f
C6760 PAD.n7715 VSS 0.036454f
C6761 PAD.n7716 VSS 0.036454f
C6762 PAD.n7717 VSS 0.036454f
C6763 PAD.n7718 VSS 0.036454f
C6764 PAD.n7719 VSS 0.036454f
C6765 PAD.n7720 VSS 0.036454f
C6766 PAD.n7721 VSS 0.036454f
C6767 PAD.n7723 VSS 0.036454f
C6768 PAD.n7724 VSS 0.036454f
C6769 PAD.n7725 VSS 0.036454f
C6770 PAD.n7727 VSS 0.036454f
C6771 PAD.n7728 VSS 0.036454f
C6772 PAD.n7729 VSS 0.036454f
C6773 PAD.n7730 VSS 0.036454f
C6774 PAD.n7731 VSS 0.036454f
C6775 PAD.n7732 VSS 0.036454f
C6776 PAD.n7733 VSS 0.036454f
C6777 PAD.n7735 VSS 0.036454f
C6778 PAD.n7736 VSS 0.036454f
C6779 PAD.n7737 VSS 0.036454f
C6780 PAD.n7739 VSS 0.036454f
C6781 PAD.n7740 VSS 0.036454f
C6782 PAD.n7741 VSS 0.036454f
C6783 PAD.n7742 VSS 0.036454f
C6784 PAD.n7743 VSS 0.036454f
C6785 PAD.n7744 VSS 0.036454f
C6786 PAD.n7745 VSS 0.036454f
C6787 PAD.n7747 VSS 0.036454f
C6788 PAD.n7748 VSS 0.036454f
C6789 PAD.n7749 VSS 0.036454f
C6790 PAD.n7751 VSS 0.036454f
C6791 PAD.n7752 VSS 0.036454f
C6792 PAD.n7753 VSS 0.036454f
C6793 PAD.n7754 VSS 0.036454f
C6794 PAD.n7755 VSS 0.036454f
C6795 PAD.n7756 VSS 0.036454f
C6796 PAD.n7757 VSS 0.036454f
C6797 PAD.n7759 VSS 0.036454f
C6798 PAD.n7760 VSS 0.036454f
C6799 PAD.n7761 VSS 0.036454f
C6800 PAD.n7763 VSS 0.036454f
C6801 PAD.n7764 VSS 0.036454f
C6802 PAD.n7765 VSS 0.036454f
C6803 PAD.n7766 VSS 0.036454f
C6804 PAD.n7767 VSS 0.036454f
C6805 PAD.n7768 VSS 0.036454f
C6806 PAD.n7769 VSS 0.036454f
C6807 PAD.n7771 VSS 0.036454f
C6808 PAD.n7772 VSS 0.036454f
C6809 PAD.n7774 VSS 0.036454f
C6810 PAD.n7775 VSS 0.036454f
C6811 PAD.n7776 VSS 0.036454f
C6812 PAD.n7777 VSS 0.036454f
C6813 PAD.n7778 VSS 0.033374f
C6814 PAD.n7779 VSS 0.023105f
C6815 PAD.n7780 VSS 0.023105f
C6816 PAD.n7782 VSS 0.611619f
C6817 PAD.n7783 VSS 0.24662f
C6818 PAD.n7784 VSS 0.061877f
C6819 PAD.n7785 VSS 0.061877f
C6820 PAD.n7786 VSS 0.055232f
C6821 PAD.n7787 VSS 0.062262f
C6822 PAD.n7788 VSS 0.04519f
C6823 PAD.n7789 VSS 0.050627f
C6824 PAD.n7790 VSS 0.050627f
C6825 PAD.n7791 VSS 0.350201f
C6826 PAD.n7792 VSS 0.611619f
C6827 PAD.n7793 VSS 0.025072f
C6828 PAD.n7794 VSS 0.025072f
C6829 PAD.n7795 VSS 0.021897f
C6830 PAD.n7796 VSS 0.033766f
C6831 PAD.n7797 VSS 0.042434f
C6832 PAD.n7798 VSS 0.039414f
C6833 PAD.n7799 VSS 0.045129f
C6834 PAD.n7800 VSS 0.045129f
C6835 PAD.n7801 VSS 0.611619f
C6836 PAD.n7802 VSS 0.221958f
C6837 PAD.n7803 VSS 0.058502f
C6838 PAD.n7804 VSS 0.058502f
C6839 PAD.n7805 VSS 0.05222f
C6840 PAD.n7806 VSS 0.041759f
C6841 PAD.n7807 VSS 1.26066f
C6842 PAD.n7808 VSS 16.0799f
C6843 PAD.n7809 VSS 19.3704f
C6844 PAD.n7810 VSS 13.142799f
C6845 PAD.n7811 VSS 14.504801f
C6846 PAD.n7812 VSS 8.7754f
C6847 PAD.n7813 VSS 0.061877f
C6848 PAD.n7814 VSS 0.034646f
C6849 PAD.n7815 VSS 0.046278f
C6850 PAD.n7816 VSS 0.038161f
C6851 PAD.n7817 VSS 0.042751f
C6852 PAD.n7818 VSS 0.042751f
C6853 PAD.n7819 VSS 0.675741f
C6854 PAD.n7820 VSS 0.187431f
C6855 PAD.n7821 VSS 0.0351f
C6856 PAD.n7822 VSS 0.0351f
C6857 PAD.n7823 VSS 0.030655f
C6858 PAD.n7824 VSS 0.033766f
C6859 PAD.n7825 VSS 0.033676f
C6860 PAD.n7826 VSS 0.038559f
C6861 PAD.n7827 VSS 0.038559f
C6862 PAD.n7828 VSS 0.098648f
C6863 PAD.n7829 VSS 0.685606f
C6864 PAD.n7871 VSS 0.036454f
C6865 PAD.n7873 VSS 0.036454f
C6866 PAD.n7874 VSS 0.036454f
C6867 PAD.n7875 VSS 0.036454f
C6868 PAD.n7876 VSS 0.036454f
C6869 PAD.n7877 VSS 0.036454f
C6870 PAD.n7879 VSS 0.036454f
C6871 PAD.n7880 VSS 0.036454f
C6872 PAD.n7881 VSS 0.036454f
C6873 PAD.n7882 VSS 0.036454f
C6874 PAD.n7884 VSS 0.036454f
C6875 PAD.n7885 VSS 0.036454f
C6876 PAD.n7886 VSS 0.036454f
C6877 PAD.n7887 VSS 0.036454f
C6878 PAD.n7889 VSS 0.036454f
C6879 PAD.n7890 VSS 0.036454f
C6880 PAD.n7891 VSS 0.036454f
C6881 PAD.n7892 VSS 0.036454f
C6882 PAD.n7894 VSS 0.036454f
C6883 PAD.n7895 VSS 0.036454f
C6884 PAD.n7896 VSS 0.036454f
C6885 PAD.n7897 VSS 0.036454f
C6886 PAD.n7899 VSS 0.036454f
C6887 PAD.n7900 VSS 0.036454f
C6888 PAD.n7901 VSS 0.036454f
C6889 PAD.n7902 VSS 0.036454f
C6890 PAD.n7904 VSS 0.036454f
C6891 PAD.n7905 VSS 0.036454f
C6892 PAD.n7906 VSS 0.036454f
C6893 PAD.n7907 VSS 0.036454f
C6894 PAD.n7909 VSS 0.036454f
C6895 PAD.n7910 VSS 0.036454f
C6896 PAD.n7911 VSS 0.036454f
C6897 PAD.n7912 VSS 0.036454f
C6898 PAD.n7914 VSS 0.036454f
C6899 PAD.n7915 VSS 0.036454f
C6900 PAD.n7916 VSS 0.036454f
C6901 PAD.n7917 VSS 0.036454f
C6902 PAD.n7919 VSS 0.036454f
C6903 PAD.n7920 VSS 0.036454f
C6904 PAD.n7921 VSS 0.036454f
C6905 PAD.n7922 VSS 0.036454f
C6906 PAD.n7924 VSS 0.036454f
C6907 PAD.n7925 VSS 0.036454f
C6908 PAD.n7926 VSS 0.036454f
C6909 PAD.n7927 VSS 0.036454f
C6910 PAD.n7929 VSS 0.036454f
C6911 PAD.n7930 VSS 0.036454f
C6912 PAD.n7931 VSS 0.036454f
C6913 PAD.n7932 VSS 0.036454f
C6914 PAD.n7934 VSS 0.036454f
C6915 PAD.n7935 VSS 0.036454f
C6916 PAD.n7936 VSS 0.036454f
C6917 PAD.n7937 VSS 0.036454f
C6918 PAD.n7939 VSS 0.036454f
C6919 PAD.n7940 VSS 0.036454f
C6920 PAD.n7941 VSS 0.036454f
C6921 PAD.n7942 VSS 0.036454f
C6922 PAD.n7944 VSS 0.036454f
C6923 PAD.n7945 VSS 0.036454f
C6924 PAD.n7946 VSS 0.036454f
C6925 PAD.n7947 VSS 0.036454f
C6926 PAD.n7949 VSS 0.036454f
C6927 PAD.n7950 VSS 0.036454f
C6928 PAD.n7951 VSS 0.036454f
C6929 PAD.n7952 VSS 0.036454f
C6930 PAD.n7954 VSS 0.036454f
C6931 PAD.n7955 VSS 0.036454f
C6932 PAD.n7956 VSS 0.036454f
C6933 PAD.n7957 VSS 0.036454f
C6934 PAD.n7959 VSS 0.036454f
C6935 PAD.n7960 VSS 0.036454f
C6936 PAD.n7961 VSS 0.036454f
C6937 PAD.n7962 VSS 0.036454f
C6938 PAD.n7964 VSS 0.036454f
C6939 PAD.n7965 VSS 0.036454f
C6940 PAD.n7966 VSS 0.036454f
C6941 PAD.n7967 VSS 0.036454f
C6942 PAD.n7969 VSS 0.036454f
C6943 PAD.n7970 VSS 0.036454f
C6944 PAD.n7971 VSS 0.023105f
C6945 PAD.n7972 VSS 0.023105f
C6946 PAD.n7973 VSS 0.036454f
C6947 PAD.n7974 VSS 0.036454f
C6948 PAD.n7976 VSS 0.036454f
C6949 PAD.n7977 VSS 0.036454f
C6950 PAD.n7978 VSS 0.036454f
C6951 PAD.n7979 VSS 0.036454f
C6952 PAD.n7980 VSS 0.036454f
C6953 PAD.n7981 VSS 0.036454f
C6954 PAD.n7983 VSS 0.036454f
C6955 PAD.n7984 VSS 0.036454f
C6956 PAD.n7985 VSS 0.036454f
C6957 PAD.n7986 VSS 0.036454f
C6958 PAD.n7987 VSS 0.036454f
C6959 PAD.n7988 VSS 0.036454f
C6960 PAD.n7989 VSS 0.036454f
C6961 PAD.n7990 VSS 0.036454f
C6962 PAD.n7992 VSS 0.036454f
C6963 PAD.n7993 VSS 0.036454f
C6964 PAD.n7994 VSS 0.036454f
C6965 PAD.n7995 VSS 0.036454f
C6966 PAD.n7996 VSS 0.036454f
C6967 PAD.n7997 VSS 0.036454f
C6968 PAD.n7998 VSS 0.036454f
C6969 PAD.n7999 VSS 0.036454f
C6970 PAD.n8001 VSS 0.036454f
C6971 PAD.n8002 VSS 0.036454f
C6972 PAD.n8003 VSS 0.036454f
C6973 PAD.n8004 VSS 0.036454f
C6974 PAD.n8005 VSS 0.036454f
C6975 PAD.n8006 VSS 0.036454f
C6976 PAD.n8007 VSS 0.036454f
C6977 PAD.n8008 VSS 0.036454f
C6978 PAD.n8010 VSS 0.036454f
C6979 PAD.n8011 VSS 0.036454f
C6980 PAD.n8012 VSS 0.036454f
C6981 PAD.n8013 VSS 0.036454f
C6982 PAD.n8014 VSS 0.036454f
C6983 PAD.n8015 VSS 0.036454f
C6984 PAD.n8016 VSS 0.036454f
C6985 PAD.n8017 VSS 0.036454f
C6986 PAD.n8019 VSS 0.036454f
C6987 PAD.n8020 VSS 0.036454f
C6988 PAD.n8021 VSS 0.036454f
C6989 PAD.n8022 VSS 0.036454f
C6990 PAD.n8023 VSS 0.036454f
C6991 PAD.n8024 VSS 0.036454f
C6992 PAD.n8025 VSS 0.036454f
C6993 PAD.n8026 VSS 0.036454f
C6994 PAD.n8028 VSS 0.036454f
C6995 PAD.n8029 VSS 0.036454f
C6996 PAD.n8030 VSS 0.036454f
C6997 PAD.n8031 VSS 0.036454f
C6998 PAD.n8032 VSS 0.036454f
C6999 PAD.n8033 VSS 0.036454f
C7000 PAD.n8034 VSS 0.036454f
C7001 PAD.n8035 VSS 0.036454f
C7002 PAD.n8037 VSS 0.036454f
C7003 PAD.n8038 VSS 0.036454f
C7004 PAD.n8039 VSS 0.036454f
C7005 PAD.n8040 VSS 0.036454f
C7006 PAD.n8041 VSS 0.036454f
C7007 PAD.n8042 VSS 0.036454f
C7008 PAD.n8043 VSS 0.036454f
C7009 PAD.n8044 VSS 0.036454f
C7010 PAD.n8046 VSS 0.036454f
C7011 PAD.n8047 VSS 0.036454f
C7012 PAD.n8048 VSS 0.036454f
C7013 PAD.n8049 VSS 0.036454f
C7014 PAD.n8050 VSS 0.036454f
C7015 PAD.n8051 VSS 0.036454f
C7016 PAD.n8052 VSS 0.036454f
C7017 PAD.n8053 VSS 0.036454f
C7018 PAD.n8055 VSS 0.036454f
C7019 PAD.n8056 VSS 0.036454f
C7020 PAD.n8057 VSS 0.036454f
C7021 PAD.n8058 VSS 0.036454f
C7022 PAD.n8059 VSS 0.036454f
C7023 PAD.n8060 VSS 0.036454f
C7024 PAD.n8061 VSS 0.036454f
C7025 PAD.n8062 VSS 0.036454f
C7026 PAD.n8064 VSS 0.036454f
C7027 PAD.n8065 VSS 0.036454f
C7028 PAD.n8066 VSS 0.036454f
C7029 PAD.n8067 VSS 0.036454f
C7030 PAD.n8068 VSS 0.036454f
C7031 PAD.n8069 VSS 0.036454f
C7032 PAD.n8070 VSS 0.036454f
C7033 PAD.n8071 VSS 0.036454f
C7034 PAD.n8073 VSS 0.036454f
C7035 PAD.n8074 VSS 0.036454f
C7036 PAD.n8075 VSS 0.036454f
C7037 PAD.n8076 VSS 0.036454f
C7038 PAD.n8077 VSS 0.036454f
C7039 PAD.n8078 VSS 0.036454f
C7040 PAD.n8079 VSS 0.036454f
C7041 PAD.n8080 VSS 0.036454f
C7042 PAD.n8082 VSS 0.036454f
C7043 PAD.n8083 VSS 0.036454f
C7044 PAD.n8084 VSS 0.036454f
C7045 PAD.n8085 VSS 0.036454f
C7046 PAD.n8086 VSS 0.036454f
C7047 PAD.n8087 VSS 0.036454f
C7048 PAD.n8088 VSS 0.036454f
C7049 PAD.n8089 VSS 0.036454f
C7050 PAD.n8091 VSS 0.036454f
C7051 PAD.n8092 VSS 0.036454f
C7052 PAD.n8093 VSS 0.036454f
C7053 PAD.n8094 VSS 0.036454f
C7054 PAD.n8095 VSS 0.036454f
C7055 PAD.n8096 VSS 0.036454f
C7056 PAD.n8097 VSS 0.036454f
C7057 PAD.n8098 VSS 0.036454f
C7058 PAD.n8100 VSS 0.036454f
C7059 PAD.n8101 VSS 0.036454f
C7060 PAD.n8102 VSS 0.036454f
C7061 PAD.n8103 VSS 0.036454f
C7062 PAD.n8104 VSS 0.036454f
C7063 PAD.n8105 VSS 0.036454f
C7064 PAD.n8106 VSS 0.036454f
C7065 PAD.n8107 VSS 0.036454f
C7066 PAD.n8109 VSS 0.036454f
C7067 PAD.n8110 VSS 0.036454f
C7068 PAD.n8111 VSS 0.036454f
C7069 PAD.n8112 VSS 0.036454f
C7070 PAD.n8113 VSS 0.036454f
C7071 PAD.n8114 VSS 0.036454f
C7072 PAD.n8115 VSS 0.036454f
C7073 PAD.n8116 VSS 0.036454f
C7074 PAD.n8118 VSS 0.036454f
C7075 PAD.n8119 VSS 0.036454f
C7076 PAD.n8120 VSS 0.036454f
C7077 PAD.n8121 VSS 0.036454f
C7078 PAD.n8122 VSS 0.036454f
C7079 PAD.n8123 VSS 0.036454f
C7080 PAD.n8124 VSS 0.036454f
C7081 PAD.n8125 VSS 0.036454f
C7082 PAD.n8127 VSS 0.036454f
C7083 PAD.n8128 VSS 0.036454f
C7084 PAD.n8129 VSS 0.036454f
C7085 PAD.n8130 VSS 0.036454f
C7086 PAD.n8131 VSS 0.036454f
C7087 PAD.n8132 VSS 0.036454f
C7088 PAD.n8133 VSS 0.036454f
C7089 PAD.n8134 VSS 0.036454f
C7090 PAD.n8136 VSS 0.036454f
C7091 PAD.n8137 VSS 0.036454f
C7092 PAD.n8138 VSS 0.036454f
C7093 PAD.n8139 VSS 0.036454f
C7094 PAD.n8140 VSS 0.036454f
C7095 PAD.n8141 VSS 0.036454f
C7096 PAD.n8142 VSS 0.036454f
C7097 PAD.n8143 VSS 0.036454f
C7098 PAD.n8145 VSS 0.036454f
C7099 PAD.n8146 VSS 0.036454f
C7100 PAD.n8147 VSS 0.036454f
C7101 PAD.n8148 VSS 0.036454f
C7102 PAD.n8149 VSS 0.036454f
C7103 PAD.n8150 VSS 0.036454f
C7104 PAD.n8151 VSS 0.036454f
C7105 PAD.n8152 VSS 0.036454f
C7106 PAD.n8154 VSS 0.036454f
C7107 PAD.n8155 VSS 0.036454f
C7108 PAD.n8156 VSS 0.036454f
C7109 PAD.n8157 VSS 0.036454f
C7110 PAD.n8158 VSS 0.036454f
C7111 PAD.n8159 VSS 0.036454f
C7112 PAD.n8160 VSS 0.023105f
C7113 PAD.n8161 VSS 0.023105f
C7114 PAD.n8163 VSS 0.596822f
C7115 PAD.n8164 VSS 0.542565f
C7116 PAD.n8165 VSS 0.626417f
C7117 PAD.n8166 VSS 0.069752f
C7118 PAD.n8167 VSS 0.050627f
C7119 PAD.n8168 VSS 0.050627f
C7120 PAD.n8169 VSS 0.04519f
C7121 PAD.n8170 VSS 0.046278f
C7122 PAD.n8171 VSS 0.048203f
C7123 PAD.n8172 VSS 0.054002f
C7124 PAD.n8173 VSS 0.054002f
C7125 PAD.n8174 VSS 0.527768f
C7126 PAD.n8175 VSS 0.611619f
C7127 PAD.n8176 VSS 0.030605f
C7128 PAD.n8177 VSS 0.030605f
C7129 PAD.n8178 VSS 0.026729f
C7130 PAD.n8179 VSS 0.033766f
C7131 PAD.n8180 VSS 0.037602f
C7132 PAD.n8181 VSS 0.043054f
C7133 PAD.n8182 VSS 0.043054f
C7134 PAD.n8183 VSS 0.591889f
C7135 PAD.n8184 VSS 0.700403f
C7136 PAD.n8185 VSS 0.611619f
C7137 PAD.n8186 VSS 0.419255f
C7138 PAD.n8187 VSS 0.058502f
C7139 PAD.n8188 VSS 0.058502f
C7140 PAD.n8189 VSS 0.05222f
C7141 PAD.n8190 VSS 0.046278f
C7142 PAD.n8191 VSS 0.041173f
C7143 PAD.n8192 VSS 0.046126f
C7144 PAD.n8193 VSS 0.046126f
C7145 PAD.n8194 VSS 0.419255f
C7146 PAD.n8195 VSS 0.522836f
C7147 PAD.n8196 VSS 0.026109f
C7148 PAD.n8197 VSS 0.026109f
C7149 PAD.n8198 VSS 0.022803f
C7150 PAD.n8199 VSS 0.033766f
C7151 PAD.n8200 VSS 0.041528f
C7152 PAD.n8201 VSS 0.04755f
C7153 PAD.n8202 VSS 0.046166f
C7154 PAD.n8203 VSS 0.046166f
C7155 PAD.n8204 VSS 0.029431f
C7156 PAD.n8205 VSS 0.300877f
C7157 PAD.n8206 VSS 0.027492f
C7158 PAD.n8207 VSS 0.027492f
C7159 PAD.n8208 VSS 0.024011f
C7160 PAD.n8209 VSS 0.033766f
C7161 PAD.n8210 VSS 0.03055f
C7162 PAD.n8211 VSS 0.036454f
C7163 PAD.n8212 VSS 0.036454f
C7164 PAD.n8213 VSS 0.036454f
C7165 PAD.n8214 VSS 0.036454f
C7166 PAD.n8215 VSS 0.036454f
C7167 PAD.n8217 VSS 0.036454f
C7168 PAD.n8218 VSS 0.036454f
C7169 PAD.n8219 VSS 0.036454f
C7170 PAD.n8220 VSS 0.036454f
C7171 PAD.n8221 VSS 0.036454f
C7172 PAD.n8222 VSS 0.036454f
C7173 PAD.n8223 VSS 0.036454f
C7174 PAD.n8224 VSS 0.036454f
C7175 PAD.n8226 VSS 0.036454f
C7176 PAD.n8227 VSS 0.036454f
C7177 PAD.n8228 VSS 0.036454f
C7178 PAD.n8229 VSS 0.036454f
C7179 PAD.n8230 VSS 0.036454f
C7180 PAD.n8231 VSS 0.036454f
C7181 PAD.n8232 VSS 0.036454f
C7182 PAD.n8233 VSS 0.036454f
C7183 PAD.n8235 VSS 0.036454f
C7184 PAD.n8236 VSS 0.036454f
C7185 PAD.n8237 VSS 0.036454f
C7186 PAD.n8238 VSS 0.036454f
C7187 PAD.n8239 VSS 0.036454f
C7188 PAD.n8240 VSS 0.036454f
C7189 PAD.n8241 VSS 0.036454f
C7190 PAD.n8242 VSS 0.036454f
C7191 PAD.n8244 VSS 0.036454f
C7192 PAD.n8245 VSS 0.036454f
C7193 PAD.n8246 VSS 0.036454f
C7194 PAD.n8247 VSS 0.036454f
C7195 PAD.n8248 VSS 0.036454f
C7196 PAD.n8249 VSS 0.036454f
C7197 PAD.n8250 VSS 0.036454f
C7198 PAD.n8251 VSS 0.036454f
C7199 PAD.n8253 VSS 0.036454f
C7200 PAD.n8254 VSS 0.036454f
C7201 PAD.n8255 VSS 0.036454f
C7202 PAD.n8256 VSS 0.036454f
C7203 PAD.n8257 VSS 0.036454f
C7204 PAD.n8258 VSS 0.036454f
C7205 PAD.n8259 VSS 0.036454f
C7206 PAD.n8260 VSS 0.036454f
C7207 PAD.n8262 VSS 0.036454f
C7208 PAD.n8263 VSS 0.036454f
C7209 PAD.n8264 VSS 0.036454f
C7210 PAD.n8265 VSS 0.036454f
C7211 PAD.n8266 VSS 0.036454f
C7212 PAD.n8267 VSS 0.036454f
C7213 PAD.n8268 VSS 0.036454f
C7214 PAD.n8269 VSS 0.036454f
C7215 PAD.n8271 VSS 0.036454f
C7216 PAD.n8272 VSS 0.036454f
C7217 PAD.n8273 VSS 0.036454f
C7218 PAD.n8274 VSS 0.036454f
C7219 PAD.n8275 VSS 0.036454f
C7220 PAD.n8276 VSS 0.036454f
C7221 PAD.n8277 VSS 0.036454f
C7222 PAD.n8278 VSS 0.036454f
C7223 PAD.n8280 VSS 0.036454f
C7224 PAD.n8281 VSS 0.036454f
C7225 PAD.n8282 VSS 0.036454f
C7226 PAD.n8283 VSS 0.036454f
C7227 PAD.n8284 VSS 0.036454f
C7228 PAD.n8285 VSS 0.036454f
C7229 PAD.n8286 VSS 0.036454f
C7230 PAD.n8287 VSS 0.036454f
C7231 PAD.n8289 VSS 0.036454f
C7232 PAD.n8290 VSS 0.036454f
C7233 PAD.n8291 VSS 0.036454f
C7234 PAD.n8292 VSS 0.036454f
C7235 PAD.n8293 VSS 0.036454f
C7236 PAD.n8294 VSS 0.036454f
C7237 PAD.n8295 VSS 0.036454f
C7238 PAD.n8296 VSS 0.036454f
C7239 PAD.n8298 VSS 0.036454f
C7240 PAD.n8299 VSS 0.036454f
C7241 PAD.n8300 VSS 0.036454f
C7242 PAD.n8301 VSS 0.036454f
C7243 PAD.n8302 VSS 0.036454f
C7244 PAD.n8303 VSS 0.036454f
C7245 PAD.n8304 VSS 0.036454f
C7246 PAD.n8305 VSS 0.036454f
C7247 PAD.n8307 VSS 0.036454f
C7248 PAD.n8308 VSS 0.036454f
C7249 PAD.n8309 VSS 0.036454f
C7250 PAD.n8310 VSS 0.036454f
C7251 PAD.n8311 VSS 0.036454f
C7252 PAD.n8312 VSS 0.036454f
C7253 PAD.n8313 VSS 0.036454f
C7254 PAD.n8314 VSS 0.036454f
C7255 PAD.n8316 VSS 0.036454f
C7256 PAD.n8317 VSS 0.036454f
C7257 PAD.n8318 VSS 0.036454f
C7258 PAD.n8319 VSS 0.036454f
C7259 PAD.n8320 VSS 0.036454f
C7260 PAD.n8321 VSS 0.036454f
C7261 PAD.n8322 VSS 0.036454f
C7262 PAD.n8323 VSS 0.036454f
C7263 PAD.n8325 VSS 0.036454f
C7264 PAD.n8326 VSS 0.036454f
C7265 PAD.n8327 VSS 0.036454f
C7266 PAD.n8328 VSS 0.036454f
C7267 PAD.n8329 VSS 0.036454f
C7268 PAD.n8330 VSS 0.036454f
C7269 PAD.n8331 VSS 0.036454f
C7270 PAD.n8332 VSS 0.036454f
C7271 PAD.n8334 VSS 0.036454f
C7272 PAD.n8335 VSS 0.036454f
C7273 PAD.n8336 VSS 0.036454f
C7274 PAD.n8337 VSS 0.036454f
C7275 PAD.n8338 VSS 0.036454f
C7276 PAD.n8339 VSS 0.036454f
C7277 PAD.n8340 VSS 0.036454f
C7278 PAD.n8341 VSS 0.036454f
C7279 PAD.n8343 VSS 0.036454f
C7280 PAD.n8344 VSS 0.036454f
C7281 PAD.n8345 VSS 0.036454f
C7282 PAD.n8346 VSS 0.036454f
C7283 PAD.n8347 VSS 0.036454f
C7284 PAD.n8348 VSS 0.036454f
C7285 PAD.n8349 VSS 0.036454f
C7286 PAD.n8350 VSS 0.036454f
C7287 PAD.n8352 VSS 0.036454f
C7288 PAD.n8353 VSS 0.036454f
C7289 PAD.n8354 VSS 0.036454f
C7290 PAD.n8355 VSS 0.036454f
C7291 PAD.n8356 VSS 0.036454f
C7292 PAD.n8357 VSS 0.036454f
C7293 PAD.n8358 VSS 0.036454f
C7294 PAD.n8359 VSS 0.036454f
C7295 PAD.n8361 VSS 0.036454f
C7296 PAD.n8362 VSS 0.036454f
C7297 PAD.n8363 VSS 0.036454f
C7298 PAD.n8364 VSS 0.036454f
C7299 PAD.n8365 VSS 0.036454f
C7300 PAD.n8366 VSS 0.036454f
C7301 PAD.n8367 VSS 0.036454f
C7302 PAD.n8368 VSS 0.036454f
C7303 PAD.n8370 VSS 0.036454f
C7304 PAD.n8371 VSS 0.036454f
C7305 PAD.n8372 VSS 0.036454f
C7306 PAD.n8373 VSS 0.036454f
C7307 PAD.n8374 VSS 0.036454f
C7308 PAD.n8375 VSS 0.036454f
C7309 PAD.n8376 VSS 0.036454f
C7310 PAD.n8377 VSS 0.036454f
C7311 PAD.n8379 VSS 0.036454f
C7312 PAD.n8380 VSS 0.036454f
C7313 PAD.n8381 VSS 0.036454f
C7314 PAD.n8382 VSS 0.036454f
C7315 PAD.n8383 VSS 0.036454f
C7316 PAD.n8384 VSS 0.036454f
C7317 PAD.n8385 VSS 0.036454f
C7318 PAD.n8386 VSS 0.036454f
C7319 PAD.n8388 VSS 0.036454f
C7320 PAD.n8389 VSS 0.036454f
C7321 PAD.n8390 VSS 0.036454f
C7322 PAD.n8391 VSS 0.036454f
C7323 PAD.n8392 VSS 0.036454f
C7324 PAD.n8393 VSS 0.036454f
C7325 PAD.n8394 VSS 0.023105f
C7326 PAD.n8395 VSS 0.023105f
C7327 PAD.n8397 VSS 0.611619f
C7328 PAD.n8398 VSS 0.276215f
C7329 PAD.n8399 VSS 0.066377f
C7330 PAD.n8400 VSS 0.066377f
C7331 PAD.n8401 VSS 0.059249f
C7332 PAD.n8402 VSS 0.046278f
C7333 PAD.n8403 VSS 0.034144f
C7334 PAD.n8404 VSS 0.062262f
C7335 PAD.n8405 VSS 0.069752f
C7336 PAD.n8406 VSS 0.069752f
C7337 PAD.n8407 VSS 0.424187f
C7338 PAD.n8408 VSS 0.611619f
C7339 PAD.n8409 VSS 0.700403f
C7340 PAD.n8410 VSS 0.335404f
C7341 PAD.n8411 VSS 0.041671f
C7342 PAD.n8412 VSS 0.041671f
C7343 PAD.n8413 VSS 0.036394f
C7344 PAD.n8414 VSS 0.033766f
C7345 PAD.n8415 VSS 0.042887f
C7346 PAD.n8416 VSS 0.027937f
C7347 PAD.n8417 VSS 0.031988f
C7348 PAD.n8418 VSS 0.031988f
C7349 PAD.n8419 VSS 0.424187f
C7350 PAD.n8420 VSS 0.567228f
C7351 PAD.n8421 VSS 0.039376f
C7352 PAD.n8422 VSS 0.039376f
C7353 PAD.n8423 VSS 0.035148f
C7354 PAD.n8424 VSS 0.046278f
C7355 PAD.n8425 VSS 0.058245f
C7356 PAD.n8426 VSS 0.042178f
C7357 PAD.n8427 VSS 0.062262f
C7358 PAD.n8428 VSS 0.069752f
C7359 PAD.n8429 VSS 0.069752f
C7360 PAD.n8430 VSS 0.700403f
C7361 PAD.n8431 VSS 0.473511f
C7362 PAD.n8432 VSS 0.037175f
C7363 PAD.n8433 VSS 0.037175f
C7364 PAD.n8434 VSS 0.029431f
C7365 PAD.n8435 VSS 0.036484f
C7366 PAD.n8436 VSS 0.031863f
C7367 PAD.n8437 VSS 0.033766f
C7368 PAD.n8438 VSS 0.03055f
C7369 PAD.n8439 VSS 0.036454f
C7370 PAD.n8440 VSS 0.036454f
C7371 PAD.n8441 VSS 0.036454f
C7372 PAD.n8443 VSS 0.023105f
C7373 PAD.n8444 VSS 0.054256f
C7374 PAD.n8445 VSS 0.660944f
C7375 PAD.n8446 VSS 0.057377f
C7376 PAD.n8447 VSS 0.057377f
C7377 PAD.n8448 VSS 0.051216f
C7378 PAD.n8449 VSS 0.062262f
C7379 PAD.n8450 VSS 0.049207f
C7380 PAD.n8451 VSS 0.055127f
C7381 PAD.n8452 VSS 0.055127f
C7382 PAD.n8453 VSS 0.582025f
C7383 PAD.n8454 VSS 0.611619f
C7384 PAD.n8455 VSS 0.049106f
C7385 PAD.n8456 VSS 0.03268f
C7386 PAD.n8457 VSS 0.03268f
C7387 PAD.n8458 VSS 0.029431f
C7388 PAD.n8459 VSS 0.040979f
C7389 PAD.n8460 VSS 0.03579f
C7390 PAD.n8461 VSS 0.033766f
C7391 PAD.n8462 VSS 0.03055f
C7392 PAD.n8463 VSS 0.036454f
C7393 PAD.n8464 VSS 0.036454f
C7394 PAD.n8465 VSS 0.036454f
C7395 PAD.n8467 VSS 0.023105f
C7396 PAD.n8468 VSS 0.212094f
C7397 PAD.n8469 VSS 0.582025f
C7398 PAD.n8470 VSS 0.049502f
C7399 PAD.n8471 VSS 0.049502f
C7400 PAD.n8472 VSS 0.02134f
C7401 PAD.n8473 VSS 8.77683f
C7402 PAD.n8474 VSS 0.053977f
C7403 PAD.n8475 VSS 0.056237f
C7404 PAD.n8476 VSS 0.063002f
C7405 PAD.n8477 VSS 0.063002f
C7406 PAD.n8478 VSS 0.424187f
C7407 PAD.n8479 VSS 0.611619f
C7408 PAD.n8480 VSS 0.049106f
C7409 PAD.n8481 VSS 0.028184f
C7410 PAD.n8482 VSS 0.028184f
C7411 PAD.n8483 VSS 0.024615f
C7412 PAD.n8484 VSS 0.039716f
C7413 PAD.n8485 VSS 0.033766f
C7414 PAD.n8486 VSS 0.03055f
C7415 PAD.n8487 VSS 0.036454f
C7416 PAD.n8488 VSS 0.036454f
C7417 PAD.n8489 VSS 0.036454f
C7418 PAD.n8491 VSS 0.023105f
C7419 PAD.n8492 VSS 0.478444f
C7420 PAD.n8493 VSS 0.424187f
C7421 PAD.n8494 VSS 0.041626f
C7422 PAD.n8495 VSS 0.041626f
C7423 PAD.n8496 VSS 0.037156f
C7424 PAD.n8497 VSS 0.062262f
C7425 PAD.n8498 VSS 0.032135f
C7426 PAD.n8499 VSS 0.062262f
C7427 PAD.n8500 VSS 0.069752f
C7428 PAD.n8501 VSS 0.069752f
C7429 PAD.n8502 VSS 0.310742f
C7430 PAD.n8503 VSS 0.611619f
C7431 PAD.n8504 VSS 0.048241f
C7432 PAD.n8505 VSS 0.048241f
C7433 PAD.n8506 VSS 0.029431f
C7434 PAD.n8507 VSS 0.025417f
C7435 PAD.n8508 VSS 0.025417f
C7436 PAD.n8509 VSS 0.022199f
C7437 PAD.n8510 VSS 0.033766f
C7438 PAD.n8511 VSS 0.03055f
C7439 PAD.n8512 VSS 0.036454f
C7440 PAD.n8513 VSS 0.036454f
C7441 PAD.n8514 VSS 0.036454f
C7442 PAD.n8516 VSS 0.023105f
C7443 PAD.n8517 VSS 0.567228f
C7444 PAD.n8518 VSS 0.611619f
C7445 PAD.n8519 VSS 0.389661f
C7446 PAD.n8520 VSS 0.068627f
C7447 PAD.n8521 VSS 0.068627f
C7448 PAD.n8522 VSS 0.061258f
C7449 PAD.n8523 VSS 0.062262f
C7450 PAD.n8524 VSS 0.039165f
C7451 PAD.n8525 VSS 0.043876f
C7452 PAD.n8526 VSS 0.043876f
C7453 PAD.n8527 VSS 0.202229f
C7454 PAD.n8528 VSS 0.036454f
C7455 PAD.n8529 VSS 0.036454f
C7456 PAD.n8530 VSS 0.036454f
C7457 PAD.n8531 VSS 0.036454f
C7458 PAD.n8532 VSS 0.036454f
C7459 PAD.n8533 VSS 0.036454f
C7460 PAD.n8534 VSS 0.036454f
C7461 PAD.n8535 VSS 0.036454f
C7462 PAD.n8536 VSS 0.036454f
C7463 PAD.n8537 VSS 0.036454f
C7464 PAD.n8538 VSS 0.036454f
C7465 PAD.n8539 VSS 0.036454f
C7466 PAD.n8540 VSS 0.036454f
C7467 PAD.n8541 VSS 0.036454f
C7468 PAD.n8542 VSS 0.036454f
C7469 PAD.n8543 VSS 0.036454f
C7470 PAD.n8544 VSS 0.036454f
C7471 PAD.n8545 VSS 0.036454f
C7472 PAD.n8546 VSS 0.036454f
C7473 PAD.n8547 VSS 0.036454f
C7474 PAD.n8548 VSS 0.036454f
C7475 PAD.n8549 VSS 0.036454f
C7476 PAD.n8550 VSS 0.036454f
C7477 PAD.n8551 VSS 0.036454f
C7478 PAD.n8552 VSS 0.036454f
C7479 PAD.n8553 VSS 0.036454f
C7480 PAD.n8554 VSS 0.036454f
C7481 PAD.n8555 VSS 0.036454f
C7482 PAD.n8556 VSS 0.036454f
C7483 PAD.n8557 VSS 0.036454f
C7484 PAD.n8558 VSS 0.036454f
C7485 PAD.n8559 VSS 0.036454f
C7486 PAD.n8560 VSS 0.036454f
C7487 PAD.n8561 VSS 0.036454f
C7488 PAD.n8562 VSS 0.036454f
C7489 PAD.n8563 VSS 0.036454f
C7490 PAD.n8564 VSS 0.036454f
C7491 PAD.n8565 VSS 0.036454f
C7492 PAD.n8566 VSS 0.036454f
C7493 PAD.n8567 VSS 0.036454f
C7494 PAD.n8568 VSS 0.036454f
C7495 PAD.n8569 VSS 0.036454f
C7496 PAD.n8570 VSS 0.023105f
C7497 PAD.n8571 VSS 0.023105f
C7498 PAD.n8572 VSS 0.036454f
C7499 PAD.n8574 VSS 0.036454f
C7500 PAD.n8575 VSS 0.036454f
C7501 PAD.n8576 VSS 0.036454f
C7502 PAD.n8577 VSS 0.036454f
C7503 PAD.n8578 VSS 0.036454f
C7504 PAD.n8579 VSS 0.036454f
C7505 PAD.n8580 VSS 0.036454f
C7506 PAD.n8582 VSS 0.036454f
C7507 PAD.n8583 VSS 0.036454f
C7508 PAD.n8584 VSS 0.036454f
C7509 PAD.n8586 VSS 0.036454f
C7510 PAD.n8587 VSS 0.036454f
C7511 PAD.n8588 VSS 0.036454f
C7512 PAD.n8589 VSS 0.036454f
C7513 PAD.n8590 VSS 0.036454f
C7514 PAD.n8591 VSS 0.036454f
C7515 PAD.n8592 VSS 0.036454f
C7516 PAD.n8594 VSS 0.036454f
C7517 PAD.n8595 VSS 0.036454f
C7518 PAD.n8596 VSS 0.036454f
C7519 PAD.n8598 VSS 0.036454f
C7520 PAD.n8599 VSS 0.036454f
C7521 PAD.n8600 VSS 0.036454f
C7522 PAD.n8601 VSS 0.036454f
C7523 PAD.n8602 VSS 0.036454f
C7524 PAD.n8603 VSS 0.036454f
C7525 PAD.n8604 VSS 0.036454f
C7526 PAD.n8606 VSS 0.036454f
C7527 PAD.n8607 VSS 0.036454f
C7528 PAD.n8608 VSS 0.036454f
C7529 PAD.n8610 VSS 0.036454f
C7530 PAD.n8611 VSS 0.036454f
C7531 PAD.n8612 VSS 0.036454f
C7532 PAD.n8613 VSS 0.036454f
C7533 PAD.n8614 VSS 0.036454f
C7534 PAD.n8615 VSS 0.036454f
C7535 PAD.n8616 VSS 0.036454f
C7536 PAD.n8618 VSS 0.036454f
C7537 PAD.n8619 VSS 0.036454f
C7538 PAD.n8620 VSS 0.036454f
C7539 PAD.n8622 VSS 0.036454f
C7540 PAD.n8623 VSS 0.036454f
C7541 PAD.n8624 VSS 0.036454f
C7542 PAD.n8625 VSS 0.036454f
C7543 PAD.n8626 VSS 0.036454f
C7544 PAD.n8627 VSS 0.036454f
C7545 PAD.n8628 VSS 0.036454f
C7546 PAD.n8630 VSS 0.036454f
C7547 PAD.n8631 VSS 0.036454f
C7548 PAD.n8632 VSS 0.036454f
C7549 PAD.n8634 VSS 0.036454f
C7550 PAD.n8635 VSS 0.036454f
C7551 PAD.n8636 VSS 0.036454f
C7552 PAD.n8637 VSS 0.036454f
C7553 PAD.n8638 VSS 0.036454f
C7554 PAD.n8639 VSS 0.036454f
C7555 PAD.n8640 VSS 0.036454f
C7556 PAD.n8642 VSS 0.036454f
C7557 PAD.n8643 VSS 0.036454f
C7558 PAD.n8644 VSS 0.036454f
C7559 PAD.n8646 VSS 0.036454f
C7560 PAD.n8647 VSS 0.036454f
C7561 PAD.n8648 VSS 0.036454f
C7562 PAD.n8649 VSS 0.036454f
C7563 PAD.n8650 VSS 0.036454f
C7564 PAD.n8651 VSS 0.036454f
C7565 PAD.n8652 VSS 0.036454f
C7566 PAD.n8654 VSS 0.036454f
C7567 PAD.n8655 VSS 0.036454f
C7568 PAD.n8656 VSS 0.036454f
C7569 PAD.n8658 VSS 0.036454f
C7570 PAD.n8659 VSS 0.036454f
C7571 PAD.n8660 VSS 0.036454f
C7572 PAD.n8661 VSS 0.036454f
C7573 PAD.n8662 VSS 0.036454f
C7574 PAD.n8663 VSS 0.036454f
C7575 PAD.n8664 VSS 0.036454f
C7576 PAD.n8666 VSS 0.036454f
C7577 PAD.n8667 VSS 0.036454f
C7578 PAD.n8668 VSS 0.036454f
C7579 PAD.n8670 VSS 0.036454f
C7580 PAD.n8671 VSS 0.036454f
C7581 PAD.n8672 VSS 0.036454f
C7582 PAD.n8673 VSS 0.036454f
C7583 PAD.n8674 VSS 0.036454f
C7584 PAD.n8675 VSS 0.036454f
C7585 PAD.n8676 VSS 0.036454f
C7586 PAD.n8678 VSS 0.036454f
C7587 PAD.n8679 VSS 0.036454f
C7588 PAD.n8680 VSS 0.036454f
C7589 PAD.n8682 VSS 0.036454f
C7590 PAD.n8683 VSS 0.036454f
C7591 PAD.n8684 VSS 0.036454f
C7592 PAD.n8685 VSS 0.036454f
C7593 PAD.n8686 VSS 0.036454f
C7594 PAD.n8687 VSS 0.036454f
C7595 PAD.n8688 VSS 0.036454f
C7596 PAD.n8690 VSS 0.036454f
C7597 PAD.n8691 VSS 0.036454f
C7598 PAD.n8692 VSS 0.036454f
C7599 PAD.n8694 VSS 0.036454f
C7600 PAD.n8695 VSS 0.036454f
C7601 PAD.n8696 VSS 0.036454f
C7602 PAD.n8697 VSS 0.036454f
C7603 PAD.n8698 VSS 0.036454f
C7604 PAD.n8699 VSS 0.036454f
C7605 PAD.n8700 VSS 0.036454f
C7606 PAD.n8702 VSS 0.036454f
C7607 PAD.n8703 VSS 0.036454f
C7608 PAD.n8704 VSS 0.036454f
C7609 PAD.n8706 VSS 0.036454f
C7610 PAD.n8707 VSS 0.036454f
C7611 PAD.n8708 VSS 0.036454f
C7612 PAD.n8709 VSS 0.036454f
C7613 PAD.n8710 VSS 0.036454f
C7614 PAD.n8711 VSS 0.036454f
C7615 PAD.n8712 VSS 0.036454f
C7616 PAD.n8714 VSS 0.036454f
C7617 PAD.n8715 VSS 0.036454f
C7618 PAD.n8716 VSS 0.036454f
C7619 PAD.n8718 VSS 0.036454f
C7620 PAD.n8719 VSS 0.036454f
C7621 PAD.n8720 VSS 0.036454f
C7622 PAD.n8721 VSS 0.036454f
C7623 PAD.n8722 VSS 0.036454f
C7624 PAD.n8723 VSS 0.036454f
C7625 PAD.n8724 VSS 0.036454f
C7626 PAD.n8726 VSS 0.036454f
C7627 PAD.n8727 VSS 0.036454f
C7628 PAD.n8728 VSS 0.036454f
C7629 PAD.n8730 VSS 0.036454f
C7630 PAD.n8731 VSS 0.036454f
C7631 PAD.n8732 VSS 0.036454f
C7632 PAD.n8733 VSS 0.036454f
C7633 PAD.n8734 VSS 0.036454f
C7634 PAD.n8735 VSS 0.036454f
C7635 PAD.n8736 VSS 0.036454f
C7636 PAD.n8738 VSS 0.036454f
C7637 PAD.n8739 VSS 0.036454f
C7638 PAD.n8740 VSS 0.036454f
C7639 PAD.n8742 VSS 0.036454f
C7640 PAD.n8743 VSS 0.036454f
C7641 PAD.n8744 VSS 0.036454f
C7642 PAD.n8745 VSS 0.036454f
C7643 PAD.n8746 VSS 0.036454f
C7644 PAD.n8747 VSS 0.036454f
C7645 PAD.n8748 VSS 0.036454f
C7646 PAD.n8750 VSS 0.036454f
C7647 PAD.n8751 VSS 0.036454f
C7648 PAD.n8752 VSS 0.036454f
C7649 PAD.n8754 VSS 0.036454f
C7650 PAD.n8755 VSS 0.036454f
C7651 PAD.n8756 VSS 0.036454f
C7652 PAD.n8757 VSS 0.036454f
C7653 PAD.n8758 VSS 0.036454f
C7654 PAD.n8759 VSS 0.036454f
C7655 PAD.n8760 VSS 0.036454f
C7656 PAD.n8762 VSS 0.036454f
C7657 PAD.n8763 VSS 0.036454f
C7658 PAD.n8764 VSS 0.036454f
C7659 PAD.n8766 VSS 0.036454f
C7660 PAD.n8767 VSS 0.036454f
C7661 PAD.n8768 VSS 0.036454f
C7662 PAD.n8769 VSS 0.036454f
C7663 PAD.n8770 VSS 0.036454f
C7664 PAD.n8771 VSS 0.036454f
C7665 PAD.n8772 VSS 0.036454f
C7666 PAD.n8774 VSS 0.036454f
C7667 PAD.n8775 VSS 0.036454f
C7668 PAD.n8776 VSS 0.036454f
C7669 PAD.n8778 VSS 0.036454f
C7670 PAD.n8779 VSS 0.036454f
C7671 PAD.n8780 VSS 0.036454f
C7672 PAD.n8781 VSS 0.036454f
C7673 PAD.n8782 VSS 0.036454f
C7674 PAD.n8783 VSS 0.036454f
C7675 PAD.n8784 VSS 0.036454f
C7676 PAD.n8786 VSS 0.036454f
C7677 PAD.n8787 VSS 0.036454f
C7678 PAD.n8788 VSS 0.036454f
C7679 PAD.n8790 VSS 0.036454f
C7680 PAD.n8791 VSS 0.036454f
C7681 PAD.n8792 VSS 0.036454f
C7682 PAD.n8793 VSS 0.036454f
C7683 PAD.n8794 VSS 0.036454f
C7684 PAD.n8795 VSS 0.036454f
C7685 PAD.n8796 VSS 0.036454f
C7686 PAD.n8798 VSS 0.036454f
C7687 PAD.n8799 VSS 0.036454f
C7688 PAD.n8800 VSS 0.036454f
C7689 PAD.n8802 VSS 0.036454f
C7690 PAD.n8803 VSS 0.036454f
C7691 PAD.n8804 VSS 0.036454f
C7692 PAD.n8805 VSS 0.036454f
C7693 PAD.n8806 VSS 0.036454f
C7694 PAD.n8807 VSS 0.036454f
C7695 PAD.n8808 VSS 0.036454f
C7696 PAD.n8810 VSS 0.036454f
C7697 PAD.n8811 VSS 0.036454f
C7698 PAD.n8813 VSS 0.036454f
C7699 PAD.n8814 VSS 0.036454f
C7700 PAD.n8815 VSS 0.036454f
C7701 PAD.n8816 VSS 0.036454f
C7702 PAD.n8817 VSS 0.033374f
C7703 PAD.n8818 VSS 0.023105f
C7704 PAD.n8819 VSS 0.023105f
C7705 PAD.n8821 VSS 0.389661f
C7706 PAD.n8822 VSS 0.414322f
C7707 PAD.n8823 VSS 0.043746f
C7708 PAD.n8824 VSS 0.043746f
C7709 PAD.n8825 VSS 0.038206f
C7710 PAD.n8826 VSS 0.033766f
C7711 PAD.n8827 VSS 0.026125f
C7712 PAD.n8828 VSS 0.042887f
C7713 PAD.n8829 VSS 0.049106f
C7714 PAD.n8830 VSS 0.049106f
C7715 PAD.n8831 VSS 0.611619f
C7716 PAD.n8832 VSS 0.508039f
C7717 PAD.n8833 VSS 0.060752f
C7718 PAD.n8834 VSS 0.060752f
C7719 PAD.n8835 VSS 0.054228f
C7720 PAD.n8836 VSS 0.062262f
C7721 PAD.n8837 VSS 0.036454f
C7722 PAD.n8838 VSS 0.036454f
C7723 PAD.n8839 VSS 0.036454f
C7724 PAD.n8841 VSS 0.036454f
C7725 PAD.n8842 VSS 0.036454f
C7726 PAD.n8843 VSS 0.036454f
C7727 PAD.n8844 VSS 0.036454f
C7728 PAD.n8846 VSS 0.036454f
C7729 PAD.n8847 VSS 0.036454f
C7730 PAD.n8848 VSS 0.036454f
C7731 PAD.n8849 VSS 0.036454f
C7732 PAD.n8851 VSS 0.036454f
C7733 PAD.n8852 VSS 0.036454f
C7734 PAD.n8853 VSS 0.036454f
C7735 PAD.n8854 VSS 0.036454f
C7736 PAD.n8856 VSS 0.036454f
C7737 PAD.n8857 VSS 0.036454f
C7738 PAD.n8858 VSS 0.036454f
C7739 PAD.n8859 VSS 0.036454f
C7740 PAD.n8861 VSS 0.036454f
C7741 PAD.n8862 VSS 0.036454f
C7742 PAD.n8863 VSS 0.036454f
C7743 PAD.n8864 VSS 0.036454f
C7744 PAD.n8866 VSS 0.036454f
C7745 PAD.n8867 VSS 0.036454f
C7746 PAD.n8868 VSS 0.036454f
C7747 PAD.n8869 VSS 0.036454f
C7748 PAD.n8871 VSS 0.036454f
C7749 PAD.n8872 VSS 0.036454f
C7750 PAD.n8873 VSS 0.036454f
C7751 PAD.n8874 VSS 0.036454f
C7752 PAD.n8876 VSS 0.036454f
C7753 PAD.n8877 VSS 0.036454f
C7754 PAD.n8878 VSS 0.036454f
C7755 PAD.n8879 VSS 0.036454f
C7756 PAD.n8881 VSS 0.036454f
C7757 PAD.n8882 VSS 0.036454f
C7758 PAD.n8883 VSS 0.036454f
C7759 PAD.n8884 VSS 0.036454f
C7760 PAD.n8886 VSS 0.036454f
C7761 PAD.n8887 VSS 0.036454f
C7762 PAD.n8888 VSS 0.036454f
C7763 PAD.n8889 VSS 0.036454f
C7764 PAD.n8891 VSS 0.036454f
C7765 PAD.n8892 VSS 0.036454f
C7766 PAD.n8893 VSS 0.036454f
C7767 PAD.n8894 VSS 0.036454f
C7768 PAD.n8896 VSS 0.036454f
C7769 PAD.n8897 VSS 0.036454f
C7770 PAD.n8898 VSS 0.036454f
C7771 PAD.n8899 VSS 0.036454f
C7772 PAD.n8901 VSS 0.036454f
C7773 PAD.n8902 VSS 0.036454f
C7774 PAD.n8903 VSS 0.036454f
C7775 PAD.n8904 VSS 0.036454f
C7776 PAD.n8906 VSS 0.036454f
C7777 PAD.n8907 VSS 0.036454f
C7778 PAD.n8908 VSS 0.036454f
C7779 PAD.n8909 VSS 0.036454f
C7780 PAD.n8911 VSS 0.036454f
C7781 PAD.n8912 VSS 0.036454f
C7782 PAD.n8913 VSS 0.036454f
C7783 PAD.n8914 VSS 0.036454f
C7784 PAD.n8916 VSS 0.036454f
C7785 PAD.n8917 VSS 0.036454f
C7786 PAD.n8918 VSS 0.036454f
C7787 PAD.n8919 VSS 0.036454f
C7788 PAD.n8921 VSS 0.036454f
C7789 PAD.n8922 VSS 0.036454f
C7790 PAD.n8923 VSS 0.036454f
C7791 PAD.n8924 VSS 0.036454f
C7792 PAD.n8926 VSS 0.036454f
C7793 PAD.n8927 VSS 0.036454f
C7794 PAD.n8928 VSS 0.036454f
C7795 PAD.n8929 VSS 0.036454f
C7796 PAD.n8931 VSS 0.036454f
C7797 PAD.n8932 VSS 0.036454f
C7798 PAD.n8933 VSS 0.036454f
C7799 PAD.n8934 VSS 0.036454f
C7800 PAD.n8936 VSS 0.036454f
C7801 PAD.n8937 VSS 0.036454f
C7802 PAD.n8939 VSS 0.036454f
C7803 PAD.n8940 VSS 0.036454f
C7804 PAD.n8941 VSS 0.036454f
C7805 PAD.n8942 VSS 0.036454f
C7806 PAD.n8943 VSS 0.036454f
C7807 PAD.n8944 VSS 0.036454f
C7808 PAD.n8945 VSS 0.036454f
C7809 PAD.n8946 VSS 0.036454f
C7810 PAD.n8948 VSS 0.036454f
C7811 PAD.n8949 VSS 0.036454f
C7812 PAD.n8950 VSS 0.036454f
C7813 PAD.n8951 VSS 0.036454f
C7814 PAD.n8952 VSS 0.036454f
C7815 PAD.n8953 VSS 0.036454f
C7816 PAD.n8954 VSS 0.036454f
C7817 PAD.n8955 VSS 0.036454f
C7818 PAD.n8957 VSS 0.036454f
C7819 PAD.n8958 VSS 0.036454f
C7820 PAD.n8959 VSS 0.036454f
C7821 PAD.n8960 VSS 0.036454f
C7822 PAD.n8961 VSS 0.036454f
C7823 PAD.n8962 VSS 0.036454f
C7824 PAD.n8963 VSS 0.036454f
C7825 PAD.n8964 VSS 0.036454f
C7826 PAD.n8966 VSS 0.036454f
C7827 PAD.n8967 VSS 0.036454f
C7828 PAD.n8968 VSS 0.036454f
C7829 PAD.n8969 VSS 0.036454f
C7830 PAD.n8970 VSS 0.036454f
C7831 PAD.n8971 VSS 0.036454f
C7832 PAD.n8972 VSS 0.036454f
C7833 PAD.n8973 VSS 0.036454f
C7834 PAD.n8975 VSS 0.036454f
C7835 PAD.n8976 VSS 0.036454f
C7836 PAD.n8977 VSS 0.036454f
C7837 PAD.n8978 VSS 0.036454f
C7838 PAD.n8979 VSS 0.036454f
C7839 PAD.n8980 VSS 0.036454f
C7840 PAD.n8981 VSS 0.036454f
C7841 PAD.n8982 VSS 0.036454f
C7842 PAD.n8984 VSS 0.036454f
C7843 PAD.n8985 VSS 0.036454f
C7844 PAD.n8986 VSS 0.036454f
C7845 PAD.n8987 VSS 0.036454f
C7846 PAD.n8988 VSS 0.036454f
C7847 PAD.n8989 VSS 0.036454f
C7848 PAD.n8990 VSS 0.036454f
C7849 PAD.n8991 VSS 0.036454f
C7850 PAD.n8993 VSS 0.036454f
C7851 PAD.n8994 VSS 0.036454f
C7852 PAD.n8995 VSS 0.036454f
C7853 PAD.n8996 VSS 0.036454f
C7854 PAD.n8997 VSS 0.036454f
C7855 PAD.n8998 VSS 0.036454f
C7856 PAD.n8999 VSS 0.036454f
C7857 PAD.n9000 VSS 0.036454f
C7858 PAD.n9002 VSS 0.036454f
C7859 PAD.n9003 VSS 0.036454f
C7860 PAD.n9004 VSS 0.036454f
C7861 PAD.n9005 VSS 0.036454f
C7862 PAD.n9006 VSS 0.036454f
C7863 PAD.n9007 VSS 0.036454f
C7864 PAD.n9008 VSS 0.036454f
C7865 PAD.n9009 VSS 0.036454f
C7866 PAD.n9011 VSS 0.036454f
C7867 PAD.n9012 VSS 0.036454f
C7868 PAD.n9013 VSS 0.036454f
C7869 PAD.n9014 VSS 0.036454f
C7870 PAD.n9015 VSS 0.036454f
C7871 PAD.n9016 VSS 0.036454f
C7872 PAD.n9017 VSS 0.036454f
C7873 PAD.n9018 VSS 0.036454f
C7874 PAD.n9020 VSS 0.036454f
C7875 PAD.n9021 VSS 0.036454f
C7876 PAD.n9022 VSS 0.036454f
C7877 PAD.n9023 VSS 0.036454f
C7878 PAD.n9024 VSS 0.036454f
C7879 PAD.n9025 VSS 0.036454f
C7880 PAD.n9026 VSS 0.036454f
C7881 PAD.n9027 VSS 0.036454f
C7882 PAD.n9029 VSS 0.036454f
C7883 PAD.n9030 VSS 0.036454f
C7884 PAD.n9031 VSS 0.036454f
C7885 PAD.n9032 VSS 0.036454f
C7886 PAD.n9033 VSS 0.036454f
C7887 PAD.n9034 VSS 0.036454f
C7888 PAD.n9035 VSS 0.036454f
C7889 PAD.n9036 VSS 0.036454f
C7890 PAD.n9038 VSS 0.036454f
C7891 PAD.n9039 VSS 0.036454f
C7892 PAD.n9040 VSS 0.036454f
C7893 PAD.n9041 VSS 0.036454f
C7894 PAD.n9042 VSS 0.036454f
C7895 PAD.n9043 VSS 0.036454f
C7896 PAD.n9044 VSS 0.036454f
C7897 PAD.n9045 VSS 0.036454f
C7898 PAD.n9047 VSS 0.036454f
C7899 PAD.n9048 VSS 0.036454f
C7900 PAD.n9049 VSS 0.036454f
C7901 PAD.n9050 VSS 0.036454f
C7902 PAD.n9051 VSS 0.036454f
C7903 PAD.n9052 VSS 0.036454f
C7904 PAD.n9053 VSS 0.036454f
C7905 PAD.n9054 VSS 0.036454f
C7906 PAD.n9056 VSS 0.036454f
C7907 PAD.n9057 VSS 0.036454f
C7908 PAD.n9058 VSS 0.036454f
C7909 PAD.n9059 VSS 0.036454f
C7910 PAD.n9060 VSS 0.036454f
C7911 PAD.n9061 VSS 0.036454f
C7912 PAD.n9062 VSS 0.036454f
C7913 PAD.n9063 VSS 0.036454f
C7914 PAD.n9065 VSS 0.036454f
C7915 PAD.n9066 VSS 0.036454f
C7916 PAD.n9067 VSS 0.036454f
C7917 PAD.n9068 VSS 0.036454f
C7918 PAD.n9069 VSS 0.036454f
C7919 PAD.n9070 VSS 0.036454f
C7920 PAD.n9071 VSS 0.036454f
C7921 PAD.n9072 VSS 0.036454f
C7922 PAD.n9074 VSS 0.036454f
C7923 PAD.n9075 VSS 0.036454f
C7924 PAD.n9076 VSS 0.036454f
C7925 PAD.n9077 VSS 0.036454f
C7926 PAD.n9078 VSS 0.036454f
C7927 PAD.n9079 VSS 0.036454f
C7928 PAD.n9080 VSS 0.036454f
C7929 PAD.n9081 VSS 0.036454f
C7930 PAD.n9083 VSS 0.036454f
C7931 PAD.n9084 VSS 0.036454f
C7932 PAD.n9085 VSS 0.036454f
C7933 PAD.n9086 VSS 0.036454f
C7934 PAD.n9087 VSS 0.036454f
C7935 PAD.n9088 VSS 0.036454f
C7936 PAD.n9089 VSS 0.036454f
C7937 PAD.n9090 VSS 0.036454f
C7938 PAD.n9092 VSS 0.036454f
C7939 PAD.n9093 VSS 0.036454f
C7940 PAD.n9094 VSS 0.036454f
C7941 PAD.n9095 VSS 0.036454f
C7942 PAD.n9096 VSS 0.036454f
C7943 PAD.n9097 VSS 0.036454f
C7944 PAD.n9098 VSS 0.036454f
C7945 PAD.n9099 VSS 0.036454f
C7946 PAD.n9101 VSS 0.036454f
C7947 PAD.n9102 VSS 0.036454f
C7948 PAD.n9103 VSS 0.036454f
C7949 PAD.n9104 VSS 0.036454f
C7950 PAD.n9105 VSS 0.036454f
C7951 PAD.n9106 VSS 0.036454f
C7952 PAD.n9107 VSS 0.036454f
C7953 PAD.n9108 VSS 0.036454f
C7954 PAD.n9110 VSS 0.036454f
C7955 PAD.n9111 VSS 0.036454f
C7956 PAD.n9112 VSS 0.036454f
C7957 PAD.n9113 VSS 0.036454f
C7958 PAD.n9114 VSS 0.036454f
C7959 PAD.n9115 VSS 0.036454f
C7960 PAD.n9117 VSS 0.036454f
C7961 PAD.n9118 VSS 0.036454f
C7962 PAD.n9119 VSS 0.023105f
C7963 PAD.n9120 VSS 0.033374f
C7964 PAD.n9121 VSS 0.052877f
C7965 PAD.n9122 VSS 0.052877f
C7966 PAD.n9123 VSS 0.047199f
C7967 PAD.n9124 VSS 0.046278f
C7968 PAD.n9125 VSS 0.046195f
C7969 PAD.n9126 VSS 0.051752f
C7970 PAD.n9127 VSS 0.051752f
C7971 PAD.n9128 VSS 0.621484f
C7972 PAD.n9129 VSS 0.611619f
C7973 PAD.n9130 VSS 0.034409f
C7974 PAD.n9131 VSS 0.034409f
C7975 PAD.n9132 VSS 0.030051f
C7976 PAD.n9133 VSS 0.033766f
C7977 PAD.n9134 VSS 0.03055f
C7978 PAD.n9135 VSS 0.036454f
C7979 PAD.n9136 VSS 0.036454f
C7980 PAD.n9137 VSS 0.036454f
C7981 PAD.n9139 VSS 0.023105f
C7982 PAD.n9140 VSS 0.611619f
C7983 PAD.n9141 VSS 0.621484f
C7984 PAD.n9142 VSS 0.611619f
C7985 PAD.n9143 VSS 0.636282f
C7986 PAD.n9144 VSS 0.059627f
C7987 PAD.n9145 VSS 0.059627f
C7988 PAD.n9146 VSS 0.053224f
C7989 PAD.n9147 VSS 0.046278f
C7990 PAD.n9148 VSS 0.040169f
C7991 PAD.n9149 VSS 0.045001f
C7992 PAD.n9150 VSS 0.045001f
C7993 PAD.n9151 VSS 0.636282f
C7994 PAD.n9152 VSS 0.5327f
C7995 PAD.n9153 VSS 0.034755f
C7996 PAD.n9154 VSS 0.034755f
C7997 PAD.n9155 VSS 0.030353f
C7998 PAD.n9156 VSS 0.033766f
C7999 PAD.n9157 VSS 0.033978f
C8000 PAD.n9158 VSS 0.038904f
C8001 PAD.n9159 VSS 0.038904f
C8002 PAD.n9160 VSS 0.443917f
C8003 PAD.n9161 VSS 0.700403f
C8004 PAD.n9162 VSS 0.611619f
C8005 PAD.n9163 VSS 0.493241f
C8006 PAD.n9164 VSS 0.067502f
C8007 PAD.n9165 VSS 0.067502f
C8008 PAD.n9166 VSS 0.060254f
C8009 PAD.n9167 VSS 0.046278f
C8010 PAD.n9168 VSS 14.504801f
C8011 PAD.n9169 VSS 0.062262f
C8012 PAD.n9170 VSS 0.055735f
C8013 PAD.n9171 VSS 8.7754f
C8014 PAD.n9172 VSS 0.008536f
C8015 PAD.n9173 VSS 0.037126f
C8016 PAD.n9174 VSS 0.037126f
C8017 PAD.n9175 VSS 0.493241f
C8018 PAD.n9176 VSS 0.40939f
C8019 PAD.n9177 VSS 0.030259f
C8020 PAD.n9178 VSS 0.030259f
C8021 PAD.n9179 VSS 0.026427f
C8022 PAD.n9180 VSS 0.033766f
C8023 PAD.n9181 VSS 0.037904f
C8024 PAD.n9182 VSS 0.0434f
C8025 PAD.n9183 VSS 0.0434f
C8026 PAD.n9184 VSS 0.320607f
C8027 PAD.n9185 VSS 0.700403f
C8028 PAD.n9186 VSS 0.611619f
C8029 PAD.n9187 VSS 0.389661f
C8030 PAD.n9188 VSS 0.069752f
C8031 PAD.n9189 VSS 0.039754f
C8032 PAD.n9190 VSS 0.040501f
C8033 PAD.n9191 VSS 0.040501f
C8034 PAD.n9192 VSS 0.043182f
C8035 PAD.n9193 VSS 0.062262f
C8036 PAD.n9194 VSS 0.057241f
C8037 PAD.n9195 VSS 0.064127f
C8038 PAD.n9196 VSS 0.039754f
C8039 PAD.n9197 VSS 0.023105f
C8040 PAD.n9198 VSS 0.033374f
C8041 PAD.n9199 VSS 0.036454f
C8042 PAD.n9200 VSS 0.036454f
C8043 PAD.n9201 VSS 0.036454f
C8044 PAD.n9202 VSS 0.036454f
C8045 PAD.n9204 VSS 0.036454f
C8046 PAD.n9205 VSS 0.036454f
C8047 PAD.n9206 VSS 0.036454f
C8048 PAD.n9208 VSS 0.036454f
C8049 PAD.n9209 VSS 0.036454f
C8050 PAD.n9210 VSS 0.036454f
C8051 PAD.n9211 VSS 0.036454f
C8052 PAD.n9212 VSS 0.036454f
C8053 PAD.n9213 VSS 0.036454f
C8054 PAD.n9214 VSS 0.036454f
C8055 PAD.n9216 VSS 0.036454f
C8056 PAD.n9217 VSS 0.036454f
C8057 PAD.n9218 VSS 0.036454f
C8058 PAD.n9220 VSS 0.036454f
C8059 PAD.n9221 VSS 0.036454f
C8060 PAD.n9222 VSS 0.036454f
C8061 PAD.n9223 VSS 0.036454f
C8062 PAD.n9224 VSS 0.036454f
C8063 PAD.n9225 VSS 0.036454f
C8064 PAD.n9226 VSS 0.036454f
C8065 PAD.n9228 VSS 0.036454f
C8066 PAD.n9229 VSS 0.036454f
C8067 PAD.n9230 VSS 0.036454f
C8068 PAD.n9232 VSS 0.036454f
C8069 PAD.n9233 VSS 0.036454f
C8070 PAD.n9234 VSS 0.036454f
C8071 PAD.n9235 VSS 0.036454f
C8072 PAD.n9236 VSS 0.036454f
C8073 PAD.n9237 VSS 0.036454f
C8074 PAD.n9238 VSS 0.036454f
C8075 PAD.n9240 VSS 0.036454f
C8076 PAD.n9241 VSS 0.036454f
C8077 PAD.n9242 VSS 0.036454f
C8078 PAD.n9244 VSS 0.036454f
C8079 PAD.n9245 VSS 0.036454f
C8080 PAD.n9246 VSS 0.036454f
C8081 PAD.n9247 VSS 0.036454f
C8082 PAD.n9248 VSS 0.036454f
C8083 PAD.n9249 VSS 0.036454f
C8084 PAD.n9250 VSS 0.036454f
C8085 PAD.n9252 VSS 0.036454f
C8086 PAD.n9253 VSS 0.036454f
C8087 PAD.n9254 VSS 0.036454f
C8088 PAD.n9256 VSS 0.036454f
C8089 PAD.n9257 VSS 0.036454f
C8090 PAD.n9258 VSS 0.036454f
C8091 PAD.n9259 VSS 0.036454f
C8092 PAD.n9260 VSS 0.036454f
C8093 PAD.n9261 VSS 0.036454f
C8094 PAD.n9262 VSS 0.036454f
C8095 PAD.n9264 VSS 0.036454f
C8096 PAD.n9265 VSS 0.036454f
C8097 PAD.n9266 VSS 0.036454f
C8098 PAD.n9268 VSS 0.036454f
C8099 PAD.n9269 VSS 0.036454f
C8100 PAD.n9270 VSS 0.036454f
C8101 PAD.n9271 VSS 0.036454f
C8102 PAD.n9272 VSS 0.036454f
C8103 PAD.n9273 VSS 0.036454f
C8104 PAD.n9274 VSS 0.036454f
C8105 PAD.n9276 VSS 0.036454f
C8106 PAD.n9277 VSS 0.036454f
C8107 PAD.n9278 VSS 0.036454f
C8108 PAD.n9280 VSS 0.036454f
C8109 PAD.n9281 VSS 0.036454f
C8110 PAD.n9282 VSS 0.036454f
C8111 PAD.n9283 VSS 0.036454f
C8112 PAD.n9284 VSS 0.036454f
C8113 PAD.n9285 VSS 0.036454f
C8114 PAD.n9286 VSS 0.036454f
C8115 PAD.n9288 VSS 0.036454f
C8116 PAD.n9289 VSS 0.036454f
C8117 PAD.n9290 VSS 0.036454f
C8118 PAD.n9292 VSS 0.036454f
C8119 PAD.n9293 VSS 0.036454f
C8120 PAD.n9294 VSS 0.036454f
C8121 PAD.n9295 VSS 0.036454f
C8122 PAD.n9296 VSS 0.036454f
C8123 PAD.n9297 VSS 0.036454f
C8124 PAD.n9298 VSS 0.036454f
C8125 PAD.n9300 VSS 0.036454f
C8126 PAD.n9301 VSS 0.036454f
C8127 PAD.n9302 VSS 0.036454f
C8128 PAD.n9304 VSS 0.036454f
C8129 PAD.n9305 VSS 0.036454f
C8130 PAD.n9306 VSS 0.036454f
C8131 PAD.n9307 VSS 0.036454f
C8132 PAD.n9308 VSS 0.036454f
C8133 PAD.n9309 VSS 0.036454f
C8134 PAD.n9310 VSS 0.036454f
C8135 PAD.n9312 VSS 0.036454f
C8136 PAD.n9313 VSS 0.036454f
C8137 PAD.n9314 VSS 0.036454f
C8138 PAD.n9316 VSS 0.036454f
C8139 PAD.n9317 VSS 0.036454f
C8140 PAD.n9318 VSS 0.036454f
C8141 PAD.n9319 VSS 0.036454f
C8142 PAD.n9320 VSS 0.036454f
C8143 PAD.n9321 VSS 0.036454f
C8144 PAD.n9322 VSS 0.036454f
C8145 PAD.n9324 VSS 0.036454f
C8146 PAD.n9325 VSS 0.036454f
C8147 PAD.n9326 VSS 0.036454f
C8148 PAD.n9328 VSS 0.036454f
C8149 PAD.n9329 VSS 0.036454f
C8150 PAD.n9330 VSS 0.036454f
C8151 PAD.n9331 VSS 0.036454f
C8152 PAD.n9332 VSS 0.036454f
C8153 PAD.n9333 VSS 0.036454f
C8154 PAD.n9334 VSS 0.036454f
C8155 PAD.n9336 VSS 0.036454f
C8156 PAD.n9337 VSS 0.036454f
C8157 PAD.n9338 VSS 0.036454f
C8158 PAD.n9340 VSS 0.036454f
C8159 PAD.n9341 VSS 0.036454f
C8160 PAD.n9342 VSS 0.036454f
C8161 PAD.n9343 VSS 0.036454f
C8162 PAD.n9344 VSS 0.036454f
C8163 PAD.n9345 VSS 0.036454f
C8164 PAD.n9346 VSS 0.036454f
C8165 PAD.n9348 VSS 0.036454f
C8166 PAD.n9349 VSS 0.036454f
C8167 PAD.n9350 VSS 0.036454f
C8168 PAD.n9352 VSS 0.036454f
C8169 PAD.n9353 VSS 0.036454f
C8170 PAD.n9354 VSS 0.036454f
C8171 PAD.n9355 VSS 0.036454f
C8172 PAD.n9356 VSS 0.036454f
C8173 PAD.n9357 VSS 0.036454f
C8174 PAD.n9358 VSS 0.036454f
C8175 PAD.n9360 VSS 0.036454f
C8176 PAD.n9361 VSS 0.036454f
C8177 PAD.n9362 VSS 0.036454f
C8178 PAD.n9364 VSS 0.036454f
C8179 PAD.n9365 VSS 0.036454f
C8180 PAD.n9366 VSS 0.036454f
C8181 PAD.n9367 VSS 0.036454f
C8182 PAD.n9368 VSS 0.036454f
C8183 PAD.n9369 VSS 0.036454f
C8184 PAD.n9370 VSS 0.036454f
C8185 PAD.n9372 VSS 0.036454f
C8186 PAD.n9373 VSS 0.036454f
C8187 PAD.n9374 VSS 0.036454f
C8188 PAD.n9376 VSS 0.036454f
C8189 PAD.n9377 VSS 0.036454f
C8190 PAD.n9378 VSS 0.036454f
C8191 PAD.n9379 VSS 0.036454f
C8192 PAD.n9380 VSS 0.036454f
C8193 PAD.n9381 VSS 0.036454f
C8194 PAD.n9382 VSS 0.036454f
C8195 PAD.n9384 VSS 0.036454f
C8196 PAD.n9385 VSS 0.036454f
C8197 PAD.n9386 VSS 0.036454f
C8198 PAD.n9388 VSS 0.036454f
C8199 PAD.n9389 VSS 0.036454f
C8200 PAD.n9390 VSS 0.036454f
C8201 PAD.n9391 VSS 0.036454f
C8202 PAD.n9392 VSS 0.036454f
C8203 PAD.n9393 VSS 0.036454f
C8204 PAD.n9394 VSS 0.036454f
C8205 PAD.n9396 VSS 0.036454f
C8206 PAD.n9397 VSS 0.036454f
C8207 PAD.n9398 VSS 0.036454f
C8208 PAD.n9400 VSS 0.036454f
C8209 PAD.n9401 VSS 0.036454f
C8210 PAD.n9402 VSS 0.036454f
C8211 PAD.n9403 VSS 0.036454f
C8212 PAD.n9404 VSS 0.036454f
C8213 PAD.n9405 VSS 0.036454f
C8214 PAD.n9406 VSS 0.036454f
C8215 PAD.n9408 VSS 0.036454f
C8216 PAD.n9409 VSS 0.036454f
C8217 PAD.n9410 VSS 0.036454f
C8218 PAD.n9412 VSS 0.036454f
C8219 PAD.n9413 VSS 0.036454f
C8220 PAD.n9414 VSS 0.036454f
C8221 PAD.n9415 VSS 0.036454f
C8222 PAD.n9416 VSS 0.036454f
C8223 PAD.n9417 VSS 0.036454f
C8224 PAD.n9418 VSS 0.036454f
C8225 PAD.n9420 VSS 0.036454f
C8226 PAD.n9421 VSS 0.036454f
C8227 PAD.n9422 VSS 0.036454f
C8228 PAD.n9424 VSS 0.036454f
C8229 PAD.n9425 VSS 0.036454f
C8230 PAD.n9426 VSS 0.036454f
C8231 PAD.n9427 VSS 0.036454f
C8232 PAD.n9428 VSS 0.036454f
C8233 PAD.n9429 VSS 0.036454f
C8234 PAD.n9430 VSS 0.036454f
C8235 PAD.n9432 VSS 0.036454f
C8236 PAD.n9433 VSS 0.036454f
C8237 PAD.n9434 VSS 0.036454f
C8238 PAD.n9436 VSS 0.036454f
C8239 PAD.n9437 VSS 0.036454f
C8240 PAD.n9438 VSS 0.036454f
C8241 PAD.n9439 VSS 0.036454f
C8242 PAD.n9440 VSS 0.036454f
C8243 PAD.n9441 VSS 0.036454f
C8244 PAD.n9442 VSS 0.036454f
C8245 PAD.n9444 VSS 0.023105f
C8246 PAD.n9445 VSS 0.547498f
C8247 PAD.n9446 VSS 0.453782f
C8248 PAD.n9447 VSS 0.025763f
C8249 PAD.n9448 VSS 0.025763f
C8250 PAD.n9449 VSS 0.022501f
C8251 PAD.n9450 VSS 0.033766f
C8252 PAD.n9451 VSS 0.04183f
C8253 PAD.n9452 VSS 0.040018f
C8254 PAD.n9453 VSS 0.045821f
C8255 PAD.n9454 VSS 0.045821f
C8256 PAD.n9455 VSS 0.503106f
C8257 PAD.n9456 VSS 0.700403f
C8258 PAD.n9457 VSS 0.069752f
C8259 PAD.n9458 VSS 0.048377f
C8260 PAD.n9459 VSS 0.039754f
C8261 PAD.n9460 VSS 0.056252f
C8262 PAD.n9461 VSS 0.056252f
C8263 PAD.n9462 VSS 0.039754f
C8264 PAD.n9463 VSS 0.023105f
C8265 PAD.n9464 VSS 0.033374f
C8266 PAD.n9465 VSS 0.036454f
C8267 PAD.n9466 VSS 0.036454f
C8268 PAD.n9467 VSS 0.036454f
C8269 PAD.n9468 VSS 0.036454f
C8270 PAD.n9470 VSS 0.036454f
C8271 PAD.n9471 VSS 0.036454f
C8272 PAD.n9472 VSS 0.036454f
C8273 PAD.n9474 VSS 0.036454f
C8274 PAD.n9475 VSS 0.036454f
C8275 PAD.n9476 VSS 0.036454f
C8276 PAD.n9477 VSS 0.036454f
C8277 PAD.n9478 VSS 0.036454f
C8278 PAD.n9479 VSS 0.036454f
C8279 PAD.n9480 VSS 0.036454f
C8280 PAD.n9482 VSS 0.036454f
C8281 PAD.n9483 VSS 0.036454f
C8282 PAD.n9484 VSS 0.036454f
C8283 PAD.n9486 VSS 0.036454f
C8284 PAD.n9487 VSS 0.036454f
C8285 PAD.n9488 VSS 0.036454f
C8286 PAD.n9489 VSS 0.036454f
C8287 PAD.n9490 VSS 0.036454f
C8288 PAD.n9491 VSS 0.036454f
C8289 PAD.n9492 VSS 0.036454f
C8290 PAD.n9494 VSS 0.036454f
C8291 PAD.n9495 VSS 0.036454f
C8292 PAD.n9496 VSS 0.036454f
C8293 PAD.n9498 VSS 0.036454f
C8294 PAD.n9499 VSS 0.036454f
C8295 PAD.n9500 VSS 0.036454f
C8296 PAD.n9501 VSS 0.036454f
C8297 PAD.n9502 VSS 0.036454f
C8298 PAD.n9503 VSS 0.036454f
C8299 PAD.n9504 VSS 0.036454f
C8300 PAD.n9506 VSS 0.036454f
C8301 PAD.n9507 VSS 0.036454f
C8302 PAD.n9508 VSS 0.036454f
C8303 PAD.n9510 VSS 0.036454f
C8304 PAD.n9511 VSS 0.036454f
C8305 PAD.n9512 VSS 0.036454f
C8306 PAD.n9513 VSS 0.036454f
C8307 PAD.n9514 VSS 0.036454f
C8308 PAD.n9515 VSS 0.036454f
C8309 PAD.n9516 VSS 0.036454f
C8310 PAD.n9518 VSS 0.036454f
C8311 PAD.n9519 VSS 0.036454f
C8312 PAD.n9520 VSS 0.036454f
C8313 PAD.n9522 VSS 0.036454f
C8314 PAD.n9523 VSS 0.036454f
C8315 PAD.n9524 VSS 0.036454f
C8316 PAD.n9525 VSS 0.036454f
C8317 PAD.n9526 VSS 0.036454f
C8318 PAD.n9527 VSS 0.036454f
C8319 PAD.n9528 VSS 0.036454f
C8320 PAD.n9530 VSS 0.036454f
C8321 PAD.n9531 VSS 0.036454f
C8322 PAD.n9532 VSS 0.036454f
C8323 PAD.n9534 VSS 0.036454f
C8324 PAD.n9535 VSS 0.036454f
C8325 PAD.n9536 VSS 0.036454f
C8326 PAD.n9537 VSS 0.036454f
C8327 PAD.n9538 VSS 0.036454f
C8328 PAD.n9539 VSS 0.036454f
C8329 PAD.n9540 VSS 0.036454f
C8330 PAD.n9542 VSS 0.036454f
C8331 PAD.n9543 VSS 0.036454f
C8332 PAD.n9544 VSS 0.036454f
C8333 PAD.n9546 VSS 0.036454f
C8334 PAD.n9547 VSS 0.036454f
C8335 PAD.n9548 VSS 0.036454f
C8336 PAD.n9549 VSS 0.036454f
C8337 PAD.n9550 VSS 0.036454f
C8338 PAD.n9551 VSS 0.036454f
C8339 PAD.n9552 VSS 0.036454f
C8340 PAD.n9554 VSS 0.036454f
C8341 PAD.n9555 VSS 0.036454f
C8342 PAD.n9556 VSS 0.036454f
C8343 PAD.n9558 VSS 0.036454f
C8344 PAD.n9559 VSS 0.036454f
C8345 PAD.n9560 VSS 0.036454f
C8346 PAD.n9561 VSS 0.036454f
C8347 PAD.n9562 VSS 0.036454f
C8348 PAD.n9563 VSS 0.036454f
C8349 PAD.n9564 VSS 0.036454f
C8350 PAD.n9566 VSS 0.036454f
C8351 PAD.n9567 VSS 0.036454f
C8352 PAD.n9568 VSS 0.036454f
C8353 PAD.n9570 VSS 0.036454f
C8354 PAD.n9571 VSS 0.036454f
C8355 PAD.n9572 VSS 0.036454f
C8356 PAD.n9573 VSS 0.036454f
C8357 PAD.n9574 VSS 0.036454f
C8358 PAD.n9575 VSS 0.036454f
C8359 PAD.n9576 VSS 0.036454f
C8360 PAD.n9578 VSS 0.036454f
C8361 PAD.n9579 VSS 0.036454f
C8362 PAD.n9580 VSS 0.036454f
C8363 PAD.n9582 VSS 0.036454f
C8364 PAD.n9583 VSS 0.036454f
C8365 PAD.n9584 VSS 0.036454f
C8366 PAD.n9585 VSS 0.036454f
C8367 PAD.n9586 VSS 0.036454f
C8368 PAD.n9587 VSS 0.036454f
C8369 PAD.n9588 VSS 0.036454f
C8370 PAD.n9590 VSS 0.036454f
C8371 PAD.n9591 VSS 0.036454f
C8372 PAD.n9592 VSS 0.036454f
C8373 PAD.n9594 VSS 0.036454f
C8374 PAD.n9595 VSS 0.036454f
C8375 PAD.n9596 VSS 0.036454f
C8376 PAD.n9597 VSS 0.036454f
C8377 PAD.n9598 VSS 0.036454f
C8378 PAD.n9599 VSS 0.036454f
C8379 PAD.n9600 VSS 0.036454f
C8380 PAD.n9602 VSS 0.036454f
C8381 PAD.n9603 VSS 0.036454f
C8382 PAD.n9604 VSS 0.036454f
C8383 PAD.n9606 VSS 0.036454f
C8384 PAD.n9607 VSS 0.036454f
C8385 PAD.n9608 VSS 0.036454f
C8386 PAD.n9609 VSS 0.036454f
C8387 PAD.n9610 VSS 0.036454f
C8388 PAD.n9611 VSS 0.036454f
C8389 PAD.n9612 VSS 0.036454f
C8390 PAD.n9614 VSS 0.036454f
C8391 PAD.n9615 VSS 0.036454f
C8392 PAD.n9616 VSS 0.036454f
C8393 PAD.n9618 VSS 0.036454f
C8394 PAD.n9619 VSS 0.036454f
C8395 PAD.n9620 VSS 0.036454f
C8396 PAD.n9621 VSS 0.036454f
C8397 PAD.n9622 VSS 0.036454f
C8398 PAD.n9623 VSS 0.036454f
C8399 PAD.n9624 VSS 0.036454f
C8400 PAD.n9626 VSS 0.036454f
C8401 PAD.n9627 VSS 0.036454f
C8402 PAD.n9628 VSS 0.036454f
C8403 PAD.n9630 VSS 0.036454f
C8404 PAD.n9631 VSS 0.036454f
C8405 PAD.n9632 VSS 0.036454f
C8406 PAD.n9633 VSS 0.036454f
C8407 PAD.n9634 VSS 0.036454f
C8408 PAD.n9635 VSS 0.036454f
C8409 PAD.n9636 VSS 0.036454f
C8410 PAD.n9638 VSS 0.036454f
C8411 PAD.n9639 VSS 0.036454f
C8412 PAD.n9640 VSS 0.036454f
C8413 PAD.n9642 VSS 0.036454f
C8414 PAD.n9643 VSS 0.036454f
C8415 PAD.n9644 VSS 0.036454f
C8416 PAD.n9645 VSS 0.036454f
C8417 PAD.n9646 VSS 0.036454f
C8418 PAD.n9647 VSS 0.036454f
C8419 PAD.n9648 VSS 0.036454f
C8420 PAD.n9650 VSS 0.036454f
C8421 PAD.n9651 VSS 0.036454f
C8422 PAD.n9652 VSS 0.036454f
C8423 PAD.n9654 VSS 0.036454f
C8424 PAD.n9655 VSS 0.036454f
C8425 PAD.n9656 VSS 0.036454f
C8426 PAD.n9657 VSS 0.036454f
C8427 PAD.n9658 VSS 0.036454f
C8428 PAD.n9659 VSS 0.036454f
C8429 PAD.n9660 VSS 0.036454f
C8430 PAD.n9662 VSS 0.036454f
C8431 PAD.n9663 VSS 0.036454f
C8432 PAD.n9664 VSS 0.036454f
C8433 PAD.n9666 VSS 0.036454f
C8434 PAD.n9667 VSS 0.036454f
C8435 PAD.n9668 VSS 0.036454f
C8436 PAD.n9669 VSS 0.036454f
C8437 PAD.n9670 VSS 0.036454f
C8438 PAD.n9671 VSS 0.036454f
C8439 PAD.n9672 VSS 0.036454f
C8440 PAD.n9674 VSS 0.036454f
C8441 PAD.n9675 VSS 0.036454f
C8442 PAD.n9676 VSS 0.036454f
C8443 PAD.n9678 VSS 0.036454f
C8444 PAD.n9679 VSS 0.036454f
C8445 PAD.n9680 VSS 0.036454f
C8446 PAD.n9681 VSS 0.036454f
C8447 PAD.n9682 VSS 0.036454f
C8448 PAD.n9683 VSS 0.036454f
C8449 PAD.n9684 VSS 0.036454f
C8450 PAD.n9686 VSS 0.036454f
C8451 PAD.n9687 VSS 0.036454f
C8452 PAD.n9688 VSS 0.036454f
C8453 PAD.n9690 VSS 0.036454f
C8454 PAD.n9691 VSS 0.036454f
C8455 PAD.n9692 VSS 0.036454f
C8456 PAD.n9693 VSS 0.036454f
C8457 PAD.n9694 VSS 0.036454f
C8458 PAD.n9695 VSS 0.036454f
C8459 PAD.n9696 VSS 0.036454f
C8460 PAD.n9698 VSS 0.036454f
C8461 PAD.n9699 VSS 0.036454f
C8462 PAD.n9700 VSS 0.036454f
C8463 PAD.n9702 VSS 0.036454f
C8464 PAD.n9703 VSS 0.036454f
C8465 PAD.n9704 VSS 0.036454f
C8466 PAD.n9705 VSS 0.036454f
C8467 PAD.n9706 VSS 0.03055f
C8468 PAD.n9707 VSS 0.036454f
C8469 PAD.n9708 VSS 0.036454f
C8470 PAD.n9709 VSS 0.036454f
C8471 PAD.n9711 VSS 0.023105f
C8472 PAD.n9712 VSS 0.281147f
C8473 PAD.n9713 VSS 0.591889f
C8474 PAD.n9714 VSS 0.027838f
C8475 PAD.n9715 VSS 0.027838f
C8476 PAD.n9716 VSS 0.024313f
C8477 PAD.n9717 VSS 0.042887f
C8478 PAD.n9718 VSS 0.036092f
C8479 PAD.n9719 VSS 0.041325f
C8480 PAD.n9720 VSS 0.041325f
C8481 PAD.n9721 VSS 0.611619f
C8482 PAD.n9722 VSS 0.157837f
C8483 PAD.n9723 VSS 0.056252f
C8484 PAD.n9724 VSS 0.056252f
C8485 PAD.n9725 VSS 0.050211f
C8486 PAD.n9726 VSS 0.046278f
C8487 PAD.n9727 VSS 0.057241f
C8488 PAD.n9728 VSS 0.062262f
C8489 PAD.n9729 VSS 0.043182f
C8490 PAD.n9730 VSS 0.048377f
C8491 PAD.n9731 VSS 0.048377f
C8492 PAD.n9732 VSS 0.157837f
C8493 PAD.n9733 VSS 0.557363f
C8494 PAD.n9734 VSS 0.032334f
C8495 PAD.n9735 VSS 0.032334f
C8496 PAD.n9736 VSS 0.028239f
C8497 PAD.n9737 VSS 0.042887f
C8498 PAD.n9738 VSS 0.032166f
C8499 PAD.n9739 VSS 0.036829f
C8500 PAD.n9740 VSS 0.036829f
C8501 PAD.n9741 VSS 0.177566f
C8502 PAD.n9742 VSS 0.700403f
C8503 PAD.n9743 VSS 0.064127f
C8504 PAD.n9744 VSS 0.039754f
C8505 PAD.n9745 VSS 0.069752f
C8506 PAD.n9746 VSS 0.040501f
C8507 PAD.n9747 VSS 0.040501f
C8508 PAD.n9748 VSS 0.039754f
C8509 PAD.n9749 VSS 0.023105f
C8510 PAD.n9750 VSS 0.033374f
C8511 PAD.n9751 VSS 0.036454f
C8512 PAD.n9752 VSS 0.036454f
C8513 PAD.n9753 VSS 0.036454f
C8514 PAD.n9754 VSS 0.036454f
C8515 PAD.n9756 VSS 0.036454f
C8516 PAD.n9757 VSS 0.036454f
C8517 PAD.n9758 VSS 0.036454f
C8518 PAD.n9760 VSS 0.036454f
C8519 PAD.n9761 VSS 0.036454f
C8520 PAD.n9762 VSS 0.036454f
C8521 PAD.n9763 VSS 0.036454f
C8522 PAD.n9764 VSS 0.036454f
C8523 PAD.n9765 VSS 0.036454f
C8524 PAD.n9766 VSS 0.036454f
C8525 PAD.n9768 VSS 0.036454f
C8526 PAD.n9769 VSS 0.036454f
C8527 PAD.n9770 VSS 0.036454f
C8528 PAD.n9772 VSS 0.036454f
C8529 PAD.n9773 VSS 0.036454f
C8530 PAD.n9774 VSS 0.036454f
C8531 PAD.n9775 VSS 0.036454f
C8532 PAD.n9776 VSS 0.036454f
C8533 PAD.n9777 VSS 0.036454f
C8534 PAD.n9778 VSS 0.036454f
C8535 PAD.n9780 VSS 0.036454f
C8536 PAD.n9781 VSS 0.036454f
C8537 PAD.n9782 VSS 0.036454f
C8538 PAD.n9784 VSS 0.036454f
C8539 PAD.n9785 VSS 0.036454f
C8540 PAD.n9786 VSS 0.036454f
C8541 PAD.n9787 VSS 0.036454f
C8542 PAD.n9788 VSS 0.036454f
C8543 PAD.n9789 VSS 0.036454f
C8544 PAD.n9790 VSS 0.036454f
C8545 PAD.n9792 VSS 0.036454f
C8546 PAD.n9793 VSS 0.036454f
C8547 PAD.n9794 VSS 0.036454f
C8548 PAD.n9796 VSS 0.036454f
C8549 PAD.n9797 VSS 0.036454f
C8550 PAD.n9798 VSS 0.036454f
C8551 PAD.n9799 VSS 0.036454f
C8552 PAD.n9800 VSS 0.036454f
C8553 PAD.n9801 VSS 0.036454f
C8554 PAD.n9802 VSS 0.036454f
C8555 PAD.n9804 VSS 0.036454f
C8556 PAD.n9805 VSS 0.036454f
C8557 PAD.n9806 VSS 0.036454f
C8558 PAD.n9808 VSS 0.036454f
C8559 PAD.n9809 VSS 0.036454f
C8560 PAD.n9810 VSS 0.036454f
C8561 PAD.n9811 VSS 0.036454f
C8562 PAD.n9812 VSS 0.036454f
C8563 PAD.n9813 VSS 0.036454f
C8564 PAD.n9814 VSS 0.036454f
C8565 PAD.n9816 VSS 0.036454f
C8566 PAD.n9817 VSS 0.036454f
C8567 PAD.n9818 VSS 0.036454f
C8568 PAD.n9820 VSS 0.036454f
C8569 PAD.n9821 VSS 0.036454f
C8570 PAD.n9822 VSS 0.036454f
C8571 PAD.n9823 VSS 0.036454f
C8572 PAD.n9824 VSS 0.036454f
C8573 PAD.n9825 VSS 0.036454f
C8574 PAD.n9826 VSS 0.036454f
C8575 PAD.n9828 VSS 0.036454f
C8576 PAD.n9829 VSS 0.036454f
C8577 PAD.n9830 VSS 0.036454f
C8578 PAD.n9832 VSS 0.036454f
C8579 PAD.n9833 VSS 0.036454f
C8580 PAD.n9834 VSS 0.036454f
C8581 PAD.n9835 VSS 0.036454f
C8582 PAD.n9836 VSS 0.036454f
C8583 PAD.n9837 VSS 0.036454f
C8584 PAD.n9838 VSS 0.036454f
C8585 PAD.n9840 VSS 0.036454f
C8586 PAD.n9841 VSS 0.036454f
C8587 PAD.n9842 VSS 0.036454f
C8588 PAD.n9844 VSS 0.036454f
C8589 PAD.n9845 VSS 0.036454f
C8590 PAD.n9846 VSS 0.036454f
C8591 PAD.n9847 VSS 0.036454f
C8592 PAD.n9848 VSS 0.036454f
C8593 PAD.n9849 VSS 0.036454f
C8594 PAD.n9850 VSS 0.036454f
C8595 PAD.n9852 VSS 0.036454f
C8596 PAD.n9853 VSS 0.036454f
C8597 PAD.n9854 VSS 0.036454f
C8598 PAD.n9856 VSS 0.036454f
C8599 PAD.n9857 VSS 0.036454f
C8600 PAD.n9858 VSS 0.036454f
C8601 PAD.n9859 VSS 0.036454f
C8602 PAD.n9860 VSS 0.036454f
C8603 PAD.n9861 VSS 0.036454f
C8604 PAD.n9862 VSS 0.036454f
C8605 PAD.n9864 VSS 0.036454f
C8606 PAD.n9865 VSS 0.036454f
C8607 PAD.n9866 VSS 0.036454f
C8608 PAD.n9868 VSS 0.036454f
C8609 PAD.n9869 VSS 0.036454f
C8610 PAD.n9870 VSS 0.036454f
C8611 PAD.n9871 VSS 0.036454f
C8612 PAD.n9872 VSS 0.036454f
C8613 PAD.n9873 VSS 0.036454f
C8614 PAD.n9874 VSS 0.036454f
C8615 PAD.n9876 VSS 0.036454f
C8616 PAD.n9877 VSS 0.036454f
C8617 PAD.n9878 VSS 0.036454f
C8618 PAD.n9880 VSS 0.036454f
C8619 PAD.n9881 VSS 0.036454f
C8620 PAD.n9882 VSS 0.036454f
C8621 PAD.n9883 VSS 0.036454f
C8622 PAD.n9884 VSS 0.036454f
C8623 PAD.n9885 VSS 0.036454f
C8624 PAD.n9886 VSS 0.036454f
C8625 PAD.n9888 VSS 0.036454f
C8626 PAD.n9889 VSS 0.036454f
C8627 PAD.n9890 VSS 0.036454f
C8628 PAD.n9892 VSS 0.036454f
C8629 PAD.n9893 VSS 0.036454f
C8630 PAD.n9894 VSS 0.036454f
C8631 PAD.n9895 VSS 0.036454f
C8632 PAD.n9896 VSS 0.036454f
C8633 PAD.n9897 VSS 0.036454f
C8634 PAD.n9898 VSS 0.036454f
C8635 PAD.n9900 VSS 0.036454f
C8636 PAD.n9901 VSS 0.036454f
C8637 PAD.n9902 VSS 0.036454f
C8638 PAD.n9904 VSS 0.036454f
C8639 PAD.n9905 VSS 0.036454f
C8640 PAD.n9906 VSS 0.036454f
C8641 PAD.n9907 VSS 0.036454f
C8642 PAD.n9908 VSS 0.036454f
C8643 PAD.n9909 VSS 0.036454f
C8644 PAD.n9910 VSS 0.036454f
C8645 PAD.n9912 VSS 0.036454f
C8646 PAD.n9913 VSS 0.036454f
C8647 PAD.n9914 VSS 0.036454f
C8648 PAD.n9916 VSS 0.036454f
C8649 PAD.n9917 VSS 0.036454f
C8650 PAD.n9918 VSS 0.036454f
C8651 PAD.n9919 VSS 0.036454f
C8652 PAD.n9920 VSS 0.036454f
C8653 PAD.n9921 VSS 0.036454f
C8654 PAD.n9922 VSS 0.036454f
C8655 PAD.n9924 VSS 0.036454f
C8656 PAD.n9925 VSS 0.036454f
C8657 PAD.n9926 VSS 0.036454f
C8658 PAD.n9928 VSS 0.036454f
C8659 PAD.n9929 VSS 0.036454f
C8660 PAD.n9930 VSS 0.036454f
C8661 PAD.n9931 VSS 0.036454f
C8662 PAD.n9932 VSS 0.036454f
C8663 PAD.n9933 VSS 0.036454f
C8664 PAD.n9934 VSS 0.036454f
C8665 PAD.n9936 VSS 0.036454f
C8666 PAD.n9937 VSS 0.036454f
C8667 PAD.n9938 VSS 0.036454f
C8668 PAD.n9940 VSS 0.036454f
C8669 PAD.n9941 VSS 0.036454f
C8670 PAD.n9942 VSS 0.036454f
C8671 PAD.n9943 VSS 0.036454f
C8672 PAD.n9944 VSS 0.036454f
C8673 PAD.n9945 VSS 0.036454f
C8674 PAD.n9946 VSS 0.036454f
C8675 PAD.n9948 VSS 0.036454f
C8676 PAD.n9949 VSS 0.036454f
C8677 PAD.n9950 VSS 0.036454f
C8678 PAD.n9952 VSS 0.036454f
C8679 PAD.n9953 VSS 0.036454f
C8680 PAD.n9954 VSS 0.036454f
C8681 PAD.n9955 VSS 0.036454f
C8682 PAD.n9956 VSS 0.036454f
C8683 PAD.n9957 VSS 0.036454f
C8684 PAD.n9958 VSS 0.036454f
C8685 PAD.n9960 VSS 0.036454f
C8686 PAD.n9961 VSS 0.036454f
C8687 PAD.n9962 VSS 0.036454f
C8688 PAD.n9964 VSS 0.036454f
C8689 PAD.n9965 VSS 0.036454f
C8690 PAD.n9966 VSS 0.036454f
C8691 PAD.n9967 VSS 0.036454f
C8692 PAD.n9968 VSS 0.036454f
C8693 PAD.n9969 VSS 0.036454f
C8694 PAD.n9970 VSS 0.036454f
C8695 PAD.n9972 VSS 0.036454f
C8696 PAD.n9973 VSS 0.036454f
C8697 PAD.n9974 VSS 0.036454f
C8698 PAD.n9976 VSS 0.036454f
C8699 PAD.n9977 VSS 0.036454f
C8700 PAD.n9978 VSS 0.036454f
C8701 PAD.n9979 VSS 0.036454f
C8702 PAD.n9980 VSS 0.036454f
C8703 PAD.n9981 VSS 0.036454f
C8704 PAD.n9982 VSS 0.036454f
C8705 PAD.n9984 VSS 0.036454f
C8706 PAD.n9985 VSS 0.036454f
C8707 PAD.n9986 VSS 0.036454f
C8708 PAD.n9988 VSS 0.036454f
C8709 PAD.n9989 VSS 0.036454f
C8710 PAD.n9990 VSS 0.036454f
C8711 PAD.n9991 VSS 0.036454f
C8712 PAD.n9992 VSS 0.03055f
C8713 PAD.n9993 VSS 0.036454f
C8714 PAD.n9994 VSS 0.036454f
C8715 PAD.n9995 VSS 0.036454f
C8716 PAD.n9997 VSS 0.023105f
C8717 PAD.n9998 VSS 0.360066f
C8718 PAD.n9999 VSS 0.26635f
C8719 PAD.n10000 VSS 0.036829f
C8720 PAD.n10001 VSS 0.036829f
C8721 PAD.n10002 VSS 0.032166f
C8722 PAD.n10003 VSS 0.042887f
C8723 PAD.n10004 VSS 0.028239f
C8724 PAD.n10005 VSS 0.032334f
C8725 PAD.n10006 VSS 0.032334f
C8726 PAD.n10007 VSS 0.295944f
C8727 PAD.n10008 VSS 0.586957f
C8728 PAD.n10009 VSS 0.037126f
C8729 PAD.n10010 VSS 0.037126f
C8730 PAD.n10011 VSS 0.03314f
C8731 PAD.n10012 VSS 0.046278f
C8732 PAD.n10013 VSS 0.060254f
C8733 PAD.n10014 VSS 0.067502f
C8734 PAD.n10015 VSS 0.067502f
C8735 PAD.n10016 VSS 0.700403f
C8736 PAD.n10017 VSS 0.207161f
C8737 PAD.n10018 VSS 0.041325f
C8738 PAD.n10019 VSS 0.041325f
C8739 PAD.n10020 VSS 0.036092f
C8740 PAD.n10021 VSS 0.042887f
C8741 PAD.n10022 VSS 0.036454f
C8742 PAD.n10023 VSS 0.036454f
C8743 PAD.n10024 VSS 0.036454f
C8744 PAD.n10026 VSS 0.036454f
C8745 PAD.n10027 VSS 0.036454f
C8746 PAD.n10028 VSS 0.036454f
C8747 PAD.n10030 VSS 0.036454f
C8748 PAD.n10031 VSS 0.036454f
C8749 PAD.n10032 VSS 0.036454f
C8750 PAD.n10034 VSS 0.036454f
C8751 PAD.n10035 VSS 0.036454f
C8752 PAD.n10036 VSS 0.036454f
C8753 PAD.n10038 VSS 0.036454f
C8754 PAD.n10039 VSS 0.036454f
C8755 PAD.n10040 VSS 0.036454f
C8756 PAD.n10042 VSS 0.036454f
C8757 PAD.n10043 VSS 0.036454f
C8758 PAD.n10044 VSS 0.036454f
C8759 PAD.n10046 VSS 0.036454f
C8760 PAD.n10047 VSS 0.036454f
C8761 PAD.n10048 VSS 0.036454f
C8762 PAD.n10050 VSS 0.036454f
C8763 PAD.n10051 VSS 0.036454f
C8764 PAD.n10052 VSS 0.036454f
C8765 PAD.n10054 VSS 0.036454f
C8766 PAD.n10055 VSS 0.036454f
C8767 PAD.n10056 VSS 0.036454f
C8768 PAD.n10058 VSS 0.036454f
C8769 PAD.n10059 VSS 0.036454f
C8770 PAD.n10060 VSS 0.036454f
C8771 PAD.n10062 VSS 0.036454f
C8772 PAD.n10063 VSS 0.036454f
C8773 PAD.n10064 VSS 0.036454f
C8774 PAD.n10066 VSS 0.036454f
C8775 PAD.n10067 VSS 0.036454f
C8776 PAD.n10068 VSS 0.036454f
C8777 PAD.n10070 VSS 0.036454f
C8778 PAD.n10071 VSS 0.036454f
C8779 PAD.n10072 VSS 0.036454f
C8780 PAD.n10074 VSS 0.036454f
C8781 PAD.n10075 VSS 0.036454f
C8782 PAD.n10076 VSS 0.036454f
C8783 PAD.n10078 VSS 0.036454f
C8784 PAD.n10079 VSS 0.036454f
C8785 PAD.n10080 VSS 0.036454f
C8786 PAD.n10082 VSS 0.036454f
C8787 PAD.n10083 VSS 0.036454f
C8788 PAD.n10084 VSS 0.036454f
C8789 PAD.n10086 VSS 0.036454f
C8790 PAD.n10087 VSS 0.036454f
C8791 PAD.n10088 VSS 0.036454f
C8792 PAD.n10090 VSS 0.036454f
C8793 PAD.n10091 VSS 0.036454f
C8794 PAD.n10092 VSS 0.036454f
C8795 PAD.n10094 VSS 0.036454f
C8796 PAD.n10095 VSS 0.036454f
C8797 PAD.n10096 VSS 0.036454f
C8798 PAD.n10098 VSS 0.036454f
C8799 PAD.n10099 VSS 0.036454f
C8800 PAD.n10100 VSS 0.036454f
C8801 PAD.n10102 VSS 0.036454f
C8802 PAD.n10103 VSS 0.036454f
C8803 PAD.n10104 VSS 0.036454f
C8804 PAD.n10105 VSS 0.023105f
C8805 PAD.n10106 VSS 0.023105f
C8806 PAD.n10108 VSS 0.036454f
C8807 PAD.n10110 VSS 0.036454f
C8808 PAD.n10112 VSS 0.036454f
C8809 PAD.n10113 VSS 0.036454f
C8810 PAD.n10114 VSS 0.036454f
C8811 PAD.n10115 VSS 0.036454f
C8812 PAD.n10116 VSS 0.036454f
C8813 PAD.n10117 VSS 0.036454f
C8814 PAD.n10118 VSS 0.036454f
C8815 PAD.n10120 VSS 0.036454f
C8816 PAD.n10122 VSS 0.036454f
C8817 PAD.n10124 VSS 0.036454f
C8818 PAD.n10125 VSS 0.036454f
C8819 PAD.n10126 VSS 0.036454f
C8820 PAD.n10127 VSS 0.036454f
C8821 PAD.n10128 VSS 0.036454f
C8822 PAD.n10129 VSS 0.036454f
C8823 PAD.n10130 VSS 0.036454f
C8824 PAD.n10132 VSS 0.036454f
C8825 PAD.n10134 VSS 0.036454f
C8826 PAD.n10136 VSS 0.036454f
C8827 PAD.n10137 VSS 0.036454f
C8828 PAD.n10138 VSS 0.036454f
C8829 PAD.n10139 VSS 0.036454f
C8830 PAD.n10140 VSS 0.036454f
C8831 PAD.n10141 VSS 0.036454f
C8832 PAD.n10142 VSS 0.036454f
C8833 PAD.n10144 VSS 0.036454f
C8834 PAD.n10146 VSS 0.036454f
C8835 PAD.n10148 VSS 0.036454f
C8836 PAD.n10149 VSS 0.036454f
C8837 PAD.n10150 VSS 0.036454f
C8838 PAD.n10151 VSS 0.036454f
C8839 PAD.n10152 VSS 0.036454f
C8840 PAD.n10153 VSS 0.036454f
C8841 PAD.n10154 VSS 0.036454f
C8842 PAD.n10156 VSS 0.036454f
C8843 PAD.n10158 VSS 0.036454f
C8844 PAD.n10160 VSS 0.036454f
C8845 PAD.n10161 VSS 0.036454f
C8846 PAD.n10162 VSS 0.036454f
C8847 PAD.n10163 VSS 0.036454f
C8848 PAD.n10164 VSS 0.036454f
C8849 PAD.n10165 VSS 0.036454f
C8850 PAD.n10166 VSS 0.036454f
C8851 PAD.n10168 VSS 0.036454f
C8852 PAD.n10170 VSS 0.036454f
C8853 PAD.n10172 VSS 0.036454f
C8854 PAD.n10173 VSS 0.036454f
C8855 PAD.n10174 VSS 0.036454f
C8856 PAD.n10175 VSS 0.036454f
C8857 PAD.n10176 VSS 0.036454f
C8858 PAD.n10177 VSS 0.036454f
C8859 PAD.n10178 VSS 0.036454f
C8860 PAD.n10180 VSS 0.036454f
C8861 PAD.n10182 VSS 0.036454f
C8862 PAD.n10184 VSS 0.036454f
C8863 PAD.n10185 VSS 0.036454f
C8864 PAD.n10186 VSS 0.036454f
C8865 PAD.n10187 VSS 0.036454f
C8866 PAD.n10188 VSS 0.036454f
C8867 PAD.n10189 VSS 0.036454f
C8868 PAD.n10190 VSS 0.036454f
C8869 PAD.n10192 VSS 0.036454f
C8870 PAD.n10194 VSS 0.036454f
C8871 PAD.n10196 VSS 0.036454f
C8872 PAD.n10197 VSS 0.036454f
C8873 PAD.n10198 VSS 0.036454f
C8874 PAD.n10199 VSS 0.036454f
C8875 PAD.n10200 VSS 0.036454f
C8876 PAD.n10201 VSS 0.036454f
C8877 PAD.n10202 VSS 0.036454f
C8878 PAD.n10204 VSS 0.036454f
C8879 PAD.n10206 VSS 0.036454f
C8880 PAD.n10208 VSS 0.036454f
C8881 PAD.n10209 VSS 0.036454f
C8882 PAD.n10210 VSS 0.036454f
C8883 PAD.n10211 VSS 0.036454f
C8884 PAD.n10212 VSS 0.036454f
C8885 PAD.n10213 VSS 0.036454f
C8886 PAD.n10214 VSS 0.036454f
C8887 PAD.n10216 VSS 0.036454f
C8888 PAD.n10218 VSS 0.036454f
C8889 PAD.n10220 VSS 0.036454f
C8890 PAD.n10221 VSS 0.036454f
C8891 PAD.n10222 VSS 0.036454f
C8892 PAD.n10223 VSS 0.036454f
C8893 PAD.n10224 VSS 0.036454f
C8894 PAD.n10225 VSS 0.036454f
C8895 PAD.n10226 VSS 0.036454f
C8896 PAD.n10228 VSS 0.036454f
C8897 PAD.n10230 VSS 0.036454f
C8898 PAD.n10232 VSS 0.036454f
C8899 PAD.n10233 VSS 0.036454f
C8900 PAD.n10234 VSS 0.036454f
C8901 PAD.n10235 VSS 0.036454f
C8902 PAD.n10236 VSS 0.036454f
C8903 PAD.n10237 VSS 0.036454f
C8904 PAD.n10238 VSS 0.036454f
C8905 PAD.n10240 VSS 0.036454f
C8906 PAD.n10242 VSS 0.036454f
C8907 PAD.n10244 VSS 0.036454f
C8908 PAD.n10245 VSS 0.036454f
C8909 PAD.n10246 VSS 0.036454f
C8910 PAD.n10247 VSS 0.036454f
C8911 PAD.n10248 VSS 0.036454f
C8912 PAD.n10249 VSS 0.036454f
C8913 PAD.n10250 VSS 0.036454f
C8914 PAD.n10252 VSS 0.036454f
C8915 PAD.n10254 VSS 0.036454f
C8916 PAD.n10256 VSS 0.036454f
C8917 PAD.n10257 VSS 0.036454f
C8918 PAD.n10258 VSS 0.036454f
C8919 PAD.n10259 VSS 0.036454f
C8920 PAD.n10260 VSS 0.036454f
C8921 PAD.n10261 VSS 0.036454f
C8922 PAD.n10262 VSS 0.036454f
C8923 PAD.n10264 VSS 0.036454f
C8924 PAD.n10266 VSS 0.036454f
C8925 PAD.n10268 VSS 0.036454f
C8926 PAD.n10269 VSS 0.036454f
C8927 PAD.n10270 VSS 0.036454f
C8928 PAD.n10271 VSS 0.036454f
C8929 PAD.n10272 VSS 0.036454f
C8930 PAD.n10273 VSS 0.036454f
C8931 PAD.n10274 VSS 0.036454f
C8932 PAD.n10276 VSS 0.036454f
C8933 PAD.n10278 VSS 0.036454f
C8934 PAD.n10280 VSS 0.036454f
C8935 PAD.n10281 VSS 0.036454f
C8936 PAD.n10282 VSS 0.036454f
C8937 PAD.n10283 VSS 0.036454f
C8938 PAD.n10284 VSS 0.036454f
C8939 PAD.n10285 VSS 0.036454f
C8940 PAD.n10286 VSS 0.036454f
C8941 PAD.n10288 VSS 0.036454f
C8942 PAD.n10290 VSS 0.036454f
C8943 PAD.n10292 VSS 0.036454f
C8944 PAD.n10293 VSS 0.036454f
C8945 PAD.n10294 VSS 0.036454f
C8946 PAD.n10295 VSS 0.036454f
C8947 PAD.n10296 VSS 0.036454f
C8948 PAD.n10297 VSS 0.036454f
C8949 PAD.n10298 VSS 0.036454f
C8950 PAD.n10300 VSS 0.036454f
C8951 PAD.n10302 VSS 0.036454f
C8952 PAD.n10304 VSS 0.036454f
C8953 PAD.n10305 VSS 0.036454f
C8954 PAD.n10306 VSS 0.036454f
C8955 PAD.n10307 VSS 0.036454f
C8956 PAD.n10308 VSS 0.036454f
C8957 PAD.n10309 VSS 0.036454f
C8958 PAD.n10310 VSS 0.036454f
C8959 PAD.n10312 VSS 0.036454f
C8960 PAD.n10314 VSS 0.036454f
C8961 PAD.n10316 VSS 0.036454f
C8962 PAD.n10317 VSS 0.036454f
C8963 PAD.n10318 VSS 0.036454f
C8964 PAD.n10319 VSS 0.036454f
C8965 PAD.n10320 VSS 0.036454f
C8966 PAD.n10321 VSS 0.036454f
C8967 PAD.n10322 VSS 0.036454f
C8968 PAD.n10324 VSS 0.036454f
C8969 PAD.n10326 VSS 0.036454f
C8970 PAD.n10328 VSS 0.036454f
C8971 PAD.n10329 VSS 0.036454f
C8972 PAD.n10330 VSS 0.036454f
C8973 PAD.n10331 VSS 0.036454f
C8974 PAD.n10332 VSS 0.036454f
C8975 PAD.n10333 VSS 0.036454f
C8976 PAD.n10334 VSS 0.036454f
C8977 PAD.n10336 VSS 0.036454f
C8978 PAD.n10338 VSS 0.036454f
C8979 PAD.n10340 VSS 0.036454f
C8980 PAD.n10341 VSS 0.036454f
C8981 PAD.n10342 VSS 0.036454f
C8982 PAD.n10343 VSS 0.036454f
C8983 PAD.n10344 VSS 0.036454f
C8984 PAD.n10345 VSS 0.036454f
C8985 PAD.n10346 VSS 0.036454f
C8986 PAD.n10347 VSS 0.036454f
C8987 PAD.n10349 VSS 0.036454f
C8988 PAD.n10351 VSS 0.036454f
C8989 PAD.n10353 VSS 0.023105f
C8990 PAD.n10354 VSS 0.023105f
C8991 PAD.n10355 VSS 0.03055f
C8992 PAD.n10356 VSS 0.040018f
C8993 PAD.n10357 VSS 0.033766f
C8994 PAD.n10358 VSS 0.024313f
C8995 PAD.n10359 VSS 0.027838f
C8996 PAD.n10360 VSS 0.027838f
C8997 PAD.n10361 VSS 0.522836f
C8998 PAD.n10362 VSS 0.261418f
C8999 PAD.n10363 VSS 0.045001f
C9000 PAD.n10364 VSS 0.045001f
C9001 PAD.n10365 VSS 0.03565f
C9002 PAD.n10366 VSS 8.753309f
C9003 PAD.n10367 VSS 0.041759f
C9004 PAD.n10368 VSS 0.053224f
C9005 PAD.n10369 VSS 0.047199f
C9006 PAD.n10370 VSS 0.062262f
C9007 PAD.n10371 VSS 0.069752f
C9008 PAD.n10372 VSS 0.069752f
C9009 PAD.n10373 VSS 0.700403f
C9010 PAD.n10374 VSS 0.591889f
C9011 PAD.n10375 VSS 0.047896f
C9012 PAD.n10376 VSS 0.047896f
C9013 PAD.n10377 VSS 0.029431f
C9014 PAD.n10378 VSS 0.025763f
C9015 PAD.n10379 VSS 0.025763f
C9016 PAD.n10380 VSS 0.022501f
C9017 PAD.n10381 VSS 0.033766f
C9018 PAD.n10382 VSS 0.03055f
C9019 PAD.n10383 VSS 0.036454f
C9020 PAD.n10384 VSS 0.036454f
C9021 PAD.n10385 VSS 0.036454f
C9022 PAD.n10387 VSS 0.023105f
C9023 PAD.n10388 VSS 0.438985f
C9024 PAD.n10389 VSS 0.330472f
C9025 PAD.n10390 VSS 0.051752f
C9026 PAD.n10391 VSS 0.051752f
C9027 PAD.n10392 VSS 0.046195f
C9028 PAD.n10393 VSS 0.062262f
C9029 PAD.n10394 VSS 0.054228f
C9030 PAD.n10395 VSS 0.060752f
C9031 PAD.n10396 VSS 0.060752f
C9032 PAD.n10397 VSS 0.187431f
C9033 PAD.n10398 VSS 0.611619f
C9034 PAD.n10399 VSS 0.0434f
C9035 PAD.n10400 VSS 0.0434f
C9036 PAD.n10401 VSS 0.037904f
C9037 PAD.n10402 VSS 0.033766f
C9038 PAD.n10403 VSS 0.042887f
C9039 PAD.n10404 VSS 0.026427f
C9040 PAD.n10405 VSS 0.030259f
C9041 PAD.n10406 VSS 0.030259f
C9042 PAD.n10407 VSS 0.192364f
C9043 PAD.n10408 VSS 0.512971f
C9044 PAD.n10409 VSS 0.043876f
C9045 PAD.n10410 VSS 0.043876f
C9046 PAD.n10411 VSS 0.039165f
C9047 PAD.n10412 VSS 0.062262f
C9048 PAD.n10413 VSS 0.036454f
C9049 PAD.n10414 VSS 0.036454f
C9050 PAD.n10415 VSS 0.036454f
C9051 PAD.n10417 VSS 0.036454f
C9052 PAD.n10418 VSS 0.036454f
C9053 PAD.n10419 VSS 0.036454f
C9054 PAD.n10420 VSS 0.036454f
C9055 PAD.n10422 VSS 0.036454f
C9056 PAD.n10423 VSS 0.036454f
C9057 PAD.n10424 VSS 0.036454f
C9058 PAD.n10425 VSS 0.036454f
C9059 PAD.n10427 VSS 0.036454f
C9060 PAD.n10428 VSS 0.036454f
C9061 PAD.n10429 VSS 0.036454f
C9062 PAD.n10430 VSS 0.036454f
C9063 PAD.n10432 VSS 0.036454f
C9064 PAD.n10433 VSS 0.036454f
C9065 PAD.n10434 VSS 0.036454f
C9066 PAD.n10435 VSS 0.036454f
C9067 PAD.n10437 VSS 0.036454f
C9068 PAD.n10438 VSS 0.036454f
C9069 PAD.n10439 VSS 0.036454f
C9070 PAD.n10440 VSS 0.036454f
C9071 PAD.n10442 VSS 0.036454f
C9072 PAD.n10443 VSS 0.036454f
C9073 PAD.n10444 VSS 0.036454f
C9074 PAD.n10445 VSS 0.036454f
C9075 PAD.n10447 VSS 0.036454f
C9076 PAD.n10448 VSS 0.036454f
C9077 PAD.n10449 VSS 0.036454f
C9078 PAD.n10450 VSS 0.036454f
C9079 PAD.n10452 VSS 0.036454f
C9080 PAD.n10453 VSS 0.036454f
C9081 PAD.n10454 VSS 0.036454f
C9082 PAD.n10455 VSS 0.036454f
C9083 PAD.n10457 VSS 0.036454f
C9084 PAD.n10458 VSS 0.036454f
C9085 PAD.n10459 VSS 0.036454f
C9086 PAD.n10460 VSS 0.036454f
C9087 PAD.n10462 VSS 0.036454f
C9088 PAD.n10463 VSS 0.036454f
C9089 PAD.n10464 VSS 0.036454f
C9090 PAD.n10465 VSS 0.036454f
C9091 PAD.n10467 VSS 0.036454f
C9092 PAD.n10468 VSS 0.036454f
C9093 PAD.n10469 VSS 0.036454f
C9094 PAD.n10470 VSS 0.036454f
C9095 PAD.n10472 VSS 0.036454f
C9096 PAD.n10473 VSS 0.036454f
C9097 PAD.n10474 VSS 0.036454f
C9098 PAD.n10475 VSS 0.036454f
C9099 PAD.n10477 VSS 0.036454f
C9100 PAD.n10478 VSS 0.036454f
C9101 PAD.n10479 VSS 0.036454f
C9102 PAD.n10480 VSS 0.036454f
C9103 PAD.n10482 VSS 0.036454f
C9104 PAD.n10483 VSS 0.036454f
C9105 PAD.n10484 VSS 0.036454f
C9106 PAD.n10485 VSS 0.036454f
C9107 PAD.n10487 VSS 0.036454f
C9108 PAD.n10488 VSS 0.036454f
C9109 PAD.n10489 VSS 0.036454f
C9110 PAD.n10490 VSS 0.036454f
C9111 PAD.n10492 VSS 0.036454f
C9112 PAD.n10493 VSS 0.036454f
C9113 PAD.n10494 VSS 0.036454f
C9114 PAD.n10495 VSS 0.036454f
C9115 PAD.n10497 VSS 0.036454f
C9116 PAD.n10498 VSS 0.036454f
C9117 PAD.n10499 VSS 0.036454f
C9118 PAD.n10500 VSS 0.036454f
C9119 PAD.n10502 VSS 0.036454f
C9120 PAD.n10503 VSS 0.036454f
C9121 PAD.n10504 VSS 0.036454f
C9122 PAD.n10505 VSS 0.036454f
C9123 PAD.n10507 VSS 0.036454f
C9124 PAD.n10508 VSS 0.036454f
C9125 PAD.n10509 VSS 0.036454f
C9126 PAD.n10510 VSS 0.036454f
C9127 PAD.n10512 VSS 0.036454f
C9128 PAD.n10513 VSS 0.036454f
C9129 PAD.n10515 VSS 0.036454f
C9130 PAD.n10516 VSS 0.036454f
C9131 PAD.n10517 VSS 0.036454f
C9132 PAD.n10518 VSS 0.036454f
C9133 PAD.n10519 VSS 0.036454f
C9134 PAD.n10520 VSS 0.036454f
C9135 PAD.n10521 VSS 0.036454f
C9136 PAD.n10522 VSS 0.036454f
C9137 PAD.n10524 VSS 0.036454f
C9138 PAD.n10525 VSS 0.036454f
C9139 PAD.n10526 VSS 0.036454f
C9140 PAD.n10527 VSS 0.036454f
C9141 PAD.n10528 VSS 0.036454f
C9142 PAD.n10529 VSS 0.036454f
C9143 PAD.n10530 VSS 0.036454f
C9144 PAD.n10531 VSS 0.036454f
C9145 PAD.n10533 VSS 0.036454f
C9146 PAD.n10534 VSS 0.036454f
C9147 PAD.n10535 VSS 0.036454f
C9148 PAD.n10536 VSS 0.036454f
C9149 PAD.n10537 VSS 0.036454f
C9150 PAD.n10538 VSS 0.036454f
C9151 PAD.n10539 VSS 0.036454f
C9152 PAD.n10540 VSS 0.036454f
C9153 PAD.n10542 VSS 0.036454f
C9154 PAD.n10543 VSS 0.036454f
C9155 PAD.n10544 VSS 0.036454f
C9156 PAD.n10545 VSS 0.036454f
C9157 PAD.n10546 VSS 0.036454f
C9158 PAD.n10547 VSS 0.036454f
C9159 PAD.n10548 VSS 0.036454f
C9160 PAD.n10549 VSS 0.036454f
C9161 PAD.n10551 VSS 0.036454f
C9162 PAD.n10552 VSS 0.036454f
C9163 PAD.n10553 VSS 0.036454f
C9164 PAD.n10554 VSS 0.036454f
C9165 PAD.n10555 VSS 0.036454f
C9166 PAD.n10556 VSS 0.036454f
C9167 PAD.n10557 VSS 0.036454f
C9168 PAD.n10558 VSS 0.036454f
C9169 PAD.n10560 VSS 0.036454f
C9170 PAD.n10561 VSS 0.036454f
C9171 PAD.n10562 VSS 0.036454f
C9172 PAD.n10563 VSS 0.036454f
C9173 PAD.n10564 VSS 0.036454f
C9174 PAD.n10565 VSS 0.036454f
C9175 PAD.n10566 VSS 0.036454f
C9176 PAD.n10567 VSS 0.036454f
C9177 PAD.n10569 VSS 0.036454f
C9178 PAD.n10570 VSS 0.036454f
C9179 PAD.n10571 VSS 0.036454f
C9180 PAD.n10572 VSS 0.036454f
C9181 PAD.n10573 VSS 0.036454f
C9182 PAD.n10574 VSS 0.036454f
C9183 PAD.n10575 VSS 0.036454f
C9184 PAD.n10576 VSS 0.036454f
C9185 PAD.n10578 VSS 0.036454f
C9186 PAD.n10579 VSS 0.036454f
C9187 PAD.n10580 VSS 0.036454f
C9188 PAD.n10581 VSS 0.036454f
C9189 PAD.n10582 VSS 0.036454f
C9190 PAD.n10583 VSS 0.036454f
C9191 PAD.n10584 VSS 0.036454f
C9192 PAD.n10585 VSS 0.036454f
C9193 PAD.n10587 VSS 0.036454f
C9194 PAD.n10588 VSS 0.036454f
C9195 PAD.n10589 VSS 0.036454f
C9196 PAD.n10590 VSS 0.036454f
C9197 PAD.n10591 VSS 0.036454f
C9198 PAD.n10592 VSS 0.036454f
C9199 PAD.n10593 VSS 0.036454f
C9200 PAD.n10594 VSS 0.036454f
C9201 PAD.n10596 VSS 0.036454f
C9202 PAD.n10597 VSS 0.036454f
C9203 PAD.n10598 VSS 0.036454f
C9204 PAD.n10599 VSS 0.036454f
C9205 PAD.n10600 VSS 0.036454f
C9206 PAD.n10601 VSS 0.036454f
C9207 PAD.n10602 VSS 0.036454f
C9208 PAD.n10603 VSS 0.036454f
C9209 PAD.n10605 VSS 0.036454f
C9210 PAD.n10606 VSS 0.036454f
C9211 PAD.n10607 VSS 0.036454f
C9212 PAD.n10608 VSS 0.036454f
C9213 PAD.n10609 VSS 0.036454f
C9214 PAD.n10610 VSS 0.036454f
C9215 PAD.n10611 VSS 0.036454f
C9216 PAD.n10612 VSS 0.036454f
C9217 PAD.n10614 VSS 0.036454f
C9218 PAD.n10615 VSS 0.036454f
C9219 PAD.n10616 VSS 0.036454f
C9220 PAD.n10617 VSS 0.036454f
C9221 PAD.n10618 VSS 0.036454f
C9222 PAD.n10619 VSS 0.036454f
C9223 PAD.n10620 VSS 0.036454f
C9224 PAD.n10621 VSS 0.036454f
C9225 PAD.n10623 VSS 0.036454f
C9226 PAD.n10624 VSS 0.036454f
C9227 PAD.n10625 VSS 0.036454f
C9228 PAD.n10626 VSS 0.036454f
C9229 PAD.n10627 VSS 0.036454f
C9230 PAD.n10628 VSS 0.036454f
C9231 PAD.n10629 VSS 0.036454f
C9232 PAD.n10630 VSS 0.036454f
C9233 PAD.n10632 VSS 0.036454f
C9234 PAD.n10633 VSS 0.036454f
C9235 PAD.n10634 VSS 0.036454f
C9236 PAD.n10635 VSS 0.036454f
C9237 PAD.n10636 VSS 0.036454f
C9238 PAD.n10637 VSS 0.036454f
C9239 PAD.n10638 VSS 0.036454f
C9240 PAD.n10639 VSS 0.036454f
C9241 PAD.n10641 VSS 0.036454f
C9242 PAD.n10642 VSS 0.036454f
C9243 PAD.n10643 VSS 0.036454f
C9244 PAD.n10644 VSS 0.036454f
C9245 PAD.n10645 VSS 0.036454f
C9246 PAD.n10646 VSS 0.036454f
C9247 PAD.n10647 VSS 0.036454f
C9248 PAD.n10648 VSS 0.036454f
C9249 PAD.n10650 VSS 0.036454f
C9250 PAD.n10651 VSS 0.036454f
C9251 PAD.n10652 VSS 0.036454f
C9252 PAD.n10653 VSS 0.036454f
C9253 PAD.n10654 VSS 0.036454f
C9254 PAD.n10655 VSS 0.036454f
C9255 PAD.n10656 VSS 0.036454f
C9256 PAD.n10657 VSS 0.036454f
C9257 PAD.n10659 VSS 0.036454f
C9258 PAD.n10660 VSS 0.036454f
C9259 PAD.n10661 VSS 0.036454f
C9260 PAD.n10662 VSS 0.036454f
C9261 PAD.n10663 VSS 0.036454f
C9262 PAD.n10664 VSS 0.036454f
C9263 PAD.n10665 VSS 0.036454f
C9264 PAD.n10666 VSS 0.036454f
C9265 PAD.n10668 VSS 0.036454f
C9266 PAD.n10669 VSS 0.036454f
C9267 PAD.n10670 VSS 0.036454f
C9268 PAD.n10671 VSS 0.036454f
C9269 PAD.n10672 VSS 0.036454f
C9270 PAD.n10673 VSS 0.036454f
C9271 PAD.n10674 VSS 0.036454f
C9272 PAD.n10675 VSS 0.036454f
C9273 PAD.n10677 VSS 0.036454f
C9274 PAD.n10678 VSS 0.036454f
C9275 PAD.n10679 VSS 0.036454f
C9276 PAD.n10680 VSS 0.036454f
C9277 PAD.n10681 VSS 0.036454f
C9278 PAD.n10682 VSS 0.036454f
C9279 PAD.n10683 VSS 0.036454f
C9280 PAD.n10684 VSS 0.036454f
C9281 PAD.n10686 VSS 0.036454f
C9282 PAD.n10687 VSS 0.036454f
C9283 PAD.n10688 VSS 0.036454f
C9284 PAD.n10689 VSS 0.036454f
C9285 PAD.n10690 VSS 0.036454f
C9286 PAD.n10691 VSS 0.036454f
C9287 PAD.n10693 VSS 0.036454f
C9288 PAD.n10694 VSS 0.036454f
C9289 PAD.n10695 VSS 0.023105f
C9290 PAD.n10696 VSS 0.033374f
C9291 PAD.n10697 VSS 0.046278f
C9292 PAD.n10698 VSS 0.061258f
C9293 PAD.n10699 VSS 0.068627f
C9294 PAD.n10700 VSS 0.068627f
C9295 PAD.n10701 VSS 0.700403f
C9296 PAD.n10702 VSS 0.22689f
C9297 PAD.n10703 VSS 0.038904f
C9298 PAD.n10704 VSS 0.038904f
C9299 PAD.n10705 VSS 0.029431f
C9300 PAD.n10706 VSS 0.034755f
C9301 PAD.n10707 VSS 0.034755f
C9302 PAD.n10708 VSS 0.030353f
C9303 PAD.n10709 VSS 0.033766f
C9304 PAD.n10710 VSS 0.03055f
C9305 PAD.n10711 VSS 0.036454f
C9306 PAD.n10712 VSS 0.036454f
C9307 PAD.n10713 VSS 0.036454f
C9308 PAD.n10715 VSS 0.023105f
C9309 PAD.n10716 VSS 0.340336f
C9310 PAD.n10717 VSS 0.616552f
C9311 PAD.n10718 VSS 0.611619f
C9312 PAD.n10719 VSS 0.656011f
C9313 PAD.n10720 VSS 0.069752f
C9314 PAD.n10721 VSS 0.069752f
C9315 PAD.n10722 VSS 0.062262f
C9316 PAD.n10723 VSS 0.062262f
C9317 PAD.n10724 VSS 0.037156f
C9318 PAD.n10725 VSS 0.041626f
C9319 PAD.n10726 VSS 0.041626f
C9320 PAD.n10727 VSS 0.616552f
C9321 PAD.n10728 VSS 0.24662f
C9322 PAD.n10729 VSS 0.034409f
C9323 PAD.n10730 VSS 0.034409f
C9324 PAD.n10731 VSS 0.030051f
C9325 PAD.n10732 VSS 0.033766f
C9326 PAD.n10733 VSS 0.03428f
C9327 PAD.n10734 VSS 0.03055f
C9328 PAD.n10735 VSS 0.042887f
C9329 PAD.n10736 VSS 0.029431f
C9330 PAD.n10737 VSS 0.049106f
C9331 PAD.n10738 VSS 0.029431f
C9332 PAD.n10739 VSS 0.049106f
C9333 PAD.n10740 VSS 0.207161f
C9334 PAD.n10741 VSS 0.611619f
C9335 PAD.n10742 VSS 0.055127f
C9336 PAD.n10743 VSS 0.068065f
C9337 PAD.n10744 VSS 0.055127f
C9338 PAD.n10745 VSS 0.068065f
C9339 PAD.n10746 VSS 0.044186f
C9340 PAD.n10747 VSS 0.036454f
C9341 PAD.n10748 VSS 0.039754f
C9342 PAD.n10749 VSS 0.036454f
C9343 PAD.n10750 VSS 0.039754f
C9344 PAD.n10751 VSS 0.049502f
C9345 PAD.n10752 VSS 0.049502f
C9346 PAD.n10753 VSS 0.207161f
C9347 PAD.n10754 VSS 0.596822f
C9348 PAD.n10755 VSS 0.508039f
C9349 PAD.n10757 VSS 0.036454f
C9350 PAD.n10758 VSS 0.036454f
C9351 PAD.n10759 VSS 0.036454f
C9352 PAD.n10761 VSS 0.036454f
C9353 PAD.n10762 VSS 0.036454f
C9354 PAD.n10763 VSS 0.036454f
C9355 PAD.n10765 VSS 0.036454f
C9356 PAD.n10766 VSS 0.036454f
C9357 PAD.n10767 VSS 0.036454f
C9358 PAD.n10769 VSS 0.036454f
C9359 PAD.n10770 VSS 0.036454f
C9360 PAD.n10771 VSS 0.036454f
C9361 PAD.n10773 VSS 0.036454f
C9362 PAD.n10774 VSS 0.036454f
C9363 PAD.n10775 VSS 0.036454f
C9364 PAD.n10777 VSS 0.036454f
C9365 PAD.n10778 VSS 0.036454f
C9366 PAD.n10779 VSS 0.036454f
C9367 PAD.n10781 VSS 0.036454f
C9368 PAD.n10782 VSS 0.036454f
C9369 PAD.n10783 VSS 0.036454f
C9370 PAD.n10785 VSS 0.036454f
C9371 PAD.n10786 VSS 0.036454f
C9372 PAD.n10787 VSS 0.036454f
C9373 PAD.n10789 VSS 0.036454f
C9374 PAD.n10790 VSS 0.036454f
C9375 PAD.n10791 VSS 0.036454f
C9376 PAD.n10793 VSS 0.036454f
C9377 PAD.n10794 VSS 0.036454f
C9378 PAD.n10795 VSS 0.036454f
C9379 PAD.n10797 VSS 0.036454f
C9380 PAD.n10798 VSS 0.036454f
C9381 PAD.n10799 VSS 0.036454f
C9382 PAD.n10801 VSS 0.036454f
C9383 PAD.n10802 VSS 0.036454f
C9384 PAD.n10803 VSS 0.036454f
C9385 PAD.n10805 VSS 0.036454f
C9386 PAD.n10806 VSS 0.036454f
C9387 PAD.n10807 VSS 0.036454f
C9388 PAD.n10809 VSS 0.036454f
C9389 PAD.n10810 VSS 0.036454f
C9390 PAD.n10811 VSS 0.036454f
C9391 PAD.n10813 VSS 0.036454f
C9392 PAD.n10814 VSS 0.036454f
C9393 PAD.n10815 VSS 0.036454f
C9394 PAD.n10817 VSS 0.036454f
C9395 PAD.n10818 VSS 0.036454f
C9396 PAD.n10819 VSS 0.036454f
C9397 PAD.n10821 VSS 0.036454f
C9398 PAD.n10822 VSS 0.036454f
C9399 PAD.n10823 VSS 0.036454f
C9400 PAD.n10825 VSS 0.036454f
C9401 PAD.n10826 VSS 0.036454f
C9402 PAD.n10827 VSS 0.036454f
C9403 PAD.n10829 VSS 0.036454f
C9404 PAD.n10830 VSS 0.036454f
C9405 PAD.n10831 VSS 0.036454f
C9406 PAD.n10833 VSS 0.036454f
C9407 PAD.n10834 VSS 0.036454f
C9408 PAD.n10835 VSS 0.036454f
C9409 PAD.n10837 VSS 0.023105f
C9410 PAD.n10838 VSS 0.023105f
C9411 PAD.n10839 VSS 0.036454f
C9412 PAD.n10840 VSS 0.036454f
C9413 PAD.n10841 VSS 0.036454f
C9414 PAD.n10843 VSS 0.036454f
C9415 PAD.n10845 VSS 0.036454f
C9416 PAD.n10847 VSS 0.036454f
C9417 PAD.n10848 VSS 0.036454f
C9418 PAD.n10849 VSS 0.036454f
C9419 PAD.n10850 VSS 0.036454f
C9420 PAD.n10851 VSS 0.036454f
C9421 PAD.n10852 VSS 0.036454f
C9422 PAD.n10853 VSS 0.036454f
C9423 PAD.n10855 VSS 0.036454f
C9424 PAD.n10857 VSS 0.036454f
C9425 PAD.n10859 VSS 0.036454f
C9426 PAD.n10860 VSS 0.036454f
C9427 PAD.n10861 VSS 0.036454f
C9428 PAD.n10862 VSS 0.036454f
C9429 PAD.n10863 VSS 0.036454f
C9430 PAD.n10864 VSS 0.036454f
C9431 PAD.n10865 VSS 0.036454f
C9432 PAD.n10867 VSS 0.036454f
C9433 PAD.n10869 VSS 0.036454f
C9434 PAD.n10871 VSS 0.036454f
C9435 PAD.n10872 VSS 0.036454f
C9436 PAD.n10873 VSS 0.036454f
C9437 PAD.n10874 VSS 0.036454f
C9438 PAD.n10875 VSS 0.036454f
C9439 PAD.n10876 VSS 0.036454f
C9440 PAD.n10877 VSS 0.036454f
C9441 PAD.n10879 VSS 0.036454f
C9442 PAD.n10881 VSS 0.036454f
C9443 PAD.n10883 VSS 0.036454f
C9444 PAD.n10884 VSS 0.036454f
C9445 PAD.n10885 VSS 0.036454f
C9446 PAD.n10886 VSS 0.036454f
C9447 PAD.n10887 VSS 0.036454f
C9448 PAD.n10888 VSS 0.036454f
C9449 PAD.n10889 VSS 0.036454f
C9450 PAD.n10891 VSS 0.036454f
C9451 PAD.n10893 VSS 0.036454f
C9452 PAD.n10895 VSS 0.036454f
C9453 PAD.n10896 VSS 0.036454f
C9454 PAD.n10897 VSS 0.036454f
C9455 PAD.n10898 VSS 0.036454f
C9456 PAD.n10899 VSS 0.036454f
C9457 PAD.n10900 VSS 0.036454f
C9458 PAD.n10901 VSS 0.036454f
C9459 PAD.n10903 VSS 0.036454f
C9460 PAD.n10905 VSS 0.036454f
C9461 PAD.n10907 VSS 0.036454f
C9462 PAD.n10908 VSS 0.036454f
C9463 PAD.n10909 VSS 0.036454f
C9464 PAD.n10910 VSS 0.036454f
C9465 PAD.n10911 VSS 0.036454f
C9466 PAD.n10912 VSS 0.036454f
C9467 PAD.n10913 VSS 0.036454f
C9468 PAD.n10915 VSS 0.036454f
C9469 PAD.n10917 VSS 0.036454f
C9470 PAD.n10919 VSS 0.036454f
C9471 PAD.n10920 VSS 0.036454f
C9472 PAD.n10921 VSS 0.036454f
C9473 PAD.n10922 VSS 0.036454f
C9474 PAD.n10923 VSS 0.036454f
C9475 PAD.n10924 VSS 0.036454f
C9476 PAD.n10925 VSS 0.036454f
C9477 PAD.n10927 VSS 0.036454f
C9478 PAD.n10929 VSS 0.036454f
C9479 PAD.n10931 VSS 0.036454f
C9480 PAD.n10932 VSS 0.036454f
C9481 PAD.n10933 VSS 0.036454f
C9482 PAD.n10934 VSS 0.036454f
C9483 PAD.n10935 VSS 0.036454f
C9484 PAD.n10936 VSS 0.036454f
C9485 PAD.n10937 VSS 0.036454f
C9486 PAD.n10939 VSS 0.036454f
C9487 PAD.n10941 VSS 0.036454f
C9488 PAD.n10943 VSS 0.036454f
C9489 PAD.n10944 VSS 0.036454f
C9490 PAD.n10945 VSS 0.036454f
C9491 PAD.n10946 VSS 0.036454f
C9492 PAD.n10947 VSS 0.036454f
C9493 PAD.n10948 VSS 0.036454f
C9494 PAD.n10949 VSS 0.036454f
C9495 PAD.n10951 VSS 0.036454f
C9496 PAD.n10953 VSS 0.036454f
C9497 PAD.n10955 VSS 0.036454f
C9498 PAD.n10956 VSS 0.036454f
C9499 PAD.n10957 VSS 0.036454f
C9500 PAD.n10958 VSS 0.036454f
C9501 PAD.n10959 VSS 0.036454f
C9502 PAD.n10960 VSS 0.036454f
C9503 PAD.n10961 VSS 0.036454f
C9504 PAD.n10963 VSS 0.036454f
C9505 PAD.n10965 VSS 0.036454f
C9506 PAD.n10967 VSS 0.036454f
C9507 PAD.n10968 VSS 0.036454f
C9508 PAD.n10969 VSS 0.036454f
C9509 PAD.n10970 VSS 0.036454f
C9510 PAD.n10971 VSS 0.036454f
C9511 PAD.n10972 VSS 0.036454f
C9512 PAD.n10973 VSS 0.036454f
C9513 PAD.n10975 VSS 0.036454f
C9514 PAD.n10977 VSS 0.036454f
C9515 PAD.n10979 VSS 0.036454f
C9516 PAD.n10980 VSS 0.036454f
C9517 PAD.n10981 VSS 0.036454f
C9518 PAD.n10982 VSS 0.036454f
C9519 PAD.n10983 VSS 0.036454f
C9520 PAD.n10984 VSS 0.036454f
C9521 PAD.n10985 VSS 0.036454f
C9522 PAD.n10987 VSS 0.036454f
C9523 PAD.n10989 VSS 0.036454f
C9524 PAD.n10991 VSS 0.036454f
C9525 PAD.n10992 VSS 0.036454f
C9526 PAD.n10993 VSS 0.036454f
C9527 PAD.n10994 VSS 0.036454f
C9528 PAD.n10995 VSS 0.036454f
C9529 PAD.n10996 VSS 0.036454f
C9530 PAD.n10997 VSS 0.036454f
C9531 PAD.n10999 VSS 0.036454f
C9532 PAD.n11001 VSS 0.036454f
C9533 PAD.n11003 VSS 0.036454f
C9534 PAD.n11004 VSS 0.036454f
C9535 PAD.n11005 VSS 0.036454f
C9536 PAD.n11006 VSS 0.036454f
C9537 PAD.n11007 VSS 0.036454f
C9538 PAD.n11008 VSS 0.036454f
C9539 PAD.n11009 VSS 0.036454f
C9540 PAD.n11011 VSS 0.036454f
C9541 PAD.n11013 VSS 0.036454f
C9542 PAD.n11015 VSS 0.036454f
C9543 PAD.n11016 VSS 0.036454f
C9544 PAD.n11017 VSS 0.036454f
C9545 PAD.n11018 VSS 0.036454f
C9546 PAD.n11019 VSS 0.036454f
C9547 PAD.n11020 VSS 0.036454f
C9548 PAD.n11021 VSS 0.036454f
C9549 PAD.n11023 VSS 0.036454f
C9550 PAD.n11025 VSS 0.036454f
C9551 PAD.n11027 VSS 0.036454f
C9552 PAD.n11028 VSS 0.036454f
C9553 PAD.n11029 VSS 0.036454f
C9554 PAD.n11030 VSS 0.036454f
C9555 PAD.n11031 VSS 0.036454f
C9556 PAD.n11032 VSS 0.036454f
C9557 PAD.n11033 VSS 0.036454f
C9558 PAD.n11035 VSS 0.036454f
C9559 PAD.n11037 VSS 0.036454f
C9560 PAD.n11039 VSS 0.036454f
C9561 PAD.n11040 VSS 0.036454f
C9562 PAD.n11041 VSS 0.036454f
C9563 PAD.n11042 VSS 0.036454f
C9564 PAD.n11043 VSS 0.036454f
C9565 PAD.n11044 VSS 0.036454f
C9566 PAD.n11045 VSS 0.036454f
C9567 PAD.n11047 VSS 0.036454f
C9568 PAD.n11049 VSS 0.036454f
C9569 PAD.n11051 VSS 0.036454f
C9570 PAD.n11052 VSS 0.036454f
C9571 PAD.n11053 VSS 0.036454f
C9572 PAD.n11054 VSS 0.036454f
C9573 PAD.n11055 VSS 0.036454f
C9574 PAD.n11056 VSS 0.036454f
C9575 PAD.n11057 VSS 0.036454f
C9576 PAD.n11059 VSS 0.036454f
C9577 PAD.n11061 VSS 0.036454f
C9578 PAD.n11063 VSS 0.036454f
C9579 PAD.n11064 VSS 0.036454f
C9580 PAD.n11065 VSS 0.036454f
C9581 PAD.n11066 VSS 0.036454f
C9582 PAD.n11067 VSS 0.036454f
C9583 PAD.n11068 VSS 0.036454f
C9584 PAD.n11069 VSS 0.036454f
C9585 PAD.n11071 VSS 0.036454f
C9586 PAD.n11073 VSS 0.036454f
C9587 PAD.n11075 VSS 0.036454f
C9588 PAD.n11076 VSS 0.036454f
C9589 PAD.n11077 VSS 0.036454f
C9590 PAD.n11078 VSS 0.036454f
C9591 PAD.n11079 VSS 0.036454f
C9592 PAD.n11080 VSS 0.036454f
C9593 PAD.n11081 VSS 0.036454f
C9594 PAD.n11083 VSS 0.036454f
C9595 PAD.n11085 VSS 0.023105f
C9596 PAD.n11086 VSS 0.023105f
C9597 PAD.n11087 VSS 0.033374f
C9598 PAD.n11088 VSS 0.046278f
C9599 PAD.n11089 VSS 0.049207f
C9600 PAD.n11090 VSS 0.128354f
C9601 PAD.n11091 VSS 0.103594f
C9602 PAD.n11092 VSS 0.07064f
C9603 PAD.n11093 VSS 0.103594f
C9604 PAD.n11094 VSS 0.07064f
C9605 PAD.n11096 VSS 0.61162f
C9606 PAD.n11097 VSS 0.853308f
C9607 PAD.n11098 VSS 0.769457f
C9608 PAD.n11099 VSS 0.61162f
C9609 PAD.n11100 VSS 0.61162f
C9610 PAD.n11101 VSS 0.069163f
C9611 PAD.n11102 VSS 0.069163f
C9612 PAD.n11104 VSS 0.103594f
C9613 PAD.n11105 VSS 1.55864f
C9614 PAD.n11106 VSS 0.103594f
C9615 PAD.n11107 VSS 0.074902f
C9616 PAD.n11108 VSS 0.074902f
C9617 PAD.n11109 VSS 0.074902f
C9618 PAD.n11110 VSS 0.074902f
C9619 PAD.n11111 VSS 0.074902f
C9620 PAD.n11112 VSS 0.074902f
C9621 PAD.n11113 VSS 0.074902f
C9622 PAD.n11114 VSS 0.074902f
C9623 PAD.n11115 VSS 0.074902f
C9624 PAD.n11116 VSS 0.074902f
C9625 PAD.n11117 VSS 0.074902f
C9626 PAD.n11118 VSS 0.074902f
C9627 PAD.n11119 VSS 0.074902f
C9628 PAD.n11120 VSS 0.074902f
C9629 PAD.n11121 VSS 0.074902f
C9630 PAD.n11122 VSS 0.074902f
C9631 PAD.n11123 VSS 0.074902f
C9632 PAD.n11124 VSS 0.074902f
C9633 PAD.n11125 VSS 0.074902f
C9634 PAD.n11126 VSS 0.074902f
C9635 PAD.n11127 VSS 0.074902f
C9636 PAD.n11128 VSS 0.074902f
C9637 PAD.n11129 VSS 0.074902f
C9638 PAD.n11130 VSS 0.074902f
C9639 PAD.n11131 VSS 0.074902f
C9640 PAD.n11132 VSS 0.074902f
C9641 PAD.n11133 VSS 0.074902f
C9642 PAD.n11134 VSS 0.074902f
C9643 PAD.n11135 VSS 0.074902f
C9644 PAD.n11136 VSS 0.074902f
C9645 PAD.n11137 VSS 0.074902f
C9646 PAD.n11138 VSS 0.074902f
C9647 PAD.n11139 VSS 0.074902f
C9648 PAD.n11140 VSS 0.074902f
C9649 PAD.n11141 VSS 0.074902f
C9650 PAD.n11142 VSS 0.074902f
C9651 PAD.n11143 VSS 0.074902f
C9652 PAD.n11144 VSS 0.074902f
C9653 PAD.n11145 VSS 0.074902f
C9654 PAD.n11146 VSS 0.074902f
C9655 PAD.n11147 VSS 0.074902f
C9656 PAD.n11148 VSS 0.074902f
C9657 PAD.n11149 VSS 0.074902f
C9658 PAD.n11150 VSS 0.074902f
C9659 PAD.n11151 VSS 0.074902f
C9660 PAD.n11152 VSS 0.074902f
C9661 PAD.n11153 VSS 0.074902f
C9662 PAD.n11154 VSS 0.074902f
C9663 PAD.n11156 VSS 0.059499f
C9664 PAD.n11158 VSS 0.074902f
C9665 PAD.n11160 VSS 0.074902f
C9666 PAD.n11162 VSS 0.074902f
C9667 PAD.n11164 VSS 0.074902f
C9668 PAD.n11166 VSS 0.074902f
C9669 PAD.n11168 VSS 0.074902f
C9670 PAD.n11170 VSS 0.074902f
C9671 PAD.n11172 VSS 0.074902f
C9672 PAD.n11174 VSS 0.074902f
C9673 PAD.n11176 VSS 0.074902f
C9674 PAD.n11178 VSS 0.074902f
C9675 PAD.n11180 VSS 0.074902f
C9676 PAD.n11182 VSS 0.074902f
C9677 PAD.n11184 VSS 0.074902f
C9678 PAD.n11186 VSS 0.074902f
C9679 PAD.n11188 VSS 0.074902f
C9680 PAD.n11190 VSS 0.074902f
C9681 PAD.n11192 VSS 0.074902f
C9682 PAD.n11194 VSS 0.074902f
C9683 PAD.n11196 VSS 0.074902f
C9684 PAD.n11198 VSS 0.074902f
C9685 PAD.n11200 VSS 0.074902f
C9686 PAD.n11202 VSS 0.074902f
C9687 PAD.n11204 VSS 0.074902f
C9688 PAD.n11206 VSS 0.074902f
C9689 PAD.n11208 VSS 0.074902f
C9690 PAD.n11210 VSS 0.074902f
C9691 PAD.n11212 VSS 0.074902f
C9692 PAD.n11214 VSS 0.074902f
C9693 PAD.n11216 VSS 0.074902f
C9694 PAD.n11218 VSS 0.074902f
C9695 PAD.n11220 VSS 0.074902f
C9696 PAD.n11222 VSS 0.074902f
C9697 PAD.n11224 VSS 0.074902f
C9698 PAD.n11226 VSS 0.074902f
C9699 PAD.n11228 VSS 0.074902f
C9700 PAD.n11230 VSS 0.074902f
C9701 PAD.n11232 VSS 0.074902f
C9702 PAD.n11234 VSS 0.074902f
C9703 PAD.n11236 VSS 0.074902f
C9704 PAD.n11238 VSS 0.074902f
C9705 PAD.n11240 VSS 0.074902f
C9706 PAD.n11242 VSS 0.074902f
C9707 PAD.n11244 VSS 0.074902f
C9708 PAD.n11246 VSS 0.074902f
C9709 PAD.n11248 VSS 0.074902f
C9710 PAD.n11250 VSS 0.074902f
C9711 PAD.n11252 VSS 0.074902f
C9712 PAD.n11253 VSS 0.044886f
C9713 PAD.n11302 VSS 0.61162f
C9714 PAD.n11303 VSS 0.044886f
C9715 PAD.n11304 VSS 0.074902f
C9716 PAD.n11305 VSS 0.074902f
C9717 PAD.n11306 VSS 0.074902f
C9718 PAD.n11307 VSS 0.074902f
C9719 PAD.n11308 VSS 0.074902f
C9720 PAD.n11309 VSS 0.074902f
C9721 PAD.n11310 VSS 0.074902f
C9722 PAD.n11311 VSS 0.074902f
C9723 PAD.n11312 VSS 0.074902f
C9724 PAD.n11313 VSS 0.074902f
C9725 PAD.n11314 VSS 0.074902f
C9726 PAD.n11315 VSS 0.074902f
C9727 PAD.n11316 VSS 0.074902f
C9728 PAD.n11317 VSS 0.074902f
C9729 PAD.n11318 VSS 0.074902f
C9730 PAD.n11319 VSS 0.074902f
C9731 PAD.n11320 VSS 0.074902f
C9732 PAD.n11321 VSS 0.074902f
C9733 PAD.n11322 VSS 0.074902f
C9734 PAD.n11323 VSS 0.074902f
C9735 PAD.n11324 VSS 0.074902f
C9736 PAD.n11325 VSS 0.074902f
C9737 PAD.n11326 VSS 0.074902f
C9738 PAD.n11327 VSS 0.074902f
C9739 PAD.n11328 VSS 0.074902f
C9740 PAD.n11329 VSS 0.074902f
C9741 PAD.n11330 VSS 0.074902f
C9742 PAD.n11331 VSS 0.074902f
C9743 PAD.n11332 VSS 0.074902f
C9744 PAD.n11333 VSS 0.074902f
C9745 PAD.n11334 VSS 0.074902f
C9746 PAD.n11335 VSS 0.074902f
C9747 PAD.n11336 VSS 0.074902f
C9748 PAD.n11337 VSS 0.074902f
C9749 PAD.n11338 VSS 0.074902f
C9750 PAD.n11339 VSS 0.074902f
C9751 PAD.n11340 VSS 0.074902f
C9752 PAD.n11341 VSS 0.074902f
C9753 PAD.n11342 VSS 0.074902f
C9754 PAD.n11343 VSS 0.074902f
C9755 PAD.n11344 VSS 0.074902f
C9756 PAD.n11345 VSS 0.074902f
C9757 PAD.n11346 VSS 0.074902f
C9758 PAD.n11347 VSS 0.074902f
C9759 PAD.n11348 VSS 0.074902f
C9760 PAD.n11349 VSS 0.074902f
C9761 PAD.n11350 VSS 0.074902f
C9762 PAD.n11351 VSS 0.074902f
C9763 PAD.n11352 VSS 0.103594f
C9764 PAD.n11353 VSS 0.103594f
C9765 PAD.n11354 VSS 0.074902f
C9766 PAD.n11355 VSS 0.074902f
C9767 PAD.n11356 VSS 0.074902f
C9768 PAD.n11357 VSS 0.074902f
C9769 PAD.n11358 VSS 0.074902f
C9770 PAD.n11359 VSS 0.074902f
C9771 PAD.n11360 VSS 0.074902f
C9772 PAD.n11361 VSS 0.074902f
C9773 PAD.n11362 VSS 0.074902f
C9774 PAD.n11363 VSS 0.074902f
C9775 PAD.n11364 VSS 0.074902f
C9776 PAD.n11365 VSS 0.074902f
C9777 PAD.n11366 VSS 0.074902f
C9778 PAD.n11367 VSS 0.074902f
C9779 PAD.n11368 VSS 0.074902f
C9780 PAD.n11369 VSS 0.074902f
C9781 PAD.n11370 VSS 0.074902f
C9782 PAD.n11371 VSS 0.074902f
C9783 PAD.n11372 VSS 0.074902f
C9784 PAD.n11373 VSS 0.074902f
C9785 PAD.n11374 VSS 0.074902f
C9786 PAD.n11375 VSS 0.074902f
C9787 PAD.n11376 VSS 0.074902f
C9788 PAD.n11377 VSS 0.074902f
C9789 PAD.n11378 VSS 0.074902f
C9790 PAD.n11379 VSS 0.074902f
C9791 PAD.n11380 VSS 0.074902f
C9792 PAD.n11381 VSS 0.074902f
C9793 PAD.n11382 VSS 0.074902f
C9794 PAD.n11383 VSS 0.074902f
C9795 PAD.n11384 VSS 0.074902f
C9796 PAD.n11385 VSS 0.074902f
C9797 PAD.n11386 VSS 0.074902f
C9798 PAD.n11387 VSS 0.074902f
C9799 PAD.n11388 VSS 0.074902f
C9800 PAD.n11389 VSS 0.074902f
C9801 PAD.n11390 VSS 0.074902f
C9802 PAD.n11391 VSS 0.074902f
C9803 PAD.n11392 VSS 0.074902f
C9804 PAD.n11393 VSS 0.074902f
C9805 PAD.n11394 VSS 0.074902f
C9806 PAD.n11395 VSS 0.074902f
C9807 PAD.n11396 VSS 0.074902f
C9808 PAD.n11397 VSS 0.074902f
C9809 PAD.n11398 VSS 0.074902f
C9810 PAD.n11399 VSS 0.074902f
C9811 PAD.n11400 VSS 0.074902f
C9812 PAD.n11401 VSS 0.074902f
C9813 PAD.n11402 VSS 0.074902f
C9814 PAD.n11403 VSS 0.074902f
C9815 PAD.n11404 VSS 0.074902f
C9816 PAD.n11405 VSS 0.074902f
C9817 PAD.n11406 VSS 0.074902f
C9818 PAD.n11407 VSS 0.074902f
C9819 PAD.n11408 VSS 0.074902f
C9820 PAD.n11409 VSS 0.074902f
C9821 PAD.n11410 VSS 0.074902f
C9822 PAD.n11411 VSS 0.074902f
C9823 PAD.n11412 VSS 0.074902f
C9824 PAD.n11413 VSS 0.074902f
C9825 PAD.n11414 VSS 0.074902f
C9826 PAD.n11415 VSS 0.074902f
C9827 PAD.n11416 VSS 0.074902f
C9828 PAD.n11417 VSS 0.074902f
C9829 PAD.n11418 VSS 0.074902f
C9830 PAD.n11419 VSS 0.074902f
C9831 PAD.n11420 VSS 0.074902f
C9832 PAD.n11421 VSS 0.074902f
C9833 PAD.n11422 VSS 0.074902f
C9834 PAD.n11423 VSS 0.074902f
C9835 PAD.n11424 VSS 0.074902f
C9836 PAD.n11425 VSS 0.074902f
C9837 PAD.n11426 VSS 0.074902f
C9838 PAD.n11427 VSS 0.074902f
C9839 PAD.n11428 VSS 0.074902f
C9840 PAD.n11429 VSS 0.074902f
C9841 PAD.n11430 VSS 0.074902f
C9842 PAD.n11431 VSS 0.074902f
C9843 PAD.n11432 VSS 0.074902f
C9844 PAD.n11433 VSS 0.074902f
C9845 PAD.n11434 VSS 0.074902f
C9846 PAD.n11435 VSS 0.074902f
C9847 PAD.n11436 VSS 0.074902f
C9848 PAD.n11437 VSS 0.074902f
C9849 PAD.n11438 VSS 0.074902f
C9850 PAD.n11439 VSS 0.074902f
C9851 PAD.n11440 VSS 0.074902f
C9852 PAD.n11441 VSS 0.074902f
C9853 PAD.n11442 VSS 0.074902f
C9854 PAD.n11443 VSS 0.074902f
C9855 PAD.n11444 VSS 0.074902f
C9856 PAD.n11445 VSS 0.074902f
C9857 PAD.n11446 VSS 0.074902f
C9858 PAD.n11447 VSS 0.074902f
C9859 PAD.n11448 VSS 0.074902f
C9860 PAD.n11449 VSS 0.074902f
C9861 PAD.n11450 VSS 0.074902f
C9862 PAD.n11451 VSS 0.074902f
C9863 PAD.n11452 VSS 0.074902f
C9864 PAD.n11453 VSS 0.074902f
C9865 PAD.n11454 VSS 0.074902f
C9866 PAD.n11455 VSS 0.074902f
C9867 PAD.n11456 VSS 0.074902f
C9868 PAD.n11457 VSS 0.074902f
C9869 PAD.n11458 VSS 0.074902f
C9870 PAD.n11459 VSS 0.074902f
C9871 PAD.n11460 VSS 0.074902f
C9872 PAD.n11461 VSS 0.074902f
C9873 PAD.n11462 VSS 0.074902f
C9874 PAD.n11463 VSS 0.074902f
C9875 PAD.n11464 VSS 0.074902f
C9876 PAD.n11465 VSS 0.074902f
C9877 PAD.n11466 VSS 0.074902f
C9878 PAD.n11467 VSS 0.074902f
C9879 PAD.n11468 VSS 0.074902f
C9880 PAD.n11469 VSS 0.074902f
C9881 PAD.n11470 VSS 0.074902f
C9882 PAD.n11471 VSS 0.074902f
C9883 PAD.n11472 VSS 0.074902f
C9884 PAD.n11473 VSS 0.074902f
C9885 PAD.n11474 VSS 0.074902f
C9886 PAD.n11475 VSS 0.074902f
C9887 PAD.n11476 VSS 0.074902f
C9888 PAD.n11477 VSS 0.074902f
C9889 PAD.n11478 VSS 0.074902f
C9890 PAD.n11479 VSS 0.074902f
C9891 PAD.n11480 VSS 0.074902f
C9892 PAD.n11481 VSS 0.074902f
C9893 PAD.n11482 VSS 0.074902f
C9894 PAD.n11483 VSS 0.074902f
C9895 PAD.n11484 VSS 0.074902f
C9896 PAD.n11485 VSS 0.074902f
C9897 PAD.n11486 VSS 0.074902f
C9898 PAD.n11487 VSS 0.074902f
C9899 PAD.n11488 VSS 0.074902f
C9900 PAD.n11489 VSS 0.074902f
C9901 PAD.n11490 VSS 0.074902f
C9902 PAD.n11491 VSS 0.074902f
C9903 PAD.n11492 VSS 0.074902f
C9904 PAD.n11493 VSS 0.074902f
C9905 PAD.n11494 VSS 0.074902f
C9906 PAD.n11495 VSS 0.074902f
C9907 PAD.n11496 VSS 0.074902f
C9908 PAD.n11497 VSS 0.074902f
C9909 PAD.n11498 VSS 0.059499f
C9910 PAD.n11499 VSS 0.068257f
C9911 PAD.n11500 VSS 0.700403f
C9912 PAD.n11501 VSS 0.611619f
C9913 PAD.n11502 VSS 0.031988f
C9914 PAD.n11503 VSS 0.031988f
C9915 PAD.n11504 VSS 0.027937f
C9916 PAD.n11505 VSS 0.157796f
C9917 PAD.n11506 VSS 0.123237f
C9918 PAD.n11507 VSS 0.61162f
C9919 PAD.n11508 VSS 0.122923f
C9920 PAD.n11509 VSS 0.61162f
C9921 PAD.n11510 VSS 0.61162f
C9922 PAD.n11512 VSS 0.1262f
C9923 PAD.n11513 VSS 0.61162f
C9924 PAD.n11514 VSS 0.043189f
C9925 PAD.n11515 VSS 0.043189f
C9926 PAD.n11516 VSS 0.05527f
C9927 PAD.n11517 VSS 0.242904f
C9928 PAD.n11518 VSS 0.060756f
C9929 PAD.n11519 VSS 0.062262f
C9930 PAD.n11520 VSS 0.069752f
C9931 PAD.n11521 VSS 0.069752f
C9932 PAD.n11522 VSS 0.700403f
C9933 PAD.n11523 VSS 0.611619f
C9934 PAD.n11524 VSS 0.043746f
C9935 PAD.n11525 VSS 0.043746f
C9936 PAD.n11526 VSS 0.038206f
C9937 PAD.n11527 VSS 0.033766f
C9938 PAD.n11528 VSS 0.026125f
C9939 PAD.n11529 VSS 0.042887f
C9940 PAD.n11530 VSS 0.049106f
C9941 PAD.n11531 VSS 0.049106f
C9942 PAD.n11532 VSS 0.508039f
C9943 PAD.n11533 VSS 0.626417f
C9944 PAD.n11534 VSS 0.685606f
C9945 PAD.n11535 VSS 0.063002f
C9946 PAD.n11536 VSS 0.063002f
C9947 PAD.n11537 VSS 0.034144f
C9948 PAD.n11538 VSS 1.33597f
C9949 PAD.n11539 VSS 16.0728f
C9950 PAD.n11540 VSS 19.3704f
C9951 PAD.n11541 VSS 10.139299f
C9952 PAD.n11542 VSS 0.182422f
C9953 GF_NI_IN_C_BASE_0.comp018green_out_predrv_1.nmos_6p0_CDNS_4066195314519_0.D.t0 VSS 1.57596f
C9954 GF_NI_IN_C_BASE_0.comp018green_out_predrv_1.nmos_6p0_CDNS_4066195314519_0.D.t1 VSS 1.51789f
C9955 GF_NI_IN_C_BASE_0.comp018green_out_predrv_1.nmos_6p0_CDNS_4066195314519_0.D.t2 VSS 1.89864f
C9956 GF_NI_IN_C_BASE_0.comp018green_out_predrv_1.nmos_6p0_CDNS_4066195314519_0.D.t7 VSS 1.25234f
C9957 GF_NI_IN_C_BASE_0.comp018green_out_predrv_1.nmos_6p0_CDNS_4066195314519_0.D.t6 VSS 1.37161f
C9958 GF_NI_IN_C_BASE_0.comp018green_out_predrv_1.nmos_6p0_CDNS_4066195314519_0.D.n0 VSS 0.981389f
C9959 GF_NI_IN_C_BASE_0.comp018green_out_predrv_1.nmos_6p0_CDNS_4066195314519_0.D.t3 VSS 1.25234f
C9960 GF_NI_IN_C_BASE_0.comp018green_out_predrv_1.nmos_6p0_CDNS_4066195314519_0.D.t4 VSS 1.37161f
C9961 GF_NI_IN_C_BASE_0.comp018green_out_predrv_1.nmos_6p0_CDNS_4066195314519_0.D.n1 VSS 0.981389f
C9962 GF_NI_IN_C_BASE_0.comp018green_out_predrv_1.nmos_6p0_CDNS_4066195314519_0.D.n2 VSS 0.25845f
C9963 GF_NI_IN_C_BASE_0.comp018green_out_predrv_1.nmos_6p0_CDNS_4066195314519_0.D.n3 VSS 1.19395f
C9964 GF_NI_IN_C_BASE_0.comp018green_out_predrv_1.nmos_6p0_CDNS_4066195314519_0.D.t5 VSS 0.631878f
C9965 GF_NI_IN_C_BASE_0.comp018green_out_predrv_1.nmos_6p0_CDNS_4066195314519_0.D.t8 VSS 0.727229f
C9966 GF_NI_IN_C_BASE_0.comp018green_out_predrv_1.nmos_6p0_CDNS_4066195314519_0.D.n4 VSS 0.820403f
C9967 GF_NI_IN_C_BASE_0.comp018green_out_predrv_0.A.t0 VSS 0.227858f
C9968 GF_NI_IN_C_BASE_0.comp018green_out_predrv_0.A.t1 VSS 0.789415f
C9969 GF_NI_IN_C_BASE_0.comp018green_out_predrv_0.A.t2 VSS 0.785268f
C9970 GF_NI_IN_C_BASE_0.comp018green_out_predrv_0.A.t8 VSS 1.58711f
C9971 GF_NI_IN_C_BASE_0.comp018green_out_predrv_0.A.t9 VSS 0.785268f
C9972 GF_NI_IN_C_BASE_0.comp018green_out_predrv_0.A.t7 VSS 1.58711f
C9973 GF_NI_IN_C_BASE_0.comp018green_out_predrv_0.A.t6 VSS 0.785268f
C9974 GF_NI_IN_C_BASE_0.comp018green_out_predrv_0.A.t5 VSS 1.58711f
C9975 GF_NI_IN_C_BASE_0.comp018green_out_predrv_0.A.n0 VSS 2.81472f
C9976 GF_NI_IN_C_BASE_0.comp018green_out_predrv_0.A.n1 VSS 2.35462f
C9977 GF_NI_IN_C_BASE_0.comp018green_out_predrv_0.A.n2 VSS 1.65739f
C9978 GF_NI_IN_C_BASE_0.comp018green_out_predrv_0.A.t4 VSS 0.785268f
C9979 GF_NI_IN_C_BASE_0.comp018green_out_predrv_0.A.t3 VSS 1.58711f
C9980 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n0 VSS 0.032995f
C9981 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n1 VSS 0.05081f
C9982 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n2 VSS 0.037555f
C9983 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n3 VSS -1.07192f
C9984 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n4 VSS 1.46073f
C9985 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n5 VSS 0.044183f
C9986 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n6 VSS 0.033137f
C9987 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.t5 VSS 0.162003f
C9988 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n7 VSS 0.044183f
C9989 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n9 VSS 0.05081f
C9990 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n10 VSS 0.02651f
C9991 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n11 VSS 0.037555f
C9992 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n12 VSS 0.05081f
C9993 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n13 VSS 0.033137f
C9994 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n14 VSS 0.05081f
C9995 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n15 VSS 0.02651f
C9996 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n16 VSS 0.037555f
C9997 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n18 VSS 0.243005f
C9998 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n19 VSS 0.388808f
C9999 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n21 VSS 0.05081f
C10000 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n22 VSS 0.05081f
C10001 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n23 VSS 0.033137f
C10002 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.t15 VSS 0.466424f
C10003 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.t10 VSS 0.504368f
C10004 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n24 VSS 0.604239f
C10005 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n25 VSS 0.492247f
C10006 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.t18 VSS 0.205409f
C10007 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n26 VSS 0.496582f
C10008 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n27 VSS 4.56226f
C10009 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.t21 VSS 0.205409f
C10010 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n28 VSS 0.231062f
C10011 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.t16 VSS 0.478595f
C10012 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.t25 VSS 0.288159f
C10013 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n29 VSS 0.507599f
C10014 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n30 VSS 4.40871f
C10015 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n31 VSS 8.20065f
C10016 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.t11 VSS 0.429912f
C10017 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.t23 VSS 0.288159f
C10018 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n32 VSS 0.458907f
C10019 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.t26 VSS 0.205325f
C10020 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n33 VSS 0.08677f
C10021 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n34 VSS 2.82266f
C10022 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.t0 VSS 0.068017f
C10023 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n35 VSS 0.836602f
C10024 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n36 VSS 0.020742f
C10025 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n37 VSS 0.05081f
C10026 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n38 VSS 0.044183f
C10027 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n39 VSS 0.388808f
C10028 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n40 VSS 0.044183f
C10029 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n41 VSS 0.044183f
C10030 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n43 VSS 0.037555f
C10031 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n44 VSS 0.02651f
C10032 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n45 VSS 0.016813f
C10033 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n46 VSS 0.037555f
C10034 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n47 VSS 0.05081f
C10035 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n48 VSS 0.05081f
C10036 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n49 VSS 0.033137f
C10037 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n50 VSS 0.033137f
C10038 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n51 VSS 0.033137f
C10039 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n52 VSS 0.05081f
C10040 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n53 VSS 0.05081f
C10041 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n54 VSS 0.037555f
C10042 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n55 VSS 0.02651f
C10043 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n56 VSS 0.02651f
C10044 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n57 VSS 0.05081f
C10045 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n58 VSS 0.05081f
C10046 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n60 VSS 0.388808f
C10047 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n61 VSS 0.243005f
C10048 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.t2 VSS 0.162003f
C10049 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n62 VSS 0.243005f
C10050 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n63 VSS 0.044183f
C10051 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n64 VSS 0.031197f
C10052 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n65 VSS 0.560119f
C10053 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.t12 VSS 0.466424f
C10054 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.t6 VSS 0.504368f
C10055 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n66 VSS 0.604239f
C10056 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n67 VSS 0.036359f
C10057 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n68 VSS 4.60813f
C10058 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n69 VSS 0.031197f
C10059 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n70 VSS 0.016813f
C10060 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n71 VSS 0.044183f
C10061 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n72 VSS 0.243005f
C10062 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n73 VSS 0.037555f
C10063 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n74 VSS 0.044183f
C10064 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n75 VSS 0.02651f
C10065 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n76 VSS 0.05081f
C10066 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n77 VSS 0.05081f
C10067 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n78 VSS 0.388808f
C10068 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.t1 VSS 0.162003f
C10069 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n79 VSS 0.05081f
C10070 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n82 VSS 0.02651f
C10071 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n83 VSS 0.037555f
C10072 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n84 VSS 0.037555f
C10073 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n85 VSS 0.02651f
C10074 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n86 VSS 0.05081f
C10075 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n87 VSS 0.033137f
C10076 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n88 VSS 0.044183f
C10077 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n89 VSS 0.243005f
C10078 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n90 VSS 0.044183f
C10079 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n91 VSS 0.033137f
C10080 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n92 VSS 0.033137f
C10081 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n93 VSS 0.05081f
C10082 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n94 VSS 0.05081f
C10083 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n95 VSS 0.388808f
C10084 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n96 VSS 0.05081f
C10085 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n97 VSS 0.020742f
C10086 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n98 VSS 0.560119f
C10087 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.t7 VSS 0.466424f
C10088 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.t24 VSS 0.504368f
C10089 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n99 VSS 0.604239f
C10090 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n100 VSS 0.036359f
C10091 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n101 VSS 4.19166f
C10092 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n102 VSS 8.449809f
C10093 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n103 VSS 2.70456f
C10094 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n104 VSS 6.35215f
C10095 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.t14 VSS 0.466424f
C10096 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.t9 VSS 0.504368f
C10097 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n105 VSS 0.604239f
C10098 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n106 VSS 0.419209f
C10099 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n107 VSS 4.81347f
C10100 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n108 VSS 0.025773f
C10101 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n109 VSS 0.032995f
C10102 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n110 VSS 0.044183f
C10103 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n111 VSS 0.388808f
C10104 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n113 VSS 0.033137f
C10105 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n114 VSS 0.044183f
C10106 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n115 VSS 0.388808f
C10107 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n116 VSS 0.05081f
C10108 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n119 VSS 0.033137f
C10109 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n120 VSS 0.05081f
C10110 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n121 VSS 0.05081f
C10111 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n122 VSS 0.02651f
C10112 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n123 VSS 0.037555f
C10113 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n124 VSS 0.037555f
C10114 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n125 VSS 0.02651f
C10115 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n126 VSS 0.05081f
C10116 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n127 VSS 0.033137f
C10117 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n128 VSS 0.044183f
C10118 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n129 VSS 0.243005f
C10119 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.t3 VSS 0.162003f
C10120 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n130 VSS 0.243005f
C10121 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n131 VSS 0.044183f
C10122 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n132 VSS 0.05081f
C10123 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n133 VSS 0.05081f
C10124 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n134 VSS 0.02651f
C10125 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n135 VSS 0.037555f
C10126 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n136 VSS 0.037555f
C10127 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n138 VSS 0.05081f
C10128 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n139 VSS 0.454776f
C10129 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.t20 VSS 0.466424f
C10130 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.t17 VSS 0.504368f
C10131 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n140 VSS 0.604239f
C10132 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n141 VSS 0.060652f
C10133 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n142 VSS 1.49197f
C10134 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n143 VSS 1.34997f
C10135 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n144 VSS 0.025773f
C10136 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n145 VSS 0.032995f
C10137 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n146 VSS 0.044183f
C10138 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n147 VSS 0.388808f
C10139 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n148 VSS 0.02651f
C10140 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n149 VSS 0.044183f
C10141 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n150 VSS 0.05081f
C10142 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n151 VSS 0.05081f
C10143 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n152 VSS 0.243005f
C10144 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.t4 VSS 0.162003f
C10145 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n153 VSS 0.388808f
C10146 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n154 VSS 0.05081f
C10147 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n155 VSS 0.02651f
C10148 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n156 VSS 0.037555f
C10149 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n158 VSS 0.037555f
C10150 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n159 VSS 0.02651f
C10151 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n160 VSS 0.05081f
C10152 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n161 VSS 0.033137f
C10153 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n162 VSS 0.044183f
C10154 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n163 VSS 0.243005f
C10155 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n164 VSS 0.044183f
C10156 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n165 VSS 0.033137f
C10157 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n166 VSS 0.033137f
C10158 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n167 VSS 0.05081f
C10159 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n168 VSS 0.05081f
C10160 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n170 VSS 0.037555f
C10161 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n171 VSS 0.037555f
C10162 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n173 VSS 0.05081f
C10163 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n174 VSS 0.454776f
C10164 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.t13 VSS 0.466424f
C10165 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.t8 VSS 0.504368f
C10166 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n175 VSS 0.604239f
C10167 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n176 VSS 0.060652f
C10168 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n177 VSS 1.49197f
C10169 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n178 VSS 1.59999f
C10170 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.t22 VSS 0.466424f
C10171 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.t19 VSS 0.504368f
C10172 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n179 VSS 0.604239f
C10173 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n180 VSS 0.060652f
C10174 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n181 VSS 1.84223f
C10175 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n182 VSS 0.454776f
C10176 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n183 VSS 0.025773f
C10177 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n184 VSS 0.044183f
C10178 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n185 VSS 0.243005f
C10179 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n186 VSS 0.044183f
C10180 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n187 VSS 0.05081f
C10181 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n189 VSS 0.037555f
C10182 GF_NI_IN_C_BASE_0.comp018green_out_sigbuf_oe_0.OE.n190 VSS 0.02651f
C10183 VDD.n0 VSS 0.125777f
C10184 VDD.n1 VSS 0.139533f
C10185 VDD.n2 VSS 0.071732f
C10186 VDD.n3 VSS 0.039867f
C10187 VDD.n4 VSS 0.039867f
C10188 VDD.n5 VSS 0.039867f
C10189 VDD.n6 VSS 0.039867f
C10190 VDD.n8 VSS 0.069767f
C10191 VDD.n9 VSS 0.129216f
C10192 VDD.n10 VSS 0.039867f
C10193 VDD.n11 VSS 0.039867f
C10194 VDD.n12 VSS 0.039867f
C10195 VDD.n13 VSS 0.039867f
C10196 VDD.n15 VSS 0.043102f
C10197 VDD.n16 VSS 0.03873f
C10198 VDD.n18 VSS 0.070005f
C10199 VDD.n19 VSS 0.042854f
C10200 VDD.n20 VSS 0.074179f
C10201 VDD.n21 VSS 2.48e-19
C10202 VDD.n22 VSS 0.355018f
C10203 VDD.t38 VSS 0.162335f
C10204 VDD.n23 VSS 0.162633f
C10205 VDD.n24 VSS 0.029672f
C10206 VDD.n25 VSS 0.004952f
C10207 VDD.n26 VSS 0.005862f
C10208 VDD.n27 VSS 0.152689f
C10209 VDD.n28 VSS 0.006772f
C10210 VDD.n29 VSS 0.173093f
C10211 VDD.n30 VSS 0.003011f
C10212 VDD.n32 VSS 0.005862f
C10213 VDD.n33 VSS 0.484412f
C10214 VDD.n35 VSS 0.003761f
C10215 VDD.n37 VSS 0.006772f
C10216 VDD.n38 VSS 0.087635f
C10217 VDD.n39 VSS 0.004952f
C10218 VDD.n40 VSS 0.036231f
C10219 VDD.n42 VSS 0.005862f
C10220 VDD.t58 VSS 0.124732f
C10221 VDD.n43 VSS 0.005862f
C10222 VDD.n44 VSS 0.005862f
C10223 VDD.n45 VSS 0.005862f
C10224 VDD.n46 VSS 0.005862f
C10225 VDD.n47 VSS 0.010815f
C10226 VDD.n48 VSS 0.005862f
C10227 VDD.n49 VSS 0.006772f
C10228 VDD.n50 VSS 0.152689f
C10229 VDD.n51 VSS 0.005862f
C10230 VDD.n52 VSS 0.005862f
C10231 VDD.n53 VSS 0.006772f
C10232 VDD.n55 VSS 0.004952f
C10233 VDD.n56 VSS 0.004952f
C10234 VDD.n57 VSS 0.004952f
C10235 VDD.n58 VSS 0.004952f
C10236 VDD.n60 VSS 0.006772f
C10237 VDD.n62 VSS 0.005862f
C10238 VDD.n63 VSS 0.006772f
C10239 VDD.n64 VSS 0.003761f
C10240 VDD.n65 VSS 0.003011f
C10241 VDD.n66 VSS 0.005862f
C10242 VDD.n67 VSS 0.004952f
C10243 VDD.n68 VSS 0.005862f
C10244 VDD.n69 VSS 0.003011f
C10245 VDD.n70 VSS 0.003761f
C10246 VDD.n71 VSS 0.004952f
C10247 VDD.n72 VSS 0.004952f
C10248 VDD.n73 VSS 0.010815f
C10249 VDD.n74 VSS 0.004952f
C10250 VDD.n75 VSS 0.004952f
C10251 VDD.n76 VSS 0.005862f
C10252 VDD.n78 VSS 0.004952f
C10253 VDD.n79 VSS 0.004952f
C10254 VDD.n80 VSS 0.016013f
C10255 VDD.t60 VSS 0.040445f
C10256 VDD.n81 VSS 0.052887f
C10257 VDD.n82 VSS 0.39691f
C10258 VDD.t19 VSS 0.029564f
C10259 VDD.n83 VSS 0.070046f
C10260 VDD.n84 VSS 0.062922f
C10261 VDD.t21 VSS 0.029564f
C10262 VDD.n85 VSS 0.070046f
C10263 VDD.n86 VSS 0.021904f
C10264 VDD.n87 VSS 0.036602f
C10265 VDD.t18 VSS 0.245152f
C10266 VDD.n88 VSS 0.070688f
C10267 VDD.n89 VSS 0.0196f
C10268 VDD.n90 VSS 0.019494f
C10269 VDD.n91 VSS 0.019409f
C10270 VDD.n92 VSS 0.021904f
C10271 VDD.n93 VSS 0.036602f
C10272 VDD.n94 VSS 0.035027f
C10273 VDD.n95 VSS 0.045956f
C10274 VDD.n96 VSS 0.309707f
C10275 VDD.t20 VSS 0.245152f
C10276 VDD.n97 VSS 0.070688f
C10277 VDD.n98 VSS 0.39691f
C10278 VDD.n99 VSS 0.021504f
C10279 VDD.n100 VSS 0.051601f
C10280 VDD.t62 VSS 0.041336f
C10281 VDD.n101 VSS 0.055147f
C10282 VDD.n102 VSS 0.032271f
C10283 VDD.n103 VSS 0.345838f
C10284 VDD.t61 VSS 0.24574f
C10285 VDD.n104 VSS 0.070688f
C10286 VDD.n105 VSS 0.503243f
C10287 VDD.n106 VSS 0.176187f
C10288 VDD.n107 VSS 0.050235f
C10289 VDD.n108 VSS 0.042804f
C10290 VDD.n109 VSS 0.050022f
C10291 VDD.n110 VSS 0.17597f
C10292 VDD.n111 VSS 0.531549f
C10293 VDD.t59 VSS 0.253741f
C10294 VDD.n112 VSS 0.118594f
C10295 VDD.n113 VSS 0.397014f
C10296 VDD.n114 VSS 0.197062f
C10297 VDD.n115 VSS 0.036231f
C10298 VDD.n116 VSS 0.005862f
C10299 VDD.n117 VSS 0.124732f
C10300 VDD.n118 VSS 0.005862f
C10301 VDD.n119 VSS 0.005862f
C10302 VDD.n120 VSS 0.005862f
C10303 VDD.n121 VSS 0.006772f
C10304 VDD.n122 VSS 0.006772f
C10305 VDD.n124 VSS 0.004952f
C10306 VDD.n125 VSS 0.004952f
C10307 VDD.n126 VSS 0.004952f
C10308 VDD.n127 VSS 0.004952f
C10309 VDD.n128 VSS 0.003761f
C10310 VDD.n129 VSS 0.003011f
C10311 VDD.n130 VSS 0.005862f
C10312 VDD.n131 VSS 0.124732f
C10313 VDD.n132 VSS 0.005862f
C10314 VDD.n133 VSS 0.006772f
C10315 VDD.n134 VSS 0.112966f
C10316 VDD.n135 VSS 0.110135f
C10317 VDD.n136 VSS 0.034588f
C10318 VDD.n137 VSS 0.224637f
C10319 VDD.n138 VSS 0.106469f
C10320 VDD.n139 VSS 0.005862f
C10321 VDD.n140 VSS 0.005862f
C10322 VDD.n141 VSS 0.005862f
C10323 VDD.n142 VSS 0.005862f
C10324 VDD.n145 VSS 0.004952f
C10325 VDD.n146 VSS 0.004952f
C10326 VDD.n147 VSS 0.006772f
C10327 VDD.n148 VSS 0.005862f
C10328 VDD.n149 VSS 0.005862f
C10329 VDD.n150 VSS 0.005862f
C10330 VDD.n151 VSS 0.006772f
C10331 VDD.n152 VSS 0.006772f
C10332 VDD.n153 VSS 0.004952f
C10333 VDD.n154 VSS 0.004952f
C10334 VDD.n155 VSS 0.005862f
C10335 VDD.n156 VSS 0.004952f
C10336 VDD.n157 VSS 0.005862f
C10337 VDD.n158 VSS 0.007403f
C10338 VDD.n159 VSS 0.006772f
C10339 VDD.n160 VSS 0.005862f
C10340 VDD.n161 VSS 0.124732f
C10341 VDD.n162 VSS 0.003011f
C10342 VDD.n163 VSS 0.005862f
C10343 VDD.n164 VSS 0.005862f
C10344 VDD.n166 VSS 0.005862f
C10345 VDD.t0 VSS 0.099463f
C10346 VDD.n167 VSS 0.005862f
C10347 VDD.n168 VSS 0.036231f
C10348 VDD.n169 VSS 0.005862f
C10349 VDD.n170 VSS 0.005467f
C10350 VDD.n171 VSS 0.004952f
C10351 VDD.n172 VSS 0.005862f
C10352 VDD.n173 VSS 0.004952f
C10353 VDD.n174 VSS 0.004952f
C10354 VDD.n175 VSS 0.006772f
C10355 VDD.n176 VSS 0.484412f
C10356 VDD.n177 VSS 0.003761f
C10357 VDD.n178 VSS 0.004952f
C10358 VDD.n179 VSS 0.005467f
C10359 VDD.n180 VSS 0.168621f
C10360 VDD.n181 VSS 0.008439f
C10361 VDD.n182 VSS 0.005862f
C10362 VDD.n183 VSS 0.004952f
C10363 VDD.n185 VSS 0.005862f
C10364 VDD.n186 VSS 0.004952f
C10365 VDD.n188 VSS 0.006772f
C10366 VDD.n189 VSS 0.078699f
C10367 VDD.n190 VSS 0.018115f
C10368 VDD.n191 VSS 0.055768f
C10369 VDD.n192 VSS 0.175498f
C10370 VDD.t22 VSS 0.179788f
C10371 VDD.n193 VSS 0.401155f
C10372 VDD.t23 VSS 0.009336f
C10373 VDD.n194 VSS 0.364823f
C10374 VDD.n195 VSS 0.024949f
C10375 VDD.n196 VSS 0.045482f
C10376 VDD.n197 VSS 0.034669f
C10377 VDD.n198 VSS 0.034813f
C10378 VDD.n200 VSS 0.110195f
C10379 VDD.n201 VSS 0.110195f
C10380 VDD.n202 VSS 0.083862f
C10381 VDD.n203 VSS 0.034813f
C10382 VDD.n205 VSS 0.435726f
C10383 VDD.n206 VSS 0.438253f
C10384 VDD.n207 VSS 0.069767f
C10385 VDD.n209 VSS 0.039867f
C10386 VDD.n211 VSS 0.039867f
C10387 VDD.n213 VSS 0.039867f
C10388 VDD.n214 VSS 0.069767f
C10389 VDD.n218 VSS 0.139533f
C10390 VDD.n219 VSS 0.137568f
C10391 VDD.n220 VSS 0.015722f
C10392 VDD.n221 VSS 0.139533f
C10393 VDD.n222 VSS 0.139533f
C10394 VDD.n223 VSS 0.139533f
C10395 VDD.n224 VSS 0.139533f
C10396 VDD.n225 VSS 0.139533f
C10397 VDD.n226 VSS 0.139533f
C10398 VDD.n227 VSS 0.139533f
C10399 VDD.n228 VSS 0.139533f
C10400 VDD.n229 VSS 0.139533f
C10401 VDD.n230 VSS 0.139533f
C10402 VDD.n231 VSS 0.139533f
C10403 VDD.n232 VSS 0.139533f
C10404 VDD.n233 VSS 0.139533f
C10405 VDD.n234 VSS 0.139533f
C10406 VDD.n235 VSS 0.139533f
C10407 VDD.n236 VSS 0.139533f
C10408 VDD.n237 VSS 0.139533f
C10409 VDD.n238 VSS 0.139533f
C10410 VDD.n239 VSS 0.139533f
C10411 VDD.n240 VSS 0.139533f
C10412 VDD.n241 VSS 0.139533f
C10413 VDD.n242 VSS 0.139533f
C10414 VDD.n243 VSS 0.139533f
C10415 VDD.n244 VSS 0.139533f
C10416 VDD.n245 VSS 0.139533f
C10417 VDD.n246 VSS 0.139533f
C10418 VDD.n247 VSS 0.139533f
C10419 VDD.n248 VSS 0.139533f
C10420 VDD.n249 VSS 0.139533f
C10421 VDD.n250 VSS 0.139533f
C10422 VDD.n251 VSS 0.139533f
C10423 VDD.n252 VSS 0.139533f
C10424 VDD.n253 VSS 0.139533f
C10425 VDD.n254 VSS 0.139533f
C10426 VDD.n255 VSS 0.139533f
C10427 VDD.n256 VSS 0.139533f
C10428 VDD.n257 VSS 0.139533f
C10429 VDD.n258 VSS 0.139533f
C10430 VDD.n259 VSS 0.139533f
C10431 VDD.n260 VSS 0.139533f
C10432 VDD.n261 VSS 0.139533f
C10433 VDD.n262 VSS 0.139533f
C10434 VDD.n263 VSS 0.139533f
C10435 VDD.n264 VSS 0.139533f
C10436 VDD.n265 VSS 0.139533f
C10437 VDD.n266 VSS 0.139533f
C10438 VDD.n267 VSS 0.139533f
C10439 VDD.n268 VSS 0.139533f
C10440 VDD.n269 VSS 0.139533f
C10441 VDD.n270 VSS 0.139533f
C10442 VDD.n271 VSS 0.139533f
C10443 VDD.n272 VSS 0.139533f
C10444 VDD.n273 VSS 0.139533f
C10445 VDD.n274 VSS 0.139533f
C10446 VDD.n275 VSS 0.139533f
C10447 VDD.n276 VSS 0.139533f
C10448 VDD.n277 VSS 0.139533f
C10449 VDD.n278 VSS 0.139533f
C10450 VDD.n279 VSS 0.139533f
C10451 VDD.n280 VSS 0.139533f
C10452 VDD.n281 VSS 0.139533f
C10453 VDD.n282 VSS 0.139533f
C10454 VDD.n283 VSS 0.139533f
C10455 VDD.n284 VSS 0.139533f
C10456 VDD.n285 VSS 0.139533f
C10457 VDD.n286 VSS 0.139533f
C10458 VDD.n287 VSS 0.139533f
C10459 VDD.n288 VSS 0.139533f
C10460 VDD.n289 VSS 0.139533f
C10461 VDD.n290 VSS 0.139533f
C10462 VDD.n291 VSS 0.139533f
C10463 VDD.n292 VSS 0.139533f
C10464 VDD.n293 VSS 0.118898f
C10465 VDD.t29 VSS 0.034261f
C10466 VDD.n294 VSS 0.072876f
C10467 VDD.t42 VSS 0.192545f
C10468 VDD.n295 VSS 0.825895f
C10469 VDD.n296 VSS 0.139533f
C10470 VDD.n297 VSS 0.139533f
C10471 VDD.n298 VSS 0.139533f
C10472 VDD.n299 VSS 0.139533f
C10473 VDD.n300 VSS 0.139533f
C10474 VDD.n301 VSS 0.139533f
C10475 VDD.n302 VSS 0.139533f
C10476 VDD.n303 VSS 0.139533f
C10477 VDD.n304 VSS 0.139533f
C10478 VDD.n305 VSS 0.139533f
C10479 VDD.n306 VSS 0.139533f
C10480 VDD.n307 VSS 0.139533f
C10481 VDD.n308 VSS 0.139533f
C10482 VDD.n309 VSS 0.139533f
C10483 VDD.n310 VSS 0.139533f
C10484 VDD.n311 VSS 0.139533f
C10485 VDD.n312 VSS 0.139533f
C10486 VDD.t41 VSS 0.037778f
C10487 VDD.n313 VSS 0.053288f
C10488 VDD.t55 VSS 0.219338f
C10489 VDD.t63 VSS 0.396283f
C10490 VDD.t56 VSS 0.03689f
C10491 VDD.n314 VSS 0.056722f
C10492 VDD.n315 VSS 0.010533f
C10493 VDD.n316 VSS 0.295985f
C10494 VDD.t54 VSS 0.03689f
C10495 VDD.n317 VSS -0.011443f
C10496 VDD.t65 VSS 0.291088f
C10497 VDD.n318 VSS 0.12669f
C10498 VDD.t57 VSS 0.275648f
C10499 VDD.t36 VSS 0.411712f
C10500 VDD.t37 VSS 0.041328f
C10501 VDD.n319 VSS 0.057501f
C10502 VDD.t35 VSS 0.03689f
C10503 VDD.n320 VSS 0.119987f
C10504 VDD.n321 VSS 0.284723f
C10505 VDD.t34 VSS 0.220861f
C10506 VDD.t53 VSS 0.219338f
C10507 VDD.n322 VSS 0.087179f
C10508 VDD.n323 VSS 0.043801f
C10509 VDD.n324 VSS 0.131433f
C10510 VDD.n325 VSS 0.049873f
C10511 VDD.n326 VSS 0.029375f
C10512 VDD.n327 VSS 0.027262f
C10513 VDD.t64 VSS 0.040443f
C10514 VDD.n328 VSS 0.062296f
C10515 VDD.n329 VSS 0.030591f
C10516 VDD.n330 VSS 0.010533f
C10517 VDD.n331 VSS 0.018241f
C10518 VDD.n332 VSS 0.327126f
C10519 VDD.n333 VSS -0.014963f
C10520 VDD.n334 VSS 0.087179f
C10521 VDD.t40 VSS 0.22094f
C10522 VDD.n335 VSS 0.437333f
C10523 VDD.n336 VSS 0.225011f
C10524 VDD.n337 VSS 0.070087f
C10525 VDD.n338 VSS 0.139533f
C10526 VDD.n339 VSS 0.139533f
C10527 VDD.n340 VSS 0.139533f
C10528 VDD.n341 VSS 0.084997f
C10529 VDD.n342 VSS 0.139533f
C10530 VDD.n343 VSS 0.139533f
C10531 VDD.n344 VSS 0.139533f
C10532 VDD.n345 VSS 0.139533f
C10533 VDD.n346 VSS 0.139533f
C10534 VDD.n347 VSS 0.139533f
C10535 VDD.n348 VSS 0.139533f
C10536 VDD.n349 VSS 0.139533f
C10537 VDD.n350 VSS 0.139533f
C10538 VDD.n351 VSS 0.139533f
C10539 VDD.n352 VSS 0.055027f
C10540 VDD.n353 VSS 0.070084f
C10541 VDD.n354 VSS 0.139042f
C10542 VDD.n355 VSS 0.139533f
C10543 VDD.n356 VSS 0.139533f
C10544 VDD.n357 VSS 0.139533f
C10545 VDD.n358 VSS 0.139533f
C10546 VDD.n359 VSS 0.139533f
C10547 VDD.n360 VSS 0.139533f
C10548 VDD.n361 VSS 0.139533f
C10549 VDD.n362 VSS 0.139533f
C10550 VDD.n363 VSS 0.139533f
C10551 VDD.n364 VSS 0.139533f
C10552 VDD.n365 VSS 0.139533f
C10553 VDD.n366 VSS 0.139533f
C10554 VDD.n367 VSS 0.139533f
C10555 VDD.n368 VSS 0.139533f
C10556 VDD.n369 VSS 0.139533f
C10557 VDD.n370 VSS 0.139533f
C10558 VDD.n371 VSS 0.139533f
C10559 VDD.n372 VSS 0.139533f
C10560 VDD.n373 VSS 0.139533f
C10561 VDD.n374 VSS 0.139533f
C10562 VDD.n375 VSS 0.139533f
C10563 VDD.n376 VSS 0.139533f
C10564 VDD.n377 VSS 0.139533f
C10565 VDD.n378 VSS 0.139533f
C10566 VDD.n379 VSS 0.139533f
C10567 VDD.n380 VSS 0.139533f
C10568 VDD.n381 VSS 0.139533f
C10569 VDD.n382 VSS 0.139533f
C10570 VDD.n383 VSS 0.966293f
C10571 VDD.n384 VSS 0.139533f
C10572 VDD.n385 VSS 0.270218f
C10573 VDD.n386 VSS 0.131181f
C10574 VDD.n387 VSS 0.806792f
C10575 VDD.t46 VSS 0.221608f
C10576 VDD.t30 VSS 0.221608f
C10577 VDD.t48 VSS 0.221608f
C10578 VDD.t32 VSS 0.296319f
C10579 VDD.n388 VSS 0.403675f
C10580 VDD.t33 VSS 0.046165f
C10581 VDD.n389 VSS 0.073267f
C10582 VDD.t49 VSS 0.012774f
C10583 VDD.t31 VSS 0.012774f
C10584 VDD.n390 VSS 0.042223f
C10585 VDD.n391 VSS 0.054145f
C10586 VDD.t47 VSS 0.012774f
C10587 VDD.t43 VSS 0.012774f
C10588 VDD.n392 VSS 0.042223f
C10589 VDD.n393 VSS 0.048394f
C10590 VDD.t45 VSS 0.046165f
C10591 VDD.t25 VSS 0.034261f
C10592 VDD.t27 VSS 0.009124f
C10593 VDD.t67 VSS 0.009124f
C10594 VDD.n394 VSS 0.032191f
C10595 VDD.n395 VSS 0.055197f
C10596 VDD.n396 VSS 0.0599f
C10597 VDD.n397 VSS 0.054049f
C10598 VDD.n398 VSS -0.08616f
C10599 VDD.n399 VSS 0.018893f
C10600 VDD.t44 VSS 0.217975f
C10601 VDD.t24 VSS 0.299716f
C10602 VDD.t26 VSS 0.221608f
C10603 VDD.t66 VSS 0.221608f
C10604 VDD.t28 VSS 0.257177f
C10605 VDD.n400 VSS 0.226166f
C10606 VDD.n401 VSS 0.082955f
C10607 VDD.n402 VSS 0.090402f
C10608 VDD.n403 VSS 0.139533f
C10609 VDD.n404 VSS 0.139533f
C10610 VDD.n405 VSS 0.139533f
C10611 VDD.n406 VSS 0.139533f
C10612 VDD.n407 VSS 0.139533f
C10613 VDD.n408 VSS 0.139533f
C10614 VDD.n409 VSS 0.139533f
C10615 VDD.n410 VSS 0.139533f
C10616 VDD.n411 VSS 0.139533f
C10617 VDD.n412 VSS 0.139533f
C10618 VDD.n413 VSS 0.139533f
C10619 VDD.n414 VSS 0.139533f
C10620 VDD.n415 VSS 0.139533f
C10621 VDD.n416 VSS 0.139533f
C10622 VDD.n417 VSS 0.139533f
C10623 VDD.n418 VSS 0.139533f
C10624 VDD.n419 VSS 0.139533f
C10625 VDD.n420 VSS 0.139533f
C10626 VDD.n421 VSS 0.139533f
C10627 VDD.n422 VSS 0.139533f
C10628 VDD.n423 VSS 0.139533f
C10629 VDD.n424 VSS 0.139533f
C10630 VDD.n425 VSS 0.139533f
C10631 VDD.n426 VSS 0.139533f
C10632 VDD.n427 VSS 0.139533f
C10633 VDD.n428 VSS 0.139533f
C10634 VDD.n429 VSS 0.139533f
C10635 VDD.n430 VSS 0.139533f
C10636 VDD.n431 VSS 0.139533f
C10637 VDD.n432 VSS 0.139533f
C10638 VDD.n433 VSS 0.139533f
C10639 VDD.n434 VSS 0.139533f
C10640 VDD.n435 VSS 0.139533f
C10641 VDD.n436 VSS 0.139533f
C10642 VDD.n437 VSS 0.139533f
C10643 VDD.n438 VSS 0.139533f
C10644 VDD.n439 VSS 0.139533f
C10645 VDD.n440 VSS 0.139533f
C10646 VDD.n441 VSS 0.139533f
C10647 VDD.n442 VSS 0.139533f
C10648 VDD.n443 VSS 0.139533f
C10649 VDD.n444 VSS 0.139533f
C10650 VDD.n445 VSS 0.139533f
C10651 VDD.n446 VSS 0.139533f
C10652 VDD.n447 VSS 0.139533f
C10653 VDD.n448 VSS 0.139533f
C10654 VDD.n449 VSS 0.139533f
C10655 VDD.n450 VSS 0.139533f
C10656 VDD.n451 VSS 0.139533f
C10657 VDD.n452 VSS 0.139533f
C10658 VDD.n453 VSS 0.139533f
C10659 VDD.n454 VSS 0.139533f
C10660 VDD.n455 VSS 0.139533f
C10661 VDD.n456 VSS 0.139533f
C10662 VDD.n457 VSS 0.139533f
C10663 VDD.n458 VSS 0.139533f
C10664 VDD.n459 VSS 0.139533f
C10665 VDD.n460 VSS 0.139533f
C10666 VDD.n461 VSS 0.139533f
C10667 VDD.n462 VSS 0.139533f
C10668 VDD.n463 VSS 0.139533f
C10669 VDD.n464 VSS 0.139533f
C10670 VDD.n465 VSS 0.139533f
C10671 VDD.n466 VSS 0.139533f
C10672 VDD.n467 VSS 0.139533f
C10673 VDD.n468 VSS 0.139533f
C10674 VDD.n469 VSS 0.139533f
C10675 VDD.n470 VSS 0.139533f
C10676 VDD.n471 VSS 0.139533f
C10677 VDD.n472 VSS 0.139533f
C10678 VDD.n473 VSS 0.139533f
C10679 VDD.n474 VSS 0.139533f
C10680 VDD.n475 VSS 0.139533f
C10681 VDD.n476 VSS 0.139533f
C10682 VDD.n477 VSS 0.139533f
C10683 VDD.n478 VSS 0.139533f
C10684 VDD.n479 VSS 0.139533f
C10685 VDD.n480 VSS 0.139533f
C10686 VDD.n481 VSS 0.139533f
C10687 VDD.n482 VSS 0.139533f
C10688 VDD.n483 VSS 0.139533f
C10689 VDD.n484 VSS 0.139533f
C10690 VDD.n485 VSS 0.139533f
C10691 VDD.n486 VSS 0.139533f
C10692 VDD.n487 VSS 0.139533f
C10693 VDD.n488 VSS 0.139533f
C10694 VDD.n489 VSS 0.139533f
C10695 VDD.n490 VSS 0.139533f
C10696 VDD.n491 VSS 0.139533f
C10697 VDD.n492 VSS 0.139533f
C10698 VDD.n493 VSS 0.139533f
C10699 VDD.n494 VSS 0.139533f
C10700 VDD.n495 VSS 0.139533f
C10701 VDD.n496 VSS 0.139533f
C10702 VDD.n497 VSS 0.139533f
C10703 VDD.n498 VSS 0.139533f
C10704 VDD.n499 VSS 0.139533f
C10705 VDD.n500 VSS 0.139533f
C10706 VDD.n501 VSS 0.139533f
C10707 VDD.n502 VSS 0.139533f
C10708 VDD.n503 VSS 0.139533f
C10709 VDD.n504 VSS 0.139533f
C10710 VDD.n505 VSS 0.139533f
C10711 VDD.n506 VSS 0.139533f
C10712 VDD.n507 VSS 0.139533f
C10713 VDD.n508 VSS 0.139533f
C10714 VDD.n509 VSS 0.139533f
C10715 VDD.n510 VSS 0.139533f
C10716 VDD.n511 VSS 0.139533f
C10717 VDD.n512 VSS 0.139533f
C10718 VDD.n513 VSS 0.139533f
C10719 VDD.n514 VSS 0.139533f
C10720 VDD.n515 VSS 0.139533f
C10721 VDD.n516 VSS 0.139533f
C10722 VDD.n517 VSS 0.139533f
C10723 VDD.n518 VSS 0.139533f
C10724 VDD.n519 VSS 0.139533f
C10725 VDD.n520 VSS 0.139533f
C10726 VDD.n521 VSS 0.139533f
C10727 VDD.n522 VSS 0.139533f
C10728 VDD.n523 VSS 0.139533f
C10729 VDD.n524 VSS 0.139533f
C10730 VDD.n525 VSS 0.139533f
C10731 VDD.n526 VSS 0.139533f
C10732 VDD.n527 VSS 0.139533f
C10733 VDD.n528 VSS 0.139533f
C10734 VDD.n529 VSS 0.139533f
C10735 VDD.n530 VSS 0.139533f
C10736 VDD.n531 VSS 0.139533f
C10737 VDD.n532 VSS 0.139533f
C10738 VDD.n533 VSS 0.139533f
C10739 VDD.n534 VSS 0.139533f
C10740 VDD.n535 VSS 0.139533f
C10741 VDD.n536 VSS 0.139533f
C10742 VDD.n537 VSS 0.139533f
C10743 VDD.n538 VSS 0.139533f
C10744 VDD.n539 VSS 0.139533f
C10745 VDD.n540 VSS 0.139533f
C10746 VDD.n541 VSS 0.139533f
C10747 VDD.n542 VSS 0.125777f
C10748 VDD.n543 VSS 0.125777f
C10749 VDD.n544 VSS 0.125777f
C10750 VDD.n545 VSS 0.083523f
C10751 VDD.n546 VSS 0.083523f
C10752 VDD.n547 VSS 0.139533f
C10753 VDD.n548 VSS 0.139533f
C10754 VDD.n549 VSS 0.520817f
C10755 VDD.n550 VSS 0.266933f
C10756 VDD.n551 VSS 0.268086f
C10757 VDD.n554 VSS 0.039867f
C10758 VDD.n555 VSS 0.069767f
C10759 VDD.n556 VSS 1.33581f
C10760 VDD.t16 VSS 0.290299f
C10761 VDD.t17 VSS 0.037778f
C10762 VDD.t2 VSS 0.037778f
C10763 VDD.n557 VSS 0.071818f
C10764 VDD.n558 VSS 0.126759f
C10765 VDD.n559 VSS 0.139533f
C10766 VDD.n560 VSS 0.139533f
C10767 VDD.n561 VSS 0.139533f
C10768 VDD.n562 VSS 0.139533f
C10769 VDD.n563 VSS 0.139533f
C10770 VDD.n564 VSS 0.139533f
C10771 VDD.n565 VSS 0.139533f
C10772 VDD.n566 VSS 0.139533f
C10773 VDD.n567 VSS 0.139533f
C10774 VDD.n568 VSS 0.139533f
C10775 VDD.n569 VSS 0.139533f
C10776 VDD.n570 VSS 0.139533f
C10777 VDD.n571 VSS 0.139533f
C10778 VDD.n572 VSS 0.139533f
C10779 VDD.n573 VSS 0.139533f
C10780 VDD.n574 VSS 0.139533f
C10781 VDD.n575 VSS 0.139533f
C10782 VDD.n576 VSS 0.139533f
C10783 VDD.n577 VSS 0.139533f
C10784 VDD.n578 VSS 0.139533f
C10785 VDD.n579 VSS 0.139533f
C10786 VDD.n580 VSS 0.139533f
C10787 VDD.n581 VSS 0.139533f
C10788 VDD.n582 VSS 0.139533f
C10789 VDD.n583 VSS 0.139533f
C10790 VDD.n584 VSS 0.104159f
C10791 VDD.t13 VSS 0.037778f
C10792 VDD.n585 VSS 0.071823f
C10793 VDD.t14 VSS 0.287817f
C10794 VDD.n586 VSS 0.114164f
C10795 VDD.t3 VSS 0.289019f
C10796 VDD.n587 VSS 0.131672f
C10797 VDD.n588 VSS 0.139533f
C10798 VDD.n589 VSS 0.139533f
C10799 VDD.n590 VSS 0.139533f
C10800 VDD.n591 VSS 0.139533f
C10801 VDD.n592 VSS 0.139533f
C10802 VDD.n593 VSS 0.139533f
C10803 VDD.n594 VSS 0.139533f
C10804 VDD.n595 VSS 0.139533f
C10805 VDD.n596 VSS 0.139533f
C10806 VDD.n597 VSS 0.139533f
C10807 VDD.n598 VSS 0.139533f
C10808 VDD.n599 VSS 0.139533f
C10809 VDD.n600 VSS 0.139533f
C10810 VDD.n601 VSS 0.139533f
C10811 VDD.n602 VSS 0.139533f
C10812 VDD.n603 VSS 0.139533f
C10813 VDD.n604 VSS 0.139533f
C10814 VDD.n605 VSS 0.139533f
C10815 VDD.n606 VSS 0.139533f
C10816 VDD.n607 VSS 0.139533f
C10817 VDD.n608 VSS 0.139533f
C10818 VDD.n609 VSS 0.139533f
C10819 VDD.n610 VSS 0.139533f
C10820 VDD.n611 VSS 0.139533f
C10821 VDD.n612 VSS 0.139533f
C10822 VDD.n613 VSS 0.109072f
C10823 VDD.t9 VSS 0.037778f
C10824 VDD.n614 VSS 0.070746f
C10825 VDD.t10 VSS 0.25981f
C10826 VDD.n615 VSS 0.004683f
C10827 VDD.n616 VSS 0.004952f
C10828 VDD.n617 VSS 0.005862f
C10829 VDD.n618 VSS 0.004952f
C10830 VDD.n619 VSS 0.089234f
C10831 VDD.n622 VSS 0.005862f
C10832 VDD.n623 VSS 0.004952f
C10833 VDD.n624 VSS 0.005862f
C10834 VDD.n625 VSS 0.004952f
C10835 VDD.n626 VSS 0.005862f
C10836 VDD.n627 VSS 0.005862f
C10837 VDD.n628 VSS 0.089234f
C10838 VDD.n629 VSS 0.005862f
C10839 VDD.n630 VSS 0.005862f
C10840 VDD.n631 VSS 0.005862f
C10841 VDD.n632 VSS 0.004952f
C10842 VDD.n633 VSS 0.004952f
C10843 VDD.n634 VSS 0.004952f
C10844 VDD.n635 VSS 0.004952f
C10845 VDD.n637 VSS 0.004952f
C10846 VDD.n638 VSS 0.005862f
C10847 VDD.n639 VSS 0.005862f
C10848 VDD.n640 VSS 0.004952f
C10849 VDD.n641 VSS 0.005862f
C10850 VDD.n642 VSS 0.006772f
C10851 VDD.n643 VSS 0.006772f
C10852 VDD.n645 VSS 0.005862f
C10853 VDD.n646 VSS 0.004952f
C10854 VDD.n647 VSS 0.004952f
C10855 VDD.n648 VSS 0.006772f
C10856 VDD.n649 VSS 0.006772f
C10857 VDD.n651 VSS 0.109235f
C10858 VDD.n653 VSS 0.008793f
C10859 VDD.n654 VSS 0.008793f
C10860 VDD.n655 VSS 0.005862f
C10861 VDD.n656 VSS 0.004952f
C10862 VDD.n657 VSS 0.004952f
C10863 VDD.n658 VSS 0.008793f
C10864 VDD.n659 VSS 0.005862f
C10865 VDD.n660 VSS 0.004952f
C10866 VDD.n661 VSS 0.004952f
C10867 VDD.n662 VSS 0.008793f
C10868 VDD.n663 VSS 0.005862f
C10869 VDD.n664 VSS 0.005862f
C10870 VDD.t5 VSS 0.089234f
C10871 VDD.n665 VSS 0.005862f
C10872 VDD.n666 VSS 0.005862f
C10873 VDD.n667 VSS 0.006772f
C10874 VDD.n668 VSS 0.006772f
C10875 VDD.n670 VSS 0.109235f
C10876 VDD.n672 VSS 0.006772f
C10877 VDD.n673 VSS 0.005382f
C10878 VDD.n674 VSS 0.03087f
C10879 VDD.n675 VSS 5.18407f
C10880 VDD.n676 VSS 0.139533f
C10881 VDD.n677 VSS 0.139533f
C10882 VDD.n678 VSS 0.139533f
C10883 VDD.n679 VSS 0.139533f
C10884 VDD.n680 VSS 0.139533f
C10885 VDD.n681 VSS 0.139533f
C10886 VDD.n682 VSS 0.139533f
C10887 VDD.n683 VSS 0.139533f
C10888 VDD.n684 VSS 0.139533f
C10889 VDD.n685 VSS 0.139533f
C10890 VDD.n686 VSS 0.139533f
C10891 VDD.n687 VSS 0.139533f
C10892 VDD.n688 VSS 3.19519f
C10893 VDD.n689 VSS 0.139533f
C10894 VDD.n690 VSS 0.472462f
C10895 VDD.n691 VSS 0.110546f
C10896 VDD.n692 VSS 2.82128f
C10897 VDD.n693 VSS 0.116991f
C10898 VDD.n694 VSS 0.052009f
C10899 VDD.t7 VSS 0.046586f
C10900 VDD.n695 VSS 0.080002f
C10901 VDD.n696 VSS 0.389119f
C10902 VDD.t6 VSS 0.412229f
C10903 VDD.n697 VSS 0.098332f
C10904 VDD.n698 VSS 0.059682f
C10905 VDD.n699 VSS 0.021281f
C10906 VDD.t11 VSS 0.037778f
C10907 VDD.n700 VSS 0.052572f
C10908 VDD.n701 VSS -0.010824f
C10909 VDD.n702 VSS 0.124742f
C10910 VDD.t8 VSS 0.261045f
C10911 VDD.n703 VSS 0.324035f
C10912 VDD.n704 VSS 0.113645f
C10913 VDD.n705 VSS 0.100228f
C10914 VDD.n706 VSS 0.139533f
C10915 VDD.n707 VSS 0.139533f
C10916 VDD.n708 VSS 0.139533f
C10917 VDD.n709 VSS 0.139533f
C10918 VDD.n710 VSS 0.139533f
C10919 VDD.n711 VSS 0.139533f
C10920 VDD.n712 VSS 0.139533f
C10921 VDD.n713 VSS 0.139533f
C10922 VDD.n714 VSS 0.139533f
C10923 VDD.n715 VSS 0.139533f
C10924 VDD.n716 VSS 0.139533f
C10925 VDD.n717 VSS 0.139533f
C10926 VDD.n718 VSS 0.139533f
C10927 VDD.n719 VSS 0.139533f
C10928 VDD.n720 VSS 0.139533f
C10929 VDD.n721 VSS 0.139533f
C10930 VDD.n722 VSS 0.139533f
C10931 VDD.n723 VSS 0.139533f
C10932 VDD.n724 VSS 0.139533f
C10933 VDD.n725 VSS 0.139533f
C10934 VDD.n726 VSS 0.139533f
C10935 VDD.n727 VSS 0.139533f
C10936 VDD.n728 VSS 0.139533f
C10937 VDD.n729 VSS 0.139533f
C10938 VDD.n730 VSS 0.139533f
C10939 VDD.n731 VSS 0.139533f
C10940 VDD.n732 VSS 0.139533f
C10941 VDD.n733 VSS 0.139533f
C10942 VDD.n734 VSS 0.139533f
C10943 VDD.n735 VSS 0.139533f
C10944 VDD.n736 VSS 0.139533f
C10945 VDD.n737 VSS 0.139533f
C10946 VDD.n738 VSS 0.139533f
C10947 VDD.n739 VSS 0.139533f
C10948 VDD.n740 VSS 0.139533f
C10949 VDD.n741 VSS 0.139533f
C10950 VDD.n742 VSS 0.139533f
C10951 VDD.n743 VSS 0.139533f
C10952 VDD.n744 VSS 0.139533f
C10953 VDD.n745 VSS 0.139533f
C10954 VDD.n746 VSS 0.139533f
C10955 VDD.n747 VSS 0.139533f
C10956 VDD.n748 VSS 0.139533f
C10957 VDD.n749 VSS 0.139533f
C10958 VDD.n750 VSS 0.139533f
C10959 VDD.n751 VSS 0.139533f
C10960 VDD.n752 VSS 0.139533f
C10961 VDD.n753 VSS 0.139533f
C10962 VDD.n754 VSS 0.139533f
C10963 VDD.n755 VSS 0.139533f
C10964 VDD.n756 VSS 0.139533f
C10965 VDD.n757 VSS 0.139533f
C10966 VDD.n758 VSS 0.139533f
C10967 VDD.n759 VSS 0.139533f
C10968 VDD.n760 VSS 0.139533f
C10969 VDD.n761 VSS 0.139533f
C10970 VDD.n762 VSS 0.139533f
C10971 VDD.n763 VSS 0.139533f
C10972 VDD.n764 VSS 0.139533f
C10973 VDD.n765 VSS 0.139533f
C10974 VDD.n766 VSS 0.139533f
C10975 VDD.n767 VSS 0.139533f
C10976 VDD.n768 VSS 0.139533f
C10977 VDD.n769 VSS 0.139533f
C10978 VDD.n770 VSS 0.139533f
C10979 VDD.n771 VSS 0.139533f
C10980 VDD.n772 VSS 0.091385f
C10981 VDD.n773 VSS 0.139533f
C10982 VDD.n774 VSS 0.117916f
C10983 VDD.n775 VSS 0.139533f
C10984 VDD.n776 VSS 0.139533f
C10985 VDD.n777 VSS 0.139533f
C10986 VDD.n778 VSS 0.139533f
C10987 VDD.n779 VSS 0.139533f
C10988 VDD.n780 VSS 0.139533f
C10989 VDD.n781 VSS 0.139533f
C10990 VDD.n782 VSS 0.139533f
C10991 VDD.n783 VSS 0.139533f
C10992 VDD.n784 VSS 0.139533f
C10993 VDD.n785 VSS 0.139533f
C10994 VDD.n786 VSS 0.139533f
C10995 VDD.n787 VSS 0.139533f
C10996 VDD.n788 VSS 0.077628f
C10997 VDD.n789 VSS 0.087471f
C10998 VDD.n790 VSS 0.305376f
C10999 VDD.t4 VSS 0.037778f
C11000 VDD.n791 VSS 0.071823f
C11001 VDD.t52 VSS 0.025443f
C11002 VDD.t50 VSS 0.064018f
C11003 VDD.t68 VSS 0.069226f
C11004 VDD.n792 VSS 0.082934f
C11005 VDD.n793 VSS 0.004282f
C11006 VDD.n794 VSS 0.002308f
C11007 VDD.n795 VSS 0.006064f
C11008 VDD.n796 VSS 0.033353f
C11009 VDD.n797 VSS 0.005155f
C11010 VDD.n798 VSS 0.006064f
C11011 VDD.n799 VSS 0.003639f
C11012 VDD.n800 VSS 0.006974f
C11013 VDD.n801 VSS 0.006974f
C11014 VDD.n802 VSS 0.053365f
C11015 VDD.t39 VSS 0.022235f
C11016 VDD.n803 VSS 0.006974f
C11017 VDD.n806 VSS 0.003639f
C11018 VDD.n807 VSS 0.005155f
C11019 VDD.n808 VSS 0.005155f
C11020 VDD.n809 VSS 0.003639f
C11021 VDD.n810 VSS 0.006974f
C11022 VDD.n811 VSS 0.004548f
C11023 VDD.n812 VSS 0.006064f
C11024 VDD.n813 VSS 0.033353f
C11025 VDD.n814 VSS 0.006064f
C11026 VDD.n815 VSS 0.004548f
C11027 VDD.n816 VSS 0.004548f
C11028 VDD.n817 VSS 0.006974f
C11029 VDD.n818 VSS 0.006974f
C11030 VDD.n819 VSS 0.053365f
C11031 VDD.n820 VSS 0.006974f
C11032 VDD.n821 VSS 0.002847f
C11033 VDD.n822 VSS 0.103872f
C11034 VDD.n823 VSS 0.059346f
C11035 VDD.n824 VSS 0.044494f
C11036 VDD.n825 VSS 0.026042f
C11037 VDD.n826 VSS -0.013793f
C11038 VDD.n827 VSS 0.121773f
C11039 VDD.t51 VSS 0.287817f
C11040 VDD.n828 VSS 0.404311f
C11041 VDD.n829 VSS 0.026716f
C11042 VDD.n830 VSS 0.017231f
C11043 VDD.t15 VSS 0.037778f
C11044 VDD.n831 VSS 0.0541f
C11045 VDD.n832 VSS -0.013793f
C11046 VDD.n833 VSS 0.121773f
C11047 VDD.t12 VSS 0.289019f
C11048 VDD.n834 VSS 0.305376f
C11049 VDD.n835 VSS 0.087471f
C11050 VDD.n836 VSS 0.105141f
C11051 VDD.n837 VSS 0.139533f
C11052 VDD.n838 VSS 0.139533f
C11053 VDD.n839 VSS 0.139533f
C11054 VDD.n840 VSS 0.139533f
C11055 VDD.n841 VSS 0.139533f
C11056 VDD.n842 VSS 0.139533f
C11057 VDD.n843 VSS 0.139533f
C11058 VDD.n844 VSS 0.139533f
C11059 VDD.n845 VSS 0.139533f
C11060 VDD.n846 VSS 0.139533f
C11061 VDD.n847 VSS 0.139533f
C11062 VDD.n848 VSS 0.139533f
C11063 VDD.n849 VSS 0.139533f
C11064 VDD.n850 VSS 0.139533f
C11065 VDD.n851 VSS 0.139533f
C11066 VDD.n852 VSS 0.139533f
C11067 VDD.n853 VSS 0.139533f
C11068 VDD.n854 VSS 0.139533f
C11069 VDD.n855 VSS 0.139533f
C11070 VDD.n856 VSS 0.139533f
C11071 VDD.n857 VSS 0.139533f
C11072 VDD.n858 VSS 0.139533f
C11073 VDD.n859 VSS 0.139533f
C11074 VDD.n860 VSS 0.139533f
C11075 VDD.n861 VSS 0.139533f
C11076 VDD.n862 VSS 0.139533f
C11077 VDD.n863 VSS 0.139533f
C11078 VDD.n864 VSS 0.139533f
C11079 VDD.n865 VSS 0.139533f
C11080 VDD.n866 VSS 0.139533f
C11081 VDD.n867 VSS 0.139533f
C11082 VDD.n868 VSS 0.139533f
C11083 VDD.n869 VSS 0.139533f
C11084 VDD.n870 VSS 0.139533f
C11085 VDD.n871 VSS 0.139533f
C11086 VDD.n872 VSS 0.139533f
C11087 VDD.n873 VSS 0.139533f
C11088 VDD.n874 VSS 0.139533f
C11089 VDD.n875 VSS 0.139533f
C11090 VDD.n876 VSS 0.139533f
C11091 VDD.n877 VSS 0.139533f
C11092 VDD.n878 VSS 0.139533f
C11093 VDD.n879 VSS 0.139533f
C11094 VDD.n880 VSS 0.139533f
C11095 VDD.n881 VSS 0.139533f
C11096 VDD.n882 VSS 0.139533f
C11097 VDD.n883 VSS 0.125777f
C11098 VDD.n884 VSS 0.139533f
C11099 VDD.n885 VSS 0.139533f
C11100 VDD.n886 VSS 0.139533f
C11101 VDD.n887 VSS 0.139533f
C11102 VDD.n888 VSS 0.139533f
C11103 VDD.n889 VSS 0.139533f
C11104 VDD.n890 VSS 0.139533f
C11105 VDD.n891 VSS 0.139533f
C11106 VDD.n892 VSS 0.139533f
C11107 VDD.n893 VSS 0.139533f
C11108 VDD.n894 VSS 0.139533f
C11109 VDD.n895 VSS 0.139533f
C11110 VDD.n896 VSS 0.139533f
C11111 VDD.n897 VSS 0.139533f
C11112 VDD.n898 VSS 0.082541f
C11113 VDD.n899 VSS 0.087821f
C11114 VDD.n900 VSS 0.303768f
C11115 VDD.t1 VSS 0.289019f
C11116 VDD.n901 VSS 0.121773f
C11117 VDD.n902 VSS -0.013793f
C11118 VDD.n903 VSS 0.0541f
C11119 VDD.n904 VSS 0.374678f
C11120 VDD.n905 VSS 1.40036f
C11121 VDD.n906 VSS 0.096859f
C11122 VDD.n907 VSS 0.069767f
C11123 VDD.n908 VSS 0.039867f
C11124 VDD.n909 VSS 0.039867f
C11125 VDD.n910 VSS 0.039867f
C11126 VDD.n911 VSS 0.039867f
C11127 VDD.n917 VSS 0.069767f
C11128 VDD.n918 VSS 0.069767f
C11129 VDD.n919 VSS 0.139533f
C11130 VDD.n920 VSS 0.137568f
C11131 VDD.n921 VSS 0.139533f
C11132 VDD.n922 VSS 0.520817f
C11133 VDD.n923 VSS 0.266933f
C11134 VDD.n928 VSS 0.268086f
C11135 VDD.n929 VSS 0.035094f
C11136 VDD.n930 VSS 0.069767f
C11137 VDD.n931 VSS 0.129216f
C11138 VDD.n932 VSS 0.083523f
C11139 VDD.n933 VSS 0.083523f
C11140 PU.t4 VSS 0.540989f
C11141 PU.t3 VSS 0.546481f
C11142 PU.n0 VSS 0.618798f
C11143 PU.n1 VSS 0.045359f
C11144 PU.t1 VSS 0.131457f
C11145 PU.n2 VSS 0.126931f
C11146 PU.t5 VSS 0.328163f
C11147 PU.t2 VSS 0.589961f
C11148 PU.n3 VSS 0.586763f
C11149 PU.n4 VSS 0.473031f
C11150 PU.t0 VSS 0.237171f
C11151 PU.n5 VSS 1.0599f
C11152 PU.n6 VSS 6.29129f
C11153 PU.t6 VSS 0.263463f
C11154 PU.n7 VSS 0.129121f
C11155 PU.n8 VSS 6.62889f
C11156 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_cms_smt_0.nmos_6p0_CDNS_4066195314540_0.S.t4 VSS 0.133903f
C11157 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_cms_smt_0.nmos_6p0_CDNS_4066195314540_0.S.t2 VSS 0.152948f
C11158 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_cms_smt_0.nmos_6p0_CDNS_4066195314540_0.S.t0 VSS 0.036976f
C11159 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_cms_smt_0.nmos_6p0_CDNS_4066195314540_0.S.t5 VSS 0.086707f
C11160 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_cms_smt_0.nmos_6p0_CDNS_4066195314540_0.S.t6 VSS 0.113596f
C11161 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_cms_smt_0.nmos_6p0_CDNS_4066195314540_0.S.t1 VSS 0.097639f
C11162 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_cms_smt_0.nmos_6p0_CDNS_4066195314540_0.S.t3 VSS 0.097738f
C11163 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_drv_0.A.n0 VSS 2.16238f
C11164 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_drv_0.A.t2 VSS 0.311005f
C11165 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_drv_0.A.t7 VSS 0.301456f
C11166 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_drv_0.A.t6 VSS 0.215035f
C11167 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_drv_0.A.n1 VSS 1.2991f
C11168 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_drv_0.A.n2 VSS 0.289908f
C11169 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_drv_0.A.t10 VSS 0.445267f
C11170 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_drv_0.A.t9 VSS 0.314023f
C11171 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_drv_0.A.n3 VSS 0.431502f
C11172 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_drv_0.A.t11 VSS 0.473114f
C11173 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_drv_0.A.t8 VSS 0.122036f
C11174 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_drv_0.A.t4 VSS 0.122044f
C11175 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_drv_0.A.t0 VSS 0.066482f
C11176 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_drv_0.A.t1 VSS 0.067162f
C11177 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_drv_0.A.t3 VSS 0.065232f
C11178 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_drv_0.A.n4 VSS 0.625782f
C11179 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_drv_0.A.t5 VSS 0.215061f
C11180 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_drv_0.A.n5 VSS 0.577838f
C11181 GF_NI_IN_C_BASE_0.comp018green_esd_cdm_0.IP_IN.n0 VSS 3.15767f
C11182 GF_NI_IN_C_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_pupd_0.ppolyf_u_CDNS_4066195314532_0.PLUS VSS 82.8841f
C11183 GF_NI_IN_C_BASE_0.comp018green_esd_cdm_0.IP_IN.t4 VSS 0.254635f
C11184 GF_NI_IN_C_BASE_0.comp018green_esd_cdm_0.IP_IN.t12 VSS 0.25282f
C11185 GF_NI_IN_C_BASE_0.comp018green_esd_cdm_0.IP_IN.t11 VSS 0.25282f
C11186 GF_NI_IN_C_BASE_0.comp018green_esd_cdm_0.IP_IN.t2 VSS 0.25282f
C11187 GF_NI_IN_C_BASE_0.comp018green_esd_cdm_0.IP_IN.t5 VSS 0.179786f
C11188 GF_NI_IN_C_BASE_0.comp018green_esd_cdm_0.IP_IN.t8 VSS 0.176741f
C11189 GF_NI_IN_C_BASE_0.comp018green_esd_cdm_0.IP_IN.t10 VSS 0.162077f
C11190 GF_NI_IN_C_BASE_0.comp018green_esd_cdm_0.IP_IN.t9 VSS 0.158929f
C11191 GF_NI_IN_C_BASE_0.comp018green_esd_cdm_0.IP_IN.t7 VSS 0.279759f
C11192 GF_NI_IN_C_BASE_0.comp018green_esd_cdm_0.IP_IN.t6 VSS 0.279759f
C11193 GF_NI_IN_C_BASE_0.comp018green_esd_cdm_0.IP_IN.t3 VSS 0.279759f
C11194 GF_NI_IN_C_BASE_0.comp018green_esd_cdm_0.IP_IN.t1 VSS 0.279759f
C11195 GF_NI_IN_C_BASE_0.comp018green_esd_cdm_0.IP_IN.t0 VSS 0.048603f
C11196 DVSS.n0 VSS 0.127092f
C11197 DVSS.n1 VSS 0.168761f
C11198 DVSS.n2 VSS 0.197235f
C11199 DVSS.n3 VSS 0.197235f
C11200 DVSS.n4 VSS 0.197235f
C11201 DVSS.n5 VSS 0.111118f
C11202 DVSS.n6 VSS 0.098618f
C11203 DVSS.n7 VSS 0.014332f
C11204 DVSS.n8 VSS 0.014332f
C11205 DVSS.n9 VSS 0.014332f
C11206 DVSS.n10 VSS 0.014332f
C11207 DVSS.n11 VSS 0.014332f
C11208 DVSS.n12 VSS 0.014332f
C11209 DVSS.n13 VSS 0.014332f
C11210 DVSS.n14 VSS 0.014332f
C11211 DVSS.n15 VSS 0.014332f
C11212 DVSS.n16 VSS 0.014332f
C11213 DVSS.n17 VSS 0.014332f
C11214 DVSS.n18 VSS 0.014332f
C11215 DVSS.n19 VSS 0.014332f
C11216 DVSS.n20 VSS 0.014332f
C11217 DVSS.n21 VSS 0.014332f
C11218 DVSS.n22 VSS 0.014332f
C11219 DVSS.n23 VSS 0.014332f
C11220 DVSS.n24 VSS 0.014332f
C11221 DVSS.n25 VSS 0.007166f
C11222 DVSS.n26 VSS 0.247275f
C11223 DVSS.n27 VSS 0.197235f
C11224 DVSS.n28 VSS 0.179178f
C11225 DVSS.n29 VSS 0.197235f
C11226 DVSS.n30 VSS 0.197235f
C11227 DVSS.n31 VSS 0.197235f
C11228 DVSS.n32 VSS 0.197235f
C11229 DVSS.n33 VSS 0.197235f
C11230 DVSS.n34 VSS 0.197235f
C11231 DVSS.n35 VSS 0.197235f
C11232 DVSS.n36 VSS 0.197235f
C11233 DVSS.n37 VSS 0.197235f
C11234 DVSS.n38 VSS 0.197235f
C11235 DVSS.n39 VSS 0.197235f
C11236 DVSS.n40 VSS 0.237516f
C11237 DVSS.n41 VSS 0.237516f
C11238 DVSS.n42 VSS 0.115285f
C11239 DVSS.n43 VSS 0.237516f
C11240 DVSS.n44 VSS 0.115285f
C11241 DVSS.n45 VSS 0.197235f
C11242 DVSS.n46 VSS 0.376414f
C11243 DVSS.n47 VSS 0.237516f
C11244 DVSS.n48 VSS 0.098618f
C11245 DVSS.n49 VSS 0.197235f
C11246 DVSS.n50 VSS 0.141676f
C11247 DVSS.n51 VSS 0.197235f
C11248 DVSS.n52 VSS 0.197235f
C11249 DVSS.n53 VSS 0.197235f
C11250 DVSS.n54 VSS 0.125703f
C11251 DVSS.n55 VSS 0.001949f
C11252 DVSS.n56 VSS 0.023022f
C11253 DVSS.n57 VSS 0.025749f
C11254 DVSS.n58 VSS 0.044438f
C11255 DVSS.t101 VSS 4.60438f
C11256 DVSS.n60 VSS 0.825745f
C11257 DVSS.n61 VSS 0.226854f
C11258 DVSS.n62 VSS 0.051498f
C11259 DVSS.n63 VSS 0.023022f
C11260 DVSS.n64 VSS 0.051498f
C11261 DVSS.n65 VSS 0.023022f
C11262 DVSS.n66 VSS 0.051498f
C11263 DVSS.n67 VSS 0.023022f
C11264 DVSS.n68 VSS 0.051498f
C11265 DVSS.n69 VSS 0.023022f
C11266 DVSS.n70 VSS 0.051498f
C11267 DVSS.n71 VSS 0.023022f
C11268 DVSS.n72 VSS 0.023022f
C11269 DVSS.n73 VSS 0.023022f
C11270 DVSS.n74 VSS 0.051498f
C11271 DVSS.n75 VSS 0.051498f
C11272 DVSS.n76 VSS 0.051498f
C11273 DVSS.n77 VSS 0.023022f
C11274 DVSS.n78 VSS 0.023022f
C11275 DVSS.n79 VSS 0.023022f
C11276 DVSS.n80 VSS 0.051498f
C11277 DVSS.n81 VSS 0.051498f
C11278 DVSS.n82 VSS 0.051498f
C11279 DVSS.n83 VSS 0.023022f
C11280 DVSS.n84 VSS 0.023022f
C11281 DVSS.n85 VSS 0.023022f
C11282 DVSS.n86 VSS 0.051498f
C11283 DVSS.n87 VSS 0.051498f
C11284 DVSS.n88 VSS 0.051498f
C11285 DVSS.n89 VSS 0.023022f
C11286 DVSS.n90 VSS 0.023022f
C11287 DVSS.n91 VSS 0.023022f
C11288 DVSS.n92 VSS 0.051498f
C11289 DVSS.n93 VSS 0.051498f
C11290 DVSS.n94 VSS 0.051498f
C11291 DVSS.n95 VSS 0.023022f
C11292 DVSS.n96 VSS 0.023022f
C11293 DVSS.n97 VSS 0.023022f
C11294 DVSS.n98 VSS 0.051498f
C11295 DVSS.n99 VSS 0.051498f
C11296 DVSS.n100 VSS 0.051498f
C11297 DVSS.n101 VSS 0.012903f
C11298 DVSS.n102 VSS 0.17015f
C11299 DVSS.n103 VSS 0.141676f
C11300 DVSS.n104 VSS 0.197235f
C11301 DVSS.n105 VSS 0.098618f
C11302 DVSS.n106 VSS 0.072227f
C11303 DVSS.n107 VSS 0.115285f
C11304 DVSS.n108 VSS 0.197235f
C11305 DVSS.n109 VSS 0.197235f
C11306 DVSS.n110 VSS 0.197235f
C11307 DVSS.n111 VSS 0.197235f
C11308 DVSS.n112 VSS 0.197235f
C11309 DVSS.n113 VSS 0.197235f
C11310 DVSS.n114 VSS 0.197235f
C11311 DVSS.n115 VSS 0.197235f
C11312 DVSS.n116 VSS 0.197235f
C11313 DVSS.n117 VSS 0.197235f
C11314 DVSS.n118 VSS 0.197235f
C11315 DVSS.n119 VSS 0.197235f
C11316 DVSS.n120 VSS 0.197235f
C11317 DVSS.n121 VSS 0.197235f
C11318 DVSS.n122 VSS 0.197235f
C11319 DVSS.n123 VSS 0.431096f
C11320 DVSS.n124 VSS 0.197235f
C11321 DVSS.n125 VSS 0.197235f
C11322 DVSS.n126 VSS 0.197235f
C11323 DVSS.n127 VSS 0.175012f
C11324 DVSS.n128 VSS 0.175012f
C11325 DVSS.n129 VSS 0.376414f
C11326 DVSS.n130 VSS 0.197235f
C11327 DVSS.n131 VSS 0.197235f
C11328 DVSS.n132 VSS 0.120841f
C11329 DVSS.n133 VSS 0.237516f
C11330 DVSS.n134 VSS 0.120841f
C11331 DVSS.n135 VSS 0.175012f
C11332 DVSS.n136 VSS 0.197235f
C11333 DVSS.n137 VSS 0.197235f
C11334 DVSS.n138 VSS 0.197235f
C11335 DVSS.n139 VSS 0.197235f
C11336 DVSS.n140 VSS 0.197235f
C11337 DVSS.n141 VSS 0.117369f
C11338 DVSS.n142 VSS 0.197235f
C11339 DVSS.n143 VSS 0.197235f
C11340 DVSS.n144 VSS 0.117369f
C11341 DVSS.n145 VSS 0.197235f
C11342 DVSS.n146 VSS 0.197235f
C11343 DVSS.n147 VSS 0.197235f
C11344 DVSS.n148 VSS 0.197235f
C11345 DVSS.n149 VSS 0.197235f
C11346 DVSS.n150 VSS 0.175012f
C11347 DVSS.n151 VSS 0.175012f
C11348 DVSS.n152 VSS 0.197235f
C11349 DVSS.n153 VSS 0.197235f
C11350 DVSS.n154 VSS 0.197235f
C11351 DVSS.n155 VSS 0.237516f
C11352 DVSS.n156 VSS 0.197235f
C11353 DVSS.n157 VSS 0.197235f
C11354 DVSS.n158 VSS 0.197235f
C11355 DVSS.n159 VSS 0.197235f
C11356 DVSS.n160 VSS 0.197235f
C11357 DVSS.n161 VSS 0.197235f
C11358 DVSS.n162 VSS 0.197235f
C11359 DVSS.n163 VSS 0.197235f
C11360 DVSS.n164 VSS 0.197235f
C11361 DVSS.n165 VSS 0.197235f
C11362 DVSS.n166 VSS 0.197235f
C11363 DVSS.n167 VSS 0.197235f
C11364 DVSS.n168 VSS 0.163205f
C11365 DVSS.n169 VSS 0.485035f
C11366 DVSS.n170 VSS 0.163205f
C11367 DVSS.n171 VSS 0.197235f
C11368 DVSS.n172 VSS 0.197235f
C11369 DVSS.n173 VSS 0.197235f
C11370 DVSS.n174 VSS 0.197235f
C11371 DVSS.n175 VSS 0.197235f
C11372 DVSS.n176 VSS 0.197235f
C11373 DVSS.n177 VSS 0.197235f
C11374 DVSS.n178 VSS 0.197235f
C11375 DVSS.n179 VSS 0.197235f
C11376 DVSS.n180 VSS 0.197235f
C11377 DVSS.n181 VSS 0.197235f
C11378 DVSS.n182 VSS 0.197235f
C11379 DVSS.n183 VSS 0.197235f
C11380 DVSS.n184 VSS 0.237516f
C11381 DVSS.n185 VSS 0.237516f
C11382 DVSS.n186 VSS 0.376414f
C11383 DVSS.n187 VSS 0.197235f
C11384 DVSS.n188 VSS 0.197235f
C11385 DVSS.n189 VSS 0.185429f
C11386 DVSS.n190 VSS 0.197235f
C11387 DVSS.n191 VSS 0.197235f
C11388 DVSS.n192 VSS 0.197235f
C11389 DVSS.n193 VSS 0.197235f
C11390 DVSS.n194 VSS 0.485035f
C11391 DVSS.n195 VSS 0.110424f
C11392 DVSS.n196 VSS 0.197235f
C11393 DVSS.n197 VSS 0.197235f
C11394 DVSS.n198 VSS 0.197235f
C11395 DVSS.n199 VSS 0.197235f
C11396 DVSS.n200 VSS 0.126397f
C11397 DVSS.n201 VSS 0.197235f
C11398 DVSS.n202 VSS 0.126397f
C11399 DVSS.n203 VSS 0.237516f
C11400 DVSS.n204 VSS 0.126397f
C11401 DVSS.n205 VSS 0.197235f
C11402 DVSS.n206 VSS 0.197235f
C11403 DVSS.n207 VSS 0.197235f
C11404 DVSS.n208 VSS 0.197235f
C11405 DVSS.n209 VSS 0.197235f
C11406 DVSS.n210 VSS 0.197235f
C11407 DVSS.n211 VSS 0.197235f
C11408 DVSS.n212 VSS 0.197235f
C11409 DVSS.n213 VSS 0.197235f
C11410 DVSS.n214 VSS 0.197235f
C11411 DVSS.n215 VSS 0.197235f
C11412 DVSS.n216 VSS 0.197235f
C11413 DVSS.n217 VSS 0.197235f
C11414 DVSS.n218 VSS 0.197235f
C11415 DVSS.n219 VSS 0.197235f
C11416 DVSS.n220 VSS 0.197235f
C11417 DVSS.n221 VSS 0.197235f
C11418 DVSS.n222 VSS 0.197235f
C11419 DVSS.n223 VSS 0.197235f
C11420 DVSS.n224 VSS 0.136815f
C11421 DVSS.n225 VSS 0.197235f
C11422 DVSS.n226 VSS 0.197235f
C11423 DVSS.n227 VSS 0.197235f
C11424 DVSS.n228 VSS 0.10834f
C11425 DVSS.n229 VSS 0.257556f
C11426 DVSS.n230 VSS 0.025376f
C11427 DVSS.n231 VSS 0.054081f
C11428 DVSS.n232 VSS 0.025376f
C11429 DVSS.n233 VSS 0.054081f
C11430 DVSS.n234 VSS 0.025376f
C11431 DVSS.n235 VSS 0.054081f
C11432 DVSS.n236 VSS 0.025376f
C11433 DVSS.n237 VSS 0.054081f
C11434 DVSS.n238 VSS 0.025376f
C11435 DVSS.n239 VSS 0.054081f
C11436 DVSS.n240 VSS 0.025376f
C11437 DVSS.n241 VSS 0.027041f
C11438 DVSS.n242 VSS 0.003274f
C11439 DVSS.n243 VSS 0.154177f
C11440 DVSS.n244 VSS 0.159038f
C11441 DVSS.n245 VSS 0.1639f
C11442 DVSS.n246 VSS 0.197235f
C11443 DVSS.n247 VSS 3.37033f
C11444 DVSS.n248 VSS 3.59901f
C11445 DVSS.n249 VSS 1.79594f
C11446 DVSS.n250 VSS 0.963609f
C11447 DVSS.n251 VSS 3.59901f
C11448 DVSS.n252 VSS 0.098618f
C11449 DVSS.n253 VSS 0.905847f
C11450 DVSS.n254 VSS 0.766949f
C11451 DVSS.n255 VSS 0.197235f
C11452 DVSS.n256 VSS 0.197235f
C11453 DVSS.n257 VSS 0.10834f
C11454 DVSS.n258 VSS 0.159038f
C11455 DVSS.n259 VSS 0.014223f
C11456 DVSS.n260 VSS 0.252796f
C11457 DVSS.n261 VSS 0.024864f
C11458 DVSS.n262 VSS 0.054081f
C11459 DVSS.n263 VSS 0.025376f
C11460 DVSS.n264 VSS 0.054081f
C11461 DVSS.n265 VSS 0.025376f
C11462 DVSS.n266 VSS 0.054081f
C11463 DVSS.n267 VSS 0.025376f
C11464 DVSS.n268 VSS 0.054081f
C11465 DVSS.n269 VSS 0.025376f
C11466 DVSS.n270 VSS 0.054081f
C11467 DVSS.n271 VSS 0.025376f
C11468 DVSS.n272 VSS 0.014734f
C11469 DVSS.n273 VSS 0.035981f
C11470 DVSS.n274 VSS 0.034455f
C11471 DVSS.t185 VSS 5.17029f
C11472 DVSS.t114 VSS 5.17029f
C11473 DVSS.t130 VSS 6.04903f
C11474 DVSS.n275 VSS 6.38652f
C11475 DVSS.n276 VSS 0.027041f
C11476 DVSS.n277 VSS 0.046667f
C11477 DVSS.n278 VSS 0.025376f
C11478 DVSS.n279 VSS 0.025376f
C11479 DVSS.n280 VSS 0.025376f
C11480 DVSS.n281 VSS 0.054081f
C11481 DVSS.n282 VSS 0.054081f
C11482 DVSS.n283 VSS 0.054081f
C11483 DVSS.n284 VSS 0.025376f
C11484 DVSS.n285 VSS 0.025376f
C11485 DVSS.n286 VSS 0.025376f
C11486 DVSS.n287 VSS 0.054081f
C11487 DVSS.n288 VSS 0.054081f
C11488 DVSS.n289 VSS 0.054081f
C11489 DVSS.n290 VSS 0.025376f
C11490 DVSS.n291 VSS 0.025376f
C11491 DVSS.n292 VSS 0.025376f
C11492 DVSS.n293 VSS 0.054081f
C11493 DVSS.n294 VSS 0.054081f
C11494 DVSS.n295 VSS 0.054081f
C11495 DVSS.n296 VSS 0.025376f
C11496 DVSS.n297 VSS 0.025376f
C11497 DVSS.n298 VSS 0.025376f
C11498 DVSS.n299 VSS 0.054081f
C11499 DVSS.n300 VSS 0.054081f
C11500 DVSS.n301 VSS 0.054081f
C11501 DVSS.n302 VSS 0.025376f
C11502 DVSS.n303 VSS 0.025376f
C11503 DVSS.n304 VSS 0.025376f
C11504 DVSS.n305 VSS 0.054081f
C11505 DVSS.n306 VSS 0.054081f
C11506 DVSS.n307 VSS 0.095171f
C11507 DVSS.n308 VSS 0.054081f
C11508 DVSS.n309 VSS 0.023841f
C11509 DVSS.n310 VSS 0.012688f
C11510 DVSS.n311 VSS 0.098618f
C11511 DVSS.n312 VSS 0.136815f
C11512 DVSS.n313 VSS 0.197235f
C11513 DVSS.n314 VSS 0.197235f
C11514 DVSS.n315 VSS 0.197235f
C11515 DVSS.n316 VSS 0.197235f
C11516 DVSS.n317 VSS 0.197235f
C11517 DVSS.n318 VSS 0.197235f
C11518 DVSS.n319 VSS 0.197235f
C11519 DVSS.n320 VSS 0.197235f
C11520 DVSS.n321 VSS 0.197235f
C11521 DVSS.n322 VSS 0.197235f
C11522 DVSS.n323 VSS 0.197235f
C11523 DVSS.n324 VSS 0.197235f
C11524 DVSS.n325 VSS 0.197235f
C11525 DVSS.n326 VSS 0.197235f
C11526 DVSS.n327 VSS 0.197235f
C11527 DVSS.n328 VSS 0.197235f
C11528 DVSS.n329 VSS 0.197235f
C11529 DVSS.n330 VSS 0.197235f
C11530 DVSS.n331 VSS 0.197235f
C11531 DVSS.n332 VSS 0.197235f
C11532 DVSS.n333 VSS 0.197235f
C11533 DVSS.n334 VSS 0.197235f
C11534 DVSS.n335 VSS 0.197235f
C11535 DVSS.n336 VSS 0.197235f
C11536 DVSS.n337 VSS 0.197235f
C11537 DVSS.n338 VSS 0.197235f
C11538 DVSS.n339 VSS 0.197235f
C11539 DVSS.n340 VSS 0.197235f
C11540 DVSS.n341 VSS 0.197235f
C11541 DVSS.n342 VSS 0.197235f
C11542 DVSS.n343 VSS 0.197235f
C11543 DVSS.n344 VSS 0.197235f
C11544 DVSS.n345 VSS 0.197235f
C11545 DVSS.n346 VSS 0.197235f
C11546 DVSS.n347 VSS 0.197235f
C11547 DVSS.n348 VSS 0.197235f
C11548 DVSS.n349 VSS 0.197235f
C11549 DVSS.n350 VSS 0.197235f
C11550 DVSS.n351 VSS 0.197235f
C11551 DVSS.n352 VSS 0.197235f
C11552 DVSS.n353 VSS 0.197235f
C11553 DVSS.n354 VSS 0.197235f
C11554 DVSS.n355 VSS 0.197235f
C11555 DVSS.n356 VSS 0.197235f
C11556 DVSS.n357 VSS 0.197235f
C11557 DVSS.n358 VSS 0.197235f
C11558 DVSS.n359 VSS 0.1639f
C11559 DVSS.n360 VSS 0.1639f
C11560 DVSS.n361 VSS 0.154177f
C11561 DVSS.n362 VSS 2.72273f
C11562 DVSS.n363 VSS 2.86163f
C11563 DVSS.n364 VSS 4.28235f
C11564 DVSS.n365 VSS 0.098618f
C11565 DVSS.n366 VSS 0.154177f
C11566 DVSS.n367 VSS 0.1639f
C11567 DVSS.n368 VSS 0.1639f
C11568 DVSS.n369 VSS 3.41712f
C11569 DVSS.n370 VSS 3.50923f
C11570 DVSS.n371 VSS 0.1639f
C11571 DVSS.n372 VSS 0.197235f
C11572 DVSS.n373 VSS 0.098618f
C11573 DVSS.n374 VSS 0.136815f
C11574 DVSS.n375 VSS 0.197235f
C11575 DVSS.n376 VSS 0.197235f
C11576 DVSS.n377 VSS 0.197235f
C11577 DVSS.n378 VSS 0.197235f
C11578 DVSS.n379 VSS 0.197235f
C11579 DVSS.n380 VSS 0.197235f
C11580 DVSS.n381 VSS 0.197235f
C11581 DVSS.n382 VSS 0.197235f
C11582 DVSS.n383 VSS 0.197235f
C11583 DVSS.n384 VSS 0.197235f
C11584 DVSS.n385 VSS 0.197235f
C11585 DVSS.n386 VSS 0.197235f
C11586 DVSS.n387 VSS 0.197235f
C11587 DVSS.n388 VSS 0.197235f
C11588 DVSS.n389 VSS 0.197235f
C11589 DVSS.n390 VSS 0.197235f
C11590 DVSS.n391 VSS 0.197235f
C11591 DVSS.n392 VSS 0.197235f
C11592 DVSS.n393 VSS 0.197235f
C11593 DVSS.n394 VSS 0.197235f
C11594 DVSS.n395 VSS 0.197235f
C11595 DVSS.n396 VSS 0.197235f
C11596 DVSS.n397 VSS 0.197235f
C11597 DVSS.n398 VSS 0.197235f
C11598 DVSS.n399 VSS 0.197235f
C11599 DVSS.n400 VSS 0.197235f
C11600 DVSS.n401 VSS 0.197235f
C11601 DVSS.n402 VSS 0.197235f
C11602 DVSS.n403 VSS 0.197235f
C11603 DVSS.n404 VSS 0.197235f
C11604 DVSS.n405 VSS 0.197235f
C11605 DVSS.n406 VSS 0.197235f
C11606 DVSS.n407 VSS 0.197235f
C11607 DVSS.n408 VSS 0.197235f
C11608 DVSS.n409 VSS 0.197235f
C11609 DVSS.n410 VSS 0.197235f
C11610 DVSS.n411 VSS 0.197235f
C11611 DVSS.n412 VSS 0.197235f
C11612 DVSS.n413 VSS 0.197235f
C11613 DVSS.n414 VSS 0.197235f
C11614 DVSS.n415 VSS 0.197235f
C11615 DVSS.n416 VSS 0.197235f
C11616 DVSS.n417 VSS 0.197235f
C11617 DVSS.n418 VSS 0.197235f
C11618 DVSS.n419 VSS 0.197235f
C11619 DVSS.n420 VSS 0.197235f
C11620 DVSS.n421 VSS 0.197235f
C11621 DVSS.n422 VSS 0.197235f
C11622 DVSS.n423 VSS 0.197235f
C11623 DVSS.n424 VSS 0.10834f
C11624 DVSS.n425 VSS 0.098618f
C11625 DVSS.n426 VSS 0.002149f
C11626 DVSS.n427 VSS 0.009414f
C11627 DVSS.n428 VSS 0.021181f
C11628 DVSS.n429 VSS 0.030668f
C11629 DVSS.n430 VSS -0.290359f
C11630 DVSS.n431 VSS 0.054081f
C11631 DVSS.n432 VSS 0.025376f
C11632 DVSS.n433 VSS 0.025376f
C11633 DVSS.n434 VSS 0.025376f
C11634 DVSS.n435 VSS 0.054081f
C11635 DVSS.n436 VSS 0.054081f
C11636 DVSS.n437 VSS 0.054081f
C11637 DVSS.n438 VSS 0.025376f
C11638 DVSS.n439 VSS 0.025376f
C11639 DVSS.n440 VSS 0.025376f
C11640 DVSS.n441 VSS 0.054081f
C11641 DVSS.n442 VSS 0.054081f
C11642 DVSS.n443 VSS 0.054081f
C11643 DVSS.n444 VSS 0.025376f
C11644 DVSS.n445 VSS 0.025376f
C11645 DVSS.n446 VSS 0.025376f
C11646 DVSS.n447 VSS 0.054081f
C11647 DVSS.n448 VSS 0.054081f
C11648 DVSS.n449 VSS 0.054081f
C11649 DVSS.n450 VSS 0.025376f
C11650 DVSS.n451 VSS 0.025376f
C11651 DVSS.n452 VSS 0.025376f
C11652 DVSS.n453 VSS 0.054081f
C11653 DVSS.n454 VSS 0.054081f
C11654 DVSS.n455 VSS 0.054081f
C11655 DVSS.n456 VSS 0.025376f
C11656 DVSS.n457 VSS 0.025376f
C11657 DVSS.n458 VSS 0.025376f
C11658 DVSS.n459 VSS 0.054081f
C11659 DVSS.n460 VSS 0.054081f
C11660 DVSS.n461 VSS 0.536664f
C11661 DVSS.n462 VSS 0.015655f
C11662 DVSS.n463 VSS 0.004298f
C11663 DVSS.n464 VSS 0.098618f
C11664 DVSS.n465 VSS 0.159038f
C11665 DVSS.n466 VSS 0.197235f
C11666 DVSS.n467 VSS 0.197235f
C11667 DVSS.n468 VSS 0.197235f
C11668 DVSS.n469 VSS 0.197235f
C11669 DVSS.n470 VSS 0.197235f
C11670 DVSS.n471 VSS 0.197235f
C11671 DVSS.n472 VSS 0.197235f
C11672 DVSS.n473 VSS 0.197235f
C11673 DVSS.n474 VSS 0.197235f
C11674 DVSS.n475 VSS 0.197235f
C11675 DVSS.n476 VSS 0.197235f
C11676 DVSS.n477 VSS 0.197235f
C11677 DVSS.n478 VSS 0.197235f
C11678 DVSS.n479 VSS 0.197235f
C11679 DVSS.n480 VSS 0.197235f
C11680 DVSS.n481 VSS 0.197235f
C11681 DVSS.n482 VSS 0.197235f
C11682 DVSS.n483 VSS 0.197235f
C11683 DVSS.n484 VSS 0.197235f
C11684 DVSS.n485 VSS 0.197235f
C11685 DVSS.n486 VSS 0.197235f
C11686 DVSS.n487 VSS 0.197235f
C11687 DVSS.n488 VSS 0.197235f
C11688 DVSS.n489 VSS 0.197235f
C11689 DVSS.n490 VSS 0.197235f
C11690 DVSS.n491 VSS 0.197235f
C11691 DVSS.n492 VSS 0.197235f
C11692 DVSS.n493 VSS 0.197235f
C11693 DVSS.n494 VSS 0.197235f
C11694 DVSS.n495 VSS 0.197235f
C11695 DVSS.n496 VSS 0.197235f
C11696 DVSS.n497 VSS 0.110424f
C11697 DVSS.n498 VSS 0.197235f
C11698 DVSS.n499 VSS 0.197235f
C11699 DVSS.n500 VSS 0.197235f
C11700 DVSS.n501 VSS 0.197235f
C11701 DVSS.n502 VSS 0.197235f
C11702 DVSS.n503 VSS 0.197235f
C11703 DVSS.n504 VSS 0.197235f
C11704 DVSS.n505 VSS 0.185429f
C11705 DVSS.n506 VSS 0.197235f
C11706 DVSS.n507 VSS 0.197235f
C11707 DVSS.n508 VSS 0.197235f
C11708 DVSS.n509 VSS 0.126397f
C11709 DVSS.n510 VSS 0.126397f
C11710 DVSS.n511 VSS 0.237516f
C11711 DVSS.n512 VSS 0.197235f
C11712 DVSS.n513 VSS 0.197235f
C11713 DVSS.n514 VSS 0.197235f
C11714 DVSS.n515 VSS 0.197235f
C11715 DVSS.n516 VSS 0.197235f
C11716 DVSS.n517 VSS 0.197235f
C11717 DVSS.n518 VSS 0.197235f
C11718 DVSS.n519 VSS 0.197235f
C11719 DVSS.n520 VSS 0.197235f
C11720 DVSS.n521 VSS 0.197235f
C11721 DVSS.n522 VSS 0.197235f
C11722 DVSS.n523 VSS 0.197235f
C11723 DVSS.n524 VSS 0.197235f
C11724 DVSS.n525 VSS 0.197235f
C11725 DVSS.n526 VSS 0.163205f
C11726 DVSS.n527 VSS 0.132648f
C11727 DVSS.n528 VSS 0.197235f
C11728 DVSS.n529 VSS 0.197235f
C11729 DVSS.n530 VSS 0.197235f
C11730 DVSS.n531 VSS 0.197235f
C11731 DVSS.n532 VSS 0.197235f
C11732 DVSS.n533 VSS 0.197235f
C11733 DVSS.n534 VSS 0.197235f
C11734 DVSS.n535 VSS 0.197235f
C11735 DVSS.n536 VSS 0.197235f
C11736 DVSS.n537 VSS 0.197235f
C11737 DVSS.n538 VSS 0.197235f
C11738 DVSS.n539 VSS 0.197235f
C11739 DVSS.n540 VSS 0.197235f
C11740 DVSS.n541 VSS 0.197235f
C11741 DVSS.n542 VSS 0.197235f
C11742 DVSS.n543 VSS 0.197235f
C11743 DVSS.n544 VSS 0.197235f
C11744 DVSS.n545 VSS 0.197235f
C11745 DVSS.n546 VSS 0.197235f
C11746 DVSS.n547 VSS 0.197235f
C11747 DVSS.n548 VSS 0.197235f
C11748 DVSS.n549 VSS 0.197235f
C11749 DVSS.n550 VSS 0.197235f
C11750 DVSS.n551 VSS 0.197235f
C11751 DVSS.n552 VSS 0.197235f
C11752 DVSS.n553 VSS 0.197235f
C11753 DVSS.n554 VSS 0.197235f
C11754 DVSS.n555 VSS 0.197235f
C11755 DVSS.n556 VSS 0.197235f
C11756 DVSS.n557 VSS 0.197235f
C11757 DVSS.n558 VSS 0.197235f
C11758 DVSS.n559 VSS 0.197235f
C11759 DVSS.n560 VSS 0.197235f
C11760 DVSS.n561 VSS 0.197235f
C11761 DVSS.n562 VSS 0.197235f
C11762 DVSS.n563 VSS 0.197235f
C11763 DVSS.n564 VSS 0.197235f
C11764 DVSS.n565 VSS 0.197235f
C11765 DVSS.n566 VSS 0.197235f
C11766 DVSS.n567 VSS 0.197235f
C11767 DVSS.n568 VSS 0.197235f
C11768 DVSS.n569 VSS 0.197235f
C11769 DVSS.n570 VSS 0.197235f
C11770 DVSS.n571 VSS 0.197235f
C11771 DVSS.n572 VSS 0.197235f
C11772 DVSS.n573 VSS 0.169456f
C11773 DVSS.n574 VSS 0.169456f
C11774 DVSS.n575 VSS 0.169456f
C11775 DVSS.n576 VSS 0.237516f
C11776 DVSS.n577 VSS 0.376414f
C11777 DVSS.n578 VSS 0.169456f
C11778 DVSS.n579 VSS 0.197235f
C11779 DVSS.n580 VSS 0.197235f
C11780 DVSS.n581 VSS 0.197235f
C11781 DVSS.n582 VSS 0.197235f
C11782 DVSS.n583 VSS 0.197235f
C11783 DVSS.n584 VSS 0.197235f
C11784 DVSS.n585 VSS 0.197235f
C11785 DVSS.n586 VSS 0.197235f
C11786 DVSS.n587 VSS 0.197235f
C11787 DVSS.n588 VSS 0.197235f
C11788 DVSS.n589 VSS 0.197235f
C11789 DVSS.n590 VSS 0.197235f
C11790 DVSS.n591 VSS 0.197235f
C11791 DVSS.n592 VSS 0.197235f
C11792 DVSS.n593 VSS 0.197235f
C11793 DVSS.n594 VSS 0.197235f
C11794 DVSS.n595 VSS 0.197235f
C11795 DVSS.n596 VSS 0.197235f
C11796 DVSS.n597 VSS 0.197235f
C11797 DVSS.n598 VSS 0.197235f
C11798 DVSS.n599 VSS 0.197235f
C11799 DVSS.n600 VSS 0.197235f
C11800 DVSS.n601 VSS 0.197235f
C11801 DVSS.n602 VSS 0.197235f
C11802 DVSS.n603 VSS 0.197235f
C11803 DVSS.n604 VSS 0.197235f
C11804 DVSS.n605 VSS 0.197235f
C11805 DVSS.n606 VSS 0.197235f
C11806 DVSS.n607 VSS 0.197235f
C11807 DVSS.n608 VSS 0.197235f
C11808 DVSS.n609 VSS 0.169456f
C11809 DVSS.n610 VSS 0.169456f
C11810 DVSS.n611 VSS 0.376414f
C11811 DVSS.n612 VSS 0.126397f
C11812 DVSS.n613 VSS 0.197235f
C11813 DVSS.n614 VSS 0.197235f
C11814 DVSS.n615 VSS 0.197235f
C11815 DVSS.n616 VSS 0.197235f
C11816 DVSS.n617 VSS 0.197235f
C11817 DVSS.n618 VSS 0.185429f
C11818 DVSS.n619 VSS 0.144307f
C11819 DVSS.n620 VSS 0.48809f
C11820 DVSS.n621 VSS 0.431096f
C11821 DVSS.n622 VSS 0.110424f
C11822 DVSS.n623 VSS 0.197235f
C11823 DVSS.n624 VSS 0.197235f
C11824 DVSS.n625 VSS 0.197235f
C11825 DVSS.n626 VSS 0.197235f
C11826 DVSS.n627 VSS 0.197235f
C11827 DVSS.n628 VSS 0.197235f
C11828 DVSS.n629 VSS 0.197235f
C11829 DVSS.n630 VSS 0.126397f
C11830 DVSS.n631 VSS 0.126397f
C11831 DVSS.n632 VSS 0.126397f
C11832 DVSS.n633 VSS 0.237516f
C11833 DVSS.n634 VSS 0.169456f
C11834 DVSS.n635 VSS 0.169456f
C11835 DVSS.n636 VSS 0.169456f
C11836 DVSS.n637 VSS 0.197235f
C11837 DVSS.n638 VSS 0.197235f
C11838 DVSS.n639 VSS 0.197235f
C11839 DVSS.n640 VSS 0.197235f
C11840 DVSS.n641 VSS 0.197235f
C11841 DVSS.n642 VSS 0.197235f
C11842 DVSS.n643 VSS 0.197235f
C11843 DVSS.n644 VSS 0.197235f
C11844 DVSS.n645 VSS 0.197235f
C11845 DVSS.n646 VSS 0.197235f
C11846 DVSS.n647 VSS 0.197235f
C11847 DVSS.n648 VSS 0.197235f
C11848 DVSS.n649 VSS 0.197235f
C11849 DVSS.n650 VSS 0.197235f
C11850 DVSS.n651 VSS 0.197235f
C11851 DVSS.n652 VSS 0.197235f
C11852 DVSS.n653 VSS 0.197235f
C11853 DVSS.n654 VSS 0.197235f
C11854 DVSS.n655 VSS 0.197235f
C11855 DVSS.n656 VSS 0.197235f
C11856 DVSS.n657 VSS 0.197235f
C11857 DVSS.n658 VSS 0.197235f
C11858 DVSS.n659 VSS 0.197235f
C11859 DVSS.n660 VSS 0.197235f
C11860 DVSS.n661 VSS 0.197235f
C11861 DVSS.n662 VSS 0.197235f
C11862 DVSS.n663 VSS 0.197235f
C11863 DVSS.n664 VSS 0.197235f
C11864 DVSS.n665 VSS 0.197235f
C11865 DVSS.n666 VSS 0.197235f
C11866 DVSS.n667 VSS 0.197235f
C11867 DVSS.n668 VSS 0.197235f
C11868 DVSS.n669 VSS 0.197235f
C11869 DVSS.n670 VSS 0.197235f
C11870 DVSS.n671 VSS 0.197235f
C11871 DVSS.n672 VSS 0.197235f
C11872 DVSS.n673 VSS 0.197235f
C11873 DVSS.n674 VSS 0.197235f
C11874 DVSS.n675 VSS 0.197235f
C11875 DVSS.n676 VSS 0.197235f
C11876 DVSS.n677 VSS 0.197235f
C11877 DVSS.n678 VSS 0.197235f
C11878 DVSS.n679 VSS 0.197235f
C11879 DVSS.n680 VSS 0.197235f
C11880 DVSS.n681 VSS 0.197235f
C11881 DVSS.n682 VSS 0.197235f
C11882 DVSS.n683 VSS 0.197235f
C11883 DVSS.n684 VSS 0.197235f
C11884 DVSS.n685 VSS 0.197235f
C11885 DVSS.n686 VSS 0.132648f
C11886 DVSS.n687 VSS 0.431096f
C11887 DVSS.n688 VSS 0.48809f
C11888 DVSS.n689 VSS 0.144307f
C11889 DVSS.n690 VSS 0.132648f
C11890 DVSS.n691 VSS 0.197235f
C11891 DVSS.n692 VSS 0.197235f
C11892 DVSS.n693 VSS 0.197235f
C11893 DVSS.n694 VSS 0.197235f
C11894 DVSS.n695 VSS 0.197235f
C11895 DVSS.n696 VSS 0.197235f
C11896 DVSS.n697 VSS 0.197235f
C11897 DVSS.n698 VSS 0.197235f
C11898 DVSS.n699 VSS 0.197235f
C11899 DVSS.n700 VSS 0.197235f
C11900 DVSS.n701 VSS 0.197235f
C11901 DVSS.n702 VSS 0.197235f
C11902 DVSS.n703 VSS 0.197235f
C11903 DVSS.n704 VSS 0.197235f
C11904 DVSS.n705 VSS 0.197235f
C11905 DVSS.n706 VSS 0.197235f
C11906 DVSS.n707 VSS 0.197235f
C11907 DVSS.n708 VSS 0.197235f
C11908 DVSS.n709 VSS 0.197235f
C11909 DVSS.n710 VSS 0.120841f
C11910 DVSS.n711 VSS 0.197235f
C11911 DVSS.n712 VSS 0.197235f
C11912 DVSS.n713 VSS 0.197235f
C11913 DVSS.n714 VSS 0.120841f
C11914 DVSS.n715 VSS 0.376414f
C11915 DVSS.n716 VSS 0.237516f
C11916 DVSS.n717 VSS 0.120841f
C11917 DVSS.n718 VSS 0.120841f
C11918 DVSS.n719 VSS 0.120841f
C11919 DVSS.n720 VSS 0.237516f
C11920 DVSS.n721 VSS 0.175012f
C11921 DVSS.n722 VSS 0.197235f
C11922 DVSS.n723 VSS 0.197235f
C11923 DVSS.n724 VSS 0.197235f
C11924 DVSS.n725 VSS 0.197235f
C11925 DVSS.n726 VSS 0.197235f
C11926 DVSS.n727 VSS 0.197235f
C11927 DVSS.n728 VSS 0.197235f
C11928 DVSS.n729 VSS 0.197235f
C11929 DVSS.n730 VSS 0.197235f
C11930 DVSS.n731 VSS 0.197235f
C11931 DVSS.n732 VSS 0.197235f
C11932 DVSS.n733 VSS 0.197235f
C11933 DVSS.n734 VSS 0.197235f
C11934 DVSS.n735 VSS 0.197235f
C11935 DVSS.n736 VSS 0.197235f
C11936 DVSS.n737 VSS 0.197235f
C11937 DVSS.n738 VSS 0.197235f
C11938 DVSS.n739 VSS 0.197235f
C11939 DVSS.n740 VSS 0.197235f
C11940 DVSS.n741 VSS 0.197235f
C11941 DVSS.n742 VSS 0.197235f
C11942 DVSS.n743 VSS 0.197235f
C11943 DVSS.n744 VSS 0.197235f
C11944 DVSS.n745 VSS 0.197235f
C11945 DVSS.n746 VSS 0.197235f
C11946 DVSS.n747 VSS 0.197235f
C11947 DVSS.n748 VSS 0.197235f
C11948 DVSS.n749 VSS 0.197235f
C11949 DVSS.n750 VSS 0.17015f
C11950 DVSS.n751 VSS 0.125703f
C11951 DVSS.n752 VSS 0.197235f
C11952 DVSS.n753 VSS 0.141676f
C11953 DVSS.n754 VSS 0.512686f
C11954 DVSS.n755 VSS 0.023022f
C11955 DVSS.n756 VSS 0.051498f
C11956 DVSS.n757 VSS 0.023022f
C11957 DVSS.n758 VSS 0.051498f
C11958 DVSS.n759 VSS 0.023022f
C11959 DVSS.n760 VSS 0.051498f
C11960 DVSS.n761 VSS 0.023022f
C11961 DVSS.n762 VSS 0.051498f
C11962 DVSS.n763 VSS 0.023022f
C11963 DVSS.n764 VSS 0.051498f
C11964 DVSS.n765 VSS 0.00854f
C11965 DVSS.n766 VSS 0.019216f
C11966 DVSS.n767 VSS 0.028511f
C11967 DVSS.n768 VSS -0.292943f
C11968 DVSS.n769 VSS 0.023022f
C11969 DVSS.n770 VSS 0.023022f
C11970 DVSS.n771 VSS 0.023022f
C11971 DVSS.n772 VSS 0.051498f
C11972 DVSS.n773 VSS 0.051498f
C11973 DVSS.n774 VSS 0.051498f
C11974 DVSS.n775 VSS 0.023022f
C11975 DVSS.n776 VSS 0.023022f
C11976 DVSS.n777 VSS 0.023022f
C11977 DVSS.n778 VSS 0.051498f
C11978 DVSS.n779 VSS 0.051498f
C11979 DVSS.n780 VSS 0.051498f
C11980 DVSS.n781 VSS 0.023022f
C11981 DVSS.n782 VSS 0.023022f
C11982 DVSS.n783 VSS 0.023022f
C11983 DVSS.n784 VSS 0.051498f
C11984 DVSS.n785 VSS 0.051498f
C11985 DVSS.n786 VSS 0.051498f
C11986 DVSS.n787 VSS 0.023022f
C11987 DVSS.n788 VSS 0.023022f
C11988 DVSS.n789 VSS 0.023022f
C11989 DVSS.n790 VSS 0.051498f
C11990 DVSS.n791 VSS 0.051498f
C11991 DVSS.n792 VSS 0.051498f
C11992 DVSS.n793 VSS 0.023022f
C11993 DVSS.n794 VSS 0.023022f
C11994 DVSS.n795 VSS 0.023022f
C11995 DVSS.n796 VSS 0.051498f
C11996 DVSS.n797 VSS 0.051498f
C11997 DVSS.n798 VSS 0.051498f
C11998 DVSS.n799 VSS 0.023022f
C11999 DVSS.n800 VSS 0.014203f
C12000 DVSS.n801 VSS 0.098618f
C12001 DVSS.n802 VSS 0.003898f
C12002 DVSS.n803 VSS 0.233037f
C12003 DVSS.n804 VSS 0.098618f
C12004 DVSS.n805 VSS 0.072227f
C12005 DVSS.n806 VSS 0.180567f
C12006 DVSS.n807 VSS 0.197235f
C12007 DVSS.n808 VSS 0.197235f
C12008 DVSS.n809 VSS 0.197235f
C12009 DVSS.n810 VSS 0.197235f
C12010 DVSS.n811 VSS 0.197235f
C12011 DVSS.n812 VSS 0.197235f
C12012 DVSS.n813 VSS 0.197235f
C12013 DVSS.n814 VSS 0.197235f
C12014 DVSS.n815 VSS 0.197235f
C12015 DVSS.n816 VSS 0.197235f
C12016 DVSS.n817 VSS 0.197235f
C12017 DVSS.n818 VSS 0.197235f
C12018 DVSS.n819 VSS 0.197235f
C12019 DVSS.n820 VSS 0.101396f
C12020 DVSS.n821 VSS 0.197235f
C12021 DVSS.n822 VSS 0.17779f
C12022 DVSS.n823 VSS 0.118063f
C12023 DVSS.n824 VSS 0.197235f
C12024 DVSS.n825 VSS 0.197235f
C12025 DVSS.n826 VSS 0.197235f
C12026 DVSS.n827 VSS 0.197235f
C12027 DVSS.n828 VSS 0.111118f
C12028 DVSS.n829 VSS 0.098618f
C12029 DVSS.n830 VSS 0.014332f
C12030 DVSS.n831 VSS 0.014332f
C12031 DVSS.n832 VSS 0.014332f
C12032 DVSS.n833 VSS 0.014332f
C12033 DVSS.n834 VSS 0.014332f
C12034 DVSS.n835 VSS 0.014332f
C12035 DVSS.n836 VSS 0.014332f
C12036 DVSS.n837 VSS 0.014332f
C12037 DVSS.n838 VSS 0.014332f
C12038 DVSS.n839 VSS 0.014332f
C12039 DVSS.n840 VSS 0.014332f
C12040 DVSS.n841 VSS 0.014332f
C12041 DVSS.n842 VSS 0.014332f
C12042 DVSS.n843 VSS 0.014332f
C12043 DVSS.n844 VSS 0.014332f
C12044 DVSS.n845 VSS 0.014332f
C12045 DVSS.n846 VSS 0.014332f
C12046 DVSS.n847 VSS 0.014332f
C12047 DVSS.n848 VSS 0.023175f
C12048 DVSS.n849 VSS 0.04635f
C12049 DVSS.n850 VSS 0.023175f
C12050 DVSS.n851 VSS 0.04635f
C12051 DVSS.n852 VSS 0.023175f
C12052 DVSS.n853 VSS 0.04635f
C12053 DVSS.n854 VSS 0.04635f
C12054 DVSS.n855 VSS 0.429254f
C12055 DVSS.n856 VSS 0.421881f
C12056 DVSS.n857 VSS 0.092043f
C12057 DVSS.n858 VSS 0.092043f
C12058 DVSS.n859 VSS 0.092043f
C12059 DVSS.n860 VSS 0.092043f
C12060 DVSS.n861 VSS 0.092043f
C12061 DVSS.n862 VSS 0.092043f
C12062 DVSS.n863 VSS 0.092043f
C12063 DVSS.n864 VSS 0.092043f
C12064 DVSS.n865 VSS 0.092043f
C12065 DVSS.n866 VSS 0.092043f
C12066 DVSS.n867 VSS 0.092043f
C12067 DVSS.n868 VSS 0.092043f
C12068 DVSS.n869 VSS 0.092043f
C12069 DVSS.n870 VSS 0.092043f
C12070 DVSS.n871 VSS 0.092043f
C12071 DVSS.n872 VSS 0.092043f
C12072 DVSS.n873 VSS 0.092043f
C12073 DVSS.n874 VSS 0.092043f
C12074 DVSS.n875 VSS 0.092043f
C12075 DVSS.n876 VSS 0.092043f
C12076 DVSS.n877 VSS 0.092043f
C12077 DVSS.n878 VSS 0.092043f
C12078 DVSS.n879 VSS 0.092043f
C12079 DVSS.n880 VSS 0.092043f
C12080 DVSS.n881 VSS 0.092043f
C12081 DVSS.n882 VSS 0.092043f
C12082 DVSS.n883 VSS 0.092043f
C12083 DVSS.n884 VSS 0.092043f
C12084 DVSS.n885 VSS 0.092043f
C12085 DVSS.n886 VSS 0.092043f
C12086 DVSS.n887 VSS 0.092043f
C12087 DVSS.n888 VSS 0.092043f
C12088 DVSS.n889 VSS 0.092043f
C12089 DVSS.n890 VSS 0.092043f
C12090 DVSS.n891 VSS 0.092043f
C12091 DVSS.n892 VSS 0.092043f
C12092 DVSS.n893 VSS 0.092043f
C12093 DVSS.n894 VSS 0.092043f
C12094 DVSS.n895 VSS 0.092043f
C12095 DVSS.n896 VSS 0.092043f
C12096 DVSS.n897 VSS 0.092043f
C12097 DVSS.n898 VSS 0.092043f
C12098 DVSS.n899 VSS 0.092043f
C12099 DVSS.n900 VSS 0.092043f
C12100 DVSS.n901 VSS 0.092043f
C12101 DVSS.n902 VSS 0.092043f
C12102 DVSS.n903 VSS 0.092043f
C12103 DVSS.n904 VSS 0.092043f
C12104 DVSS.n905 VSS 0.092043f
C12105 DVSS.n906 VSS 0.092043f
C12106 DVSS.n907 VSS 0.092043f
C12107 DVSS.n908 VSS 0.092043f
C12108 DVSS.n909 VSS 0.092043f
C12109 DVSS.n910 VSS 0.092043f
C12110 DVSS.n911 VSS 0.092043f
C12111 DVSS.n912 VSS 0.092043f
C12112 DVSS.n913 VSS 0.092043f
C12113 DVSS.n914 VSS 0.092043f
C12114 DVSS.n915 VSS 0.092043f
C12115 DVSS.n916 VSS 0.092043f
C12116 DVSS.n917 VSS 0.092043f
C12117 DVSS.n918 VSS 0.092043f
C12118 DVSS.n919 VSS 0.092043f
C12119 DVSS.n920 VSS 0.092043f
C12120 DVSS.n921 VSS 0.092043f
C12121 DVSS.n922 VSS 0.092043f
C12122 DVSS.n923 VSS 0.092043f
C12123 DVSS.n924 VSS 0.092043f
C12124 DVSS.n925 VSS 0.092043f
C12125 DVSS.n926 VSS 0.092043f
C12126 DVSS.n927 VSS 0.092043f
C12127 DVSS.n928 VSS 0.092043f
C12128 DVSS.n929 VSS 0.092043f
C12129 DVSS.n930 VSS 0.092043f
C12130 DVSS.n931 VSS 0.092043f
C12131 DVSS.n932 VSS 0.092043f
C12132 DVSS.n933 VSS 0.092043f
C12133 DVSS.n934 VSS 0.092043f
C12134 DVSS.n935 VSS 0.092043f
C12135 DVSS.n936 VSS 0.092043f
C12136 DVSS.n937 VSS 0.092043f
C12137 DVSS.n938 VSS 0.092043f
C12138 DVSS.n939 VSS 0.092043f
C12139 DVSS.n940 VSS 0.092043f
C12140 DVSS.n941 VSS 0.092043f
C12141 DVSS.n942 VSS 0.092043f
C12142 DVSS.n943 VSS 0.092043f
C12143 DVSS.n944 VSS 0.092043f
C12144 DVSS.n945 VSS 0.092043f
C12145 DVSS.n946 VSS 0.092043f
C12146 DVSS.n947 VSS 0.092043f
C12147 DVSS.n948 VSS 0.092043f
C12148 DVSS.n949 VSS 0.569373f
C12149 DVSS.n950 VSS 0.092043f
C12150 DVSS.n951 VSS 0.046022f
C12151 DVSS.n952 VSS 0.047263f
C12152 DVSS.n953 VSS 0.158112f
C12153 DVSS.n954 VSS 0.442649f
C12154 DVSS.n955 VSS 0.448111f
C12155 DVSS.n956 VSS 2.40579f
C12156 DVSS.n957 VSS 2.06753f
C12157 DVSS.n958 VSS 3.45621f
C12158 DVSS.n959 VSS 4.38413f
C12159 DVSS.n960 VSS 6.06821f
C12160 DVSS.n961 VSS 4.18995f
C12161 DVSS.n962 VSS 1.5391f
C12162 DVSS.n963 VSS 0.835931f
C12163 DVSS.n964 VSS 0.029222f
C12164 DVSS.n965 VSS 0.012286f
C12165 DVSS.n966 VSS 0.789346f
C12166 DVSS.n967 VSS 0.012286f
C12167 DVSS.n968 VSS 0.029222f
C12168 DVSS.n969 VSS 0.012286f
C12169 DVSS.n970 VSS 0.789346f
C12170 DVSS.n971 VSS 0.012286f
C12171 DVSS.n972 VSS 0.029222f
C12172 DVSS.n973 VSS 0.012286f
C12173 DVSS.n974 VSS 0.789346f
C12174 DVSS.n975 VSS 0.012286f
C12175 DVSS.n976 VSS 0.029222f
C12176 DVSS.n977 VSS 0.012286f
C12177 DVSS.n978 VSS 0.789346f
C12178 DVSS.n979 VSS 0.012286f
C12179 DVSS.n980 VSS 0.029222f
C12180 DVSS.n981 VSS 0.012286f
C12181 DVSS.n982 VSS 0.789346f
C12182 DVSS.n983 VSS 0.012286f
C12183 DVSS.n984 VSS 0.029222f
C12184 DVSS.n985 VSS 0.012286f
C12185 DVSS.n986 VSS 0.789346f
C12186 DVSS.n987 VSS 0.012286f
C12187 DVSS.n988 VSS 0.029222f
C12188 DVSS.n989 VSS 0.012286f
C12189 DVSS.n990 VSS 0.789346f
C12190 DVSS.n991 VSS 0.012286f
C12191 DVSS.n992 VSS 0.029222f
C12192 DVSS.n993 VSS 0.012286f
C12193 DVSS.n994 VSS 0.789346f
C12194 DVSS.n995 VSS 0.012286f
C12195 DVSS.n996 VSS 0.029222f
C12196 DVSS.n997 VSS 0.012286f
C12197 DVSS.n998 VSS 0.789346f
C12198 DVSS.n999 VSS 0.012286f
C12199 DVSS.n1000 VSS 0.029222f
C12200 DVSS.n1001 VSS 0.012286f
C12201 DVSS.n1002 VSS 0.789346f
C12202 DVSS.n1003 VSS 0.012286f
C12203 DVSS.n1004 VSS 0.029222f
C12204 DVSS.n1005 VSS 0.012286f
C12205 DVSS.n1006 VSS 0.789346f
C12206 DVSS.n1007 VSS 0.012286f
C12207 DVSS.n1008 VSS 0.029222f
C12208 DVSS.n1009 VSS 0.012286f
C12209 DVSS.n1010 VSS 0.789346f
C12210 DVSS.n1011 VSS 0.012286f
C12211 DVSS.n1012 VSS 0.029222f
C12212 DVSS.n1013 VSS 0.012286f
C12213 DVSS.n1014 VSS 0.789346f
C12214 DVSS.n1015 VSS 0.012286f
C12215 DVSS.n1016 VSS 0.029222f
C12216 DVSS.n1017 VSS 0.012286f
C12217 DVSS.n1018 VSS 0.789346f
C12218 DVSS.n1019 VSS 0.012286f
C12219 DVSS.n1020 VSS 0.022034f
C12220 DVSS.n1021 VSS 0.012286f
C12221 DVSS.n1022 VSS 0.588827f
C12222 DVSS.n1023 VSS 1.59219f
C12223 DVSS.n1024 VSS 1.59455f
C12224 DVSS.n1025 VSS 0.029222f
C12225 DVSS.n1026 VSS 0.012286f
C12226 DVSS.n1027 VSS 0.789346f
C12227 DVSS.n1028 VSS 0.012286f
C12228 DVSS.n1029 VSS 0.029222f
C12229 DVSS.n1030 VSS 0.012286f
C12230 DVSS.n1031 VSS 0.789346f
C12231 DVSS.n1032 VSS 0.012286f
C12232 DVSS.n1033 VSS 0.029222f
C12233 DVSS.n1034 VSS 0.012286f
C12234 DVSS.n1035 VSS 0.789346f
C12235 DVSS.n1036 VSS 0.012286f
C12236 DVSS.n1037 VSS 0.029222f
C12237 DVSS.n1038 VSS 0.012286f
C12238 DVSS.n1039 VSS 0.789346f
C12239 DVSS.n1040 VSS 0.012286f
C12240 DVSS.n1041 VSS 0.029222f
C12241 DVSS.n1042 VSS 0.012286f
C12242 DVSS.n1043 VSS 0.789346f
C12243 DVSS.n1044 VSS 0.012286f
C12244 DVSS.n1045 VSS 0.029222f
C12245 DVSS.n1046 VSS 0.012286f
C12246 DVSS.n1047 VSS 0.789346f
C12247 DVSS.n1048 VSS 0.012286f
C12248 DVSS.n1049 VSS 0.029222f
C12249 DVSS.n1050 VSS 0.012286f
C12250 DVSS.n1051 VSS 0.789346f
C12251 DVSS.n1052 VSS 0.012286f
C12252 DVSS.n1053 VSS 0.029222f
C12253 DVSS.n1054 VSS 0.012286f
C12254 DVSS.n1055 VSS 0.789346f
C12255 DVSS.n1056 VSS 0.012286f
C12256 DVSS.n1057 VSS 0.029222f
C12257 DVSS.n1058 VSS 0.012286f
C12258 DVSS.n1059 VSS 0.789346f
C12259 DVSS.n1060 VSS 0.012286f
C12260 DVSS.n1061 VSS 0.029222f
C12261 DVSS.n1062 VSS 0.012286f
C12262 DVSS.n1063 VSS 0.789346f
C12263 DVSS.n1064 VSS 0.012286f
C12264 DVSS.n1065 VSS 0.029222f
C12265 DVSS.n1066 VSS 0.012286f
C12266 DVSS.n1067 VSS 0.789346f
C12267 DVSS.n1068 VSS 0.012286f
C12268 DVSS.n1069 VSS 0.029222f
C12269 DVSS.n1070 VSS 0.012286f
C12270 DVSS.n1071 VSS 0.789346f
C12271 DVSS.n1072 VSS 0.012286f
C12272 DVSS.n1073 VSS 0.029222f
C12273 DVSS.n1074 VSS 0.012286f
C12274 DVSS.n1075 VSS 0.789346f
C12275 DVSS.n1076 VSS 0.012286f
C12276 DVSS.n1077 VSS 0.029222f
C12277 DVSS.n1078 VSS 0.012286f
C12278 DVSS.n1079 VSS 0.690678f
C12279 DVSS.n1080 VSS 0.012286f
C12280 DVSS.n1081 VSS 0.81518f
C12281 DVSS.n1082 VSS 0.092043f
C12282 DVSS.n1083 VSS 0.092043f
C12283 DVSS.n1084 VSS 0.092043f
C12284 DVSS.n1085 VSS 0.092043f
C12285 DVSS.n1086 VSS 0.092043f
C12286 DVSS.n1087 VSS 0.092043f
C12287 DVSS.n1088 VSS 0.092043f
C12288 DVSS.n1089 VSS 0.092043f
C12289 DVSS.n1090 VSS 0.092043f
C12290 DVSS.n1091 VSS 0.092043f
C12291 DVSS.n1092 VSS 0.092043f
C12292 DVSS.n1093 VSS 0.092043f
C12293 DVSS.n1094 VSS 0.092043f
C12294 DVSS.n1095 VSS 0.092043f
C12295 DVSS.n1096 VSS 0.092043f
C12296 DVSS.n1097 VSS 0.092043f
C12297 DVSS.n1098 VSS 0.538002f
C12298 DVSS.n1099 VSS 0.058279f
C12299 DVSS.n1100 VSS 0.092043f
C12300 DVSS.n1101 VSS 0.092043f
C12301 DVSS.n1102 VSS 0.092043f
C12302 DVSS.n1103 VSS 0.049587f
C12303 DVSS.n1104 VSS 0.092043f
C12304 DVSS.n1105 VSS 0.092043f
C12305 DVSS.n1106 VSS 0.092043f
C12306 DVSS.n1107 VSS 0.092043f
C12307 DVSS.n1108 VSS 0.046022f
C12308 DVSS.n1109 VSS 0.004997f
C12309 DVSS.n1110 VSS 0.046022f
C12310 DVSS.n1111 VSS 0.092043f
C12311 DVSS.n1112 VSS 0.092043f
C12312 DVSS.n1113 VSS 0.092043f
C12313 DVSS.n1114 VSS 0.092043f
C12314 DVSS.n1115 VSS 0.092043f
C12315 DVSS.n1116 VSS 0.046022f
C12316 DVSS.n1117 VSS 0.046022f
C12317 DVSS.n1118 VSS 0.046022f
C12318 DVSS.n1119 VSS 0.004082f
C12319 DVSS.n1120 VSS 0.002498f
C12320 DVSS.n1121 VSS 0.011882f
C12321 DVSS.n1122 VSS 0.046022f
C12322 DVSS.n1123 VSS 0.092043f
C12323 DVSS.n1124 VSS 0.092043f
C12324 DVSS.n1125 VSS 0.092043f
C12325 DVSS.n1126 VSS 0.046022f
C12326 DVSS.n1127 VSS 0.046279f
C12327 DVSS.n1128 VSS 0.092043f
C12328 DVSS.n1129 VSS 0.092043f
C12329 DVSS.n1130 VSS 0.092043f
C12330 DVSS.n1131 VSS 0.092043f
C12331 DVSS.n1132 VSS 0.092043f
C12332 DVSS.n1133 VSS 0.092043f
C12333 DVSS.n1134 VSS 0.092043f
C12334 DVSS.n1135 VSS 0.092043f
C12335 DVSS.n1136 VSS 0.092043f
C12336 DVSS.n1137 VSS 0.092043f
C12337 DVSS.n1138 VSS 0.092043f
C12338 DVSS.n1139 VSS 0.092043f
C12339 DVSS.n1140 VSS 0.092043f
C12340 DVSS.n1141 VSS 0.092043f
C12341 DVSS.n1142 VSS 0.092043f
C12342 DVSS.n1143 VSS 0.092043f
C12343 DVSS.n1144 VSS 0.092043f
C12344 DVSS.n1145 VSS 0.092043f
C12345 DVSS.n1146 VSS 0.092043f
C12346 DVSS.n1147 VSS 0.092043f
C12347 DVSS.n1148 VSS 0.092043f
C12348 DVSS.n1149 VSS 0.092043f
C12349 DVSS.n1150 VSS 0.092043f
C12350 DVSS.n1151 VSS 0.092043f
C12351 DVSS.n1152 VSS 0.092043f
C12352 DVSS.n1153 VSS 0.092043f
C12353 DVSS.n1154 VSS 0.092043f
C12354 DVSS.n1155 VSS 0.092043f
C12355 DVSS.n1156 VSS 0.080621f
C12356 DVSS.n1157 VSS 0.092043f
C12357 DVSS.n1158 VSS 0.092043f
C12358 DVSS.n1159 VSS 0.092043f
C12359 DVSS.n1160 VSS 0.060282f
C12360 DVSS.n1161 VSS 0.092043f
C12361 DVSS.n1162 VSS 0.092043f
C12362 DVSS.n1163 VSS 0.092043f
C12363 DVSS.n1164 VSS 0.092043f
C12364 DVSS.n1165 VSS 0.092043f
C12365 DVSS.n1166 VSS 0.092043f
C12366 DVSS.n1167 VSS 0.092043f
C12367 DVSS.n1168 VSS 0.092043f
C12368 DVSS.n1169 VSS 0.092043f
C12369 DVSS.n1170 VSS 0.092043f
C12370 DVSS.n1171 VSS 0.092043f
C12371 DVSS.n1172 VSS 0.092043f
C12372 DVSS.n1173 VSS 0.092043f
C12373 DVSS.n1174 VSS 0.092043f
C12374 DVSS.n1175 VSS 0.092043f
C12375 DVSS.n1176 VSS 0.092043f
C12376 DVSS.n1177 VSS 0.092043f
C12377 DVSS.n1178 VSS 0.092043f
C12378 DVSS.n1179 VSS 0.092043f
C12379 DVSS.n1180 VSS 0.092043f
C12380 DVSS.n1181 VSS 0.092043f
C12381 DVSS.n1182 VSS 0.092043f
C12382 DVSS.n1183 VSS 0.092043f
C12383 DVSS.n1184 VSS 0.092043f
C12384 DVSS.n1185 VSS 0.092043f
C12385 DVSS.n1186 VSS 0.092043f
C12386 DVSS.n1187 VSS 0.092043f
C12387 DVSS.n1188 VSS 0.092043f
C12388 DVSS.n1189 VSS 0.092043f
C12389 DVSS.n1190 VSS 0.092043f
C12390 DVSS.n1191 VSS 0.092043f
C12391 DVSS.n1192 VSS 0.092043f
C12392 DVSS.n1193 VSS 0.046022f
C12393 DVSS.n1194 VSS 0.082968f
C12394 DVSS.n1195 VSS 0.092043f
C12395 DVSS.n1196 VSS 1.22564f
C12396 DVSS.n1197 VSS 0.026298f
C12397 DVSS.n1198 VSS 0.026298f
C12398 DVSS.n1199 VSS 0.083292f
C12399 DVSS.n1201 VSS 0.026298f
C12400 DVSS.n1202 VSS 2.23352f
C12401 DVSS.n1203 VSS 0.400772f
C12402 DVSS.n1204 VSS 0.478809f
C12403 DVSS.n1205 VSS 0.159008f
C12404 DVSS.t198 VSS 0.17128f
C12405 DVSS.t166 VSS 0.007223f
C12406 DVSS.t199 VSS 0.007223f
C12407 DVSS.n1206 VSS 0.015027f
C12408 DVSS.n1207 VSS 0.006767f
C12409 DVSS.n1208 VSS 0.010533f
C12410 DVSS.n1209 VSS 0.3096f
C12411 DVSS.t72 VSS 0.17128f
C12412 DVSS.n1210 VSS 0.076841f
C12413 DVSS.t84 VSS 0.007223f
C12414 DVSS.t73 VSS 0.007223f
C12415 DVSS.n1211 VSS 0.015027f
C12416 DVSS.n1212 VSS 0.006767f
C12417 DVSS.n1213 VSS 0.323888f
C12418 DVSS.n1214 VSS 0.463646f
C12419 DVSS.n1215 VSS 0.296597f
C12420 DVSS.n1216 VSS 0.317423f
C12421 DVSS.n1217 VSS 0.740632f
C12422 DVSS.n1218 VSS 0.286047f
C12423 DVSS.t146 VSS 0.144516f
C12424 DVSS.t189 VSS 0.007223f
C12425 DVSS.t147 VSS 0.007223f
C12426 DVSS.n1219 VSS 0.015027f
C12427 DVSS.n1220 VSS 0.006767f
C12428 DVSS.n1221 VSS 0.010533f
C12429 DVSS.n1222 VSS 0.19732f
C12430 DVSS.n1223 VSS 0.04967f
C12431 DVSS.t163 VSS 0.014445f
C12432 DVSS.n1224 VSS 0.038498f
C12433 DVSS.n1225 VSS 0.012005f
C12434 DVSS.n1226 VSS 0.010866f
C12435 DVSS.t71 VSS 0.014445f
C12436 DVSS.t37 VSS 0.014445f
C12437 DVSS.n1227 VSS 0.032942f
C12438 DVSS.n1228 VSS 0.012058f
C12439 DVSS.n1229 VSS 0.02551f
C12440 DVSS.t65 VSS 0.014445f
C12441 DVSS.t206 VSS 0.01434f
C12442 DVSS.n1230 VSS 0.683214f
C12443 DVSS.t9 VSS 0.014445f
C12444 DVSS.t168 VSS 0.014445f
C12445 DVSS.n1231 VSS 0.032684f
C12446 DVSS.n1232 VSS 0.020331f
C12447 DVSS.n1233 VSS 0.021032f
C12448 DVSS.t82 VSS 0.207452f
C12449 DVSS.n1234 VSS 0.049402f
C12450 DVSS.n1235 VSS 0.18404f
C12451 DVSS.n1236 VSS 0.197235f
C12452 DVSS.n1237 VSS 0.197235f
C12453 DVSS.n1238 VSS 0.197235f
C12454 DVSS.n1239 VSS 0.197235f
C12455 DVSS.n1240 VSS 0.197235f
C12456 DVSS.n1241 VSS 0.197235f
C12457 DVSS.n1242 VSS 0.197235f
C12458 DVSS.n1243 VSS 0.197235f
C12459 DVSS.n1244 VSS 0.197235f
C12460 DVSS.n1245 VSS 0.197235f
C12461 DVSS.n1246 VSS 0.197235f
C12462 DVSS.n1247 VSS 0.197235f
C12463 DVSS.n1248 VSS 0.178484f
C12464 DVSS.n1249 VSS 0.078841f
C12465 DVSS.n1250 VSS 0.025192f
C12466 DVSS.n1251 VSS 0.024059f
C12467 DVSS.t129 VSS 0.014445f
C12468 DVSS.t18 VSS 0.014445f
C12469 DVSS.n1252 VSS 0.032684f
C12470 DVSS.n1253 VSS 0.020331f
C12471 DVSS.t34 VSS 0.55148f
C12472 DVSS.n1254 VSS 0.082172f
C12473 DVSS.n1255 VSS 0.024059f
C12474 DVSS.t29 VSS 0.251375f
C12475 DVSS.n1256 VSS 0.643209f
C12476 DVSS.t35 VSS 0.579185f
C12477 DVSS.n1257 VSS 0.124391f
C12478 DVSS.n1258 VSS 0.032165f
C12479 DVSS.n1259 VSS 0.060171f
C12480 DVSS.n1260 VSS 0.032165f
C12481 DVSS.n1261 VSS 0.124391f
C12482 DVSS.n1262 VSS 0.683214f
C12483 DVSS.n1263 VSS 0.070246f
C12484 DVSS.t31 VSS 0.308812f
C12485 DVSS.t126 VSS 0.345302f
C12486 DVSS.n1264 VSS 0.018424f
C12487 DVSS.n1265 VSS 0.002551f
C12488 DVSS.t127 VSS 0.014445f
C12489 DVSS.n1266 VSS 0.038498f
C12490 DVSS.n1267 VSS 0.009596f
C12491 DVSS.n1268 VSS 0.035876f
C12492 DVSS.t157 VSS 0.014445f
C12493 DVSS.t153 VSS 0.014445f
C12494 DVSS.n1269 VSS 0.032942f
C12495 DVSS.n1270 VSS 0.012058f
C12496 DVSS.t155 VSS 0.014445f
C12497 DVSS.t207 VSS 0.01434f
C12498 DVSS.n1271 VSS 0.026861f
C12499 DVSS.n1272 VSS 0.018385f
C12500 DVSS.t121 VSS 0.014445f
C12501 DVSS.n1273 VSS 0.028891f
C12502 DVSS.n1274 VSS 0.012058f
C12503 DVSS.n1275 VSS 0.075164f
C12504 DVSS.n1276 VSS 0.165289f
C12505 DVSS.n1277 VSS 0.247165f
C12506 DVSS.n1278 VSS 0.197235f
C12507 DVSS.n1279 VSS 0.197235f
C12508 DVSS.n1280 VSS 0.197235f
C12509 DVSS.n1281 VSS 0.197235f
C12510 DVSS.n1282 VSS 0.197235f
C12511 DVSS.n1283 VSS 0.197235f
C12512 DVSS.n1284 VSS 0.197235f
C12513 DVSS.n1285 VSS 0.197235f
C12514 DVSS.n1286 VSS 0.197235f
C12515 DVSS.n1287 VSS 0.197235f
C12516 DVSS.n1288 VSS 0.197235f
C12517 DVSS.n1289 VSS 0.197235f
C12518 DVSS.n1290 VSS 0.197235f
C12519 DVSS.n1291 VSS 0.197235f
C12520 DVSS.n1292 VSS 0.197235f
C12521 DVSS.n1293 VSS 0.197235f
C12522 DVSS.n1294 VSS 0.197235f
C12523 DVSS.n1295 VSS 0.197235f
C12524 DVSS.n1296 VSS 0.197235f
C12525 DVSS.n1297 VSS 0.197235f
C12526 DVSS.n1298 VSS 0.197235f
C12527 DVSS.n1299 VSS 0.197235f
C12528 DVSS.n1300 VSS 0.197235f
C12529 DVSS.n1301 VSS 0.197235f
C12530 DVSS.n1302 VSS 0.197235f
C12531 DVSS.n1303 VSS 0.197235f
C12532 DVSS.n1304 VSS 0.197235f
C12533 DVSS.n1305 VSS 0.197235f
C12534 DVSS.n1306 VSS 0.197235f
C12535 DVSS.n1307 VSS 0.197235f
C12536 DVSS.n1308 VSS 0.197235f
C12537 DVSS.n1309 VSS 0.197235f
C12538 DVSS.n1310 VSS 0.149315f
C12539 DVSS.n1311 VSS 0.105248f
C12540 DVSS.n1312 VSS 0.146537f
C12541 DVSS.n1313 VSS 0.197235f
C12542 DVSS.n1314 VSS 0.197235f
C12543 DVSS.n1315 VSS 0.197235f
C12544 DVSS.n1316 VSS 0.197235f
C12545 DVSS.n1317 VSS 0.197235f
C12546 DVSS.n1318 VSS 0.197235f
C12547 DVSS.n1319 VSS 0.197235f
C12548 DVSS.n1320 VSS 0.197235f
C12549 DVSS.n1321 VSS 0.197235f
C12550 DVSS.n1322 VSS 0.197235f
C12551 DVSS.n1323 VSS 0.197235f
C12552 DVSS.n1324 VSS 0.197235f
C12553 DVSS.n1325 VSS 0.197235f
C12554 DVSS.n1326 VSS 0.197235f
C12555 DVSS.n1327 VSS 0.197235f
C12556 DVSS.n1328 VSS 0.197235f
C12557 DVSS.n1329 VSS 0.197235f
C12558 DVSS.n1330 VSS 0.197235f
C12559 DVSS.n1331 VSS 0.197235f
C12560 DVSS.n1332 VSS 0.197235f
C12561 DVSS.n1333 VSS 0.197235f
C12562 DVSS.n1334 VSS 0.197235f
C12563 DVSS.n1335 VSS 0.197235f
C12564 DVSS.n1336 VSS 0.197235f
C12565 DVSS.n1337 VSS 0.197235f
C12566 DVSS.n1338 VSS 0.197235f
C12567 DVSS.n1339 VSS 0.197235f
C12568 DVSS.n1340 VSS 0.197235f
C12569 DVSS.n1341 VSS 0.17779f
C12570 DVSS.n1342 VSS 0.17779f
C12571 DVSS.n1343 VSS 0.17779f
C12572 DVSS.n1344 VSS 0.009557f
C12573 DVSS.t98 VSS 0.014445f
C12574 DVSS.n1345 VSS 0.038498f
C12575 DVSS.n1346 VSS 0.002551f
C12576 DVSS.n1347 VSS 0.032017f
C12577 DVSS.n1348 VSS 0.126367f
C12578 DVSS.n1349 VSS 0.038197f
C12579 DVSS.n1350 VSS 0.118063f
C12580 DVSS.n1351 VSS 0.022224f
C12581 DVSS.n1352 VSS 0.194457f
C12582 DVSS.n1353 VSS 0.736605f
C12583 DVSS.n1354 VSS 0.046022f
C12584 DVSS.n1355 VSS 0.046022f
C12585 DVSS.n1356 VSS 0.02426f
C12586 DVSS.n1357 VSS 0.116674f
C12587 DVSS.n1358 VSS 0.079403f
C12588 DVSS.n1359 VSS 0.018451f
C12589 DVSS.n1360 VSS 0.018451f
C12590 DVSS.n1361 VSS 0.018451f
C12591 DVSS.n1362 VSS 0.018451f
C12592 DVSS.n1363 VSS 0.018451f
C12593 DVSS.n1364 VSS 0.018451f
C12594 DVSS.n1365 VSS 0.018451f
C12595 DVSS.n1366 VSS 0.018451f
C12596 DVSS.n1367 VSS 0.034602f
C12597 DVSS.n1368 VSS 0.023175f
C12598 DVSS.n1369 VSS 0.056768f
C12599 DVSS.n1370 VSS 3.35583f
C12600 DVSS.n1371 VSS 1.30625f
C12601 DVSS.n1372 VSS 0.02033f
C12602 DVSS.n1373 VSS 0.022381f
C12603 DVSS.n1374 VSS 0.034602f
C12604 DVSS.n1375 VSS 0.02426f
C12605 DVSS.n1376 VSS 0.034602f
C12606 DVSS.n1377 VSS 0.02426f
C12607 DVSS.n1378 VSS 0.034602f
C12608 DVSS.n1379 VSS 0.034602f
C12609 DVSS.n1380 VSS 0.021356f
C12610 DVSS.n1381 VSS 0.021356f
C12611 DVSS.n1382 VSS 0.034602f
C12612 DVSS.n1383 VSS 0.02426f
C12613 DVSS.n1384 VSS 0.034602f
C12614 DVSS.n1385 VSS 0.02426f
C12615 DVSS.n1386 VSS 0.034602f
C12616 DVSS.n1387 VSS 0.034602f
C12617 DVSS.n1388 VSS 0.022381f
C12618 DVSS.n1389 VSS 0.02033f
C12619 DVSS.n1390 VSS 0.034602f
C12620 DVSS.n1391 VSS 0.119037f
C12621 DVSS.n1392 VSS 0.188185f
C12622 DVSS.n1393 VSS 2.06082f
C12623 DVSS.n1394 VSS 1.33188f
C12624 DVSS.n1395 VSS 0.068967f
C12625 DVSS.n1396 VSS 0.259592f
C12626 DVSS.n1397 VSS 0.023539f
C12627 DVSS.n1398 VSS 0.026956f
C12628 DVSS.n1399 VSS 0.046022f
C12629 DVSS.n1400 VSS 0.046022f
C12630 DVSS.n1401 VSS 0.092043f
C12631 DVSS.n1402 VSS 0.092043f
C12632 DVSS.n1403 VSS 0.092043f
C12633 DVSS.n1404 VSS 0.092043f
C12634 DVSS.n1405 VSS 0.046022f
C12635 DVSS.n1406 VSS 0.042497f
C12636 DVSS.n1407 VSS 0.051531f
C12637 DVSS.n1408 VSS 0.046022f
C12638 DVSS.n1409 VSS 0.092043f
C12639 DVSS.n1410 VSS 0.092043f
C12640 DVSS.n1411 VSS 0.092043f
C12641 DVSS.n1412 VSS 0.092043f
C12642 DVSS.n1413 VSS 0.092043f
C12643 DVSS.n1414 VSS 0.092043f
C12644 DVSS.n1415 VSS 0.092043f
C12645 DVSS.n1416 VSS 0.046022f
C12646 DVSS.n1417 VSS 0.042497f
C12647 DVSS.n1418 VSS 0.066064f
C12648 DVSS.n1419 VSS 0.026956f
C12649 DVSS.n1420 VSS 0.046022f
C12650 DVSS.n1421 VSS 0.046022f
C12651 DVSS.n1422 VSS 0.092043f
C12652 DVSS.n1423 VSS 0.092043f
C12653 DVSS.n1424 VSS 0.092043f
C12654 DVSS.n1425 VSS 0.092043f
C12655 DVSS.n1426 VSS 0.046022f
C12656 DVSS.n1427 VSS 0.023539f
C12657 DVSS.n1428 VSS 0.051772f
C12658 DVSS.n1429 VSS 0.046205f
C12659 DVSS.n1430 VSS 0.092043f
C12660 DVSS.n1431 VSS 0.092043f
C12661 DVSS.n1432 VSS 0.092043f
C12662 DVSS.n1433 VSS 0.092043f
C12663 DVSS.n1434 VSS 0.092043f
C12664 DVSS.n1435 VSS 0.092043f
C12665 DVSS.n1436 VSS 0.092043f
C12666 DVSS.n1437 VSS 0.046022f
C12667 DVSS.n1438 VSS 0.042497f
C12668 DVSS.n1439 VSS 0.066064f
C12669 DVSS.n1440 VSS 0.026956f
C12670 DVSS.n1441 VSS 0.046022f
C12671 DVSS.n1442 VSS 0.046022f
C12672 DVSS.n1443 VSS 0.092043f
C12673 DVSS.n1444 VSS 0.092043f
C12674 DVSS.n1445 VSS 0.092043f
C12675 DVSS.n1446 VSS 0.046022f
C12676 DVSS.n1447 VSS 0.023539f
C12677 DVSS.n1448 VSS 0.253973f
C12678 DVSS.n1449 VSS 1.33226f
C12679 DVSS.n1450 VSS 4.18995f
C12680 DVSS.n1451 VSS 1.46105f
C12681 DVSS.t200 VSS 0.658108f
C12682 DVSS.n1452 VSS 0.070246f
C12683 DVSS.t201 VSS 0.014445f
C12684 DVSS.n1453 VSS 0.038498f
C12685 DVSS.n1454 VSS 0.012005f
C12686 DVSS.n1455 VSS 0.137761f
C12687 DVSS.t123 VSS 0.014445f
C12688 DVSS.t204 VSS 0.01434f
C12689 DVSS.n1456 VSS 0.026861f
C12690 DVSS.n1457 VSS 0.018385f
C12691 DVSS.t125 VSS 0.014445f
C12692 DVSS.n1458 VSS 0.028891f
C12693 DVSS.n1459 VSS 0.012058f
C12694 DVSS.t203 VSS 0.014445f
C12695 DVSS.t161 VSS 0.014445f
C12696 DVSS.n1460 VSS 0.032942f
C12697 DVSS.n1461 VSS 0.012058f
C12698 DVSS.n1462 VSS 0.035876f
C12699 DVSS.t118 VSS 0.192835f
C12700 DVSS.n1463 VSS 0.86139f
C12701 DVSS.t11 VSS 0.257861f
C12702 DVSS.n1464 VSS 0.683214f
C12703 DVSS.t6 VSS 0.014445f
C12704 DVSS.t1 VSS 0.014445f
C12705 DVSS.n1465 VSS 0.032684f
C12706 DVSS.n1466 VSS 0.020331f
C12707 DVSS.n1467 VSS 0.024059f
C12708 DVSS.n1468 VSS 0.02356f
C12709 DVSS.n1469 VSS 0.024059f
C12710 DVSS.t107 VSS 0.014445f
C12711 DVSS.t24 VSS 0.014445f
C12712 DVSS.n1470 VSS 0.032684f
C12713 DVSS.n1471 VSS 0.020331f
C12714 DVSS.n1472 VSS 0.683214f
C12715 DVSS.n1473 VSS 0.049774f
C12716 DVSS.t112 VSS 0.163686f
C12717 DVSS.t23 VSS 0.526935f
C12718 DVSS.t43 VSS 0.007223f
C12719 DVSS.t172 VSS 0.007223f
C12720 DVSS.n1474 VSS 0.015027f
C12721 DVSS.n1475 VSS 0.006767f
C12722 DVSS.n1476 VSS 0.011305f
C12723 DVSS.t42 VSS 0.273557f
C12724 DVSS.n1477 VSS -0.001195f
C12725 DVSS.t188 VSS 0.136778f
C12726 DVSS.t40 VSS 0.301586f
C12727 DVSS.t38 VSS 0.368854f
C12728 DVSS.t41 VSS 0.014445f
C12729 DVSS.t205 VSS 0.01434f
C12730 DVSS.n1478 VSS 0.026861f
C12731 DVSS.n1479 VSS 0.018385f
C12732 DVSS.t75 VSS 0.014445f
C12733 DVSS.n1480 VSS 0.028891f
C12734 DVSS.n1481 VSS 0.012058f
C12735 DVSS.n1482 VSS 0.023245f
C12736 DVSS.n1483 VSS 0.007702f
C12737 DVSS.n1484 VSS 0.120841f
C12738 DVSS.n1485 VSS 0.197235f
C12739 DVSS.n1486 VSS 0.197235f
C12740 DVSS.n1487 VSS 0.197235f
C12741 DVSS.n1488 VSS 0.197235f
C12742 DVSS.n1489 VSS 0.197235f
C12743 DVSS.n1490 VSS 0.197235f
C12744 DVSS.n1491 VSS 0.197235f
C12745 DVSS.n1492 VSS 0.197235f
C12746 DVSS.n1493 VSS 0.197235f
C12747 DVSS.n1494 VSS 0.197235f
C12748 DVSS.n1495 VSS 0.197235f
C12749 DVSS.n1496 VSS 0.197235f
C12750 DVSS.n1497 VSS 0.114591f
C12751 DVSS.t47 VSS 0.014445f
C12752 DVSS.t39 VSS 0.014445f
C12753 DVSS.n1498 VSS 0.032942f
C12754 DVSS.n1499 VSS 0.01122f
C12755 DVSS.n1500 VSS 0.019546f
C12756 DVSS.n1501 VSS -0.047203f
C12757 DVSS.n1502 VSS 0.060171f
C12758 DVSS.n1503 VSS 0.018785f
C12759 DVSS.n1504 VSS 0.032165f
C12760 DVSS.n1505 VSS 0.124391f
C12761 DVSS.t30 VSS 0.584739f
C12762 DVSS.n1506 VSS 0.435595f
C12763 DVSS.n1507 VSS 0.504893f
C12764 DVSS.t33 VSS 0.383429f
C12765 DVSS.n1508 VSS 0.032165f
C12766 DVSS.n1509 VSS 0.124391f
C12767 DVSS.t32 VSS 0.554468f
C12768 DVSS.n1510 VSS 0.273557f
C12769 DVSS.n1511 VSS 0.033005f
C12770 DVSS.n1512 VSS 0.033796f
C12771 DVSS.n1513 VSS 0.014344f
C12772 DVSS.n1514 VSS 0.02426f
C12773 DVSS.n1515 VSS 0.016369f
C12774 DVSS.n1516 VSS 0.003835f
C12775 DVSS.t28 VSS 0.348674f
C12776 DVSS.n1517 VSS 0.08583f
C12777 DVSS.n1518 VSS 0.251518f
C12778 DVSS.n1519 VSS 0.052887f
C12779 DVSS.n1520 VSS 0.04732f
C12780 DVSS.n1521 VSS 0.051726f
C12781 DVSS.n1522 VSS -0.17564f
C12782 DVSS.n1523 VSS 0.696328f
C12783 DVSS.n1524 VSS 1.42696f
C12784 DVSS.n1525 VSS 0.018401f
C12785 DVSS.n1526 VSS 0.01116f
C12786 DVSS.n1527 VSS 0.046022f
C12787 DVSS.n1528 VSS 0.046022f
C12788 DVSS.n1529 VSS 0.046022f
C12789 DVSS.n1530 VSS 0.011671f
C12790 DVSS.n1531 VSS 0.009201f
C12791 DVSS.n1532 VSS 0.009201f
C12792 DVSS.n1533 VSS 0.009201f
C12793 DVSS.n1534 VSS 0.050235f
C12794 DVSS.n1535 VSS 0.009201f
C12795 DVSS.n1536 VSS 0.009201f
C12796 DVSS.n1537 VSS 0.01116f
C12797 DVSS.n1538 VSS 0.010267f
C12798 DVSS.n1539 VSS 0.234615f
C12799 DVSS.n1540 VSS 0.68664f
C12800 DVSS.n1541 VSS 0.170167f
C12801 DVSS.n1542 VSS 0.052887f
C12802 DVSS.n1543 VSS 0.051726f
C12803 DVSS.n1544 VSS 0.052887f
C12804 DVSS.n1545 VSS 0.068934f
C12805 DVSS.n1546 VSS 0.052887f
C12806 DVSS.n1547 VSS 0.127793f
C12807 DVSS.n1548 VSS 0.305067f
C12808 DVSS.n1549 VSS 0.689543f
C12809 DVSS.n1550 VSS 0.01735f
C12810 DVSS.t57 VSS 0.037108f
C12811 DVSS.n1551 VSS 0.071349f
C12812 DVSS.t53 VSS 0.037108f
C12813 DVSS.n1552 VSS 0.184323f
C12814 DVSS.n1553 VSS 0.647257f
C12815 DVSS.n1554 VSS 0.421806f
C12816 DVSS.n1555 VSS 0.035931f
C12817 DVSS.n1556 VSS 0.007344f
C12818 DVSS.n1557 VSS 0.068384f
C12819 DVSS.n1558 VSS 0.092043f
C12820 DVSS.n1559 VSS 0.092043f
C12821 DVSS.n1560 VSS 0.092043f
C12822 DVSS.n1561 VSS 0.092043f
C12823 DVSS.n1562 VSS 0.092043f
C12824 DVSS.n1563 VSS 0.092043f
C12825 DVSS.n1564 VSS 0.092043f
C12826 DVSS.n1565 VSS 0.092043f
C12827 DVSS.n1566 VSS 0.092043f
C12828 DVSS.n1567 VSS 0.092043f
C12829 DVSS.n1568 VSS 0.092043f
C12830 DVSS.n1569 VSS 0.341066f
C12831 DVSS.n1570 VSS 0.092043f
C12832 DVSS.n1571 VSS 0.195546f
C12833 DVSS.n1572 VSS 0.173028f
C12834 DVSS.n1573 VSS 0.092043f
C12835 DVSS.n1574 VSS 0.092043f
C12836 DVSS.n1575 VSS 0.092043f
C12837 DVSS.n1576 VSS 0.092043f
C12838 DVSS.n1577 VSS 0.092043f
C12839 DVSS.n1578 VSS 0.092043f
C12840 DVSS.n1579 VSS 0.092043f
C12841 DVSS.n1580 VSS 0.092043f
C12842 DVSS.n1581 VSS 0.092043f
C12843 DVSS.n1582 VSS 0.092043f
C12844 DVSS.n1583 VSS 0.092043f
C12845 DVSS.n1584 VSS 0.092043f
C12846 DVSS.n1585 VSS 0.092043f
C12847 DVSS.n1586 VSS 0.092043f
C12848 DVSS.n1587 VSS 0.092043f
C12849 DVSS.n1588 VSS 0.092043f
C12850 DVSS.n1589 VSS 0.092043f
C12851 DVSS.n1590 VSS 0.092043f
C12852 DVSS.n1591 VSS 0.092043f
C12853 DVSS.n1592 VSS 0.092043f
C12854 DVSS.n1593 VSS 0.092043f
C12855 DVSS.n1594 VSS 0.092043f
C12856 DVSS.n1595 VSS 0.092043f
C12857 DVSS.n1596 VSS 0.092043f
C12858 DVSS.n1597 VSS 0.092043f
C12859 DVSS.n1598 VSS 0.092043f
C12860 DVSS.n1599 VSS 0.092043f
C12861 DVSS.n1600 VSS 0.092043f
C12862 DVSS.n1601 VSS 0.092043f
C12863 DVSS.n1602 VSS 0.092043f
C12864 DVSS.n1603 VSS 0.092043f
C12865 DVSS.n1604 VSS 0.092043f
C12866 DVSS.n1605 VSS 0.092043f
C12867 DVSS.n1606 VSS 0.092043f
C12868 DVSS.n1607 VSS 0.092043f
C12869 DVSS.n1608 VSS 0.092043f
C12870 DVSS.n1609 VSS 0.092043f
C12871 DVSS.n1610 VSS 0.059634f
C12872 DVSS.t133 VSS 0.35047f
C12873 DVSS.t176 VSS 0.272754f
C12874 DVSS.n1611 VSS 0.021956f
C12875 DVSS.t136 VSS 0.003611f
C12876 DVSS.t177 VSS 0.003611f
C12877 DVSS.n1612 VSS 0.007291f
C12878 DVSS.n1613 VSS 8.12e-19
C12879 DVSS.n1614 VSS 0.021061f
C12880 DVSS.t134 VSS 0.009309f
C12881 DVSS.n1615 VSS 0.003795f
C12882 DVSS.n1616 VSS 0.021061f
C12883 DVSS.n1617 VSS 0.018248f
C12884 DVSS.t111 VSS 0.009309f
C12885 DVSS.n1618 VSS 0.003795f
C12886 DVSS.n1619 VSS 0.021061f
C12887 DVSS.t145 VSS 0.003611f
C12888 DVSS.t109 VSS 0.003611f
C12889 DVSS.n1620 VSS 0.007291f
C12890 DVSS.n1621 VSS 8.12e-19
C12891 DVSS.n1622 VSS 0.021061f
C12892 DVSS.n1623 VSS 0.432321f
C12893 DVSS.t110 VSS 0.409505f
C12894 DVSS.t108 VSS 0.274249f
C12895 DVSS.n1624 VSS 0.158916f
C12896 DVSS.n1625 VSS 0.016916f
C12897 DVSS.t143 VSS 0.009309f
C12898 DVSS.n1626 VSS 0.003795f
C12899 DVSS.n1627 VSS 0.058661f
C12900 DVSS.n1628 VSS 0.092043f
C12901 DVSS.n1629 VSS 0.092043f
C12902 DVSS.n1630 VSS 0.092043f
C12903 DVSS.n1631 VSS 1.13868f
C12904 DVSS.n1632 VSS 0.04829f
C12905 DVSS.n1633 VSS 0.291792f
C12906 DVSS.n1634 VSS 1.97868f
C12907 DVSS.n1635 VSS 1.29089f
C12908 DVSS.n1636 VSS 0.092043f
C12909 DVSS.n1637 VSS 0.092043f
C12910 DVSS.n1638 VSS 0.092043f
C12911 DVSS.n1639 VSS 0.092043f
C12912 DVSS.n1640 VSS 0.092043f
C12913 DVSS.n1641 VSS 0.092043f
C12914 DVSS.n1642 VSS 0.06048f
C12915 DVSS.n1643 VSS 0.092043f
C12916 DVSS.n1644 VSS 0.092043f
C12917 DVSS.n1645 VSS 0.092043f
C12918 DVSS.n1646 VSS 0.059309f
C12919 DVSS.n1647 VSS 0.06048f
C12920 DVSS.n1648 VSS 0.092043f
C12921 DVSS.n1649 VSS 0.092043f
C12922 DVSS.n1650 VSS 0.092043f
C12923 DVSS.n1651 VSS 0.085237f
C12924 DVSS.n1652 VSS 0.062562f
C12925 DVSS.n1653 VSS 0.092043f
C12926 DVSS.n1654 VSS 0.092043f
C12927 DVSS.n1655 VSS 0.092043f
C12928 DVSS.n1656 VSS 0.050235f
C12929 DVSS.n1657 VSS 0.046022f
C12930 DVSS.n1658 VSS 0.092043f
C12931 DVSS.n1659 VSS 0.092043f
C12932 DVSS.n1660 VSS 0.092043f
C12933 DVSS.n1661 VSS 0.046022f
C12934 DVSS.n1662 VSS 0.046022f
C12935 DVSS.n1663 VSS 0.026298f
C12936 DVSS.n1664 VSS 0.026298f
C12937 DVSS.n1665 VSS 0.026298f
C12938 DVSS.n1666 VSS 0.026298f
C12939 DVSS.n1668 VSS 0.026298f
C12940 DVSS.n1670 VSS 0.092043f
C12941 DVSS.n1671 VSS 0.092043f
C12942 DVSS.n1672 VSS 0.092043f
C12943 DVSS.n1673 VSS 0.092043f
C12944 DVSS.n1674 VSS 0.092043f
C12945 DVSS.n1675 VSS 0.092043f
C12946 DVSS.n1676 VSS 0.092043f
C12947 DVSS.n1677 VSS 0.092043f
C12948 DVSS.n1678 VSS 0.092043f
C12949 DVSS.n1679 VSS 0.092043f
C12950 DVSS.n1680 VSS 0.092043f
C12951 DVSS.n1681 VSS 0.092043f
C12952 DVSS.n1682 VSS 0.051531f
C12953 DVSS.n1683 VSS 0.162256f
C12954 DVSS.n1684 VSS -0.005479f
C12955 DVSS.t194 VSS 0.009309f
C12956 DVSS.n1685 VSS 0.003795f
C12957 DVSS.n1686 VSS 0.042888f
C12958 DVSS.n1687 VSS 0.05542f
C12959 DVSS.n1688 VSS 0.092043f
C12960 DVSS.n1689 VSS 0.092043f
C12961 DVSS.n1690 VSS 0.092043f
C12962 DVSS.n1691 VSS 0.092043f
C12963 DVSS.n1692 VSS 0.092043f
C12964 DVSS.n1693 VSS 0.092043f
C12965 DVSS.n1694 VSS 0.06255f
C12966 DVSS.n1695 VSS 0.047774f
C12967 DVSS.n1696 VSS 0.10121f
C12968 DVSS.t91 VSS 0.056793f
C12969 DVSS.t191 VSS 0.216709f
C12970 DVSS.n1697 VSS 0.021956f
C12971 DVSS.t94 VSS 0.003611f
C12972 DVSS.t192 VSS 0.003611f
C12973 DVSS.n1698 VSS 0.007291f
C12974 DVSS.n1699 VSS 8.12e-19
C12975 DVSS.n1700 VSS 0.021061f
C12976 DVSS.t92 VSS 0.009309f
C12977 DVSS.n1701 VSS 0.003795f
C12978 DVSS.n1702 VSS 0.021061f
C12979 DVSS.t10 VSS 0.228665f
C12980 DVSS.t193 VSS 0.182334f
C12981 DVSS.t7 VSS 0.182334f
C12982 DVSS.t99 VSS 0.158422f
C12983 DVSS.n1703 VSS 0.090914f
C12984 DVSS.t13 VSS 0.091914f
C12985 DVSS.t140 VSS 0.250336f
C12986 DVSS.t148 VSS 0.22194f
C12987 DVSS.t15 VSS 0.22194f
C12988 DVSS.t4 VSS 0.187565f
C12989 DVSS.t2 VSS 0.227171f
C12990 DVSS.n1704 VSS 0.160314f
C12991 DVSS.n1705 VSS 0.018248f
C12992 DVSS.t149 VSS 0.009309f
C12993 DVSS.n1706 VSS 0.003795f
C12994 DVSS.n1707 VSS 0.049587f
C12995 DVSS.n1708 VSS 0.063581f
C12996 DVSS.n1709 VSS 0.092043f
C12997 DVSS.n1710 VSS 0.092043f
C12998 DVSS.n1711 VSS 0.092043f
C12999 DVSS.n1712 VSS 0.092043f
C13000 DVSS.n1713 VSS 0.092043f
C13001 DVSS.n1714 VSS 0.092043f
C13002 DVSS.n1715 VSS 0.092043f
C13003 DVSS.n1716 VSS 0.092043f
C13004 DVSS.n1717 VSS 0.092043f
C13005 DVSS.n1718 VSS 0.092043f
C13006 DVSS.n1719 VSS 0.092043f
C13007 DVSS.n1720 VSS 0.058985f
C13008 DVSS.n1721 VSS 0.06048f
C13009 DVSS.n1722 VSS 0.049587f
C13010 DVSS.n1723 VSS 0.092043f
C13011 DVSS.n1724 VSS 0.092043f
C13012 DVSS.n1725 VSS 0.092043f
C13013 DVSS.n1726 VSS 0.06048f
C13014 DVSS.t88 VSS 0.009309f
C13015 DVSS.n1727 VSS 0.003795f
C13016 DVSS.n1728 VSS 0.01033f
C13017 DVSS.n1729 VSS 0.045313f
C13018 DVSS.n1730 VSS 0.047349f
C13019 DVSS.n1731 VSS 0.092043f
C13020 DVSS.n1732 VSS 0.092043f
C13021 DVSS.n1733 VSS 0.092043f
C13022 DVSS.n1734 VSS 0.06093f
C13023 DVSS.n1735 VSS 0.062562f
C13024 DVSS.n1736 VSS 0.092043f
C13025 DVSS.n1737 VSS 0.092043f
C13026 DVSS.n1738 VSS 0.092043f
C13027 DVSS.n1739 VSS 0.092043f
C13028 DVSS.n1740 VSS 0.092043f
C13029 DVSS.n1741 VSS 0.092043f
C13030 DVSS.n1742 VSS 0.092043f
C13031 DVSS.n1743 VSS 0.092043f
C13032 DVSS.n1744 VSS 0.092043f
C13033 DVSS.n1745 VSS 0.092043f
C13034 DVSS.n1746 VSS 0.092043f
C13035 DVSS.n1747 VSS 0.092043f
C13036 DVSS.n1748 VSS 0.092043f
C13037 DVSS.n1749 VSS 0.092043f
C13038 DVSS.n1750 VSS 0.092043f
C13039 DVSS.n1751 VSS 0.092043f
C13040 DVSS.n1752 VSS 0.092043f
C13041 DVSS.n1753 VSS 0.092043f
C13042 DVSS.n1754 VSS 0.092043f
C13043 DVSS.n1755 VSS 0.092043f
C13044 DVSS.n1756 VSS 0.092043f
C13045 DVSS.n1757 VSS 0.092043f
C13046 DVSS.n1758 VSS 0.092043f
C13047 DVSS.n1759 VSS 0.092043f
C13048 DVSS.n1760 VSS 0.082968f
C13049 DVSS.n1761 VSS 0.082968f
C13050 DVSS.n1762 VSS 0.443616f
C13051 DVSS.n1763 VSS 0.121157f
C13052 DVSS.n1764 VSS 0.047318f
C13053 DVSS.n1765 VSS 0.092043f
C13054 DVSS.n1766 VSS 0.092043f
C13055 DVSS.n1767 VSS 0.092043f
C13056 DVSS.n1768 VSS 0.092043f
C13057 DVSS.n1769 VSS 0.092043f
C13058 DVSS.n1770 VSS 0.092043f
C13059 DVSS.n1771 VSS 0.092043f
C13060 DVSS.n1772 VSS 0.092043f
C13061 DVSS.n1773 VSS 0.092043f
C13062 DVSS.n1774 VSS 0.092043f
C13063 DVSS.n1775 VSS 0.092043f
C13064 DVSS.n1776 VSS 0.092043f
C13065 DVSS.n1777 VSS 0.091719f
C13066 DVSS.n1778 VSS 0.042307f
C13067 DVSS.n1779 VSS 0.084022f
C13068 DVSS.n1780 VSS 0.084022f
C13069 DVSS.n1781 VSS 0.084022f
C13070 DVSS.n1782 VSS 0.084022f
C13071 DVSS.n1783 VSS 0.052366f
C13072 DVSS.n1784 VSS 0.084022f
C13073 DVSS.n1785 VSS 0.084022f
C13074 DVSS.n1786 VSS 0.084022f
C13075 DVSS.n1787 VSS 0.042011f
C13076 DVSS.n1788 VSS 0.019808f
C13077 DVSS.n1789 VSS 0.010334f
C13078 DVSS.n1790 VSS 0.023309f
C13079 DVSS.n1791 VSS 0.051455f
C13080 DVSS.n1792 VSS 0.277464f
C13081 DVSS.n1793 VSS 0.277464f
C13082 DVSS.n1794 VSS 1.9283f
C13083 DVSS.t104 VSS 0.323604f
C13084 DVSS.n1795 VSS 0.098622f
C13085 DVSS.n1796 VSS 0.044396f
C13086 DVSS.n1797 VSS 0.044396f
C13087 DVSS.n1798 VSS 0.044396f
C13088 DVSS.n1799 VSS 0.044396f
C13089 DVSS.n1800 VSS 0.044396f
C13090 DVSS.n1801 VSS 0.044396f
C13091 DVSS.n1804 VSS 0.044396f
C13092 DVSS.n1806 VSS 0.044396f
C13093 DVSS.n1808 VSS 0.044396f
C13094 DVSS.n1810 VSS 0.044396f
C13095 DVSS.n1812 VSS 0.044396f
C13096 DVSS.n1813 VSS 0.1146f
C13097 DVSS.n1814 VSS 0.1146f
C13098 DVSS.n1815 VSS 0.1146f
C13099 DVSS.n1822 VSS 1.72114f
C13100 DVSS.n1824 VSS 0.1146f
C13101 DVSS.n1826 VSS 0.1146f
C13102 DVSS.t151 VSS 0.007612f
C13103 DVSS.n1827 VSS 0.006851f
C13104 DVSS.t105 VSS 0.007612f
C13105 DVSS.n1828 VSS 0.006851f
C13106 DVSS.t77 VSS 0.003611f
C13107 DVSS.n1829 VSS 0.00868f
C13108 DVSS.n1830 VSS 0.007358f
C13109 DVSS.t86 VSS 0.00812f
C13110 DVSS.t90 VSS 0.007704f
C13111 DVSS.t182 VSS 0.007704f
C13112 DVSS.n1831 VSS 0.016246f
C13113 DVSS.n1832 VSS 0.009892f
C13114 DVSS.t184 VSS 0.007704f
C13115 DVSS.t96 VSS 0.007704f
C13116 DVSS.n1833 VSS 0.016246f
C13117 DVSS.n1834 VSS 0.007586f
C13118 DVSS.n1835 VSS 0.0832f
C13119 DVSS.n1836 VSS 0.01908f
C13120 DVSS.n1837 VSS 0.011857f
C13121 DVSS.n1838 VSS 0.025736f
C13122 DVSS.n1839 VSS 0.018738f
C13123 DVSS.n1840 VSS 0.019893f
C13124 DVSS.n1841 VSS 0.013911f
C13125 DVSS.n1842 VSS 0.064155f
C13126 DVSS.n1843 VSS 0.044795f
C13127 DVSS.n1845 VSS 0.122954f
C13128 DVSS.n1846 VSS 0.034039f
C13129 DVSS.t138 VSS 0.003611f
C13130 DVSS.n1847 VSS 0.008681f
C13131 DVSS.n1848 VSS 0.006598f
C13132 DVSS.n1849 VSS 3.80907f
C13133 DVSS.n1850 VSS 0.06968f
C13134 DVSS.n1851 VSS 0.092043f
C13135 DVSS.n1852 VSS 0.092043f
C13136 DVSS.n1853 VSS 0.092043f
C13137 DVSS.n1854 VSS 0.068384f
C13138 DVSS.n1855 VSS 0.046022f
C13139 DVSS.n1856 VSS 0.092043f
C13140 DVSS.n1857 VSS 0.092043f
C13141 DVSS.n1858 VSS 0.092043f
C13142 DVSS.n1859 VSS 0.045373f
C13143 DVSS.n1860 VSS 0.046022f
C13144 DVSS.n1861 VSS 0.004491f
C13145 DVSS.n1862 VSS 0.004491f
C13146 DVSS.n1863 VSS 0.009456f
C13147 DVSS.n1864 VSS 0.006575f
C13148 DVSS.n1865 VSS 0.006575f
C13149 DVSS.n1866 VSS 0.011101f
C13150 DVSS.n1867 VSS 0.014694f
C13151 DVSS.n1868 VSS 0.006308f
C13152 DVSS.n1869 VSS 0.007331f
C13153 DVSS.n1870 VSS 0.00555f
C13154 DVSS.n1871 VSS 0.011101f
C13155 DVSS.n1872 VSS 0.00555f
C13156 DVSS.n1873 VSS 0.025928f
C13157 DVSS.n1874 VSS 0.025928f
C13158 DVSS.n1875 VSS 0.035827f
C13159 DVSS.n1876 VSS 0.025928f
C13160 DVSS.n1877 VSS 0.020742f
C13161 DVSS.n1878 VSS 0.046022f
C13162 DVSS.n1879 VSS 0.092043f
C13163 DVSS.n1880 VSS 0.092043f
C13164 DVSS.n1881 VSS 0.092043f
C13165 DVSS.n1882 VSS 0.092043f
C13166 DVSS.n1883 VSS 0.092043f
C13167 DVSS.n1884 VSS 0.046022f
C13168 DVSS.n1885 VSS 0.046022f
C13169 DVSS.n1886 VSS 0.046022f
C13170 DVSS.n1887 VSS 0.007166f
C13171 DVSS.n1888 VSS 0.00545f
C13172 DVSS.n1889 VSS 0.011101f
C13173 DVSS.n1890 VSS 0.011101f
C13174 DVSS.n1891 VSS 0.011101f
C13175 DVSS.n1892 VSS 0.00545f
C13176 DVSS.n1893 VSS 0.005703f
C13177 DVSS.n1894 VSS 0.00545f
C13178 DVSS.n1895 VSS 0.006914f
C13179 DVSS.n1896 VSS 0.011101f
C13180 DVSS.n1897 VSS 0.011101f
C13181 DVSS.n1898 VSS 0.011101f
C13182 DVSS.n1899 VSS 0.003945f
C13183 DVSS.n1901 VSS 0.019426f
C13184 DVSS.n1902 VSS 0.036299f
C13185 DVSS.n1903 VSS 0.019279f
C13186 DVSS.n1904 VSS 0.010371f
C13187 DVSS.n1905 VSS 0.092043f
C13188 DVSS.n1906 VSS 0.092043f
C13189 DVSS.n1907 VSS 0.092043f
C13190 DVSS.n1908 VSS 0.092043f
C13191 DVSS.n1909 VSS 0.092043f
C13192 DVSS.n1910 VSS 0.092043f
C13193 DVSS.n1911 VSS 0.012334f
C13194 DVSS.n1912 VSS 0.045373f
C13195 DVSS.n1913 VSS 0.035975f
C13196 DVSS.n1914 VSS 0.010695f
C13197 DVSS.n1916 VSS 0.003129f
C13198 DVSS.n1917 VSS 0.011101f
C13199 DVSS.n1918 VSS 0.171951f
C13200 DVSS.t14 VSS 2.19675f
C13201 DVSS.n1919 VSS 0.248361f
C13202 DVSS.n1920 VSS 0.00555f
C13203 DVSS.n1921 VSS 0.17198f
C13204 DVSS.n1922 VSS 0.027748f
C13205 DVSS.n1923 VSS 0.007298f
C13206 DVSS.n1924 VSS 0.045373f
C13207 DVSS.n1925 VSS 0.045373f
C13208 DVSS.n1926 VSS 0.110631f
C13209 DVSS.n1927 VSS 0.030664f
C13210 DVSS.n1928 VSS 0.07864f
C13211 DVSS.n1929 VSS 0.248361f
C13212 DVSS.n1930 VSS 0.090023f
C13213 DVSS.n1931 VSS 0.027748f
C13214 DVSS.n1932 VSS 0.00545f
C13215 DVSS.n1933 VSS 0.00555f
C13216 DVSS.n1934 VSS 0.00545f
C13217 DVSS.n1935 VSS 0.008171f
C13218 DVSS.n1936 VSS 0.016723f
C13219 DVSS.n1937 VSS 0.005834f
C13220 DVSS.n1938 VSS 0.040836f
C13221 DVSS.n1939 VSS 0.008409f
C13222 DVSS.n1940 VSS 0.008075f
C13223 DVSS.n1941 VSS 0.008125f
C13224 DVSS.n1942 VSS 0.005753f
C13225 DVSS.n1943 VSS 0.011101f
C13226 DVSS.n1944 VSS 0.006321f
C13227 DVSS.n1945 VSS 0.007166f
C13228 DVSS.n1946 VSS 0.00545f
C13229 DVSS.n1947 VSS 0.007166f
C13230 DVSS.n1948 VSS 0.01033f
C13231 DVSS.n1949 VSS 0.009405f
C13232 DVSS.n1950 VSS 0.007166f
C13233 DVSS.n1951 VSS 0.02002f
C13234 DVSS.n1952 VSS 0.018926f
C13235 DVSS.n1954 VSS 0.024884f
C13236 DVSS.n1955 VSS 0.018926f
C13237 DVSS.n1957 VSS 0.046022f
C13238 DVSS.n1958 VSS 0.024359f
C13239 DVSS.n1959 VSS 0.046022f
C13240 DVSS.n1960 VSS 0.051531f
C13241 DVSS.n1961 VSS 0.018926f
C13242 DVSS.n1962 VSS 0.018926f
C13243 DVSS.n1963 VSS 0.018926f
C13244 DVSS.n1964 VSS 0.092043f
C13245 DVSS.n1965 VSS 0.046022f
C13246 DVSS.n1966 VSS 0.092043f
C13247 DVSS.n1967 VSS 0.092043f
C13248 DVSS.n1968 VSS 0.092043f
C13249 DVSS.n1969 VSS 0.046022f
C13250 DVSS.n1970 VSS 0.312003f
C13251 DVSS.n1971 VSS 0.041808f
C13252 DVSS.n1972 VSS 0.071513f
C13253 DVSS.n1973 VSS 0.009596f
C13254 DVSS.t12 VSS 0.014445f
C13255 DVSS.n1974 VSS 0.038498f
C13256 DVSS.n1975 VSS 0.002551f
C13257 DVSS.n1976 VSS 0.024934f
C13258 DVSS.n1977 VSS 5.33422f
C13259 DVSS.n1978 VSS 0.197235f
C13260 DVSS.n1979 VSS 3.99643f
C13261 DVSS.n1980 VSS 0.197235f
C13262 DVSS.n1981 VSS 0.197235f
C13263 DVSS.n1982 VSS 0.181262f
C13264 DVSS.n1983 VSS 0.197235f
C13265 DVSS.n1984 VSS 0.197235f
C13266 DVSS.n1985 VSS 0.197235f
C13267 DVSS.n1986 VSS 0.197235f
C13268 DVSS.n1987 VSS 0.197235f
C13269 DVSS.n1988 VSS 0.129078f
C13270 DVSS.n1989 VSS 0.197235f
C13271 DVSS.n1990 VSS 0.197235f
C13272 DVSS.n1991 VSS 0.197235f
C13273 DVSS.n1992 VSS 0.197235f
C13274 DVSS.n1993 VSS 0.197235f
C13275 DVSS.n1994 VSS 0.197235f
C13276 DVSS.n1995 VSS 0.197235f
C13277 DVSS.n1996 VSS 0.197235f
C13278 DVSS.n1997 VSS 0.197235f
C13279 DVSS.n1998 VSS 0.197235f
C13280 DVSS.n1999 VSS 0.197235f
C13281 DVSS.n2000 VSS 0.197235f
C13282 DVSS.n2001 VSS 0.197235f
C13283 DVSS.n2002 VSS 0.197235f
C13284 DVSS.n2003 VSS 0.114591f
C13285 DVSS.n2004 VSS 0.197235f
C13286 DVSS.n2005 VSS 0.197235f
C13287 DVSS.n2006 VSS 0.197235f
C13288 DVSS.n2007 VSS 0.197235f
C13289 DVSS.n2008 VSS 0.197235f
C13290 DVSS.n2009 VSS 0.197235f
C13291 DVSS.n2010 VSS 0.197235f
C13292 DVSS.n2011 VSS 0.197235f
C13293 DVSS.n2012 VSS 0.699965f
C13294 DVSS.n2013 VSS 0.146537f
C13295 DVSS.n2014 VSS 3.52082f
C13296 DVSS.n2015 VSS 0.590127f
C13297 DVSS.n2016 VSS 0.362971f
C13298 DVSS.n2017 VSS 1.86223f
C13299 DVSS.n2018 VSS 3.62392f
C13300 DVSS.n2019 VSS 2.18756f
C13301 DVSS.n2020 VSS 0.092043f
C13302 DVSS.n2021 VSS 0.063847f
C13303 DVSS.n2022 VSS 0.092043f
C13304 DVSS.n2023 VSS 0.092043f
C13305 DVSS.n2024 VSS 0.092043f
C13306 DVSS.n2025 VSS 0.092043f
C13307 DVSS.n2026 VSS 0.092043f
C13308 DVSS.n2027 VSS 0.092043f
C13309 DVSS.n2028 VSS 0.092043f
C13310 DVSS.n2029 VSS 0.092043f
C13311 DVSS.n2030 VSS 0.092043f
C13312 DVSS.n2031 VSS 0.092043f
C13313 DVSS.n2032 VSS 0.092043f
C13314 DVSS.n2033 VSS 0.092043f
C13315 DVSS.n2034 VSS 0.092043f
C13316 DVSS.n2035 VSS 0.092043f
C13317 DVSS.n2036 VSS 0.092043f
C13318 DVSS.n2037 VSS 0.092043f
C13319 DVSS.n2038 VSS 0.092043f
C13320 DVSS.n2039 VSS 0.092043f
C13321 DVSS.n2040 VSS 0.092043f
C13322 DVSS.n2041 VSS 0.092043f
C13323 DVSS.n2042 VSS 0.092043f
C13324 DVSS.n2043 VSS 0.092043f
C13325 DVSS.n2044 VSS 0.092043f
C13326 DVSS.n2045 VSS 0.092043f
C13327 DVSS.n2046 VSS 0.092043f
C13328 DVSS.n2047 VSS 0.092043f
C13329 DVSS.n2048 VSS 0.092043f
C13330 DVSS.n2049 VSS 0.092043f
C13331 DVSS.n2050 VSS 0.092043f
C13332 DVSS.n2051 VSS 0.092043f
C13333 DVSS.n2052 VSS 0.092043f
C13334 DVSS.n2053 VSS 0.092043f
C13335 DVSS.n2054 VSS 0.092043f
C13336 DVSS.n2055 VSS 0.092043f
C13337 DVSS.n2056 VSS 0.092043f
C13338 DVSS.n2057 VSS 0.092043f
C13339 DVSS.n2058 VSS 0.092043f
C13340 DVSS.n2059 VSS 0.092043f
C13341 DVSS.n2060 VSS 0.092043f
C13342 DVSS.n2061 VSS 0.08783f
C13343 DVSS.n2062 VSS 0.092043f
C13344 DVSS.n2063 VSS 0.092043f
C13345 DVSS.n2064 VSS 0.092043f
C13346 DVSS.n2065 VSS 0.092043f
C13347 DVSS.n2066 VSS 0.092043f
C13348 DVSS.n2067 VSS 0.092043f
C13349 DVSS.n2068 VSS 0.092043f
C13350 DVSS.n2069 VSS 0.092043f
C13351 DVSS.n2070 VSS 0.092043f
C13352 DVSS.n2071 VSS 0.092043f
C13353 DVSS.n2072 VSS 0.092043f
C13354 DVSS.n2073 VSS 0.092043f
C13355 DVSS.n2074 VSS 0.092043f
C13356 DVSS.n2075 VSS 0.092043f
C13357 DVSS.n2076 VSS 0.092043f
C13358 DVSS.n2077 VSS 0.092043f
C13359 DVSS.n2078 VSS 0.092043f
C13360 DVSS.n2079 VSS 0.092043f
C13361 DVSS.n2080 VSS 0.092043f
C13362 DVSS.n2081 VSS 0.092043f
C13363 DVSS.n2082 VSS 0.092043f
C13364 DVSS.n2083 VSS 0.092043f
C13365 DVSS.n2084 VSS 0.092043f
C13366 DVSS.n2085 VSS 0.092043f
C13367 DVSS.n2086 VSS 0.092043f
C13368 DVSS.n2087 VSS 0.092043f
C13369 DVSS.n2088 VSS 0.092043f
C13370 DVSS.n2089 VSS 0.092043f
C13371 DVSS.n2090 VSS 0.047318f
C13372 DVSS.n2091 VSS 0.121165f
C13373 DVSS.n2092 VSS 0.443501f
C13374 DVSS.n2093 VSS 0.082968f
C13375 DVSS.n2094 VSS 0.082968f
C13376 DVSS.n2095 VSS 0.092043f
C13377 DVSS.n2096 VSS 0.092043f
C13378 DVSS.n2097 VSS 0.092043f
C13379 DVSS.n2098 VSS 0.092043f
C13380 DVSS.n2099 VSS 0.092043f
C13381 DVSS.n2100 VSS 0.092043f
C13382 DVSS.n2101 VSS 0.092043f
C13383 DVSS.n2102 VSS 0.092043f
C13384 DVSS.n2103 VSS 0.092043f
C13385 DVSS.n2104 VSS 0.092043f
C13386 DVSS.n2105 VSS 0.092043f
C13387 DVSS.n2106 VSS 0.092043f
C13388 DVSS.n2107 VSS 0.092043f
C13389 DVSS.n2108 VSS 0.092043f
C13390 DVSS.n2109 VSS 0.092043f
C13391 DVSS.n2110 VSS 0.092043f
C13392 DVSS.n2111 VSS 0.092043f
C13393 DVSS.n2112 VSS 0.092043f
C13394 DVSS.n2113 VSS 0.092043f
C13395 DVSS.n2114 VSS 0.092043f
C13396 DVSS.n2115 VSS 0.092043f
C13397 DVSS.n2116 VSS 0.092043f
C13398 DVSS.n2117 VSS 0.092043f
C13399 DVSS.n2118 VSS 0.092043f
C13400 DVSS.n2119 VSS 0.092043f
C13401 DVSS.n2120 VSS 0.092043f
C13402 DVSS.n2121 VSS 0.092043f
C13403 DVSS.n2122 VSS 0.092043f
C13404 DVSS.n2123 VSS 0.092043f
C13405 DVSS.n2124 VSS 0.092043f
C13406 DVSS.n2125 VSS 0.092043f
C13407 DVSS.n2126 VSS 0.092043f
C13408 DVSS.n2127 VSS 0.092043f
C13409 DVSS.n2128 VSS 0.092043f
C13410 DVSS.n2129 VSS 0.092043f
C13411 DVSS.n2130 VSS 0.092043f
C13412 DVSS.n2131 VSS 0.092043f
C13413 DVSS.n2132 VSS 0.092043f
C13414 DVSS.n2133 VSS 0.092043f
C13415 DVSS.n2134 VSS 0.092043f
C13416 DVSS.n2135 VSS 0.092043f
C13417 DVSS.n2136 VSS 0.092043f
C13418 DVSS.n2137 VSS 0.092043f
C13419 DVSS.n2138 VSS 0.092043f
C13420 DVSS.n2139 VSS 0.092043f
C13421 DVSS.n2140 VSS 0.092043f
C13422 DVSS.n2141 VSS 0.092043f
C13423 DVSS.n2142 VSS 0.092043f
C13424 DVSS.n2143 VSS 0.092043f
C13425 DVSS.n2144 VSS 0.092043f
C13426 DVSS.n2145 VSS 0.092043f
C13427 DVSS.n2146 VSS 0.092043f
C13428 DVSS.n2147 VSS 0.092043f
C13429 DVSS.n2148 VSS 0.046022f
C13430 DVSS.n2149 VSS 0.092043f
C13431 DVSS.n2150 VSS 0.092043f
C13432 DVSS.n2151 VSS 0.092043f
C13433 DVSS.n2152 VSS 0.092043f
C13434 DVSS.n2153 VSS 0.092043f
C13435 DVSS.n2154 VSS 0.092043f
C13436 DVSS.n2155 VSS 0.092043f
C13437 DVSS.n2156 VSS 0.092043f
C13438 DVSS.n2157 VSS 0.092043f
C13439 DVSS.n2158 VSS 0.092043f
C13440 DVSS.n2159 VSS 0.092043f
C13441 DVSS.n2160 VSS 0.092043f
C13442 DVSS.n2161 VSS 0.092043f
C13443 DVSS.n2162 VSS 0.092043f
C13444 DVSS.n2163 VSS 0.092043f
C13445 DVSS.n2164 VSS 0.092043f
C13446 DVSS.n2165 VSS 0.092043f
C13447 DVSS.n2166 VSS 0.092043f
C13448 DVSS.n2167 VSS 0.092043f
C13449 DVSS.n2168 VSS 0.092043f
C13450 DVSS.n2169 VSS 0.092043f
C13451 DVSS.n2170 VSS 0.092043f
C13452 DVSS.n2171 VSS 0.092043f
C13453 DVSS.n2172 VSS 0.092043f
C13454 DVSS.n2173 VSS 0.092043f
C13455 DVSS.n2174 VSS 0.092043f
C13456 DVSS.n2175 VSS 0.092043f
C13457 DVSS.n2176 VSS 0.092043f
C13458 DVSS.n2177 VSS 0.092043f
C13459 DVSS.n2178 VSS 0.092043f
C13460 DVSS.n2179 VSS 0.092043f
C13461 DVSS.n2180 VSS 0.092043f
C13462 DVSS.n2181 VSS 0.092043f
C13463 DVSS.n2182 VSS 0.092043f
C13464 DVSS.n2183 VSS 0.092043f
C13465 DVSS.n2184 VSS 0.092043f
C13466 DVSS.n2185 VSS 0.092043f
C13467 DVSS.n2186 VSS 0.092043f
C13468 DVSS.n2187 VSS 0.092043f
C13469 DVSS.n2188 VSS 0.092043f
C13470 DVSS.n2189 VSS 0.092043f
C13471 DVSS.n2190 VSS 0.092043f
C13472 DVSS.n2191 VSS 0.092043f
C13473 DVSS.n2192 VSS 0.092043f
C13474 DVSS.n2193 VSS 0.092043f
C13475 DVSS.n2194 VSS 0.092043f
C13476 DVSS.n2195 VSS 0.092043f
C13477 DVSS.n2196 VSS 0.092043f
C13478 DVSS.n2197 VSS 0.092043f
C13479 DVSS.n2198 VSS 0.092043f
C13480 DVSS.n2199 VSS 0.092043f
C13481 DVSS.n2200 VSS 0.092043f
C13482 DVSS.n2201 VSS 0.092043f
C13483 DVSS.n2202 VSS 0.092043f
C13484 DVSS.n2203 VSS 0.092043f
C13485 DVSS.n2204 VSS 0.092043f
C13486 DVSS.n2205 VSS 0.092043f
C13487 DVSS.n2206 VSS 0.092043f
C13488 DVSS.n2207 VSS 0.092043f
C13489 DVSS.n2208 VSS 0.092043f
C13490 DVSS.n2209 VSS 0.092043f
C13491 DVSS.n2210 VSS 0.092043f
C13492 DVSS.n2211 VSS 0.092043f
C13493 DVSS.n2212 VSS 0.092043f
C13494 DVSS.n2213 VSS 0.092043f
C13495 DVSS.n2214 VSS 0.092043f
C13496 DVSS.n2215 VSS 0.092043f
C13497 DVSS.n2216 VSS 0.092043f
C13498 DVSS.n2217 VSS 0.092043f
C13499 DVSS.n2218 VSS 0.092043f
C13500 DVSS.n2219 VSS 0.092043f
C13501 DVSS.n2220 VSS 0.086534f
C13502 DVSS.n2221 VSS 0.092043f
C13503 DVSS.n2222 VSS 0.092043f
C13504 DVSS.n2223 VSS 0.092043f
C13505 DVSS.n2224 VSS 0.092043f
C13506 DVSS.n2225 VSS 0.092043f
C13507 DVSS.n2226 VSS 0.046022f
C13508 DVSS.n2227 VSS 0.018926f
C13509 DVSS.n2228 VSS 0.018926f
C13510 DVSS.n2229 VSS 0.018926f
C13511 DVSS.n2230 VSS 0.024884f
C13512 DVSS.n2231 VSS 0.010819f
C13513 DVSS.n2232 VSS 0.019452f
C13514 DVSS.n2233 VSS 0.018401f
C13515 DVSS.n2234 VSS 0.024884f
C13516 DVSS.n2235 VSS 0.018401f
C13517 DVSS.n2236 VSS 0.024884f
C13518 DVSS.n2237 VSS 0.018401f
C13519 DVSS.n2238 VSS 0.024884f
C13520 DVSS.n2239 VSS 0.018401f
C13521 DVSS.n2240 VSS 0.018401f
C13522 DVSS.n2241 VSS 0.019452f
C13523 DVSS.n2242 VSS 0.024359f
C13524 DVSS.n2243 VSS 0.018401f
C13525 DVSS.n2244 VSS 0.024884f
C13526 DVSS.n2245 VSS 0.018401f
C13527 DVSS.n2246 VSS 0.018401f
C13528 DVSS.n2247 VSS 0.024123f
C13529 DVSS.n2248 VSS 0.038714f
C13530 DVSS.n2249 VSS 0.046022f
C13531 DVSS.n2250 VSS 0.018926f
C13532 DVSS.n2251 VSS 0.024884f
C13533 DVSS.n2252 VSS 0.02215f
C13534 DVSS.n2253 VSS 0.113302f
C13535 DVSS.n2254 VSS 0.421982f
C13536 DVSS.n2255 VSS 0.054924f
C13537 DVSS.n2256 VSS 0.007889f
C13538 DVSS.n2257 VSS 0.036299f
C13539 DVSS.n2258 VSS 0.092043f
C13540 DVSS.n2259 VSS 0.092043f
C13541 DVSS.n2260 VSS 0.010371f
C13542 DVSS.n2261 VSS 0.045373f
C13543 DVSS.n2262 VSS 0.007889f
C13544 DVSS.n2263 VSS 0.015779f
C13545 DVSS.n2264 VSS 0.045373f
C13546 DVSS.n2265 VSS 0.016501f
C13547 DVSS.n2266 VSS 0.102854f
C13548 DVSS.n2267 VSS 0.110631f
C13549 DVSS.n2269 VSS 0.045373f
C13550 DVSS.n2270 VSS 0.029322f
C13551 DVSS.n2271 VSS 0.020742f
C13552 DVSS.n2272 VSS 0.092043f
C13553 DVSS.n2273 VSS 0.092043f
C13554 DVSS.n2274 VSS 0.092043f
C13555 DVSS.n2275 VSS 0.046022f
C13556 DVSS.n2276 VSS 0.008612f
C13557 DVSS.n2277 VSS 0.288091f
C13558 DVSS.n2278 VSS 0.046022f
C13559 DVSS.n2279 VSS 0.046022f
C13560 DVSS.n2280 VSS 0.046022f
C13561 DVSS.n2281 VSS 0.092043f
C13562 DVSS.n2282 VSS 0.092043f
C13563 DVSS.n2283 VSS 0.092043f
C13564 DVSS.n2284 VSS 0.092043f
C13565 DVSS.n2285 VSS 0.046022f
C13566 DVSS.n2286 VSS 0.046022f
C13567 DVSS.n2287 VSS 0.382838f
C13568 DVSS.n2288 VSS 0.046022f
C13569 DVSS.n2289 VSS 0.046022f
C13570 DVSS.n2290 VSS 0.092043f
C13571 DVSS.n2291 VSS 0.092043f
C13572 DVSS.n2292 VSS 0.092043f
C13573 DVSS.n2293 VSS 0.092043f
C13574 DVSS.n2294 VSS 0.092043f
C13575 DVSS.n2295 VSS 0.020742f
C13576 DVSS.n2296 VSS 0.045373f
C13577 DVSS.n2299 VSS 0.029322f
C13578 DVSS.n2300 VSS 0.045373f
C13579 DVSS.n2301 VSS 0.030664f
C13580 DVSS.n2302 VSS 0.144261f
C13581 DVSS.n2303 VSS 0.189694f
C13582 DVSS.n2304 VSS 0.167296f
C13583 DVSS.n2305 VSS 0.088697f
C13584 DVSS.n2306 VSS 0.100594f
C13585 DVSS.n2307 VSS 0.014483f
C13586 DVSS.n2308 VSS 0.199919f
C13587 DVSS.n2309 VSS 1.17505f
C13588 DVSS.n2310 VSS 0.17198f
C13589 DVSS.n2311 VSS 0.291498f
C13590 DVSS.n2312 VSS 0.032428f
C13591 DVSS.n2313 VSS 0.046022f
C13592 DVSS.n2314 VSS 0.092043f
C13593 DVSS.n2315 VSS 0.092043f
C13594 DVSS.n2316 VSS 0.092043f
C13595 DVSS.n2317 VSS 0.046022f
C13596 DVSS.n2318 VSS 0.046022f
C13597 DVSS.n2319 VSS 0.046022f
C13598 DVSS.n2320 VSS 0.007166f
C13599 DVSS.n2321 VSS 0.005703f
C13600 DVSS.n2322 VSS 0.011101f
C13601 DVSS.n2323 VSS 0.00545f
C13602 DVSS.n2324 VSS 0.00545f
C13603 DVSS.n2325 VSS 0.007166f
C13604 DVSS.n2326 VSS 0.011101f
C13605 DVSS.n2327 VSS 0.011101f
C13606 DVSS.n2328 VSS 0.011101f
C13607 DVSS.n2329 VSS 0.00545f
C13608 DVSS.n2330 VSS 0.007331f
C13609 DVSS.n2331 VSS 0.007331f
C13610 DVSS.n2332 VSS 0.00545f
C13611 DVSS.n2333 VSS 0.00555f
C13612 DVSS.n2334 VSS 0.011101f
C13613 DVSS.n2335 VSS 0.00555f
C13614 DVSS.n2336 VSS 0.011101f
C13615 DVSS.n2337 VSS 0.011101f
C13616 DVSS.n2338 VSS 0.005804f
C13617 DVSS.n2339 VSS 0.046022f
C13618 DVSS.n2340 VSS 0.046022f
C13619 DVSS.n2341 VSS 0.092043f
C13620 DVSS.n2342 VSS 0.092043f
C13621 DVSS.n2343 VSS 0.092043f
C13622 DVSS.n2344 VSS 0.092043f
C13623 DVSS.n2345 VSS 0.025279f
C13624 DVSS.n2346 VSS 0.022921f
C13625 DVSS.n2347 VSS 0.02139f
C13626 DVSS.n2348 VSS 0.02139f
C13627 DVSS.n2349 VSS 0.046022f
C13628 DVSS.n2350 VSS 0.046022f
C13629 DVSS.n2351 VSS 0.029322f
C13630 DVSS.n2352 VSS 0.035827f
C13631 DVSS.n2353 VSS 0.025279f
C13632 DVSS.n2354 VSS 0.092043f
C13633 DVSS.n2355 VSS 0.092043f
C13634 DVSS.n2356 VSS 0.092043f
C13635 DVSS.n2357 VSS 0.092043f
C13636 DVSS.n2358 VSS 0.092043f
C13637 DVSS.n2359 VSS 0.092043f
C13638 DVSS.n2360 VSS 0.025279f
C13639 DVSS.n2362 VSS 0.045373f
C13640 DVSS.n2364 VSS 0.045373f
C13641 DVSS.n2366 VSS 0.029322f
C13642 DVSS.n2367 VSS 0.045373f
C13643 DVSS.n2368 VSS 0.02139f
C13644 DVSS.n2369 VSS 0.009602f
C13645 DVSS.n2370 VSS 0.046022f
C13646 DVSS.n2371 VSS 0.046022f
C13647 DVSS.n2372 VSS 0.046022f
C13648 DVSS.n2373 VSS 0.092043f
C13649 DVSS.n2374 VSS 0.092043f
C13650 DVSS.n2375 VSS 0.092043f
C13651 DVSS.n2376 VSS 0.092043f
C13652 DVSS.n2377 VSS 0.092043f
C13653 DVSS.n2378 VSS 0.092043f
C13654 DVSS.n2379 VSS 0.092043f
C13655 DVSS.n2380 VSS 0.092043f
C13656 DVSS.n2381 VSS 0.092043f
C13657 DVSS.n2382 VSS 0.092043f
C13658 DVSS.n2383 VSS 0.092043f
C13659 DVSS.n2384 VSS 0.092043f
C13660 DVSS.n2385 VSS 0.092043f
C13661 DVSS.n2386 VSS 0.092043f
C13662 DVSS.n2387 VSS 0.092043f
C13663 DVSS.n2388 VSS 0.092043f
C13664 DVSS.n2389 VSS 0.092043f
C13665 DVSS.n2390 VSS 0.092043f
C13666 DVSS.n2391 VSS 0.092043f
C13667 DVSS.n2392 VSS 0.092043f
C13668 DVSS.n2393 VSS 0.092043f
C13669 DVSS.n2394 VSS 0.092043f
C13670 DVSS.n2395 VSS 0.092043f
C13671 DVSS.n2396 VSS 0.092043f
C13672 DVSS.n2397 VSS 0.092043f
C13673 DVSS.n2398 VSS 0.092043f
C13674 DVSS.n2399 VSS 0.092043f
C13675 DVSS.n2400 VSS 0.092043f
C13676 DVSS.n2401 VSS 0.092043f
C13677 DVSS.n2402 VSS 0.092043f
C13678 DVSS.n2403 VSS 0.092043f
C13679 DVSS.n2404 VSS 0.092043f
C13680 DVSS.n2405 VSS 0.092043f
C13681 DVSS.n2406 VSS 0.092043f
C13682 DVSS.n2407 VSS 0.082968f
C13683 DVSS.n2408 VSS 0.047318f
C13684 DVSS.n2409 VSS 0.121157f
C13685 DVSS.n2410 VSS 0.443616f
C13686 DVSS.n2411 VSS 0.082968f
C13687 DVSS.n2412 VSS 0.092043f
C13688 DVSS.n2413 VSS 0.092043f
C13689 DVSS.n2414 VSS 0.092043f
C13690 DVSS.n2415 VSS 0.092043f
C13691 DVSS.n2416 VSS 0.092043f
C13692 DVSS.n2417 VSS 0.092043f
C13693 DVSS.n2418 VSS 0.092043f
C13694 DVSS.n2419 VSS 0.092043f
C13695 DVSS.n2420 VSS 0.092043f
C13696 DVSS.n2421 VSS 0.092043f
C13697 DVSS.n2422 VSS 0.092043f
C13698 DVSS.n2423 VSS 0.092043f
C13699 DVSS.n2424 VSS 0.092043f
C13700 DVSS.n2425 VSS 0.092043f
C13701 DVSS.n2426 VSS 0.092043f
C13702 DVSS.n2427 VSS 0.092043f
C13703 DVSS.n2428 VSS 0.092043f
C13704 DVSS.n2429 VSS 0.092043f
C13705 DVSS.n2430 VSS 0.092043f
C13706 DVSS.n2431 VSS 0.092043f
C13707 DVSS.n2432 VSS 0.092043f
C13708 DVSS.n2433 VSS 0.092043f
C13709 DVSS.n2434 VSS 0.092043f
C13710 DVSS.n2435 VSS 0.092043f
C13711 DVSS.n2436 VSS 0.092043f
C13712 DVSS.n2437 VSS 0.092043f
C13713 DVSS.n2438 VSS 0.092043f
C13714 DVSS.n2439 VSS 0.092043f
C13715 DVSS.n2440 VSS 0.092043f
C13716 DVSS.n2441 VSS 0.092043f
C13717 DVSS.n2442 VSS 0.092043f
C13718 DVSS.n2443 VSS 0.092043f
C13719 DVSS.n2444 VSS 0.092043f
C13720 DVSS.n2445 VSS 0.092043f
C13721 DVSS.n2446 VSS 0.092043f
C13722 DVSS.n2447 VSS 0.092043f
C13723 DVSS.n2448 VSS 0.092043f
C13724 DVSS.n2449 VSS 0.092043f
C13725 DVSS.n2450 VSS 0.092043f
C13726 DVSS.n2451 VSS 0.092043f
C13727 DVSS.n2452 VSS 0.092043f
C13728 DVSS.n2453 VSS 0.092043f
C13729 DVSS.n2454 VSS 0.092043f
C13730 DVSS.n2455 VSS 0.092043f
C13731 DVSS.n2456 VSS 0.092043f
C13732 DVSS.n2457 VSS 0.092043f
C13733 DVSS.n2458 VSS 0.092043f
C13734 DVSS.n2459 VSS 0.092043f
C13735 DVSS.n2460 VSS 0.092043f
C13736 DVSS.n2461 VSS 0.092043f
C13737 DVSS.n2462 VSS 0.092043f
C13738 DVSS.n2463 VSS 0.092043f
C13739 DVSS.n2464 VSS 0.092043f
C13740 DVSS.n2465 VSS 0.092043f
C13741 DVSS.n2466 VSS 0.092043f
C13742 DVSS.n2467 VSS 0.092043f
C13743 DVSS.n2468 VSS 0.085561f
C13744 DVSS.n2469 VSS 0.092043f
C13745 DVSS.n2470 VSS 0.092043f
C13746 DVSS.n2471 VSS 0.046022f
C13747 DVSS.n2472 VSS 0.046022f
C13748 DVSS.n2473 VSS 0.00555f
C13749 DVSS.n2474 VSS 0.040188f
C13750 DVSS.n2475 VSS 0.006482f
C13751 DVSS.n2476 VSS 0.009456f
C13752 DVSS.n2477 VSS 0.00545f
C13753 DVSS.n2478 VSS 0.011101f
C13754 DVSS.n2479 VSS 0.006813f
C13755 DVSS.n2480 VSS 0.00545f
C13756 DVSS.n2481 VSS 0.007166f
C13757 DVSS.n2482 VSS 0.011101f
C13758 DVSS.n2483 VSS 0.012231f
C13759 DVSS.n2484 VSS 0.006056f
C13760 DVSS.n2485 VSS 0.009234f
C13761 DVSS.n2486 VSS 0.010227f
C13762 DVSS.n2487 VSS 0.006321f
C13763 DVSS.n2488 VSS 0.00555f
C13764 DVSS.n2489 VSS 0.009405f
C13765 DVSS.n2490 VSS 0.01033f
C13766 DVSS.n2491 VSS 0.007298f
C13767 DVSS.n2492 VSS 0.00555f
C13768 DVSS.n2493 VSS 0.007298f
C13769 DVSS.n2494 VSS 0.00555f
C13770 DVSS.n2495 VSS 0.005859f
C13771 DVSS.n2496 VSS 0.011101f
C13772 DVSS.n2497 VSS 0.008171f
C13773 DVSS.n2498 VSS 0.008171f
C13774 DVSS.n2499 VSS 0.003649f
C13775 DVSS.n2500 VSS 0.008634f
C13776 DVSS.n2501 VSS 0.003649f
C13777 DVSS.n2502 VSS 0.004779f
C13778 DVSS.n2503 VSS 0.006482f
C13779 DVSS.n2504 VSS 0.046022f
C13780 DVSS.n2505 VSS 0.092043f
C13781 DVSS.n2506 VSS 0.092043f
C13782 DVSS.n2507 VSS 0.092043f
C13783 DVSS.n2508 VSS 0.092043f
C13784 DVSS.n2509 VSS 0.092043f
C13785 DVSS.n2510 VSS 0.046022f
C13786 DVSS.n2511 VSS 0.046022f
C13787 DVSS.n2512 VSS 0.00545f
C13788 DVSS.n2513 VSS 0.007166f
C13789 DVSS.n2514 VSS 0.011101f
C13790 DVSS.n2515 VSS 0.011101f
C13791 DVSS.n2516 VSS 0.007015f
C13792 DVSS.n2517 VSS 0.015895f
C13793 DVSS.n2518 VSS 0.006308f
C13794 DVSS.n2519 VSS 0.011101f
C13795 DVSS.n2520 VSS 0.011101f
C13796 DVSS.n2521 VSS 0.011101f
C13797 DVSS.n2522 VSS 0.006914f
C13798 DVSS.n2523 VSS 0.00545f
C13799 DVSS.n2524 VSS 0.046022f
C13800 DVSS.n2525 VSS 0.046022f
C13801 DVSS.n2526 VSS 0.092043f
C13802 DVSS.n2527 VSS 0.092043f
C13803 DVSS.n2528 VSS 0.092043f
C13804 DVSS.n2529 VSS 0.092043f
C13805 DVSS.n2530 VSS 0.092043f
C13806 DVSS.n2531 VSS 0.035975f
C13807 DVSS.n2532 VSS 0.045373f
C13808 DVSS.n2533 VSS 0.019279f
C13809 DVSS.n2534 VSS 0.007889f
C13810 DVSS.n2535 VSS 0.015779f
C13811 DVSS.n2536 VSS 0.007889f
C13812 DVSS.n2537 VSS 0.016501f
C13813 DVSS.n2538 VSS 0.102854f
C13814 DVSS.n2539 VSS 0.07864f
C13815 DVSS.n2540 VSS 0.090023f
C13816 DVSS.n2541 VSS 0.144312f
C13817 DVSS.n2542 VSS 0.189694f
C13818 DVSS.n2543 VSS 0.167035f
C13819 DVSS.n2544 VSS 0.088697f
C13820 DVSS.n2545 VSS 0.009456f
C13821 DVSS.n2546 VSS 0.014483f
C13822 DVSS.n2547 VSS 0.199919f
C13823 DVSS.n2548 VSS 1.17505f
C13824 DVSS.n2549 VSS 0.171951f
C13825 DVSS.n2550 VSS 0.292234f
C13826 DVSS.n2551 VSS 0.027752f
C13827 DVSS.n2552 VSS 0.019426f
C13828 DVSS.n2553 VSS 0.003945f
C13829 DVSS.n2554 VSS 0.006556f
C13830 DVSS.n2555 VSS 0.003945f
C13831 DVSS.n2556 VSS 0.005167f
C13832 DVSS.n2557 VSS 0.010695f
C13833 DVSS.n2558 VSS 0.04667f
C13834 DVSS.n2559 VSS 0.092043f
C13835 DVSS.n2560 VSS 0.092043f
C13836 DVSS.n2561 VSS 0.092043f
C13837 DVSS.n2562 VSS 0.092043f
C13838 DVSS.n2563 VSS 0.092043f
C13839 DVSS.n2564 VSS 0.091395f
C13840 DVSS.n2565 VSS 0.005167f
C13841 DVSS.n2566 VSS 0.046022f
C13842 DVSS.n2567 VSS 0.012334f
C13843 DVSS.n2568 VSS 0.003945f
C13844 DVSS.n2569 VSS 0.006404f
C13845 DVSS.n2570 VSS 0.003078f
C13846 DVSS.n2571 VSS 0.011101f
C13847 DVSS.n2572 VSS 0.011101f
C13848 DVSS.n2573 VSS 0.007166f
C13849 DVSS.n2574 VSS 0.00545f
C13850 DVSS.n2575 VSS 0.046022f
C13851 DVSS.n2576 VSS 0.046022f
C13852 DVSS.n2577 VSS 0.092043f
C13853 DVSS.n2578 VSS 0.092043f
C13854 DVSS.n2579 VSS 0.092043f
C13855 DVSS.n2580 VSS 0.092043f
C13856 DVSS.n2581 VSS 0.092043f
C13857 DVSS.n2582 VSS 0.046022f
C13858 DVSS.n2583 VSS 0.009602f
C13859 DVSS.n2584 VSS 0.046022f
C13860 DVSS.n2585 VSS 0.022921f
C13861 DVSS.n2586 VSS 0.007331f
C13862 DVSS.n2587 VSS 0.015895f
C13863 DVSS.n2588 VSS 0.006207f
C13864 DVSS.n2589 VSS 0.011101f
C13865 DVSS.n2590 VSS 0.011101f
C13866 DVSS.n2591 VSS 0.00555f
C13867 DVSS.n2592 VSS 0.011101f
C13868 DVSS.n2593 VSS 0.00555f
C13869 DVSS.n2594 VSS 0.011101f
C13870 DVSS.n2595 VSS 0.012231f
C13871 DVSS.n2596 VSS 0.007166f
C13872 DVSS.n2597 VSS 0.006561f
C13873 DVSS.n2598 VSS 0.046022f
C13874 DVSS.n2599 VSS 0.005834f
C13875 DVSS.n2600 VSS 0.092043f
C13876 DVSS.n2601 VSS 0.092043f
C13877 DVSS.n2602 VSS 0.092043f
C13878 DVSS.n2603 VSS 0.092043f
C13879 DVSS.n2604 VSS 0.092043f
C13880 DVSS.n2605 VSS 0.086858f
C13881 DVSS.n2606 VSS 0.092043f
C13882 DVSS.n2607 VSS 0.092043f
C13883 DVSS.n2608 VSS 0.092043f
C13884 DVSS.n2609 VSS 0.092043f
C13885 DVSS.n2610 VSS 0.092043f
C13886 DVSS.n2611 VSS 2.35092f
C13887 DVSS.n2612 VSS 0.092043f
C13888 DVSS.n2613 VSS 0.312388f
C13889 DVSS.n2614 VSS 0.075514f
C13890 DVSS.n2615 VSS 2.06844f
C13891 DVSS.n2616 VSS 0.02462f
C13892 DVSS.t137 VSS 0.112435f
C13893 DVSS.n2617 VSS 0.318115f
C13894 DVSS.n2618 VSS 0.048117f
C13895 DVSS.n2619 VSS 0.03317f
C13896 DVSS.n2620 VSS 0.306187f
C13897 DVSS.n2621 VSS 0.411753f
C13898 DVSS.n2622 VSS 1.20071f
C13899 DVSS.n2623 VSS 0.016916f
C13900 DVSS.n2624 VSS 0.201862f
C13901 DVSS.n2625 VSS 0.172093f
C13902 DVSS.t20 VSS 0.00963f
C13903 DVSS.t22 VSS 0.00963f
C13904 DVSS.n2626 VSS 0.020417f
C13905 DVSS.n2627 VSS 0.006797f
C13906 DVSS.t169 VSS 0.204005f
C13907 DVSS.n2628 VSS 0.209143f
C13908 DVSS.n2629 VSS 0.029493f
C13909 DVSS.n2630 VSS 0.211534f
C13910 DVSS.n2631 VSS 0.320579f
C13911 DVSS.n2632 VSS 0.023106f
C13912 DVSS.t21 VSS 0.222687f
C13913 DVSS.n2633 VSS 0.319474f
C13914 DVSS.n2634 VSS 0.123472f
C13915 DVSS.n2635 VSS 0.04066f
C13916 DVSS.n2636 VSS 0.094244f
C13917 DVSS.n2637 VSS 0.036474f
C13918 DVSS.n2638 VSS 0.071185f
C13919 DVSS.n2639 VSS 0.038276f
C13920 DVSS.t117 VSS 0.255567f
C13921 DVSS.n2640 VSS 0.012655f
C13922 DVSS.t139 VSS 0.255567f
C13923 DVSS.n2641 VSS 0.289941f
C13924 DVSS.n2642 VSS 0.023111f
C13925 DVSS.n2643 VSS 0.036474f
C13926 DVSS.n2644 VSS 0.289941f
C13927 DVSS.t63 VSS 0.222687f
C13928 DVSS.t16 VSS 0.222687f
C13929 DVSS.n2645 VSS 0.391791f
C13930 DVSS.t144 VSS 0.272754f
C13931 DVSS.t142 VSS 0.226423f
C13932 DVSS.n2646 VSS 0.017444f
C13933 DVSS.n2647 VSS 0.016457f
C13934 DVSS.n2648 VSS 0.020503f
C13935 DVSS.n2649 VSS 0.0172f
C13936 DVSS.n2650 VSS -0.054143f
C13937 DVSS.n2651 VSS 0.168036f
C13938 DVSS.n2652 VSS 0.387185f
C13939 DVSS.n2653 VSS 0.547223f
C13940 DVSS.n2654 VSS 0.511134f
C13941 DVSS.n2655 VSS 0.478254f
C13942 DVSS.n2656 VSS 0.036474f
C13943 DVSS.n2657 VSS 0.033005f
C13944 DVSS.n2658 VSS 0.012655f
C13945 DVSS.n2659 VSS 0.054676f
C13946 DVSS.n2660 VSS 0.283216f
C13947 DVSS.n2661 VSS 0.017649f
C13948 DVSS.n2662 VSS 0.030479f
C13949 DVSS.n2663 VSS 0.426987f
C13950 DVSS.n2664 VSS 2.08413f
C13951 DVSS.t58 VSS 0.061846f
C13952 DVSS.n2665 VSS 0.163721f
C13953 DVSS.n2666 VSS 0.023309f
C13954 DVSS.n2667 VSS 0.71504f
C13955 DVSS.n2668 VSS 0.010501f
C13956 DVSS.n2669 VSS 0.042011f
C13957 DVSS.n2670 VSS 0.042011f
C13958 DVSS.n2671 VSS 0.019808f
C13959 DVSS.n2672 VSS 0.011667f
C13960 DVSS.n2673 VSS 0.011749f
C13961 DVSS.n2674 VSS 0.018986f
C13962 DVSS.n2675 VSS 0.010334f
C13963 DVSS.n2676 VSS 0.011834f
C13964 DVSS.n2677 VSS 0.042011f
C13965 DVSS.n2678 VSS 0.010334f
C13966 DVSS.n2679 VSS 0.042011f
C13967 DVSS.n2680 VSS 0.084022f
C13968 DVSS.n2681 VSS 1.00462f
C13969 DVSS.n2682 VSS 0.220678f
C13970 DVSS.n2683 VSS 0.084022f
C13971 DVSS.n2684 VSS 0.814397f
C13972 DVSS.n2685 VSS 0.084022f
C13973 DVSS.n2686 VSS 0.084022f
C13974 DVSS.n2687 VSS 0.084022f
C13975 DVSS.n2688 VSS 0.084022f
C13976 DVSS.n2689 VSS 0.010334f
C13977 DVSS.n2690 VSS 0.042011f
C13978 DVSS.n2691 VSS 0.010334f
C13979 DVSS.n2692 VSS 0.011834f
C13980 DVSS.n2693 VSS 0.010334f
C13981 DVSS.n2694 VSS 0.015978f
C13982 DVSS.n2695 VSS 0.023309f
C13983 DVSS.n2696 VSS 0.011834f
C13984 DVSS.n2697 VSS 0.042011f
C13985 DVSS.n2698 VSS 0.010334f
C13986 DVSS.n2699 VSS 0.042011f
C13987 DVSS.n2700 VSS 0.084022f
C13988 DVSS.n2701 VSS 0.084022f
C13989 DVSS.n2702 VSS 0.084022f
C13990 DVSS.n2703 VSS 0.084022f
C13991 DVSS.n2704 VSS 0.084022f
C13992 DVSS.n2705 VSS 0.084022f
C13993 DVSS.n2706 VSS 0.010334f
C13994 DVSS.n2707 VSS 0.042011f
C13995 DVSS.n2708 VSS 0.011834f
C13996 DVSS.n2709 VSS 0.010334f
C13997 DVSS.n2710 VSS 0.020668f
C13998 DVSS.n2711 VSS 0.023309f
C13999 DVSS.n2712 VSS 0.019549f
C14000 DVSS.t49 VSS 0.061846f
C14001 DVSS.n2713 VSS 0.021475f
C14002 DVSS.n2714 VSS 0.011834f
C14003 DVSS.n2715 VSS 0.042011f
C14004 DVSS.n2716 VSS 0.010334f
C14005 DVSS.n2717 VSS 0.042011f
C14006 DVSS.n2718 VSS 0.084022f
C14007 DVSS.n2719 VSS 0.084022f
C14008 DVSS.n2720 VSS 0.084022f
C14009 DVSS.n2721 VSS 0.084022f
C14010 DVSS.n2722 VSS 0.084022f
C14011 DVSS.n2723 VSS 0.084022f
C14012 DVSS.n2724 VSS 0.010334f
C14013 DVSS.n2725 VSS 0.042011f
C14014 DVSS.n2726 VSS 0.010334f
C14015 DVSS.n2727 VSS 0.011834f
C14016 DVSS.n2728 VSS 0.010334f
C14017 DVSS.n2729 VSS 0.022275f
C14018 DVSS.n2730 VSS 0.023309f
C14019 DVSS.n2731 VSS 0.019433f
C14020 DVSS.n2732 VSS 0.010334f
C14021 DVSS.n2733 VSS 0.023309f
C14022 DVSS.n2734 VSS 0.011834f
C14023 DVSS.n2735 VSS 0.042011f
C14024 DVSS.n2736 VSS 0.010334f
C14025 DVSS.n2737 VSS 0.042011f
C14026 DVSS.n2738 VSS 0.084022f
C14027 DVSS.n2739 VSS 0.084022f
C14028 DVSS.n2740 VSS 0.084022f
C14029 DVSS.n2741 VSS 0.084022f
C14030 DVSS.n2742 VSS 0.010334f
C14031 DVSS.n2743 VSS 0.042011f
C14032 DVSS.n2744 VSS 0.010334f
C14033 DVSS.n2745 VSS 0.011834f
C14034 DVSS.n2746 VSS 0.010334f
C14035 DVSS.n2747 VSS 0.023309f
C14036 DVSS.t55 VSS 0.061846f
C14037 DVSS.n2748 VSS 0.021475f
C14038 DVSS.n2749 VSS 0.011834f
C14039 DVSS.n2750 VSS 0.042011f
C14040 DVSS.n2751 VSS 0.010334f
C14041 DVSS.n2752 VSS 0.042011f
C14042 DVSS.n2753 VSS 0.084022f
C14043 DVSS.n2754 VSS 0.084022f
C14044 DVSS.n2755 VSS 0.084022f
C14045 DVSS.n2756 VSS 0.084022f
C14046 DVSS.n2757 VSS 0.084022f
C14047 DVSS.n2758 VSS 0.084022f
C14048 DVSS.n2759 VSS 0.010334f
C14049 DVSS.n2760 VSS 0.042011f
C14050 DVSS.n2761 VSS 0.010667f
C14051 DVSS.n2762 VSS 0.010334f
C14052 DVSS.n2763 VSS 0.014286f
C14053 DVSS.n2764 VSS 0.010334f
C14054 DVSS.n2765 VSS 0.011501f
C14055 DVSS.n2766 VSS 0.013816f
C14056 DVSS.n2767 VSS 0.021147f
C14057 DVSS.n2768 VSS 0.021241f
C14058 DVSS.n2769 VSS 0.011834f
C14059 DVSS.n2770 VSS 0.042011f
C14060 DVSS.n2771 VSS 0.010334f
C14061 DVSS.n2772 VSS 0.042011f
C14062 DVSS.n2773 VSS 0.084022f
C14063 DVSS.n2774 VSS 0.084022f
C14064 DVSS.n2775 VSS 0.084022f
C14065 DVSS.n2776 VSS 0.084022f
C14066 DVSS.n2777 VSS 0.084022f
C14067 DVSS.n2778 VSS 0.084022f
C14068 DVSS.n2779 VSS 0.010334f
C14069 DVSS.n2780 VSS 0.042011f
C14070 DVSS.n2781 VSS 0.010334f
C14071 DVSS.n2782 VSS 0.011834f
C14072 DVSS.n2783 VSS 0.010334f
C14073 DVSS.n2784 VSS 0.013722f
C14074 DVSS.n2785 VSS 0.023309f
C14075 DVSS.n2786 VSS 0.011334f
C14076 DVSS.n2787 VSS 0.042011f
C14077 DVSS.n2788 VSS 0.010334f
C14078 DVSS.n2789 VSS 0.042011f
C14079 DVSS.n2790 VSS 0.084022f
C14080 DVSS.n2791 VSS 0.084022f
C14081 DVSS.n2792 VSS 0.084022f
C14082 DVSS.n2793 VSS 0.084022f
C14083 DVSS.n2794 VSS 0.084022f
C14084 DVSS.n2795 VSS 0.084022f
C14085 DVSS.n2796 VSS 0.010334f
C14086 DVSS.n2797 VSS 0.042011f
C14087 DVSS.n2798 VSS 0.011834f
C14088 DVSS.n2799 VSS 0.010334f
C14089 DVSS.n2800 VSS 0.010334f
C14090 DVSS.n2801 VSS 0.010834f
C14091 DVSS.n2802 VSS 0.023309f
C14092 DVSS.n2803 VSS 0.021805f
C14093 DVSS.t51 VSS 0.061846f
C14094 DVSS.n2804 VSS 0.021475f
C14095 DVSS.n2805 VSS 0.011834f
C14096 DVSS.n2806 VSS 0.042011f
C14097 DVSS.n2807 VSS 0.010334f
C14098 DVSS.n2808 VSS 0.042011f
C14099 DVSS.n2809 VSS 0.084022f
C14100 DVSS.n2810 VSS 0.084022f
C14101 DVSS.n2811 VSS 0.084022f
C14102 DVSS.n2812 VSS 0.084022f
C14103 DVSS.n2813 VSS 0.084022f
C14104 DVSS.n2814 VSS 0.084022f
C14105 DVSS.n2815 VSS 0.010334f
C14106 DVSS.n2816 VSS 0.042011f
C14107 DVSS.n2817 VSS 0.010334f
C14108 DVSS.n2818 VSS 0.011834f
C14109 DVSS.n2819 VSS 0.010334f
C14110 DVSS.n2820 VSS 0.020019f
C14111 DVSS.n2821 VSS 0.023309f
C14112 DVSS.n2822 VSS 0.010715f
C14113 DVSS.n2823 VSS 0.010334f
C14114 DVSS.n2824 VSS 0.01088f
C14115 DVSS.n2825 VSS 0.023309f
C14116 DVSS.n2826 VSS 0.011834f
C14117 DVSS.n2827 VSS 0.042011f
C14118 DVSS.n2828 VSS 0.010334f
C14119 DVSS.n2829 VSS 0.042011f
C14120 DVSS.n2830 VSS 0.084022f
C14121 DVSS.n2831 VSS 0.084022f
C14122 DVSS.n2832 VSS 0.084022f
C14123 DVSS.n2833 VSS 0.084022f
C14124 DVSS.n2834 VSS 0.010334f
C14125 DVSS.n2835 VSS 0.042011f
C14126 DVSS.n2836 VSS 0.010334f
C14127 DVSS.n2837 VSS 0.011834f
C14128 DVSS.n2838 VSS 0.010334f
C14129 DVSS.n2839 VSS 0.023309f
C14130 DVSS.t59 VSS 0.061846f
C14131 DVSS.n2840 VSS 0.021475f
C14132 DVSS.n2841 VSS 0.011834f
C14133 DVSS.n2842 VSS 0.042011f
C14134 DVSS.n2843 VSS 0.010334f
C14135 DVSS.n2844 VSS 0.042011f
C14136 DVSS.n2845 VSS 0.084022f
C14137 DVSS.n2846 VSS 0.084022f
C14138 DVSS.n2847 VSS 0.084022f
C14139 DVSS.n2848 VSS 0.084022f
C14140 DVSS.n2849 VSS 0.084022f
C14141 DVSS.n2850 VSS 0.084022f
C14142 DVSS.n2851 VSS 0.010334f
C14143 DVSS.n2852 VSS 0.042011f
C14144 DVSS.n2853 VSS 0.011167f
C14145 DVSS.n2854 VSS 0.010334f
C14146 DVSS.n2855 VSS 0.01203f
C14147 DVSS.n2856 VSS 0.010334f
C14148 DVSS.n2857 VSS 0.011001f
C14149 DVSS.n2858 VSS 0.016072f
C14150 DVSS.n2859 VSS 0.018892f
C14151 DVSS.n2860 VSS 0.023309f
C14152 DVSS.n2861 VSS 0.011834f
C14153 DVSS.n2862 VSS 0.042011f
C14154 DVSS.n2863 VSS 0.010334f
C14155 DVSS.n2864 VSS 0.042011f
C14156 DVSS.n2865 VSS 0.084022f
C14157 DVSS.n2866 VSS 0.084022f
C14158 DVSS.n2867 VSS 0.084022f
C14159 DVSS.n2868 VSS 0.084022f
C14160 DVSS.n2869 VSS 0.084022f
C14161 DVSS.n2870 VSS 0.084022f
C14162 DVSS.n2871 VSS 0.010334f
C14163 DVSS.n2872 VSS 0.042011f
C14164 DVSS.n2873 VSS 0.010334f
C14165 DVSS.n2874 VSS 0.011834f
C14166 DVSS.n2875 VSS 0.010334f
C14167 DVSS.n2876 VSS 0.011842f
C14168 DVSS.n2877 VSS 0.019433f
C14169 DVSS.n2878 VSS 0.023309f
C14170 DVSS.n2879 VSS 0.010834f
C14171 DVSS.n2880 VSS 0.042011f
C14172 DVSS.n2881 VSS 0.010334f
C14173 DVSS.n2882 VSS 0.042011f
C14174 DVSS.n2883 VSS 0.084022f
C14175 DVSS.n2884 VSS 0.084022f
C14176 DVSS.n2885 VSS 0.084022f
C14177 DVSS.n2886 VSS 0.084022f
C14178 DVSS.n2887 VSS 0.084022f
C14179 DVSS.n2888 VSS 0.084022f
C14180 DVSS.n2889 VSS 0.010334f
C14181 DVSS.n2890 VSS 0.042011f
C14182 DVSS.n2891 VSS 0.011834f
C14183 DVSS.n2892 VSS 0.010334f
C14184 DVSS.n2893 VSS 0.010334f
C14185 DVSS.n2894 VSS 0.011334f
C14186 DVSS.n2895 VSS 0.023309f
C14187 DVSS.n2896 VSS 0.023309f
C14188 DVSS.n2897 VSS 0.011834f
C14189 DVSS.n2898 VSS 0.042011f
C14190 DVSS.n2899 VSS 0.010334f
C14191 DVSS.n2900 VSS 0.042011f
C14192 DVSS.n2901 VSS 0.084022f
C14193 DVSS.n2902 VSS 0.084022f
C14194 DVSS.n2903 VSS 0.084022f
C14195 DVSS.n2904 VSS 0.084022f
C14196 DVSS.n2905 VSS 0.084022f
C14197 DVSS.n2906 VSS 0.084022f
C14198 DVSS.n2907 VSS 0.010334f
C14199 DVSS.n2908 VSS 0.042011f
C14200 DVSS.n2909 VSS 0.010334f
C14201 DVSS.n2910 VSS 0.011834f
C14202 DVSS.n2911 VSS 0.010334f
C14203 DVSS.n2912 VSS 0.017764f
C14204 DVSS.n2913 VSS 0.023309f
C14205 DVSS.n2914 VSS 0.01297f
C14206 DVSS.n2915 VSS 0.011834f
C14207 DVSS.n2916 VSS 0.042011f
C14208 DVSS.n2917 VSS 0.010334f
C14209 DVSS.n2918 VSS 0.042011f
C14210 DVSS.n2919 VSS 0.084022f
C14211 DVSS.n2920 VSS 0.084022f
C14212 DVSS.n2921 VSS 0.084022f
C14213 DVSS.n2922 VSS 0.084022f
C14214 DVSS.n2923 VSS 0.084022f
C14215 DVSS.n2924 VSS 0.084022f
C14216 DVSS.n2925 VSS 0.010334f
C14217 DVSS.n2926 VSS 0.042011f
C14218 DVSS.n2927 VSS 0.010334f
C14219 DVSS.n2928 VSS 0.011834f
C14220 DVSS.n2929 VSS 0.010334f
C14221 DVSS.n2930 VSS 0.023309f
C14222 DVSS.n2931 VSS 0.023309f
C14223 DVSS.n2932 VSS 0.011834f
C14224 DVSS.n2933 VSS 0.042011f
C14225 DVSS.n2934 VSS 0.010334f
C14226 DVSS.n2935 VSS 0.042011f
C14227 DVSS.n2936 VSS 0.084022f
C14228 DVSS.n2937 VSS 0.084022f
C14229 DVSS.n2938 VSS 0.084022f
C14230 DVSS.n2939 VSS 0.084022f
C14231 DVSS.n2940 VSS 0.084022f
C14232 DVSS.n2941 VSS 0.084022f
C14233 DVSS.n2942 VSS 0.010334f
C14234 DVSS.n2943 VSS 0.042011f
C14235 DVSS.n2944 VSS 0.010334f
C14236 DVSS.n2945 VSS 0.011834f
C14237 DVSS.n2946 VSS 0.011667f
C14238 DVSS.n2947 VSS 0.013534f
C14239 DVSS.t56 VSS 0.061846f
C14240 DVSS.n2948 VSS 0.021475f
C14241 DVSS.n2949 VSS 0.023309f
C14242 DVSS.n2950 VSS 0.010334f
C14243 DVSS.n2951 VSS 0.011834f
C14244 DVSS.n2952 VSS 0.042011f
C14245 DVSS.n2953 VSS 0.010334f
C14246 DVSS.n2954 VSS 0.042011f
C14247 DVSS.n2955 VSS 0.084022f
C14248 DVSS.n2956 VSS 0.084022f
C14249 DVSS.n2957 VSS 0.084022f
C14250 DVSS.n2958 VSS 0.084022f
C14251 DVSS.n2959 VSS 0.084022f
C14252 DVSS.n2960 VSS 0.084022f
C14253 DVSS.n2961 VSS 0.010334f
C14254 DVSS.n2962 VSS 0.042011f
C14255 DVSS.n2963 VSS 0.010334f
C14256 DVSS.n2964 VSS 0.011834f
C14257 DVSS.n2965 VSS 0.010334f
C14258 DVSS.n2966 VSS 0.023309f
C14259 DVSS.n2967 VSS 0.023309f
C14260 DVSS.n2968 VSS 0.011834f
C14261 DVSS.n2969 VSS 0.042011f
C14262 DVSS.n2970 VSS 0.010334f
C14263 DVSS.n2971 VSS 0.042011f
C14264 DVSS.n2972 VSS 0.084022f
C14265 DVSS.n2973 VSS 0.084022f
C14266 DVSS.n2974 VSS 0.084022f
C14267 DVSS.n2975 VSS 0.084022f
C14268 DVSS.n2976 VSS 0.084022f
C14269 DVSS.n2977 VSS 0.084022f
C14270 DVSS.n2978 VSS 0.010334f
C14271 DVSS.n2979 VSS 0.042011f
C14272 DVSS.n2980 VSS 0.011834f
C14273 DVSS.n2981 VSS 0.010334f
C14274 DVSS.n2982 VSS 0.020668f
C14275 DVSS.n2983 VSS 0.023309f
C14276 DVSS.n2984 VSS 0.023309f
C14277 DVSS.t48 VSS 0.061846f
C14278 DVSS.n2985 VSS 0.021475f
C14279 DVSS.n2986 VSS 0.011834f
C14280 DVSS.n2987 VSS 0.042011f
C14281 DVSS.n2988 VSS 0.010334f
C14282 DVSS.n2989 VSS 0.042011f
C14283 DVSS.n2990 VSS 0.084022f
C14284 DVSS.n2991 VSS 0.084022f
C14285 DVSS.n2992 VSS 0.084022f
C14286 DVSS.n2993 VSS 0.084022f
C14287 DVSS.n2994 VSS 0.084022f
C14288 DVSS.n2995 VSS 0.084022f
C14289 DVSS.n2996 VSS 0.084022f
C14290 DVSS.n2997 VSS 0.010334f
C14291 DVSS.n2998 VSS 0.042011f
C14292 DVSS.n2999 VSS 0.010334f
C14293 DVSS.n3000 VSS 0.011834f
C14294 DVSS.n3001 VSS 0.011834f
C14295 DVSS.n3002 VSS 0.010334f
C14296 DVSS.n3003 VSS 0.010501f
C14297 DVSS.n3004 VSS 0.023309f
C14298 DVSS.n3005 VSS 0.019433f
C14299 DVSS.n3006 VSS 0.016636f
C14300 DVSS.n3007 VSS 0.021993f
C14301 DVSS.n3008 VSS 0.019433f
C14302 DVSS.n3009 VSS 0.023309f
C14303 DVSS.n3010 VSS 0.021475f
C14304 DVSS.n3011 VSS 0.023309f
C14305 DVSS.n3012 VSS 0.010334f
C14306 DVSS.n3013 VSS 0.012594f
C14307 DVSS.n3014 VSS 0.011001f
C14308 DVSS.n3015 VSS 0.011834f
C14309 DVSS.n3016 VSS 0.023309f
C14310 DVSS.n3017 VSS 0.019433f
C14311 DVSS.n3018 VSS 0.019433f
C14312 DVSS.n3019 VSS 0.010334f
C14313 DVSS.n3020 VSS 0.01485f
C14314 DVSS.n3021 VSS 0.010501f
C14315 DVSS.n3022 VSS 0.011834f
C14316 DVSS.n3023 VSS 0.023309f
C14317 DVSS.n3024 VSS 0.019433f
C14318 DVSS.n3025 VSS 0.019433f
C14319 DVSS.n3026 VSS 0.023309f
C14320 DVSS.n3027 VSS 0.011667f
C14321 DVSS.n3028 VSS 0.042011f
C14322 DVSS.n3029 VSS 0.010334f
C14323 DVSS.n3030 VSS 0.011834f
C14324 DVSS.n3031 VSS 0.023309f
C14325 DVSS.n3032 VSS 0.018986f
C14326 DVSS.n3033 VSS 0.011834f
C14327 DVSS.n3034 VSS 0.010334f
C14328 DVSS.n3035 VSS 0.011834f
C14329 DVSS.n3036 VSS 0.015978f
C14330 DVSS.n3037 VSS 0.023309f
C14331 DVSS.n3038 VSS 0.011834f
C14332 DVSS.n3039 VSS 0.042011f
C14333 DVSS.n3040 VSS 0.010334f
C14334 DVSS.n3041 VSS 0.011834f
C14335 DVSS.n3042 VSS 0.023309f
C14336 DVSS.n3043 VSS 0.023309f
C14337 DVSS.n3044 VSS 0.011834f
C14338 DVSS.n3045 VSS 0.020668f
C14339 DVSS.n3046 VSS 0.011834f
C14340 DVSS.n3047 VSS 0.019549f
C14341 DVSS.n3048 VSS 0.021475f
C14342 DVSS.n3049 VSS 0.015414f
C14343 DVSS.n3050 VSS 0.011834f
C14344 DVSS.n3051 VSS 0.042011f
C14345 DVSS.n3052 VSS 0.010334f
C14346 DVSS.n3053 VSS 0.011834f
C14347 DVSS.n3054 VSS 0.012688f
C14348 DVSS.n3055 VSS 0.022275f
C14349 DVSS.n3056 VSS 0.011834f
C14350 DVSS.n3057 VSS 0.010334f
C14351 DVSS.n3058 VSS 0.011834f
C14352 DVSS.n3059 VSS 0.023309f
C14353 DVSS.n3060 VSS 0.023309f
C14354 DVSS.n3061 VSS 0.019433f
C14355 DVSS.n3062 VSS 0.020113f
C14356 DVSS.n3063 VSS 0.011667f
C14357 DVSS.n3064 VSS 0.010334f
C14358 DVSS.n3065 VSS 0.042011f
C14359 DVSS.n3066 VSS 0.084022f
C14360 DVSS.n3067 VSS 0.084022f
C14361 DVSS.n3068 VSS 0.084022f
C14362 DVSS.n3069 VSS 0.084022f
C14363 DVSS.n3070 VSS 0.042011f
C14364 DVSS.n3071 VSS 0.042011f
C14365 DVSS.n3072 VSS 0.010334f
C14366 DVSS.n3073 VSS 0.011834f
C14367 DVSS.n3074 VSS 0.023309f
C14368 DVSS.n3075 VSS 0.023309f
C14369 DVSS.n3076 VSS 0.011834f
C14370 DVSS.n3077 VSS 0.010334f
C14371 DVSS.n3078 VSS 0.011834f
C14372 DVSS.n3079 VSS 0.023309f
C14373 DVSS.n3080 VSS 0.023309f
C14374 DVSS.n3081 VSS 0.011834f
C14375 DVSS.n3082 VSS 0.042011f
C14376 DVSS.n3083 VSS 0.010334f
C14377 DVSS.n3084 VSS 0.011834f
C14378 DVSS.n3085 VSS 0.020677f
C14379 DVSS.n3086 VSS 0.021475f
C14380 DVSS.n3087 VSS 0.011834f
C14381 DVSS.n3088 VSS 0.014286f
C14382 DVSS.n3089 VSS 0.013816f
C14383 DVSS.n3090 VSS 0.011501f
C14384 DVSS.n3091 VSS 0.010667f
C14385 DVSS.n3092 VSS 0.021147f
C14386 DVSS.n3093 VSS 0.023309f
C14387 DVSS.n3094 VSS 0.011834f
C14388 DVSS.n3095 VSS 0.042011f
C14389 DVSS.n3096 VSS 0.010334f
C14390 DVSS.n3097 VSS 0.011834f
C14391 DVSS.n3098 VSS 0.023309f
C14392 DVSS.n3099 VSS 0.021241f
C14393 DVSS.n3100 VSS 0.011834f
C14394 DVSS.n3101 VSS 0.010334f
C14395 DVSS.n3102 VSS 0.011834f
C14396 DVSS.n3103 VSS 0.013722f
C14397 DVSS.n3104 VSS 0.023309f
C14398 DVSS.n3105 VSS 0.011834f
C14399 DVSS.n3106 VSS 0.042011f
C14400 DVSS.n3107 VSS 0.010334f
C14401 DVSS.n3108 VSS 0.011834f
C14402 DVSS.n3109 VSS 0.023309f
C14403 DVSS.n3110 VSS 0.023309f
C14404 DVSS.n3111 VSS 0.011334f
C14405 DVSS.n3112 VSS 0.010834f
C14406 DVSS.n3113 VSS 0.010334f
C14407 DVSS.n3114 VSS 0.011834f
C14408 DVSS.n3115 VSS 0.021805f
C14409 DVSS.n3116 VSS 0.021475f
C14410 DVSS.n3117 VSS 0.013158f
C14411 DVSS.n3118 VSS 0.011834f
C14412 DVSS.n3119 VSS 0.042011f
C14413 DVSS.n3120 VSS 0.010334f
C14414 DVSS.n3121 VSS 0.011834f
C14415 DVSS.n3122 VSS 0.014944f
C14416 DVSS.n3123 VSS 0.020019f
C14417 DVSS.n3124 VSS 0.011834f
C14418 DVSS.n3125 VSS 0.010334f
C14419 DVSS.n3126 VSS 0.011834f
C14420 DVSS.n3127 VSS 0.023309f
C14421 DVSS.n3128 VSS 0.023309f
C14422 DVSS.n3129 VSS 0.01088f
C14423 DVSS.n3130 VSS 0.010715f
C14424 DVSS.n3131 VSS 0.020207f
C14425 DVSS.n3132 VSS 0.011167f
C14426 DVSS.n3133 VSS 0.010334f
C14427 DVSS.n3134 VSS 0.042011f
C14428 DVSS.n3135 VSS 0.084022f
C14429 DVSS.n3136 VSS 0.084022f
C14430 DVSS.n3137 VSS 0.084022f
C14431 DVSS.n3138 VSS 0.084022f
C14432 DVSS.n3139 VSS 0.042011f
C14433 DVSS.n3140 VSS 0.042011f
C14434 DVSS.n3141 VSS 0.010334f
C14435 DVSS.n3142 VSS 0.011834f
C14436 DVSS.n3143 VSS 0.023309f
C14437 DVSS.n3144 VSS 0.023309f
C14438 DVSS.n3145 VSS 0.011834f
C14439 DVSS.n3146 VSS 0.010334f
C14440 DVSS.n3147 VSS 0.011834f
C14441 DVSS.n3148 VSS 0.023309f
C14442 DVSS.n3149 VSS 0.023309f
C14443 DVSS.n3150 VSS 0.011834f
C14444 DVSS.n3151 VSS 0.042011f
C14445 DVSS.n3152 VSS 0.010334f
C14446 DVSS.n3153 VSS 0.011834f
C14447 DVSS.n3154 VSS 0.022933f
C14448 DVSS.n3155 VSS 0.021475f
C14449 DVSS.n3156 VSS 0.011834f
C14450 DVSS.n3157 VSS 0.01203f
C14451 DVSS.n3158 VSS 0.016072f
C14452 DVSS.n3159 VSS 0.011001f
C14453 DVSS.n3160 VSS 0.011167f
C14454 DVSS.n3161 VSS 0.018892f
C14455 DVSS.n3162 VSS 0.023309f
C14456 DVSS.n3163 VSS 0.011834f
C14457 DVSS.n3164 VSS 0.042011f
C14458 DVSS.n3165 VSS 0.010334f
C14459 DVSS.n3166 VSS 0.011834f
C14460 DVSS.n3167 VSS 0.023309f
C14461 DVSS.n3168 VSS 0.023309f
C14462 DVSS.n3169 VSS 0.011834f
C14463 DVSS.n3170 VSS 0.010334f
C14464 DVSS.n3171 VSS 0.011834f
C14465 DVSS.n3172 VSS 0.011842f
C14466 DVSS.n3173 VSS 0.019433f
C14467 DVSS.n3174 VSS 0.023121f
C14468 DVSS.n3175 VSS 0.011834f
C14469 DVSS.n3176 VSS 0.042011f
C14470 DVSS.n3177 VSS 0.010334f
C14471 DVSS.n3178 VSS 0.011834f
C14472 DVSS.n3179 VSS 0.023309f
C14473 DVSS.n3180 VSS 0.023309f
C14474 DVSS.n3181 VSS 0.010834f
C14475 DVSS.n3182 VSS 0.011334f
C14476 DVSS.n3183 VSS 0.010334f
C14477 DVSS.n3184 VSS 0.011834f
C14478 DVSS.n3185 VSS 0.023309f
C14479 DVSS.n3186 VSS 0.012406f
C14480 DVSS.n3187 VSS 0.011834f
C14481 DVSS.n3188 VSS 0.042011f
C14482 DVSS.n3189 VSS 0.010334f
C14483 DVSS.n3190 VSS 0.011834f
C14484 DVSS.n3191 VSS 0.016448f
C14485 DVSS.n3192 VSS 0.017764f
C14486 DVSS.n3193 VSS 0.011834f
C14487 DVSS.n3194 VSS 0.010334f
C14488 DVSS.n3195 VSS 0.011834f
C14489 DVSS.n3196 VSS 0.023309f
C14490 DVSS.n3197 VSS 0.023309f
C14491 DVSS.n3198 VSS 0.011834f
C14492 DVSS.n3199 VSS 0.042011f
C14493 DVSS.n3200 VSS 0.010334f
C14494 DVSS.n3201 VSS 0.010667f
C14495 DVSS.n3202 VSS 0.011501f
C14496 DVSS.n3203 VSS 0.01297f
C14497 DVSS.n3204 VSS 0.019433f
C14498 DVSS.n3205 VSS 0.021993f
C14499 DVSS.n3206 VSS 0.011834f
C14500 DVSS.n3207 VSS 0.010334f
C14501 DVSS.n3208 VSS 0.011834f
C14502 DVSS.n3209 VSS 0.023309f
C14503 DVSS.n3210 VSS 0.023309f
C14504 DVSS.n3211 VSS 0.011834f
C14505 DVSS.n3212 VSS 0.042011f
C14506 DVSS.n3213 VSS 0.010334f
C14507 DVSS.n3214 VSS 0.011834f
C14508 DVSS.n3215 VSS 0.023309f
C14509 DVSS.n3216 VSS 0.023309f
C14510 DVSS.n3217 VSS 0.011834f
C14511 DVSS.n3218 VSS 0.010334f
C14512 DVSS.n3219 VSS 0.011834f
C14513 DVSS.n3220 VSS 0.013534f
C14514 DVSS.n3221 VSS 0.021475f
C14515 DVSS.n3222 VSS 0.016448f
C14516 DVSS.n3223 VSS 0.010501f
C14517 DVSS.n3224 VSS 0.011667f
C14518 DVSS.n3225 VSS 0.042011f
C14519 DVSS.n3226 VSS 0.010334f
C14520 DVSS.n3227 VSS 0.011834f
C14521 DVSS.n3228 VSS 0.023309f
C14522 DVSS.n3229 VSS 0.023309f
C14523 DVSS.n3230 VSS 0.011834f
C14524 DVSS.n3231 VSS 0.010334f
C14525 DVSS.n3232 VSS 0.011834f
C14526 DVSS.n3233 VSS 0.023309f
C14527 DVSS.n3234 VSS 0.014098f
C14528 DVSS.n3235 VSS 0.011834f
C14529 DVSS.n3236 VSS 0.042011f
C14530 DVSS.n3237 VSS 0.010334f
C14531 DVSS.n3238 VSS 0.011834f
C14532 DVSS.n3239 VSS 0.020865f
C14533 DVSS.n3240 VSS 0.023309f
C14534 DVSS.n3241 VSS 0.011834f
C14535 DVSS.n3242 VSS 0.020668f
C14536 DVSS.n3243 VSS 0.011834f
C14537 DVSS.n3244 VSS 0.023309f
C14538 DVSS.n3245 VSS 0.023309f
C14539 DVSS.n3246 VSS 0.011834f
C14540 DVSS.n3247 VSS 0.042011f
C14541 DVSS.n3248 VSS 0.010334f
C14542 DVSS.n3249 VSS 0.011834f
C14543 DVSS.n3250 VSS 0.014662f
C14544 DVSS.n3251 VSS 0.021475f
C14545 DVSS.n3252 VSS 0.016448f
C14546 DVSS.n3253 VSS 0.011834f
C14547 DVSS.n3254 VSS 0.010334f
C14548 DVSS.n3255 VSS 0.011834f
C14549 DVSS.n3256 VSS 0.015508f
C14550 DVSS.n3257 VSS 0.023309f
C14551 DVSS.n3258 VSS 0.023309f
C14552 DVSS.n3259 VSS 0.023309f
C14553 DVSS.n3260 VSS 0.011667f
C14554 DVSS.n3261 VSS 0.010334f
C14555 DVSS.n3262 VSS 0.042011f
C14556 DVSS.n3263 VSS 0.042011f
C14557 DVSS.n3264 VSS 0.010334f
C14558 DVSS.n3265 VSS 0.016448f
C14559 DVSS.n3266 VSS 0.015508f
C14560 DVSS.n3267 VSS 0.010501f
C14561 DVSS.n3268 VSS 0.011667f
C14562 DVSS.n3269 VSS 0.023309f
C14563 DVSS.n3270 VSS 0.023309f
C14564 DVSS.n3271 VSS 0.011834f
C14565 DVSS.n3272 VSS 0.010334f
C14566 DVSS.n3273 VSS 0.042011f
C14567 DVSS.n3274 VSS 0.042011f
C14568 DVSS.n3275 VSS 0.084022f
C14569 DVSS.n3276 VSS 0.084022f
C14570 DVSS.n3277 VSS 0.042011f
C14571 DVSS.n3278 VSS 0.042011f
C14572 DVSS.n3279 VSS 0.010334f
C14573 DVSS.n3280 VSS 0.011834f
C14574 DVSS.n3281 VSS 0.014662f
C14575 DVSS.n3282 VSS 0.023309f
C14576 DVSS.n3283 VSS 0.011834f
C14577 DVSS.n3284 VSS 0.010334f
C14578 DVSS.n3285 VSS 0.042011f
C14579 DVSS.n3286 VSS 0.042011f
C14580 DVSS.n3287 VSS 0.084022f
C14581 DVSS.n3288 VSS 0.084022f
C14582 DVSS.n3289 VSS 0.042011f
C14583 DVSS.n3290 VSS 0.042011f
C14584 DVSS.n3291 VSS 0.010334f
C14585 DVSS.n3292 VSS 0.011834f
C14586 DVSS.n3293 VSS 0.020865f
C14587 DVSS.n3294 VSS 0.019433f
C14588 DVSS.n3295 VSS 0.014098f
C14589 DVSS.n3296 VSS 0.011834f
C14590 DVSS.n3297 VSS 0.010334f
C14591 DVSS.n3298 VSS 0.042011f
C14592 DVSS.n3299 VSS 0.042011f
C14593 DVSS.n3300 VSS 0.084022f
C14594 DVSS.n3301 VSS 0.084022f
C14595 DVSS.n3302 VSS 0.042011f
C14596 DVSS.n3303 VSS 0.042011f
C14597 DVSS.n3304 VSS 0.010334f
C14598 DVSS.n3305 VSS 0.011834f
C14599 DVSS.n3306 VSS 0.023309f
C14600 DVSS.n3307 VSS 0.016636f
C14601 DVSS.n3308 VSS 0.016448f
C14602 DVSS.n3309 VSS 0.010501f
C14603 DVSS.n3310 VSS 0.010334f
C14604 DVSS.n3311 VSS 0.042011f
C14605 DVSS.n3312 VSS 0.042011f
C14606 DVSS.n3313 VSS 0.084022f
C14607 DVSS.n3314 VSS 0.084022f
C14608 DVSS.n3315 VSS 0.042011f
C14609 DVSS.n3316 VSS 0.042011f
C14610 DVSS.n3317 VSS 0.010334f
C14611 DVSS.n3318 VSS 0.011834f
C14612 DVSS.n3319 VSS 0.023309f
C14613 DVSS.n3320 VSS 0.023309f
C14614 DVSS.n3321 VSS 0.011834f
C14615 DVSS.n3322 VSS 0.010334f
C14616 DVSS.n3323 VSS 0.042011f
C14617 DVSS.n3324 VSS 0.042011f
C14618 DVSS.n3325 VSS 0.084022f
C14619 DVSS.n3326 VSS 0.084022f
C14620 DVSS.n3327 VSS 0.042011f
C14621 DVSS.n3328 VSS 0.042011f
C14622 DVSS.n3329 VSS 0.010334f
C14623 DVSS.n3330 VSS 0.011501f
C14624 DVSS.n3331 VSS 0.010667f
C14625 DVSS.n3332 VSS 0.023309f
C14626 DVSS.n3333 VSS 0.023309f
C14627 DVSS.n3334 VSS 0.011834f
C14628 DVSS.n3335 VSS 0.010334f
C14629 DVSS.n3336 VSS 0.042011f
C14630 DVSS.n3337 VSS 0.042011f
C14631 DVSS.n3338 VSS 0.084022f
C14632 DVSS.n3339 VSS 0.084022f
C14633 DVSS.n3340 VSS 0.042011f
C14634 DVSS.n3341 VSS 0.042011f
C14635 DVSS.n3342 VSS 0.010334f
C14636 DVSS.n3343 VSS 0.011834f
C14637 DVSS.n3344 VSS 0.016448f
C14638 DVSS.t50 VSS 0.061846f
C14639 DVSS.n3345 VSS 0.021475f
C14640 DVSS.n3346 VSS 0.012406f
C14641 DVSS.n3347 VSS 0.011834f
C14642 DVSS.n3348 VSS 0.010334f
C14643 DVSS.n3349 VSS 0.042011f
C14644 DVSS.n3350 VSS 0.042011f
C14645 DVSS.n3351 VSS 0.084022f
C14646 DVSS.n3352 VSS 0.084022f
C14647 DVSS.n3353 VSS 0.042011f
C14648 DVSS.n3354 VSS 0.042011f
C14649 DVSS.n3355 VSS 0.010334f
C14650 DVSS.n3356 VSS 0.011834f
C14651 DVSS.n3357 VSS 0.023309f
C14652 DVSS.n3358 VSS 0.023121f
C14653 DVSS.n3359 VSS 0.011834f
C14654 DVSS.n3360 VSS 0.010334f
C14655 DVSS.n3361 VSS 0.042011f
C14656 DVSS.n3362 VSS 0.042011f
C14657 DVSS.n3363 VSS 0.084022f
C14658 DVSS.n3364 VSS 0.084022f
C14659 DVSS.n3365 VSS 0.042011f
C14660 DVSS.n3366 VSS 0.042011f
C14661 DVSS.n3367 VSS 0.010334f
C14662 DVSS.n3368 VSS 0.011834f
C14663 DVSS.n3369 VSS 0.023309f
C14664 DVSS.n3370 VSS 0.023309f
C14665 DVSS.n3371 VSS 0.011834f
C14666 DVSS.n3372 VSS 0.010334f
C14667 DVSS.n3373 VSS 0.042011f
C14668 DVSS.n3374 VSS 0.042011f
C14669 DVSS.n3375 VSS 0.084022f
C14670 DVSS.n3376 VSS 0.084022f
C14671 DVSS.n3377 VSS 0.042011f
C14672 DVSS.n3378 VSS 0.042011f
C14673 DVSS.n3379 VSS 0.010334f
C14674 DVSS.n3380 VSS 0.011834f
C14675 DVSS.n3381 VSS 0.022933f
C14676 DVSS.n3382 VSS 0.023309f
C14677 DVSS.n3383 VSS 0.011834f
C14678 DVSS.n3384 VSS 0.010334f
C14679 DVSS.n3385 VSS 0.042011f
C14680 DVSS.n3386 VSS 0.042011f
C14681 DVSS.n3387 VSS 0.084022f
C14682 DVSS.n3388 VSS 0.084022f
C14683 DVSS.n3389 VSS 0.042011f
C14684 DVSS.n3390 VSS 0.042011f
C14685 DVSS.n3391 VSS 0.010334f
C14686 DVSS.n3392 VSS 0.011834f
C14687 DVSS.n3393 VSS 0.023309f
C14688 DVSS.n3394 VSS 0.012594f
C14689 DVSS.n3395 VSS 0.011001f
C14690 DVSS.n3396 VSS 0.011167f
C14691 DVSS.n3397 VSS 0.020207f
C14692 DVSS.n3398 VSS 0.023309f
C14693 DVSS.n3399 VSS 0.011834f
C14694 DVSS.n3400 VSS 0.010334f
C14695 DVSS.n3401 VSS 0.042011f
C14696 DVSS.n3402 VSS 0.042011f
C14697 DVSS.n3403 VSS 0.084022f
C14698 DVSS.n3404 VSS 0.084022f
C14699 DVSS.n3405 VSS 0.042011f
C14700 DVSS.n3406 VSS 0.042011f
C14701 DVSS.n3407 VSS 0.010334f
C14702 DVSS.n3408 VSS 0.011834f
C14703 DVSS.n3409 VSS 0.014944f
C14704 DVSS.n3410 VSS 0.013158f
C14705 DVSS.n3411 VSS 0.011834f
C14706 DVSS.n3412 VSS 0.010334f
C14707 DVSS.n3413 VSS 0.042011f
C14708 DVSS.n3414 VSS 0.042011f
C14709 DVSS.n3415 VSS 0.084022f
C14710 DVSS.n3416 VSS 0.084022f
C14711 DVSS.n3417 VSS 0.042011f
C14712 DVSS.n3418 VSS 0.042011f
C14713 DVSS.n3419 VSS 0.010334f
C14714 DVSS.n3420 VSS 0.011834f
C14715 DVSS.n3421 VSS 0.023309f
C14716 DVSS.n3422 VSS 0.023309f
C14717 DVSS.n3423 VSS 0.011834f
C14718 DVSS.n3424 VSS 0.010334f
C14719 DVSS.n3425 VSS 0.042011f
C14720 DVSS.n3426 VSS 0.042011f
C14721 DVSS.n3427 VSS 0.084022f
C14722 DVSS.n3428 VSS 0.084022f
C14723 DVSS.n3429 VSS 0.042011f
C14724 DVSS.n3430 VSS 0.042011f
C14725 DVSS.n3431 VSS 0.010334f
C14726 DVSS.n3432 VSS 0.011834f
C14727 DVSS.n3433 VSS 0.023309f
C14728 DVSS.n3434 VSS 0.023309f
C14729 DVSS.n3435 VSS 0.011834f
C14730 DVSS.n3436 VSS 0.010334f
C14731 DVSS.n3437 VSS 0.042011f
C14732 DVSS.n3438 VSS 0.042011f
C14733 DVSS.n3439 VSS 0.084022f
C14734 DVSS.n3440 VSS 0.084022f
C14735 DVSS.n3441 VSS 0.042011f
C14736 DVSS.n3442 VSS 0.042011f
C14737 DVSS.n3443 VSS 0.010334f
C14738 DVSS.n3444 VSS 0.011834f
C14739 DVSS.n3445 VSS 0.020677f
C14740 DVSS.n3446 VSS 0.023309f
C14741 DVSS.n3447 VSS 0.011834f
C14742 DVSS.n3448 VSS 0.010334f
C14743 DVSS.n3449 VSS 0.042011f
C14744 DVSS.n3450 VSS 0.042011f
C14745 DVSS.n3451 VSS 0.084022f
C14746 DVSS.n3452 VSS 0.084022f
C14747 DVSS.n3453 VSS 0.042011f
C14748 DVSS.n3454 VSS 0.042011f
C14749 DVSS.n3455 VSS 0.010334f
C14750 DVSS.n3456 VSS 0.011834f
C14751 DVSS.n3457 VSS 0.023309f
C14752 DVSS.n3458 VSS 0.01485f
C14753 DVSS.n3459 VSS 0.010501f
C14754 DVSS.n3460 VSS 0.011667f
C14755 DVSS.n3461 VSS 0.020113f
C14756 DVSS.n3462 VSS 0.023309f
C14757 DVSS.n3463 VSS 0.011834f
C14758 DVSS.n3464 VSS 0.010334f
C14759 DVSS.n3465 VSS 0.042011f
C14760 DVSS.n3466 VSS 0.042011f
C14761 DVSS.n3467 VSS 0.084022f
C14762 DVSS.n3468 VSS 0.084022f
C14763 DVSS.n3469 VSS 0.042011f
C14764 DVSS.n3470 VSS 0.042011f
C14765 DVSS.n3471 VSS 0.010334f
C14766 DVSS.n3472 VSS 0.011834f
C14767 DVSS.n3473 VSS 0.012688f
C14768 DVSS.n3474 VSS 0.015414f
C14769 DVSS.n3475 VSS 0.011834f
C14770 DVSS.n3476 VSS 0.010334f
C14771 DVSS.n3477 VSS 0.042011f
C14772 DVSS.n3478 VSS 0.042011f
C14773 DVSS.n3479 VSS 0.084022f
C14774 DVSS.n3480 VSS 0.084022f
C14775 DVSS.n3481 VSS 0.042011f
C14776 DVSS.n3482 VSS 0.042011f
C14777 DVSS.n3483 VSS 0.010334f
C14778 DVSS.n3484 VSS 0.011834f
C14779 DVSS.n3485 VSS 0.023309f
C14780 DVSS.n3486 VSS 0.023309f
C14781 DVSS.n3487 VSS 0.011834f
C14782 DVSS.n3488 VSS 0.010334f
C14783 DVSS.n3489 VSS 0.042011f
C14784 DVSS.n3490 VSS 0.042011f
C14785 DVSS.n3491 VSS 0.084022f
C14786 DVSS.n3492 VSS 0.084022f
C14787 DVSS.n3493 VSS 0.042011f
C14788 DVSS.n3494 VSS 0.042011f
C14789 DVSS.n3495 VSS 0.010334f
C14790 DVSS.n3496 VSS 0.011834f
C14791 DVSS.n3497 VSS 0.023309f
C14792 DVSS.n3498 VSS 0.023309f
C14793 DVSS.n3499 VSS 0.023309f
C14794 DVSS.n3500 VSS 0.010501f
C14795 DVSS.n3501 VSS 0.010334f
C14796 DVSS.n3502 VSS 0.042011f
C14797 DVSS.n3503 VSS 0.010334f
C14798 DVSS.n3504 VSS 0.019808f
C14799 DVSS.n3505 VSS 0.011749f
C14800 DVSS.n3506 VSS 0.163721f
C14801 DVSS.n3507 VSS 0.098089f
C14802 DVSS.n3508 VSS 0.60418f
C14803 DVSS.n3509 VSS 0.925863f
C14804 DVSS.n3510 VSS 1.97433f
C14805 DVSS.n3511 VSS 1.83056f
C14806 DVSS.n3512 VSS 0.757008f
C14807 DVSS.n3513 VSS 0.474957f
C14808 DVSS.n3514 VSS 0.092043f
C14809 DVSS.n3515 VSS 0.092043f
C14810 DVSS.n3516 VSS 0.090747f
C14811 DVSS.n3517 VSS 0.092043f
C14812 DVSS.n3518 VSS 0.092043f
C14813 DVSS.n3519 VSS 0.343557f
C14814 DVSS.n3520 VSS 0.175694f
C14815 DVSS.n3521 VSS 0.198754f
C14816 DVSS.n3522 VSS 0.673063f
C14817 DVSS.n3523 VSS 0.092043f
C14818 DVSS.n3524 VSS 0.092043f
C14819 DVSS.n3525 VSS 0.090747f
C14820 DVSS.n3526 VSS 0.092043f
C14821 DVSS.n3527 VSS 0.017825f
C14822 DVSS.n3528 VSS 0.139132f
C14823 DVSS.n3534 VSS 0.054772f
C14824 DVSS.n3535 VSS 0.026298f
C14825 DVSS.n3536 VSS 0.026298f
C14826 DVSS.n3537 VSS 0.026298f
C14827 DVSS.n3538 VSS 0.026298f
C14828 DVSS.n3539 VSS 0.092043f
C14829 DVSS.n3540 VSS 0.092043f
C14830 DVSS.n3541 VSS 0.092043f
C14831 DVSS.n3542 VSS 0.092043f
C14832 DVSS.n3543 VSS 0.092043f
C14833 DVSS.n3544 VSS 0.092043f
C14834 DVSS.n3545 VSS 0.092043f
C14835 DVSS.n3546 VSS 0.092043f
C14836 DVSS.n3547 VSS 0.092043f
C14837 DVSS.n3548 VSS 0.092043f
C14838 DVSS.n3549 VSS 0.092043f
C14839 DVSS.n3550 VSS 0.092043f
C14840 DVSS.n3551 VSS 0.092043f
C14841 DVSS.n3552 VSS 0.092043f
C14842 DVSS.n3553 VSS 0.092043f
C14843 DVSS.n3554 VSS 0.092043f
C14844 DVSS.n3555 VSS 0.092043f
C14845 DVSS.n3556 VSS 0.092043f
C14846 DVSS.n3557 VSS 0.092043f
C14847 DVSS.n3558 VSS 0.092043f
C14848 DVSS.n3559 VSS 0.092043f
C14849 DVSS.n3560 VSS 0.092043f
C14850 DVSS.n3561 VSS 0.092043f
C14851 DVSS.n3562 VSS 0.092043f
C14852 DVSS.n3563 VSS 0.092043f
C14853 DVSS.n3564 VSS 0.092043f
C14854 DVSS.n3565 VSS 0.092043f
C14855 DVSS.n3566 VSS 0.092043f
C14856 DVSS.n3567 VSS 0.092043f
C14857 DVSS.n3568 VSS 0.092043f
C14858 DVSS.n3569 VSS 0.092043f
C14859 DVSS.n3570 VSS 0.092043f
C14860 DVSS.n3571 VSS 0.092043f
C14861 DVSS.n3572 VSS 0.092043f
C14862 DVSS.n3573 VSS 0.092043f
C14863 DVSS.n3574 VSS 0.092043f
C14864 DVSS.n3575 VSS 0.092043f
C14865 DVSS.n3576 VSS 0.092043f
C14866 DVSS.n3577 VSS 0.092043f
C14867 DVSS.n3578 VSS 0.092043f
C14868 DVSS.n3579 VSS 0.092043f
C14869 DVSS.n3580 VSS 0.092043f
C14870 DVSS.n3581 VSS 0.092043f
C14871 DVSS.n3582 VSS 0.092043f
C14872 DVSS.n3583 VSS 0.092043f
C14873 DVSS.n3584 VSS 0.092043f
C14874 DVSS.n3585 VSS 0.092043f
C14875 DVSS.n3586 VSS 0.092043f
C14876 DVSS.n3587 VSS 0.092043f
C14877 DVSS.n3588 VSS 0.092043f
C14878 DVSS.n3589 VSS 0.092043f
C14879 DVSS.n3590 VSS 0.092043f
C14880 DVSS.n3591 VSS 0.092043f
C14881 DVSS.n3592 VSS 0.092043f
C14882 DVSS.n3593 VSS 0.092043f
C14883 DVSS.n3594 VSS 0.092043f
C14884 DVSS.n3595 VSS 0.092043f
C14885 DVSS.n3596 VSS 0.092043f
C14886 DVSS.n3597 VSS 0.092043f
C14887 DVSS.n3598 VSS 0.092043f
C14888 DVSS.n3599 VSS 0.092043f
C14889 DVSS.n3600 VSS 0.092043f
C14890 DVSS.n3601 VSS 0.092043f
C14891 DVSS.n3602 VSS 0.092043f
C14892 DVSS.n3603 VSS 0.092043f
C14893 DVSS.n3604 VSS 0.092043f
C14894 DVSS.n3605 VSS 0.092043f
C14895 DVSS.n3606 VSS 0.092043f
C14896 DVSS.n3607 VSS 0.092043f
C14897 DVSS.n3608 VSS 0.092043f
C14898 DVSS.n3609 VSS 0.092043f
C14899 DVSS.n3610 VSS 0.092043f
C14900 DVSS.n3611 VSS 0.092043f
C14901 DVSS.n3612 VSS 0.092043f
C14902 DVSS.n3613 VSS 0.092043f
C14903 DVSS.n3614 VSS 0.092043f
C14904 DVSS.n3615 VSS 0.092043f
C14905 DVSS.n3616 VSS 0.092043f
C14906 DVSS.n3617 VSS 0.092043f
C14907 DVSS.n3618 VSS 0.092043f
C14908 DVSS.n3619 VSS 0.092043f
C14909 DVSS.n3620 VSS 0.092043f
C14910 DVSS.n3621 VSS 0.092043f
C14911 DVSS.n3622 VSS 0.092043f
C14912 DVSS.n3623 VSS 0.092043f
C14913 DVSS.n3624 VSS 0.092043f
C14914 DVSS.n3625 VSS 0.092043f
C14915 DVSS.n3626 VSS 0.092043f
C14916 DVSS.n3627 VSS 0.092043f
C14917 DVSS.n3628 VSS 0.092043f
C14918 DVSS.n3629 VSS 0.092043f
C14919 DVSS.n3630 VSS 0.092043f
C14920 DVSS.n3631 VSS 0.092043f
C14921 DVSS.n3632 VSS 0.092043f
C14922 DVSS.n3633 VSS 0.092043f
C14923 DVSS.n3634 VSS 0.092043f
C14924 DVSS.n3635 VSS 0.092043f
C14925 DVSS.n3636 VSS 0.092043f
C14926 DVSS.n3637 VSS 0.092043f
C14927 DVSS.n3638 VSS 0.092043f
C14928 DVSS.n3639 VSS 0.092043f
C14929 DVSS.n3640 VSS 0.092043f
C14930 DVSS.n3641 VSS 0.092043f
C14931 DVSS.n3642 VSS 0.092043f
C14932 DVSS.n3643 VSS 0.092043f
C14933 DVSS.n3644 VSS 0.092043f
C14934 DVSS.n3645 VSS 0.092043f
C14935 DVSS.n3646 VSS 0.092043f
C14936 DVSS.n3647 VSS 0.092043f
C14937 DVSS.n3648 VSS 0.092043f
C14938 DVSS.n3649 VSS 0.092043f
C14939 DVSS.n3650 VSS 0.092043f
C14940 DVSS.n3651 VSS 0.092043f
C14941 DVSS.n3652 VSS 0.092043f
C14942 DVSS.n3653 VSS 0.092043f
C14943 DVSS.n3654 VSS 0.092043f
C14944 DVSS.n3655 VSS 0.092043f
C14945 DVSS.n3656 VSS 0.092043f
C14946 DVSS.n3657 VSS 0.092043f
C14947 DVSS.n3658 VSS 0.092043f
C14948 DVSS.n3659 VSS 0.092043f
C14949 DVSS.n3660 VSS 0.092043f
C14950 DVSS.n3661 VSS 0.092043f
C14951 DVSS.n3662 VSS 0.092043f
C14952 DVSS.n3663 VSS 0.092043f
C14953 DVSS.n3664 VSS 0.092043f
C14954 DVSS.n3665 VSS 0.092043f
C14955 DVSS.n3666 VSS 0.092043f
C14956 DVSS.n3667 VSS 0.092043f
C14957 DVSS.n3668 VSS 0.092043f
C14958 DVSS.n3669 VSS 0.092043f
C14959 DVSS.n3670 VSS 0.092043f
C14960 DVSS.n3671 VSS 0.092043f
C14961 DVSS.n3672 VSS 0.092043f
C14962 DVSS.n3673 VSS 0.092043f
C14963 DVSS.n3674 VSS 0.092043f
C14964 DVSS.n3675 VSS 0.092043f
C14965 DVSS.n3676 VSS 0.092043f
C14966 DVSS.n3677 VSS 0.092043f
C14967 DVSS.n3678 VSS 0.092043f
C14968 DVSS.n3679 VSS 0.092043f
C14969 DVSS.n3680 VSS 0.092043f
C14970 DVSS.n3681 VSS 0.092043f
C14971 DVSS.n3682 VSS 0.092043f
C14972 DVSS.n3683 VSS 0.092043f
C14973 DVSS.n3684 VSS 0.092043f
C14974 DVSS.n3685 VSS 0.092043f
C14975 DVSS.n3686 VSS 0.092043f
C14976 DVSS.n3687 VSS 0.092043f
C14977 DVSS.n3688 VSS 0.092043f
C14978 DVSS.n3689 VSS 0.092043f
C14979 DVSS.n3690 VSS 0.092043f
C14980 DVSS.n3691 VSS 0.092043f
C14981 DVSS.n3692 VSS 0.092043f
C14982 DVSS.n3693 VSS 0.092043f
C14983 DVSS.n3694 VSS 0.092043f
C14984 DVSS.n3695 VSS 0.092043f
C14985 DVSS.n3696 VSS 0.092043f
C14986 DVSS.n3697 VSS 0.092043f
C14987 DVSS.n3698 VSS 0.092043f
C14988 DVSS.n3699 VSS 0.092043f
C14989 DVSS.n3700 VSS 0.092043f
C14990 DVSS.n3701 VSS 0.092043f
C14991 DVSS.n3702 VSS 0.092043f
C14992 DVSS.n3703 VSS 0.092043f
C14993 DVSS.n3704 VSS 0.092043f
C14994 DVSS.n3705 VSS 0.092043f
C14995 DVSS.n3706 VSS 0.092043f
C14996 DVSS.n3707 VSS 0.092043f
C14997 DVSS.n3708 VSS 0.092043f
C14998 DVSS.n3709 VSS 0.092043f
C14999 DVSS.n3710 VSS 0.092043f
C15000 DVSS.n3711 VSS 0.092043f
C15001 DVSS.n3712 VSS 0.092043f
C15002 DVSS.n3713 VSS 0.092043f
C15003 DVSS.n3714 VSS 0.092043f
C15004 DVSS.n3715 VSS 0.092043f
C15005 DVSS.n3716 VSS 0.092043f
C15006 DVSS.n3717 VSS 0.092043f
C15007 DVSS.n3718 VSS 0.092043f
C15008 DVSS.n3719 VSS 0.092043f
C15009 DVSS.n3720 VSS 0.092043f
C15010 DVSS.n3721 VSS 0.092043f
C15011 DVSS.n3722 VSS 0.092043f
C15012 DVSS.n3723 VSS 0.092043f
C15013 DVSS.n3724 VSS 0.092043f
C15014 DVSS.n3725 VSS 0.092043f
C15015 DVSS.n3726 VSS 0.092043f
C15016 DVSS.n3727 VSS 0.092043f
C15017 DVSS.n3728 VSS 0.092043f
C15018 DVSS.n3729 VSS 0.092043f
C15019 DVSS.n3730 VSS 0.092043f
C15020 DVSS.n3731 VSS 0.092043f
C15021 DVSS.n3732 VSS 0.092043f
C15022 DVSS.n3733 VSS 0.092043f
C15023 DVSS.n3734 VSS 0.092043f
C15024 DVSS.n3735 VSS 0.092043f
C15025 DVSS.n3736 VSS 0.092043f
C15026 DVSS.n3737 VSS 0.092043f
C15027 DVSS.n3738 VSS 0.092043f
C15028 DVSS.n3739 VSS 0.092043f
C15029 DVSS.n3740 VSS 0.092043f
C15030 DVSS.n3741 VSS 0.092043f
C15031 DVSS.n3742 VSS 0.092043f
C15032 DVSS.n3743 VSS 0.092043f
C15033 DVSS.n3744 VSS 0.092043f
C15034 DVSS.n3745 VSS 0.055096f
C15035 DVSS.n3746 VSS 0.047318f
C15036 DVSS.n3747 VSS 0.092043f
C15037 DVSS.n3748 VSS 0.082968f
C15038 DVSS.n3749 VSS 0.046022f
C15039 DVSS.n3750 VSS 0.026298f
C15040 DVSS.n3751 VSS 0.026298f
C15041 DVSS.n3752 VSS 0.026298f
C15042 DVSS.n3756 VSS 0.036947f
C15043 DVSS.n3758 VSS 0.026298f
C15044 DVSS.n3759 VSS 0.046022f
C15045 DVSS.n3760 VSS 1.22823f
C15046 DVSS.n3761 VSS 0.046022f
C15047 DVSS.n3762 VSS 0.083292f
C15048 DVSS.n3763 VSS 0.092043f
C15049 DVSS.n3764 VSS 0.092043f
C15050 DVSS.n3765 VSS 0.343557f
C15051 DVSS.n3766 VSS 0.175694f
C15052 DVSS.n3767 VSS 0.19875f
C15053 DVSS.n3768 VSS 0.816868f
C15054 DVSS.n3769 VSS 1.03455f
C15055 DVSS.n3770 VSS 2.32106f
C15056 DVSS.n3771 VSS 1.26425f
C15057 DVSS.n3772 VSS 1.71338f
C15058 DVSS.t89 VSS 0.182334f
C15059 DVSS.t87 VSS 0.182334f
C15060 DVSS.t181 VSS 0.228665f
C15061 DVSS.n3773 VSS 0.016916f
C15062 DVSS.n3774 VSS 0.162256f
C15063 DVSS.t183 VSS 0.222687f
C15064 DVSS.n3775 VSS 0.284184f
C15065 DVSS.t95 VSS 0.22194f
C15066 DVSS.t85 VSS 0.183082f
C15067 DVSS.n3776 VSS 0.256314f
C15068 DVSS.n3777 VSS 0.346634f
C15069 DVSS.t76 VSS 0.255567f
C15070 DVSS.n3778 VSS 0.430428f
C15071 DVSS.n3779 VSS 0.033005f
C15072 DVSS.n3780 VSS 0.012655f
C15073 DVSS.n3781 VSS 0.022126f
C15074 DVSS.n3782 VSS 0.053985f
C15075 DVSS.n3783 VSS 0.158917f
C15076 DVSS.n3784 VSS 0.105432f
C15077 DVSS.n3785 VSS 0.146129f
C15078 DVSS.n3786 VSS 0.030315f
C15079 DVSS.n3787 VSS 0.058762f
C15080 DVSS.n3788 VSS 0.013968f
C15081 DVSS.n3789 VSS 0.03233f
C15082 DVSS.n3790 VSS 0.023111f
C15083 DVSS.n3791 VSS 0.274996f
C15084 DVSS.n3792 VSS 0.167282f
C15085 DVSS.t173 VSS 0.004574f
C15086 DVSS.t178 VSS 0.004574f
C15087 DVSS.n3793 VSS 0.082418f
C15088 DVSS.n3794 VSS 0.098351f
C15089 DVSS.n3795 VSS 0.015019f
C15090 DVSS.n3796 VSS 0.021357f
C15091 DVSS.n3797 VSS -0.009133f
C15092 DVSS.n3798 VSS 0.155824f
C15093 DVSS.t19 VSS 0.146465f
C15094 DVSS.n3799 VSS 0.279456f
C15095 DVSS.n3800 VSS 1.31875f
C15096 DVSS.n3801 VSS 1.89449f
C15097 DVSS.n3802 VSS 2.53162f
C15098 DVSS.n3806 VSS 0.043336f
C15099 DVSS.n3807 VSS 0.043336f
C15100 DVSS.n3808 VSS 0.043336f
C15101 DVSS.n3809 VSS 0.043336f
C15102 DVSS.n3810 VSS 0.043336f
C15103 DVSS.n3811 VSS 0.043336f
C15104 DVSS.n3812 VSS 0.043336f
C15105 DVSS.n3813 VSS 0.043336f
C15106 DVSS.n3814 VSS 0.043336f
C15107 DVSS.n3815 VSS 0.043336f
C15108 DVSS.n3816 VSS 0.078538f
C15109 DVSS.n3817 VSS 0.042041f
C15110 DVSS.n3819 VSS 0.854875f
C15111 DVSS.n3820 VSS 0.041407f
C15112 DVSS.n3821 VSS 0.073278f
C15113 DVSS.n3822 VSS 0.11357f
C15114 DVSS.n3823 VSS 0.223447f
C15115 DVSS.t150 VSS 0.389389f
C15116 DVSS.n3824 VSS 0.781718f
C15117 DVSS.n3825 VSS 0.953727f
C15118 DVSS.n3826 VSS 0.280656f
C15119 DVSS.n3827 VSS 0.051455f
C15120 DVSS.n3828 VSS 0.019808f
C15121 DVSS.n3829 VSS 0.042064f
C15122 DVSS.n3830 VSS 0.042011f
C15123 DVSS.n3831 VSS 0.084022f
C15124 DVSS.n3832 VSS 0.084022f
C15125 DVSS.n3833 VSS 0.084022f
C15126 DVSS.n3834 VSS 0.084022f
C15127 DVSS.n3835 VSS 0.084022f
C15128 DVSS.n3836 VSS 0.084022f
C15129 DVSS.n3837 VSS 0.084022f
C15130 DVSS.n3838 VSS 0.084022f
C15131 DVSS.n3839 VSS 0.084022f
C15132 DVSS.n3840 VSS 0.084022f
C15133 DVSS.n3841 VSS 0.084022f
C15134 DVSS.n3842 VSS 0.084022f
C15135 DVSS.n3843 VSS 0.084022f
C15136 DVSS.n3844 VSS 0.084022f
C15137 DVSS.n3845 VSS 0.084022f
C15138 DVSS.n3846 VSS 0.084022f
C15139 DVSS.n3847 VSS 0.084022f
C15140 DVSS.n3848 VSS 0.084022f
C15141 DVSS.n3849 VSS 0.084022f
C15142 DVSS.n3850 VSS 0.084022f
C15143 DVSS.n3851 VSS 0.043195f
C15144 DVSS.n3852 VSS 0.109963f
C15145 DVSS.n3853 VSS 0.405581f
C15146 DVSS.n3854 VSS 0.075738f
C15147 DVSS.n3855 VSS 0.075738f
C15148 DVSS.n3856 VSS 0.084022f
C15149 DVSS.n3857 VSS 0.084022f
C15150 DVSS.n3858 VSS 0.084022f
C15151 DVSS.n3859 VSS 0.084022f
C15152 DVSS.n3860 VSS 0.084022f
C15153 DVSS.n3861 VSS 0.084022f
C15154 DVSS.n3862 VSS 0.084022f
C15155 DVSS.n3863 VSS 0.084022f
C15156 DVSS.n3864 VSS 0.083726f
C15157 DVSS.n3865 VSS 0.11738f
C15158 DVSS.n3866 VSS 0.126498f
C15159 DVSS.n3867 VSS 0.046346f
C15160 DVSS.n3868 VSS 0.092043f
C15161 DVSS.n3869 VSS 0.092043f
C15162 DVSS.n3870 VSS 0.092043f
C15163 DVSS.n3871 VSS 0.092043f
C15164 DVSS.n3872 VSS 0.092043f
C15165 DVSS.n3873 VSS 0.092043f
C15166 DVSS.n3874 VSS 0.092043f
C15167 DVSS.n3875 VSS 0.092043f
C15168 DVSS.n3876 VSS 0.092043f
C15169 DVSS.n3877 VSS 0.092043f
C15170 DVSS.n3878 VSS 0.092043f
C15171 DVSS.n3879 VSS 0.092043f
C15172 DVSS.n3880 VSS 0.092043f
C15173 DVSS.n3881 VSS 0.092043f
C15174 DVSS.n3882 VSS 0.092043f
C15175 DVSS.n3883 VSS 0.092043f
C15176 DVSS.n3884 VSS 0.092043f
C15177 DVSS.n3885 VSS 0.092043f
C15178 DVSS.n3886 VSS 0.092043f
C15179 DVSS.n3887 VSS 0.092043f
C15180 DVSS.n3888 VSS 0.092043f
C15181 DVSS.n3889 VSS 0.092043f
C15182 DVSS.n3890 VSS 0.092043f
C15183 DVSS.n3891 VSS 0.092043f
C15184 DVSS.n3892 VSS 0.092043f
C15185 DVSS.n3893 VSS 0.092043f
C15186 DVSS.n3894 VSS 0.092043f
C15187 DVSS.n3895 VSS 0.092043f
C15188 DVSS.n3896 VSS 0.092043f
C15189 DVSS.n3897 VSS 0.092043f
C15190 DVSS.n3898 VSS 0.092043f
C15191 DVSS.n3899 VSS 0.092043f
C15192 DVSS.n3900 VSS 0.092043f
C15193 DVSS.n3901 VSS 0.092043f
C15194 DVSS.n3902 VSS 0.092043f
C15195 DVSS.n3903 VSS 0.092043f
C15196 DVSS.n3904 VSS 0.092043f
C15197 DVSS.n3905 VSS 0.092043f
C15198 DVSS.n3906 VSS 0.092043f
C15199 DVSS.n3907 VSS 0.053476f
C15200 DVSS.n3908 VSS 0.092043f
C15201 DVSS.n3909 VSS 0.092043f
C15202 DVSS.n3910 VSS 0.092043f
C15203 DVSS.n3911 VSS 0.092043f
C15204 DVSS.n3912 VSS 0.092043f
C15205 DVSS.n3913 VSS 0.06968f
C15206 DVSS.n3914 VSS 0.092043f
C15207 DVSS.n3915 VSS 0.088478f
C15208 DVSS.n3916 VSS 0.092043f
C15209 DVSS.n3917 VSS 0.092043f
C15210 DVSS.n3918 VSS 0.092043f
C15211 DVSS.n3919 VSS 0.092043f
C15212 DVSS.n3920 VSS 0.092043f
C15213 DVSS.n3921 VSS 0.092043f
C15214 DVSS.n3922 VSS 0.092043f
C15215 DVSS.n3923 VSS 0.06255f
C15216 DVSS.n3924 VSS 0.092043f
C15217 DVSS.n3925 VSS 0.092043f
C15218 DVSS.n3926 VSS 0.092043f
C15219 DVSS.n3927 VSS 0.092043f
C15220 DVSS.n3928 VSS 0.092043f
C15221 DVSS.n3929 VSS 0.058985f
C15222 DVSS.n3930 VSS 0.06048f
C15223 DVSS.n3931 VSS 0.021061f
C15224 DVSS.n3932 VSS 0.010037f
C15225 DVSS.n3933 VSS 0.011923f
C15226 DVSS.n3934 VSS 0.010037f
C15227 DVSS.n3935 VSS -0.005479f
C15228 DVSS.n3936 VSS 0.158916f
C15229 DVSS.t93 VSS 0.141982f
C15230 DVSS.t3 VSS 0.175609f
C15231 DVSS.n3937 VSS 0.132267f
C15232 DVSS.n3938 VSS 0.211185f
C15233 DVSS.n3939 VSS 0.026469f
C15234 DVSS.n3940 VSS 0.043595f
C15235 DVSS.t100 VSS 0.003611f
C15236 DVSS.t141 VSS 0.003611f
C15237 DVSS.n3941 VSS 0.007291f
C15238 DVSS.n3942 VSS 8.12e-19
C15239 DVSS.n3943 VSS 0.01033f
C15240 DVSS.n3944 VSS 0.045791f
C15241 DVSS.n3945 VSS 0.047349f
C15242 DVSS.n3946 VSS 0.075514f
C15243 DVSS.n3947 VSS 0.092043f
C15244 DVSS.n3948 VSS 0.092043f
C15245 DVSS.n3949 VSS 0.092043f
C15246 DVSS.n3950 VSS 0.092043f
C15247 DVSS.n3951 VSS 0.092043f
C15248 DVSS.n3952 VSS 0.082644f
C15249 DVSS.n3953 VSS 0.047352f
C15250 DVSS.n3954 VSS 0.04528f
C15251 DVSS.n3955 VSS 0.010322f
C15252 DVSS.n3956 VSS 0.021956f
C15253 DVSS.n3957 VSS 0.016916f
C15254 DVSS.n3958 VSS 0.062562f
C15255 DVSS.n3959 VSS 0.086534f
C15256 DVSS.n3960 VSS 0.092043f
C15257 DVSS.n3961 VSS 0.092043f
C15258 DVSS.n3962 VSS 0.092043f
C15259 DVSS.n3963 VSS 0.092043f
C15260 DVSS.n3964 VSS 0.092043f
C15261 DVSS.n3965 VSS 0.092043f
C15262 DVSS.n3966 VSS 0.092043f
C15263 DVSS.n3967 VSS 0.092043f
C15264 DVSS.n3968 VSS 0.092043f
C15265 DVSS.n3969 VSS 0.092043f
C15266 DVSS.n3970 VSS 0.092043f
C15267 DVSS.n3971 VSS 0.092043f
C15268 DVSS.n3972 VSS 0.092043f
C15269 DVSS.n3973 VSS 0.092043f
C15270 DVSS.n3974 VSS 0.092043f
C15271 DVSS.n3975 VSS 0.092043f
C15272 DVSS.n3976 VSS 0.092043f
C15273 DVSS.n3977 VSS 0.092043f
C15274 DVSS.n3978 VSS 0.092043f
C15275 DVSS.n3979 VSS 0.092043f
C15276 DVSS.n3980 VSS 0.092043f
C15277 DVSS.n3981 VSS 0.092043f
C15278 DVSS.n3982 VSS 0.058985f
C15279 DVSS.n3985 VSS 0.026298f
C15280 DVSS.n3988 VSS 0.026298f
C15281 DVSS.n3991 VSS 0.026298f
C15282 DVSS.n3993 VSS 0.025742f
C15283 DVSS.n3994 VSS 0.046022f
C15284 DVSS.n3995 VSS 0.046022f
C15285 DVSS.n3996 VSS 0.092043f
C15286 DVSS.n3997 VSS 0.092043f
C15287 DVSS.n3998 VSS 0.092043f
C15288 DVSS.n3999 VSS 0.092043f
C15289 DVSS.n4000 VSS 0.092043f
C15290 DVSS.n4001 VSS 0.079079f
C15291 DVSS.n4002 VSS 0.092043f
C15292 DVSS.n4003 VSS 0.092043f
C15293 DVSS.n4004 VSS 0.092043f
C15294 DVSS.n4005 VSS 0.092043f
C15295 DVSS.n4006 VSS 0.092043f
C15296 DVSS.n4007 VSS 0.092043f
C15297 DVSS.n4008 VSS 0.092043f
C15298 DVSS.n4009 VSS 0.06093f
C15299 DVSS.t170 VSS 0.009309f
C15300 DVSS.n4010 VSS 0.003795f
C15301 DVSS.n4011 VSS 0.021061f
C15302 DVSS.n4012 VSS 0.06048f
C15303 DVSS.n4013 VSS 0.072921f
C15304 DVSS.n4014 VSS 0.092043f
C15305 DVSS.n4015 VSS 0.092043f
C15306 DVSS.n4016 VSS 0.092043f
C15307 DVSS.n4017 VSS 0.092043f
C15308 DVSS.n4018 VSS 0.092043f
C15309 DVSS.n4019 VSS 0.092043f
C15310 DVSS.n4020 VSS 0.052828f
C15311 DVSS.n4021 VSS 0.092043f
C15312 DVSS.n4022 VSS 0.092043f
C15313 DVSS.n4023 VSS 0.092043f
C15314 DVSS.n4024 VSS 0.092043f
C15315 DVSS.n4025 VSS 0.092043f
C15316 DVSS.n4026 VSS 0.092043f
C15317 DVSS.n4027 VSS 0.092043f
C15318 DVSS.n4028 VSS 0.058985f
C15319 DVSS.n4029 VSS 0.063581f
C15320 DVSS.n4030 VSS 0.058985f
C15321 DVSS.n4031 VSS 0.06048f
C15322 DVSS.n4032 VSS 0.052828f
C15323 DVSS.n4033 VSS 0.092043f
C15324 DVSS.n4034 VSS 0.092043f
C15325 DVSS.n4035 VSS 0.092043f
C15326 DVSS.n4036 VSS 0.092043f
C15327 DVSS.n4037 VSS 0.092043f
C15328 DVSS.n4038 VSS 0.092043f
C15329 DVSS.n4039 VSS 0.059309f
C15330 DVSS.n4040 VSS 0.06048f
C15331 DVSS.n4041 VSS 0.078755f
C15332 DVSS.n4042 VSS 0.092043f
C15333 DVSS.n4043 VSS 0.092043f
C15334 DVSS.n4044 VSS 0.092043f
C15335 DVSS.n4045 VSS 0.092043f
C15336 DVSS.n4046 VSS 0.092043f
C15337 DVSS.n4047 VSS 0.079403f
C15338 DVSS.n4048 VSS 0.06048f
C15339 DVSS.n4049 VSS 0.021061f
C15340 DVSS.n4050 VSS 0.021956f
C15341 DVSS.n4051 VSS -0.005479f
C15342 DVSS.n4052 VSS 0.010037f
C15343 DVSS.n4053 VSS 0.011923f
C15344 DVSS.n4054 VSS 0.010037f
C15345 DVSS.n4055 VSS -0.005479f
C15346 DVSS.n4056 VSS 0.158916f
C15347 DVSS.t135 VSS 0.150949f
C15348 DVSS.n4057 VSS 0.160874f
C15349 DVSS.n4058 VSS 0.014254f
C15350 DVSS.n4059 VSS 0.058027f
C15351 DVSS.n4060 VSS 0.078431f
C15352 DVSS.n4061 VSS 0.092043f
C15353 DVSS.n4062 VSS 0.092043f
C15354 DVSS.n4063 VSS 0.092043f
C15355 DVSS.n4064 VSS 0.092043f
C15356 DVSS.n4065 VSS 0.092043f
C15357 DVSS.n4066 VSS 0.092043f
C15358 DVSS.n4067 VSS 0.092043f
C15359 DVSS.n4068 VSS 0.092043f
C15360 DVSS.n4069 VSS 0.092043f
C15361 DVSS.n4070 VSS 0.092043f
C15362 DVSS.n4071 VSS 0.092043f
C15363 DVSS.n4072 VSS 0.092043f
C15364 DVSS.n4073 VSS 0.092043f
C15365 DVSS.n4074 VSS 0.092043f
C15366 DVSS.n4075 VSS 0.092043f
C15367 DVSS.n4076 VSS 0.092043f
C15368 DVSS.n4077 VSS 0.092043f
C15369 DVSS.n4078 VSS 0.092043f
C15370 DVSS.n4079 VSS 0.092043f
C15371 DVSS.n4080 VSS 0.092043f
C15372 DVSS.n4081 VSS 0.092043f
C15373 DVSS.n4082 VSS 0.092043f
C15374 DVSS.n4083 VSS 0.092043f
C15375 DVSS.n4084 VSS 0.092043f
C15376 DVSS.n4085 VSS 0.092043f
C15377 DVSS.n4086 VSS 0.092043f
C15378 DVSS.n4087 VSS 0.092043f
C15379 DVSS.n4088 VSS 0.092043f
C15380 DVSS.n4089 VSS 0.092043f
C15381 DVSS.n4090 VSS 0.06968f
C15382 DVSS.n4091 VSS 0.046022f
C15383 DVSS.n4092 VSS 0.224373f
C15384 DVSS.n4093 VSS 0.067808f
C15385 DVSS.n4094 VSS -0.029005f
C15386 DVSS.n4095 VSS 0.023111f
C15387 DVSS.n4096 VSS 1.02392f
C15388 DVSS.n4097 VSS 0.956897f
C15389 DVSS.n4098 VSS 1.27256f
C15390 DVSS.n4099 VSS 0.800055f
C15391 DVSS.n4100 VSS 0.18454f
C15392 DVSS.t54 VSS 0.037108f
C15393 DVSS.n4101 VSS 0.071349f
C15394 DVSS.n4102 VSS 0.041247f
C15395 DVSS.n4103 VSS 0.082356f
C15396 DVSS.n4104 VSS 0.423086f
C15397 DVSS.n4105 VSS 0.013184f
C15398 DVSS.n4106 VSS 0.05833f
C15399 DVSS.n4107 VSS 0.073639f
C15400 DVSS.n4108 VSS 0.058234f
C15401 DVSS.t52 VSS 0.037108f
C15402 DVSS.n4109 VSS 0.082194f
C15403 DVSS.n4110 VSS 0.01313f
C15404 DVSS.n4111 VSS 0.263841f
C15405 DVSS.n4112 VSS 0.556116f
C15406 DVSS.n4113 VSS -0.004788f
C15407 DVSS.n4114 VSS 0.016403f
C15408 DVSS.n4115 VSS 0.174237f
C15409 DVSS.n4116 VSS 0.01735f
C15410 DVSS.n4117 VSS 0.00676f
C15411 DVSS.n4118 VSS 0.197124f
C15412 DVSS.n4119 VSS 0.158225f
C15413 DVSS.n4120 VSS 0.287343f
C15414 DVSS.n4121 VSS 0.04732f
C15415 DVSS.n4122 VSS 0.033576f
C15416 DVSS.n4123 VSS 0.051726f
C15417 DVSS.n4124 VSS 0.051726f
C15418 DVSS.n4125 VSS 0.052887f
C15419 DVSS.n4126 VSS 0.097025f
C15420 DVSS.n4127 VSS 0.170167f
C15421 DVSS.n4128 VSS 0.170167f
C15422 DVSS.n4129 VSS 0.052887f
C15423 DVSS.n4130 VSS 0.051726f
C15424 DVSS.n4131 VSS 0.051726f
C15425 DVSS.n4132 VSS 0.051726f
C15426 DVSS.n4133 VSS 0.052887f
C15427 DVSS.n4134 VSS 0.167928f
C15428 DVSS.n4135 VSS 0.192192f
C15429 DVSS.n4136 VSS -0.078956f
C15430 DVSS.n4137 VSS 0.856609f
C15431 DVSS.n4138 VSS 0.217692f
C15432 DVSS.n4139 VSS 0.006899f
C15433 DVSS.n4140 VSS 0.263943f
C15434 DVSS.n4141 VSS 0.031599f
C15435 DVSS.n4142 VSS 0.012097f
C15436 DVSS.n4143 VSS 0.018401f
C15437 DVSS.n4144 VSS 0.012097f
C15438 DVSS.n4145 VSS 0.018401f
C15439 DVSS.n4146 VSS 0.018401f
C15440 DVSS.n4147 VSS 0.010649f
C15441 DVSS.n4148 VSS 0.010649f
C15442 DVSS.n4149 VSS 0.018401f
C15443 DVSS.n4150 VSS 0.012097f
C15444 DVSS.n4151 VSS 0.018401f
C15445 DVSS.n4152 VSS 0.018401f
C15446 DVSS.n4153 VSS 0.012097f
C15447 DVSS.n4154 VSS 0.009201f
C15448 DVSS.n4155 VSS 0.046022f
C15449 DVSS.n4156 VSS 0.011671f
C15450 DVSS.n4157 VSS 0.010138f
C15451 DVSS.n4158 VSS 0.025983f
C15452 DVSS.n4159 VSS -0.130991f
C15453 DVSS.n4160 VSS 0.501971f
C15454 DVSS.n4161 VSS 0.748387f
C15455 DVSS.n4162 VSS 1.24092f
C15456 DVSS.n4163 VSS 0.304048f
C15457 DVSS.n4164 VSS -0.010323f
C15458 DVSS.n4165 VSS 0.393316f
C15459 DVSS.n4166 VSS 0.092732f
C15460 DVSS.n4167 VSS 0.051726f
C15461 DVSS.n4168 VSS 0.052887f
C15462 DVSS.n4169 VSS 0.086576f
C15463 DVSS.n4170 VSS 0.29917f
C15464 DVSS.n4171 VSS 0.461959f
C15465 DVSS.n4172 VSS 0.508959f
C15466 DVSS.n4173 VSS 0.524925f
C15467 DVSS.n4174 VSS 0.393954f
C15468 DVSS.n4175 VSS 0.34247f
C15469 DVSS.n4176 VSS 0.055783f
C15470 DVSS.n4177 VSS 0.645493f
C15471 DVSS.n4178 VSS 0.082172f
C15472 DVSS.n4179 VSS 0.078841f
C15473 DVSS.n4180 VSS 0.049402f
C15474 DVSS.n4181 VSS 0.035876f
C15475 DVSS.n4182 VSS 0.009596f
C15476 DVSS.t113 VSS 0.014445f
C15477 DVSS.n4183 VSS 0.038498f
C15478 DVSS.n4184 VSS 0.002551f
C15479 DVSS.n4185 VSS 0.032017f
C15480 DVSS.n4186 VSS 0.126367f
C15481 DVSS.n4187 VSS 0.181262f
C15482 DVSS.n4188 VSS 0.197235f
C15483 DVSS.n4189 VSS 0.197235f
C15484 DVSS.n4190 VSS 0.197235f
C15485 DVSS.n4191 VSS 0.197235f
C15486 DVSS.n4192 VSS 0.197235f
C15487 DVSS.n4193 VSS 0.197235f
C15488 DVSS.n4194 VSS 0.197235f
C15489 DVSS.n4195 VSS 0.197235f
C15490 DVSS.n4196 VSS 0.197235f
C15491 DVSS.n4197 VSS 0.197235f
C15492 DVSS.n4198 VSS 0.197235f
C15493 DVSS.n4199 VSS 0.197235f
C15494 DVSS.n4200 VSS 0.197235f
C15495 DVSS.n4201 VSS 0.197235f
C15496 DVSS.n4202 VSS 0.197235f
C15497 DVSS.n4203 VSS 0.197235f
C15498 DVSS.n4204 VSS 0.197235f
C15499 DVSS.n4205 VSS 0.197235f
C15500 DVSS.n4206 VSS 0.197235f
C15501 DVSS.n4207 VSS 0.197235f
C15502 DVSS.n4208 VSS 0.197235f
C15503 DVSS.n4209 VSS 0.197235f
C15504 DVSS.n4210 VSS 0.197235f
C15505 DVSS.n4211 VSS 0.197235f
C15506 DVSS.n4212 VSS 0.197235f
C15507 DVSS.n4213 VSS 0.197235f
C15508 DVSS.n4214 VSS 0.197235f
C15509 DVSS.n4215 VSS 0.197235f
C15510 DVSS.n4216 VSS 0.197235f
C15511 DVSS.n4217 VSS 0.197235f
C15512 DVSS.n4218 VSS 0.197235f
C15513 DVSS.n4219 VSS 0.197235f
C15514 DVSS.n4220 VSS 0.197235f
C15515 DVSS.n4221 VSS 0.197235f
C15516 DVSS.n4222 VSS 0.197235f
C15517 DVSS.n4223 VSS 0.197235f
C15518 DVSS.n4224 VSS 0.197235f
C15519 DVSS.n4225 VSS 0.197235f
C15520 DVSS.n4226 VSS 0.197235f
C15521 DVSS.n4227 VSS 0.197235f
C15522 DVSS.n4228 VSS 0.197235f
C15523 DVSS.n4229 VSS 0.197235f
C15524 DVSS.n4230 VSS 0.197235f
C15525 DVSS.n4231 VSS 0.197235f
C15526 DVSS.n4232 VSS 0.197235f
C15527 DVSS.n4233 VSS 0.197235f
C15528 DVSS.n4234 VSS 0.197235f
C15529 DVSS.n4235 VSS 0.197235f
C15530 DVSS.n4236 VSS 0.197235f
C15531 DVSS.n4237 VSS 0.197235f
C15532 DVSS.n4238 VSS 0.197235f
C15533 DVSS.n4239 VSS 0.197235f
C15534 DVSS.n4240 VSS 0.197235f
C15535 DVSS.n4241 VSS 0.197235f
C15536 DVSS.n4242 VSS 0.197235f
C15537 DVSS.n4243 VSS 0.197235f
C15538 DVSS.n4244 VSS 0.197235f
C15539 DVSS.n4245 VSS 0.197235f
C15540 DVSS.n4246 VSS 0.197235f
C15541 DVSS.n4247 VSS 0.197235f
C15542 DVSS.n4248 VSS 0.197235f
C15543 DVSS.n4249 VSS 0.197235f
C15544 DVSS.n4250 VSS 0.197235f
C15545 DVSS.n4251 VSS 0.197235f
C15546 DVSS.n4252 VSS 0.197235f
C15547 DVSS.n4253 VSS 0.197235f
C15548 DVSS.n4254 VSS 0.197235f
C15549 DVSS.n4255 VSS 0.197235f
C15550 DVSS.n4256 VSS 0.197235f
C15551 DVSS.n4257 VSS 0.197235f
C15552 DVSS.n4258 VSS 0.197235f
C15553 DVSS.n4259 VSS 0.197235f
C15554 DVSS.n4260 VSS 0.197235f
C15555 DVSS.n4261 VSS 0.197235f
C15556 DVSS.n4262 VSS 0.197235f
C15557 DVSS.n4263 VSS 0.197235f
C15558 DVSS.n4264 VSS 0.197235f
C15559 DVSS.n4265 VSS 0.197235f
C15560 DVSS.n4266 VSS 0.197235f
C15561 DVSS.n4267 VSS 0.197235f
C15562 DVSS.n4268 VSS 0.197235f
C15563 DVSS.n4269 VSS 0.197235f
C15564 DVSS.n4270 VSS 0.197235f
C15565 DVSS.n4271 VSS 0.197235f
C15566 DVSS.n4272 VSS 0.197235f
C15567 DVSS.n4273 VSS 0.197235f
C15568 DVSS.n4274 VSS 0.197235f
C15569 DVSS.n4275 VSS 0.197235f
C15570 DVSS.n4276 VSS 0.197235f
C15571 DVSS.n4277 VSS 0.197235f
C15572 DVSS.n4278 VSS 0.197235f
C15573 DVSS.n4279 VSS 0.197235f
C15574 DVSS.n4280 VSS 0.197235f
C15575 DVSS.n4281 VSS 0.175012f
C15576 DVSS.n4282 VSS 0.123472f
C15577 DVSS.n4283 VSS 0.074656f
C15578 DVSS.n4284 VSS 0.019367f
C15579 DVSS.n4285 VSS 0.050526f
C15580 DVSS.n4286 VSS 0.252098f
C15581 DVSS.t46 VSS 0.387914f
C15582 DVSS.t171 VSS 0.273557f
C15583 DVSS.t81 VSS 0.206289f
C15584 DVSS.n4287 VSS 0.175293f
C15585 DVSS.n4288 VSS 0.002351f
C15586 DVSS.n4289 VSS 0.259431f
C15587 DVSS.t106 VSS 0.170413f
C15588 DVSS.n4290 VSS 0.273557f
C15589 DVSS.n4291 VSS 0.04679f
C15590 DVSS.n4292 VSS 0.021032f
C15591 DVSS.n4293 VSS 0.025192f
C15592 DVSS.n4294 VSS 0.093193f
C15593 DVSS.n4295 VSS 0.025192f
C15594 DVSS.n4296 VSS 0.021032f
C15595 DVSS.n4297 VSS 0.04679f
C15596 DVSS.n4298 VSS 0.182745f
C15597 DVSS.n4299 VSS 0.300697f
C15598 DVSS.t0 VSS 0.334099f
C15599 DVSS.t119 VSS 0.009309f
C15600 DVSS.n4300 VSS 0.009615f
C15601 DVSS.t175 VSS 0.003611f
C15602 DVSS.t159 VSS 0.003611f
C15603 DVSS.n4301 VSS 0.007291f
C15604 DVSS.n4302 VSS 0.006632f
C15605 DVSS.n4303 VSS 0.260684f
C15606 DVSS.t122 VSS 0.155838f
C15607 DVSS.n4304 VSS 0.273558f
C15608 DVSS.t124 VSS 0.241045f
C15609 DVSS.t44 VSS 0.273557f
C15610 DVSS.t202 VSS 0.273557f
C15611 DVSS.t174 VSS 0.238802f
C15612 DVSS.t190 VSS 0.273557f
C15613 DVSS.t158 VSS 0.273557f
C15614 DVSS.t160 VSS 0.139021f
C15615 DVSS.n4305 VSS 0.143915f
C15616 DVSS.t45 VSS 0.009309f
C15617 DVSS.n4306 VSS 0.009615f
C15618 DVSS.n4307 VSS 0.012141f
C15619 DVSS.n4308 VSS -0.004609f
C15620 DVSS.n4309 VSS 0.027535f
C15621 DVSS.n4310 VSS 0.255903f
C15622 DVSS.t5 VSS 0.303828f
C15623 DVSS.n4311 VSS 0.293665f
C15624 DVSS.n4312 VSS -0.047747f
C15625 DVSS.n4313 VSS 0.02551f
C15626 DVSS.n4314 VSS 0.018694f
C15627 DVSS.n4315 VSS 0.081583f
C15628 DVSS.n4316 VSS 0.02826f
C15629 DVSS.n4317 VSS 0.113302f
C15630 DVSS.n4318 VSS 0.439486f
C15631 DVSS.n4319 VSS 2.20853f
C15632 DVSS.n4320 VSS 0.710505f
C15633 DVSS.n4321 VSS 2.8251f
C15634 DVSS.n4322 VSS 1.42228f
C15635 DVSS.n4323 VSS 2.359f
C15636 DVSS.n4324 VSS 0.068967f
C15637 DVSS.n4325 VSS 0.259592f
C15638 DVSS.n4326 VSS 0.023539f
C15639 DVSS.n4327 VSS 0.026956f
C15640 DVSS.n4328 VSS 0.046022f
C15641 DVSS.n4329 VSS 0.046022f
C15642 DVSS.n4330 VSS 0.092043f
C15643 DVSS.n4331 VSS 0.092043f
C15644 DVSS.n4332 VSS 0.092043f
C15645 DVSS.n4333 VSS 0.092043f
C15646 DVSS.n4334 VSS 0.046022f
C15647 DVSS.n4335 VSS 0.042497f
C15648 DVSS.n4336 VSS 0.061578f
C15649 DVSS.n4337 VSS 0.046022f
C15650 DVSS.n4338 VSS 0.092043f
C15651 DVSS.n4339 VSS 0.092043f
C15652 DVSS.n4340 VSS 0.092043f
C15653 DVSS.n4341 VSS 0.046022f
C15654 DVSS.n4342 VSS 0.092043f
C15655 DVSS.n4343 VSS 0.986707f
C15656 DVSS.n4345 VSS 0.026298f
C15657 DVSS.n4347 VSS 0.026298f
C15658 DVSS.n4349 VSS 0.026298f
C15659 DVSS.n4351 VSS 0.026298f
C15660 DVSS.n4353 VSS 0.026298f
C15661 DVSS.n4355 VSS 0.026298f
C15662 DVSS.n4357 VSS 0.016853f
C15663 DVSS.n4359 VSS 0.020187f
C15664 DVSS.n4360 VSS 1.49051f
C15665 DVSS.n4361 VSS 0.038351f
C15666 DVSS.n4364 VSS 0.022965f
C15667 DVSS.n4366 VSS 0.022965f
C15668 DVSS.n4367 VSS 0.066495f
C15669 DVSS.n4368 VSS 0.028706f
C15670 DVSS.n4369 VSS 0.086134f
C15671 DVSS.n4370 VSS 0.013149f
C15672 DVSS.n4371 VSS 0.011482f
C15673 DVSS.n4372 VSS 0.046022f
C15674 DVSS.n4373 VSS 0.026298f
C15675 DVSS.n4375 VSS 0.024446f
C15676 DVSS.n4376 VSS 0.046022f
C15677 DVSS.n4377 VSS 0.046022f
C15678 DVSS.n4378 VSS 0.273386f
C15679 DVSS.n4379 VSS 1.47934f
C15680 DVSS.n4380 VSS 1.09008f
C15681 DVSS.n4381 VSS 0.092043f
C15682 DVSS.n4382 VSS 0.092043f
C15683 DVSS.n4383 VSS 0.073894f
C15684 DVSS.n4384 VSS 0.092043f
C15685 DVSS.n4385 VSS 0.092043f
C15686 DVSS.n4386 VSS 0.092043f
C15687 DVSS.n4387 VSS 0.092043f
C15688 DVSS.n4388 VSS 0.092043f
C15689 DVSS.n4389 VSS 0.092043f
C15690 DVSS.n4390 VSS 0.092043f
C15691 DVSS.n4391 VSS 0.046022f
C15692 DVSS.n4392 VSS 0.046205f
C15693 DVSS.n4393 VSS 0.051772f
C15694 DVSS.n4394 VSS 0.253973f
C15695 DVSS.n4395 VSS 0.026956f
C15696 DVSS.n4396 VSS 0.026956f
C15697 DVSS.n4397 VSS 0.023539f
C15698 DVSS.n4398 VSS 0.046022f
C15699 DVSS.n4399 VSS 0.046022f
C15700 DVSS.n4400 VSS 0.046022f
C15701 DVSS.n4401 VSS 0.092043f
C15702 DVSS.n4402 VSS 0.092043f
C15703 DVSS.n4403 VSS 0.092043f
C15704 DVSS.n4404 VSS 0.092043f
C15705 DVSS.n4405 VSS 0.092043f
C15706 DVSS.n4406 VSS 0.046022f
C15707 DVSS.n4407 VSS 0.042497f
C15708 DVSS.n4408 VSS 0.05196f
C15709 DVSS.n4409 VSS 0.046205f
C15710 DVSS.n4410 VSS 0.092043f
C15711 DVSS.n4411 VSS 0.092043f
C15712 DVSS.n4412 VSS 0.092043f
C15713 DVSS.n4413 VSS 0.092043f
C15714 DVSS.n4414 VSS 0.046022f
C15715 DVSS.n4415 VSS 0.253973f
C15716 DVSS.n4416 VSS 0.026956f
C15717 DVSS.n4417 VSS 0.046022f
C15718 DVSS.n4418 VSS 0.092043f
C15719 DVSS.n4419 VSS 0.092043f
C15720 DVSS.n4420 VSS 0.092043f
C15721 DVSS.n4421 VSS 0.092043f
C15722 DVSS.n4422 VSS 0.092043f
C15723 DVSS.n4423 VSS 0.046022f
C15724 DVSS.n4424 VSS 0.046022f
C15725 DVSS.n4425 VSS 0.046022f
C15726 DVSS.n4426 VSS 0.026956f
C15727 DVSS.n4427 VSS 0.042497f
C15728 DVSS.n4428 VSS 0.023539f
C15729 DVSS.n4429 VSS 0.023539f
C15730 DVSS.n4430 VSS 0.026956f
C15731 DVSS.n4431 VSS 0.068967f
C15732 DVSS.n4432 VSS 0.04501f
C15733 DVSS.n4433 VSS 0.066064f
C15734 DVSS.n4434 VSS 0.046022f
C15735 DVSS.n4435 VSS 0.046022f
C15736 DVSS.n4436 VSS 0.092043f
C15737 DVSS.n4437 VSS 0.092043f
C15738 DVSS.n4438 VSS 0.092043f
C15739 DVSS.n4439 VSS 0.092043f
C15740 DVSS.n4440 VSS 0.092043f
C15741 DVSS.n4441 VSS 0.092043f
C15742 DVSS.n4442 VSS 0.092043f
C15743 DVSS.n4443 VSS 0.092043f
C15744 DVSS.n4444 VSS 0.092043f
C15745 DVSS.n4445 VSS 0.092043f
C15746 DVSS.n4446 VSS 0.046022f
C15747 DVSS.n4447 VSS 0.026956f
C15748 DVSS.n4448 VSS 0.046022f
C15749 DVSS.n4449 VSS 0.046022f
C15750 DVSS.n4450 VSS 0.042497f
C15751 DVSS.n4451 VSS 0.051772f
C15752 DVSS.n4452 VSS 0.046205f
C15753 DVSS.n4453 VSS 0.056717f
C15754 DVSS.n4454 VSS 0.092043f
C15755 DVSS.n4455 VSS 0.092043f
C15756 DVSS.n4456 VSS 0.092043f
C15757 DVSS.n4457 VSS 0.092043f
C15758 DVSS.n4458 VSS 0.092043f
C15759 DVSS.n4459 VSS 0.092043f
C15760 DVSS.n4460 VSS 0.092043f
C15761 DVSS.n4461 VSS 0.092043f
C15762 DVSS.n4462 VSS 0.092043f
C15763 DVSS.n4463 VSS 0.092043f
C15764 DVSS.n4464 VSS 0.092043f
C15765 DVSS.n4465 VSS 0.092043f
C15766 DVSS.n4466 VSS 0.092043f
C15767 DVSS.n4467 VSS 0.056393f
C15768 DVSS.n4468 VSS 0.046205f
C15769 DVSS.n4469 VSS 0.05196f
C15770 DVSS.n4470 VSS 0.259592f
C15771 DVSS.n4471 VSS 0.026956f
C15772 DVSS.n4472 VSS 0.023539f
C15773 DVSS.n4473 VSS 0.046022f
C15774 DVSS.n4474 VSS 0.046022f
C15775 DVSS.n4475 VSS 0.092043f
C15776 DVSS.n4476 VSS 0.092043f
C15777 DVSS.n4477 VSS 0.092043f
C15778 DVSS.n4478 VSS 0.092043f
C15779 DVSS.n4479 VSS 0.092043f
C15780 DVSS.n4480 VSS 0.046022f
C15781 DVSS.n4481 VSS 0.046022f
C15782 DVSS.n4482 VSS 0.042497f
C15783 DVSS.n4483 VSS 0.051772f
C15784 DVSS.n4484 VSS 0.046205f
C15785 DVSS.n4485 VSS 0.081672f
C15786 DVSS.n4486 VSS 0.092043f
C15787 DVSS.n4487 VSS 0.092043f
C15788 DVSS.n4488 VSS 0.092043f
C15789 DVSS.n4489 VSS 0.092043f
C15790 DVSS.n4490 VSS 0.092043f
C15791 DVSS.n4491 VSS 0.092043f
C15792 DVSS.n4492 VSS 0.092043f
C15793 DVSS.n4493 VSS 0.092043f
C15794 DVSS.n4494 VSS 0.076487f
C15795 DVSS.n4495 VSS 0.092043f
C15796 DVSS.n4496 VSS 0.092043f
C15797 DVSS.n4497 VSS 0.092043f
C15798 DVSS.n4498 VSS 0.092043f
C15799 DVSS.n4499 VSS 0.092043f
C15800 DVSS.n4500 VSS 0.046022f
C15801 DVSS.n4501 VSS 0.046022f
C15802 DVSS.n4502 VSS 0.023539f
C15803 DVSS.n4503 VSS 0.026956f
C15804 DVSS.n4504 VSS 0.066064f
C15805 DVSS.n4505 VSS 0.04501f
C15806 DVSS.n4506 VSS 1.30211f
C15807 DVSS.n4507 VSS 2.01475f
C15808 DVSS.n4508 VSS 2.0614f
C15809 DVSS.n4509 VSS 2.06315f
C15810 DVSS.n4510 VSS 1.33339f
C15811 DVSS.n4511 VSS 0.04501f
C15812 DVSS.n4512 VSS 0.068967f
C15813 DVSS.n4513 VSS 0.026956f
C15814 DVSS.n4514 VSS 0.023539f
C15815 DVSS.n4515 VSS 0.046022f
C15816 DVSS.n4516 VSS 0.046022f
C15817 DVSS.n4517 VSS 0.092043f
C15818 DVSS.n4518 VSS 0.092043f
C15819 DVSS.n4519 VSS 0.092043f
C15820 DVSS.n4520 VSS 0.092043f
C15821 DVSS.n4521 VSS 0.092043f
C15822 DVSS.n4522 VSS 0.046022f
C15823 DVSS.n4523 VSS 0.046022f
C15824 DVSS.n4524 VSS 0.023539f
C15825 DVSS.n4525 VSS 0.026956f
C15826 DVSS.n4526 VSS 0.259592f
C15827 DVSS.n4527 VSS 0.05196f
C15828 DVSS.n4528 VSS 0.046205f
C15829 DVSS.n4529 VSS 0.081348f
C15830 DVSS.n4530 VSS 0.092043f
C15831 DVSS.n4531 VSS 0.092043f
C15832 DVSS.n4532 VSS 0.092043f
C15833 DVSS.n4533 VSS 0.092043f
C15834 DVSS.n4534 VSS 0.092043f
C15835 DVSS.n4535 VSS 0.092043f
C15836 DVSS.n4536 VSS 0.092043f
C15837 DVSS.n4537 VSS 0.077783f
C15838 DVSS.n4538 VSS 0.092043f
C15839 DVSS.n4539 VSS 0.092043f
C15840 DVSS.n4540 VSS 0.092043f
C15841 DVSS.n4541 VSS 0.092043f
C15842 DVSS.n4542 VSS 0.092043f
C15843 DVSS.n4543 VSS 0.092043f
C15844 DVSS.n4544 VSS 0.046022f
C15845 DVSS.n4545 VSS 0.046022f
C15846 DVSS.n4546 VSS 0.046022f
C15847 DVSS.n4547 VSS 0.042497f
C15848 DVSS.n4548 VSS 0.026956f
C15849 DVSS.n4549 VSS 0.253973f
C15850 DVSS.n4550 VSS 0.04501f
C15851 DVSS.n4551 VSS 0.068967f
C15852 DVSS.n4552 VSS 0.026956f
C15853 DVSS.n4553 VSS 0.023539f
C15854 DVSS.n4554 VSS 0.046022f
C15855 DVSS.n4555 VSS 0.046022f
C15856 DVSS.n4556 VSS 0.092043f
C15857 DVSS.n4557 VSS 0.092043f
C15858 DVSS.n4558 VSS 0.092043f
C15859 DVSS.n4559 VSS 0.092043f
C15860 DVSS.n4560 VSS 0.092043f
C15861 DVSS.n4561 VSS 0.092043f
C15862 DVSS.n4562 VSS 0.046022f
C15863 DVSS.n4563 VSS 0.046022f
C15864 DVSS.n4564 VSS 0.023539f
C15865 DVSS.n4565 VSS 0.026956f
C15866 DVSS.n4566 VSS 0.259592f
C15867 DVSS.n4567 VSS 0.05196f
C15868 DVSS.n4568 VSS 0.046205f
C15869 DVSS.n4569 VSS 0.060282f
C15870 DVSS.n4570 VSS 0.092043f
C15871 DVSS.n4571 VSS 0.092043f
C15872 DVSS.n4572 VSS 0.092043f
C15873 DVSS.n4573 VSS 0.092043f
C15874 DVSS.n4574 VSS 0.092043f
C15875 DVSS.n4575 VSS 0.092043f
C15876 DVSS.n4576 VSS 0.092043f
C15877 DVSS.n4577 VSS 0.092043f
C15878 DVSS.n4578 VSS 0.092043f
C15879 DVSS.n4579 VSS 0.092043f
C15880 DVSS.n4580 VSS 0.092043f
C15881 DVSS.n4581 VSS 0.092043f
C15882 DVSS.n4582 VSS 0.092043f
C15883 DVSS.n4583 VSS 0.092043f
C15884 DVSS.n4584 VSS 0.046022f
C15885 DVSS.n4585 VSS 0.046205f
C15886 DVSS.n4586 VSS 0.051772f
C15887 DVSS.n4587 VSS 0.253973f
C15888 DVSS.n4588 VSS 0.026956f
C15889 DVSS.n4589 VSS 0.026956f
C15890 DVSS.n4590 VSS 0.023539f
C15891 DVSS.n4591 VSS 0.046022f
C15892 DVSS.n4592 VSS 0.046022f
C15893 DVSS.n4593 VSS 0.046022f
C15894 DVSS.n4594 VSS 0.092043f
C15895 DVSS.n4595 VSS 0.092043f
C15896 DVSS.n4596 VSS 0.092043f
C15897 DVSS.n4597 VSS 0.092043f
C15898 DVSS.n4598 VSS 0.092043f
C15899 DVSS.n4599 VSS 0.046022f
C15900 DVSS.n4600 VSS 0.042497f
C15901 DVSS.n4601 VSS 0.05196f
C15902 DVSS.n4602 VSS 0.046205f
C15903 DVSS.n4603 VSS 0.092043f
C15904 DVSS.n4604 VSS 0.092043f
C15905 DVSS.n4605 VSS 0.092043f
C15906 DVSS.n4606 VSS 0.092043f
C15907 DVSS.n4607 VSS 0.046022f
C15908 DVSS.n4608 VSS 0.253973f
C15909 DVSS.n4609 VSS 0.026956f
C15910 DVSS.n4610 VSS 0.046022f
C15911 DVSS.n4611 VSS 0.092043f
C15912 DVSS.n4612 VSS 0.092043f
C15913 DVSS.n4613 VSS 0.092043f
C15914 DVSS.n4614 VSS 0.092043f
C15915 DVSS.n4615 VSS 0.092043f
C15916 DVSS.n4616 VSS 0.046022f
C15917 DVSS.n4617 VSS 0.046022f
C15918 DVSS.n4618 VSS 0.046022f
C15919 DVSS.n4619 VSS 0.026956f
C15920 DVSS.n4620 VSS 0.042497f
C15921 DVSS.n4621 VSS 0.023539f
C15922 DVSS.n4622 VSS 0.023539f
C15923 DVSS.n4623 VSS 0.026956f
C15924 DVSS.n4624 VSS 0.068967f
C15925 DVSS.n4625 VSS 0.04501f
C15926 DVSS.n4626 VSS 0.066064f
C15927 DVSS.n4627 VSS 0.046022f
C15928 DVSS.n4628 VSS 0.046022f
C15929 DVSS.n4629 VSS 0.092043f
C15930 DVSS.n4630 VSS 0.092043f
C15931 DVSS.n4631 VSS 0.092043f
C15932 DVSS.n4632 VSS 0.092043f
C15933 DVSS.n4633 VSS 0.092043f
C15934 DVSS.n4634 VSS 0.092043f
C15935 DVSS.n4635 VSS 0.026298f
C15936 DVSS.n4636 VSS 0.026298f
C15937 DVSS.n4637 VSS 0.026298f
C15938 DVSS.n4638 VSS 0.026298f
C15939 DVSS.n4639 VSS 0.011482f
C15940 DVSS.n4640 VSS 0.046022f
C15941 DVSS.n4642 VSS 0.022965f
C15942 DVSS.n4644 VSS 0.022965f
C15943 DVSS.n4646 VSS 0.038351f
C15944 DVSS.n4647 VSS 0.016853f
C15945 DVSS.n4649 VSS 0.072371f
C15946 DVSS.n4651 VSS 0.028706f
C15947 DVSS.n4652 VSS 0.083196f
C15948 DVSS.n4653 VSS 0.013149f
C15949 DVSS.n4654 VSS 0.020187f
C15950 DVSS.n4655 VSS 0.026298f
C15951 DVSS.n4656 VSS 0.026298f
C15952 DVSS.n4657 VSS 0.026298f
C15953 DVSS.n4662 VSS 0.046022f
C15954 DVSS.n4663 VSS 0.046022f
C15955 DVSS.n4667 VSS 0.092043f
C15956 DVSS.n4668 VSS 0.092043f
C15957 DVSS.n4669 VSS 0.092043f
C15958 DVSS.n4670 VSS 0.092043f
C15959 DVSS.n4671 VSS 0.092043f
C15960 DVSS.n4672 VSS 0.092043f
C15961 DVSS.n4673 VSS 0.092043f
C15962 DVSS.n4674 VSS 0.092043f
C15963 DVSS.n4675 VSS 0.092043f
C15964 DVSS.n4676 VSS 0.092043f
C15965 DVSS.n4677 VSS 0.092043f
C15966 DVSS.n4678 VSS 0.047917f
C15967 DVSS.n4679 VSS 0.175694f
C15968 DVSS.n4680 VSS 0.092043f
C15969 DVSS.n4681 VSS 0.058661f
C15970 DVSS.n4682 VSS 0.051855f
C15971 DVSS.n4683 VSS 0.092043f
C15972 DVSS.n4684 VSS 0.092043f
C15973 DVSS.n4685 VSS 0.343557f
C15974 DVSS.n4686 VSS 0.090747f
C15975 DVSS.n4687 VSS 0.010371f
C15976 DVSS.n4688 VSS 0.042457f
C15977 DVSS.n4689 VSS 0.055096f
C15978 DVSS.n4690 VSS 0.082968f
C15979 DVSS.n4691 VSS 0.082968f
C15980 DVSS.n4692 VSS 0.092043f
C15981 DVSS.n4693 VSS 0.092043f
C15982 DVSS.n4694 VSS 0.092043f
C15983 DVSS.n4695 VSS 0.092043f
C15984 DVSS.n4696 VSS 0.092043f
C15985 DVSS.n4697 VSS 0.092043f
C15986 DVSS.n4698 VSS 0.092043f
C15987 DVSS.n4699 VSS 0.092043f
C15988 DVSS.n4700 VSS 0.092043f
C15989 DVSS.n4701 VSS 0.092043f
C15990 DVSS.n4702 VSS 0.092043f
C15991 DVSS.n4703 VSS 0.056717f
C15992 DVSS.n4704 VSS 0.046022f
C15993 DVSS.n4706 VSS 0.024446f
C15994 DVSS.n4707 VSS 0.046022f
C15995 DVSS.n4708 VSS 0.081348f
C15996 DVSS.n4709 VSS 0.092043f
C15997 DVSS.n4710 VSS 0.092043f
C15998 DVSS.n4711 VSS 0.092043f
C15999 DVSS.n4712 VSS 0.092043f
C16000 DVSS.n4713 VSS 0.092043f
C16001 DVSS.n4714 VSS 0.092043f
C16002 DVSS.n4715 VSS 0.064495f
C16003 DVSS.n4716 VSS 0.046205f
C16004 DVSS.n4717 VSS 0.05196f
C16005 DVSS.n4718 VSS 0.259592f
C16006 DVSS.n4719 VSS 0.026956f
C16007 DVSS.n4720 VSS 0.023539f
C16008 DVSS.n4721 VSS 0.046022f
C16009 DVSS.n4722 VSS 0.046022f
C16010 DVSS.n4723 VSS 0.092043f
C16011 DVSS.n4724 VSS 0.092043f
C16012 DVSS.n4725 VSS 0.092043f
C16013 DVSS.n4726 VSS 0.092043f
C16014 DVSS.n4727 VSS 0.092043f
C16015 DVSS.n4728 VSS 0.046022f
C16016 DVSS.n4729 VSS 0.046022f
C16017 DVSS.n4730 VSS 0.042497f
C16018 DVSS.n4731 VSS 0.051772f
C16019 DVSS.n4732 VSS 0.046205f
C16020 DVSS.n4733 VSS 0.07357f
C16021 DVSS.n4734 VSS 0.092043f
C16022 DVSS.n4735 VSS 0.092043f
C16023 DVSS.n4736 VSS 0.092043f
C16024 DVSS.n4737 VSS 0.092043f
C16025 DVSS.n4738 VSS 0.092043f
C16026 DVSS.n4739 VSS 0.092043f
C16027 DVSS.n4740 VSS 0.092043f
C16028 DVSS.n4741 VSS 0.092043f
C16029 DVSS.n4742 VSS 0.086534f
C16030 DVSS.n4743 VSS 0.092043f
C16031 DVSS.n4744 VSS 0.092043f
C16032 DVSS.n4745 VSS 0.092043f
C16033 DVSS.n4746 VSS 0.092043f
C16034 DVSS.n4747 VSS 0.092043f
C16035 DVSS.n4748 VSS 0.046022f
C16036 DVSS.n4749 VSS 0.046022f
C16037 DVSS.n4750 VSS 0.023539f
C16038 DVSS.n4751 VSS 0.026956f
C16039 DVSS.n4752 VSS 0.066064f
C16040 DVSS.n4753 VSS 0.04501f
C16041 DVSS.n4754 VSS 1.33301f
C16042 DVSS.n4755 VSS 2.06257f
C16043 DVSS.n4756 VSS 2.02116f
C16044 DVSS.t164 VSS 0.209479f
C16045 DVSS.t156 VSS 0.320854f
C16046 DVSS.t152 VSS 0.338667f
C16047 DVSS.t154 VSS 0.24732f
C16048 DVSS.n4757 VSS 0.16488f
C16049 DVSS.t120 VSS 0.24732f
C16050 DVSS.t97 VSS 0.266917f
C16051 DVSS.n4758 VSS 0.500008f
C16052 DVSS.n4759 VSS 1.19949f
C16053 DVSS.n4760 VSS 0.713052f
C16054 DVSS.n4761 VSS 2.8251f
C16055 DVSS.n4762 VSS 1.42519f
C16056 DVSS.n4763 VSS 2.36089f
C16057 DVSS.n4764 VSS 3.45644f
C16058 DVSS.n4765 VSS 2.15335f
C16059 DVSS.n4766 VSS 1.08837f
C16060 DVSS.n4767 VSS 0.02426f
C16061 DVSS.n4768 VSS 0.698357f
C16062 DVSS.n4769 VSS 0.682325f
C16063 DVSS.n4770 VSS 0.036947f
C16064 DVSS.n4771 VSS 0.341018f
C16065 DVSS.n4772 VSS 0.813798f
C16066 DVSS.n4773 VSS 0.38022f
C16067 DVSS.n4774 VSS 0.197235f
C16068 DVSS.n4775 VSS 0.197235f
C16069 DVSS.n4776 VSS 0.111813f
C16070 DVSS.n4777 VSS 0.136849f
C16071 DVSS.n4778 VSS 0.079717f
C16072 DVSS.n4779 VSS 0.026357f
C16073 DVSS.n4780 VSS 0.024125f
C16074 DVSS.n4781 VSS 0.02551f
C16075 DVSS.n4782 VSS -0.047747f
C16076 DVSS.n4783 VSS 0.168046f
C16077 DVSS.t17 VSS 0.329761f
C16078 DVSS.t128 VSS 0.265565f
C16079 DVSS.n4784 VSS 0.16488f
C16080 DVSS.n4785 VSS 0.04679f
C16081 DVSS.n4786 VSS 0.021032f
C16082 DVSS.n4787 VSS 0.025192f
C16083 DVSS.n4788 VSS 0.093193f
C16084 DVSS.n4789 VSS 0.02356f
C16085 DVSS.n4790 VSS 0.129078f
C16086 DVSS.n4791 VSS 0.117369f
C16087 DVSS.n4792 VSS 0.197235f
C16088 DVSS.n4793 VSS 0.197235f
C16089 DVSS.n4794 VSS 0.197235f
C16090 DVSS.n4795 VSS 0.197235f
C16091 DVSS.n4796 VSS 0.197235f
C16092 DVSS.n4797 VSS 0.197235f
C16093 DVSS.n4798 VSS 0.197235f
C16094 DVSS.n4799 VSS 0.197235f
C16095 DVSS.n4800 VSS 0.197235f
C16096 DVSS.n4801 VSS 0.111813f
C16097 DVSS.n4802 VSS 0.126367f
C16098 DVSS.n4803 VSS 0.032017f
C16099 DVSS.t180 VSS 0.014445f
C16100 DVSS.n4804 VSS 0.002551f
C16101 DVSS.n4805 VSS 0.038498f
C16102 DVSS.n4806 VSS 0.009596f
C16103 DVSS.n4807 VSS 0.035876f
C16104 DVSS.n4808 VSS -0.047747f
C16105 DVSS.n4809 VSS 0.212645f
C16106 DVSS.t8 VSS 0.329761f
C16107 DVSS.t167 VSS 0.265565f
C16108 DVSS.t179 VSS 0.258808f
C16109 DVSS.n4810 VSS 0.16488f
C16110 DVSS.n4811 VSS 0.04679f
C16111 DVSS.t68 VSS 0.328409f
C16112 DVSS.t64 VSS 0.24732f
C16113 DVSS.t36 VSS 0.238536f
C16114 DVSS.t70 VSS 0.329761f
C16115 DVSS.t66 VSS 0.24732f
C16116 DVSS.n4812 VSS 0.16488f
C16117 DVSS.n4813 VSS 0.049774f
C16118 DVSS.n4814 VSS 0.026861f
C16119 DVSS.n4815 VSS 0.018385f
C16120 DVSS.t67 VSS 0.014445f
C16121 DVSS.n4816 VSS 0.028891f
C16122 DVSS.n4817 VSS 0.012058f
C16123 DVSS.n4818 VSS 0.024125f
C16124 DVSS.t69 VSS 0.014445f
C16125 DVSS.n4819 VSS 0.038498f
C16126 DVSS.n4820 VSS 0.012005f
C16127 DVSS.n4821 VSS 0.010866f
C16128 DVSS.n4822 VSS 0.027768f
C16129 DVSS.n4823 VSS 0.093262f
C16130 DVSS.n4824 VSS 0.323003f
C16131 DVSS.t162 VSS 0.395307f
C16132 DVSS.n4825 VSS 0.194847f
C16133 DVSS.t74 VSS 0.056671f
C16134 DVSS.n4826 VSS 0.119236f
C16135 DVSS.n4827 VSS 0.002225f
C16136 DVSS.n4828 VSS 0.211123f
C16137 DVSS.n4829 VSS 0.139085f
C16138 DVSS.n4830 VSS 0.250312f
C16139 DVSS.n4831 VSS 0.233544f
C16140 DVSS.n4832 VSS 0.004267f
C16141 DVSS.n4833 VSS 0.004267f
C16142 DVSS.n4834 VSS 0.069463f
C16143 DVSS.n4835 VSS 0.019351f
C16144 DVSS.n4836 VSS 0.017161f
C16145 DVSS.n4837 VSS -0.005991f
C16146 DVSS.n4838 VSS 0.296597f
C16147 DVSS.n4839 VSS 0.443265f
C16148 DVSS.n4840 VSS 0.030185f
C16149 DVSS.n4841 VSS 0.014912f
C16150 DVSS.n4842 VSS 0.017161f
C16151 DVSS.n4843 VSS -0.005991f
C16152 DVSS.n4844 VSS 0.004267f
C16153 DVSS.n4845 VSS 0.004267f
C16154 DVSS.n4846 VSS 0.069463f
C16155 DVSS.n4847 VSS 0.019351f
C16156 DVSS.n4848 VSS 0.233544f
C16157 DVSS.n4849 VSS 0.250312f
C16158 DVSS.n4850 VSS 0.139085f
C16159 DVSS.n4851 VSS 0.211123f
C16160 DVSS.t83 VSS 0.17128f
C16161 DVSS.n4852 VSS 0.06131f
C16162 DVSS.n4853 VSS 0.002225f
C16163 DVSS.n4854 VSS 0.010533f
C16164 DVSS.n4855 VSS 0.020138f
C16165 DVSS.n4856 VSS 0.063438f
C16166 DVSS.n4857 VSS 0.352065f
C16167 DVSS.t165 VSS 0.17128f
C16168 DVSS.n4858 VSS 0.06131f
C16169 DVSS.n4859 VSS 0.002225f
C16170 DVSS.n4860 VSS 0.211123f
C16171 DVSS.n4861 VSS 0.139085f
C16172 DVSS.n4862 VSS 0.250312f
C16173 DVSS.n4863 VSS 0.017161f
C16174 DVSS.n4864 VSS -0.005991f
C16175 DVSS.n4865 VSS 0.004267f
C16176 DVSS.n4866 VSS 0.004267f
C16177 DVSS.n4867 VSS 0.069463f
C16178 DVSS.n4868 VSS 0.019351f
C16179 DVSS.n4869 VSS 0.187977f
C16180 DVSS.n4870 VSS 0.958555f
C16181 DVSS.n4871 VSS 0.008144f
C16182 DVSS.n4872 VSS 0.013242f
C16183 DVSS.n4874 VSS 0.015742f
C16184 DVSS.n4877 VSS 0.026298f
C16185 DVSS.n4878 VSS 0.046022f
C16186 DVSS.n4879 VSS 0.026298f
C16187 DVSS.n4880 VSS 0.026298f
C16188 DVSS.n4882 VSS 0.026298f
C16189 DVSS.n4885 VSS 0.036947f
C16190 DVSS.n4887 VSS 0.02315f
C16191 DVSS.n4888 VSS 0.046022f
C16192 DVSS.n4889 VSS 0.017825f
C16193 DVSS.n4890 VSS 0.055096f
C16194 DVSS.n4891 VSS 0.047318f
C16195 DVSS.n4892 VSS 0.092043f
C16196 DVSS.n4893 VSS 0.092043f
C16197 DVSS.n4894 VSS 0.092043f
C16198 DVSS.n4895 VSS 0.054772f
C16199 DVSS.n4896 VSS 0.092043f
C16200 DVSS.n4897 VSS 0.092043f
C16201 DVSS.n4898 VSS 0.092043f
C16202 DVSS.n4899 VSS 0.092043f
C16203 DVSS.n4900 VSS 0.092043f
C16204 DVSS.n4901 VSS 0.092043f
C16205 DVSS.n4902 VSS 0.092043f
C16206 DVSS.n4903 VSS 0.092043f
C16207 DVSS.n4904 VSS 0.092043f
C16208 DVSS.n4905 VSS 0.092043f
C16209 DVSS.n4906 VSS 0.092043f
C16210 DVSS.n4907 VSS 0.092043f
C16211 DVSS.n4908 VSS 0.092043f
C16212 DVSS.n4909 VSS 0.092043f
C16213 DVSS.n4910 VSS 0.092043f
C16214 DVSS.n4911 VSS 0.092043f
C16215 DVSS.n4912 VSS 0.092043f
C16216 DVSS.n4913 VSS 0.092043f
C16217 DVSS.n4914 VSS 0.092043f
C16218 DVSS.n4915 VSS 0.092043f
C16219 DVSS.n4916 VSS 0.092043f
C16220 DVSS.n4917 VSS 0.092043f
C16221 DVSS.n4918 VSS 0.092043f
C16222 DVSS.n4919 VSS 0.092043f
C16223 DVSS.n4920 VSS 0.092043f
C16224 DVSS.n4921 VSS 0.092043f
C16225 DVSS.n4922 VSS 0.092043f
C16226 DVSS.n4923 VSS 0.092043f
C16227 DVSS.n4924 VSS 0.092043f
C16228 DVSS.n4925 VSS 0.092043f
C16229 DVSS.n4926 VSS 0.092043f
C16230 DVSS.n4927 VSS 0.092043f
C16231 DVSS.n4928 VSS 0.092043f
C16232 DVSS.n4929 VSS 0.092043f
C16233 DVSS.n4930 VSS 0.092043f
C16234 DVSS.n4931 VSS 0.092043f
C16235 DVSS.n4932 VSS 0.092043f
C16236 DVSS.n4933 VSS 0.092043f
C16237 DVSS.n4934 VSS 0.092043f
C16238 DVSS.n4935 VSS 0.092043f
C16239 DVSS.n4936 VSS 0.092043f
C16240 DVSS.n4937 VSS 0.092043f
C16241 DVSS.n4938 VSS 0.092043f
C16242 DVSS.n4939 VSS 0.092043f
C16243 DVSS.n4940 VSS 0.092043f
C16244 DVSS.n4941 VSS 0.092043f
C16245 DVSS.n4942 VSS 0.092043f
C16246 DVSS.n4943 VSS 0.092043f
C16247 DVSS.n4944 VSS 0.092043f
C16248 DVSS.n4945 VSS 0.092043f
C16249 DVSS.n4946 VSS 0.092043f
C16250 DVSS.n4947 VSS 0.092043f
C16251 DVSS.n4948 VSS 0.092043f
C16252 DVSS.n4949 VSS 0.092043f
C16253 DVSS.n4950 VSS 0.092043f
C16254 DVSS.n4951 VSS 0.092043f
C16255 DVSS.n4952 VSS 0.092043f
C16256 DVSS.n4953 VSS 0.092043f
C16257 DVSS.n4954 VSS 0.092043f
C16258 DVSS.n4955 VSS 0.092043f
C16259 DVSS.n4956 VSS 0.092043f
C16260 DVSS.n4957 VSS 0.092043f
C16261 DVSS.n4958 VSS 0.092043f
C16262 DVSS.n4959 VSS 0.092043f
C16263 DVSS.n4960 VSS 0.092043f
C16264 DVSS.n4961 VSS 0.092043f
C16265 DVSS.n4962 VSS 0.092043f
C16266 DVSS.n4963 VSS 0.092043f
C16267 DVSS.n4964 VSS 0.092043f
C16268 DVSS.n4965 VSS 0.092043f
C16269 DVSS.n4966 VSS 0.092043f
C16270 DVSS.n4967 VSS 0.077783f
C16271 DVSS.n4968 VSS 0.092043f
C16272 DVSS.n4969 VSS 0.092043f
C16273 DVSS.n4970 VSS 0.092043f
C16274 DVSS.n4971 VSS 0.092043f
C16275 DVSS.n4972 VSS 0.092043f
C16276 DVSS.n4973 VSS 0.092043f
C16277 DVSS.n4974 VSS 0.092043f
C16278 DVSS.n4975 VSS 0.092043f
C16279 DVSS.n4976 VSS 0.092043f
C16280 DVSS.n4977 VSS 0.092043f
C16281 DVSS.n4978 VSS 0.092043f
C16282 DVSS.n4979 VSS 0.092043f
C16283 DVSS.n4980 VSS 0.092043f
C16284 DVSS.n4981 VSS 0.092043f
C16285 DVSS.n4982 VSS 0.092043f
C16286 DVSS.n4983 VSS 0.092043f
C16287 DVSS.n4984 VSS 0.092043f
C16288 DVSS.n4985 VSS 0.092043f
C16289 DVSS.n4986 VSS 0.092043f
C16290 DVSS.n4987 VSS 0.092043f
C16291 DVSS.n4988 VSS 0.092043f
C16292 DVSS.n4989 VSS 0.092043f
C16293 DVSS.n4990 VSS 0.092043f
C16294 DVSS.n4991 VSS 0.092043f
C16295 DVSS.n4992 VSS 0.092043f
C16296 DVSS.n4993 VSS 0.092043f
C16297 DVSS.n4994 VSS 0.092043f
C16298 DVSS.n4995 VSS 0.092043f
C16299 DVSS.n4996 VSS 0.092043f
C16300 DVSS.n4997 VSS 0.092043f
C16301 DVSS.n4998 VSS 0.092043f
C16302 DVSS.n4999 VSS 0.092043f
C16303 DVSS.n5000 VSS 0.092043f
C16304 DVSS.n5001 VSS 0.092043f
C16305 DVSS.n5002 VSS 0.092043f
C16306 DVSS.n5003 VSS 0.092043f
C16307 DVSS.n5004 VSS 0.092043f
C16308 DVSS.n5005 VSS 0.092043f
C16309 DVSS.n5006 VSS 0.092043f
C16310 DVSS.n5007 VSS 0.092043f
C16311 DVSS.n5008 VSS 0.092043f
C16312 DVSS.n5009 VSS 0.092043f
C16313 DVSS.n5010 VSS 0.092043f
C16314 DVSS.n5011 VSS 0.092043f
C16315 DVSS.n5012 VSS 0.092043f
C16316 DVSS.n5013 VSS 0.092043f
C16317 DVSS.n5014 VSS 0.092043f
C16318 DVSS.n5015 VSS 0.092043f
C16319 DVSS.n5016 VSS 0.092043f
C16320 DVSS.n5017 VSS 0.092043f
C16321 DVSS.n5018 VSS 0.092043f
C16322 DVSS.n5019 VSS 0.092043f
C16323 DVSS.n5020 VSS 0.092043f
C16324 DVSS.n5021 VSS 0.092043f
C16325 DVSS.n5022 VSS 0.092043f
C16326 DVSS.n5023 VSS 0.092043f
C16327 DVSS.n5024 VSS 0.092043f
C16328 DVSS.n5025 VSS 0.051855f
C16329 DVSS.n5026 VSS 0.092043f
C16330 DVSS.n5027 VSS 0.092043f
C16331 DVSS.n5028 VSS 0.092043f
C16332 DVSS.n5029 VSS 0.092043f
C16333 DVSS.n5030 VSS 0.092043f
C16334 DVSS.n5031 VSS 0.046022f
C16335 DVSS.n5032 VSS 0.046022f
C16336 DVSS.n5033 VSS 0.004997f
C16337 DVSS.n5034 VSS 0.003413f
C16338 DVSS.n5035 VSS 0.046022f
C16339 DVSS.n5036 VSS 0.046022f
C16340 DVSS.n5037 VSS 0.092043f
C16341 DVSS.n5038 VSS 0.092043f
C16342 DVSS.n5039 VSS 0.092043f
C16343 DVSS.n5040 VSS 0.092043f
C16344 DVSS.n5041 VSS 0.092043f
C16345 DVSS.n5042 VSS 0.046022f
C16346 DVSS.n5043 VSS 0.046022f
C16347 DVSS.n5044 VSS 0.010593f
C16348 DVSS.n5045 VSS 0.046231f
C16349 DVSS.n5046 VSS 0.086209f
C16350 DVSS.n5047 VSS 0.092043f
C16351 DVSS.n5048 VSS 0.092043f
C16352 DVSS.n5049 VSS 0.092043f
C16353 DVSS.n5050 VSS 0.092043f
C16354 DVSS.n5051 VSS 0.092043f
C16355 DVSS.n5052 VSS 0.092043f
C16356 DVSS.n5053 VSS 0.092043f
C16357 DVSS.n5054 VSS 0.092043f
C16358 DVSS.n5055 VSS 0.092043f
C16359 DVSS.n5056 VSS 0.092043f
C16360 DVSS.n5057 VSS 0.092043f
C16361 DVSS.n5058 VSS 0.092043f
C16362 DVSS.n5059 VSS 0.092043f
C16363 DVSS.n5060 VSS 0.092043f
C16364 DVSS.n5061 VSS 0.046022f
C16365 DVSS.n5062 VSS 0.058329f
C16366 DVSS.n5063 VSS 0.088478f
C16367 DVSS.n5064 VSS 0.092043f
C16368 DVSS.n5065 VSS 0.092043f
C16369 DVSS.n5066 VSS 0.092043f
C16370 DVSS.n5067 VSS 0.092043f
C16371 DVSS.n5068 VSS 0.092043f
C16372 DVSS.n5069 VSS 0.092043f
C16373 DVSS.n5070 VSS 0.092043f
C16374 DVSS.n5071 VSS 0.092043f
C16375 DVSS.n5072 VSS 0.092043f
C16376 DVSS.n5073 VSS 0.092043f
C16377 DVSS.n5074 VSS 0.092043f
C16378 DVSS.n5075 VSS 0.092043f
C16379 DVSS.n5076 VSS 0.092043f
C16380 DVSS.n5077 VSS 0.092043f
C16381 DVSS.n5078 VSS 0.092043f
C16382 DVSS.n5079 VSS 0.092043f
C16383 DVSS.n5080 VSS 0.092043f
C16384 DVSS.n5081 VSS 0.092043f
C16385 DVSS.n5082 VSS 0.092043f
C16386 DVSS.n5083 VSS 0.092043f
C16387 DVSS.n5084 VSS 0.092043f
C16388 DVSS.n5085 VSS 0.092043f
C16389 DVSS.n5086 VSS 0.092043f
C16390 DVSS.n5087 VSS 0.092043f
C16391 DVSS.n5088 VSS 0.092043f
C16392 DVSS.n5089 VSS 0.092043f
C16393 DVSS.n5090 VSS 0.341066f
C16394 DVSS.n5091 VSS 0.173028f
C16395 DVSS.n5092 VSS 0.196174f
C16396 DVSS.n5093 VSS 0.673022f
C16397 DVSS.n5094 VSS 0.827135f
C16398 DVSS.n5095 VSS 1.35909f
C16399 DVSS.n5096 VSS 1.88682f
C16400 DVSS.n5097 VSS 1.93316f
C16401 DVSS.n5098 VSS 1.8219f
C16402 DVSS.n5099 VSS 0.468957f
C16403 DVSS.n5100 VSS 0.029222f
C16404 DVSS.n5101 VSS 0.029222f
C16405 DVSS.n5102 VSS 0.012286f
C16406 DVSS.n5103 VSS 0.789346f
C16407 DVSS.n5104 VSS 0.789346f
C16408 DVSS.n5105 VSS 0.789346f
C16409 DVSS.n5106 VSS 0.012286f
C16410 DVSS.n5107 VSS 0.029222f
C16411 DVSS.n5108 VSS 0.029222f
C16412 DVSS.n5109 VSS 0.029222f
C16413 DVSS.n5110 VSS 0.012286f
C16414 DVSS.n5111 VSS 0.789346f
C16415 DVSS.n5112 VSS 0.789346f
C16416 DVSS.n5113 VSS 0.789346f
C16417 DVSS.n5114 VSS 0.012286f
C16418 DVSS.n5115 VSS 0.029222f
C16419 DVSS.n5116 VSS 0.029222f
C16420 DVSS.n5117 VSS 0.029222f
C16421 DVSS.n5118 VSS 0.012286f
C16422 DVSS.n5119 VSS 0.789346f
C16423 DVSS.n5120 VSS 0.789346f
C16424 DVSS.n5121 VSS 0.789346f
C16425 DVSS.n5122 VSS 0.012286f
C16426 DVSS.n5123 VSS 0.029222f
C16427 DVSS.n5124 VSS 0.029222f
C16428 DVSS.n5125 VSS 0.029222f
C16429 DVSS.n5126 VSS 0.012286f
C16430 DVSS.n5127 VSS 0.789346f
C16431 DVSS.n5128 VSS 0.789346f
C16432 DVSS.n5129 VSS 0.789346f
C16433 DVSS.n5130 VSS 0.012286f
C16434 DVSS.n5131 VSS 0.029222f
C16435 DVSS.n5132 VSS 0.029222f
C16436 DVSS.n5133 VSS 0.029222f
C16437 DVSS.n5134 VSS 0.012286f
C16438 DVSS.n5135 VSS 0.789346f
C16439 DVSS.n5136 VSS 0.789346f
C16440 DVSS.n5137 VSS 0.789346f
C16441 DVSS.n5138 VSS 0.012286f
C16442 DVSS.n5139 VSS 0.029222f
C16443 DVSS.n5140 VSS 0.029222f
C16444 DVSS.n5141 VSS 0.029222f
C16445 DVSS.n5142 VSS 0.012286f
C16446 DVSS.n5143 VSS 0.789346f
C16447 DVSS.n5144 VSS 0.789346f
C16448 DVSS.n5145 VSS 0.789346f
C16449 DVSS.n5146 VSS 0.012286f
C16450 DVSS.n5147 VSS 0.029222f
C16451 DVSS.n5148 VSS 0.029222f
C16452 DVSS.n5149 VSS 0.029222f
C16453 DVSS.n5150 VSS 0.012286f
C16454 DVSS.n5151 VSS 0.789346f
C16455 DVSS.n5152 VSS 0.789346f
C16456 DVSS.n5153 VSS 0.789346f
C16457 DVSS.n5154 VSS 0.012286f
C16458 DVSS.n5155 VSS 0.029222f
C16459 DVSS.n5156 VSS 0.029222f
C16460 DVSS.n5157 VSS 0.029222f
C16461 DVSS.n5158 VSS 0.012286f
C16462 DVSS.n5159 VSS 0.789346f
C16463 DVSS.n5160 VSS 0.789346f
C16464 DVSS.n5161 VSS 0.789346f
C16465 DVSS.n5162 VSS 0.012286f
C16466 DVSS.n5163 VSS 0.029222f
C16467 DVSS.n5164 VSS 0.029222f
C16468 DVSS.n5165 VSS 0.029222f
C16469 DVSS.n5166 VSS 0.012286f
C16470 DVSS.n5167 VSS 0.789346f
C16471 DVSS.n5168 VSS 0.789346f
C16472 DVSS.n5169 VSS 0.789346f
C16473 DVSS.n5170 VSS 0.012286f
C16474 DVSS.n5171 VSS 0.029222f
C16475 DVSS.n5172 VSS 0.029222f
C16476 DVSS.n5173 VSS 0.029222f
C16477 DVSS.n5174 VSS 0.012286f
C16478 DVSS.n5175 VSS 0.789346f
C16479 DVSS.n5176 VSS 0.789346f
C16480 DVSS.n5177 VSS 0.789346f
C16481 DVSS.n5178 VSS 0.012286f
C16482 DVSS.n5179 VSS 0.029222f
C16483 DVSS.n5180 VSS 0.029222f
C16484 DVSS.n5181 VSS 0.029222f
C16485 DVSS.n5182 VSS 0.012286f
C16486 DVSS.n5183 VSS 0.789346f
C16487 DVSS.n5184 VSS 0.789346f
C16488 DVSS.n5185 VSS 0.789346f
C16489 DVSS.n5186 VSS 0.012286f
C16490 DVSS.n5187 VSS 0.029222f
C16491 DVSS.n5188 VSS 0.029222f
C16492 DVSS.n5189 VSS 0.029222f
C16493 DVSS.n5190 VSS 0.012286f
C16494 DVSS.n5191 VSS 0.789346f
C16495 DVSS.n5192 VSS 0.789346f
C16496 DVSS.n5193 VSS 0.789346f
C16497 DVSS.n5194 VSS 0.012286f
C16498 DVSS.n5195 VSS 0.029222f
C16499 DVSS.n5196 VSS 0.029222f
C16500 DVSS.n5197 VSS 0.029222f
C16501 DVSS.n5198 VSS 0.012286f
C16502 DVSS.n5199 VSS 0.789346f
C16503 DVSS.n5200 VSS 0.789346f
C16504 DVSS.n5201 VSS 0.789346f
C16505 DVSS.n5202 VSS 0.012286f
C16506 DVSS.n5203 VSS 0.029222f
C16507 DVSS.n5204 VSS 0.029222f
C16508 DVSS.n5205 VSS 0.029222f
C16509 DVSS.n5206 VSS 0.029222f
C16510 DVSS.n5207 VSS 0.012286f
C16511 DVSS.n5208 VSS 0.789346f
C16512 DVSS.n5209 VSS 0.789346f
C16513 DVSS.n5210 VSS 0.789346f
C16514 DVSS.n5211 VSS 0.012286f
C16515 DVSS.n5212 VSS 0.012286f
C16516 DVSS.n5213 VSS 0.021799f
C16517 DVSS.n5214 VSS 0.014611f
C16518 DVSS.n5215 VSS 2.3203f
C16519 DVSS.n5216 VSS 0.394673f
C16520 DVSS.n5217 VSS 0.595193f
C16521 DVSS.n5218 VSS 0.789346f
C16522 DVSS.n5219 VSS 0.012286f
C16523 DVSS.n5220 VSS 0.029222f
C16524 DVSS.n5221 VSS 0.029222f
C16525 DVSS.n5222 VSS 0.029222f
C16526 DVSS.n5223 VSS 0.012286f
C16527 DVSS.n5224 VSS 0.789346f
C16528 DVSS.n5225 VSS 0.789346f
C16529 DVSS.n5226 VSS 0.789346f
C16530 DVSS.n5227 VSS 0.012286f
C16531 DVSS.n5228 VSS 0.029222f
C16532 DVSS.n5229 VSS 0.029222f
C16533 DVSS.n5230 VSS 0.029222f
C16534 DVSS.n5231 VSS 0.012286f
C16535 DVSS.n5232 VSS 0.789346f
C16536 DVSS.n5233 VSS 0.789346f
C16537 DVSS.n5234 VSS 0.789346f
C16538 DVSS.n5235 VSS 0.012286f
C16539 DVSS.n5236 VSS 0.029222f
C16540 DVSS.n5237 VSS 0.029222f
C16541 DVSS.n5238 VSS 0.029222f
C16542 DVSS.n5239 VSS 0.012286f
C16543 DVSS.n5240 VSS 0.789346f
C16544 DVSS.n5241 VSS 0.789346f
C16545 DVSS.n5242 VSS 0.789346f
C16546 DVSS.n5243 VSS 0.012286f
C16547 DVSS.n5244 VSS 0.029222f
C16548 DVSS.n5245 VSS 0.029222f
C16549 DVSS.n5246 VSS 0.029222f
C16550 DVSS.n5247 VSS 0.012286f
C16551 DVSS.n5248 VSS 0.789346f
C16552 DVSS.n5249 VSS 0.789346f
C16553 DVSS.n5250 VSS 0.789346f
C16554 DVSS.n5251 VSS 0.012286f
C16555 DVSS.n5252 VSS 0.029222f
C16556 DVSS.n5253 VSS 0.029222f
C16557 DVSS.n5254 VSS 0.029222f
C16558 DVSS.n5255 VSS 0.012286f
C16559 DVSS.n5256 VSS 0.789346f
C16560 DVSS.n5257 VSS 0.789346f
C16561 DVSS.n5258 VSS 0.789346f
C16562 DVSS.n5259 VSS 0.012286f
C16563 DVSS.n5260 VSS 0.029222f
C16564 DVSS.n5261 VSS 0.029222f
C16565 DVSS.n5262 VSS 0.029222f
C16566 DVSS.n5263 VSS 0.012286f
C16567 DVSS.n5264 VSS 0.789346f
C16568 DVSS.n5265 VSS 0.789346f
C16569 DVSS.n5266 VSS 0.789346f
C16570 DVSS.n5267 VSS 0.012286f
C16571 DVSS.n5268 VSS 0.029222f
C16572 DVSS.n5269 VSS 0.029222f
C16573 DVSS.n5270 VSS 0.029222f
C16574 DVSS.n5271 VSS 0.012286f
C16575 DVSS.n5272 VSS 0.789346f
C16576 DVSS.n5273 VSS 0.789346f
C16577 DVSS.n5274 VSS 0.789346f
C16578 DVSS.n5275 VSS 0.012286f
C16579 DVSS.n5276 VSS 0.029222f
C16580 DVSS.n5277 VSS 0.029222f
C16581 DVSS.n5278 VSS 0.029222f
C16582 DVSS.n5279 VSS 0.012286f
C16583 DVSS.n5280 VSS 0.789346f
C16584 DVSS.n5281 VSS 0.789346f
C16585 DVSS.n5282 VSS 0.789346f
C16586 DVSS.n5283 VSS 0.012286f
C16587 DVSS.n5284 VSS 0.029222f
C16588 DVSS.n5285 VSS 0.029222f
C16589 DVSS.n5286 VSS 0.029222f
C16590 DVSS.n5287 VSS 0.012286f
C16591 DVSS.n5288 VSS 0.789346f
C16592 DVSS.n5289 VSS 0.789346f
C16593 DVSS.n5290 VSS 0.789346f
C16594 DVSS.n5291 VSS 0.012286f
C16595 DVSS.n5292 VSS 0.029222f
C16596 DVSS.n5293 VSS 0.029222f
C16597 DVSS.n5294 VSS 0.029222f
C16598 DVSS.n5295 VSS 0.012286f
C16599 DVSS.n5296 VSS 0.789346f
C16600 DVSS.n5297 VSS 0.789346f
C16601 DVSS.n5298 VSS 0.789346f
C16602 DVSS.n5299 VSS 0.012286f
C16603 DVSS.n5300 VSS 0.029222f
C16604 DVSS.n5301 VSS 0.029222f
C16605 DVSS.n5302 VSS 0.029222f
C16606 DVSS.n5303 VSS 0.012286f
C16607 DVSS.n5304 VSS 0.789346f
C16608 DVSS.n5305 VSS 0.789346f
C16609 DVSS.n5306 VSS 0.789346f
C16610 DVSS.n5307 VSS 0.012286f
C16611 DVSS.n5308 VSS 0.029222f
C16612 DVSS.n5309 VSS 0.029222f
C16613 DVSS.n5310 VSS 0.029222f
C16614 DVSS.n5311 VSS 0.012286f
C16615 DVSS.n5312 VSS 0.789346f
C16616 DVSS.n5313 VSS 0.789346f
C16617 DVSS.n5314 VSS 0.789346f
C16618 DVSS.n5315 VSS 0.012286f
C16619 DVSS.n5316 VSS 0.029222f
C16620 DVSS.n5317 VSS 0.029222f
C16621 DVSS.n5318 VSS 0.029222f
C16622 DVSS.n5319 VSS 0.012286f
C16623 DVSS.n5320 VSS 0.789346f
C16624 DVSS.n5321 VSS 0.789346f
C16625 DVSS.n5322 VSS 0.789346f
C16626 DVSS.n5323 VSS 0.012286f
C16627 DVSS.n5324 VSS 0.029222f
C16628 DVSS.n5325 VSS 0.029222f
C16629 DVSS.n5326 VSS 0.029222f
C16630 DVSS.n5327 VSS 0.029222f
C16631 DVSS.n5328 VSS 0.012286f
C16632 DVSS.n5329 VSS 0.789346f
C16633 DVSS.n5330 VSS 0.789346f
C16634 DVSS.n5331 VSS 0.556998f
C16635 DVSS.n5332 VSS 0.012286f
C16636 DVSS.n5333 VSS 1.92749f
C16637 DVSS.n5334 VSS 0.388601f
C16638 DVSS.n5335 VSS 1.13563f
C16639 DVSS.n5336 VSS 1.79392f
C16640 DVSS.n5337 VSS 6.01726f
C16641 DVSS.n5338 VSS 2.39903f
C16642 DVSS.n5339 VSS 2.39868f
C16643 DVSS.n5340 VSS 4.38371f
C16644 DVSS.n5341 VSS 2.06722f
C16645 DVSS.n5342 VSS 3.35559f
C16646 DVSS.n5343 VSS 0.045844f
C16647 DVSS.n5344 VSS 0.047323f
C16648 DVSS.n5345 VSS 0.049319f
C16649 DVSS.n5346 VSS 0.079403f
C16650 DVSS.n5347 VSS 0.092043f
C16651 DVSS.n5348 VSS 0.092043f
C16652 DVSS.n5349 VSS 0.092043f
C16653 DVSS.n5350 VSS 0.092043f
C16654 DVSS.n5351 VSS 0.092043f
C16655 DVSS.n5352 VSS 0.092043f
C16656 DVSS.n5353 VSS 0.092043f
C16657 DVSS.n5354 VSS 0.092043f
C16658 DVSS.n5355 VSS 0.092043f
C16659 DVSS.n5356 VSS 0.092043f
C16660 DVSS.n5357 VSS 0.092043f
C16661 DVSS.n5358 VSS 0.092043f
C16662 DVSS.n5359 VSS 0.092043f
C16663 DVSS.n5360 VSS 0.092043f
C16664 DVSS.n5361 VSS 0.092043f
C16665 DVSS.n5362 VSS 0.092043f
C16666 DVSS.n5363 VSS 0.092043f
C16667 DVSS.n5364 VSS 0.092043f
C16668 DVSS.n5365 VSS 0.092043f
C16669 DVSS.n5366 VSS 0.092043f
C16670 DVSS.n5367 VSS 0.092043f
C16671 DVSS.n5368 VSS 0.092043f
C16672 DVSS.n5369 VSS 0.092043f
C16673 DVSS.n5370 VSS 0.092043f
C16674 DVSS.n5371 VSS 0.092043f
C16675 DVSS.n5372 VSS 0.092043f
C16676 DVSS.n5373 VSS 0.092043f
C16677 DVSS.n5374 VSS 0.092043f
C16678 DVSS.n5375 VSS 0.092043f
C16679 DVSS.n5376 VSS 0.092043f
C16680 DVSS.n5377 VSS 0.092043f
C16681 DVSS.n5378 VSS 0.092043f
C16682 DVSS.n5379 VSS 0.092043f
C16683 DVSS.n5380 VSS 0.092043f
C16684 DVSS.n5381 VSS 0.092043f
C16685 DVSS.n5382 VSS 0.092043f
C16686 DVSS.n5383 VSS 0.092043f
C16687 DVSS.n5384 VSS 0.092043f
C16688 DVSS.n5385 VSS 0.092043f
C16689 DVSS.n5386 VSS 0.092043f
C16690 DVSS.n5387 VSS 0.092043f
C16691 DVSS.n5388 VSS 0.092043f
C16692 DVSS.n5389 VSS 0.092043f
C16693 DVSS.n5390 VSS 0.092043f
C16694 DVSS.n5391 VSS 0.092043f
C16695 DVSS.n5392 VSS 0.092043f
C16696 DVSS.n5393 VSS 0.092043f
C16697 DVSS.n5394 VSS 0.092043f
C16698 DVSS.n5395 VSS 0.092043f
C16699 DVSS.n5396 VSS 0.092043f
C16700 DVSS.n5397 VSS 0.092043f
C16701 DVSS.n5398 VSS 0.092043f
C16702 DVSS.n5399 VSS 0.092043f
C16703 DVSS.n5400 VSS 0.092043f
C16704 DVSS.n5401 VSS 0.092043f
C16705 DVSS.n5402 VSS 0.092043f
C16706 DVSS.n5403 VSS 0.092043f
C16707 DVSS.n5404 VSS 0.092043f
C16708 DVSS.n5405 VSS 0.092043f
C16709 DVSS.n5406 VSS 0.092043f
C16710 DVSS.n5407 VSS 0.092043f
C16711 DVSS.n5408 VSS 0.092043f
C16712 DVSS.n5409 VSS 0.092043f
C16713 DVSS.n5410 VSS 0.092043f
C16714 DVSS.n5411 VSS 0.092043f
C16715 DVSS.n5412 VSS 0.092043f
C16716 DVSS.n5413 VSS 0.092043f
C16717 DVSS.n5414 VSS 0.092043f
C16718 DVSS.n5415 VSS 0.092043f
C16719 DVSS.n5416 VSS 0.092043f
C16720 DVSS.n5417 VSS 0.092043f
C16721 DVSS.n5418 VSS 0.092043f
C16722 DVSS.n5419 VSS 0.092043f
C16723 DVSS.n5420 VSS 0.092043f
C16724 DVSS.n5421 VSS 0.092043f
C16725 DVSS.n5422 VSS 0.092043f
C16726 DVSS.n5423 VSS 0.092043f
C16727 DVSS.n5424 VSS 0.092043f
C16728 DVSS.n5425 VSS 0.092043f
C16729 DVSS.n5426 VSS 0.092043f
C16730 DVSS.n5427 VSS 0.092043f
C16731 DVSS.n5428 VSS 0.092043f
C16732 DVSS.n5429 VSS 0.092043f
C16733 DVSS.n5430 VSS 0.092043f
C16734 DVSS.n5431 VSS 0.092043f
C16735 DVSS.n5432 VSS 0.092043f
C16736 DVSS.n5433 VSS 0.092043f
C16737 DVSS.n5434 VSS 0.092043f
C16738 DVSS.n5435 VSS 0.092043f
C16739 DVSS.n5436 VSS 0.092043f
C16740 DVSS.n5437 VSS 0.092043f
C16741 DVSS.n5438 VSS 0.092043f
C16742 DVSS.n5439 VSS 0.092043f
C16743 DVSS.n5440 VSS 0.092043f
C16744 DVSS.n5441 VSS 0.092043f
C16745 DVSS.n5442 VSS 0.092043f
C16746 DVSS.n5443 VSS 0.092043f
C16747 DVSS.n5444 VSS 0.092043f
C16748 DVSS.n5445 VSS 0.092043f
C16749 DVSS.n5446 VSS 0.092043f
C16750 DVSS.n5447 VSS 0.092043f
C16751 DVSS.n5448 VSS 0.092043f
C16752 DVSS.n5449 VSS 0.092043f
C16753 DVSS.n5450 VSS 0.092043f
C16754 DVSS.n5451 VSS 0.092043f
C16755 DVSS.n5452 VSS 0.092043f
C16756 DVSS.n5453 VSS 0.092043f
C16757 DVSS.n5454 VSS 0.092043f
C16758 DVSS.n5455 VSS 0.092043f
C16759 DVSS.n5456 VSS 0.092043f
C16760 DVSS.n5457 VSS 0.092043f
C16761 DVSS.n5458 VSS 0.092043f
C16762 DVSS.n5459 VSS 0.092043f
C16763 DVSS.n5460 VSS 0.092043f
C16764 DVSS.n5461 VSS 0.092043f
C16765 DVSS.n5462 VSS 0.092043f
C16766 DVSS.n5463 VSS 0.092043f
C16767 DVSS.n5464 VSS 0.092043f
C16768 DVSS.n5465 VSS 0.092043f
C16769 DVSS.n5466 VSS 0.092043f
C16770 DVSS.n5467 VSS 0.092043f
C16771 DVSS.n5468 VSS 0.092043f
C16772 DVSS.n5469 VSS 0.092043f
C16773 DVSS.n5470 VSS 0.092043f
C16774 DVSS.n5471 VSS 0.092043f
C16775 DVSS.n5472 VSS 0.092043f
C16776 DVSS.n5473 VSS 0.092043f
C16777 DVSS.n5474 VSS 0.092043f
C16778 DVSS.n5475 VSS 0.092043f
C16779 DVSS.n5476 VSS 0.092043f
C16780 DVSS.n5477 VSS 0.092043f
C16781 DVSS.n5478 VSS 0.092043f
C16782 DVSS.n5479 VSS 0.092043f
C16783 DVSS.n5480 VSS 0.092043f
C16784 DVSS.n5481 VSS 0.092043f
C16785 DVSS.n5482 VSS 0.092043f
C16786 DVSS.n5483 VSS 0.092043f
C16787 DVSS.n5484 VSS 0.092043f
C16788 DVSS.n5485 VSS 0.092043f
C16789 DVSS.n5486 VSS 0.092043f
C16790 DVSS.n5487 VSS 0.092043f
C16791 DVSS.n5488 VSS 0.092043f
C16792 DVSS.n5489 VSS 0.092043f
C16793 DVSS.n5490 VSS 0.092043f
C16794 DVSS.n5491 VSS 0.092043f
C16795 DVSS.n5492 VSS 0.092043f
C16796 DVSS.n5493 VSS 0.092043f
C16797 DVSS.n5494 VSS 0.092043f
C16798 DVSS.n5495 VSS 0.092043f
C16799 DVSS.n5496 VSS 0.092043f
C16800 DVSS.n5497 VSS 0.092043f
C16801 DVSS.n5498 VSS 0.092043f
C16802 DVSS.n5499 VSS 0.092043f
C16803 DVSS.n5500 VSS 0.092043f
C16804 DVSS.n5501 VSS 0.092043f
C16805 DVSS.n5502 VSS 0.092043f
C16806 DVSS.n5503 VSS 0.092043f
C16807 DVSS.n5504 VSS 0.092043f
C16808 DVSS.n5505 VSS 0.092043f
C16809 DVSS.n5506 VSS 0.092043f
C16810 DVSS.n5507 VSS 0.092043f
C16811 DVSS.n5508 VSS 0.092043f
C16812 DVSS.n5509 VSS 0.092043f
C16813 DVSS.n5510 VSS 0.092043f
C16814 DVSS.n5511 VSS 0.092043f
C16815 DVSS.n5512 VSS 0.092043f
C16816 DVSS.n5513 VSS 0.092043f
C16817 DVSS.n5514 VSS 0.092043f
C16818 DVSS.n5515 VSS 0.092043f
C16819 DVSS.n5516 VSS 0.092043f
C16820 DVSS.n5517 VSS 0.092043f
C16821 DVSS.n5518 VSS 0.092043f
C16822 DVSS.n5519 VSS 0.092043f
C16823 DVSS.n5520 VSS 0.092043f
C16824 DVSS.n5521 VSS 0.092043f
C16825 DVSS.n5522 VSS 0.092043f
C16826 DVSS.n5523 VSS 0.092043f
C16827 DVSS.n5524 VSS 0.092043f
C16828 DVSS.n5525 VSS 0.092043f
C16829 DVSS.n5526 VSS 0.092043f
C16830 DVSS.n5527 VSS 0.092043f
C16831 DVSS.n5528 VSS 0.092043f
C16832 DVSS.n5529 VSS 0.092043f
C16833 DVSS.n5530 VSS 0.092043f
C16834 DVSS.n5531 VSS 0.082968f
C16835 DVSS.n5532 VSS 0.082968f
C16836 DVSS.n5533 VSS 0.082968f
C16837 DVSS.n5534 VSS 0.010371f
C16838 DVSS.n5535 VSS 0.121165f
C16839 DVSS.n5536 VSS 0.046022f
C16840 DVSS.n5537 VSS 0.009075f
C16841 DVSS.n5538 VSS 0.135809f
C16842 DVSS.n5539 VSS 0.107483f
C16843 DVSS.n5540 VSS 0.007166f
C16844 DVSS.n5541 VSS 0.025334f
C16845 DVSS.n5542 VSS 0.007166f
C16846 DVSS.n5543 VSS 0.025334f
C16847 DVSS.n5544 VSS 0.250016f
C16848 DVSS.n5545 VSS 0.122809f
C16849 DVSS.n5546 VSS 0.355436f
C16850 DVSS.n5547 VSS 0.737113f
C16851 DVSS.n5548 VSS 0.194457f
C16852 DVSS.n5549 VSS 0.197235f
C16853 DVSS.n5550 VSS 0.118063f
C16854 DVSS.n5551 VSS 0.17779f
C16855 DVSS.n5552 VSS 0.197235f
C16856 DVSS.n5553 VSS 0.197235f
C16857 DVSS.n5554 VSS 0.197235f
C16858 DVSS.n5555 VSS 0.197235f
C16859 DVSS.n5556 VSS 0.197235f
C16860 DVSS.n5557 VSS 0.197235f
C16861 DVSS.n5558 VSS 0.197235f
C16862 DVSS.n5559 VSS 0.197235f
C16863 DVSS.n5560 VSS 0.197235f
C16864 DVSS.n5561 VSS 0.197235f
C16865 DVSS.n5562 VSS 0.197235f
C16866 DVSS.n5563 VSS 0.197235f
C16867 DVSS.n5564 VSS 0.197235f
C16868 DVSS.n5565 VSS 0.197235f
C16869 DVSS.n5566 VSS 0.180567f
C16870 DVSS.n5567 VSS 0.180567f
C16871 DVSS.n5568 VSS 0.237516f
C16872 DVSS.n5569 VSS 0.115285f
C16873 DVSS.n5570 VSS 0.115285f
C16874 DVSS.n5571 VSS 0.197235f
C16875 DVSS.n5572 VSS 0.197235f
C16876 DVSS.n5573 VSS 0.197235f
C16877 DVSS.n5574 VSS 0.197235f
C16878 DVSS.n5575 VSS 0.197235f
C16879 DVSS.n5576 VSS 0.197235f
C16880 DVSS.n5577 VSS 0.197235f
C16881 DVSS.n5578 VSS 0.197235f
C16882 DVSS.n5579 VSS 0.197235f
C16883 DVSS.n5580 VSS 0.197235f
C16884 DVSS.n5581 VSS 0.197235f
C16885 DVSS.n5582 VSS 0.197235f
C16886 DVSS.n5583 VSS 0.197235f
C16887 DVSS.n5584 VSS 0.197235f
C16888 DVSS.n5585 VSS 0.197235f
C16889 DVSS.n5586 VSS 0.197235f
C16890 DVSS.n5587 VSS 0.197235f
C16891 DVSS.n5588 VSS 0.197235f
C16892 DVSS.n5589 VSS 0.197235f
C16893 DVSS.n5590 VSS 0.197235f
C16894 DVSS.n5591 VSS 0.197235f
C16895 DVSS.n5592 VSS 0.197235f
C16896 DVSS.n5593 VSS 0.197235f
C16897 DVSS.n5594 VSS 0.197235f
C16898 DVSS.n5595 VSS 0.197235f
C16899 DVSS.n5596 VSS 0.197235f
C16900 DVSS.n5597 VSS 0.197235f
C16901 DVSS.n5598 VSS 0.178484f
C16902 DVSS.n5599 VSS 0.485035f
C16903 DVSS.n5600 VSS 0.48809f
C16904 DVSS.n5601 VSS 0.144307f
C16905 DVSS.n5602 VSS 0.178484f
C16906 DVSS.n5603 VSS 0.197235f
C16907 DVSS.n5604 VSS 0.197235f
C16908 DVSS.n5605 VSS 0.197235f
C16909 DVSS.n5606 VSS 0.197235f
C16910 DVSS.n5607 VSS 0.197235f
C16911 DVSS.n5608 VSS 0.197235f
C16912 DVSS.n5609 VSS 0.197235f
C16913 DVSS.n5610 VSS 0.197235f
C16914 DVSS.n5611 VSS 0.197235f
C16915 DVSS.n5612 VSS 0.197235f
C16916 DVSS.n5613 VSS 0.197235f
C16917 DVSS.n5614 VSS 0.197235f
C16918 DVSS.n5615 VSS 0.197235f
C16919 DVSS.n5616 VSS 0.197235f
C16920 DVSS.n5617 VSS 0.197235f
C16921 DVSS.n5618 VSS 0.197235f
C16922 DVSS.n5619 VSS 0.197235f
C16923 DVSS.n5620 VSS 0.197235f
C16924 DVSS.n5621 VSS 0.197235f
C16925 DVSS.n5622 VSS 0.197235f
C16926 DVSS.n5623 VSS 0.197235f
C16927 DVSS.n5624 VSS 0.197235f
C16928 DVSS.n5625 VSS 0.197235f
C16929 DVSS.n5626 VSS 0.197235f
C16930 DVSS.n5627 VSS 0.197235f
C16931 DVSS.n5628 VSS 0.197235f
C16932 DVSS.n5629 VSS 0.197235f
C16933 DVSS.n5630 VSS 0.197235f
C16934 DVSS.n5631 VSS 0.197235f
C16935 DVSS.n5632 VSS 0.197235f
C16936 DVSS.n5633 VSS 0.197235f
C16937 DVSS.n5634 VSS 0.197235f
C16938 DVSS.n5635 VSS 0.197235f
C16939 DVSS.n5636 VSS 0.197235f
C16940 DVSS.n5637 VSS 0.197235f
C16941 DVSS.n5638 VSS 0.197235f
C16942 DVSS.n5639 VSS 0.197235f
C16943 DVSS.n5640 VSS 0.197235f
C16944 DVSS.n5641 VSS 0.197235f
C16945 DVSS.n5642 VSS 0.197235f
C16946 DVSS.n5643 VSS 0.197235f
C16947 DVSS.n5644 VSS 0.197235f
C16948 DVSS.n5645 VSS 0.197235f
C16949 DVSS.n5646 VSS 0.197235f
C16950 DVSS.n5647 VSS 0.197235f
C16951 DVSS.n5648 VSS 0.175012f
C16952 DVSS.n5649 VSS 0.175012f
C16953 DVSS.n5650 VSS 0.376414f
C16954 DVSS.n5651 VSS 0.237516f
C16955 DVSS.n5652 VSS 0.120841f
C16956 DVSS.n5653 VSS 0.120841f
C16957 DVSS.n5654 VSS 0.237516f
C16958 DVSS.n5655 VSS 0.175012f
C16959 DVSS.n5656 VSS 0.197235f
C16960 DVSS.n5657 VSS 0.197235f
C16961 DVSS.n5658 VSS 0.197235f
C16962 DVSS.n5659 VSS 0.197235f
C16963 DVSS.n5660 VSS 0.117369f
C16964 DVSS.n5661 VSS 0.197235f
C16965 DVSS.n5662 VSS 0.197235f
C16966 DVSS.n5663 VSS 0.197235f
C16967 DVSS.n5664 VSS 0.197235f
C16968 DVSS.n5665 VSS 0.197235f
C16969 DVSS.n5666 VSS 0.197235f
C16970 DVSS.n5667 VSS 0.178484f
C16971 DVSS.n5668 VSS 0.197235f
C16972 DVSS.n5669 VSS 0.197235f
C16973 DVSS.n5670 VSS 0.197235f
C16974 DVSS.n5671 VSS 0.197235f
C16975 DVSS.n5672 VSS 0.197235f
C16976 DVSS.n5673 VSS 0.197235f
C16977 DVSS.n5674 VSS 0.197235f
C16978 DVSS.n5675 VSS 0.197235f
C16979 DVSS.n5676 VSS 0.197235f
C16980 DVSS.n5677 VSS 0.197235f
C16981 DVSS.n5678 VSS 0.197235f
C16982 DVSS.n5679 VSS 0.197235f
C16983 DVSS.n5680 VSS 0.197235f
C16984 DVSS.n5681 VSS 0.197235f
C16985 DVSS.n5682 VSS 0.197235f
C16986 DVSS.n5683 VSS 0.197235f
C16987 DVSS.n5684 VSS 0.197235f
C16988 DVSS.n5685 VSS 0.197235f
C16989 DVSS.n5686 VSS 0.197235f
C16990 DVSS.n5687 VSS 0.197235f
C16991 DVSS.n5688 VSS 0.197235f
C16992 DVSS.n5689 VSS 0.197235f
C16993 DVSS.n5690 VSS 0.197235f
C16994 DVSS.n5691 VSS 0.197235f
C16995 DVSS.n5692 VSS 0.197235f
C16996 DVSS.n5693 VSS 0.197235f
C16997 DVSS.n5694 VSS 0.197235f
C16998 DVSS.n5695 VSS 0.197235f
C16999 DVSS.n5696 VSS 0.197235f
C17000 DVSS.n5697 VSS 0.197235f
C17001 DVSS.n5698 VSS 0.197235f
C17002 DVSS.n5699 VSS 0.197235f
C17003 DVSS.n5700 VSS 0.125703f
C17004 DVSS.n5701 VSS 0.098618f
C17005 DVSS.n5702 VSS 0.011511f
C17006 DVSS.n5703 VSS 0.021629f
C17007 DVSS.n5704 VSS 0.022558f
C17008 DVSS.n5705 VSS 0.090209f
C17009 DVSS.n5706 VSS 0.80403f
C17010 DVSS.n5707 VSS 0.649156f
C17011 DVSS.n5708 VSS 1.22973f
C17012 DVSS.n5709 VSS 1.04375f
C17013 DVSS.t78 VSS 4.69246f
C17014 DVSS.t195 VSS 5.17029f
C17015 DVSS.t60 VSS 5.17029f
C17016 DVSS.t25 VSS 5.94999f
C17017 DVSS.n5710 VSS 5.90508f
C17018 DVSS.n5711 VSS 0.025749f
C17019 DVSS.n5712 VSS 0.032809f
C17020 DVSS.n5713 VSS 0.034262f
C17021 DVSS.n5714 VSS 0.013368f
C17022 DVSS.n5715 VSS 0.002971f
C17023 DVSS.n5716 VSS 0.098618f
C17024 DVSS.n5717 VSS 0.17015f
C17025 DVSS.n5718 VSS 0.197235f
C17026 DVSS.n5719 VSS 0.197235f
C17027 DVSS.n5720 VSS 0.197235f
C17028 DVSS.n5721 VSS 0.197235f
C17029 DVSS.n5722 VSS 0.197235f
C17030 DVSS.n5723 VSS 0.115285f
C17031 DVSS.n5724 VSS 0.072227f
C17032 DVSS.n5725 VSS 0.376414f
C17033 DVSS.n5726 VSS 0.180567f
C17034 DVSS.n5727 VSS 0.197235f
C17035 DVSS.n5728 VSS 0.197235f
C17036 DVSS.n5729 VSS 0.197235f
C17037 DVSS.n5730 VSS 0.197235f
C17038 DVSS.n5731 VSS 0.197235f
C17039 DVSS.n5732 VSS 0.197235f
C17040 DVSS.n5733 VSS 0.197235f
C17041 DVSS.n5734 VSS 0.197235f
C17042 DVSS.n5735 VSS 0.197235f
C17043 DVSS.n5736 VSS 0.197235f
C17044 DVSS.n5737 VSS 0.197235f
C17045 DVSS.n5738 VSS 0.197235f
C17046 DVSS.n5739 VSS 0.197235f
C17047 DVSS.n5740 VSS 0.127092f
C17048 DVSS.n5741 VSS 0.197235f
C17049 DVSS.n5742 VSS 0.149315f
C17050 DVSS.n5743 VSS 0.197235f
C17051 DVSS.n5744 VSS 0.197235f
C17052 DVSS.n5745 VSS 0.197235f
C17053 DVSS.n5746 VSS 0.197235f
C17054 DVSS.n5747 VSS 0.197235f
C17055 DVSS.n5748 VSS 0.197235f
C17056 DVSS.n5749 VSS 0.197235f
C17057 DVSS.n5750 VSS 0.197235f
C17058 DVSS.n5751 VSS 0.197235f
C17059 DVSS.n5752 VSS 0.197235f
C17060 DVSS.n5753 VSS 0.197235f
C17061 DVSS.n5754 VSS 0.197235f
C17062 DVSS.n5755 VSS 0.197235f
C17063 DVSS.n5756 VSS 0.197235f
C17064 DVSS.n5757 VSS 0.197235f
C17065 DVSS.n5758 VSS 0.180567f
C17066 DVSS.n5759 VSS 0.180567f
C17067 DVSS.n5760 VSS 0.376414f
C17068 DVSS.n5761 VSS 0.237516f
C17069 DVSS.n5762 VSS 0.180567f
C17070 DVSS.n5763 VSS 0.180567f
C17071 DVSS.n5764 VSS 0.180567f
C17072 DVSS.n5765 VSS 0.197235f
C17073 DVSS.n5766 VSS 0.197235f
C17074 DVSS.n5767 VSS 0.197235f
C17075 DVSS.n5768 VSS 0.197235f
C17076 DVSS.n5769 VSS 0.197235f
C17077 DVSS.n5770 VSS 0.197235f
C17078 DVSS.n5771 VSS 0.197235f
C17079 DVSS.n5772 VSS 0.197235f
C17080 DVSS.n5773 VSS 0.197235f
C17081 DVSS.n5774 VSS 0.197235f
C17082 DVSS.n5775 VSS 0.197235f
C17083 DVSS.n5776 VSS 0.197235f
C17084 DVSS.n5777 VSS 0.197235f
C17085 DVSS.n5778 VSS 0.197235f
C17086 DVSS.n5779 VSS 0.197235f
C17087 DVSS.n5780 VSS 0.197235f
C17088 DVSS.n5781 VSS 0.197235f
C17089 DVSS.n5782 VSS 0.193068f
C17090 DVSS.n5783 VSS 0.193068f
C17091 DVSS.n5784 VSS 0.197235f
C17092 DVSS.n5785 VSS 0.116674f
C17093 DVSS.n5786 VSS 0.102785f
C17094 DVSS.n5787 VSS 0.102785f
C17095 DVSS.n5788 VSS 0.197235f
C17096 DVSS.n5789 VSS 0.197235f
C17097 DVSS.n5790 VSS 0.197235f
C17098 DVSS.n5791 VSS 0.737113f
C17099 DVSS.n5792 VSS 0.359898f
C17100 DVSS.n5793 VSS 0.569501f
C17101 DVSS.n5794 VSS 0.007166f
C17102 DVSS.n5795 VSS 0.099549f
C17103 DVSS.n5796 VSS 0.250016f
C17104 DVSS.n5797 VSS 0.122809f
C17105 DVSS.n5798 VSS 0.355436f
C17106 DVSS.n5799 VSS 0.737113f
C17107 DVSS.n5800 VSS 0.146537f
C17108 DVSS.n5801 VSS 0.168761f
C17109 GF_NI_IN_C_BASE_0.pdrive_y_<1>.t3 VSS 4.07002f
C17110 GF_NI_IN_C_BASE_0.pdrive_y_<1>.n0 VSS 2.16219f
C17111 GF_NI_IN_C_BASE_0.pdrive_y_<1>.t0 VSS 0.90553f
C17112 GF_NI_IN_C_BASE_0.pdrive_y_<1>.t2 VSS 0.905248f
C17113 GF_NI_IN_C_BASE_0.pdrive_y_<1>.t1 VSS 0.134451f
C17114 GF_NI_IN_C_BASE_0.pdrive_y_<1>.t4 VSS 6.29957f
C17115 GF_NI_IN_C_BASE_0.pdrive_x_<1>.t1 VSS 2.30771f
C17116 GF_NI_IN_C_BASE_0.pdrive_x_<1>.t3 VSS 3.87089f
C17117 GF_NI_IN_C_BASE_0.pdrive_x_<1>.n0 VSS 1.83972f
C17118 GF_NI_IN_C_BASE_0.pdrive_x_<1>.t0 VSS 0.782923f
C17119 GF_NI_IN_C_BASE_0.pdrive_x_<1>.t2 VSS 0.132551f
C17120 GF_NI_IN_C_BASE_0.pdrive_x_<1>.t5 VSS 5.83096f
C17121 GF_NI_IN_C_BASE_0.pdrive_x_<1>.t4 VSS 5.94093f
C17122 GF_NI_IN_C_BASE_0.pdrive_x_<1>.n1 VSS 32.1564f
C17123 GF_NI_IN_C_BASE_0.comp018green_out_predrv_0.SLB.n0 VSS 4.47641f
C17124 GF_NI_IN_C_BASE_0.comp018green_out_predrv_0.SLB.t1 VSS 2.03366f
C17125 GF_NI_IN_C_BASE_0.comp018green_out_predrv_0.SLB.t0 VSS 0.742022f
C17126 GF_NI_IN_C_BASE_0.comp018green_out_predrv_0.SLB.t6 VSS 0.975903f
C17127 GF_NI_IN_C_BASE_0.comp018green_out_predrv_0.SLB.t3 VSS 1.12317f
C17128 GF_NI_IN_C_BASE_0.comp018green_out_predrv_0.SLB.n1 VSS 1.10814f
C17129 GF_NI_IN_C_BASE_0.comp018green_out_predrv_0.SLB.t8 VSS 0.975903f
C17130 GF_NI_IN_C_BASE_0.comp018green_out_predrv_0.SLB.t2 VSS 1.12317f
C17131 GF_NI_IN_C_BASE_0.comp018green_out_predrv_0.SLB.n2 VSS 1.10814f
C17132 GF_NI_IN_C_BASE_0.comp018green_out_predrv_0.SLB.n3 VSS 2.87718f
C17133 GF_NI_IN_C_BASE_0.comp018green_out_predrv_0.SLB.t9 VSS 0.975903f
C17134 GF_NI_IN_C_BASE_0.comp018green_out_predrv_0.SLB.t7 VSS 1.12317f
C17135 GF_NI_IN_C_BASE_0.comp018green_out_predrv_0.SLB.n4 VSS 1.10814f
C17136 GF_NI_IN_C_BASE_0.comp018green_out_predrv_0.SLB.t4 VSS 0.975903f
C17137 GF_NI_IN_C_BASE_0.comp018green_out_predrv_0.SLB.t5 VSS 1.12317f
C17138 GF_NI_IN_C_BASE_0.comp018green_out_predrv_0.SLB.n5 VSS 1.10814f
C17139 GF_NI_IN_C_BASE_0.comp018green_out_predrv_1.ENB.t1 VSS 0.239584f
C17140 GF_NI_IN_C_BASE_0.comp018green_out_predrv_1.ENB.t0 VSS 0.830038f
C17141 GF_NI_IN_C_BASE_0.comp018green_out_predrv_1.ENB.t2 VSS 0.825677f
C17142 GF_NI_IN_C_BASE_0.comp018green_out_predrv_1.ENB.t3 VSS 1.67106f
C17143 DVDD.n0 VSS 0.251684f
C17144 DVDD.n1 VSS 0.279212f
C17145 DVDD.n2 VSS 0.279212f
C17146 DVDD.n3 VSS 0.279212f
C17147 DVDD.n4 VSS 0.279212f
C17148 DVDD.n5 VSS 0.279212f
C17149 DVDD.n6 VSS 0.279212f
C17150 DVDD.n7 VSS 0.139606f
C17151 DVDD.n8 VSS 0.02361f
C17152 DVDD.n9 VSS 0.02361f
C17153 DVDD.n10 VSS 0.02361f
C17154 DVDD.n11 VSS 0.02361f
C17155 DVDD.n12 VSS 0.02361f
C17156 DVDD.n13 VSS 0.02361f
C17157 DVDD.n14 VSS 0.02361f
C17158 DVDD.n15 VSS 0.02361f
C17159 DVDD.n16 VSS 0.02361f
C17160 DVDD.n17 VSS 0.02361f
C17161 DVDD.n18 VSS 0.02361f
C17162 DVDD.n19 VSS 0.02361f
C17163 DVDD.n20 VSS 0.02361f
C17164 DVDD.n21 VSS 0.02361f
C17165 DVDD.n22 VSS 0.02361f
C17166 DVDD.n23 VSS 0.02361f
C17167 DVDD.n24 VSS 0.02361f
C17168 DVDD.n25 VSS 0.02361f
C17169 DVDD.n26 VSS 0.02361f
C17170 DVDD.n27 VSS 0.02361f
C17171 DVDD.n28 VSS 0.024841f
C17172 DVDD.n29 VSS 0.139606f
C17173 DVDD.n30 VSS 0.026275f
C17174 DVDD.n31 VSS 0.139606f
C17175 DVDD.n32 VSS 0.166151f
C17176 DVDD.n33 VSS 0.255617f
C17177 DVDD.n34 VSS 0.336235f
C17178 DVDD.n35 VSS 0.532863f
C17179 DVDD.n36 VSS 0.279212f
C17180 DVDD.n37 VSS 0.279212f
C17181 DVDD.n38 VSS 0.532863f
C17182 DVDD.n39 VSS 0.279212f
C17183 DVDD.n40 VSS 0.336235f
C17184 DVDD.n41 VSS 0.336235f
C17185 DVDD.n42 VSS 0.163202f
C17186 DVDD.n43 VSS 0.139606f
C17187 DVDD.n44 VSS 0.532863f
C17188 DVDD.n45 VSS 0.255617f
C17189 DVDD.n46 VSS 0.279212f
C17190 DVDD.n47 VSS 0.279212f
C17191 DVDD.n48 VSS 0.012947f
C17192 DVDD.n49 VSS 0.007235f
C17193 DVDD.n50 VSS 0.023609f
C17194 DVDD.n51 VSS 0.017135f
C17195 DVDD.n52 VSS 0.010281f
C17196 DVDD.n53 VSS 0.003427f
C17197 DVDD.n54 VSS 0.020182f
C17198 DVDD.n55 VSS 0.013327f
C17199 DVDD.n56 VSS 0.006473f
C17200 DVDD.n57 VSS 0.023228f
C17201 DVDD.n58 VSS 0.17205f
C17202 DVDD.n59 VSS 0.019801f
C17203 DVDD.n60 VSS 0.003046f
C17204 DVDD.n61 VSS 0.0099f
C17205 DVDD.n62 VSS 0.016755f
C17206 DVDD.n63 VSS 0.023609f
C17207 DVDD.n64 VSS 0.006854f
C17208 DVDD.n65 VSS 0.013708f
C17209 DVDD.n66 VSS 0.020563f
C17210 DVDD.n67 VSS 0.003807f
C17211 DVDD.n68 VSS 0.010662f
C17212 DVDD.n69 VSS 0.008187f
C17213 DVDD.n70 VSS 0.011614f
C17214 DVDD.n71 VSS 0.026085f
C17215 DVDD.n72 VSS 0.070464f
C17216 DVDD.n73 VSS 0.070464f
C17217 DVDD.n74 VSS 0.02361f
C17218 DVDD.n75 VSS 0.045744f
C17219 DVDD.n76 VSS 0.101264f
C17220 DVDD.n77 VSS 0.101264f
C17221 DVDD.n78 VSS 0.015422f
C17222 DVDD.n79 VSS 0.101264f
C17223 DVDD.n80 VSS 0.166151f
C17224 DVDD.n81 VSS 0.016565f
C17225 DVDD.n82 VSS 0.139606f
C17226 DVDD.n83 VSS 0.027037f
C17227 DVDD.n84 VSS 0.018659f
C17228 DVDD.n85 VSS 0.035231f
C17229 DVDD.n86 VSS 0.059951f
C17230 DVDD.n88 VSS 0.017929f
C17231 DVDD.n89 VSS 0.018056f
C17232 DVDD.n90 VSS 0.015894f
C17233 DVDD.n91 VSS 0.018056f
C17234 DVDD.n92 VSS 0.018056f
C17235 DVDD.n93 VSS 0.018056f
C17236 DVDD.n94 VSS 0.018056f
C17237 DVDD.n95 VSS 0.018056f
C17238 DVDD.n96 VSS 0.018056f
C17239 DVDD.n97 VSS 0.018056f
C17240 DVDD.n98 VSS 0.017929f
C17241 DVDD.n99 VSS 0.018056f
C17242 DVDD.n100 VSS 0.020726f
C17243 DVDD.n102 VSS 0.015767f
C17244 DVDD.n103 VSS 3.87242f
C17245 DVDD.n105 VSS 0.175794f
C17246 DVDD.n107 VSS 0.057022f
C17247 DVDD.n108 VSS 0.089466f
C17248 DVDD.n109 VSS 0.015767f
C17249 DVDD.n110 VSS 0.015767f
C17250 DVDD.n111 VSS 0.015767f
C17251 DVDD.n112 VSS 0.015767f
C17252 DVDD.n113 VSS 0.015767f
C17253 DVDD.n114 VSS 0.015767f
C17254 DVDD.n115 VSS 0.279212f
C17255 DVDD.n116 VSS 0.120926f
C17256 DVDD.n117 VSS 0.279212f
C17257 DVDD.n118 VSS 0.279212f
C17258 DVDD.n119 VSS 0.336235f
C17259 DVDD.n120 VSS 0.279212f
C17260 DVDD.n121 VSS 0.279212f
C17261 DVDD.n122 VSS 0.279212f
C17262 DVDD.n123 VSS 0.279212f
C17263 DVDD.n124 VSS 0.279212f
C17264 DVDD.n125 VSS 0.279212f
C17265 DVDD.n126 VSS 0.279212f
C17266 DVDD.n127 VSS 0.279212f
C17267 DVDD.n128 VSS 0.279212f
C17268 DVDD.n129 VSS 0.279212f
C17269 DVDD.n130 VSS 0.139606f
C17270 DVDD.n131 VSS 0.279212f
C17271 DVDD.n132 VSS 0.279212f
C17272 DVDD.n133 VSS 0.279212f
C17273 DVDD.n134 VSS 0.279212f
C17274 DVDD.n135 VSS 0.017764f
C17275 DVDD.n136 VSS 0.009915f
C17276 DVDD.n137 VSS 0.139606f
C17277 DVDD.n138 VSS 0.009915f
C17278 DVDD.n139 VSS 0.019831f
C17279 DVDD.n140 VSS 0.009915f
C17280 DVDD.n141 VSS 0.019831f
C17281 DVDD.n142 VSS 0.011355f
C17282 DVDD.n143 VSS 0.139606f
C17283 DVDD.n144 VSS 0.139606f
C17284 DVDD.n145 VSS 0.009915f
C17285 DVDD.n146 VSS 0.009915f
C17286 DVDD.n147 VSS 0.009915f
C17287 DVDD.n148 VSS 0.009915f
C17288 DVDD.n149 VSS 0.009915f
C17289 DVDD.n150 VSS 0.009915f
C17290 DVDD.n151 VSS 0.009915f
C17291 DVDD.n152 VSS 0.009915f
C17292 DVDD.n153 VSS 0.009915f
C17293 DVDD.n154 VSS 0.009915f
C17294 DVDD.n155 VSS 0.152387f
C17295 DVDD.n156 VSS 0.009915f
C17296 DVDD.n157 VSS 0.009915f
C17297 DVDD.n158 VSS 0.009915f
C17298 DVDD.n159 VSS 0.009915f
C17299 DVDD.n160 VSS 0.009915f
C17300 DVDD.n161 VSS 0.009915f
C17301 DVDD.n162 VSS 0.009915f
C17302 DVDD.n163 VSS 0.009915f
C17303 DVDD.n164 VSS 0.011355f
C17304 DVDD.n165 VSS -0.292745f
C17305 DVDD.n166 VSS 0.009915f
C17306 DVDD.n167 VSS 0.019831f
C17307 DVDD.n168 VSS 0.011355f
C17308 DVDD.n169 VSS 0.139606f
C17309 DVDD.n170 VSS 0.266432f
C17310 DVDD.n171 VSS 0.009915f
C17311 DVDD.n172 VSS 0.009915f
C17312 DVDD.n173 VSS 0.009915f
C17313 DVDD.n174 VSS 0.009915f
C17314 DVDD.n175 VSS 0.009915f
C17315 DVDD.n176 VSS 0.009915f
C17316 DVDD.n177 VSS 0.009915f
C17317 DVDD.n178 VSS 0.009915f
C17318 DVDD.n179 VSS 0.009915f
C17319 DVDD.n180 VSS 0.139606f
C17320 DVDD.n181 VSS 0.009915f
C17321 DVDD.n182 VSS 0.009915f
C17322 DVDD.n183 VSS 0.009915f
C17323 DVDD.n184 VSS 0.009915f
C17324 DVDD.n185 VSS 0.009915f
C17325 DVDD.n186 VSS 0.009915f
C17326 DVDD.n187 VSS 0.009915f
C17327 DVDD.n188 VSS 0.009915f
C17328 DVDD.n189 VSS 0.009915f
C17329 DVDD.n190 VSS 0.011355f
C17330 DVDD.n191 VSS 0.010555f
C17331 DVDD.n192 VSS 0.019831f
C17332 DVDD.n193 VSS 0.009915f
C17333 DVDD.n194 VSS 0.019831f
C17334 DVDD.n195 VSS 0.011355f
C17335 DVDD.n196 VSS 0.139606f
C17336 DVDD.n197 VSS 0.139606f
C17337 DVDD.n198 VSS 0.017212f
C17338 DVDD.n199 VSS 0.279212f
C17339 DVDD.n200 VSS 0.279212f
C17340 DVDD.n201 VSS 0.279212f
C17341 DVDD.n202 VSS 0.279212f
C17342 DVDD.n203 VSS 0.279212f
C17343 DVDD.n204 VSS 0.279212f
C17344 DVDD.n205 VSS 0.279212f
C17345 DVDD.n206 VSS 0.279212f
C17346 DVDD.n207 VSS 0.279212f
C17347 DVDD.n208 VSS 0.279212f
C17348 DVDD.n209 VSS 0.279212f
C17349 DVDD.n210 VSS 0.279212f
C17350 DVDD.n211 VSS 0.279212f
C17351 DVDD.n212 VSS 0.279212f
C17352 DVDD.n213 VSS 0.279212f
C17353 DVDD.n214 VSS 0.279212f
C17354 DVDD.n215 VSS 0.163202f
C17355 DVDD.n216 VSS 0.255617f
C17356 DVDD.n217 VSS 0.279212f
C17357 DVDD.n218 VSS 0.023609f
C17358 DVDD.n219 VSS 0.023609f
C17359 DVDD.n220 VSS 0.139606f
C17360 DVDD.n221 VSS 0.023609f
C17361 DVDD.n222 VSS 0.023609f
C17362 DVDD.n223 VSS 0.14022f
C17363 DVDD.n224 VSS 0.101264f
C17364 DVDD.n225 VSS 0.027036f
C17365 DVDD.n226 VSS 0.101264f
C17366 DVDD.n227 VSS 0.120926f
C17367 DVDD.n228 VSS 0.026575f
C17368 DVDD.n229 VSS 0.015767f
C17369 DVDD.n230 VSS 0.015767f
C17370 DVDD.n231 VSS 0.015767f
C17371 DVDD.n232 VSS 0.015767f
C17372 DVDD.n233 VSS 0.015767f
C17373 DVDD.n234 VSS 0.177949f
C17374 DVDD.n235 VSS 0.021998f
C17375 DVDD.n236 VSS 0.015767f
C17376 DVDD.n237 VSS 0.015767f
C17377 DVDD.n238 VSS 0.015767f
C17378 DVDD.n239 VSS 0.015767f
C17379 DVDD.n240 VSS 0.018056f
C17380 DVDD.n241 VSS 0.057022f
C17381 DVDD.n242 VSS 0.017929f
C17382 DVDD.n243 VSS 0.060711f
C17383 DVDD.n244 VSS 0.018056f
C17384 DVDD.n245 VSS 0.107987f
C17385 DVDD.n246 VSS 0.018056f
C17386 DVDD.n247 VSS 0.060711f
C17387 DVDD.n248 VSS 0.060711f
C17388 DVDD.n249 VSS 0.015894f
C17389 DVDD.n250 VSS 0.017929f
C17390 DVDD.n251 VSS 0.060711f
C17391 DVDD.n252 VSS 0.018056f
C17392 DVDD.n253 VSS 0.060711f
C17393 DVDD.n254 VSS 0.018056f
C17394 DVDD.n255 VSS 0.045533f
C17395 DVDD.n256 VSS 0.534473f
C17396 DVDD.n257 VSS 0.018056f
C17397 DVDD.n258 VSS 0.198575f
C17398 DVDD.n259 VSS 1.25266f
C17399 DVDD.t99 VSS 4.647759f
C17400 DVDD.n260 VSS 8.39546f
C17401 DVDD.n261 VSS 0.849875f
C17402 DVDD.t21 VSS 4.69202f
C17403 DVDD.n262 VSS 0.879805f
C17404 DVDD.t143 VSS 4.647759f
C17405 DVDD.n263 VSS 1.24841f
C17406 DVDD.n264 VSS 0.030071f
C17407 DVDD.n265 VSS 0.065482f
C17408 DVDD.n266 VSS -0.171235f
C17409 DVDD.n267 VSS 0.02361f
C17410 DVDD.n268 VSS 0.013899f
C17411 DVDD.n269 VSS 0.070301f
C17412 DVDD.n270 VSS 0.010662f
C17413 DVDD.n271 VSS 0.139606f
C17414 DVDD.n272 VSS 0.007235f
C17415 DVDD.n273 VSS 0.139606f
C17416 DVDD.n274 VSS 0.026085f
C17417 DVDD.n275 VSS 0.020753f
C17418 DVDD.n276 VSS 0.003998f
C17419 DVDD.n277 VSS 0.010853f
C17420 DVDD.n278 VSS 0.017707f
C17421 DVDD.n279 VSS 0.003237f
C17422 DVDD.n280 VSS 0.007806f
C17423 DVDD.n281 VSS 0.014661f
C17424 DVDD.n282 VSS 0.021515f
C17425 DVDD.n283 VSS 0.00476f
C17426 DVDD.n284 VSS 0.17205f
C17427 DVDD.n285 VSS 0.008187f
C17428 DVDD.n286 VSS 0.001332f
C17429 DVDD.n287 VSS 0.018088f
C17430 DVDD.n288 VSS 0.011233f
C17431 DVDD.n289 VSS 0.004379f
C17432 DVDD.n290 VSS 0.021134f
C17433 DVDD.n291 VSS 0.01428f
C17434 DVDD.n292 VSS 0.007425f
C17435 DVDD.n293 VSS 0.02361f
C17436 DVDD.n294 VSS 0.026085f
C17437 DVDD.n295 VSS 0.139606f
C17438 DVDD.n296 VSS 0.026039f
C17439 DVDD.n297 VSS 0.139606f
C17440 DVDD.n298 VSS 0.003807f
C17441 DVDD.n299 VSS 0.020563f
C17442 DVDD.n300 VSS 0.013708f
C17443 DVDD.n301 VSS 0.006854f
C17444 DVDD.n302 VSS 0.023609f
C17445 DVDD.n303 VSS 0.016755f
C17446 DVDD.n304 VSS 0.0099f
C17447 DVDD.n305 VSS 0.003046f
C17448 DVDD.n306 VSS 0.019801f
C17449 DVDD.n307 VSS 0.095365f
C17450 DVDD.n308 VSS 0.016374f
C17451 DVDD.n309 VSS 0.023228f
C17452 DVDD.n310 VSS 0.006473f
C17453 DVDD.n311 VSS 0.013327f
C17454 DVDD.n312 VSS 0.020182f
C17455 DVDD.n313 VSS 0.003427f
C17456 DVDD.n314 VSS 0.010281f
C17457 DVDD.n315 VSS 0.017135f
C17458 DVDD.n316 VSS 9.52e-19
C17459 DVDD.n317 VSS 0.026085f
C17460 DVDD.n318 VSS 0.070301f
C17461 DVDD.n319 VSS 0.070301f
C17462 DVDD.n320 VSS 0.070301f
C17463 DVDD.n321 VSS 0.090449f
C17464 DVDD.n322 VSS 0.139606f
C17465 DVDD.n323 VSS 0.027037f
C17466 DVDD.n324 VSS 0.090449f
C17467 DVDD.n325 VSS 0.058989f
C17468 DVDD.n326 VSS 0.02361f
C17469 DVDD.n327 VSS 0.058624f
C17470 DVDD.n328 VSS 0.129775f
C17471 DVDD.n329 VSS 0.018659f
C17472 DVDD.n330 VSS 0.070301f
C17473 DVDD.n331 VSS 0.015422f
C17474 DVDD.n332 VSS 0.045639f
C17475 DVDD.n333 VSS 0.03515f
C17476 DVDD.n334 VSS 0.017929f
C17477 DVDD.n335 VSS 0.018056f
C17478 DVDD.n336 VSS 0.018056f
C17479 DVDD.n337 VSS 0.017929f
C17480 DVDD.n338 VSS 0.018056f
C17481 DVDD.n339 VSS 0.020726f
C17482 DVDD.n341 VSS 0.020726f
C17483 DVDD.n342 VSS 0.018056f
C17484 DVDD.n343 VSS 0.018056f
C17485 DVDD.n344 VSS 0.015894f
C17486 DVDD.n345 VSS 0.018056f
C17487 DVDD.n346 VSS 0.018056f
C17488 DVDD.n347 VSS 0.018056f
C17489 DVDD.n349 VSS 0.015767f
C17490 DVDD.n350 VSS 0.175794f
C17491 DVDD.n352 VSS 0.015767f
C17492 DVDD.n353 VSS 0.058989f
C17493 DVDD.n354 VSS 0.279212f
C17494 DVDD.n355 VSS 0.279212f
C17495 DVDD.n356 VSS 0.279212f
C17496 DVDD.n357 VSS 0.186797f
C17497 DVDD.n358 VSS 0.336235f
C17498 DVDD.n359 VSS 0.532863f
C17499 DVDD.n360 VSS 0.279212f
C17500 DVDD.n361 VSS 0.232022f
C17501 DVDD.n362 VSS 0.279212f
C17502 DVDD.n363 VSS 0.279212f
C17503 DVDD.n364 VSS 0.279212f
C17504 DVDD.n365 VSS 0.279212f
C17505 DVDD.n366 VSS 0.279212f
C17506 DVDD.n367 VSS 0.279212f
C17507 DVDD.n368 VSS 0.279212f
C17508 DVDD.n369 VSS 0.279212f
C17509 DVDD.n370 VSS 0.279212f
C17510 DVDD.n371 VSS 0.279212f
C17511 DVDD.n372 VSS 0.279212f
C17512 DVDD.n373 VSS 0.279212f
C17513 DVDD.n374 VSS 0.279212f
C17514 DVDD.n375 VSS 0.279212f
C17515 DVDD.n376 VSS 0.279212f
C17516 DVDD.n377 VSS 0.017764f
C17517 DVDD.n378 VSS 0.009915f
C17518 DVDD.n379 VSS 0.139606f
C17519 DVDD.n380 VSS 0.009915f
C17520 DVDD.n381 VSS 0.005197f
C17521 DVDD.n382 VSS 0.279212f
C17522 DVDD.n383 VSS 0.279212f
C17523 DVDD.n384 VSS 0.279212f
C17524 DVDD.n385 VSS 0.279212f
C17525 DVDD.n386 VSS 0.279212f
C17526 DVDD.n387 VSS 0.279212f
C17527 DVDD.n388 VSS 0.279212f
C17528 DVDD.n389 VSS 0.279212f
C17529 DVDD.n390 VSS 0.279212f
C17530 DVDD.n391 VSS 0.279212f
C17531 DVDD.n392 VSS 0.279212f
C17532 DVDD.n393 VSS 0.279212f
C17533 DVDD.n394 VSS 0.279212f
C17534 DVDD.n395 VSS 0.279212f
C17535 DVDD.n396 VSS 0.279212f
C17536 DVDD.n397 VSS 0.279212f
C17537 DVDD.n398 VSS 0.279212f
C17538 DVDD.n399 VSS 0.178932f
C17539 DVDD.n400 VSS 0.017764f
C17540 DVDD.n401 VSS 0.009915f
C17541 DVDD.n402 VSS 0.101264f
C17542 DVDD.n403 VSS 0.009915f
C17543 DVDD.n404 VSS 0.005197f
C17544 DVDD.n405 VSS 0.274297f
C17545 DVDD.n406 VSS 0.279212f
C17546 DVDD.n407 VSS 0.336235f
C17547 DVDD.n408 VSS 0.239887f
C17548 DVDD.n409 VSS 0.279212f
C17549 DVDD.n410 VSS 0.279212f
C17550 DVDD.n411 VSS 0.279212f
C17551 DVDD.n412 VSS 0.279212f
C17552 DVDD.n413 VSS 0.279212f
C17553 DVDD.n414 VSS 0.279212f
C17554 DVDD.n415 VSS 0.279212f
C17555 DVDD.n416 VSS 0.279212f
C17556 DVDD.n417 VSS 0.279212f
C17557 DVDD.n418 VSS 0.279212f
C17558 DVDD.n419 VSS 0.279212f
C17559 DVDD.n420 VSS 0.279212f
C17560 DVDD.n421 VSS 0.279212f
C17561 DVDD.n422 VSS 0.279212f
C17562 DVDD.n423 VSS 0.279212f
C17563 DVDD.n424 VSS 0.017764f
C17564 DVDD.n425 VSS 0.009915f
C17565 DVDD.n426 VSS 0.139606f
C17566 DVDD.n427 VSS 0.009915f
C17567 DVDD.n428 VSS 0.005197f
C17568 DVDD.n429 VSS 0.279212f
C17569 DVDD.n430 VSS 0.279212f
C17570 DVDD.n431 VSS 0.279212f
C17571 DVDD.n432 VSS 0.279212f
C17572 DVDD.n433 VSS 0.279212f
C17573 DVDD.n434 VSS 0.279212f
C17574 DVDD.n435 VSS 0.279212f
C17575 DVDD.n436 VSS 0.279212f
C17576 DVDD.n437 VSS 0.279212f
C17577 DVDD.n438 VSS 0.279212f
C17578 DVDD.n439 VSS 0.279212f
C17579 DVDD.n440 VSS 0.279212f
C17580 DVDD.n441 VSS 0.279212f
C17581 DVDD.n442 VSS 0.279212f
C17582 DVDD.n443 VSS 0.279212f
C17583 DVDD.n444 VSS 0.279212f
C17584 DVDD.n445 VSS 0.279212f
C17585 DVDD.n446 VSS 0.279212f
C17586 DVDD.n447 VSS 0.171067f
C17587 DVDD.n448 VSS 0.336235f
C17588 DVDD.n449 VSS 0.108146f
C17589 DVDD.n450 VSS 0.457161f
C17590 DVDD.n451 VSS 0.171067f
C17591 DVDD.n452 VSS 0.009915f
C17592 DVDD.n453 VSS 0.009915f
C17593 DVDD.n454 VSS 0.009915f
C17594 DVDD.n455 VSS 0.009915f
C17595 DVDD.n456 VSS 0.009915f
C17596 DVDD.n457 VSS 0.009915f
C17597 DVDD.n458 VSS 0.009915f
C17598 DVDD.n459 VSS 0.009915f
C17599 DVDD.n460 VSS 0.009915f
C17600 DVDD.n461 VSS 0.009915f
C17601 DVDD.n462 VSS 0.139606f
C17602 DVDD.n463 VSS 0.009915f
C17603 DVDD.n464 VSS 0.009915f
C17604 DVDD.n465 VSS 0.009915f
C17605 DVDD.n466 VSS 0.009915f
C17606 DVDD.n467 VSS 0.009915f
C17607 DVDD.n468 VSS 0.009915f
C17608 DVDD.n469 VSS 0.009915f
C17609 DVDD.n470 VSS 0.009915f
C17610 DVDD.n471 VSS 0.009915f
C17611 DVDD.n472 VSS 0.009915f
C17612 DVDD.n473 VSS 0.011355f
C17613 DVDD.n474 VSS 0.011355f
C17614 DVDD.n475 VSS 0.279212f
C17615 DVDD.n476 VSS 0.247752f
C17616 DVDD.n477 VSS 0.532863f
C17617 DVDD.n478 VSS 0.336235f
C17618 DVDD.n479 VSS 0.279212f
C17619 DVDD.n480 VSS 0.279212f
C17620 DVDD.n481 VSS 0.336235f
C17621 DVDD.n482 VSS 0.171067f
C17622 DVDD.n483 VSS 0.247752f
C17623 DVDD.n484 VSS 0.279212f
C17624 DVDD.n485 VSS 0.108146f
C17625 DVDD.n486 VSS 0.009915f
C17626 DVDD.n487 VSS 0.009915f
C17627 DVDD.n488 VSS 0.009915f
C17628 DVDD.n489 VSS 0.009915f
C17629 DVDD.n490 VSS 0.009915f
C17630 DVDD.n491 VSS 0.009915f
C17631 DVDD.n492 VSS 0.009915f
C17632 DVDD.n493 VSS 0.009915f
C17633 DVDD.n494 VSS 0.009915f
C17634 DVDD.n495 VSS 0.009915f
C17635 DVDD.n496 VSS 0.279212f
C17636 DVDD.n497 VSS 0.279212f
C17637 DVDD.n498 VSS 0.279212f
C17638 DVDD.n499 VSS 0.279212f
C17639 DVDD.n500 VSS 0.279212f
C17640 DVDD.n501 VSS 0.279212f
C17641 DVDD.n502 VSS 0.279212f
C17642 DVDD.n503 VSS 0.279212f
C17643 DVDD.n504 VSS 0.279212f
C17644 DVDD.n505 VSS 0.279212f
C17645 DVDD.n506 VSS 0.279212f
C17646 DVDD.n507 VSS 0.279212f
C17647 DVDD.n508 VSS 0.279212f
C17648 DVDD.n509 VSS 0.279212f
C17649 DVDD.n510 VSS 0.279212f
C17650 DVDD.n511 VSS 0.279212f
C17651 DVDD.n512 VSS 0.279212f
C17652 DVDD.n513 VSS 0.279212f
C17653 DVDD.n514 VSS 0.279212f
C17654 DVDD.n515 VSS 0.279212f
C17655 DVDD.n516 VSS 0.279212f
C17656 DVDD.n517 VSS 0.279212f
C17657 DVDD.n518 VSS 0.279212f
C17658 DVDD.n519 VSS 0.279212f
C17659 DVDD.n520 VSS 0.279212f
C17660 DVDD.n521 VSS 0.279212f
C17661 DVDD.n522 VSS 0.279212f
C17662 DVDD.n523 VSS 0.279212f
C17663 DVDD.n524 VSS 0.279212f
C17664 DVDD.n525 VSS 0.279212f
C17665 DVDD.n526 VSS 0.279212f
C17666 DVDD.n527 VSS 0.279212f
C17667 DVDD.n528 VSS 0.279212f
C17668 DVDD.n529 VSS 0.279212f
C17669 DVDD.n530 VSS 0.279212f
C17670 DVDD.n531 VSS 0.279212f
C17671 DVDD.n532 VSS 0.279212f
C17672 DVDD.n533 VSS 0.279212f
C17673 DVDD.n534 VSS 0.279212f
C17674 DVDD.n535 VSS 0.279212f
C17675 DVDD.n536 VSS 0.279212f
C17676 DVDD.n537 VSS 0.152387f
C17677 DVDD.n538 VSS 0.279212f
C17678 DVDD.n539 VSS 0.279212f
C17679 DVDD.n540 VSS 0.279212f
C17680 DVDD.n541 VSS 0.279212f
C17681 DVDD.n542 VSS 0.279212f
C17682 DVDD.n543 VSS 0.279212f
C17683 DVDD.n544 VSS 0.279212f
C17684 DVDD.n545 VSS 0.279212f
C17685 DVDD.n546 VSS 0.279212f
C17686 DVDD.n547 VSS 0.279212f
C17687 DVDD.n548 VSS 0.279212f
C17688 DVDD.n549 VSS 0.279212f
C17689 DVDD.n550 VSS 0.279212f
C17690 DVDD.n551 VSS 0.279212f
C17691 DVDD.n552 VSS 0.279212f
C17692 DVDD.n553 VSS 0.279212f
C17693 DVDD.n554 VSS 0.279212f
C17694 DVDD.n555 VSS 0.215308f
C17695 DVDD.n556 VSS 0.009915f
C17696 DVDD.n557 VSS 0.009915f
C17697 DVDD.n558 VSS 0.009915f
C17698 DVDD.n559 VSS 0.009915f
C17699 DVDD.n560 VSS 0.009915f
C17700 DVDD.n561 VSS 0.009915f
C17701 DVDD.n562 VSS 0.009915f
C17702 DVDD.n563 VSS 0.009915f
C17703 DVDD.n564 VSS 0.009915f
C17704 DVDD.n565 VSS 0.009915f
C17705 DVDD.n566 VSS 0.018711f
C17706 DVDD.n567 VSS 0.010235f
C17707 DVDD.n568 VSS 0.019831f
C17708 DVDD.n569 VSS 0.011355f
C17709 DVDD.n570 VSS 0.139606f
C17710 DVDD.n571 VSS 0.260533f
C17711 DVDD.n572 VSS 0.027427f
C17712 DVDD.n573 VSS 0.009915f
C17713 DVDD.n574 VSS 0.279212f
C17714 DVDD.n575 VSS 0.279212f
C17715 DVDD.n576 VSS 0.279212f
C17716 DVDD.n577 VSS 0.279212f
C17717 DVDD.n578 VSS 0.279212f
C17718 DVDD.n579 VSS 0.279212f
C17719 DVDD.n580 VSS 0.279212f
C17720 DVDD.n581 VSS 0.279212f
C17721 DVDD.n582 VSS 0.279212f
C17722 DVDD.n583 VSS 0.279212f
C17723 DVDD.n584 VSS 0.139606f
C17724 DVDD.n585 VSS 0.279212f
C17725 DVDD.n586 VSS 0.279212f
C17726 DVDD.n587 VSS 0.279212f
C17727 DVDD.n588 VSS 0.279212f
C17728 DVDD.n589 VSS 0.027427f
C17729 DVDD.n590 VSS 0.009915f
C17730 DVDD.n591 VSS 0.139606f
C17731 DVDD.n592 VSS 0.009915f
C17732 DVDD.n593 VSS 0.017212f
C17733 DVDD.n594 VSS 0.011355f
C17734 DVDD.n595 VSS 0.019831f
C17735 DVDD.n596 VSS 0.005821f
C17736 DVDD.n597 VSS 0.011355f
C17737 DVDD.n598 VSS 0.063326f
C17738 DVDD.n599 VSS 0.011355f
C17739 DVDD.n600 VSS 0.019831f
C17740 DVDD.n601 VSS 0.019831f
C17741 DVDD.n602 VSS 0.019831f
C17742 DVDD.n603 VSS 0.139606f
C17743 DVDD.n604 VSS 0.011035f
C17744 DVDD.n605 VSS 0.140589f
C17745 DVDD.n606 VSS 0.009915f
C17746 DVDD.n607 VSS 0.009915f
C17747 DVDD.n608 VSS 0.009915f
C17748 DVDD.n609 VSS 0.009915f
C17749 DVDD.n610 VSS 0.009915f
C17750 DVDD.n611 VSS 0.009915f
C17751 DVDD.n612 VSS 0.009915f
C17752 DVDD.n613 VSS 0.009915f
C17753 DVDD.n614 VSS 0.009915f
C17754 DVDD.n615 VSS 0.009915f
C17755 DVDD.n616 VSS 0.139606f
C17756 DVDD.n617 VSS 0.009915f
C17757 DVDD.n618 VSS 0.009915f
C17758 DVDD.n619 VSS 0.009915f
C17759 DVDD.n620 VSS 0.009915f
C17760 DVDD.n621 VSS 0.009915f
C17761 DVDD.n622 VSS 0.009915f
C17762 DVDD.n623 VSS 0.009915f
C17763 DVDD.n624 VSS 0.009915f
C17764 DVDD.n625 VSS 0.009915f
C17765 DVDD.n626 VSS 0.011355f
C17766 DVDD.n627 VSS 0.019831f
C17767 DVDD.n628 VSS 0.010235f
C17768 DVDD.n629 VSS 0.019831f
C17769 DVDD.n630 VSS 0.011355f
C17770 DVDD.n631 VSS 0.019831f
C17771 DVDD.n632 VSS 0.011355f
C17772 DVDD.n633 VSS 0.019831f
C17773 DVDD.n634 VSS 0.011355f
C17774 DVDD.n635 VSS 0.019831f
C17775 DVDD.n636 VSS 0.011355f
C17776 DVDD.n637 VSS 0.019831f
C17777 DVDD.n638 VSS 0.011355f
C17778 DVDD.n639 VSS 0.019831f
C17779 DVDD.n640 VSS 0.011355f
C17780 DVDD.n641 VSS 0.019831f
C17781 DVDD.n642 VSS 0.019831f
C17782 DVDD.n643 VSS 0.010875f
C17783 DVDD.n644 VSS 0.010395f
C17784 DVDD.n645 VSS 0.019831f
C17785 DVDD.n646 VSS 0.011355f
C17786 DVDD.n647 VSS 0.019831f
C17787 DVDD.n648 VSS 0.011355f
C17788 DVDD.n649 VSS 0.019831f
C17789 DVDD.n650 VSS 0.011355f
C17790 DVDD.n651 VSS 0.019831f
C17791 DVDD.n652 VSS 0.011355f
C17792 DVDD.n653 VSS 0.019831f
C17793 DVDD.n654 VSS 0.011355f
C17794 DVDD.n655 VSS 0.019831f
C17795 DVDD.n656 VSS 0.011355f
C17796 DVDD.n657 VSS 0.019831f
C17797 DVDD.n658 VSS 0.019831f
C17798 DVDD.n659 VSS 0.010715f
C17799 DVDD.n660 VSS 0.010555f
C17800 DVDD.n661 VSS 0.019831f
C17801 DVDD.n662 VSS 0.011355f
C17802 DVDD.n663 VSS 0.019831f
C17803 DVDD.n664 VSS 0.011355f
C17804 DVDD.n665 VSS 0.019831f
C17805 DVDD.n666 VSS 0.011355f
C17806 DVDD.n667 VSS 0.019831f
C17807 DVDD.n668 VSS 0.011355f
C17808 DVDD.n669 VSS 0.019831f
C17809 DVDD.n670 VSS 0.019831f
C17810 DVDD.n671 VSS 0.019831f
C17811 DVDD.n672 VSS 0.139606f
C17812 DVDD.n673 VSS 0.011355f
C17813 DVDD.n674 VSS 0.140589f
C17814 DVDD.n675 VSS 0.009915f
C17815 DVDD.n676 VSS 0.009915f
C17816 DVDD.n677 VSS 0.009915f
C17817 DVDD.n678 VSS 0.009915f
C17818 DVDD.n679 VSS 0.009915f
C17819 DVDD.n680 VSS 0.009915f
C17820 DVDD.n681 VSS 0.009915f
C17821 DVDD.n682 VSS 0.009915f
C17822 DVDD.n683 VSS 0.009915f
C17823 DVDD.n684 VSS 0.279212f
C17824 DVDD.n685 VSS 0.279212f
C17825 DVDD.n686 VSS 0.279212f
C17826 DVDD.n687 VSS 0.279212f
C17827 DVDD.n688 VSS 0.279212f
C17828 DVDD.n689 VSS 0.279212f
C17829 DVDD.n690 VSS 0.279212f
C17830 DVDD.n691 VSS 0.279212f
C17831 DVDD.n692 VSS 0.279212f
C17832 DVDD.n693 VSS 0.279212f
C17833 DVDD.n694 VSS 0.279212f
C17834 DVDD.n695 VSS 0.100281f
C17835 DVDD.n696 VSS 0.532863f
C17836 DVDD.n697 VSS 0.532863f
C17837 DVDD.n698 VSS 0.178932f
C17838 DVDD.n699 VSS 0.336235f
C17839 DVDD.n700 VSS 0.279212f
C17840 DVDD.n701 VSS 0.279212f
C17841 DVDD.n702 VSS 0.139606f
C17842 DVDD.n703 VSS 0.274297f
C17843 DVDD.n704 VSS 0.101264f
C17844 DVDD.n705 VSS 0.009915f
C17845 DVDD.n706 VSS 0.009915f
C17846 DVDD.n707 VSS 0.009915f
C17847 DVDD.n708 VSS 0.009915f
C17848 DVDD.n709 VSS 0.009915f
C17849 DVDD.n710 VSS 0.009915f
C17850 DVDD.n711 VSS 0.009915f
C17851 DVDD.n712 VSS 0.009915f
C17852 DVDD.n713 VSS 0.009915f
C17853 DVDD.n714 VSS 0.009915f
C17854 DVDD.n715 VSS 0.201544f
C17855 DVDD.n716 VSS 0.009915f
C17856 DVDD.n717 VSS 0.009915f
C17857 DVDD.n718 VSS 0.009915f
C17858 DVDD.n719 VSS 0.009915f
C17859 DVDD.n720 VSS 0.009915f
C17860 DVDD.n721 VSS 0.009915f
C17861 DVDD.n722 VSS 0.009915f
C17862 DVDD.n723 VSS 0.009915f
C17863 DVDD.n724 VSS 0.009915f
C17864 DVDD.n725 VSS 0.009915f
C17865 DVDD.n726 VSS 0.018711f
C17866 DVDD.n727 VSS 0.011035f
C17867 DVDD.n728 VSS 0.279212f
C17868 DVDD.n729 VSS 0.279212f
C17869 DVDD.n730 VSS 0.279212f
C17870 DVDD.n731 VSS 0.178932f
C17871 DVDD.n732 VSS 0.178932f
C17872 DVDD.n733 VSS 0.239887f
C17873 DVDD.n734 VSS 0.279212f
C17874 DVDD.n735 VSS 0.017212f
C17875 DVDD.n736 VSS 0.009915f
C17876 DVDD.n737 VSS 0.009915f
C17877 DVDD.n738 VSS 0.009915f
C17878 DVDD.n739 VSS -0.292745f
C17879 DVDD.n740 VSS 0.009915f
C17880 DVDD.n741 VSS 0.019831f
C17881 DVDD.n742 VSS 0.010155f
C17882 DVDD.n743 VSS 0.019831f
C17883 DVDD.n744 VSS 0.009915f
C17884 DVDD.n745 VSS 0.009915f
C17885 DVDD.n746 VSS 0.019831f
C17886 DVDD.n747 VSS 0.009915f
C17887 DVDD.n748 VSS 0.019831f
C17888 DVDD.n749 VSS 0.009915f
C17889 DVDD.n750 VSS 0.019831f
C17890 DVDD.n751 VSS 0.009915f
C17891 DVDD.n752 VSS 0.019831f
C17892 DVDD.n753 VSS 0.010475f
C17893 DVDD.n754 VSS 0.019831f
C17894 DVDD.n755 VSS 0.009915f
C17895 DVDD.n756 VSS 0.009915f
C17896 DVDD.n757 VSS 0.019831f
C17897 DVDD.n758 VSS 0.011355f
C17898 DVDD.n759 VSS 0.0615f
C17899 DVDD.n760 VSS 0.011355f
C17900 DVDD.n761 VSS 0.019831f
C17901 DVDD.n762 VSS 0.019831f
C17902 DVDD.n763 VSS 0.014873f
C17903 DVDD.n764 VSS 0.019831f
C17904 DVDD.n765 VSS 0.014953f
C17905 DVDD.n766 VSS 0.019831f
C17906 DVDD.n767 VSS 0.019831f
C17907 DVDD.n768 VSS 0.011355f
C17908 DVDD.n769 VSS 0.009915f
C17909 DVDD.n770 VSS 0.011355f
C17910 DVDD.n771 VSS 0.009915f
C17911 DVDD.n772 VSS 0.011355f
C17912 DVDD.n773 VSS 0.019831f
C17913 DVDD.n774 VSS 0.019831f
C17914 DVDD.n775 VSS 0.019831f
C17915 DVDD.n776 VSS 0.010795f
C17916 DVDD.n777 VSS 0.009915f
C17917 DVDD.n778 VSS 0.011355f
C17918 DVDD.n779 VSS 0.009915f
C17919 DVDD.n780 VSS 0.011355f
C17920 DVDD.n781 VSS 0.019831f
C17921 DVDD.n782 VSS 0.019831f
C17922 DVDD.n783 VSS 0.011355f
C17923 DVDD.n784 VSS 0.009915f
C17924 DVDD.n785 VSS 0.011355f
C17925 DVDD.n786 VSS 0.009915f
C17926 DVDD.n787 VSS 0.011355f
C17927 DVDD.n788 VSS 0.019831f
C17928 DVDD.n789 VSS 0.019831f
C17929 DVDD.n790 VSS 0.011355f
C17930 DVDD.n791 VSS 0.009915f
C17931 DVDD.n792 VSS 0.010315f
C17932 DVDD.n793 VSS 0.010955f
C17933 DVDD.n794 VSS 0.019831f
C17934 DVDD.n795 VSS 0.019831f
C17935 DVDD.n796 VSS 0.011355f
C17936 DVDD.n797 VSS 0.009915f
C17937 DVDD.n798 VSS 0.011355f
C17938 DVDD.n799 VSS 0.009915f
C17939 DVDD.n800 VSS 0.011355f
C17940 DVDD.n801 VSS 0.019831f
C17941 DVDD.n802 VSS 0.019831f
C17942 DVDD.n803 VSS 0.011355f
C17943 DVDD.n804 VSS 0.009915f
C17944 DVDD.n805 VSS 0.011355f
C17945 DVDD.n806 VSS 0.009915f
C17946 DVDD.n807 VSS 0.011355f
C17947 DVDD.n808 VSS 0.019831f
C17948 DVDD.n809 VSS 0.019831f
C17949 DVDD.n810 VSS 0.019831f
C17950 DVDD.n811 VSS 0.011115f
C17951 DVDD.n812 VSS 0.009915f
C17952 DVDD.n813 VSS 0.011355f
C17953 DVDD.n814 VSS 0.009915f
C17954 DVDD.n815 VSS 0.011355f
C17955 DVDD.n816 VSS 0.019831f
C17956 DVDD.n817 VSS 0.019831f
C17957 DVDD.n818 VSS 0.015753f
C17958 DVDD.n819 VSS 0.019831f
C17959 DVDD.n820 VSS 0.011994f
C17960 DVDD.n821 VSS -0.359726f
C17961 DVDD.n822 VSS 0.011355f
C17962 DVDD.n823 VSS 0.019831f
C17963 DVDD.n824 VSS 0.011355f
C17964 DVDD.n825 VSS 0.019831f
C17965 DVDD.n826 VSS 0.011355f
C17966 DVDD.n827 VSS 0.019831f
C17967 DVDD.n828 VSS 0.011355f
C17968 DVDD.n829 VSS 0.019831f
C17969 DVDD.n830 VSS 0.011355f
C17970 DVDD.n831 VSS 0.019831f
C17971 DVDD.n832 VSS 0.019831f
C17972 DVDD.n833 VSS 0.010555f
C17973 DVDD.n834 VSS 0.010715f
C17974 DVDD.n835 VSS 0.019831f
C17975 DVDD.n836 VSS 0.011355f
C17976 DVDD.n837 VSS 0.019831f
C17977 DVDD.n838 VSS 0.011355f
C17978 DVDD.n839 VSS 0.019831f
C17979 DVDD.n840 VSS 0.011355f
C17980 DVDD.n841 VSS 0.019831f
C17981 DVDD.n842 VSS 0.011355f
C17982 DVDD.n843 VSS 0.019831f
C17983 DVDD.n844 VSS 0.011355f
C17984 DVDD.n845 VSS 0.019831f
C17985 DVDD.n846 VSS 0.011355f
C17986 DVDD.n847 VSS 0.019831f
C17987 DVDD.n848 VSS 0.019831f
C17988 DVDD.n849 VSS 0.010395f
C17989 DVDD.n850 VSS 0.010875f
C17990 DVDD.n851 VSS 0.019831f
C17991 DVDD.n852 VSS 0.011355f
C17992 DVDD.n853 VSS 0.019831f
C17993 DVDD.n854 VSS 0.011355f
C17994 DVDD.n855 VSS 0.019831f
C17995 DVDD.n856 VSS 0.011355f
C17996 DVDD.n857 VSS 0.019831f
C17997 DVDD.n858 VSS 0.011355f
C17998 DVDD.n859 VSS 0.019831f
C17999 DVDD.n860 VSS 0.011355f
C18000 DVDD.n861 VSS 0.019831f
C18001 DVDD.n862 VSS 0.011355f
C18002 DVDD.n863 VSS 0.019831f
C18003 DVDD.n864 VSS 0.010235f
C18004 DVDD.n865 VSS 0.019831f
C18005 DVDD.n866 VSS 0.019831f
C18006 DVDD.n867 VSS 0.019831f
C18007 DVDD.n868 VSS 0.019831f
C18008 DVDD.n869 VSS 0.019831f
C18009 DVDD.n870 VSS 0.013034f
C18010 DVDD.n871 VSS 0.019831f
C18011 DVDD.n872 VSS 0.011355f
C18012 DVDD.n873 VSS 0.019831f
C18013 DVDD.n874 VSS 0.011355f
C18014 DVDD.n875 VSS 0.019831f
C18015 DVDD.n876 VSS 0.011355f
C18016 DVDD.n877 VSS 0.063326f
C18017 DVDD.n878 VSS 0.005821f
C18018 DVDD.n879 VSS 0.279212f
C18019 DVDD.n880 VSS 0.279212f
C18020 DVDD.n881 VSS 0.279212f
C18021 DVDD.n882 VSS 0.279212f
C18022 DVDD.n883 VSS 0.279212f
C18023 DVDD.n884 VSS 0.279212f
C18024 DVDD.n885 VSS 0.279212f
C18025 DVDD.n886 VSS 0.279212f
C18026 DVDD.n887 VSS 0.279212f
C18027 DVDD.n888 VSS 0.279212f
C18028 DVDD.n889 VSS 0.279212f
C18029 DVDD.n890 VSS 0.279212f
C18030 DVDD.n891 VSS 0.139606f
C18031 DVDD.n892 VSS 0.017212f
C18032 DVDD.n893 VSS 0.009915f
C18033 DVDD.n894 VSS 0.009915f
C18034 DVDD.n895 VSS 0.009915f
C18035 DVDD.n896 VSS 0.005821f
C18036 DVDD.n897 VSS 0.279212f
C18037 DVDD.n898 VSS 0.279212f
C18038 DVDD.n899 VSS 0.279212f
C18039 DVDD.n900 VSS 0.279212f
C18040 DVDD.n901 VSS 0.279212f
C18041 DVDD.n902 VSS 0.279212f
C18042 DVDD.n903 VSS 0.279212f
C18043 DVDD.n904 VSS 0.279212f
C18044 DVDD.n905 VSS 0.279212f
C18045 DVDD.n906 VSS 0.279212f
C18046 DVDD.n907 VSS 0.336235f
C18047 DVDD.n908 VSS 0.336235f
C18048 DVDD.n909 VSS 0.532863f
C18049 DVDD.n910 VSS 0.139606f
C18050 DVDD.n911 VSS 0.279212f
C18051 DVDD.n912 VSS 0.279212f
C18052 DVDD.n913 VSS 0.279212f
C18053 DVDD.n914 VSS 0.090449f
C18054 DVDD.n915 VSS 0.021998f
C18055 DVDD.n916 VSS 0.015767f
C18056 DVDD.n917 VSS 0.015767f
C18057 DVDD.n918 VSS 0.015767f
C18058 DVDD.n919 VSS 0.015767f
C18059 DVDD.n920 VSS 0.015767f
C18060 DVDD.n921 VSS 0.139606f
C18061 DVDD.n922 VSS 0.090449f
C18062 DVDD.n923 VSS 0.015767f
C18063 DVDD.n924 VSS 0.015767f
C18064 DVDD.n925 VSS 0.015767f
C18065 DVDD.n926 VSS 0.015767f
C18066 DVDD.n927 VSS 0.018056f
C18067 DVDD.n928 VSS 0.196455f
C18068 DVDD.n929 VSS 0.018056f
C18069 DVDD.n930 VSS 0.045107f
C18070 DVDD.n931 VSS 0.018056f
C18071 DVDD.n932 VSS 0.060142f
C18072 DVDD.n933 VSS 0.018056f
C18073 DVDD.n934 VSS 0.060142f
C18074 DVDD.n935 VSS 0.060142f
C18075 DVDD.n936 VSS 0.017929f
C18076 DVDD.n937 VSS 0.015894f
C18077 DVDD.n938 VSS 0.060142f
C18078 DVDD.n939 VSS 0.060142f
C18079 DVDD.n940 VSS 0.018056f
C18080 DVDD.n941 VSS 0.015767f
C18081 DVDD.n942 VSS 0.018056f
C18082 DVDD.n943 VSS 0.058989f
C18083 DVDD.n944 VSS 0.064128f
C18084 DVDD.n945 VSS 0.023609f
C18085 DVDD.n946 VSS 0.023609f
C18086 DVDD.n947 VSS 0.023609f
C18087 DVDD.n948 VSS 0.027036f
C18088 DVDD.n949 VSS 0.019967f
C18089 DVDD.n950 VSS 0.018056f
C18090 DVDD.n951 VSS 0.045107f
C18091 DVDD.n952 VSS 0.018056f
C18092 DVDD.n953 VSS 0.060142f
C18093 DVDD.n954 VSS 0.060142f
C18094 DVDD.n955 VSS 0.017929f
C18095 DVDD.n956 VSS 0.015894f
C18096 DVDD.n957 VSS 0.060142f
C18097 DVDD.n958 VSS 0.018056f
C18098 DVDD.n959 VSS 0.060142f
C18099 DVDD.n960 VSS 0.107455f
C18100 DVDD.n961 VSS 0.140017f
C18101 DVDD.n962 VSS 0.027036f
C18102 DVDD.n963 VSS 0.070301f
C18103 DVDD.n964 VSS 0.027036f
C18104 DVDD.n965 VSS 0.04904f
C18105 DVDD.n966 VSS 0.03515f
C18106 DVDD.n967 VSS 0.027036f
C18107 DVDD.n968 VSS 0.056411f
C18108 DVDD.n969 VSS 0.070301f
C18109 DVDD.n970 VSS 0.070301f
C18110 DVDD.n971 VSS 0.139606f
C18111 DVDD.n972 VSS 0.139606f
C18112 DVDD.n973 VSS 0.026275f
C18113 DVDD.n974 VSS 0.139606f
C18114 DVDD.n975 VSS 0.198595f
C18115 DVDD.n976 VSS 0.02361f
C18116 DVDD.n977 VSS 0.02361f
C18117 DVDD.n978 VSS 0.02361f
C18118 DVDD.n979 VSS 0.02361f
C18119 DVDD.n980 VSS 0.02361f
C18120 DVDD.n981 VSS 0.02361f
C18121 DVDD.n982 VSS 0.02361f
C18122 DVDD.n983 VSS 0.02361f
C18123 DVDD.n984 VSS 0.02361f
C18124 DVDD.n985 VSS 0.279212f
C18125 DVDD.n986 VSS 0.279212f
C18126 DVDD.n987 VSS 0.279212f
C18127 DVDD.n988 VSS 0.279212f
C18128 DVDD.n989 VSS 0.186797f
C18129 DVDD.n990 VSS 0.532863f
C18130 DVDD.n991 VSS 0.232022f
C18131 DVDD.n992 VSS 0.279212f
C18132 DVDD.n993 VSS 0.279212f
C18133 DVDD.n994 VSS 0.279212f
C18134 DVDD.n995 VSS 0.279212f
C18135 DVDD.n996 VSS 0.279212f
C18136 DVDD.n997 VSS 0.279212f
C18137 DVDD.n998 VSS 0.279212f
C18138 DVDD.n999 VSS 0.279212f
C18139 DVDD.n1000 VSS 0.279212f
C18140 DVDD.n1001 VSS 0.279212f
C18141 DVDD.n1002 VSS 0.279212f
C18142 DVDD.n1003 VSS 0.279212f
C18143 DVDD.n1004 VSS 0.279212f
C18144 DVDD.n1005 VSS 0.139606f
C18145 DVDD.n1006 VSS 0.279212f
C18146 DVDD.n1007 VSS 0.279212f
C18147 DVDD.n1008 VSS 0.279212f
C18148 DVDD.n1009 VSS 0.279212f
C18149 DVDD.n1010 VSS 0.009915f
C18150 DVDD.n1011 VSS 0.009915f
C18151 DVDD.n1012 VSS 0.009915f
C18152 DVDD.n1013 VSS 0.009915f
C18153 DVDD.n1014 VSS 0.009915f
C18154 DVDD.n1015 VSS 0.009915f
C18155 DVDD.n1016 VSS 0.009915f
C18156 DVDD.n1017 VSS 0.009915f
C18157 DVDD.n1018 VSS 0.009915f
C18158 DVDD.n1019 VSS 0.009915f
C18159 DVDD.n1020 VSS 0.279212f
C18160 DVDD.n1021 VSS 0.279212f
C18161 DVDD.n1022 VSS 0.279212f
C18162 DVDD.n1023 VSS 0.279212f
C18163 DVDD.n1024 VSS 0.279212f
C18164 DVDD.n1025 VSS 0.279212f
C18165 DVDD.n1026 VSS 0.279212f
C18166 DVDD.n1027 VSS 0.279212f
C18167 DVDD.n1028 VSS 0.279212f
C18168 DVDD.n1029 VSS 0.279212f
C18169 DVDD.n1030 VSS 0.279212f
C18170 DVDD.n1031 VSS 0.279212f
C18171 DVDD.n1032 VSS 0.279212f
C18172 DVDD.n1033 VSS 0.279212f
C18173 DVDD.n1034 VSS 0.279212f
C18174 DVDD.n1035 VSS 0.279212f
C18175 DVDD.n1036 VSS 0.279212f
C18176 DVDD.n1037 VSS 0.279212f
C18177 DVDD.n1038 VSS 0.279212f
C18178 DVDD.n1039 VSS 0.279212f
C18179 DVDD.n1040 VSS 0.279212f
C18180 DVDD.n1041 VSS 0.279212f
C18181 DVDD.n1042 VSS 0.279212f
C18182 DVDD.n1043 VSS 0.279212f
C18183 DVDD.n1044 VSS 0.279212f
C18184 DVDD.n1045 VSS 0.279212f
C18185 DVDD.n1046 VSS 0.264465f
C18186 DVDD.n1047 VSS 0.009915f
C18187 DVDD.n1048 VSS 0.009915f
C18188 DVDD.n1049 VSS 0.009915f
C18189 DVDD.n1050 VSS 0.009915f
C18190 DVDD.n1051 VSS 0.009915f
C18191 DVDD.n1052 VSS 0.009915f
C18192 DVDD.n1053 VSS 0.009915f
C18193 DVDD.n1054 VSS 0.009915f
C18194 DVDD.n1055 VSS 0.009915f
C18195 DVDD.n1056 VSS 0.009915f
C18196 DVDD.n1057 VSS 0.018711f
C18197 DVDD.n1058 VSS 0.010235f
C18198 DVDD.n1059 VSS 0.011355f
C18199 DVDD.n1060 VSS 0.063326f
C18200 DVDD.n1061 VSS 0.011355f
C18201 DVDD.n1062 VSS 0.019831f
C18202 DVDD.n1063 VSS 0.011355f
C18203 DVDD.n1064 VSS 0.019831f
C18204 DVDD.n1065 VSS 0.019831f
C18205 DVDD.n1066 VSS 0.013034f
C18206 DVDD.n1067 VSS 0.019831f
C18207 DVDD.n1068 VSS 0.019831f
C18208 DVDD.n1069 VSS 0.019831f
C18209 DVDD.n1070 VSS -0.292745f
C18210 DVDD.n1071 VSS 0.009915f
C18211 DVDD.n1072 VSS 0.019831f
C18212 DVDD.n1073 VSS 0.139606f
C18213 DVDD.n1074 VSS 0.011355f
C18214 DVDD.n1075 VSS 0.154353f
C18215 DVDD.n1076 VSS 0.009915f
C18216 DVDD.n1077 VSS 0.009915f
C18217 DVDD.n1078 VSS 0.009915f
C18218 DVDD.n1079 VSS 0.009915f
C18219 DVDD.n1080 VSS 0.009915f
C18220 DVDD.n1081 VSS 0.009915f
C18221 DVDD.n1082 VSS 0.009915f
C18222 DVDD.n1083 VSS 0.009915f
C18223 DVDD.n1084 VSS 0.009915f
C18224 DVDD.n1085 VSS 0.279212f
C18225 DVDD.n1086 VSS 0.279212f
C18226 DVDD.n1087 VSS 0.279212f
C18227 DVDD.n1088 VSS 0.279212f
C18228 DVDD.n1089 VSS 0.279212f
C18229 DVDD.n1090 VSS 0.279212f
C18230 DVDD.n1091 VSS 0.279212f
C18231 DVDD.n1092 VSS 0.279212f
C18232 DVDD.n1093 VSS 0.279212f
C18233 DVDD.n1094 VSS 0.532863f
C18234 DVDD.n1095 VSS 0.336235f
C18235 DVDD.n1096 VSS 0.279212f
C18236 DVDD.n1097 VSS 0.279212f
C18237 DVDD.n1098 VSS 0.279212f
C18238 DVDD.n1099 VSS 0.279212f
C18239 DVDD.n1100 VSS 0.279212f
C18240 DVDD.n1101 VSS 0.279212f
C18241 DVDD.n1102 VSS 0.279212f
C18242 DVDD.n1103 VSS 0.279212f
C18243 DVDD.n1104 VSS 0.279212f
C18244 DVDD.n1105 VSS 0.279212f
C18245 DVDD.n1106 VSS 1.0352f
C18246 DVDD.n1107 VSS 0.279212f
C18247 DVDD.n1108 VSS 0.139606f
C18248 DVDD.n1109 VSS 0.037228f
C18249 DVDD.n1110 VSS 0.037228f
C18250 DVDD.n1111 VSS 0.037228f
C18251 DVDD.n1112 VSS 0.037228f
C18252 DVDD.n1113 VSS 0.037228f
C18253 DVDD.n1114 VSS 0.037228f
C18254 DVDD.n1115 VSS 0.037228f
C18255 DVDD.n1116 VSS 0.037228f
C18256 DVDD.n1117 VSS 0.037228f
C18257 DVDD.n1118 VSS 0.037228f
C18258 DVDD.n1120 VSS 0.624053f
C18259 DVDD.n1121 VSS 0.139606f
C18260 DVDD.n1122 VSS 0.042254f
C18261 DVDD.n1123 VSS 0.042254f
C18262 DVDD.n1124 VSS 0.042254f
C18263 DVDD.n1125 VSS 0.042254f
C18264 DVDD.n1126 VSS 0.042254f
C18265 DVDD.n1127 VSS 0.042254f
C18266 DVDD.n1128 VSS 0.042254f
C18267 DVDD.n1129 VSS 0.042254f
C18268 DVDD.n1130 VSS 0.042254f
C18269 DVDD.n1131 VSS 0.15632f
C18270 DVDD.n1134 VSS 0.042254f
C18271 DVDD.n1136 VSS 0.042254f
C18272 DVDD.n1138 VSS 0.042254f
C18273 DVDD.n1140 VSS 0.042254f
C18274 DVDD.n1142 VSS 0.042254f
C18275 DVDD.n1144 VSS 0.042254f
C18276 DVDD.n1146 VSS 0.042254f
C18277 DVDD.n1148 VSS 0.042254f
C18278 DVDD.n1150 VSS 0.532172f
C18279 DVDD.n1151 VSS 1.0352f
C18280 DVDD.n1152 VSS 0.279212f
C18281 DVDD.n1153 VSS 0.279212f
C18282 DVDD.n1154 VSS 0.279212f
C18283 DVDD.n1155 VSS 0.279212f
C18284 DVDD.n1156 VSS 0.279212f
C18285 DVDD.n1157 VSS 0.279212f
C18286 DVDD.n1158 VSS 0.279212f
C18287 DVDD.n1159 VSS 0.279212f
C18288 DVDD.n1160 VSS 0.279212f
C18289 DVDD.n1161 VSS 0.188763f
C18290 DVDD.n1162 VSS 0.279212f
C18291 DVDD.n1163 VSS 0.279212f
C18292 DVDD.n1164 VSS 0.279212f
C18293 DVDD.n1165 VSS 0.279212f
C18294 DVDD.n1166 VSS 0.279212f
C18295 DVDD.n1167 VSS 0.279212f
C18296 DVDD.n1168 VSS 0.279212f
C18297 DVDD.n1169 VSS 0.279212f
C18298 DVDD.n1170 VSS 0.279212f
C18299 DVDD.n1171 VSS 0.279212f
C18300 DVDD.n1172 VSS 0.279212f
C18301 DVDD.n1173 VSS 0.279212f
C18302 DVDD.n1174 VSS 0.279212f
C18303 DVDD.n1175 VSS 0.279212f
C18304 DVDD.n1176 VSS 0.279212f
C18305 DVDD.n1177 VSS 0.279212f
C18306 DVDD.n1178 VSS 0.279212f
C18307 DVDD.n1179 VSS 0.279212f
C18308 DVDD.n1180 VSS 0.279212f
C18309 DVDD.n1181 VSS 0.139606f
C18310 DVDD.n1189 VSS 0.042254f
C18311 DVDD.n1192 VSS 0.06515f
C18312 DVDD.n1193 VSS 0.486474f
C18313 DVDD.n1194 VSS 0.061892f
C18314 DVDD.n1195 VSS 0.041407f
C18315 DVDD.n1196 VSS 0.061892f
C18316 DVDD.n1197 VSS 0.06515f
C18317 DVDD.n1199 VSS 0.061892f
C18318 DVDD.n1200 VSS 0.051431f
C18319 DVDD.n1202 VSS 0.061892f
C18320 DVDD.n1205 VSS 0.193533f
C18321 DVDD.n1206 VSS 0.130299f
C18322 DVDD.n1207 VSS 0.130299f
C18323 DVDD.n1208 VSS 0.130299f
C18324 DVDD.n1209 VSS 0.112406f
C18325 DVDD.n1210 VSS 0.130299f
C18326 DVDD.n1211 VSS 0.130299f
C18327 DVDD.n1212 VSS 0.130299f
C18328 DVDD.n1213 VSS 0.130299f
C18329 DVDD.n1214 VSS 0.016758f
C18330 DVDD.n1215 VSS 0.008859f
C18331 DVDD.n1216 VSS 0.008859f
C18332 DVDD.n1217 VSS 0.008859f
C18333 DVDD.n1218 VSS 0.06515f
C18334 DVDD.n1219 VSS 0.008859f
C18335 DVDD.n1220 VSS 0.005501f
C18336 DVDD.n1221 VSS 0.008859f
C18337 DVDD.n1222 VSS 0.003689f
C18338 DVDD.n1223 VSS 0.130299f
C18339 DVDD.n1224 VSS 0.130299f
C18340 DVDD.n1225 VSS 0.130299f
C18341 DVDD.n1226 VSS 0.130299f
C18342 DVDD.n1227 VSS 0.130299f
C18343 DVDD.n1228 VSS 0.130299f
C18344 DVDD.n1229 VSS 0.130299f
C18345 DVDD.n1230 VSS 0.130299f
C18346 DVDD.n1231 VSS 0.130299f
C18347 DVDD.n1232 VSS 0.130299f
C18348 DVDD.n1233 VSS 0.130299f
C18349 DVDD.n1234 VSS 0.130299f
C18350 DVDD.n1235 VSS 0.130299f
C18351 DVDD.n1236 VSS 0.130299f
C18352 DVDD.n1237 VSS 0.130299f
C18353 DVDD.n1238 VSS 0.130299f
C18354 DVDD.n1239 VSS 0.130299f
C18355 DVDD.n1240 VSS 0.130299f
C18356 DVDD.n1241 VSS 0.130299f
C18357 DVDD.n1242 VSS 0.130299f
C18358 DVDD.n1243 VSS 0.130299f
C18359 DVDD.n1244 VSS 0.130299f
C18360 DVDD.n1245 VSS 0.130299f
C18361 DVDD.n1246 VSS 0.130299f
C18362 DVDD.n1247 VSS 0.130299f
C18363 DVDD.n1248 VSS 0.130299f
C18364 DVDD.n1249 VSS 0.130299f
C18365 DVDD.n1250 VSS 0.130299f
C18366 DVDD.n1251 VSS 0.130299f
C18367 DVDD.n1252 VSS 0.130299f
C18368 DVDD.n1253 VSS 0.130299f
C18369 DVDD.n1254 VSS 0.130299f
C18370 DVDD.n1255 VSS 0.130299f
C18371 DVDD.n1256 VSS 0.130299f
C18372 DVDD.n1257 VSS 0.130299f
C18373 DVDD.n1258 VSS 0.130299f
C18374 DVDD.n1259 VSS 0.130299f
C18375 DVDD.n1260 VSS 0.130299f
C18376 DVDD.n1261 VSS 0.130299f
C18377 DVDD.n1262 VSS 0.130299f
C18378 DVDD.n1263 VSS 0.130299f
C18379 DVDD.n1264 VSS 0.130299f
C18380 DVDD.n1265 VSS 0.130299f
C18381 DVDD.n1266 VSS 0.130299f
C18382 DVDD.n1267 VSS 0.130299f
C18383 DVDD.n1268 VSS 0.130299f
C18384 DVDD.n1269 VSS 0.130299f
C18385 DVDD.n1270 VSS 0.130299f
C18386 DVDD.n1271 VSS 0.130299f
C18387 DVDD.n1272 VSS 0.130299f
C18388 DVDD.n1273 VSS 0.130299f
C18389 DVDD.n1274 VSS 0.130299f
C18390 DVDD.n1275 VSS 0.130299f
C18391 DVDD.n1276 VSS 0.130299f
C18392 DVDD.n1277 VSS 0.130299f
C18393 DVDD.n1278 VSS 0.130299f
C18394 DVDD.n1279 VSS 0.130299f
C18395 DVDD.n1280 VSS 0.130299f
C18396 DVDD.n1281 VSS 0.130299f
C18397 DVDD.n1282 VSS 0.130299f
C18398 DVDD.n1283 VSS 0.130299f
C18399 DVDD.n1284 VSS 0.130299f
C18400 DVDD.n1285 VSS 0.130299f
C18401 DVDD.n1286 VSS 0.130299f
C18402 DVDD.n1287 VSS 0.130299f
C18403 DVDD.n1288 VSS 0.130299f
C18404 DVDD.n1289 VSS 0.130299f
C18405 DVDD.n1290 VSS 0.130299f
C18406 DVDD.n1291 VSS 0.130299f
C18407 DVDD.n1292 VSS 0.130299f
C18408 DVDD.n1293 VSS 0.130299f
C18409 DVDD.n1294 VSS 0.130299f
C18410 DVDD.n1295 VSS 0.130299f
C18411 DVDD.n1296 VSS 0.130299f
C18412 DVDD.n1297 VSS 0.130299f
C18413 DVDD.n1298 VSS 0.130299f
C18414 DVDD.n1299 VSS 0.130299f
C18415 DVDD.n1300 VSS 0.130299f
C18416 DVDD.n1301 VSS 0.116994f
C18417 DVDD.n1302 VSS 0.130299f
C18418 DVDD.n1303 VSS 0.130299f
C18419 DVDD.n1304 VSS 0.130299f
C18420 DVDD.n1305 VSS 0.06515f
C18421 DVDD.n1306 VSS 0.005501f
C18422 DVDD.n1307 VSS 0.008859f
C18423 DVDD.n1308 VSS 0.008859f
C18424 DVDD.n1309 VSS 0.016758f
C18425 DVDD.n1310 VSS 0.078455f
C18426 DVDD.n1311 VSS 0.008859f
C18427 DVDD.n1312 VSS 0.008859f
C18428 DVDD.n1313 VSS 0.008859f
C18429 DVDD.n1314 VSS 0.010145f
C18430 DVDD.n1315 VSS 0.036655f
C18431 DVDD.n1316 VSS 0.033199f
C18432 DVDD.n1317 VSS 0.010145f
C18433 DVDD.n1318 VSS 0.010145f
C18434 DVDD.n1320 VSS 0.010145f
C18435 DVDD.n1321 VSS 0.00893f
C18436 DVDD.n1322 VSS 0.010073f
C18437 DVDD.n1323 VSS 0.137213f
C18438 DVDD.n1324 VSS 0.010145f
C18439 DVDD.n1325 VSS 1.47856f
C18440 DVDD.n1326 VSS 8.54052f
C18441 DVDD.n1327 VSS 3.61626f
C18442 DVDD.n1328 VSS 2.53032f
C18443 DVDD.n1329 VSS 0.027843f
C18444 DVDD.n1331 VSS 0.06515f
C18445 DVDD.n1332 VSS 0.033505f
C18446 DVDD.n1335 VSS 0.033505f
C18447 DVDD.n1336 VSS 0.025719f
C18448 DVDD.n1337 VSS 0.06515f
C18449 DVDD.n1339 VSS 0.033505f
C18450 DVDD.n1340 VSS 0.06515f
C18451 DVDD.n1342 VSS 0.130299f
C18452 DVDD.n1343 VSS 0.130299f
C18453 DVDD.n1344 VSS 0.130299f
C18454 DVDD.n1345 VSS 0.130299f
C18455 DVDD.n1346 VSS 0.130299f
C18456 DVDD.n1347 VSS 0.130299f
C18457 DVDD.n1348 VSS 0.130299f
C18458 DVDD.n1349 VSS 0.130299f
C18459 DVDD.n1350 VSS 0.130299f
C18460 DVDD.n1351 VSS 0.130299f
C18461 DVDD.n1352 VSS 0.130299f
C18462 DVDD.n1353 VSS 0.130299f
C18463 DVDD.n1354 VSS 0.130299f
C18464 DVDD.n1355 VSS 0.130299f
C18465 DVDD.n1356 VSS 0.130299f
C18466 DVDD.n1357 VSS 0.117453f
C18467 DVDD.n1358 VSS 0.117453f
C18468 DVDD.n1359 VSS 0.130299f
C18469 DVDD.n1360 VSS 0.066985f
C18470 DVDD.n1361 VSS 0.077996f
C18471 DVDD.n1362 VSS 0.212852f
C18472 DVDD.n1363 VSS 0.450198f
C18473 DVDD.n1364 VSS 0.504402f
C18474 DVDD.n1365 VSS 0.033505f
C18475 DVDD.n1367 VSS 0.025719f
C18476 DVDD.n1368 VSS 0.012846f
C18477 DVDD.n1369 VSS 0.022416f
C18478 DVDD.n1370 VSS 1.13814f
C18479 DVDD.n1371 VSS 1.15753f
C18480 DVDD.n1372 VSS 7.58992f
C18481 DVDD.n1373 VSS 5.61607f
C18482 DVDD.n1374 VSS 2.38892f
C18483 DVDD.n1375 VSS 5.62423f
C18484 DVDD.n1376 VSS 7.85556f
C18485 DVDD.n1377 VSS 8.80625f
C18486 DVDD.n1378 VSS 10.8381f
C18487 DVDD.n1379 VSS 5.84562f
C18488 DVDD.n1380 VSS 1.47386f
C18489 DVDD.n1381 VSS 0.010145f
C18490 DVDD.n1382 VSS 0.010145f
C18491 DVDD.n1383 VSS 0.00893f
C18492 DVDD.n1385 VSS 0.010073f
C18493 DVDD.n1386 VSS 0.010145f
C18494 DVDD.n1387 VSS 0.010145f
C18495 DVDD.n1388 VSS 0.11217f
C18496 DVDD.n1389 VSS 0.033199f
C18497 DVDD.n1390 VSS 0.010145f
C18498 DVDD.n1391 VSS 0.036655f
C18499 DVDD.n1392 VSS 0.003689f
C18500 DVDD.n1393 VSS 0.014605f
C18501 DVDD.n1394 VSS 0.06515f
C18502 DVDD.n1395 VSS 0.06515f
C18503 DVDD.n1396 VSS 0.130299f
C18504 DVDD.n1397 VSS 0.130299f
C18505 DVDD.n1398 VSS 0.130299f
C18506 DVDD.n1399 VSS 0.130299f
C18507 DVDD.n1400 VSS 0.130299f
C18508 DVDD.n1401 VSS 0.130299f
C18509 DVDD.n1402 VSS 0.130299f
C18510 DVDD.n1403 VSS 0.130299f
C18511 DVDD.n1404 VSS 0.130299f
C18512 DVDD.n1405 VSS 0.130299f
C18513 DVDD.n1406 VSS 0.130299f
C18514 DVDD.n1407 VSS 0.130299f
C18515 DVDD.n1408 VSS 0.130299f
C18516 DVDD.n1409 VSS 0.130299f
C18517 DVDD.n1410 VSS 0.130299f
C18518 DVDD.n1411 VSS 0.130299f
C18519 DVDD.n1412 VSS 0.130299f
C18520 DVDD.n1413 VSS 0.130299f
C18521 DVDD.n1414 VSS 0.130299f
C18522 DVDD.n1415 VSS 0.130299f
C18523 DVDD.n1416 VSS 0.130299f
C18524 DVDD.n1417 VSS 0.130299f
C18525 DVDD.n1418 VSS 0.130299f
C18526 DVDD.n1419 VSS 0.130299f
C18527 DVDD.n1420 VSS 0.130299f
C18528 DVDD.n1421 VSS 0.130299f
C18529 DVDD.n1422 VSS 0.130299f
C18530 DVDD.n1423 VSS 0.130299f
C18531 DVDD.n1424 VSS 0.130299f
C18532 DVDD.n1425 VSS 0.130299f
C18533 DVDD.n1426 VSS 0.130299f
C18534 DVDD.n1427 VSS 0.130299f
C18535 DVDD.n1428 VSS 0.130299f
C18536 DVDD.n1429 VSS 0.130299f
C18537 DVDD.n1430 VSS 0.130299f
C18538 DVDD.n1431 VSS 0.130299f
C18539 DVDD.n1432 VSS 0.130299f
C18540 DVDD.n1433 VSS 0.130299f
C18541 DVDD.n1434 VSS 0.130299f
C18542 DVDD.n1435 VSS 0.130299f
C18543 DVDD.n1436 VSS 0.130299f
C18544 DVDD.n1437 VSS 0.130299f
C18545 DVDD.n1438 VSS 0.130299f
C18546 DVDD.n1439 VSS 0.130299f
C18547 DVDD.n1440 VSS 0.130299f
C18548 DVDD.n1441 VSS 0.130299f
C18549 DVDD.n1442 VSS 0.130299f
C18550 DVDD.n1443 VSS 0.130299f
C18551 DVDD.n1444 VSS 0.130299f
C18552 DVDD.n1445 VSS 0.130299f
C18553 DVDD.n1446 VSS 0.130299f
C18554 DVDD.n1447 VSS 0.130299f
C18555 DVDD.n1448 VSS 0.130299f
C18556 DVDD.n1449 VSS 0.130299f
C18557 DVDD.n1450 VSS 0.130299f
C18558 DVDD.n1451 VSS 0.130299f
C18559 DVDD.n1452 VSS 0.130299f
C18560 DVDD.n1453 VSS 0.130299f
C18561 DVDD.n1454 VSS 0.130299f
C18562 DVDD.n1455 VSS 0.130299f
C18563 DVDD.n1456 VSS 0.130299f
C18564 DVDD.n1457 VSS 0.130299f
C18565 DVDD.n1458 VSS 0.130299f
C18566 DVDD.n1459 VSS 0.130299f
C18567 DVDD.n1460 VSS 0.130299f
C18568 DVDD.n1461 VSS 0.130299f
C18569 DVDD.n1462 VSS 0.130299f
C18570 DVDD.n1463 VSS 0.130299f
C18571 DVDD.n1464 VSS 0.130299f
C18572 DVDD.n1465 VSS 0.130299f
C18573 DVDD.n1466 VSS 0.130299f
C18574 DVDD.n1467 VSS 0.130299f
C18575 DVDD.n1468 VSS 0.130299f
C18576 DVDD.n1469 VSS 0.130299f
C18577 DVDD.n1470 VSS 0.130299f
C18578 DVDD.n1471 VSS 0.130299f
C18579 DVDD.n1472 VSS 0.130299f
C18580 DVDD.n1473 VSS 0.130299f
C18581 DVDD.n1474 VSS 0.130299f
C18582 DVDD.n1475 VSS 0.130299f
C18583 DVDD.n1476 VSS 0.130299f
C18584 DVDD.n1477 VSS 0.130299f
C18585 DVDD.n1478 VSS 0.130299f
C18586 DVDD.n1479 VSS 0.130299f
C18587 DVDD.n1480 VSS 0.130299f
C18588 DVDD.n1481 VSS 0.130299f
C18589 DVDD.n1482 VSS 0.130299f
C18590 DVDD.n1483 VSS 0.130299f
C18591 DVDD.n1484 VSS 0.130299f
C18592 DVDD.n1485 VSS 0.130299f
C18593 DVDD.n1486 VSS 0.130299f
C18594 DVDD.n1487 VSS 0.130299f
C18595 DVDD.n1488 VSS 0.130299f
C18596 DVDD.n1489 VSS 0.130299f
C18597 DVDD.n1490 VSS 0.130299f
C18598 DVDD.n1491 VSS 0.130299f
C18599 DVDD.n1492 VSS 0.130299f
C18600 DVDD.n1493 VSS 0.130299f
C18601 DVDD.n1494 VSS 0.130299f
C18602 DVDD.n1495 VSS 0.130299f
C18603 DVDD.n1496 VSS 0.130299f
C18604 DVDD.n1497 VSS 0.130299f
C18605 DVDD.n1498 VSS 0.130299f
C18606 DVDD.n1499 VSS 0.130299f
C18607 DVDD.n1500 VSS 0.130299f
C18608 DVDD.n1501 VSS 0.130299f
C18609 DVDD.n1502 VSS 0.130299f
C18610 DVDD.n1503 VSS 0.130299f
C18611 DVDD.n1504 VSS 0.130299f
C18612 DVDD.n1505 VSS 0.130299f
C18613 DVDD.n1506 VSS 0.130299f
C18614 DVDD.n1507 VSS 0.130299f
C18615 DVDD.n1508 VSS 0.130299f
C18616 DVDD.n1509 VSS 0.130299f
C18617 DVDD.n1510 VSS 0.130299f
C18618 DVDD.n1511 VSS 0.130299f
C18619 DVDD.n1512 VSS 0.130299f
C18620 DVDD.n1513 VSS 0.130299f
C18621 DVDD.n1514 VSS 0.130299f
C18622 DVDD.n1515 VSS 0.130299f
C18623 DVDD.n1516 VSS 0.130299f
C18624 DVDD.n1517 VSS 0.130299f
C18625 DVDD.n1518 VSS 0.130299f
C18626 DVDD.n1519 VSS 0.130299f
C18627 DVDD.n1520 VSS 0.130299f
C18628 DVDD.n1521 VSS 0.130299f
C18629 DVDD.n1522 VSS 0.130299f
C18630 DVDD.n1523 VSS 0.130299f
C18631 DVDD.n1524 VSS 0.130299f
C18632 DVDD.n1525 VSS 0.130299f
C18633 DVDD.n1526 VSS 0.130299f
C18634 DVDD.n1527 VSS 0.130299f
C18635 DVDD.n1528 VSS 0.130299f
C18636 DVDD.n1529 VSS 0.130299f
C18637 DVDD.n1530 VSS 0.130299f
C18638 DVDD.n1531 VSS 0.130299f
C18639 DVDD.n1532 VSS 0.130299f
C18640 DVDD.n1533 VSS 0.130299f
C18641 DVDD.n1534 VSS 0.130299f
C18642 DVDD.n1535 VSS 0.130299f
C18643 DVDD.n1536 VSS 0.130299f
C18644 DVDD.n1537 VSS 0.130299f
C18645 DVDD.n1538 VSS 0.130299f
C18646 DVDD.n1539 VSS 0.130299f
C18647 DVDD.n1540 VSS 0.130299f
C18648 DVDD.n1541 VSS 0.130299f
C18649 DVDD.n1542 VSS 0.130299f
C18650 DVDD.n1543 VSS 0.130299f
C18651 DVDD.n1544 VSS 0.130299f
C18652 DVDD.n1545 VSS 0.130299f
C18653 DVDD.n1546 VSS 0.130299f
C18654 DVDD.n1547 VSS 0.130299f
C18655 DVDD.n1548 VSS 0.130299f
C18656 DVDD.n1549 VSS 0.130299f
C18657 DVDD.n1550 VSS 0.130299f
C18658 DVDD.n1551 VSS 0.130299f
C18659 DVDD.n1552 VSS 0.130299f
C18660 DVDD.n1553 VSS 0.124335f
C18661 DVDD.n1554 VSS 0.06515f
C18662 DVDD.n1555 VSS 0.014605f
C18663 DVDD.n1556 VSS 0.06515f
C18664 DVDD.n1557 VSS 0.071114f
C18665 DVDD.n1558 VSS 0.130299f
C18666 DVDD.n1559 VSS 0.130299f
C18667 DVDD.n1560 VSS 0.130299f
C18668 DVDD.n1561 VSS 0.130299f
C18669 DVDD.n1562 VSS 0.130299f
C18670 DVDD.n1563 VSS 0.130299f
C18671 DVDD.n1564 VSS 0.130299f
C18672 DVDD.n1565 VSS 0.130299f
C18673 DVDD.n1566 VSS 0.130299f
C18674 DVDD.n1567 VSS 0.130299f
C18675 DVDD.n1568 VSS 0.130299f
C18676 DVDD.n1569 VSS 0.130299f
C18677 DVDD.n1570 VSS 0.705551f
C18678 DVDD.n1571 VSS 0.130299f
C18679 DVDD.n1572 VSS 0.06515f
C18680 DVDD.n1573 VSS 0.06515f
C18681 DVDD.n1575 VSS 0.047509f
C18682 DVDD.n1576 VSS 0.509743f
C18683 DVDD.n1577 VSS 0.187285f
C18684 DVDD.n1578 VSS 0.181353f
C18685 DVDD.n1579 VSS 0.139606f
C18686 DVDD.n1581 VSS 0.042254f
C18687 DVDD.n1582 VSS 0.139606f
C18688 DVDD.n1583 VSS 0.071861f
C18689 DVDD.n1584 VSS 0.065093f
C18690 DVDD.n1585 VSS 0.037228f
C18691 DVDD.n1586 VSS 0.037228f
C18692 DVDD.n1587 VSS 0.037228f
C18693 DVDD.n1588 VSS 0.037228f
C18694 DVDD.n1589 VSS 0.037228f
C18695 DVDD.n1590 VSS 0.037228f
C18696 DVDD.n1591 VSS 0.037228f
C18697 DVDD.n1592 VSS 0.037228f
C18698 DVDD.n1593 VSS 0.037228f
C18699 DVDD.n1595 VSS 0.624053f
C18700 DVDD.n1596 VSS 0.139606f
C18701 DVDD.n1597 VSS 0.037228f
C18702 DVDD.n1598 VSS 0.037228f
C18703 DVDD.n1599 VSS 0.037228f
C18704 DVDD.n1600 VSS 0.037228f
C18705 DVDD.n1601 VSS 0.037228f
C18706 DVDD.n1602 VSS 0.037228f
C18707 DVDD.n1603 VSS 0.037228f
C18708 DVDD.n1604 VSS 0.037228f
C18709 DVDD.n1605 VSS 0.037228f
C18710 DVDD.n1606 VSS 0.037228f
C18711 DVDD.n1607 VSS 0.15632f
C18712 DVDD.n1609 VSS 0.037228f
C18713 DVDD.n1611 VSS 0.037228f
C18714 DVDD.n1613 VSS 0.037228f
C18715 DVDD.n1615 VSS 0.037228f
C18716 DVDD.n1617 VSS 0.037228f
C18717 DVDD.n1619 VSS 0.037228f
C18718 DVDD.n1621 VSS 0.037228f
C18719 DVDD.n1623 VSS 0.037228f
C18720 DVDD.n1625 VSS 0.037228f
C18721 DVDD.n1627 VSS 0.624053f
C18722 DVDD.n1628 VSS 0.139606f
C18723 DVDD.n1629 VSS 0.037228f
C18724 DVDD.n1630 VSS 0.037228f
C18725 DVDD.n1631 VSS 0.037228f
C18726 DVDD.n1632 VSS 0.037228f
C18727 DVDD.n1633 VSS 0.037228f
C18728 DVDD.n1634 VSS 0.037228f
C18729 DVDD.n1635 VSS 0.037228f
C18730 DVDD.n1636 VSS 0.037228f
C18731 DVDD.n1637 VSS 0.037228f
C18732 DVDD.n1638 VSS 0.037228f
C18733 DVDD.n1639 VSS 0.15632f
C18734 DVDD.n1641 VSS 0.037228f
C18735 DVDD.n1643 VSS 0.037228f
C18736 DVDD.n1645 VSS 0.037228f
C18737 DVDD.n1647 VSS 0.037228f
C18738 DVDD.n1649 VSS 0.037228f
C18739 DVDD.n1651 VSS 0.037228f
C18740 DVDD.n1653 VSS 0.037228f
C18741 DVDD.n1655 VSS 0.037228f
C18742 DVDD.n1657 VSS 0.037228f
C18743 DVDD.n1658 VSS 0.037228f
C18744 DVDD.n1659 VSS 0.04016f
C18745 DVDD.n1660 VSS 0.08032f
C18746 DVDD.n1661 VSS 0.08032f
C18747 DVDD.n1662 VSS 0.08032f
C18748 DVDD.n1663 VSS 0.04016f
C18749 DVDD.n1664 VSS 0.037228f
C18750 DVDD.n1665 VSS 0.021211f
C18751 DVDD.n1666 VSS 0.056938f
C18752 DVDD.n1667 VSS 0.059108f
C18753 DVDD.n1668 VSS 0.148913f
C18754 DVDD.n1669 VSS 0.148913f
C18755 DVDD.n1670 VSS 0.055807f
C18756 DVDD.n1671 VSS 0.148913f
C18757 DVDD.n1672 VSS 0.148913f
C18758 DVDD.n1673 VSS 0.148913f
C18759 DVDD.n1674 VSS 0.148913f
C18760 DVDD.n1675 VSS 0.074652f
C18761 DVDD.n1676 VSS 0.148913f
C18762 DVDD.n1677 VSS 0.148913f
C18763 DVDD.n1678 VSS 0.148913f
C18764 DVDD.n1679 VSS 0.074457f
C18765 DVDD.n1680 VSS 0.074457f
C18766 DVDD.n1681 VSS 0.074457f
C18767 DVDD.n1682 VSS 0.012307f
C18768 DVDD.n1683 VSS 0.005305f
C18769 DVDD.n1684 VSS 0.025168f
C18770 DVDD.n1685 VSS 0.214063f
C18771 DVDD.n1686 VSS 0.123745f
C18772 DVDD.n1687 VSS 0.186797f
C18773 DVDD.n1688 VSS 0.279212f
C18774 DVDD.n1689 VSS 0.279212f
C18775 DVDD.n1690 VSS 0.169458f
C18776 DVDD.n1691 VSS 0.216649f
C18777 DVDD.n1692 VSS 0.279212f
C18778 DVDD.n1693 VSS 0.279212f
C18779 DVDD.n1694 VSS 0.279212f
C18780 DVDD.n1695 VSS 0.214611f
C18781 DVDD.n1696 VSS 0.279212f
C18782 DVDD.n1697 VSS 0.279212f
C18783 DVDD.n1698 VSS 0.279212f
C18784 DVDD.n1699 VSS 0.279212f
C18785 DVDD.n1700 VSS 0.162218f
C18786 DVDD.n1701 VSS 0.279212f
C18787 DVDD.n1702 VSS 0.279212f
C18788 DVDD.n1703 VSS 0.279212f
C18789 DVDD.n1704 VSS 0.279212f
C18790 DVDD.n1705 VSS 0.279212f
C18791 DVDD.n1706 VSS 0.151362f
C18792 DVDD.n1707 VSS 0.162218f
C18793 DVDD.n1708 VSS 0.038174f
C18794 DVDD.t0 VSS 0.590255f
C18795 DVDD.n1709 VSS -0.067592f
C18796 DVDD.t202 VSS 0.432504f
C18797 DVDD.t203 VSS 0.432504f
C18798 DVDD.n1710 VSS 0.054923f
C18799 DVDD.n1711 VSS -0.067592f
C18800 DVDD.t169 VSS 0.590255f
C18801 DVDD.n1712 VSS 0.236283f
C18802 DVDD.n1713 VSS 0.050823f
C18803 DVDD.t170 VSS 0.0973f
C18804 DVDD.n1714 VSS 0.124781f
C18805 DVDD.t133 VSS 0.040899f
C18806 DVDD.t147 VSS 0.040899f
C18807 DVDD.n1715 VSS 0.081797f
C18808 DVDD.n1716 VSS 0.100809f
C18809 DVDD.t172 VSS 0.0973f
C18810 DVDD.n1717 VSS 0.17088f
C18811 DVDD.n1718 VSS 0.044059f
C18812 DVDD.n1719 VSS 0.005305f
C18813 DVDD.n1720 VSS 0.007073f
C18814 DVDD.n1721 VSS 0.074457f
C18815 DVDD.n1722 VSS 0.11647f
C18816 DVDD.n1723 VSS 0.148913f
C18817 DVDD.n1724 VSS 0.214063f
C18818 DVDD.n1725 VSS 0.148913f
C18819 DVDD.n1726 VSS 0.148913f
C18820 DVDD.n1727 VSS 0.148913f
C18821 DVDD.n1728 VSS 0.061872f
C18822 DVDD.n1729 VSS 0.074457f
C18823 DVDD.n1730 VSS 0.074652f
C18824 DVDD.n1731 VSS 0.148913f
C18825 DVDD.n1732 VSS 0.148913f
C18826 DVDD.n1733 VSS 0.148913f
C18827 DVDD.n1734 VSS 0.125842f
C18828 DVDD.n1735 VSS 0.148913f
C18829 DVDD.n1736 VSS 0.148913f
C18830 DVDD.n1737 VSS 0.128988f
C18831 DVDD.n1738 VSS 0.128988f
C18832 DVDD.n1739 VSS 0.374604f
C18833 DVDD.n1740 VSS 0.46953f
C18834 DVDD.n1741 VSS 0.169753f
C18835 DVDD.n1742 VSS 0.369017f
C18836 DVDD.n1743 VSS 0.450446f
C18837 DVDD.n1744 VSS 0.128988f
C18838 DVDD.n1745 VSS 0.148913f
C18839 DVDD.n1746 VSS 0.148913f
C18840 DVDD.n1747 VSS 0.148913f
C18841 DVDD.n1748 VSS 0.148913f
C18842 DVDD.n1749 VSS 0.148913f
C18843 DVDD.n1750 VSS 0.148913f
C18844 DVDD.n1751 VSS 0.148913f
C18845 DVDD.n1752 VSS 0.148913f
C18846 DVDD.n1753 VSS 0.148913f
C18847 DVDD.n1754 VSS 0.148913f
C18848 DVDD.n1755 VSS 0.148913f
C18849 DVDD.n1756 VSS 0.148913f
C18850 DVDD.n1757 VSS 0.148913f
C18851 DVDD.n1758 VSS 0.148913f
C18852 DVDD.n1759 VSS 0.074457f
C18853 DVDD.n1760 VSS 0.074457f
C18854 DVDD.n1761 VSS 0.012307f
C18855 DVDD.n1762 VSS 0.007073f
C18856 DVDD.n1763 VSS 0.074457f
C18857 DVDD.n1764 VSS 0.074457f
C18858 DVDD.n1765 VSS 0.136329f
C18859 DVDD.n1766 VSS 0.136329f
C18860 DVDD.n1767 VSS 0.279212f
C18861 DVDD.n1768 VSS 0.279212f
C18862 DVDD.n1769 VSS 0.216649f
C18863 DVDD.n1770 VSS 0.279212f
C18864 DVDD.n1771 VSS 0.279212f
C18865 DVDD.n1772 VSS 0.279212f
C18866 DVDD.n1773 VSS 0.279212f
C18867 DVDD.n1774 VSS 0.279212f
C18868 DVDD.n1775 VSS 0.279212f
C18869 DVDD.n1776 VSS 0.279212f
C18870 DVDD.n1777 VSS 0.279212f
C18871 DVDD.n1778 VSS 0.279212f
C18872 DVDD.n1779 VSS 0.279212f
C18873 DVDD.n1780 VSS 0.268398f
C18874 DVDD.n1781 VSS 0.279212f
C18875 DVDD.n1782 VSS 0.279212f
C18876 DVDD.n1783 VSS 0.279212f
C18877 DVDD.n1784 VSS 0.279212f
C18878 DVDD.t184 VSS 0.0973f
C18879 DVDD.n1785 VSS 0.142981f
C18880 DVDD.n1786 VSS 0.207443f
C18881 DVDD.n1787 VSS 0.279212f
C18882 DVDD.n1788 VSS 0.247752f
C18883 DVDD.n1789 VSS 0.171067f
C18884 DVDD.n1790 VSS 0.091236f
C18885 DVDD.n1791 VSS 0.148913f
C18886 DVDD.n1792 VSS 0.214063f
C18887 DVDD.n1793 VSS 0.148913f
C18888 DVDD.n1794 VSS 0.091236f
C18889 DVDD.n1795 VSS 0.279212f
C18890 DVDD.n1796 VSS 0.279212f
C18891 DVDD.n1797 VSS 0.279212f
C18892 DVDD.n1798 VSS 0.279212f
C18893 DVDD.n1799 VSS 0.279212f
C18894 DVDD.n1800 VSS 0.279212f
C18895 DVDD.n1801 VSS 0.279212f
C18896 DVDD.n1802 VSS 0.279212f
C18897 DVDD.n1803 VSS 0.279212f
C18898 DVDD.n1804 VSS 0.279212f
C18899 DVDD.n1805 VSS 0.279212f
C18900 DVDD.n1806 VSS 0.279212f
C18901 DVDD.n1807 VSS 0.262499f
C18902 DVDD.n1808 VSS 0.279212f
C18903 DVDD.n1809 VSS 0.279212f
C18904 DVDD.n1810 VSS 0.279212f
C18905 DVDD.n1811 VSS 0.279212f
C18906 DVDD.n1812 VSS 0.279212f
C18907 DVDD.n1813 VSS 0.279212f
C18908 DVDD.n1814 VSS 0.279212f
C18909 DVDD.n1815 VSS 0.279212f
C18910 DVDD.n1816 VSS 0.279212f
C18911 DVDD.n1817 VSS 0.214063f
C18912 DVDD.n1818 VSS 0.214063f
C18913 DVDD.n1819 VSS 0.148913f
C18914 DVDD.n1820 VSS 0.148913f
C18915 DVDD.n1821 VSS 0.148913f
C18916 DVDD.n1822 VSS 0.148913f
C18917 DVDD.n1823 VSS 0.148913f
C18918 DVDD.n1824 VSS 0.148913f
C18919 DVDD.n1825 VSS 0.148913f
C18920 DVDD.n1826 VSS 0.148913f
C18921 DVDD.n1827 VSS 0.148913f
C18922 DVDD.n1828 VSS 0.148913f
C18923 DVDD.n1829 VSS 0.434269f
C18924 DVDD.n1830 VSS 0.177581f
C18925 DVDD.n1831 VSS 0.168103f
C18926 DVDD.n1832 VSS 0.148913f
C18927 DVDD.n1833 VSS 0.148913f
C18928 DVDD.n1834 VSS 0.148913f
C18929 DVDD.n1835 VSS 0.148913f
C18930 DVDD.n1836 VSS 0.074652f
C18931 DVDD.n1837 VSS 0.148913f
C18932 DVDD.n1838 VSS 0.148913f
C18933 DVDD.n1839 VSS 0.148913f
C18934 DVDD.n1840 VSS 0.074457f
C18935 DVDD.n1841 VSS 0.074457f
C18936 DVDD.n1842 VSS 0.005305f
C18937 DVDD.n1843 VSS 0.074457f
C18938 DVDD.n1844 VSS 0.279212f
C18939 DVDD.n1845 VSS 0.279212f
C18940 DVDD.n1846 VSS 0.279212f
C18941 DVDD.n1847 VSS 0.279212f
C18942 DVDD.n1848 VSS 0.279212f
C18943 DVDD.n1849 VSS 0.279212f
C18944 DVDD.n1850 VSS 0.279212f
C18945 DVDD.n1851 VSS 0.279212f
C18946 DVDD.n1852 VSS 0.216649f
C18947 DVDD.n1853 VSS 0.279212f
C18948 DVDD.n1854 VSS 0.279212f
C18949 DVDD.n1855 VSS 0.279212f
C18950 DVDD.n1856 VSS 0.139606f
C18951 DVDD.n1861 VSS 0.030281f
C18952 DVDD.t201 VSS 0.513692f
C18953 DVDD.t130 VSS 0.040899f
C18954 DVDD.t139 VSS 0.040899f
C18955 DVDD.n1867 VSS 0.081797f
C18956 DVDD.n1868 VSS 0.1308f
C18957 DVDD.n1869 VSS 0.06758f
C18958 DVDD.t192 VSS 0.040899f
C18959 DVDD.t3 VSS 0.040899f
C18960 DVDD.n1870 VSS 0.081797f
C18961 DVDD.n1871 VSS 0.129754f
C18962 DVDD.t35 VSS 0.0973f
C18963 DVDD.n1872 VSS 0.17088f
C18964 DVDD.t207 VSS 0.031969f
C18965 DVDD.n1873 VSS 0.162851f
C18966 DVDD.t1 VSS 0.0973f
C18967 DVDD.n1874 VSS 0.124781f
C18968 DVDD.n1875 VSS 0.050823f
C18969 DVDD.t17 VSS 0.040899f
C18970 DVDD.t8 VSS 0.040899f
C18971 DVDD.n1876 VSS 0.081797f
C18972 DVDD.n1877 VSS 0.101855f
C18973 DVDD.n1878 VSS 0.056704f
C18974 DVDD.n1879 VSS 0.054497f
C18975 DVDD.n1880 VSS 0.003537f
C18976 DVDD.n1881 VSS 0.010361f
C18977 DVDD.n1882 VSS 0.039153f
C18978 DVDD.n1883 VSS -0.063676f
C18979 DVDD.t7 VSS 0.476895f
C18980 DVDD.t16 VSS 0.476895f
C18981 DVDD.t34 VSS 0.644981f
C18982 DVDD.t2 VSS 0.644981f
C18983 DVDD.t191 VSS 0.379977f
C18984 DVDD.t18 VSS 0.644981f
C18985 DVDD.t48 VSS 0.644981f
C18986 DVDD.t52 VSS 0.476895f
C18987 DVDD.t138 VSS 0.341058f
C18988 DVDD.n1884 VSS 0.497348f
C18989 DVDD.t129 VSS 0.488923f
C18990 DVDD.n1885 VSS 0.501011f
C18991 DVDD.n1886 VSS 0.047009f
C18992 DVDD.n1887 VSS 0.025562f
C18993 DVDD.n1888 VSS 0.037228f
C18994 DVDD.n1889 VSS 0.040159f
C18995 DVDD.n1890 VSS 0.08032f
C18996 DVDD.n1891 VSS 0.08032f
C18997 DVDD.n1892 VSS 0.08032f
C18998 DVDD.n1893 VSS 0.040159f
C18999 DVDD.n1894 VSS 0.040159f
C19000 DVDD.n1895 VSS 0.037228f
C19001 DVDD.n1896 VSS 1.8305f
C19002 DVDD.n1897 VSS 0.951996f
C19003 DVDD.n1898 VSS 0.168643f
C19004 DVDD.n1899 VSS 0.378085f
C19005 DVDD.n1900 VSS 0.346456f
C19006 DVDD.n1901 VSS 0.205477f
C19007 DVDD.n1902 VSS 0.213342f
C19008 DVDD.n1903 VSS 0.027397f
C19009 DVDD.n1904 VSS 0.167294f
C19010 DVDD.n1905 VSS 1.06162f
C19011 DVDD.n1906 VSS 0.279212f
C19012 DVDD.n1907 VSS 0.02661f
C19013 DVDD.n1908 VSS 0.140884f
C19014 DVDD.n1909 VSS 0.027397f
C19015 DVDD.n1910 VSS 0.027397f
C19016 DVDD.n1911 VSS 0.037228f
C19017 DVDD.n1912 VSS 0.037228f
C19018 DVDD.n1913 VSS 0.044999f
C19019 DVDD.n1914 VSS 0.072209f
C19020 DVDD.n1915 VSS 0.082862f
C19021 DVDD.n1916 VSS 0.026381f
C19022 DVDD.t110 VSS 0.020449f
C19023 DVDD.t200 VSS 0.020449f
C19024 DVDD.n1917 VSS 0.077026f
C19025 DVDD.t199 VSS 0.298009f
C19026 DVDD.t68 VSS 0.298001f
C19027 DVDD.t69 VSS 0.020449f
C19028 DVDD.t66 VSS 0.020449f
C19029 DVDD.n1918 VSS 0.077026f
C19030 DVDD.n1919 VSS 0.393109f
C19031 DVDD.n1920 VSS 0.129477f
C19032 DVDD.t65 VSS 0.295113f
C19033 DVDD.n1921 VSS 0.351665f
C19034 DVDD.t109 VSS 0.295113f
C19035 DVDD.n1922 VSS 0.12948f
C19036 DVDD.n1923 VSS 0.39316f
C19037 DVDD.n1924 VSS 0.0253f
C19038 DVDD.n1925 VSS 0.199578f
C19039 DVDD.n1926 VSS 1.06025f
C19040 DVDD.n1927 VSS 0.205477f
C19041 DVDD.n1928 VSS 0.205477f
C19042 DVDD.n1929 VSS 0.279212f
C19043 DVDD.n1930 VSS 0.279212f
C19044 DVDD.n1931 VSS 0.361182f
C19045 DVDD.n1932 VSS 0.509923f
C19046 DVDD.n1933 VSS 0.647968f
C19047 DVDD.n1934 VSS 0.037471f
C19048 DVDD.n1935 VSS 0.032863f
C19049 DVDD.n1936 VSS 0.626283f
C19050 DVDD.n1937 VSS 0.509735f
C19051 DVDD.n1938 VSS 0.361156f
C19052 DVDD.n1939 VSS 0.199578f
C19053 DVDD.n1940 VSS 0.279212f
C19054 DVDD.n1941 VSS 0.205477f
C19055 DVDD.n1942 VSS 0.205477f
C19056 DVDD.n1943 VSS 0.205477f
C19057 DVDD.n1944 VSS 0.213342f
C19058 DVDD.n1945 VSS 0.168096f
C19059 DVDD.n1946 VSS 0.167294f
C19060 DVDD.n1947 VSS 1.06025f
C19061 DVDD.n1948 VSS 0.205477f
C19062 DVDD.n1949 VSS 0.279212f
C19063 DVDD.n1950 VSS 0.199578f
C19064 DVDD.t45 VSS 0.297985f
C19065 DVDD.t46 VSS 0.020449f
C19066 DVDD.t174 VSS 0.020449f
C19067 DVDD.n1951 VSS 0.077026f
C19068 DVDD.n1952 VSS 0.396871f
C19069 DVDD.n1953 VSS 0.132045f
C19070 DVDD.t173 VSS 0.295084f
C19071 DVDD.n1954 VSS 0.347213f
C19072 DVDD.t194 VSS 0.020449f
C19073 DVDD.t156 VSS 0.020449f
C19074 DVDD.n1955 VSS 0.077026f
C19075 DVDD.t155 VSS 0.298037f
C19076 DVDD.t193 VSS 0.295113f
C19077 DVDD.n1956 VSS 0.129423f
C19078 DVDD.n1957 VSS 0.392083f
C19079 DVDD.n1958 VSS 0.028747f
C19080 DVDD.n1959 VSS 0.050484f
C19081 DVDD.n1960 VSS 0.676854f
C19082 DVDD.n1961 VSS 0.509923f
C19083 DVDD.n1962 VSS 0.361182f
C19084 DVDD.n1963 VSS 0.279212f
C19085 DVDD.n1964 VSS 0.205477f
C19086 DVDD.n1965 VSS 0.205477f
C19087 DVDD.n1966 VSS 0.213342f
C19088 DVDD.n1967 VSS 0.168096f
C19089 DVDD.n1968 VSS 0.061371f
C19090 DVDD.n1969 VSS 0.279212f
C19091 DVDD.n1970 VSS 0.279212f
C19092 DVDD.n1971 VSS 0.279212f
C19093 DVDD.n1972 VSS 0.279212f
C19094 DVDD.n1973 VSS 0.448313f
C19095 DVDD.n1974 VSS 0.448313f
C19096 DVDD.n1975 VSS 0.130873f
C19097 DVDD.n1976 VSS 0.279212f
C19098 DVDD.n1977 VSS 0.213342f
C19099 DVDD.n1978 VSS 0.213342f
C19100 DVDD.n1979 VSS 0.139606f
C19101 DVDD.n1980 VSS 0.110112f
C19102 DVDD.n1981 VSS 0.037585f
C19103 DVDD.n1982 VSS 0.168098f
C19104 DVDD.n1983 VSS 0.078651f
C19105 DVDD.n1984 VSS 0.342823f
C19106 DVDD.n1985 VSS 0.344401f
C19107 DVDD.n1986 VSS 0.168635f
C19108 DVDD.n1987 VSS 0.168098f
C19109 DVDD.n1988 VSS 0.168635f
C19110 DVDD.n1989 VSS 0.168098f
C19111 DVDD.n1990 VSS 0.078651f
C19112 DVDD.n1991 VSS 0.06587f
C19113 DVDD.n1992 VSS 0.078651f
C19114 DVDD.n1993 VSS 0.06587f
C19115 DVDD.n1994 VSS 0.168635f
C19116 DVDD.n1995 VSS 0.06587f
C19117 DVDD.n1996 VSS 0.076685f
C19118 DVDD.n1997 VSS 0.378077f
C19119 DVDD.n1998 VSS 1.16281f
C19120 DVDD.n1999 VSS 0.213342f
C19121 DVDD.n2000 VSS 0.205477f
C19122 DVDD.n2001 VSS 0.205477f
C19123 DVDD.n2002 VSS 0.213342f
C19124 DVDD.n2003 VSS 0.213342f
C19125 DVDD.n2004 VSS 0.205477f
C19126 DVDD.n2005 VSS 0.279212f
C19127 DVDD.n2006 VSS 0.279212f
C19128 DVDD.n2007 VSS 0.139606f
C19129 DVDD.n2008 VSS 0.122893f
C19130 DVDD.n2009 VSS 0.009001f
C19131 DVDD.n2010 VSS 0.069733f
C19132 DVDD.t213 VSS 0.155477f
C19133 DVDD.n2011 VSS 0.1204f
C19134 DVDD.n2012 VSS 0.009001f
C19135 DVDD.n2013 VSS 0.069733f
C19136 DVDD.t215 VSS 0.155477f
C19137 DVDD.n2014 VSS 0.1204f
C19138 DVDD.n2015 VSS 0.018792f
C19139 DVDD.n2016 VSS 0.139606f
C19140 DVDD.n2017 VSS 0.464043f
C19141 DVDD.n2018 VSS 0.279212f
C19142 DVDD.n2019 VSS 0.279212f
C19143 DVDD.n2020 VSS 0.279212f
C19144 DVDD.n2021 VSS 0.279212f
C19145 DVDD.n2022 VSS 3.86077f
C19146 DVDD.n2023 VSS 1.3987f
C19147 DVDD.n2024 VSS 0.350073f
C19148 DVDD.n2025 VSS 0.37809f
C19149 DVDD.n2026 VSS 0.073736f
C19150 DVDD.n2027 VSS 0.139606f
C19151 DVDD.n2028 VSS 0.279212f
C19152 DVDD.n2029 VSS 0.279212f
C19153 DVDD.n2030 VSS 0.139606f
C19154 DVDD.n2031 VSS 0.139606f
C19155 DVDD.n2032 VSS 0.139606f
C19156 DVDD.n2033 VSS 0.464043f
C19157 DVDD.n2034 VSS 0.279212f
C19158 DVDD.n2035 VSS 0.139606f
C19159 DVDD.n2036 VSS 0.139606f
C19160 DVDD.n2037 VSS 0.139606f
C19161 DVDD.n2038 VSS 0.139606f
C19162 DVDD.n2039 VSS 0.007073f
C19163 DVDD.n2040 VSS 0.005305f
C19164 DVDD.n2041 VSS 0.007073f
C19165 DVDD.n2042 VSS 0.139606f
C19166 DVDD.n2043 VSS 0.279212f
C19167 DVDD.n2044 VSS 0.26569f
C19168 DVDD.n2045 VSS 0.279212f
C19169 DVDD.n2046 VSS 0.139606f
C19170 DVDD.n2047 VSS 0.265587f
C19171 DVDD.n2048 VSS 0.012307f
C19172 DVDD.n2049 VSS 0.139606f
C19173 DVDD.n2050 VSS 0.139606f
C19174 DVDD.n2051 VSS 0.139606f
C19175 DVDD.n2052 VSS 0.279212f
C19176 DVDD.n2053 VSS 0.793212f
C19177 DVDD.n2054 VSS 0.279212f
C19178 DVDD.n2055 VSS 0.213342f
C19179 DVDD.n2056 VSS 0.213342f
C19180 DVDD.n2057 VSS 0.139606f
C19181 DVDD.n2058 VSS 0.139606f
C19182 DVDD.n2059 VSS 0.007073f
C19183 DVDD.n2060 VSS 0.005305f
C19184 DVDD.n2061 VSS 0.139606f
C19185 DVDD.n2062 VSS 0.012307f
C19186 DVDD.n2063 VSS 0.139802f
C19187 DVDD.n2064 VSS 0.316572f
C19188 DVDD.n2065 VSS 0.324633f
C19189 DVDD.n2066 VSS 0.139606f
C19190 DVDD.n2067 VSS 0.012307f
C19191 DVDD.n2068 VSS 0.139606f
C19192 DVDD.n2069 VSS 0.007073f
C19193 DVDD.n2070 VSS 0.139606f
C19194 DVDD.n2071 VSS 0.139606f
C19195 DVDD.n2072 VSS 0.007073f
C19196 DVDD.n2073 VSS 0.005305f
C19197 DVDD.n2074 VSS 0.003537f
C19198 DVDD.n2075 VSS 0.071443f
C19199 DVDD.n2076 VSS 0.603443f
C19200 DVDD.n2077 VSS 4.68694f
C19201 DVDD.n2078 VSS 0.1225f
C19202 DVDD.n2079 VSS 0.130299f
C19203 DVDD.n2080 VSS 0.130299f
C19204 DVDD.n2081 VSS 0.130299f
C19205 DVDD.n2082 VSS 0.130299f
C19206 DVDD.n2083 VSS 0.130299f
C19207 DVDD.n2084 VSS 0.130299f
C19208 DVDD.n2085 VSS 0.130299f
C19209 DVDD.n2086 VSS 0.130299f
C19210 DVDD.n2087 VSS 0.130299f
C19211 DVDD.n2088 VSS 0.06515f
C19212 DVDD.n2089 VSS 0.031535f
C19213 DVDD.n2090 VSS 0.014157f
C19214 DVDD.n2091 VSS 0.014157f
C19215 DVDD.n2092 VSS 0.014157f
C19216 DVDD.n2093 VSS 0.014157f
C19217 DVDD.n2094 VSS 0.014157f
C19218 DVDD.n2095 VSS 0.014157f
C19219 DVDD.n2096 VSS 0.027266f
C19220 DVDD.n2097 VSS 0.06515f
C19221 DVDD.n2098 VSS 0.018614f
C19222 DVDD.n2099 VSS 0.124335f
C19223 DVDD.n2100 VSS 0.130299f
C19224 DVDD.n2101 VSS 0.130299f
C19225 DVDD.n2102 VSS 0.130299f
C19226 DVDD.n2103 VSS 0.130299f
C19227 DVDD.n2104 VSS 0.130299f
C19228 DVDD.n2105 VSS 0.130299f
C19229 DVDD.n2106 VSS 0.130299f
C19230 DVDD.n2107 VSS 0.130299f
C19231 DVDD.n2108 VSS 0.130299f
C19232 DVDD.n2109 VSS 0.130299f
C19233 DVDD.n2110 VSS 0.130299f
C19234 DVDD.n2111 VSS 0.130299f
C19235 DVDD.n2112 VSS 0.130299f
C19236 DVDD.n2113 VSS 0.130299f
C19237 DVDD.n2114 VSS 0.130299f
C19238 DVDD.n2115 VSS 0.130299f
C19239 DVDD.n2116 VSS 0.130299f
C19240 DVDD.n2117 VSS 0.130299f
C19241 DVDD.n2118 VSS 0.130299f
C19242 DVDD.n2119 VSS 0.130299f
C19243 DVDD.n2120 VSS 0.130299f
C19244 DVDD.n2121 VSS 0.130299f
C19245 DVDD.n2122 VSS 0.130299f
C19246 DVDD.n2123 VSS 0.130299f
C19247 DVDD.n2124 VSS 0.130299f
C19248 DVDD.n2125 VSS 0.130299f
C19249 DVDD.n2126 VSS 0.130299f
C19250 DVDD.n2127 VSS 0.130299f
C19251 DVDD.n2128 VSS 0.130299f
C19252 DVDD.n2129 VSS 0.130299f
C19253 DVDD.n2130 VSS 0.130299f
C19254 DVDD.n2131 VSS 0.130299f
C19255 DVDD.n2132 VSS 0.130299f
C19256 DVDD.n2133 VSS 0.130299f
C19257 DVDD.n2134 VSS 0.130299f
C19258 DVDD.n2135 VSS 0.130299f
C19259 DVDD.n2136 VSS 0.06515f
C19260 DVDD.n2137 VSS 0.130299f
C19261 DVDD.n2138 VSS 0.130299f
C19262 DVDD.n2139 VSS 0.130299f
C19263 DVDD.n2140 VSS 0.130299f
C19264 DVDD.n2141 VSS 0.130299f
C19265 DVDD.n2142 VSS 0.130299f
C19266 DVDD.n2143 VSS 0.130299f
C19267 DVDD.n2144 VSS 0.130299f
C19268 DVDD.n2145 VSS 0.130299f
C19269 DVDD.n2146 VSS 0.130299f
C19270 DVDD.n2147 VSS 0.130299f
C19271 DVDD.n2148 VSS 0.130299f
C19272 DVDD.n2149 VSS 0.130299f
C19273 DVDD.n2150 VSS 0.130299f
C19274 DVDD.n2151 VSS 0.130299f
C19275 DVDD.n2152 VSS 0.130299f
C19276 DVDD.n2153 VSS 0.130299f
C19277 DVDD.n2154 VSS 0.130299f
C19278 DVDD.n2155 VSS 0.130299f
C19279 DVDD.n2156 VSS 0.130299f
C19280 DVDD.n2157 VSS 0.130299f
C19281 DVDD.n2158 VSS 0.130299f
C19282 DVDD.n2159 VSS 0.130299f
C19283 DVDD.n2160 VSS 0.130299f
C19284 DVDD.n2161 VSS 0.130299f
C19285 DVDD.n2162 VSS 0.130299f
C19286 DVDD.n2163 VSS 0.130299f
C19287 DVDD.n2164 VSS 0.130299f
C19288 DVDD.n2165 VSS 0.130299f
C19289 DVDD.n2166 VSS 0.130299f
C19290 DVDD.n2167 VSS 0.130299f
C19291 DVDD.n2168 VSS 0.06515f
C19292 DVDD.n2169 VSS 0.037228f
C19293 DVDD.n2170 VSS 0.037228f
C19294 DVDD.n2171 VSS 0.037228f
C19295 DVDD.n2172 VSS 0.037228f
C19296 DVDD.n2173 VSS 0.037228f
C19297 DVDD.n2174 VSS 0.075864f
C19298 DVDD.n2175 VSS 0.040159f
C19299 DVDD.n2176 VSS 0.228989f
C19300 DVDD.n2177 VSS 0.08032f
C19301 DVDD.n2178 VSS 0.08032f
C19302 DVDD.n2179 VSS 0.040159f
C19303 DVDD.n2180 VSS 0.021211f
C19304 DVDD.n2181 VSS 0.061371f
C19305 DVDD.n2182 VSS 0.040159f
C19306 DVDD.n2183 VSS 0.040159f
C19307 DVDD.n2184 VSS 0.037228f
C19308 DVDD.n2185 VSS 0.037228f
C19309 DVDD.n2186 VSS 0.040159f
C19310 DVDD.n2187 VSS 0.040159f
C19311 DVDD.n2188 VSS 0.08032f
C19312 DVDD.n2189 VSS 0.08032f
C19313 DVDD.n2190 VSS 0.040159f
C19314 DVDD.n2191 VSS 0.076101f
C19315 DVDD.n2192 VSS 0.690035f
C19316 DVDD.n2193 VSS 0.690035f
C19317 DVDD.n2194 VSS 0.037228f
C19318 DVDD.n2195 VSS 0.037228f
C19319 DVDD.n2196 VSS 0.037228f
C19320 DVDD.n2197 VSS 0.037228f
C19321 DVDD.n2198 VSS 0.06515f
C19322 DVDD.n2200 VSS 0.06515f
C19323 DVDD.n2201 VSS 0.037228f
C19324 DVDD.n2202 VSS 0.037228f
C19325 DVDD.n2203 VSS 0.037228f
C19326 DVDD.n2204 VSS 0.037228f
C19327 DVDD.n2205 VSS 0.072949f
C19328 DVDD.n2207 VSS 0.037228f
C19329 DVDD.n2209 VSS 0.037228f
C19330 DVDD.n2211 VSS 0.037228f
C19331 DVDD.n2213 VSS 0.037228f
C19332 DVDD.t220 VSS 0.142962f
C19333 DVDD.n2214 VSS 0.064841f
C19334 DVDD.n2215 VSS 0.22817f
C19335 DVDD.t210 VSS 0.142962f
C19336 DVDD.n2216 VSS 0.07475f
C19337 DVDD.n2217 VSS 0.07475f
C19338 DVDD.n2218 VSS 0.106179f
C19339 DVDD.n2219 VSS 0.106179f
C19340 DVDD.t217 VSS 0.142962f
C19341 DVDD.n2220 VSS 0.07475f
C19342 DVDD.n2221 VSS 0.07475f
C19343 DVDD.n2222 VSS 0.106179f
C19344 DVDD.n2223 VSS 0.106179f
C19345 DVDD.t206 VSS 0.142962f
C19346 DVDD.n2224 VSS 0.07475f
C19347 DVDD.n2225 VSS 0.07475f
C19348 DVDD.n2226 VSS 0.106179f
C19349 DVDD.n2227 VSS 0.106179f
C19350 DVDD.t216 VSS 0.142962f
C19351 DVDD.n2228 VSS 0.07475f
C19352 DVDD.n2229 VSS 0.07475f
C19353 DVDD.n2230 VSS 0.106179f
C19354 DVDD.n2231 VSS 0.106179f
C19355 DVDD.t211 VSS 0.142962f
C19356 DVDD.n2232 VSS 0.07475f
C19357 DVDD.n2233 VSS 0.07475f
C19358 DVDD.n2234 VSS 0.106179f
C19359 DVDD.n2235 VSS 0.106179f
C19360 DVDD.t218 VSS 0.142962f
C19361 DVDD.n2236 VSS 0.07475f
C19362 DVDD.n2237 VSS 0.07475f
C19363 DVDD.n2238 VSS 0.146793f
C19364 DVDD.n2239 VSS 0.086235f
C19365 DVDD.t208 VSS 0.142962f
C19366 DVDD.n2240 VSS 0.248931f
C19367 DVDD.n2244 VSS 0.130299f
C19368 DVDD.n2245 VSS 0.130299f
C19369 DVDD.n2246 VSS 0.130299f
C19370 DVDD.n2247 VSS 0.130299f
C19371 DVDD.n2248 VSS 0.130299f
C19372 DVDD.n2249 VSS 0.130299f
C19373 DVDD.n2250 VSS 0.130299f
C19374 DVDD.n2251 VSS 0.130299f
C19375 DVDD.n2252 VSS 0.130299f
C19376 DVDD.n2253 VSS 0.130299f
C19377 DVDD.n2254 VSS 0.130299f
C19378 DVDD.n2255 VSS 0.089384f
C19379 DVDD.n2256 VSS 0.130299f
C19380 DVDD.n2257 VSS 0.130299f
C19381 DVDD.n2258 VSS 0.130299f
C19382 DVDD.n2259 VSS 0.068361f
C19383 DVDD.n2260 VSS 0.112406f
C19384 DVDD.n2261 VSS -0.005423f
C19385 DVDD.t136 VSS 0.232386f
C19386 DVDD.n2262 VSS 0.018124f
C19387 DVDD.n2263 VSS 0.083502f
C19388 DVDD.n2264 VSS 0.085002f
C19389 DVDD.n2265 VSS 0.130299f
C19390 DVDD.n2266 VSS 0.130299f
C19391 DVDD.n2267 VSS 0.130299f
C19392 DVDD.n2268 VSS 0.130299f
C19393 DVDD.n2269 VSS 0.08396f
C19394 DVDD.n2270 VSS 0.130299f
C19395 DVDD.n2271 VSS 0.130299f
C19396 DVDD.n2272 VSS 0.130299f
C19397 DVDD.n2273 VSS 0.130299f
C19398 DVDD.t89 VSS 0.010225f
C19399 DVDD.t93 VSS 0.010225f
C19400 DVDD.n2274 VSS 0.02257f
C19401 DVDD.n2275 VSS 0.049642f
C19402 DVDD.n2276 VSS 0.085002f
C19403 DVDD.n2277 VSS 0.111488f
C19404 DVDD.n2278 VSS 0.130299f
C19405 DVDD.n2279 VSS 0.130299f
C19406 DVDD.n2280 VSS 0.130299f
C19407 DVDD.n2281 VSS 0.130299f
C19408 DVDD.n2282 VSS 0.130299f
C19409 DVDD.n2283 VSS 0.130299f
C19410 DVDD.n2284 VSS 0.130299f
C19411 DVDD.n2285 VSS 0.01614f
C19412 DVDD.t95 VSS 0.026048f
C19413 DVDD.n2286 VSS 0.060321f
C19414 DVDD.n2287 VSS 0.085002f
C19415 DVDD.n2288 VSS 0.074784f
C19416 DVDD.n2289 VSS 0.130299f
C19417 DVDD.n2290 VSS 0.130299f
C19418 DVDD.n2291 VSS 0.130299f
C19419 DVDD.n2292 VSS 0.130299f
C19420 DVDD.n2293 VSS 0.130299f
C19421 DVDD.n2294 VSS 0.08396f
C19422 DVDD.n2295 VSS 0.085002f
C19423 DVDD.n2296 VSS 0.130299f
C19424 DVDD.n2297 VSS 0.130299f
C19425 DVDD.n2298 VSS 0.130299f
C19426 DVDD.n2299 VSS 0.120664f
C19427 DVDD.n2300 VSS 0.086254f
C19428 DVDD.n2301 VSS 0.130299f
C19429 DVDD.n2302 VSS 0.130299f
C19430 DVDD.n2303 VSS 0.130299f
C19431 DVDD.n2304 VSS 0.130299f
C19432 DVDD.n2305 VSS 0.130299f
C19433 DVDD.n2306 VSS 0.130299f
C19434 DVDD.n2307 VSS 0.130299f
C19435 DVDD.n2308 VSS 0.130299f
C19436 DVDD.n2309 VSS 0.130299f
C19437 DVDD.n2310 VSS 0.130299f
C19438 DVDD.n2311 VSS 0.130299f
C19439 DVDD.n2312 VSS 0.130299f
C19440 DVDD.n2313 VSS 0.130299f
C19441 DVDD.n2314 VSS 0.130299f
C19442 DVDD.n2315 VSS 0.130299f
C19443 DVDD.n2316 VSS 0.130299f
C19444 DVDD.n2317 VSS 0.130299f
C19445 DVDD.n2318 VSS 0.130299f
C19446 DVDD.n2319 VSS 0.1225f
C19447 DVDD.n2320 VSS 0.130299f
C19448 DVDD.n2321 VSS 0.130299f
C19449 DVDD.n2322 VSS 0.130299f
C19450 DVDD.n2323 VSS 0.089384f
C19451 DVDD.n2324 VSS 0.116994f
C19452 DVDD.n2325 VSS -0.005423f
C19453 DVDD.t187 VSS 0.232386f
C19454 DVDD.n2326 VSS 0.018124f
C19455 DVDD.n2327 VSS 0.083502f
C19456 DVDD.n2328 VSS 0.085002f
C19457 DVDD.n2329 VSS 0.130299f
C19458 DVDD.n2330 VSS 0.130299f
C19459 DVDD.n2331 VSS 0.130299f
C19460 DVDD.n2332 VSS 0.130299f
C19461 DVDD.n2333 VSS 0.088548f
C19462 DVDD.n2334 VSS 0.130299f
C19463 DVDD.n2335 VSS 0.130299f
C19464 DVDD.n2336 VSS 0.130299f
C19465 DVDD.n2337 VSS 0.130299f
C19466 DVDD.n2338 VSS 0.130299f
C19467 DVDD.n2339 VSS 0.130299f
C19468 DVDD.t77 VSS 0.010225f
C19469 DVDD.t119 VSS 0.010225f
C19470 DVDD.n2340 VSS 0.02257f
C19471 DVDD.n2341 VSS 0.049642f
C19472 DVDD.n2342 VSS 0.085002f
C19473 DVDD.n2343 VSS 0.1069f
C19474 DVDD.n2344 VSS 0.130299f
C19475 DVDD.n2345 VSS 0.130299f
C19476 DVDD.n2346 VSS 0.130299f
C19477 DVDD.n2347 VSS 0.130299f
C19478 DVDD.n2348 VSS 0.130299f
C19479 DVDD.n2349 VSS 0.130299f
C19480 DVDD.n2350 VSS 0.130299f
C19481 DVDD.n2351 VSS 0.01614f
C19482 DVDD.t85 VSS 0.026048f
C19483 DVDD.n2352 VSS 0.060321f
C19484 DVDD.n2353 VSS 0.085002f
C19485 DVDD.n2354 VSS 0.070196f
C19486 DVDD.n2355 VSS 0.130299f
C19487 DVDD.n2356 VSS 0.130299f
C19488 DVDD.n2357 VSS 0.130299f
C19489 DVDD.n2358 VSS 0.130299f
C19490 DVDD.n2359 VSS 0.130299f
C19491 DVDD.n2360 VSS 0.088548f
C19492 DVDD.n2361 VSS 0.085002f
C19493 DVDD.n2362 VSS 0.130299f
C19494 DVDD.n2363 VSS 0.130299f
C19495 DVDD.n2364 VSS 0.130299f
C19496 DVDD.n2365 VSS 0.125252f
C19497 DVDD.n2366 VSS 0.086254f
C19498 DVDD.n2367 VSS 0.130299f
C19499 DVDD.n2368 VSS 0.130299f
C19500 DVDD.n2369 VSS 0.130299f
C19501 DVDD.n2370 VSS 0.130299f
C19502 DVDD.n2371 VSS 0.130299f
C19503 DVDD.n2372 VSS 0.130299f
C19504 DVDD.n2373 VSS 0.130299f
C19505 DVDD.n2374 VSS 0.130299f
C19506 DVDD.n2375 VSS 0.130299f
C19507 DVDD.n2376 VSS 0.130299f
C19508 DVDD.n2377 VSS 0.130299f
C19509 DVDD.n2378 VSS 0.130299f
C19510 DVDD.n2379 VSS 0.130299f
C19511 DVDD.n2380 VSS 0.130299f
C19512 DVDD.n2381 VSS 0.130299f
C19513 DVDD.n2382 VSS 0.130299f
C19514 DVDD.n2383 VSS 0.130299f
C19515 DVDD.n2384 VSS 0.130299f
C19516 DVDD.n2385 VSS 0.130299f
C19517 DVDD.n2386 VSS 0.130299f
C19518 DVDD.n2387 VSS 0.130299f
C19519 DVDD.n2388 VSS 0.130299f
C19520 DVDD.n2389 VSS 0.130299f
C19521 DVDD.n2390 VSS 0.130299f
C19522 DVDD.n2391 VSS 0.130299f
C19523 DVDD.n2392 VSS 0.130299f
C19524 DVDD.n2393 VSS 0.130299f
C19525 DVDD.n2394 VSS 0.130299f
C19526 DVDD.n2395 VSS 0.117453f
C19527 DVDD.n2396 VSS 0.117453f
C19528 DVDD.n2397 VSS 0.014682f
C19529 DVDD.n2398 VSS 0.171513f
C19530 DVDD.n2399 VSS 0.627997f
C19531 DVDD.n2400 VSS 0.117453f
C19532 DVDD.n2401 VSS 0.130299f
C19533 DVDD.n2402 VSS 0.130299f
C19534 DVDD.n2403 VSS 0.130299f
C19535 DVDD.n2404 VSS 0.130299f
C19536 DVDD.n2405 VSS 0.130299f
C19537 DVDD.n2406 VSS 0.130299f
C19538 DVDD.n2407 VSS 0.130299f
C19539 DVDD.n2408 VSS 0.130299f
C19540 DVDD.n2409 VSS 0.130299f
C19541 DVDD.n2410 VSS 0.130299f
C19542 DVDD.n2411 VSS 0.130299f
C19543 DVDD.n2412 VSS 0.130299f
C19544 DVDD.n2413 VSS 0.130299f
C19545 DVDD.n2414 VSS 0.130299f
C19546 DVDD.n2415 VSS 0.130299f
C19547 DVDD.n2416 VSS 0.130299f
C19548 DVDD.n2417 VSS 0.130299f
C19549 DVDD.n2418 VSS 0.130299f
C19550 DVDD.n2419 VSS 0.130299f
C19551 DVDD.n2420 VSS 0.130299f
C19552 DVDD.n2421 VSS 0.130299f
C19553 DVDD.n2422 VSS 0.130299f
C19554 DVDD.n2423 VSS 0.130299f
C19555 DVDD.n2424 VSS 0.130299f
C19556 DVDD.n2425 VSS 0.130299f
C19557 DVDD.n2426 VSS 0.130299f
C19558 DVDD.n2427 VSS 0.130299f
C19559 DVDD.n2428 VSS 0.130299f
C19560 DVDD.n2429 VSS 0.130299f
C19561 DVDD.n2430 VSS 0.130299f
C19562 DVDD.n2431 VSS 0.130299f
C19563 DVDD.n2432 VSS 0.130299f
C19564 DVDD.n2433 VSS 0.130299f
C19565 DVDD.n2434 VSS 0.130299f
C19566 DVDD.n2435 VSS 0.130299f
C19567 DVDD.n2436 VSS 0.130299f
C19568 DVDD.n2437 VSS 0.130299f
C19569 DVDD.n2438 VSS 0.130299f
C19570 DVDD.n2439 VSS 0.130299f
C19571 DVDD.n2440 VSS 0.130299f
C19572 DVDD.n2441 VSS 0.130299f
C19573 DVDD.n2442 VSS 0.130299f
C19574 DVDD.n2443 VSS 0.130299f
C19575 DVDD.n2444 VSS 0.130299f
C19576 DVDD.n2445 VSS 0.130299f
C19577 DVDD.n2446 VSS 0.130299f
C19578 DVDD.n2447 VSS 0.130299f
C19579 DVDD.n2448 VSS 0.130299f
C19580 DVDD.n2449 VSS 0.130299f
C19581 DVDD.n2450 VSS 0.130299f
C19582 DVDD.n2451 VSS 0.130299f
C19583 DVDD.n2452 VSS 0.130299f
C19584 DVDD.n2453 VSS 0.130299f
C19585 DVDD.n2454 VSS 0.130299f
C19586 DVDD.n2455 VSS 0.075702f
C19587 DVDD.n2456 VSS 0.089384f
C19588 DVDD.n2457 VSS 0.238761f
C19589 DVDD.t189 VSS 0.155631f
C19590 DVDD.t61 VSS 0.234237f
C19591 DVDD.t195 VSS 0.154783f
C19592 DVDD.n2458 VSS 0.07032f
C19593 DVDD.t190 VSS 0.010225f
C19594 DVDD.t196 VSS 0.010225f
C19595 DVDD.n2459 VSS 0.02257f
C19596 DVDD.n2460 VSS 0.049642f
C19597 DVDD.t188 VSS 0.026048f
C19598 DVDD.n2461 VSS 0.060321f
C19599 DVDD.n2462 VSS 0.01614f
C19600 DVDD.n2463 VSS -0.005423f
C19601 DVDD.n2464 VSS 0.035393f
C19602 DVDD.t62 VSS 0.025964f
C19603 DVDD.n2465 VSS 0.060581f
C19604 DVDD.n2466 VSS 0.085106f
C19605 DVDD.n2467 VSS 0.098642f
C19606 DVDD.n2468 VSS 0.130299f
C19607 DVDD.n2469 VSS 0.130299f
C19608 DVDD.n2470 VSS 0.130299f
C19609 DVDD.n2471 VSS 0.130299f
C19610 DVDD.n2472 VSS 0.130299f
C19611 DVDD.n2473 VSS 0.130299f
C19612 DVDD.n2474 VSS 0.070196f
C19613 DVDD.n2475 VSS 0.130299f
C19614 DVDD.n2476 VSS 0.130299f
C19615 DVDD.n2477 VSS 0.130299f
C19616 DVDD.n2478 VSS 0.130299f
C19617 DVDD.n2479 VSS 0.130299f
C19618 DVDD.n2480 VSS 0.130299f
C19619 DVDD.n2481 VSS 0.130299f
C19620 DVDD.n2482 VSS 0.083502f
C19621 DVDD.n2483 VSS 0.089384f
C19622 DVDD.n2484 VSS 0.028424f
C19623 DVDD.n2485 VSS 0.227451f
C19624 DVDD.t84 VSS 0.232386f
C19625 DVDD.t118 VSS 0.155631f
C19626 DVDD.n2486 VSS 0.07032f
C19627 DVDD.t76 VSS 0.154783f
C19628 DVDD.t78 VSS 0.234237f
C19629 DVDD.n2487 VSS 0.238761f
C19630 DVDD.n2488 VSS 0.035225f
C19631 DVDD.t79 VSS 0.026048f
C19632 DVDD.n2489 VSS 0.060321f
C19633 DVDD.n2490 VSS 0.085002f
C19634 DVDD.n2491 VSS 0.078455f
C19635 DVDD.n2492 VSS 0.072949f
C19636 DVDD.n2493 VSS 0.130299f
C19637 DVDD.n2494 VSS 0.130299f
C19638 DVDD.n2495 VSS 0.130299f
C19639 DVDD.n2496 VSS 0.130299f
C19640 DVDD.n2497 VSS 0.130299f
C19641 DVDD.n2498 VSS 0.130299f
C19642 DVDD.n2499 VSS 0.130299f
C19643 DVDD.n2500 VSS 0.130299f
C19644 DVDD.n2501 VSS 0.130299f
C19645 DVDD.n2502 VSS 0.130299f
C19646 DVDD.n2503 VSS 0.130299f
C19647 DVDD.n2504 VSS 0.130299f
C19648 DVDD.n2505 VSS 0.130299f
C19649 DVDD.n2506 VSS 0.130299f
C19650 DVDD.n2507 VSS 0.130299f
C19651 DVDD.n2508 VSS 0.130299f
C19652 DVDD.n2509 VSS 0.130299f
C19653 DVDD.n2510 VSS 0.130299f
C19654 DVDD.n2511 VSS 0.130299f
C19655 DVDD.n2512 VSS 0.130299f
C19656 DVDD.n2513 VSS 0.130299f
C19657 DVDD.n2514 VSS 0.130299f
C19658 DVDD.n2515 VSS 0.130299f
C19659 DVDD.n2516 VSS 0.130299f
C19660 DVDD.n2517 VSS 0.130299f
C19661 DVDD.n2518 VSS 0.130299f
C19662 DVDD.n2519 VSS 0.130299f
C19663 DVDD.n2520 VSS 0.130299f
C19664 DVDD.n2521 VSS 0.130299f
C19665 DVDD.n2522 VSS 0.130299f
C19666 DVDD.n2523 VSS 0.130299f
C19667 DVDD.n2524 VSS 0.130299f
C19668 DVDD.n2525 VSS 0.130299f
C19669 DVDD.n2526 VSS 0.130299f
C19670 DVDD.n2527 VSS 0.130299f
C19671 DVDD.n2528 VSS 0.130299f
C19672 DVDD.n2529 VSS 0.130299f
C19673 DVDD.n2530 VSS 0.071114f
C19674 DVDD.n2531 VSS 0.089384f
C19675 DVDD.n2532 VSS 0.238761f
C19676 DVDD.t134 VSS 0.155631f
C19677 DVDD.t178 VSS 0.234237f
C19678 DVDD.t180 VSS 0.154783f
C19679 DVDD.n2533 VSS 0.07032f
C19680 DVDD.t135 VSS 0.010225f
C19681 DVDD.t181 VSS 0.010225f
C19682 DVDD.n2534 VSS 0.02257f
C19683 DVDD.n2535 VSS 0.049642f
C19684 DVDD.t137 VSS 0.026048f
C19685 DVDD.n2536 VSS 0.060321f
C19686 DVDD.n2537 VSS 0.01614f
C19687 DVDD.n2538 VSS -0.005423f
C19688 DVDD.n2539 VSS 0.035225f
C19689 DVDD.t179 VSS 0.026048f
C19690 DVDD.n2540 VSS 0.060321f
C19691 DVDD.n2541 VSS 0.085002f
C19692 DVDD.n2542 VSS 0.10323f
C19693 DVDD.n2543 VSS 0.130299f
C19694 DVDD.n2544 VSS 0.130299f
C19695 DVDD.n2545 VSS 0.130299f
C19696 DVDD.n2546 VSS 0.130299f
C19697 DVDD.n2547 VSS 0.130299f
C19698 DVDD.n2548 VSS 0.130299f
C19699 DVDD.n2549 VSS 0.074784f
C19700 DVDD.n2550 VSS 0.130299f
C19701 DVDD.n2551 VSS 0.130299f
C19702 DVDD.n2552 VSS 0.130299f
C19703 DVDD.n2553 VSS 0.130299f
C19704 DVDD.n2554 VSS 0.130299f
C19705 DVDD.n2555 VSS 0.130299f
C19706 DVDD.n2556 VSS 0.130299f
C19707 DVDD.n2557 VSS 0.083502f
C19708 DVDD.n2558 VSS 0.089384f
C19709 DVDD.n2559 VSS 0.028424f
C19710 DVDD.n2560 VSS 0.227451f
C19711 DVDD.t94 VSS 0.232386f
C19712 DVDD.t92 VSS 0.155631f
C19713 DVDD.n2561 VSS 0.07032f
C19714 DVDD.t88 VSS 0.154783f
C19715 DVDD.t167 VSS 0.234237f
C19716 DVDD.n2562 VSS 0.238761f
C19717 DVDD.n2563 VSS 0.035225f
C19718 DVDD.t168 VSS 0.026048f
C19719 DVDD.n2564 VSS 0.060321f
C19720 DVDD.n2565 VSS 0.085002f
C19721 DVDD.n2566 VSS 0.083043f
C19722 DVDD.n2567 VSS 0.130299f
C19723 DVDD.n2568 VSS 0.130299f
C19724 DVDD.n2569 VSS 0.130299f
C19725 DVDD.n2570 VSS 0.130299f
C19726 DVDD.n2571 VSS 0.130299f
C19727 DVDD.n2572 VSS 0.127088f
C19728 DVDD.n2573 VSS 0.130299f
C19729 DVDD.n2574 VSS 0.130299f
C19730 DVDD.n2575 VSS 0.130299f
C19731 DVDD.n2576 VSS 0.130299f
C19732 DVDD.n2577 VSS 0.130299f
C19733 DVDD.n2578 VSS 0.130299f
C19734 DVDD.n2579 VSS 0.130299f
C19735 DVDD.n2580 VSS 0.130299f
C19736 DVDD.n2581 VSS 0.130299f
C19737 DVDD.n2582 VSS 0.130299f
C19738 DVDD.n2583 VSS 0.130299f
C19739 DVDD.n2584 VSS 0.130299f
C19740 DVDD.n2585 VSS 0.130299f
C19741 DVDD.n2586 VSS 0.130299f
C19742 DVDD.n2587 VSS 0.130299f
C19743 DVDD.n2588 VSS 0.130299f
C19744 DVDD.n2589 VSS 0.130299f
C19745 DVDD.n2590 VSS 0.130299f
C19746 DVDD.n2591 VSS 0.130299f
C19747 DVDD.n2592 VSS 0.130299f
C19748 DVDD.n2593 VSS 0.130299f
C19749 DVDD.n2594 VSS 0.482824f
C19750 DVDD.n2595 VSS 0.130299f
C19751 DVDD.n2596 VSS 0.130299f
C19752 DVDD.n2597 VSS 0.06515f
C19753 DVDD.n2598 VSS 0.29091f
C19754 DVDD.n2600 VSS 0.262689f
C19755 DVDD.n2601 VSS 0.06515f
C19756 DVDD.n2602 VSS 0.918001f
C19757 DVDD.n2604 VSS 0.248931f
C19758 DVDD.n2609 VSS 0.06515f
C19759 DVDD.n2610 VSS 0.482824f
C19760 DVDD.n2611 VSS 0.130299f
C19761 DVDD.n2612 VSS 0.130299f
C19762 DVDD.n2613 VSS 0.06515f
C19763 DVDD.n2618 VSS 0.29091f
C19764 DVDD.n2619 VSS 1.00427f
C19765 DVDD.n2620 VSS 0.06515f
C19766 DVDD.n2621 VSS 0.072949f
C19767 DVDD.n2622 VSS 0.130299f
C19768 DVDD.n2623 VSS 0.130299f
C19769 DVDD.n2624 VSS 0.130299f
C19770 DVDD.n2625 VSS 0.130299f
C19771 DVDD.n2626 VSS 0.130299f
C19772 DVDD.n2627 VSS 0.130299f
C19773 DVDD.n2628 VSS 0.130299f
C19774 DVDD.n2629 VSS 0.130299f
C19775 DVDD.n2630 VSS 0.130299f
C19776 DVDD.n2631 VSS 0.130299f
C19777 DVDD.n2632 VSS 0.130299f
C19778 DVDD.n2633 VSS 0.130299f
C19779 DVDD.n2634 VSS 0.130299f
C19780 DVDD.n2635 VSS 0.130299f
C19781 DVDD.n2636 VSS 0.130299f
C19782 DVDD.n2637 VSS 0.130299f
C19783 DVDD.n2638 VSS 0.130299f
C19784 DVDD.n2639 VSS 0.130299f
C19785 DVDD.n2640 VSS 0.130299f
C19786 DVDD.n2641 VSS 0.130299f
C19787 DVDD.n2642 VSS 0.130299f
C19788 DVDD.n2643 VSS 0.130299f
C19789 DVDD.n2644 VSS 0.130299f
C19790 DVDD.n2645 VSS 0.130299f
C19791 DVDD.n2646 VSS 0.130299f
C19792 DVDD.n2647 VSS 0.130299f
C19793 DVDD.n2648 VSS 0.130299f
C19794 DVDD.n2649 VSS 0.130299f
C19795 DVDD.n2650 VSS 0.130299f
C19796 DVDD.n2651 VSS 0.130299f
C19797 DVDD.n2652 VSS 0.130299f
C19798 DVDD.n2653 VSS 0.130299f
C19799 DVDD.n2654 VSS 0.130299f
C19800 DVDD.n2655 VSS 0.130299f
C19801 DVDD.n2656 VSS 0.130299f
C19802 DVDD.n2657 VSS 0.130299f
C19803 DVDD.n2658 VSS 0.130299f
C19804 DVDD.n2659 VSS 0.130299f
C19805 DVDD.n2660 VSS 0.130299f
C19806 DVDD.n2661 VSS 0.130299f
C19807 DVDD.n2662 VSS 0.130299f
C19808 DVDD.n2663 VSS 0.130299f
C19809 DVDD.n2664 VSS 0.130299f
C19810 DVDD.n2665 VSS 0.130299f
C19811 DVDD.n2666 VSS 0.130299f
C19812 DVDD.n2667 VSS 0.130299f
C19813 DVDD.n2668 VSS 0.11837f
C19814 DVDD.t91 VSS 0.026661f
C19815 DVDD.t90 VSS 0.295845f
C19816 DVDD.n2669 VSS 0.2723f
C19817 DVDD.n2670 VSS 0.053935f
C19818 DVDD.n2671 VSS 0.056205f
C19819 DVDD.n2672 VSS 0.081014f
C19820 DVDD.n2673 VSS 0.077078f
C19821 DVDD.n2674 VSS 0.130299f
C19822 DVDD.n2675 VSS 0.130299f
C19823 DVDD.n2676 VSS 0.130299f
C19824 DVDD.n2677 VSS 0.130299f
C19825 DVDD.n2678 VSS 0.130299f
C19826 DVDD.n2679 VSS 0.130299f
C19827 DVDD.n2680 VSS 0.130299f
C19828 DVDD.n2681 VSS 0.072949f
C19829 DVDD.n2682 VSS 0.06515f
C19830 DVDD.n2683 VSS 0.013025f
C19831 DVDD.n2684 VSS 0.013025f
C19832 DVDD.n2685 VSS 0.013025f
C19833 DVDD.n2686 VSS 0.013025f
C19834 DVDD.n2687 VSS 0.013025f
C19835 DVDD.n2688 VSS 0.06515f
C19836 DVDD.n2689 VSS 0.013025f
C19837 DVDD.n2690 VSS 0.013025f
C19838 DVDD.n2691 VSS 0.013025f
C19839 DVDD.n2692 VSS 0.013025f
C19840 DVDD.n2693 VSS -0.346392f
C19841 DVDD.n2695 VSS 0.017125f
C19842 DVDD.n2696 VSS 0.004429f
C19843 DVDD.n2697 VSS 0.032509f
C19844 DVDD.n2698 VSS 0.029909f
C19845 DVDD.n2699 VSS 0.032509f
C19846 DVDD.n2700 VSS 0.021467f
C19847 DVDD.n2702 VSS 0.17926f
C19848 DVDD.n2703 VSS 0.021467f
C19849 DVDD.n2704 VSS 0.032509f
C19850 DVDD.n2705 VSS 0.111895f
C19851 DVDD.n2706 VSS 0.651329f
C19852 DVDD.t55 VSS 0.010134f
C19853 DVDD.n2707 VSS 0.032098f
C19854 DVDD.n2708 VSS 0.115362f
C19855 DVDD.t12 VSS 0.006476f
C19856 DVDD.t10 VSS 0.006476f
C19857 DVDD.n2709 VSS 0.019733f
C19858 DVDD.t71 VSS 0.009347f
C19859 DVDD.t73 VSS 0.006816f
C19860 DVDD.t75 VSS 0.006816f
C19861 DVDD.n2710 VSS 0.029157f
C19862 DVDD.n2711 VSS 0.049055f
C19863 DVDD.t154 VSS 0.016089f
C19864 DVDD.n2712 VSS 0.028852f
C19865 DVDD.n2713 VSS 0.043311f
C19866 DVDD.n2714 VSS 0.142981f
C19867 DVDD.t29 VSS 0.180818f
C19868 DVDD.n2715 VSS 0.110895f
C19869 DVDD.t30 VSS 0.013014f
C19870 DVDD.n2716 VSS 0.322657f
C19871 DVDD.n2717 VSS 0.277723f
C19872 DVDD.n2718 VSS 0.303782f
C19873 DVDD.t60 VSS 0.358809f
C19874 DVDD.t67 VSS 0.491912f
C19875 DVDD.t175 VSS 0.430847f
C19876 DVDD.t182 VSS 0.268007f
C19877 DVDD.t4 VSS 0.268007f
C19878 DVDD.t13 VSS 0.368086f
C19879 DVDD.t11 VSS 0.344338f
C19880 DVDD.n2719 VSS 0.074163f
C19881 DVDD.n2720 VSS 0.047033f
C19882 DVDD.n2721 VSS 0.047033f
C19883 DVDD.n2722 VSS 0.034823f
C19884 DVDD.n2723 VSS 0.047033f
C19885 DVDD.n2725 VSS 0.047033f
C19886 DVDD.n2726 VSS 0.023517f
C19887 DVDD.n2727 VSS 0.088896f
C19888 DVDD.n2728 VSS 0.047033f
C19889 DVDD.n2733 VSS 0.062848f
C19890 DVDD.t152 VSS 0.051574f
C19891 DVDD.t83 VSS 0.051574f
C19892 DVDD.t117 VSS 0.016089f
C19893 DVDD.n2734 VSS 0.046162f
C19894 DVDD.n2735 VSS 0.045326f
C19895 DVDD.n2736 VSS 0.045095f
C19896 DVDD.n2737 VSS 0.062848f
C19897 DVDD.n2740 VSS 0.03408f
C19898 DVDD.n2742 VSS 0.074163f
C19899 DVDD.n2743 VSS 0.053168f
C19900 DVDD.n2744 VSS 0.053168f
C19901 DVDD.n2745 VSS 0.053168f
C19902 DVDD.n2746 VSS 0.053168f
C19903 DVDD.n2748 VSS 0.053168f
C19904 DVDD.n2749 VSS 0.053168f
C19905 DVDD.n2751 VSS 0.062848f
C19906 DVDD.n2752 VSS 0.062848f
C19907 DVDD.n2755 VSS 0.062848f
C19908 DVDD.n2759 VSS 0.062848f
C19909 DVDD.n2764 VSS 0.186043f
C19910 DVDD.n2768 VSS 0.043966f
C19911 DVDD.n2769 VSS 0.062848f
C19912 DVDD.n2770 VSS 0.075096f
C19913 DVDD.n2771 VSS 0.074163f
C19914 DVDD.n2772 VSS 0.074163f
C19915 DVDD.n2773 VSS 0.074163f
C19916 DVDD.n2774 VSS 0.074163f
C19917 DVDD.n2775 VSS 0.062848f
C19918 DVDD.n2776 VSS 0.043966f
C19919 DVDD.n2777 VSS 0.062848f
C19920 DVDD.n2778 VSS 0.074163f
C19921 DVDD.n2779 VSS 0.074163f
C19922 DVDD.n2783 VSS 0.062848f
C19923 DVDD.n2784 VSS 0.074163f
C19924 DVDD.n2785 VSS 0.074163f
C19925 DVDD.n2786 VSS 0.062848f
C19926 DVDD.n2787 VSS 0.04857f
C19927 DVDD.n2788 VSS 0.058618f
C19928 DVDD.n2789 VSS 0.097537f
C19929 DVDD.n2790 VSS 0.236694f
C19930 DVDD.t151 VSS 0.256217f
C19931 DVDD.t82 VSS 0.495812f
C19932 DVDD.t116 VSS 0.513115f
C19933 DVDD.t153 VSS 0.295147f
C19934 DVDD.t70 VSS 0.295147f
C19935 DVDD.t74 VSS 0.206942f
C19936 DVDD.t72 VSS 0.299388f
C19937 DVDD.t9 VSS 0.219664f
C19938 DVDD.n2791 VSS 0.103471f
C19939 DVDD.n2792 VSS 0.298961f
C19940 DVDD.n2793 VSS 0.029614f
C19941 DVDD.n2794 VSS 0.078728f
C19942 DVDD.n2795 VSS 0.063047f
C19943 DVDD.n2796 VSS 0.319863f
C19944 DVDD.n2797 VSS -0.568215f
C19945 DVDD.n2798 VSS 0.520631f
C19946 DVDD.n2799 VSS 0.31862f
C19947 DVDD.n2800 VSS 0.016884f
C19948 DVDD.n2802 VSS 0.127022f
C19949 DVDD.n2803 VSS 0.031356f
C19950 DVDD.n2804 VSS 0.032509f
C19951 DVDD.n2805 VSS 0.032509f
C19952 DVDD.n2806 VSS 0.032509f
C19953 DVDD.n2807 VSS 0.029909f
C19954 DVDD.n2808 VSS 0.029909f
C19955 DVDD.n2809 VSS 0.029909f
C19956 DVDD.n2810 VSS 0.032509f
C19957 DVDD.n2811 VSS 0.032509f
C19958 DVDD.n2812 VSS 0.032509f
C19959 DVDD.n2813 VSS 0.029909f
C19960 DVDD.n2814 VSS 0.029909f
C19961 DVDD.n2815 VSS 0.029909f
C19962 DVDD.n2816 VSS 0.032509f
C19963 DVDD.n2817 VSS 0.032509f
C19964 DVDD.n2818 VSS 0.038015f
C19965 DVDD.n2819 VSS -0.729404f
C19966 DVDD.n2820 VSS 0.033044f
C19967 DVDD.n2821 VSS 0.026049f
C19968 DVDD.n2822 VSS 0.026049f
C19969 DVDD.n2823 VSS 0.018352f
C19970 DVDD.n2824 VSS 0.014419f
C19971 DVDD.n2825 VSS 0.026049f
C19972 DVDD.n2826 VSS 0.018614f
C19973 DVDD.n2827 VSS 0.026049f
C19974 DVDD.n2828 VSS 0.018614f
C19975 DVDD.n2829 VSS 0.026049f
C19976 DVDD.n2830 VSS 0.018614f
C19977 DVDD.n2831 VSS 0.026049f
C19978 DVDD.n2832 VSS 0.026049f
C19979 DVDD.n2833 VSS 0.014682f
C19980 DVDD.n2834 VSS 0.01809f
C19981 DVDD.n2835 VSS 0.026049f
C19982 DVDD.n2836 VSS 0.018614f
C19983 DVDD.n2837 VSS 0.052755f
C19984 DVDD.n2838 VSS 0.036673f
C19985 DVDD.n2839 VSS 0.017125f
C19986 DVDD.n2840 VSS 0.013654f
C19987 DVDD.n2841 VSS 0.031356f
C19988 DVDD.n2842 VSS 0.012783f
C19989 DVDD.n2844 VSS 0.029426f
C19990 DVDD.n2845 VSS 0.017125f
C19991 DVDD.n2846 VSS 0.016401f
C19992 DVDD.n2847 VSS 0.026049f
C19993 DVDD.n2848 VSS 0.013507f
C19994 DVDD.n2849 VSS 0.016643f
C19995 DVDD.n2850 VSS 0.026049f
C19996 DVDD.n2851 VSS 0.017125f
C19997 DVDD.n2852 VSS 0.026049f
C19998 DVDD.n2853 VSS 0.017125f
C19999 DVDD.n2854 VSS 0.026049f
C20000 DVDD.n2855 VSS 0.026049f
C20001 DVDD.n2856 VSS 0.014231f
C20002 DVDD.n2857 VSS 0.015919f
C20003 DVDD.n2858 VSS 0.026049f
C20004 DVDD.n2859 VSS 0.017125f
C20005 DVDD.n2860 VSS 0.026049f
C20006 DVDD.n2861 VSS 0.026049f
C20007 DVDD.n2862 VSS 0.017125f
C20008 DVDD.n2863 VSS 0.027459f
C20009 DVDD.n2864 VSS 0.06515f
C20010 DVDD.n2865 VSS 0.06515f
C20011 DVDD.n2866 VSS 0.130299f
C20012 DVDD.n2867 VSS 0.130299f
C20013 DVDD.n2868 VSS 0.130299f
C20014 DVDD.n2869 VSS 0.130299f
C20015 DVDD.n2870 VSS 0.130299f
C20016 DVDD.n2871 VSS 0.1225f
C20017 DVDD.n2872 VSS 0.130299f
C20018 DVDD.n2873 VSS 0.130299f
C20019 DVDD.n2874 VSS 0.130299f
C20020 DVDD.n2875 VSS 0.130299f
C20021 DVDD.n2876 VSS 0.130299f
C20022 DVDD.n2877 VSS 0.130299f
C20023 DVDD.n2878 VSS 0.130299f
C20024 DVDD.n2879 VSS 0.130299f
C20025 DVDD.n2880 VSS 0.130299f
C20026 DVDD.n2881 VSS 0.130299f
C20027 DVDD.n2882 VSS 0.130299f
C20028 DVDD.n2883 VSS 0.130299f
C20029 DVDD.n2884 VSS 0.130299f
C20030 DVDD.n2885 VSS 0.130299f
C20031 DVDD.n2886 VSS 0.130299f
C20032 DVDD.n2887 VSS 0.130299f
C20033 DVDD.n2888 VSS 0.130299f
C20034 DVDD.n2889 VSS 0.130299f
C20035 DVDD.n2890 VSS 0.130299f
C20036 DVDD.n2891 VSS 0.130299f
C20037 DVDD.n2892 VSS 0.130299f
C20038 DVDD.n2893 VSS 0.130299f
C20039 DVDD.n2894 VSS 0.130299f
C20040 DVDD.n2895 VSS 0.130299f
C20041 DVDD.n2896 VSS 0.130299f
C20042 DVDD.n2897 VSS 0.130299f
C20043 DVDD.n2898 VSS 0.130299f
C20044 DVDD.n2899 VSS 0.130299f
C20045 DVDD.n2900 VSS 0.130299f
C20046 DVDD.n2901 VSS 0.130299f
C20047 DVDD.n2902 VSS 0.130299f
C20048 DVDD.n2903 VSS 0.130299f
C20049 DVDD.n2904 VSS 0.130299f
C20050 DVDD.n2905 VSS 0.130299f
C20051 DVDD.n2906 VSS 0.130299f
C20052 DVDD.n2907 VSS 0.130299f
C20053 DVDD.n2908 VSS 0.130299f
C20054 DVDD.n2909 VSS 0.130299f
C20055 DVDD.n2910 VSS 0.130299f
C20056 DVDD.n2911 VSS 0.130299f
C20057 DVDD.n2912 VSS 0.130299f
C20058 DVDD.n2913 VSS 0.130299f
C20059 DVDD.n2914 VSS 0.130299f
C20060 DVDD.n2915 VSS 0.130299f
C20061 DVDD.n2916 VSS 0.130299f
C20062 DVDD.n2917 VSS 0.130299f
C20063 DVDD.n2918 VSS 0.130299f
C20064 DVDD.n2919 VSS 0.130299f
C20065 DVDD.n2920 VSS 0.130299f
C20066 DVDD.n2921 VSS 0.130299f
C20067 DVDD.n2922 VSS 0.130299f
C20068 DVDD.n2923 VSS 0.130299f
C20069 DVDD.n2924 VSS 0.130299f
C20070 DVDD.n2925 VSS 0.130299f
C20071 DVDD.n2926 VSS 0.130299f
C20072 DVDD.n2927 VSS 0.130299f
C20073 DVDD.n2928 VSS 0.130299f
C20074 DVDD.n2929 VSS 0.130299f
C20075 DVDD.n2930 VSS 0.130299f
C20076 DVDD.n2931 VSS 0.130299f
C20077 DVDD.n2932 VSS 0.130299f
C20078 DVDD.n2933 VSS 0.130299f
C20079 DVDD.n2934 VSS 0.130299f
C20080 DVDD.n2935 VSS 0.130299f
C20081 DVDD.n2936 VSS 0.130299f
C20082 DVDD.n2937 VSS 0.130299f
C20083 DVDD.n2938 VSS 0.130299f
C20084 DVDD.n2939 VSS 0.130299f
C20085 DVDD.n2940 VSS 0.130299f
C20086 DVDD.n2941 VSS 0.130299f
C20087 DVDD.n2942 VSS 0.130299f
C20088 DVDD.n2943 VSS 0.130299f
C20089 DVDD.n2944 VSS 0.06515f
C20090 DVDD.n2945 VSS 0.06515f
C20091 DVDD.n2946 VSS 0.014157f
C20092 DVDD.n2947 VSS 0.06515f
C20093 DVDD.n2948 VSS 0.071114f
C20094 DVDD.n2949 VSS 0.130299f
C20095 DVDD.n2950 VSS 0.130299f
C20096 DVDD.n2951 VSS 0.130299f
C20097 DVDD.n2952 VSS 0.130299f
C20098 DVDD.n2953 VSS 0.130299f
C20099 DVDD.n2954 VSS 0.130299f
C20100 DVDD.n2955 VSS 0.130299f
C20101 DVDD.n2956 VSS 0.130299f
C20102 DVDD.n2957 VSS 0.130299f
C20103 DVDD.n2958 VSS 0.130299f
C20104 DVDD.n2959 VSS 0.130299f
C20105 DVDD.n2960 VSS 0.130299f
C20106 DVDD.n2961 VSS 0.130299f
C20107 DVDD.n2962 VSS 0.130299f
C20108 DVDD.n2963 VSS 0.130299f
C20109 DVDD.n2964 VSS 0.130299f
C20110 DVDD.n2965 VSS 0.130299f
C20111 DVDD.n2966 VSS 0.130299f
C20112 DVDD.n2967 VSS 0.130299f
C20113 DVDD.n2968 VSS 0.130299f
C20114 DVDD.n2969 VSS 0.130299f
C20115 DVDD.n2970 VSS 0.130299f
C20116 DVDD.n2971 VSS 0.130299f
C20117 DVDD.n2972 VSS 0.130299f
C20118 DVDD.n2973 VSS 0.130299f
C20119 DVDD.n2974 VSS 0.130299f
C20120 DVDD.n2975 VSS 0.130299f
C20121 DVDD.n2976 VSS 0.130299f
C20122 DVDD.n2977 VSS 0.130299f
C20123 DVDD.n2978 VSS 0.117453f
C20124 DVDD.n2979 VSS 0.066985f
C20125 DVDD.n2980 VSS 0.171513f
C20126 DVDD.n2981 VSS 0.627997f
C20127 DVDD.n2982 VSS 0.117453f
C20128 DVDD.n2983 VSS 0.130299f
C20129 DVDD.n2984 VSS 0.130299f
C20130 DVDD.n2985 VSS 0.130299f
C20131 DVDD.n2986 VSS 0.130299f
C20132 DVDD.n2987 VSS 0.130299f
C20133 DVDD.n2988 VSS 0.130299f
C20134 DVDD.n2989 VSS 0.130299f
C20135 DVDD.n2990 VSS 0.130299f
C20136 DVDD.n2991 VSS 0.130299f
C20137 DVDD.n2992 VSS 0.130299f
C20138 DVDD.n2993 VSS 0.130299f
C20139 DVDD.n2994 VSS 0.130299f
C20140 DVDD.n2995 VSS 0.130299f
C20141 DVDD.n2996 VSS 0.130299f
C20142 DVDD.n2997 VSS 0.130299f
C20143 DVDD.n2998 VSS 0.130299f
C20144 DVDD.n2999 VSS 0.130299f
C20145 DVDD.n3000 VSS 0.130299f
C20146 DVDD.n3001 VSS 0.130299f
C20147 DVDD.n3002 VSS 0.130299f
C20148 DVDD.n3003 VSS 0.130299f
C20149 DVDD.n3004 VSS 0.130299f
C20150 DVDD.n3005 VSS 0.130299f
C20151 DVDD.n3006 VSS 0.130299f
C20152 DVDD.n3007 VSS 0.130299f
C20153 DVDD.n3008 VSS 0.130299f
C20154 DVDD.n3009 VSS 0.130299f
C20155 DVDD.n3010 VSS 0.130299f
C20156 DVDD.n3011 VSS 0.130299f
C20157 DVDD.n3012 VSS 0.130299f
C20158 DVDD.n3013 VSS 0.130299f
C20159 DVDD.n3014 VSS 0.130299f
C20160 DVDD.n3015 VSS 0.130299f
C20161 DVDD.n3016 VSS 0.130299f
C20162 DVDD.n3017 VSS 0.130299f
C20163 DVDD.n3018 VSS 0.130299f
C20164 DVDD.n3019 VSS 0.130299f
C20165 DVDD.n3020 VSS 0.130299f
C20166 DVDD.n3021 VSS 0.072949f
C20167 DVDD.n3022 VSS 0.091678f
C20168 DVDD.n3023 VSS 0.159245f
C20169 DVDD.n3024 VSS 0.074051f
C20170 DVDD.n3025 VSS 0.390389f
C20171 DVDD.n3026 VSS 4.34929f
C20172 DVDD.t40 VSS 1.35641f
C20173 DVDD.t131 VSS 3.94057f
C20174 DVDD.n3027 VSS 2.91939f
C20175 DVDD.n3028 VSS 0.154353f
C20176 DVDD.n3029 VSS 0.213342f
C20177 DVDD.n3030 VSS 0.279212f
C20178 DVDD.n3031 VSS 0.213342f
C20179 DVDD.n3032 VSS 0.448313f
C20180 DVDD.n3033 VSS 0.448313f
C20181 DVDD.n3034 VSS 0.139606f
C20182 DVDD.n3035 VSS 0.007073f
C20183 DVDD.n3036 VSS 0.139606f
C20184 DVDD.n3037 VSS 0.279212f
C20185 DVDD.n3038 VSS 0.448313f
C20186 DVDD.n3039 VSS 0.213342f
C20187 DVDD.n3040 VSS 0.139606f
C20188 DVDD.n3041 VSS 0.139606f
C20189 DVDD.n3042 VSS 0.007073f
C20190 DVDD.n3043 VSS 0.139606f
C20191 DVDD.n3044 VSS 0.139606f
C20192 DVDD.n3045 VSS 0.279212f
C20193 DVDD.n3046 VSS 0.279212f
C20194 DVDD.n3047 VSS 0.279212f
C20195 DVDD.n3048 VSS 0.448313f
C20196 DVDD.n3049 VSS 0.279212f
C20197 DVDD.n3050 VSS 0.279212f
C20198 DVDD.n3051 VSS 0.139606f
C20199 DVDD.n3052 VSS 0.139606f
C20200 DVDD.n3053 VSS 0.012307f
C20201 DVDD.n3054 VSS 0.308902f
C20202 DVDD.n3055 VSS 0.445363f
C20203 DVDD.n3056 VSS 0.279212f
C20204 DVDD.n3057 VSS 0.279212f
C20205 DVDD.n3058 VSS 0.279212f
C20206 DVDD.n3059 VSS 0.279212f
C20207 DVDD.n3060 VSS 0.279212f
C20208 DVDD.n3061 VSS 0.279212f
C20209 DVDD.n3062 VSS 0.264465f
C20210 DVDD.n3063 VSS 0.19367f
C20211 DVDD.n3064 VSS 0.105662f
C20212 DVDD.n3065 VSS 0.090342f
C20213 DVDD.n3066 VSS 0.003537f
C20214 DVDD.n3067 VSS 0.005305f
C20215 DVDD.n3068 VSS 0.007073f
C20216 DVDD.n3069 VSS 0.139606f
C20217 DVDD.n3070 VSS 0.139606f
C20218 DVDD.n3071 VSS 0.205477f
C20219 DVDD.n3072 VSS 0.279212f
C20220 DVDD.n3073 VSS 0.279212f
C20221 DVDD.n3074 VSS 0.279212f
C20222 DVDD.n3075 VSS 0.279212f
C20223 DVDD.n3076 VSS 0.279212f
C20224 DVDD.n3077 VSS 0.464043f
C20225 DVDD.n3078 VSS 0.464043f
C20226 DVDD.n3079 VSS 0.464043f
C20227 DVDD.n3080 VSS 0.279212f
C20228 DVDD.n3081 VSS 0.279212f
C20229 DVDD.n3082 VSS 0.279212f
C20230 DVDD.n3083 VSS 0.279212f
C20231 DVDD.n3084 VSS 0.205477f
C20232 DVDD.n3085 VSS 0.205477f
C20233 DVDD.n3086 VSS 0.076685f
C20234 DVDD.n3087 VSS 0.168643f
C20235 DVDD.n3088 VSS 0.168103f
C20236 DVDD.n3089 VSS 0.009831f
C20237 DVDD.n3090 VSS 1.15156f
C20238 DVDD.n3091 VSS 0.344417f
C20239 DVDD.n3092 VSS 0.34515f
C20240 DVDD.n3093 VSS 0.168103f
C20241 DVDD.n3094 VSS 0.168643f
C20242 DVDD.n3095 VSS 0.099297f
C20243 DVDD.n3096 VSS 0.073736f
C20244 DVDD.n3097 VSS 0.01324f
C20245 DVDD.n3098 VSS 0.073736f
C20246 DVDD.n3099 VSS 0.139689f
C20247 DVDD.n3100 VSS 0.205477f
C20248 DVDD.n3101 VSS 0.279212f
C20249 DVDD.n3102 VSS 0.279212f
C20250 DVDD.n3103 VSS 0.464043f
C20251 DVDD.n3104 VSS 0.279212f
C20252 DVDD.n3105 VSS 0.279212f
C20253 DVDD.n3106 VSS 0.464043f
C20254 DVDD.n3107 VSS 0.464043f
C20255 DVDD.n3108 VSS 0.279212f
C20256 DVDD.n3109 VSS 0.139606f
C20257 DVDD.n3111 VSS 0.013469f
C20258 DVDD.n3113 VSS 0.017125f
C20259 DVDD.n3114 VSS 0.139606f
C20260 DVDD.n3115 VSS 0.279212f
C20261 DVDD.n3116 VSS 0.279212f
C20262 DVDD.n3117 VSS 0.279212f
C20263 DVDD.n3118 VSS 0.205477f
C20264 DVDD.n3119 VSS 0.139606f
C20265 DVDD.n3120 VSS 0.013025f
C20266 DVDD.n3121 VSS 0.017125f
C20267 DVDD.n3122 VSS 0.013748f
C20268 DVDD.n3123 VSS 0.028702f
C20269 DVDD.n3124 VSS 0.015678f
C20270 DVDD.n3125 VSS 0.026049f
C20271 DVDD.n3126 VSS 0.013025f
C20272 DVDD.n3127 VSS 0.017125f
C20273 DVDD.n3128 VSS 0.139606f
C20274 DVDD.n3129 VSS 0.213342f
C20275 DVDD.n3130 VSS 0.279212f
C20276 DVDD.n3131 VSS 0.279212f
C20277 DVDD.n3132 VSS 0.279212f
C20278 DVDD.n3133 VSS 0.139606f
C20279 DVDD.n3134 VSS 0.013025f
C20280 DVDD.n3135 VSS 0.017125f
C20281 DVDD.n3136 VSS -0.22829f
C20282 DVDD.n3137 VSS -0.22829f
C20283 DVDD.n3138 VSS 0.013025f
C20284 DVDD.n3139 VSS 0.026049f
C20285 DVDD.n3140 VSS 0.017849f
C20286 DVDD.n3141 VSS 0.139606f
C20287 DVDD.n3142 VSS 0.139606f
C20288 DVDD.n3143 VSS 0.139606f
C20289 DVDD.n3144 VSS 0.448313f
C20290 DVDD.n3145 VSS 0.279212f
C20291 DVDD.n3146 VSS 0.448313f
C20292 DVDD.n3147 VSS 0.448313f
C20293 DVDD.n3148 VSS 0.279212f
C20294 DVDD.n3149 VSS 0.279212f
C20295 DVDD.n3150 VSS 0.013025f
C20296 DVDD.n3151 VSS 0.013025f
C20297 DVDD.n3152 VSS 0.013025f
C20298 DVDD.n3153 VSS 0.013025f
C20299 DVDD.n3154 VSS 0.013025f
C20300 DVDD.n3155 VSS 0.013025f
C20301 DVDD.n3156 VSS 0.013025f
C20302 DVDD.n3157 VSS 0.025227f
C20303 DVDD.n3158 VSS 0.021225f
C20304 DVDD.n3159 VSS 0.139606f
C20305 DVDD.n3160 VSS 0.028702f
C20306 DVDD.n3161 VSS 0.031247f
C20307 DVDD.n3162 VSS 0.013025f
C20308 DVDD.n3163 VSS 0.013025f
C20309 DVDD.n3164 VSS 0.013025f
C20310 DVDD.n3165 VSS 0.013025f
C20311 DVDD.n3166 VSS 0.013025f
C20312 DVDD.n3167 VSS 0.013025f
C20313 DVDD.n3168 VSS 0.015557f
C20314 DVDD.n3169 VSS 0.026049f
C20315 DVDD.n3170 VSS 0.016763f
C20316 DVDD.n3171 VSS 0.139606f
C20317 DVDD.n3172 VSS 0.139606f
C20318 DVDD.n3173 VSS 0.139606f
C20319 DVDD.n3174 VSS 0.013025f
C20320 DVDD.n3175 VSS 0.013025f
C20321 DVDD.n3176 VSS 0.013025f
C20322 DVDD.n3177 VSS 0.013025f
C20323 DVDD.n3178 VSS 0.013025f
C20324 DVDD.n3179 VSS 0.013025f
C20325 DVDD.n3180 VSS 0.013025f
C20326 DVDD.n3181 VSS 0.021225f
C20327 DVDD.n3182 VSS 0.025227f
C20328 DVDD.n3183 VSS 0.268398f
C20329 DVDD.n3184 VSS 0.028702f
C20330 DVDD.n3186 VSS 0.018693f
C20331 DVDD.n3187 VSS 0.013025f
C20332 DVDD.n3188 VSS 0.013025f
C20333 DVDD.n3189 VSS 0.013025f
C20334 DVDD.n3190 VSS 0.013025f
C20335 DVDD.n3191 VSS 0.013025f
C20336 DVDD.n3192 VSS 0.017125f
C20337 DVDD.n3193 VSS 0.026049f
C20338 DVDD.n3194 VSS 0.013025f
C20339 DVDD.n3195 VSS 0.026049f
C20340 DVDD.n3196 VSS 0.017125f
C20341 DVDD.n3197 VSS 0.139606f
C20342 DVDD.n3198 VSS 0.308707f
C20343 DVDD.n3199 VSS 0.279212f
C20344 DVDD.n3200 VSS 0.314606f
C20345 DVDD.n3201 VSS 0.448313f
C20346 DVDD.n3202 VSS 0.279212f
C20347 DVDD.n3203 VSS 0.213342f
C20348 DVDD.n3204 VSS 0.279212f
C20349 DVDD.n3205 VSS 0.139606f
C20350 DVDD.n3206 VSS 0.017125f
C20351 DVDD.n3207 VSS 0.026049f
C20352 DVDD.n3208 VSS 0.016401f
C20353 DVDD.n3209 VSS 0.028702f
C20354 DVDD.n3210 VSS 0.013025f
C20355 DVDD.n3211 VSS 0.139606f
C20356 DVDD.n3212 VSS 0.279212f
C20357 DVDD.n3213 VSS 0.464043f
C20358 DVDD.n3214 VSS 0.464043f
C20359 DVDD.n3215 VSS 0.279212f
C20360 DVDD.n3216 VSS 0.279212f
C20361 DVDD.n3217 VSS 0.279212f
C20362 DVDD.n3218 VSS 0.205477f
C20363 DVDD.n3219 VSS 0.205477f
C20364 DVDD.n3220 VSS 0.279212f
C20365 DVDD.n3221 VSS 0.029378f
C20366 DVDD.n3222 VSS 0.05005f
C20367 DVDD.n3223 VSS 0.010331f
C20368 DVDD.n3224 VSS 0.012222f
C20369 DVDD.n3225 VSS 0.012368f
C20370 DVDD.n3226 VSS 0.037686f
C20371 DVDD.n3227 VSS 0.04151f
C20372 DVDD.n3228 VSS 0.018614f
C20373 DVDD.n3229 VSS 0.139606f
C20374 DVDD.n3230 VSS 0.139606f
C20375 DVDD.n3231 VSS 0.03844f
C20376 DVDD.n3232 VSS 0.04151f
C20377 DVDD.n3233 VSS 0.009167f
C20378 DVDD.n3234 VSS 0.007857f
C20379 DVDD.n3235 VSS 0.008003f
C20380 DVDD.n3236 VSS 0.023055f
C20381 DVDD.n3237 VSS 0.41539f
C20382 DVDD.n3238 VSS 0.109896f
C20383 DVDD.n3239 VSS 0.004874f
C20384 DVDD.n3240 VSS 0.080044f
C20385 DVDD.n3241 VSS 0.022477f
C20386 DVDD.n3242 VSS 0.038044f
C20387 DVDD.n3243 VSS 0.007857f
C20388 DVDD.n3244 VSS 0.156613f
C20389 DVDD.n3245 VSS 0.208862f
C20390 DVDD.n3246 VSS 0.04151f
C20391 DVDD.n3247 VSS 0.266194f
C20392 DVDD.n3248 VSS 0.139606f
C20393 DVDD.n3249 VSS 0.270437f
C20394 DVDD.n3250 VSS 0.279212f
C20395 DVDD.n3251 VSS 0.279212f
C20396 DVDD.n3252 VSS 0.213342f
C20397 DVDD.n3253 VSS 0.213342f
C20398 DVDD.n3254 VSS 0.279212f
C20399 DVDD.n3255 VSS 0.793212f
C20400 DVDD.n3256 VSS 0.279212f
C20401 DVDD.n3257 VSS 0.139606f
C20402 DVDD.n3258 VSS 0.010331f
C20403 DVDD.n3259 VSS 0.009021f
C20404 DVDD.n3260 VSS 0.04151f
C20405 DVDD.n3261 VSS 0.139606f
C20406 DVDD.n3262 VSS 0.007857f
C20407 DVDD.n3263 VSS 0.012513f
C20408 DVDD.n3264 VSS 0.015715f
C20409 DVDD.n3265 VSS 0.010331f
C20410 DVDD.n3266 VSS 0.007857f
C20411 DVDD.n3267 VSS 0.139606f
C20412 DVDD.n3268 VSS 0.04151f
C20413 DVDD.n3269 VSS 0.035706f
C20414 DVDD.n3270 VSS 0.018614f
C20415 DVDD.n3271 VSS 0.270437f
C20416 DVDD.n3272 VSS 0.04151f
C20417 DVDD.n3273 VSS 0.266194f
C20418 DVDD.n3274 VSS 0.139606f
C20419 DVDD.n3275 VSS 0.04531f
C20420 DVDD.n3276 VSS 0.011495f
C20421 DVDD.n3277 VSS 0.007857f
C20422 DVDD.n3278 VSS 0.038044f
C20423 DVDD.n3279 VSS 0.008003f
C20424 DVDD.n3280 VSS 0.009021f
C20425 DVDD.n3281 VSS 0.139606f
C20426 DVDD.n3282 VSS 0.018614f
C20427 DVDD.n3283 VSS 0.018614f
C20428 DVDD.n3284 VSS 0.037228f
C20429 DVDD.n3285 VSS 0.037228f
C20430 DVDD.n3286 VSS 0.105598f
C20431 DVDD.n3287 VSS 0.037228f
C20432 DVDD.n3288 VSS 0.028446f
C20433 DVDD.n3289 VSS 0.018614f
C20434 DVDD.n3290 VSS 0.028446f
C20435 DVDD.n3291 VSS 0.037228f
C20436 DVDD.n3292 VSS 0.018614f
C20437 DVDD.n3293 VSS 0.018614f
C20438 DVDD.n3294 VSS 0.04151f
C20439 DVDD.n3295 VSS 0.139606f
C20440 DVDD.n3296 VSS 0.139606f
C20441 DVDD.n3297 VSS 0.04151f
C20442 DVDD.n3298 VSS 0.03844f
C20443 DVDD.n3299 VSS 0.04151f
C20444 DVDD.n3300 VSS 0.279212f
C20445 DVDD.n3301 VSS 0.279212f
C20446 DVDD.n3302 VSS 0.279212f
C20447 DVDD.n3303 VSS 0.793212f
C20448 DVDD.n3304 VSS 0.279212f
C20449 DVDD.n3305 VSS 0.213342f
C20450 DVDD.n3306 VSS 0.213342f
C20451 DVDD.n3307 VSS 0.139606f
C20452 DVDD.n3308 VSS 0.009167f
C20453 DVDD.n3309 VSS 0.007857f
C20454 DVDD.n3310 VSS 0.037283f
C20455 DVDD.n3311 VSS 0.004971f
C20456 DVDD.n3312 VSS 0.022477f
C20457 DVDD.n3313 VSS 0.020537f
C20458 DVDD.n3314 VSS 0.082786f
C20459 DVDD.n3315 VSS 0.109897f
C20460 DVDD.n3316 VSS 0.040036f
C20461 DVDD.n3317 VSS 0.127381f
C20462 DVDD.n3318 VSS 0.24914f
C20463 DVDD.n3319 VSS 0.414431f
C20464 DVDD.n3320 VSS 0.129553f
C20465 DVDD.n3321 VSS 0.037686f
C20466 DVDD.n3322 VSS 0.129553f
C20467 DVDD.n3323 VSS 0.560908f
C20468 DVDD.n3324 VSS 0.063828f
C20469 DVDD.n3325 VSS 0.156613f
C20470 DVDD.n3326 VSS 0.125562f
C20471 DVDD.n3327 VSS 0.243607f
C20472 DVDD.n3328 VSS 0.270437f
C20473 DVDD.n3329 VSS 0.208862f
C20474 DVDD.n3330 VSS 0.127381f
C20475 DVDD.n3331 VSS 0.249148f
C20476 DVDD.n3332 VSS 0.010193f
C20477 DVDD.n3333 VSS 0.004844f
C20478 DVDD.n3334 VSS 0.070963f
C20479 DVDD.n3335 VSS 0.013368f
C20480 DVDD.n3336 VSS 0.023055f
C20481 DVDD.n3337 VSS 0.247868f
C20482 DVDD.n3338 VSS 0.007857f
C20483 DVDD.n3339 VSS 0.015569f
C20484 DVDD.n3340 VSS 0.03844f
C20485 DVDD.n3341 VSS 0.051457f
C20486 DVDD.n3342 VSS 0.147497f
C20487 DVDD.n3343 VSS 0.152164f
C20488 DVDD.n3344 VSS 0.029378f
C20489 DVDD.n3345 VSS 0.020755f
C20490 DVDD.n3346 VSS 0.092468f
C20491 DVDD.n3347 VSS 0.05005f
C20492 DVDD.n3348 VSS 0.143832f
C20493 DVDD.n3349 VSS 0.074135f
C20494 DVDD.n3350 VSS 0.010331f
C20495 DVDD.n3351 VSS 0.007857f
C20496 DVDD.n3352 VSS 0.011495f
C20497 DVDD.n3353 VSS 0.012222f
C20498 DVDD.n3354 VSS 0.012368f
C20499 DVDD.n3355 VSS 0.012368f
C20500 DVDD.n3356 VSS 0.010331f
C20501 DVDD.n3357 VSS 0.007857f
C20502 DVDD.n3358 VSS 0.139606f
C20503 DVDD.n3359 VSS 0.04151f
C20504 DVDD.n3360 VSS 0.04151f
C20505 DVDD.n3361 VSS 0.139606f
C20506 DVDD.n3362 VSS 0.007857f
C20507 DVDD.n3363 VSS 0.010331f
C20508 DVDD.n3364 VSS 0.015715f
C20509 DVDD.n3365 VSS 0.012513f
C20510 DVDD.n3366 VSS 0.010331f
C20511 DVDD.n3367 VSS 0.007857f
C20512 DVDD.n3368 VSS 0.287499f
C20513 DVDD.n3369 VSS 0.04531f
C20514 DVDD.n3370 VSS 0.038284f
C20515 DVDD.n3371 VSS 0.04531f
C20516 DVDD.n3372 VSS 0.287499f
C20517 DVDD.n3373 VSS 0.04531f
C20518 DVDD.n3374 VSS 0.270437f
C20519 DVDD.n3375 VSS 0.243607f
C20520 DVDD.n3376 VSS 0.125562f
C20521 DVDD.n3377 VSS 0.011495f
C20522 DVDD.n3378 VSS 0.020537f
C20523 DVDD.n3379 VSS 0.013397f
C20524 DVDD.n3380 VSS 0.071025f
C20525 DVDD.n3381 VSS 0.005003f
C20526 DVDD.n3382 VSS 0.010158f
C20527 DVDD.n3383 VSS 0.247859f
C20528 DVDD.n3384 VSS 0.007857f
C20529 DVDD.n3385 VSS 0.015569f
C20530 DVDD.n3386 VSS 0.012368f
C20531 DVDD.n3387 VSS 0.010331f
C20532 DVDD.n3388 VSS 0.007857f
C20533 DVDD.n3389 VSS 0.139606f
C20534 DVDD.n3390 VSS 0.04151f
C20535 DVDD.n3391 VSS 0.03844f
C20536 DVDD.n3392 VSS 0.020755f
C20537 DVDD.n3393 VSS 0.092468f
C20538 DVDD.n3394 VSS 0.143832f
C20539 DVDD.n3395 VSS 0.074135f
C20540 DVDD.n3396 VSS 0.011495f
C20541 DVDD.n3397 VSS 0.007857f
C20542 DVDD.n3398 VSS 0.139689f
C20543 DVDD.n3399 VSS 0.245786f
C20544 DVDD.n3400 VSS 0.279212f
C20545 DVDD.n3401 VSS 0.279212f
C20546 DVDD.n3402 VSS 0.279212f
C20547 DVDD.n3403 VSS 0.279212f
C20548 DVDD.n3404 VSS 0.464043f
C20549 DVDD.n3405 VSS 0.464043f
C20550 DVDD.n3406 VSS 0.464043f
C20551 DVDD.n3407 VSS 0.329353f
C20552 DVDD.n3408 VSS 0.139654f
C20553 DVDD.n3409 VSS 0.139606f
C20554 DVDD.n3410 VSS 0.139606f
C20555 DVDD.n3411 VSS 0.014472f
C20556 DVDD.n3414 VSS 0.013469f
C20557 DVDD.n3415 VSS 0.028896f
C20558 DVDD.n3416 VSS 0.031356f
C20559 DVDD.n3417 VSS 0.017125f
C20560 DVDD.n3418 VSS 0.013025f
C20561 DVDD.n3419 VSS 0.139606f
C20562 DVDD.n3420 VSS 0.139606f
C20563 DVDD.n3421 VSS 0.279212f
C20564 DVDD.n3422 VSS 0.279212f
C20565 DVDD.n3423 VSS 0.279212f
C20566 DVDD.n3424 VSS 0.279212f
C20567 DVDD.n3425 VSS 0.279212f
C20568 DVDD.n3426 VSS 0.205477f
C20569 DVDD.n3427 VSS 0.139606f
C20570 DVDD.n3428 VSS 0.139606f
C20571 DVDD.n3429 VSS 0.013025f
C20572 DVDD.n3430 VSS 0.017125f
C20573 DVDD.n3431 VSS 0.015678f
C20574 DVDD.n3432 VSS 0.026049f
C20575 DVDD.n3433 VSS 0.026049f
C20576 DVDD.n3434 VSS 0.013748f
C20577 DVDD.n3435 VSS 0.013025f
C20578 DVDD.n3436 VSS 0.017125f
C20579 DVDD.n3437 VSS 0.139606f
C20580 DVDD.n3438 VSS 0.139606f
C20581 DVDD.n3439 VSS 0.013025f
C20582 DVDD.n3440 VSS 0.013025f
C20583 DVDD.n3441 VSS 0.017125f
C20584 DVDD.n3442 VSS 0.026049f
C20585 DVDD.n3443 VSS -0.22829f
C20586 DVDD.n3444 VSS -0.22829f
C20587 DVDD.n3445 VSS 0.026049f
C20588 DVDD.n3446 VSS 0.139606f
C20589 DVDD.n3447 VSS 0.139606f
C20590 DVDD.n3448 VSS 0.279212f
C20591 DVDD.n3449 VSS 0.279212f
C20592 DVDD.n3450 VSS 0.279212f
C20593 DVDD.n3451 VSS 0.279212f
C20594 DVDD.n3452 VSS 0.139606f
C20595 DVDD.n3453 VSS 0.213342f
C20596 DVDD.n3454 VSS 0.213342f
C20597 DVDD.n3455 VSS 0.279212f
C20598 DVDD.n3456 VSS 0.279212f
C20599 DVDD.n3457 VSS 0.279212f
C20600 DVDD.n3458 VSS 0.279212f
C20601 DVDD.n3459 VSS 0.279212f
C20602 DVDD.n3460 VSS 0.448313f
C20603 DVDD.n3461 VSS 0.448313f
C20604 DVDD.n3462 VSS 0.448313f
C20605 DVDD.n3463 VSS 0.139606f
C20606 DVDD.n3464 VSS 0.139606f
C20607 DVDD.n3465 VSS 0.013025f
C20608 DVDD.n3466 VSS 0.017125f
C20609 DVDD.n3467 VSS 0.026049f
C20610 DVDD.n3468 VSS 0.026049f
C20611 DVDD.n3469 VSS 0.017849f
C20612 DVDD.n3470 VSS 0.026049f
C20613 DVDD.n3471 VSS 0.015678f
C20614 DVDD.n3472 VSS 0.015678f
C20615 DVDD.n3473 VSS 0.006671f
C20616 DVDD.n3474 VSS 0.059516f
C20617 DVDD.n3475 VSS 0.017125f
C20618 DVDD.n3476 VSS 0.035818f
C20619 DVDD.n3477 VSS 0.035818f
C20620 DVDD.n3478 VSS 0.014593f
C20621 DVDD.n3479 VSS 0.015557f
C20622 DVDD.n3480 VSS 0.026049f
C20623 DVDD.n3481 VSS 0.017125f
C20624 DVDD.n3482 VSS 0.026049f
C20625 DVDD.n3483 VSS 0.017125f
C20626 DVDD.n3484 VSS 0.026049f
C20627 DVDD.n3485 VSS 0.026049f
C20628 DVDD.n3486 VSS 0.015316f
C20629 DVDD.n3487 VSS 0.014834f
C20630 DVDD.n3488 VSS 0.026049f
C20631 DVDD.n3489 VSS 0.017125f
C20632 DVDD.n3490 VSS 0.026049f
C20633 DVDD.n3491 VSS 0.017125f
C20634 DVDD.n3492 VSS 0.026049f
C20635 DVDD.n3493 VSS 0.026049f
C20636 DVDD.n3494 VSS 0.01604f
C20637 DVDD.n3495 VSS 0.01411f
C20638 DVDD.n3496 VSS 0.026049f
C20639 DVDD.n3497 VSS 0.017125f
C20640 DVDD.n3498 VSS 0.026049f
C20641 DVDD.n3499 VSS 0.017125f
C20642 DVDD.n3500 VSS 0.026049f
C20643 DVDD.n3501 VSS 0.026049f
C20644 DVDD.n3502 VSS 0.016763f
C20645 DVDD.n3503 VSS 0.013387f
C20646 DVDD.n3504 VSS 0.026049f
C20647 DVDD.n3505 VSS 0.017125f
C20648 DVDD.n3506 VSS 0.026049f
C20649 DVDD.n3507 VSS 0.026049f
C20650 DVDD.n3508 VSS 0.013387f
C20651 DVDD.n3509 VSS 0.026049f
C20652 DVDD.n3510 VSS 0.026049f
C20653 DVDD.n3511 VSS 0.017125f
C20654 DVDD.n3512 VSS 0.013025f
C20655 DVDD.n3513 VSS 0.139606f
C20656 DVDD.n3514 VSS 0.031247f
C20657 DVDD.n3515 VSS -0.526826f
C20658 DVDD.n3516 VSS -0.526826f
C20659 DVDD.n3517 VSS 0.026049f
C20660 DVDD.n3518 VSS 0.016763f
C20661 DVDD.n3519 VSS 0.013387f
C20662 DVDD.n3520 VSS 0.026049f
C20663 DVDD.n3521 VSS 0.017125f
C20664 DVDD.n3522 VSS 0.026049f
C20665 DVDD.n3523 VSS 0.017125f
C20666 DVDD.n3524 VSS 0.026049f
C20667 DVDD.n3525 VSS 0.017125f
C20668 DVDD.n3526 VSS 0.026049f
C20669 DVDD.n3527 VSS 0.026049f
C20670 DVDD.n3528 VSS 0.013387f
C20671 DVDD.n3529 VSS 0.016763f
C20672 DVDD.n3530 VSS 0.026049f
C20673 DVDD.n3531 VSS 0.017125f
C20674 DVDD.n3532 VSS 0.026049f
C20675 DVDD.n3533 VSS 0.017125f
C20676 DVDD.n3534 VSS 0.026049f
C20677 DVDD.n3535 VSS 0.026049f
C20678 DVDD.n3536 VSS 0.01411f
C20679 DVDD.n3537 VSS 0.01604f
C20680 DVDD.n3538 VSS 0.026049f
C20681 DVDD.n3539 VSS 0.017125f
C20682 DVDD.n3540 VSS 0.026049f
C20683 DVDD.n3541 VSS 0.017125f
C20684 DVDD.n3542 VSS 0.026049f
C20685 DVDD.n3543 VSS 0.026049f
C20686 DVDD.n3544 VSS 0.014834f
C20687 DVDD.n3545 VSS 0.015316f
C20688 DVDD.n3546 VSS 0.026049f
C20689 DVDD.n3547 VSS 0.017125f
C20690 DVDD.n3548 VSS 0.026049f
C20691 DVDD.n3549 VSS 0.017125f
C20692 DVDD.n3550 VSS 0.026049f
C20693 DVDD.n3551 VSS 0.025808f
C20694 DVDD.n3552 VSS 0.026049f
C20695 DVDD.n3553 VSS 0.026049f
C20696 DVDD.n3554 VSS 0.015678f
C20697 DVDD.n3555 VSS 0.015678f
C20698 DVDD.n3556 VSS 0.006671f
C20699 DVDD.n3557 VSS 0.059516f
C20700 DVDD.n3558 VSS 0.017125f
C20701 DVDD.n3559 VSS 0.035818f
C20702 DVDD.n3560 VSS 0.023034f
C20703 DVDD.n3561 VSS 0.014593f
C20704 DVDD.n3562 VSS 0.213342f
C20705 DVDD.n3563 VSS 0.279212f
C20706 DVDD.n3564 VSS 0.279212f
C20707 DVDD.n3565 VSS 0.213342f
C20708 DVDD.n3566 VSS 0.279212f
C20709 DVDD.n3567 VSS 0.268398f
C20710 DVDD.n3568 VSS 0.139606f
C20711 DVDD.n3570 VSS 0.018693f
C20712 DVDD.n3571 VSS 0.139606f
C20713 DVDD.n3572 VSS 0.139606f
C20714 DVDD.n3573 VSS 0.279212f
C20715 DVDD.n3574 VSS 0.448313f
C20716 DVDD.n3575 VSS 0.314606f
C20717 DVDD.n3576 VSS 0.308707f
C20718 DVDD.n3577 VSS 0.013025f
C20719 DVDD.n3578 VSS 0.017125f
C20720 DVDD.n3579 VSS 0.026049f
C20721 DVDD.n3580 VSS 0.026049f
C20722 DVDD.n3581 VSS 0.017125f
C20723 DVDD.n3582 VSS 0.026049f
C20724 DVDD.n3583 VSS 0.139606f
C20725 DVDD.n3584 VSS 0.139606f
C20726 DVDD.n3585 VSS 0.279212f
C20727 DVDD.n3586 VSS 0.279212f
C20728 DVDD.n3587 VSS 0.139606f
C20729 DVDD.n3588 VSS 0.139606f
C20730 DVDD.n3589 VSS 0.013025f
C20731 DVDD.n3590 VSS 0.017125f
C20732 DVDD.n3591 VSS 0.026049f
C20733 DVDD.n3592 VSS 0.026049f
C20734 DVDD.n3593 VSS 0.026049f
C20735 DVDD.n3594 VSS 0.016401f
C20736 DVDD.n3595 VSS 0.013025f
C20737 DVDD.n3596 VSS 0.139606f
C20738 DVDD.n3597 VSS 0.139606f
C20739 DVDD.n3598 VSS 0.279212f
C20740 DVDD.n3599 VSS 0.279212f
C20741 DVDD.n3600 VSS 0.139606f
C20742 DVDD.n3601 VSS 0.139606f
C20743 DVDD.n3602 VSS 0.013025f
C20744 DVDD.n3603 VSS 0.014472f
C20745 DVDD.n3604 VSS 0.031356f
C20746 DVDD.n3605 VSS 0.028896f
C20747 DVDD.n3606 VSS 0.139654f
C20748 DVDD.n3607 VSS 0.329353f
C20749 DVDD.n3608 VSS 0.464043f
C20750 DVDD.n3609 VSS 0.464043f
C20751 DVDD.n3610 VSS 0.279212f
C20752 DVDD.n3611 VSS 0.279212f
C20753 DVDD.n3612 VSS 0.279212f
C20754 DVDD.n3613 VSS 0.245786f
C20755 DVDD.n3614 VSS 0.279212f
C20756 DVDD.n3615 VSS 0.205477f
C20757 DVDD.n3616 VSS 0.099297f
C20758 DVDD.n3617 VSS 3.46356f
C20759 DVDD.n3618 VSS 0.205477f
C20760 DVDD.n3619 VSS 0.205477f
C20761 DVDD.n3620 VSS 0.205477f
C20762 DVDD.n3621 VSS 0.279212f
C20763 DVDD.n3622 VSS 0.279212f
C20764 DVDD.n3623 VSS 0.279212f
C20765 DVDD.n3624 VSS 0.279212f
C20766 DVDD.n3625 VSS 0.279212f
C20767 DVDD.n3626 VSS 0.110112f
C20768 DVDD.n3627 VSS 0.062266f
C20769 DVDD.n3628 VSS 0.324924f
C20770 DVDD.n3629 VSS 0.459127f
C20771 DVDD.n3630 VSS 0.464043f
C20772 DVDD.n3631 VSS 0.464043f
C20773 DVDD.n3632 VSS 0.464043f
C20774 DVDD.n3633 VSS 0.279212f
C20775 DVDD.n3634 VSS 0.279212f
C20776 DVDD.n3635 VSS 0.279212f
C20777 DVDD.n3636 VSS 0.110112f
C20778 DVDD.n3637 VSS 0.110112f
C20779 DVDD.n3638 VSS 0.139606f
C20780 DVDD.n3639 VSS 0.031209f
C20781 DVDD.n3640 VSS 0.037585f
C20782 DVDD.n3641 VSS 0.037585f
C20783 DVDD.n3642 VSS 0.126825f
C20784 DVDD.n3643 VSS 0.110112f
C20785 DVDD.n3644 VSS 0.279212f
C20786 DVDD.n3645 VSS 0.205477f
C20787 DVDD.n3646 VSS 0.205477f
C20788 DVDD.n3647 VSS 2.78569f
C20789 DVDD.n3648 VSS 0.293381f
C20790 DVDD.n3649 VSS 0.040226f
C20791 DVDD.n3650 VSS 0.040226f
C20792 DVDD.n3651 VSS 0.040226f
C20793 DVDD.n3652 VSS 2.63401f
C20794 DVDD.n3653 VSS 0.110112f
C20795 DVDD.n3654 VSS 0.073736f
C20796 DVDD.n3655 VSS 0.037585f
C20797 DVDD.n3656 VSS 0.037585f
C20798 DVDD.n3657 VSS 0.009001f
C20799 DVDD.n3658 VSS 0.069733f
C20800 DVDD.t209 VSS 0.155477f
C20801 DVDD.n3659 VSS 0.1204f
C20802 DVDD.n3660 VSS 0.009001f
C20803 DVDD.n3661 VSS 0.069733f
C20804 DVDD.t212 VSS 0.155477f
C20805 DVDD.n3662 VSS 0.1204f
C20806 DVDD.n3663 VSS 0.041664f
C20807 DVDD.n3664 VSS 0.11896f
C20808 DVDD.n3665 VSS 0.03037f
C20809 DVDD.n3666 VSS 0.037585f
C20810 DVDD.n3667 VSS 0.139606f
C20811 DVDD.n3668 VSS 0.110112f
C20812 DVDD.n3669 VSS 0.279212f
C20813 DVDD.n3670 VSS 0.279212f
C20814 DVDD.n3671 VSS 0.279212f
C20815 DVDD.n3672 VSS 0.279212f
C20816 DVDD.n3673 VSS 0.279212f
C20817 DVDD.n3674 VSS 0.160252f
C20818 DVDD.n3675 VSS 0.448313f
C20819 DVDD.n3676 VSS 0.448313f
C20820 DVDD.n3677 VSS 0.448313f
C20821 DVDD.n3678 VSS 0.448313f
C20822 DVDD.n3679 VSS 0.279212f
C20823 DVDD.n3680 VSS 0.279212f
C20824 DVDD.n3681 VSS 0.279212f
C20825 DVDD.n3682 VSS 0.279212f
C20826 DVDD.n3683 VSS 0.279212f
C20827 DVDD.n3684 VSS 0.213342f
C20828 DVDD.n3685 VSS 0.213342f
C20829 DVDD.n3686 VSS 0.213342f
C20830 DVDD.n3687 VSS 1.06162f
C20831 DVDD.n3688 VSS 0.279212f
C20832 DVDD.t39 VSS 0.010225f
C20833 DVDD.t121 VSS 0.010225f
C20834 DVDD.n3689 VSS 0.039995f
C20835 DVDD.n3690 VSS 0.047512f
C20836 DVDD.t177 VSS 0.042669f
C20837 DVDD.n3691 VSS 0.372837f
C20838 DVDD.t176 VSS 0.335595f
C20839 DVDD.t38 VSS 0.202551f
C20840 DVDD.t123 VSS 0.042669f
C20841 DVDD.n3692 VSS 0.379366f
C20842 DVDD.t122 VSS 0.333372f
C20843 DVDD.t120 VSS 0.204777f
C20844 DVDD.n3693 VSS 0.099852f
C20845 DVDD.n3694 VSS -0.034921f
C20846 DVDD.n3695 VSS 0.030556f
C20847 DVDD.n3696 VSS 0.650969f
C20848 DVDD.n3697 VSS 0.509735f
C20849 DVDD.n3698 VSS 0.361156f
C20850 DVDD.n3699 VSS 0.199578f
C20851 DVDD.n3700 VSS 0.279212f
C20852 DVDD.n3701 VSS 0.205477f
C20853 DVDD.n3702 VSS 0.205477f
C20854 DVDD.n3703 VSS 0.205477f
C20855 DVDD.n3704 VSS 1.89279f
C20856 DVDD.n3705 VSS 0.059108f
C20857 DVDD.n3706 VSS 0.059108f
C20858 DVDD.n3707 VSS 0.022059f
C20859 DVDD.n3708 VSS 0.040159f
C20860 DVDD.n3709 VSS 0.040159f
C20861 DVDD.n3710 VSS 0.037228f
C20862 DVDD.n3711 VSS 0.037228f
C20863 DVDD.n3712 VSS 0.037228f
C20864 DVDD.n3713 VSS 0.040159f
C20865 DVDD.n3714 VSS 0.040159f
C20866 DVDD.n3715 VSS 0.08032f
C20867 DVDD.n3716 VSS 0.233369f
C20868 DVDD.n3717 VSS 0.080449f
C20869 DVDD.n3718 VSS 0.074464f
C20870 DVDD.n3719 VSS 0.901371f
C20871 DVDD.n3721 VSS 0.532172f
C20872 DVDD.n3722 VSS 0.037228f
C20873 DVDD.n3723 VSS 0.037228f
C20874 DVDD.n3724 VSS 0.037228f
C20875 DVDD.n3725 VSS 0.037228f
C20876 DVDD.n3726 VSS 0.037228f
C20877 DVDD.n3727 VSS 0.037228f
C20878 DVDD.n3728 VSS 0.037228f
C20879 DVDD.n3729 VSS 0.037228f
C20880 DVDD.n3730 VSS 0.037228f
C20881 DVDD.n3731 VSS 1.0352f
C20882 DVDD.n3732 VSS 0.279212f
C20883 DVDD.n3733 VSS 0.279212f
C20884 DVDD.n3734 VSS 0.139606f
C20885 DVDD.n3735 VSS 0.037228f
C20886 DVDD.n3736 VSS 0.037228f
C20887 DVDD.n3737 VSS 0.037228f
C20888 DVDD.n3738 VSS 0.037228f
C20889 DVDD.n3739 VSS 0.037228f
C20890 DVDD.n3740 VSS 0.037228f
C20891 DVDD.n3741 VSS 0.037228f
C20892 DVDD.n3742 VSS 0.037228f
C20893 DVDD.n3752 VSS 0.139606f
C20894 DVDD.n3753 VSS 0.037228f
C20895 DVDD.n3754 VSS 0.04016f
C20896 DVDD.n3755 VSS 0.08032f
C20897 DVDD.n3756 VSS 0.08032f
C20898 DVDD.n3757 VSS 0.08032f
C20899 DVDD.n3758 VSS 0.04016f
C20900 DVDD.n3759 VSS 0.04016f
C20901 DVDD.n3760 VSS 0.04016f
C20902 DVDD.n3761 VSS 0.037228f
C20903 DVDD.n3762 VSS 0.059108f
C20904 DVDD.n3763 VSS 0.02008f
C20905 DVDD.n3764 VSS 0.04016f
C20906 DVDD.n3765 VSS 0.037228f
C20907 DVDD.n3766 VSS 0.037228f
C20908 DVDD.n3767 VSS 0.04016f
C20909 DVDD.n3768 VSS 0.04016f
C20910 DVDD.n3769 VSS 0.08032f
C20911 DVDD.n3770 VSS 0.233369f
C20912 DVDD.n3771 VSS 0.080449f
C20913 DVDD.n3772 VSS 0.07646f
C20914 DVDD.n3773 VSS 0.063324f
C20915 DVDD.n3774 VSS 0.063314f
C20916 DVDD.n3775 VSS 0.624053f
C20917 DVDD.n3776 VSS 0.901345f
C20918 DVDD.n3777 VSS 0.139606f
C20919 DVDD.n3778 VSS 0.15632f
C20920 DVDD.n3779 VSS 0.217274f
C20921 DVDD.n3780 VSS 0.279212f
C20922 DVDD.n3781 VSS 0.279212f
C20923 DVDD.n3782 VSS 0.279212f
C20924 DVDD.n3783 VSS 0.279212f
C20925 DVDD.n3784 VSS 0.279212f
C20926 DVDD.n3785 VSS 0.279212f
C20927 DVDD.n3786 VSS 0.201544f
C20928 DVDD.n3787 VSS 0.279212f
C20929 DVDD.n3788 VSS 0.279212f
C20930 DVDD.n3789 VSS 0.279212f
C20931 DVDD.n3790 VSS 0.279212f
C20932 DVDD.n3791 VSS 0.279212f
C20933 DVDD.n3792 VSS 0.279212f
C20934 DVDD.n3793 VSS 0.279212f
C20935 DVDD.n3794 VSS 0.279212f
C20936 DVDD.n3795 VSS 0.279212f
C20937 DVDD.n3796 VSS 0.279212f
C20938 DVDD.n3797 VSS 0.279212f
C20939 DVDD.n3798 VSS 0.279212f
C20940 DVDD.n3799 VSS 0.279212f
C20941 DVDD.n3800 VSS 0.279212f
C20942 DVDD.n3801 VSS 0.279212f
C20943 DVDD.n3802 VSS 0.279212f
C20944 DVDD.n3803 VSS 0.186797f
C20945 DVDD.n3804 VSS 0.186797f
C20946 DVDD.n3805 VSS 0.099953f
C20947 DVDD.n3806 VSS 0.073932f
C20948 DVDD.n3807 VSS 0.123745f
C20949 DVDD.n3808 VSS 0.148913f
C20950 DVDD.n3809 VSS 0.148913f
C20951 DVDD.n3810 VSS 0.074457f
C20952 DVDD.n3811 VSS 0.074457f
C20953 DVDD.n3812 VSS 0.074457f
C20954 DVDD.n3813 VSS 0.007073f
C20955 DVDD.n3814 VSS 0.007073f
C20956 DVDD.n3815 VSS 0.012307f
C20957 DVDD.n3816 VSS 0.074457f
C20958 DVDD.n3817 VSS 0.074457f
C20959 DVDD.n3818 VSS 0.148913f
C20960 DVDD.n3819 VSS 0.148913f
C20961 DVDD.n3820 VSS 0.148913f
C20962 DVDD.n3821 VSS 0.148913f
C20963 DVDD.n3822 VSS 0.148913f
C20964 DVDD.n3823 VSS 0.124269f
C20965 DVDD.n3824 VSS 0.148913f
C20966 DVDD.n3825 VSS 0.148913f
C20967 DVDD.n3826 VSS 0.148913f
C20968 DVDD.n3827 VSS 0.148913f
C20969 DVDD.n3828 VSS 0.148913f
C20970 DVDD.n3829 VSS 0.141572f
C20971 DVDD.n3830 VSS 0.141572f
C20972 DVDD.n3831 VSS 0.141572f
C20973 DVDD.n3832 VSS 0.168643f
C20974 DVDD.n3833 VSS 0.416792f
C20975 DVDD.n3834 VSS 0.09543f
C20976 DVDD.n3835 VSS 0.09543f
C20977 DVDD.n3836 VSS 0.09543f
C20978 DVDD.n3837 VSS 0.148913f
C20979 DVDD.n3838 VSS 0.148913f
C20980 DVDD.n3839 VSS 0.148913f
C20981 DVDD.n3840 VSS 0.148913f
C20982 DVDD.n3841 VSS 0.148913f
C20983 DVDD.n3842 VSS 0.148913f
C20984 DVDD.n3843 VSS 0.148913f
C20985 DVDD.n3844 VSS 0.148913f
C20986 DVDD.n3845 VSS 0.148913f
C20987 DVDD.n3846 VSS 0.148913f
C20988 DVDD.n3847 VSS 0.148913f
C20989 DVDD.n3848 VSS 0.148913f
C20990 DVDD.n3849 VSS 0.148913f
C20991 DVDD.n3850 VSS 0.148913f
C20992 DVDD.n3851 VSS 0.148913f
C20993 DVDD.n3852 VSS 0.148913f
C20994 DVDD.n3853 VSS 0.148913f
C20995 DVDD.n3854 VSS 0.09543f
C20996 DVDD.n3855 VSS 0.09543f
C20997 DVDD.n3856 VSS 0.09543f
C20998 DVDD.n3857 VSS 0.148913f
C20999 DVDD.n3858 VSS 0.148913f
C21000 DVDD.n3859 VSS 0.148913f
C21001 DVDD.n3860 VSS 0.148913f
C21002 DVDD.n3861 VSS 0.148913f
C21003 DVDD.n3862 VSS 0.148913f
C21004 DVDD.n3863 VSS 0.148913f
C21005 DVDD.n3864 VSS 0.148913f
C21006 DVDD.n3865 VSS 0.137378f
C21007 DVDD.n3866 VSS 0.137378f
C21008 DVDD.n3867 VSS 0.099625f
C21009 DVDD.n3868 VSS 0.166652f
C21010 DVDD.n3869 VSS 0.417595f
C21011 DVDD.n3870 VSS 0.148913f
C21012 DVDD.n3871 VSS 0.148913f
C21013 DVDD.n3872 VSS 0.148913f
C21014 DVDD.n3873 VSS 0.148913f
C21015 DVDD.n3874 VSS 0.148913f
C21016 DVDD.n3875 VSS 0.148913f
C21017 DVDD.n3876 VSS 0.148913f
C21018 DVDD.n3877 VSS 0.148913f
C21019 DVDD.n3878 VSS 0.148913f
C21020 DVDD.n3879 VSS 0.091236f
C21021 DVDD.n3880 VSS 0.148913f
C21022 DVDD.n3881 VSS 0.148913f
C21023 DVDD.n3882 VSS 0.148913f
C21024 DVDD.n3883 VSS 0.148913f
C21025 DVDD.n3884 VSS 0.148913f
C21026 DVDD.n3885 VSS 0.148913f
C21027 DVDD.n3886 VSS 0.148913f
C21028 DVDD.n3887 VSS 0.148913f
C21029 DVDD.n3888 VSS 0.148913f
C21030 DVDD.n3889 VSS 0.148913f
C21031 DVDD.n3890 VSS 0.148913f
C21032 DVDD.n3891 VSS 0.148913f
C21033 DVDD.n3892 VSS 0.148913f
C21034 DVDD.n3893 VSS 0.148913f
C21035 DVDD.n3894 VSS 0.148913f
C21036 DVDD.n3895 VSS 0.148913f
C21037 DVDD.n3896 VSS 0.148913f
C21038 DVDD.n3897 VSS 0.148913f
C21039 DVDD.n3898 VSS 0.099625f
C21040 DVDD.n3899 VSS 0.099625f
C21041 DVDD.n3900 VSS 0.1784f
C21042 DVDD.n3901 VSS 0.168635f
C21043 DVDD.n3902 VSS 0.434106f
C21044 DVDD.n3903 VSS 0.137378f
C21045 DVDD.n3904 VSS 0.148913f
C21046 DVDD.n3905 VSS 0.148913f
C21047 DVDD.n3906 VSS 0.148913f
C21048 DVDD.n3907 VSS 0.148913f
C21049 DVDD.n3908 VSS 0.148913f
C21050 DVDD.n3909 VSS 0.148913f
C21051 DVDD.n3910 VSS 0.148913f
C21052 DVDD.n3911 VSS 0.148913f
C21053 DVDD.n3912 VSS 0.148913f
C21054 DVDD.n3913 VSS 0.148913f
C21055 DVDD.n3914 VSS 0.148913f
C21056 DVDD.n3915 VSS 0.148913f
C21057 DVDD.n3916 VSS 0.148913f
C21058 DVDD.n3917 VSS 0.148913f
C21059 DVDD.n3918 VSS 0.148913f
C21060 DVDD.n3919 VSS 0.148913f
C21061 DVDD.n3920 VSS 0.12794f
C21062 DVDD.n3921 VSS 0.12794f
C21063 DVDD.n3922 VSS 0.12794f
C21064 DVDD.n3923 VSS 0.214611f
C21065 DVDD.n3924 VSS 0.279212f
C21066 DVDD.n3925 VSS 0.279212f
C21067 DVDD.n3926 VSS 0.279212f
C21068 DVDD.n3927 VSS 0.193679f
C21069 DVDD.t6 VSS 0.040899f
C21070 DVDD.t198 VSS 0.040899f
C21071 DVDD.n3928 VSS 0.081797f
C21072 DVDD.n3929 VSS 0.101855f
C21073 DVDD.n3930 VSS 0.046634f
C21074 DVDD.t87 VSS 0.040899f
C21075 DVDD.t81 VSS 0.040899f
C21076 DVDD.n3931 VSS 0.081797f
C21077 DVDD.n3932 VSS 0.101855f
C21078 DVDD.t214 VSS 0.031969f
C21079 DVDD.n3933 VSS 0.211376f
C21080 DVDD.n3934 VSS 0.279212f
C21081 DVDD.n3935 VSS 0.279212f
C21082 DVDD.n3936 VSS 0.279212f
C21083 DVDD.n3937 VSS 0.279212f
C21084 DVDD.n3938 VSS 0.279212f
C21085 DVDD.n3939 VSS 0.279212f
C21086 DVDD.n3940 VSS 0.279212f
C21087 DVDD.n3941 VSS 0.279212f
C21088 DVDD.n3942 VSS 0.279212f
C21089 DVDD.n3943 VSS 0.279212f
C21090 DVDD.n3944 VSS 0.279212f
C21091 DVDD.n3945 VSS 0.279212f
C21092 DVDD.n3946 VSS 0.279212f
C21093 DVDD.n3947 VSS 0.279212f
C21094 DVDD.n3948 VSS 0.279212f
C21095 DVDD.n3949 VSS 0.279212f
C21096 DVDD.n3950 VSS 0.279212f
C21097 DVDD.n3951 VSS 0.146488f
C21098 DVDD.n3952 VSS 0.214611f
C21099 DVDD.n3953 VSS 0.27233f
C21100 DVDD.n3954 VSS 0.279212f
C21101 DVDD.n3955 VSS 0.279212f
C21102 DVDD.n3956 VSS 0.279212f
C21103 DVDD.n3957 VSS 0.207443f
C21104 DVDD.n3958 VSS 0.151362f
C21105 DVDD.n3959 VSS 0.162851f
C21106 DVDD.t108 VSS 0.0973f
C21107 DVDD.n3960 VSS 0.124781f
C21108 DVDD.n3961 VSS 0.050823f
C21109 DVDD.n3962 VSS 0.055548f
C21110 DVDD.n3963 VSS 0.053943f
C21111 DVDD.t106 VSS 0.0973f
C21112 DVDD.n3964 VSS 0.142981f
C21113 DVDD.n3965 VSS 0.214611f
C21114 DVDD.n3966 VSS 0.22514f
C21115 DVDD.n3967 VSS 0.183848f
C21116 DVDD.n3968 VSS 0.279212f
C21117 DVDD.n3969 VSS 0.279212f
C21118 DVDD.n3970 VSS 0.279212f
C21119 DVDD.n3971 VSS 0.279212f
C21120 DVDD.n3972 VSS 0.178932f
C21121 DVDD.n3973 VSS 0.178932f
C21122 DVDD.n3974 VSS 0.13469f
C21123 DVDD.n3975 VSS 0.214063f
C21124 DVDD.n3976 VSS 0.239887f
C21125 DVDD.n3977 VSS 0.239887f
C21126 DVDD.n3978 VSS 0.239887f
C21127 DVDD.n3979 VSS 0.279212f
C21128 DVDD.n3980 VSS 0.279212f
C21129 DVDD.n3981 VSS 0.279212f
C21130 DVDD.n3982 VSS 0.279212f
C21131 DVDD.n3983 VSS 0.279212f
C21132 DVDD.n3984 VSS 0.279212f
C21133 DVDD.n3985 VSS 0.279212f
C21134 DVDD.n3986 VSS 0.279212f
C21135 DVDD.n3987 VSS 0.279212f
C21136 DVDD.n3988 VSS 0.279212f
C21137 DVDD.n3989 VSS 0.279212f
C21138 DVDD.n3990 VSS 0.279212f
C21139 DVDD.n3991 VSS 0.279212f
C21140 DVDD.n3992 VSS 0.067849f
C21141 DVDD.t42 VSS 0.040899f
C21142 DVDD.t44 VSS 0.040899f
C21143 DVDD.n3993 VSS 0.081797f
C21144 DVDD.n3994 VSS 0.1308f
C21145 DVDD.n3995 VSS 0.216649f
C21146 DVDD.n3996 VSS 0.15632f
C21147 DVDD.n3997 VSS 0.279212f
C21148 DVDD.n3998 VSS 0.279212f
C21149 DVDD.n3999 VSS 0.279212f
C21150 DVDD.n4000 VSS 0.279212f
C21151 DVDD.n4001 VSS 0.279212f
C21152 DVDD.n4002 VSS 0.279212f
C21153 DVDD.n4003 VSS 0.279212f
C21154 DVDD.n4004 VSS 0.279212f
C21155 DVDD.n4005 VSS 0.279212f
C21156 DVDD.n4006 VSS 0.279212f
C21157 DVDD.n4007 VSS 0.279212f
C21158 DVDD.n4008 VSS 0.279212f
C21159 DVDD.n4009 VSS 0.279212f
C21160 DVDD.n4010 VSS 0.266432f
C21161 DVDD.n4011 VSS 0.067849f
C21162 DVDD.t57 VSS 0.040899f
C21163 DVDD.t59 VSS 0.040899f
C21164 DVDD.n4012 VSS 0.081797f
C21165 DVDD.n4013 VSS 0.1308f
C21166 DVDD.n4014 VSS 0.216649f
C21167 DVDD.n4015 VSS 0.152387f
C21168 DVDD.n4016 VSS 0.279212f
C21169 DVDD.n4017 VSS 0.279212f
C21170 DVDD.n4018 VSS 0.279212f
C21171 DVDD.n4019 VSS 0.279212f
C21172 DVDD.n4020 VSS 0.279212f
C21173 DVDD.n4021 VSS 0.279212f
C21174 DVDD.n4022 VSS 0.279212f
C21175 DVDD.n4023 VSS 0.279212f
C21176 DVDD.n4024 VSS 0.279212f
C21177 DVDD.n4025 VSS 0.279212f
C21178 DVDD.n4026 VSS 0.279212f
C21179 DVDD.n4027 VSS 0.279212f
C21180 DVDD.n4028 VSS 0.279212f
C21181 DVDD.n4029 VSS 0.279212f
C21182 DVDD.n4030 VSS 0.279212f
C21183 DVDD.n4031 VSS 0.171067f
C21184 DVDD.n4032 VSS 0.171067f
C21185 DVDD.n4033 VSS 0.214063f
C21186 DVDD.n4034 VSS 0.148913f
C21187 DVDD.n4035 VSS 0.148913f
C21188 DVDD.n4036 VSS 0.148913f
C21189 DVDD.n4037 VSS 0.148913f
C21190 DVDD.n4038 VSS 0.148913f
C21191 DVDD.n4039 VSS 0.148913f
C21192 DVDD.n4040 VSS 0.133183f
C21193 DVDD.n4041 VSS 0.133183f
C21194 DVDD.n4042 VSS 0.10382f
C21195 DVDD.n4043 VSS 0.166758f
C21196 DVDD.n4044 VSS 0.178144f
C21197 DVDD.n4045 VSS 0.148913f
C21198 DVDD.n4046 VSS 0.148913f
C21199 DVDD.n4047 VSS 0.097528f
C21200 DVDD.n4048 VSS 0.148913f
C21201 DVDD.n4049 VSS 0.148913f
C21202 DVDD.n4050 VSS 0.148913f
C21203 DVDD.n4051 VSS 0.148913f
C21204 DVDD.n4052 VSS 0.074652f
C21205 DVDD.n4053 VSS 0.074457f
C21206 DVDD.n4054 VSS 0.007073f
C21207 DVDD.n4055 VSS 0.074457f
C21208 DVDD.n4056 VSS 0.074457f
C21209 DVDD.n4057 VSS 0.074457f
C21210 DVDD.n4058 VSS 0.148913f
C21211 DVDD.n4059 VSS 0.148913f
C21212 DVDD.n4060 VSS 0.148913f
C21213 DVDD.n4061 VSS 0.148913f
C21214 DVDD.n4062 VSS 0.074457f
C21215 DVDD.n4063 VSS 0.074457f
C21216 DVDD.n4064 VSS 0.007073f
C21217 DVDD.n4065 VSS 0.012307f
C21218 DVDD.n4066 VSS 0.074457f
C21219 DVDD.n4067 VSS 0.074457f
C21220 DVDD.n4068 VSS 0.148913f
C21221 DVDD.n4069 VSS 0.148913f
C21222 DVDD.n4070 VSS 0.148913f
C21223 DVDD.n4071 VSS 0.148913f
C21224 DVDD.n4072 VSS 0.148913f
C21225 DVDD.n4073 VSS 0.148913f
C21226 DVDD.n4074 VSS 0.148913f
C21227 DVDD.n4075 VSS 0.148913f
C21228 DVDD.n4076 VSS 0.148913f
C21229 DVDD.n4077 VSS 0.10382f
C21230 DVDD.n4078 VSS 0.10382f
C21231 DVDD.n4079 VSS 0.434046f
C21232 DVDD.n4080 VSS 0.168635f
C21233 DVDD.n4081 VSS 0.417805f
C21234 DVDD.n4082 VSS 0.133183f
C21235 DVDD.n4083 VSS 0.148913f
C21236 DVDD.n4084 VSS 0.148913f
C21237 DVDD.n4085 VSS 0.148913f
C21238 DVDD.n4086 VSS 0.148913f
C21239 DVDD.n4087 VSS 0.148913f
C21240 DVDD.n4088 VSS 0.148913f
C21241 DVDD.n4089 VSS 0.148913f
C21242 DVDD.n4090 VSS 0.148913f
C21243 DVDD.n4091 VSS 0.148913f
C21244 DVDD.n4092 VSS 0.148913f
C21245 DVDD.n4093 VSS 0.148913f
C21246 DVDD.n4094 VSS 0.148913f
C21247 DVDD.n4095 VSS 0.148913f
C21248 DVDD.n4096 VSS 0.148913f
C21249 DVDD.n4097 VSS 0.148913f
C21250 DVDD.n4098 VSS 0.148913f
C21251 DVDD.n4099 VSS 0.132134f
C21252 DVDD.n4100 VSS 0.132134f
C21253 DVDD.n4101 VSS 0.132134f
C21254 DVDD.n4102 VSS 0.214063f
C21255 DVDD.n4103 VSS 0.247752f
C21256 DVDD.n4104 VSS 0.279212f
C21257 DVDD.n4105 VSS 0.279212f
C21258 DVDD.n4106 VSS 0.279212f
C21259 DVDD.n4107 VSS 0.279212f
C21260 DVDD.n4108 VSS 0.279212f
C21261 DVDD.n4109 VSS 0.279212f
C21262 DVDD.n4110 VSS 0.279212f
C21263 DVDD.n4111 VSS 0.279212f
C21264 DVDD.n4112 VSS 0.189746f
C21265 DVDD.n4113 VSS 0.214611f
C21266 DVDD.n4114 VSS 0.229072f
C21267 DVDD.n4115 VSS 0.279212f
C21268 DVDD.n4116 VSS 0.279212f
C21269 DVDD.n4117 VSS 0.279212f
C21270 DVDD.n4118 VSS 0.179915f
C21271 DVDD.n4119 VSS 0.214611f
C21272 DVDD.t64 VSS 0.040899f
C21273 DVDD.t28 VSS 0.040899f
C21274 DVDD.n4120 VSS 0.081797f
C21275 DVDD.n4121 VSS 0.101855f
C21276 DVDD.n4122 VSS 0.046634f
C21277 DVDD.n4123 VSS 0.053943f
C21278 DVDD.n4124 VSS 0.055548f
C21279 DVDD.t186 VSS 0.040899f
C21280 DVDD.t164 VSS 0.040899f
C21281 DVDD.n4125 VSS 0.081797f
C21282 DVDD.n4126 VSS 0.101855f
C21283 DVDD.n4127 VSS 0.214611f
C21284 DVDD.n4128 VSS 0.150421f
C21285 DVDD.n4129 VSS 0.279212f
C21286 DVDD.n4130 VSS 0.279212f
C21287 DVDD.n4131 VSS 0.279212f
C21288 DVDD.n4132 VSS 0.279212f
C21289 DVDD.n4133 VSS 0.279212f
C21290 DVDD.n4134 VSS 0.279212f
C21291 DVDD.n4135 VSS 0.211376f
C21292 DVDD.t166 VSS 0.0973f
C21293 DVDD.n4136 VSS 0.124781f
C21294 DVDD.t219 VSS 0.031969f
C21295 DVDD.n4137 VSS 0.162851f
C21296 DVDD.n4138 VSS 0.151362f
C21297 DVDD.n4139 VSS 0.166151f
C21298 DVDD.n4140 VSS 0.207443f
C21299 DVDD.n4141 VSS 0.279212f
C21300 DVDD.n4142 VSS 0.279212f
C21301 DVDD.n4143 VSS 0.279212f
C21302 DVDD.n4144 VSS 0.279212f
C21303 DVDD.n4145 VSS 0.279212f
C21304 DVDD.n4146 VSS 0.233988f
C21305 DVDD.t205 VSS 0.031969f
C21306 DVDD.n4147 VSS 0.162851f
C21307 DVDD.n4148 VSS 0.151362f
C21308 DVDD.n4149 VSS 0.158286f
C21309 DVDD.n4150 VSS 0.279212f
C21310 DVDD.n4151 VSS 0.279212f
C21311 DVDD.n4152 VSS 0.279212f
C21312 DVDD.n4153 VSS 0.279212f
C21313 DVDD.n4154 VSS 0.279212f
C21314 DVDD.n4155 VSS 0.279212f
C21315 DVDD.n4156 VSS 0.181881f
C21316 DVDD.n4157 VSS 0.214611f
C21317 DVDD.n4158 VSS 0.236937f
C21318 DVDD.n4159 VSS 0.242836f
C21319 DVDD.n4160 VSS 0.279212f
C21320 DVDD.n4161 VSS 0.279212f
C21321 DVDD.n4162 VSS 0.279212f
C21322 DVDD.n4163 VSS 0.279212f
C21323 DVDD.n4164 VSS 0.279212f
C21324 DVDD.n4165 VSS 0.279212f
C21325 DVDD.n4166 VSS 0.175982f
C21326 DVDD.n4167 VSS 0.279212f
C21327 DVDD.n4168 VSS 0.163202f
C21328 DVDD.n4169 VSS 0.163202f
C21329 DVDD.n4170 VSS 0.163202f
C21330 DVDD.n4171 VSS 0.279212f
C21331 DVDD.n4172 VSS 0.279212f
C21332 DVDD.t20 VSS 0.040899f
C21333 DVDD.t112 VSS 0.040899f
C21334 DVDD.n4173 VSS 0.081797f
C21335 DVDD.n4174 VSS 0.129754f
C21336 DVDD.n4175 VSS 0.193053f
C21337 DVDD.n4176 VSS 0.279212f
C21338 DVDD.n4177 VSS 0.279212f
C21339 DVDD.n4178 VSS 0.279212f
C21340 DVDD.n4179 VSS 0.279212f
C21341 DVDD.n4180 VSS 0.279212f
C21342 DVDD.n4181 VSS 0.279212f
C21343 DVDD.n4182 VSS 0.279212f
C21344 DVDD.n4183 VSS 0.279212f
C21345 DVDD.n4184 VSS 0.279212f
C21346 DVDD.n4185 VSS 0.279212f
C21347 DVDD.n4186 VSS 0.279212f
C21348 DVDD.n4187 VSS 0.185814f
C21349 DVDD.n4188 VSS -0.064612f
C21350 DVDD.n4189 VSS 0.260533f
C21351 DVDD.n4190 VSS 0.437245f
C21352 DVDD.n4191 VSS 0.279212f
C21353 DVDD.n4192 VSS 0.279212f
C21354 DVDD.n4193 VSS 0.251684f
C21355 DVDD.n4194 VSS 0.167134f
C21356 DVDD.n4195 VSS 0.167134f
C21357 DVDD.n4196 VSS 0.143539f
C21358 DVDD.n4197 VSS 1.00328f
C21359 DVDD.n4198 VSS 1.23402f
C21360 DVDD.t204 VSS 0.513692f
C21361 DVDD.t132 VSS 0.476895f
C21362 DVDD.t146 VSS 0.476895f
C21363 DVDD.t171 VSS 0.644981f
C21364 DVDD.t19 VSS 0.644981f
C21365 DVDD.t111 VSS 0.379977f
C21366 DVDD.t128 VSS 0.644981f
C21367 DVDD.t36 VSS 0.644981f
C21368 DVDD.t37 VSS 0.476895f
C21369 DVDD.t124 VSS 0.341058f
C21370 DVDD.n4199 VSS 0.497348f
C21371 DVDD.t126 VSS 0.488923f
C21372 DVDD.n4200 VSS 0.581089f
C21373 DVDD.n4201 VSS 0.067483f
C21374 DVDD.t125 VSS 0.040899f
C21375 DVDD.t127 VSS 0.040899f
C21376 DVDD.n4202 VSS 0.081797f
C21377 DVDD.n4203 VSS 0.1308f
C21378 DVDD.n4204 VSS 0.216649f
C21379 DVDD.n4205 VSS 0.205477f
C21380 DVDD.n4206 VSS 0.279212f
C21381 DVDD.n4207 VSS 0.279212f
C21382 DVDD.n4208 VSS 0.279212f
C21383 DVDD.n4209 VSS 0.279212f
C21384 DVDD.n4210 VSS 0.279212f
C21385 DVDD.n4211 VSS 0.279212f
C21386 DVDD.n4212 VSS 0.279212f
C21387 DVDD.n4213 VSS 0.279212f
C21388 DVDD.n4214 VSS 0.279212f
C21389 DVDD.n4215 VSS 0.279212f
C21390 DVDD.n4216 VSS 0.279212f
C21391 DVDD.n4217 VSS 0.279212f
C21392 DVDD.n4218 VSS 0.185814f
C21393 DVDD.n4219 VSS 0.255617f
C21394 DVDD.n4220 VSS 0.255617f
C21395 DVDD.n4221 VSS 0.214063f
C21396 DVDD.n4222 VSS 0.087041f
C21397 DVDD.n4223 VSS 0.087041f
C21398 DVDD.n4224 VSS 0.06397f
C21399 DVDD.n4225 VSS 0.074457f
C21400 DVDD.n4226 VSS 0.005305f
C21401 DVDD.n4227 VSS 0.003537f
C21402 DVDD.n4228 VSS 0.010361f
C21403 DVDD.n4229 VSS 0.050385f
C21404 DVDD.n4230 VSS 0.056902f
C21405 DVDD.n4231 VSS 0.051595f
C21406 DVDD.n4232 VSS 0.038174f
C21407 DVDD.n4233 VSS 0.017911f
C21408 DVDD.n4234 VSS 0.620559f
C21409 DVDD.t165 VSS 0.590255f
C21410 DVDD.t163 VSS 0.476895f
C21411 DVDD.t185 VSS 0.476895f
C21412 DVDD.t183 VSS 0.644981f
C21413 DVDD.t27 VSS 0.644981f
C21414 DVDD.t63 VSS 0.379977f
C21415 DVDD.t51 VSS 0.644981f
C21416 DVDD.t54 VSS 0.644981f
C21417 DVDD.t49 VSS 0.476895f
C21418 DVDD.t58 VSS 0.476895f
C21419 DVDD.t56 VSS 0.590255f
C21420 DVDD.n4235 VSS 1.12635f
C21421 DVDD.t43 VSS 0.590255f
C21422 DVDD.t41 VSS 0.476895f
C21423 DVDD.t47 VSS 0.476895f
C21424 DVDD.t53 VSS 0.644981f
C21425 DVDD.t50 VSS 0.644981f
C21426 DVDD.t197 VSS 0.379977f
C21427 DVDD.t5 VSS 0.644981f
C21428 DVDD.t105 VSS 0.644981f
C21429 DVDD.t80 VSS 0.476895f
C21430 DVDD.t86 VSS 0.476895f
C21431 DVDD.t107 VSS 0.590255f
C21432 DVDD.n4236 VSS 0.620559f
C21433 DVDD.n4237 VSS 0.017911f
C21434 DVDD.n4238 VSS 0.236283f
C21435 DVDD.n4239 VSS 0.233988f
C21436 DVDD.n4240 VSS 0.279212f
C21437 DVDD.n4241 VSS 0.279212f
C21438 DVDD.n4242 VSS 0.279212f
C21439 DVDD.n4243 VSS 0.279212f
C21440 DVDD.n4244 VSS 0.279212f
C21441 DVDD.n4245 VSS 0.177949f
C21442 DVDD.n4246 VSS 0.279212f
C21443 DVDD.n4247 VSS 0.279212f
C21444 DVDD.n4248 VSS 0.24087f
C21445 DVDD.n4249 VSS 0.279212f
C21446 DVDD.n4250 VSS 0.238904f
C21447 DVDD.n4251 VSS 0.279212f
C21448 DVDD.n4252 VSS 0.279212f
C21449 DVDD.n4253 VSS 0.179915f
C21450 DVDD.n4254 VSS 0.279212f
C21451 DVDD.n4255 VSS 0.229072f
C21452 DVDD.n4256 VSS 0.232022f
C21453 DVDD.n4257 VSS 0.232022f
C21454 DVDD.n4258 VSS 0.214063f
C21455 DVDD.n4259 VSS 0.099625f
C21456 DVDD.n4260 VSS 0.099625f
C21457 DVDD.n4261 VSS 0.074457f
C21458 DVDD.n4262 VSS 0.074457f
C21459 DVDD.n4263 VSS 0.007073f
C21460 DVDD.n4264 VSS 0.007073f
C21461 DVDD.n4265 VSS 0.074457f
C21462 DVDD.n4266 VSS 0.074457f
C21463 DVDD.n4267 VSS 0.148913f
C21464 DVDD.n4268 VSS 0.148913f
C21465 DVDD.n4269 VSS 0.148913f
C21466 DVDD.n4270 VSS 0.148913f
C21467 DVDD.n4271 VSS 0.148913f
C21468 DVDD.n4272 VSS 0.099101f
C21469 DVDD.n4273 VSS 0.148913f
C21470 DVDD.n4274 VSS 0.148913f
C21471 DVDD.n4275 VSS 0.148913f
C21472 DVDD.n4276 VSS 0.148913f
C21473 DVDD.n4277 VSS 0.148913f
C21474 DVDD.n4278 VSS 0.148913f
C21475 DVDD.n4279 VSS 0.148913f
C21476 DVDD.n4280 VSS 0.148913f
C21477 DVDD.n4281 VSS 0.148913f
C21478 DVDD.n4282 VSS 0.091236f
C21479 DVDD.n4283 VSS 0.091236f
C21480 DVDD.n4284 VSS 0.091236f
C21481 DVDD.n4285 VSS 0.056938f
C21482 DVDD.n4286 VSS 0.061371f
C21483 DVDD.n4287 VSS 0.061371f
C21484 DVDD.n4288 VSS 0.04016f
C21485 DVDD.n4289 VSS 0.04016f
C21486 DVDD.n4290 VSS 0.037228f
C21487 DVDD.n4291 VSS 0.037228f
C21488 DVDD.n4292 VSS 0.04016f
C21489 DVDD.n4293 VSS 0.04016f
C21490 DVDD.n4294 VSS 0.04016f
C21491 DVDD.n4295 VSS 0.08032f
C21492 DVDD.n4296 VSS 0.228989f
C21493 DVDD.n4297 VSS 0.075834f
C21494 DVDD.n4298 VSS 0.074152f
C21495 DVDD.n4299 VSS 0.273051f
C21496 DVDD.n4300 VSS 0.532172f
C21497 DVDD.n4301 VSS 1.0352f
C21498 DVDD.n4302 VSS 0.279212f
C21499 DVDD.n4303 VSS 0.279212f
C21500 DVDD.n4304 VSS 0.279212f
C21501 DVDD.n4305 VSS 0.279212f
C21502 DVDD.n4306 VSS 0.279212f
C21503 DVDD.n4307 VSS 0.279212f
C21504 DVDD.n4308 VSS 0.279212f
C21505 DVDD.n4309 VSS 0.279212f
C21506 DVDD.n4310 VSS 0.279212f
C21507 DVDD.n4311 VSS 0.188763f
C21508 DVDD.n4312 VSS 0.279212f
C21509 DVDD.n4313 VSS 0.279212f
C21510 DVDD.n4314 VSS 0.279212f
C21511 DVDD.n4315 VSS 0.279212f
C21512 DVDD.n4316 VSS 0.279212f
C21513 DVDD.n4317 VSS 0.279212f
C21514 DVDD.n4318 VSS 0.279212f
C21515 DVDD.n4319 VSS 0.279212f
C21516 DVDD.n4320 VSS 0.279212f
C21517 DVDD.n4321 VSS 0.279212f
C21518 DVDD.n4322 VSS 0.279212f
C21519 DVDD.n4323 VSS 0.279212f
C21520 DVDD.n4324 VSS 0.279212f
C21521 DVDD.n4325 VSS 0.279212f
C21522 DVDD.n4326 VSS 0.279212f
C21523 DVDD.n4327 VSS 0.279212f
C21524 DVDD.n4328 VSS 0.279212f
C21525 DVDD.n4329 VSS 0.279212f
C21526 DVDD.n4330 VSS 0.139606f
C21527 DVDD.n4340 VSS 0.139606f
C21528 DVDD.n4342 VSS 0.273051f
C21529 DVDD.n4343 VSS 0.139606f
C21530 DVDD.n4344 VSS 0.065805f
C21531 DVDD.n4345 VSS 0.532172f
C21532 DVDD.n4346 VSS 1.0352f
C21533 DVDD.n4347 VSS 0.279212f
C21534 DVDD.n4348 VSS 0.279212f
C21535 DVDD.n4349 VSS 0.279212f
C21536 DVDD.n4350 VSS 0.279212f
C21537 DVDD.n4351 VSS 0.279212f
C21538 DVDD.n4352 VSS 0.279212f
C21539 DVDD.n4353 VSS 0.279212f
C21540 DVDD.n4354 VSS 0.279212f
C21541 DVDD.n4355 VSS 0.279212f
C21542 DVDD.n4356 VSS 0.279212f
C21543 DVDD.n4357 VSS 0.279212f
C21544 DVDD.n4358 VSS 0.279212f
C21545 DVDD.n4359 VSS 0.279212f
C21546 DVDD.n4360 VSS 0.279212f
C21547 DVDD.n4361 VSS 0.279212f
C21548 DVDD.n4362 VSS 0.279212f
C21549 DVDD.n4363 VSS 0.279212f
C21550 DVDD.n4364 VSS 0.279212f
C21551 DVDD.n4365 VSS 0.279212f
C21552 DVDD.n4366 VSS 0.279212f
C21553 DVDD.n4367 VSS 0.279212f
C21554 DVDD.n4368 VSS 0.279212f
C21555 DVDD.n4369 VSS 0.279212f
C21556 DVDD.n4370 VSS 0.279212f
C21557 DVDD.n4371 VSS 0.279212f
C21558 DVDD.n4372 VSS 0.279212f
C21559 DVDD.n4373 VSS 0.139606f
C21560 DVDD.n4383 VSS 0.139606f
C21561 DVDD.n4385 VSS 0.065805f
C21562 DVDD.n4386 VSS 0.139606f
C21563 DVDD.n4387 VSS 0.065805f
C21564 DVDD.n4398 VSS 0.139606f
C21565 DVDD.n4399 VSS 0.532172f
C21566 DVDD.n4409 VSS 0.279212f
C21567 DVDD.n4410 VSS 0.139606f
C21568 DVDD.n4411 VSS 0.624053f
C21569 DVDD.n4413 VSS 0.065805f
C21570 DVDD.n4414 VSS 0.139606f
C21571 DVDD.n4415 VSS 0.15632f
C21572 DVDD.n4416 VSS 0.279212f
C21573 DVDD.n4417 VSS 0.279212f
C21574 DVDD.n4418 VSS 0.279212f
C21575 DVDD.n4419 VSS 0.279212f
C21576 DVDD.n4420 VSS 0.279212f
C21577 DVDD.n4421 VSS 0.279212f
C21578 DVDD.n4422 VSS 0.279212f
C21579 DVDD.n4423 VSS 0.279212f
C21580 DVDD.n4424 VSS 0.279212f
C21581 DVDD.n4425 VSS 0.279212f
C21582 DVDD.n4426 VSS 0.279212f
C21583 DVDD.n4427 VSS 0.279212f
C21584 DVDD.n4428 VSS 0.279212f
C21585 DVDD.n4429 VSS 0.279212f
C21586 DVDD.n4430 VSS 0.279212f
C21587 DVDD.n4431 VSS 0.198595f
C21588 DVDD.n4432 VSS 0.279212f
C21589 DVDD.n4433 VSS 0.279212f
C21590 DVDD.n4434 VSS 0.279212f
C21591 DVDD.n4435 VSS 0.279212f
C21592 DVDD.n4436 VSS 0.279212f
C21593 DVDD.n4437 VSS 0.279212f
C21594 DVDD.n4438 VSS 0.186797f
C21595 DVDD.n4439 VSS 0.186797f
C21596 DVDD.n4440 VSS 0.532863f
C21597 DVDD.n4441 VSS 0.232022f
C21598 DVDD.n4442 VSS 0.232022f
C21599 DVDD.n4443 VSS 0.232022f
C21600 DVDD.n4444 VSS 0.279212f
C21601 DVDD.n4445 VSS 0.279212f
C21602 DVDD.n4446 VSS 0.279212f
C21603 DVDD.n4447 VSS 0.279212f
C21604 DVDD.n4448 VSS 0.279212f
C21605 DVDD.n4449 VSS 0.279212f
C21606 DVDD.n4450 VSS 0.279212f
C21607 DVDD.n4451 VSS 0.279212f
C21608 DVDD.n4452 VSS 0.279212f
C21609 DVDD.n4453 VSS 0.279212f
C21610 DVDD.n4454 VSS 0.279212f
C21611 DVDD.n4455 VSS 0.279212f
C21612 DVDD.n4456 VSS 0.279212f
C21613 DVDD.n4457 VSS 0.279212f
C21614 DVDD.n4458 VSS 0.279212f
C21615 DVDD.n4459 VSS 0.279212f
C21616 DVDD.n4460 VSS 0.279212f
C21617 DVDD.n4461 VSS 0.279212f
C21618 DVDD.n4462 VSS 0.279212f
C21619 DVDD.n4463 VSS 0.279212f
C21620 DVDD.n4464 VSS 0.279212f
C21621 DVDD.n4465 VSS 0.279212f
C21622 DVDD.n4466 VSS 0.279212f
C21623 DVDD.n4467 VSS 0.279212f
C21624 DVDD.n4468 VSS 0.279212f
C21625 DVDD.n4469 VSS 0.279212f
C21626 DVDD.n4470 VSS 0.279212f
C21627 DVDD.n4471 VSS 0.279212f
C21628 DVDD.n4472 VSS 0.279212f
C21629 DVDD.n4473 VSS 0.279212f
C21630 DVDD.n4474 VSS 0.279212f
C21631 DVDD.n4475 VSS 0.279212f
C21632 DVDD.n4476 VSS 0.279212f
C21633 DVDD.n4477 VSS 0.279212f
C21634 DVDD.n4478 VSS 0.279212f
C21635 DVDD.n4479 VSS 0.279212f
C21636 DVDD.n4480 VSS 0.217274f
C21637 DVDD.n4481 VSS 0.279212f
C21638 DVDD.n4482 VSS 0.279212f
C21639 DVDD.n4483 VSS 0.279212f
C21640 DVDD.n4484 VSS 0.279212f
C21641 DVDD.n4485 VSS 0.279212f
C21642 DVDD.n4486 VSS 0.279212f
C21643 DVDD.n4487 VSS 0.279212f
C21644 DVDD.n4488 VSS 0.279212f
C21645 DVDD.n4489 VSS 0.279212f
C21646 DVDD.n4490 VSS 0.279212f
C21647 DVDD.n4491 VSS 0.279212f
C21648 DVDD.n4492 VSS 0.279212f
C21649 DVDD.n4493 VSS 0.279212f
C21650 DVDD.n4494 VSS 0.264465f
C21651 DVDD.n4495 VSS 0.279212f
C21652 DVDD.n4496 VSS 0.279212f
C21653 DVDD.n4497 VSS 0.139606f
C21654 DVDD.n4498 VSS 0.009915f
C21655 DVDD.n4499 VSS 0.009915f
C21656 DVDD.n4500 VSS 0.009915f
C21657 DVDD.n4501 VSS 0.009915f
C21658 DVDD.n4502 VSS 0.009915f
C21659 DVDD.n4503 VSS 0.009915f
C21660 DVDD.n4504 VSS 0.009915f
C21661 DVDD.n4505 VSS 0.009915f
C21662 DVDD.n4506 VSS 0.009915f
C21663 DVDD.n4507 VSS 0.011355f
C21664 DVDD.n4508 VSS 0.019831f
C21665 DVDD.n4509 VSS 0.011115f
C21666 DVDD.n4510 VSS 0.010155f
C21667 DVDD.n4511 VSS 0.019831f
C21668 DVDD.n4512 VSS 0.011355f
C21669 DVDD.n4513 VSS 0.019831f
C21670 DVDD.n4514 VSS 0.011355f
C21671 DVDD.n4515 VSS 0.019831f
C21672 DVDD.n4516 VSS 0.011355f
C21673 DVDD.n4517 VSS 0.019831f
C21674 DVDD.n4518 VSS 0.011355f
C21675 DVDD.n4519 VSS 0.019831f
C21676 DVDD.n4520 VSS 0.011355f
C21677 DVDD.n4521 VSS 0.019831f
C21678 DVDD.n4522 VSS 0.011355f
C21679 DVDD.n4523 VSS 0.019831f
C21680 DVDD.n4524 VSS 0.019831f
C21681 DVDD.n4525 VSS 0.010955f
C21682 DVDD.n4526 VSS 0.010315f
C21683 DVDD.n4527 VSS 0.019831f
C21684 DVDD.n4528 VSS 0.011355f
C21685 DVDD.n4529 VSS 0.019831f
C21686 DVDD.n4530 VSS 0.011355f
C21687 DVDD.n4531 VSS 0.019831f
C21688 DVDD.n4532 VSS 0.011355f
C21689 DVDD.n4533 VSS 0.019831f
C21690 DVDD.n4534 VSS 0.011355f
C21691 DVDD.n4535 VSS 0.019831f
C21692 DVDD.n4536 VSS 0.011355f
C21693 DVDD.n4537 VSS 0.019831f
C21694 DVDD.n4538 VSS 0.011355f
C21695 DVDD.n4539 VSS 0.019831f
C21696 DVDD.n4540 VSS 0.019831f
C21697 DVDD.n4541 VSS 0.010795f
C21698 DVDD.n4542 VSS 0.010475f
C21699 DVDD.n4543 VSS 0.019831f
C21700 DVDD.n4544 VSS 0.011355f
C21701 DVDD.n4545 VSS 0.019831f
C21702 DVDD.n4546 VSS 0.019831f
C21703 DVDD.n4547 VSS 0.019831f
C21704 DVDD.n4548 VSS 0.011355f
C21705 DVDD.n4549 VSS 0.0615f
C21706 DVDD.n4550 VSS 0.011355f
C21707 DVDD.n4551 VSS 0.019831f
C21708 DVDD.n4552 VSS 0.019831f
C21709 DVDD.n4553 VSS 0.014873f
C21710 DVDD.n4554 VSS 0.019831f
C21711 DVDD.n4555 VSS 0.014953f
C21712 DVDD.n4556 VSS 0.019831f
C21713 DVDD.n4557 VSS 0.019831f
C21714 DVDD.n4558 VSS 0.011355f
C21715 DVDD.n4559 VSS 0.009915f
C21716 DVDD.n4560 VSS 0.139606f
C21717 DVDD.n4561 VSS 0.009915f
C21718 DVDD.n4562 VSS 0.011355f
C21719 DVDD.n4563 VSS 0.019831f
C21720 DVDD.n4564 VSS 0.019831f
C21721 DVDD.n4565 VSS 0.015753f
C21722 DVDD.n4566 VSS 0.019831f
C21723 DVDD.n4567 VSS 0.011994f
C21724 DVDD.n4568 VSS -0.359726f
C21725 DVDD.n4569 VSS 0.011355f
C21726 DVDD.n4570 VSS 0.019831f
C21727 DVDD.n4571 VSS 0.011355f
C21728 DVDD.n4572 VSS 0.019831f
C21729 DVDD.n4573 VSS 0.011355f
C21730 DVDD.n4574 VSS 0.019831f
C21731 DVDD.n4575 VSS 0.011355f
C21732 DVDD.n4576 VSS 0.019831f
C21733 DVDD.n4577 VSS 0.011355f
C21734 DVDD.n4578 VSS 0.019831f
C21735 DVDD.n4579 VSS 0.019831f
C21736 DVDD.n4580 VSS 0.010555f
C21737 DVDD.n4581 VSS 0.010715f
C21738 DVDD.n4582 VSS 0.019831f
C21739 DVDD.n4583 VSS 0.011355f
C21740 DVDD.n4584 VSS 0.019831f
C21741 DVDD.n4585 VSS 0.011355f
C21742 DVDD.n4586 VSS 0.019831f
C21743 DVDD.n4587 VSS 0.011355f
C21744 DVDD.n4588 VSS 0.019831f
C21745 DVDD.n4589 VSS 0.011355f
C21746 DVDD.n4590 VSS 0.019831f
C21747 DVDD.n4591 VSS 0.011355f
C21748 DVDD.n4592 VSS 0.019831f
C21749 DVDD.n4593 VSS 0.011355f
C21750 DVDD.n4594 VSS 0.019831f
C21751 DVDD.n4595 VSS 0.019831f
C21752 DVDD.n4596 VSS 0.010395f
C21753 DVDD.n4597 VSS 0.010875f
C21754 DVDD.n4598 VSS 0.019831f
C21755 DVDD.n4599 VSS 0.011355f
C21756 DVDD.n4600 VSS 0.019831f
C21757 DVDD.n4601 VSS 0.011355f
C21758 DVDD.n4602 VSS 0.019831f
C21759 DVDD.n4603 VSS 0.011355f
C21760 DVDD.n4604 VSS 0.019831f
C21761 DVDD.n4605 VSS 0.011355f
C21762 DVDD.n4606 VSS 0.019831f
C21763 DVDD.n4607 VSS 0.011355f
C21764 DVDD.n4608 VSS 0.019831f
C21765 DVDD.n4609 VSS 0.011355f
C21766 DVDD.n4610 VSS 0.019831f
C21767 DVDD.n4611 VSS 0.019831f
C21768 DVDD.n4612 VSS 0.019831f
C21769 DVDD.n4613 VSS 0.011035f
C21770 DVDD.n4614 VSS 0.009915f
C21771 DVDD.n4615 VSS 0.139606f
C21772 DVDD.n4616 VSS 0.139606f
C21773 DVDD.n4617 VSS 0.279212f
C21774 DVDD.n4618 VSS 0.279212f
C21775 DVDD.n4619 VSS 0.154353f
C21776 DVDD.n4620 VSS 0.279212f
C21777 DVDD.n4621 VSS 0.279212f
C21778 DVDD.n4622 VSS 0.279212f
C21779 DVDD.n4623 VSS 0.279212f
C21780 DVDD.n4624 VSS 0.279212f
C21781 DVDD.n4625 VSS 0.279212f
C21782 DVDD.n4626 VSS 0.279212f
C21783 DVDD.n4627 VSS 0.279212f
C21784 DVDD.n4628 VSS 0.279212f
C21785 DVDD.n4629 VSS 0.279212f
C21786 DVDD.n4630 VSS 0.279212f
C21787 DVDD.n4631 VSS 0.279212f
C21788 DVDD.n4632 VSS 0.279212f
C21789 DVDD.n4633 VSS 0.232022f
C21790 DVDD.n4634 VSS 0.232022f
C21791 DVDD.n4635 VSS 0.532863f
C21792 DVDD.n4636 VSS 0.095365f
C21793 DVDD.n4637 VSS 0.186797f
C21794 DVDD.n4638 VSS 0.139606f
C21795 DVDD.n4639 VSS 0.279212f
C21796 DVDD.n4640 VSS 0.17205f
C21797 DVDD.n4641 VSS 0.279212f
C21798 DVDD.n4642 VSS 0.279212f
C21799 DVDD.n4643 VSS 0.139606f
C21800 DVDD.n4644 VSS 0.027037f
C21801 DVDD.n4645 VSS 0.02361f
C21802 DVDD.n4646 VSS 0.02361f
C21803 DVDD.n4647 VSS 0.02361f
C21804 DVDD.n4648 VSS 0.02361f
C21805 DVDD.n4649 VSS 0.02361f
C21806 DVDD.n4650 VSS 0.02361f
C21807 DVDD.n4651 VSS 0.02361f
C21808 DVDD.n4652 VSS 0.02361f
C21809 DVDD.n4653 VSS 0.02361f
C21810 DVDD.n4654 VSS 0.024371f
C21811 DVDD.n4655 VSS 0.070301f
C21812 DVDD.n4656 VSS 0.027037f
C21813 DVDD.n4657 VSS 0.070301f
C21814 DVDD.n4658 VSS 0.027037f
C21815 DVDD.n4659 VSS 0.070301f
C21816 DVDD.n4660 VSS 0.027037f
C21817 DVDD.n4661 VSS 0.070301f
C21818 DVDD.n4662 VSS 0.027037f
C21819 DVDD.n4663 VSS 0.070301f
C21820 DVDD.n4664 VSS 0.070301f
C21821 DVDD.n4665 VSS 0.025133f
C21822 DVDD.n4666 VSS 0.025514f
C21823 DVDD.n4667 VSS 0.070301f
C21824 DVDD.n4668 VSS 0.027037f
C21825 DVDD.n4669 VSS 0.070301f
C21826 DVDD.n4670 VSS 0.027037f
C21827 DVDD.n4671 VSS 0.070301f
C21828 DVDD.n4672 VSS 0.027037f
C21829 DVDD.n4673 VSS 0.070301f
C21830 DVDD.n4674 VSS 0.027037f
C21831 DVDD.n4675 VSS 0.058395f
C21832 DVDD.n4676 VSS 0.035151f
C21833 DVDD.n4677 VSS 0.027037f
C21834 DVDD.n4678 VSS 0.047056f
C21835 DVDD.n4679 VSS 0.027037f
C21836 DVDD.n4680 VSS 0.070301f
C21837 DVDD.n4681 VSS 0.070301f
C21838 DVDD.n4682 VSS 0.024752f
C21839 DVDD.n4683 VSS 0.025895f
C21840 DVDD.n4684 VSS 0.070301f
C21841 DVDD.n4685 VSS 0.027037f
C21842 DVDD.n4686 VSS 0.070301f
C21843 DVDD.n4687 VSS 0.027037f
C21844 DVDD.n4688 VSS 0.070301f
C21845 DVDD.n4689 VSS 0.027037f
C21846 DVDD.n4690 VSS 0.070301f
C21847 DVDD.n4691 VSS 0.027037f
C21848 DVDD.n4692 VSS 0.070301f
C21849 DVDD.n4693 VSS 0.027037f
C21850 DVDD.n4694 VSS 0.070301f
C21851 DVDD.n4695 VSS 0.070301f
C21852 DVDD.n4696 VSS 0.027037f
C21853 DVDD.n4697 VSS 0.02361f
C21854 DVDD.n4698 VSS 0.139606f
C21855 DVDD.n4699 VSS 0.026094f
C21856 DVDD.n4700 VSS 0.024841f
C21857 DVDD.n4701 VSS 0.070301f
C21858 DVDD.n4702 VSS 0.070301f
C21859 DVDD.n4703 VSS 0.070301f
C21860 DVDD.n4704 VSS 0.03134f
C21861 DVDD.n4705 VSS 0.023609f
C21862 DVDD.n4706 VSS 0.090449f
C21863 DVDD.n4707 VSS 0.129775f
C21864 DVDD.n4708 VSS 0.058989f
C21865 DVDD.n4709 VSS 0.026575f
C21866 DVDD.n4710 VSS 0.091432f
C21867 DVDD.n4711 VSS 0.129775f
C21868 DVDD.n4712 VSS 0.279212f
C21869 DVDD.n4713 VSS 0.279212f
C21870 DVDD.n4714 VSS 0.279212f
C21871 DVDD.n4715 VSS 0.186797f
C21872 DVDD.n4716 VSS 0.186797f
C21873 DVDD.n4717 VSS 0.095365f
C21874 DVDD.n4718 VSS 0.336235f
C21875 DVDD.n4719 VSS 0.232022f
C21876 DVDD.n4720 VSS 0.232022f
C21877 DVDD.n4721 VSS 0.232022f
C21878 DVDD.n4722 VSS 0.279212f
C21879 DVDD.n4723 VSS 0.279212f
C21880 DVDD.n4724 VSS 0.279212f
C21881 DVDD.n4725 VSS 0.279212f
C21882 DVDD.n4726 VSS 0.279212f
C21883 DVDD.n4727 VSS 0.279212f
C21884 DVDD.n4728 VSS 0.279212f
C21885 DVDD.n4729 VSS 0.279212f
C21886 DVDD.n4730 VSS 0.279212f
C21887 DVDD.n4731 VSS 0.279212f
C21888 DVDD.n4732 VSS 0.279212f
C21889 DVDD.n4733 VSS 0.279212f
C21890 DVDD.n4734 VSS 0.279212f
C21891 DVDD.n4735 VSS 0.279212f
C21892 DVDD.n4736 VSS 0.279212f
C21893 DVDD.n4737 VSS 0.279212f
C21894 DVDD.n4738 VSS 0.279212f
C21895 DVDD.n4739 VSS 0.279212f
C21896 DVDD.n4740 VSS 0.279212f
C21897 DVDD.n4741 VSS 0.154353f
C21898 DVDD.n4742 VSS 0.139606f
C21899 DVDD.n4743 VSS 0.027427f
C21900 DVDD.n4744 VSS 0.139606f
C21901 DVDD.n4745 VSS 0.264465f
C21902 DVDD.n4746 VSS 0.279212f
C21903 DVDD.n4747 VSS 0.279212f
C21904 DVDD.n4748 VSS 0.279212f
C21905 DVDD.n4749 VSS 0.279212f
C21906 DVDD.n4750 VSS 0.279212f
C21907 DVDD.n4751 VSS 0.279212f
C21908 DVDD.n4752 VSS 0.279212f
C21909 DVDD.n4753 VSS 0.279212f
C21910 DVDD.n4754 VSS 0.279212f
C21911 DVDD.n4755 VSS 0.279212f
C21912 DVDD.n4756 VSS 0.279212f
C21913 DVDD.n4757 VSS 0.279212f
C21914 DVDD.n4758 VSS 0.279212f
C21915 DVDD.n4759 VSS 0.279212f
C21916 DVDD.n4760 VSS 0.279212f
C21917 DVDD.n4761 VSS 0.279212f
C21918 DVDD.n4762 VSS 0.279212f
C21919 DVDD.n4763 VSS 0.279212f
C21920 DVDD.n4764 VSS 0.279212f
C21921 DVDD.n4765 VSS 0.336235f
C21922 DVDD.n4766 VSS 0.178932f
C21923 DVDD.n4767 VSS 0.279212f
C21924 DVDD.n4768 VSS 0.279212f
C21925 DVDD.n4769 VSS 0.217274f
C21926 DVDD.n4770 VSS 0.101264f
C21927 DVDD.n4771 VSS 0.139606f
C21928 DVDD.n4772 VSS 0.027427f
C21929 DVDD.n4773 VSS 0.100281f
C21930 DVDD.n4774 VSS 0.279212f
C21931 DVDD.n4775 VSS 0.279212f
C21932 DVDD.n4776 VSS 0.279212f
C21933 DVDD.n4777 VSS 0.279212f
C21934 DVDD.n4778 VSS 0.279212f
C21935 DVDD.n4779 VSS 0.279212f
C21936 DVDD.n4780 VSS 0.279212f
C21937 DVDD.n4781 VSS 0.279212f
C21938 DVDD.n4782 VSS 0.279212f
C21939 DVDD.n4783 VSS 0.279212f
C21940 DVDD.n4784 VSS 0.279212f
C21941 DVDD.n4785 VSS 0.279212f
C21942 DVDD.n4786 VSS 0.279212f
C21943 DVDD.n4787 VSS 0.279212f
C21944 DVDD.n4788 VSS 0.279212f
C21945 DVDD.n4789 VSS 0.279212f
C21946 DVDD.n4790 VSS 0.279212f
C21947 DVDD.n4791 VSS 0.279212f
C21948 DVDD.n4792 VSS 0.279212f
C21949 DVDD.n4793 VSS 0.279212f
C21950 DVDD.n4794 VSS 0.279212f
C21951 DVDD.n4795 VSS 0.279212f
C21952 DVDD.n4796 VSS 0.279212f
C21953 DVDD.n4797 VSS 0.279212f
C21954 DVDD.n4798 VSS 0.279212f
C21955 DVDD.n4799 VSS 0.279212f
C21956 DVDD.n4800 VSS 0.201544f
C21957 DVDD.n4801 VSS 0.239887f
C21958 DVDD.n4802 VSS 0.336235f
C21959 DVDD.n4803 VSS 0.239887f
C21960 DVDD.n4804 VSS 0.279212f
C21961 DVDD.n4805 VSS 0.279212f
C21962 DVDD.n4806 VSS 0.279212f
C21963 DVDD.n4807 VSS 0.279212f
C21964 DVDD.n4808 VSS 0.279212f
C21965 DVDD.n4809 VSS 0.279212f
C21966 DVDD.n4810 VSS 0.279212f
C21967 DVDD.n4811 VSS 0.279212f
C21968 DVDD.n4812 VSS 0.279212f
C21969 DVDD.n4813 VSS 0.279212f
C21970 DVDD.n4814 VSS 0.279212f
C21971 DVDD.n4815 VSS 0.279212f
C21972 DVDD.n4816 VSS 0.279212f
C21973 DVDD.n4817 VSS 0.279212f
C21974 DVDD.n4818 VSS 0.279212f
C21975 DVDD.n4819 VSS 0.279212f
C21976 DVDD.n4820 VSS 0.279212f
C21977 DVDD.n4821 VSS 0.279212f
C21978 DVDD.n4822 VSS 0.279212f
C21979 DVDD.n4823 VSS 0.279212f
C21980 DVDD.n4824 VSS 0.279212f
C21981 DVDD.n4825 VSS 0.279212f
C21982 DVDD.n4826 VSS 0.279212f
C21983 DVDD.n4827 VSS 0.279212f
C21984 DVDD.n4828 VSS 0.279212f
C21985 DVDD.n4829 VSS 0.279212f
C21986 DVDD.n4830 VSS 0.279212f
C21987 DVDD.n4831 VSS 0.279212f
C21988 DVDD.n4832 VSS 0.279212f
C21989 DVDD.n4833 VSS 0.171067f
C21990 DVDD.n4834 VSS 0.279212f
C21991 DVDD.n4835 VSS 0.279212f
C21992 DVDD.n4836 VSS 0.171067f
C21993 DVDD.n4837 VSS 0.279212f
C21994 DVDD.n4838 VSS 0.279212f
C21995 DVDD.n4839 VSS 0.279212f
C21996 DVDD.n4840 VSS 0.279212f
C21997 DVDD.n4841 VSS 0.279212f
C21998 DVDD.n4842 VSS 0.279212f
C21999 DVDD.n4843 VSS 0.279212f
C22000 DVDD.n4844 VSS 0.279212f
C22001 DVDD.n4845 VSS 0.279212f
C22002 DVDD.n4846 VSS 0.279212f
C22003 DVDD.n4847 VSS 0.279212f
C22004 DVDD.n4848 VSS 0.279212f
C22005 DVDD.n4849 VSS 0.279212f
C22006 DVDD.n4850 VSS 0.278229f
C22007 DVDD.n4851 VSS 0.279212f
C22008 DVDD.n4852 VSS 0.279212f
C22009 DVDD.n4853 VSS 0.279212f
C22010 DVDD.n4854 VSS 0.279212f
C22011 DVDD.n4855 VSS 0.279212f
C22012 DVDD.n4856 VSS 0.279212f
C22013 DVDD.n4857 VSS 0.279212f
C22014 DVDD.n4858 VSS 0.279212f
C22015 DVDD.n4859 VSS 0.279212f
C22016 DVDD.n4860 VSS 0.279212f
C22017 DVDD.n4861 VSS 0.279212f
C22018 DVDD.n4862 VSS 0.279212f
C22019 DVDD.n4863 VSS 0.279212f
C22020 DVDD.n4864 VSS 0.279212f
C22021 DVDD.n4865 VSS 0.279212f
C22022 DVDD.n4866 VSS 0.279212f
C22023 DVDD.n4867 VSS 0.279212f
C22024 DVDD.n4868 VSS 0.279212f
C22025 DVDD.n4869 VSS 0.279212f
C22026 DVDD.n4870 VSS 0.239887f
C22027 DVDD.n4871 VSS 0.532863f
C22028 DVDD.n4872 VSS 0.178932f
C22029 DVDD.n4873 VSS 0.279212f
C22030 DVDD.n4874 VSS 0.217274f
C22031 DVDD.n4875 VSS 0.139606f
C22032 DVDD.n4876 VSS 0.009915f
C22033 DVDD.n4877 VSS 0.100281f
C22034 DVDD.n4878 VSS 0.470925f
C22035 DVDD.n4879 VSS 0.470925f
C22036 DVDD.n4880 VSS 0.101264f
C22037 DVDD.n4881 VSS 0.178932f
C22038 DVDD.n4882 VSS 0.178932f
C22039 DVDD.n4883 VSS 0.532863f
C22040 DVDD.n4884 VSS 0.239887f
C22041 DVDD.n4885 VSS 0.239887f
C22042 DVDD.n4886 VSS 0.201544f
C22043 DVDD.n4887 VSS 0.279212f
C22044 DVDD.n4888 VSS 0.279212f
C22045 DVDD.n4889 VSS 0.279212f
C22046 DVDD.n4890 VSS 0.279212f
C22047 DVDD.n4891 VSS 0.279212f
C22048 DVDD.n4892 VSS 0.279212f
C22049 DVDD.n4893 VSS 0.279212f
C22050 DVDD.n4894 VSS 0.279212f
C22051 DVDD.n4895 VSS 0.279212f
C22052 DVDD.n4896 VSS 0.279212f
C22053 DVDD.n4897 VSS 0.279212f
C22054 DVDD.n4898 VSS 0.279212f
C22055 DVDD.n4899 VSS 0.279212f
C22056 DVDD.n4900 VSS 0.279212f
C22057 DVDD.n4901 VSS 0.279212f
C22058 DVDD.n4902 VSS 0.279212f
C22059 DVDD.n4903 VSS 0.279212f
C22060 DVDD.n4904 VSS 0.279212f
C22061 DVDD.n4905 VSS 0.279212f
C22062 DVDD.n4906 VSS 0.279212f
C22063 DVDD.n4907 VSS 0.279212f
C22064 DVDD.n4908 VSS 0.279212f
C22065 DVDD.n4909 VSS 0.279212f
C22066 DVDD.n4910 VSS 0.279212f
C22067 DVDD.n4911 VSS 0.279212f
C22068 DVDD.n4912 VSS 0.279212f
C22069 DVDD.n4913 VSS 0.279212f
C22070 DVDD.n4914 VSS 0.279212f
C22071 DVDD.n4915 VSS 0.279212f
C22072 DVDD.n4916 VSS 0.279212f
C22073 DVDD.n4917 VSS 0.279212f
C22074 DVDD.n4918 VSS 0.279212f
C22075 DVDD.n4919 VSS 0.279212f
C22076 DVDD.n4920 VSS 0.279212f
C22077 DVDD.n4921 VSS 0.279212f
C22078 DVDD.n4922 VSS 0.279212f
C22079 DVDD.n4923 VSS 0.279212f
C22080 DVDD.n4924 VSS 0.279212f
C22081 DVDD.n4925 VSS 0.279212f
C22082 DVDD.n4926 VSS 0.279212f
C22083 DVDD.n4927 VSS 0.279212f
C22084 DVDD.n4928 VSS 0.279212f
C22085 DVDD.n4929 VSS 0.279212f
C22086 DVDD.n4930 VSS 0.279212f
C22087 DVDD.n4931 VSS 0.279212f
C22088 DVDD.n4932 VSS 0.279212f
C22089 DVDD.n4933 VSS 0.279212f
C22090 DVDD.n4934 VSS 0.279212f
C22091 DVDD.n4935 VSS 0.278229f
C22092 DVDD.n4936 VSS 0.279212f
C22093 DVDD.n4937 VSS 0.279212f
C22094 DVDD.n4938 VSS 0.139606f
C22095 DVDD.n4939 VSS 0.009915f
C22096 DVDD.n4940 VSS 0.009915f
C22097 DVDD.n4941 VSS 0.009915f
C22098 DVDD.n4942 VSS 0.009915f
C22099 DVDD.n4943 VSS 0.009915f
C22100 DVDD.n4944 VSS 0.009915f
C22101 DVDD.n4945 VSS 0.009915f
C22102 DVDD.n4946 VSS 0.009915f
C22103 DVDD.n4947 VSS 0.009915f
C22104 DVDD.n4948 VSS 0.009915f
C22105 DVDD.n4949 VSS 0.011355f
C22106 DVDD.n4950 VSS 0.011355f
C22107 DVDD.n4951 VSS 0.019831f
C22108 DVDD.n4952 VSS 0.019831f
C22109 DVDD.n4953 VSS 0.011115f
C22110 DVDD.n4954 VSS 0.010155f
C22111 DVDD.n4955 VSS 0.019831f
C22112 DVDD.n4956 VSS 0.011355f
C22113 DVDD.n4957 VSS 0.019831f
C22114 DVDD.n4958 VSS 0.011355f
C22115 DVDD.n4959 VSS 0.019831f
C22116 DVDD.n4960 VSS 0.011355f
C22117 DVDD.n4961 VSS 0.019831f
C22118 DVDD.n4962 VSS 0.011355f
C22119 DVDD.n4963 VSS 0.019831f
C22120 DVDD.n4964 VSS 0.011355f
C22121 DVDD.n4965 VSS 0.019831f
C22122 DVDD.n4966 VSS 0.011355f
C22123 DVDD.n4967 VSS 0.019831f
C22124 DVDD.n4968 VSS 0.019831f
C22125 DVDD.n4969 VSS 0.010955f
C22126 DVDD.n4970 VSS 0.010315f
C22127 DVDD.n4971 VSS 0.019831f
C22128 DVDD.n4972 VSS 0.011355f
C22129 DVDD.n4973 VSS 0.019831f
C22130 DVDD.n4974 VSS 0.011355f
C22131 DVDD.n4975 VSS 0.019831f
C22132 DVDD.n4976 VSS 0.011355f
C22133 DVDD.n4977 VSS 0.019831f
C22134 DVDD.n4978 VSS 0.011355f
C22135 DVDD.n4979 VSS 0.019831f
C22136 DVDD.n4980 VSS 0.011355f
C22137 DVDD.n4981 VSS 0.019831f
C22138 DVDD.n4982 VSS 0.011355f
C22139 DVDD.n4983 VSS 0.019831f
C22140 DVDD.n4984 VSS 0.019831f
C22141 DVDD.n4985 VSS 0.010795f
C22142 DVDD.n4986 VSS 0.010475f
C22143 DVDD.n4987 VSS 0.019831f
C22144 DVDD.n4988 VSS 0.011355f
C22145 DVDD.n4989 VSS 0.019831f
C22146 DVDD.n4990 VSS 0.019831f
C22147 DVDD.n4991 VSS 0.019831f
C22148 DVDD.n4992 VSS 0.011355f
C22149 DVDD.n4993 VSS 0.0615f
C22150 DVDD.n4994 VSS 0.011355f
C22151 DVDD.n4995 VSS 0.019831f
C22152 DVDD.n4996 VSS 0.019831f
C22153 DVDD.n4997 VSS 0.014873f
C22154 DVDD.n4998 VSS 0.019831f
C22155 DVDD.n4999 VSS 0.014953f
C22156 DVDD.n5000 VSS 0.019831f
C22157 DVDD.n5001 VSS 0.019831f
C22158 DVDD.n5002 VSS 0.011355f
C22159 DVDD.n5003 VSS 0.009915f
C22160 DVDD.n5004 VSS 0.139606f
C22161 DVDD.n5005 VSS 0.009915f
C22162 DVDD.n5006 VSS 0.015753f
C22163 DVDD.n5007 VSS 0.019831f
C22164 DVDD.n5008 VSS -0.292745f
C22165 DVDD.n5009 VSS -0.359726f
C22166 DVDD.n5010 VSS 0.011994f
C22167 DVDD.n5011 VSS 0.009915f
C22168 DVDD.n5012 VSS 0.139606f
C22169 DVDD.n5013 VSS 0.009915f
C22170 DVDD.n5014 VSS 0.018711f
C22171 DVDD.n5015 VSS 0.019831f
C22172 DVDD.n5016 VSS 0.019831f
C22173 DVDD.n5017 VSS 0.019831f
C22174 DVDD.n5018 VSS 0.013034f
C22175 DVDD.n5019 VSS 0.009915f
C22176 DVDD.n5020 VSS 0.139606f
C22177 DVDD.n5021 VSS 0.140589f
C22178 DVDD.n5022 VSS 0.279212f
C22179 DVDD.n5023 VSS 0.279212f
C22180 DVDD.n5024 VSS 0.279212f
C22181 DVDD.n5025 VSS 0.279212f
C22182 DVDD.n5026 VSS 0.279212f
C22183 DVDD.n5027 VSS 0.278229f
C22184 DVDD.n5028 VSS 0.279212f
C22185 DVDD.n5029 VSS 0.279212f
C22186 DVDD.n5030 VSS 0.279212f
C22187 DVDD.n5031 VSS 0.279212f
C22188 DVDD.n5032 VSS 0.279212f
C22189 DVDD.n5033 VSS 0.279212f
C22190 DVDD.n5034 VSS 0.279212f
C22191 DVDD.n5035 VSS 0.279212f
C22192 DVDD.n5036 VSS 0.279212f
C22193 DVDD.n5037 VSS 0.279212f
C22194 DVDD.n5038 VSS 0.279212f
C22195 DVDD.n5039 VSS 0.279212f
C22196 DVDD.n5040 VSS 0.279212f
C22197 DVDD.n5041 VSS 0.279212f
C22198 DVDD.n5042 VSS 0.279212f
C22199 DVDD.n5043 VSS 0.279212f
C22200 DVDD.n5044 VSS 0.279212f
C22201 DVDD.n5045 VSS 0.171067f
C22202 DVDD.n5046 VSS 0.171067f
C22203 DVDD.n5047 VSS 0.171067f
C22204 DVDD.n5048 VSS 0.336235f
C22205 DVDD.n5049 VSS 0.247752f
C22206 DVDD.n5050 VSS 0.279212f
C22207 DVDD.n5051 VSS 0.279212f
C22208 DVDD.n5052 VSS 0.279212f
C22209 DVDD.n5053 VSS 0.279212f
C22210 DVDD.n5054 VSS 0.279212f
C22211 DVDD.n5055 VSS 0.279212f
C22212 DVDD.n5056 VSS 0.279212f
C22213 DVDD.n5057 VSS 0.279212f
C22214 DVDD.n5058 VSS 0.279212f
C22215 DVDD.n5059 VSS 0.279212f
C22216 DVDD.n5060 VSS 0.279212f
C22217 DVDD.n5061 VSS 0.279212f
C22218 DVDD.n5062 VSS 0.279212f
C22219 DVDD.n5063 VSS 0.279212f
C22220 DVDD.n5064 VSS 0.279212f
C22221 DVDD.n5065 VSS 0.279212f
C22222 DVDD.n5066 VSS 0.279212f
C22223 DVDD.n5067 VSS 0.279212f
C22224 DVDD.n5068 VSS 0.266432f
C22225 DVDD.n5069 VSS 0.279212f
C22226 DVDD.n5070 VSS 0.279212f
C22227 DVDD.n5071 VSS 0.279212f
C22228 DVDD.n5072 VSS 0.279212f
C22229 DVDD.n5073 VSS 0.279212f
C22230 DVDD.n5074 VSS 0.279212f
C22231 DVDD.n5075 VSS 0.279212f
C22232 DVDD.n5076 VSS 0.279212f
C22233 DVDD.n5077 VSS 0.279212f
C22234 DVDD.n5078 VSS 0.279212f
C22235 DVDD.n5079 VSS 0.279212f
C22236 DVDD.n5080 VSS 0.279212f
C22237 DVDD.n5081 VSS 0.279212f
C22238 DVDD.n5082 VSS 0.215308f
C22239 DVDD.n5083 VSS 0.279212f
C22240 DVDD.n5084 VSS 0.247752f
C22241 DVDD.n5085 VSS 0.139606f
C22242 DVDD.n5086 VSS 0.009915f
C22243 DVDD.n5087 VSS 0.005821f
C22244 DVDD.n5088 VSS 0.019831f
C22245 DVDD.n5089 VSS 0.011355f
C22246 DVDD.n5090 VSS 0.019831f
C22247 DVDD.n5091 VSS 0.063326f
C22248 DVDD.n5092 VSS 0.011355f
C22249 DVDD.n5093 VSS 0.017212f
C22250 DVDD.n5094 VSS 0.108146f
C22251 DVDD.n5095 VSS 0.009915f
C22252 DVDD.n5096 VSS 0.013034f
C22253 DVDD.n5097 VSS 0.019831f
C22254 DVDD.n5098 VSS 0.019831f
C22255 DVDD.n5099 VSS 0.019831f
C22256 DVDD.n5100 VSS -0.292745f
C22257 DVDD.n5101 VSS 0.019831f
C22258 DVDD.n5102 VSS 0.009915f
C22259 DVDD.n5103 VSS 0.0615f
C22260 DVDD.n5104 VSS 0.139606f
C22261 DVDD.n5105 VSS 0.279212f
C22262 DVDD.n5106 VSS 0.247752f
C22263 DVDD.n5107 VSS 0.247752f
C22264 DVDD.n5108 VSS 0.279212f
C22265 DVDD.n5109 VSS 0.279212f
C22266 DVDD.n5110 VSS 0.279212f
C22267 DVDD.n5111 VSS 0.279212f
C22268 DVDD.n5112 VSS 0.279212f
C22269 DVDD.n5113 VSS 0.279212f
C22270 DVDD.n5114 VSS 0.279212f
C22271 DVDD.n5115 VSS 0.279212f
C22272 DVDD.n5116 VSS 0.279212f
C22273 DVDD.n5117 VSS 0.279212f
C22274 DVDD.n5118 VSS 0.279212f
C22275 DVDD.n5119 VSS 0.279212f
C22276 DVDD.n5120 VSS 0.279212f
C22277 DVDD.n5121 VSS 0.279212f
C22278 DVDD.n5122 VSS 0.279212f
C22279 DVDD.n5123 VSS 0.279212f
C22280 DVDD.n5124 VSS 0.279212f
C22281 DVDD.n5125 VSS 0.279212f
C22282 DVDD.n5126 VSS 0.279212f
C22283 DVDD.n5127 VSS 0.279212f
C22284 DVDD.n5128 VSS 0.279212f
C22285 DVDD.n5129 VSS 0.279212f
C22286 DVDD.n5130 VSS 0.279212f
C22287 DVDD.n5131 VSS 0.279212f
C22288 DVDD.n5132 VSS 0.279212f
C22289 DVDD.n5133 VSS 0.215308f
C22290 DVDD.n5134 VSS 0.139606f
C22291 DVDD.n5135 VSS 0.025087f
C22292 DVDD.n5136 VSS 0.005197f
C22293 DVDD.n5137 VSS 0.017764f
C22294 DVDD.n5138 VSS 0.011355f
C22295 DVDD.n5139 VSS 0.009915f
C22296 DVDD.n5140 VSS 0.011355f
C22297 DVDD.n5141 VSS 0.019831f
C22298 DVDD.n5142 VSS 0.019831f
C22299 DVDD.n5143 VSS 0.014873f
C22300 DVDD.n5144 VSS 0.019831f
C22301 DVDD.n5145 VSS 0.014953f
C22302 DVDD.n5146 VSS 0.019831f
C22303 DVDD.n5147 VSS 0.019831f
C22304 DVDD.n5148 VSS 0.019831f
C22305 DVDD.n5149 VSS 0.011355f
C22306 DVDD.n5150 VSS 0.019831f
C22307 DVDD.n5151 VSS 0.019831f
C22308 DVDD.n5152 VSS 0.010475f
C22309 DVDD.n5153 VSS 0.010795f
C22310 DVDD.n5154 VSS 0.019831f
C22311 DVDD.n5155 VSS 0.011355f
C22312 DVDD.n5156 VSS 0.019831f
C22313 DVDD.n5157 VSS 0.011355f
C22314 DVDD.n5158 VSS 0.019831f
C22315 DVDD.n5159 VSS 0.011355f
C22316 DVDD.n5160 VSS 0.019831f
C22317 DVDD.n5161 VSS 0.011355f
C22318 DVDD.n5162 VSS 0.019831f
C22319 DVDD.n5163 VSS 0.011355f
C22320 DVDD.n5164 VSS 0.019831f
C22321 DVDD.n5165 VSS 0.011355f
C22322 DVDD.n5166 VSS 0.019831f
C22323 DVDD.n5167 VSS 0.019831f
C22324 DVDD.n5168 VSS 0.010315f
C22325 DVDD.n5169 VSS 0.010955f
C22326 DVDD.n5170 VSS 0.019831f
C22327 DVDD.n5171 VSS 0.011355f
C22328 DVDD.n5172 VSS 0.019831f
C22329 DVDD.n5173 VSS 0.011355f
C22330 DVDD.n5174 VSS 0.019831f
C22331 DVDD.n5175 VSS 0.011355f
C22332 DVDD.n5176 VSS 0.019831f
C22333 DVDD.n5177 VSS 0.011355f
C22334 DVDD.n5178 VSS 0.019831f
C22335 DVDD.n5179 VSS 0.011355f
C22336 DVDD.n5180 VSS 0.019831f
C22337 DVDD.n5181 VSS 0.011355f
C22338 DVDD.n5182 VSS 0.019831f
C22339 DVDD.n5183 VSS 0.019831f
C22340 DVDD.n5184 VSS 0.010155f
C22341 DVDD.n5185 VSS 0.011115f
C22342 DVDD.n5186 VSS 0.019831f
C22343 DVDD.n5187 VSS 0.011355f
C22344 DVDD.n5188 VSS 0.019831f
C22345 DVDD.n5189 VSS 0.011355f
C22346 DVDD.n5190 VSS 0.019831f
C22347 DVDD.n5191 VSS 0.019831f
C22348 DVDD.n5192 VSS 0.015753f
C22349 DVDD.n5193 VSS 0.019831f
C22350 DVDD.n5194 VSS 0.011994f
C22351 DVDD.n5195 VSS -0.359726f
C22352 DVDD.n5196 VSS 0.011355f
C22353 DVDD.n5197 VSS 0.019831f
C22354 DVDD.n5198 VSS 0.011355f
C22355 DVDD.n5199 VSS 0.019831f
C22356 DVDD.n5200 VSS 0.011355f
C22357 DVDD.n5201 VSS 0.019831f
C22358 DVDD.n5202 VSS 0.011355f
C22359 DVDD.n5203 VSS 0.019831f
C22360 DVDD.n5204 VSS 0.011355f
C22361 DVDD.n5205 VSS 0.019831f
C22362 DVDD.n5206 VSS 0.019831f
C22363 DVDD.n5207 VSS 0.010555f
C22364 DVDD.n5208 VSS 0.010715f
C22365 DVDD.n5209 VSS 0.019831f
C22366 DVDD.n5210 VSS 0.011355f
C22367 DVDD.n5211 VSS 0.019831f
C22368 DVDD.n5212 VSS 0.011355f
C22369 DVDD.n5213 VSS 0.019831f
C22370 DVDD.n5214 VSS 0.011355f
C22371 DVDD.n5215 VSS 0.019831f
C22372 DVDD.n5216 VSS 0.011355f
C22373 DVDD.n5217 VSS 0.019831f
C22374 DVDD.n5218 VSS 0.011355f
C22375 DVDD.n5219 VSS 0.019831f
C22376 DVDD.n5220 VSS 0.011355f
C22377 DVDD.n5221 VSS 0.019831f
C22378 DVDD.n5222 VSS 0.019831f
C22379 DVDD.n5223 VSS 0.010395f
C22380 DVDD.n5224 VSS 0.010875f
C22381 DVDD.n5225 VSS 0.019831f
C22382 DVDD.n5226 VSS 0.011355f
C22383 DVDD.n5227 VSS 0.019831f
C22384 DVDD.n5228 VSS 0.011355f
C22385 DVDD.n5229 VSS 0.019831f
C22386 DVDD.n5230 VSS 0.011355f
C22387 DVDD.n5231 VSS 0.019831f
C22388 DVDD.n5232 VSS 0.011355f
C22389 DVDD.n5233 VSS 0.019831f
C22390 DVDD.n5234 VSS 0.011355f
C22391 DVDD.n5235 VSS 0.019831f
C22392 DVDD.n5236 VSS 0.011355f
C22393 DVDD.n5237 VSS 0.019831f
C22394 DVDD.n5238 VSS 0.019831f
C22395 DVDD.n5239 VSS 0.019831f
C22396 DVDD.n5240 VSS 0.011035f
C22397 DVDD.n5241 VSS 0.009915f
C22398 DVDD.n5242 VSS 0.139606f
C22399 DVDD.n5243 VSS 0.139606f
C22400 DVDD.n5244 VSS 0.247752f
C22401 DVDD.n5245 VSS 0.532863f
C22402 DVDD.n5246 VSS 0.532863f
C22403 DVDD.n5247 VSS 0.171067f
C22404 DVDD.n5248 VSS 0.171067f
C22405 DVDD.n5249 VSS 0.532863f
C22406 DVDD.n5250 VSS 0.247752f
C22407 DVDD.n5251 VSS 0.279212f
C22408 DVDD.n5252 VSS 0.279212f
C22409 DVDD.n5253 VSS 0.279212f
C22410 DVDD.n5254 VSS 0.279212f
C22411 DVDD.n5255 VSS 0.279212f
C22412 DVDD.n5256 VSS 0.279212f
C22413 DVDD.n5257 VSS 0.279212f
C22414 DVDD.n5258 VSS 0.279212f
C22415 DVDD.n5259 VSS 0.279212f
C22416 DVDD.n5260 VSS 0.279212f
C22417 DVDD.n5261 VSS 0.279212f
C22418 DVDD.n5262 VSS 0.279212f
C22419 DVDD.n5263 VSS 0.279212f
C22420 DVDD.n5264 VSS 0.279212f
C22421 DVDD.n5265 VSS 0.279212f
C22422 DVDD.n5266 VSS 0.279212f
C22423 DVDD.n5267 VSS 0.279212f
C22424 DVDD.n5268 VSS 0.279212f
C22425 DVDD.n5269 VSS 0.279212f
C22426 DVDD.n5270 VSS 0.279212f
C22427 DVDD.n5271 VSS 0.279212f
C22428 DVDD.n5272 VSS 0.279212f
C22429 DVDD.n5273 VSS 0.279212f
C22430 DVDD.n5274 VSS 0.279212f
C22431 DVDD.n5275 VSS 0.279212f
C22432 DVDD.n5276 VSS 0.279212f
C22433 DVDD.n5277 VSS 0.279212f
C22434 DVDD.n5278 VSS 0.279212f
C22435 DVDD.n5279 VSS 0.279212f
C22436 DVDD.n5280 VSS 0.279212f
C22437 DVDD.n5281 VSS 0.163202f
C22438 DVDD.n5282 VSS 0.163202f
C22439 DVDD.n5283 VSS 0.279212f
C22440 DVDD.n5284 VSS 0.279212f
C22441 DVDD.n5285 VSS 0.279212f
C22442 DVDD.n5286 VSS 0.279212f
C22443 DVDD.n5287 VSS 0.279212f
C22444 DVDD.n5288 VSS 0.279212f
C22445 DVDD.n5289 VSS 0.279212f
C22446 DVDD.n5290 VSS 0.279212f
C22447 DVDD.n5291 VSS 0.279212f
C22448 DVDD.n5292 VSS 0.279212f
C22449 DVDD.n5293 VSS 0.279212f
C22450 DVDD.n5294 VSS 0.279212f
C22451 DVDD.n5295 VSS 0.279212f
C22452 DVDD.n5296 VSS 0.279212f
C22453 DVDD.n5297 VSS 0.279212f
C22454 DVDD.n5298 VSS 0.279212f
C22455 DVDD.n5299 VSS 0.266432f
C22456 DVDD.n5300 VSS 0.279212f
C22457 DVDD.n5301 VSS 0.279212f
C22458 DVDD.n5302 VSS 0.279212f
C22459 DVDD.n5303 VSS 0.279212f
C22460 DVDD.n5304 VSS 0.279212f
C22461 DVDD.n5305 VSS 0.279212f
C22462 DVDD.n5306 VSS 0.279212f
C22463 DVDD.n5307 VSS 0.279212f
C22464 DVDD.n5308 VSS 0.279212f
C22465 DVDD.n5309 VSS 0.279212f
C22466 DVDD.n5310 VSS 0.279212f
C22467 DVDD.n5311 VSS 0.279212f
C22468 DVDD.n5312 VSS 0.279212f
C22469 DVDD.n5313 VSS 0.279212f
C22470 DVDD.n5314 VSS 0.279212f
C22471 DVDD.n5315 VSS 0.215308f
C22472 DVDD.n5316 VSS 0.139606f
C22473 DVDD.n5317 VSS 0.009915f
C22474 DVDD.n5318 VSS 0.108146f
C22475 DVDD.n5319 VSS 0.457161f
C22476 DVDD.n5320 VSS 0.260533f
C22477 DVDD.n5321 VSS 0.171067f
C22478 DVDD.n5322 VSS 0.171067f
C22479 DVDD.n5323 VSS 0.279212f
C22480 DVDD.n5324 VSS 0.279212f
C22481 DVDD.n5325 VSS 0.279212f
C22482 DVDD.n5326 VSS 0.279212f
C22483 DVDD.n5327 VSS 0.279212f
C22484 DVDD.n5328 VSS 0.279212f
C22485 DVDD.n5329 VSS 0.279212f
C22486 DVDD.n5330 VSS 0.279212f
C22487 DVDD.n5331 VSS 0.279212f
C22488 DVDD.n5332 VSS 0.279212f
C22489 DVDD.n5333 VSS 0.279212f
C22490 DVDD.n5334 VSS 0.279212f
C22491 DVDD.n5335 VSS 0.279212f
C22492 DVDD.n5336 VSS 0.279212f
C22493 DVDD.n5337 VSS 0.278229f
C22494 DVDD.n5338 VSS 0.139606f
C22495 DVDD.n5339 VSS 0.025087f
C22496 DVDD.n5340 VSS 0.139606f
C22497 DVDD.n5341 VSS 0.140589f
C22498 DVDD.n5342 VSS 0.279212f
C22499 DVDD.n5343 VSS 0.279212f
C22500 DVDD.n5344 VSS 0.279212f
C22501 DVDD.n5345 VSS 0.279212f
C22502 DVDD.n5346 VSS 0.279212f
C22503 DVDD.n5347 VSS 0.279212f
C22504 DVDD.n5348 VSS 0.279212f
C22505 DVDD.n5349 VSS 0.279212f
C22506 DVDD.n5350 VSS 0.279212f
C22507 DVDD.n5351 VSS 0.279212f
C22508 DVDD.n5352 VSS 0.279212f
C22509 DVDD.n5353 VSS 0.279212f
C22510 DVDD.n5354 VSS 0.279212f
C22511 DVDD.n5355 VSS 0.279212f
C22512 DVDD.n5356 VSS 0.279212f
C22513 DVDD.n5357 VSS 0.239887f
C22514 DVDD.n5358 VSS 0.201544f
C22515 DVDD.n5359 VSS 0.100281f
C22516 DVDD.n5360 VSS 0.025087f
C22517 DVDD.n5361 VSS 0.139606f
C22518 DVDD.n5362 VSS 0.217274f
C22519 DVDD.n5363 VSS 0.279212f
C22520 DVDD.n5364 VSS 0.279212f
C22521 DVDD.n5365 VSS 0.279212f
C22522 DVDD.n5366 VSS 0.279212f
C22523 DVDD.n5367 VSS 0.279212f
C22524 DVDD.n5368 VSS 0.279212f
C22525 DVDD.n5369 VSS 0.279212f
C22526 DVDD.n5370 VSS 0.279212f
C22527 DVDD.n5371 VSS 0.279212f
C22528 DVDD.n5372 VSS 0.279212f
C22529 DVDD.n5373 VSS 0.279212f
C22530 DVDD.n5374 VSS 0.279212f
C22531 DVDD.n5375 VSS 0.279212f
C22532 DVDD.n5376 VSS 0.279212f
C22533 DVDD.n5377 VSS 0.279212f
C22534 DVDD.n5378 VSS 0.264465f
C22535 DVDD.n5379 VSS 0.139606f
C22536 DVDD.n5380 VSS 0.025087f
C22537 DVDD.n5381 VSS 0.139606f
C22538 DVDD.n5382 VSS 0.154353f
C22539 DVDD.n5383 VSS 0.279212f
C22540 DVDD.n5384 VSS 0.279212f
C22541 DVDD.n5385 VSS 0.279212f
C22542 DVDD.n5386 VSS 0.279212f
C22543 DVDD.n5387 VSS 0.279212f
C22544 DVDD.n5388 VSS 0.279212f
C22545 DVDD.n5389 VSS 0.279212f
C22546 DVDD.n5390 VSS 0.279212f
C22547 DVDD.n5391 VSS 0.279212f
C22548 DVDD.n5392 VSS 0.279212f
C22549 DVDD.n5393 VSS 0.279212f
C22550 DVDD.n5394 VSS 0.279212f
C22551 DVDD.n5395 VSS 0.279212f
C22552 DVDD.n5396 VSS 0.279212f
C22553 DVDD.n5397 VSS 0.232022f
C22554 DVDD.n5398 VSS 0.232022f
C22555 DVDD.n5399 VSS 0.336235f
C22556 DVDD.n5400 VSS 0.095365f
C22557 DVDD.n5401 VSS 0.186797f
C22558 DVDD.n5402 VSS 0.139606f
C22559 DVDD.n5403 VSS 0.279212f
C22560 DVDD.n5404 VSS 0.279212f
C22561 DVDD.n5405 VSS 0.129775f
C22562 DVDD.n5406 VSS 0.015767f
C22563 DVDD.n5407 VSS 0.015767f
C22564 DVDD.n5408 VSS 0.015767f
C22565 DVDD.n5409 VSS 0.015767f
C22566 DVDD.n5410 VSS 0.015767f
C22567 DVDD.n5411 VSS 0.015767f
C22568 DVDD.n5412 VSS 0.015767f
C22569 DVDD.n5413 VSS 0.015767f
C22570 DVDD.n5414 VSS 0.015767f
C22571 DVDD.n5415 VSS 0.091432f
C22572 DVDD.n5416 VSS 0.015767f
C22573 DVDD.n5417 VSS 0.018056f
C22574 DVDD.n5418 VSS 3.85328f
C22575 DVDD.n5420 VSS 3.92842f
C22576 DVDD.n5421 VSS 0.015894f
C22577 DVDD.n5422 VSS 0.610461f
C22578 DVDD.n5423 VSS 0.147731f
C22579 DVDD.n5424 VSS 0.059812f
C22580 DVDD.n5425 VSS 0.027037f
C22581 DVDD.n5426 VSS 0.016565f
C22582 DVDD.n5427 VSS 0.090449f
C22583 DVDD.n5428 VSS 0.02361f
C22584 DVDD.n5429 VSS 0.029633f
C22585 DVDD.n5430 VSS 0.018391f
C22586 DVDD.n5431 VSS 0.070301f
C22587 DVDD.n5432 VSS 0.070301f
C22588 DVDD.n5433 VSS 0.070301f
C22589 DVDD.n5434 VSS 0.026085f
C22590 DVDD.n5435 VSS 0.070301f
C22591 DVDD.n5436 VSS 0.026085f
C22592 DVDD.n5437 VSS 0.070301f
C22593 DVDD.n5438 VSS 0.070301f
C22594 DVDD.n5439 VSS 0.023991f
C22595 DVDD.n5440 VSS 0.025704f
C22596 DVDD.n5441 VSS 0.070301f
C22597 DVDD.n5442 VSS 0.026085f
C22598 DVDD.n5443 VSS 0.070301f
C22599 DVDD.n5444 VSS 0.026085f
C22600 DVDD.n5445 VSS 0.070301f
C22601 DVDD.n5446 VSS 0.026085f
C22602 DVDD.n5447 VSS 0.070301f
C22603 DVDD.n5448 VSS 0.026085f
C22604 DVDD.n5449 VSS 0.070301f
C22605 DVDD.n5450 VSS 0.026085f
C22606 DVDD.n5451 VSS 0.070301f
C22607 DVDD.n5452 VSS 0.026085f
C22608 DVDD.n5453 VSS 0.070301f
C22609 DVDD.n5454 VSS 0.038552f
C22610 DVDD.n5455 VSS 0.035151f
C22611 DVDD.n5456 VSS 0.02361f
C22612 DVDD.n5457 VSS 0.0238f
C22613 DVDD.n5458 VSS 0.0669f
C22614 DVDD.n5459 VSS 0.026085f
C22615 DVDD.n5460 VSS 0.070301f
C22616 DVDD.n5461 VSS 0.026085f
C22617 DVDD.n5462 VSS 0.070301f
C22618 DVDD.n5463 VSS 0.026085f
C22619 DVDD.n5464 VSS 0.070301f
C22620 DVDD.n5465 VSS 0.026085f
C22621 DVDD.n5466 VSS 0.070301f
C22622 DVDD.n5467 VSS 0.026085f
C22623 DVDD.n5468 VSS 0.070301f
C22624 DVDD.n5469 VSS 0.070301f
C22625 DVDD.n5470 VSS 0.026085f
C22626 DVDD.n5471 VSS 0.023609f
C22627 DVDD.n5472 VSS 0.139606f
C22628 DVDD.n5473 VSS 0.012947f
C22629 DVDD.n5474 VSS 0.011614f
C22630 DVDD.n5475 VSS 0.139606f
C22631 DVDD.n5476 VSS 0.017326f
C22632 DVDD.n5477 VSS 0.026085f
C22633 DVDD.n5478 VSS 0.070301f
C22634 DVDD.n5479 VSS 0.070301f
C22635 DVDD.n5480 VSS 0.024965f
C22636 DVDD.n5481 VSS 0.018685f
C22637 DVDD.n5482 VSS 0.024511f
C22638 DVDD.n5483 VSS -0.253324f
C22639 DVDD.n5484 VSS 0.03515f
C22640 DVDD.n5485 VSS 5.34011f
C22641 DVDD.n5486 VSS 2.04978f
C22642 DVDD.n5487 VSS 2.66368f
C22643 DVDD.n5488 VSS 0.876068f
C22644 DVDD.n5489 VSS 0.525311f
C22645 DVDD.n5490 VSS 6.12618f
C22646 DVDD.t140 VSS 4.67431f
C22647 DVDD.t96 VSS 4.7717f
C22648 DVDD.n5491 VSS 6.12618f
C22649 DVDD.t148 VSS 4.75399f
C22650 DVDD.t157 VSS 4.69202f
C22651 DVDD.t160 VSS 3.90411f
C22652 DVDD.n5492 VSS 6.12618f
C22653 DVDD.n5493 VSS 1.01395f
C22654 DVDD.t31 VSS 4.75399f
C22655 DVDD.n5494 VSS 6.12618f
C22656 DVDD.t102 VSS 4.67431f
C22657 DVDD.t113 VSS 4.7717f
C22658 DVDD.n5495 VSS 6.12618f
C22659 DVDD.n5496 VSS 0.882423f
C22660 DVDD.n5497 VSS 1.01919f
C22661 DVDD.n5498 VSS 6.12618f
C22662 DVDD.t24 VSS 3.98379f
C22663 DVDD.n5499 VSS 0.929551f
C22664 DVDD.n5500 VSS 8.41752f
C22665 DVDD.n5501 VSS 0.070464f
C22666 DVDD.n5502 VSS 0.027036f
C22667 DVDD.n5503 VSS 0.049154f
C22668 DVDD.n5504 VSS 0.035231f
C22669 DVDD.n5505 VSS 0.027036f
C22670 DVDD.n5506 VSS 0.056541f
C22671 DVDD.n5507 VSS 0.027036f
C22672 DVDD.n5508 VSS 0.070464f
C22673 DVDD.n5509 VSS 0.070464f
C22674 DVDD.n5510 VSS 0.03134f
C22675 DVDD.n5511 VSS 0.019967f
C22676 DVDD.n5512 VSS 0.070464f
C22677 DVDD.n5513 VSS 0.070464f
C22678 DVDD.n5514 VSS 0.070464f
C22679 DVDD.n5515 VSS 0.024371f
C22680 DVDD.n5516 VSS 0.070464f
C22681 DVDD.n5517 VSS 0.027037f
C22682 DVDD.n5518 VSS 0.070464f
C22683 DVDD.n5519 VSS 0.027037f
C22684 DVDD.n5520 VSS 0.070464f
C22685 DVDD.n5521 VSS 0.027037f
C22686 DVDD.n5522 VSS 0.070464f
C22687 DVDD.n5523 VSS 0.027037f
C22688 DVDD.n5524 VSS 0.070464f
C22689 DVDD.n5525 VSS 0.027037f
C22690 DVDD.n5526 VSS 0.070464f
C22691 DVDD.n5527 VSS 0.027037f
C22692 DVDD.n5528 VSS 0.070464f
C22693 DVDD.n5529 VSS 0.070464f
C22694 DVDD.n5530 VSS 0.025895f
C22695 DVDD.n5531 VSS 0.024752f
C22696 DVDD.n5532 VSS 0.070464f
C22697 DVDD.n5533 VSS 0.027037f
C22698 DVDD.n5534 VSS 0.070464f
C22699 DVDD.n5535 VSS 0.027037f
C22700 DVDD.n5536 VSS 0.047165f
C22701 DVDD.n5537 VSS 0.035232f
C22702 DVDD.n5538 VSS 0.027037f
C22703 DVDD.n5539 VSS 0.05853f
C22704 DVDD.n5540 VSS 0.027037f
C22705 DVDD.n5541 VSS 0.070464f
C22706 DVDD.n5542 VSS 0.027037f
C22707 DVDD.n5543 VSS 0.070464f
C22708 DVDD.n5544 VSS 0.027037f
C22709 DVDD.n5545 VSS 0.070464f
C22710 DVDD.n5546 VSS 0.070464f
C22711 DVDD.n5547 VSS 0.025514f
C22712 DVDD.n5548 VSS 0.025133f
C22713 DVDD.n5549 VSS 0.070464f
C22714 DVDD.n5550 VSS 0.027037f
C22715 DVDD.n5551 VSS 0.070464f
C22716 DVDD.n5552 VSS 0.027037f
C22717 DVDD.n5553 VSS 0.070464f
C22718 DVDD.n5554 VSS 0.027037f
C22719 DVDD.n5555 VSS 0.070464f
C22720 DVDD.n5556 VSS 0.027037f
C22721 DVDD.n5557 VSS 0.070464f
C22722 DVDD.n5558 VSS 0.027037f
C22723 DVDD.n5559 VSS 0.065633f
C22724 DVDD.n5560 VSS -0.171072f
C22725 DVDD.n5561 VSS 0.013899f
C22726 DVDD.n5562 VSS 0.070464f
C22727 DVDD.n5563 VSS 0.139606f
C22728 DVDD.n5564 VSS 0.139606f
C22729 DVDD.n5565 VSS 0.026085f
C22730 DVDD.n5566 VSS 0.020753f
C22731 DVDD.n5567 VSS 0.003998f
C22732 DVDD.n5568 VSS 0.010853f
C22733 DVDD.n5569 VSS 0.017707f
C22734 DVDD.n5570 VSS 0.003237f
C22735 DVDD.n5571 VSS 0.007806f
C22736 DVDD.n5572 VSS 0.014661f
C22737 DVDD.n5573 VSS 0.021515f
C22738 DVDD.n5574 VSS 0.00476f
C22739 DVDD.n5575 VSS 0.279212f
C22740 DVDD.n5576 VSS 0.279212f
C22741 DVDD.n5577 VSS 0.279212f
C22742 DVDD.n5578 VSS 0.279212f
C22743 DVDD.n5579 VSS 0.279212f
C22744 DVDD.n5580 VSS 0.279212f
C22745 DVDD.n5581 VSS 0.279212f
C22746 DVDD.n5582 VSS 0.279212f
C22747 DVDD.n5583 VSS 0.279212f
C22748 DVDD.n5584 VSS 0.279212f
C22749 DVDD.n5585 VSS 0.279212f
C22750 DVDD.n5586 VSS 0.279212f
C22751 DVDD.n5587 VSS 0.251684f
C22752 DVDD.n5588 VSS 0.031461f
C22753 DVDD.n5589 VSS 0.396686f
C22754 DVDD.n5590 VSS 1.28646f
C22755 DVDD.n5591 VSS 0.251684f
C22756 DVDD.n5592 VSS 0.251684f
C22757 DVDD.n5593 VSS 0.279212f
C22758 DVDD.n5594 VSS 0.279212f
C22759 DVDD.n5595 VSS 0.279212f
C22760 DVDD.n5596 VSS 0.279212f
C22761 DVDD.n5597 VSS 0.279212f
C22762 DVDD.n5598 VSS 0.279212f
C22763 DVDD.n5599 VSS 0.279212f
C22764 DVDD.n5600 VSS 0.279212f
C22765 DVDD.n5601 VSS 0.196628f
C22766 DVDD.n5602 VSS 0.001332f
C22767 DVDD.n5603 VSS 0.018088f
C22768 DVDD.n5604 VSS 0.011233f
C22769 DVDD.n5605 VSS 0.004379f
C22770 DVDD.n5606 VSS 0.021134f
C22771 DVDD.n5607 VSS 0.01428f
C22772 DVDD.n5608 VSS 0.007425f
C22773 DVDD.n5609 VSS 0.026085f
C22774 DVDD.n5610 VSS 0.070464f
C22775 DVDD.n5611 VSS 0.026085f
C22776 DVDD.n5612 VSS 0.070464f
C22777 DVDD.n5613 VSS 0.070464f
C22778 DVDD.n5614 VSS 0.023991f
C22779 DVDD.n5615 VSS 0.025704f
C22780 DVDD.n5616 VSS 0.070464f
C22781 DVDD.n5617 VSS 0.026085f
C22782 DVDD.n5618 VSS 0.070464f
C22783 DVDD.n5619 VSS 0.026085f
C22784 DVDD.n5620 VSS 0.070464f
C22785 DVDD.n5621 VSS 0.026085f
C22786 DVDD.n5622 VSS 0.070464f
C22787 DVDD.n5623 VSS 0.026085f
C22788 DVDD.n5624 VSS 0.070464f
C22789 DVDD.n5625 VSS 0.026085f
C22790 DVDD.n5626 VSS 0.070464f
C22791 DVDD.n5627 VSS 0.026085f
C22792 DVDD.n5628 VSS 0.070464f
C22793 DVDD.n5629 VSS 0.038641f
C22794 DVDD.n5630 VSS 0.035232f
C22795 DVDD.n5631 VSS 0.02361f
C22796 DVDD.n5632 VSS 0.0238f
C22797 DVDD.n5633 VSS 0.067054f
C22798 DVDD.n5634 VSS 0.026085f
C22799 DVDD.n5635 VSS 0.070464f
C22800 DVDD.n5636 VSS 0.026085f
C22801 DVDD.n5637 VSS 0.070464f
C22802 DVDD.n5638 VSS 0.026085f
C22803 DVDD.n5639 VSS 0.070464f
C22804 DVDD.n5640 VSS 0.026085f
C22805 DVDD.n5641 VSS 0.070464f
C22806 DVDD.n5642 VSS 0.026085f
C22807 DVDD.n5643 VSS 0.070464f
C22808 DVDD.n5644 VSS 0.026085f
C22809 DVDD.n5645 VSS 0.070464f
C22810 DVDD.n5646 VSS 0.070464f
C22811 DVDD.n5647 VSS 9.52e-19
C22812 DVDD.n5648 VSS 0.02361f
C22813 DVDD.n5649 VSS 0.139606f
C22814 DVDD.n5650 VSS 0.017326f
C22815 DVDD.n5651 VSS 0.026085f
C22816 DVDD.n5652 VSS 0.070464f
C22817 DVDD.n5653 VSS 0.070464f
C22818 DVDD.n5654 VSS 0.024965f
C22819 DVDD.n5655 VSS 0.018685f
C22820 DVDD.n5656 VSS 0.024511f
C22821 DVDD.n5657 VSS -0.253232f
C22822 DVDD.n5658 VSS 0.035231f
C22823 DVDD.n5659 VSS 5.35569f
C22824 DVDD.n5660 VSS 2.05863f
C22825 DVDD.n5661 VSS 2.67254f
C22826 DVDD.n5662 VSS 0.877402f
C22827 DVDD.n5663 VSS 0.030356f
C22828 DVDD.n5664 VSS 0.018056f
C22829 DVDD.n5665 VSS 0.045533f
C22830 DVDD.n5666 VSS 0.018056f
C22831 DVDD.n5667 VSS 0.060711f
C22832 DVDD.n5668 VSS 0.018056f
C22833 DVDD.n5669 VSS 0.060711f
C22834 DVDD.n5670 VSS 0.060711f
C22835 DVDD.n5671 VSS 0.060711f
C22836 DVDD.n5672 VSS 0.015894f
C22837 DVDD.n5673 VSS 0.279212f
C22838 DVDD.n5674 VSS 0.279212f
C22839 DVDD.n5675 VSS 0.279212f
C22840 DVDD.n5676 VSS 0.279212f
C22841 DVDD.n5677 VSS 0.279212f
C22842 DVDD.n5678 VSS 0.279212f
C22843 DVDD.n5679 VSS 0.279212f
C22844 DVDD.n5680 VSS 0.279212f
C22845 DVDD.n5681 VSS 0.279212f
C22846 DVDD.n5682 VSS 0.279212f
C22847 DVDD.n5683 VSS 0.279212f
C22848 DVDD.n5684 VSS 0.251684f
C22849 DVDD.n5685 VSS 0.279212f
C22850 DVDD.n5686 VSS 0.143539f
C22851 DVDD.n5687 VSS 0.396686f
C22852 DVDD.n5688 VSS 1.28646f
C22853 DVDD.n5689 VSS 0.251684f
C22854 DVDD.n5690 VSS 0.279212f
C22855 DVDD.n5691 VSS 0.279212f
C22856 DVDD.n5692 VSS 0.279212f
C22857 DVDD.n5693 VSS 0.279212f
C22858 DVDD.n5694 VSS 0.279212f
C22859 DVDD.n5695 VSS 0.279212f
C22860 DVDD.n5696 VSS 0.279212f
C22861 DVDD.n5697 VSS 0.279212f
C22862 DVDD.n5698 VSS 0.279212f
C22863 DVDD.n5699 VSS 0.279212f
C22864 DVDD.n5700 VSS 0.279212f
C22865 DVDD.n5701 VSS 0.120926f
C22866 DVDD.n5702 VSS 0.089466f
C22867 DVDD.n5703 VSS 0.015767f
C22868 DVDD.n5704 VSS 0.057022f
C22869 DVDD.n5705 VSS 0.101264f
C22870 DVDD.n5706 VSS 0.064128f
C22871 DVDD.n5707 VSS 0.139606f
C22872 DVDD.n5708 VSS 0.166151f
C22873 DVDD.n5709 VSS 0.255617f
C22874 DVDD.n5710 VSS 0.336235f
C22875 DVDD.n5711 VSS 0.163202f
C22876 DVDD.n5712 VSS 0.163202f
C22877 DVDD.n5713 VSS 0.279212f
C22878 DVDD.n5714 VSS 0.279212f
C22879 DVDD.n5715 VSS 0.279212f
C22880 DVDD.n5716 VSS 0.279212f
C22881 DVDD.n5717 VSS 0.279212f
C22882 DVDD.n5718 VSS 0.279212f
C22883 DVDD.n5719 VSS 0.279212f
C22884 DVDD.n5720 VSS 0.279212f
C22885 DVDD.n5721 VSS 0.279212f
C22886 DVDD.n5722 VSS 0.279212f
C22887 DVDD.n5723 VSS 0.279212f
C22888 DVDD.n5724 VSS 0.279212f
C22889 DVDD.n5725 VSS 0.279212f
C22890 DVDD.n5726 VSS 0.279212f
C22891 DVDD.n5727 VSS 0.152387f
C22892 DVDD.n5728 VSS 0.009915f
C22893 DVDD.n5729 VSS 0.011355f
C22894 DVDD.n5730 VSS 0.063326f
C22895 DVDD.n5731 VSS 0.005821f
C22896 DVDD.n5732 VSS 0.027427f
C22897 DVDD.n5733 VSS 0.139606f
C22898 DVDD.n5734 VSS 0.009915f
C22899 DVDD.n5735 VSS 0.011355f
C22900 DVDD.n5736 VSS 0.019831f
C22901 DVDD.n5737 VSS 0.019831f
C22902 DVDD.n5738 VSS 0.013034f
C22903 DVDD.n5739 VSS 0.019831f
C22904 DVDD.n5740 VSS 0.018711f
C22905 DVDD.n5741 VSS 0.019831f
C22906 DVDD.n5742 VSS 0.019831f
C22907 DVDD.n5743 VSS 0.011035f
C22908 DVDD.n5744 VSS 0.010235f
C22909 DVDD.n5745 VSS 0.019831f
C22910 DVDD.n5746 VSS 0.011355f
C22911 DVDD.n5747 VSS 0.019831f
C22912 DVDD.n5748 VSS 0.011355f
C22913 DVDD.n5749 VSS 0.019831f
C22914 DVDD.n5750 VSS 0.011355f
C22915 DVDD.n5751 VSS 0.019831f
C22916 DVDD.n5752 VSS 0.011355f
C22917 DVDD.n5753 VSS 0.019831f
C22918 DVDD.n5754 VSS 0.011355f
C22919 DVDD.n5755 VSS 0.019831f
C22920 DVDD.n5756 VSS 0.011355f
C22921 DVDD.n5757 VSS 0.019831f
C22922 DVDD.n5758 VSS 0.019831f
C22923 DVDD.n5759 VSS 0.010875f
C22924 DVDD.n5760 VSS 0.010395f
C22925 DVDD.n5761 VSS 0.019831f
C22926 DVDD.n5762 VSS 0.011355f
C22927 DVDD.n5763 VSS 0.019831f
C22928 DVDD.n5764 VSS 0.011355f
C22929 DVDD.n5765 VSS 0.019831f
C22930 DVDD.n5766 VSS 0.011355f
C22931 DVDD.n5767 VSS 0.019831f
C22932 DVDD.n5768 VSS 0.011355f
C22933 DVDD.n5769 VSS 0.019831f
C22934 DVDD.n5770 VSS 0.011355f
C22935 DVDD.n5771 VSS 0.019831f
C22936 DVDD.n5772 VSS 0.019831f
C22937 DVDD.n5773 VSS 0.011355f
C22938 DVDD.n5774 VSS 0.019831f
C22939 DVDD.n5775 VSS 0.011355f
C22940 DVDD.n5776 VSS 0.019831f
C22941 DVDD.n5777 VSS 0.011355f
C22942 DVDD.n5778 VSS 0.019831f
C22943 DVDD.n5779 VSS 0.019831f
C22944 DVDD.n5780 VSS 0.019831f
C22945 DVDD.n5781 VSS 0.010715f
C22946 DVDD.n5782 VSS 0.009915f
C22947 DVDD.n5783 VSS 0.139606f
C22948 DVDD.n5784 VSS 0.009915f
C22949 DVDD.n5785 VSS 0.011355f
C22950 DVDD.n5786 VSS 0.019831f
C22951 DVDD.n5787 VSS -0.359726f
C22952 DVDD.n5788 VSS 0.011994f
C22953 DVDD.n5789 VSS 0.019831f
C22954 DVDD.n5790 VSS 0.015753f
C22955 DVDD.n5791 VSS 0.019831f
C22956 DVDD.n5792 VSS 0.019831f
C22957 DVDD.n5793 VSS 0.011355f
C22958 DVDD.n5794 VSS 0.019831f
C22959 DVDD.n5795 VSS 0.019831f
C22960 DVDD.n5796 VSS 0.010475f
C22961 DVDD.n5797 VSS 0.010795f
C22962 DVDD.n5798 VSS 0.019831f
C22963 DVDD.n5799 VSS 0.011355f
C22964 DVDD.n5800 VSS 0.019831f
C22965 DVDD.n5801 VSS 0.011355f
C22966 DVDD.n5802 VSS 0.019831f
C22967 DVDD.n5803 VSS 0.011355f
C22968 DVDD.n5804 VSS 0.019831f
C22969 DVDD.n5805 VSS 0.011355f
C22970 DVDD.n5806 VSS 0.019831f
C22971 DVDD.n5807 VSS 0.011355f
C22972 DVDD.n5808 VSS 0.019831f
C22973 DVDD.n5809 VSS 0.011355f
C22974 DVDD.n5810 VSS 0.019831f
C22975 DVDD.n5811 VSS 0.019831f
C22976 DVDD.n5812 VSS 0.010315f
C22977 DVDD.n5813 VSS 0.010955f
C22978 DVDD.n5814 VSS 0.019831f
C22979 DVDD.n5815 VSS 0.011355f
C22980 DVDD.n5816 VSS 0.019831f
C22981 DVDD.n5817 VSS 0.011355f
C22982 DVDD.n5818 VSS 0.019831f
C22983 DVDD.n5819 VSS 0.011355f
C22984 DVDD.n5820 VSS 0.019831f
C22985 DVDD.n5821 VSS 0.011355f
C22986 DVDD.n5822 VSS 0.019831f
C22987 DVDD.n5823 VSS 0.011355f
C22988 DVDD.n5824 VSS 0.019831f
C22989 DVDD.n5825 VSS 0.011355f
C22990 DVDD.n5826 VSS 0.019831f
C22991 DVDD.n5827 VSS 0.019831f
C22992 DVDD.n5828 VSS 0.010155f
C22993 DVDD.n5829 VSS 0.011115f
C22994 DVDD.n5830 VSS 0.019831f
C22995 DVDD.n5831 VSS 0.019831f
C22996 DVDD.n5832 VSS 0.011355f
C22997 DVDD.n5833 VSS 0.009915f
C22998 DVDD.n5834 VSS 0.139606f
C22999 DVDD.n5835 VSS 0.009915f
C23000 DVDD.n5836 VSS 0.011355f
C23001 DVDD.n5837 VSS 0.019831f
C23002 DVDD.n5838 VSS 0.019831f
C23003 DVDD.n5839 VSS 0.014953f
C23004 DVDD.n5840 VSS 0.019831f
C23005 DVDD.n5841 VSS 0.014873f
C23006 DVDD.n5842 VSS 0.019831f
C23007 DVDD.n5843 VSS 0.011355f
C23008 DVDD.n5844 VSS 0.019831f
C23009 DVDD.n5845 VSS 0.011355f
C23010 DVDD.n5846 VSS 0.0615f
C23011 DVDD.n5847 VSS 0.005197f
C23012 DVDD.n5848 VSS 0.025087f
C23013 DVDD.n5849 VSS 0.139606f
C23014 DVDD.n5850 VSS 0.266432f
C23015 DVDD.n5851 VSS 0.279212f
C23016 DVDD.n5852 VSS 0.279212f
C23017 DVDD.n5853 VSS 0.279212f
C23018 DVDD.n5854 VSS 0.279212f
C23019 DVDD.n5855 VSS 0.279212f
C23020 DVDD.n5856 VSS 0.152387f
C23021 DVDD.n5857 VSS 0.279212f
C23022 DVDD.n5858 VSS 0.279212f
C23023 DVDD.n5859 VSS 0.279212f
C23024 DVDD.n5860 VSS 0.279212f
C23025 DVDD.n5861 VSS 0.279212f
C23026 DVDD.n5862 VSS 0.279212f
C23027 DVDD.n5863 VSS 0.279212f
C23028 DVDD.n5864 VSS 0.279212f
C23029 DVDD.n5865 VSS 0.279212f
C23030 DVDD.n5866 VSS 0.279212f
C23031 DVDD.n5867 VSS 0.279212f
C23032 DVDD.n5868 VSS 0.279212f
C23033 DVDD.n5869 VSS 0.279212f
C23034 DVDD.n5870 VSS 0.279212f
C23035 DVDD.n5871 VSS 0.279212f
C23036 DVDD.n5872 VSS 0.279212f
C23037 DVDD.n5873 VSS 0.279212f
C23038 DVDD.n5874 VSS 0.163202f
C23039 DVDD.n5875 VSS 0.163202f
C23040 DVDD.n5876 VSS 0.163202f
C23041 DVDD.n5877 VSS 0.336235f
C23042 DVDD.n5878 VSS 0.255617f
C23043 DVDD.n5879 VSS 0.255617f
C23044 DVDD.n5880 VSS 0.279212f
C23045 DVDD.n5881 VSS 0.120926f
C23046 DVDD.n5882 VSS 0.279212f
C23047 DVDD.n5883 VSS 0.279212f
C23048 DVDD.n5884 VSS 0.279212f
C23049 DVDD.n5885 VSS 0.279212f
C23050 DVDD.n5886 VSS 0.279212f
C23051 DVDD.n5887 VSS 0.279212f
C23052 DVDD.n5888 VSS 0.279212f
C23053 DVDD.n5889 VSS 0.279212f
C23054 DVDD.n5890 VSS 0.279212f
C23055 DVDD.n5891 VSS 0.279212f
C23056 DVDD.n5892 VSS 0.279212f
C23057 DVDD.n5893 VSS 0.251684f
C23058 DVDD.n5894 VSS 0.031461f
C23059 DVDD.n5895 VSS 0.396686f
C23060 DVDD.n5896 VSS 1.28646f
C23061 DVDD.n5897 VSS 0.251684f
C23062 DVDD.n5898 VSS 0.251684f
C23063 DVDD.n5899 VSS 0.279212f
C23064 DVDD.n5900 VSS 0.279212f
C23065 DVDD.n5901 VSS 0.279212f
C23066 DVDD.n5902 VSS 0.279212f
C23067 DVDD.n5903 VSS 0.279212f
C23068 DVDD.n5904 VSS 0.279212f
C23069 DVDD.n5905 VSS 0.279212f
C23070 DVDD.n5906 VSS 0.279212f
C23071 DVDD.n5907 VSS 0.177949f
C23072 DVDD.n5908 VSS 0.015767f
C23073 DVDD.n5909 VSS 0.015767f
C23074 DVDD.n5910 VSS 0.015767f
C23075 DVDD.n5911 VSS 0.015767f
C23076 DVDD.n5912 VSS 0.057022f
C23077 DVDD.n5913 VSS 0.015767f
C23078 DVDD.n5914 VSS 0.020726f
C23079 DVDD.n5915 VSS 3.94756f
C23080 DVDD.n5916 VSS 0.015894f
C23081 DVDD.n5917 VSS 0.601272f
C23082 DVDD.n5918 VSS 0.147194f
C23083 DVDD.n5919 VSS 0.058624f
C23084 DVDD.n5920 VSS 0.139606f
C23085 DVDD.n5921 VSS 0.02361f
C23086 DVDD.n5922 VSS 0.027037f
C23087 DVDD.n5923 VSS 0.070464f
C23088 DVDD.n5924 VSS 0.070464f
C23089 DVDD.n5925 VSS 0.029633f
C23090 DVDD.n5926 VSS 0.018391f
C23091 DVDD.n5927 VSS 0.026039f
C23092 DVDD.n5928 VSS 0.070464f
C23093 DVDD.n5929 VSS 0.070464f
C23094 DVDD.n5930 VSS 0.026085f
C23095 DVDD.n5931 VSS 0.016374f
C23096 DVDD.n5932 VSS 0.139606f
C23097 DVDD.n5933 VSS 0.139606f
C23098 DVDD.n5934 VSS 0.279212f
C23099 DVDD.n5935 VSS 0.255617f
C23100 DVDD.n5936 VSS 0.166151f
C23101 DVDD.n5937 VSS 0.532863f
C23102 DVDD.n5938 VSS 0.532863f
C23103 DVDD.n5939 VSS 0.163202f
C23104 DVDD.n5940 VSS 0.163202f
C23105 DVDD.n5941 VSS 0.163202f
C23106 DVDD.n5942 VSS 0.532863f
C23107 DVDD.n5943 VSS 0.255617f
C23108 DVDD.n5944 VSS 0.279212f
C23109 DVDD.n5945 VSS 0.279212f
C23110 DVDD.n5946 VSS 0.279212f
C23111 DVDD.n5947 VSS 0.279212f
C23112 DVDD.n5948 VSS 0.17205f
C23113 DVDD.n5949 VSS 0.279212f
C23114 DVDD.n5950 VSS 0.279212f
C23115 DVDD.n5951 VSS 0.139606f
C23116 DVDD.n5952 VSS 0.139606f
C23117 DVDD.n5953 VSS 0.026094f
C23118 DVDD.n5954 VSS 0.139606f
C23119 DVDD.n5955 VSS 0.196628f
C23120 DVDD.n5956 VSS 0.279212f
C23121 DVDD.n5957 VSS 0.279212f
C23122 DVDD.n5958 VSS 0.279212f
C23123 DVDD.n5959 VSS 0.279212f
C23124 DVDD.n5960 VSS 0.279212f
C23125 DVDD.n5961 VSS 0.279212f
C23126 DVDD.n5962 VSS 0.279212f
C23127 DVDD.n5963 VSS 0.279212f
C23128 DVDD.n5964 VSS 0.279212f
C23129 DVDD.n5965 VSS 0.279212f
C23130 DVDD.n5966 VSS 0.279212f
C23131 DVDD.n5967 VSS 0.251684f
C23132 DVDD.n5968 VSS 0.279212f
C23133 DVDD.n5969 VSS 0.143539f
C23134 DVDD.n5970 VSS 0.396686f
C23135 DVDD.n5971 VSS 1.28646f
C23136 GF_NI_IN_C_BASE_0.comp018green_out_predrv_1.EN.t1 VSS 0.811404f
C23137 GF_NI_IN_C_BASE_0.comp018green_out_predrv_1.EN.t4 VSS 0.434237f
C23138 GF_NI_IN_C_BASE_0.comp018green_out_predrv_1.EN.n0 VSS 0.574127f
C23139 GF_NI_IN_C_BASE_0.comp018green_out_predrv_1.EN.t3 VSS 0.798807f
C23140 GF_NI_IN_C_BASE_0.comp018green_out_predrv_1.EN.t2 VSS 1.61653f
C23141 GF_NI_IN_C_BASE_0.comp018green_out_predrv_1.EN.t0 VSS 0.763937f
.ends

