* NGSPICE file created from gf180mcu_fd_io__bi_t_flat.ext - technology: gf180mcuD

.subckt gf180mcu_fd_io__bi_t_flat DVSS DVDD PAD SL A Y PDRV1 PDRV0 PD CS OE IE PU
+ VDD VSS
X0 GF_NI_BI_T_BASE_0.comp018green_sigbuf_1_0.pmos_6p0_CDNS_4066195314512_0.D SL VSS VSS nfet_06v0 ad=0.66p pd=3.88u as=0.66p ps=3.88u w=1.5u l=0.7u
D0 CS VDD diode_pd2nw_06v0 pj=4u area=1p
X1 DVSS GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.A GF_NI_BI_T_BASE_0.comp018green_out_predrv_2.pmos_6p0_CDNS_4066195314515_0.D DVSS nfet_06v0 ad=1.56p pd=6.52u as=2.64p ps=12.879999u w=6u l=0.7u
X2 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_cms_smt_0.pmos_6p0_CDNS_4066195314534_0.D GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_3.Z DVDD DVDD pfet_06v0 ad=0.39p pd=2.02u as=0.66p ps=3.88u w=1.5u l=0.7u
X3 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_logic_pupd_0.comp018green_std_nand2_1.nmos_6p0_CDNS_4066195314511_0.D GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_logic_pupd_0.comp018green_std_nand2_0.A GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_logic_pupd_0.PUB_OUT VSS nfet_06v0 ad=0.78p pd=3.52u as=1.32p ps=6.88u w=3u l=0.7u
X4 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_pupd_0.ppolyf_u_CDNS_4066195314533_3.MINUS GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_pupd_0.ppolyf_u_CDNS_4066195314533_0.MINUS DVDD ppolyf_u r_width=0.8u r_length=35.7u
X5 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_logic_pupd_0.PUB_OUT GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_logic_pupd_0.comp018green_std_nand2_0.A VDD VDD pfet_06v0 ad=0.78p pd=3.52u as=1.32p ps=6.88u w=3u l=0.7u
X6 DVSS GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.SL GF_NI_BI_T_BASE_0.ndrive_x_<0> DVDD pfet_06v0 ad=5.28p pd=24.88u as=3.12p ps=12.52u w=11.999999u l=0.7u
X7 DVDD GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_1.Z GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_1.ZB DVDD pfet_06v0 ad=1.32p pd=6.88u as=0.78p ps=3.52u w=3u l=0.7u
X8 GF_NI_BI_T_BASE_0.ndrive_x_<0> GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.SL DVSS DVDD pfet_06v0 ad=3.12p pd=12.52u as=3.12p ps=12.52u w=11.999999u l=0.7u
X9 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_1.ZB GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_1.Z DVDD DVDD pfet_06v0 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.7u
X10 GF_NI_BI_T_BASE_0.comp018green_esd_cdm_0.IP_IN PAD w_4468_53342# ppolyf_u r_width=2.5u r_length=2.8u
X11 PAD GF_NI_BI_T_BASE_0.pdrive_y_<0> DVDD DVDD pfet_06v0_dss d_sab=2.78u s_sab=0.28u ad=0.1112n pd=85.56u as=11.199999p ps=80.56u w=40u l=0.7u
X12 GF_NI_BI_T_BASE_0.pdrive_y_<1> DVDD GF_NI_BI_T_BASE_0.pdrive_x_<1> DVSS nfet_06v0 ad=0.528p pd=3.28u as=0.528p ps=3.28u w=1.2u l=0.7u
X13 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_cms_smt_0.nmos_6p0_CDNS_4066195314540_0.S GF_NI_BI_T_BASE_0.comp018green_esd_cdm_0.IP_IN GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_cms_smt_0.nmos_6p0_CDNS_4066195314537_0.D DVSS nfet_06v0 ad=0.689p pd=3.17u as=0.689p ps=3.17u w=2.65u l=0.7u
X14 DVSS DVSS GF_NI_BI_T_BASE_0.ndrive_x_<0> DVDD pfet_06v0 ad=0.528p pd=3.28u as=0.528p ps=3.28u w=1.2u l=0.7u
X15 PAD GF_NI_BI_T_BASE_0.ndrive_x_<1> DVSS DVSS nfet_06v0_dss d_sab=3.78u s_sab=0.28u ad=0.14364n pd=83.56u as=10.639999p ps=76.56u w=38u l=1.15u
X16 DVSS GF_NI_BI_T_BASE_0.comp018green_out_predrv_1.ENB GF_NI_BI_T_BASE_0.comp018green_out_predrv_1.pmos_6p0_CDNS_4066195314515_0.D DVSS nfet_06v0 ad=1.56p pd=6.52u as=1.56p ps=6.52u w=6u l=0.7u
X17 DVDD DVSS cap_nmos_06v0 c_width=5u c_length=1.5u
X18 GF_NI_BI_T_BASE_0.pdrive_x_<0> GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.SLB GF_NI_BI_T_BASE_0.pdrive_y_<0> DVSS nfet_06v0 ad=2.64p pd=12.879999u as=1.56p ps=6.52u w=6u l=0.7u
X19 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_cms_smt_0.nmos_6p0_CDNS_4066195314540_0.S GF_NI_BI_T_BASE_0.comp018green_esd_cdm_0.IP_IN GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_drv_0.A DVSS nfet_06v0 ad=1.32p pd=6.88u as=0.78p ps=3.52u w=3u l=0.7u
X20 PU GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_logic_pupd_0.comp018green_std_xor2_0.pmos_6p0_CDNS_4066195314512_2.D GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_logic_pupd_0.comp018green_std_nand2_0.A VSS nfet_06v0 ad=0.66p pd=3.88u as=0.66p ps=3.88u w=1.5u l=0.7u
X21 GF_NI_BI_T_BASE_0.comp018green_out_predrv_1.ENB GF_NI_BI_T_BASE_0.comp018green_out_predrv_1.EN DVDD DVDD pfet_06v0 ad=2.64p pd=12.879999u as=1.56p ps=6.52u w=6u l=0.7u
X22 VDD PU GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_logic_pupd_0.comp018green_std_xor2_0.pmos_6p0_CDNS_4066195314512_1.D VDD pfet_06v0 ad=1.32p pd=6.88u as=1.32p ps=6.88u w=3u l=0.7u
X23 GF_NI_BI_T_BASE_0.comp018green_esd_cdm_0.IP_IN PAD w_4468_53342# ppolyf_u r_width=2.5u r_length=2.8u
X24 DVSS GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_1.pmos_6p0_CDNS_4066195314512_0.D GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_1.Z DVSS nfet_06v0 ad=0.39p pd=2.02u as=0.39p ps=2.02u w=1.5u l=0.7u
X25 PAD GF_NI_BI_T_BASE_0.pdrive_x_<2> DVDD DVDD pfet_06v0_dss d_sab=2.78u s_sab=0.28u ad=0.1112n pd=85.56u as=11.199999p ps=80.56u w=40u l=0.7u
X26 GF_NI_BI_T_BASE_0.ndrive_x_<3> GF_NI_BI_T_BASE_0.comp018green_out_predrv_1.pmos_6p0_CDNS_4066195314515_0.S DVSS DVSS nfet_06v0 ad=1.56p pd=6.52u as=1.56p ps=6.52u w=6u l=0.7u
X27 DVSS GF_NI_BI_T_BASE_0.comp018green_out_predrv_3.pmos_6p0_CDNS_4066195314515_0.S DVDD DVDD pfet_06v0 ad=5.28p pd=24.88u as=3.12p ps=12.52u w=11.999999u l=0.7u
X28 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_drv_0.A GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_1.Z DVDD DVDD pfet_06v0 ad=0.88p pd=4.88u as=0.52p ps=2.52u w=2u l=0.7u
X29 Y GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_drv_0.Z VSS VSS nfet_06v0 ad=0.39p pd=2.02u as=0.39p ps=2.02u w=1.5u l=0.7u
D1 GF_NI_BI_T_BASE_0.comp018green_esd_cdm_0.IP_IN DVDD diode_pd2nw_06v0 pj=42u area=20p
X30 GF_NI_BI_T_BASE_0.comp018green_out_sigbuf_oe_0.nmos_6p0_CDNS_4066195314511_1.S PDRV0 VDD VDD pfet_06v0 ad=0.78p pd=3.52u as=1.32p ps=6.88u w=3u l=0.7u
X31 GF_NI_BI_T_BASE_0.comp018green_out_predrv_2.pmos_6p0_CDNS_4066195314515_0.S GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.A DVDD DVDD pfet_06v0 ad=5.28p pd=24.88u as=3.12p ps=12.52u w=11.999999u l=0.7u
X32 DVSS GF_NI_BI_T_BASE_0.comp018green_out_predrv_1.pmos_6p0_CDNS_4066195314515_0.D GF_NI_BI_T_BASE_0.pdrive_y_<3> DVSS nfet_06v0 ad=1.56p pd=6.52u as=1.56p ps=6.52u w=6u l=0.7u
X33 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_cms_smt_0.pmos_6p0_CDNS_4066195314538_0.S GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_cms_smt_0.pmos_6p0_CDNS_4066195314534_0.D DVSS DVDD pfet_06v0 ad=0.836p pd=4.68u as=0.494p ps=2.42u w=1.9u l=0.7u
X34 PAD GF_NI_BI_T_BASE_0.ndrive_x_<0> DVSS DVSS nfet_06v0_dss d_sab=3.78u s_sab=0.28u ad=0.14364n pd=83.56u as=10.639999p ps=76.56u w=38u l=1.15u
X35 DVSS GF_NI_BI_T_BASE_0.comp018green_out_predrv_1.pmos_6p0_CDNS_4066195314515_0.S DVSS DVSS nfet_06v0 ad=1.56p pd=6.52u as=0.266236n ps=1.1062m w=6u l=0.7u
X36 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_0.pmos_6p0_CDNS_4066195314512_0.D GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_logic_pupd_0.PDB_OUT VDD VDD pfet_06v0 ad=1.32p pd=6.88u as=1.32p ps=6.88u w=3u l=0.7u
X37 DVSS GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_cms_smt_0.pmos_6p0_CDNS_4066195314534_0.D GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_cms_smt_0.pmos_6p0_CDNS_4066195314538_0.S DVDD pfet_06v0 ad=0.494p pd=2.42u as=0.836p ps=4.68u w=1.9u l=0.7u
X38 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_pupd_0.ppolyf_u_CDNS_4066195314533_0.PLUS GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_pupd_0.ppolyf_u_CDNS_4066195314533_0.MINUS DVDD ppolyf_u r_width=0.8u r_length=35.7u
X39 GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.SLB GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.SL DVDD DVDD pfet_06v0 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.7u
X40 DVDD GF_NI_BI_T_BASE_0.comp018green_out_sigbuf_oe_1.EN GF_NI_BI_T_BASE_0.comp018green_out_predrv_2.pmos_6p0_CDNS_4066195314515_0.S DVDD pfet_06v0 ad=3.12p pd=12.52u as=3.12p ps=12.52u w=11.999999u l=0.7u
X41 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_3.Z GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_3.pmos_6p0_CDNS_4066195314512_0.D DVDD DVDD pfet_06v0 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.7u
X42 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_pupd_0.PD GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_0.Z DVDD DVDD pfet_06v0 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.7u
X43 DVSS GF_NI_BI_T_BASE_0.comp018green_out_predrv_2.pmos_6p0_CDNS_4066195314515_0.S DVSS DVSS nfet_06v0 ad=1.56p pd=6.52u as=0 ps=0 w=6u l=0.7u
X44 DVDD GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_3.Z GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_3.ZB DVDD pfet_06v0 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.7u
X45 DVDD GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_0.pmos_6p0_CDNS_4066195314512_0.D GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_0.Z DVDD pfet_06v0 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.7u
X46 PAD GF_NI_BI_T_BASE_0.pdrive_x_<3> DVDD DVDD pfet_06v0_dss d_sab=2.78u s_sab=0.28u ad=0.1112n pd=85.56u as=11.199999p ps=80.56u w=40u l=0.7u
X47 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_1.pmos_6p0_CDNS_4066195314512_0.D IE VSS VSS nfet_06v0 ad=0.66p pd=3.88u as=0.66p ps=3.88u w=1.5u l=0.7u
X48 VDD GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_drv_0.Z Y VDD pfet_06v0 ad=0.91p pd=4.02u as=0.91p ps=4.02u w=3.5u l=0.7u
X49 Y GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_drv_0.Z VDD VDD pfet_06v0 ad=0.91p pd=4.02u as=1.54p ps=7.88u w=3.5u l=0.7u
X50 DVDD DVSS cap_nmos_06v0 c_width=5u c_length=1.5u
X51 DVSS GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_2.pmos_6p0_CDNS_4066195314512_0.D GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_pupd_0.PU_B DVSS nfet_06v0 ad=0.66p pd=3.88u as=0.39p ps=2.02u w=1.5u l=0.7u
D2 DVSS GF_NI_BI_T_BASE_0.comp018green_esd_cdm_0.IP_IN diode_nd2ps_06v0 pj=42u area=20p
X52 GF_NI_BI_T_BASE_0.pdrive_y_<1> GF_NI_BI_T_BASE_0.comp018green_out_predrv_3.pmos_6p0_CDNS_4066195314515_0.D DVSS DVSS nfet_06v0 ad=1.56p pd=6.52u as=2.64p ps=12.879999u w=6u l=0.7u
X53 DVDD GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.pmos_6p0_CDNS_4066195314515_0.D GF_NI_BI_T_BASE_0.pdrive_x_<0> DVDD pfet_06v0 ad=5.28p pd=24.88u as=3.12p ps=12.52u w=11.999999u l=0.7u
X54 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_0.Z GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_0.pmos_6p0_CDNS_4066195314512_0.D DVSS DVSS nfet_06v0 ad=0.39p pd=2.02u as=0.66p ps=3.88u w=1.5u l=0.7u
X55 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_pupd_0.pmos_6p0_CDNS_4066195314512_0.D GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_pupd_0.PU_B DVDD DVDD pfet_06v0 ad=1.32p pd=6.88u as=1.32p ps=6.88u w=3u l=0.7u
X56 DVDD GF_NI_BI_T_BASE_0.comp018green_out_predrv_2.pmos_6p0_CDNS_4066195314515_0.D GF_NI_BI_T_BASE_0.pdrive_y_<2> DVDD pfet_06v0 ad=3.12p pd=12.52u as=3.12p ps=12.52u w=11.999999u l=0.7u
X57 DVSS GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_cms_smt_0.nmos_6p0_CDNS_4066195314535_0.D GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_cms_smt_0.nmos_6p0_CDNS_4066195314530_0.D DVSS nfet_06v0 ad=0.66p pd=3.88u as=0.66p ps=3.88u w=1.5u l=0.7u
X58 DVSS GF_NI_BI_T_BASE_0.comp018green_out_sigbuf_a_0.nmos_6p0_CDNS_4066195314511_3.S GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.A DVSS nfet_06v0 ad=0.78p pd=3.52u as=1.32p ps=6.88u w=3u l=0.7u
X59 DVSS GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.pmos_6p0_CDNS_4066195314515_0.D GF_NI_BI_T_BASE_0.pdrive_y_<0> DVSS nfet_06v0 ad=2.64p pd=12.879999u as=1.56p ps=6.52u w=6u l=0.7u
X60 GF_NI_BI_T_BASE_0.pdrive_y_<0> GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.pmos_6p0_CDNS_4066195314515_0.D DVSS DVSS nfet_06v0 ad=1.56p pd=6.52u as=1.56p ps=6.52u w=6u l=0.7u
X61 GF_NI_BI_T_BASE_0.comp018green_out_predrv_3.pmos_6p0_CDNS_4066195314515_0.S GF_NI_BI_T_BASE_0.comp018green_out_sigbuf_oe_1.EN DVDD DVDD pfet_06v0 ad=3.12p pd=12.52u as=3.12p ps=12.52u w=11.999999u l=0.7u
X62 DVDD GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_pupd_0.PU_B GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_2.ZB DVDD pfet_06v0 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.7u
X63 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_drv_0.A GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_3.Z GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_cms_smt_0.pmos_6p0_CDNS_4066195314534_0.D DVSS nfet_06v0 ad=0.66p pd=3.88u as=0.66p ps=3.88u w=1.5u l=0.7u
X64 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_pupd_0.ppolyf_u_CDNS_4066195314533_1.PLUS GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_pupd_0.ppolyf_u_CDNS_4066195314533_1.MINUS DVDD ppolyf_u r_width=0.8u r_length=35.7u
X65 GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.pmos_6p0_CDNS_4066195314515_0.S GF_NI_BI_T_BASE_0.comp018green_out_sigbuf_oe_0.EN GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.pmos_6p0_CDNS_4066195314515_0.D DVSS nfet_06v0 ad=2.64p pd=12.879999u as=1.56p ps=6.52u w=6u l=0.7u
X66 DVDD GF_NI_BI_T_BASE_0.comp018green_out_predrv_1.pmos_6p0_CDNS_4066195314515_0.S DVSS DVDD pfet_06v0 ad=3.12p pd=12.52u as=3.12p ps=12.52u w=11.999999u l=0.7u
X67 DVDD GF_NI_BI_T_BASE_0.comp018green_out_predrv_3.pmos_6p0_CDNS_4066195314515_0.D GF_NI_BI_T_BASE_0.pdrive_y_<1> DVDD pfet_06v0 ad=5.28p pd=24.88u as=3.12p ps=12.52u w=11.999999u l=0.7u
X68 VDD CS GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_3.pmos_6p0_CDNS_4066195314512_0.D VDD pfet_06v0 ad=1.32p pd=6.88u as=1.32p ps=6.88u w=3u l=0.7u
X69 DVSS GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_0.Z GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_pupd_0.PD DVSS nfet_06v0 ad=0.66p pd=3.88u as=0.39p ps=2.02u w=1.5u l=0.7u
X70 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_cms_smt_0.nmos_6p0_CDNS_4066195314540_0.S GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_cms_smt_0.nmos_6p0_CDNS_4066195314530_0.D DVDD DVSS nfet_06v0 ad=0.572p pd=3.48u as=0.572p ps=3.48u w=1.3u l=0.7u
X71 DVSS GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.SL GF_NI_BI_T_BASE_0.ndrive_x_<3> DVDD pfet_06v0 ad=3.12p pd=12.52u as=3.12p ps=12.52u w=11.999999u l=0.7u
D3 IE VDD diode_pd2nw_06v0 pj=4u area=1p
X72 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_2.ZB GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_pupd_0.PU_B DVDD DVDD pfet_06v0 ad=0.78p pd=3.52u as=1.32p ps=6.88u w=3u l=0.7u
X73 GF_NI_BI_T_BASE_0.comp018green_out_sigbuf_oe_2.nmos_6p0_CDNS_4066195314511_1.S OE GF_NI_BI_T_BASE_0.comp018green_out_sigbuf_oe_2.nmos_6p0_CDNS_4066195314511_0.S VSS nfet_06v0 ad=1.32p pd=6.88u as=0.78p ps=3.52u w=3u l=0.7u
X74 PAD GF_NI_BI_T_BASE_0.pdrive_y_<2> DVDD DVDD pfet_06v0_dss d_sab=2.78u s_sab=0.28u ad=0.1112n pd=85.56u as=11.199999p ps=80.56u w=40u l=0.7u
X75 GF_NI_BI_T_BASE_0.pdrive_x_<3> GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.SLB GF_NI_BI_T_BASE_0.pdrive_y_<3> DVSS nfet_06v0 ad=2.64p pd=12.879999u as=1.56p ps=6.52u w=6u l=0.7u
X76 DVDD DVSS cap_nmos_06v0 c_width=5u c_length=1.5u
X77 GF_NI_BI_T_BASE_0.ndrive_x_<3> DVSS DVSS DVDD pfet_06v0 ad=0.528p pd=3.28u as=0.528p ps=3.28u w=1.2u l=0.7u
X78 GF_NI_BI_T_BASE_0.pdrive_y_<3> GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.SLB GF_NI_BI_T_BASE_0.pdrive_x_<3> DVSS nfet_06v0 ad=1.56p pd=6.52u as=2.64p ps=12.879999u w=6u l=0.7u
X79 DVDD DVSS cap_nmos_06v0 c_width=5u c_length=1.5u
X80 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_cms_smt_0.nmos_6p0_CDNS_4066195314537_0.D GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_1.Z DVSS DVSS nfet_06v0 ad=1.408p pd=7.28u as=0.832p ps=3.72u w=3.2u l=0.7u
X81 GF_NI_BI_T_BASE_0.comp018green_out_sigbuf_oe_2.nmos_6p0_CDNS_4066195314511_0.S VDD VSS VSS nfet_06v0 ad=0.78p pd=3.52u as=1.32p ps=6.88u w=3u l=0.7u
X82 DVSS GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.SL GF_NI_BI_T_BASE_0.ndrive_x_<2> DVDD pfet_06v0 ad=5.28p pd=24.88u as=3.12p ps=12.52u w=11.999999u l=0.7u
X83 VDD PDRV1 GF_NI_BI_T_BASE_0.comp018green_out_sigbuf_oe_1.nmos_6p0_CDNS_4066195314511_1.S VDD pfet_06v0 ad=1.32p pd=6.88u as=0.78p ps=3.52u w=3u l=0.7u
X84 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_logic_pupd_0.comp018green_std_nand2_0.A GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_logic_pupd_0.comp018green_std_xor2_0.pmos_6p0_CDNS_4066195314512_2.D GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_logic_pupd_0.comp018green_std_xor2_0.pmos_6p0_CDNS_4066195314512_1.D VDD pfet_06v0 ad=1.32p pd=6.88u as=1.32p ps=6.88u w=3u l=0.7u
X85 DVSS GF_NI_BI_T_BASE_0.comp018green_out_sigbuf_oe_1.EN GF_NI_BI_T_BASE_0.comp018green_out_sigbuf_oe_1.ENB DVSS nfet_06v0 ad=0.78p pd=3.52u as=1.32p ps=6.88u w=3u l=0.7u
X86 GF_NI_BI_T_BASE_0.pdrive_y_<0> GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.pmos_6p0_CDNS_4066195314515_0.D DVDD DVDD pfet_06v0 ad=3.12p pd=12.52u as=5.28p ps=24.88u w=11.999999u l=0.7u
X87 GF_NI_BI_T_BASE_0.comp018green_out_sigbuf_oe_1.nmos_6p0_CDNS_4066195314511_1.S OE VDD VDD pfet_06v0 ad=0.78p pd=3.52u as=1.32p ps=6.88u w=3u l=0.7u
X88 VDD OE GF_NI_BI_T_BASE_0.comp018green_out_sigbuf_a_0.nmos_6p0_CDNS_4066195314511_1.D VDD pfet_06v0 ad=1.32p pd=6.88u as=0.78p ps=3.52u w=3u l=0.7u
X89 GF_NI_BI_T_BASE_0.comp018green_out_sigbuf_a_0.nmos_6p0_CDNS_4066195314511_1.D A VDD VDD pfet_06v0 ad=0.78p pd=3.52u as=1.32p ps=6.88u w=3u l=0.7u
X90 GF_NI_BI_T_BASE_0.pdrive_x_<0> DVDD GF_NI_BI_T_BASE_0.pdrive_y_<0> DVSS nfet_06v0 ad=0.528p pd=3.28u as=0.528p ps=3.28u w=1.2u l=0.7u
X91 DVDD DVSS cap_nmos_06v0 c_width=5u c_length=1.5u
X92 VSS PU GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_logic_pupd_0.comp018green_std_nand2_1.nmos_6p0_CDNS_4066195314511_0.D VSS nfet_06v0 ad=1.32p pd=6.88u as=0.78p ps=3.52u w=3u l=0.7u
X93 GF_NI_BI_T_BASE_0.comp018green_sigbuf_1_0.pmos_6p0_CDNS_4066195314512_0.D SL VDD VDD pfet_06v0 ad=1.32p pd=6.88u as=1.32p ps=6.88u w=3u l=0.7u
X94 DVSS DVSS PAD DVSS nfet_06v0_dss d_sab=0.28u s_sab=3.78u ad=10.639999p pd=76.56u as=0.14364n ps=83.56u w=38u l=1.15u
X95 VDD PU GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_logic_pupd_0.PUB_OUT VDD pfet_06v0 ad=1.32p pd=6.88u as=0.78p ps=3.52u w=3u l=0.7u
X96 DVSS GF_NI_BI_T_BASE_0.comp018green_out_predrv_3.pmos_6p0_CDNS_4066195314515_0.S DVSS DVSS nfet_06v0 ad=1.56p pd=6.52u as=0 ps=0 w=6u l=0.7u
X97 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_drv_0.Z GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_drv_0.nmos_6p0_CDNS_4066195314547_0.S VDD VDD pfet_06v0 ad=0.65p pd=3.02u as=1.1p ps=5.88u w=2.5u l=0.7u
X98 DVDD GF_NI_BI_T_BASE_0.pdrive_y_<3> PAD DVDD pfet_06v0_dss d_sab=0.28u s_sab=2.78u ad=11.199999p pd=80.56u as=0.1112n ps=85.56u w=40u l=0.7u
X99 DVDD GF_NI_BI_T_BASE_0.comp018green_out_predrv_1.pmos_6p0_CDNS_4066195314515_0.D GF_NI_BI_T_BASE_0.pdrive_x_<3> DVDD pfet_06v0 ad=3.12p pd=12.52u as=3.12p ps=12.52u w=11.999999u l=0.7u
X100 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_drv_0.nmos_6p0_CDNS_4066195314547_0.S GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_drv_0.A DVSS DVSS nfet_06v0 ad=1.76p pd=8.88u as=1.04p ps=4.52u w=4u l=0.7u
X101 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_pupd_0.ppolyf_u_CDNS_4066195314533_0.PLUS GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_pupd_0.ppolyf_u_CDNS_4066195314533_1.MINUS DVDD ppolyf_u r_width=0.8u r_length=35.7u
X102 DVSS GF_NI_BI_T_BASE_0.comp018green_out_sigbuf_oe_1.ENB GF_NI_BI_T_BASE_0.comp018green_out_predrv_3.pmos_6p0_CDNS_4066195314515_0.D DVSS nfet_06v0 ad=1.56p pd=6.52u as=1.56p ps=6.52u w=6u l=0.7u
X103 GF_NI_BI_T_BASE_0.comp018green_out_predrv_1.pmos_6p0_CDNS_4066195314515_0.D GF_NI_BI_T_BASE_0.comp018green_out_predrv_1.ENB GF_NI_BI_T_BASE_0.comp018green_out_predrv_1.pmos_6p0_CDNS_4066195314515_0.S DVDD pfet_06v0 ad=5.28p pd=24.88u as=3.12p ps=12.52u w=11.999999u l=0.7u
X104 GF_NI_BI_T_BASE_0.pdrive_y_<1> GF_NI_BI_T_BASE_0.comp018green_out_predrv_3.pmos_6p0_CDNS_4066195314515_0.D DVDD DVDD pfet_06v0 ad=3.12p pd=12.52u as=3.12p ps=12.52u w=11.999999u l=0.7u
X105 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_cms_smt_0.nmos_6p0_CDNS_4066195314540_0.S GF_NI_BI_T_BASE_0.comp018green_esd_cdm_0.IP_IN GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_cms_smt_0.nmos_6p0_CDNS_4066195314537_0.D DVSS nfet_06v0 ad=1.166p pd=6.18u as=0.689p ps=3.17u w=2.65u l=0.7u
X106 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_drv_0.A GF_NI_BI_T_BASE_0.comp018green_esd_cdm_0.IP_IN GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_cms_smt_0.nmos_6p0_CDNS_4066195314540_0.S DVSS nfet_06v0 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.7u
X107 GF_NI_BI_T_BASE_0.pdrive_x_<3> GF_NI_BI_T_BASE_0.comp018green_out_predrv_1.pmos_6p0_CDNS_4066195314515_0.D DVDD DVDD pfet_06v0 ad=3.12p pd=12.52u as=5.28p ps=24.88u w=11.999999u l=0.7u
X108 GF_NI_BI_T_BASE_0.comp018green_out_sigbuf_oe_0.nmos_6p0_CDNS_4066195314511_1.S OE GF_NI_BI_T_BASE_0.comp018green_out_sigbuf_oe_0.nmos_6p0_CDNS_4066195314511_0.S VSS nfet_06v0 ad=1.32p pd=6.88u as=0.78p ps=3.52u w=3u l=0.7u
X109 DVSS DVSS PAD DVSS nfet_06v0_dss d_sab=0.28u s_sab=3.78u ad=10.639999p pd=76.56u as=0.14364n ps=83.56u w=38u l=1.15u
X110 DVDD DVSS cap_nmos_06v0 c_width=5u c_length=1.5u
X111 DVSS GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_3.pmos_6p0_CDNS_4066195314512_0.D GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_3.Z DVSS nfet_06v0 ad=0.66p pd=3.88u as=0.39p ps=2.02u w=1.5u l=0.7u
X112 VDD GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_drv_0.nmos_6p0_CDNS_4066195314547_0.S GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_drv_0.Z VDD pfet_06v0 ad=1.1p pd=5.88u as=0.65p ps=3.02u w=2.5u l=0.7u
D4 VSS OE diode_pd2nw_06v0 pj=1.92u area=0.2304p
X113 GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.pmos_6p0_CDNS_4066195314515_0.S GF_NI_BI_T_BASE_0.comp018green_out_sigbuf_oe_0.ENB GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.pmos_6p0_CDNS_4066195314515_0.D DVDD pfet_06v0 ad=3.12p pd=12.52u as=5.28p ps=24.88u w=11.999999u l=0.7u
X114 DVSS GF_NI_BI_T_BASE_0.comp018green_out_predrv_2.pmos_6p0_CDNS_4066195314515_0.D GF_NI_BI_T_BASE_0.pdrive_y_<2> DVSS nfet_06v0 ad=2.64p pd=12.879999u as=1.56p ps=6.52u w=6u l=0.7u
X115 DVSS GF_NI_BI_T_BASE_0.comp018green_out_predrv_2.pmos_6p0_CDNS_4066195314515_0.S DVSS DVSS nfet_06v0 ad=1.56p pd=6.52u as=0 ps=0 w=6u l=0.7u
X116 DVDD GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_1.pmos_6p0_CDNS_4066195314512_0.D GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_1.Z DVDD pfet_06v0 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.7u
X117 GF_NI_BI_T_BASE_0.pdrive_y_<2> GF_NI_BI_T_BASE_0.comp018green_out_predrv_2.pmos_6p0_CDNS_4066195314515_0.D DVSS DVSS nfet_06v0 ad=1.56p pd=6.52u as=1.56p ps=6.52u w=6u l=0.7u
X118 GF_NI_BI_T_BASE_0.comp018green_out_predrv_2.pmos_6p0_CDNS_4066195314515_0.S GF_NI_BI_T_BASE_0.comp018green_out_sigbuf_oe_1.EN GF_NI_BI_T_BASE_0.comp018green_out_predrv_2.pmos_6p0_CDNS_4066195314515_0.D DVSS nfet_06v0 ad=2.64p pd=12.879999u as=1.56p ps=6.52u w=6u l=0.7u
X119 DVDD GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_3.Z GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_cms_smt_0.pmos_6p0_CDNS_4066195314534_0.D DVDD pfet_06v0 ad=0.66p pd=3.88u as=0.39p ps=2.02u w=1.5u l=0.7u
X120 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_cms_smt_0.nmos_6p0_CDNS_4066195314530_0.D GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_cms_smt_0.nmos_6p0_CDNS_4066195314535_0.D GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_drv_0.A DVDD pfet_06v0 ad=0.88p pd=4.88u as=0.88p ps=4.88u w=2u l=0.7u
X121 DVSS GF_NI_BI_T_BASE_0.comp018green_sigbuf_1_0.pmos_6p0_CDNS_4066195314512_0.D GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.SL DVSS nfet_06v0 ad=0.39p pd=2.02u as=0.39p ps=2.02u w=1.5u l=0.7u
X122 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_cms_smt_0.nmos_6p0_CDNS_4066195314537_0.D GF_NI_BI_T_BASE_0.comp018green_esd_cdm_0.IP_IN GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_cms_smt_0.nmos_6p0_CDNS_4066195314540_0.S DVSS nfet_06v0 ad=0.689p pd=3.17u as=1.166p ps=6.18u w=2.65u l=0.7u
X123 VDD GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_drv_0.Z Y VDD pfet_06v0 ad=0.91p pd=4.02u as=0.91p ps=4.02u w=3.5u l=0.7u
X124 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_pupd_0.ppolyf_u_CDNS_4066195314533_1.PLUS GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_pupd_0.ppolyf_u_CDNS_4066195314533_2.PLUS DVDD ppolyf_u r_width=0.8u r_length=35.7u
X125 VSS PU GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_logic_pupd_0.comp018green_std_xor2_0.pmos_6p0_CDNS_4066195314512_1.D VSS nfet_06v0 ad=0.66p pd=3.88u as=0.66p ps=3.88u w=1.5u l=0.7u
X126 DVSS GF_NI_BI_T_BASE_0.comp018green_out_sigbuf_oe_2.nmos_6p0_CDNS_4066195314511_1.S GF_NI_BI_T_BASE_0.comp018green_out_predrv_1.EN DVSS nfet_06v0 ad=0.78p pd=3.52u as=1.32p ps=6.88u w=3u l=0.7u
X127 GF_NI_BI_T_BASE_0.pdrive_y_<0> GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.SLB GF_NI_BI_T_BASE_0.pdrive_x_<0> DVSS nfet_06v0 ad=1.56p pd=6.52u as=2.64p ps=12.879999u w=6u l=0.7u
X128 DVDD GF_NI_BI_T_BASE_0.pdrive_x_<1> PAD DVDD pfet_06v0_dss d_sab=0.28u s_sab=2.78u ad=11.199999p pd=80.56u as=0.1112n ps=85.56u w=40u l=0.7u
X129 GF_NI_BI_T_BASE_0.ndrive_x_<1> GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.SL DVSS DVDD pfet_06v0 ad=3.12p pd=12.52u as=5.28p ps=24.88u w=11.999999u l=0.7u
X130 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_3.ZB GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_3.Z DVSS DVSS nfet_06v0 ad=0.39p pd=2.02u as=0.66p ps=3.88u w=1.5u l=0.7u
X131 VSS GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_drv_0.Z Y VSS nfet_06v0 ad=0.39p pd=2.02u as=0.39p ps=2.02u w=1.5u l=0.7u
X132 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_pupd_0.PU_B GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_2.pmos_6p0_CDNS_4066195314512_0.D DVSS DVSS nfet_06v0 ad=0.39p pd=2.02u as=0.39p ps=2.02u w=1.5u l=0.7u
X133 Y GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_drv_0.Z VSS VSS nfet_06v0 ad=0.39p pd=2.02u as=0.66p ps=3.88u w=1.5u l=0.7u
X134 DVDD GF_NI_BI_T_BASE_0.comp018green_out_sigbuf_a_0.nmos_6p0_CDNS_4066195314511_3.S GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.A DVDD pfet_06v0 ad=1.56p pd=6.52u as=2.64p ps=12.879999u w=6u l=0.7u
X135 GF_NI_BI_T_BASE_0.comp018green_out_predrv_1.pmos_6p0_CDNS_4066195314515_0.D GF_NI_BI_T_BASE_0.comp018green_out_predrv_1.EN GF_NI_BI_T_BASE_0.comp018green_out_predrv_1.pmos_6p0_CDNS_4066195314515_0.S DVSS nfet_06v0 ad=1.56p pd=6.52u as=2.64p ps=12.879999u w=6u l=0.7u
X136 GF_NI_BI_T_BASE_0.comp018green_out_predrv_3.pmos_6p0_CDNS_4066195314515_0.D GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.A DVSS DVSS nfet_06v0 ad=2.64p pd=12.879999u as=1.56p ps=6.52u w=6u l=0.7u
X137 GF_NI_BI_T_BASE_0.pdrive_y_<3> DVDD GF_NI_BI_T_BASE_0.pdrive_x_<3> DVSS nfet_06v0 ad=0.528p pd=3.28u as=0.528p ps=3.28u w=1.2u l=0.7u
X138 DVSS GF_NI_BI_T_BASE_0.comp018green_out_predrv_3.pmos_6p0_CDNS_4066195314515_0.D GF_NI_BI_T_BASE_0.pdrive_y_<1> DVSS nfet_06v0 ad=1.56p pd=6.52u as=1.56p ps=6.52u w=6u l=0.7u
X139 GF_NI_BI_T_BASE_0.pdrive_y_<2> GF_NI_BI_T_BASE_0.comp018green_out_predrv_2.pmos_6p0_CDNS_4066195314515_0.D DVDD DVDD pfet_06v0 ad=3.12p pd=12.52u as=5.28p ps=24.88u w=11.999999u l=0.7u
X140 DVDD DVSS cap_nmos_06v0 c_width=3u c_length=3u
X141 DVSS GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.SL GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.SLB DVSS nfet_06v0 ad=0.66p pd=3.88u as=0.39p ps=2.02u w=1.5u l=0.7u
X142 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_1.Z GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_1.pmos_6p0_CDNS_4066195314512_0.D DVSS DVSS nfet_06v0 ad=0.39p pd=2.02u as=0.66p ps=3.88u w=1.5u l=0.7u
X143 VDD GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_drv_0.Z Y VDD pfet_06v0 ad=1.54p pd=7.88u as=0.91p ps=4.02u w=3.5u l=0.7u
X144 PAD GF_NI_BI_T_BASE_0.ndrive_x_<2> DVSS DVSS nfet_06v0_dss d_sab=3.78u s_sab=0.28u ad=0.14364n pd=83.56u as=10.639999p ps=76.56u w=38u l=1.15u
X145 GF_NI_BI_T_BASE_0.pdrive_x_<2> GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.SLB GF_NI_BI_T_BASE_0.pdrive_y_<2> DVSS nfet_06v0 ad=2.64p pd=12.879999u as=1.56p ps=6.52u w=6u l=0.7u
X146 DVDD GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_2.pmos_6p0_CDNS_4066195314512_0.D GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_pupd_0.PU_B DVDD pfet_06v0 ad=1.32p pd=6.88u as=0.78p ps=3.52u w=3u l=0.7u
X147 DVDD GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_1.Z GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_drv_0.A DVDD pfet_06v0 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=0.7u
X148 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_cms_smt_0.pmos_6p0_CDNS_4066195314538_0.S GF_NI_BI_T_BASE_0.comp018green_esd_cdm_0.IP_IN GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_drv_0.A DVDD pfet_06v0 ad=0.946p pd=5.18u as=0.559p ps=2.67u w=2.15u l=0.7u
X149 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_0.Z GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_0.pmos_6p0_CDNS_4066195314512_0.D DVDD DVDD pfet_06v0 ad=0.78p pd=3.52u as=1.32p ps=6.88u w=3u l=0.7u
D5 VSS VDD diode_pd2nw_06v0 pj=1.92u area=0.2304p
X150 GF_NI_BI_T_BASE_0.ndrive_x_<2> GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.SL DVSS DVDD pfet_06v0 ad=3.12p pd=12.52u as=3.12p ps=12.52u w=11.999999u l=0.7u
X151 VSS GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_logic_pupd_0.PUB_OUT GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_2.pmos_6p0_CDNS_4066195314512_0.D VSS nfet_06v0 ad=0.66p pd=3.88u as=0.66p ps=3.88u w=1.5u l=0.7u
D6 VSS OE diode_pd2nw_06v0 pj=1.92u area=0.2304p
X152 DVDD GF_NI_BI_T_BASE_0.comp018green_out_sigbuf_oe_1.EN GF_NI_BI_T_BASE_0.comp018green_out_sigbuf_oe_1.ENB DVDD pfet_06v0 ad=1.56p pd=6.52u as=2.64p ps=12.879999u w=6u l=0.7u
X153 DVSS DVSS GF_NI_BI_T_BASE_0.ndrive_x_<2> DVDD pfet_06v0 ad=0.528p pd=3.28u as=0.528p ps=3.28u w=1.2u l=0.7u
X154 GF_NI_BI_T_BASE_0.comp018green_esd_cdm_0.IP_IN GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_pupd_0.ppolyf_u_CDNS_4066195314533_2.PLUS DVDD ppolyf_u r_width=0.8u r_length=22.999998u
X155 DVDD GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_0.Z GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_pupd_0.PD DVDD pfet_06v0 ad=1.32p pd=6.88u as=0.78p ps=3.52u w=3u l=0.7u
X156 GF_NI_BI_T_BASE_0.pdrive_x_<0> GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.pmos_6p0_CDNS_4066195314515_0.D DVDD DVDD pfet_06v0 ad=3.12p pd=12.52u as=3.12p ps=12.52u w=11.999999u l=0.7u
X157 GF_NI_BI_T_BASE_0.comp018green_out_sigbuf_oe_0.ENB GF_NI_BI_T_BASE_0.comp018green_out_sigbuf_oe_0.EN DVSS DVSS nfet_06v0 ad=1.32p pd=6.88u as=0.78p ps=3.52u w=3u l=0.7u
X158 GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.SL GF_NI_BI_T_BASE_0.comp018green_sigbuf_1_0.pmos_6p0_CDNS_4066195314512_0.D DVSS DVSS nfet_06v0 ad=0.39p pd=2.02u as=0.66p ps=3.88u w=1.5u l=0.7u
X159 DVSS GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.pmos_6p0_CDNS_4066195314515_0.S GF_NI_BI_T_BASE_0.ndrive_x_<0> DVSS nfet_06v0 ad=1.56p pd=6.52u as=1.56p ps=6.52u w=6u l=0.7u
X160 Y GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_drv_0.Z VDD VDD pfet_06v0 ad=0.91p pd=4.02u as=0.91p ps=4.02u w=3.5u l=0.7u
X161 DVDD DVSS cap_nmos_06v0 c_width=3u c_length=3u
X162 DVDD GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.A GF_NI_BI_T_BASE_0.comp018green_out_predrv_3.pmos_6p0_CDNS_4066195314515_0.S DVDD pfet_06v0 ad=3.12p pd=12.52u as=5.28p ps=24.88u w=11.999999u l=0.7u
X163 DVSS GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_1.Z GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_cms_smt_0.nmos_6p0_CDNS_4066195314537_0.D DVSS nfet_06v0 ad=0.832p pd=3.72u as=0.832p ps=3.72u w=3.2u l=0.7u
X164 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_logic_pupd_0.comp018green_std_xor2_0.pmos_6p0_CDNS_4066195314512_2.D PD VDD VDD pfet_06v0 ad=1.32p pd=6.88u as=1.32p ps=6.88u w=3u l=0.7u
X165 GF_NI_BI_T_BASE_0.pdrive_y_<3> GF_NI_BI_T_BASE_0.comp018green_out_predrv_1.pmos_6p0_CDNS_4066195314515_0.D DVSS DVSS nfet_06v0 ad=1.56p pd=6.52u as=2.64p ps=12.879999u w=6u l=0.7u
D7 A VDD diode_pd2nw_06v0 pj=4u area=1p
X166 GF_NI_BI_T_BASE_0.pdrive_x_<1> GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.SLB GF_NI_BI_T_BASE_0.pdrive_y_<1> DVSS nfet_06v0 ad=2.64p pd=12.879999u as=1.56p ps=6.52u w=6u l=0.7u
X167 DVDD GF_NI_BI_T_BASE_0.comp018green_out_predrv_2.pmos_6p0_CDNS_4066195314515_0.D GF_NI_BI_T_BASE_0.pdrive_x_<2> DVDD pfet_06v0 ad=5.28p pd=24.88u as=3.12p ps=12.52u w=11.999999u l=0.7u
X168 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_cms_smt_0.nmos_6p0_CDNS_4066195314537_0.D GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_1.Z DVSS DVSS nfet_06v0 ad=0.832p pd=3.72u as=1.408p ps=7.28u w=3.2u l=0.7u
X169 GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.pmos_6p0_CDNS_4066195314515_0.D GF_NI_BI_T_BASE_0.comp018green_out_sigbuf_oe_0.ENB DVSS DVSS nfet_06v0 ad=1.56p pd=6.52u as=1.56p ps=6.52u w=6u l=0.7u
X170 DVDD GF_NI_BI_T_BASE_0.pdrive_x_<0> PAD DVDD pfet_06v0_dss d_sab=0.28u s_sab=2.78u ad=11.199999p pd=80.56u as=0.1112n ps=85.56u w=40u l=0.7u
X171 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_1.pmos_6p0_CDNS_4066195314512_0.D IE VDD VDD pfet_06v0 ad=1.32p pd=6.88u as=1.32p ps=6.88u w=3u l=0.7u
X172 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_pupd_0.pmos_6p0_CDNS_4066195314512_0.D GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_pupd_0.ppolyf_u_CDNS_4066195314533_4.PLUS DVDD ppolyf_u r_width=0.8u r_length=35.7u
X173 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_logic_pupd_0.comp018green_std_nand2_0.A PD GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_logic_pupd_0.comp018green_std_xor2_0.pmos_6p0_CDNS_4066195314512_1.D VSS nfet_06v0 ad=0.66p pd=3.88u as=0.66p ps=3.88u w=1.5u l=0.7u
X174 GF_NI_BI_T_BASE_0.comp018green_out_predrv_1.pmos_6p0_CDNS_4066195314515_0.S GF_NI_BI_T_BASE_0.comp018green_out_predrv_1.EN DVDD DVDD pfet_06v0 ad=3.12p pd=12.52u as=3.12p ps=12.52u w=11.999999u l=0.7u
X175 DVDD GF_NI_BI_T_BASE_0.comp018green_out_predrv_1.pmos_6p0_CDNS_4066195314515_0.D GF_NI_BI_T_BASE_0.pdrive_y_<3> DVDD pfet_06v0 ad=5.28p pd=24.88u as=3.12p ps=12.52u w=11.999999u l=0.7u
X176 VDD OE GF_NI_BI_T_BASE_0.comp018green_out_sigbuf_oe_2.nmos_6p0_CDNS_4066195314511_1.S VDD pfet_06v0 ad=1.32p pd=6.88u as=0.78p ps=3.52u w=3u l=0.7u
X177 PAD GF_NI_BI_T_BASE_0.pdrive_x_<1> DVDD DVDD pfet_06v0_dss d_sab=2.78u s_sab=0.28u ad=0.1112n pd=85.56u as=11.199999p ps=80.56u w=40u l=0.7u
X178 GF_NI_BI_T_BASE_0.comp018green_out_sigbuf_oe_2.nmos_6p0_CDNS_4066195314511_1.S VDD VDD VDD pfet_06v0 ad=0.78p pd=3.52u as=1.32p ps=6.88u w=3u l=0.7u
X179 DVSS GF_NI_BI_T_BASE_0.comp018green_out_predrv_1.pmos_6p0_CDNS_4066195314515_0.S GF_NI_BI_T_BASE_0.ndrive_x_<3> DVSS nfet_06v0 ad=2.64p pd=12.879999u as=1.56p ps=6.52u w=6u l=0.7u
X180 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_cms_smt_0.nmos_6p0_CDNS_4066195314535_0.D GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_3.Z DVSS DVSS nfet_06v0 ad=0.52p pd=2.52u as=0.88p ps=4.88u w=2u l=0.7u
X181 DVSS DVSS PAD DVSS nfet_06v0_dss d_sab=0.28u s_sab=3.78u ad=10.639999p pd=76.56u as=0.14364n ps=83.56u w=38u l=1.15u
X182 GF_NI_BI_T_BASE_0.comp018green_out_sigbuf_oe_1.EN GF_NI_BI_T_BASE_0.comp018green_out_sigbuf_oe_1.nmos_6p0_CDNS_4066195314511_1.S DVSS DVSS nfet_06v0 ad=1.32p pd=6.88u as=0.78p ps=3.52u w=3u l=0.7u
D8 VSS OE diode_pd2nw_06v0 pj=1.92u area=0.2304p
X183 DVSS GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.pmos_6p0_CDNS_4066195314515_0.S DVDD DVDD pfet_06v0 ad=3.12p pd=12.52u as=3.12p ps=12.52u w=11.999999u l=0.7u
X184 DVDD GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_3.pmos_6p0_CDNS_4066195314512_0.D GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_3.Z DVDD pfet_06v0 ad=1.32p pd=6.88u as=0.78p ps=3.52u w=3u l=0.7u
X185 DVSS GF_NI_BI_T_BASE_0.comp018green_out_sigbuf_oe_0.nmos_6p0_CDNS_4066195314511_1.S GF_NI_BI_T_BASE_0.comp018green_out_sigbuf_oe_0.EN DVSS nfet_06v0 ad=0.78p pd=3.52u as=1.32p ps=6.88u w=3u l=0.7u
X186 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_cms_smt_0.nmos_6p0_CDNS_4066195314535_0.D GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_3.Z DVDD DVDD pfet_06v0 ad=1.04p pd=4.52u as=1.76p ps=8.88u w=4u l=0.7u
D9 SL VDD diode_pd2nw_06v0 pj=4u area=1p
X187 DVDD DVSS cap_nmos_06v0 c_width=3u c_length=3u
X188 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_0.pmos_6p0_CDNS_4066195314512_0.D GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_logic_pupd_0.PDB_OUT VSS VSS nfet_06v0 ad=0.66p pd=3.88u as=0.66p ps=3.88u w=1.5u l=0.7u
X189 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_cms_smt_0.nmos_6p0_CDNS_4066195314530_0.D GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_3.Z GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_drv_0.A DVSS nfet_06v0 ad=0.66p pd=3.88u as=0.66p ps=3.88u w=1.5u l=0.7u
X190 DVSS GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_drv_0.A GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_drv_0.nmos_6p0_CDNS_4066195314547_0.S DVSS nfet_06v0 ad=1.04p pd=4.52u as=1.76p ps=8.88u w=4u l=0.7u
X191 DVDD GF_NI_BI_T_BASE_0.comp018green_out_sigbuf_oe_2.nmos_6p0_CDNS_4066195314511_1.S GF_NI_BI_T_BASE_0.comp018green_out_predrv_1.EN DVDD pfet_06v0 ad=1.56p pd=6.52u as=2.64p ps=12.879999u w=6u l=0.7u
X192 GF_NI_BI_T_BASE_0.pdrive_x_<2> DVDD GF_NI_BI_T_BASE_0.pdrive_y_<2> DVSS nfet_06v0 ad=0.528p pd=3.28u as=0.528p ps=3.28u w=1.2u l=0.7u
X193 DVDD GF_NI_BI_T_BASE_0.comp018green_out_predrv_3.pmos_6p0_CDNS_4066195314515_0.D GF_NI_BI_T_BASE_0.pdrive_x_<1> DVDD pfet_06v0 ad=3.12p pd=12.52u as=3.12p ps=12.52u w=11.999999u l=0.7u
X194 DVDD DVSS cap_nmos_06v0 c_width=5u c_length=1.5u
X195 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_cms_smt_0.pmos_6p0_CDNS_4066195314538_0.S GF_NI_BI_T_BASE_0.comp018green_esd_cdm_0.IP_IN DVDD DVDD pfet_06v0 ad=0.836p pd=4.68u as=0.494p ps=2.42u w=1.9u l=0.7u
X196 GF_NI_BI_T_BASE_0.comp018green_out_sigbuf_oe_0.nmos_6p0_CDNS_4066195314511_0.S PDRV0 VSS VSS nfet_06v0 ad=0.78p pd=3.52u as=1.32p ps=6.88u w=3u l=0.7u
X197 VSS GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_drv_0.Z Y VSS nfet_06v0 ad=0.39p pd=2.02u as=0.39p ps=2.02u w=1.5u l=0.7u
X198 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_drv_0.Z GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_drv_0.nmos_6p0_CDNS_4066195314547_0.S VDD VDD pfet_06v0 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.7u
X199 DVSS DVSS PAD DVSS nfet_06v0_dss d_sab=0.28u s_sab=3.78u ad=10.639999p pd=76.56u as=0.14364n ps=83.56u w=38u l=1.15u
X200 DVDD GF_NI_BI_T_BASE_0.pdrive_y_<1> PAD DVDD pfet_06v0_dss d_sab=0.28u s_sab=2.78u ad=11.199999p pd=80.56u as=0.1112n ps=85.56u w=40u l=0.7u
X201 GF_NI_BI_T_BASE_0.ndrive_x_<1> GF_NI_BI_T_BASE_0.comp018green_out_predrv_3.pmos_6p0_CDNS_4066195314515_0.S DVSS DVSS nfet_06v0 ad=1.56p pd=6.52u as=1.56p ps=6.52u w=6u l=0.7u
X202 DVDD GF_NI_BI_T_BASE_0.comp018green_esd_cdm_0.IP_IN GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_cms_smt_0.pmos_6p0_CDNS_4066195314538_0.S DVDD pfet_06v0 ad=0.494p pd=2.42u as=0.836p ps=4.68u w=1.9u l=0.7u
X203 DVSS GF_NI_BI_T_BASE_0.comp018green_out_predrv_1.pmos_6p0_CDNS_4066195314515_0.S DVSS DVSS nfet_06v0 ad=1.56p pd=6.52u as=0 ps=0 w=6u l=0.7u
X204 DVSS GF_NI_BI_T_BASE_0.comp018green_out_predrv_3.pmos_6p0_CDNS_4066195314515_0.S DVSS DVSS nfet_06v0 ad=1.56p pd=6.52u as=0 ps=0 w=6u l=0.7u
X205 VDD GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_drv_0.nmos_6p0_CDNS_4066195314547_0.S GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_drv_0.Z VDD pfet_06v0 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.7u
X206 GF_NI_BI_T_BASE_0.comp018green_out_sigbuf_a_0.nmos_6p0_CDNS_4066195314511_3.S GF_NI_BI_T_BASE_0.comp018green_out_sigbuf_a_0.nmos_6p0_CDNS_4066195314511_1.D DVSS DVSS nfet_06v0 ad=1.32p pd=6.88u as=0.78p ps=3.52u w=3u l=0.7u
X207 DVDD GF_NI_BI_T_BASE_0.comp018green_sigbuf_1_0.pmos_6p0_CDNS_4066195314512_0.D GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.SL DVDD pfet_06v0 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.7u
X208 GF_NI_BI_T_BASE_0.pdrive_y_<3> GF_NI_BI_T_BASE_0.comp018green_out_predrv_1.pmos_6p0_CDNS_4066195314515_0.D DVDD DVDD pfet_06v0 ad=3.12p pd=12.52u as=3.12p ps=12.52u w=11.999999u l=0.7u
D10 PU VDD diode_pd2nw_06v0 pj=4u area=1p
X209 VSS GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_logic_pupd_0.comp018green_std_nand2_0.A GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_logic_pupd_0.comp018green_std_nand2_0.nmos_6p0_CDNS_4066195314511_0.D VSS nfet_06v0 ad=1.32p pd=6.88u as=0.78p ps=3.52u w=3u l=0.7u
X210 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_3.ZB GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_3.Z DVDD DVDD pfet_06v0 ad=0.78p pd=3.52u as=1.32p ps=6.88u w=3u l=0.7u
X211 DVSS GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_1.Z GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_1.ZB DVSS nfet_06v0 ad=0.66p pd=3.88u as=0.39p ps=2.02u w=1.5u l=0.7u
X212 PU PD GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_logic_pupd_0.comp018green_std_nand2_0.A VDD pfet_06v0 ad=1.32p pd=6.88u as=1.32p ps=6.88u w=3u l=0.7u
X213 DVSS GF_NI_BI_T_BASE_0.comp018green_out_predrv_1.pmos_6p0_CDNS_4066195314515_0.S DVDD DVDD pfet_06v0 ad=5.28p pd=24.88u as=3.12p ps=12.52u w=11.999999u l=0.7u
X214 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_1.ZB GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_1.Z DVSS DVSS nfet_06v0 ad=0.39p pd=2.02u as=0.39p ps=2.02u w=1.5u l=0.7u
X215 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_pupd_0.PU_B GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_2.pmos_6p0_CDNS_4066195314512_0.D DVDD DVDD pfet_06v0 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.7u
X216 GF_NI_BI_T_BASE_0.ndrive_x_<0> GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.pmos_6p0_CDNS_4066195314515_0.S DVSS DVSS nfet_06v0 ad=1.56p pd=6.52u as=2.64p ps=12.879999u w=6u l=0.7u
X217 DVSS GF_NI_BI_T_BASE_0.comp018green_out_predrv_2.pmos_6p0_CDNS_4066195314515_0.S GF_NI_BI_T_BASE_0.ndrive_x_<2> DVSS nfet_06v0 ad=1.56p pd=6.52u as=1.56p ps=6.52u w=6u l=0.7u
X218 VSS GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_drv_0.Z Y VSS nfet_06v0 ad=0.66p pd=3.88u as=0.39p ps=2.02u w=1.5u l=0.7u
X219 VDD GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_logic_pupd_0.comp018green_std_nand2_0.A GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_logic_pupd_0.PDB_OUT VDD pfet_06v0 ad=1.32p pd=6.88u as=0.78p ps=3.52u w=3u l=0.7u
X220 VDD OE GF_NI_BI_T_BASE_0.comp018green_out_sigbuf_oe_0.nmos_6p0_CDNS_4066195314511_1.S VDD pfet_06v0 ad=1.32p pd=6.88u as=0.78p ps=3.52u w=3u l=0.7u
X221 DVDD DVSS cap_nmos_06v0 c_width=5u c_length=1.5u
X222 DVDD DVSS cap_nmos_06v0 c_width=3u c_length=3u
X223 VSS CS GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_3.pmos_6p0_CDNS_4066195314512_0.D VSS nfet_06v0 ad=0.66p pd=3.88u as=0.66p ps=3.88u w=1.5u l=0.7u
X224 GF_NI_BI_T_BASE_0.comp018green_esd_cdm_0.IP_IN PAD w_4468_53342# ppolyf_u r_width=2.5u r_length=2.8u
X225 DVDD GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.SL GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.SLB DVDD pfet_06v0 ad=1.32p pd=6.88u as=0.78p ps=3.52u w=3u l=0.7u
X226 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_1.Z GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_1.pmos_6p0_CDNS_4066195314512_0.D DVDD DVDD pfet_06v0 ad=0.78p pd=3.52u as=1.32p ps=6.88u w=3u l=0.7u
X227 GF_NI_BI_T_BASE_0.comp018green_out_predrv_2.pmos_6p0_CDNS_4066195314515_0.D GF_NI_BI_T_BASE_0.comp018green_out_sigbuf_oe_1.ENB DVSS DVSS nfet_06v0 ad=1.56p pd=6.52u as=1.56p ps=6.52u w=6u l=0.7u
X228 VSS GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_drv_0.nmos_6p0_CDNS_4066195314547_0.S GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_drv_0.Z VSS nfet_06v0 ad=0.55p pd=3.38u as=0.325p ps=1.77u w=1.25u l=0.7u
X229 PAD GF_NI_BI_T_BASE_0.ndrive_x_<3> DVSS DVSS nfet_06v0_dss d_sab=3.78u s_sab=0.28u ad=0.14364n pd=83.56u as=10.639999p ps=76.56u w=38u l=1.15u
X230 DVDD GF_NI_BI_T_BASE_0.pdrive_x_<3> PAD DVDD pfet_06v0_dss d_sab=0.28u s_sab=2.78u ad=11.199999p pd=80.56u as=0.1112n ps=85.56u w=40u l=0.7u
X231 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_drv_0.Z GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_drv_0.nmos_6p0_CDNS_4066195314547_0.S VSS VSS nfet_06v0 ad=0.325p pd=1.77u as=0.55p ps=3.38u w=1.25u l=0.7u
X232 GF_NI_BI_T_BASE_0.comp018green_out_sigbuf_oe_0.ENB GF_NI_BI_T_BASE_0.comp018green_out_sigbuf_oe_0.EN DVDD DVDD pfet_06v0 ad=2.64p pd=12.879999u as=1.56p ps=6.52u w=6u l=0.7u
X233 GF_NI_BI_T_BASE_0.comp018green_out_predrv_3.pmos_6p0_CDNS_4066195314515_0.D GF_NI_BI_T_BASE_0.comp018green_out_sigbuf_oe_1.EN GF_NI_BI_T_BASE_0.comp018green_out_predrv_3.pmos_6p0_CDNS_4066195314515_0.S DVSS nfet_06v0 ad=1.56p pd=6.52u as=2.64p ps=12.879999u w=6u l=0.7u
X234 DVDD GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.pmos_6p0_CDNS_4066195314515_0.D GF_NI_BI_T_BASE_0.pdrive_y_<0> DVDD pfet_06v0 ad=3.12p pd=12.52u as=3.12p ps=12.52u w=11.999999u l=0.7u
X235 DVSS GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.A GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.pmos_6p0_CDNS_4066195314515_0.D DVSS nfet_06v0 ad=1.56p pd=6.52u as=2.64p ps=12.879999u w=6u l=0.7u
X236 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_cms_smt_0.nmos_6p0_CDNS_4066195314540_0.S GF_NI_BI_T_BASE_0.comp018green_esd_cdm_0.IP_IN GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_drv_0.A DVSS nfet_06v0 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.7u
X237 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_pupd_0.ppolyf_u_CDNS_4066195314533_3.MINUS GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_pupd_0.ppolyf_u_CDNS_4066195314533_4.PLUS DVDD ppolyf_u r_width=0.8u r_length=35.7u
X238 GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.SLB GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.SL DVSS DVSS nfet_06v0 ad=0.39p pd=2.02u as=0.39p ps=2.02u w=1.5u l=0.7u
X239 DVDD GF_NI_BI_T_BASE_0.comp018green_out_predrv_3.pmos_6p0_CDNS_4066195314515_0.S DVSS DVDD pfet_06v0 ad=3.12p pd=12.52u as=3.12p ps=12.52u w=11.999999u l=0.7u
X240 DVDD DVSS cap_nmos_06v0 c_width=5u c_length=1.5u
X241 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_3.Z GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_3.pmos_6p0_CDNS_4066195314512_0.D DVSS DVSS nfet_06v0 ad=0.39p pd=2.02u as=0.39p ps=2.02u w=1.5u l=0.7u
X242 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_pupd_0.PD GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_0.Z DVSS DVSS nfet_06v0 ad=0.39p pd=2.02u as=0.39p ps=2.02u w=1.5u l=0.7u
X243 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_drv_0.A GF_NI_BI_T_BASE_0.comp018green_esd_cdm_0.IP_IN GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_cms_smt_0.nmos_6p0_CDNS_4066195314540_0.S DVSS nfet_06v0 ad=0.78p pd=3.52u as=1.32p ps=6.88u w=3u l=0.7u
D11 GF_NI_BI_T_BASE_0.comp018green_esd_cdm_0.IP_IN DVDD diode_pd2nw_06v0 pj=42u area=20p
X244 GF_NI_BI_T_BASE_0.ndrive_x_<3> GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.SL DVSS DVDD pfet_06v0 ad=3.12p pd=12.52u as=5.28p ps=24.88u w=11.999999u l=0.7u
X245 GF_NI_BI_T_BASE_0.pdrive_y_<2> GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.SLB GF_NI_BI_T_BASE_0.pdrive_x_<2> DVSS nfet_06v0 ad=1.56p pd=6.52u as=2.64p ps=12.879999u w=6u l=0.7u
X246 DVDD DVSS cap_nmos_06v0 c_width=5u c_length=1.5u
X247 Y GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_drv_0.Z VDD VDD pfet_06v0 ad=0.91p pd=4.02u as=0.91p ps=4.02u w=3.5u l=0.7u
X248 GF_NI_BI_T_BASE_0.comp018green_out_predrv_1.ENB GF_NI_BI_T_BASE_0.comp018green_out_predrv_1.EN DVSS DVSS nfet_06v0 ad=1.32p pd=6.88u as=0.78p ps=3.52u w=3u l=0.7u
X249 DVSS GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.SL GF_NI_BI_T_BASE_0.ndrive_x_<1> DVDD pfet_06v0 ad=3.12p pd=12.52u as=3.12p ps=12.52u w=11.999999u l=0.7u
X250 DVSS GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_3.Z GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_3.ZB DVSS nfet_06v0 ad=0.39p pd=2.02u as=0.39p ps=2.02u w=1.5u l=0.7u
X251 DVSS GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_0.pmos_6p0_CDNS_4066195314512_0.D GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_0.Z DVSS nfet_06v0 ad=0.39p pd=2.02u as=0.39p ps=2.02u w=1.5u l=0.7u
X252 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_drv_0.A GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_1.Z DVDD DVDD pfet_06v0 ad=0.52p pd=2.52u as=0.88p ps=4.88u w=2u l=0.7u
X253 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_drv_0.A GF_NI_BI_T_BASE_0.comp018green_esd_cdm_0.IP_IN GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_cms_smt_0.pmos_6p0_CDNS_4066195314538_0.S DVDD pfet_06v0 ad=0.559p pd=2.67u as=0.946p ps=5.18u w=2.15u l=0.7u
X254 Y GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_drv_0.Z VSS VSS nfet_06v0 ad=0.39p pd=2.02u as=0.39p ps=2.02u w=1.5u l=0.7u
X255 GF_NI_BI_T_BASE_0.comp018green_out_predrv_2.pmos_6p0_CDNS_4066195314515_0.S GF_NI_BI_T_BASE_0.comp018green_out_sigbuf_oe_1.ENB GF_NI_BI_T_BASE_0.comp018green_out_predrv_2.pmos_6p0_CDNS_4066195314515_0.D DVDD pfet_06v0 ad=3.12p pd=12.52u as=5.28p ps=24.88u w=11.999999u l=0.7u
X256 GF_NI_BI_T_BASE_0.pdrive_y_<1> GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.SLB GF_NI_BI_T_BASE_0.pdrive_x_<1> DVSS nfet_06v0 ad=1.56p pd=6.52u as=2.64p ps=12.879999u w=6u l=0.7u
X257 GF_NI_BI_T_BASE_0.comp018green_out_predrv_1.pmos_6p0_CDNS_4066195314515_0.D GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.A DVSS DVSS nfet_06v0 ad=2.64p pd=12.879999u as=1.56p ps=6.52u w=6u l=0.7u
X258 GF_NI_BI_T_BASE_0.ndrive_x_<1> DVSS DVSS DVDD pfet_06v0 ad=0.528p pd=3.28u as=0.528p ps=3.28u w=1.2u l=0.7u
X259 VSS PDRV1 GF_NI_BI_T_BASE_0.comp018green_out_sigbuf_oe_1.nmos_6p0_CDNS_4066195314511_0.S VSS nfet_06v0 ad=1.32p pd=6.88u as=0.78p ps=3.52u w=3u l=0.7u
X260 GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.SL GF_NI_BI_T_BASE_0.comp018green_sigbuf_1_0.pmos_6p0_CDNS_4066195314512_0.D DVDD DVDD pfet_06v0 ad=0.78p pd=3.52u as=1.32p ps=6.88u w=3u l=0.7u
X261 DVSS GF_NI_BI_T_BASE_0.comp018green_out_predrv_2.pmos_6p0_CDNS_4066195314515_0.S DVDD DVDD pfet_06v0 ad=3.12p pd=12.52u as=3.12p ps=12.52u w=11.999999u l=0.7u
X262 DVDD GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.pmos_6p0_CDNS_4066195314515_0.S DVSS DVDD pfet_06v0 ad=3.12p pd=12.52u as=5.28p ps=24.88u w=11.999999u l=0.7u
X263 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_logic_pupd_0.comp018green_std_nand2_0.nmos_6p0_CDNS_4066195314511_0.D PD GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_logic_pupd_0.PDB_OUT VSS nfet_06v0 ad=0.78p pd=3.52u as=1.32p ps=6.88u w=3u l=0.7u
X264 GF_NI_BI_T_BASE_0.comp018green_out_sigbuf_oe_1.nmos_6p0_CDNS_4066195314511_0.S OE GF_NI_BI_T_BASE_0.comp018green_out_sigbuf_oe_1.nmos_6p0_CDNS_4066195314511_1.S VSS nfet_06v0 ad=0.78p pd=3.52u as=1.32p ps=6.88u w=3u l=0.7u
X265 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_drv_0.nmos_6p0_CDNS_4066195314547_0.S GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_drv_0.A DVDD DVDD pfet_06v0 ad=0.88p pd=4.88u as=0.88p ps=4.88u w=2u l=0.7u
X266 VSS OE GF_NI_BI_T_BASE_0.comp018green_out_sigbuf_a_0.nmos_6p0_CDNS_4066195314511_1.S VSS nfet_06v0 ad=1.32p pd=6.88u as=0.78p ps=3.52u w=3u l=0.7u
D12 DVSS GF_NI_BI_T_BASE_0.comp018green_esd_cdm_0.IP_IN diode_nd2ps_06v0 pj=42u area=20p
X267 GF_NI_BI_T_BASE_0.comp018green_out_sigbuf_a_0.nmos_6p0_CDNS_4066195314511_1.S A GF_NI_BI_T_BASE_0.comp018green_out_sigbuf_a_0.nmos_6p0_CDNS_4066195314511_1.D VSS nfet_06v0 ad=0.78p pd=3.52u as=1.32p ps=6.88u w=3u l=0.7u
X268 GF_NI_BI_T_BASE_0.ndrive_x_<2> GF_NI_BI_T_BASE_0.comp018green_out_predrv_2.pmos_6p0_CDNS_4066195314515_0.S DVSS DVSS nfet_06v0 ad=1.56p pd=6.52u as=2.64p ps=12.879999u w=6u l=0.7u
X269 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_logic_pupd_0.PDB_OUT PD VDD VDD pfet_06v0 ad=0.78p pd=3.52u as=1.32p ps=6.88u w=3u l=0.7u
X270 DVDD GF_NI_BI_T_BASE_0.pdrive_x_<2> PAD DVDD pfet_06v0_dss d_sab=0.28u s_sab=2.78u ad=11.199999p pd=80.56u as=0.1112n ps=85.56u w=40u l=0.7u
X271 DVSS GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_pupd_0.PU_B GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_2.ZB DVSS nfet_06v0 ad=0.39p pd=2.02u as=0.39p ps=2.02u w=1.5u l=0.7u
D13 VSS PDRV1 diode_pd2nw_06v0 pj=1.92u area=0.2304p
X272 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_logic_pupd_0.comp018green_std_xor2_0.pmos_6p0_CDNS_4066195314512_2.D PD VSS VSS nfet_06v0 ad=0.66p pd=3.88u as=0.66p ps=3.88u w=1.5u l=0.7u
X273 GF_NI_BI_T_BASE_0.comp018green_esd_cdm_0.IP_IN PAD w_4468_53342# ppolyf_u r_width=2.5u r_length=2.8u
X274 GF_NI_BI_T_BASE_0.comp018green_out_sigbuf_oe_1.EN GF_NI_BI_T_BASE_0.comp018green_out_sigbuf_oe_1.nmos_6p0_CDNS_4066195314511_1.S DVDD DVDD pfet_06v0 ad=2.64p pd=12.879999u as=1.56p ps=6.52u w=6u l=0.7u
X275 GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.pmos_6p0_CDNS_4066195314515_0.S GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.A DVDD DVDD pfet_06v0 ad=5.28p pd=24.88u as=3.12p ps=12.52u w=11.999999u l=0.7u
X276 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_2.ZB GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_pupd_0.PU_B DVSS DVSS nfet_06v0 ad=0.39p pd=2.02u as=0.66p ps=3.88u w=1.5u l=0.7u
X277 DVDD GF_NI_BI_T_BASE_0.comp018green_out_sigbuf_oe_0.nmos_6p0_CDNS_4066195314511_1.S GF_NI_BI_T_BASE_0.comp018green_out_sigbuf_oe_0.EN DVDD pfet_06v0 ad=1.56p pd=6.52u as=2.64p ps=12.879999u w=6u l=0.7u
X278 DVDD GF_NI_BI_T_BASE_0.comp018green_out_sigbuf_oe_0.EN GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.pmos_6p0_CDNS_4066195314515_0.S DVDD pfet_06v0 ad=3.12p pd=12.52u as=3.12p ps=12.52u w=11.999999u l=0.7u
X279 DVSS GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_3.Z GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_cms_smt_0.nmos_6p0_CDNS_4066195314535_0.D DVSS nfet_06v0 ad=0.88p pd=4.88u as=0.52p ps=2.52u w=2u l=0.7u
X280 PAD GF_NI_BI_T_BASE_0.pdrive_x_<0> DVDD DVDD pfet_06v0_dss d_sab=2.78u s_sab=0.28u ad=0.1112n pd=85.56u as=11.199999p ps=80.56u w=40u l=0.7u
X281 GF_NI_BI_T_BASE_0.pdrive_x_<2> GF_NI_BI_T_BASE_0.comp018green_out_predrv_2.pmos_6p0_CDNS_4066195314515_0.D DVDD DVDD pfet_06v0 ad=3.12p pd=12.52u as=3.12p ps=12.52u w=11.999999u l=0.7u
X282 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_drv_0.A GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_cms_smt_0.nmos_6p0_CDNS_4066195314535_0.D GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_cms_smt_0.pmos_6p0_CDNS_4066195314534_0.D DVDD pfet_06v0 ad=0.88p pd=4.88u as=0.88p ps=4.88u w=2u l=0.7u
X283 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_pupd_0.pmos_6p0_CDNS_4066195314512_0.D GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_pupd_0.PD DVSS DVSS nfet_06v0 ad=0.66p pd=3.88u as=0.66p ps=3.88u w=1.5u l=0.7u
X284 DVSS GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.pmos_6p0_CDNS_4066195314515_0.S DVSS DVSS nfet_06v0 ad=1.56p pd=6.52u as=0 ps=0 w=6u l=0.7u
X285 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_cms_smt_0.nmos_6p0_CDNS_4066195314537_0.D GF_NI_BI_T_BASE_0.comp018green_esd_cdm_0.IP_IN GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_cms_smt_0.nmos_6p0_CDNS_4066195314540_0.S DVSS nfet_06v0 ad=0.689p pd=3.17u as=0.689p ps=3.17u w=2.65u l=0.7u
X286 DVSS GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.pmos_6p0_CDNS_4066195314515_0.S DVSS DVSS nfet_06v0 ad=1.56p pd=6.52u as=0 ps=0 w=6u l=0.7u
X287 GF_NI_BI_T_BASE_0.comp018green_out_predrv_3.pmos_6p0_CDNS_4066195314515_0.D GF_NI_BI_T_BASE_0.comp018green_out_sigbuf_oe_1.ENB GF_NI_BI_T_BASE_0.comp018green_out_predrv_3.pmos_6p0_CDNS_4066195314515_0.S DVDD pfet_06v0 ad=5.28p pd=24.88u as=3.12p ps=12.52u w=11.999999u l=0.7u
X288 GF_NI_BI_T_BASE_0.pdrive_x_<1> GF_NI_BI_T_BASE_0.comp018green_out_predrv_3.pmos_6p0_CDNS_4066195314515_0.D DVDD DVDD pfet_06v0 ad=3.12p pd=12.52u as=5.28p ps=24.88u w=11.999999u l=0.7u
D14 PD VDD diode_pd2nw_06v0 pj=4u area=1p
X289 VDD GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_logic_pupd_0.PUB_OUT GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_2.pmos_6p0_CDNS_4066195314512_0.D VDD pfet_06v0 ad=1.32p pd=6.88u as=1.32p ps=6.88u w=3u l=0.7u
X290 DVDD GF_NI_BI_T_BASE_0.comp018green_out_predrv_0.A GF_NI_BI_T_BASE_0.comp018green_out_predrv_1.pmos_6p0_CDNS_4066195314515_0.S DVDD pfet_06v0 ad=3.12p pd=12.52u as=5.28p ps=24.88u w=11.999999u l=0.7u
X291 DVSS GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_1.Z GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_cms_smt_0.nmos_6p0_CDNS_4066195314537_0.D DVSS nfet_06v0 ad=0.832p pd=3.72u as=0.832p ps=3.72u w=3.2u l=0.7u
X292 DVDD GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_3.Z GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_cms_smt_0.nmos_6p0_CDNS_4066195314535_0.D DVDD pfet_06v0 ad=1.76p pd=8.88u as=1.04p ps=4.52u w=4u l=0.7u
X293 GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_in_cms_smt_0.nmos_6p0_CDNS_4066195314537_0.D GF_NI_BI_T_BASE_0.comp018green_inpath_cms_smt_0.comp018green_sigbuf_1.Z DVSS DVSS nfet_06v0 ad=0.832p pd=3.72u as=0.832p ps=3.72u w=3.2u l=0.7u
D15 VSS PDRV0 diode_pd2nw_06v0 pj=1.92u area=0.2304p
X294 DVDD GF_NI_BI_T_BASE_0.comp018green_out_predrv_2.pmos_6p0_CDNS_4066195314515_0.S DVSS DVDD pfet_06v0 ad=3.12p pd=12.52u as=5.28p ps=24.88u w=11.999999u l=0.7u
X295 GF_NI_BI_T_BASE_0.comp018green_out_sigbuf_a_0.nmos_6p0_CDNS_4066195314511_3.S GF_NI_BI_T_BASE_0.comp018green_out_sigbuf_a_0.nmos_6p0_CDNS_4066195314511_1.D DVDD DVDD pfet_06v0 ad=2.64p pd=12.879999u as=1.56p ps=6.52u w=6u l=0.7u
X296 DVSS GF_NI_BI_T_BASE_0.comp018green_out_predrv_3.pmos_6p0_CDNS_4066195314515_0.S GF_NI_BI_T_BASE_0.ndrive_x_<1> DVSS nfet_06v0 ad=2.64p pd=12.879999u as=1.56p ps=6.52u w=6u l=0.7u
.ends

