** sch_path: /workspaces/gf180-io-verification/test/digital_io_switching_pex/digital_io_switching_pex.sch
**.subckt digital_io_switching_pex
V1 DVDD GND 3
V2 VDD GND 3
V3 DVSS GND 0
V4 VSS GND 0
V5 A GND PULSE(0 3 10n 100p 100p 10n 20n)
V7 IE GND 3
V8 OE GND 3
V9 PU GND 0
V10 PD GND 0
V11 SL GND 0
V13 CS GND 3.3
**** begin user architecture code


.tran 100p 100n
.save all
.control
run
display
plot A PAD0 Y0
plot PAD0 PAD1
.endc



.include /home/designer/.volare/gf180mcuD/libs.tech/ngspice/design.ngspice
.lib /home/designer/.volare/gf180mcuD/libs.tech/ngspice/sm141064.ngspice typical
.lib /home/designer/.volare/gf180mcuD/libs.tech/ngspice/sm141064.ngspice diode_typical
.lib /home/designer/.volare/gf180mcuD/libs.tech/ngspice/sm141064.ngspice res_typical
.lib /home/designer/.volare/gf180mcuD/libs.tech/ngspice/sm141064.ngspice mimcap_typical
.lib /home/designer/.volare/gf180mcuD/libs.tech/ngspice/sm141064.ngspice moscap_typical


.include ./gf180mcu_fd_io.spice
.include ./gf180mcu_fd_io__bi_t_extracted.spice
XDUT0 A CS DVDD DVSS IE OE PAD0 PD VSS VSS PU SL VDD VSS Y0 gf180mcu_fd_io__bi_t
XDUT1 A CS DVDD DVSS IE OE PAD1 PD VSS VSS PU SL VDD VSS Y1 gf180mcu_fd_io__bi_t_extracted

**** end user architecture code
**.ends
.GLOBAL GND
.end
