* NGSPICE file created from gf180mcu_fd_io__in_c.ext - technology: gf180mcuD

.subckt x5LM_METAL_RAIL_PAD_60 Bondpad_5LM_0/m5_n400_0# 5LM_METAL_RAIL_0/VSS 5LM_METAL_RAIL_0/VDD
+ 5LM_METAL_RAIL_0/DVSS 5LM_METAL_RAIL_0/DVDD VSUBS
.ends

.subckt nmoscap_6p0_CDNS_4066195314523 G D
X0 G D cap_nmos_06v0 c_width=5u c_length=1.5u
.ends

.subckt comp018green_out_drv_pleg_4T_Y w_0_12# a_278_44# a_974_132# a_222_132#
X0 a_974_132# a_278_44# a_222_132# w_0_12# pfet_06v0_dss d_sab=2.78u s_sab=0.28u ad=0.1112n pd=85.56u as=11.199999p ps=80.56u w=40u l=0.7u
.ends

.subckt comp018green_out_drv_pleg_4T_X a_1662_44# w_0_12# a_278_44# a_1858_132# a_974_132#
+ a_222_132#
X0 a_974_132# a_278_44# a_222_132# w_0_12# pfet_06v0_dss d_sab=2.78u s_sab=0.28u ad=0.1112n pd=85.56u as=11.199999p ps=80.56u w=40u l=0.7u
X1 a_1858_132# a_1662_44# a_974_132# w_0_12# pfet_06v0_dss d_sab=0.28u s_sab=2.78u ad=11.199999p pd=80.56u as=0.1112n ps=85.56u w=40u l=0.7u
.ends

.subckt comp018green_out_paddrv_4T_PMOS_GROUP a_2360_2800# a_4511_2800# PMOS_4T_metal_stack_5/m2_340_0#
+ PMOS_4T_metal_stack_1/m2_340_0# PMOS_4T_metal_stack_6/m2_340_0# a_n767_13534# PMOS_4T_metal_stack_2/m2_340_0#
+ a_9428_2800# a_7662_2800# a_11201_2800# a_9815_2800# PMOS_4T_metal_stack_3/m2_340_0#
+ a_6280_2800# a_2746_2800# a_974_2800# a_8049_2800# a_5892_2800# PMOS_4T_metal_stack_1/m2_n44_0#
+ w_n2_111# PMOS_4T_metal_stack_4/m2_340_0# PMOS_4T_metal_stack_2/m2_n44_0# a_4120_2800#
+ PMOS_4T_metal_stack_6/VSUBS PMOS_4T_metal_stack_3/m2_n44_0# PMOS_4T_metal_stack_4/m2_n44_0#
+ PMOS_4T_metal_stack_5/m2_n44_0#
Xcomp018green_out_drv_pleg_4T_Y_0 w_n2_111# a_4120_2800# PMOS_4T_metal_stack_1/m2_340_0#
+ PMOS_4T_metal_stack_2/m2_n44_0# comp018green_out_drv_pleg_4T_Y
Xcomp018green_out_drv_pleg_4T_Y_1 w_n2_111# a_9428_2800# PMOS_4T_metal_stack_4/m2_340_0#
+ PMOS_4T_metal_stack_5/m2_n44_0# comp018green_out_drv_pleg_4T_Y
Xcomp018green_out_drv_pleg_4T_Y_2 w_n2_111# a_2746_2800# PMOS_4T_metal_stack_1/m2_340_0#
+ PMOS_4T_metal_stack_1/m2_n44_0# comp018green_out_drv_pleg_4T_Y
Xcomp018green_out_drv_pleg_4T_Y_3 w_n2_111# a_8049_2800# PMOS_4T_metal_stack_4/m2_340_0#
+ PMOS_4T_metal_stack_4/m2_n44_0# comp018green_out_drv_pleg_4T_Y
Xcomp018green_out_drv_pleg_4T_X_0 a_4511_2800# w_n2_111# a_5892_2800# PMOS_4T_metal_stack_2/m2_n44_0#
+ PMOS_4T_metal_stack_2/m2_340_0# PMOS_4T_metal_stack_3/m2_n44_0# comp018green_out_drv_pleg_4T_X
Xcomp018green_out_drv_pleg_4T_X_1 a_9815_2800# w_n2_111# a_11201_2800# PMOS_4T_metal_stack_5/m2_n44_0#
+ PMOS_4T_metal_stack_5/m2_340_0# w_n2_111# comp018green_out_drv_pleg_4T_X
Xcomp018green_out_drv_pleg_4T_X_2 a_7662_2800# w_n2_111# a_6280_2800# PMOS_4T_metal_stack_4/m2_n44_0#
+ PMOS_4T_metal_stack_3/m2_340_0# PMOS_4T_metal_stack_3/m2_n44_0# comp018green_out_drv_pleg_4T_X
Xcomp018green_out_drv_pleg_4T_X_3 a_2360_2800# w_n2_111# a_974_2800# PMOS_4T_metal_stack_1/m2_n44_0#
+ PMOS_4T_metal_stack_6/m2_340_0# w_n2_111# comp018green_out_drv_pleg_4T_X
.ends

.subckt comp018green_out_drv_nleg_4T a_206_444# a_2080_444# a_2366_532# a_48_532#
+ a_436_532# VSUBS
X0 a_436_532# a_206_444# a_48_532# VSUBS nfet_06v0_dss d_sab=3.78u s_sab=0.28u ad=0.14364n pd=83.56u as=10.639999p ps=76.56u w=38u l=1.15u
X1 a_2366_532# a_2080_444# a_436_532# VSUBS nfet_06v0_dss d_sab=0.28u s_sab=3.78u ad=10.639999p pd=76.56u as=0.14364n ps=83.56u w=38u l=1.15u
.ends

.subckt comp018green_out_paddrv_4T_NMOS_GROUP a_7847_1028# a_7373_1028# GR_NMOS_4T_0/w_n1730_n583#
+ a_803_1028# a_2677_1028# nmos_4T_metal_stack_1/m2_430_401# a_9721_1028# nmos_4T_metal_stack_2/m2_430_401#
+ nmos_4T_metal_stack_4/m2_430_401# nmos_4T_metal_stack_3/m2_430_401# a_5499_1028#
+ nmos_4T_metal_stack_0/m2_n44_400# a_3151_1028# VSUBS a_5025_1028# nmos_4T_metal_stack_4/m2_n44_400#
+ nmos_4T_metal_stack_1/m2_n44_400# nmos_4T_metal_stack_2/m2_n44_400# nmos_4T_metal_stack_3/m2_n44_400#
Xcomp018green_out_drv_nleg_4T_0 a_7847_1028# a_9721_1028# nmos_4T_metal_stack_0/m2_n44_400#
+ nmos_4T_metal_stack_3/m2_n44_400# nmos_4T_metal_stack_3/m2_430_401# VSUBS comp018green_out_drv_nleg_4T
Xcomp018green_out_drv_nleg_4T_1 a_5499_1028# a_7373_1028# nmos_4T_metal_stack_3/m2_n44_400#
+ nmos_4T_metal_stack_2/m2_n44_400# nmos_4T_metal_stack_2/m2_430_401# VSUBS comp018green_out_drv_nleg_4T
Xcomp018green_out_drv_nleg_4T_2 a_3151_1028# a_5025_1028# nmos_4T_metal_stack_2/m2_n44_400#
+ nmos_4T_metal_stack_1/m2_n44_400# nmos_4T_metal_stack_1/m2_430_401# VSUBS comp018green_out_drv_nleg_4T
Xcomp018green_out_drv_nleg_4T_3 a_803_1028# a_2677_1028# nmos_4T_metal_stack_1/m2_n44_400#
+ nmos_4T_metal_stack_4/m2_n44_400# nmos_4T_metal_stack_4/m2_430_401# VSUBS comp018green_out_drv_nleg_4T
.ends

.subckt comp018green_out_paddrv_16T comp018green_out_paddrv_4T_PMOS_GROUP_0/a_7662_2800#
+ comp018green_out_paddrv_4T_PMOS_GROUP_0/a_11201_2800# comp018green_out_paddrv_4T_PMOS_GROUP_0/a_9428_2800#
+ comp018green_out_paddrv_4T_PMOS_GROUP_0/a_9815_2800# m1_12305_8954# comp018green_out_paddrv_4T_PMOS_GROUP_0/a_974_2800#
+ comp018green_out_paddrv_4T_PMOS_GROUP_0/a_6280_2800# comp018green_out_paddrv_4T_PMOS_GROUP_0/a_2746_2800#
+ m1_1026_8954# m1_12305_9280# comp018green_out_paddrv_4T_PMOS_GROUP_0/a_8049_2800#
+ comp018green_out_paddrv_4T_PMOS_GROUP_0/a_5892_2800# m1_12305_9120# comp018green_out_paddrv_4T_PMOS_GROUP_0/a_4120_2800#
+ m1_1026_9280# m1_1026_9120# comp018green_out_paddrv_4T_PMOS_GROUP_0/a_2360_2800#
+ m1_12305_9446# comp018green_out_paddrv_4T_NMOS_GROUP_0/nmos_4T_metal_stack_2/m2_n44_400#
+ comp018green_out_paddrv_4T_PMOS_GROUP_0/a_4511_2800# comp018green_out_paddrv_4T_NMOS_GROUP_0/nmos_4T_metal_stack_3/m2_n44_400#
+ m2_1697_23319# comp018green_out_paddrv_4T_PMOS_GROUP_0/PMOS_4T_metal_stack_5/m2_n44_0#
+ comp018green_out_paddrv_4T_PMOS_GROUP_0/w_n2_111# m1_1026_9446# comp018green_out_paddrv_4T_NMOS_GROUP_0/nmos_4T_metal_stack_1/m2_n44_400#
+ m1_n360_8434# comp018green_out_paddrv_4T_PMOS_GROUP_0/PMOS_4T_metal_stack_1/m2_n44_0#
+ comp018green_out_paddrv_4T_PMOS_GROUP_0/PMOS_4T_metal_stack_4/m2_n44_0# comp018green_out_paddrv_4T_PMOS_GROUP_0/PMOS_4T_metal_stack_2/m2_n44_0#
+ comp018green_out_paddrv_4T_NMOS_GROUP_0/VSUBS comp018green_out_paddrv_4T_PMOS_GROUP_0/PMOS_4T_metal_stack_3/m2_n44_0#
Xcomp018green_out_paddrv_4T_PMOS_GROUP_0 comp018green_out_paddrv_4T_PMOS_GROUP_0/a_2360_2800#
+ comp018green_out_paddrv_4T_PMOS_GROUP_0/a_4511_2800# m2_1697_23319# m2_1697_23319#
+ m2_1697_23319# comp018green_out_paddrv_4T_NMOS_GROUP_0/VSUBS m2_1697_23319# comp018green_out_paddrv_4T_PMOS_GROUP_0/a_9428_2800#
+ comp018green_out_paddrv_4T_PMOS_GROUP_0/a_7662_2800# comp018green_out_paddrv_4T_PMOS_GROUP_0/a_11201_2800#
+ comp018green_out_paddrv_4T_PMOS_GROUP_0/a_9815_2800# m2_1697_23319# comp018green_out_paddrv_4T_PMOS_GROUP_0/a_6280_2800#
+ comp018green_out_paddrv_4T_PMOS_GROUP_0/a_2746_2800# comp018green_out_paddrv_4T_PMOS_GROUP_0/a_974_2800#
+ comp018green_out_paddrv_4T_PMOS_GROUP_0/a_8049_2800# comp018green_out_paddrv_4T_PMOS_GROUP_0/a_5892_2800#
+ comp018green_out_paddrv_4T_PMOS_GROUP_0/PMOS_4T_metal_stack_1/m2_n44_0# comp018green_out_paddrv_4T_PMOS_GROUP_0/w_n2_111#
+ m2_1697_23319# comp018green_out_paddrv_4T_PMOS_GROUP_0/PMOS_4T_metal_stack_2/m2_n44_0#
+ comp018green_out_paddrv_4T_PMOS_GROUP_0/a_4120_2800# comp018green_out_paddrv_4T_NMOS_GROUP_0/VSUBS
+ comp018green_out_paddrv_4T_PMOS_GROUP_0/PMOS_4T_metal_stack_3/m2_n44_0# comp018green_out_paddrv_4T_PMOS_GROUP_0/PMOS_4T_metal_stack_4/m2_n44_0#
+ comp018green_out_paddrv_4T_PMOS_GROUP_0/PMOS_4T_metal_stack_5/m2_n44_0# comp018green_out_paddrv_4T_PMOS_GROUP
Xcomp018green_out_paddrv_4T_NMOS_GROUP_0 m1_12305_9120# m1_12305_9280# m1_n360_8434#
+ m1_1026_8954# m1_1026_9120# m2_1697_23319# m1_12305_8954# m2_1697_23319# m2_1697_23319#
+ m2_1697_23319# m1_12305_9446# comp018green_out_paddrv_4T_NMOS_GROUP_0/VSUBS m1_1026_9280#
+ comp018green_out_paddrv_4T_NMOS_GROUP_0/VSUBS m1_1026_9446# comp018green_out_paddrv_4T_NMOS_GROUP_0/VSUBS
+ comp018green_out_paddrv_4T_NMOS_GROUP_0/nmos_4T_metal_stack_1/m2_n44_400# comp018green_out_paddrv_4T_NMOS_GROUP_0/nmos_4T_metal_stack_2/m2_n44_400#
+ comp018green_out_paddrv_4T_NMOS_GROUP_0/nmos_4T_metal_stack_3/m2_n44_400# comp018green_out_paddrv_4T_NMOS_GROUP
.ends

.subckt nmos_6p0_CDNS_4066195314531 D a_0_n44# S a_244_n44#
X0 S a_244_n44# D VSUBS nfet_06v0 ad=0.66p pd=3.88u as=0.39p ps=2.02u w=1.5u l=0.7u
X1 D a_0_n44# S VSUBS nfet_06v0 ad=0.39p pd=2.02u as=0.66p ps=3.88u w=1.5u l=0.7u
.ends

.subckt nmos_6p0_CDNS_4066195314530 D a_0_n44# S VSUBS
X0 D a_0_n44# S VSUBS nfet_06v0 ad=0.66p pd=3.88u as=0.66p ps=3.88u w=1.5u l=0.7u
.ends

.subckt comp018green_sigbuf_1 Z VSS A VDD ZB DVSS DVDD
Xnmos_6p0_CDNS_4066195314531_0 ZB Z DVSS Z nmos_6p0_CDNS_4066195314531
Xnmos_6p0_CDNS_4066195314531_1 Z nmos_6p0_CDNS_4066195314530_0/D DVSS nmos_6p0_CDNS_4066195314530_0/D
+ nmos_6p0_CDNS_4066195314531
Xnmos_6p0_CDNS_4066195314530_0 nmos_6p0_CDNS_4066195314530_0/D A VSS VSS nmos_6p0_CDNS_4066195314530
X0 Z nmos_6p0_CDNS_4066195314530_0/D DVDD DVDD pfet_06v0 ad=0.78p pd=3.52u as=1.32p ps=6.88u w=3u l=0.7u
X1 ZB Z DVDD DVDD pfet_06v0 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.7u
X2 DVDD Z ZB DVDD pfet_06v0 ad=1.32p pd=6.88u as=0.78p ps=3.52u w=3u l=0.7u
X3 DVDD nmos_6p0_CDNS_4066195314530_0/D Z DVDD pfet_06v0 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.7u
X4 nmos_6p0_CDNS_4066195314530_0/D A VDD VDD pfet_06v0 ad=1.32p pd=6.88u as=1.32p ps=6.88u w=3u l=0.7u
.ends

.subckt nmos_6p0_CDNS_4066195314514 D a_0_n44# S
X0 D a_0_n44# S VSUBS nfet_06v0 ad=0.528p pd=3.28u as=0.528p ps=3.28u w=1.2u l=0.7u
.ends

.subckt nmos_6p0_CDNS_4066195314519 D a_0_n44# S
X0 D a_0_n44# S VSUBS nfet_06v0 ad=2.64p pd=12.879999u as=2.64p ps=12.879999u w=6u l=0.7u
.ends

.subckt nmos_6p0_CDNS_4066195314520 D a_0_n44# S a_244_n44#
X0 S a_244_n44# D VSUBS nfet_06v0 ad=2.64p pd=12.879999u as=1.56p ps=6.52u w=6u l=0.7u
X1 D a_0_n44# S VSUBS nfet_06v0 ad=1.56p pd=6.52u as=2.64p ps=12.879999u w=6u l=0.7u
.ends

.subckt nmos_6p0_CDNS_4066195314518 D a_0_n44# S a_244_n44#
X0 S a_244_n44# D VSUBS nfet_06v0 ad=2.64p pd=12.879999u as=1.56p ps=6.52u w=6u l=0.7u
X1 D a_0_n44# S VSUBS nfet_06v0 ad=1.56p pd=6.52u as=2.64p ps=12.879999u w=6u l=0.7u
.ends

.subckt comp018green_out_predrv SL SLB NDRIVE_X ENB A NDRIVE_Y PDRIVE_Y PDRIVE_X EN
+ DVDD DVSS
Xnmos_6p0_CDNS_4066195314514_0 PDRIVE_X DVDD PDRIVE_Y nmos_6p0_CDNS_4066195314514
Xnmos_6p0_CDNS_4066195314519_0 nmos_6p0_CDNS_4066195314519_2/D A DVSS nmos_6p0_CDNS_4066195314519
Xnmos_6p0_CDNS_4066195314519_1 DVSS ENB nmos_6p0_CDNS_4066195314519_2/D nmos_6p0_CDNS_4066195314519
Xnmos_6p0_CDNS_4066195314519_2 nmos_6p0_CDNS_4066195314519_2/D EN nmos_6p0_CDNS_4066195314519_2/S
+ nmos_6p0_CDNS_4066195314519
Xnmos_6p0_CDNS_4066195314520_0 NDRIVE_X nmos_6p0_CDNS_4066195314519_2/S DVSS nmos_6p0_CDNS_4066195314519_2/S
+ nmos_6p0_CDNS_4066195314520
Xnmos_6p0_CDNS_4066195314520_1 PDRIVE_Y SLB PDRIVE_X SLB nmos_6p0_CDNS_4066195314520
Xnmos_6p0_CDNS_4066195314518_0 PDRIVE_Y nmos_6p0_CDNS_4066195314519_2/D DVSS nmos_6p0_CDNS_4066195314519_2/D
+ nmos_6p0_CDNS_4066195314518
Xnmos_6p0_CDNS_4066195314518_1 NDRIVE_Y nmos_6p0_CDNS_4066195314519_2/S DVSS nmos_6p0_CDNS_4066195314519_2/S
+ nmos_6p0_CDNS_4066195314518
X0 DVDD nmos_6p0_CDNS_4066195314519_2/D PDRIVE_Y DVDD pfet_06v0 ad=3.12p pd=12.52u as=3.12p ps=12.52u w=11.999999u l=0.7u
X1 NDRIVE_Y SL NDRIVE_X DVDD pfet_06v0 ad=5.28p pd=24.88u as=3.12p ps=12.52u w=11.999999u l=0.7u
X2 nmos_6p0_CDNS_4066195314519_2/S A DVDD DVDD pfet_06v0 ad=5.28p pd=24.88u as=3.12p ps=12.52u w=11.999999u l=0.7u
X3 DVDD nmos_6p0_CDNS_4066195314519_2/S NDRIVE_Y DVDD pfet_06v0 ad=3.12p pd=12.52u as=5.28p ps=24.88u w=11.999999u l=0.7u
X4 PDRIVE_X nmos_6p0_CDNS_4066195314519_2/D DVDD DVDD pfet_06v0 ad=3.12p pd=12.52u as=3.12p ps=12.52u w=11.999999u l=0.7u
X5 NDRIVE_Y nmos_6p0_CDNS_4066195314519_2/S DVDD DVDD pfet_06v0 ad=3.12p pd=12.52u as=3.12p ps=12.52u w=11.999999u l=0.7u
X6 nmos_6p0_CDNS_4066195314519_2/S ENB nmos_6p0_CDNS_4066195314519_2/D DVDD pfet_06v0 ad=3.12p pd=12.52u as=5.28p ps=24.88u w=11.999999u l=0.7u
X7 DVDD EN nmos_6p0_CDNS_4066195314519_2/S DVDD pfet_06v0 ad=3.12p pd=12.52u as=3.12p ps=12.52u w=11.999999u l=0.7u
X8 NDRIVE_Y DVSS NDRIVE_X DVDD pfet_06v0 ad=0.528p pd=3.28u as=0.528p ps=3.28u w=1.2u l=0.7u
X9 PDRIVE_Y nmos_6p0_CDNS_4066195314519_2/D DVDD DVDD pfet_06v0 ad=3.12p pd=12.52u as=5.28p ps=24.88u w=11.999999u l=0.7u
X10 DVDD nmos_6p0_CDNS_4066195314519_2/D PDRIVE_X DVDD pfet_06v0 ad=5.28p pd=24.88u as=3.12p ps=12.52u w=11.999999u l=0.7u
X11 NDRIVE_X SL NDRIVE_Y DVDD pfet_06v0 ad=3.12p pd=12.52u as=3.12p ps=12.52u w=11.999999u l=0.7u
.ends

.subckt nmos_6p0_CDNS_4066195314511 D a_0_n44# S VSUBS
X0 D a_0_n44# S VSUBS nfet_06v0 ad=1.32p pd=6.88u as=1.32p ps=6.88u w=3u l=0.7u
.ends

.subckt comp018green_out_sigbuf_a AB A OE VDD DVSS DVDD VSS
Xnmos_6p0_CDNS_4066195314511_0 AB nmos_6p0_CDNS_4066195314511_3/S DVSS nmos_6p0_CDNS_4066195314511_0/VSUBS
+ nmos_6p0_CDNS_4066195314511
Xnmos_6p0_CDNS_4066195314511_1 nmos_6p0_CDNS_4066195314511_1/D A nmos_6p0_CDNS_4066195314511_2/D
+ VSS nmos_6p0_CDNS_4066195314511
Xnmos_6p0_CDNS_4066195314511_2 nmos_6p0_CDNS_4066195314511_2/D OE VSS VSS nmos_6p0_CDNS_4066195314511
Xnmos_6p0_CDNS_4066195314511_3 DVSS nmos_6p0_CDNS_4066195314511_1/D nmos_6p0_CDNS_4066195314511_3/S
+ nmos_6p0_CDNS_4066195314511_3/VSUBS nmos_6p0_CDNS_4066195314511
X0 nmos_6p0_CDNS_4066195314511_1/D OE VDD VDD pfet_06v0 ad=0.78p pd=3.52u as=1.32p ps=6.88u w=3u l=0.7u
X1 AB nmos_6p0_CDNS_4066195314511_3/S DVDD DVDD pfet_06v0 ad=2.64p pd=12.879999u as=1.56p ps=6.52u w=6u l=0.7u
X2 VDD A nmos_6p0_CDNS_4066195314511_1/D VDD pfet_06v0 ad=1.32p pd=6.88u as=0.78p ps=3.52u w=3u l=0.7u
X3 DVDD nmos_6p0_CDNS_4066195314511_1/D nmos_6p0_CDNS_4066195314511_3/S DVDD pfet_06v0 ad=1.56p pd=6.52u as=2.64p ps=12.879999u w=6u l=0.7u
.ends

.subckt ppolyf_u_CDNS_4066195314551 PLUS MINUS VSUBS
X0 PLUS MINUS VSUBS ppolyf_u r_width=0.8u r_length=3.9u
.ends

.subckt pn_6p0_CDNS_4066195314510 PLUS MINUS
D0 PLUS MINUS diode_pd2nw_06v0 pj=1.92u area=0.2304p
.ends

.subckt comp018green_out_sigbuf_oe PDRV ENB DVDD OE EN VDD DVSS VSS
Xnmos_6p0_CDNS_4066195314511_0 VSS PDRV nmos_6p0_CDNS_4066195314511_1/D VSS nmos_6p0_CDNS_4066195314511
Xnmos_6p0_CDNS_4066195314511_1 nmos_6p0_CDNS_4066195314511_1/D OE nmos_6p0_CDNS_4066195314511_1/S
+ VSS nmos_6p0_CDNS_4066195314511
Xnmos_6p0_CDNS_4066195314511_2 ENB EN DVSS nmos_6p0_CDNS_4066195314511_2/VSUBS nmos_6p0_CDNS_4066195314511
Xnmos_6p0_CDNS_4066195314511_3 DVSS nmos_6p0_CDNS_4066195314511_1/S EN nmos_6p0_CDNS_4066195314511_3/VSUBS
+ nmos_6p0_CDNS_4066195314511
Xpn_6p0_CDNS_4066195314510_0 VSS PDRV pn_6p0_CDNS_4066195314510
Xpn_6p0_CDNS_4066195314510_1 VSS OE pn_6p0_CDNS_4066195314510
X0 DVDD nmos_6p0_CDNS_4066195314511_1/S EN DVDD pfet_06v0 ad=1.56p pd=6.52u as=2.64p ps=12.879999u w=6u l=0.7u
X1 nmos_6p0_CDNS_4066195314511_1/S PDRV VDD VDD pfet_06v0 ad=0.78p pd=3.52u as=1.32p ps=6.88u w=3u l=0.7u
X2 ENB EN DVDD DVDD pfet_06v0 ad=2.64p pd=12.879999u as=1.56p ps=6.52u w=6u l=0.7u
X3 VDD OE nmos_6p0_CDNS_4066195314511_1/S VDD pfet_06v0 ad=1.32p pd=6.88u as=0.78p ps=3.52u w=3u l=0.7u
.ends

.subckt ppolyf_u_CDNS_4066195314532 PLUS MINUS VSUBS
X0 PLUS MINUS VSUBS ppolyf_u r_width=0.8u r_length=22.999998u
.ends

.subckt ppolyf_u_CDNS_4066195314533 PLUS MINUS VSUBS
X0 PLUS MINUS VSUBS ppolyf_u r_width=0.8u r_length=35.7u
.ends

.subckt comp018green_in_pupd A DVDD DVSS PU_B PD w_n83_53# a_6234_n7404# VSUBS
Xppolyf_u_CDNS_4066195314532_0 A ppolyf_u_CDNS_4066195314533_2/PLUS VSUBS ppolyf_u_CDNS_4066195314532
Xppolyf_u_CDNS_4066195314533_0 ppolyf_u_CDNS_4066195314533_0/PLUS ppolyf_u_CDNS_4066195314533_3/PLUS
+ VSUBS ppolyf_u_CDNS_4066195314533
Xppolyf_u_CDNS_4066195314533_1 ppolyf_u_CDNS_4066195314533_1/PLUS ppolyf_u_CDNS_4066195314533_6/PLUS
+ VSUBS ppolyf_u_CDNS_4066195314533
Xppolyf_u_CDNS_4066195314533_2 ppolyf_u_CDNS_4066195314533_2/PLUS ppolyf_u_CDNS_4066195314533_1/PLUS
+ VSUBS ppolyf_u_CDNS_4066195314533
Xppolyf_u_CDNS_4066195314533_3 ppolyf_u_CDNS_4066195314533_3/PLUS ppolyf_u_CDNS_4066195314533_4/MINUS
+ VSUBS ppolyf_u_CDNS_4066195314533
Xppolyf_u_CDNS_4066195314533_4 ppolyf_u_CDNS_4066195314533_5/PLUS ppolyf_u_CDNS_4066195314533_4/MINUS
+ VSUBS ppolyf_u_CDNS_4066195314533
Xppolyf_u_CDNS_4066195314533_5 ppolyf_u_CDNS_4066195314533_5/PLUS nmos_6p0_CDNS_4066195314530_0/D
+ VSUBS ppolyf_u_CDNS_4066195314533
Xppolyf_u_CDNS_4066195314533_6 ppolyf_u_CDNS_4066195314533_6/PLUS ppolyf_u_CDNS_4066195314533_0/PLUS
+ VSUBS ppolyf_u_CDNS_4066195314533
Xnmos_6p0_CDNS_4066195314530_0 nmos_6p0_CDNS_4066195314530_0/D PD DVSS nmos_6p0_CDNS_4066195314530_0/VSUBS
+ nmos_6p0_CDNS_4066195314530
X0 DVDD a_6234_n7404# nmos_6p0_CDNS_4066195314530_0/D DVDD pfet_06v0 ad=1.32p pd=6.88u as=1.32p ps=6.88u w=3u l=0.7u
.ends

.subckt comp018green_std_xor2 B Z VDD VSS A
Xnmos_6p0_CDNS_4066195314530_2 nmos_6p0_CDNS_4066195314530_3/D B Z VSS nmos_6p0_CDNS_4066195314530
Xnmos_6p0_CDNS_4066195314530_3 nmos_6p0_CDNS_4066195314530_3/D A VSS VSS nmos_6p0_CDNS_4066195314530
Xnmos_6p0_CDNS_4066195314530_0 nmos_6p0_CDNS_4066195314530_0/D B VSS VSS nmos_6p0_CDNS_4066195314530
Xnmos_6p0_CDNS_4066195314530_1 A nmos_6p0_CDNS_4066195314530_0/D Z VSS nmos_6p0_CDNS_4066195314530
X0 nmos_6p0_CDNS_4066195314530_3/D nmos_6p0_CDNS_4066195314530_0/D Z VDD pfet_06v0 ad=1.32p pd=6.88u as=1.32p ps=6.88u w=3u l=0.7u
X1 VDD B nmos_6p0_CDNS_4066195314530_0/D VDD pfet_06v0 ad=1.32p pd=6.88u as=1.32p ps=6.88u w=3u l=0.7u
X2 nmos_6p0_CDNS_4066195314530_3/D A VDD VDD pfet_06v0 ad=1.32p pd=6.88u as=1.32p ps=6.88u w=3u l=0.7u
X3 Z B A VDD pfet_06v0 ad=1.32p pd=6.88u as=1.32p ps=6.88u w=3u l=0.7u
.ends

.subckt comp018green_std_nand2 VDD A B Z VSS
Xnmos_6p0_CDNS_4066195314511_0 nmos_6p0_CDNS_4066195314511_1/S A VSS VSS nmos_6p0_CDNS_4066195314511
Xnmos_6p0_CDNS_4066195314511_1 Z B nmos_6p0_CDNS_4066195314511_1/S VSS nmos_6p0_CDNS_4066195314511
X0 VDD B Z VDD pfet_06v0 ad=1.32p pd=6.88u as=0.78p ps=3.52u w=3u l=0.7u
X1 Z A VDD VDD pfet_06v0 ad=0.78p pd=3.52u as=1.32p ps=6.88u w=3u l=0.7u
.ends

.subckt comp018green_in_logic_pupd PDB_OUT VDD comp018green_std_nand2_1/VDD comp018green_std_xor2_0/A
+ PUB_OUT PD_IN VSS
Xcomp018green_std_xor2_0 PD_IN comp018green_std_xor2_0/Z VDD VSS comp018green_std_xor2_0/A
+ comp018green_std_xor2
Xcomp018green_std_nand2_0 comp018green_std_nand2_1/VDD comp018green_std_xor2_0/Z PD_IN
+ PDB_OUT VSS comp018green_std_nand2
Xcomp018green_std_nand2_1 comp018green_std_nand2_1/VDD comp018green_std_xor2_0/A comp018green_std_xor2_0/Z
+ PUB_OUT VSS comp018green_std_nand2
.ends

.subckt comp018green_sigbuf Z VSS DVDD A ZB VDD DVSS
Xnmos_6p0_CDNS_4066195314531_0 ZB Z DVSS Z nmos_6p0_CDNS_4066195314531
Xnmos_6p0_CDNS_4066195314531_1 Z nmos_6p0_CDNS_4066195314530_0/D DVSS nmos_6p0_CDNS_4066195314530_0/D
+ nmos_6p0_CDNS_4066195314531
Xnmos_6p0_CDNS_4066195314530_0 nmos_6p0_CDNS_4066195314530_0/D A VSS VSS nmos_6p0_CDNS_4066195314530
X0 DVDD Z ZB DVDD pfet_06v0 ad=1.32p pd=6.88u as=0.78p ps=3.52u w=3u l=0.7u
X1 nmos_6p0_CDNS_4066195314530_0/D A VDD VDD pfet_06v0 ad=1.32p pd=6.88u as=1.32p ps=6.88u w=3u l=0.7u
X2 ZB Z DVDD DVDD pfet_06v0 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.7u
X3 Z nmos_6p0_CDNS_4066195314530_0/D DVDD DVDD pfet_06v0 ad=0.78p pd=3.52u as=1.32p ps=6.88u w=3u l=0.7u
X4 DVDD nmos_6p0_CDNS_4066195314530_0/D Z DVDD pfet_06v0 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.7u
.ends

.subckt nmos_6p0_CDNS_4066195314549 D a_732_n44# a_976_n44# a_0_n44# S a_1220_n44#
+ a_244_n44# a_488_n44# VSUBS
X0 D a_976_n44# S VSUBS nfet_06v0 ad=0.39p pd=2.02u as=0.39p ps=2.02u w=1.5u l=0.7u
X1 S a_732_n44# D VSUBS nfet_06v0 ad=0.39p pd=2.02u as=0.39p ps=2.02u w=1.5u l=0.7u
X2 S a_1220_n44# D VSUBS nfet_06v0 ad=0.66p pd=3.88u as=0.39p ps=2.02u w=1.5u l=0.7u
X3 S a_244_n44# D VSUBS nfet_06v0 ad=0.39p pd=2.02u as=0.39p ps=2.02u w=1.5u l=0.7u
X4 D a_488_n44# S VSUBS nfet_06v0 ad=0.39p pd=2.02u as=0.39p ps=2.02u w=1.5u l=0.7u
X5 D a_0_n44# S VSUBS nfet_06v0 ad=0.39p pd=2.02u as=0.66p ps=3.88u w=1.5u l=0.7u
.ends

.subckt nmos_6p0_CDNS_4066195314547 D a_0_n44# S a_244_n44#
X0 S a_244_n44# D VSUBS nfet_06v0 ad=1.76p pd=8.88u as=1.04p ps=4.52u w=4u l=0.7u
X1 D a_0_n44# S VSUBS nfet_06v0 ad=1.04p pd=4.52u as=1.76p ps=8.88u w=4u l=0.7u
.ends

.subckt nmos_6p0_CDNS_4066195314550 D a_0_n44# S a_244_n44# VSUBS
X0 S a_244_n44# D VSUBS nfet_06v0 ad=0.55p pd=3.38u as=0.325p ps=1.77u w=1.25u l=0.7u
X1 D a_0_n44# S VSUBS nfet_06v0 ad=0.325p pd=1.77u as=0.55p ps=3.38u w=1.25u l=0.7u
.ends

.subckt comp018green_in_drv DVDD A VDD Z DVSS nmos_6p0_CDNS_4066195314549_0/D VSS
Xnmos_6p0_CDNS_4066195314549_0 nmos_6p0_CDNS_4066195314549_0/D Z Z Z VSS Z Z Z VSS
+ nmos_6p0_CDNS_4066195314549
Xnmos_6p0_CDNS_4066195314547_0 DVSS A nmos_6p0_CDNS_4066195314547_0/S A nmos_6p0_CDNS_4066195314547
Xnmos_6p0_CDNS_4066195314550_0 Z nmos_6p0_CDNS_4066195314547_0/S VSS nmos_6p0_CDNS_4066195314547_0/S
+ VSS nmos_6p0_CDNS_4066195314550
X0 VDD nmos_6p0_CDNS_4066195314547_0/S Z VDD pfet_06v0 ad=1.1p pd=5.88u as=0.65p ps=3.02u w=2.5u l=0.7u
X1 VDD Z nmos_6p0_CDNS_4066195314549_0/D VDD pfet_06v0 ad=1.54p pd=7.88u as=0.91p ps=4.02u w=3.5u l=0.7u
X2 VDD nmos_6p0_CDNS_4066195314547_0/S Z VDD pfet_06v0 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.7u
X3 nmos_6p0_CDNS_4066195314549_0/D Z VDD VDD pfet_06v0 ad=0.91p pd=4.02u as=0.91p ps=4.02u w=3.5u l=0.7u
X4 nmos_6p0_CDNS_4066195314549_0/D Z VDD VDD pfet_06v0 ad=0.91p pd=4.02u as=1.54p ps=7.88u w=3.5u l=0.7u
X5 Z nmos_6p0_CDNS_4066195314547_0/S VDD VDD pfet_06v0 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.7u
X6 VDD Z nmos_6p0_CDNS_4066195314549_0/D VDD pfet_06v0 ad=0.91p pd=4.02u as=0.91p ps=4.02u w=3.5u l=0.7u
X7 nmos_6p0_CDNS_4066195314547_0/S A DVDD DVDD pfet_06v0 ad=0.88p pd=4.88u as=0.88p ps=4.88u w=2u l=0.7u
X8 VDD Z nmos_6p0_CDNS_4066195314549_0/D VDD pfet_06v0 ad=0.91p pd=4.02u as=0.91p ps=4.02u w=3.5u l=0.7u
X9 nmos_6p0_CDNS_4066195314549_0/D Z VDD VDD pfet_06v0 ad=0.91p pd=4.02u as=0.91p ps=4.02u w=3.5u l=0.7u
X10 Z nmos_6p0_CDNS_4066195314547_0/S VDD VDD pfet_06v0 ad=0.65p pd=3.02u as=1.1p ps=5.88u w=2.5u l=0.7u
.ends

.subckt nmos_6p0_CDNS_4066195314537 D a_732_n44# a_976_n44# a_0_n44# S a_244_n44#
+ a_488_n44#
X0 D a_976_n44# S VSUBS nfet_06v0 ad=1.408p pd=7.28u as=0.832p ps=3.72u w=3.2u l=0.7u
X1 S a_732_n44# D VSUBS nfet_06v0 ad=0.832p pd=3.72u as=0.832p ps=3.72u w=3.2u l=0.7u
X2 S a_244_n44# D VSUBS nfet_06v0 ad=0.832p pd=3.72u as=0.832p ps=3.72u w=3.2u l=0.7u
X3 D a_488_n44# S VSUBS nfet_06v0 ad=0.832p pd=3.72u as=0.832p ps=3.72u w=3.2u l=0.7u
X4 D a_0_n44# S VSUBS nfet_06v0 ad=0.832p pd=3.72u as=1.408p ps=7.28u w=3.2u l=0.7u
.ends

.subckt nmos_6p0_CDNS_4066195314542 D a_732_n44# a_0_n44# S a_244_n44# a_488_n44#
X0 D a_732_n44# S VSUBS nfet_06v0 ad=1.32p pd=6.88u as=0.78p ps=3.52u w=3u l=0.7u
X1 D a_244_n44# S VSUBS nfet_06v0 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.7u
X2 S a_488_n44# D VSUBS nfet_06v0 ad=0.78p pd=3.52u as=0.78p ps=3.52u w=3u l=0.7u
X3 S a_0_n44# D VSUBS nfet_06v0 ad=0.78p pd=3.52u as=1.32p ps=6.88u w=3u l=0.7u
.ends

.subckt nmos_6p0_CDNS_4066195314535 D a_0_n44# S a_244_n44#
X0 S a_244_n44# D VSUBS nfet_06v0 ad=0.88p pd=4.88u as=0.52p ps=2.52u w=2u l=0.7u
X1 D a_0_n44# S VSUBS nfet_06v0 ad=0.52p pd=2.52u as=0.88p ps=4.88u w=2u l=0.7u
.ends

.subckt nmos_6p0_CDNS_4066195314540 D a_0_n44# S
X0 S a_0_n44# D VSUBS nfet_06v0 ad=0.572p pd=3.48u as=0.572p ps=3.48u w=1.3u l=0.7u
.ends

.subckt nmos_6p0_CDNS_4066195314536 D a_0_n44# S
X0 D a_0_n44# S VSUBS nfet_06v0 ad=0.66p pd=3.88u as=0.66p ps=3.88u w=1.5u l=0.7u
.ends

.subckt nmos_6p0_CDNS_4066195314541 D a_732_n44# a_0_n44# S a_244_n44# a_488_n44#
X0 S a_732_n44# D VSUBS nfet_06v0 ad=1.166p pd=6.18u as=0.689p ps=3.17u w=2.65u l=0.7u
X1 S a_244_n44# D VSUBS nfet_06v0 ad=0.689p pd=3.17u as=0.689p ps=3.17u w=2.65u l=0.7u
X2 D a_488_n44# S VSUBS nfet_06v0 ad=0.689p pd=3.17u as=0.689p ps=3.17u w=2.65u l=0.7u
X3 D a_0_n44# S VSUBS nfet_06v0 ad=0.689p pd=3.17u as=1.166p ps=6.18u w=2.65u l=0.7u
.ends

.subckt comp018green_in_cms_smt IE CS A Z nmos_6p0_CDNS_4066195314540_0/D m2_5364_1052#
+ a_459_724# DVSS DVDD
Xnmos_6p0_CDNS_4066195314537_0 nmos_6p0_CDNS_4066195314541_0/D IE IE IE DVSS IE IE
+ nmos_6p0_CDNS_4066195314537
Xnmos_6p0_CDNS_4066195314542_0 nmos_6p0_CDNS_4066195314542_0/D A A Z A A nmos_6p0_CDNS_4066195314542
Xnmos_6p0_CDNS_4066195314535_0 nmos_6p0_CDNS_4066195314535_0/D a_459_724# DVSS a_459_724#
+ nmos_6p0_CDNS_4066195314535
Xnmos_6p0_CDNS_4066195314540_0 nmos_6p0_CDNS_4066195314540_0/D nmos_6p0_CDNS_4066195314536_0/D
+ nmos_6p0_CDNS_4066195314542_0/D nmos_6p0_CDNS_4066195314540
Xnmos_6p0_CDNS_4066195314536_1 Z CS nmos_6p0_CDNS_4066195314536_1/S nmos_6p0_CDNS_4066195314536
Xnmos_6p0_CDNS_4066195314536_0 nmos_6p0_CDNS_4066195314536_0/D nmos_6p0_CDNS_4066195314535_0/D
+ DVSS nmos_6p0_CDNS_4066195314536
Xnmos_6p0_CDNS_4066195314541_0 nmos_6p0_CDNS_4066195314541_0/D A A nmos_6p0_CDNS_4066195314542_0/D
+ A A nmos_6p0_CDNS_4066195314541
Xnmos_6p0_CDNS_4066195314530_0 nmos_6p0_CDNS_4066195314536_0/D CS Z nmos_6p0_CDNS_4066195314530_0/VSUBS
+ nmos_6p0_CDNS_4066195314530
X0 DVSS nmos_6p0_CDNS_4066195314536_1/S a_3227_1730# DVDD pfet_06v0 ad=0.494p pd=2.42u as=0.836p ps=4.68u w=1.9u l=0.7u
X1 Z IE DVDD DVDD pfet_06v0 ad=0.88p pd=4.88u as=0.52p ps=2.52u w=2u l=0.7u
X2 Z nmos_6p0_CDNS_4066195314535_0/D nmos_6p0_CDNS_4066195314536_1/S DVDD pfet_06v0 ad=0.88p pd=4.88u as=0.88p ps=4.88u w=2u l=0.7u
X3 DVDD CS nmos_6p0_CDNS_4066195314536_1/S DVDD pfet_06v0 ad=0.66p pd=3.88u as=0.39p ps=2.02u w=1.5u l=0.7u
X4 Z A a_3227_1730# DVDD pfet_06v0 ad=0.559p pd=2.67u as=0.946p ps=5.18u w=2.15u l=0.7u
X5 a_3227_1730# A Z DVDD pfet_06v0 ad=0.946p pd=5.18u as=0.559p ps=2.67u w=2.15u l=0.7u
X6 DVDD A a_3227_1730# DVDD pfet_06v0 ad=0.494p pd=2.42u as=0.836p ps=4.68u w=1.9u l=0.7u
X7 nmos_6p0_CDNS_4066195314535_0/D a_459_724# DVDD DVDD pfet_06v0 ad=1.04p pd=4.52u as=1.76p ps=8.88u w=4u l=0.7u
X8 Z IE DVDD DVDD pfet_06v0 ad=0.52p pd=2.52u as=0.88p ps=4.88u w=2u l=0.7u
X9 DVDD IE Z DVDD pfet_06v0 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=0.7u
X10 a_3227_1730# A DVDD DVDD pfet_06v0 ad=0.836p pd=4.68u as=0.494p ps=2.42u w=1.9u l=0.7u
X11 a_3227_1730# nmos_6p0_CDNS_4066195314536_1/S DVSS DVDD pfet_06v0 ad=0.836p pd=4.68u as=0.494p ps=2.42u w=1.9u l=0.7u
X12 DVDD a_459_724# nmos_6p0_CDNS_4066195314535_0/D DVDD pfet_06v0 ad=1.76p pd=8.88u as=1.04p ps=4.52u w=4u l=0.7u
X13 nmos_6p0_CDNS_4066195314536_1/S CS DVDD DVDD pfet_06v0 ad=0.39p pd=2.02u as=0.66p ps=3.88u w=1.5u l=0.7u
X14 nmos_6p0_CDNS_4066195314536_0/D nmos_6p0_CDNS_4066195314535_0/D Z DVDD pfet_06v0 ad=0.88p pd=4.88u as=0.88p ps=4.88u w=2u l=0.7u
.ends

.subckt pn_6p0_CDNS_4066195314528 PLUS MINUS
D0 PLUS MINUS diode_pd2nw_06v0 pj=4u area=1p
.ends

.subckt comp018green_inpath_cms_smt PAD IE CS PD PU VDD comp018green_in_pupd_0/w_n83_53#
+ comp018green_in_pupd_0/A comp018green_in_pupd_0/DVDD comp018green_in_pupd_0/DVSS
+ comp018green_in_cms_smt_0/nmos_6p0_CDNS_4066195314540_0/D comp018green_sigbuf_2/VDD
+ comp018green_sigbuf_3/DVDD comp018green_in_drv_0/nmos_6p0_CDNS_4066195314549_0/D
+ comp018green_sigbuf_1/VDD comp018green_in_logic_pupd_0/VDD comp018green_in_drv_0/DVDD
+ comp018green_sigbuf_3/VDD comp018green_sigbuf_3/DVSS comp018green_in_drv_0/DVSS
+ comp018green_sigbuf_2/DVDD VSUBS comp018green_in_logic_pupd_0/comp018green_std_nand2_1/VDD
+ comp018green_sigbuf_2/DVSS
Xcomp018green_in_pupd_0 comp018green_in_pupd_0/A comp018green_in_pupd_0/DVDD comp018green_in_pupd_0/DVSS
+ comp018green_in_pupd_0/PU_B comp018green_sigbuf_0/ZB comp018green_in_pupd_0/w_n83_53#
+ comp018green_sigbuf_2/Z VSUBS comp018green_in_pupd
Xcomp018green_in_logic_pupd_0 comp018green_sigbuf_0/A comp018green_in_logic_pupd_0/VDD
+ comp018green_in_logic_pupd_0/comp018green_std_nand2_1/VDD PU comp018green_sigbuf_2/A
+ PD VSUBS comp018green_in_logic_pupd
Xcomp018green_sigbuf_0 comp018green_sigbuf_0/Z VSUBS comp018green_sigbuf_2/DVDD comp018green_sigbuf_0/A
+ comp018green_sigbuf_0/ZB comp018green_sigbuf_3/VDD comp018green_sigbuf_2/DVSS comp018green_sigbuf
Xcomp018green_sigbuf_1 comp018green_sigbuf_1/Z VSUBS comp018green_sigbuf_3/DVDD IE
+ comp018green_sigbuf_1/ZB comp018green_sigbuf_1/VDD comp018green_sigbuf_3/DVSS comp018green_sigbuf
Xcomp018green_sigbuf_2 comp018green_sigbuf_2/Z VSUBS comp018green_sigbuf_2/DVDD comp018green_sigbuf_2/A
+ comp018green_sigbuf_2/ZB comp018green_sigbuf_2/VDD comp018green_sigbuf_2/DVSS comp018green_sigbuf
Xcomp018green_sigbuf_3 comp018green_sigbuf_3/Z VSUBS comp018green_sigbuf_3/DVDD CS
+ comp018green_sigbuf_3/ZB comp018green_sigbuf_3/VDD comp018green_sigbuf_3/DVSS comp018green_sigbuf
Xcomp018green_in_drv_0 comp018green_in_drv_0/DVDD comp018green_in_drv_0/A VDD comp018green_in_drv_0/Z
+ comp018green_in_drv_0/DVSS comp018green_in_drv_0/nmos_6p0_CDNS_4066195314549_0/D
+ VSUBS comp018green_in_drv
Xcomp018green_in_cms_smt_0 comp018green_sigbuf_1/Z comp018green_sigbuf_3/Z PAD comp018green_in_drv_0/A
+ comp018green_in_cms_smt_0/nmos_6p0_CDNS_4066195314540_0/D PAD comp018green_sigbuf_3/Z
+ comp018green_in_drv_0/DVSS comp018green_in_drv_0/DVDD comp018green_in_cms_smt
Xpn_6p0_CDNS_4066195314528_0 PD comp018green_sigbuf_1/VDD pn_6p0_CDNS_4066195314528
Xpn_6p0_CDNS_4066195314528_1 CS comp018green_sigbuf_1/VDD pn_6p0_CDNS_4066195314528
Xpn_6p0_CDNS_4066195314528_2 IE comp018green_sigbuf_1/VDD pn_6p0_CDNS_4066195314528
Xpn_6p0_CDNS_4066195314528_3 PU comp018green_sigbuf_1/VDD pn_6p0_CDNS_4066195314528
.ends

.subckt nmoscap_6p0_CDNS_4066195314522 G D
X0 G D cap_nmos_06v0 c_width=3u c_length=3u
.ends

.subckt np_6p0_CDNS_4066195314526 MINUS
D0 VSUBS MINUS diode_nd2ps_06v0 pj=42u area=20p
.ends

.subckt ppolyf_u_CDNS_4066195314525 PLUS MINUS
X0 PLUS MINUS VSUBS ppolyf_u r_width=2.5u r_length=2.8u
.ends

.subckt pn_6p0_CDNS_4066195314527 w_n120_n120# PLUS
D0 PLUS w_n120_n120# diode_pd2nw_06v0 pj=42u area=20p
.ends

.subckt comp018green_esd_cdm PAD w_n83_n83# DVSS w_454_3720# IP_IN m1_379_11# DVDD
Xnp_6p0_CDNS_4066195314526_1 IP_IN np_6p0_CDNS_4066195314526
Xppolyf_u_CDNS_4066195314525_0 PAD IP_IN ppolyf_u_CDNS_4066195314525
Xppolyf_u_CDNS_4066195314525_1 PAD IP_IN ppolyf_u_CDNS_4066195314525
Xppolyf_u_CDNS_4066195314525_2 PAD IP_IN ppolyf_u_CDNS_4066195314525
Xppolyf_u_CDNS_4066195314525_3 PAD IP_IN ppolyf_u_CDNS_4066195314525
Xpn_6p0_CDNS_4066195314527_0 w_454_3720# IP_IN pn_6p0_CDNS_4066195314527
Xpn_6p0_CDNS_4066195314527_1 w_454_3720# IP_IN pn_6p0_CDNS_4066195314527
Xnp_6p0_CDNS_4066195314526_0 IP_IN np_6p0_CDNS_4066195314526
.ends

.subckt GF_NI_IN_C_BASE pdrive_x_<3> pdrive_y_<3> pdrive_y_<2> pdrive_x_<2> pdrive_x_<1>
+ pdrive_y_<1> pdrive_y_<0> pdrive_x_<0> ndrive_Y_<3> ndrive_x_<3> ndrive_y_<2> ndrive_x_<2>
+ ndrive_Y_<1> ndrive_x_<1> ndrive_y_<0> ndrive_x_<0> Y PU PD comp018green_out_sigbuf_oe_1/DVDD
+ m2_1886_53031# PAD comp018green_out_sigbuf_oe_0/VDD comp018green_out_paddrv_16T_0/comp018green_out_paddrv_4T_NMOS_GROUP_0/nmos_4T_metal_stack_2/m2_n44_400#
+ comp018green_out_paddrv_16T_0/comp018green_out_paddrv_4T_NMOS_GROUP_0/nmos_4T_metal_stack_3/m2_n44_400#
+ comp018green_out_paddrv_16T_0/comp018green_out_paddrv_4T_PMOS_GROUP_0/PMOS_4T_metal_stack_1/m2_n44_0#
+ comp018green_out_paddrv_16T_0/comp018green_out_paddrv_4T_PMOS_GROUP_0/PMOS_4T_metal_stack_2/m2_n44_0#
+ comp018green_out_paddrv_16T_0/comp018green_out_paddrv_4T_NMOS_GROUP_0/nmos_4T_metal_stack_1/m2_n44_400#
+ comp018green_sigbuf_1_0/VDD comp018green_out_paddrv_16T_0/comp018green_out_paddrv_4T_PMOS_GROUP_0/PMOS_4T_metal_stack_3/m2_n44_0#
+ comp018green_out_sigbuf_oe_2/VDD comp018green_out_paddrv_16T_0/comp018green_out_paddrv_4T_PMOS_GROUP_0/PMOS_4T_metal_stack_5/m2_n44_0#
+ comp018green_out_sigbuf_a_0/DVDD comp018green_inpath_cms_smt_0/comp018green_in_logic_pupd_0/VDD
+ comp018green_out_paddrv_16T_0/comp018green_out_paddrv_4T_PMOS_GROUP_0/PMOS_4T_metal_stack_4/m2_n44_0#
+ comp018green_esd_cdm_0/DVDD comp018green_inpath_cms_smt_0/comp018green_in_pupd_0/DVDD
+ comp018green_inpath_cms_smt_0/VDD M3_M2_CDNS_40661953145188_0/m2_n961_n38# comp018green_esd_cdm_0/w_454_3720#
+ nmoscap_6p0_CDNS_4066195314522_3/G comp018green_out_paddrv_16T_0/comp018green_out_paddrv_4T_NMOS_GROUP_0/VSUBS
+ nmoscap_6p0_CDNS_4066195314523_7/D comp018green_out_predrv_3/DVDD comp018green_inpath_cms_smt_0/comp018green_in_drv_0/DVDD
+ comp018green_inpath_cms_smt_0/comp018green_sigbuf_2/DVDD VSUBS comp018green_sigbuf_1_0/DVSS
+ comp018green_sigbuf_1_0/DVDD comp018green_esd_cdm_0/DVSS comp018green_out_paddrv_16T_0/comp018green_out_paddrv_4T_PMOS_GROUP_0/w_n2_111#
+ comp018green_inpath_cms_smt_0/comp018green_sigbuf_3/DVDD
Xnmoscap_6p0_CDNS_4066195314523_7 comp018green_out_predrv_3/DVDD nmoscap_6p0_CDNS_4066195314523_7/D
+ nmoscap_6p0_CDNS_4066195314523
Xcomp018green_out_paddrv_16T_0 pdrive_x_<2> pdrive_x_<3> pdrive_y_<3> pdrive_x_<3>
+ ndrive_Y_<3> pdrive_x_<0> pdrive_x_<2> pdrive_y_<0> ndrive_x_<0> ndrive_y_<2> pdrive_y_<2>
+ pdrive_x_<1> ndrive_x_<3> pdrive_y_<1> ndrive_x_<1> ndrive_y_<0> pdrive_x_<0> ndrive_x_<2>
+ comp018green_out_paddrv_16T_0/comp018green_out_paddrv_4T_NMOS_GROUP_0/nmos_4T_metal_stack_2/m2_n44_400#
+ pdrive_x_<1> comp018green_out_paddrv_16T_0/comp018green_out_paddrv_4T_NMOS_GROUP_0/nmos_4T_metal_stack_3/m2_n44_400#
+ PAD comp018green_out_paddrv_16T_0/comp018green_out_paddrv_4T_PMOS_GROUP_0/PMOS_4T_metal_stack_5/m2_n44_0#
+ comp018green_out_paddrv_16T_0/comp018green_out_paddrv_4T_PMOS_GROUP_0/w_n2_111#
+ ndrive_Y_<1> comp018green_out_paddrv_16T_0/comp018green_out_paddrv_4T_NMOS_GROUP_0/nmos_4T_metal_stack_1/m2_n44_400#
+ comp018green_out_predrv_3/DVDD comp018green_out_paddrv_16T_0/comp018green_out_paddrv_4T_PMOS_GROUP_0/PMOS_4T_metal_stack_1/m2_n44_0#
+ comp018green_out_paddrv_16T_0/comp018green_out_paddrv_4T_PMOS_GROUP_0/PMOS_4T_metal_stack_4/m2_n44_0#
+ comp018green_out_paddrv_16T_0/comp018green_out_paddrv_4T_PMOS_GROUP_0/PMOS_4T_metal_stack_2/m2_n44_0#
+ comp018green_out_paddrv_16T_0/comp018green_out_paddrv_4T_NMOS_GROUP_0/VSUBS comp018green_out_paddrv_16T_0/comp018green_out_paddrv_4T_PMOS_GROUP_0/PMOS_4T_metal_stack_3/m2_n44_0#
+ comp018green_out_paddrv_16T
Xcomp018green_sigbuf_1_0 comp018green_sigbuf_1_0/Z VSUBS comp018green_sigbuf_1_0/A
+ comp018green_sigbuf_1_0/VDD comp018green_sigbuf_1_0/ZB comp018green_sigbuf_1_0/DVSS
+ comp018green_sigbuf_1_0/DVDD comp018green_sigbuf_1
Xcomp018green_out_predrv_0 comp018green_sigbuf_1_0/Z comp018green_sigbuf_1_0/ZB ndrive_x_<0>
+ comp018green_out_predrv_0/ENB comp018green_out_predrv_3/A ndrive_y_<0> pdrive_y_<0>
+ pdrive_x_<0> comp018green_out_predrv_0/EN comp018green_out_predrv_3/DVDD comp018green_sigbuf_1_0/DVSS
+ comp018green_out_predrv
Xcomp018green_out_predrv_1 comp018green_sigbuf_1_0/Z comp018green_sigbuf_1_0/ZB ndrive_x_<3>
+ comp018green_out_predrv_1/ENB comp018green_out_predrv_3/A ndrive_Y_<3> pdrive_y_<3>
+ pdrive_x_<3> comp018green_out_predrv_1/EN comp018green_out_predrv_3/DVDD comp018green_sigbuf_1_0/DVSS
+ comp018green_out_predrv
Xcomp018green_out_sigbuf_a_0 comp018green_out_predrv_3/A comp018green_sigbuf_1_0/A
+ comp018green_sigbuf_1_0/A comp018green_sigbuf_1_0/VDD comp018green_sigbuf_1_0/DVSS
+ comp018green_out_sigbuf_a_0/DVDD VSUBS comp018green_out_sigbuf_a
Xppolyf_u_CDNS_4066195314551_0 comp018green_out_sigbuf_oe_0/VDD comp018green_inpath_cms_smt_0/IE
+ VSUBS ppolyf_u_CDNS_4066195314551
Xcomp018green_out_predrv_2 comp018green_sigbuf_1_0/Z comp018green_sigbuf_1_0/ZB ndrive_x_<2>
+ comp018green_out_predrv_3/ENB comp018green_out_predrv_3/A ndrive_y_<2> pdrive_y_<2>
+ pdrive_x_<2> comp018green_out_predrv_3/EN comp018green_out_predrv_3/DVDD comp018green_sigbuf_1_0/DVSS
+ comp018green_out_predrv
Xcomp018green_out_sigbuf_oe_0 comp018green_sigbuf_1_0/A comp018green_out_predrv_0/ENB
+ comp018green_out_sigbuf_oe_1/DVDD comp018green_sigbuf_1_0/A comp018green_out_predrv_0/EN
+ comp018green_out_sigbuf_oe_0/VDD comp018green_sigbuf_1_0/DVSS VSUBS comp018green_out_sigbuf_oe
Xppolyf_u_CDNS_4066195314551_1 VSUBS comp018green_sigbuf_1_0/A VSUBS ppolyf_u_CDNS_4066195314551
Xcomp018green_out_predrv_3 comp018green_sigbuf_1_0/Z comp018green_sigbuf_1_0/ZB ndrive_x_<1>
+ comp018green_out_predrv_3/ENB comp018green_out_predrv_3/A ndrive_Y_<1> pdrive_y_<1>
+ pdrive_x_<1> comp018green_out_predrv_3/EN comp018green_out_predrv_3/DVDD comp018green_sigbuf_1_0/DVSS
+ comp018green_out_predrv
Xcomp018green_out_sigbuf_oe_1 comp018green_sigbuf_1_0/A comp018green_out_predrv_3/ENB
+ comp018green_out_sigbuf_oe_1/DVDD comp018green_sigbuf_1_0/A comp018green_out_predrv_3/EN
+ comp018green_out_sigbuf_oe_2/VDD comp018green_sigbuf_1_0/DVSS VSUBS comp018green_out_sigbuf_oe
Xcomp018green_inpath_cms_smt_0 comp018green_esd_cdm_0/IP_IN comp018green_inpath_cms_smt_0/IE
+ comp018green_sigbuf_1_0/A PD PU comp018green_inpath_cms_smt_0/VDD M3_M2_CDNS_40661953145188_0/m2_n961_n38#
+ comp018green_esd_cdm_0/IP_IN comp018green_inpath_cms_smt_0/comp018green_in_pupd_0/DVDD
+ comp018green_esd_cdm_0/DVSS comp018green_inpath_cms_smt_0/comp018green_in_drv_0/DVDD
+ comp018green_out_sigbuf_oe_0/VDD comp018green_inpath_cms_smt_0/comp018green_sigbuf_3/DVDD
+ Y comp018green_out_sigbuf_oe_0/VDD comp018green_inpath_cms_smt_0/comp018green_in_logic_pupd_0/VDD
+ comp018green_inpath_cms_smt_0/comp018green_in_drv_0/DVDD comp018green_out_sigbuf_oe_0/VDD
+ nmoscap_6p0_CDNS_4066195314523_7/D nmoscap_6p0_CDNS_4066195314523_7/D comp018green_inpath_cms_smt_0/comp018green_sigbuf_2/DVDD
+ VSUBS comp018green_inpath_cms_smt_0/comp018green_in_logic_pupd_0/VDD nmoscap_6p0_CDNS_4066195314523_7/D
+ comp018green_inpath_cms_smt
Xcomp018green_out_sigbuf_oe_2 comp018green_out_sigbuf_oe_2/VDD comp018green_out_predrv_1/ENB
+ comp018green_out_sigbuf_a_0/DVDD comp018green_sigbuf_1_0/A comp018green_out_predrv_1/EN
+ comp018green_out_sigbuf_oe_2/VDD comp018green_sigbuf_1_0/DVSS VSUBS comp018green_out_sigbuf_oe
Xnmoscap_6p0_CDNS_4066195314522_0 nmoscap_6p0_CDNS_4066195314522_3/G comp018green_esd_cdm_0/DVSS
+ nmoscap_6p0_CDNS_4066195314522
Xnmoscap_6p0_CDNS_4066195314522_1 nmoscap_6p0_CDNS_4066195314522_3/G comp018green_esd_cdm_0/DVSS
+ nmoscap_6p0_CDNS_4066195314522
Xnmoscap_6p0_CDNS_4066195314522_2 nmoscap_6p0_CDNS_4066195314522_3/G comp018green_esd_cdm_0/DVSS
+ nmoscap_6p0_CDNS_4066195314522
Xnmoscap_6p0_CDNS_4066195314522_3 nmoscap_6p0_CDNS_4066195314522_3/G comp018green_esd_cdm_0/DVSS
+ nmoscap_6p0_CDNS_4066195314522
Xnmoscap_6p0_CDNS_4066195314523_0 comp018green_out_predrv_3/DVDD nmoscap_6p0_CDNS_4066195314523_7/D
+ nmoscap_6p0_CDNS_4066195314523
Xnmoscap_6p0_CDNS_4066195314523_1 comp018green_out_predrv_3/DVDD nmoscap_6p0_CDNS_4066195314523_7/D
+ nmoscap_6p0_CDNS_4066195314523
Xnmoscap_6p0_CDNS_4066195314523_2 comp018green_out_predrv_3/DVDD nmoscap_6p0_CDNS_4066195314523_7/D
+ nmoscap_6p0_CDNS_4066195314523
Xnmoscap_6p0_CDNS_4066195314523_3 comp018green_out_predrv_3/DVDD nmoscap_6p0_CDNS_4066195314523_7/D
+ nmoscap_6p0_CDNS_4066195314523
Xpn_6p0_CDNS_4066195314528_0 comp018green_sigbuf_1_0/A comp018green_sigbuf_1_0/VDD
+ pn_6p0_CDNS_4066195314528
Xnmoscap_6p0_CDNS_4066195314523_4 comp018green_out_predrv_3/DVDD nmoscap_6p0_CDNS_4066195314523_7/D
+ nmoscap_6p0_CDNS_4066195314523
Xcomp018green_esd_cdm_0 PAD comp018green_inpath_cms_smt_0/comp018green_in_pupd_0/DVDD
+ comp018green_esd_cdm_0/DVSS comp018green_esd_cdm_0/w_454_3720# comp018green_esd_cdm_0/IP_IN
+ comp018green_inpath_cms_smt_0/comp018green_in_drv_0/DVDD comp018green_esd_cdm_0/DVDD
+ comp018green_esd_cdm
Xpn_6p0_CDNS_4066195314528_1 comp018green_sigbuf_1_0/A comp018green_sigbuf_1_0/VDD
+ pn_6p0_CDNS_4066195314528
Xnmoscap_6p0_CDNS_4066195314523_5 comp018green_out_predrv_3/DVDD nmoscap_6p0_CDNS_4066195314523_7/D
+ nmoscap_6p0_CDNS_4066195314523
Xnmoscap_6p0_CDNS_4066195314523_6 comp018green_out_predrv_3/DVDD nmoscap_6p0_CDNS_4066195314523_7/D
+ nmoscap_6p0_CDNS_4066195314523
.ends

.subckt gf180mcu_fd_io__in_c VSS VDD DVSS DVDD PAD PU PD Y
X5LM_METAL_RAIL_PAD_60_0 GF_NI_IN_C_BASE_0/PAD VSS VDD DVSS DVDD VSS x5LM_METAL_RAIL_PAD_60
XGF_NI_IN_C_BASE_0 GF_NI_IN_C_BASE_0/pdrive_x_<3> GF_NI_IN_C_BASE_0/pdrive_y_<3> GF_NI_IN_C_BASE_0/pdrive_y_<2>
+ GF_NI_IN_C_BASE_0/pdrive_x_<2> GF_NI_IN_C_BASE_0/pdrive_x_<1> GF_NI_IN_C_BASE_0/pdrive_y_<1>
+ GF_NI_IN_C_BASE_0/pdrive_y_<0> GF_NI_IN_C_BASE_0/pdrive_x_<0> GF_NI_IN_C_BASE_0/ndrive_Y_<3>
+ GF_NI_IN_C_BASE_0/ndrive_x_<3> GF_NI_IN_C_BASE_0/ndrive_y_<2> GF_NI_IN_C_BASE_0/ndrive_x_<2>
+ GF_NI_IN_C_BASE_0/ndrive_Y_<1> GF_NI_IN_C_BASE_0/ndrive_x_<1> GF_NI_IN_C_BASE_0/ndrive_y_<0>
+ GF_NI_IN_C_BASE_0/ndrive_x_<0> Y PU PD DVDD DVSS GF_NI_IN_C_BASE_0/PAD VDD DVSS
+ DVSS DVDD DVDD DVSS VDD DVDD VDD DVDD DVDD VDD DVDD DVDD DVDD VDD DVDD DVDD DVDD
+ DVSS DVSS DVDD DVDD DVDD VSS DVSS DVDD DVSS DVDD DVDD GF_NI_IN_C_BASE
.ends

