* NGSPICE file created from gf180mcu_fd_io__dvss_flat.ext - technology: gf180mcuD

.subckt gf180mcu_fd_io__dvss_flat VDD DVDD DVSS
X0 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/comp018green_esd_rc_v5p0_0.ppolyf_u_CDNS_406619531453_5.MINUS GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/comp018green_esd_rc_v5p0_0.ppolyf_u_CDNS_406619531453_5.PLUS DVDD ppolyf_u r_width=0.8u r_length=63.854996u
X1 DVDD GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/pmos_6p0_CDNS_406619531455_0.D DVSS DVSS nfet_06v0 ad=12.999999p pd=50.52u as=12.999999p ps=50.52u w=50u l=0.7u
X2 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/pmos_6p0_CDNS_406619531455_0.D GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/pmos_6p0_CDNS_406619531456_0.D DVSS DVSS nfet_06v0 ad=1.3p pd=5.52u as=1.3p ps=5.52u w=5u l=0.7u
X3 DVDD GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/pmos_6p0_CDNS_406619531455_0.D DVSS DVSS nfet_06v0 ad=12.999999p pd=50.52u as=12.999999p ps=50.52u w=50u l=0.7u
X4 DVDD GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/pmos_6p0_CDNS_406619531455_0.D DVSS DVSS nfet_06v0 ad=12.999999p pd=50.52u as=21.999998p ps=0.10088m w=50u l=0.7u
X5 DVSS GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/pmos_6p0_CDNS_406619531452_0.D GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/pmos_6p0_CDNS_406619531456_0.D DVSS nfet_06v0 ad=1.3p pd=5.52u as=1.3p ps=5.52u w=5u l=0.7u
X6 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/comp018green_esd_rc_v5p0_0.ppolyf_u_CDNS_406619531453_2.MINUS GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/comp018green_esd_rc_v5p0_0.ppolyf_u_CDNS_406619531453_2.PLUS DVDD ppolyf_u r_width=0.8u r_length=63.854996u
X7 DVSS GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/pmos_6p0_CDNS_406619531455_0.D DVDD DVSS nfet_06v0 ad=21.999998p pd=0.10088m as=12.999999p ps=50.52u w=50u l=0.7u
X8 DVSS GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/pmos_6p0_CDNS_406619531455_0.D DVDD DVSS nfet_06v0 ad=12.999999p pd=50.52u as=12.999999p ps=50.52u w=50u l=0.7u
X9 DVDD GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/comp018green_esd_rc_v5p0_0.VRC GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/pmos_6p0_CDNS_406619531452_0.D DVDD pfet_06v0 ad=1.3p pd=5.52u as=1.3p ps=5.52u w=5u l=0.7u
X10 DVSS GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/pmos_6p0_CDNS_406619531455_0.D DVDD DVSS nfet_06v0 ad=12.999999p pd=50.52u as=12.999999p ps=50.52u w=50u l=0.7u
X11 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/pmos_6p0_CDNS_406619531452_0.D GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/comp018green_esd_rc_v5p0_0.VRC DVDD DVDD pfet_06v0 ad=1.3p pd=5.52u as=1.3p ps=5.52u w=5u l=0.7u
X12 DVDD GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/pmos_6p0_CDNS_406619531455_0.D DVSS DVSS nfet_06v0 ad=12.999999p pd=50.52u as=12.999999p ps=50.52u w=50u l=0.7u
X13 DVSS GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/pmos_6p0_CDNS_406619531455_0.D DVDD DVSS nfet_06v0 ad=12.999999p pd=50.52u as=12.999999p ps=50.52u w=50u l=0.7u
X14 DVDD GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/pmos_6p0_CDNS_406619531455_0.D DVSS DVSS nfet_06v0 ad=12.999999p pd=50.52u as=12.999999p ps=50.52u w=50u l=0.7u
X15 DVDD DVSS cap_nmos_06v0 c_width=15u c_length=15u
X16 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/comp018green_esd_rc_v5p0_0.ppolyf_u_CDNS_406619531453_2.MINUS GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/comp018green_esd_rc_v5p0_0.ppolyf_u_CDNS_406619531453_4.PLUS DVDD ppolyf_u r_width=0.8u r_length=63.854996u
X17 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/pmos_6p0_CDNS_406619531455_0.D GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/pmos_6p0_CDNS_406619531456_0.D DVDD DVDD pfet_06v0 ad=1.3p pd=5.52u as=1.3p ps=5.52u w=5u l=0.7u
X18 DVSS GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/pmos_6p0_CDNS_406619531455_0.D DVDD DVSS nfet_06v0 ad=12.999999p pd=50.52u as=12.999999p ps=50.52u w=50u l=0.7u
X19 DVSS GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/pmos_6p0_CDNS_406619531455_0.D DVDD DVSS nfet_06v0 ad=12.999999p pd=50.52u as=12.999999p ps=50.52u w=50u l=0.7u
X20 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/pmos_6p0_CDNS_406619531455_0.D GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/pmos_6p0_CDNS_406619531456_0.D DVDD DVDD pfet_06v0 ad=1.3p pd=5.52u as=1.3p ps=5.52u w=5u l=0.7u
X21 DVDD GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/pmos_6p0_CDNS_406619531455_0.D DVSS DVSS nfet_06v0 ad=12.999999p pd=50.52u as=12.999999p ps=50.52u w=50u l=0.7u
X22 DVDD GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/pmos_6p0_CDNS_406619531455_0.D DVSS DVSS nfet_06v0 ad=12.999999p pd=50.52u as=12.999999p ps=50.52u w=50u l=0.7u
X23 DVDD GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/pmos_6p0_CDNS_406619531455_0.D DVSS DVSS nfet_06v0 ad=12.999999p pd=50.52u as=12.999999p ps=50.52u w=50u l=0.7u
X24 DVDD GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/pmos_6p0_CDNS_406619531455_0.D DVSS DVSS nfet_06v0 ad=12.999999p pd=50.52u as=12.999999p ps=50.52u w=50u l=0.7u
D0 DVSS DVDD diode_nd2ps_06v0 pj=82u area=40p
X25 DVDD GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/pmos_6p0_CDNS_406619531456_0.D GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/pmos_6p0_CDNS_406619531455_0.D DVDD pfet_06v0 ad=1.3p pd=5.52u as=1.3p ps=5.52u w=5u l=0.7u
X26 DVSS GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/pmos_6p0_CDNS_406619531455_0.D DVDD DVSS nfet_06v0 ad=12.999999p pd=50.52u as=12.999999p ps=50.52u w=50u l=0.7u
X27 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/pmos_6p0_CDNS_406619531455_0.D GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/pmos_6p0_CDNS_406619531456_0.D DVDD DVDD pfet_06v0 ad=1.3p pd=5.52u as=1.3p ps=5.52u w=5u l=0.7u
X28 DVSS GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/pmos_6p0_CDNS_406619531455_0.D DVDD DVSS nfet_06v0 ad=12.999999p pd=50.52u as=12.999999p ps=50.52u w=50u l=0.7u
X29 DVSS GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/pmos_6p0_CDNS_406619531455_0.D DVDD DVSS nfet_06v0 ad=12.999999p pd=50.52u as=12.999999p ps=50.52u w=50u l=0.7u
X30 DVDD DVSS cap_nmos_06v0 c_width=15u c_length=15u
X31 DVDD DVSS cap_nmos_06v0 c_width=15u c_length=15u
X32 DVDD GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/pmos_6p0_CDNS_406619531456_0.D GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/pmos_6p0_CDNS_406619531455_0.D DVDD pfet_06v0 ad=1.3p pd=5.52u as=1.3p ps=5.52u w=5u l=0.7u
X33 DVDD GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/pmos_6p0_CDNS_406619531455_0.D DVSS DVSS nfet_06v0 ad=12.999999p pd=50.52u as=12.999999p ps=50.52u w=50u l=0.7u
X34 DVDD GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/pmos_6p0_CDNS_406619531455_0.D DVSS DVSS nfet_06v0 ad=12.999999p pd=50.52u as=12.999999p ps=50.52u w=50u l=0.7u
X35 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/comp018green_esd_rc_v5p0_0.ppolyf_u_CDNS_406619531453_1.MINUS GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/comp018green_esd_rc_v5p0_0.ppolyf_u_CDNS_406619531453_0.PLUS DVDD ppolyf_u r_width=0.8u r_length=63.854996u
X36 DVSS GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/pmos_6p0_CDNS_406619531455_0.D DVDD DVSS nfet_06v0 ad=21.999998p pd=0.10088m as=12.999999p ps=50.52u w=50u l=0.7u
X37 DVDD GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/pmos_6p0_CDNS_406619531456_0.D GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/pmos_6p0_CDNS_406619531455_0.D DVDD pfet_06v0 ad=1.3p pd=5.52u as=1.3p ps=5.52u w=5u l=0.7u
X38 DVDD GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/pmos_6p0_CDNS_406619531455_0.D DVSS DVSS nfet_06v0 ad=12.999999p pd=50.52u as=12.999999p ps=50.52u w=50u l=0.7u
X39 DVSS GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/pmos_6p0_CDNS_406619531455_0.D DVDD DVSS nfet_06v0 ad=12.999999p pd=50.52u as=12.999999p ps=50.52u w=50u l=0.7u
X40 DVDD GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/pmos_6p0_CDNS_406619531456_0.D GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/pmos_6p0_CDNS_406619531455_0.D DVDD pfet_06v0 ad=1.3p pd=5.52u as=1.3p ps=5.52u w=5u l=0.7u
X41 DVDD GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/pmos_6p0_CDNS_406619531455_0.D DVSS DVSS nfet_06v0 ad=12.999999p pd=50.52u as=12.999999p ps=50.52u w=50u l=0.7u
X42 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/comp018green_esd_rc_v5p0_0.ppolyf_u_CDNS_406619531453_5.MINUS GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/comp018green_esd_rc_v5p0_0.ppolyf_u_CDNS_406619531453_3.PLUS DVDD ppolyf_u r_width=0.8u r_length=63.854996u
X43 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/pmos_6p0_CDNS_406619531455_0.D GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/pmos_6p0_CDNS_406619531456_0.D DVDD DVDD pfet_06v0 ad=1.3p pd=5.52u as=2.2p ps=10.879999u w=5u l=0.7u
X44 DVDD GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/pmos_6p0_CDNS_406619531455_0.D DVSS DVSS nfet_06v0 ad=12.999999p pd=50.52u as=12.999999p ps=50.52u w=50u l=0.7u
X45 DVDD GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/pmos_6p0_CDNS_406619531456_0.D GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/pmos_6p0_CDNS_406619531455_0.D DVDD pfet_06v0 ad=1.3p pd=5.52u as=1.3p ps=5.52u w=5u l=0.7u
X46 DVSS GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/pmos_6p0_CDNS_406619531456_0.D GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/pmos_6p0_CDNS_406619531455_0.D DVSS nfet_06v0 ad=1.3p pd=5.52u as=1.3p ps=5.52u w=5u l=0.7u
X47 DVSS GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/pmos_6p0_CDNS_406619531455_0.D DVDD DVSS nfet_06v0 ad=12.999999p pd=50.52u as=12.999999p ps=50.52u w=50u l=0.7u
X48 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/pmos_6p0_CDNS_406619531455_0.D GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/pmos_6p0_CDNS_406619531456_0.D DVSS DVSS nfet_06v0 ad=1.3p pd=5.52u as=1.3p ps=5.52u w=5u l=0.7u
X49 DVSS GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/pmos_6p0_CDNS_406619531455_0.D DVDD DVSS nfet_06v0 ad=12.999999p pd=50.52u as=12.999999p ps=50.52u w=50u l=0.7u
X50 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/pmos_6p0_CDNS_406619531455_0.D GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/pmos_6p0_CDNS_406619531456_0.D DVDD DVDD pfet_06v0 ad=1.3p pd=5.52u as=1.3p ps=5.52u w=5u l=0.7u
X51 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/pmos_6p0_CDNS_406619531452_0.D GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/comp018green_esd_rc_v5p0_0.VRC DVSS DVSS nfet_06v0 ad=2.2p pd=10.879999u as=2.2p ps=10.879999u w=5u l=0.7u
X52 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/comp018green_esd_rc_v5p0_0.ppolyf_u_CDNS_406619531453_3.MINUS GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/comp018green_esd_rc_v5p0_0.ppolyf_u_CDNS_406619531453_3.PLUS DVDD ppolyf_u r_width=0.8u r_length=63.854996u
X53 DVDD GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/pmos_6p0_CDNS_406619531455_0.D DVSS DVSS nfet_06v0 ad=12.999999p pd=50.52u as=12.999999p ps=50.52u w=50u l=0.7u
X54 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/pmos_6p0_CDNS_406619531456_0.D GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/pmos_6p0_CDNS_406619531452_0.D DVSS DVSS nfet_06v0 ad=1.3p pd=5.52u as=2.2p ps=10.879999u w=5u l=0.7u
X55 DVDD GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/pmos_6p0_CDNS_406619531455_0.D DVSS DVSS nfet_06v0 ad=12.999999p pd=50.52u as=12.999999p ps=50.52u w=50u l=0.7u
X56 DVDD GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/pmos_6p0_CDNS_406619531455_0.D DVSS DVSS nfet_06v0 ad=12.999999p pd=50.52u as=12.999999p ps=50.52u w=50u l=0.7u
X57 DVDD GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/pmos_6p0_CDNS_406619531455_0.D DVSS DVSS nfet_06v0 ad=12.999999p pd=50.52u as=12.999999p ps=50.52u w=50u l=0.7u
X58 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/comp018green_esd_rc_v5p0_0.ppolyf_u_CDNS_406619531453_4.MINUS GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/comp018green_esd_rc_v5p0_0.ppolyf_u_CDNS_406619531453_4.PLUS DVDD ppolyf_u r_width=0.8u r_length=63.854996u
X59 DVSS GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/pmos_6p0_CDNS_406619531455_0.D DVDD DVSS nfet_06v0 ad=12.999999p pd=50.52u as=12.999999p ps=50.52u w=50u l=0.7u
X60 DVSS GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/pmos_6p0_CDNS_406619531452_0.D GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/pmos_6p0_CDNS_406619531456_0.D DVSS nfet_06v0 ad=1.3p pd=5.52u as=1.3p ps=5.52u w=5u l=0.7u
X61 DVDD GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/pmos_6p0_CDNS_406619531452_0.D GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/pmos_6p0_CDNS_406619531456_0.D DVDD pfet_06v0 ad=1.3p pd=5.52u as=1.3p ps=5.52u w=5u l=0.7u
X62 DVSS GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/pmos_6p0_CDNS_406619531455_0.D DVDD DVSS nfet_06v0 ad=12.999999p pd=50.52u as=12.999999p ps=50.52u w=50u l=0.7u
X63 DVSS GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/pmos_6p0_CDNS_406619531455_0.D DVDD DVSS nfet_06v0 ad=12.999999p pd=50.52u as=12.999999p ps=50.52u w=50u l=0.7u
X64 DVSS GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/pmos_6p0_CDNS_406619531455_0.D DVDD DVSS nfet_06v0 ad=12.999999p pd=50.52u as=12.999999p ps=50.52u w=50u l=0.7u
X65 DVSS GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/pmos_6p0_CDNS_406619531455_0.D DVDD DVSS nfet_06v0 ad=12.999999p pd=50.52u as=12.999999p ps=50.52u w=50u l=0.7u
X66 DVSS GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/pmos_6p0_CDNS_406619531455_0.D DVDD DVSS nfet_06v0 ad=12.999999p pd=50.52u as=12.999999p ps=50.52u w=50u l=0.7u
X67 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/pmos_6p0_CDNS_406619531456_0.D GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/pmos_6p0_CDNS_406619531452_0.D DVDD DVDD pfet_06v0 ad=1.3p pd=5.52u as=1.3p ps=5.52u w=5u l=0.7u
X68 DVDD GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/pmos_6p0_CDNS_406619531456_0.D GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/pmos_6p0_CDNS_406619531455_0.D DVDD pfet_06v0 ad=1.3p pd=5.52u as=1.3p ps=5.52u w=5u l=0.7u
X69 DVDD GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/pmos_6p0_CDNS_406619531455_0.D DVSS DVSS nfet_06v0 ad=12.999999p pd=50.52u as=12.999999p ps=50.52u w=50u l=0.7u
X70 DVDD GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/pmos_6p0_CDNS_406619531455_0.D DVSS DVSS nfet_06v0 ad=12.999999p pd=50.52u as=12.999999p ps=50.52u w=50u l=0.7u
X71 DVSS GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/pmos_6p0_CDNS_406619531455_0.D DVDD DVSS nfet_06v0 ad=12.999999p pd=50.52u as=12.999999p ps=50.52u w=50u l=0.7u
X72 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/pmos_6p0_CDNS_406619531455_0.D GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/pmos_6p0_CDNS_406619531456_0.D DVDD DVDD pfet_06v0 ad=1.3p pd=5.52u as=1.3p ps=5.52u w=5u l=0.7u
X73 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/comp018green_esd_rc_v5p0_0.VRC DVSS cap_nmos_06v0 c_width=25u c_length=10u
X74 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/pmos_6p0_CDNS_406619531455_0.D GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/pmos_6p0_CDNS_406619531456_0.D DVDD DVDD pfet_06v0 ad=1.3p pd=5.52u as=1.3p ps=5.52u w=5u l=0.7u
X75 DVSS GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/pmos_6p0_CDNS_406619531455_0.D DVDD DVSS nfet_06v0 ad=12.999999p pd=50.52u as=12.999999p ps=50.52u w=50u l=0.7u
X76 DVSS GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/pmos_6p0_CDNS_406619531455_0.D DVDD DVSS nfet_06v0 ad=12.999999p pd=50.52u as=12.999999p ps=50.52u w=50u l=0.7u
X77 DVSS GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/pmos_6p0_CDNS_406619531455_0.D DVDD DVSS nfet_06v0 ad=12.999999p pd=50.52u as=12.999999p ps=50.52u w=50u l=0.7u
X78 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/comp018green_esd_rc_v5p0_0.VRC GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/comp018green_esd_rc_v5p0_0.ppolyf_u_CDNS_406619531453_0.PLUS DVDD ppolyf_u r_width=0.8u r_length=63.854996u
X79 DVDD GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/pmos_6p0_CDNS_406619531455_0.D DVSS DVSS nfet_06v0 ad=12.999999p pd=50.52u as=12.999999p ps=50.52u w=50u l=0.7u
X80 DVDD GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/pmos_6p0_CDNS_406619531455_0.D DVSS DVSS nfet_06v0 ad=12.999999p pd=50.52u as=12.999999p ps=50.52u w=50u l=0.7u
X81 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/comp018green_esd_rc_v5p0_0.VRC DVSS cap_nmos_06v0 c_width=25u c_length=10u
X82 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/comp018green_esd_rc_v5p0_0.VRC DVSS cap_nmos_06v0 c_width=25u c_length=10u
X83 DVDD GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/pmos_6p0_CDNS_406619531455_0.D DVSS DVSS nfet_06v0 ad=12.999999p pd=50.52u as=12.999999p ps=50.52u w=50u l=0.7u
X84 DVSS GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/pmos_6p0_CDNS_406619531455_0.D DVDD DVSS nfet_06v0 ad=12.999999p pd=50.52u as=12.999999p ps=50.52u w=50u l=0.7u
X85 DVDD GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/pmos_6p0_CDNS_406619531455_0.D DVSS DVSS nfet_06v0 ad=12.999999p pd=50.52u as=21.999998p ps=0.10088m w=50u l=0.7u
X86 DVSS GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/pmos_6p0_CDNS_406619531455_0.D DVDD DVSS nfet_06v0 ad=21.999998p pd=0.10088m as=12.999999p ps=50.52u w=50u l=0.7u
X87 DVSS GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/pmos_6p0_CDNS_406619531455_0.D DVDD DVSS nfet_06v0 ad=12.999999p pd=50.52u as=12.999999p ps=50.52u w=50u l=0.7u
X88 DVSS GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/pmos_6p0_CDNS_406619531455_0.D DVDD DVSS nfet_06v0 ad=21.999998p pd=0.10088m as=12.999999p ps=50.52u w=50u l=0.7u
X89 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/pmos_6p0_CDNS_406619531455_0.D GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/pmos_6p0_CDNS_406619531456_0.D DVDD DVDD pfet_06v0 ad=1.3p pd=5.52u as=1.3p ps=5.52u w=5u l=0.7u
X90 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/pmos_6p0_CDNS_406619531455_0.D GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/pmos_6p0_CDNS_406619531456_0.D DVDD DVDD pfet_06v0 ad=1.3p pd=5.52u as=1.3p ps=5.52u w=5u l=0.7u
X91 DVSS GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/pmos_6p0_CDNS_406619531455_0.D DVDD DVSS nfet_06v0 ad=12.999999p pd=50.52u as=12.999999p ps=50.52u w=50u l=0.7u
X92 DVSS GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/pmos_6p0_CDNS_406619531455_0.D DVDD DVSS nfet_06v0 ad=12.999999p pd=50.52u as=12.999999p ps=50.52u w=50u l=0.7u
X93 DVSS GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/pmos_6p0_CDNS_406619531456_0.D GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/pmos_6p0_CDNS_406619531455_0.D DVSS nfet_06v0 ad=1.3p pd=5.52u as=1.3p ps=5.52u w=5u l=0.7u
X94 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/pmos_6p0_CDNS_406619531455_0.D GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/pmos_6p0_CDNS_406619531456_0.D DVSS DVSS nfet_06v0 ad=1.3p pd=5.52u as=1.3p ps=5.52u w=5u l=0.7u
X95 DVDD GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/pmos_6p0_CDNS_406619531456_0.D GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/pmos_6p0_CDNS_406619531455_0.D DVDD pfet_06v0 ad=1.3p pd=5.52u as=1.3p ps=5.52u w=5u l=0.7u
X96 DVDD GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/pmos_6p0_CDNS_406619531455_0.D DVSS DVSS nfet_06v0 ad=12.999999p pd=50.52u as=12.999999p ps=50.52u w=50u l=0.7u
X97 DVDD GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/pmos_6p0_CDNS_406619531456_0.D GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/pmos_6p0_CDNS_406619531455_0.D DVDD pfet_06v0 ad=1.3p pd=5.52u as=1.3p ps=5.52u w=5u l=0.7u
X98 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/comp018green_esd_rc_v5p0_0.ppolyf_u_CDNS_406619531453_3.MINUS GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/comp018green_esd_rc_v5p0_0.ppolyf_u_CDNS_406619531453_1.PLUS DVDD ppolyf_u r_width=0.8u r_length=63.854996u
X99 DVDD GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/pmos_6p0_CDNS_406619531455_0.D DVSS DVSS nfet_06v0 ad=12.999999p pd=50.52u as=21.999998p ps=0.10088m w=50u l=0.7u
X100 DVDD GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/pmos_6p0_CDNS_406619531455_0.D DVSS DVSS nfet_06v0 ad=12.999999p pd=50.52u as=12.999999p ps=50.52u w=50u l=0.7u
X101 DVSS GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/pmos_6p0_CDNS_406619531455_0.D DVDD DVSS nfet_06v0 ad=12.999999p pd=50.52u as=12.999999p ps=50.52u w=50u l=0.7u
X102 DVSS GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/pmos_6p0_CDNS_406619531455_0.D DVDD DVSS nfet_06v0 ad=12.999999p pd=50.52u as=12.999999p ps=50.52u w=50u l=0.7u
X103 DVSS GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/pmos_6p0_CDNS_406619531455_0.D DVDD DVSS nfet_06v0 ad=12.999999p pd=50.52u as=12.999999p ps=50.52u w=50u l=0.7u
X104 DVSS GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/pmos_6p0_CDNS_406619531456_0.D GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/pmos_6p0_CDNS_406619531455_0.D DVSS nfet_06v0 ad=2.2p pd=10.879999u as=1.3p ps=5.52u w=5u l=0.7u
X105 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/comp018green_esd_rc_v5p0_0.VRC DVSS cap_nmos_06v0 c_width=25u c_length=10u
X106 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/comp018green_esd_rc_v5p0_0.VRC DVSS cap_nmos_06v0 c_width=25u c_length=10u
X107 DVSS GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/pmos_6p0_CDNS_406619531455_0.D DVDD DVSS nfet_06v0 ad=12.999999p pd=50.52u as=12.999999p ps=50.52u w=50u l=0.7u
X108 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/comp018green_esd_rc_v5p0_0.ppolyf_u_CDNS_406619531453_4.MINUS GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/comp018green_esd_rc_v5p0_0.ppolyf_u_CDNS_406619531453_5.PLUS DVDD ppolyf_u r_width=0.8u r_length=63.854996u
X109 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/pmos_6p0_CDNS_406619531456_0.D GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/pmos_6p0_CDNS_406619531452_0.D DVSS DVSS nfet_06v0 ad=1.3p pd=5.52u as=1.3p ps=5.52u w=5u l=0.7u
X110 DVDD GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/pmos_6p0_CDNS_406619531455_0.D DVSS DVSS nfet_06v0 ad=12.999999p pd=50.52u as=12.999999p ps=50.52u w=50u l=0.7u
X111 DVDD GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/pmos_6p0_CDNS_406619531455_0.D DVSS DVSS nfet_06v0 ad=12.999999p pd=50.52u as=12.999999p ps=50.52u w=50u l=0.7u
X112 DVSS GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/pmos_6p0_CDNS_406619531452_0.D GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/pmos_6p0_CDNS_406619531456_0.D DVSS nfet_06v0 ad=1.3p pd=5.52u as=1.3p ps=5.52u w=5u l=0.7u
X113 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/comp018green_esd_rc_v5p0_0.VRC DVSS cap_nmos_06v0 c_width=25u c_length=10u
D1 DVSS DVDD diode_nd2ps_06v0 pj=82u area=40p
X114 DVDD GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/comp018green_esd_rc_v5p0_0.ppolyf_u_CDNS_406619531453_2.PLUS DVDD ppolyf_u r_width=0.8u r_length=63.854996u
X115 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/comp018green_esd_rc_v5p0_0.VRC DVSS cap_nmos_06v0 c_width=25u c_length=10u
X116 DVSS GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/pmos_6p0_CDNS_406619531455_0.D DVDD DVSS nfet_06v0 ad=12.999999p pd=50.52u as=12.999999p ps=50.52u w=50u l=0.7u
X117 DVDD GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/pmos_6p0_CDNS_406619531455_0.D DVSS DVSS nfet_06v0 ad=12.999999p pd=50.52u as=12.999999p ps=50.52u w=50u l=0.7u
D2 DVSS DVDD diode_nd2ps_06v0 pj=82u area=40p
X118 DVDD GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/comp018green_esd_rc_v5p0_0.VRC GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/pmos_6p0_CDNS_406619531452_0.D DVDD pfet_06v0 ad=1.3p pd=5.52u as=1.3p ps=5.52u w=5u l=0.7u
X119 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/pmos_6p0_CDNS_406619531452_0.D GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/comp018green_esd_rc_v5p0_0.VRC DVDD DVDD pfet_06v0 ad=1.3p pd=5.52u as=2.2p ps=10.879999u w=5u l=0.7u
X120 DVDD GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/pmos_6p0_CDNS_406619531455_0.D DVSS DVSS nfet_06v0 ad=12.999999p pd=50.52u as=12.999999p ps=50.52u w=50u l=0.7u
X121 DVDD GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/pmos_6p0_CDNS_406619531455_0.D DVSS DVSS nfet_06v0 ad=12.999999p pd=50.52u as=12.999999p ps=50.52u w=50u l=0.7u
X122 DVSS GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/pmos_6p0_CDNS_406619531455_0.D DVDD DVSS nfet_06v0 ad=12.999999p pd=50.52u as=12.999999p ps=50.52u w=50u l=0.7u
X123 DVDD GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/pmos_6p0_CDNS_406619531456_0.D GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/pmos_6p0_CDNS_406619531455_0.D DVDD pfet_06v0 ad=1.3p pd=5.52u as=1.3p ps=5.52u w=5u l=0.7u
X124 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/comp018green_esd_rc_v5p0_0.VRC DVSS cap_nmos_06v0 c_width=25u c_length=10u
X125 DVDD DVSS cap_nmos_06v0 c_width=15u c_length=15u
X126 DVDD GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/pmos_6p0_CDNS_406619531455_0.D DVSS DVSS nfet_06v0 ad=12.999999p pd=50.52u as=12.999999p ps=50.52u w=50u l=0.7u
X127 DVDD GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/pmos_6p0_CDNS_406619531455_0.D DVSS DVSS nfet_06v0 ad=12.999999p pd=50.52u as=12.999999p ps=50.52u w=50u l=0.7u
X128 DVDD GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/pmos_6p0_CDNS_406619531456_0.D GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/pmos_6p0_CDNS_406619531455_0.D DVDD pfet_06v0 ad=1.3p pd=5.52u as=1.3p ps=5.52u w=5u l=0.7u
X129 DVDD GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/pmos_6p0_CDNS_406619531455_0.D DVSS DVSS nfet_06v0 ad=12.999999p pd=50.52u as=12.999999p ps=50.52u w=50u l=0.7u
X130 DVDD GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/pmos_6p0_CDNS_406619531455_0.D DVSS DVSS nfet_06v0 ad=12.999999p pd=50.52u as=21.999998p ps=0.10088m w=50u l=0.7u
X131 DVSS GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/pmos_6p0_CDNS_406619531455_0.D DVDD DVSS nfet_06v0 ad=12.999999p pd=50.52u as=12.999999p ps=50.52u w=50u l=0.7u
X132 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/pmos_6p0_CDNS_406619531455_0.D GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/pmos_6p0_CDNS_406619531456_0.D DVDD DVDD pfet_06v0 ad=1.3p pd=5.52u as=1.3p ps=5.52u w=5u l=0.7u
X133 DVDD GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/pmos_6p0_CDNS_406619531456_0.D GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/pmos_6p0_CDNS_406619531455_0.D DVDD pfet_06v0 ad=1.3p pd=5.52u as=1.3p ps=5.52u w=5u l=0.7u
X134 DVSS GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/pmos_6p0_CDNS_406619531455_0.D DVDD DVSS nfet_06v0 ad=12.999999p pd=50.52u as=12.999999p ps=50.52u w=50u l=0.7u
X135 DVDD GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/pmos_6p0_CDNS_406619531456_0.D GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/pmos_6p0_CDNS_406619531455_0.D DVDD pfet_06v0 ad=2.2p pd=10.879999u as=1.3p ps=5.52u w=5u l=0.7u
D3 DVSS DVDD diode_nd2ps_06v0 pj=82u area=40p
X136 DVSS GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/pmos_6p0_CDNS_406619531455_0.D DVDD DVSS nfet_06v0 ad=12.999999p pd=50.52u as=12.999999p ps=50.52u w=50u l=0.7u
X137 DVDD GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/pmos_6p0_CDNS_406619531455_0.D DVSS DVSS nfet_06v0 ad=12.999999p pd=50.52u as=12.999999p ps=50.52u w=50u l=0.7u
X138 DVDD GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/pmos_6p0_CDNS_406619531455_0.D DVSS DVSS nfet_06v0 ad=12.999999p pd=50.52u as=12.999999p ps=50.52u w=50u l=0.7u
X139 DVDD GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/pmos_6p0_CDNS_406619531455_0.D DVSS DVSS nfet_06v0 ad=12.999999p pd=50.52u as=12.999999p ps=50.52u w=50u l=0.7u
X140 DVDD GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/pmos_6p0_CDNS_406619531455_0.D DVSS DVSS nfet_06v0 ad=12.999999p pd=50.52u as=12.999999p ps=50.52u w=50u l=0.7u
X141 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/comp018green_esd_rc_v5p0_0.ppolyf_u_CDNS_406619531453_1.MINUS GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/comp018green_esd_rc_v5p0_0.ppolyf_u_CDNS_406619531453_1.PLUS DVDD ppolyf_u r_width=0.8u r_length=63.854996u
X142 DVSS GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/pmos_6p0_CDNS_406619531455_0.D DVDD DVSS nfet_06v0 ad=12.999999p pd=50.52u as=12.999999p ps=50.52u w=50u l=0.7u
X143 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/pmos_6p0_CDNS_406619531456_0.D GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/pmos_6p0_CDNS_406619531452_0.D DVSS DVSS nfet_06v0 ad=1.3p pd=5.52u as=1.3p ps=5.52u w=5u l=0.7u
X144 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/pmos_6p0_CDNS_406619531456_0.D GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/pmos_6p0_CDNS_406619531452_0.D DVDD DVDD pfet_06v0 ad=2.2p pd=10.879999u as=1.3p ps=5.52u w=5u l=0.7u
X145 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/pmos_6p0_CDNS_406619531455_0.D GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/pmos_6p0_CDNS_406619531456_0.D DVDD DVDD pfet_06v0 ad=1.3p pd=5.52u as=1.3p ps=5.52u w=5u l=0.7u
X146 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/pmos_6p0_CDNS_406619531455_0.D GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/pmos_6p0_CDNS_406619531456_0.D DVDD DVDD pfet_06v0 ad=1.3p pd=5.52u as=1.3p ps=5.52u w=5u l=0.7u
X147 DVSS GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/pmos_6p0_CDNS_406619531455_0.D DVDD DVSS nfet_06v0 ad=12.999999p pd=50.52u as=12.999999p ps=50.52u w=50u l=0.7u
.ends

