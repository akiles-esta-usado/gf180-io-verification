* NGSPICE file created from gf180mcu_fd_io__asig_5p0.ext - technology: gf180mcuD

.subckt x5LM_METAL_RAIL_PAD_60 Bondpad_5LM_0/m5_n400_0# 5LM_METAL_RAIL_0/VDD 5LM_METAL_RAIL_0/VSS
+ 5LM_METAL_RAIL_0/DVDD 5LM_METAL_RAIL_0/DVSS VSUBS
.ends

.subckt nmoscap_6p0_CDNS_406619531450 G D
X0 G D cap_nmos_06v0 c_width=15u c_length=15u
.ends

.subckt np_6p0_CDNS_406619531451 MINUS
D0 VSUBS MINUS diode_nd2ps_06v0 pj=82u area=40p
.ends

.subckt pn_6p0_CDNS_4066195314552 w_n120_n120# PLUS
D0 PLUS w_n120_n120# diode_pd2nw_06v0 pj=0.106m area=0.15n
.ends

.subckt np_6p0_CDNS_4066195314553 MINUS
D0 VSUBS MINUS diode_nd2ps_06v0 pj=0.106m area=0.15n
.ends

.subckt comp018green_esd_hbm pn_6p0_CDNS_4066195314552_3/PLUS m2_n5_43# w_601_591#
Xpn_6p0_CDNS_4066195314552_0 w_601_591# pn_6p0_CDNS_4066195314552_3/PLUS pn_6p0_CDNS_4066195314552
Xpn_6p0_CDNS_4066195314552_1 w_601_591# pn_6p0_CDNS_4066195314552_3/PLUS pn_6p0_CDNS_4066195314552
Xpn_6p0_CDNS_4066195314552_2 w_601_591# pn_6p0_CDNS_4066195314552_3/PLUS pn_6p0_CDNS_4066195314552
Xpn_6p0_CDNS_4066195314552_3 w_601_591# pn_6p0_CDNS_4066195314552_3/PLUS pn_6p0_CDNS_4066195314552
Xnp_6p0_CDNS_4066195314553_0 pn_6p0_CDNS_4066195314552_3/PLUS np_6p0_CDNS_4066195314553
Xnp_6p0_CDNS_4066195314553_1 pn_6p0_CDNS_4066195314552_3/PLUS np_6p0_CDNS_4066195314553
Xnp_6p0_CDNS_4066195314553_2 pn_6p0_CDNS_4066195314552_3/PLUS np_6p0_CDNS_4066195314553
Xnp_6p0_CDNS_4066195314553_3 pn_6p0_CDNS_4066195314552_3/PLUS np_6p0_CDNS_4066195314553
.ends

.subckt GF_NI_ASIG_5P0_BASE m2_828_38097# VSUBS m2_13160_36497# comp018green_esd_hbm_0/pn_6p0_CDNS_4066195314552_3/PLUS
+ nmoscap_6p0_CDNS_406619531450_9/D np_6p0_CDNS_406619531451_3/MINUS
Xnmoscap_6p0_CDNS_406619531450_30 np_6p0_CDNS_406619531451_3/MINUS nmoscap_6p0_CDNS_406619531450_9/D
+ nmoscap_6p0_CDNS_406619531450
Xnmoscap_6p0_CDNS_406619531450_31 np_6p0_CDNS_406619531451_3/MINUS nmoscap_6p0_CDNS_406619531450_9/D
+ nmoscap_6p0_CDNS_406619531450
Xnmoscap_6p0_CDNS_406619531450_20 np_6p0_CDNS_406619531451_3/MINUS nmoscap_6p0_CDNS_406619531450_9/D
+ nmoscap_6p0_CDNS_406619531450
Xnmoscap_6p0_CDNS_406619531450_32 np_6p0_CDNS_406619531451_3/MINUS nmoscap_6p0_CDNS_406619531450_9/D
+ nmoscap_6p0_CDNS_406619531450
Xnmoscap_6p0_CDNS_406619531450_10 np_6p0_CDNS_406619531451_3/MINUS nmoscap_6p0_CDNS_406619531450_9/D
+ nmoscap_6p0_CDNS_406619531450
Xnmoscap_6p0_CDNS_406619531450_21 np_6p0_CDNS_406619531451_3/MINUS nmoscap_6p0_CDNS_406619531450_9/D
+ nmoscap_6p0_CDNS_406619531450
Xnmoscap_6p0_CDNS_406619531450_11 np_6p0_CDNS_406619531451_3/MINUS nmoscap_6p0_CDNS_406619531450_9/D
+ nmoscap_6p0_CDNS_406619531450
Xnmoscap_6p0_CDNS_406619531450_22 np_6p0_CDNS_406619531451_3/MINUS nmoscap_6p0_CDNS_406619531450_9/D
+ nmoscap_6p0_CDNS_406619531450
Xnmoscap_6p0_CDNS_406619531450_33 np_6p0_CDNS_406619531451_3/MINUS nmoscap_6p0_CDNS_406619531450_9/D
+ nmoscap_6p0_CDNS_406619531450
Xnmoscap_6p0_CDNS_406619531450_12 np_6p0_CDNS_406619531451_3/MINUS nmoscap_6p0_CDNS_406619531450_9/D
+ nmoscap_6p0_CDNS_406619531450
Xnmoscap_6p0_CDNS_406619531450_23 np_6p0_CDNS_406619531451_3/MINUS nmoscap_6p0_CDNS_406619531450_9/D
+ nmoscap_6p0_CDNS_406619531450
Xnmoscap_6p0_CDNS_406619531450_34 np_6p0_CDNS_406619531451_3/MINUS nmoscap_6p0_CDNS_406619531450_9/D
+ nmoscap_6p0_CDNS_406619531450
Xnmoscap_6p0_CDNS_406619531450_35 np_6p0_CDNS_406619531451_3/MINUS nmoscap_6p0_CDNS_406619531450_9/D
+ nmoscap_6p0_CDNS_406619531450
Xnmoscap_6p0_CDNS_406619531450_24 np_6p0_CDNS_406619531451_3/MINUS nmoscap_6p0_CDNS_406619531450_9/D
+ nmoscap_6p0_CDNS_406619531450
Xnmoscap_6p0_CDNS_406619531450_13 np_6p0_CDNS_406619531451_3/MINUS nmoscap_6p0_CDNS_406619531450_9/D
+ nmoscap_6p0_CDNS_406619531450
Xnmoscap_6p0_CDNS_406619531450_0 np_6p0_CDNS_406619531451_3/MINUS nmoscap_6p0_CDNS_406619531450_9/D
+ nmoscap_6p0_CDNS_406619531450
Xnmoscap_6p0_CDNS_406619531450_14 np_6p0_CDNS_406619531451_3/MINUS nmoscap_6p0_CDNS_406619531450_9/D
+ nmoscap_6p0_CDNS_406619531450
Xnmoscap_6p0_CDNS_406619531450_25 np_6p0_CDNS_406619531451_3/MINUS nmoscap_6p0_CDNS_406619531450_9/D
+ nmoscap_6p0_CDNS_406619531450
Xnmoscap_6p0_CDNS_406619531450_1 np_6p0_CDNS_406619531451_3/MINUS nmoscap_6p0_CDNS_406619531450_9/D
+ nmoscap_6p0_CDNS_406619531450
Xnmoscap_6p0_CDNS_406619531450_26 np_6p0_CDNS_406619531451_3/MINUS nmoscap_6p0_CDNS_406619531450_9/D
+ nmoscap_6p0_CDNS_406619531450
Xnmoscap_6p0_CDNS_406619531450_15 np_6p0_CDNS_406619531451_3/MINUS nmoscap_6p0_CDNS_406619531450_9/D
+ nmoscap_6p0_CDNS_406619531450
Xnp_6p0_CDNS_406619531451_0 np_6p0_CDNS_406619531451_3/MINUS np_6p0_CDNS_406619531451
Xnmoscap_6p0_CDNS_406619531450_27 np_6p0_CDNS_406619531451_3/MINUS nmoscap_6p0_CDNS_406619531450_9/D
+ nmoscap_6p0_CDNS_406619531450
Xnmoscap_6p0_CDNS_406619531450_16 np_6p0_CDNS_406619531451_3/MINUS nmoscap_6p0_CDNS_406619531450_9/D
+ nmoscap_6p0_CDNS_406619531450
Xnmoscap_6p0_CDNS_406619531450_2 np_6p0_CDNS_406619531451_3/MINUS nmoscap_6p0_CDNS_406619531450_9/D
+ nmoscap_6p0_CDNS_406619531450
Xnp_6p0_CDNS_406619531451_1 np_6p0_CDNS_406619531451_3/MINUS np_6p0_CDNS_406619531451
Xnmoscap_6p0_CDNS_406619531450_17 np_6p0_CDNS_406619531451_3/MINUS nmoscap_6p0_CDNS_406619531450_9/D
+ nmoscap_6p0_CDNS_406619531450
Xnmoscap_6p0_CDNS_406619531450_3 np_6p0_CDNS_406619531451_3/MINUS nmoscap_6p0_CDNS_406619531450_9/D
+ nmoscap_6p0_CDNS_406619531450
Xnmoscap_6p0_CDNS_406619531450_28 np_6p0_CDNS_406619531451_3/MINUS nmoscap_6p0_CDNS_406619531450_9/D
+ nmoscap_6p0_CDNS_406619531450
Xnp_6p0_CDNS_406619531451_2 np_6p0_CDNS_406619531451_3/MINUS np_6p0_CDNS_406619531451
Xnmoscap_6p0_CDNS_406619531450_18 np_6p0_CDNS_406619531451_3/MINUS nmoscap_6p0_CDNS_406619531450_9/D
+ nmoscap_6p0_CDNS_406619531450
Xnmoscap_6p0_CDNS_406619531450_4 np_6p0_CDNS_406619531451_3/MINUS nmoscap_6p0_CDNS_406619531450_9/D
+ nmoscap_6p0_CDNS_406619531450
Xnmoscap_6p0_CDNS_406619531450_29 np_6p0_CDNS_406619531451_3/MINUS nmoscap_6p0_CDNS_406619531450_9/D
+ nmoscap_6p0_CDNS_406619531450
Xnp_6p0_CDNS_406619531451_3 np_6p0_CDNS_406619531451_3/MINUS np_6p0_CDNS_406619531451
Xcomp018green_esd_hbm_0 comp018green_esd_hbm_0/pn_6p0_CDNS_4066195314552_3/PLUS nmoscap_6p0_CDNS_406619531450_9/D
+ np_6p0_CDNS_406619531451_3/MINUS comp018green_esd_hbm
Xnmoscap_6p0_CDNS_406619531450_19 np_6p0_CDNS_406619531451_3/MINUS nmoscap_6p0_CDNS_406619531450_9/D
+ nmoscap_6p0_CDNS_406619531450
Xnmoscap_6p0_CDNS_406619531450_5 np_6p0_CDNS_406619531451_3/MINUS nmoscap_6p0_CDNS_406619531450_9/D
+ nmoscap_6p0_CDNS_406619531450
Xnmoscap_6p0_CDNS_406619531450_6 np_6p0_CDNS_406619531451_3/MINUS nmoscap_6p0_CDNS_406619531450_9/D
+ nmoscap_6p0_CDNS_406619531450
Xnmoscap_6p0_CDNS_406619531450_7 np_6p0_CDNS_406619531451_3/MINUS nmoscap_6p0_CDNS_406619531450_9/D
+ nmoscap_6p0_CDNS_406619531450
Xnmoscap_6p0_CDNS_406619531450_8 np_6p0_CDNS_406619531451_3/MINUS nmoscap_6p0_CDNS_406619531450_9/D
+ nmoscap_6p0_CDNS_406619531450
Xnmoscap_6p0_CDNS_406619531450_9 np_6p0_CDNS_406619531451_3/MINUS nmoscap_6p0_CDNS_406619531450_9/D
+ nmoscap_6p0_CDNS_406619531450
.ends

.subckt gf180mcu_fd_io__asig_5p0 DVSS VDD DVDD VSS ASIG5V
X5LM_METAL_RAIL_PAD_60_0 ASIG5V VDD VSS DVDD DVSS VSS x5LM_METAL_RAIL_PAD_60
XGF_NI_ASIG_5P0_BASE_0 VDD VSS VSS ASIG5V DVSS DVDD GF_NI_ASIG_5P0_BASE
.ends

