* NGSPICE file created from gf180mcu_fd_io__dvss_pex.ext - technology: gf180mcuD

.subckt gf180mcu_fd_io__dvss_pex VDD DVDD DVSS
X0 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/comp018green_esd_rc_v5p0_0.ppolyf_u_CDNS_406619531453_5.MINUS.t1 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/comp018green_esd_rc_v5p0_0.ppolyf_u_CDNS_406619531453_5.PLUS.t1 DVDD.t72 ppolyf_u r_width=0.8u r_length=63.854996u
X1 DVDD.t148 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.t17 DVSS.t161 DVSS.t160 nfet_06v0 ad=12.999999p pd=50.52u as=12.999999p ps=50.52u w=50u l=0.7u
X2 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.t8 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_1.D.t4 DVSS.t196 DVSS.t195 nfet_06v0 ad=1.3p pd=5.52u as=1.3p ps=5.52u w=5u l=0.7u
X3 DVDD.t141 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.t18 DVSS.t159 DVSS.t158 nfet_06v0 ad=12.999999p pd=50.52u as=12.999999p ps=50.52u w=50u l=0.7u
X4 DVDD.t132 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.t19 DVSS.t157 DVSS.t156 nfet_06v0 ad=12.999999p pd=50.52u as=21.999998p ps=0.10088m w=50u l=0.7u
X5 DVSS.t171 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531459_0.D.t3 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_1.D.t1 DVSS.t170 nfet_06v0 ad=1.3p pd=5.52u as=1.3p ps=5.52u w=5u l=0.7u
X6 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/comp018green_esd_rc_v5p0_0.ppolyf_u_CDNS_406619531453_2.MINUS.t1 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/comp018green_esd_rc_v5p0_0.ppolyf_u_CDNS_406619531453_2.PLUS.t1 DVDD.t70 ppolyf_u r_width=0.8u r_length=63.854996u
X7 DVSS.t155 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.t20 DVDD.t142 DVSS.t154 nfet_06v0 ad=21.999998p pd=0.10088m as=12.999999p ps=50.52u w=50u l=0.7u
X8 DVSS.t153 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.t21 DVDD.t139 DVSS.t152 nfet_06v0 ad=12.999999p pd=50.52u as=12.999999p ps=50.52u w=50u l=0.7u
X9 DVDD.t47 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/comp018green_esd_rc_v5p0_0.VRC.t1 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531459_0.D.t1 DVDD.t46 pfet_06v0 ad=1.3p pd=5.52u as=1.3p ps=5.52u w=5u l=0.7u
X10 DVSS.t151 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.t22 DVDD.t137 DVSS.t150 nfet_06v0 ad=12.999999p pd=50.52u as=12.999999p ps=50.52u w=50u l=0.7u
X11 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531459_0.D.t1 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/comp018green_esd_rc_v5p0_0.VRC.t2 DVDD.t63 DVDD.t62 pfet_06v0 ad=1.3p pd=5.52u as=1.3p ps=5.52u w=5u l=0.7u
X12 DVDD.t134 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.t23 DVSS.t149 DVSS.t148 nfet_06v0 ad=12.999999p pd=50.52u as=12.999999p ps=50.52u w=50u l=0.7u
X13 DVSS.t147 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.t24 DVDD.t143 DVSS.t146 nfet_06v0 ad=12.999999p pd=50.52u as=12.999999p ps=50.52u w=50u l=0.7u
X14 DVDD.t140 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.t25 DVSS.t145 DVSS.t144 nfet_06v0 ad=12.999999p pd=50.52u as=12.999999p ps=50.52u w=50u l=0.7u
X15 DVDD.t155 DVSS.t194 cap_nmos_06v0 c_width=15u c_length=15u
X16 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/comp018green_esd_rc_v5p0_0.ppolyf_u_CDNS_406619531453_2.MINUS.t0 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/comp018green_esd_rc_v5p0_0.ppolyf_u_CDNS_406619531453_4.PLUS.t0 DVDD.t61 ppolyf_u r_width=0.8u r_length=63.854996u
X17 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.t0 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_1.D.t5 DVDD.t11 DVDD.t10 pfet_06v0 ad=1.3p pd=5.52u as=1.3p ps=5.52u w=5u l=0.7u
X18 DVSS.t143 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.t26 DVDD.t136 DVSS.t142 nfet_06v0 ad=12.999999p pd=50.52u as=12.999999p ps=50.52u w=50u l=0.7u
X19 DVSS.t141 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.t27 DVDD.t150 DVSS.t140 nfet_06v0 ad=12.999999p pd=50.52u as=12.999999p ps=50.52u w=50u l=0.7u
X20 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.t9 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_1.D.t6 DVDD.t29 DVDD.t28 pfet_06v0 ad=1.3p pd=5.52u as=1.3p ps=5.52u w=5u l=0.7u
X21 DVDD.t154 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.t28 DVSS.t139 DVSS.t138 nfet_06v0 ad=12.999999p pd=50.52u as=12.999999p ps=50.52u w=50u l=0.7u
X22 DVDD.t151 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.t29 DVSS.t137 DVSS.t136 nfet_06v0 ad=12.999999p pd=50.52u as=12.999999p ps=50.52u w=50u l=0.7u
X23 DVDD.t144 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.t30 DVSS.t135 DVSS.t134 nfet_06v0 ad=12.999999p pd=50.52u as=12.999999p ps=50.52u w=50u l=0.7u
X24 DVDD.t145 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.t31 DVSS.t133 DVSS.t132 nfet_06v0 ad=12.999999p pd=50.52u as=12.999999p ps=50.52u w=50u l=0.7u
D0 DVSS.t190 DVDD.t156 diode_nd2ps_06v0 pj=82u area=40p
X25 DVDD.t31 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_1.D.t7 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.t10 DVDD.t30 pfet_06v0 ad=1.3p pd=5.52u as=1.3p ps=5.52u w=5u l=0.7u
X26 DVSS.t131 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.t32 DVDD.t133 DVSS.t130 nfet_06v0 ad=12.999999p pd=50.52u as=12.999999p ps=50.52u w=50u l=0.7u
X27 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.t10 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_1.D.t8 DVDD.t54 DVDD.t53 pfet_06v0 ad=1.3p pd=5.52u as=1.3p ps=5.52u w=5u l=0.7u
X28 DVSS.t129 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.t33 DVDD.t88 DVSS.t128 nfet_06v0 ad=12.999999p pd=50.52u as=12.999999p ps=50.52u w=50u l=0.7u
X29 DVSS.t127 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.t34 DVDD.t117 DVSS.t126 nfet_06v0 ad=12.999999p pd=50.52u as=12.999999p ps=50.52u w=50u l=0.7u
X30 DVDD.t157 DVSS.t193 cap_nmos_06v0 c_width=15u c_length=15u
X31 DVDD.t158 DVSS.t192 cap_nmos_06v0 c_width=15u c_length=15u
X32 DVDD.t49 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_1.D.t9 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.t12 DVDD.t48 pfet_06v0 ad=1.3p pd=5.52u as=1.3p ps=5.52u w=5u l=0.7u
X33 DVDD.t94 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.t35 DVSS.t125 DVSS.t124 nfet_06v0 ad=12.999999p pd=50.52u as=12.999999p ps=50.52u w=50u l=0.7u
X34 DVDD.t147 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.t36 DVSS.t123 DVSS.t122 nfet_06v0 ad=12.999999p pd=50.52u as=12.999999p ps=50.52u w=50u l=0.7u
X35 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/comp018green_esd_rc_v5p0_0.ppolyf_u_CDNS_406619531453_1.MINUS.t1 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/comp018green_esd_rc_v5p0_0.ppolyf_u_CDNS_406619531453_0.PLUS.t1 DVDD.t27 ppolyf_u r_width=0.8u r_length=63.854996u
X36 DVSS.t121 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.t37 DVDD.t153 DVSS.t120 nfet_06v0 ad=21.999998p pd=0.10088m as=12.999999p ps=50.52u w=50u l=0.7u
X37 DVDD.t51 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_1.D.t10 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.t1 DVDD.t50 pfet_06v0 ad=1.3p pd=5.52u as=1.3p ps=5.52u w=5u l=0.7u
X38 DVDD.t152 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.t38 DVSS.t119 DVSS.t118 nfet_06v0 ad=12.999999p pd=50.52u as=12.999999p ps=50.52u w=50u l=0.7u
X39 DVSS.t117 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.t39 DVDD.t131 DVSS.t116 nfet_06v0 ad=12.999999p pd=50.52u as=12.999999p ps=50.52u w=50u l=0.7u
X40 DVDD.t45 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_1.D.t11 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.t4 DVDD.t44 pfet_06v0 ad=1.3p pd=5.52u as=1.3p ps=5.52u w=5u l=0.7u
X41 DVDD.t87 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.t40 DVSS.t115 DVSS.t114 nfet_06v0 ad=12.999999p pd=50.52u as=12.999999p ps=50.52u w=50u l=0.7u
X42 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/comp018green_esd_rc_v5p0_0.ppolyf_u_CDNS_406619531453_5.MINUS.t0 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/comp018green_esd_rc_v5p0_0.ppolyf_u_CDNS_406619531453_3.PLUS.t1 DVDD.t52 ppolyf_u r_width=0.8u r_length=63.854996u
X43 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.t4 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_1.D.t12 DVDD.t20 DVDD.t19 pfet_06v0 ad=1.3p pd=5.52u as=2.2p ps=10.879999u w=5u l=0.7u
X44 DVDD.t92 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.t41 DVSS.t113 DVSS.t112 nfet_06v0 ad=12.999999p pd=50.52u as=12.999999p ps=50.52u w=50u l=0.7u
X45 DVDD.t22 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_1.D.t13 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.t5 DVDD.t21 pfet_06v0 ad=1.3p pd=5.52u as=1.3p ps=5.52u w=5u l=0.7u
X46 DVSS.t198 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_1.D.t14 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.t16 DVSS.t197 nfet_06v0 ad=1.3p pd=5.52u as=1.3p ps=5.52u w=5u l=0.7u
X47 DVSS.t111 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.t42 DVDD.t84 DVSS.t110 nfet_06v0 ad=12.999999p pd=50.52u as=12.999999p ps=50.52u w=50u l=0.7u
X48 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.t6 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_1.D.t15 DVSS.t163 DVSS.t162 nfet_06v0 ad=1.3p pd=5.52u as=1.3p ps=5.52u w=5u l=0.7u
X49 DVSS.t109 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.t43 DVDD.t76 DVSS.t108 nfet_06v0 ad=12.999999p pd=50.52u as=12.999999p ps=50.52u w=50u l=0.7u
X50 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.t3 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_1.D.t16 DVDD.t24 DVDD.t23 pfet_06v0 ad=1.3p pd=5.52u as=1.3p ps=5.52u w=5u l=0.7u
X51 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531459_0.D.t2 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/comp018green_esd_rc_v5p0_0.VRC.t3 DVSS.t188 DVSS.t187 nfet_06v0 ad=2.2p pd=10.879999u as=2.2p ps=10.879999u w=5u l=0.7u
X52 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/comp018green_esd_rc_v5p0_0.ppolyf_u_CDNS_406619531453_3.MINUS.t1 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/comp018green_esd_rc_v5p0_0.ppolyf_u_CDNS_406619531453_3.PLUS.t0 DVDD.t9 ppolyf_u r_width=0.8u r_length=63.854996u
X53 DVDD.t95 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.t44 DVSS.t107 DVSS.t106 nfet_06v0 ad=12.999999p pd=50.52u as=12.999999p ps=50.52u w=50u l=0.7u
X54 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_1.D.t1 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531459_0.D.t4 DVSS.t173 DVSS.t172 nfet_06v0 ad=1.3p pd=5.52u as=2.2p ps=10.879999u w=5u l=0.7u
X55 DVDD.t85 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.t45 DVSS.t105 DVSS.t104 nfet_06v0 ad=12.999999p pd=50.52u as=12.999999p ps=50.52u w=50u l=0.7u
X56 DVDD.t104 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.t46 DVSS.t103 DVSS.t102 nfet_06v0 ad=12.999999p pd=50.52u as=12.999999p ps=50.52u w=50u l=0.7u
X57 DVDD.t77 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.t47 DVSS.t101 DVSS.t100 nfet_06v0 ad=12.999999p pd=50.52u as=12.999999p ps=50.52u w=50u l=0.7u
X58 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/comp018green_esd_rc_v5p0_0.ppolyf_u_CDNS_406619531453_4.MINUS.t1 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/comp018green_esd_rc_v5p0_0.ppolyf_u_CDNS_406619531453_4.PLUS.t1 DVDD.t71 ppolyf_u r_width=0.8u r_length=63.854996u
X59 DVSS.t99 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.t48 DVDD.t75 DVSS.t98 nfet_06v0 ad=12.999999p pd=50.52u as=12.999999p ps=50.52u w=50u l=0.7u
X60 DVSS.t177 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531459_0.D.t5 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_1.D.t0 DVSS.t176 nfet_06v0 ad=1.3p pd=5.52u as=1.3p ps=5.52u w=5u l=0.7u
X61 DVDD.t37 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531459_0.D.t6 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_1.D.t2 DVDD.t36 pfet_06v0 ad=1.3p pd=5.52u as=1.3p ps=5.52u w=5u l=0.7u
X62 DVSS.t97 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.t49 DVDD.t115 DVSS.t96 nfet_06v0 ad=12.999999p pd=50.52u as=12.999999p ps=50.52u w=50u l=0.7u
X63 DVSS.t95 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.t50 DVDD.t82 DVSS.t94 nfet_06v0 ad=12.999999p pd=50.52u as=12.999999p ps=50.52u w=50u l=0.7u
X64 DVSS.t93 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.t51 DVDD.t97 DVSS.t92 nfet_06v0 ad=12.999999p pd=50.52u as=12.999999p ps=50.52u w=50u l=0.7u
X65 DVSS.t91 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.t52 DVDD.t98 DVSS.t90 nfet_06v0 ad=12.999999p pd=50.52u as=12.999999p ps=50.52u w=50u l=0.7u
X66 DVSS.t89 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.t53 DVDD.t100 DVSS.t88 nfet_06v0 ad=12.999999p pd=50.52u as=12.999999p ps=50.52u w=50u l=0.7u
X67 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_1.D.t2 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531459_0.D.t7 DVDD.t39 DVDD.t38 pfet_06v0 ad=1.3p pd=5.52u as=1.3p ps=5.52u w=5u l=0.7u
X68 DVDD.t26 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_1.D.t17 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.t7 DVDD.t25 pfet_06v0 ad=1.3p pd=5.52u as=1.3p ps=5.52u w=5u l=0.7u
X69 DVDD.t91 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.t54 DVSS.t87 DVSS.t86 nfet_06v0 ad=12.999999p pd=50.52u as=12.999999p ps=50.52u w=50u l=0.7u
X70 DVDD.t108 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.t55 DVSS.t85 DVSS.t84 nfet_06v0 ad=12.999999p pd=50.52u as=12.999999p ps=50.52u w=50u l=0.7u
X71 DVSS.t83 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.t56 DVDD.t125 DVSS.t82 nfet_06v0 ad=12.999999p pd=50.52u as=12.999999p ps=50.52u w=50u l=0.7u
X72 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.t2 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_1.D.t18 DVDD.t41 DVDD.t40 pfet_06v0 ad=1.3p pd=5.52u as=1.3p ps=5.52u w=5u l=0.7u
X73 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/comp018green_esd_rc_v5p0_0.VRC.t4 DVSS.t174 cap_nmos_06v0 c_width=25u c_length=10u
X74 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.t5 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_1.D.t19 DVDD.t43 DVDD.t42 pfet_06v0 ad=1.3p pd=5.52u as=1.3p ps=5.52u w=5u l=0.7u
X75 DVSS.t81 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.t57 DVDD.t93 DVSS.t80 nfet_06v0 ad=12.999999p pd=50.52u as=12.999999p ps=50.52u w=50u l=0.7u
X76 DVSS.t79 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.t58 DVDD.t109 DVSS.t78 nfet_06v0 ad=12.999999p pd=50.52u as=12.999999p ps=50.52u w=50u l=0.7u
X77 DVSS.t77 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.t59 DVDD.t130 DVSS.t76 nfet_06v0 ad=12.999999p pd=50.52u as=12.999999p ps=50.52u w=50u l=0.7u
X78 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/comp018green_esd_rc_v5p0_0.VRC.t0 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/comp018green_esd_rc_v5p0_0.ppolyf_u_CDNS_406619531453_0.PLUS.t0 DVDD.t7 ppolyf_u r_width=0.8u r_length=63.854996u
X79 DVDD.t124 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.t60 DVSS.t75 DVSS.t74 nfet_06v0 ad=12.999999p pd=50.52u as=12.999999p ps=50.52u w=50u l=0.7u
X80 DVDD.t128 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.t61 DVSS.t73 DVSS.t72 nfet_06v0 ad=12.999999p pd=50.52u as=12.999999p ps=50.52u w=50u l=0.7u
X81 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/comp018green_esd_rc_v5p0_0.VRC.t5 DVSS.t175 cap_nmos_06v0 c_width=25u c_length=10u
X82 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/comp018green_esd_rc_v5p0_0.VRC.t6 DVSS.t168 cap_nmos_06v0 c_width=25u c_length=10u
X83 DVDD.t129 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.t62 DVSS.t71 DVSS.t70 nfet_06v0 ad=12.999999p pd=50.52u as=12.999999p ps=50.52u w=50u l=0.7u
X84 DVSS.t69 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.t63 DVDD.t127 DVSS.t68 nfet_06v0 ad=12.999999p pd=50.52u as=12.999999p ps=50.52u w=50u l=0.7u
X85 DVDD.t86 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.t64 DVSS.t67 DVSS.t66 nfet_06v0 ad=12.999999p pd=50.52u as=21.999998p ps=0.10088m w=50u l=0.7u
X86 DVSS.t65 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.t65 DVDD.t121 DVSS.t64 nfet_06v0 ad=21.999998p pd=0.10088m as=12.999999p ps=50.52u w=50u l=0.7u
X87 DVSS.t63 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.t66 DVDD.t79 DVSS.t62 nfet_06v0 ad=12.999999p pd=50.52u as=12.999999p ps=50.52u w=50u l=0.7u
X88 DVSS.t61 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.t67 DVDD.t126 DVSS.t60 nfet_06v0 ad=21.999998p pd=0.10088m as=12.999999p ps=50.52u w=50u l=0.7u
X89 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.t12 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_1.D.t20 DVDD.t35 DVDD.t34 pfet_06v0 ad=1.3p pd=5.52u as=1.3p ps=5.52u w=5u l=0.7u
X90 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.t7 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_1.D.t21 DVDD.t60 DVDD.t59 pfet_06v0 ad=1.3p pd=5.52u as=1.3p ps=5.52u w=5u l=0.7u
X91 DVSS.t59 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.t68 DVDD.t96 DVSS.t58 nfet_06v0 ad=12.999999p pd=50.52u as=12.999999p ps=50.52u w=50u l=0.7u
X92 DVSS.t57 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.t69 DVDD.t112 DVSS.t56 nfet_06v0 ad=12.999999p pd=50.52u as=12.999999p ps=50.52u w=50u l=0.7u
X93 DVSS.t186 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_1.D.t22 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.t13 DVSS.t185 nfet_06v0 ad=1.3p pd=5.52u as=1.3p ps=5.52u w=5u l=0.7u
X94 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.t13 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_1.D.t23 DVSS.t179 DVSS.t178 nfet_06v0 ad=1.3p pd=5.52u as=1.3p ps=5.52u w=5u l=0.7u
X95 DVDD.t56 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_1.D.t24 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.t14 DVDD.t55 pfet_06v0 ad=1.3p pd=5.52u as=1.3p ps=5.52u w=5u l=0.7u
X96 DVDD.t111 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.t70 DVSS.t55 DVSS.t54 nfet_06v0 ad=12.999999p pd=50.52u as=12.999999p ps=50.52u w=50u l=0.7u
X97 DVDD.t58 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_1.D.t25 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.t11 DVDD.t57 pfet_06v0 ad=1.3p pd=5.52u as=1.3p ps=5.52u w=5u l=0.7u
X98 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/comp018green_esd_rc_v5p0_0.ppolyf_u_CDNS_406619531453_3.MINUS.t0 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/comp018green_esd_rc_v5p0_0.ppolyf_u_CDNS_406619531453_1.PLUS.t0 DVDD.t8 ppolyf_u r_width=0.8u r_length=63.854996u
X99 DVDD.t110 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.t71 DVSS.t53 DVSS.t52 nfet_06v0 ad=12.999999p pd=50.52u as=21.999998p ps=0.10088m w=50u l=0.7u
X100 DVDD.t99 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.t72 DVSS.t51 DVSS.t50 nfet_06v0 ad=12.999999p pd=50.52u as=12.999999p ps=50.52u w=50u l=0.7u
X101 DVSS.t49 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.t73 DVDD.t116 DVSS.t48 nfet_06v0 ad=12.999999p pd=50.52u as=12.999999p ps=50.52u w=50u l=0.7u
X102 DVSS.t47 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.t74 DVDD.t101 DVSS.t46 nfet_06v0 ad=12.999999p pd=50.52u as=12.999999p ps=50.52u w=50u l=0.7u
X103 DVSS.t45 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.t75 DVDD.t120 DVSS.t44 nfet_06v0 ad=12.999999p pd=50.52u as=12.999999p ps=50.52u w=50u l=0.7u
X104 DVSS.t167 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_1.D.t26 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.t8 DVSS.t166 nfet_06v0 ad=2.2p pd=10.879999u as=1.3p ps=5.52u w=5u l=0.7u
X105 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/comp018green_esd_rc_v5p0_0.VRC.t7 DVSS.t169 cap_nmos_06v0 c_width=25u c_length=10u
X106 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/comp018green_esd_rc_v5p0_0.VRC.t8 DVSS.t1 cap_nmos_06v0 c_width=25u c_length=10u
X107 DVSS.t43 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.t76 DVDD.t119 DVSS.t42 nfet_06v0 ad=12.999999p pd=50.52u as=12.999999p ps=50.52u w=50u l=0.7u
X108 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/comp018green_esd_rc_v5p0_0.ppolyf_u_CDNS_406619531453_4.MINUS.t0 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/comp018green_esd_rc_v5p0_0.ppolyf_u_CDNS_406619531453_5.PLUS.t0 DVDD.t6 ppolyf_u r_width=0.8u r_length=63.854996u
X109 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_1.D.t0 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531459_0.D.t8 DVSS.t165 DVSS.t164 nfet_06v0 ad=1.3p pd=5.52u as=1.3p ps=5.52u w=5u l=0.7u
X110 DVDD.t123 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.t77 DVSS.t41 DVSS.t40 nfet_06v0 ad=12.999999p pd=50.52u as=12.999999p ps=50.52u w=50u l=0.7u
X111 DVDD.t118 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.t78 DVSS.t39 DVSS.t38 nfet_06v0 ad=12.999999p pd=50.52u as=12.999999p ps=50.52u w=50u l=0.7u
X112 DVSS.t181 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531459_0.D.t9 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_1.D.t0 DVSS.t180 nfet_06v0 ad=1.3p pd=5.52u as=1.3p ps=5.52u w=5u l=0.7u
X113 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/comp018green_esd_rc_v5p0_0.VRC.t9 DVSS.t184 cap_nmos_06v0 c_width=25u c_length=10u
D1 DVSS.t190 DVDD.t159 diode_nd2ps_06v0 pj=82u area=40p
X114 DVDD.t5 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/comp018green_esd_rc_v5p0_0.ppolyf_u_CDNS_406619531453_2.PLUS.t0 DVDD.t4 ppolyf_u r_width=0.8u r_length=63.854996u
X115 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/comp018green_esd_rc_v5p0_0.VRC.t10 DVSS.t189 cap_nmos_06v0 c_width=25u c_length=10u
X116 DVSS.t37 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.t79 DVDD.t122 DVSS.t36 nfet_06v0 ad=12.999999p pd=50.52u as=12.999999p ps=50.52u w=50u l=0.7u
X117 DVDD.t78 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.t80 DVSS.t35 DVSS.t34 nfet_06v0 ad=12.999999p pd=50.52u as=12.999999p ps=50.52u w=50u l=0.7u
D2 DVSS.t190 DVDD.t160 diode_nd2ps_06v0 pj=82u area=40p
X118 DVDD.t1 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/comp018green_esd_rc_v5p0_0.VRC.t11 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531459_0.D.t0 DVDD.t0 pfet_06v0 ad=1.3p pd=5.52u as=1.3p ps=5.52u w=5u l=0.7u
X119 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531459_0.D.t0 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/comp018green_esd_rc_v5p0_0.VRC.t12 DVDD.t3 DVDD.t2 pfet_06v0 ad=1.3p pd=5.52u as=2.2p ps=10.879999u w=5u l=0.7u
X120 DVDD.t81 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.t81 DVSS.t33 DVSS.t32 nfet_06v0 ad=12.999999p pd=50.52u as=12.999999p ps=50.52u w=50u l=0.7u
X121 DVDD.t102 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.t82 DVSS.t31 DVSS.t30 nfet_06v0 ad=12.999999p pd=50.52u as=12.999999p ps=50.52u w=50u l=0.7u
X122 DVSS.t29 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.t83 DVDD.t80 DVSS.t28 nfet_06v0 ad=12.999999p pd=50.52u as=12.999999p ps=50.52u w=50u l=0.7u
X123 DVDD.t67 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_1.D.t27 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.t9 DVDD.t66 pfet_06v0 ad=1.3p pd=5.52u as=1.3p ps=5.52u w=5u l=0.7u
X124 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/comp018green_esd_rc_v5p0_0.VRC.t13 DVSS.t0 cap_nmos_06v0 c_width=25u c_length=10u
X125 DVDD.t161 DVSS.t191 cap_nmos_06v0 c_width=15u c_length=15u
X126 DVDD.t90 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.t84 DVSS.t27 DVSS.t26 nfet_06v0 ad=12.999999p pd=50.52u as=12.999999p ps=50.52u w=50u l=0.7u
X127 DVDD.t106 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.t85 DVSS.t25 DVSS.t24 nfet_06v0 ad=12.999999p pd=50.52u as=12.999999p ps=50.52u w=50u l=0.7u
X128 DVDD.t69 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_1.D.t28 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.t15 DVDD.t68 pfet_06v0 ad=1.3p pd=5.52u as=1.3p ps=5.52u w=5u l=0.7u
X129 DVDD.t107 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.t86 DVSS.t23 DVSS.t22 nfet_06v0 ad=12.999999p pd=50.52u as=12.999999p ps=50.52u w=50u l=0.7u
X130 DVDD.t114 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.t87 DVSS.t21 DVSS.t20 nfet_06v0 ad=12.999999p pd=50.52u as=21.999998p ps=0.10088m w=50u l=0.7u
X131 DVSS.t19 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.t88 DVDD.t103 DVSS.t18 nfet_06v0 ad=12.999999p pd=50.52u as=12.999999p ps=50.52u w=50u l=0.7u
X132 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.t1 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_1.D.t29 DVDD.t14 DVDD.t13 pfet_06v0 ad=1.3p pd=5.52u as=1.3p ps=5.52u w=5u l=0.7u
X133 DVDD.t16 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_1.D.t30 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.t2 DVDD.t15 pfet_06v0 ad=1.3p pd=5.52u as=1.3p ps=5.52u w=5u l=0.7u
X134 DVSS.t17 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.t89 DVDD.t135 DVSS.t16 nfet_06v0 ad=12.999999p pd=50.52u as=12.999999p ps=50.52u w=50u l=0.7u
X135 DVDD.t18 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_1.D.t31 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.t3 DVDD.t17 pfet_06v0 ad=2.2p pd=10.879999u as=1.3p ps=5.52u w=5u l=0.7u
D3 DVSS.t190 DVDD.t162 diode_nd2ps_06v0 pj=82u area=40p
X136 DVSS.t15 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.t90 DVDD.t89 DVSS.t14 nfet_06v0 ad=12.999999p pd=50.52u as=12.999999p ps=50.52u w=50u l=0.7u
X137 DVDD.t138 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.t91 DVSS.t13 DVSS.t12 nfet_06v0 ad=12.999999p pd=50.52u as=12.999999p ps=50.52u w=50u l=0.7u
X138 DVDD.t105 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.t92 DVSS.t11 DVSS.t10 nfet_06v0 ad=12.999999p pd=50.52u as=12.999999p ps=50.52u w=50u l=0.7u
X139 DVDD.t149 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.t93 DVSS.t9 DVSS.t8 nfet_06v0 ad=12.999999p pd=50.52u as=12.999999p ps=50.52u w=50u l=0.7u
X140 DVDD.t83 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.t94 DVSS.t7 DVSS.t6 nfet_06v0 ad=12.999999p pd=50.52u as=12.999999p ps=50.52u w=50u l=0.7u
X141 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/comp018green_esd_rc_v5p0_0.ppolyf_u_CDNS_406619531453_1.MINUS.t0 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/comp018green_esd_rc_v5p0_0.ppolyf_u_CDNS_406619531453_1.PLUS.t1 DVDD.t12 ppolyf_u r_width=0.8u r_length=63.854996u
X142 DVSS.t5 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.t95 DVDD.t113 DVSS.t4 nfet_06v0 ad=12.999999p pd=50.52u as=12.999999p ps=50.52u w=50u l=0.7u
X143 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_1.D.t0 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531459_0.D.t10 DVSS.t183 DVSS.t182 nfet_06v0 ad=1.3p pd=5.52u as=1.3p ps=5.52u w=5u l=0.7u
X144 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_1.D.t3 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531459_0.D.t11 DVDD.t65 DVDD.t64 pfet_06v0 ad=2.2p pd=10.879999u as=1.3p ps=5.52u w=5u l=0.7u
X145 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.t14 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_1.D.t32 DVDD.t74 DVDD.t73 pfet_06v0 ad=1.3p pd=5.52u as=1.3p ps=5.52u w=5u l=0.7u
X146 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.t11 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_1.D.t33 DVDD.t33 DVDD.t32 pfet_06v0 ad=1.3p pd=5.52u as=1.3p ps=5.52u w=5u l=0.7u
X147 DVSS.t3 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.t96 DVDD.t146 DVSS.t2 nfet_06v0 ad=12.999999p pd=50.52u as=12.999999p ps=50.52u w=50u l=0.7u
R0 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/comp018green_esd_rc_v5p0_0.ppolyf_u_CDNS_406619531453_5.MINUS GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/comp018green_esd_rc_v5p0_0.ppolyf_u_CDNS_406619531453_5.MINUS.t0 11.0117
R1 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/comp018green_esd_rc_v5p0_0.ppolyf_u_CDNS_406619531453_5.MINUS GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/comp018green_esd_rc_v5p0_0.ppolyf_u_CDNS_406619531453_5.MINUS.t1 11.0117
R2 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/comp018green_esd_rc_v5p0_0.ppolyf_u_CDNS_406619531453_5.PLUS.t0 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/comp018green_esd_rc_v5p0_0.ppolyf_u_CDNS_406619531453_5.PLUS.t1 22.3936
R3 DVDD.n546 DVDD.n545 33140.3
R4 DVDD.n5528 DVDD.n545 33140.3
R5 DVDD.n5528 DVDD.n5527 33140.3
R6 DVDD.n5527 DVDD.n546 33140.3
R7 DVDD.n3846 DVDD.n3831 12187
R8 DVDD.n3846 DVDD.n3845 12187
R9 DVDD.n3845 DVDD.n3844 12187
R10 DVDD.n3844 DVDD.n3831 12187
R11 DVDD.n5710 DVDD.t17 286
R12 DVDD.n5481 DVDD.t2 286
R13 DVDD.t64 DVDD.t19 270.481
R14 DVDD.t23 DVDD.t17 158.649
R15 DVDD.t57 DVDD.t23 158.649
R16 DVDD.t32 DVDD.t57 158.649
R17 DVDD.t21 DVDD.t32 158.649
R18 DVDD.t42 DVDD.t21 158.649
R19 DVDD.t68 DVDD.t42 158.649
R20 DVDD.t10 DVDD.t68 158.649
R21 DVDD.t25 DVDD.t10 158.649
R22 DVDD.t59 DVDD.t25 158.649
R23 DVDD.t30 DVDD.t59 158.649
R24 DVDD.t53 DVDD.t30 158.649
R25 DVDD.t66 DVDD.t53 158.649
R26 DVDD.t28 DVDD.t66 158.649
R27 DVDD.t50 DVDD.t28 158.649
R28 DVDD.t13 DVDD.t50 158.649
R29 DVDD.t40 DVDD.t15 158.649
R30 DVDD.t55 DVDD.t40 158.649
R31 DVDD.t73 DVDD.t55 158.649
R32 DVDD.t48 DVDD.t73 158.649
R33 DVDD.t34 DVDD.t48 158.649
R34 DVDD.t44 DVDD.t34 158.649
R35 DVDD.t19 DVDD.t44 158.649
R36 DVDD.t36 DVDD.t64 158.649
R37 DVDD.t38 DVDD.t36 158.649
R38 DVDD.t46 DVDD.t38 158.649
R39 DVDD.t62 DVDD.t46 158.649
R40 DVDD.t0 DVDD.t62 158.649
R41 DVDD.t2 DVDD.t0 158.649
R42 DVDD.t15 DVDD.n5480 102.731
R43 DVDD.n5480 DVDD.t13 55.9173
R44 DVDD.n5876 DVDD.n5875 29.1205
R45 DVDD.n5948 DVDD.n31 11.1794
R46 DVDD.n5877 DVDD.n102 11.1794
R47 DVDD DVDD.t5 11.0117
R48 DVDD.n5952 DVDD.n5951 8.60804
R49 DVDD.n5872 DVDD.n5833 7.6305
R50 DVDD.n5879 DVDD.n103 7.6305
R51 DVDD.n5948 DVDD.n45 7.54986
R52 DVDD.n5942 DVDD.n5941 7.54986
R53 DVDD.n5941 DVDD.n5940 7.54986
R54 DVDD.n5934 DVDD.n56 7.54986
R55 DVDD.n5934 DVDD.n5933 7.54986
R56 DVDD.n5932 DVDD.n60 7.54986
R57 DVDD.n5926 DVDD.n5925 7.54986
R58 DVDD.n5925 DVDD.n5924 7.54986
R59 DVDD.n5918 DVDD.n70 7.54986
R60 DVDD.n5918 DVDD.n5917 7.54986
R61 DVDD.n5916 DVDD.n74 7.54986
R62 DVDD.n5910 DVDD.n5909 7.54986
R63 DVDD.n5909 DVDD.n5908 7.54986
R64 DVDD.n5902 DVDD.n84 7.54986
R65 DVDD.n5902 DVDD.n5901 7.54986
R66 DVDD.n5900 DVDD.n88 7.54986
R67 DVDD.n5894 DVDD.n5893 7.54986
R68 DVDD.n5893 DVDD.n5892 7.54986
R69 DVDD.n5886 DVDD.n98 7.54986
R70 DVDD.n5886 DVDD.n5885 7.54986
R71 DVDD.n5884 DVDD.n102 7.54986
R72 DVDD.n4228 DVDD.n4226 7.2805
R73 DVDD.n4232 DVDD.n4230 7.2805
R74 DVDD.n4236 DVDD.n4224 7.2805
R75 DVDD.n4240 DVDD.n4238 7.2805
R76 DVDD.n4244 DVDD.n4222 7.2805
R77 DVDD.n4248 DVDD.n4246 7.2805
R78 DVDD.n4252 DVDD.n4220 7.2805
R79 DVDD.n4255 DVDD.n4254 7.2805
R80 DVDD.n4259 DVDD.n4258 7.2805
R81 DVDD.n4317 DVDD.n4316 7.2805
R82 DVDD.n4314 DVDD.n4262 7.2805
R83 DVDD.n4310 DVDD.n4309 7.2805
R84 DVDD.n4307 DVDD.n4265 7.2805
R85 DVDD.n4303 DVDD.n4302 7.2805
R86 DVDD.n4300 DVDD.n4268 7.2805
R87 DVDD.n4296 DVDD.n4295 7.2805
R88 DVDD.n4293 DVDD.n4271 7.2805
R89 DVDD.n4289 DVDD.n4288 7.2805
R90 DVDD.n4286 DVDD.n4274 7.2805
R91 DVDD.n4282 DVDD.n4281 7.2805
R92 DVDD.n4279 DVDD.n4277 7.2805
R93 DVDD.n4681 DVDD.n4680 7.2805
R94 DVDD.n4678 DVDD.n3380 7.2805
R95 DVDD.n4674 DVDD.n4673 7.2805
R96 DVDD.n4671 DVDD.n3383 7.2805
R97 DVDD.n4667 DVDD.n4666 7.2805
R98 DVDD.n4664 DVDD.n3386 7.2805
R99 DVDD.n4660 DVDD.n4659 7.2805
R100 DVDD.n4657 DVDD.n3389 7.2805
R101 DVDD.n4653 DVDD.n4652 7.2805
R102 DVDD.n4650 DVDD.n3392 7.2805
R103 DVDD.n4646 DVDD.n4645 7.2805
R104 DVDD.n4643 DVDD.n3396 7.2805
R105 DVDD.n3406 DVDD.n3405 7.2805
R106 DVDD.n4637 DVDD.n4636 7.2805
R107 DVDD.n4634 DVDD.n3408 7.2805
R108 DVDD.n4630 DVDD.n4629 7.2805
R109 DVDD.n4627 DVDD.n3411 7.2805
R110 DVDD.n4623 DVDD.n4622 7.2805
R111 DVDD.n4620 DVDD.n3414 7.2805
R112 DVDD.n4616 DVDD.n4615 7.2805
R113 DVDD.n4613 DVDD.n3417 7.2805
R114 DVDD.n4609 DVDD.n4608 7.2805
R115 DVDD.n4606 DVDD.n3420 7.2805
R116 DVDD.n4602 DVDD.n4601 7.2805
R117 DVDD.n4599 DVDD.n3424 7.2805
R118 DVDD.n4595 DVDD.n4594 7.2805
R119 DVDD.n4592 DVDD.n4548 7.2805
R120 DVDD.n4588 DVDD.n4587 7.2805
R121 DVDD.n4585 DVDD.n4551 7.2805
R122 DVDD.n4581 DVDD.n4580 7.2805
R123 DVDD.n4578 DVDD.n4554 7.2805
R124 DVDD.n4574 DVDD.n4573 7.2805
R125 DVDD.n4571 DVDD.n4557 7.2805
R126 DVDD.n4567 DVDD.n4566 7.2805
R127 DVDD.n4564 DVDD.n4561 7.2805
R128 DVDD.n5981 DVDD.n30 7.2805
R129 DVDD.n5979 DVDD.n5978 7.2805
R130 DVDD.n5976 DVDD.n33 7.2805
R131 DVDD.n5972 DVDD.n5971 7.2805
R132 DVDD.n5969 DVDD.n36 7.2805
R133 DVDD.n5965 DVDD.n5964 7.2805
R134 DVDD.n5962 DVDD.n39 7.2805
R135 DVDD.n5958 DVDD.n5957 7.2805
R136 DVDD.n5955 DVDD.n42 7.2805
R137 DVDD.n5949 DVDD.n44 7.2805
R138 DVDD.n50 DVDD.n44 7.2805
R139 DVDD.n51 DVDD.n50 7.2805
R140 DVDD.n52 DVDD.n51 7.2805
R141 DVDD.n5837 DVDD.n52 7.2805
R142 DVDD.n5837 DVDD.n57 7.2805
R143 DVDD.n58 DVDD.n57 7.2805
R144 DVDD.n59 DVDD.n58 7.2805
R145 DVDD.n5842 DVDD.n59 7.2805
R146 DVDD.n5842 DVDD.n64 7.2805
R147 DVDD.n65 DVDD.n64 7.2805
R148 DVDD.n66 DVDD.n65 7.2805
R149 DVDD.n5847 DVDD.n66 7.2805
R150 DVDD.n5847 DVDD.n71 7.2805
R151 DVDD.n72 DVDD.n71 7.2805
R152 DVDD.n73 DVDD.n72 7.2805
R153 DVDD.n5852 DVDD.n73 7.2805
R154 DVDD.n5852 DVDD.n78 7.2805
R155 DVDD.n79 DVDD.n78 7.2805
R156 DVDD.n80 DVDD.n79 7.2805
R157 DVDD.n5857 DVDD.n80 7.2805
R158 DVDD.n5857 DVDD.n85 7.2805
R159 DVDD.n86 DVDD.n85 7.2805
R160 DVDD.n87 DVDD.n86 7.2805
R161 DVDD.n5862 DVDD.n87 7.2805
R162 DVDD.n5862 DVDD.n92 7.2805
R163 DVDD.n93 DVDD.n92 7.2805
R164 DVDD.n94 DVDD.n93 7.2805
R165 DVDD.n5867 DVDD.n94 7.2805
R166 DVDD.n5867 DVDD.n99 7.2805
R167 DVDD.n100 DVDD.n99 7.2805
R168 DVDD.n101 DVDD.n100 7.2805
R169 DVDD.n5872 DVDD.n101 7.2805
R170 DVDD.n5947 DVDD.n46 7.2805
R171 DVDD.n5943 DVDD.n46 7.2805
R172 DVDD.n5943 DVDD.n49 7.2805
R173 DVDD.n5939 DVDD.n49 7.2805
R174 DVDD.n5939 DVDD.n53 7.2805
R175 DVDD.n5935 DVDD.n53 7.2805
R176 DVDD.n5935 DVDD.n55 7.2805
R177 DVDD.n5931 DVDD.n55 7.2805
R178 DVDD.n5931 DVDD.n61 7.2805
R179 DVDD.n5927 DVDD.n61 7.2805
R180 DVDD.n5927 DVDD.n63 7.2805
R181 DVDD.n5923 DVDD.n63 7.2805
R182 DVDD.n5923 DVDD.n67 7.2805
R183 DVDD.n5919 DVDD.n67 7.2805
R184 DVDD.n5919 DVDD.n69 7.2805
R185 DVDD.n5915 DVDD.n69 7.2805
R186 DVDD.n5915 DVDD.n75 7.2805
R187 DVDD.n5911 DVDD.n75 7.2805
R188 DVDD.n5911 DVDD.n77 7.2805
R189 DVDD.n5907 DVDD.n77 7.2805
R190 DVDD.n5907 DVDD.n81 7.2805
R191 DVDD.n5903 DVDD.n81 7.2805
R192 DVDD.n5903 DVDD.n83 7.2805
R193 DVDD.n5899 DVDD.n83 7.2805
R194 DVDD.n5899 DVDD.n89 7.2805
R195 DVDD.n5895 DVDD.n89 7.2805
R196 DVDD.n5895 DVDD.n91 7.2805
R197 DVDD.n5891 DVDD.n91 7.2805
R198 DVDD.n5891 DVDD.n95 7.2805
R199 DVDD.n5887 DVDD.n95 7.2805
R200 DVDD.n5887 DVDD.n97 7.2805
R201 DVDD.n5883 DVDD.n97 7.2805
R202 DVDD.n5883 DVDD.n103 7.2805
R203 DVDD.n4812 DVDD.n105 7.2805
R204 DVDD.n4816 DVDD.n4815 7.2805
R205 DVDD.n4820 DVDD.n4819 7.2805
R206 DVDD.n4824 DVDD.n4823 7.2805
R207 DVDD.n4828 DVDD.n4827 7.2805
R208 DVDD.n4832 DVDD.n4831 7.2805
R209 DVDD.n4836 DVDD.n4835 7.2805
R210 DVDD.n4840 DVDD.n4839 7.2805
R211 DVDD.n4844 DVDD.n4843 7.2805
R212 DVDD.n4784 DVDD.n4783 7.2805
R213 DVDD.n4780 DVDD.n4779 7.2805
R214 DVDD.n4776 DVDD.n4775 7.2805
R215 DVDD.n4772 DVDD.n4771 7.2805
R216 DVDD.n4768 DVDD.n4767 7.2805
R217 DVDD.n4764 DVDD.n4763 7.2805
R218 DVDD.n4760 DVDD.n4759 7.2805
R219 DVDD.n4756 DVDD.n4755 7.2805
R220 DVDD.n4752 DVDD.n4751 7.2805
R221 DVDD.n4748 DVDD.n4747 7.2805
R222 DVDD.n4744 DVDD.n4743 7.2805
R223 DVDD.n3353 DVDD.n3352 7.2805
R224 DVDD.n3350 DVDD.n3349 7.2805
R225 DVDD.n3346 DVDD.n3345 7.2805
R226 DVDD.n3342 DVDD.n3341 7.2805
R227 DVDD.n3338 DVDD.n3337 7.2805
R228 DVDD.n3334 DVDD.n3333 7.2805
R229 DVDD.n3330 DVDD.n3329 7.2805
R230 DVDD.n3326 DVDD.n3325 7.2805
R231 DVDD.n3322 DVDD.n3321 7.2805
R232 DVDD.n3318 DVDD.n3317 7.2805
R233 DVDD.n3314 DVDD.n3313 7.2805
R234 DVDD.n3309 DVDD.n3308 7.2805
R235 DVDD.n3304 DVDD.n3258 7.2805
R236 DVDD.n3301 DVDD.n3300 7.2805
R237 DVDD.n3297 DVDD.n3296 7.2805
R238 DVDD.n3293 DVDD.n3292 7.2805
R239 DVDD.n3289 DVDD.n3288 7.2805
R240 DVDD.n3285 DVDD.n3284 7.2805
R241 DVDD.n3281 DVDD.n3280 7.2805
R242 DVDD.n3277 DVDD.n3276 7.2805
R243 DVDD.n3273 DVDD.n3272 7.2805
R244 DVDD.n3269 DVDD.n3268 7.2805
R245 DVDD.n3265 DVDD.n3264 7.2805
R246 DVDD.n3261 DVDD.n3260 7.2805
R247 DVDD.n5762 DVDD.n5761 7.2805
R248 DVDD.n5766 DVDD.n5765 7.2805
R249 DVDD.n5770 DVDD.n5769 7.2805
R250 DVDD.n5774 DVDD.n5773 7.2805
R251 DVDD.n5778 DVDD.n5777 7.2805
R252 DVDD.n5782 DVDD.n5781 7.2805
R253 DVDD.n5786 DVDD.n5785 7.2805
R254 DVDD.n5790 DVDD.n5789 7.2805
R255 DVDD.n5794 DVDD.n5793 7.2805
R256 DVDD.n5798 DVDD.n5797 7.2805
R257 DVDD.n5802 DVDD.n5801 7.2805
R258 DVDD.n5805 DVDD.n5804 7.2805
R259 DVDD.n5812 DVDD.n5811 7.2805
R260 DVDD.n5816 DVDD.n5815 7.2805
R261 DVDD.n5820 DVDD.n5819 7.2805
R262 DVDD.n5824 DVDD.n5823 7.2805
R263 DVDD.n5828 DVDD.n5827 7.2805
R264 DVDD.n5830 DVDD.n167 7.2805
R265 DVDD.t61 DVDD.n5932 6.96914
R266 DVDD.t12 DVDD.n88 6.96914
R267 DVDD.n5875 DVDD.n5874 6.43815
R268 DVDD.t72 DVDD.n5916 6.38842
R269 DVDD.t52 DVDD.n74 6.38842
R270 DVDD.n5881 DVDD.n103 6.3005
R271 DVDD.n103 DVDD.n102 6.3005
R272 DVDD.n5883 DVDD.n5882 6.3005
R273 DVDD.n5884 DVDD.n5883 6.3005
R274 DVDD.n97 DVDD.n96 6.3005
R275 DVDD.n5885 DVDD.n97 6.3005
R276 DVDD.n5888 DVDD.n5887 6.3005
R277 DVDD.n5887 DVDD.n5886 6.3005
R278 DVDD.n5889 DVDD.n95 6.3005
R279 DVDD.n98 DVDD.n95 6.3005
R280 DVDD.n5891 DVDD.n5890 6.3005
R281 DVDD.n5892 DVDD.n5891 6.3005
R282 DVDD.n91 DVDD.n90 6.3005
R283 DVDD.n5893 DVDD.n91 6.3005
R284 DVDD.n5896 DVDD.n5895 6.3005
R285 DVDD.n5895 DVDD.n5894 6.3005
R286 DVDD.n5897 DVDD.n89 6.3005
R287 DVDD.n89 DVDD.n88 6.3005
R288 DVDD.n5899 DVDD.n5898 6.3005
R289 DVDD.n5900 DVDD.n5899 6.3005
R290 DVDD.n83 DVDD.n82 6.3005
R291 DVDD.n5901 DVDD.n83 6.3005
R292 DVDD.n5904 DVDD.n5903 6.3005
R293 DVDD.n5903 DVDD.n5902 6.3005
R294 DVDD.n5905 DVDD.n81 6.3005
R295 DVDD.n84 DVDD.n81 6.3005
R296 DVDD.n5907 DVDD.n5906 6.3005
R297 DVDD.n5908 DVDD.n5907 6.3005
R298 DVDD.n77 DVDD.n76 6.3005
R299 DVDD.n5909 DVDD.n77 6.3005
R300 DVDD.n5912 DVDD.n5911 6.3005
R301 DVDD.n5911 DVDD.n5910 6.3005
R302 DVDD.n5913 DVDD.n75 6.3005
R303 DVDD.n75 DVDD.n74 6.3005
R304 DVDD.n5915 DVDD.n5914 6.3005
R305 DVDD.n5916 DVDD.n5915 6.3005
R306 DVDD.n69 DVDD.n68 6.3005
R307 DVDD.n5917 DVDD.n69 6.3005
R308 DVDD.n5920 DVDD.n5919 6.3005
R309 DVDD.n5919 DVDD.n5918 6.3005
R310 DVDD.n5921 DVDD.n67 6.3005
R311 DVDD.n70 DVDD.n67 6.3005
R312 DVDD.n5923 DVDD.n5922 6.3005
R313 DVDD.n5924 DVDD.n5923 6.3005
R314 DVDD.n63 DVDD.n62 6.3005
R315 DVDD.n5925 DVDD.n63 6.3005
R316 DVDD.n5928 DVDD.n5927 6.3005
R317 DVDD.n5927 DVDD.n5926 6.3005
R318 DVDD.n5929 DVDD.n61 6.3005
R319 DVDD.n61 DVDD.n60 6.3005
R320 DVDD.n5931 DVDD.n5930 6.3005
R321 DVDD.n5932 DVDD.n5931 6.3005
R322 DVDD.n55 DVDD.n54 6.3005
R323 DVDD.n5933 DVDD.n55 6.3005
R324 DVDD.n5936 DVDD.n5935 6.3005
R325 DVDD.n5935 DVDD.n5934 6.3005
R326 DVDD.n5937 DVDD.n53 6.3005
R327 DVDD.n56 DVDD.n53 6.3005
R328 DVDD.n5939 DVDD.n5938 6.3005
R329 DVDD.n5940 DVDD.n5939 6.3005
R330 DVDD.n49 DVDD.n48 6.3005
R331 DVDD.n5941 DVDD.n49 6.3005
R332 DVDD.n5944 DVDD.n5943 6.3005
R333 DVDD.n5943 DVDD.n5942 6.3005
R334 DVDD.n5945 DVDD.n46 6.3005
R335 DVDD.n46 DVDD.n45 6.3005
R336 DVDD.n5947 DVDD.n5946 6.3005
R337 DVDD.n5948 DVDD.n5947 6.3005
R338 DVDD.n5877 DVDD.n5876 6.3005
R339 DVDD.n5877 DVDD.n167 6.3005
R340 DVDD.n5831 DVDD.n5830 6.3005
R341 DVDD.n5829 DVDD.n5828 6.3005
R342 DVDD.n5827 DVDD.n5826 6.3005
R343 DVDD.n5825 DVDD.n5824 6.3005
R344 DVDD.n5823 DVDD.n5822 6.3005
R345 DVDD.n5821 DVDD.n5820 6.3005
R346 DVDD.n5819 DVDD.n5818 6.3005
R347 DVDD.n5817 DVDD.n5816 6.3005
R348 DVDD.n5815 DVDD.n5814 6.3005
R349 DVDD.n5813 DVDD.n5812 6.3005
R350 DVDD.n5811 DVDD.n5810 6.3005
R351 DVDD.n5804 DVDD.n169 6.3005
R352 DVDD.n5806 DVDD.n5805 6.3005
R353 DVDD.n5803 DVDD.n5802 6.3005
R354 DVDD.n5801 DVDD.n5800 6.3005
R355 DVDD.n5799 DVDD.n5798 6.3005
R356 DVDD.n5797 DVDD.n5796 6.3005
R357 DVDD.n5795 DVDD.n5794 6.3005
R358 DVDD.n5793 DVDD.n5792 6.3005
R359 DVDD.n5791 DVDD.n5790 6.3005
R360 DVDD.n5789 DVDD.n5788 6.3005
R361 DVDD.n5787 DVDD.n5786 6.3005
R362 DVDD.n5785 DVDD.n5784 6.3005
R363 DVDD.n5783 DVDD.n5782 6.3005
R364 DVDD.n5781 DVDD.n5780 6.3005
R365 DVDD.n5779 DVDD.n5778 6.3005
R366 DVDD.n5777 DVDD.n5776 6.3005
R367 DVDD.n5775 DVDD.n5774 6.3005
R368 DVDD.n5773 DVDD.n5772 6.3005
R369 DVDD.n5771 DVDD.n5770 6.3005
R370 DVDD.n5769 DVDD.n5768 6.3005
R371 DVDD.n5767 DVDD.n5766 6.3005
R372 DVDD.n5765 DVDD.n5764 6.3005
R373 DVDD.n5763 DVDD.n5762 6.3005
R374 DVDD.n5761 DVDD.n5760 6.3005
R375 DVDD.n3260 DVDD.n173 6.3005
R376 DVDD.n3262 DVDD.n3261 6.3005
R377 DVDD.n3264 DVDD.n3263 6.3005
R378 DVDD.n3266 DVDD.n3265 6.3005
R379 DVDD.n3268 DVDD.n3267 6.3005
R380 DVDD.n3270 DVDD.n3269 6.3005
R381 DVDD.n3272 DVDD.n3271 6.3005
R382 DVDD.n3274 DVDD.n3273 6.3005
R383 DVDD.n3276 DVDD.n3275 6.3005
R384 DVDD.n3278 DVDD.n3277 6.3005
R385 DVDD.n3280 DVDD.n3279 6.3005
R386 DVDD.n3282 DVDD.n3281 6.3005
R387 DVDD.n3284 DVDD.n3283 6.3005
R388 DVDD.n3286 DVDD.n3285 6.3005
R389 DVDD.n3288 DVDD.n3287 6.3005
R390 DVDD.n3290 DVDD.n3289 6.3005
R391 DVDD.n3292 DVDD.n3291 6.3005
R392 DVDD.n3294 DVDD.n3293 6.3005
R393 DVDD.n3296 DVDD.n3295 6.3005
R394 DVDD.n3298 DVDD.n3297 6.3005
R395 DVDD.n3300 DVDD.n3299 6.3005
R396 DVDD.n3302 DVDD.n3301 6.3005
R397 DVDD.n3305 DVDD.n3304 6.3005
R398 DVDD.n3306 DVDD.n3258 6.3005
R399 DVDD.n3308 DVDD.n3307 6.3005
R400 DVDD.n3310 DVDD.n3309 6.3005
R401 DVDD.n3313 DVDD.n3312 6.3005
R402 DVDD.n3315 DVDD.n3314 6.3005
R403 DVDD.n3317 DVDD.n3316 6.3005
R404 DVDD.n3319 DVDD.n3318 6.3005
R405 DVDD.n3321 DVDD.n3320 6.3005
R406 DVDD.n3323 DVDD.n3322 6.3005
R407 DVDD.n3325 DVDD.n3324 6.3005
R408 DVDD.n3327 DVDD.n3326 6.3005
R409 DVDD.n3329 DVDD.n3328 6.3005
R410 DVDD.n3331 DVDD.n3330 6.3005
R411 DVDD.n3333 DVDD.n3332 6.3005
R412 DVDD.n3335 DVDD.n3334 6.3005
R413 DVDD.n3337 DVDD.n3336 6.3005
R414 DVDD.n3339 DVDD.n3338 6.3005
R415 DVDD.n3341 DVDD.n3340 6.3005
R416 DVDD.n3343 DVDD.n3342 6.3005
R417 DVDD.n3345 DVDD.n3344 6.3005
R418 DVDD.n3347 DVDD.n3346 6.3005
R419 DVDD.n3349 DVDD.n3348 6.3005
R420 DVDD.n3351 DVDD.n3350 6.3005
R421 DVDD.n3354 DVDD.n3353 6.3005
R422 DVDD.n3352 DVDD.n3255 6.3005
R423 DVDD.n4743 DVDD.n4742 6.3005
R424 DVDD.n4745 DVDD.n4744 6.3005
R425 DVDD.n4747 DVDD.n4746 6.3005
R426 DVDD.n4749 DVDD.n4748 6.3005
R427 DVDD.n4751 DVDD.n4750 6.3005
R428 DVDD.n4753 DVDD.n4752 6.3005
R429 DVDD.n4755 DVDD.n4754 6.3005
R430 DVDD.n4757 DVDD.n4756 6.3005
R431 DVDD.n4759 DVDD.n4758 6.3005
R432 DVDD.n4761 DVDD.n4760 6.3005
R433 DVDD.n4763 DVDD.n4762 6.3005
R434 DVDD.n4765 DVDD.n4764 6.3005
R435 DVDD.n4767 DVDD.n4766 6.3005
R436 DVDD.n4769 DVDD.n4768 6.3005
R437 DVDD.n4771 DVDD.n4770 6.3005
R438 DVDD.n4773 DVDD.n4772 6.3005
R439 DVDD.n4775 DVDD.n4774 6.3005
R440 DVDD.n4777 DVDD.n4776 6.3005
R441 DVDD.n4779 DVDD.n4778 6.3005
R442 DVDD.n4781 DVDD.n4780 6.3005
R443 DVDD.n4783 DVDD.n4782 6.3005
R444 DVDD.n4785 DVDD.n4784 6.3005
R445 DVDD.n4845 DVDD.n4844 6.3005
R446 DVDD.n4843 DVDD.n4842 6.3005
R447 DVDD.n4841 DVDD.n4840 6.3005
R448 DVDD.n4839 DVDD.n4838 6.3005
R449 DVDD.n4837 DVDD.n4836 6.3005
R450 DVDD.n4835 DVDD.n4834 6.3005
R451 DVDD.n4833 DVDD.n4832 6.3005
R452 DVDD.n4831 DVDD.n4830 6.3005
R453 DVDD.n4829 DVDD.n4828 6.3005
R454 DVDD.n4827 DVDD.n4826 6.3005
R455 DVDD.n4825 DVDD.n4824 6.3005
R456 DVDD.n4823 DVDD.n4822 6.3005
R457 DVDD.n4821 DVDD.n4820 6.3005
R458 DVDD.n4819 DVDD.n4818 6.3005
R459 DVDD.n4817 DVDD.n4816 6.3005
R460 DVDD.n4815 DVDD.n4814 6.3005
R461 DVDD.n4813 DVDD.n4812 6.3005
R462 DVDD.n105 DVDD.n104 6.3005
R463 DVDD.n5880 DVDD.n5879 6.3005
R464 DVDD.n5874 DVDD.n5833 6.3005
R465 DVDD.n5950 DVDD.n5949 6.3005
R466 DVDD.n5949 DVDD.n5948 6.3005
R467 DVDD.n44 DVDD.n43 6.3005
R468 DVDD.n45 DVDD.n44 6.3005
R469 DVDD.n5834 DVDD.n50 6.3005
R470 DVDD.n5942 DVDD.n50 6.3005
R471 DVDD.n5835 DVDD.n51 6.3005
R472 DVDD.n5941 DVDD.n51 6.3005
R473 DVDD.n5836 DVDD.n52 6.3005
R474 DVDD.n5940 DVDD.n52 6.3005
R475 DVDD.n5838 DVDD.n5837 6.3005
R476 DVDD.n5837 DVDD.n56 6.3005
R477 DVDD.n5839 DVDD.n57 6.3005
R478 DVDD.n5934 DVDD.n57 6.3005
R479 DVDD.n5840 DVDD.n58 6.3005
R480 DVDD.n5933 DVDD.n58 6.3005
R481 DVDD.n5841 DVDD.n59 6.3005
R482 DVDD.n5932 DVDD.n59 6.3005
R483 DVDD.n5843 DVDD.n5842 6.3005
R484 DVDD.n5842 DVDD.n60 6.3005
R485 DVDD.n5844 DVDD.n64 6.3005
R486 DVDD.n5926 DVDD.n64 6.3005
R487 DVDD.n5845 DVDD.n65 6.3005
R488 DVDD.n5925 DVDD.n65 6.3005
R489 DVDD.n5846 DVDD.n66 6.3005
R490 DVDD.n5924 DVDD.n66 6.3005
R491 DVDD.n5848 DVDD.n5847 6.3005
R492 DVDD.n5847 DVDD.n70 6.3005
R493 DVDD.n5849 DVDD.n71 6.3005
R494 DVDD.n5918 DVDD.n71 6.3005
R495 DVDD.n5850 DVDD.n72 6.3005
R496 DVDD.n5917 DVDD.n72 6.3005
R497 DVDD.n5851 DVDD.n73 6.3005
R498 DVDD.n5916 DVDD.n73 6.3005
R499 DVDD.n5853 DVDD.n5852 6.3005
R500 DVDD.n5852 DVDD.n74 6.3005
R501 DVDD.n5854 DVDD.n78 6.3005
R502 DVDD.n5910 DVDD.n78 6.3005
R503 DVDD.n5855 DVDD.n79 6.3005
R504 DVDD.n5909 DVDD.n79 6.3005
R505 DVDD.n5856 DVDD.n80 6.3005
R506 DVDD.n5908 DVDD.n80 6.3005
R507 DVDD.n5858 DVDD.n5857 6.3005
R508 DVDD.n5857 DVDD.n84 6.3005
R509 DVDD.n5859 DVDD.n85 6.3005
R510 DVDD.n5902 DVDD.n85 6.3005
R511 DVDD.n5860 DVDD.n86 6.3005
R512 DVDD.n5901 DVDD.n86 6.3005
R513 DVDD.n5861 DVDD.n87 6.3005
R514 DVDD.n5900 DVDD.n87 6.3005
R515 DVDD.n5863 DVDD.n5862 6.3005
R516 DVDD.n5862 DVDD.n88 6.3005
R517 DVDD.n5864 DVDD.n92 6.3005
R518 DVDD.n5894 DVDD.n92 6.3005
R519 DVDD.n5865 DVDD.n93 6.3005
R520 DVDD.n5893 DVDD.n93 6.3005
R521 DVDD.n5866 DVDD.n94 6.3005
R522 DVDD.n5892 DVDD.n94 6.3005
R523 DVDD.n5868 DVDD.n5867 6.3005
R524 DVDD.n5867 DVDD.n98 6.3005
R525 DVDD.n5869 DVDD.n99 6.3005
R526 DVDD.n5886 DVDD.n99 6.3005
R527 DVDD.n5870 DVDD.n100 6.3005
R528 DVDD.n5885 DVDD.n100 6.3005
R529 DVDD.n5871 DVDD.n101 6.3005
R530 DVDD.n5884 DVDD.n101 6.3005
R531 DVDD.n5873 DVDD.n5872 6.3005
R532 DVDD.n5872 DVDD.n102 6.3005
R533 DVDD.n5953 DVDD.n42 6.3005
R534 DVDD.n5955 DVDD.n5954 6.3005
R535 DVDD.n5957 DVDD.n41 6.3005
R536 DVDD.n5959 DVDD.n5958 6.3005
R537 DVDD.n5960 DVDD.n39 6.3005
R538 DVDD.n5962 DVDD.n5961 6.3005
R539 DVDD.n5964 DVDD.n37 6.3005
R540 DVDD.n5966 DVDD.n5965 6.3005
R541 DVDD.n5967 DVDD.n36 6.3005
R542 DVDD.n5969 DVDD.n5968 6.3005
R543 DVDD.n5971 DVDD.n34 6.3005
R544 DVDD.n5973 DVDD.n5972 6.3005
R545 DVDD.n5974 DVDD.n33 6.3005
R546 DVDD.n5976 DVDD.n5975 6.3005
R547 DVDD.n5978 DVDD.n32 6.3005
R548 DVDD.n5979 DVDD.n29 6.3005
R549 DVDD.n5982 DVDD.n5981 6.3005
R550 DVDD.n30 DVDD.n28 6.3005
R551 DVDD.n4562 DVDD.n4561 6.3005
R552 DVDD.n4564 DVDD.n4563 6.3005
R553 DVDD.n4566 DVDD.n4558 6.3005
R554 DVDD.n4568 DVDD.n4567 6.3005
R555 DVDD.n4569 DVDD.n4557 6.3005
R556 DVDD.n4571 DVDD.n4570 6.3005
R557 DVDD.n4573 DVDD.n4555 6.3005
R558 DVDD.n4575 DVDD.n4574 6.3005
R559 DVDD.n4576 DVDD.n4554 6.3005
R560 DVDD.n4578 DVDD.n4577 6.3005
R561 DVDD.n4580 DVDD.n4552 6.3005
R562 DVDD.n4582 DVDD.n4581 6.3005
R563 DVDD.n4583 DVDD.n4551 6.3005
R564 DVDD.n4585 DVDD.n4584 6.3005
R565 DVDD.n4587 DVDD.n4549 6.3005
R566 DVDD.n4589 DVDD.n4588 6.3005
R567 DVDD.n4590 DVDD.n4548 6.3005
R568 DVDD.n4592 DVDD.n4591 6.3005
R569 DVDD.n4594 DVDD.n4546 6.3005
R570 DVDD.n4596 DVDD.n4595 6.3005
R571 DVDD.n4597 DVDD.n3424 6.3005
R572 DVDD.n4599 DVDD.n4598 6.3005
R573 DVDD.n4601 DVDD.n3423 6.3005
R574 DVDD.n4603 DVDD.n4602 6.3005
R575 DVDD.n4604 DVDD.n3420 6.3005
R576 DVDD.n4606 DVDD.n4605 6.3005
R577 DVDD.n4608 DVDD.n3418 6.3005
R578 DVDD.n4610 DVDD.n4609 6.3005
R579 DVDD.n4611 DVDD.n3417 6.3005
R580 DVDD.n4613 DVDD.n4612 6.3005
R581 DVDD.n4615 DVDD.n3415 6.3005
R582 DVDD.n4617 DVDD.n4616 6.3005
R583 DVDD.n4618 DVDD.n3414 6.3005
R584 DVDD.n4620 DVDD.n4619 6.3005
R585 DVDD.n4622 DVDD.n3412 6.3005
R586 DVDD.n4624 DVDD.n4623 6.3005
R587 DVDD.n4625 DVDD.n3411 6.3005
R588 DVDD.n4627 DVDD.n4626 6.3005
R589 DVDD.n4629 DVDD.n3409 6.3005
R590 DVDD.n4631 DVDD.n4630 6.3005
R591 DVDD.n4632 DVDD.n3408 6.3005
R592 DVDD.n4634 DVDD.n4633 6.3005
R593 DVDD.n4636 DVDD.n3403 6.3005
R594 DVDD.n4638 DVDD.n4637 6.3005
R595 DVDD.n3406 DVDD.n3402 6.3005
R596 DVDD.n3405 DVDD.n3398 6.3005
R597 DVDD.n4641 DVDD.n3396 6.3005
R598 DVDD.n4643 DVDD.n4642 6.3005
R599 DVDD.n4645 DVDD.n3395 6.3005
R600 DVDD.n4647 DVDD.n4646 6.3005
R601 DVDD.n4648 DVDD.n3392 6.3005
R602 DVDD.n4650 DVDD.n4649 6.3005
R603 DVDD.n4652 DVDD.n3390 6.3005
R604 DVDD.n4654 DVDD.n4653 6.3005
R605 DVDD.n4655 DVDD.n3389 6.3005
R606 DVDD.n4657 DVDD.n4656 6.3005
R607 DVDD.n4659 DVDD.n3387 6.3005
R608 DVDD.n4661 DVDD.n4660 6.3005
R609 DVDD.n4662 DVDD.n3386 6.3005
R610 DVDD.n4664 DVDD.n4663 6.3005
R611 DVDD.n4666 DVDD.n3384 6.3005
R612 DVDD.n4668 DVDD.n4667 6.3005
R613 DVDD.n4669 DVDD.n3383 6.3005
R614 DVDD.n4671 DVDD.n4670 6.3005
R615 DVDD.n4673 DVDD.n3381 6.3005
R616 DVDD.n4675 DVDD.n4674 6.3005
R617 DVDD.n4676 DVDD.n3380 6.3005
R618 DVDD.n4678 DVDD.n4677 6.3005
R619 DVDD.n4680 DVDD.n3378 6.3005
R620 DVDD.n4682 DVDD.n4681 6.3005
R621 DVDD.n4277 DVDD.n3377 6.3005
R622 DVDD.n4279 DVDD.n4278 6.3005
R623 DVDD.n4281 DVDD.n4275 6.3005
R624 DVDD.n4283 DVDD.n4282 6.3005
R625 DVDD.n4284 DVDD.n4274 6.3005
R626 DVDD.n4286 DVDD.n4285 6.3005
R627 DVDD.n4288 DVDD.n4272 6.3005
R628 DVDD.n4290 DVDD.n4289 6.3005
R629 DVDD.n4291 DVDD.n4271 6.3005
R630 DVDD.n4293 DVDD.n4292 6.3005
R631 DVDD.n4295 DVDD.n4269 6.3005
R632 DVDD.n4297 DVDD.n4296 6.3005
R633 DVDD.n4298 DVDD.n4268 6.3005
R634 DVDD.n4300 DVDD.n4299 6.3005
R635 DVDD.n4302 DVDD.n4266 6.3005
R636 DVDD.n4304 DVDD.n4303 6.3005
R637 DVDD.n4305 DVDD.n4265 6.3005
R638 DVDD.n4307 DVDD.n4306 6.3005
R639 DVDD.n4309 DVDD.n4263 6.3005
R640 DVDD.n4311 DVDD.n4310 6.3005
R641 DVDD.n4312 DVDD.n4262 6.3005
R642 DVDD.n4314 DVDD.n4313 6.3005
R643 DVDD.n4316 DVDD.n4261 6.3005
R644 DVDD.n4318 DVDD.n4317 6.3005
R645 DVDD.n4259 DVDD.n4217 6.3005
R646 DVDD.n4258 DVDD.n4257 6.3005
R647 DVDD.n4256 DVDD.n4255 6.3005
R648 DVDD.n4254 DVDD.n4219 6.3005
R649 DVDD.n4252 DVDD.n4251 6.3005
R650 DVDD.n4250 DVDD.n4220 6.3005
R651 DVDD.n4249 DVDD.n4248 6.3005
R652 DVDD.n4246 DVDD.n4221 6.3005
R653 DVDD.n4244 DVDD.n4243 6.3005
R654 DVDD.n4242 DVDD.n4222 6.3005
R655 DVDD.n4241 DVDD.n4240 6.3005
R656 DVDD.n4238 DVDD.n4223 6.3005
R657 DVDD.n4236 DVDD.n4235 6.3005
R658 DVDD.n4234 DVDD.n4224 6.3005
R659 DVDD.n4233 DVDD.n4232 6.3005
R660 DVDD.n4230 DVDD.n4225 6.3005
R661 DVDD.n4228 DVDD.n4227 6.3005
R662 DVDD.n4226 DVDD.n47 6.3005
R663 DVDD.n4226 DVDD.n31 6.3005
R664 DVDD.t71 DVDD.n60 5.8077
R665 DVDD.t8 DVDD.n5900 5.8077
R666 DVDD.t4 DVDD.n45 5.22698
R667 DVDD.t7 DVDD.n5884 5.22698
R668 DVDD.n5543 DVDD.n541 5.02526
R669 DVDD.n5542 DVDD.n540 5.02526
R670 DVDD.n5541 DVDD.n539 5.02526
R671 DVDD.n5540 DVDD.n538 5.02526
R672 DVDD.n5539 DVDD.n537 5.02526
R673 DVDD.n5538 DVDD.n536 5.02526
R674 DVDD.n5537 DVDD.n535 5.02526
R675 DVDD.n5536 DVDD.n534 5.02526
R676 DVDD.n5535 DVDD.n533 5.02526
R677 DVDD.n5534 DVDD.n532 5.02526
R678 DVDD.n5533 DVDD.n531 5.02526
R679 DVDD.n5532 DVDD.n530 5.02526
R680 DVDD.n5531 DVDD.n529 5.02526
R681 DVDD.n5530 DVDD.n528 5.02526
R682 DVDD.n5563 DVDD.n526 5.02526
R683 DVDD.n2922 DVDD.n2921 5.02526
R684 DVDD.n2757 DVDD.n2604 5.02526
R685 DVDD.n2932 DVDD.n2573 5.02526
R686 DVDD.n2933 DVDD.n1007 5.02526
R687 DVDD.n1011 DVDD.n997 5.02526
R688 DVDD.n5629 DVDD.n443 5.02526
R689 DVDD.n2939 DVDD.n2937 5.02526
R690 DVDD.n2556 DVDD.n2554 5.02526
R691 DVDD.n2538 DVDD.n2536 5.02526
R692 DVDD.n2523 DVDD.n2521 5.02526
R693 DVDD.n2453 DVDD.n411 5.02526
R694 DVDD.n1261 DVDD.n1260 5.02526
R695 DVDD.n2449 DVDD.n2448 5.02526
R696 DVDD.n1249 DVDD.n1247 5.02526
R697 DVDD.n1231 DVDD.n1229 5.02526
R698 DVDD.n2232 DVDD.n381 5.02526
R699 DVDD.n2228 DVDD.n2227 5.02526
R700 DVDD.n1533 DVDD.n1531 5.02526
R701 DVDD.n1519 DVDD.n1517 5.02526
R702 DVDD.n1505 DVDD.n1503 5.02526
R703 DVDD.n1491 DVDD.n1489 5.02526
R704 DVDD.n5649 DVDD.n359 5.02526
R705 DVDD.n2045 DVDD.n1713 5.02526
R706 DVDD.n1735 DVDD.n1733 5.02526
R707 DVDD.n5544 DVDD.n542 5.02526
R708 DVDD.n1740 DVDD.n1739 5.02426
R709 DVDD.n2041 DVDD.n2040 5.02426
R710 DVDD.n2967 DVDD.n2966 5.02426
R711 DVDD.n1485 DVDD.n1484 5.02426
R712 DVDD.n1499 DVDD.n1498 5.02426
R713 DVDD.n1513 DVDD.n1512 5.02426
R714 DVDD.n1527 DVDD.n1526 5.02426
R715 DVDD.n2223 DVDD.n2222 5.02426
R716 DVDD.n2218 DVDD.n920 5.02426
R717 DVDD.n1225 DVDD.n1224 5.02426
R718 DVDD.n1243 DVDD.n1242 5.02426
R719 DVDD.n2444 DVDD.n2443 5.02426
R720 DVDD.n1257 DVDD.n1138 5.02426
R721 DVDD.n2436 DVDD.n950 5.02426
R722 DVDD.n2517 DVDD.n2516 5.02426
R723 DVDD.n2533 DVDD.n2532 5.02426
R724 DVDD.n2551 DVDD.n2550 5.02426
R725 DVDD.n2944 DVDD.n2943 5.02426
R726 DVDD.n5625 DVDD.n5624 5.02426
R727 DVDD.n1009 DVDD.n463 5.02426
R728 DVDD.n5620 DVDD.n5619 5.02426
R729 DVDD.n476 DVDD.n473 5.02426
R730 DVDD.n2763 DVDD.n2762 5.02426
R731 DVDD.n2917 DVDD.n2916 5.02426
R732 DVDD.n2863 DVDD.n2862 5.02426
R733 DVDD.n2770 DVDD.n2766 5.02426
R734 DVDD.n2830 DVDD.n2771 5.02426
R735 DVDD.n2831 DVDD.n2772 5.02426
R736 DVDD.n2832 DVDD.n2773 5.02426
R737 DVDD.n2833 DVDD.n2774 5.02426
R738 DVDD.n2834 DVDD.n2775 5.02426
R739 DVDD.n2835 DVDD.n2776 5.02426
R740 DVDD.n2836 DVDD.n2777 5.02426
R741 DVDD.n2837 DVDD.n2778 5.02426
R742 DVDD.n2838 DVDD.n2779 5.02426
R743 DVDD.n2839 DVDD.n2780 5.02426
R744 DVDD.n2840 DVDD.n2781 5.02426
R745 DVDD.n2842 DVDD.n2841 5.02426
R746 DVDD.n2846 DVDD.n557 5.02426
R747 DVDD.n5518 DVDD.n5517 5.02426
R748 DVDD.n56 DVDD.t70 4.64626
R749 DVDD.n5892 DVDD.t27 4.64626
R750 DVDD.n5984 DVDD.n27 4.5005
R751 DVDD.n4112 DVDD.n3550 4.5005
R752 DVDD.n4116 DVDD.n4115 4.5005
R753 DVDD.n5391 DVDD.n5367 4.5005
R754 DVDD.n5391 DVDD.n606 4.5005
R755 DVDD.n5483 DVDD.n605 4.5005
R756 DVDD.n5494 DVDD.n604 4.5005
R757 DVDD.n5497 DVDD.n5496 4.5005
R758 DVDD.n580 DVDD.n579 4.5005
R759 DVDD.n5498 DVDD.n580 4.5005
R760 DVDD.n5498 DVDD.n5497 4.5005
R761 DVDD.n599 DVDD.n580 4.5005
R762 DVDD.n5497 DVDD.n599 4.5005
R763 DVDD.n5497 DVDD.n597 4.5005
R764 DVDD.n1731 DVDD.n580 4.5005
R765 DVDD.n1732 DVDD.n580 4.5005
R766 DVDD.n1711 DVDD.n580 4.5005
R767 DVDD.n1712 DVDD.n580 4.5005
R768 DVDD.n582 DVDD.n580 4.5005
R769 DVDD.n1371 DVDD.n1370 4.5005
R770 DVDD.n1487 DVDD.n1370 4.5005
R771 DVDD.n1488 DVDD.n1370 4.5005
R772 DVDD.n1501 DVDD.n1370 4.5005
R773 DVDD.n1502 DVDD.n1370 4.5005
R774 DVDD.n1515 DVDD.n1370 4.5005
R775 DVDD.n1516 DVDD.n1370 4.5005
R776 DVDD.n1529 DVDD.n1370 4.5005
R777 DVDD.n1530 DVDD.n1370 4.5005
R778 DVDD.n1387 DVDD.n1370 4.5005
R779 DVDD.n2229 DVDD.n1370 4.5005
R780 DVDD.n2233 DVDD.n1370 4.5005
R781 DVDD.n2231 DVDD.n1093 4.5005
R782 DVDD.n1227 DVDD.n1093 4.5005
R783 DVDD.n1228 DVDD.n1093 4.5005
R784 DVDD.n1245 DVDD.n1093 4.5005
R785 DVDD.n1246 DVDD.n1093 4.5005
R786 DVDD.n1117 DVDD.n1093 4.5005
R787 DVDD.n2450 DVDD.n1093 4.5005
R788 DVDD.n2456 DVDD.n1099 4.5005
R789 DVDD.n1259 DVDD.n1093 4.5005
R790 DVDD.n2456 DVDD.n2455 4.5005
R791 DVDD.n2452 DVDD.n1006 4.5005
R792 DVDD.n2519 DVDD.n1006 4.5005
R793 DVDD.n2520 DVDD.n1006 4.5005
R794 DVDD.n2935 DVDD.n987 4.5005
R795 DVDD.n2535 DVDD.n1006 4.5005
R796 DVDD.n2553 DVDD.n1006 4.5005
R797 DVDD.n2935 DVDD.n992 4.5005
R798 DVDD.n2935 DVDD.n980 4.5005
R799 DVDD.n2936 DVDD.n2935 4.5005
R800 DVDD.n2935 DVDD.n984 4.5005
R801 DVDD.n2935 DVDD.n995 4.5005
R802 DVDD.n2935 DVDD.n983 4.5005
R803 DVDD.n2934 DVDD.n1006 4.5005
R804 DVDD.n2935 DVDD.n2934 4.5005
R805 DVDD.n2931 DVDD.n2930 4.5005
R806 DVDD.n2930 DVDD.n2577 4.5005
R807 DVDD.n2930 DVDD.n2580 4.5005
R808 DVDD.n2930 DVDD.n2576 4.5005
R809 DVDD.n2927 DVDD.n2923 4.5005
R810 DVDD.n2930 DVDD.n2929 4.5005
R811 DVDD.n5984 DVDD.n5983 4.5005
R812 DVDD.n5809 DVDD.n5808 4.5005
R813 DVDD.n5808 DVDD.n5807 4.5005
R814 DVDD.n4544 DVDD.n3421 4.5005
R815 DVDD.n4035 DVDD.n3581 4.5005
R816 DVDD.n4037 DVDD.n3581 4.5005
R817 DVDD.n4035 DVDD.n3580 4.5005
R818 DVDD.n4037 DVDD.n3580 4.5005
R819 DVDD.n4037 DVDD.n3582 4.5005
R820 DVDD.n4037 DVDD.n3579 4.5005
R821 DVDD.n4037 DVDD.n3583 4.5005
R822 DVDD.n4037 DVDD.n3578 4.5005
R823 DVDD.n4035 DVDD.n3584 4.5005
R824 DVDD.n4037 DVDD.n3584 4.5005
R825 DVDD.n4035 DVDD.n3577 4.5005
R826 DVDD.n4037 DVDD.n3577 4.5005
R827 DVDD.n4035 DVDD.n3585 4.5005
R828 DVDD.n4037 DVDD.n3585 4.5005
R829 DVDD.n4037 DVDD.n3576 4.5005
R830 DVDD.n4037 DVDD.n4036 4.5005
R831 DVDD.n4036 DVDD.n4035 4.5005
R832 DVDD.n4035 DVDD.n3576 4.5005
R833 DVDD.n4035 DVDD.n3578 4.5005
R834 DVDD.n4035 DVDD.n3583 4.5005
R835 DVDD.n4035 DVDD.n3579 4.5005
R836 DVDD.n4035 DVDD.n3582 4.5005
R837 DVDD.n5215 DVDD.n5142 4.5005
R838 DVDD.n5215 DVDD.n626 4.5005
R839 DVDD.n5470 DVDD.n5469 4.5005
R840 DVDD.n1597 DVDD.n638 4.5005
R841 DVDD.n2048 DVDD.n1598 4.5005
R842 DVDD.n1709 DVDD.n575 4.5005
R843 DVDD.n2048 DVDD.n576 4.5005
R844 DVDD.n1709 DVDD.n576 4.5005
R845 DVDD.n2048 DVDD.n1596 4.5005
R846 DVDD.n1709 DVDD.n1596 4.5005
R847 DVDD.n1709 DVDD.n1701 4.5005
R848 DVDD.n2048 DVDD.n1606 4.5005
R849 DVDD.n2048 DVDD.n1594 4.5005
R850 DVDD.n2048 DVDD.n2047 4.5005
R851 DVDD.n2048 DVDD.n1593 4.5005
R852 DVDD.n2048 DVDD.n360 4.5005
R853 DVDD.n5647 DVDD.n5646 4.5005
R854 DVDD.n5646 DVDD.n370 4.5005
R855 DVDD.n5646 DVDD.n367 4.5005
R856 DVDD.n5646 DVDD.n372 4.5005
R857 DVDD.n5646 DVDD.n366 4.5005
R858 DVDD.n5646 DVDD.n374 4.5005
R859 DVDD.n5646 DVDD.n365 4.5005
R860 DVDD.n5646 DVDD.n376 4.5005
R861 DVDD.n5646 DVDD.n364 4.5005
R862 DVDD.n5646 DVDD.n378 4.5005
R863 DVDD.n5646 DVDD.n363 4.5005
R864 DVDD.n5646 DVDD.n5645 4.5005
R865 DVDD.n5643 DVDD.n5642 4.5005
R866 DVDD.n5642 DVDD.n389 4.5005
R867 DVDD.n5642 DVDD.n387 4.5005
R868 DVDD.n5642 DVDD.n395 4.5005
R869 DVDD.n5642 DVDD.n386 4.5005
R870 DVDD.n5642 DVDD.n397 4.5005
R871 DVDD.n5642 DVDD.n385 4.5005
R872 DVDD.n5639 DVDD.n400 4.5005
R873 DVDD.n5642 DVDD.n5641 4.5005
R874 DVDD.n5639 DVDD.n5638 4.5005
R875 DVDD.n5636 DVDD.n5635 4.5005
R876 DVDD.n5635 DVDD.n422 4.5005
R877 DVDD.n5635 DVDD.n419 4.5005
R878 DVDD.n5633 DVDD.n435 4.5005
R879 DVDD.n5635 DVDD.n424 4.5005
R880 DVDD.n5635 DVDD.n417 4.5005
R881 DVDD.n5633 DVDD.n439 4.5005
R882 DVDD.n5633 DVDD.n432 4.5005
R883 DVDD.n5633 DVDD.n441 4.5005
R884 DVDD.n5633 DVDD.n431 4.5005
R885 DVDD.n5633 DVDD.n5631 4.5005
R886 DVDD.n5633 DVDD.n430 4.5005
R887 DVDD.n5635 DVDD.n5634 4.5005
R888 DVDD.n5634 DVDD.n5633 4.5005
R889 DVDD.n2754 DVDD.n2611 4.5005
R890 DVDD.n2754 DVDD.n2605 4.5005
R891 DVDD.n2755 DVDD.n2754 4.5005
R892 DVDD.n2754 DVDD.n2608 4.5005
R893 DVDD.n2754 DVDD.n2614 4.5005
R894 DVDD.n2751 DVDD.n527 4.5005
R895 DVDD.n4545 DVDD.n4544 4.5005
R896 DVDD.n5758 DVDD.n172 4.5005
R897 DVDD.n5759 DVDD.n5758 4.5005
R898 DVDD.n3894 DVDD.n3682 4.5005
R899 DVDD.n3893 DVDD.n3892 4.5005
R900 DVDD.n4181 DVDD.n3528 4.5005
R901 DVDD.n4180 DVDD.n4179 4.5005
R902 DVDD.n4178 DVDD.n3529 4.5005
R903 DVDD.n4177 DVDD.n4176 4.5005
R904 DVDD.n4175 DVDD.n3530 4.5005
R905 DVDD.n4174 DVDD.n4173 4.5005
R906 DVDD.n4172 DVDD.n3531 4.5005
R907 DVDD.n4171 DVDD.n4170 4.5005
R908 DVDD.n4169 DVDD.n3532 4.5005
R909 DVDD.n4168 DVDD.n4167 4.5005
R910 DVDD.n4166 DVDD.n3533 4.5005
R911 DVDD.n4165 DVDD.n4164 4.5005
R912 DVDD.n4163 DVDD.n3534 4.5005
R913 DVDD.n4162 DVDD.n4161 4.5005
R914 DVDD.n4160 DVDD.n3535 4.5005
R915 DVDD.n4159 DVDD.n4158 4.5005
R916 DVDD.n4157 DVDD.n3536 4.5005
R917 DVDD.n4156 DVDD.n4155 4.5005
R918 DVDD.n4154 DVDD.n3537 4.5005
R919 DVDD.n4153 DVDD.n4152 4.5005
R920 DVDD.n4151 DVDD.n4150 4.5005
R921 DVDD.n4149 DVDD.n3539 4.5005
R922 DVDD.n4148 DVDD.n4147 4.5005
R923 DVDD.n4146 DVDD.n3540 4.5005
R924 DVDD.n4145 DVDD.n4144 4.5005
R925 DVDD.n4143 DVDD.n3541 4.5005
R926 DVDD.n4142 DVDD.n4141 4.5005
R927 DVDD.n4140 DVDD.n3542 4.5005
R928 DVDD.n4139 DVDD.n4138 4.5005
R929 DVDD.n4137 DVDD.n3543 4.5005
R930 DVDD.n4136 DVDD.n4135 4.5005
R931 DVDD.n4134 DVDD.n3544 4.5005
R932 DVDD.n4133 DVDD.n4132 4.5005
R933 DVDD.n4131 DVDD.n3545 4.5005
R934 DVDD.n4130 DVDD.n4129 4.5005
R935 DVDD.n4128 DVDD.n3546 4.5005
R936 DVDD.n4127 DVDD.n4126 4.5005
R937 DVDD.n4125 DVDD.n3547 4.5005
R938 DVDD.n4124 DVDD.n4123 4.5005
R939 DVDD.n4122 DVDD.n3548 4.5005
R940 DVDD.n4193 DVDD.n4186 4.5005
R941 DVDD.n4196 DVDD.n3527 4.5005
R942 DVDD.n4184 DVDD.n4183 4.5005
R943 DVDD.n3843 DVDD.n3842 4.5005
R944 DVDD.n3842 DVDD.n3841 4.5005
R945 DVDD.n3841 DVDD.n3840 4.5005
R946 DVDD.n3835 DVDD.n3523 4.5005
R947 DVDD.n3841 DVDD.n3523 4.5005
R948 DVDD.n3525 DVDD 4.5005
R949 DVDD.n4198 DVDD.n3525 4.5005
R950 DVDD.n4199 DVDD.n4198 4.5005
R951 DVDD.n4200 DVDD.n4199 4.5005
R952 DVDD.n3679 DVDD 4.5005
R953 DVDD.n3679 DVDD.n3678 4.5005
R954 DVDD.n3678 DVDD.n3677 4.5005
R955 DVDD.n3677 DVDD.n3676 4.5005
R956 DVDD.n3681 DVDD 4.5005
R957 DVDD.n3910 DVDD.n3681 4.5005
R958 DVDD.n3911 DVDD.n3910 4.5005
R959 DVDD.n3912 DVDD.n3911 4.5005
R960 DVDD DVDD.n3902 4.5005
R961 DVDD.n3907 DVDD.n3902 4.5005
R962 DVDD.n3907 DVDD.n3906 4.5005
R963 DVDD.n3906 DVDD.n3668 4.5005
R964 DVDD.n3901 DVDD.n3847 4.5005
R965 DVDD.n3901 DVDD.n3900 4.5005
R966 DVDD.n3897 DVDD.n3849 4.5005
R967 DVDD.n3849 DVDD.n3847 4.5005
R968 DVDD.n3900 DVDD.n3849 4.5005
R969 DVDD.n3899 DVDD.n3897 4.5005
R970 DVDD.n3900 DVDD.n3899 4.5005
R971 DVDD.n4640 DVDD.n3393 4.5005
R972 DVDD.n3627 DVDD.n3611 4.5005
R973 DVDD.n3998 DVDD.n3611 4.5005
R974 DVDD.n4001 DVDD.n3611 4.5005
R975 DVDD.n3998 DVDD.n3610 4.5005
R976 DVDD.n4001 DVDD.n3610 4.5005
R977 DVDD.n3998 DVDD.n3612 4.5005
R978 DVDD.n4001 DVDD.n3612 4.5005
R979 DVDD.n3998 DVDD.n3609 4.5005
R980 DVDD.n4001 DVDD.n3609 4.5005
R981 DVDD.n3998 DVDD.n3613 4.5005
R982 DVDD.n4001 DVDD.n3613 4.5005
R983 DVDD.n3998 DVDD.n3608 4.5005
R984 DVDD.n4001 DVDD.n3608 4.5005
R985 DVDD.n3998 DVDD.n3614 4.5005
R986 DVDD.n4001 DVDD.n3614 4.5005
R987 DVDD.n3998 DVDD.n3607 4.5005
R988 DVDD.n4001 DVDD.n3607 4.5005
R989 DVDD.n3998 DVDD.n3615 4.5005
R990 DVDD.n4001 DVDD.n3615 4.5005
R991 DVDD.n3998 DVDD.n3606 4.5005
R992 DVDD.n4001 DVDD.n3606 4.5005
R993 DVDD.n4001 DVDD.n4000 4.5005
R994 DVDD.n4536 DVDD.n4535 4.5005
R995 DVDD.n4504 DVDD.n4495 4.5005
R996 DVDD.n4507 DVDD.n4506 4.5005
R997 DVDD.n4514 DVDD.n4501 4.5005
R998 DVDD.n4525 DVDD.n4519 4.5005
R999 DVDD.n4523 DVDD.n3150 4.5005
R1000 DVDD.n4870 DVDD.n3147 4.5005
R1001 DVDD.n4876 DVDD.n4875 4.5005
R1002 DVDD.n3140 DVDD.n3139 4.5005
R1003 DVDD.n4884 DVDD.n4883 4.5005
R1004 DVDD.n5756 DVDD.n5755 4.5005
R1005 DVDD.n179 DVDD.n177 4.5005
R1006 DVDD.n3133 DVDD.n3132 4.5005
R1007 DVDD.n4895 DVDD.n3129 4.5005
R1008 DVDD.n4902 DVDD.n4898 4.5005
R1009 DVDD.n5319 DVDD.n4903 4.5005
R1010 DVDD.n5088 DVDD.n4904 4.5005
R1011 DVDD.n5103 DVDD.n4911 4.5005
R1012 DVDD.n5309 DVDD.n4912 4.5005
R1013 DVDD.n5308 DVDD.n4913 4.5005
R1014 DVDD.n5307 DVDD.n4914 4.5005
R1015 DVDD.n5112 DVDD.n4915 4.5005
R1016 DVDD.n5111 DVDD.n5110 4.5005
R1017 DVDD.n5120 DVDD.n4921 4.5005
R1018 DVDD.n5296 DVDD.n4922 4.5005
R1019 DVDD.n5294 DVDD.n4923 4.5005
R1020 DVDD.n5130 DVDD.n4924 4.5005
R1021 DVDD.n5138 DVDD.n4932 4.5005
R1022 DVDD.n5284 DVDD.n4933 4.5005
R1023 DVDD.n5283 DVDD.n4934 4.5005
R1024 DVDD.n5282 DVDD.n4936 4.5005
R1025 DVDD.n5282 DVDD.n4937 4.5005
R1026 DVDD.n5282 DVDD.n5281 4.5005
R1027 DVDD.n5247 DVDD.n4937 4.5005
R1028 DVDD.n5281 DVDD.n5247 4.5005
R1029 DVDD.n4949 DVDD.n4937 4.5005
R1030 DVDD.n5281 DVDD.n4949 4.5005
R1031 DVDD.n5249 DVDD.n4937 4.5005
R1032 DVDD.n5281 DVDD.n5249 4.5005
R1033 DVDD.n4948 DVDD.n4937 4.5005
R1034 DVDD.n5281 DVDD.n4948 4.5005
R1035 DVDD.n5251 DVDD.n4937 4.5005
R1036 DVDD.n5281 DVDD.n5251 4.5005
R1037 DVDD.n4947 DVDD.n4937 4.5005
R1038 DVDD.n5281 DVDD.n4947 4.5005
R1039 DVDD.n5253 DVDD.n4937 4.5005
R1040 DVDD.n5281 DVDD.n5253 4.5005
R1041 DVDD.n4946 DVDD.n4937 4.5005
R1042 DVDD.n5281 DVDD.n4946 4.5005
R1043 DVDD.n5255 DVDD.n4937 4.5005
R1044 DVDD.n5281 DVDD.n5255 4.5005
R1045 DVDD.n4945 DVDD.n4937 4.5005
R1046 DVDD.n5281 DVDD.n4945 4.5005
R1047 DVDD.n5257 DVDD.n4937 4.5005
R1048 DVDD.n5281 DVDD.n5257 4.5005
R1049 DVDD.n4944 DVDD.n4937 4.5005
R1050 DVDD.n5281 DVDD.n4944 4.5005
R1051 DVDD.n5259 DVDD.n4937 4.5005
R1052 DVDD.n5281 DVDD.n5259 4.5005
R1053 DVDD.n4943 DVDD.n4937 4.5005
R1054 DVDD.n5281 DVDD.n4943 4.5005
R1055 DVDD.n5261 DVDD.n4937 4.5005
R1056 DVDD.n5281 DVDD.n5261 4.5005
R1057 DVDD.n4942 DVDD.n4937 4.5005
R1058 DVDD.n5281 DVDD.n4942 4.5005
R1059 DVDD.n5263 DVDD.n4937 4.5005
R1060 DVDD.n5281 DVDD.n5263 4.5005
R1061 DVDD.n4941 DVDD.n4937 4.5005
R1062 DVDD.n5281 DVDD.n4941 4.5005
R1063 DVDD.n5265 DVDD.n4937 4.5005
R1064 DVDD.n5281 DVDD.n5265 4.5005
R1065 DVDD.n4940 DVDD.n4937 4.5005
R1066 DVDD.n5281 DVDD.n4940 4.5005
R1067 DVDD.n5267 DVDD.n4937 4.5005
R1068 DVDD.n5281 DVDD.n5267 4.5005
R1069 DVDD.n4939 DVDD.n4937 4.5005
R1070 DVDD.n5281 DVDD.n4939 4.5005
R1071 DVDD.n5280 DVDD.n4936 4.5005
R1072 DVDD.n5280 DVDD.n4937 4.5005
R1073 DVDD.n5281 DVDD.n5280 4.5005
R1074 DVDD.n5656 DVDD.n296 4.5005
R1075 DVDD.n5655 DVDD.n312 4.5005
R1076 DVDD.n5655 DVDD.n313 4.5005
R1077 DVDD.n5655 DVDD.n5654 4.5005
R1078 DVDD.n328 DVDD.n313 4.5005
R1079 DVDD.n5654 DVDD.n328 4.5005
R1080 DVDD.n325 DVDD.n313 4.5005
R1081 DVDD.n5654 DVDD.n325 4.5005
R1082 DVDD.n330 DVDD.n313 4.5005
R1083 DVDD.n5654 DVDD.n330 4.5005
R1084 DVDD.n5654 DVDD.n324 4.5005
R1085 DVDD.n5654 DVDD.n331 4.5005
R1086 DVDD.n355 DVDD.n331 4.5005
R1087 DVDD.n331 DVDD.n313 4.5005
R1088 DVDD.n331 DVDD.n312 4.5005
R1089 DVDD.n5654 DVDD.n323 4.5005
R1090 DVDD.n355 DVDD.n323 4.5005
R1091 DVDD.n323 DVDD.n313 4.5005
R1092 DVDD.n323 DVDD.n312 4.5005
R1093 DVDD.n5654 DVDD.n333 4.5005
R1094 DVDD.n355 DVDD.n333 4.5005
R1095 DVDD.n333 DVDD.n312 4.5005
R1096 DVDD.n322 DVDD.n312 4.5005
R1097 DVDD.n5654 DVDD.n322 4.5005
R1098 DVDD.n335 DVDD.n313 4.5005
R1099 DVDD.n5654 DVDD.n335 4.5005
R1100 DVDD.n321 DVDD.n313 4.5005
R1101 DVDD.n5654 DVDD.n321 4.5005
R1102 DVDD.n337 DVDD.n313 4.5005
R1103 DVDD.n5654 DVDD.n337 4.5005
R1104 DVDD.n320 DVDD.n313 4.5005
R1105 DVDD.n5654 DVDD.n320 4.5005
R1106 DVDD.n339 DVDD.n313 4.5005
R1107 DVDD.n5654 DVDD.n339 4.5005
R1108 DVDD.n319 DVDD.n313 4.5005
R1109 DVDD.n5654 DVDD.n319 4.5005
R1110 DVDD.n341 DVDD.n313 4.5005
R1111 DVDD.n5654 DVDD.n341 4.5005
R1112 DVDD.n318 DVDD.n313 4.5005
R1113 DVDD.n5654 DVDD.n318 4.5005
R1114 DVDD.n342 DVDD.n312 4.5005
R1115 DVDD.n342 DVDD.n313 4.5005
R1116 DVDD.n5654 DVDD.n342 4.5005
R1117 DVDD.n317 DVDD.n312 4.5005
R1118 DVDD.n317 DVDD.n313 4.5005
R1119 DVDD.n5654 DVDD.n317 4.5005
R1120 DVDD.n344 DVDD.n313 4.5005
R1121 DVDD.n5654 DVDD.n344 4.5005
R1122 DVDD.n316 DVDD.n313 4.5005
R1123 DVDD.n5654 DVDD.n316 4.5005
R1124 DVDD.n345 DVDD.n312 4.5005
R1125 DVDD.n345 DVDD.n313 4.5005
R1126 DVDD.n5654 DVDD.n345 4.5005
R1127 DVDD.n315 DVDD.n312 4.5005
R1128 DVDD.n315 DVDD.n313 4.5005
R1129 DVDD.n5654 DVDD.n315 4.5005
R1130 DVDD.n5653 DVDD.n312 4.5005
R1131 DVDD.n5653 DVDD.n313 4.5005
R1132 DVDD.n5654 DVDD.n5653 4.5005
R1133 DVDD.n1548 DVDD.n357 4.5005
R1134 DVDD.n2152 DVDD.n357 4.5005
R1135 DVDD.n2154 DVDD.n357 4.5005
R1136 DVDD.n2152 DVDD.n1482 4.5005
R1137 DVDD.n2154 DVDD.n1482 4.5005
R1138 DVDD.n2152 DVDD.n1480 4.5005
R1139 DVDD.n2154 DVDD.n1480 4.5005
R1140 DVDD.n1548 DVDD.n1495 4.5005
R1141 DVDD.n2152 DVDD.n1495 4.5005
R1142 DVDD.n2154 DVDD.n1495 4.5005
R1143 DVDD.n1548 DVDD.n1479 4.5005
R1144 DVDD.n2152 DVDD.n1479 4.5005
R1145 DVDD.n2154 DVDD.n1479 4.5005
R1146 DVDD.n2152 DVDD.n1496 4.5005
R1147 DVDD.n2154 DVDD.n1496 4.5005
R1148 DVDD.n2152 DVDD.n1478 4.5005
R1149 DVDD.n2154 DVDD.n1478 4.5005
R1150 DVDD.n1548 DVDD.n1509 4.5005
R1151 DVDD.n2152 DVDD.n1509 4.5005
R1152 DVDD.n2154 DVDD.n1509 4.5005
R1153 DVDD.n1548 DVDD.n1477 4.5005
R1154 DVDD.n2152 DVDD.n1477 4.5005
R1155 DVDD.n2154 DVDD.n1477 4.5005
R1156 DVDD.n2152 DVDD.n1510 4.5005
R1157 DVDD.n2154 DVDD.n1510 4.5005
R1158 DVDD.n2152 DVDD.n1476 4.5005
R1159 DVDD.n2154 DVDD.n1476 4.5005
R1160 DVDD.n1548 DVDD.n1523 4.5005
R1161 DVDD.n2152 DVDD.n1523 4.5005
R1162 DVDD.n2154 DVDD.n1523 4.5005
R1163 DVDD.n1548 DVDD.n1475 4.5005
R1164 DVDD.n2152 DVDD.n1475 4.5005
R1165 DVDD.n2154 DVDD.n1475 4.5005
R1166 DVDD.n2152 DVDD.n1524 4.5005
R1167 DVDD.n2154 DVDD.n1524 4.5005
R1168 DVDD.n2152 DVDD.n1474 4.5005
R1169 DVDD.n2154 DVDD.n1474 4.5005
R1170 DVDD.n1548 DVDD.n1537 4.5005
R1171 DVDD.n2152 DVDD.n1537 4.5005
R1172 DVDD.n2154 DVDD.n1537 4.5005
R1173 DVDD.n1548 DVDD.n1473 4.5005
R1174 DVDD.n2152 DVDD.n1473 4.5005
R1175 DVDD.n2154 DVDD.n1473 4.5005
R1176 DVDD.n2152 DVDD.n1538 4.5005
R1177 DVDD.n2154 DVDD.n1538 4.5005
R1178 DVDD.n2152 DVDD.n1472 4.5005
R1179 DVDD.n2154 DVDD.n1472 4.5005
R1180 DVDD.n1548 DVDD.n1539 4.5005
R1181 DVDD.n2152 DVDD.n1539 4.5005
R1182 DVDD.n2154 DVDD.n1539 4.5005
R1183 DVDD.n1548 DVDD.n1471 4.5005
R1184 DVDD.n2152 DVDD.n1471 4.5005
R1185 DVDD.n2154 DVDD.n1471 4.5005
R1186 DVDD.n2152 DVDD.n1540 4.5005
R1187 DVDD.n2154 DVDD.n1540 4.5005
R1188 DVDD.n2152 DVDD.n1470 4.5005
R1189 DVDD.n2154 DVDD.n1470 4.5005
R1190 DVDD.n2153 DVDD.n1548 4.5005
R1191 DVDD.n2153 DVDD.n2152 4.5005
R1192 DVDD.n2154 DVDD.n2153 4.5005
R1193 DVDD.n2369 DVDD.n1221 4.5005
R1194 DVDD.n2371 DVDD.n1221 4.5005
R1195 DVDD.n1221 DVDD.n1189 4.5005
R1196 DVDD.n2369 DVDD.n1235 4.5005
R1197 DVDD.n2371 DVDD.n1235 4.5005
R1198 DVDD.n1235 DVDD.n1189 4.5005
R1199 DVDD.n2369 DVDD.n1220 4.5005
R1200 DVDD.n2371 DVDD.n1220 4.5005
R1201 DVDD.n1220 DVDD.n1189 4.5005
R1202 DVDD.n2371 DVDD.n1236 4.5005
R1203 DVDD.n1236 DVDD.n1189 4.5005
R1204 DVDD.n2371 DVDD.n1219 4.5005
R1205 DVDD.n1219 DVDD.n1189 4.5005
R1206 DVDD.n2371 DVDD.n1237 4.5005
R1207 DVDD.n1237 DVDD.n1189 4.5005
R1208 DVDD.n2371 DVDD.n1218 4.5005
R1209 DVDD.n1218 DVDD.n1189 4.5005
R1210 DVDD.n2371 DVDD.n1238 4.5005
R1211 DVDD.n1238 DVDD.n1189 4.5005
R1212 DVDD.n2371 DVDD.n1217 4.5005
R1213 DVDD.n1217 DVDD.n1189 4.5005
R1214 DVDD.n2371 DVDD.n1239 4.5005
R1215 DVDD.n1239 DVDD.n1189 4.5005
R1216 DVDD.n2371 DVDD.n1216 4.5005
R1217 DVDD.n1216 DVDD.n1189 4.5005
R1218 DVDD.n2371 DVDD.n1240 4.5005
R1219 DVDD.n1240 DVDD.n1189 4.5005
R1220 DVDD.n2371 DVDD.n1215 4.5005
R1221 DVDD.n1215 DVDD.n1189 4.5005
R1222 DVDD.n2369 DVDD.n1253 4.5005
R1223 DVDD.n2371 DVDD.n1253 4.5005
R1224 DVDD.n1253 DVDD.n1189 4.5005
R1225 DVDD.n2369 DVDD.n1214 4.5005
R1226 DVDD.n2371 DVDD.n1214 4.5005
R1227 DVDD.n1214 DVDD.n1189 4.5005
R1228 DVDD.n2371 DVDD.n1254 4.5005
R1229 DVDD.n1254 DVDD.n1189 4.5005
R1230 DVDD.n2371 DVDD.n1213 4.5005
R1231 DVDD.n1213 DVDD.n1189 4.5005
R1232 DVDD.n2369 DVDD.n1255 4.5005
R1233 DVDD.n2371 DVDD.n1255 4.5005
R1234 DVDD.n1255 DVDD.n1189 4.5005
R1235 DVDD.n2369 DVDD.n1212 4.5005
R1236 DVDD.n2371 DVDD.n1212 4.5005
R1237 DVDD.n1212 DVDD.n1189 4.5005
R1238 DVDD.n2371 DVDD.n1256 4.5005
R1239 DVDD.n1256 DVDD.n1189 4.5005
R1240 DVDD.n1265 DVDD.n1189 4.5005
R1241 DVDD.n2370 DVDD.n2369 4.5005
R1242 DVDD.n2371 DVDD.n2370 4.5005
R1243 DVDD.n2370 DVDD.n1189 4.5005
R1244 DVDD.n2371 DVDD.n1211 4.5005
R1245 DVDD.n1211 DVDD.n1189 4.5005
R1246 DVDD.n2372 DVDD.n2371 4.5005
R1247 DVDD.n2373 DVDD.n2372 4.5005
R1248 DVDD.n2372 DVDD.n1189 4.5005
R1249 DVDD.n2564 DVDD.n1042 4.5005
R1250 DVDD.n1042 DVDD.n1015 4.5005
R1251 DVDD.n1042 DVDD.n1016 4.5005
R1252 DVDD.n1040 DVDD.n1015 4.5005
R1253 DVDD.n1040 DVDD.n1016 4.5005
R1254 DVDD.n2511 DVDD.n1015 4.5005
R1255 DVDD.n2511 DVDD.n1016 4.5005
R1256 DVDD.n2564 DVDD.n2527 4.5005
R1257 DVDD.n2527 DVDD.n1015 4.5005
R1258 DVDD.n2527 DVDD.n1016 4.5005
R1259 DVDD.n2564 DVDD.n1038 4.5005
R1260 DVDD.n1038 DVDD.n1015 4.5005
R1261 DVDD.n1038 DVDD.n1016 4.5005
R1262 DVDD.n1036 DVDD.n1015 4.5005
R1263 DVDD.n1036 DVDD.n1016 4.5005
R1264 DVDD.n2529 DVDD.n1016 4.5005
R1265 DVDD.n2564 DVDD.n2542 4.5005
R1266 DVDD.n2542 DVDD.n1015 4.5005
R1267 DVDD.n2542 DVDD.n1016 4.5005
R1268 DVDD.n2546 DVDD.n1015 4.5005
R1269 DVDD.n2546 DVDD.n1016 4.5005
R1270 DVDD.n2544 DVDD.n1015 4.5005
R1271 DVDD.n2544 DVDD.n1016 4.5005
R1272 DVDD.n2564 DVDD.n1034 4.5005
R1273 DVDD.n1034 DVDD.n1015 4.5005
R1274 DVDD.n1034 DVDD.n1016 4.5005
R1275 DVDD.n2561 DVDD.n1016 4.5005
R1276 DVDD.n2561 DVDD.n1017 4.5005
R1277 DVDD.n2564 DVDD.n2561 4.5005
R1278 DVDD.n2564 DVDD.n1033 4.5005
R1279 DVDD.n1033 DVDD.n1016 4.5005
R1280 DVDD.n1031 DVDD.n1015 4.5005
R1281 DVDD.n1031 DVDD.n1016 4.5005
R1282 DVDD.n1015 DVDD.n978 4.5005
R1283 DVDD.n1017 DVDD.n978 4.5005
R1284 DVDD.n1016 DVDD.n978 4.5005
R1285 DVDD.n1016 DVDD.n979 4.5005
R1286 DVDD.n1017 DVDD.n979 4.5005
R1287 DVDD.n2564 DVDD.n979 4.5005
R1288 DVDD.n2564 DVDD.n1029 4.5005
R1289 DVDD.n1029 DVDD.n1016 4.5005
R1290 DVDD.n1027 DVDD.n1015 4.5005
R1291 DVDD.n1027 DVDD.n1016 4.5005
R1292 DVDD.n1024 DVDD.n1015 4.5005
R1293 DVDD.n1024 DVDD.n1017 4.5005
R1294 DVDD.n1024 DVDD.n1016 4.5005
R1295 DVDD.n2563 DVDD.n1016 4.5005
R1296 DVDD.n2563 DVDD.n1017 4.5005
R1297 DVDD.n2564 DVDD.n2563 4.5005
R1298 DVDD.n2564 DVDD.n1023 4.5005
R1299 DVDD.n1023 DVDD.n1016 4.5005
R1300 DVDD.n1021 DVDD.n1015 4.5005
R1301 DVDD.n1021 DVDD.n1016 4.5005
R1302 DVDD.n1019 DVDD.n1015 4.5005
R1303 DVDD.n1019 DVDD.n1017 4.5005
R1304 DVDD.n1019 DVDD.n1016 4.5005
R1305 DVDD.n2565 DVDD.n1016 4.5005
R1306 DVDD.n2565 DVDD.n1017 4.5005
R1307 DVDD.n2565 DVDD.n1015 4.5005
R1308 DVDD.n2565 DVDD.n2564 4.5005
R1309 DVDD.n518 DVDD.n506 4.5005
R1310 DVDD.n2601 DVDD.n518 4.5005
R1311 DVDD.n5568 DVDD.n518 4.5005
R1312 DVDD.n5568 DVDD.n515 4.5005
R1313 DVDD.n515 DVDD.n506 4.5005
R1314 DVDD.n2597 DVDD.n510 4.5005
R1315 DVDD.n2597 DVDD.n506 4.5005
R1316 DVDD.n2603 DVDD.n506 4.5005
R1317 DVDD.n520 DVDD.n506 4.5005
R1318 DVDD.n2601 DVDD.n520 4.5005
R1319 DVDD.n5568 DVDD.n520 4.5005
R1320 DVDD.n5568 DVDD.n513 4.5005
R1321 DVDD.n513 DVDD.n506 4.5005
R1322 DVDD.n2599 DVDD.n510 4.5005
R1323 DVDD.n2599 DVDD.n506 4.5005
R1324 DVDD.n2596 DVDD.n510 4.5005
R1325 DVDD.n2601 DVDD.n2596 4.5005
R1326 DVDD.n2596 DVDD.n506 4.5005
R1327 DVDD.n522 DVDD.n506 4.5005
R1328 DVDD.n2601 DVDD.n522 4.5005
R1329 DVDD.n5568 DVDD.n522 4.5005
R1330 DVDD.n5568 DVDD.n511 4.5005
R1331 DVDD.n511 DVDD.n506 4.5005
R1332 DVDD.n5568 DVDD.n5567 4.5005
R1333 DVDD.n5567 DVDD.n510 4.5005
R1334 DVDD.n5567 DVDD.n506 4.5005
R1335 DVDD.n4640 DVDD.n3397 4.5005
R1336 DVDD.n4641 DVDD.n4640 4.5005
R1337 DVDD.n4640 DVDD.n3400 4.5005
R1338 DVDD.n4640 DVDD.n4639 4.5005
R1339 DVDD.n3259 DVDD.n178 4.5005
R1340 DVDD.n3303 DVDD.n178 4.5005
R1341 DVDD.n3306 DVDD.n178 4.5005
R1342 DVDD.n3257 DVDD.n178 4.5005
R1343 DVDD.n3311 DVDD.n178 4.5005
R1344 DVDD.n3517 DVDD.n3510 4.5005
R1345 DVDD.n4204 DVDD.n4203 4.5005
R1346 DVDD.n3915 DVDD.n3667 4.5005
R1347 DVDD.n3918 DVDD.n3666 4.5005
R1348 DVDD.n4684 DVDD.n3376 4.5005
R1349 DVDD.n3956 DVDD.n3655 4.5005
R1350 DVDD.n3655 DVDD.n3644 4.5005
R1351 DVDD.n3956 DVDD.n3653 4.5005
R1352 DVDD.n3653 DVDD.n3644 4.5005
R1353 DVDD.n3955 DVDD.n3644 4.5005
R1354 DVDD.n3649 DVDD.n3644 4.5005
R1355 DVDD.n3659 DVDD.n3644 4.5005
R1356 DVDD.n3650 DVDD.n3644 4.5005
R1357 DVDD.n3956 DVDD.n3656 4.5005
R1358 DVDD.n3656 DVDD.n3644 4.5005
R1359 DVDD.n3956 DVDD.n3652 4.5005
R1360 DVDD.n3652 DVDD.n3644 4.5005
R1361 DVDD.n3956 DVDD.n3657 4.5005
R1362 DVDD.n3657 DVDD.n3644 4.5005
R1363 DVDD.n3658 DVDD.n3644 4.5005
R1364 DVDD.n3651 DVDD.n3644 4.5005
R1365 DVDD.n3956 DVDD.n3651 4.5005
R1366 DVDD.n3956 DVDD.n3658 4.5005
R1367 DVDD.n3956 DVDD.n3650 4.5005
R1368 DVDD.n3956 DVDD.n3659 4.5005
R1369 DVDD.n3956 DVDD.n3649 4.5005
R1370 DVDD.n3956 DVDD.n3955 4.5005
R1371 DVDD.n3041 DVDD.n3040 4.5005
R1372 DVDD.n3040 DVDD.n261 4.5005
R1373 DVDD.n5704 DVDD.n5703 4.5005
R1374 DVDD.n1721 DVDD.n273 4.5005
R1375 DVDD.n2037 DVDD.n1722 4.5005
R1376 DVDD.n2034 DVDD.n564 4.5005
R1377 DVDD.n2037 DVDD.n565 4.5005
R1378 DVDD.n2034 DVDD.n565 4.5005
R1379 DVDD.n2037 DVDD.n1720 4.5005
R1380 DVDD.n2034 DVDD.n1720 4.5005
R1381 DVDD.n2034 DVDD.n2028 4.5005
R1382 DVDD.n2037 DVDD.n1742 4.5005
R1383 DVDD.n2037 DVDD.n1718 4.5005
R1384 DVDD.n2037 DVDD.n1715 4.5005
R1385 DVDD.n2038 DVDD.n2037 4.5005
R1386 DVDD.n2037 DVDD.n899 4.5005
R1387 DVDD.n2964 DVDD.n2963 4.5005
R1388 DVDD.n2963 DVDD.n909 4.5005
R1389 DVDD.n2963 DVDD.n906 4.5005
R1390 DVDD.n2963 DVDD.n911 4.5005
R1391 DVDD.n2963 DVDD.n905 4.5005
R1392 DVDD.n2963 DVDD.n913 4.5005
R1393 DVDD.n2963 DVDD.n904 4.5005
R1394 DVDD.n2963 DVDD.n915 4.5005
R1395 DVDD.n2963 DVDD.n903 4.5005
R1396 DVDD.n2963 DVDD.n917 4.5005
R1397 DVDD.n2963 DVDD.n902 4.5005
R1398 DVDD.n2963 DVDD.n2962 4.5005
R1399 DVDD.n2960 DVDD.n2959 4.5005
R1400 DVDD.n2959 DVDD.n928 4.5005
R1401 DVDD.n2959 DVDD.n926 4.5005
R1402 DVDD.n2959 DVDD.n934 4.5005
R1403 DVDD.n2959 DVDD.n925 4.5005
R1404 DVDD.n2959 DVDD.n936 4.5005
R1405 DVDD.n2959 DVDD.n924 4.5005
R1406 DVDD.n2956 DVDD.n939 4.5005
R1407 DVDD.n2959 DVDD.n2958 4.5005
R1408 DVDD.n2956 DVDD.n2955 4.5005
R1409 DVDD.n2953 DVDD.n2952 4.5005
R1410 DVDD.n2952 DVDD.n961 4.5005
R1411 DVDD.n2952 DVDD.n958 4.5005
R1412 DVDD.n2949 DVDD.n971 4.5005
R1413 DVDD.n2952 DVDD.n963 4.5005
R1414 DVDD.n2952 DVDD.n956 4.5005
R1415 DVDD.n2949 DVDD.n975 4.5005
R1416 DVDD.n2949 DVDD.n968 4.5005
R1417 DVDD.n2949 DVDD.n2946 4.5005
R1418 DVDD.n2949 DVDD.n967 4.5005
R1419 DVDD.n2949 DVDD.n2948 4.5005
R1420 DVDD.n2949 DVDD.n966 4.5005
R1421 DVDD.n2952 DVDD.n475 4.5005
R1422 DVDD.n2949 DVDD.n475 4.5005
R1423 DVDD.n5616 DVDD.n5615 4.5005
R1424 DVDD.n5615 DVDD.n480 4.5005
R1425 DVDD.n5615 DVDD.n483 4.5005
R1426 DVDD.n5615 DVDD.n479 4.5005
R1427 DVDD.n5615 DVDD.n485 4.5005
R1428 DVDD.n5612 DVDD.n486 4.5005
R1429 DVDD.n4684 DVDD.n4683 4.5005
R1430 DVDD.n4740 DVDD.n3355 4.5005
R1431 DVDD.n4741 DVDD.n4740 4.5005
R1432 DVDD.n5506 DVDD.n5505 4.5005
R1433 DVDD.n5511 DVDD.n562 4.5005
R1434 DVDD.n5509 DVDD.n562 4.5005
R1435 DVDD.n5508 DVDD.n566 4.5005
R1436 DVDD.n5503 DVDD.n573 4.5005
R1437 DVDD.n5501 DVDD.n573 4.5005
R1438 DVDD.n5500 DVDD.n577 4.5005
R1439 DVDD.n577 DVDD.n544 4.5005
R1440 DVDD.n5511 DVDD.n5510 4.5005
R1441 DVDD.n5510 DVDD.n5509 4.5005
R1442 DVDD.n5508 DVDD.n5507 4.5005
R1443 DVDD.n5507 DVDD.n569 4.5005
R1444 DVDD.n5507 DVDD.n571 4.5005
R1445 DVDD.n5507 DVDD.n568 4.5005
R1446 DVDD.n5507 DVDD.n5506 4.5005
R1447 DVDD.n5503 DVDD.n5502 4.5005
R1448 DVDD.n5502 DVDD.n5501 4.5005
R1449 DVDD.n5500 DVDD.n5499 4.5005
R1450 DVDD.n5499 DVDD.n544 4.5005
R1451 DVDD.n5526 DVDD.n549 4.5005
R1452 DVDD.n549 DVDD.n543 4.5005
R1453 DVDD.n5525 DVDD.n5524 4.5005
R1454 DVDD.n5526 DVDD.n5525 4.5005
R1455 DVDD.n5525 DVDD.n543 4.5005
R1456 DVDD.n5524 DVDD.n5523 4.5005
R1457 DVDD.n5523 DVDD.n543 4.5005
R1458 DVDD.n5514 DVDD.n558 4.5005
R1459 DVDD.n5512 DVDD.n558 4.5005
R1460 DVDD.n5514 DVDD.n5513 4.5005
R1461 DVDD.n5513 DVDD.n5512 4.5005
R1462 DVDD.n4207 DVDD.n4206 4.5005
R1463 DVDD.n3800 DVDD.n3509 4.5005
R1464 DVDD.n3802 DVDD.n3801 4.5005
R1465 DVDD.n3803 DVDD.n3799 4.5005
R1466 DVDD.n3805 DVDD.n3804 4.5005
R1467 DVDD.n3806 DVDD.n3798 4.5005
R1468 DVDD.n3808 DVDD.n3807 4.5005
R1469 DVDD.n3809 DVDD.n3797 4.5005
R1470 DVDD.n3811 DVDD.n3810 4.5005
R1471 DVDD.n3812 DVDD.n3796 4.5005
R1472 DVDD.n3814 DVDD.n3813 4.5005
R1473 DVDD.n3815 DVDD.n3795 4.5005
R1474 DVDD.n3817 DVDD.n3816 4.5005
R1475 DVDD.n3818 DVDD.n3794 4.5005
R1476 DVDD.n3820 DVDD.n3819 4.5005
R1477 DVDD.n3821 DVDD.n3793 4.5005
R1478 DVDD.n3823 DVDD.n3822 4.5005
R1479 DVDD.n3824 DVDD.n3792 4.5005
R1480 DVDD.n3826 DVDD.n3825 4.5005
R1481 DVDD.n3827 DVDD.n3687 4.5005
R1482 DVDD.n3829 DVDD.n3828 4.5005
R1483 DVDD.n3791 DVDD.n3686 4.5005
R1484 DVDD.n3790 DVDD.n3789 4.5005
R1485 DVDD.n3788 DVDD.n3688 4.5005
R1486 DVDD.n3787 DVDD.n3786 4.5005
R1487 DVDD.n3785 DVDD.n3689 4.5005
R1488 DVDD.n3784 DVDD.n3783 4.5005
R1489 DVDD.n3782 DVDD.n3690 4.5005
R1490 DVDD.n3781 DVDD.n3780 4.5005
R1491 DVDD.n3779 DVDD.n3691 4.5005
R1492 DVDD.n3778 DVDD.n3777 4.5005
R1493 DVDD.n3776 DVDD.n3692 4.5005
R1494 DVDD.n3775 DVDD.n3774 4.5005
R1495 DVDD.n3773 DVDD.n3693 4.5005
R1496 DVDD.n3772 DVDD.n3771 4.5005
R1497 DVDD.n3770 DVDD.n3694 4.5005
R1498 DVDD.n3769 DVDD.n3768 4.5005
R1499 DVDD.n3767 DVDD.n3695 4.5005
R1500 DVDD.n3766 DVDD.n3765 4.5005
R1501 DVDD.n3764 DVDD.n3696 4.5005
R1502 DVDD.n3763 DVDD.n3762 4.5005
R1503 DVDD.n3745 DVDD.n3698 4.5005
R1504 DVDD.n3756 DVDD.n3699 4.5005
R1505 DVDD.n5714 DVDD.n5713 4.5005
R1506 DVDD.n5713 DVDD.n5712 4.5005
R1507 DVDD.n2974 DVDD.n256 4.5005
R1508 DVDD.n2972 DVDD.n2971 4.5005
R1509 DVDD.n2970 DVDD.n2969 4.5005
R1510 DVDD.n1798 DVDD.n560 4.5005
R1511 DVDD.n2969 DVDD.n561 4.5005
R1512 DVDD.n1798 DVDD.n561 4.5005
R1513 DVDD.n2969 DVDD.n886 4.5005
R1514 DVDD.n1798 DVDD.n886 4.5005
R1515 DVDD.n1798 DVDD.n1790 4.5005
R1516 DVDD.n2969 DVDD.n894 4.5005
R1517 DVDD.n2969 DVDD.n884 4.5005
R1518 DVDD.n2969 DVDD.n896 4.5005
R1519 DVDD.n2969 DVDD.n883 4.5005
R1520 DVDD.n2969 DVDD.n2968 4.5005
R1521 DVDD.n2220 DVDD.n898 4.5005
R1522 DVDD.n2220 DVDD.n1400 4.5005
R1523 DVDD.n2220 DVDD.n1397 4.5005
R1524 DVDD.n2220 DVDD.n1402 4.5005
R1525 DVDD.n2220 DVDD.n1396 4.5005
R1526 DVDD.n2220 DVDD.n1404 4.5005
R1527 DVDD.n2220 DVDD.n1395 4.5005
R1528 DVDD.n2220 DVDD.n1406 4.5005
R1529 DVDD.n2220 DVDD.n1394 4.5005
R1530 DVDD.n2220 DVDD.n1391 4.5005
R1531 DVDD.n2221 DVDD.n2220 4.5005
R1532 DVDD.n2220 DVDD.n2219 4.5005
R1533 DVDD.n2441 DVDD.n1127 4.5005
R1534 DVDD.n2441 DVDD.n1129 4.5005
R1535 DVDD.n2441 DVDD.n1126 4.5005
R1536 DVDD.n2441 DVDD.n1135 4.5005
R1537 DVDD.n2441 DVDD.n1125 4.5005
R1538 DVDD.n2441 DVDD.n1121 4.5005
R1539 DVDD.n2442 DVDD.n2441 4.5005
R1540 DVDD.n2438 DVDD.n1139 4.5005
R1541 DVDD.n2441 DVDD.n2440 4.5005
R1542 DVDD.n2438 DVDD.n2437 4.5005
R1543 DVDD.n2435 DVDD.n472 4.5005
R1544 DVDD.n2514 DVDD.n472 4.5005
R1545 DVDD.n2515 DVDD.n472 4.5005
R1546 DVDD.n5622 DVDD.n453 4.5005
R1547 DVDD.n2531 DVDD.n472 4.5005
R1548 DVDD.n2549 DVDD.n472 4.5005
R1549 DVDD.n5622 DVDD.n458 4.5005
R1550 DVDD.n5622 DVDD.n450 4.5005
R1551 DVDD.n5622 DVDD.n460 4.5005
R1552 DVDD.n5622 DVDD.n446 4.5005
R1553 DVDD.n5623 DVDD.n5622 4.5005
R1554 DVDD.n5622 DVDD.n449 4.5005
R1555 DVDD.n5621 DVDD.n472 4.5005
R1556 DVDD.n5622 DVDD.n5621 4.5005
R1557 DVDD.n2914 DVDD.n2592 4.5005
R1558 DVDD.n2914 DVDD.n2590 4.5005
R1559 DVDD.n2914 DVDD.n2764 4.5005
R1560 DVDD.n2914 DVDD.n2587 4.5005
R1561 DVDD.n2915 DVDD.n2914 4.5005
R1562 DVDD.n2912 DVDD.n2911 4.5005
R1563 DVDD.n4320 DVDD.n4216 4.5005
R1564 DVDD.n4847 DVDD.n4786 4.5005
R1565 DVDD.n4847 DVDD.n4846 4.5005
R1566 DVDD.n4320 DVDD.n4319 4.5005
R1567 DVDD.n4322 DVDD.n4215 4.5005
R1568 DVDD.n4325 DVDD.n4208 4.5005
R1569 DVDD.n4325 DVDD.n3505 4.5005
R1570 DVDD.n4322 DVDD.n3505 4.5005
R1571 DVDD.n4325 DVDD.n3504 4.5005
R1572 DVDD.n4322 DVDD.n4321 4.5005
R1573 DVDD.n3375 DVDD.n3373 4.5005
R1574 DVDD.n3516 DVDD.n3373 4.5005
R1575 DVDD.n4690 DVDD.n3373 4.5005
R1576 DVDD.n4685 DVDD.n3374 4.5005
R1577 DVDD.n4493 DVDD.n3399 4.5005
R1578 DVDD.n3445 DVDD.n3399 4.5005
R1579 DVDD.n4488 DVDD.n3399 4.5005
R1580 DVDD.n3447 DVDD.n3445 4.5005
R1581 DVDD.n4488 DVDD.n3447 4.5005
R1582 DVDD.n4486 DVDD.n3445 4.5005
R1583 DVDD.n4488 DVDD.n4486 4.5005
R1584 DVDD.n3446 DVDD.n3445 4.5005
R1585 DVDD.n4488 DVDD.n3446 4.5005
R1586 DVDD.n4489 DVDD.n3445 4.5005
R1587 DVDD.n4489 DVDD.n4488 4.5005
R1588 DVDD.n4493 DVDD.n3435 4.5005
R1589 DVDD.n3445 DVDD.n3435 4.5005
R1590 DVDD.n4488 DVDD.n3435 4.5005
R1591 DVDD.n4491 DVDD.n3401 4.5005
R1592 DVDD.n4488 DVDD.n3401 4.5005
R1593 DVDD.n4491 DVDD.n3439 4.5005
R1594 DVDD.n4493 DVDD.n3439 4.5005
R1595 DVDD.n4491 DVDD.n3434 4.5005
R1596 DVDD.n4493 DVDD.n3434 4.5005
R1597 DVDD.n4492 DVDD.n4491 4.5005
R1598 DVDD.n4493 DVDD.n4492 4.5005
R1599 DVDD.n4494 DVDD.n4493 4.5005
R1600 DVDD.n4493 DVDD.n3401 4.5005
R1601 DVDD.n3427 DVDD.n3425 4.5005
R1602 DVDD.n4192 DVDD.n3427 4.5005
R1603 DVDD.n4538 DVDD.n3427 4.5005
R1604 DVDD.n4543 DVDD.n3426 4.5005
R1605 DVDD.n26 DVDD.n11 4.5005
R1606 DVDD.n5987 DVDD.n22 4.5005
R1607 DVDD.n16 DVDD.n11 4.5005
R1608 DVDD.n5987 DVDD.n16 4.5005
R1609 DVDD.n3184 DVDD.n11 4.5005
R1610 DVDD.n5987 DVDD.n5986 4.5005
R1611 DVDD.n70 DVDD.t6 4.06554
R1612 DVDD.n5908 DVDD.t9 4.06554
R1613 DVDD.n5924 DVDD.t6 3.48482
R1614 DVDD.n84 DVDD.t9 3.48482
R1615 DVDD.n5516 DVDD.n5515 3.3314
R1616 DVDD.n5545 DVDD.n5529 3.33081
R1617 DVDD.n5515 DVDD.n5514 3.31632
R1618 DVDD.n5529 DVDD.n544 3.31632
R1619 DVDD.n5482 DVDD.n5481 3.10905
R1620 DVDD.n5711 DVDD.n5710 3.10905
R1621 DVDD.n5367 DVDD.n5366 3.0398
R1622 DVDD.n5142 DVDD.n5141 3.0398
R1623 DVDD.n3042 DVDD.n3041 3.0398
R1624 DVDD.n5715 DVDD.n5714 3.0398
R1625 DVDD.n5940 DVDD.t70 2.9041
R1626 DVDD.n98 DVDD.t27 2.9041
R1627 DVDD.n1736 DVDD.n1735 2.87501
R1628 DVDD.n2045 DVDD.n2044 2.87501
R1629 DVDD.n5651 DVDD.n5649 2.87501
R1630 DVDD.n1493 DVDD.n1491 2.87501
R1631 DVDD.n1507 DVDD.n1505 2.87501
R1632 DVDD.n1521 DVDD.n1519 2.87501
R1633 DVDD.n1535 DVDD.n1533 2.87501
R1634 DVDD.n2227 DVDD.n2226 2.87501
R1635 DVDD.n1551 DVDD.n381 2.87501
R1636 DVDD.n1233 DVDD.n1231 2.87501
R1637 DVDD.n1251 DVDD.n1249 2.87501
R1638 DVDD.n2448 DVDD.n2447 2.87501
R1639 DVDD.n1263 DVDD.n1261 2.87501
R1640 DVDD.n1209 DVDD.n411 2.87501
R1641 DVDD.n2525 DVDD.n2523 2.87501
R1642 DVDD.n2540 DVDD.n2538 2.87501
R1643 DVDD.n2558 DVDD.n2556 2.87501
R1644 DVDD.n2940 DVDD.n2939 2.87501
R1645 DVDD.n5629 DVDD.n5628 2.87501
R1646 DVDD.n1013 DVDD.n1011 2.87501
R1647 DVDD.n2567 DVDD.n1007 2.87501
R1648 DVDD.n2573 DVDD.n2572 2.87501
R1649 DVDD.n2758 DVDD.n2757 2.87501
R1650 DVDD.n2921 DVDD.n2920 2.87501
R1651 DVDD.n5565 DVDD.n5563 2.87501
R1652 DVDD.n2768 DVDD.n528 2.87501
R1653 DVDD.n2785 DVDD.n529 2.87501
R1654 DVDD.n2789 DVDD.n530 2.87501
R1655 DVDD.n2793 DVDD.n531 2.87501
R1656 DVDD.n2797 DVDD.n532 2.87501
R1657 DVDD.n2801 DVDD.n533 2.87501
R1658 DVDD.n2805 DVDD.n534 2.87501
R1659 DVDD.n2809 DVDD.n535 2.87501
R1660 DVDD.n2813 DVDD.n536 2.87501
R1661 DVDD.n2817 DVDD.n537 2.87501
R1662 DVDD.n2821 DVDD.n538 2.87501
R1663 DVDD.n2825 DVDD.n539 2.87501
R1664 DVDD.n2827 DVDD.n540 2.87501
R1665 DVDD.n2844 DVDD.n541 2.87501
R1666 DVDD.n5521 DVDD.n542 2.87501
R1667 DVDD.n1740 DVDD.n1738 2.81339
R1668 DVDD.n2042 DVDD.n2041 2.81339
R1669 DVDD.n2966 DVDD.n358 2.81339
R1670 DVDD.n1486 DVDD.n1485 2.81339
R1671 DVDD.n1500 DVDD.n1499 2.81339
R1672 DVDD.n1514 DVDD.n1513 2.81339
R1673 DVDD.n1528 DVDD.n1527 2.81339
R1674 DVDD.n2224 DVDD.n2223 2.81339
R1675 DVDD.n1549 DVDD.n920 2.81339
R1676 DVDD.n1226 DVDD.n1225 2.81339
R1677 DVDD.n1244 DVDD.n1243 2.81339
R1678 DVDD.n2445 DVDD.n2444 2.81339
R1679 DVDD.n1258 DVDD.n1257 2.81339
R1680 DVDD.n1207 DVDD.n950 2.81339
R1681 DVDD.n2518 DVDD.n2517 2.81339
R1682 DVDD.n2534 DVDD.n2533 2.81339
R1683 DVDD.n2552 DVDD.n2551 2.81339
R1684 DVDD.n2944 DVDD.n2942 2.81339
R1685 DVDD.n5626 DVDD.n5625 2.81339
R1686 DVDD.n1010 DVDD.n1009 2.81339
R1687 DVDD.n5619 DVDD.n474 2.81339
R1688 DVDD.n2570 DVDD.n476 2.81339
R1689 DVDD.n2762 DVDD.n2760 2.81339
R1690 DVDD.n2918 DVDD.n2917 2.81339
R1691 DVDD.n2862 DVDD.n525 2.81339
R1692 DVDD.n2770 DVDD.n2769 2.81339
R1693 DVDD.n2783 DVDD.n2771 2.81339
R1694 DVDD.n2787 DVDD.n2772 2.81339
R1695 DVDD.n2791 DVDD.n2773 2.81339
R1696 DVDD.n2795 DVDD.n2774 2.81339
R1697 DVDD.n2799 DVDD.n2775 2.81339
R1698 DVDD.n2803 DVDD.n2776 2.81339
R1699 DVDD.n2807 DVDD.n2777 2.81339
R1700 DVDD.n2811 DVDD.n2778 2.81339
R1701 DVDD.n2815 DVDD.n2779 2.81339
R1702 DVDD.n2819 DVDD.n2780 2.81339
R1703 DVDD.n2823 DVDD.n2781 2.81339
R1704 DVDD.n2842 DVDD.n2829 2.81339
R1705 DVDD.n2846 DVDD.n2845 2.81339
R1706 DVDD.n5519 DVDD.n5518 2.81339
R1707 DVDD.n4118 DVDD.n4116 2.66722
R1708 DVDD.n3757 DVDD.n3756 2.66722
R1709 DVDD.n5876 DVDD.n5832 2.33866
R1710 DVDD.n5942 DVDD.t4 2.32338
R1711 DVDD.n5885 DVDD.t7 2.32338
R1712 DVDD.n4230 DVDD.n4229 2.30804
R1713 DVDD.n4231 DVDD.n4224 2.30804
R1714 DVDD.n4238 DVDD.n4237 2.30804
R1715 DVDD.n4239 DVDD.n4222 2.30804
R1716 DVDD.n4246 DVDD.n4245 2.30804
R1717 DVDD.n4247 DVDD.n4220 2.30804
R1718 DVDD.n4254 DVDD.n4253 2.30804
R1719 DVDD.n4258 DVDD.n4218 2.30804
R1720 DVDD.n4317 DVDD.n4260 2.30804
R1721 DVDD.n4315 DVDD.n4314 2.30804
R1722 DVDD.n4310 DVDD.n4264 2.30804
R1723 DVDD.n4308 DVDD.n4307 2.30804
R1724 DVDD.n4303 DVDD.n4267 2.30804
R1725 DVDD.n4301 DVDD.n4300 2.30804
R1726 DVDD.n4296 DVDD.n4270 2.30804
R1727 DVDD.n4294 DVDD.n4293 2.30804
R1728 DVDD.n4289 DVDD.n4273 2.30804
R1729 DVDD.n4287 DVDD.n4286 2.30804
R1730 DVDD.n4282 DVDD.n4276 2.30804
R1731 DVDD.n4280 DVDD.n4279 2.30804
R1732 DVDD.n4681 DVDD.n3379 2.30804
R1733 DVDD.n4679 DVDD.n4678 2.30804
R1734 DVDD.n4674 DVDD.n3382 2.30804
R1735 DVDD.n4672 DVDD.n4671 2.30804
R1736 DVDD.n4667 DVDD.n3385 2.30804
R1737 DVDD.n4665 DVDD.n4664 2.30804
R1738 DVDD.n4660 DVDD.n3388 2.30804
R1739 DVDD.n4658 DVDD.n4657 2.30804
R1740 DVDD.n4653 DVDD.n3391 2.30804
R1741 DVDD.n4651 DVDD.n4650 2.30804
R1742 DVDD.n4646 DVDD.n3394 2.30804
R1743 DVDD.n4644 DVDD.n4643 2.30804
R1744 DVDD.n3405 DVDD.n3404 2.30804
R1745 DVDD.n4637 DVDD.n3407 2.30804
R1746 DVDD.n4635 DVDD.n4634 2.30804
R1747 DVDD.n4630 DVDD.n3410 2.30804
R1748 DVDD.n4628 DVDD.n4627 2.30804
R1749 DVDD.n4623 DVDD.n3413 2.30804
R1750 DVDD.n4621 DVDD.n4620 2.30804
R1751 DVDD.n4616 DVDD.n3416 2.30804
R1752 DVDD.n4614 DVDD.n4613 2.30804
R1753 DVDD.n4609 DVDD.n3419 2.30804
R1754 DVDD.n4607 DVDD.n4606 2.30804
R1755 DVDD.n4602 DVDD.n3422 2.30804
R1756 DVDD.n4600 DVDD.n4599 2.30804
R1757 DVDD.n4595 DVDD.n4547 2.30804
R1758 DVDD.n4593 DVDD.n4592 2.30804
R1759 DVDD.n4588 DVDD.n4550 2.30804
R1760 DVDD.n4586 DVDD.n4585 2.30804
R1761 DVDD.n4581 DVDD.n4553 2.30804
R1762 DVDD.n4579 DVDD.n4578 2.30804
R1763 DVDD.n4574 DVDD.n4556 2.30804
R1764 DVDD.n4572 DVDD.n4571 2.30804
R1765 DVDD.n4567 DVDD.n4559 2.30804
R1766 DVDD.n4565 DVDD.n4564 2.30804
R1767 DVDD.n4560 DVDD.n30 2.30804
R1768 DVDD.n5980 DVDD.n5979 2.30804
R1769 DVDD.n5977 DVDD.n5976 2.30804
R1770 DVDD.n5972 DVDD.n35 2.30804
R1771 DVDD.n5970 DVDD.n5969 2.30804
R1772 DVDD.n5965 DVDD.n38 2.30804
R1773 DVDD.n5963 DVDD.n5962 2.30804
R1774 DVDD.n5958 DVDD.n40 2.30804
R1775 DVDD.n5956 DVDD.n5955 2.30804
R1776 DVDD.n5879 DVDD.n5878 2.30804
R1777 DVDD.n4812 DVDD.n106 2.30804
R1778 DVDD.n4816 DVDD.n107 2.30804
R1779 DVDD.n4820 DVDD.n108 2.30804
R1780 DVDD.n4824 DVDD.n109 2.30804
R1781 DVDD.n4828 DVDD.n110 2.30804
R1782 DVDD.n4832 DVDD.n111 2.30804
R1783 DVDD.n4836 DVDD.n112 2.30804
R1784 DVDD.n4840 DVDD.n113 2.30804
R1785 DVDD.n4844 DVDD.n114 2.30804
R1786 DVDD.n4783 DVDD.n115 2.30804
R1787 DVDD.n4779 DVDD.n116 2.30804
R1788 DVDD.n4775 DVDD.n117 2.30804
R1789 DVDD.n4771 DVDD.n118 2.30804
R1790 DVDD.n4767 DVDD.n119 2.30804
R1791 DVDD.n4763 DVDD.n120 2.30804
R1792 DVDD.n4759 DVDD.n121 2.30804
R1793 DVDD.n4755 DVDD.n122 2.30804
R1794 DVDD.n4751 DVDD.n123 2.30804
R1795 DVDD.n4747 DVDD.n124 2.30804
R1796 DVDD.n4743 DVDD.n125 2.30804
R1797 DVDD.n3353 DVDD.n126 2.30804
R1798 DVDD.n3349 DVDD.n127 2.30804
R1799 DVDD.n3345 DVDD.n128 2.30804
R1800 DVDD.n3341 DVDD.n129 2.30804
R1801 DVDD.n3337 DVDD.n130 2.30804
R1802 DVDD.n3333 DVDD.n131 2.30804
R1803 DVDD.n3329 DVDD.n132 2.30804
R1804 DVDD.n3325 DVDD.n133 2.30804
R1805 DVDD.n3321 DVDD.n134 2.30804
R1806 DVDD.n3317 DVDD.n135 2.30804
R1807 DVDD.n3313 DVDD.n136 2.30804
R1808 DVDD.n3308 DVDD.n137 2.30804
R1809 DVDD.n3304 DVDD.n138 2.30804
R1810 DVDD.n3300 DVDD.n139 2.30804
R1811 DVDD.n3296 DVDD.n140 2.30804
R1812 DVDD.n3292 DVDD.n141 2.30804
R1813 DVDD.n3288 DVDD.n142 2.30804
R1814 DVDD.n3284 DVDD.n143 2.30804
R1815 DVDD.n3280 DVDD.n144 2.30804
R1816 DVDD.n3276 DVDD.n145 2.30804
R1817 DVDD.n3272 DVDD.n146 2.30804
R1818 DVDD.n3268 DVDD.n147 2.30804
R1819 DVDD.n3264 DVDD.n148 2.30804
R1820 DVDD.n3260 DVDD.n149 2.30804
R1821 DVDD.n5762 DVDD.n150 2.30804
R1822 DVDD.n5766 DVDD.n151 2.30804
R1823 DVDD.n5770 DVDD.n152 2.30804
R1824 DVDD.n5774 DVDD.n153 2.30804
R1825 DVDD.n5778 DVDD.n154 2.30804
R1826 DVDD.n5782 DVDD.n155 2.30804
R1827 DVDD.n5786 DVDD.n156 2.30804
R1828 DVDD.n5790 DVDD.n157 2.30804
R1829 DVDD.n5794 DVDD.n158 2.30804
R1830 DVDD.n5798 DVDD.n159 2.30804
R1831 DVDD.n5802 DVDD.n160 2.30804
R1832 DVDD.n5804 DVDD.n161 2.30804
R1833 DVDD.n5812 DVDD.n162 2.30804
R1834 DVDD.n5816 DVDD.n163 2.30804
R1835 DVDD.n5820 DVDD.n164 2.30804
R1836 DVDD.n5824 DVDD.n165 2.30804
R1837 DVDD.n5828 DVDD.n166 2.30804
R1838 DVDD.n5875 DVDD.n168 2.30804
R1839 DVDD.n5830 DVDD.n166 2.30804
R1840 DVDD.n5827 DVDD.n165 2.30804
R1841 DVDD.n5823 DVDD.n164 2.30804
R1842 DVDD.n5819 DVDD.n163 2.30804
R1843 DVDD.n5815 DVDD.n162 2.30804
R1844 DVDD.n5811 DVDD.n161 2.30804
R1845 DVDD.n5805 DVDD.n160 2.30804
R1846 DVDD.n5801 DVDD.n159 2.30804
R1847 DVDD.n5797 DVDD.n158 2.30804
R1848 DVDD.n5793 DVDD.n157 2.30804
R1849 DVDD.n5789 DVDD.n156 2.30804
R1850 DVDD.n5785 DVDD.n155 2.30804
R1851 DVDD.n5781 DVDD.n154 2.30804
R1852 DVDD.n5777 DVDD.n153 2.30804
R1853 DVDD.n5773 DVDD.n152 2.30804
R1854 DVDD.n5769 DVDD.n151 2.30804
R1855 DVDD.n5765 DVDD.n150 2.30804
R1856 DVDD.n5761 DVDD.n149 2.30804
R1857 DVDD.n3261 DVDD.n148 2.30804
R1858 DVDD.n3265 DVDD.n147 2.30804
R1859 DVDD.n3269 DVDD.n146 2.30804
R1860 DVDD.n3273 DVDD.n145 2.30804
R1861 DVDD.n3277 DVDD.n144 2.30804
R1862 DVDD.n3281 DVDD.n143 2.30804
R1863 DVDD.n3285 DVDD.n142 2.30804
R1864 DVDD.n3289 DVDD.n141 2.30804
R1865 DVDD.n3293 DVDD.n140 2.30804
R1866 DVDD.n3297 DVDD.n139 2.30804
R1867 DVDD.n3301 DVDD.n138 2.30804
R1868 DVDD.n3258 DVDD.n137 2.30804
R1869 DVDD.n3309 DVDD.n136 2.30804
R1870 DVDD.n3314 DVDD.n135 2.30804
R1871 DVDD.n3318 DVDD.n134 2.30804
R1872 DVDD.n3322 DVDD.n133 2.30804
R1873 DVDD.n3326 DVDD.n132 2.30804
R1874 DVDD.n3330 DVDD.n131 2.30804
R1875 DVDD.n3334 DVDD.n130 2.30804
R1876 DVDD.n3338 DVDD.n129 2.30804
R1877 DVDD.n3342 DVDD.n128 2.30804
R1878 DVDD.n3346 DVDD.n127 2.30804
R1879 DVDD.n3350 DVDD.n126 2.30804
R1880 DVDD.n3352 DVDD.n125 2.30804
R1881 DVDD.n4744 DVDD.n124 2.30804
R1882 DVDD.n4748 DVDD.n123 2.30804
R1883 DVDD.n4752 DVDD.n122 2.30804
R1884 DVDD.n4756 DVDD.n121 2.30804
R1885 DVDD.n4760 DVDD.n120 2.30804
R1886 DVDD.n4764 DVDD.n119 2.30804
R1887 DVDD.n4768 DVDD.n118 2.30804
R1888 DVDD.n4772 DVDD.n117 2.30804
R1889 DVDD.n4776 DVDD.n116 2.30804
R1890 DVDD.n4780 DVDD.n115 2.30804
R1891 DVDD.n4784 DVDD.n114 2.30804
R1892 DVDD.n4843 DVDD.n113 2.30804
R1893 DVDD.n4839 DVDD.n112 2.30804
R1894 DVDD.n4835 DVDD.n111 2.30804
R1895 DVDD.n4831 DVDD.n110 2.30804
R1896 DVDD.n4827 DVDD.n109 2.30804
R1897 DVDD.n4823 DVDD.n108 2.30804
R1898 DVDD.n4819 DVDD.n107 2.30804
R1899 DVDD.n4815 DVDD.n106 2.30804
R1900 DVDD.n5878 DVDD.n105 2.30804
R1901 DVDD.n5833 DVDD.n168 2.30804
R1902 DVDD.n5951 DVDD.n42 2.30804
R1903 DVDD.n5957 DVDD.n5956 2.30804
R1904 DVDD.n40 DVDD.n39 2.30804
R1905 DVDD.n5964 DVDD.n5963 2.30804
R1906 DVDD.n38 DVDD.n36 2.30804
R1907 DVDD.n5971 DVDD.n5970 2.30804
R1908 DVDD.n35 DVDD.n33 2.30804
R1909 DVDD.n5978 DVDD.n5977 2.30804
R1910 DVDD.n5981 DVDD.n5980 2.30804
R1911 DVDD.n4561 DVDD.n4560 2.30804
R1912 DVDD.n4566 DVDD.n4565 2.30804
R1913 DVDD.n4559 DVDD.n4557 2.30804
R1914 DVDD.n4573 DVDD.n4572 2.30804
R1915 DVDD.n4556 DVDD.n4554 2.30804
R1916 DVDD.n4580 DVDD.n4579 2.30804
R1917 DVDD.n4553 DVDD.n4551 2.30804
R1918 DVDD.n4587 DVDD.n4586 2.30804
R1919 DVDD.n4550 DVDD.n4548 2.30804
R1920 DVDD.n4594 DVDD.n4593 2.30804
R1921 DVDD.n4547 DVDD.n3424 2.30804
R1922 DVDD.n4601 DVDD.n4600 2.30804
R1923 DVDD.n3422 DVDD.n3420 2.30804
R1924 DVDD.n4608 DVDD.n4607 2.30804
R1925 DVDD.n3419 DVDD.n3417 2.30804
R1926 DVDD.n4615 DVDD.n4614 2.30804
R1927 DVDD.n3416 DVDD.n3414 2.30804
R1928 DVDD.n4622 DVDD.n4621 2.30804
R1929 DVDD.n3413 DVDD.n3411 2.30804
R1930 DVDD.n4629 DVDD.n4628 2.30804
R1931 DVDD.n3410 DVDD.n3408 2.30804
R1932 DVDD.n4636 DVDD.n4635 2.30804
R1933 DVDD.n3407 DVDD.n3406 2.30804
R1934 DVDD.n3404 DVDD.n3396 2.30804
R1935 DVDD.n4645 DVDD.n4644 2.30804
R1936 DVDD.n3394 DVDD.n3392 2.30804
R1937 DVDD.n4652 DVDD.n4651 2.30804
R1938 DVDD.n3391 DVDD.n3389 2.30804
R1939 DVDD.n4659 DVDD.n4658 2.30804
R1940 DVDD.n3388 DVDD.n3386 2.30804
R1941 DVDD.n4666 DVDD.n4665 2.30804
R1942 DVDD.n3385 DVDD.n3383 2.30804
R1943 DVDD.n4673 DVDD.n4672 2.30804
R1944 DVDD.n3382 DVDD.n3380 2.30804
R1945 DVDD.n4680 DVDD.n4679 2.30804
R1946 DVDD.n4277 DVDD.n3379 2.30804
R1947 DVDD.n4281 DVDD.n4280 2.30804
R1948 DVDD.n4276 DVDD.n4274 2.30804
R1949 DVDD.n4288 DVDD.n4287 2.30804
R1950 DVDD.n4273 DVDD.n4271 2.30804
R1951 DVDD.n4295 DVDD.n4294 2.30804
R1952 DVDD.n4270 DVDD.n4268 2.30804
R1953 DVDD.n4302 DVDD.n4301 2.30804
R1954 DVDD.n4267 DVDD.n4265 2.30804
R1955 DVDD.n4309 DVDD.n4308 2.30804
R1956 DVDD.n4264 DVDD.n4262 2.30804
R1957 DVDD.n4316 DVDD.n4315 2.30804
R1958 DVDD.n4260 DVDD.n4259 2.30804
R1959 DVDD.n4255 DVDD.n4218 2.30804
R1960 DVDD.n4253 DVDD.n4252 2.30804
R1961 DVDD.n4248 DVDD.n4247 2.30804
R1962 DVDD.n4245 DVDD.n4244 2.30804
R1963 DVDD.n4240 DVDD.n4239 2.30804
R1964 DVDD.n4237 DVDD.n4236 2.30804
R1965 DVDD.n4232 DVDD.n4231 2.30804
R1966 DVDD.n4229 DVDD.n4228 2.30804
R1967 DVDD.n5832 DVDD.n167 2.29384
R1968 DVDD.n3185 DVDD.n3181 2.2505
R1969 DVDD.n3188 DVDD.n3187 2.2505
R1970 DVDD.n3186 DVDD.n3183 2.2505
R1971 DVDD.n3179 DVDD.n3178 2.2505
R1972 DVDD.n3198 DVDD.n3197 2.2505
R1973 DVDD.n3199 DVDD.n3169 2.2505
R1974 DVDD.n3240 DVDD.n3239 2.2505
R1975 DVDD.n3238 DVDD.n3237 2.2505
R1976 DVDD.n3201 DVDD.n3200 2.2505
R1977 DVDD.n3232 DVDD.n3231 2.2505
R1978 DVDD.n3230 DVDD.n170 2.2505
R1979 DVDD.n3206 DVDD.n171 2.2505
R1980 DVDD.n3213 DVDD.n3211 2.2505
R1981 DVDD.n3224 DVDD.n3223 2.2505
R1982 DVDD.n3222 DVDD.n3221 2.2505
R1983 DVDD.n3215 DVDD.n3214 2.2505
R1984 DVDD.n5321 DVDD.n725 2.2505
R1985 DVDD.n5325 DVDD.n5324 2.2505
R1986 DVDD.n5326 DVDD.n723 2.2505
R1987 DVDD.n5328 DVDD.n5327 2.2505
R1988 DVDD.n724 DVDD.n716 2.2505
R1989 DVDD.n5337 DVDD.n5336 2.2505
R1990 DVDD.n5338 DVDD.n712 2.2505
R1991 DVDD.n5341 DVDD.n5340 2.2505
R1992 DVDD.n5339 DVDD.n715 2.2505
R1993 DVDD.n713 DVDD.n707 2.2505
R1994 DVDD.n5351 DVDD.n5350 2.2505
R1995 DVDD.n5352 DVDD.n233 2.2505
R1996 DVDD.n5357 DVDD.n5356 2.2505
R1997 DVDD.n5358 DVDD.n705 2.2505
R1998 DVDD.n5360 DVDD.n5359 2.2505
R1999 DVDD.n701 DVDD.n700 2.2505
R2000 DVDD.n5366 DVDD.n5365 2.2505
R2001 DVDD.n3888 DVDD.n3852 2.2505
R2002 DVDD.n3887 DVDD.n3886 2.2505
R2003 DVDD.n3885 DVDD.n3853 2.2505
R2004 DVDD.n3884 DVDD.n3883 2.2505
R2005 DVDD.n3882 DVDD.n3854 2.2505
R2006 DVDD.n3881 DVDD.n3880 2.2505
R2007 DVDD.n3879 DVDD.n3878 2.2505
R2008 DVDD.n3877 DVDD.n3876 2.2505
R2009 DVDD.n3875 DVDD.n3874 2.2505
R2010 DVDD.n3873 DVDD.n3872 2.2505
R2011 DVDD.n3871 DVDD.n3870 2.2505
R2012 DVDD.n3869 DVDD.n3868 2.2505
R2013 DVDD.n3867 DVDD.n3866 2.2505
R2014 DVDD.n3865 DVDD.n3864 2.2505
R2015 DVDD.n3863 DVDD.n3862 2.2505
R2016 DVDD.n3861 DVDD.n3860 2.2505
R2017 DVDD.n3859 DVDD.n3858 2.2505
R2018 DVDD.n3857 DVDD.n3856 2.2505
R2019 DVDD.n3855 DVDD.n3587 2.2505
R2020 DVDD.n3891 DVDD.n3890 2.2505
R2021 DVDD.n4537 DVDD.n4536 2.2505
R2022 DVDD.n4504 DVDD.n3428 2.2505
R2023 DVDD.n4507 DVDD.n4503 2.2505
R2024 DVDD.n4515 DVDD.n4514 2.2505
R2025 DVDD.n4519 DVDD.n4517 2.2505
R2026 DVDD.n4516 DVDD.n3169 2.2505
R2027 DVDD.n3150 DVDD.n3149 2.2505
R2028 DVDD.n4871 DVDD.n4870 2.2505
R2029 DVDD.n4875 DVDD.n4873 2.2505
R2030 DVDD.n4872 DVDD.n3139 2.2505
R2031 DVDD.n4884 DVDD.n174 2.2505
R2032 DVDD.n5757 DVDD.n5756 2.2505
R2033 DVDD.n177 DVDD.n175 2.2505
R2034 DVDD.n3133 DVDD.n3131 2.2505
R2035 DVDD.n4896 DVDD.n4895 2.2505
R2036 DVDD.n4898 DVDD.n4897 2.2505
R2037 DVDD.n5321 DVDD.n727 2.2505
R2038 DVDD.n5086 DVDD.n4903 2.2505
R2039 DVDD.n5088 DVDD.n5087 2.2505
R2040 DVDD.n5104 DVDD.n5103 2.2505
R2041 DVDD.n5105 DVDD.n4912 2.2505
R2042 DVDD.n5106 DVDD.n4913 2.2505
R2043 DVDD.n5107 DVDD.n4914 2.2505
R2044 DVDD.n5112 DVDD.n5108 2.2505
R2045 DVDD.n5111 DVDD.n5079 2.2505
R2046 DVDD.n5121 DVDD.n5120 2.2505
R2047 DVDD.n5122 DVDD.n4922 2.2505
R2048 DVDD.n5123 DVDD.n233 2.2505
R2049 DVDD.n5124 DVDD.n4923 2.2505
R2050 DVDD.n5130 DVDD.n5125 2.2505
R2051 DVDD.n5139 DVDD.n5138 2.2505
R2052 DVDD.n5140 DVDD.n4933 2.2505
R2053 DVDD.n5141 DVDD.n4934 2.2505
R2054 DVDD.n5472 DVDD.n5471 2.2505
R2055 DVDD.n5706 DVDD.n5705 2.2505
R2056 DVDD.n3935 DVDD.n3934 2.2505
R2057 DVDD.n3933 DVDD.n3932 2.2505
R2058 DVDD.n3931 DVDD.n3930 2.2505
R2059 DVDD.n3929 DVDD.n3928 2.2505
R2060 DVDD.n3927 DVDD.n3926 2.2505
R2061 DVDD.n3925 DVDD.n3924 2.2505
R2062 DVDD.n3923 DVDD.n3922 2.2505
R2063 DVDD.n3921 DVDD.n3920 2.2505
R2064 DVDD.n3662 DVDD.n3660 2.2505
R2065 DVDD.n3954 DVDD.n3953 2.2505
R2066 DVDD.n3952 DVDD.n3661 2.2505
R2067 DVDD.n3951 DVDD.n3950 2.2505
R2068 DVDD.n3949 DVDD.n3948 2.2505
R2069 DVDD.n3947 DVDD.n3663 2.2505
R2070 DVDD.n3946 DVDD.n3945 2.2505
R2071 DVDD.n3944 DVDD.n3664 2.2505
R2072 DVDD.n3943 DVDD.n3942 2.2505
R2073 DVDD.n3941 DVDD.n3665 2.2505
R2074 DVDD.n3940 DVDD.n3939 2.2505
R2075 DVDD.n3938 DVDD.n3919 2.2505
R2076 DVDD.n4691 DVDD.n3370 2.2505
R2077 DVDD.n4694 DVDD.n4693 2.2505
R2078 DVDD.n4692 DVDD.n3372 2.2505
R2079 DVDD.n3368 DVDD.n3367 2.2505
R2080 DVDD.n4704 DVDD.n4703 2.2505
R2081 DVDD.n4705 DVDD.n3169 2.2505
R2082 DVDD.n4707 DVDD.n4706 2.2505
R2083 DVDD.n3365 DVDD.n3364 2.2505
R2084 DVDD.n4715 DVDD.n4714 2.2505
R2085 DVDD.n4717 DVDD.n4716 2.2505
R2086 DVDD.n4718 DVDD.n3256 2.2505
R2087 DVDD.n4739 DVDD.n4738 2.2505
R2088 DVDD.n4737 DVDD.n3356 2.2505
R2089 DVDD.n4726 DVDD.n3358 2.2505
R2090 DVDD.n4727 DVDD.n4725 2.2505
R2091 DVDD.n4729 DVDD.n4728 2.2505
R2092 DVDD.n5321 DVDD.n3078 2.2505
R2093 DVDD.n3077 DVDD.n3076 2.2505
R2094 DVDD.n3074 DVDD.n3073 2.2505
R2095 DVDD.n3072 DVDD.n3071 2.2505
R2096 DVDD.n3070 DVDD.n3069 2.2505
R2097 DVDD.n3068 DVDD.n3067 2.2505
R2098 DVDD.n3066 DVDD.n3065 2.2505
R2099 DVDD.n3063 DVDD.n3062 2.2505
R2100 DVDD.n3061 DVDD.n3060 2.2505
R2101 DVDD.n3059 DVDD.n3058 2.2505
R2102 DVDD.n3057 DVDD.n3056 2.2505
R2103 DVDD.n3054 DVDD.n233 2.2505
R2104 DVDD.n3053 DVDD.n3052 2.2505
R2105 DVDD.n737 DVDD.n735 2.2505
R2106 DVDD.n743 DVDD.n742 2.2505
R2107 DVDD.n3044 DVDD.n3043 2.2505
R2108 DVDD.n3042 DVDD.n740 2.2505
R2109 DVDD.n3503 DVDD.n3502 2.2505
R2110 DVDD.n3486 DVDD.n3484 2.2505
R2111 DVDD.n3492 DVDD.n3490 2.2505
R2112 DVDD.n3497 DVDD.n3496 2.2505
R2113 DVDD.n3495 DVDD.n3494 2.2505
R2114 DVDD.n3247 DVDD.n3169 2.2505
R2115 DVDD.n4858 DVDD.n4857 2.2505
R2116 DVDD.n4856 DVDD.n4855 2.2505
R2117 DVDD.n3249 DVDD.n3248 2.2505
R2118 DVDD.n4850 DVDD.n4849 2.2505
R2119 DVDD.n4848 DVDD.n3254 2.2505
R2120 DVDD.n4811 DVDD.n4810 2.2505
R2121 DVDD.n4809 DVDD.n4787 2.2505
R2122 DVDD.n4800 DVDD.n4790 2.2505
R2123 DVDD.n4804 DVDD.n4803 2.2505
R2124 DVDD.n4802 DVDD.n4801 2.2505
R2125 DVDD.n5321 DVDD.n3128 2.2505
R2126 DVDD.n3127 DVDD.n3126 2.2505
R2127 DVDD.n3082 DVDD.n3081 2.2505
R2128 DVDD.n3121 DVDD.n3120 2.2505
R2129 DVDD.n3119 DVDD.n3087 2.2505
R2130 DVDD.n3118 DVDD.n3117 2.2505
R2131 DVDD.n3096 DVDD.n3088 2.2505
R2132 DVDD.n3111 DVDD.n3110 2.2505
R2133 DVDD.n3109 DVDD.n3097 2.2505
R2134 DVDD.n3108 DVDD.n3107 2.2505
R2135 DVDD.n3100 DVDD.n3098 2.2505
R2136 DVDD.n235 DVDD.n233 2.2505
R2137 DVDD.n5725 DVDD.n5724 2.2505
R2138 DVDD.n5723 DVDD.n5722 2.2505
R2139 DVDD.n237 DVDD.n236 2.2505
R2140 DVDD.n5717 DVDD.n5716 2.2505
R2141 DVDD.n5715 DVDD.n240 2.2505
R2142 DVDD.n346 DVDD.n324 2.25007
R2143 DVDD.n1265 DVDD.n1195 2.25007
R2144 DVDD.n2529 DVDD.n2528 2.25007
R2145 DVDD.n4000 DVDD.n3999 2.24901
R2146 DVDD.n4494 DVDD.n3432 2.24901
R2147 DVDD.n2603 DVDD.n2602 2.24901
R2148 DVDD.n3837 DVDD.n3834 2.24648
R2149 DVDD.n3839 DVDD.n3838 2.24648
R2150 DVDD.n3524 DVDD.n3521 2.24648
R2151 DVDD.n3674 DVDD.n3672 2.24648
R2152 DVDD.n3680 DVDD.n3670 2.24648
R2153 DVDD.n3903 DVDD.n3683 2.24648
R2154 DVDD.n3848 DVDD.n3684 2.24648
R2155 DVDD.n3896 DVDD.n3895 2.24648
R2156 DVDD.n552 DVDD.n551 2.24648
R2157 DVDD.n550 DVDD.n547 2.24648
R2158 DVDD.n3622 DVDD.n3617 2.24581
R2159 DVDD.n3627 DVDD.n3626 2.24581
R2160 DVDD.n3622 DVDD.n3618 2.24581
R2161 DVDD.n3627 DVDD.n3625 2.24581
R2162 DVDD.n3622 DVDD.n3619 2.24581
R2163 DVDD.n3627 DVDD.n3624 2.24581
R2164 DVDD.n3622 DVDD.n3620 2.24581
R2165 DVDD.n3627 DVDD.n3623 2.24581
R2166 DVDD.n3622 DVDD.n3621 2.24581
R2167 DVDD.n3627 DVDD.n3616 2.24581
R2168 DVDD.n5278 DVDD.n4935 2.24581
R2169 DVDD.n5246 DVDD.n4936 2.24581
R2170 DVDD.n5278 DVDD.n5268 2.24581
R2171 DVDD.n5248 DVDD.n4936 2.24581
R2172 DVDD.n5278 DVDD.n5269 2.24581
R2173 DVDD.n5250 DVDD.n4936 2.24581
R2174 DVDD.n5278 DVDD.n5270 2.24581
R2175 DVDD.n5252 DVDD.n4936 2.24581
R2176 DVDD.n5278 DVDD.n5271 2.24581
R2177 DVDD.n5254 DVDD.n4936 2.24581
R2178 DVDD.n5278 DVDD.n5272 2.24581
R2179 DVDD.n5256 DVDD.n4936 2.24581
R2180 DVDD.n5278 DVDD.n5273 2.24581
R2181 DVDD.n5258 DVDD.n4936 2.24581
R2182 DVDD.n5278 DVDD.n5274 2.24581
R2183 DVDD.n5260 DVDD.n4936 2.24581
R2184 DVDD.n5278 DVDD.n5275 2.24581
R2185 DVDD.n5262 DVDD.n4936 2.24581
R2186 DVDD.n5278 DVDD.n5276 2.24581
R2187 DVDD.n5264 DVDD.n4936 2.24581
R2188 DVDD.n5278 DVDD.n5277 2.24581
R2189 DVDD.n5266 DVDD.n4936 2.24581
R2190 DVDD.n5279 DVDD.n5278 2.24581
R2191 DVDD.n5016 DVDD.n296 2.24581
R2192 DVDD.n5023 DVDD.n296 2.24581
R2193 DVDD.n299 DVDD.n296 2.24581
R2194 DVDD.n300 DVDD.n296 2.24581
R2195 DVDD.n310 DVDD.n296 2.24581
R2196 DVDD.n355 DVDD.n311 2.24581
R2197 DVDD.n327 DVDD.n312 2.24581
R2198 DVDD.n355 DVDD.n347 2.24581
R2199 DVDD.n329 DVDD.n312 2.24581
R2200 DVDD.n332 DVDD.n313 2.24581
R2201 DVDD.n355 DVDD.n348 2.24581
R2202 DVDD.n334 DVDD.n312 2.24581
R2203 DVDD.n355 DVDD.n349 2.24581
R2204 DVDD.n336 DVDD.n312 2.24581
R2205 DVDD.n355 DVDD.n350 2.24581
R2206 DVDD.n338 DVDD.n312 2.24581
R2207 DVDD.n355 DVDD.n351 2.24581
R2208 DVDD.n340 DVDD.n312 2.24581
R2209 DVDD.n355 DVDD.n352 2.24581
R2210 DVDD.n355 DVDD.n353 2.24581
R2211 DVDD.n343 DVDD.n312 2.24581
R2212 DVDD.n355 DVDD.n354 2.24581
R2213 DVDD.n356 DVDD.n355 2.24581
R2214 DVDD.n1564 DVDD.n1553 2.24581
R2215 DVDD.n1548 DVDD.n1547 2.24581
R2216 DVDD.n1564 DVDD.n1554 2.24581
R2217 DVDD.n1564 DVDD.n1555 2.24581
R2218 DVDD.n1548 DVDD.n1546 2.24581
R2219 DVDD.n1564 DVDD.n1556 2.24581
R2220 DVDD.n1564 DVDD.n1557 2.24581
R2221 DVDD.n1548 DVDD.n1545 2.24581
R2222 DVDD.n1564 DVDD.n1558 2.24581
R2223 DVDD.n1564 DVDD.n1559 2.24581
R2224 DVDD.n1548 DVDD.n1544 2.24581
R2225 DVDD.n1564 DVDD.n1560 2.24581
R2226 DVDD.n1564 DVDD.n1561 2.24581
R2227 DVDD.n1548 DVDD.n1543 2.24581
R2228 DVDD.n1564 DVDD.n1562 2.24581
R2229 DVDD.n1564 DVDD.n1563 2.24581
R2230 DVDD.n1548 DVDD.n1542 2.24581
R2231 DVDD.n1564 DVDD.n1541 2.24581
R2232 DVDD.n2373 DVDD.n1196 2.24581
R2233 DVDD.n2373 DVDD.n1197 2.24581
R2234 DVDD.n2369 DVDD.n1272 2.24581
R2235 DVDD.n2373 DVDD.n1198 2.24581
R2236 DVDD.n2369 DVDD.n1271 2.24581
R2237 DVDD.n2373 DVDD.n1199 2.24581
R2238 DVDD.n2369 DVDD.n1270 2.24581
R2239 DVDD.n2373 DVDD.n1200 2.24581
R2240 DVDD.n2369 DVDD.n1269 2.24581
R2241 DVDD.n2373 DVDD.n1201 2.24581
R2242 DVDD.n2369 DVDD.n1268 2.24581
R2243 DVDD.n2373 DVDD.n1202 2.24581
R2244 DVDD.n2373 DVDD.n1203 2.24581
R2245 DVDD.n2369 DVDD.n1267 2.24581
R2246 DVDD.n2373 DVDD.n1204 2.24581
R2247 DVDD.n2373 DVDD.n1205 2.24581
R2248 DVDD.n2369 DVDD.n1266 2.24581
R2249 DVDD.n2373 DVDD.n1194 2.24581
R2250 DVDD.n2369 DVDD.n1206 2.24581
R2251 DVDD.n1041 DVDD.n1017 2.24581
R2252 DVDD.n2564 DVDD.n1039 2.24581
R2253 DVDD.n2512 DVDD.n1017 2.24581
R2254 DVDD.n1037 DVDD.n1017 2.24581
R2255 DVDD.n2564 DVDD.n1035 2.24581
R2256 DVDD.n2545 DVDD.n1017 2.24581
R2257 DVDD.n2564 DVDD.n2547 2.24581
R2258 DVDD.n2543 DVDD.n1017 2.24581
R2259 DVDD.n2560 DVDD.n1015 2.24581
R2260 DVDD.n1032 DVDD.n1017 2.24581
R2261 DVDD.n2564 DVDD.n1030 2.24581
R2262 DVDD.n1026 DVDD.n1015 2.24581
R2263 DVDD.n1028 DVDD.n1017 2.24581
R2264 DVDD.n2564 DVDD.n1025 2.24581
R2265 DVDD.n2562 DVDD.n1015 2.24581
R2266 DVDD.n1022 DVDD.n1017 2.24581
R2267 DVDD.n2564 DVDD.n1020 2.24581
R2268 DVDD.n517 DVDD.n510 2.24581
R2269 DVDD.n2601 DVDD.n2598 2.24581
R2270 DVDD.n5568 DVDD.n514 2.24581
R2271 DVDD.n519 DVDD.n510 2.24581
R2272 DVDD.n2601 DVDD.n2600 2.24581
R2273 DVDD.n5568 DVDD.n512 2.24581
R2274 DVDD.n521 DVDD.n510 2.24581
R2275 DVDD.n2601 DVDD.n523 2.24581
R2276 DVDD.n4491 DVDD.n3442 2.24581
R2277 DVDD.n4493 DVDD.n3437 2.24581
R2278 DVDD.n4491 DVDD.n3443 2.24581
R2279 DVDD.n4493 DVDD.n3436 2.24581
R2280 DVDD.n4491 DVDD.n4490 2.24581
R2281 DVDD.n3445 DVDD.n3444 2.24581
R2282 DVDD.n4488 DVDD.n4487 2.24581
R2283 DVDD.n3445 DVDD.n3440 2.24581
R2284 DVDD.n4488 DVDD.n3431 2.24581
R2285 DVDD.n3842 DVDD.n3836 2.24442
R2286 DVDD.n3840 DVDD.n3832 2.24442
R2287 DVDD.n3833 DVDD.n3523 2.24442
R2288 DVDD.n3901 DVDD.n3685 2.24442
R2289 DVDD.n3899 DVDD.n3898 2.24442
R2290 DVDD.n2027 DVDD.n563 2.24442
R2291 DVDD.n5505 DVDD.n567 2.24442
R2292 DVDD.n5505 DVDD.n5504 2.24442
R2293 DVDD.n1700 DVDD.n574 2.24442
R2294 DVDD.n598 DVDD.n578 2.24442
R2295 DVDD.n570 DVDD.n566 2.24442
R2296 DVDD.n572 DVDD.n566 2.24442
R2297 DVDD.n554 DVDD.n549 2.24442
R2298 DVDD.n5523 DVDD.n548 2.24442
R2299 DVDD.n1789 DVDD.n559 2.24442
R2300 DVDD.n3893 DVDD.n3851 2.23892
R2301 DVDD.n3894 DVDD.n3850 2.23892
R2302 DVDD.n4194 DVDD.n3527 2.23892
R2303 DVDD.n4195 DVDD.n4186 2.23892
R2304 DVDD.n4184 DVDD.n4182 2.23892
R2305 DVDD.n3525 DVDD.n3520 2.23892
R2306 DVDD.n4199 DVDD.n3522 2.23892
R2307 DVDD.n3679 DVDD.n3673 2.23892
R2308 DVDD.n3677 DVDD.n3675 2.23892
R2309 DVDD.n3681 DVDD.n3669 2.23892
R2310 DVDD.n3911 DVDD.n3671 2.23892
R2311 DVDD.n3904 DVDD.n3902 2.23892
R2312 DVDD.n3906 DVDD.n3905 2.23892
R2313 DVDD.n4204 DVDD.n3518 2.23892
R2314 DVDD.n4202 DVDD.n3510 2.23892
R2315 DVDD.n3916 DVDD.n3666 2.23892
R2316 DVDD.n3917 DVDD.n3667 2.23892
R2317 DVDD.n4206 DVDD.n3508 2.23892
R2318 DVDD.n4115 DVDD.n3554 2.23714
R2319 DVDD.n4112 DVDD.n4111 2.23714
R2320 DVDD.n4115 DVDD.n3555 2.23714
R2321 DVDD.n4112 DVDD.n4110 2.23714
R2322 DVDD.n4115 DVDD.n3556 2.23714
R2323 DVDD.n4112 DVDD.n4109 2.23714
R2324 DVDD.n4115 DVDD.n3557 2.23714
R2325 DVDD.n4113 DVDD.n4112 2.23714
R2326 DVDD.n4115 DVDD.n4114 2.23714
R2327 DVDD.n4112 DVDD.n3551 2.23714
R2328 DVDD.n5368 DVDD.n696 2.23714
R2329 DVDD.n5391 DVDD.n5369 2.23714
R2330 DVDD.n5370 DVDD.n696 2.23714
R2331 DVDD.n5391 DVDD.n5371 2.23714
R2332 DVDD.n5372 DVDD.n696 2.23714
R2333 DVDD.n5391 DVDD.n5373 2.23714
R2334 DVDD.n5374 DVDD.n696 2.23714
R2335 DVDD.n5391 DVDD.n5375 2.23714
R2336 DVDD.n5376 DVDD.n696 2.23714
R2337 DVDD.n5391 DVDD.n5377 2.23714
R2338 DVDD.n5378 DVDD.n696 2.23714
R2339 DVDD.n5391 DVDD.n5379 2.23714
R2340 DVDD.n5380 DVDD.n696 2.23714
R2341 DVDD.n5391 DVDD.n5381 2.23714
R2342 DVDD.n5382 DVDD.n696 2.23714
R2343 DVDD.n5391 DVDD.n5383 2.23714
R2344 DVDD.n5384 DVDD.n696 2.23714
R2345 DVDD.n5391 DVDD.n5385 2.23714
R2346 DVDD.n5386 DVDD.n696 2.23714
R2347 DVDD.n5391 DVDD.n5387 2.23714
R2348 DVDD.n5389 DVDD.n696 2.23714
R2349 DVDD.n5391 DVDD.n5390 2.23714
R2350 DVDD.n5388 DVDD.n696 2.23714
R2351 DVDD.n5484 DVDD.n604 2.23714
R2352 DVDD.n5485 DVDD.n605 2.23714
R2353 DVDD.n5486 DVDD.n604 2.23714
R2354 DVDD.n5487 DVDD.n605 2.23714
R2355 DVDD.n5488 DVDD.n604 2.23714
R2356 DVDD.n5489 DVDD.n605 2.23714
R2357 DVDD.n5490 DVDD.n604 2.23714
R2358 DVDD.n5491 DVDD.n605 2.23714
R2359 DVDD.n5492 DVDD.n604 2.23714
R2360 DVDD.n5493 DVDD.n605 2.23714
R2361 DVDD.n5495 DVDD.n580 2.23714
R2362 DVDD.n5497 DVDD.n602 2.23714
R2363 DVDD.n601 DVDD.n580 2.23714
R2364 DVDD.n5497 DVDD.n600 2.23714
R2365 DVDD.n596 DVDD.n580 2.23714
R2366 DVDD.n5497 DVDD.n595 2.23714
R2367 DVDD.n594 DVDD.n580 2.23714
R2368 DVDD.n5497 DVDD.n593 2.23714
R2369 DVDD.n592 DVDD.n580 2.23714
R2370 DVDD.n5497 DVDD.n591 2.23714
R2371 DVDD.n590 DVDD.n580 2.23714
R2372 DVDD.n5497 DVDD.n589 2.23714
R2373 DVDD.n588 DVDD.n580 2.23714
R2374 DVDD.n5497 DVDD.n587 2.23714
R2375 DVDD.n5497 DVDD.n586 2.23714
R2376 DVDD.n585 DVDD.n580 2.23714
R2377 DVDD.n5497 DVDD.n584 2.23714
R2378 DVDD.n5497 DVDD.n583 2.23714
R2379 DVDD.n2236 DVDD.n1372 2.23714
R2380 DVDD.n1373 DVDD.n1370 2.23714
R2381 DVDD.n2236 DVDD.n1374 2.23714
R2382 DVDD.n2236 DVDD.n1375 2.23714
R2383 DVDD.n1376 DVDD.n1370 2.23714
R2384 DVDD.n2236 DVDD.n1377 2.23714
R2385 DVDD.n2236 DVDD.n1378 2.23714
R2386 DVDD.n1379 DVDD.n1370 2.23714
R2387 DVDD.n2236 DVDD.n1380 2.23714
R2388 DVDD.n2236 DVDD.n1381 2.23714
R2389 DVDD.n1382 DVDD.n1370 2.23714
R2390 DVDD.n2236 DVDD.n1383 2.23714
R2391 DVDD.n2236 DVDD.n1384 2.23714
R2392 DVDD.n1385 DVDD.n1370 2.23714
R2393 DVDD.n2236 DVDD.n1386 2.23714
R2394 DVDD.n2236 DVDD.n2230 2.23714
R2395 DVDD.n2234 DVDD.n1370 2.23714
R2396 DVDD.n2236 DVDD.n2235 2.23714
R2397 DVDD.n2456 DVDD.n1101 2.23714
R2398 DVDD.n2456 DVDD.n1102 2.23714
R2399 DVDD.n1103 DVDD.n1093 2.23714
R2400 DVDD.n2456 DVDD.n1104 2.23714
R2401 DVDD.n1105 DVDD.n1093 2.23714
R2402 DVDD.n2456 DVDD.n1106 2.23714
R2403 DVDD.n1107 DVDD.n1093 2.23714
R2404 DVDD.n2456 DVDD.n1108 2.23714
R2405 DVDD.n1109 DVDD.n1093 2.23714
R2406 DVDD.n2456 DVDD.n1110 2.23714
R2407 DVDD.n1111 DVDD.n1093 2.23714
R2408 DVDD.n2456 DVDD.n1112 2.23714
R2409 DVDD.n2456 DVDD.n1113 2.23714
R2410 DVDD.n1114 DVDD.n1093 2.23714
R2411 DVDD.n2456 DVDD.n1115 2.23714
R2412 DVDD.n2456 DVDD.n2451 2.23714
R2413 DVDD.n1116 DVDD.n1093 2.23714
R2414 DVDD.n2456 DVDD.n1098 2.23714
R2415 DVDD.n2454 DVDD.n1093 2.23714
R2416 DVDD.n2935 DVDD.n989 2.23714
R2417 DVDD.n1006 DVDD.n1001 2.23714
R2418 DVDD.n2935 DVDD.n990 2.23714
R2419 DVDD.n2935 DVDD.n991 2.23714
R2420 DVDD.n1006 DVDD.n1002 2.23714
R2421 DVDD.n2935 DVDD.n986 2.23714
R2422 DVDD.n1006 DVDD.n1000 2.23714
R2423 DVDD.n2935 DVDD.n985 2.23714
R2424 DVDD.n1006 DVDD.n999 2.23714
R2425 DVDD.n2935 DVDD.n993 2.23714
R2426 DVDD.n1006 DVDD.n1003 2.23714
R2427 DVDD.n1006 DVDD.n981 2.23714
R2428 DVDD.n2935 DVDD.n994 2.23714
R2429 DVDD.n1006 DVDD.n1004 2.23714
R2430 DVDD.n1006 DVDD.n998 2.23714
R2431 DVDD.n2935 DVDD.n996 2.23714
R2432 DVDD.n1006 DVDD.n1005 2.23714
R2433 DVDD.n2927 DVDD.n2574 2.23714
R2434 DVDD.n2930 DVDD.n2579 2.23714
R2435 DVDD.n2927 DVDD.n2926 2.23714
R2436 DVDD.n2927 DVDD.n2925 2.23714
R2437 DVDD.n2930 DVDD.n2581 2.23714
R2438 DVDD.n2927 DVDD.n2924 2.23714
R2439 DVDD.n2930 DVDD.n2582 2.23714
R2440 DVDD.n2928 DVDD.n2927 2.23714
R2441 DVDD.n5212 DVDD.n5202 2.23714
R2442 DVDD.n5215 DVDD.n5144 2.23714
R2443 DVDD.n5212 DVDD.n5203 2.23714
R2444 DVDD.n5215 DVDD.n5145 2.23714
R2445 DVDD.n5212 DVDD.n5204 2.23714
R2446 DVDD.n5215 DVDD.n5146 2.23714
R2447 DVDD.n5212 DVDD.n5205 2.23714
R2448 DVDD.n5215 DVDD.n5147 2.23714
R2449 DVDD.n5212 DVDD.n5206 2.23714
R2450 DVDD.n5215 DVDD.n5148 2.23714
R2451 DVDD.n5212 DVDD.n5207 2.23714
R2452 DVDD.n5215 DVDD.n5149 2.23714
R2453 DVDD.n5212 DVDD.n5208 2.23714
R2454 DVDD.n5215 DVDD.n5150 2.23714
R2455 DVDD.n5212 DVDD.n5209 2.23714
R2456 DVDD.n5215 DVDD.n5151 2.23714
R2457 DVDD.n5212 DVDD.n5210 2.23714
R2458 DVDD.n5215 DVDD.n5152 2.23714
R2459 DVDD.n5212 DVDD.n5211 2.23714
R2460 DVDD.n5215 DVDD.n5153 2.23714
R2461 DVDD.n5213 DVDD.n5212 2.23714
R2462 DVDD.n5215 DVDD.n5214 2.23714
R2463 DVDD.n5212 DVDD.n5154 2.23714
R2464 DVDD.n638 DVDD.n627 2.23714
R2465 DVDD.n5469 DVDD.n633 2.23714
R2466 DVDD.n638 DVDD.n637 2.23714
R2467 DVDD.n5469 DVDD.n632 2.23714
R2468 DVDD.n638 DVDD.n636 2.23714
R2469 DVDD.n5469 DVDD.n631 2.23714
R2470 DVDD.n638 DVDD.n635 2.23714
R2471 DVDD.n5469 DVDD.n630 2.23714
R2472 DVDD.n638 DVDD.n634 2.23714
R2473 DVDD.n5469 DVDD.n629 2.23714
R2474 DVDD.n1709 DVDD.n1698 2.23714
R2475 DVDD.n2048 DVDD.n1600 2.23714
R2476 DVDD.n1709 DVDD.n1699 2.23714
R2477 DVDD.n2048 DVDD.n1601 2.23714
R2478 DVDD.n2048 DVDD.n1595 2.23714
R2479 DVDD.n1709 DVDD.n1702 2.23714
R2480 DVDD.n2048 DVDD.n1602 2.23714
R2481 DVDD.n1709 DVDD.n1703 2.23714
R2482 DVDD.n2048 DVDD.n1603 2.23714
R2483 DVDD.n1709 DVDD.n1704 2.23714
R2484 DVDD.n2048 DVDD.n1604 2.23714
R2485 DVDD.n1709 DVDD.n1705 2.23714
R2486 DVDD.n2048 DVDD.n1605 2.23714
R2487 DVDD.n1709 DVDD.n1706 2.23714
R2488 DVDD.n1709 DVDD.n1707 2.23714
R2489 DVDD.n2048 DVDD.n1607 2.23714
R2490 DVDD.n1710 DVDD.n1709 2.23714
R2491 DVDD.n1709 DVDD.n1708 2.23714
R2492 DVDD.n2078 DVDD.n361 2.23714
R2493 DVDD.n5646 DVDD.n369 2.23714
R2494 DVDD.n2078 DVDD.n2068 2.23714
R2495 DVDD.n2078 DVDD.n2069 2.23714
R2496 DVDD.n5646 DVDD.n371 2.23714
R2497 DVDD.n2078 DVDD.n2070 2.23714
R2498 DVDD.n2078 DVDD.n2071 2.23714
R2499 DVDD.n5646 DVDD.n373 2.23714
R2500 DVDD.n2078 DVDD.n2072 2.23714
R2501 DVDD.n2078 DVDD.n2073 2.23714
R2502 DVDD.n5646 DVDD.n375 2.23714
R2503 DVDD.n2078 DVDD.n2074 2.23714
R2504 DVDD.n2078 DVDD.n2075 2.23714
R2505 DVDD.n5646 DVDD.n377 2.23714
R2506 DVDD.n2078 DVDD.n2076 2.23714
R2507 DVDD.n2078 DVDD.n2077 2.23714
R2508 DVDD.n5646 DVDD.n379 2.23714
R2509 DVDD.n2078 DVDD.n380 2.23714
R2510 DVDD.n5639 DVDD.n382 2.23714
R2511 DVDD.n5639 DVDD.n402 2.23714
R2512 DVDD.n5642 DVDD.n390 2.23714
R2513 DVDD.n5639 DVDD.n403 2.23714
R2514 DVDD.n5642 DVDD.n391 2.23714
R2515 DVDD.n5639 DVDD.n404 2.23714
R2516 DVDD.n5642 DVDD.n392 2.23714
R2517 DVDD.n5639 DVDD.n405 2.23714
R2518 DVDD.n5642 DVDD.n393 2.23714
R2519 DVDD.n5639 DVDD.n406 2.23714
R2520 DVDD.n5642 DVDD.n394 2.23714
R2521 DVDD.n5639 DVDD.n407 2.23714
R2522 DVDD.n5639 DVDD.n408 2.23714
R2523 DVDD.n5642 DVDD.n396 2.23714
R2524 DVDD.n5639 DVDD.n409 2.23714
R2525 DVDD.n5639 DVDD.n410 2.23714
R2526 DVDD.n5642 DVDD.n398 2.23714
R2527 DVDD.n5640 DVDD.n5639 2.23714
R2528 DVDD.n5642 DVDD.n384 2.23714
R2529 DVDD.n5633 DVDD.n412 2.23714
R2530 DVDD.n5635 DVDD.n421 2.23714
R2531 DVDD.n5633 DVDD.n437 2.23714
R2532 DVDD.n5633 DVDD.n438 2.23714
R2533 DVDD.n5635 DVDD.n423 2.23714
R2534 DVDD.n5633 DVDD.n434 2.23714
R2535 DVDD.n5635 DVDD.n418 2.23714
R2536 DVDD.n5633 DVDD.n433 2.23714
R2537 DVDD.n5635 DVDD.n416 2.23714
R2538 DVDD.n5633 DVDD.n440 2.23714
R2539 DVDD.n5635 DVDD.n425 2.23714
R2540 DVDD.n5635 DVDD.n415 2.23714
R2541 DVDD.n5633 DVDD.n442 2.23714
R2542 DVDD.n5635 DVDD.n426 2.23714
R2543 DVDD.n5635 DVDD.n414 2.23714
R2544 DVDD.n5633 DVDD.n5632 2.23714
R2545 DVDD.n5635 DVDD.n427 2.23714
R2546 DVDD.n2751 DVDD.n2748 2.23714
R2547 DVDD.n2754 DVDD.n2612 2.23714
R2548 DVDD.n2751 DVDD.n2749 2.23714
R2549 DVDD.n2751 DVDD.n2606 2.23714
R2550 DVDD.n2754 DVDD.n2613 2.23714
R2551 DVDD.n2751 DVDD.n2750 2.23714
R2552 DVDD.n2752 DVDD.n2751 2.23714
R2553 DVDD.n2754 DVDD.n2753 2.23714
R2554 DVDD.n3037 DVDD.n744 2.23714
R2555 DVDD.n3040 DVDD.n747 2.23714
R2556 DVDD.n3037 DVDD.n3028 2.23714
R2557 DVDD.n3040 DVDD.n748 2.23714
R2558 DVDD.n3037 DVDD.n3029 2.23714
R2559 DVDD.n3040 DVDD.n749 2.23714
R2560 DVDD.n3037 DVDD.n3030 2.23714
R2561 DVDD.n3040 DVDD.n750 2.23714
R2562 DVDD.n3037 DVDD.n3031 2.23714
R2563 DVDD.n3040 DVDD.n751 2.23714
R2564 DVDD.n3037 DVDD.n3032 2.23714
R2565 DVDD.n3040 DVDD.n752 2.23714
R2566 DVDD.n3037 DVDD.n3033 2.23714
R2567 DVDD.n3040 DVDD.n753 2.23714
R2568 DVDD.n3037 DVDD.n3034 2.23714
R2569 DVDD.n3040 DVDD.n754 2.23714
R2570 DVDD.n3037 DVDD.n3035 2.23714
R2571 DVDD.n3040 DVDD.n755 2.23714
R2572 DVDD.n3037 DVDD.n3036 2.23714
R2573 DVDD.n3040 DVDD.n756 2.23714
R2574 DVDD.n3038 DVDD.n3037 2.23714
R2575 DVDD.n3040 DVDD.n3039 2.23714
R2576 DVDD.n3037 DVDD.n757 2.23714
R2577 DVDD.n273 DVDD.n262 2.23714
R2578 DVDD.n5703 DVDD.n268 2.23714
R2579 DVDD.n273 DVDD.n272 2.23714
R2580 DVDD.n5703 DVDD.n267 2.23714
R2581 DVDD.n273 DVDD.n271 2.23714
R2582 DVDD.n5703 DVDD.n266 2.23714
R2583 DVDD.n273 DVDD.n270 2.23714
R2584 DVDD.n5703 DVDD.n265 2.23714
R2585 DVDD.n273 DVDD.n269 2.23714
R2586 DVDD.n5703 DVDD.n264 2.23714
R2587 DVDD.n2034 DVDD.n2025 2.23714
R2588 DVDD.n2037 DVDD.n1724 2.23714
R2589 DVDD.n2034 DVDD.n2026 2.23714
R2590 DVDD.n2037 DVDD.n1725 2.23714
R2591 DVDD.n2037 DVDD.n1719 2.23714
R2592 DVDD.n2034 DVDD.n2029 2.23714
R2593 DVDD.n2037 DVDD.n1726 2.23714
R2594 DVDD.n2034 DVDD.n2030 2.23714
R2595 DVDD.n2037 DVDD.n1727 2.23714
R2596 DVDD.n2034 DVDD.n2031 2.23714
R2597 DVDD.n2037 DVDD.n1728 2.23714
R2598 DVDD.n2034 DVDD.n2032 2.23714
R2599 DVDD.n2037 DVDD.n1729 2.23714
R2600 DVDD.n2034 DVDD.n2033 2.23714
R2601 DVDD.n2035 DVDD.n2034 2.23714
R2602 DVDD.n2037 DVDD.n2036 2.23714
R2603 DVDD.n2034 DVDD.n1743 2.23714
R2604 DVDD.n2034 DVDD.n1716 2.23714
R2605 DVDD.n1446 DVDD.n900 2.23714
R2606 DVDD.n2963 DVDD.n908 2.23714
R2607 DVDD.n1446 DVDD.n1436 2.23714
R2608 DVDD.n1446 DVDD.n1437 2.23714
R2609 DVDD.n2963 DVDD.n910 2.23714
R2610 DVDD.n1446 DVDD.n1438 2.23714
R2611 DVDD.n1446 DVDD.n1439 2.23714
R2612 DVDD.n2963 DVDD.n912 2.23714
R2613 DVDD.n1446 DVDD.n1440 2.23714
R2614 DVDD.n1446 DVDD.n1441 2.23714
R2615 DVDD.n2963 DVDD.n914 2.23714
R2616 DVDD.n1446 DVDD.n1442 2.23714
R2617 DVDD.n1446 DVDD.n1443 2.23714
R2618 DVDD.n2963 DVDD.n916 2.23714
R2619 DVDD.n1446 DVDD.n1444 2.23714
R2620 DVDD.n1446 DVDD.n1445 2.23714
R2621 DVDD.n2963 DVDD.n918 2.23714
R2622 DVDD.n1446 DVDD.n919 2.23714
R2623 DVDD.n2956 DVDD.n921 2.23714
R2624 DVDD.n2956 DVDD.n941 2.23714
R2625 DVDD.n2959 DVDD.n929 2.23714
R2626 DVDD.n2956 DVDD.n942 2.23714
R2627 DVDD.n2959 DVDD.n930 2.23714
R2628 DVDD.n2956 DVDD.n943 2.23714
R2629 DVDD.n2959 DVDD.n931 2.23714
R2630 DVDD.n2956 DVDD.n944 2.23714
R2631 DVDD.n2959 DVDD.n932 2.23714
R2632 DVDD.n2956 DVDD.n945 2.23714
R2633 DVDD.n2959 DVDD.n933 2.23714
R2634 DVDD.n2956 DVDD.n946 2.23714
R2635 DVDD.n2956 DVDD.n947 2.23714
R2636 DVDD.n2959 DVDD.n935 2.23714
R2637 DVDD.n2956 DVDD.n948 2.23714
R2638 DVDD.n2956 DVDD.n949 2.23714
R2639 DVDD.n2959 DVDD.n937 2.23714
R2640 DVDD.n2957 DVDD.n2956 2.23714
R2641 DVDD.n2959 DVDD.n923 2.23714
R2642 DVDD.n2949 DVDD.n951 2.23714
R2643 DVDD.n2952 DVDD.n960 2.23714
R2644 DVDD.n2949 DVDD.n973 2.23714
R2645 DVDD.n2949 DVDD.n974 2.23714
R2646 DVDD.n2952 DVDD.n962 2.23714
R2647 DVDD.n2949 DVDD.n970 2.23714
R2648 DVDD.n2952 DVDD.n957 2.23714
R2649 DVDD.n2949 DVDD.n969 2.23714
R2650 DVDD.n2952 DVDD.n955 2.23714
R2651 DVDD.n2949 DVDD.n976 2.23714
R2652 DVDD.n2952 DVDD.n964 2.23714
R2653 DVDD.n2952 DVDD.n954 2.23714
R2654 DVDD.n2949 DVDD.n2947 2.23714
R2655 DVDD.n2952 DVDD.n965 2.23714
R2656 DVDD.n2952 DVDD.n953 2.23714
R2657 DVDD.n2950 DVDD.n2949 2.23714
R2658 DVDD.n2952 DVDD.n2951 2.23714
R2659 DVDD.n5612 DVDD.n477 2.23714
R2660 DVDD.n5615 DVDD.n482 2.23714
R2661 DVDD.n5612 DVDD.n5610 2.23714
R2662 DVDD.n5612 DVDD.n5609 2.23714
R2663 DVDD.n5615 DVDD.n484 2.23714
R2664 DVDD.n5612 DVDD.n5611 2.23714
R2665 DVDD.n5613 DVDD.n5612 2.23714
R2666 DVDD.n5615 DVDD.n5614 2.23714
R2667 DVDD.n3746 DVDD.n3699 2.23714
R2668 DVDD.n3747 DVDD.n3745 2.23714
R2669 DVDD.n3748 DVDD.n3699 2.23714
R2670 DVDD.n3749 DVDD.n3745 2.23714
R2671 DVDD.n3750 DVDD.n3699 2.23714
R2672 DVDD.n3751 DVDD.n3745 2.23714
R2673 DVDD.n3752 DVDD.n3699 2.23714
R2674 DVDD.n3753 DVDD.n3745 2.23714
R2675 DVDD.n3754 DVDD.n3699 2.23714
R2676 DVDD.n3755 DVDD.n3745 2.23714
R2677 DVDD.n784 DVDD.n241 2.23714
R2678 DVDD.n5713 DVDD.n244 2.23714
R2679 DVDD.n784 DVDD.n774 2.23714
R2680 DVDD.n5713 DVDD.n245 2.23714
R2681 DVDD.n784 DVDD.n775 2.23714
R2682 DVDD.n5713 DVDD.n246 2.23714
R2683 DVDD.n784 DVDD.n776 2.23714
R2684 DVDD.n5713 DVDD.n247 2.23714
R2685 DVDD.n784 DVDD.n777 2.23714
R2686 DVDD.n5713 DVDD.n248 2.23714
R2687 DVDD.n784 DVDD.n778 2.23714
R2688 DVDD.n5713 DVDD.n249 2.23714
R2689 DVDD.n784 DVDD.n779 2.23714
R2690 DVDD.n5713 DVDD.n250 2.23714
R2691 DVDD.n784 DVDD.n780 2.23714
R2692 DVDD.n5713 DVDD.n251 2.23714
R2693 DVDD.n784 DVDD.n781 2.23714
R2694 DVDD.n5713 DVDD.n252 2.23714
R2695 DVDD.n784 DVDD.n782 2.23714
R2696 DVDD.n5713 DVDD.n253 2.23714
R2697 DVDD.n784 DVDD.n783 2.23714
R2698 DVDD.n5713 DVDD.n254 2.23714
R2699 DVDD.n784 DVDD.n255 2.23714
R2700 DVDD.n2972 DVDD.n838 2.23714
R2701 DVDD.n2974 DVDD.n833 2.23714
R2702 DVDD.n2972 DVDD.n837 2.23714
R2703 DVDD.n2974 DVDD.n832 2.23714
R2704 DVDD.n2972 DVDD.n836 2.23714
R2705 DVDD.n2974 DVDD.n831 2.23714
R2706 DVDD.n2972 DVDD.n835 2.23714
R2707 DVDD.n2974 DVDD.n830 2.23714
R2708 DVDD.n2972 DVDD.n834 2.23714
R2709 DVDD.n2974 DVDD.n829 2.23714
R2710 DVDD.n1798 DVDD.n881 2.23714
R2711 DVDD.n2969 DVDD.n888 2.23714
R2712 DVDD.n1798 DVDD.n1788 2.23714
R2713 DVDD.n2969 DVDD.n889 2.23714
R2714 DVDD.n2969 DVDD.n885 2.23714
R2715 DVDD.n1798 DVDD.n1791 2.23714
R2716 DVDD.n2969 DVDD.n890 2.23714
R2717 DVDD.n1798 DVDD.n1792 2.23714
R2718 DVDD.n2969 DVDD.n891 2.23714
R2719 DVDD.n1798 DVDD.n1793 2.23714
R2720 DVDD.n2969 DVDD.n892 2.23714
R2721 DVDD.n1798 DVDD.n1794 2.23714
R2722 DVDD.n2969 DVDD.n893 2.23714
R2723 DVDD.n1798 DVDD.n1795 2.23714
R2724 DVDD.n1798 DVDD.n1796 2.23714
R2725 DVDD.n2969 DVDD.n895 2.23714
R2726 DVDD.n1798 DVDD.n1797 2.23714
R2727 DVDD.n1798 DVDD.n897 2.23714
R2728 DVDD.n2216 DVDD.n2206 2.23714
R2729 DVDD.n2220 DVDD.n1399 2.23714
R2730 DVDD.n2216 DVDD.n2207 2.23714
R2731 DVDD.n2216 DVDD.n2208 2.23714
R2732 DVDD.n2220 DVDD.n1401 2.23714
R2733 DVDD.n2216 DVDD.n2209 2.23714
R2734 DVDD.n2216 DVDD.n2210 2.23714
R2735 DVDD.n2220 DVDD.n1403 2.23714
R2736 DVDD.n2216 DVDD.n2211 2.23714
R2737 DVDD.n2216 DVDD.n2212 2.23714
R2738 DVDD.n2220 DVDD.n1405 2.23714
R2739 DVDD.n2216 DVDD.n2213 2.23714
R2740 DVDD.n2216 DVDD.n2214 2.23714
R2741 DVDD.n2220 DVDD.n1407 2.23714
R2742 DVDD.n2216 DVDD.n2215 2.23714
R2743 DVDD.n2216 DVDD.n1392 2.23714
R2744 DVDD.n2220 DVDD.n1408 2.23714
R2745 DVDD.n2217 DVDD.n2216 2.23714
R2746 DVDD.n2438 DVDD.n2426 2.23714
R2747 DVDD.n2438 DVDD.n2427 2.23714
R2748 DVDD.n2441 DVDD.n1130 2.23714
R2749 DVDD.n2438 DVDD.n2428 2.23714
R2750 DVDD.n2441 DVDD.n1131 2.23714
R2751 DVDD.n2438 DVDD.n2429 2.23714
R2752 DVDD.n2441 DVDD.n1132 2.23714
R2753 DVDD.n2438 DVDD.n2430 2.23714
R2754 DVDD.n2441 DVDD.n1133 2.23714
R2755 DVDD.n2438 DVDD.n2431 2.23714
R2756 DVDD.n2441 DVDD.n1134 2.23714
R2757 DVDD.n2438 DVDD.n2432 2.23714
R2758 DVDD.n2438 DVDD.n2433 2.23714
R2759 DVDD.n2441 DVDD.n1136 2.23714
R2760 DVDD.n2438 DVDD.n2434 2.23714
R2761 DVDD.n2438 DVDD.n1122 2.23714
R2762 DVDD.n2441 DVDD.n1137 2.23714
R2763 DVDD.n2439 DVDD.n2438 2.23714
R2764 DVDD.n2441 DVDD.n1124 2.23714
R2765 DVDD.n5622 DVDD.n455 2.23714
R2766 DVDD.n472 DVDD.n467 2.23714
R2767 DVDD.n5622 DVDD.n456 2.23714
R2768 DVDD.n5622 DVDD.n457 2.23714
R2769 DVDD.n472 DVDD.n468 2.23714
R2770 DVDD.n5622 DVDD.n452 2.23714
R2771 DVDD.n472 DVDD.n466 2.23714
R2772 DVDD.n5622 DVDD.n451 2.23714
R2773 DVDD.n472 DVDD.n465 2.23714
R2774 DVDD.n5622 DVDD.n459 2.23714
R2775 DVDD.n472 DVDD.n469 2.23714
R2776 DVDD.n472 DVDD.n464 2.23714
R2777 DVDD.n5622 DVDD.n461 2.23714
R2778 DVDD.n472 DVDD.n470 2.23714
R2779 DVDD.n472 DVDD.n447 2.23714
R2780 DVDD.n5622 DVDD.n462 2.23714
R2781 DVDD.n472 DVDD.n471 2.23714
R2782 DVDD.n2911 DVDD.n2908 2.23714
R2783 DVDD.n2914 DVDD.n2593 2.23714
R2784 DVDD.n2911 DVDD.n2909 2.23714
R2785 DVDD.n2911 DVDD.n2907 2.23714
R2786 DVDD.n2914 DVDD.n2765 2.23714
R2787 DVDD.n2911 DVDD.n2910 2.23714
R2788 DVDD.n2911 DVDD.n2588 2.23714
R2789 DVDD.n2914 DVDD.n2913 2.23714
R2790 DVDD.n4325 DVDD.n3506 2.23714
R2791 DVDD.n4322 DVDD.n4214 2.23714
R2792 DVDD.n4325 DVDD.n3507 2.23714
R2793 DVDD.n4322 DVDD.n4213 2.23714
R2794 DVDD.n4325 DVDD.n4209 2.23714
R2795 DVDD.n4323 DVDD.n4322 2.23714
R2796 DVDD.n4325 DVDD.n4324 2.23714
R2797 DVDD.n4322 DVDD.n4210 2.23714
R2798 DVDD.n3511 DVDD.n3374 2.23714
R2799 DVDD.n3512 DVDD.n3373 2.23714
R2800 DVDD.n3513 DVDD.n3374 2.23714
R2801 DVDD.n3514 DVDD.n3373 2.23714
R2802 DVDD.n3515 DVDD.n3374 2.23714
R2803 DVDD.n4686 DVDD.n3373 2.23714
R2804 DVDD.n4687 DVDD.n3374 2.23714
R2805 DVDD.n4688 DVDD.n3373 2.23714
R2806 DVDD.n4689 DVDD.n3374 2.23714
R2807 DVDD.n4187 DVDD.n3426 2.23714
R2808 DVDD.n4188 DVDD.n3427 2.23714
R2809 DVDD.n4189 DVDD.n3426 2.23714
R2810 DVDD.n4190 DVDD.n3427 2.23714
R2811 DVDD.n4191 DVDD.n3426 2.23714
R2812 DVDD.n4542 DVDD.n3427 2.23714
R2813 DVDD.n4541 DVDD.n3426 2.23714
R2814 DVDD.n4540 DVDD.n3427 2.23714
R2815 DVDD.n4539 DVDD.n3426 2.23714
R2816 DVDD.n5987 DVDD.n18 2.23714
R2817 DVDD.n19 DVDD.n11 2.23714
R2818 DVDD.n5987 DVDD.n20 2.23714
R2819 DVDD.n21 DVDD.n11 2.23714
R2820 DVDD.n5985 DVDD.n11 2.23714
R2821 DVDD.n5987 DVDD.n23 2.23714
R2822 DVDD.n24 DVDD.n11 2.23714
R2823 DVDD.n5987 DVDD.n25 2.23714
R2824 DVDD.n4120 DVDD.n4119 2.21947
R2825 DVDD.n5547 DVDD.n542 2.21947
R2826 DVDD.n5548 DVDD.n541 2.21947
R2827 DVDD.n5549 DVDD.n540 2.21947
R2828 DVDD.n5550 DVDD.n539 2.21947
R2829 DVDD.n5551 DVDD.n538 2.21947
R2830 DVDD.n5552 DVDD.n537 2.21947
R2831 DVDD.n5553 DVDD.n536 2.21947
R2832 DVDD.n5554 DVDD.n535 2.21947
R2833 DVDD.n5555 DVDD.n534 2.21947
R2834 DVDD.n5556 DVDD.n533 2.21947
R2835 DVDD.n5557 DVDD.n532 2.21947
R2836 DVDD.n5558 DVDD.n531 2.21947
R2837 DVDD.n5559 DVDD.n530 2.21947
R2838 DVDD.n5560 DVDD.n529 2.21947
R2839 DVDD.n5561 DVDD.n528 2.21947
R2840 DVDD.n5563 DVDD.n5562 2.21947
R2841 DVDD.n2921 DVDD.n2584 2.21947
R2842 DVDD.n2757 DVDD.n2756 2.21947
R2843 DVDD.n2610 DVDD.n2573 2.21947
R2844 DVDD.n1007 DVDD.n429 2.21947
R2845 DVDD.n1011 DVDD.n428 2.21947
R2846 DVDD.n5630 DVDD.n5629 2.21947
R2847 DVDD.n2939 DVDD.n2938 2.21947
R2848 DVDD.n2556 DVDD.n2555 2.21947
R2849 DVDD.n2538 DVDD.n2537 2.21947
R2850 DVDD.n2523 DVDD.n2522 2.21947
R2851 DVDD.n5637 DVDD.n411 2.21947
R2852 DVDD.n1261 DVDD.n399 2.21947
R2853 DVDD.n2448 DVDD.n1118 2.21947
R2854 DVDD.n1249 DVDD.n1248 2.21947
R2855 DVDD.n1231 DVDD.n1230 2.21947
R2856 DVDD.n5644 DVDD.n381 2.21947
R2857 DVDD.n2227 DVDD.n1388 2.21947
R2858 DVDD.n1533 DVDD.n1532 2.21947
R2859 DVDD.n1519 DVDD.n1518 2.21947
R2860 DVDD.n1505 DVDD.n1504 2.21947
R2861 DVDD.n1491 DVDD.n1490 2.21947
R2862 DVDD.n5649 DVDD.n5648 2.21947
R2863 DVDD.n2046 DVDD.n2045 2.21947
R2864 DVDD.n1735 DVDD.n1734 2.21947
R2865 DVDD.n5522 DVDD.n5519 2.21947
R2866 DVDD.n2845 DVDD.n555 2.21947
R2867 DVDD.n2829 DVDD.n2828 2.21947
R2868 DVDD.n2826 DVDD.n2823 2.21947
R2869 DVDD.n2822 DVDD.n2819 2.21947
R2870 DVDD.n2818 DVDD.n2815 2.21947
R2871 DVDD.n2814 DVDD.n2811 2.21947
R2872 DVDD.n2810 DVDD.n2807 2.21947
R2873 DVDD.n2806 DVDD.n2803 2.21947
R2874 DVDD.n2802 DVDD.n2799 2.21947
R2875 DVDD.n2798 DVDD.n2795 2.21947
R2876 DVDD.n2794 DVDD.n2791 2.21947
R2877 DVDD.n2790 DVDD.n2787 2.21947
R2878 DVDD.n2786 DVDD.n2783 2.21947
R2879 DVDD.n2769 DVDD.n524 2.21947
R2880 DVDD.n5566 DVDD.n525 2.21947
R2881 DVDD.n2918 DVDD.n2585 2.21947
R2882 DVDD.n2760 DVDD.n2759 2.21947
R2883 DVDD.n2570 DVDD.n2569 2.21947
R2884 DVDD.n2568 DVDD.n474 2.21947
R2885 DVDD.n1014 DVDD.n1010 2.21947
R2886 DVDD.n5626 DVDD.n444 2.21947
R2887 DVDD.n2942 DVDD.n2941 2.21947
R2888 DVDD.n2559 DVDD.n2552 2.21947
R2889 DVDD.n2541 DVDD.n2534 2.21947
R2890 DVDD.n2526 DVDD.n2518 2.21947
R2891 DVDD.n1210 DVDD.n1207 2.21947
R2892 DVDD.n1264 DVDD.n1258 2.21947
R2893 DVDD.n2445 DVDD.n1119 2.21947
R2894 DVDD.n1252 DVDD.n1244 2.21947
R2895 DVDD.n1234 DVDD.n1226 2.21947
R2896 DVDD.n1552 DVDD.n1549 2.21947
R2897 DVDD.n2224 DVDD.n1389 2.21947
R2898 DVDD.n1536 DVDD.n1528 2.21947
R2899 DVDD.n1522 DVDD.n1514 2.21947
R2900 DVDD.n1508 DVDD.n1500 2.21947
R2901 DVDD.n1494 DVDD.n1486 2.21947
R2902 DVDD.n5652 DVDD.n358 2.21947
R2903 DVDD.n2042 DVDD.n1714 2.21947
R2904 DVDD.n1738 DVDD.n1737 2.21947
R2905 DVDD.n5518 DVDD.n556 2.21947
R2906 DVDD.n2847 DVDD.n2846 2.21947
R2907 DVDD.n2848 DVDD.n2842 2.21947
R2908 DVDD.n2849 DVDD.n2781 2.21947
R2909 DVDD.n2850 DVDD.n2780 2.21947
R2910 DVDD.n2851 DVDD.n2779 2.21947
R2911 DVDD.n2852 DVDD.n2778 2.21947
R2912 DVDD.n2853 DVDD.n2777 2.21947
R2913 DVDD.n2854 DVDD.n2776 2.21947
R2914 DVDD.n2855 DVDD.n2775 2.21947
R2915 DVDD.n2856 DVDD.n2774 2.21947
R2916 DVDD.n2857 DVDD.n2773 2.21947
R2917 DVDD.n2858 DVDD.n2772 2.21947
R2918 DVDD.n2859 DVDD.n2771 2.21947
R2919 DVDD.n2860 DVDD.n2770 2.21947
R2920 DVDD.n2862 DVDD.n2861 2.21947
R2921 DVDD.n2917 DVDD.n2586 2.21947
R2922 DVDD.n2762 DVDD.n2761 2.21947
R2923 DVDD.n5617 DVDD.n476 2.21947
R2924 DVDD.n5619 DVDD.n5618 2.21947
R2925 DVDD.n1009 DVDD.n1008 2.21947
R2926 DVDD.n5625 DVDD.n445 2.21947
R2927 DVDD.n2945 DVDD.n2944 2.21947
R2928 DVDD.n2551 DVDD.n2548 2.21947
R2929 DVDD.n2533 DVDD.n2530 2.21947
R2930 DVDD.n2517 DVDD.n2513 2.21947
R2931 DVDD.n2954 DVDD.n950 2.21947
R2932 DVDD.n1257 DVDD.n938 2.21947
R2933 DVDD.n2444 DVDD.n1120 2.21947
R2934 DVDD.n1243 DVDD.n1241 2.21947
R2935 DVDD.n1225 DVDD.n1223 2.21947
R2936 DVDD.n2961 DVDD.n920 2.21947
R2937 DVDD.n2223 DVDD.n1390 2.21947
R2938 DVDD.n1527 DVDD.n1525 2.21947
R2939 DVDD.n1513 DVDD.n1511 2.21947
R2940 DVDD.n1499 DVDD.n1497 2.21947
R2941 DVDD.n1485 DVDD.n1483 2.21947
R2942 DVDD.n2966 DVDD.n2965 2.21947
R2943 DVDD.n2041 DVDD.n2039 2.21947
R2944 DVDD.n1741 DVDD.n1740 2.21947
R2945 DVDD.n3760 DVDD.n3759 2.21947
R2946 DVDD.n3908 DVDD.n3907 2.14722
R2947 DVDD.n3910 DVDD.n3909 2.14722
R2948 DVDD.n3678 DVDD.n3526 2.14722
R2949 DVDD.n4198 DVDD.n4197 2.14722
R2950 DVDD.n5832 DVDD.n5831 2.14713
R2951 DVDD.n3914 DVDD.n3668 2.14672
R2952 DVDD.n3913 DVDD.n3912 2.14672
R2953 DVDD.n3676 DVDD.n3519 2.14672
R2954 DVDD.n4201 DVDD.n4200 2.14672
R2955 DVDD.n5877 DVDD.n166 1.99748
R2956 DVDD.n5877 DVDD.n165 1.99748
R2957 DVDD.n5877 DVDD.n164 1.99748
R2958 DVDD.n5877 DVDD.n163 1.99748
R2959 DVDD.n5877 DVDD.n162 1.99748
R2960 DVDD.n5877 DVDD.n161 1.99748
R2961 DVDD.n5877 DVDD.n160 1.99748
R2962 DVDD.n5877 DVDD.n159 1.99748
R2963 DVDD.n5877 DVDD.n158 1.99748
R2964 DVDD.n5877 DVDD.n157 1.99748
R2965 DVDD.n5877 DVDD.n156 1.99748
R2966 DVDD.n5877 DVDD.n155 1.99748
R2967 DVDD.n5877 DVDD.n154 1.99748
R2968 DVDD.n5877 DVDD.n153 1.99748
R2969 DVDD.n5877 DVDD.n152 1.99748
R2970 DVDD.n5877 DVDD.n151 1.99748
R2971 DVDD.n5877 DVDD.n150 1.99748
R2972 DVDD.n5877 DVDD.n149 1.99748
R2973 DVDD.n5877 DVDD.n148 1.99748
R2974 DVDD.n5877 DVDD.n147 1.99748
R2975 DVDD.n5877 DVDD.n146 1.99748
R2976 DVDD.n5877 DVDD.n145 1.99748
R2977 DVDD.n5877 DVDD.n144 1.99748
R2978 DVDD.n5877 DVDD.n143 1.99748
R2979 DVDD.n5877 DVDD.n142 1.99748
R2980 DVDD.n5877 DVDD.n141 1.99748
R2981 DVDD.n5877 DVDD.n140 1.99748
R2982 DVDD.n5877 DVDD.n139 1.99748
R2983 DVDD.n5877 DVDD.n138 1.99748
R2984 DVDD.n5877 DVDD.n137 1.99748
R2985 DVDD.n5877 DVDD.n136 1.99748
R2986 DVDD.n5877 DVDD.n135 1.99748
R2987 DVDD.n5877 DVDD.n134 1.99748
R2988 DVDD.n5877 DVDD.n133 1.99748
R2989 DVDD.n5877 DVDD.n132 1.99748
R2990 DVDD.n5877 DVDD.n131 1.99748
R2991 DVDD.n5877 DVDD.n130 1.99748
R2992 DVDD.n5877 DVDD.n129 1.99748
R2993 DVDD.n5877 DVDD.n128 1.99748
R2994 DVDD.n5877 DVDD.n127 1.99748
R2995 DVDD.n5877 DVDD.n126 1.99748
R2996 DVDD.n5877 DVDD.n125 1.99748
R2997 DVDD.n5877 DVDD.n124 1.99748
R2998 DVDD.n5877 DVDD.n123 1.99748
R2999 DVDD.n5877 DVDD.n122 1.99748
R3000 DVDD.n5877 DVDD.n121 1.99748
R3001 DVDD.n5877 DVDD.n120 1.99748
R3002 DVDD.n5877 DVDD.n119 1.99748
R3003 DVDD.n5877 DVDD.n118 1.99748
R3004 DVDD.n5877 DVDD.n117 1.99748
R3005 DVDD.n5877 DVDD.n116 1.99748
R3006 DVDD.n5877 DVDD.n115 1.99748
R3007 DVDD.n5877 DVDD.n114 1.99748
R3008 DVDD.n5877 DVDD.n113 1.99748
R3009 DVDD.n5877 DVDD.n112 1.99748
R3010 DVDD.n5877 DVDD.n111 1.99748
R3011 DVDD.n5877 DVDD.n110 1.99748
R3012 DVDD.n5877 DVDD.n109 1.99748
R3013 DVDD.n5877 DVDD.n108 1.99748
R3014 DVDD.n5877 DVDD.n107 1.99748
R3015 DVDD.n5877 DVDD.n106 1.99748
R3016 DVDD.n5878 DVDD.n5877 1.99748
R3017 DVDD.n5877 DVDD.n168 1.99748
R3018 DVDD.n5951 DVDD.n31 1.99748
R3019 DVDD.n5956 DVDD.n31 1.99748
R3020 DVDD.n40 DVDD.n31 1.99748
R3021 DVDD.n5963 DVDD.n31 1.99748
R3022 DVDD.n38 DVDD.n31 1.99748
R3023 DVDD.n5970 DVDD.n31 1.99748
R3024 DVDD.n35 DVDD.n31 1.99748
R3025 DVDD.n5977 DVDD.n31 1.99748
R3026 DVDD.n5980 DVDD.n31 1.99748
R3027 DVDD.n4560 DVDD.n31 1.99748
R3028 DVDD.n4565 DVDD.n31 1.99748
R3029 DVDD.n4559 DVDD.n31 1.99748
R3030 DVDD.n4572 DVDD.n31 1.99748
R3031 DVDD.n4556 DVDD.n31 1.99748
R3032 DVDD.n4579 DVDD.n31 1.99748
R3033 DVDD.n4553 DVDD.n31 1.99748
R3034 DVDD.n4586 DVDD.n31 1.99748
R3035 DVDD.n4550 DVDD.n31 1.99748
R3036 DVDD.n4593 DVDD.n31 1.99748
R3037 DVDD.n4547 DVDD.n31 1.99748
R3038 DVDD.n4600 DVDD.n31 1.99748
R3039 DVDD.n3422 DVDD.n31 1.99748
R3040 DVDD.n4607 DVDD.n31 1.99748
R3041 DVDD.n3419 DVDD.n31 1.99748
R3042 DVDD.n4614 DVDD.n31 1.99748
R3043 DVDD.n3416 DVDD.n31 1.99748
R3044 DVDD.n4621 DVDD.n31 1.99748
R3045 DVDD.n3413 DVDD.n31 1.99748
R3046 DVDD.n4628 DVDD.n31 1.99748
R3047 DVDD.n3410 DVDD.n31 1.99748
R3048 DVDD.n4635 DVDD.n31 1.99748
R3049 DVDD.n3407 DVDD.n31 1.99748
R3050 DVDD.n3404 DVDD.n31 1.99748
R3051 DVDD.n4644 DVDD.n31 1.99748
R3052 DVDD.n3394 DVDD.n31 1.99748
R3053 DVDD.n4651 DVDD.n31 1.99748
R3054 DVDD.n3391 DVDD.n31 1.99748
R3055 DVDD.n4658 DVDD.n31 1.99748
R3056 DVDD.n3388 DVDD.n31 1.99748
R3057 DVDD.n4665 DVDD.n31 1.99748
R3058 DVDD.n3385 DVDD.n31 1.99748
R3059 DVDD.n4672 DVDD.n31 1.99748
R3060 DVDD.n3382 DVDD.n31 1.99748
R3061 DVDD.n4679 DVDD.n31 1.99748
R3062 DVDD.n3379 DVDD.n31 1.99748
R3063 DVDD.n4280 DVDD.n31 1.99748
R3064 DVDD.n4276 DVDD.n31 1.99748
R3065 DVDD.n4287 DVDD.n31 1.99748
R3066 DVDD.n4273 DVDD.n31 1.99748
R3067 DVDD.n4294 DVDD.n31 1.99748
R3068 DVDD.n4270 DVDD.n31 1.99748
R3069 DVDD.n4301 DVDD.n31 1.99748
R3070 DVDD.n4267 DVDD.n31 1.99748
R3071 DVDD.n4308 DVDD.n31 1.99748
R3072 DVDD.n4264 DVDD.n31 1.99748
R3073 DVDD.n4315 DVDD.n31 1.99748
R3074 DVDD.n4260 DVDD.n31 1.99748
R3075 DVDD.n4218 DVDD.n31 1.99748
R3076 DVDD.n4253 DVDD.n31 1.99748
R3077 DVDD.n4247 DVDD.n31 1.99748
R3078 DVDD.n4245 DVDD.n31 1.99748
R3079 DVDD.n4239 DVDD.n31 1.99748
R3080 DVDD.n4237 DVDD.n31 1.99748
R3081 DVDD.n4231 DVDD.n31 1.99748
R3082 DVDD.n4229 DVDD.n31 1.99748
R3083 DVDD.n5926 DVDD.t71 1.74266
R3084 DVDD.n5901 DVDD.t8 1.74266
R3085 DVDD.n3758 DVDD.t155 1.70818
R3086 DVDD.n3937 DVDD.t157 1.70818
R3087 DVDD.n4117 DVDD.t158 1.70818
R3088 DVDD.n3889 DVDD.t161 1.70818
R3089 DVDD.n5661 DVDD.n305 1.52209
R3090 DVDD.n4534 DVDD.n4496 1.52209
R3091 DVDD.n5313 DVDD.n4908 1.52209
R3092 DVDD.n5306 DVDD.n4916 1.52209
R3093 DVDD.n5474 DVDD.t20 1.52141
R3094 DVDD.n607 DVDD.t3 1.52141
R3095 DVDD.n5709 DVDD.t18 1.52141
R3096 DVDD.n5018 DVDD.n5012 1.52029
R3097 DVDD.n5754 DVDD.n180 1.52029
R3098 DVDD.n5288 DVDD.n4929 1.52029
R3099 DVDD.n4882 DVDD.n4881 1.52029
R3100 DVDD.n3761 DVDD.n3697 1.50887
R3101 DVDD.n4121 DVDD.n3549 1.50887
R3102 DVDD.n5660 DVDD.n5659 1.5005
R3103 DVDD.n5034 DVDD.n297 1.5005
R3104 DVDD.n5015 DVDD.n5011 1.5005
R3105 DVDD.n5029 DVDD.n5028 1.5005
R3106 DVDD.n5019 DVDD.n5013 1.5005
R3107 DVDD.n302 DVDD.n298 1.5005
R3108 DVDD.n5665 DVDD.n5664 1.5005
R3109 DVDD.n306 DVDD.n303 1.5005
R3110 DVDD.n5662 DVDD.n303 1.5005
R3111 DVDD.n5664 DVDD.n5663 1.5005
R3112 DVDD.n304 DVDD.n302 1.5005
R3113 DVDD.n5034 DVDD.n5033 1.5005
R3114 DVDD.n5031 DVDD.n5011 1.5005
R3115 DVDD.n5030 DVDD.n5029 1.5005
R3116 DVDD.n5312 DVDD.n5311 1.5005
R3117 DVDD.n5746 DVDD.n185 1.5005
R3118 DVDD.n4900 DVDD.n183 1.5005
R3119 DVDD.n5750 DVDD.n182 1.5005
R3120 DVDD.n5752 DVDD.n5751 1.5005
R3121 DVDD.n733 DVDD.n200 1.5005
R3122 DVDD.n5317 DVDD.n5316 1.5005
R3123 DVDD.n4909 DVDD.n4906 1.5005
R3124 DVDD.n5314 DVDD.n4906 1.5005
R3125 DVDD.n5316 DVDD.n5315 1.5005
R3126 DVDD.n4907 DVDD.n200 1.5005
R3127 DVDD.n5747 DVDD.n5746 1.5005
R3128 DVDD.n5748 DVDD.n183 1.5005
R3129 DVDD.n5750 DVDD.n5749 1.5005
R3130 DVDD.n4927 DVDD.n4925 1.5005
R3131 DVDD.n5299 DVDD.n5298 1.5005
R3132 DVDD.n5300 DVDD.n4919 1.5005
R3133 DVDD.n5303 DVDD.n4918 1.5005
R3134 DVDD.n5305 DVDD.n5304 1.5005
R3135 DVDD.n5292 DVDD.n5291 1.5005
R3136 DVDD.n4930 DVDD.n4928 1.5005
R3137 DVDD.n5287 DVDD.n5286 1.5005
R3138 DVDD.n5289 DVDD.n4928 1.5005
R3139 DVDD.n5291 DVDD.n5290 1.5005
R3140 DVDD.n4927 DVDD.n222 1.5005
R3141 DVDD.n5299 DVDD.n223 1.5005
R3142 DVDD.n5301 DVDD.n5300 1.5005
R3143 DVDD.n5303 DVDD.n5302 1.5005
R3144 DVDD.n4520 DVDD.n3170 1.5005
R3145 DVDD.n4500 DVDD.n3171 1.5005
R3146 DVDD.n4528 DVDD.n4527 1.5005
R3147 DVDD.n4531 DVDD.n4498 1.5005
R3148 DVDD.n4533 DVDD.n4532 1.5005
R3149 DVDD.n4521 DVDD.n3144 1.5005
R3150 DVDD.n4879 DVDD.n4878 1.5005
R3151 DVDD.n3146 DVDD.n3142 1.5005
R3152 DVDD.n4880 DVDD.n4879 1.5005
R3153 DVDD.n3144 DVDD.n3143 1.5005
R3154 DVDD.n3170 DVDD.n3157 1.5005
R3155 DVDD.n3171 DVDD.n3158 1.5005
R3156 DVDD.n4529 DVDD.n4528 1.5005
R3157 DVDD.n4531 DVDD.n4530 1.5005
R3158 DVDD.n4535 DVDD.n4534 1.5005
R3159 DVDD.n4497 DVDD.n4495 1.5005
R3160 DVDD.n4506 DVDD.n4505 1.5005
R3161 DVDD.n4501 DVDD.n4499 1.5005
R3162 DVDD.n4526 DVDD.n4525 1.5005
R3163 DVDD.n4523 DVDD.n4522 1.5005
R3164 DVDD.n3147 DVDD.n3145 1.5005
R3165 DVDD.n4877 DVDD.n4876 1.5005
R3166 DVDD.n3141 DVDD.n3140 1.5005
R3167 DVDD.n4883 DVDD.n4882 1.5005
R3168 DVDD.n5755 DVDD.n5754 1.5005
R3169 DVDD.n5753 DVDD.n179 1.5005
R3170 DVDD.n3132 DVDD.n181 1.5005
R3171 DVDD.n4899 DVDD.n3129 1.5005
R3172 DVDD.n4902 DVDD.n4901 1.5005
R3173 DVDD.n5319 DVDD.n5318 1.5005
R3174 DVDD.n4905 DVDD.n4904 1.5005
R3175 DVDD.n4911 DVDD.n4910 1.5005
R3176 DVDD.n5310 DVDD.n5309 1.5005
R3177 DVDD.n5308 DVDD.n4908 1.5005
R3178 DVDD.n5307 DVDD.n5306 1.5005
R3179 DVDD.n4917 DVDD.n4915 1.5005
R3180 DVDD.n5110 DVDD.n5109 1.5005
R3181 DVDD.n4921 DVDD.n4920 1.5005
R3182 DVDD.n5297 DVDD.n5296 1.5005
R3183 DVDD.n5294 DVDD.n5293 1.5005
R3184 DVDD.n4926 DVDD.n4924 1.5005
R3185 DVDD.n4932 DVDD.n4931 1.5005
R3186 DVDD.n5285 DVDD.n5284 1.5005
R3187 DVDD.n5283 DVDD.n4929 1.5005
R3188 DVDD.n5018 DVDD.n5017 1.5005
R3189 DVDD.n5021 DVDD.n5020 1.5005
R3190 DVDD.n5022 DVDD.n5014 1.5005
R3191 DVDD.n5027 DVDD.n5026 1.5005
R3192 DVDD.n5025 DVDD.n5024 1.5005
R3193 DVDD.n5669 DVDD.n5668 1.5005
R3194 DVDD.n5667 DVDD.n5666 1.5005
R3195 DVDD.n308 DVDD.n301 1.5005
R3196 DVDD.n309 DVDD.n307 1.5005
R3197 DVDD.n5658 DVDD.n5657 1.5005
R3198 DVDD.n5656 DVDD.n305 1.5005
R3199 DVDD.n5522 DVDD.n5521 1.44597
R3200 DVDD.n2844 DVDD.n555 1.44597
R3201 DVDD.n2828 DVDD.n2827 1.44597
R3202 DVDD.n2826 DVDD.n2825 1.44597
R3203 DVDD.n2822 DVDD.n2821 1.44597
R3204 DVDD.n2818 DVDD.n2817 1.44597
R3205 DVDD.n2814 DVDD.n2813 1.44597
R3206 DVDD.n2810 DVDD.n2809 1.44597
R3207 DVDD.n2806 DVDD.n2805 1.44597
R3208 DVDD.n2802 DVDD.n2801 1.44597
R3209 DVDD.n2798 DVDD.n2797 1.44597
R3210 DVDD.n2794 DVDD.n2793 1.44597
R3211 DVDD.n2790 DVDD.n2789 1.44597
R3212 DVDD.n2786 DVDD.n2785 1.44597
R3213 DVDD.n2768 DVDD.n524 1.44597
R3214 DVDD.n5566 DVDD.n5565 1.44597
R3215 DVDD.n2920 DVDD.n2585 1.44597
R3216 DVDD.n2759 DVDD.n2758 1.44597
R3217 DVDD.n2572 DVDD.n2569 1.44597
R3218 DVDD.n2568 DVDD.n2567 1.44597
R3219 DVDD.n1014 DVDD.n1013 1.44597
R3220 DVDD.n5628 DVDD.n444 1.44597
R3221 DVDD.n2941 DVDD.n2940 1.44597
R3222 DVDD.n2559 DVDD.n2558 1.44597
R3223 DVDD.n2541 DVDD.n2540 1.44597
R3224 DVDD.n2526 DVDD.n2525 1.44597
R3225 DVDD.n1210 DVDD.n1209 1.44597
R3226 DVDD.n1264 DVDD.n1263 1.44597
R3227 DVDD.n2447 DVDD.n1119 1.44597
R3228 DVDD.n1252 DVDD.n1251 1.44597
R3229 DVDD.n1234 DVDD.n1233 1.44597
R3230 DVDD.n1552 DVDD.n1551 1.44597
R3231 DVDD.n2226 DVDD.n1389 1.44597
R3232 DVDD.n1536 DVDD.n1535 1.44597
R3233 DVDD.n1522 DVDD.n1521 1.44597
R3234 DVDD.n1508 DVDD.n1507 1.44597
R3235 DVDD.n1494 DVDD.n1493 1.44597
R3236 DVDD.n5652 DVDD.n5651 1.44597
R3237 DVDD.n2044 DVDD.n1714 1.44597
R3238 DVDD.n1737 DVDD.n1736 1.44597
R3239 DVDD.n5545 DVDD.n5544 1.37387
R3240 DVDD.n5547 DVDD.n5546 1.37387
R3241 DVDD.n556 DVDD.n553 1.37387
R3242 DVDD.n5517 DVDD.n5516 1.37358
R3243 DVDD.n5917 DVDD.t72 1.16194
R3244 DVDD.n5910 DVDD.t52 1.16194
R3245 DVDD.n609 DVDD.n608 1.15801
R3246 DVDD.n611 DVDD.n610 1.15801
R3247 DVDD.n613 DVDD.n612 1.15801
R3248 DVDD.n615 DVDD.n614 1.15801
R3249 DVDD.n5477 DVDD.n618 1.15801
R3250 DVDD.n5476 DVDD.n619 1.15801
R3251 DVDD.n5475 DVDD.n620 1.15801
R3252 DVDD.n625 DVDD.n622 1.15801
R3253 DVDD.n624 DVDD.n623 1.15801
R3254 DVDD.n5708 DVDD.n257 1.15801
R3255 DVDD.n5707 DVDD.n258 1.15801
R3256 DVDD.n5283 DVDD.n5282 1.13457
R3257 DVDD.n4524 DVDD.n3169 1.1255
R3258 DVDD.n5321 DVDD.n5320 1.1255
R3259 DVDD.n5295 DVDD.n233 1.1255
R3260 DVDD.n5478 DVDD.n617 1.10828
R3261 DVDD.n5473 DVDD.n621 1.10828
R3262 DVDD.n260 DVDD.n259 1.10828
R3263 DVDD.n5479 DVDD.n616 0.9005
R3264 DVDD.n3185 DVDD.n3184 0.8825
R3265 DVDD.n4538 DVDD.n4537 0.8825
R3266 DVDD.n4691 DVDD.n4690 0.8825
R3267 DVDD.n3504 DVDD.n3503 0.8825
R3268 DVDD.n5496 DVDD.n5494 0.8798
R3269 DVDD.n1598 DVDD.n1597 0.8798
R3270 DVDD.n1722 DVDD.n1721 0.8798
R3271 DVDD.n2971 DVDD.n2970 0.8798
R3272 DVDD.n3759 DVDD.n3757 0.81533
R3273 DVDD.n4119 DVDD.n4118 0.81533
R3274 DVDD.n5030 DVDD.n5012 0.769684
R3275 DVDD.n5662 DVDD.n5661 0.769684
R3276 DVDD.n5749 DVDD.n180 0.769684
R3277 DVDD.n5314 DVDD.n5313 0.769684
R3278 DVDD.n5302 DVDD.n4916 0.769684
R3279 DVDD.n5289 DVDD.n5288 0.769684
R3280 DVDD.n4530 DVDD.n4496 0.769684
R3281 DVDD.n4881 DVDD.n4880 0.769684
R3282 DVDD.n731 DVDD.n194 0.7505
R3283 DVDD.n729 DVDD.n194 0.7505
R3284 DVDD.n5535 DVDD.n5534 0.6665
R3285 DVDD.n5557 DVDD.n5556 0.6665
R3286 DVDD.n2856 DVDD.n2855 0.6665
R3287 DVDD.n2834 DVDD.n2833 0.6665
R3288 DVDD DVDD.n3936 0.66035
R3289 DVDD DVDD.n3586 0.659428
R3290 DVDD.n2934 DVDD.n2933 0.65165
R3291 DVDD.n5634 DVDD.n429 0.65165
R3292 DVDD.n5618 DVDD.n475 0.65165
R3293 DVDD.n5621 DVDD.n5620 0.65165
R3294 DVDD DVDD.n3758 0.630979
R3295 DVDD.n3758 DVDD 0.630979
R3296 DVDD DVDD.n3937 0.630979
R3297 DVDD.n3937 DVDD 0.630979
R3298 DVDD.n4117 DVDD 0.630979
R3299 DVDD DVDD.n4117 0.630979
R3300 DVDD DVDD.n3889 0.630979
R3301 DVDD.n3889 DVDD 0.630979
R3302 DVDD.n3938 DVDD 0.610636
R3303 DVDD.n3890 DVDD 0.610636
R3304 DVDD.n609 DVDD.n260 0.590794
R3305 DVDD.n5516 DVDD.n553 0.583456
R3306 DVDD.n5546 DVDD.n5545 0.58288
R3307 DVDD.n5933 DVDD.t61 0.58122
R3308 DVDD.n5894 DVDD.t12 0.58122
R3309 DVDD.n5546 DVDD.n543 0.56985
R3310 DVDD.n5524 DVDD.n553 0.569671
R3311 DVDD.n5478 DVDD.n5477 0.566831
R3312 DVDD.n3897 DVDD.n3667 0.555174
R3313 DVDD.n3900 DVDD.n3894 0.555174
R3314 DVDD.n3838 DVDD.n3510 0.555174
R3315 DVDD.n3841 DVDD.n3527 0.555174
R3316 DVDD.n5509 DVDD.n5508 0.555174
R3317 DVDD.n5506 DVDD.n5503 0.555174
R3318 DVDD.n5512 DVDD.n5511 0.553707
R3319 DVDD.n5501 DVDD.n5500 0.553707
R3320 DVDD.n611 DVDD.n609 0.545794
R3321 DVDD.n613 DVDD.n611 0.545794
R3322 DVDD.n615 DVDD.n613 0.545794
R3323 DVDD.n5477 DVDD.n5476 0.545794
R3324 DVDD.n5476 DVDD.n5475 0.545794
R3325 DVDD.n5475 DVDD.n5474 0.545794
R3326 DVDD.n625 DVDD.n624 0.545794
R3327 DVDD.n624 DVDD.n607 0.545794
R3328 DVDD.n5709 DVDD.n5708 0.545794
R3329 DVDD.n5708 DVDD.n5707 0.545794
R3330 DVDD.n3697 DVDD.n3666 0.52925
R3331 DVDD.n3893 DVDD.n3549 0.52925
R3332 DVDD.n4205 DVDD.n4204 0.52925
R3333 DVDD.n4186 DVDD.n4185 0.52925
R3334 DVDD.n5479 DVDD.n615 0.514169
R3335 DVDD.n4121 DVDD.n4120 0.511554
R3336 DVDD.n3761 DVDD.n3760 0.511554
R3337 DVDD.n5474 DVDD.n5473 0.4955
R3338 DVDD.n3892 DVDD.n3891 0.49415
R3339 DVDD.n3919 DVDD.n3918 0.49415
R3340 DVDD.n2710 DVDD.n2709 0.4505
R3341 DVDD.n2708 DVDD.n2673 0.4505
R3342 DVDD.n2677 DVDD.n2674 0.4505
R3343 DVDD.n2704 DVDD.n2703 0.4505
R3344 DVDD.n2702 DVDD.n2676 0.4505
R3345 DVDD.n2701 DVDD.n2700 0.4505
R3346 DVDD.n2679 DVDD.n2678 0.4505
R3347 DVDD.n2696 DVDD.n2695 0.4505
R3348 DVDD.n2694 DVDD.n2681 0.4505
R3349 DVDD.n2693 DVDD.n2692 0.4505
R3350 DVDD.n2683 DVDD.n2682 0.4505
R3351 DVDD.n2688 DVDD.n2687 0.4505
R3352 DVDD.n2686 DVDD.n2685 0.4505
R3353 DVDD.n2904 DVDD.n2864 0.4505
R3354 DVDD.n2903 DVDD.n2866 0.4505
R3355 DVDD.n2869 DVDD.n2865 0.4505
R3356 DVDD.n2899 DVDD.n2898 0.4505
R3357 DVDD.n2897 DVDD.n2868 0.4505
R3358 DVDD.n2896 DVDD.n2895 0.4505
R3359 DVDD.n2871 DVDD.n2870 0.4505
R3360 DVDD.n2891 DVDD.n2890 0.4505
R3361 DVDD.n2889 DVDD.n2873 0.4505
R3362 DVDD.n2888 DVDD.n2887 0.4505
R3363 DVDD.n2875 DVDD.n2874 0.4505
R3364 DVDD.n2883 DVDD.n2882 0.4505
R3365 DVDD.n2881 DVDD.n2877 0.4505
R3366 DVDD.n2880 DVDD.n2879 0.4505
R3367 DVDD.n490 DVDD.n488 0.4505
R3368 DVDD.n5607 DVDD.n5606 0.4505
R3369 DVDD.n5605 DVDD.n489 0.4505
R3370 DVDD.n5604 DVDD.n5603 0.4505
R3371 DVDD.n5602 DVDD.n491 0.4505
R3372 DVDD.n495 DVDD.n492 0.4505
R3373 DVDD.n5598 DVDD.n5597 0.4505
R3374 DVDD.n5596 DVDD.n494 0.4505
R3375 DVDD.n5595 DVDD.n5594 0.4505
R3376 DVDD.n497 DVDD.n496 0.4505
R3377 DVDD.n5590 DVDD.n5589 0.4505
R3378 DVDD.n5588 DVDD.n499 0.4505
R3379 DVDD.n5587 DVDD.n5586 0.4505
R3380 DVDD.n501 DVDD.n500 0.4505
R3381 DVDD.n5582 DVDD.n5581 0.4505
R3382 DVDD.n5580 DVDD.n503 0.4505
R3383 DVDD.n5579 DVDD.n5578 0.4505
R3384 DVDD.n505 DVDD.n504 0.4505
R3385 DVDD.n5574 DVDD.n5573 0.4505
R3386 DVDD.n5572 DVDD.n507 0.4505
R3387 DVDD.n5571 DVDD.n5570 0.4505
R3388 DVDD.n509 DVDD.n508 0.4505
R3389 DVDD.n2632 DVDD.n2631 0.4505
R3390 DVDD.n2633 DVDD.n2629 0.4505
R3391 DVDD.n2635 DVDD.n2634 0.4505
R3392 DVDD.n2627 DVDD.n2626 0.4505
R3393 DVDD.n2640 DVDD.n2639 0.4505
R3394 DVDD.n2641 DVDD.n2625 0.4505
R3395 DVDD.n2643 DVDD.n2642 0.4505
R3396 DVDD.n2623 DVDD.n2622 0.4505
R3397 DVDD.n2648 DVDD.n2647 0.4505
R3398 DVDD.n2649 DVDD.n2621 0.4505
R3399 DVDD.n2651 DVDD.n2650 0.4505
R3400 DVDD.n2619 DVDD.n2618 0.4505
R3401 DVDD.n2656 DVDD.n2655 0.4505
R3402 DVDD.n2657 DVDD.n2616 0.4505
R3403 DVDD.n2746 DVDD.n2745 0.4505
R3404 DVDD.n2744 DVDD.n2617 0.4505
R3405 DVDD.n2743 DVDD.n2742 0.4505
R3406 DVDD.n2741 DVDD.n2658 0.4505
R3407 DVDD.n2662 DVDD.n2659 0.4505
R3408 DVDD.n2737 DVDD.n2736 0.4505
R3409 DVDD.n2735 DVDD.n2661 0.4505
R3410 DVDD.n2734 DVDD.n2733 0.4505
R3411 DVDD.n2664 DVDD.n2663 0.4505
R3412 DVDD.n2729 DVDD.n2728 0.4505
R3413 DVDD.n2727 DVDD.n2666 0.4505
R3414 DVDD.n2726 DVDD.n2725 0.4505
R3415 DVDD.n2668 DVDD.n2667 0.4505
R3416 DVDD.n2721 DVDD.n2720 0.4505
R3417 DVDD.n2719 DVDD.n2670 0.4505
R3418 DVDD.n2718 DVDD.n2717 0.4505
R3419 DVDD.n2714 DVDD.n2671 0.4505
R3420 DVDD.n2713 DVDD.n2712 0.4505
R3421 DVDD.n2711 DVDD.n2672 0.4505
R3422 DVDD.n2689 DVDD.n2688 0.4505
R3423 DVDD.n2690 DVDD.n2683 0.4505
R3424 DVDD.n2692 DVDD.n2691 0.4505
R3425 DVDD.n2681 DVDD.n2680 0.4505
R3426 DVDD.n2697 DVDD.n2696 0.4505
R3427 DVDD.n2698 DVDD.n2679 0.4505
R3428 DVDD.n2700 DVDD.n2699 0.4505
R3429 DVDD.n2676 DVDD.n2675 0.4505
R3430 DVDD.n2705 DVDD.n2704 0.4505
R3431 DVDD.n2706 DVDD.n2674 0.4505
R3432 DVDD.n2708 DVDD.n2707 0.4505
R3433 DVDD.n2709 DVDD.n2578 0.4505
R3434 DVDD.n2905 DVDD.n2589 0.4505
R3435 DVDD.n2904 DVDD.n2591 0.4505
R3436 DVDD.n2903 DVDD.n2902 0.4505
R3437 DVDD.n2901 DVDD.n2865 0.4505
R3438 DVDD.n2900 DVDD.n2899 0.4505
R3439 DVDD.n2868 DVDD.n2867 0.4505
R3440 DVDD.n2895 DVDD.n2894 0.4505
R3441 DVDD.n2893 DVDD.n2871 0.4505
R3442 DVDD.n2892 DVDD.n2891 0.4505
R3443 DVDD.n2873 DVDD.n2872 0.4505
R3444 DVDD.n2887 DVDD.n2886 0.4505
R3445 DVDD.n2885 DVDD.n2875 0.4505
R3446 DVDD.n2884 DVDD.n2883 0.4505
R3447 DVDD.n2877 DVDD.n2876 0.4505
R3448 DVDD.n2879 DVDD.n2878 0.4505
R3449 DVDD.n488 DVDD.n487 0.4505
R3450 DVDD.n5608 DVDD.n5607 0.4505
R3451 DVDD.n489 DVDD.n478 0.4505
R3452 DVDD.n5603 DVDD.n481 0.4505
R3453 DVDD.n5602 DVDD.n5601 0.4505
R3454 DVDD.n5600 DVDD.n492 0.4505
R3455 DVDD.n5599 DVDD.n5598 0.4505
R3456 DVDD.n494 DVDD.n493 0.4505
R3457 DVDD.n5594 DVDD.n5593 0.4505
R3458 DVDD.n5592 DVDD.n497 0.4505
R3459 DVDD.n5591 DVDD.n5590 0.4505
R3460 DVDD.n499 DVDD.n498 0.4505
R3461 DVDD.n5586 DVDD.n5585 0.4505
R3462 DVDD.n5584 DVDD.n501 0.4505
R3463 DVDD.n5583 DVDD.n5582 0.4505
R3464 DVDD.n503 DVDD.n502 0.4505
R3465 DVDD.n5578 DVDD.n5577 0.4505
R3466 DVDD.n5576 DVDD.n505 0.4505
R3467 DVDD.n5575 DVDD.n5574 0.4505
R3468 DVDD.n2595 DVDD.n507 0.4505
R3469 DVDD.n5570 DVDD.n5569 0.4505
R3470 DVDD.n516 DVDD.n509 0.4505
R3471 DVDD.n2631 DVDD.n2630 0.4505
R3472 DVDD.n2629 DVDD.n2628 0.4505
R3473 DVDD.n2636 DVDD.n2635 0.4505
R3474 DVDD.n2637 DVDD.n2627 0.4505
R3475 DVDD.n2639 DVDD.n2638 0.4505
R3476 DVDD.n2625 DVDD.n2624 0.4505
R3477 DVDD.n2644 DVDD.n2643 0.4505
R3478 DVDD.n2645 DVDD.n2623 0.4505
R3479 DVDD.n2647 DVDD.n2646 0.4505
R3480 DVDD.n2621 DVDD.n2620 0.4505
R3481 DVDD.n2652 DVDD.n2651 0.4505
R3482 DVDD.n2653 DVDD.n2619 0.4505
R3483 DVDD.n2655 DVDD.n2654 0.4505
R3484 DVDD.n2616 DVDD.n2615 0.4505
R3485 DVDD.n2747 DVDD.n2746 0.4505
R3486 DVDD.n2617 DVDD.n2607 0.4505
R3487 DVDD.n2742 DVDD.n2609 0.4505
R3488 DVDD.n2741 DVDD.n2740 0.4505
R3489 DVDD.n2739 DVDD.n2659 0.4505
R3490 DVDD.n2738 DVDD.n2737 0.4505
R3491 DVDD.n2661 DVDD.n2660 0.4505
R3492 DVDD.n2733 DVDD.n2732 0.4505
R3493 DVDD.n2731 DVDD.n2664 0.4505
R3494 DVDD.n2730 DVDD.n2729 0.4505
R3495 DVDD.n2666 DVDD.n2665 0.4505
R3496 DVDD.n2725 DVDD.n2724 0.4505
R3497 DVDD.n2723 DVDD.n2668 0.4505
R3498 DVDD.n2722 DVDD.n2721 0.4505
R3499 DVDD.n2670 DVDD.n2669 0.4505
R3500 DVDD.n2717 DVDD.n2716 0.4505
R3501 DVDD.n2715 DVDD.n2714 0.4505
R3502 DVDD.n2713 DVDD.n2583 0.4505
R3503 DVDD.n2672 DVDD.n2575 0.4505
R3504 DVDD.n678 DVDD.n677 0.4505
R3505 DVDD.n679 DVDD.n670 0.4505
R3506 DVDD.n681 DVDD.n680 0.4505
R3507 DVDD.n668 DVDD.n667 0.4505
R3508 DVDD.n686 DVDD.n685 0.4505
R3509 DVDD.n687 DVDD.n665 0.4505
R3510 DVDD.n689 DVDD.n688 0.4505
R3511 DVDD.n666 DVDD.n663 0.4505
R3512 DVDD.n693 DVDD.n662 0.4505
R3513 DVDD.n695 DVDD.n694 0.4505
R3514 DVDD.n5433 DVDD.n657 0.4505
R3515 DVDD.n5453 DVDD.n5452 0.4505
R3516 DVDD.n5451 DVDD.n648 0.4505
R3517 DVDD.n5450 DVDD.n5449 0.4505
R3518 DVDD.n650 DVDD.n649 0.4505
R3519 DVDD.n5445 DVDD.n5444 0.4505
R3520 DVDD.n5443 DVDD.n652 0.4505
R3521 DVDD.n5442 DVDD.n5441 0.4505
R3522 DVDD.n654 DVDD.n653 0.4505
R3523 DVDD.n5437 DVDD.n5436 0.4505
R3524 DVDD.n5433 DVDD.n5432 0.4505
R3525 DVDD.n694 DVDD.n658 0.4505
R3526 DVDD.n693 DVDD.n692 0.4505
R3527 DVDD.n691 DVDD.n663 0.4505
R3528 DVDD.n690 DVDD.n689 0.4505
R3529 DVDD.n665 DVDD.n664 0.4505
R3530 DVDD.n685 DVDD.n684 0.4505
R3531 DVDD.n683 DVDD.n668 0.4505
R3532 DVDD.n682 DVDD.n681 0.4505
R3533 DVDD.n670 DVDD.n669 0.4505
R3534 DVDD.n677 DVDD.n676 0.4505
R3535 DVDD.n5454 DVDD.n5453 0.4505
R3536 DVDD.n648 DVDD.n647 0.4505
R3537 DVDD.n5449 DVDD.n5448 0.4505
R3538 DVDD.n5447 DVDD.n650 0.4505
R3539 DVDD.n5446 DVDD.n5445 0.4505
R3540 DVDD.n652 DVDD.n651 0.4505
R3541 DVDD.n5441 DVDD.n5440 0.4505
R3542 DVDD.n5439 DVDD.n654 0.4505
R3543 DVDD.n5438 DVDD.n5437 0.4505
R3544 DVDD.n5435 DVDD.n655 0.4505
R3545 DVDD.n5435 DVDD.n5434 0.4505
R3546 DVDD.n5037 DVDD.n5036 0.4505
R3547 DVDD.n5039 DVDD.n5038 0.4505
R3548 DVDD.n5009 DVDD.n5008 0.4505
R3549 DVDD.n5044 DVDD.n5043 0.4505
R3550 DVDD.n5045 DVDD.n5007 0.4505
R3551 DVDD.n5047 DVDD.n5046 0.4505
R3552 DVDD.n5005 DVDD.n5004 0.4505
R3553 DVDD.n5052 DVDD.n5051 0.4505
R3554 DVDD.n5053 DVDD.n5003 0.4505
R3555 DVDD.n5056 DVDD.n5055 0.4505
R3556 DVDD.n5054 DVDD.n5000 0.4505
R3557 DVDD.n5061 DVDD.n5001 0.4505
R3558 DVDD.n5067 DVDD.n5066 0.4505
R3559 DVDD.n5065 DVDD.n5060 0.4505
R3560 DVDD.n5064 DVDD.n5063 0.4505
R3561 DVDD.n639 DVDD.n628 0.4505
R3562 DVDD.n5468 DVDD.n5467 0.4505
R3563 DVDD.n644 DVDD.n640 0.4505
R3564 DVDD.n5463 DVDD.n5462 0.4505
R3565 DVDD.n5461 DVDD.n643 0.4505
R3566 DVDD.n5460 DVDD.n5459 0.4505
R3567 DVDD.n5036 DVDD.n5010 0.4505
R3568 DVDD.n5040 DVDD.n5039 0.4505
R3569 DVDD.n5041 DVDD.n5009 0.4505
R3570 DVDD.n5043 DVDD.n5042 0.4505
R3571 DVDD.n5007 DVDD.n5006 0.4505
R3572 DVDD.n5048 DVDD.n5047 0.4505
R3573 DVDD.n5049 DVDD.n5005 0.4505
R3574 DVDD.n5051 DVDD.n5050 0.4505
R3575 DVDD.n5003 DVDD.n5002 0.4505
R3576 DVDD.n5057 DVDD.n5056 0.4505
R3577 DVDD.n5058 DVDD.n5000 0.4505
R3578 DVDD.n5069 DVDD.n5001 0.4505
R3579 DVDD.n5068 DVDD.n5067 0.4505
R3580 DVDD.n5060 DVDD.n5059 0.4505
R3581 DVDD.n5063 DVDD.n5062 0.4505
R3582 DVDD.n641 DVDD.n639 0.4505
R3583 DVDD.n5467 DVDD.n5466 0.4505
R3584 DVDD.n5465 DVDD.n640 0.4505
R3585 DVDD.n5464 DVDD.n5463 0.4505
R3586 DVDD.n643 DVDD.n642 0.4505
R3587 DVDD.n5459 DVDD.n5458 0.4505
R3588 DVDD.n860 DVDD.n848 0.4505
R3589 DVDD.n859 DVDD.n858 0.4505
R3590 DVDD.n857 DVDD.n852 0.4505
R3591 DVDD.n856 DVDD.n855 0.4505
R3592 DVDD.n274 DVDD.n263 0.4505
R3593 DVDD.n5702 DVDD.n5701 0.4505
R3594 DVDD.n279 DVDD.n275 0.4505
R3595 DVDD.n5697 DVDD.n5696 0.4505
R3596 DVDD.n5695 DVDD.n278 0.4505
R3597 DVDD.n5694 DVDD.n5693 0.4505
R3598 DVDD.n281 DVDD.n280 0.4505
R3599 DVDD.n5688 DVDD.n5687 0.4505
R3600 DVDD.n5686 DVDD.n286 0.4505
R3601 DVDD.n5685 DVDD.n5684 0.4505
R3602 DVDD.n289 DVDD.n288 0.4505
R3603 DVDD.n5680 DVDD.n5679 0.4505
R3604 DVDD.n5678 DVDD.n291 0.4505
R3605 DVDD.n5677 DVDD.n5676 0.4505
R3606 DVDD.n293 DVDD.n292 0.4505
R3607 DVDD.n5672 DVDD.n5671 0.4505
R3608 DVDD.n5670 DVDD.n295 0.4505
R3609 DVDD.n861 DVDD.n860 0.4505
R3610 DVDD.n859 DVDD.n851 0.4505
R3611 DVDD.n853 DVDD.n852 0.4505
R3612 DVDD.n855 DVDD.n854 0.4505
R3613 DVDD.n276 DVDD.n274 0.4505
R3614 DVDD.n5701 DVDD.n5700 0.4505
R3615 DVDD.n5699 DVDD.n275 0.4505
R3616 DVDD.n5698 DVDD.n5697 0.4505
R3617 DVDD.n278 DVDD.n277 0.4505
R3618 DVDD.n5693 DVDD.n5692 0.4505
R3619 DVDD.n5691 DVDD.n281 0.4505
R3620 DVDD.n5689 DVDD.n5688 0.4505
R3621 DVDD.n286 DVDD.n284 0.4505
R3622 DVDD.n5684 DVDD.n5683 0.4505
R3623 DVDD.n5682 DVDD.n289 0.4505
R3624 DVDD.n5681 DVDD.n5680 0.4505
R3625 DVDD.n291 DVDD.n290 0.4505
R3626 DVDD.n5676 DVDD.n5675 0.4505
R3627 DVDD.n5674 DVDD.n293 0.4505
R3628 DVDD.n5673 DVDD.n5672 0.4505
R3629 DVDD.n295 DVDD.n294 0.4505
R3630 DVDD.n806 DVDD.n800 0.4505
R3631 DVDD.n808 DVDD.n807 0.4505
R3632 DVDD.n798 DVDD.n797 0.4505
R3633 DVDD.n813 DVDD.n812 0.4505
R3634 DVDD.n814 DVDD.n796 0.4505
R3635 DVDD.n816 DVDD.n815 0.4505
R3636 DVDD.n794 DVDD.n793 0.4505
R3637 DVDD.n821 DVDD.n820 0.4505
R3638 DVDD.n822 DVDD.n792 0.4505
R3639 DVDD.n825 DVDD.n824 0.4505
R3640 DVDD.n823 DVDD.n788 0.4505
R3641 DVDD.n2976 DVDD.n790 0.4505
R3642 DVDD.n841 DVDD.n789 0.4505
R3643 DVDD.n879 DVDD.n878 0.4505
R3644 DVDD.n877 DVDD.n840 0.4505
R3645 DVDD.n876 DVDD.n875 0.4505
R3646 DVDD.n843 DVDD.n842 0.4505
R3647 DVDD.n871 DVDD.n870 0.4505
R3648 DVDD.n869 DVDD.n845 0.4505
R3649 DVDD.n868 DVDD.n867 0.4505
R3650 DVDD.n847 DVDD.n846 0.4505
R3651 DVDD.n800 DVDD.n799 0.4505
R3652 DVDD.n809 DVDD.n808 0.4505
R3653 DVDD.n810 DVDD.n798 0.4505
R3654 DVDD.n812 DVDD.n811 0.4505
R3655 DVDD.n796 DVDD.n795 0.4505
R3656 DVDD.n817 DVDD.n816 0.4505
R3657 DVDD.n818 DVDD.n794 0.4505
R3658 DVDD.n820 DVDD.n819 0.4505
R3659 DVDD.n792 DVDD.n791 0.4505
R3660 DVDD.n826 DVDD.n825 0.4505
R3661 DVDD.n827 DVDD.n788 0.4505
R3662 DVDD.n2976 DVDD.n2975 0.4505
R3663 DVDD.n2973 DVDD.n789 0.4505
R3664 DVDD.n880 DVDD.n879 0.4505
R3665 DVDD.n840 DVDD.n839 0.4505
R3666 DVDD.n875 DVDD.n874 0.4505
R3667 DVDD.n873 DVDD.n843 0.4505
R3668 DVDD.n872 DVDD.n871 0.4505
R3669 DVDD.n845 DVDD.n844 0.4505
R3670 DVDD.n867 DVDD.n866 0.4505
R3671 DVDD.n865 DVDD.n847 0.4505
R3672 DVDD.n4080 DVDD.n4079 0.4505
R3673 DVDD.n4082 DVDD.n4081 0.4505
R3674 DVDD.n4077 DVDD.n4076 0.4505
R3675 DVDD.n4087 DVDD.n4086 0.4505
R3676 DVDD.n4088 DVDD.n4075 0.4505
R3677 DVDD.n4090 DVDD.n4089 0.4505
R3678 DVDD.n4073 DVDD.n4072 0.4505
R3679 DVDD.n4095 DVDD.n4094 0.4505
R3680 DVDD.n4096 DVDD.n4070 0.4505
R3681 DVDD.n4098 DVDD.n4097 0.4505
R3682 DVDD.n4071 DVDD.n4068 0.4505
R3683 DVDD.n4102 DVDD.n4067 0.4505
R3684 DVDD.n4104 DVDD.n4103 0.4505
R3685 DVDD.n3743 DVDD.n3742 0.4505
R3686 DVDD.n3741 DVDD.n3703 0.4505
R3687 DVDD.n3740 DVDD.n3739 0.4505
R3688 DVDD.n3706 DVDD.n3705 0.4505
R3689 DVDD.n3735 DVDD.n3734 0.4505
R3690 DVDD.n3733 DVDD.n3708 0.4505
R3691 DVDD.n3732 DVDD.n3731 0.4505
R3692 DVDD.n3710 DVDD.n3709 0.4505
R3693 DVDD.n3727 DVDD.n3726 0.4505
R3694 DVDD.n3725 DVDD.n3712 0.4505
R3695 DVDD.n3724 DVDD.n3723 0.4505
R3696 DVDD.n3714 DVDD.n3713 0.4505
R3697 DVDD.n3719 DVDD.n3718 0.4505
R3698 DVDD.n3717 DVDD.n3716 0.4505
R3699 DVDD.n3647 DVDD.n3646 0.4505
R3700 DVDD.n3959 DVDD.n3958 0.4505
R3701 DVDD.n3960 DVDD.n3645 0.4505
R3702 DVDD.n3962 DVDD.n3961 0.4505
R3703 DVDD.n3643 DVDD.n3642 0.4505
R3704 DVDD.n3967 DVDD.n3966 0.4505
R3705 DVDD.n3968 DVDD.n3641 0.4505
R3706 DVDD.n3970 DVDD.n3969 0.4505
R3707 DVDD.n3639 DVDD.n3638 0.4505
R3708 DVDD.n3975 DVDD.n3974 0.4505
R3709 DVDD.n3976 DVDD.n3637 0.4505
R3710 DVDD.n3978 DVDD.n3977 0.4505
R3711 DVDD.n3635 DVDD.n3634 0.4505
R3712 DVDD.n3983 DVDD.n3982 0.4505
R3713 DVDD.n3984 DVDD.n3633 0.4505
R3714 DVDD.n3986 DVDD.n3985 0.4505
R3715 DVDD.n3631 DVDD.n3630 0.4505
R3716 DVDD.n3992 DVDD.n3991 0.4505
R3717 DVDD.n3993 DVDD.n3628 0.4505
R3718 DVDD.n3996 DVDD.n3995 0.4505
R3719 DVDD.n3994 DVDD.n3629 0.4505
R3720 DVDD.n3604 DVDD.n3603 0.4505
R3721 DVDD.n4005 DVDD.n4004 0.4505
R3722 DVDD.n4006 DVDD.n3602 0.4505
R3723 DVDD.n4008 DVDD.n4007 0.4505
R3724 DVDD.n3600 DVDD.n3599 0.4505
R3725 DVDD.n4013 DVDD.n4012 0.4505
R3726 DVDD.n4014 DVDD.n3598 0.4505
R3727 DVDD.n4016 DVDD.n4015 0.4505
R3728 DVDD.n3596 DVDD.n3595 0.4505
R3729 DVDD.n4021 DVDD.n4020 0.4505
R3730 DVDD.n4022 DVDD.n3594 0.4505
R3731 DVDD.n4024 DVDD.n4023 0.4505
R3732 DVDD.n3592 DVDD.n3591 0.4505
R3733 DVDD.n4029 DVDD.n4028 0.4505
R3734 DVDD.n4030 DVDD.n3589 0.4505
R3735 DVDD.n4033 DVDD.n4032 0.4505
R3736 DVDD.n4031 DVDD.n3590 0.4505
R3737 DVDD.n3574 DVDD.n3573 0.4505
R3738 DVDD.n4041 DVDD.n4040 0.4505
R3739 DVDD.n4042 DVDD.n3572 0.4505
R3740 DVDD.n4044 DVDD.n4043 0.4505
R3741 DVDD.n3570 DVDD.n3569 0.4505
R3742 DVDD.n4049 DVDD.n4048 0.4505
R3743 DVDD.n4050 DVDD.n3568 0.4505
R3744 DVDD.n4052 DVDD.n4051 0.4505
R3745 DVDD.n3566 DVDD.n3565 0.4505
R3746 DVDD.n4057 DVDD.n4056 0.4505
R3747 DVDD.n4058 DVDD.n3564 0.4505
R3748 DVDD.n4060 DVDD.n4059 0.4505
R3749 DVDD.n3562 DVDD.n3561 0.4505
R3750 DVDD.n4065 DVDD.n4064 0.4505
R3751 DVDD.n4066 DVDD.n3559 0.4505
R3752 DVDD.n4107 DVDD.n4106 0.4505
R3753 DVDD.n4105 DVDD.n3560 0.4505
R3754 DVDD.n4083 DVDD.n4082 0.4505
R3755 DVDD.n4084 DVDD.n4077 0.4505
R3756 DVDD.n4086 DVDD.n4085 0.4505
R3757 DVDD.n4075 DVDD.n4074 0.4505
R3758 DVDD.n4091 DVDD.n4090 0.4505
R3759 DVDD.n4092 DVDD.n4073 0.4505
R3760 DVDD.n4094 DVDD.n4093 0.4505
R3761 DVDD.n4070 DVDD.n4069 0.4505
R3762 DVDD.n4099 DVDD.n4098 0.4505
R3763 DVDD.n4100 DVDD.n4068 0.4505
R3764 DVDD.n4102 DVDD.n4101 0.4505
R3765 DVDD.n4103 DVDD.n3553 0.4505
R3766 DVDD.n3702 DVDD.n3700 0.4505
R3767 DVDD.n3744 DVDD.n3743 0.4505
R3768 DVDD.n3703 DVDD.n3701 0.4505
R3769 DVDD.n3739 DVDD.n3738 0.4505
R3770 DVDD.n3737 DVDD.n3706 0.4505
R3771 DVDD.n3736 DVDD.n3735 0.4505
R3772 DVDD.n3708 DVDD.n3707 0.4505
R3773 DVDD.n3731 DVDD.n3730 0.4505
R3774 DVDD.n3729 DVDD.n3710 0.4505
R3775 DVDD.n3728 DVDD.n3727 0.4505
R3776 DVDD.n3712 DVDD.n3711 0.4505
R3777 DVDD.n3723 DVDD.n3722 0.4505
R3778 DVDD.n3721 DVDD.n3714 0.4505
R3779 DVDD.n3720 DVDD.n3719 0.4505
R3780 DVDD.n3716 DVDD.n3715 0.4505
R3781 DVDD.n3648 DVDD.n3647 0.4505
R3782 DVDD.n3958 DVDD.n3957 0.4505
R3783 DVDD.n3654 DVDD.n3645 0.4505
R3784 DVDD.n3963 DVDD.n3962 0.4505
R3785 DVDD.n3964 DVDD.n3643 0.4505
R3786 DVDD.n3966 DVDD.n3965 0.4505
R3787 DVDD.n3641 DVDD.n3640 0.4505
R3788 DVDD.n3971 DVDD.n3970 0.4505
R3789 DVDD.n3972 DVDD.n3639 0.4505
R3790 DVDD.n3974 DVDD.n3973 0.4505
R3791 DVDD.n3637 DVDD.n3636 0.4505
R3792 DVDD.n3979 DVDD.n3978 0.4505
R3793 DVDD.n3980 DVDD.n3635 0.4505
R3794 DVDD.n3982 DVDD.n3981 0.4505
R3795 DVDD.n3633 DVDD.n3632 0.4505
R3796 DVDD.n3987 DVDD.n3986 0.4505
R3797 DVDD.n3988 DVDD.n3631 0.4505
R3798 DVDD.n3991 DVDD.n3990 0.4505
R3799 DVDD.n3989 DVDD.n3628 0.4505
R3800 DVDD.n3997 DVDD.n3996 0.4505
R3801 DVDD.n3629 DVDD.n3605 0.4505
R3802 DVDD.n4002 DVDD.n3604 0.4505
R3803 DVDD.n4004 DVDD.n4003 0.4505
R3804 DVDD.n3602 DVDD.n3601 0.4505
R3805 DVDD.n4009 DVDD.n4008 0.4505
R3806 DVDD.n4010 DVDD.n3600 0.4505
R3807 DVDD.n4012 DVDD.n4011 0.4505
R3808 DVDD.n3598 DVDD.n3597 0.4505
R3809 DVDD.n4017 DVDD.n4016 0.4505
R3810 DVDD.n4018 DVDD.n3596 0.4505
R3811 DVDD.n4020 DVDD.n4019 0.4505
R3812 DVDD.n3594 DVDD.n3593 0.4505
R3813 DVDD.n4025 DVDD.n4024 0.4505
R3814 DVDD.n4026 DVDD.n3592 0.4505
R3815 DVDD.n4028 DVDD.n4027 0.4505
R3816 DVDD.n3589 DVDD.n3588 0.4505
R3817 DVDD.n4034 DVDD.n4033 0.4505
R3818 DVDD.n3590 DVDD.n3575 0.4505
R3819 DVDD.n4038 DVDD.n3574 0.4505
R3820 DVDD.n4040 DVDD.n4039 0.4505
R3821 DVDD.n3572 DVDD.n3571 0.4505
R3822 DVDD.n4045 DVDD.n4044 0.4505
R3823 DVDD.n4046 DVDD.n3570 0.4505
R3824 DVDD.n4048 DVDD.n4047 0.4505
R3825 DVDD.n3568 DVDD.n3567 0.4505
R3826 DVDD.n4053 DVDD.n4052 0.4505
R3827 DVDD.n4054 DVDD.n3566 0.4505
R3828 DVDD.n4056 DVDD.n4055 0.4505
R3829 DVDD.n3564 DVDD.n3563 0.4505
R3830 DVDD.n4061 DVDD.n4060 0.4505
R3831 DVDD.n4062 DVDD.n3562 0.4505
R3832 DVDD.n4064 DVDD.n4063 0.4505
R3833 DVDD.n3559 DVDD.n3558 0.4505
R3834 DVDD.n4108 DVDD.n4107 0.4505
R3835 DVDD.n3560 DVDD.n3552 0.4505
R3836 DVDD.n5994 DVDD.n5993 0.4505
R3837 DVDD.n6015 DVDD.n0 0.4505
R3838 DVDD.n6014 DVDD.n6013 0.4505
R3839 DVDD.n6012 DVDD.n2 0.4505
R3840 DVDD.n6011 DVDD.n6010 0.4505
R3841 DVDD.n4 DVDD.n3 0.4505
R3842 DVDD.n6005 DVDD.n6004 0.4505
R3843 DVDD.n6003 DVDD.n6 0.4505
R3844 DVDD.n6002 DVDD.n6001 0.4505
R3845 DVDD.n8 DVDD.n7 0.4505
R3846 DVDD.n5997 DVDD.n5996 0.4505
R3847 DVDD.n5995 DVDD.n10 0.4505
R3848 DVDD.n4211 DVDD.n3483 0.4505
R3849 DVDD.n4326 DVDD.n3482 0.4505
R3850 DVDD.n4328 DVDD.n4327 0.4505
R3851 DVDD.n3480 DVDD.n3479 0.4505
R3852 DVDD.n4333 DVDD.n4332 0.4505
R3853 DVDD.n4334 DVDD.n3478 0.4505
R3854 DVDD.n4336 DVDD.n4335 0.4505
R3855 DVDD.n3476 DVDD.n3475 0.4505
R3856 DVDD.n4341 DVDD.n4340 0.4505
R3857 DVDD.n4342 DVDD.n3474 0.4505
R3858 DVDD.n4344 DVDD.n4343 0.4505
R3859 DVDD.n3472 DVDD.n3471 0.4505
R3860 DVDD.n4349 DVDD.n4348 0.4505
R3861 DVDD.n4350 DVDD.n3470 0.4505
R3862 DVDD.n4353 DVDD.n4352 0.4505
R3863 DVDD.n4351 DVDD.n3467 0.4505
R3864 DVDD.n4357 DVDD.n3468 0.4505
R3865 DVDD.n4359 DVDD.n4358 0.4505
R3866 DVDD.n4361 DVDD.n4360 0.4505
R3867 DVDD.n3465 DVDD.n3464 0.4505
R3868 DVDD.n4366 DVDD.n4365 0.4505
R3869 DVDD.n4367 DVDD.n3463 0.4505
R3870 DVDD.n4369 DVDD.n4368 0.4505
R3871 DVDD.n3461 DVDD.n3460 0.4505
R3872 DVDD.n4374 DVDD.n4373 0.4505
R3873 DVDD.n4375 DVDD.n3459 0.4505
R3874 DVDD.n4377 DVDD.n4376 0.4505
R3875 DVDD.n3457 DVDD.n3456 0.4505
R3876 DVDD.n4382 DVDD.n4381 0.4505
R3877 DVDD.n4383 DVDD.n3455 0.4505
R3878 DVDD.n4386 DVDD.n4385 0.4505
R3879 DVDD.n4384 DVDD.n3452 0.4505
R3880 DVDD.n4390 DVDD.n3453 0.4505
R3881 DVDD.n4391 DVDD.n3433 0.4505
R3882 DVDD.n4392 DVDD.n3438 0.4505
R3883 DVDD.n3449 DVDD.n3441 0.4505
R3884 DVDD.n4485 DVDD.n4484 0.4505
R3885 DVDD.n3450 DVDD.n3448 0.4505
R3886 DVDD.n4480 DVDD.n4479 0.4505
R3887 DVDD.n4478 DVDD.n4396 0.4505
R3888 DVDD.n4477 DVDD.n4476 0.4505
R3889 DVDD.n4398 DVDD.n4397 0.4505
R3890 DVDD.n4472 DVDD.n4471 0.4505
R3891 DVDD.n4470 DVDD.n4400 0.4505
R3892 DVDD.n4469 DVDD.n4468 0.4505
R3893 DVDD.n4402 DVDD.n4401 0.4505
R3894 DVDD.n4464 DVDD.n4463 0.4505
R3895 DVDD.n4462 DVDD.n4404 0.4505
R3896 DVDD.n4461 DVDD.n4460 0.4505
R3897 DVDD.n4406 DVDD.n4405 0.4505
R3898 DVDD.n4456 DVDD.n4455 0.4505
R3899 DVDD.n4454 DVDD.n4453 0.4505
R3900 DVDD.n4452 DVDD.n4409 0.4505
R3901 DVDD.n4412 DVDD.n4408 0.4505
R3902 DVDD.n4448 DVDD.n4447 0.4505
R3903 DVDD.n4446 DVDD.n4411 0.4505
R3904 DVDD.n4445 DVDD.n4444 0.4505
R3905 DVDD.n4414 DVDD.n4413 0.4505
R3906 DVDD.n4440 DVDD.n4439 0.4505
R3907 DVDD.n4438 DVDD.n4416 0.4505
R3908 DVDD.n4437 DVDD.n4436 0.4505
R3909 DVDD.n4418 DVDD.n4417 0.4505
R3910 DVDD.n4432 DVDD.n4431 0.4505
R3911 DVDD.n4430 DVDD.n4420 0.4505
R3912 DVDD.n4429 DVDD.n4428 0.4505
R3913 DVDD.n4422 DVDD.n4421 0.4505
R3914 DVDD.n4424 DVDD.n4423 0.4505
R3915 DVDD.n15 DVDD.n14 0.4505
R3916 DVDD.n5989 DVDD.n5988 0.4505
R3917 DVDD.n5993 DVDD.n5992 0.4505
R3918 DVDD.n10 DVDD.n9 0.4505
R3919 DVDD.n5998 DVDD.n5997 0.4505
R3920 DVDD.n5999 DVDD.n8 0.4505
R3921 DVDD.n6001 DVDD.n6000 0.4505
R3922 DVDD.n6 DVDD.n5 0.4505
R3923 DVDD.n6006 DVDD.n6005 0.4505
R3924 DVDD.n6007 DVDD.n4 0.4505
R3925 DVDD.n6010 DVDD.n6009 0.4505
R3926 DVDD.n6008 DVDD.n2 0.4505
R3927 DVDD.n6014 DVDD.n1 0.4505
R3928 DVDD.n6016 DVDD.n6015 0.4505
R3929 DVDD.n6018 DVDD.n6017 0.4505
R3930 DVDD.n3482 DVDD.n3481 0.4505
R3931 DVDD.n4329 DVDD.n4328 0.4505
R3932 DVDD.n4330 DVDD.n3480 0.4505
R3933 DVDD.n4332 DVDD.n4331 0.4505
R3934 DVDD.n3478 DVDD.n3477 0.4505
R3935 DVDD.n4337 DVDD.n4336 0.4505
R3936 DVDD.n4338 DVDD.n3476 0.4505
R3937 DVDD.n4340 DVDD.n4339 0.4505
R3938 DVDD.n3474 DVDD.n3473 0.4505
R3939 DVDD.n4345 DVDD.n4344 0.4505
R3940 DVDD.n4346 DVDD.n3472 0.4505
R3941 DVDD.n4348 DVDD.n4347 0.4505
R3942 DVDD.n3470 DVDD.n3469 0.4505
R3943 DVDD.n4354 DVDD.n4353 0.4505
R3944 DVDD.n4355 DVDD.n3467 0.4505
R3945 DVDD.n4357 DVDD.n4356 0.4505
R3946 DVDD.n4359 DVDD.n3466 0.4505
R3947 DVDD.n4362 DVDD.n4361 0.4505
R3948 DVDD.n4363 DVDD.n3465 0.4505
R3949 DVDD.n4365 DVDD.n4364 0.4505
R3950 DVDD.n3463 DVDD.n3462 0.4505
R3951 DVDD.n4370 DVDD.n4369 0.4505
R3952 DVDD.n4371 DVDD.n3461 0.4505
R3953 DVDD.n4373 DVDD.n4372 0.4505
R3954 DVDD.n3459 DVDD.n3458 0.4505
R3955 DVDD.n4378 DVDD.n4377 0.4505
R3956 DVDD.n4379 DVDD.n3457 0.4505
R3957 DVDD.n4381 DVDD.n4380 0.4505
R3958 DVDD.n3455 DVDD.n3454 0.4505
R3959 DVDD.n4387 DVDD.n4386 0.4505
R3960 DVDD.n4388 DVDD.n3452 0.4505
R3961 DVDD.n4390 DVDD.n4389 0.4505
R3962 DVDD.n4391 DVDD.n3451 0.4505
R3963 DVDD.n4393 DVDD.n4392 0.4505
R3964 DVDD.n4394 DVDD.n3449 0.4505
R3965 DVDD.n4484 DVDD.n4483 0.4505
R3966 DVDD.n4482 DVDD.n3450 0.4505
R3967 DVDD.n4481 DVDD.n4480 0.4505
R3968 DVDD.n4396 DVDD.n4395 0.4505
R3969 DVDD.n4476 DVDD.n4475 0.4505
R3970 DVDD.n4474 DVDD.n4398 0.4505
R3971 DVDD.n4473 DVDD.n4472 0.4505
R3972 DVDD.n4400 DVDD.n4399 0.4505
R3973 DVDD.n4468 DVDD.n4467 0.4505
R3974 DVDD.n4466 DVDD.n4402 0.4505
R3975 DVDD.n4465 DVDD.n4464 0.4505
R3976 DVDD.n4404 DVDD.n4403 0.4505
R3977 DVDD.n4460 DVDD.n4459 0.4505
R3978 DVDD.n4458 DVDD.n4406 0.4505
R3979 DVDD.n4457 DVDD.n4456 0.4505
R3980 DVDD.n4453 DVDD.n4407 0.4505
R3981 DVDD.n4452 DVDD.n4451 0.4505
R3982 DVDD.n4450 DVDD.n4408 0.4505
R3983 DVDD.n4449 DVDD.n4448 0.4505
R3984 DVDD.n4411 DVDD.n4410 0.4505
R3985 DVDD.n4444 DVDD.n4443 0.4505
R3986 DVDD.n4442 DVDD.n4414 0.4505
R3987 DVDD.n4441 DVDD.n4440 0.4505
R3988 DVDD.n4416 DVDD.n4415 0.4505
R3989 DVDD.n4436 DVDD.n4435 0.4505
R3990 DVDD.n4434 DVDD.n4418 0.4505
R3991 DVDD.n4433 DVDD.n4432 0.4505
R3992 DVDD.n4420 DVDD.n4419 0.4505
R3993 DVDD.n4428 DVDD.n4427 0.4505
R3994 DVDD.n4426 DVDD.n4422 0.4505
R3995 DVDD.n4425 DVDD.n4424 0.4505
R3996 DVDD.n14 DVDD.n13 0.4505
R3997 DVDD.n5990 DVDD.n5989 0.4505
R3998 DVDD.n5991 DVDD.n12 0.4505
R3999 DVDD.n17 DVDD.n12 0.4505
R4000 DVDD.n3914 DVDD.n3913 0.423265
R4001 DVDD.n3913 DVDD.n3519 0.423265
R4002 DVDD.n4201 DVDD.n3519 0.423265
R4003 DVDD.n3909 DVDD.n3908 0.422275
R4004 DVDD.n3909 DVDD.n3526 0.422275
R4005 DVDD.n4197 DVDD.n3526 0.422275
R4006 DVDD.n5472 DVDD.n625 0.406197
R4007 DVDD.n5707 DVDD.n5706 0.406197
R4008 DVDD.n4120 DVDD.n3550 0.39875
R4009 DVDD.n3760 DVDD.n3698 0.39875
R4010 DVDD.n41 DVDD 0.386971
R4011 DVDD.n4036 DVDD.n3586 0.382843
R4012 DVDD.n3936 DVDD.n3651 0.3828
R4013 DVDD.n608 DVDD.t11 0.3645
R4014 DVDD.n608 DVDD.t26 0.3645
R4015 DVDD.n610 DVDD.t60 0.3645
R4016 DVDD.n610 DVDD.t31 0.3645
R4017 DVDD.n612 DVDD.t54 0.3645
R4018 DVDD.n612 DVDD.t67 0.3645
R4019 DVDD.n614 DVDD.t29 0.3645
R4020 DVDD.n614 DVDD.t51 0.3645
R4021 DVDD.n617 DVDD.t14 0.3645
R4022 DVDD.n617 DVDD.t16 0.3645
R4023 DVDD.n618 DVDD.t41 0.3645
R4024 DVDD.n618 DVDD.t56 0.3645
R4025 DVDD.n619 DVDD.t74 0.3645
R4026 DVDD.n619 DVDD.t49 0.3645
R4027 DVDD.n620 DVDD.t35 0.3645
R4028 DVDD.n620 DVDD.t45 0.3645
R4029 DVDD.n621 DVDD.t65 0.3645
R4030 DVDD.n621 DVDD.t37 0.3645
R4031 DVDD.n622 DVDD.t39 0.3645
R4032 DVDD.n622 DVDD.t47 0.3645
R4033 DVDD.n623 DVDD.t63 0.3645
R4034 DVDD.n623 DVDD.t1 0.3645
R4035 DVDD.n257 DVDD.t24 0.3645
R4036 DVDD.n257 DVDD.t58 0.3645
R4037 DVDD.n258 DVDD.t33 0.3645
R4038 DVDD.n258 DVDD.t22 0.3645
R4039 DVDD.n259 DVDD.t43 0.3645
R4040 DVDD.n259 DVDD.t69 0.3645
R4041 DVDD.n5481 DVDD.n607 0.362381
R4042 DVDD.n5710 DVDD.n5709 0.362381
R4043 DVDD.n3915 DVDD.n3914 0.357811
R4044 DVDD.n4203 DVDD.n4201 0.357553
R4045 DVDD.n4197 DVDD.n4196 0.357321
R4046 DVDD.n3908 DVDD.n3682 0.357055
R4047 DVDD.n5456 DVDD.n645 0.35585
R4048 DVDD.n864 DVDD.n863 0.35585
R4049 DVDD.n3169 DVDD.n3163 0.355277
R4050 DVDD.n3169 DVDD.n3167 0.355277
R4051 DVDD.n233 DVDD.n215 0.355277
R4052 DVDD.n233 DVDD.n221 0.355277
R4053 DVDD.n5321 DVDD.n191 0.35501
R4054 DVDD.n5321 DVDD.n196 0.35501
R4055 DVDD.n233 DVDD.n225 0.35405
R4056 DVDD.n233 DVDD.n218 0.35405
R4057 DVDD.n5455 DVDD.n645 0.353477
R4058 DVDD.n864 DVDD.n849 0.353477
R4059 DVDD.n5321 DVDD.n188 0.353477
R4060 DVDD.n5321 DVDD.n197 0.353477
R4061 DVDD.n3169 DVDD.n3159 0.353373
R4062 DVDD.n4862 DVDD.n3169 0.353373
R4063 DVDD.n191 DVDD.n184 0.339299
R4064 DVDD.n196 DVDD.n184 0.339299
R4065 DVDD.n4863 DVDD.n3167 0.339029
R4066 DVDD.n5729 DVDD.n215 0.339029
R4067 DVDD.n5729 DVDD.n221 0.339029
R4068 DVDD.n4863 DVDD.n3163 0.339029
R4069 DVDD.n5457 DVDD.n5456 0.338454
R4070 DVDD.n863 DVDD.n862 0.338454
R4071 DVDD.n4863 DVDD.n4862 0.338164
R4072 DVDD.n4863 DVDD.n3159 0.338164
R4073 DVDD.n5457 DVDD.n5455 0.337829
R4074 DVDD.n862 DVDD.n849 0.337829
R4075 DVDD.n188 DVDD.n184 0.337829
R4076 DVDD.n197 DVDD.n184 0.337829
R4077 DVDD.n5729 DVDD.n225 0.337254
R4078 DVDD.n5729 DVDD.n218 0.337254
R4079 DVDD.n4535 DVDD.n4494 0.329604
R4080 DVDD.n5656 DVDD.n5655 0.328597
R4081 DVDD.n3899 DVDD.n3611 0.325239
R4082 DVDD.n3759 DVDD 0.312875
R4083 DVDD DVDD.n3757 0.312875
R4084 DVDD.n4118 DVDD 0.312875
R4085 DVDD.n4119 DVDD 0.312875
R4086 DVDD.n2802 DVDD.n2798 0.249007
R4087 DVDD.n2568 DVDD.n2565 0.243466
R4088 DVDD.n5523 DVDD.n5522 0.225164
R4089 DVDD.n2933 DVDD.n2932 0.2201
R4090 DVDD.n5530 DVDD.n526 0.2201
R4091 DVDD.n5531 DVDD.n5530 0.2201
R4092 DVDD.n5532 DVDD.n5531 0.2201
R4093 DVDD.n5533 DVDD.n5532 0.2201
R4094 DVDD.n5534 DVDD.n5533 0.2201
R4095 DVDD.n5536 DVDD.n5535 0.2201
R4096 DVDD.n5537 DVDD.n5536 0.2201
R4097 DVDD.n5538 DVDD.n5537 0.2201
R4098 DVDD.n5539 DVDD.n5538 0.2201
R4099 DVDD.n5540 DVDD.n5539 0.2201
R4100 DVDD.n5541 DVDD.n5540 0.2201
R4101 DVDD.n5542 DVDD.n5541 0.2201
R4102 DVDD.n5543 DVDD.n5542 0.2201
R4103 DVDD.n5544 DVDD.n5543 0.2201
R4104 DVDD.n2610 DVDD.n429 0.2201
R4105 DVDD.n5562 DVDD.n5561 0.2201
R4106 DVDD.n5561 DVDD.n5560 0.2201
R4107 DVDD.n5560 DVDD.n5559 0.2201
R4108 DVDD.n5559 DVDD.n5558 0.2201
R4109 DVDD.n5558 DVDD.n5557 0.2201
R4110 DVDD.n5556 DVDD.n5555 0.2201
R4111 DVDD.n5555 DVDD.n5554 0.2201
R4112 DVDD.n5554 DVDD.n5553 0.2201
R4113 DVDD.n5553 DVDD.n5552 0.2201
R4114 DVDD.n5552 DVDD.n5551 0.2201
R4115 DVDD.n5551 DVDD.n5550 0.2201
R4116 DVDD.n5550 DVDD.n5549 0.2201
R4117 DVDD.n5549 DVDD.n5548 0.2201
R4118 DVDD.n5548 DVDD.n5547 0.2201
R4119 DVDD.n5618 DVDD.n5617 0.2201
R4120 DVDD.n2861 DVDD.n2860 0.2201
R4121 DVDD.n2860 DVDD.n2859 0.2201
R4122 DVDD.n2859 DVDD.n2858 0.2201
R4123 DVDD.n2858 DVDD.n2857 0.2201
R4124 DVDD.n2857 DVDD.n2856 0.2201
R4125 DVDD.n2855 DVDD.n2854 0.2201
R4126 DVDD.n2854 DVDD.n2853 0.2201
R4127 DVDD.n2853 DVDD.n2852 0.2201
R4128 DVDD.n2852 DVDD.n2851 0.2201
R4129 DVDD.n2851 DVDD.n2850 0.2201
R4130 DVDD.n2850 DVDD.n2849 0.2201
R4131 DVDD.n2849 DVDD.n2848 0.2201
R4132 DVDD.n2848 DVDD.n2847 0.2201
R4133 DVDD.n2847 DVDD.n556 0.2201
R4134 DVDD.n5620 DVDD.n473 0.2201
R4135 DVDD.n2863 DVDD.n2766 0.2201
R4136 DVDD.n2830 DVDD.n2766 0.2201
R4137 DVDD.n2831 DVDD.n2830 0.2201
R4138 DVDD.n2832 DVDD.n2831 0.2201
R4139 DVDD.n2833 DVDD.n2832 0.2201
R4140 DVDD.n2835 DVDD.n2834 0.2201
R4141 DVDD.n2836 DVDD.n2835 0.2201
R4142 DVDD.n2837 DVDD.n2836 0.2201
R4143 DVDD.n2838 DVDD.n2837 0.2201
R4144 DVDD.n2839 DVDD.n2838 0.2201
R4145 DVDD.n2840 DVDD.n2839 0.2201
R4146 DVDD.n2841 DVDD.n2840 0.2201
R4147 DVDD.n2841 DVDD.n557 0.2201
R4148 DVDD.n5517 DVDD.n557 0.2201
R4149 DVDD.n4536 DVDD.n3429 0.218099
R4150 DVDD.n4697 DVDD.n3370 0.218099
R4151 DVDD.n3502 DVDD.n3485 0.218099
R4152 DVDD.n3191 DVDD.n3181 0.218099
R4153 DVDD.n240 DVDD.n239 0.217859
R4154 DVDD.n5135 DVDD.n4934 0.217859
R4155 DVDD.n3047 DVDD.n740 0.217859
R4156 DVDD.n5365 DVDD.n5364 0.217859
R4157 DVDD.n1847 DVDD.n1846 0.214786
R4158 DVDD.n1845 DVDD.n1782 0.214786
R4159 DVDD.n1844 DVDD.n1786 0.214786
R4160 DVDD.n1800 DVDD.n1787 0.214786
R4161 DVDD.n1840 DVDD.n1801 0.214786
R4162 DVDD.n1839 DVDD.n1802 0.214786
R4163 DVDD.n1838 DVDD.n1803 0.214786
R4164 DVDD.n1806 DVDD.n1804 0.214786
R4165 DVDD.n1834 DVDD.n1807 0.214786
R4166 DVDD.n1833 DVDD.n1808 0.214786
R4167 DVDD.n1832 DVDD.n1809 0.214786
R4168 DVDD.n1812 DVDD.n1810 0.214786
R4169 DVDD.n1828 DVDD.n1813 0.214786
R4170 DVDD.n1827 DVDD.n1814 0.214786
R4171 DVDD.n1826 DVDD.n1815 0.214786
R4172 DVDD.n1817 DVDD.n1816 0.214786
R4173 DVDD.n1822 DVDD.n1818 0.214786
R4174 DVDD.n1821 DVDD.n1820 0.214786
R4175 DVDD.n1819 DVDD.n1745 0.214786
R4176 DVDD.n2023 DVDD.n1746 0.214786
R4177 DVDD.n2022 DVDD.n1747 0.214786
R4178 DVDD.n2021 DVDD.n1748 0.214786
R4179 DVDD.n1750 DVDD.n1749 0.214786
R4180 DVDD.n2017 DVDD.n1751 0.214786
R4181 DVDD.n2015 DVDD.n1946 0.214786
R4182 DVDD.n1949 DVDD.n1947 0.214786
R4183 DVDD.n2011 DVDD.n1950 0.214786
R4184 DVDD.n2010 DVDD.n1951 0.214786
R4185 DVDD.n2009 DVDD.n1952 0.214786
R4186 DVDD.n1955 DVDD.n1953 0.214786
R4187 DVDD.n2005 DVDD.n1956 0.214786
R4188 DVDD.n2004 DVDD.n1957 0.214786
R4189 DVDD.n2003 DVDD.n1958 0.214786
R4190 DVDD.n2000 DVDD.n1959 0.214786
R4191 DVDD.n1999 DVDD.n1960 0.214786
R4192 DVDD.n1998 DVDD.n1961 0.214786
R4193 DVDD.n1997 DVDD.n1962 0.214786
R4194 DVDD.n1995 DVDD.n1963 0.214786
R4195 DVDD.n1966 DVDD.n1964 0.214786
R4196 DVDD.n1991 DVDD.n1967 0.214786
R4197 DVDD.n1990 DVDD.n1968 0.214786
R4198 DVDD.n1989 DVDD.n1969 0.214786
R4199 DVDD.n1972 DVDD.n1970 0.214786
R4200 DVDD.n1985 DVDD.n1973 0.214786
R4201 DVDD.n1984 DVDD.n1974 0.214786
R4202 DVDD.n1983 DVDD.n1975 0.214786
R4203 DVDD.n1979 DVDD.n1978 0.214786
R4204 DVDD.n1977 DVDD.n1583 0.214786
R4205 DVDD.n2056 DVDD.n1584 0.214786
R4206 DVDD.n1588 DVDD.n1585 0.214786
R4207 DVDD.n2052 DVDD.n1589 0.214786
R4208 DVDD.n2051 DVDD.n1590 0.214786
R4209 DVDD.n2050 DVDD.n1591 0.214786
R4210 DVDD.n1609 DVDD.n1592 0.214786
R4211 DVDD.n1696 DVDD.n1610 0.214786
R4212 DVDD.n1695 DVDD.n1611 0.214786
R4213 DVDD.n1694 DVDD.n1612 0.214786
R4214 DVDD.n1615 DVDD.n1613 0.214786
R4215 DVDD.n1690 DVDD.n1616 0.214786
R4216 DVDD.n1689 DVDD.n1617 0.214786
R4217 DVDD.n1688 DVDD.n1618 0.214786
R4218 DVDD.n1621 DVDD.n1619 0.214786
R4219 DVDD.n1684 DVDD.n1622 0.214786
R4220 DVDD.n1683 DVDD.n1623 0.214786
R4221 DVDD.n1682 DVDD.n1624 0.214786
R4222 DVDD.n1627 DVDD.n1625 0.214786
R4223 DVDD.n1678 DVDD.n1628 0.214786
R4224 DVDD.n1677 DVDD.n1629 0.214786
R4225 DVDD.n1676 DVDD.n1630 0.214786
R4226 DVDD.n1673 DVDD.n1631 0.214786
R4227 DVDD.n1672 DVDD.n1632 0.214786
R4228 DVDD.n1671 DVDD.n1633 0.214786
R4229 DVDD.n1669 DVDD.n1634 0.214786
R4230 DVDD.n1637 DVDD.n1635 0.214786
R4231 DVDD.n1665 DVDD.n1638 0.214786
R4232 DVDD.n1664 DVDD.n1639 0.214786
R4233 DVDD.n1663 DVDD.n1640 0.214786
R4234 DVDD.n1643 DVDD.n1641 0.214786
R4235 DVDD.n1659 DVDD.n1644 0.214786
R4236 DVDD.n1658 DVDD.n1645 0.214786
R4237 DVDD.n1657 DVDD.n1646 0.214786
R4238 DVDD.n1648 DVDD.n1647 0.214786
R4239 DVDD.n1653 DVDD.n1649 0.214786
R4240 DVDD.n1652 DVDD.n1650 0.214786
R4241 DVDD.n1783 DVDD.n1779 0.214786
R4242 DVDD.n1778 DVDD.n1410 0.214786
R4243 DVDD.n2204 DVDD.n1411 0.214786
R4244 DVDD.n2203 DVDD.n1412 0.214786
R4245 DVDD.n2202 DVDD.n1413 0.214786
R4246 DVDD.n1416 DVDD.n1414 0.214786
R4247 DVDD.n2198 DVDD.n1417 0.214786
R4248 DVDD.n2197 DVDD.n1418 0.214786
R4249 DVDD.n2196 DVDD.n1419 0.214786
R4250 DVDD.n1422 DVDD.n1420 0.214786
R4251 DVDD.n2192 DVDD.n1423 0.214786
R4252 DVDD.n2191 DVDD.n1424 0.214786
R4253 DVDD.n2190 DVDD.n1425 0.214786
R4254 DVDD.n1428 DVDD.n1426 0.214786
R4255 DVDD.n2186 DVDD.n1429 0.214786
R4256 DVDD.n2185 DVDD.n1430 0.214786
R4257 DVDD.n2184 DVDD.n1431 0.214786
R4258 DVDD.n2182 DVDD.n1432 0.214786
R4259 DVDD.n2181 DVDD.n1433 0.214786
R4260 DVDD.n2180 DVDD.n1434 0.214786
R4261 DVDD.n1448 DVDD.n1435 0.214786
R4262 DVDD.n2176 DVDD.n1449 0.214786
R4263 DVDD.n2175 DVDD.n1450 0.214786
R4264 DVDD.n2174 DVDD.n1451 0.214786
R4265 DVDD.n2170 DVDD.n1454 0.214786
R4266 DVDD.n2169 DVDD.n1455 0.214786
R4267 DVDD.n2168 DVDD.n1456 0.214786
R4268 DVDD.n1459 DVDD.n1457 0.214786
R4269 DVDD.n2164 DVDD.n1460 0.214786
R4270 DVDD.n2163 DVDD.n1461 0.214786
R4271 DVDD.n2162 DVDD.n1462 0.214786
R4272 DVDD.n1465 DVDD.n1463 0.214786
R4273 DVDD.n2158 DVDD.n1466 0.214786
R4274 DVDD.n2157 DVDD.n1467 0.214786
R4275 DVDD.n2156 DVDD.n1468 0.214786
R4276 DVDD.n1565 DVDD.n1469 0.214786
R4277 DVDD.n2150 DVDD.n1566 0.214786
R4278 DVDD.n2149 DVDD.n1567 0.214786
R4279 DVDD.n1570 DVDD.n1568 0.214786
R4280 DVDD.n2145 DVDD.n1571 0.214786
R4281 DVDD.n2144 DVDD.n1572 0.214786
R4282 DVDD.n2143 DVDD.n1573 0.214786
R4283 DVDD.n1576 DVDD.n1574 0.214786
R4284 DVDD.n2139 DVDD.n1577 0.214786
R4285 DVDD.n2138 DVDD.n1578 0.214786
R4286 DVDD.n2137 DVDD.n1579 0.214786
R4287 DVDD.n1581 DVDD.n1580 0.214786
R4288 DVDD.n2133 DVDD.n1582 0.214786
R4289 DVDD.n2131 DVDD.n2058 0.214786
R4290 DVDD.n2061 DVDD.n2059 0.214786
R4291 DVDD.n2127 DVDD.n2062 0.214786
R4292 DVDD.n2126 DVDD.n2063 0.214786
R4293 DVDD.n2125 DVDD.n2064 0.214786
R4294 DVDD.n2124 DVDD.n2065 0.214786
R4295 DVDD.n2123 DVDD.n2066 0.214786
R4296 DVDD.n2080 DVDD.n2067 0.214786
R4297 DVDD.n2119 DVDD.n2081 0.214786
R4298 DVDD.n2118 DVDD.n2082 0.214786
R4299 DVDD.n2117 DVDD.n2083 0.214786
R4300 DVDD.n2086 DVDD.n2084 0.214786
R4301 DVDD.n2113 DVDD.n2087 0.214786
R4302 DVDD.n2112 DVDD.n2088 0.214786
R4303 DVDD.n2111 DVDD.n2089 0.214786
R4304 DVDD.n2092 DVDD.n2090 0.214786
R4305 DVDD.n2107 DVDD.n2093 0.214786
R4306 DVDD.n2106 DVDD.n2094 0.214786
R4307 DVDD.n2105 DVDD.n2095 0.214786
R4308 DVDD.n2098 DVDD.n2096 0.214786
R4309 DVDD.n2101 DVDD.n2100 0.214786
R4310 DVDD.n2099 DVDD.n1369 0.214786
R4311 DVDD.n2238 DVDD.n1368 0.214786
R4312 DVDD.n2240 DVDD.n2239 0.214786
R4313 DVDD.n2275 DVDD.n2242 0.214786
R4314 DVDD.n2274 DVDD.n2243 0.214786
R4315 DVDD.n2273 DVDD.n2244 0.214786
R4316 DVDD.n2247 DVDD.n2245 0.214786
R4317 DVDD.n2269 DVDD.n2248 0.214786
R4318 DVDD.n2268 DVDD.n2249 0.214786
R4319 DVDD.n2267 DVDD.n2250 0.214786
R4320 DVDD.n2253 DVDD.n2251 0.214786
R4321 DVDD.n2263 DVDD.n2254 0.214786
R4322 DVDD.n2262 DVDD.n2255 0.214786
R4323 DVDD.n2261 DVDD.n2256 0.214786
R4324 DVDD.n2258 DVDD.n2257 0.214786
R4325 DVDD.n1852 DVDD.n1851 0.214786
R4326 DVDD.n1850 DVDD.n1141 0.214786
R4327 DVDD.n2424 DVDD.n1142 0.214786
R4328 DVDD.n2423 DVDD.n1143 0.214786
R4329 DVDD.n2422 DVDD.n1144 0.214786
R4330 DVDD.n1147 DVDD.n1145 0.214786
R4331 DVDD.n2418 DVDD.n1148 0.214786
R4332 DVDD.n2417 DVDD.n1149 0.214786
R4333 DVDD.n2416 DVDD.n1150 0.214786
R4334 DVDD.n1153 DVDD.n1151 0.214786
R4335 DVDD.n2412 DVDD.n1154 0.214786
R4336 DVDD.n2411 DVDD.n1155 0.214786
R4337 DVDD.n2410 DVDD.n1156 0.214786
R4338 DVDD.n1159 DVDD.n1157 0.214786
R4339 DVDD.n2406 DVDD.n1160 0.214786
R4340 DVDD.n2405 DVDD.n1161 0.214786
R4341 DVDD.n2404 DVDD.n1162 0.214786
R4342 DVDD.n2402 DVDD.n1163 0.214786
R4343 DVDD.n2401 DVDD.n1164 0.214786
R4344 DVDD.n2400 DVDD.n1165 0.214786
R4345 DVDD.n2399 DVDD.n1166 0.214786
R4346 DVDD.n1169 DVDD.n1167 0.214786
R4347 DVDD.n2395 DVDD.n1170 0.214786
R4348 DVDD.n2394 DVDD.n1171 0.214786
R4349 DVDD.n2392 DVDD.n1174 0.214786
R4350 DVDD.n1178 DVDD.n1175 0.214786
R4351 DVDD.n2388 DVDD.n1179 0.214786
R4352 DVDD.n2387 DVDD.n1180 0.214786
R4353 DVDD.n2386 DVDD.n1181 0.214786
R4354 DVDD.n1184 DVDD.n1182 0.214786
R4355 DVDD.n2382 DVDD.n1185 0.214786
R4356 DVDD.n2381 DVDD.n1186 0.214786
R4357 DVDD.n2380 DVDD.n1187 0.214786
R4358 DVDD.n1190 DVDD.n1188 0.214786
R4359 DVDD.n2376 DVDD.n1191 0.214786
R4360 DVDD.n2375 DVDD.n1192 0.214786
R4361 DVDD.n1274 DVDD.n1193 0.214786
R4362 DVDD.n2367 DVDD.n1275 0.214786
R4363 DVDD.n2366 DVDD.n1276 0.214786
R4364 DVDD.n2365 DVDD.n1277 0.214786
R4365 DVDD.n1280 DVDD.n1278 0.214786
R4366 DVDD.n2361 DVDD.n1281 0.214786
R4367 DVDD.n2360 DVDD.n1282 0.214786
R4368 DVDD.n2359 DVDD.n1283 0.214786
R4369 DVDD.n1286 DVDD.n1284 0.214786
R4370 DVDD.n2355 DVDD.n1287 0.214786
R4371 DVDD.n2354 DVDD.n1288 0.214786
R4372 DVDD.n2353 DVDD.n2352 0.214786
R4373 DVDD.n2490 DVDD.n1066 0.214786
R4374 DVDD.n2489 DVDD.n1067 0.214786
R4375 DVDD.n2488 DVDD.n1068 0.214786
R4376 DVDD.n2485 DVDD.n1069 0.214786
R4377 DVDD.n2484 DVDD.n1070 0.214786
R4378 DVDD.n2483 DVDD.n1071 0.214786
R4379 DVDD.n2482 DVDD.n1072 0.214786
R4380 DVDD.n2481 DVDD.n1073 0.214786
R4381 DVDD.n1076 DVDD.n1074 0.214786
R4382 DVDD.n2477 DVDD.n1077 0.214786
R4383 DVDD.n2476 DVDD.n1078 0.214786
R4384 DVDD.n2475 DVDD.n1079 0.214786
R4385 DVDD.n1082 DVDD.n1080 0.214786
R4386 DVDD.n2471 DVDD.n1083 0.214786
R4387 DVDD.n2470 DVDD.n1084 0.214786
R4388 DVDD.n2469 DVDD.n1085 0.214786
R4389 DVDD.n1088 DVDD.n1086 0.214786
R4390 DVDD.n2465 DVDD.n1089 0.214786
R4391 DVDD.n2464 DVDD.n1090 0.214786
R4392 DVDD.n2463 DVDD.n1091 0.214786
R4393 DVDD.n1094 DVDD.n1092 0.214786
R4394 DVDD.n2459 DVDD.n1095 0.214786
R4395 DVDD.n2458 DVDD.n1096 0.214786
R4396 DVDD.n1331 DVDD.n1097 0.214786
R4397 DVDD.n1366 DVDD.n1365 0.214786
R4398 DVDD.n1364 DVDD.n1332 0.214786
R4399 DVDD.n1335 DVDD.n1333 0.214786
R4400 DVDD.n1360 DVDD.n1336 0.214786
R4401 DVDD.n1359 DVDD.n1337 0.214786
R4402 DVDD.n1358 DVDD.n1338 0.214786
R4403 DVDD.n1341 DVDD.n1339 0.214786
R4404 DVDD.n1354 DVDD.n1342 0.214786
R4405 DVDD.n1353 DVDD.n1343 0.214786
R4406 DVDD.n1352 DVDD.n1344 0.214786
R4407 DVDD.n1346 DVDD.n1345 0.214786
R4408 DVDD.n1348 DVDD.n1347 0.214786
R4409 DVDD.n2315 DVDD.n1320 0.214786
R4410 DVDD.n2313 DVDD.n1322 0.214786
R4411 DVDD.n2281 DVDD.n1323 0.214786
R4412 DVDD.n2309 DVDD.n2282 0.214786
R4413 DVDD.n2308 DVDD.n2283 0.214786
R4414 DVDD.n2307 DVDD.n2284 0.214786
R4415 DVDD.n2287 DVDD.n2285 0.214786
R4416 DVDD.n2303 DVDD.n2288 0.214786
R4417 DVDD.n2302 DVDD.n2289 0.214786
R4418 DVDD.n2301 DVDD.n2290 0.214786
R4419 DVDD.n2292 DVDD.n2291 0.214786
R4420 DVDD.n2297 DVDD.n2293 0.214786
R4421 DVDD.n2296 DVDD.n2294 0.214786
R4422 DVDD.n1860 DVDD.n1859 0.214786
R4423 DVDD.n1861 DVDD.n1772 0.214786
R4424 DVDD.n1863 DVDD.n1862 0.214786
R4425 DVDD.n1864 DVDD.n1771 0.214786
R4426 DVDD.n1868 DVDD.n1867 0.214786
R4427 DVDD.n1869 DVDD.n1770 0.214786
R4428 DVDD.n1871 DVDD.n1870 0.214786
R4429 DVDD.n1768 DVDD.n1767 0.214786
R4430 DVDD.n1876 DVDD.n1875 0.214786
R4431 DVDD.n1877 DVDD.n1766 0.214786
R4432 DVDD.n1879 DVDD.n1878 0.214786
R4433 DVDD.n1764 DVDD.n1763 0.214786
R4434 DVDD.n1884 DVDD.n1883 0.214786
R4435 DVDD.n1885 DVDD.n1762 0.214786
R4436 DVDD.n1887 DVDD.n1886 0.214786
R4437 DVDD.n1760 DVDD.n1759 0.214786
R4438 DVDD.n1892 DVDD.n1891 0.214786
R4439 DVDD.n1893 DVDD.n1758 0.214786
R4440 DVDD.n1895 DVDD.n1894 0.214786
R4441 DVDD.n1896 DVDD.n1757 0.214786
R4442 DVDD.n1900 DVDD.n1899 0.214786
R4443 DVDD.n1901 DVDD.n1756 0.214786
R4444 DVDD.n1903 DVDD.n1902 0.214786
R4445 DVDD.n1904 DVDD.n1752 0.214786
R4446 DVDD.n1941 DVDD.n1940 0.214786
R4447 DVDD.n1754 DVDD.n1753 0.214786
R4448 DVDD.n1936 DVDD.n1908 0.214786
R4449 DVDD.n1935 DVDD.n1909 0.214786
R4450 DVDD.n1934 DVDD.n1910 0.214786
R4451 DVDD.n1913 DVDD.n1911 0.214786
R4452 DVDD.n1930 DVDD.n1914 0.214786
R4453 DVDD.n1929 DVDD.n1915 0.214786
R4454 DVDD.n1928 DVDD.n1916 0.214786
R4455 DVDD.n1918 DVDD.n1917 0.214786
R4456 DVDD.n1924 DVDD.n1919 0.214786
R4457 DVDD.n1923 DVDD.n1921 0.214786
R4458 DVDD.n1920 DVDD.n1044 0.214786
R4459 DVDD.n2509 DVDD.n1045 0.214786
R4460 DVDD.n2508 DVDD.n1046 0.214786
R4461 DVDD.n2507 DVDD.n1047 0.214786
R4462 DVDD.n1050 DVDD.n1048 0.214786
R4463 DVDD.n2503 DVDD.n1051 0.214786
R4464 DVDD.n2502 DVDD.n1052 0.214786
R4465 DVDD.n2501 DVDD.n1053 0.214786
R4466 DVDD.n1056 DVDD.n1054 0.214786
R4467 DVDD.n2497 DVDD.n1057 0.214786
R4468 DVDD.n2496 DVDD.n1058 0.214786
R4469 DVDD.n2495 DVDD.n1059 0.214786
R4470 DVDD.n2349 DVDD.n2348 0.214786
R4471 DVDD.n2347 DVDD.n1290 0.214786
R4472 DVDD.n1292 DVDD.n1291 0.214786
R4473 DVDD.n2343 DVDD.n1293 0.214786
R4474 DVDD.n2342 DVDD.n1294 0.214786
R4475 DVDD.n2341 DVDD.n1295 0.214786
R4476 DVDD.n2340 DVDD.n1296 0.214786
R4477 DVDD.n2339 DVDD.n1297 0.214786
R4478 DVDD.n1300 DVDD.n1298 0.214786
R4479 DVDD.n2335 DVDD.n1301 0.214786
R4480 DVDD.n2334 DVDD.n1302 0.214786
R4481 DVDD.n2333 DVDD.n1303 0.214786
R4482 DVDD.n1306 DVDD.n1304 0.214786
R4483 DVDD.n2329 DVDD.n1307 0.214786
R4484 DVDD.n2328 DVDD.n1308 0.214786
R4485 DVDD.n2327 DVDD.n1309 0.214786
R4486 DVDD.n1312 DVDD.n1310 0.214786
R4487 DVDD.n2323 DVDD.n1313 0.214786
R4488 DVDD.n2322 DVDD.n1314 0.214786
R4489 DVDD.n2321 DVDD.n1315 0.214786
R4490 DVDD.n1317 DVDD.n1316 0.214786
R4491 DVDD.n2317 DVDD.n1318 0.214786
R4492 DVDD.n2316 DVDD.n1319 0.214786
R4493 DVDD.n2315 DVDD.n988 0.214786
R4494 DVDD.n2298 DVDD.n2297 0.214786
R4495 DVDD.n2299 DVDD.n2291 0.214786
R4496 DVDD.n2301 DVDD.n2300 0.214786
R4497 DVDD.n2302 DVDD.n2286 0.214786
R4498 DVDD.n2304 DVDD.n2303 0.214786
R4499 DVDD.n2305 DVDD.n2285 0.214786
R4500 DVDD.n2307 DVDD.n2306 0.214786
R4501 DVDD.n2308 DVDD.n2280 0.214786
R4502 DVDD.n2310 DVDD.n2309 0.214786
R4503 DVDD.n2311 DVDD.n1323 0.214786
R4504 DVDD.n2313 DVDD.n2312 0.214786
R4505 DVDD.n1859 DVDD.n1858 0.214786
R4506 DVDD.n1772 DVDD.n448 0.214786
R4507 DVDD.n1863 DVDD.n454 0.214786
R4508 DVDD.n1865 DVDD.n1864 0.214786
R4509 DVDD.n1867 DVDD.n1866 0.214786
R4510 DVDD.n1770 DVDD.n1769 0.214786
R4511 DVDD.n1872 DVDD.n1871 0.214786
R4512 DVDD.n1873 DVDD.n1768 0.214786
R4513 DVDD.n1875 DVDD.n1874 0.214786
R4514 DVDD.n1766 DVDD.n1765 0.214786
R4515 DVDD.n1880 DVDD.n1879 0.214786
R4516 DVDD.n1881 DVDD.n1764 0.214786
R4517 DVDD.n1883 DVDD.n1882 0.214786
R4518 DVDD.n1762 DVDD.n1761 0.214786
R4519 DVDD.n1888 DVDD.n1887 0.214786
R4520 DVDD.n1889 DVDD.n1760 0.214786
R4521 DVDD.n1891 DVDD.n1890 0.214786
R4522 DVDD.n1758 DVDD.n952 0.214786
R4523 DVDD.n1895 DVDD.n959 0.214786
R4524 DVDD.n1896 DVDD.n972 0.214786
R4525 DVDD.n1899 DVDD.n1898 0.214786
R4526 DVDD.n1897 DVDD.n1756 0.214786
R4527 DVDD.n1903 DVDD.n1755 0.214786
R4528 DVDD.n1905 DVDD.n1904 0.214786
R4529 DVDD.n1940 DVDD.n1939 0.214786
R4530 DVDD.n1938 DVDD.n1754 0.214786
R4531 DVDD.n1937 DVDD.n1936 0.214786
R4532 DVDD.n1935 DVDD.n1907 0.214786
R4533 DVDD.n1934 DVDD.n1933 0.214786
R4534 DVDD.n1932 DVDD.n1911 0.214786
R4535 DVDD.n1931 DVDD.n1930 0.214786
R4536 DVDD.n1929 DVDD.n1912 0.214786
R4537 DVDD.n1928 DVDD.n1927 0.214786
R4538 DVDD.n1926 DVDD.n1917 0.214786
R4539 DVDD.n1925 DVDD.n1924 0.214786
R4540 DVDD.n1923 DVDD.n1922 0.214786
R4541 DVDD.n1044 DVDD.n1018 0.214786
R4542 DVDD.n2510 DVDD.n2509 0.214786
R4543 DVDD.n2508 DVDD.n1043 0.214786
R4544 DVDD.n2507 DVDD.n2506 0.214786
R4545 DVDD.n2505 DVDD.n1048 0.214786
R4546 DVDD.n2504 DVDD.n2503 0.214786
R4547 DVDD.n2502 DVDD.n1049 0.214786
R4548 DVDD.n2501 DVDD.n2500 0.214786
R4549 DVDD.n2499 DVDD.n1054 0.214786
R4550 DVDD.n2498 DVDD.n2497 0.214786
R4551 DVDD.n2496 DVDD.n1055 0.214786
R4552 DVDD.n2495 DVDD.n2494 0.214786
R4553 DVDD.n2348 DVDD.n1061 0.214786
R4554 DVDD.n2347 DVDD.n2346 0.214786
R4555 DVDD.n2345 DVDD.n1291 0.214786
R4556 DVDD.n2344 DVDD.n2343 0.214786
R4557 DVDD.n2342 DVDD.n413 0.214786
R4558 DVDD.n2341 DVDD.n420 0.214786
R4559 DVDD.n2340 DVDD.n436 0.214786
R4560 DVDD.n2339 DVDD.n2338 0.214786
R4561 DVDD.n2337 DVDD.n1298 0.214786
R4562 DVDD.n2336 DVDD.n2335 0.214786
R4563 DVDD.n2334 DVDD.n1299 0.214786
R4564 DVDD.n2333 DVDD.n2332 0.214786
R4565 DVDD.n2331 DVDD.n1304 0.214786
R4566 DVDD.n2330 DVDD.n2329 0.214786
R4567 DVDD.n2328 DVDD.n1305 0.214786
R4568 DVDD.n2327 DVDD.n2326 0.214786
R4569 DVDD.n2325 DVDD.n1310 0.214786
R4570 DVDD.n2324 DVDD.n2323 0.214786
R4571 DVDD.n2322 DVDD.n1311 0.214786
R4572 DVDD.n2321 DVDD.n2320 0.214786
R4573 DVDD.n2319 DVDD.n1316 0.214786
R4574 DVDD.n2318 DVDD.n2317 0.214786
R4575 DVDD.n2316 DVDD.n982 0.214786
R4576 DVDD.n1100 DVDD.n1097 0.214786
R4577 DVDD.n1365 DVDD.n1324 0.214786
R4578 DVDD.n1364 DVDD.n1363 0.214786
R4579 DVDD.n1362 DVDD.n1333 0.214786
R4580 DVDD.n1361 DVDD.n1360 0.214786
R4581 DVDD.n1359 DVDD.n1334 0.214786
R4582 DVDD.n1358 DVDD.n1357 0.214786
R4583 DVDD.n1356 DVDD.n1339 0.214786
R4584 DVDD.n1355 DVDD.n1354 0.214786
R4585 DVDD.n1353 DVDD.n1340 0.214786
R4586 DVDD.n1352 DVDD.n1351 0.214786
R4587 DVDD.n1350 DVDD.n1345 0.214786
R4588 DVDD.n2458 DVDD.n2457 0.214786
R4589 DVDD.n2460 DVDD.n2459 0.214786
R4590 DVDD.n2461 DVDD.n1092 0.214786
R4591 DVDD.n2463 DVDD.n2462 0.214786
R4592 DVDD.n2464 DVDD.n1087 0.214786
R4593 DVDD.n2466 DVDD.n2465 0.214786
R4594 DVDD.n2467 DVDD.n1086 0.214786
R4595 DVDD.n2469 DVDD.n2468 0.214786
R4596 DVDD.n2470 DVDD.n1081 0.214786
R4597 DVDD.n2472 DVDD.n2471 0.214786
R4598 DVDD.n2473 DVDD.n1080 0.214786
R4599 DVDD.n2475 DVDD.n2474 0.214786
R4600 DVDD.n2476 DVDD.n1075 0.214786
R4601 DVDD.n2478 DVDD.n2477 0.214786
R4602 DVDD.n2479 DVDD.n1074 0.214786
R4603 DVDD.n2481 DVDD.n2480 0.214786
R4604 DVDD.n2482 DVDD.n401 0.214786
R4605 DVDD.n2483 DVDD.n388 0.214786
R4606 DVDD.n2484 DVDD.n383 0.214786
R4607 DVDD.n2486 DVDD.n2485 0.214786
R4608 DVDD.n2488 DVDD.n2487 0.214786
R4609 DVDD.n2489 DVDD.n1064 0.214786
R4610 DVDD.n2491 DVDD.n2490 0.214786
R4611 DVDD.n2353 DVDD.n1063 0.214786
R4612 DVDD.n2354 DVDD.n1285 0.214786
R4613 DVDD.n2356 DVDD.n2355 0.214786
R4614 DVDD.n2357 DVDD.n1284 0.214786
R4615 DVDD.n2359 DVDD.n2358 0.214786
R4616 DVDD.n2360 DVDD.n1279 0.214786
R4617 DVDD.n2362 DVDD.n2361 0.214786
R4618 DVDD.n2363 DVDD.n1278 0.214786
R4619 DVDD.n2365 DVDD.n2364 0.214786
R4620 DVDD.n2366 DVDD.n1273 0.214786
R4621 DVDD.n2368 DVDD.n2367 0.214786
R4622 DVDD.n1222 DVDD.n1193 0.214786
R4623 DVDD.n2375 DVDD.n2374 0.214786
R4624 DVDD.n2377 DVDD.n2376 0.214786
R4625 DVDD.n2378 DVDD.n1188 0.214786
R4626 DVDD.n2380 DVDD.n2379 0.214786
R4627 DVDD.n2381 DVDD.n1183 0.214786
R4628 DVDD.n2383 DVDD.n2382 0.214786
R4629 DVDD.n2384 DVDD.n1182 0.214786
R4630 DVDD.n2386 DVDD.n2385 0.214786
R4631 DVDD.n2387 DVDD.n1177 0.214786
R4632 DVDD.n2389 DVDD.n2388 0.214786
R4633 DVDD.n2390 DVDD.n1175 0.214786
R4634 DVDD.n2392 DVDD.n2391 0.214786
R4635 DVDD.n2394 DVDD.n1168 0.214786
R4636 DVDD.n2396 DVDD.n2395 0.214786
R4637 DVDD.n2397 DVDD.n1167 0.214786
R4638 DVDD.n2399 DVDD.n2398 0.214786
R4639 DVDD.n2400 DVDD.n940 0.214786
R4640 DVDD.n2401 DVDD.n927 0.214786
R4641 DVDD.n2402 DVDD.n922 0.214786
R4642 DVDD.n2404 DVDD.n2403 0.214786
R4643 DVDD.n2405 DVDD.n1158 0.214786
R4644 DVDD.n2407 DVDD.n2406 0.214786
R4645 DVDD.n2408 DVDD.n1157 0.214786
R4646 DVDD.n2410 DVDD.n2409 0.214786
R4647 DVDD.n2411 DVDD.n1152 0.214786
R4648 DVDD.n2413 DVDD.n2412 0.214786
R4649 DVDD.n2414 DVDD.n1151 0.214786
R4650 DVDD.n2416 DVDD.n2415 0.214786
R4651 DVDD.n2417 DVDD.n1146 0.214786
R4652 DVDD.n2419 DVDD.n2418 0.214786
R4653 DVDD.n2420 DVDD.n1145 0.214786
R4654 DVDD.n2422 DVDD.n2421 0.214786
R4655 DVDD.n2423 DVDD.n1140 0.214786
R4656 DVDD.n2425 DVDD.n2424 0.214786
R4657 DVDD.n1141 DVDD.n1128 0.214786
R4658 DVDD.n1851 DVDD.n1123 0.214786
R4659 DVDD.n2239 DVDD.n1326 0.214786
R4660 DVDD.n2276 DVDD.n2275 0.214786
R4661 DVDD.n2274 DVDD.n1327 0.214786
R4662 DVDD.n2273 DVDD.n2272 0.214786
R4663 DVDD.n2271 DVDD.n2245 0.214786
R4664 DVDD.n2270 DVDD.n2269 0.214786
R4665 DVDD.n2268 DVDD.n2246 0.214786
R4666 DVDD.n2267 DVDD.n2266 0.214786
R4667 DVDD.n2265 DVDD.n2251 0.214786
R4668 DVDD.n2264 DVDD.n2263 0.214786
R4669 DVDD.n2262 DVDD.n2252 0.214786
R4670 DVDD.n2261 DVDD.n2260 0.214786
R4671 DVDD.n2238 DVDD.n2237 0.214786
R4672 DVDD.n2097 DVDD.n1369 0.214786
R4673 DVDD.n2102 DVDD.n2101 0.214786
R4674 DVDD.n2103 DVDD.n2096 0.214786
R4675 DVDD.n2105 DVDD.n2104 0.214786
R4676 DVDD.n2106 DVDD.n2091 0.214786
R4677 DVDD.n2108 DVDD.n2107 0.214786
R4678 DVDD.n2109 DVDD.n2090 0.214786
R4679 DVDD.n2111 DVDD.n2110 0.214786
R4680 DVDD.n2112 DVDD.n2085 0.214786
R4681 DVDD.n2114 DVDD.n2113 0.214786
R4682 DVDD.n2115 DVDD.n2084 0.214786
R4683 DVDD.n2117 DVDD.n2116 0.214786
R4684 DVDD.n2118 DVDD.n2079 0.214786
R4685 DVDD.n2120 DVDD.n2119 0.214786
R4686 DVDD.n2121 DVDD.n2067 0.214786
R4687 DVDD.n2123 DVDD.n2122 0.214786
R4688 DVDD.n2124 DVDD.n368 0.214786
R4689 DVDD.n2125 DVDD.n362 0.214786
R4690 DVDD.n2126 DVDD.n2060 0.214786
R4691 DVDD.n2128 DVDD.n2127 0.214786
R4692 DVDD.n2129 DVDD.n2059 0.214786
R4693 DVDD.n2131 DVDD.n2130 0.214786
R4694 DVDD.n2134 DVDD.n2133 0.214786
R4695 DVDD.n2135 DVDD.n1580 0.214786
R4696 DVDD.n2137 DVDD.n2136 0.214786
R4697 DVDD.n2138 DVDD.n1575 0.214786
R4698 DVDD.n2140 DVDD.n2139 0.214786
R4699 DVDD.n2141 DVDD.n1574 0.214786
R4700 DVDD.n2143 DVDD.n2142 0.214786
R4701 DVDD.n2144 DVDD.n1569 0.214786
R4702 DVDD.n2146 DVDD.n2145 0.214786
R4703 DVDD.n2147 DVDD.n1568 0.214786
R4704 DVDD.n2149 DVDD.n2148 0.214786
R4705 DVDD.n2151 DVDD.n2150 0.214786
R4706 DVDD.n1481 DVDD.n1469 0.214786
R4707 DVDD.n2156 DVDD.n2155 0.214786
R4708 DVDD.n2157 DVDD.n1464 0.214786
R4709 DVDD.n2159 DVDD.n2158 0.214786
R4710 DVDD.n2160 DVDD.n1463 0.214786
R4711 DVDD.n2162 DVDD.n2161 0.214786
R4712 DVDD.n2163 DVDD.n1458 0.214786
R4713 DVDD.n2165 DVDD.n2164 0.214786
R4714 DVDD.n2166 DVDD.n1457 0.214786
R4715 DVDD.n2168 DVDD.n2167 0.214786
R4716 DVDD.n2169 DVDD.n1453 0.214786
R4717 DVDD.n2171 DVDD.n2170 0.214786
R4718 DVDD.n2174 DVDD.n2173 0.214786
R4719 DVDD.n2175 DVDD.n1447 0.214786
R4720 DVDD.n2177 DVDD.n2176 0.214786
R4721 DVDD.n2178 DVDD.n1435 0.214786
R4722 DVDD.n2180 DVDD.n2179 0.214786
R4723 DVDD.n2181 DVDD.n907 0.214786
R4724 DVDD.n2182 DVDD.n901 0.214786
R4725 DVDD.n2184 DVDD.n2183 0.214786
R4726 DVDD.n2185 DVDD.n1427 0.214786
R4727 DVDD.n2187 DVDD.n2186 0.214786
R4728 DVDD.n2188 DVDD.n1426 0.214786
R4729 DVDD.n2190 DVDD.n2189 0.214786
R4730 DVDD.n2191 DVDD.n1421 0.214786
R4731 DVDD.n2193 DVDD.n2192 0.214786
R4732 DVDD.n2194 DVDD.n1420 0.214786
R4733 DVDD.n2196 DVDD.n2195 0.214786
R4734 DVDD.n2197 DVDD.n1415 0.214786
R4735 DVDD.n2199 DVDD.n2198 0.214786
R4736 DVDD.n2200 DVDD.n1414 0.214786
R4737 DVDD.n2202 DVDD.n2201 0.214786
R4738 DVDD.n2203 DVDD.n1409 0.214786
R4739 DVDD.n2205 DVDD.n2204 0.214786
R4740 DVDD.n1410 DVDD.n1398 0.214786
R4741 DVDD.n1783 DVDD.n1393 0.214786
R4742 DVDD.n1671 DVDD.n603 0.214786
R4743 DVDD.n1669 DVDD.n1668 0.214786
R4744 DVDD.n1667 DVDD.n1635 0.214786
R4745 DVDD.n1666 DVDD.n1665 0.214786
R4746 DVDD.n1664 DVDD.n1636 0.214786
R4747 DVDD.n1663 DVDD.n1662 0.214786
R4748 DVDD.n1661 DVDD.n1641 0.214786
R4749 DVDD.n1660 DVDD.n1659 0.214786
R4750 DVDD.n1658 DVDD.n1642 0.214786
R4751 DVDD.n1657 DVDD.n1656 0.214786
R4752 DVDD.n1655 DVDD.n1647 0.214786
R4753 DVDD.n1654 DVDD.n1653 0.214786
R4754 DVDD.n1672 DVDD.n581 0.214786
R4755 DVDD.n1674 DVDD.n1673 0.214786
R4756 DVDD.n1676 DVDD.n1675 0.214786
R4757 DVDD.n1677 DVDD.n1626 0.214786
R4758 DVDD.n1679 DVDD.n1678 0.214786
R4759 DVDD.n1680 DVDD.n1625 0.214786
R4760 DVDD.n1682 DVDD.n1681 0.214786
R4761 DVDD.n1683 DVDD.n1620 0.214786
R4762 DVDD.n1685 DVDD.n1684 0.214786
R4763 DVDD.n1686 DVDD.n1619 0.214786
R4764 DVDD.n1688 DVDD.n1687 0.214786
R4765 DVDD.n1689 DVDD.n1614 0.214786
R4766 DVDD.n1691 DVDD.n1690 0.214786
R4767 DVDD.n1692 DVDD.n1613 0.214786
R4768 DVDD.n1694 DVDD.n1693 0.214786
R4769 DVDD.n1695 DVDD.n1608 0.214786
R4770 DVDD.n1697 DVDD.n1696 0.214786
R4771 DVDD.n1599 DVDD.n1592 0.214786
R4772 DVDD.n2050 DVDD.n2049 0.214786
R4773 DVDD.n2051 DVDD.n1587 0.214786
R4774 DVDD.n2053 DVDD.n2052 0.214786
R4775 DVDD.n2054 DVDD.n1585 0.214786
R4776 DVDD.n2056 DVDD.n2055 0.214786
R4777 DVDD.n1980 DVDD.n1583 0.214786
R4778 DVDD.n1981 DVDD.n1979 0.214786
R4779 DVDD.n1983 DVDD.n1982 0.214786
R4780 DVDD.n1984 DVDD.n1971 0.214786
R4781 DVDD.n1986 DVDD.n1985 0.214786
R4782 DVDD.n1987 DVDD.n1970 0.214786
R4783 DVDD.n1989 DVDD.n1988 0.214786
R4784 DVDD.n1990 DVDD.n1965 0.214786
R4785 DVDD.n1992 DVDD.n1991 0.214786
R4786 DVDD.n1993 DVDD.n1964 0.214786
R4787 DVDD.n1995 DVDD.n1994 0.214786
R4788 DVDD.n1997 DVDD.n1996 0.214786
R4789 DVDD.n1998 DVDD.n326 0.214786
R4790 DVDD.n1999 DVDD.n314 0.214786
R4791 DVDD.n2001 DVDD.n2000 0.214786
R4792 DVDD.n2003 DVDD.n2002 0.214786
R4793 DVDD.n2004 DVDD.n1954 0.214786
R4794 DVDD.n2006 DVDD.n2005 0.214786
R4795 DVDD.n2007 DVDD.n1953 0.214786
R4796 DVDD.n2009 DVDD.n2008 0.214786
R4797 DVDD.n2010 DVDD.n1948 0.214786
R4798 DVDD.n2012 DVDD.n2011 0.214786
R4799 DVDD.n2013 DVDD.n1947 0.214786
R4800 DVDD.n2015 DVDD.n2014 0.214786
R4801 DVDD.n2018 DVDD.n2017 0.214786
R4802 DVDD.n2019 DVDD.n1749 0.214786
R4803 DVDD.n2021 DVDD.n2020 0.214786
R4804 DVDD.n2022 DVDD.n1744 0.214786
R4805 DVDD.n2024 DVDD.n2023 0.214786
R4806 DVDD.n1745 DVDD.n1723 0.214786
R4807 DVDD.n1821 DVDD.n1717 0.214786
R4808 DVDD.n1823 DVDD.n1822 0.214786
R4809 DVDD.n1824 DVDD.n1816 0.214786
R4810 DVDD.n1826 DVDD.n1825 0.214786
R4811 DVDD.n1827 DVDD.n1811 0.214786
R4812 DVDD.n1829 DVDD.n1828 0.214786
R4813 DVDD.n1830 DVDD.n1810 0.214786
R4814 DVDD.n1832 DVDD.n1831 0.214786
R4815 DVDD.n1833 DVDD.n1805 0.214786
R4816 DVDD.n1835 DVDD.n1834 0.214786
R4817 DVDD.n1836 DVDD.n1804 0.214786
R4818 DVDD.n1838 DVDD.n1837 0.214786
R4819 DVDD.n1839 DVDD.n1799 0.214786
R4820 DVDD.n1841 DVDD.n1840 0.214786
R4821 DVDD.n1842 DVDD.n1787 0.214786
R4822 DVDD.n1844 DVDD.n1843 0.214786
R4823 DVDD.n1845 DVDD.n887 0.214786
R4824 DVDD.n1846 DVDD.n882 0.214786
R4825 DVDD.n2979 DVDD.n2978 0.214786
R4826 DVDD.n2980 DVDD.n785 0.214786
R4827 DVDD.n2982 DVDD.n2981 0.214786
R4828 DVDD.n773 DVDD.n772 0.214786
R4829 DVDD.n2987 DVDD.n2986 0.214786
R4830 DVDD.n2988 DVDD.n771 0.214786
R4831 DVDD.n2990 DVDD.n2989 0.214786
R4832 DVDD.n769 DVDD.n768 0.214786
R4833 DVDD.n2995 DVDD.n2994 0.214786
R4834 DVDD.n2996 DVDD.n767 0.214786
R4835 DVDD.n2998 DVDD.n2997 0.214786
R4836 DVDD.n765 DVDD.n764 0.214786
R4837 DVDD.n3003 DVDD.n3002 0.214786
R4838 DVDD.n3004 DVDD.n763 0.214786
R4839 DVDD.n3007 DVDD.n3006 0.214786
R4840 DVDD.n3005 DVDD.n761 0.214786
R4841 DVDD.n3011 DVDD.n760 0.214786
R4842 DVDD.n3013 DVDD.n3012 0.214786
R4843 DVDD.n3014 DVDD.n759 0.214786
R4844 DVDD.n3026 DVDD.n3015 0.214786
R4845 DVDD.n3025 DVDD.n3016 0.214786
R4846 DVDD.n3024 DVDD.n3017 0.214786
R4847 DVDD.n3019 DVDD.n3018 0.214786
R4848 DVDD.n3020 DVDD.n282 0.214786
R4849 DVDD.n4959 DVDD.n283 0.214786
R4850 DVDD.n4963 DVDD.n4962 0.214786
R4851 DVDD.n4964 DVDD.n4958 0.214786
R4852 DVDD.n4966 DVDD.n4965 0.214786
R4853 DVDD.n4956 DVDD.n4955 0.214786
R4854 DVDD.n4971 DVDD.n4970 0.214786
R4855 DVDD.n4972 DVDD.n4954 0.214786
R4856 DVDD.n4974 DVDD.n4973 0.214786
R4857 DVDD.n4952 DVDD.n4951 0.214786
R4858 DVDD.n4979 DVDD.n4978 0.214786
R4859 DVDD.n4980 DVDD.n4950 0.214786
R4860 DVDD.n5244 DVDD.n4981 0.214786
R4861 DVDD.n5243 DVDD.n4982 0.214786
R4862 DVDD.n5241 DVDD.n4983 0.214786
R4863 DVDD.n4986 DVDD.n4984 0.214786
R4864 DVDD.n5237 DVDD.n4987 0.214786
R4865 DVDD.n5236 DVDD.n4988 0.214786
R4866 DVDD.n5235 DVDD.n4989 0.214786
R4867 DVDD.n4992 DVDD.n4990 0.214786
R4868 DVDD.n5231 DVDD.n4993 0.214786
R4869 DVDD.n5230 DVDD.n4994 0.214786
R4870 DVDD.n5229 DVDD.n4995 0.214786
R4871 DVDD.n4998 DVDD.n4996 0.214786
R4872 DVDD.n5225 DVDD.n4999 0.214786
R4873 DVDD.n5223 DVDD.n5071 0.214786
R4874 DVDD.n5074 DVDD.n5072 0.214786
R4875 DVDD.n5219 DVDD.n5075 0.214786
R4876 DVDD.n5218 DVDD.n5076 0.214786
R4877 DVDD.n5217 DVDD.n5077 0.214786
R4878 DVDD.n5156 DVDD.n5078 0.214786
R4879 DVDD.n5200 DVDD.n5157 0.214786
R4880 DVDD.n5199 DVDD.n5158 0.214786
R4881 DVDD.n5198 DVDD.n5159 0.214786
R4882 DVDD.n5162 DVDD.n5160 0.214786
R4883 DVDD.n5194 DVDD.n5163 0.214786
R4884 DVDD.n5193 DVDD.n5164 0.214786
R4885 DVDD.n5192 DVDD.n5165 0.214786
R4886 DVDD.n5168 DVDD.n5166 0.214786
R4887 DVDD.n5188 DVDD.n5169 0.214786
R4888 DVDD.n5187 DVDD.n5170 0.214786
R4889 DVDD.n5186 DVDD.n5171 0.214786
R4890 DVDD.n5174 DVDD.n5172 0.214786
R4891 DVDD.n5182 DVDD.n5175 0.214786
R4892 DVDD.n5181 DVDD.n5176 0.214786
R4893 DVDD.n5180 DVDD.n5178 0.214786
R4894 DVDD.n5177 DVDD.n697 0.214786
R4895 DVDD.n5393 DVDD.n698 0.214786
R4896 DVDD.n5394 DVDD.n659 0.214786
R4897 DVDD.n5430 DVDD.n5429 0.214786
R4898 DVDD.n661 DVDD.n660 0.214786
R4899 DVDD.n5425 DVDD.n5398 0.214786
R4900 DVDD.n5424 DVDD.n5399 0.214786
R4901 DVDD.n5423 DVDD.n5400 0.214786
R4902 DVDD.n5403 DVDD.n5401 0.214786
R4903 DVDD.n5419 DVDD.n5404 0.214786
R4904 DVDD.n5418 DVDD.n5405 0.214786
R4905 DVDD.n5417 DVDD.n5406 0.214786
R4906 DVDD.n5408 DVDD.n5407 0.214786
R4907 DVDD.n5413 DVDD.n5409 0.214786
R4908 DVDD.n5412 DVDD.n5410 0.214786
R4909 DVDD.n5395 DVDD.n5394 0.214786
R4910 DVDD.n5429 DVDD.n5428 0.214786
R4911 DVDD.n5427 DVDD.n661 0.214786
R4912 DVDD.n5426 DVDD.n5425 0.214786
R4913 DVDD.n5424 DVDD.n5397 0.214786
R4914 DVDD.n5423 DVDD.n5422 0.214786
R4915 DVDD.n5421 DVDD.n5401 0.214786
R4916 DVDD.n5420 DVDD.n5419 0.214786
R4917 DVDD.n5418 DVDD.n5402 0.214786
R4918 DVDD.n5417 DVDD.n5416 0.214786
R4919 DVDD.n5415 DVDD.n5407 0.214786
R4920 DVDD.n5414 DVDD.n5413 0.214786
R4921 DVDD.n5393 DVDD.n5392 0.214786
R4922 DVDD.n699 DVDD.n697 0.214786
R4923 DVDD.n5180 DVDD.n5179 0.214786
R4924 DVDD.n5181 DVDD.n5173 0.214786
R4925 DVDD.n5183 DVDD.n5182 0.214786
R4926 DVDD.n5184 DVDD.n5172 0.214786
R4927 DVDD.n5186 DVDD.n5185 0.214786
R4928 DVDD.n5187 DVDD.n5167 0.214786
R4929 DVDD.n5189 DVDD.n5188 0.214786
R4930 DVDD.n5190 DVDD.n5166 0.214786
R4931 DVDD.n5192 DVDD.n5191 0.214786
R4932 DVDD.n5193 DVDD.n5161 0.214786
R4933 DVDD.n5195 DVDD.n5194 0.214786
R4934 DVDD.n5196 DVDD.n5160 0.214786
R4935 DVDD.n5198 DVDD.n5197 0.214786
R4936 DVDD.n5199 DVDD.n5155 0.214786
R4937 DVDD.n5201 DVDD.n5200 0.214786
R4938 DVDD.n5143 DVDD.n5078 0.214786
R4939 DVDD.n5217 DVDD.n5216 0.214786
R4940 DVDD.n5218 DVDD.n5073 0.214786
R4941 DVDD.n5220 DVDD.n5219 0.214786
R4942 DVDD.n5221 DVDD.n5072 0.214786
R4943 DVDD.n5223 DVDD.n5222 0.214786
R4944 DVDD.n5226 DVDD.n5225 0.214786
R4945 DVDD.n5227 DVDD.n4996 0.214786
R4946 DVDD.n5229 DVDD.n5228 0.214786
R4947 DVDD.n5230 DVDD.n4991 0.214786
R4948 DVDD.n5232 DVDD.n5231 0.214786
R4949 DVDD.n5233 DVDD.n4990 0.214786
R4950 DVDD.n5235 DVDD.n5234 0.214786
R4951 DVDD.n5236 DVDD.n4985 0.214786
R4952 DVDD.n5238 DVDD.n5237 0.214786
R4953 DVDD.n5239 DVDD.n4984 0.214786
R4954 DVDD.n5241 DVDD.n5240 0.214786
R4955 DVDD.n5243 DVDD.n5242 0.214786
R4956 DVDD.n5245 DVDD.n5244 0.214786
R4957 DVDD.n4950 DVDD.n4938 0.214786
R4958 DVDD.n4978 DVDD.n4977 0.214786
R4959 DVDD.n4976 DVDD.n4952 0.214786
R4960 DVDD.n4975 DVDD.n4974 0.214786
R4961 DVDD.n4954 DVDD.n4953 0.214786
R4962 DVDD.n4970 DVDD.n4969 0.214786
R4963 DVDD.n4968 DVDD.n4956 0.214786
R4964 DVDD.n4967 DVDD.n4966 0.214786
R4965 DVDD.n4958 DVDD.n4957 0.214786
R4966 DVDD.n4962 DVDD.n4961 0.214786
R4967 DVDD.n4960 DVDD.n4959 0.214786
R4968 DVDD.n3021 DVDD.n3020 0.214786
R4969 DVDD.n3022 DVDD.n3019 0.214786
R4970 DVDD.n3024 DVDD.n3023 0.214786
R4971 DVDD.n3025 DVDD.n758 0.214786
R4972 DVDD.n3027 DVDD.n3026 0.214786
R4973 DVDD.n759 DVDD.n746 0.214786
R4974 DVDD.n3012 DVDD.n745 0.214786
R4975 DVDD.n3011 DVDD.n3010 0.214786
R4976 DVDD.n3009 DVDD.n761 0.214786
R4977 DVDD.n3008 DVDD.n3007 0.214786
R4978 DVDD.n763 DVDD.n762 0.214786
R4979 DVDD.n3002 DVDD.n3001 0.214786
R4980 DVDD.n3000 DVDD.n765 0.214786
R4981 DVDD.n2999 DVDD.n2998 0.214786
R4982 DVDD.n767 DVDD.n766 0.214786
R4983 DVDD.n2994 DVDD.n2993 0.214786
R4984 DVDD.n2992 DVDD.n769 0.214786
R4985 DVDD.n2991 DVDD.n2990 0.214786
R4986 DVDD.n771 DVDD.n770 0.214786
R4987 DVDD.n2986 DVDD.n2985 0.214786
R4988 DVDD.n2984 DVDD.n773 0.214786
R4989 DVDD.n2983 DVDD.n2982 0.214786
R4990 DVDD.n785 DVDD.n243 0.214786
R4991 DVDD.n2978 DVDD.n242 0.214786
R4992 DVDD.n5720 DVDD.n238 0.214786
R4993 DVDD.n231 DVDD.n229 0.214786
R4994 DVDD.n5728 DVDD.n5727 0.214786
R4995 DVDD.n3104 DVDD.n228 0.214786
R4996 DVDD.n3105 DVDD.n3102 0.214786
R4997 DVDD.n3101 DVDD.n3095 0.214786
R4998 DVDD.n3113 DVDD.n3094 0.214786
R4999 DVDD.n3114 DVDD.n3093 0.214786
R5000 DVDD.n3115 DVDD.n3092 0.214786
R5001 DVDD.n3091 DVDD.n3086 0.214786
R5002 DVDD.n3123 DVDD.n3085 0.214786
R5003 DVDD.n3124 DVDD.n3084 0.214786
R5004 DVDD.n3083 DVDD.n189 0.214786
R5005 DVDD.n4796 DVDD.n190 0.214786
R5006 DVDD.n4798 DVDD.n4797 0.214786
R5007 DVDD.n4806 DVDD.n4795 0.214786
R5008 DVDD.n4807 DVDD.n4794 0.214786
R5009 DVDD.n4793 DVDD.n4791 0.214786
R5010 DVDD.n4792 DVDD.n3253 0.214786
R5011 DVDD.n4852 DVDD.n3252 0.214786
R5012 DVDD.n4853 DVDD.n3251 0.214786
R5013 DVDD.n3250 DVDD.n3245 0.214786
R5014 DVDD.n4860 DVDD.n3166 0.214786
R5015 DVDD.n3244 DVDD.n3165 0.214786
R5016 DVDD.n3489 DVDD.n3488 0.214786
R5017 DVDD.n3499 DVDD.n3487 0.214786
R5018 DVDD.n5727 DVDD.n5726 0.214786
R5019 DVDD.n3104 DVDD.n3103 0.214786
R5020 DVDD.n3106 DVDD.n3105 0.214786
R5021 DVDD.n3099 DVDD.n3095 0.214786
R5022 DVDD.n3116 DVDD.n3115 0.214786
R5023 DVDD.n3089 DVDD.n3086 0.214786
R5024 DVDD.n3079 DVDD.n190 0.214786
R5025 DVDD.n4799 DVDD.n4798 0.214786
R5026 DVDD.n4806 DVDD.n4805 0.214786
R5027 DVDD.n4808 DVDD.n4807 0.214786
R5028 DVDD.n4788 DVDD.n3253 0.214786
R5029 DVDD.n4860 DVDD.n4859 0.214786
R5030 DVDD.n3493 DVDD.n3244 0.214786
R5031 DVDD.n3491 DVDD.n3489 0.214786
R5032 DVDD.n3499 DVDD.n3498 0.214786
R5033 DVDD.n3501 DVDD.n3500 0.214786
R5034 DVDD.n3246 DVDD.n3245 0.214786
R5035 DVDD.n4854 DVDD.n4853 0.214786
R5036 DVDD.n4852 DVDD.n4851 0.214786
R5037 DVDD.n4791 DVDD.n4789 0.214786
R5038 DVDD.n3080 DVDD.n189 0.214786
R5039 DVDD.n3125 DVDD.n3124 0.214786
R5040 DVDD.n3123 DVDD.n3122 0.214786
R5041 DVDD.n3114 DVDD.n3090 0.214786
R5042 DVDD.n3113 DVDD.n3112 0.214786
R5043 DVDD.n234 DVDD.n231 0.214786
R5044 DVDD.n5721 DVDD.n5720 0.214786
R5045 DVDD.n5719 DVDD.n5718 0.214786
R5046 DVDD.n5129 DVDD.n5128 0.214786
R5047 DVDD.n5083 DVDD.n5082 0.214786
R5048 DVDD.n5119 DVDD.n5118 0.214786
R5049 DVDD.n5081 DVDD.n5080 0.214786
R5050 DVDD.n5097 DVDD.n5096 0.214786
R5051 DVDD.n5092 DVDD.n5091 0.214786
R5052 DVDD.n726 DVDD.n199 0.214786
R5053 DVDD.n3136 DVDD.n3130 0.214786
R5054 DVDD.n4894 DVDD.n4893 0.214786
R5055 DVDD.n3135 DVDD.n3134 0.214786
R5056 DVDD.n4886 DVDD.n4885 0.214786
R5057 DVDD.n3168 DVDD.n3151 0.214786
R5058 DVDD.n4518 DVDD.n3243 0.214786
R5059 DVDD.n4509 DVDD.n4502 0.214786
R5060 DVDD.n4513 DVDD.n4512 0.214786
R5061 DVDD.n4508 DVDD.n3430 0.214786
R5062 DVDD.n4869 DVDD.n4868 0.214786
R5063 DVDD.n3152 DVDD.n3148 0.214786
R5064 DVDD.n4874 DVDD.n3138 0.214786
R5065 DVDD.n4887 DVDD.n176 0.214786
R5066 DVDD.n732 DVDD.n198 0.214786
R5067 DVDD.n5090 DVDD.n5089 0.214786
R5068 DVDD.n5102 DVDD.n5101 0.214786
R5069 DVDD.n5095 DVDD.n5085 0.214786
R5070 DVDD.n5114 DVDD.n5113 0.214786
R5071 DVDD.n5132 DVDD.n5131 0.214786
R5072 DVDD.n5127 DVDD.n5126 0.214786
R5073 DVDD.n5137 DVDD.n5136 0.214786
R5074 DVDD.n738 DVDD.n736 0.214786
R5075 DVDD.n3055 DVDD.n213 0.214786
R5076 DVDD.n5732 DVDD.n212 0.214786
R5077 DVDD.n5733 DVDD.n211 0.214786
R5078 DVDD.n5738 DVDD.n207 0.214786
R5079 DVDD.n5739 DVDD.n206 0.214786
R5080 DVDD.n734 DVDD.n201 0.214786
R5081 DVDD.n4731 DVDD.n4730 0.214786
R5082 DVDD.n4724 DVDD.n3360 0.214786
R5083 DVDD.n4736 DVDD.n4735 0.214786
R5084 DVDD.n4720 DVDD.n4719 0.214786
R5085 DVDD.n3366 DVDD.n3172 0.214786
R5086 DVDD.n4702 DVDD.n3173 0.214786
R5087 DVDD.n4701 DVDD.n4700 0.214786
R5088 DVDD.n3371 DVDD.n3369 0.214786
R5089 DVDD.n4696 DVDD.n4695 0.214786
R5090 DVDD.n4709 DVDD.n4708 0.214786
R5091 DVDD.n4713 DVDD.n4712 0.214786
R5092 DVDD.n3363 DVDD.n3362 0.214786
R5093 DVDD.n3359 DVDD.n3357 0.214786
R5094 DVDD.n5744 DVDD.n202 0.214786
R5095 DVDD.n3075 DVDD.n203 0.214786
R5096 DVDD.n5740 DVDD.n205 0.214786
R5097 DVDD.n3064 DVDD.n208 0.214786
R5098 DVDD.n5734 DVDD.n210 0.214786
R5099 DVDD.n3051 DVDD.n3050 0.214786
R5100 DVDD.n741 DVDD.n739 0.214786
R5101 DVDD.n3046 DVDD.n3045 0.214786
R5102 DVDD.n3048 DVDD.n739 0.214786
R5103 DVDD.n3050 DVDD.n3049 0.214786
R5104 DVDD.n738 DVDD.n224 0.214786
R5105 DVDD.n5730 DVDD.n213 0.214786
R5106 DVDD.n5732 DVDD.n5731 0.214786
R5107 DVDD.n5733 DVDD.n209 0.214786
R5108 DVDD.n5735 DVDD.n5734 0.214786
R5109 DVDD.n5736 DVDD.n208 0.214786
R5110 DVDD.n5738 DVDD.n5737 0.214786
R5111 DVDD.n5739 DVDD.n204 0.214786
R5112 DVDD.n5741 DVDD.n5740 0.214786
R5113 DVDD.n5742 DVDD.n203 0.214786
R5114 DVDD.n5744 DVDD.n5743 0.214786
R5115 DVDD.n4723 DVDD.n201 0.214786
R5116 DVDD.n4732 DVDD.n4731 0.214786
R5117 DVDD.n4733 DVDD.n3360 0.214786
R5118 DVDD.n4735 DVDD.n4734 0.214786
R5119 DVDD.n4722 DVDD.n3359 0.214786
R5120 DVDD.n4721 DVDD.n4720 0.214786
R5121 DVDD.n3362 DVDD.n3361 0.214786
R5122 DVDD.n4712 DVDD.n4711 0.214786
R5123 DVDD.n4710 DVDD.n4709 0.214786
R5124 DVDD.n3172 DVDD.n3164 0.214786
R5125 DVDD.n3173 DVDD.n3155 0.214786
R5126 DVDD.n4700 DVDD.n4699 0.214786
R5127 DVDD.n4698 DVDD.n3369 0.214786
R5128 DVDD.n5134 DVDD.n5127 0.214786
R5129 DVDD.n5133 DVDD.n5132 0.214786
R5130 DVDD.n5129 DVDD.n220 0.214786
R5131 DVDD.n5083 DVDD.n219 0.214786
R5132 DVDD.n5118 DVDD.n5117 0.214786
R5133 DVDD.n5116 DVDD.n5081 0.214786
R5134 DVDD.n5115 DVDD.n5114 0.214786
R5135 DVDD.n5085 DVDD.n5084 0.214786
R5136 DVDD.n5098 DVDD.n5097 0.214786
R5137 DVDD.n5099 DVDD.n5092 0.214786
R5138 DVDD.n5101 DVDD.n5100 0.214786
R5139 DVDD.n5094 DVDD.n5090 0.214786
R5140 DVDD.n5093 DVDD.n198 0.214786
R5141 DVDD.n4890 DVDD.n199 0.214786
R5142 DVDD.n4891 DVDD.n3136 0.214786
R5143 DVDD.n4893 DVDD.n4892 0.214786
R5144 DVDD.n4889 DVDD.n3135 0.214786
R5145 DVDD.n4888 DVDD.n4887 0.214786
R5146 DVDD.n4886 DVDD.n3137 0.214786
R5147 DVDD.n4865 DVDD.n3138 0.214786
R5148 DVDD.n4866 DVDD.n3152 0.214786
R5149 DVDD.n4868 DVDD.n4867 0.214786
R5150 DVDD.n4864 DVDD.n3151 0.214786
R5151 DVDD.n3243 DVDD.n3156 0.214786
R5152 DVDD.n4510 DVDD.n4509 0.214786
R5153 DVDD.n4512 DVDD.n4511 0.214786
R5154 DVDD.n5363 DVDD.n5362 0.214786
R5155 DVDD.n704 DVDD.n703 0.214786
R5156 DVDD.n5353 DVDD.n216 0.214786
R5157 DVDD.n5348 DVDD.n217 0.214786
R5158 DVDD.n5347 DVDD.n5346 0.214786
R5159 DVDD.n5345 DVDD.n709 0.214786
R5160 DVDD.n5344 DVDD.n5343 0.214786
R5161 DVDD.n711 DVDD.n710 0.214786
R5162 DVDD.n5334 DVDD.n5333 0.214786
R5163 DVDD.n5332 DVDD.n719 0.214786
R5164 DVDD.n5331 DVDD.n5330 0.214786
R5165 DVDD.n722 DVDD.n721 0.214786
R5166 DVDD.n720 DVDD.n192 0.214786
R5167 DVDD.n3217 DVDD.n193 0.214786
R5168 DVDD.n3219 DVDD.n3218 0.214786
R5169 DVDD.n3216 DVDD.n3210 0.214786
R5170 DVDD.n3226 DVDD.n3209 0.214786
R5171 DVDD.n3227 DVDD.n3208 0.214786
R5172 DVDD.n3207 DVDD.n3205 0.214786
R5173 DVDD.n3234 DVDD.n3204 0.214786
R5174 DVDD.n3235 DVDD.n3203 0.214786
R5175 DVDD.n3202 DVDD.n3176 0.214786
R5176 DVDD.n3242 DVDD.n3161 0.214786
R5177 DVDD.n3175 DVDD.n3160 0.214786
R5178 DVDD.n3194 DVDD.n3193 0.214786
R5179 DVDD.n3192 DVDD.n3180 0.214786
R5180 DVDD.n706 DVDD.n702 0.214786
R5181 DVDD.n5354 DVDD.n5353 0.214786
R5182 DVDD.n5349 DVDD.n5348 0.214786
R5183 DVDD.n5347 DVDD.n708 0.214786
R5184 DVDD.n714 DVDD.n709 0.214786
R5185 DVDD.n5335 DVDD.n5334 0.214786
R5186 DVDD.n719 DVDD.n717 0.214786
R5187 DVDD.n728 DVDD.n193 0.214786
R5188 DVDD.n3220 DVDD.n3219 0.214786
R5189 DVDD.n3212 DVDD.n3210 0.214786
R5190 DVDD.n3226 DVDD.n3225 0.214786
R5191 DVDD.n3229 DVDD.n3205 0.214786
R5192 DVDD.n3242 DVDD.n3241 0.214786
R5193 DVDD.n3196 DVDD.n3175 0.214786
R5194 DVDD.n3195 DVDD.n3194 0.214786
R5195 DVDD.n3182 DVDD.n3180 0.214786
R5196 DVDD.n3190 DVDD.n3189 0.214786
R5197 DVDD.n3177 DVDD.n3176 0.214786
R5198 DVDD.n3236 DVDD.n3235 0.214786
R5199 DVDD.n3234 DVDD.n3233 0.214786
R5200 DVDD.n3228 DVDD.n3227 0.214786
R5201 DVDD.n5322 DVDD.n192 0.214786
R5202 DVDD.n5323 DVDD.n722 0.214786
R5203 DVDD.n5330 DVDD.n5329 0.214786
R5204 DVDD.n718 DVDD.n711 0.214786
R5205 DVDD.n5343 DVDD.n5342 0.214786
R5206 DVDD.n5355 DVDD.n704 0.214786
R5207 DVDD.n5362 DVDD.n5361 0.214786
R5208 DVDD DVDD.n730 0.209062
R5209 DVDD.n3169 DVDD.n3153 0.207064
R5210 DVDD.n233 DVDD.n226 0.207064
R5211 DVDD.n233 DVDD.n227 0.2068
R5212 DVDD.n5321 DVDD.n187 0.206795
R5213 DVDD.n804 DVDD.n802 0.2067
R5214 DVDD.n802 DVDD.n801 0.206533
R5215 DVDD.n3169 DVDD.n3154 0.206298
R5216 DVDD.n5321 DVDD.n186 0.206229
R5217 DVDD.n730 DVDD 0.203317
R5218 DVDD.n805 DVDD.n804 0.19985
R5219 DVDD.n187 DVDD.n184 0.199751
R5220 DVDD.n5729 DVDD.n226 0.19948
R5221 DVDD.n4863 DVDD.n3153 0.19948
R5222 DVDD.n4863 DVDD.n3154 0.199329
R5223 DVDD.n186 DVDD.n184 0.198923
R5224 DVDD.n805 DVDD.n801 0.198626
R5225 DVDD.n5729 DVDD.n227 0.198351
R5226 DVDD.n1738 DVDD 0.191946
R5227 DVDD DVDD.n2042 0.191946
R5228 DVDD DVDD.n358 0.191946
R5229 DVDD DVDD.n1486 0.191946
R5230 DVDD DVDD.n1500 0.191946
R5231 DVDD DVDD.n1514 0.191946
R5232 DVDD DVDD.n1528 0.191946
R5233 DVDD DVDD.n2224 0.191946
R5234 DVDD DVDD.n1549 0.191946
R5235 DVDD DVDD.n1226 0.191946
R5236 DVDD DVDD.n1244 0.191946
R5237 DVDD DVDD.n2445 0.191946
R5238 DVDD DVDD.n1258 0.191946
R5239 DVDD DVDD.n1207 0.191946
R5240 DVDD DVDD.n2518 0.191946
R5241 DVDD DVDD.n2534 0.191946
R5242 DVDD DVDD.n2552 0.191946
R5243 DVDD.n2942 DVDD 0.191946
R5244 DVDD DVDD.n5626 0.191946
R5245 DVDD DVDD.n1010 0.191946
R5246 DVDD DVDD.n474 0.191946
R5247 DVDD DVDD.n2570 0.191946
R5248 DVDD.n2760 DVDD 0.191946
R5249 DVDD DVDD.n2918 0.191946
R5250 DVDD DVDD.n525 0.191946
R5251 DVDD.n2769 DVDD 0.191946
R5252 DVDD DVDD.n2783 0.191946
R5253 DVDD DVDD.n2787 0.191946
R5254 DVDD DVDD.n2791 0.191946
R5255 DVDD DVDD.n2795 0.191946
R5256 DVDD DVDD.n2799 0.191946
R5257 DVDD DVDD.n2803 0.191946
R5258 DVDD DVDD.n2807 0.191946
R5259 DVDD DVDD.n2811 0.191946
R5260 DVDD DVDD.n2815 0.191946
R5261 DVDD DVDD.n2819 0.191946
R5262 DVDD DVDD.n2823 0.191946
R5263 DVDD.n2829 DVDD 0.191946
R5264 DVDD.n2845 DVDD 0.191946
R5265 DVDD DVDD.n5519 0.191946
R5266 DVDD.n673 DVDD.n671 0.174559
R5267 DVDD.n233 DVDD.n214 0.174559
R5268 DVDD.n5321 DVDD.n195 0.174559
R5269 DVDD.n3169 DVDD.n3162 0.174401
R5270 DVDD.n674 DVDD 0.174175
R5271 DVDD DVDD.n232 0.172062
R5272 DVDD.n3174 DVDD 0.172062
R5273 DVDD.n4863 DVDD.n3162 0.168052
R5274 DVDD.n675 DVDD.n673 0.16731
R5275 DVDD.n5729 DVDD.n214 0.16731
R5276 DVDD.n195 DVDD.n184 0.16731
R5277 DVDD DVDD.n674 0.167054
R5278 DVDD.n232 DVDD 0.165645
R5279 DVDD.n3174 DVDD 0.165645
R5280 DVDD.n5338 DVDD.n5337 0.1625
R5281 DVDD.n5107 DVDD.n5106 0.1625
R5282 DVDD.n3068 DVDD.n3066 0.1625
R5283 DVDD.n3118 DVDD.n3088 0.1625
R5284 DVDD.n5874 DVDD.n5873 0.159324
R5285 DVDD.n5473 DVDD.n5472 0.159184
R5286 DVDD.n5706 DVDD.n260 0.159184
R5287 DVDD.n5946 DVDD.n47 0.154029
R5288 DVDD.n5881 DVDD.n5880 0.154029
R5289 DVDD.n5952 DVDD.n5950 0.154029
R5290 DVDD.n2232 DVDD.n2231 0.15395
R5291 DVDD.n5644 DVDD.n5643 0.15395
R5292 DVDD.n2961 DVDD.n2960 0.15395
R5293 DVDD.n2218 DVDD.n1127 0.15395
R5294 DVDD.n5808 DVDD.n171 0.1436
R5295 DVDD.n5758 DVDD.n5757 0.1436
R5296 DVDD.n4740 DVDD.n4739 0.1436
R5297 DVDD.n4847 DVDD.n4811 0.1436
R5298 DVDD.n5480 DVDD.n5479 0.1405
R5299 DVDD.n3906 DVDD.n3681 0.139194
R5300 DVDD.n3911 DVDD.n3679 0.139194
R5301 DVDD.n3677 DVDD.n3525 0.139194
R5302 DVDD.n5946 DVDD.n5945 0.138147
R5303 DVDD.n5945 DVDD.n5944 0.138147
R5304 DVDD.n5944 DVDD.n48 0.138147
R5305 DVDD.n5938 DVDD.n48 0.138147
R5306 DVDD.n5938 DVDD.n5937 0.138147
R5307 DVDD.n5937 DVDD.n5936 0.138147
R5308 DVDD.n5936 DVDD.n54 0.138147
R5309 DVDD.n5930 DVDD.n54 0.138147
R5310 DVDD.n5930 DVDD.n5929 0.138147
R5311 DVDD.n5929 DVDD.n5928 0.138147
R5312 DVDD.n5928 DVDD.n62 0.138147
R5313 DVDD.n5922 DVDD.n62 0.138147
R5314 DVDD.n5922 DVDD.n5921 0.138147
R5315 DVDD.n5921 DVDD.n5920 0.138147
R5316 DVDD.n5920 DVDD.n68 0.138147
R5317 DVDD.n5914 DVDD.n68 0.138147
R5318 DVDD.n5914 DVDD.n5913 0.138147
R5319 DVDD.n5913 DVDD.n5912 0.138147
R5320 DVDD.n5912 DVDD.n76 0.138147
R5321 DVDD.n5906 DVDD.n76 0.138147
R5322 DVDD.n5906 DVDD.n5905 0.138147
R5323 DVDD.n5905 DVDD.n5904 0.138147
R5324 DVDD.n5904 DVDD.n82 0.138147
R5325 DVDD.n5898 DVDD.n82 0.138147
R5326 DVDD.n5898 DVDD.n5897 0.138147
R5327 DVDD.n5897 DVDD.n5896 0.138147
R5328 DVDD.n5896 DVDD.n90 0.138147
R5329 DVDD.n5890 DVDD.n90 0.138147
R5330 DVDD.n5890 DVDD.n5889 0.138147
R5331 DVDD.n5889 DVDD.n5888 0.138147
R5332 DVDD.n5888 DVDD.n96 0.138147
R5333 DVDD.n5882 DVDD.n96 0.138147
R5334 DVDD.n5882 DVDD.n5881 0.138147
R5335 DVDD.n5950 DVDD.n43 0.138147
R5336 DVDD.n5834 DVDD.n43 0.138147
R5337 DVDD.n5835 DVDD.n5834 0.138147
R5338 DVDD.n5836 DVDD.n5835 0.138147
R5339 DVDD.n5838 DVDD.n5836 0.138147
R5340 DVDD.n5839 DVDD.n5838 0.138147
R5341 DVDD.n5840 DVDD.n5839 0.138147
R5342 DVDD.n5841 DVDD.n5840 0.138147
R5343 DVDD.n5843 DVDD.n5841 0.138147
R5344 DVDD.n5844 DVDD.n5843 0.138147
R5345 DVDD.n5845 DVDD.n5844 0.138147
R5346 DVDD.n5846 DVDD.n5845 0.138147
R5347 DVDD.n5848 DVDD.n5846 0.138147
R5348 DVDD.n5849 DVDD.n5848 0.138147
R5349 DVDD.n5850 DVDD.n5849 0.138147
R5350 DVDD.n5851 DVDD.n5850 0.138147
R5351 DVDD.n5853 DVDD.n5851 0.138147
R5352 DVDD.n5854 DVDD.n5853 0.138147
R5353 DVDD.n5855 DVDD.n5854 0.138147
R5354 DVDD.n5856 DVDD.n5855 0.138147
R5355 DVDD.n5858 DVDD.n5856 0.138147
R5356 DVDD.n5859 DVDD.n5858 0.138147
R5357 DVDD.n5860 DVDD.n5859 0.138147
R5358 DVDD.n5861 DVDD.n5860 0.138147
R5359 DVDD.n5863 DVDD.n5861 0.138147
R5360 DVDD.n5864 DVDD.n5863 0.138147
R5361 DVDD.n5865 DVDD.n5864 0.138147
R5362 DVDD.n5866 DVDD.n5865 0.138147
R5363 DVDD.n5868 DVDD.n5866 0.138147
R5364 DVDD.n5869 DVDD.n5868 0.138147
R5365 DVDD.n5870 DVDD.n5869 0.138147
R5366 DVDD.n5871 DVDD.n5870 0.138147
R5367 DVDD.n5873 DVDD.n5871 0.138147
R5368 DVDD.n2684 DVDD 0.130618
R5369 DVDD.n4078 DVDD 0.130618
R5370 DVDD.n6019 DVDD 0.13017
R5371 DVDD.n582 DVDD.n359 0.12605
R5372 DVDD.n5648 DVDD.n360 0.12605
R5373 DVDD.n2965 DVDD.n899 0.12605
R5374 DVDD.n2968 DVDD.n2967 0.12605
R5375 DVDD.n5521 DVDD 0.126026
R5376 DVDD DVDD.n2844 0.126026
R5377 DVDD.n2827 DVDD 0.126026
R5378 DVDD.n2825 DVDD 0.126026
R5379 DVDD.n2821 DVDD 0.126026
R5380 DVDD.n2817 DVDD 0.126026
R5381 DVDD.n2813 DVDD 0.126026
R5382 DVDD.n2809 DVDD 0.126026
R5383 DVDD.n2805 DVDD 0.126026
R5384 DVDD.n2801 DVDD 0.126026
R5385 DVDD.n2797 DVDD 0.126026
R5386 DVDD.n2793 DVDD 0.126026
R5387 DVDD.n2789 DVDD 0.126026
R5388 DVDD.n2785 DVDD 0.126026
R5389 DVDD DVDD.n2768 0.126026
R5390 DVDD.n5565 DVDD 0.126026
R5391 DVDD.n2920 DVDD 0.126026
R5392 DVDD.n2758 DVDD 0.126026
R5393 DVDD.n2572 DVDD 0.126026
R5394 DVDD.n2567 DVDD 0.126026
R5395 DVDD.n1013 DVDD 0.126026
R5396 DVDD.n5628 DVDD 0.126026
R5397 DVDD.n2940 DVDD 0.126026
R5398 DVDD.n2558 DVDD 0.126026
R5399 DVDD.n2540 DVDD 0.126026
R5400 DVDD.n2525 DVDD 0.126026
R5401 DVDD.n1209 DVDD 0.126026
R5402 DVDD.n1263 DVDD 0.126026
R5403 DVDD.n2447 DVDD 0.126026
R5404 DVDD.n1251 DVDD 0.126026
R5405 DVDD.n1233 DVDD 0.126026
R5406 DVDD.n1551 DVDD 0.126026
R5407 DVDD.n2226 DVDD 0.126026
R5408 DVDD.n1535 DVDD 0.126026
R5409 DVDD.n1521 DVDD 0.126026
R5410 DVDD.n1507 DVDD 0.126026
R5411 DVDD.n1493 DVDD 0.126026
R5412 DVDD.n5651 DVDD 0.126026
R5413 DVDD.n2044 DVDD 0.126026
R5414 DVDD.n1736 DVDD 0.126026
R5415 DVDD.n3902 DVDD.n3901 0.12425
R5416 DVDD.n4199 DVDD.n3523 0.12425
R5417 DVDD.n5880 DVDD.n104 0.123658
R5418 DVDD.n4813 DVDD.n104 0.123658
R5419 DVDD.n4814 DVDD.n4813 0.123658
R5420 DVDD.n4817 DVDD.n4814 0.123658
R5421 DVDD.n4818 DVDD.n4817 0.123658
R5422 DVDD.n4821 DVDD.n4818 0.123658
R5423 DVDD.n4822 DVDD.n4821 0.123658
R5424 DVDD.n4825 DVDD.n4822 0.123658
R5425 DVDD.n4826 DVDD.n4825 0.123658
R5426 DVDD.n4829 DVDD.n4826 0.123658
R5427 DVDD.n4830 DVDD.n4829 0.123658
R5428 DVDD.n4833 DVDD.n4830 0.123658
R5429 DVDD.n4834 DVDD.n4833 0.123658
R5430 DVDD.n4837 DVDD.n4834 0.123658
R5431 DVDD.n4838 DVDD.n4837 0.123658
R5432 DVDD.n4841 DVDD.n4838 0.123658
R5433 DVDD.n4842 DVDD.n4841 0.123658
R5434 DVDD.n4785 DVDD.n4782 0.123658
R5435 DVDD.n4782 DVDD.n4781 0.123658
R5436 DVDD.n4781 DVDD.n4778 0.123658
R5437 DVDD.n4778 DVDD.n4777 0.123658
R5438 DVDD.n4777 DVDD.n4774 0.123658
R5439 DVDD.n4774 DVDD.n4773 0.123658
R5440 DVDD.n4773 DVDD.n4770 0.123658
R5441 DVDD.n4770 DVDD.n4769 0.123658
R5442 DVDD.n4769 DVDD.n4766 0.123658
R5443 DVDD.n4766 DVDD.n4765 0.123658
R5444 DVDD.n4765 DVDD.n4762 0.123658
R5445 DVDD.n4762 DVDD.n4761 0.123658
R5446 DVDD.n4761 DVDD.n4758 0.123658
R5447 DVDD.n4758 DVDD.n4757 0.123658
R5448 DVDD.n4757 DVDD.n4754 0.123658
R5449 DVDD.n4754 DVDD.n4753 0.123658
R5450 DVDD.n4753 DVDD.n4750 0.123658
R5451 DVDD.n4750 DVDD.n4749 0.123658
R5452 DVDD.n4749 DVDD.n4746 0.123658
R5453 DVDD.n4746 DVDD.n4745 0.123658
R5454 DVDD.n4745 DVDD.n4742 0.123658
R5455 DVDD.n3354 DVDD.n3351 0.123658
R5456 DVDD.n3351 DVDD.n3348 0.123658
R5457 DVDD.n3348 DVDD.n3347 0.123658
R5458 DVDD.n3347 DVDD.n3344 0.123658
R5459 DVDD.n3344 DVDD.n3343 0.123658
R5460 DVDD.n3343 DVDD.n3340 0.123658
R5461 DVDD.n3340 DVDD.n3339 0.123658
R5462 DVDD.n3339 DVDD.n3336 0.123658
R5463 DVDD.n3336 DVDD.n3335 0.123658
R5464 DVDD.n3335 DVDD.n3332 0.123658
R5465 DVDD.n3332 DVDD.n3331 0.123658
R5466 DVDD.n3331 DVDD.n3328 0.123658
R5467 DVDD.n3328 DVDD.n3327 0.123658
R5468 DVDD.n3327 DVDD.n3324 0.123658
R5469 DVDD.n3324 DVDD.n3323 0.123658
R5470 DVDD.n3323 DVDD.n3320 0.123658
R5471 DVDD.n3320 DVDD.n3319 0.123658
R5472 DVDD.n3319 DVDD.n3316 0.123658
R5473 DVDD.n3316 DVDD.n3315 0.123658
R5474 DVDD.n3315 DVDD.n3312 0.123658
R5475 DVDD.n3307 DVDD.n3306 0.123658
R5476 DVDD.n3306 DVDD.n3305 0.123658
R5477 DVDD.n3299 DVDD.n3298 0.123658
R5478 DVDD.n3298 DVDD.n3295 0.123658
R5479 DVDD.n3295 DVDD.n3294 0.123658
R5480 DVDD.n3294 DVDD.n3291 0.123658
R5481 DVDD.n3291 DVDD.n3290 0.123658
R5482 DVDD.n3290 DVDD.n3287 0.123658
R5483 DVDD.n3287 DVDD.n3286 0.123658
R5484 DVDD.n3286 DVDD.n3283 0.123658
R5485 DVDD.n3283 DVDD.n3282 0.123658
R5486 DVDD.n3282 DVDD.n3279 0.123658
R5487 DVDD.n3279 DVDD.n3278 0.123658
R5488 DVDD.n3278 DVDD.n3275 0.123658
R5489 DVDD.n3275 DVDD.n3274 0.123658
R5490 DVDD.n3274 DVDD.n3271 0.123658
R5491 DVDD.n3271 DVDD.n3270 0.123658
R5492 DVDD.n3270 DVDD.n3267 0.123658
R5493 DVDD.n3267 DVDD.n3266 0.123658
R5494 DVDD.n3266 DVDD.n3263 0.123658
R5495 DVDD.n3263 DVDD.n3262 0.123658
R5496 DVDD.n3262 DVDD.n173 0.123658
R5497 DVDD.n5764 DVDD.n5763 0.123658
R5498 DVDD.n5767 DVDD.n5764 0.123658
R5499 DVDD.n5768 DVDD.n5767 0.123658
R5500 DVDD.n5771 DVDD.n5768 0.123658
R5501 DVDD.n5772 DVDD.n5771 0.123658
R5502 DVDD.n5775 DVDD.n5772 0.123658
R5503 DVDD.n5776 DVDD.n5775 0.123658
R5504 DVDD.n5779 DVDD.n5776 0.123658
R5505 DVDD.n5780 DVDD.n5779 0.123658
R5506 DVDD.n5783 DVDD.n5780 0.123658
R5507 DVDD.n5784 DVDD.n5783 0.123658
R5508 DVDD.n5787 DVDD.n5784 0.123658
R5509 DVDD.n5788 DVDD.n5787 0.123658
R5510 DVDD.n5791 DVDD.n5788 0.123658
R5511 DVDD.n5792 DVDD.n5791 0.123658
R5512 DVDD.n5795 DVDD.n5792 0.123658
R5513 DVDD.n5796 DVDD.n5795 0.123658
R5514 DVDD.n5799 DVDD.n5796 0.123658
R5515 DVDD.n5800 DVDD.n5799 0.123658
R5516 DVDD.n5803 DVDD.n5800 0.123658
R5517 DVDD.n5806 DVDD.n5803 0.123658
R5518 DVDD.n5813 DVDD.n5810 0.123658
R5519 DVDD.n5814 DVDD.n5813 0.123658
R5520 DVDD.n5817 DVDD.n5814 0.123658
R5521 DVDD.n5818 DVDD.n5817 0.123658
R5522 DVDD.n5821 DVDD.n5818 0.123658
R5523 DVDD.n5822 DVDD.n5821 0.123658
R5524 DVDD.n5825 DVDD.n5822 0.123658
R5525 DVDD.n5826 DVDD.n5825 0.123658
R5526 DVDD.n5829 DVDD.n5826 0.123658
R5527 DVDD.n5831 DVDD.n5829 0.123658
R5528 DVDD.n4227 DVDD.n47 0.123658
R5529 DVDD.n4227 DVDD.n4225 0.123658
R5530 DVDD.n4233 DVDD.n4225 0.123658
R5531 DVDD.n4234 DVDD.n4233 0.123658
R5532 DVDD.n4235 DVDD.n4234 0.123658
R5533 DVDD.n4235 DVDD.n4223 0.123658
R5534 DVDD.n4241 DVDD.n4223 0.123658
R5535 DVDD.n4242 DVDD.n4241 0.123658
R5536 DVDD.n4243 DVDD.n4242 0.123658
R5537 DVDD.n4243 DVDD.n4221 0.123658
R5538 DVDD.n4249 DVDD.n4221 0.123658
R5539 DVDD.n4250 DVDD.n4249 0.123658
R5540 DVDD.n4251 DVDD.n4250 0.123658
R5541 DVDD.n4251 DVDD.n4219 0.123658
R5542 DVDD.n4256 DVDD.n4219 0.123658
R5543 DVDD.n4257 DVDD.n4256 0.123658
R5544 DVDD.n4257 DVDD.n4217 0.123658
R5545 DVDD.n4313 DVDD.n4261 0.123658
R5546 DVDD.n4313 DVDD.n4312 0.123658
R5547 DVDD.n4312 DVDD.n4311 0.123658
R5548 DVDD.n4311 DVDD.n4263 0.123658
R5549 DVDD.n4306 DVDD.n4263 0.123658
R5550 DVDD.n4306 DVDD.n4305 0.123658
R5551 DVDD.n4305 DVDD.n4304 0.123658
R5552 DVDD.n4304 DVDD.n4266 0.123658
R5553 DVDD.n4299 DVDD.n4266 0.123658
R5554 DVDD.n4299 DVDD.n4298 0.123658
R5555 DVDD.n4298 DVDD.n4297 0.123658
R5556 DVDD.n4297 DVDD.n4269 0.123658
R5557 DVDD.n4292 DVDD.n4269 0.123658
R5558 DVDD.n4292 DVDD.n4291 0.123658
R5559 DVDD.n4291 DVDD.n4290 0.123658
R5560 DVDD.n4290 DVDD.n4272 0.123658
R5561 DVDD.n4285 DVDD.n4272 0.123658
R5562 DVDD.n4285 DVDD.n4284 0.123658
R5563 DVDD.n4284 DVDD.n4283 0.123658
R5564 DVDD.n4283 DVDD.n4275 0.123658
R5565 DVDD.n4278 DVDD.n4275 0.123658
R5566 DVDD.n4682 DVDD.n3378 0.123658
R5567 DVDD.n4677 DVDD.n3378 0.123658
R5568 DVDD.n4677 DVDD.n4676 0.123658
R5569 DVDD.n4676 DVDD.n4675 0.123658
R5570 DVDD.n4675 DVDD.n3381 0.123658
R5571 DVDD.n4670 DVDD.n3381 0.123658
R5572 DVDD.n4670 DVDD.n4669 0.123658
R5573 DVDD.n4669 DVDD.n4668 0.123658
R5574 DVDD.n4668 DVDD.n3384 0.123658
R5575 DVDD.n4663 DVDD.n3384 0.123658
R5576 DVDD.n4663 DVDD.n4662 0.123658
R5577 DVDD.n4662 DVDD.n4661 0.123658
R5578 DVDD.n4661 DVDD.n3387 0.123658
R5579 DVDD.n4656 DVDD.n3387 0.123658
R5580 DVDD.n4656 DVDD.n4655 0.123658
R5581 DVDD.n4655 DVDD.n4654 0.123658
R5582 DVDD.n4654 DVDD.n3390 0.123658
R5583 DVDD.n4649 DVDD.n3390 0.123658
R5584 DVDD.n4649 DVDD.n4648 0.123658
R5585 DVDD.n4648 DVDD.n4647 0.123658
R5586 DVDD.n4642 DVDD.n4641 0.123658
R5587 DVDD.n4641 DVDD.n3398 0.123658
R5588 DVDD.n4638 DVDD.n3403 0.123658
R5589 DVDD.n4633 DVDD.n3403 0.123658
R5590 DVDD.n4633 DVDD.n4632 0.123658
R5591 DVDD.n4632 DVDD.n4631 0.123658
R5592 DVDD.n4631 DVDD.n3409 0.123658
R5593 DVDD.n4626 DVDD.n3409 0.123658
R5594 DVDD.n4626 DVDD.n4625 0.123658
R5595 DVDD.n4625 DVDD.n4624 0.123658
R5596 DVDD.n4624 DVDD.n3412 0.123658
R5597 DVDD.n4619 DVDD.n3412 0.123658
R5598 DVDD.n4619 DVDD.n4618 0.123658
R5599 DVDD.n4618 DVDD.n4617 0.123658
R5600 DVDD.n4617 DVDD.n3415 0.123658
R5601 DVDD.n4612 DVDD.n3415 0.123658
R5602 DVDD.n4612 DVDD.n4611 0.123658
R5603 DVDD.n4611 DVDD.n4610 0.123658
R5604 DVDD.n4610 DVDD.n3418 0.123658
R5605 DVDD.n4605 DVDD.n3418 0.123658
R5606 DVDD.n4605 DVDD.n4604 0.123658
R5607 DVDD.n4604 DVDD.n4603 0.123658
R5608 DVDD.n4598 DVDD.n4597 0.123658
R5609 DVDD.n4597 DVDD.n4596 0.123658
R5610 DVDD.n4596 DVDD.n4546 0.123658
R5611 DVDD.n4591 DVDD.n4546 0.123658
R5612 DVDD.n4591 DVDD.n4590 0.123658
R5613 DVDD.n4590 DVDD.n4589 0.123658
R5614 DVDD.n4589 DVDD.n4549 0.123658
R5615 DVDD.n4584 DVDD.n4549 0.123658
R5616 DVDD.n4584 DVDD.n4583 0.123658
R5617 DVDD.n4583 DVDD.n4582 0.123658
R5618 DVDD.n4582 DVDD.n4552 0.123658
R5619 DVDD.n4577 DVDD.n4552 0.123658
R5620 DVDD.n4577 DVDD.n4576 0.123658
R5621 DVDD.n4576 DVDD.n4575 0.123658
R5622 DVDD.n4575 DVDD.n4555 0.123658
R5623 DVDD.n4570 DVDD.n4555 0.123658
R5624 DVDD.n4570 DVDD.n4569 0.123658
R5625 DVDD.n4569 DVDD.n4568 0.123658
R5626 DVDD.n4568 DVDD.n4558 0.123658
R5627 DVDD.n4563 DVDD.n4558 0.123658
R5628 DVDD.n4563 DVDD.n4562 0.123658
R5629 DVDD.n5982 DVDD.n29 0.123658
R5630 DVDD.n32 DVDD.n29 0.123658
R5631 DVDD.n5975 DVDD.n32 0.123658
R5632 DVDD.n5975 DVDD.n5974 0.123658
R5633 DVDD.n5974 DVDD.n5973 0.123658
R5634 DVDD.n5973 DVDD.n34 0.123658
R5635 DVDD.n5968 DVDD.n34 0.123658
R5636 DVDD.n5968 DVDD.n5967 0.123658
R5637 DVDD.n5967 DVDD.n5966 0.123658
R5638 DVDD.n5966 DVDD.n37 0.123658
R5639 DVDD.n5961 DVDD.n37 0.123658
R5640 DVDD.n5961 DVDD.n5960 0.123658
R5641 DVDD.n5960 DVDD.n5959 0.123658
R5642 DVDD.n5954 DVDD.n41 0.123658
R5643 DVDD.n5954 DVDD.n5953 0.123658
R5644 DVDD.n5953 DVDD.n5952 0.123658
R5645 DVDD.n3310 DVDD.n3257 0.118921
R5646 DVDD.n3303 DVDD.n3302 0.118921
R5647 DVDD.n3397 DVDD.n3395 0.118921
R5648 DVDD.n3402 DVDD.n3400 0.118921
R5649 DVDD.n4741 DVDD.n3255 0.114184
R5650 DVDD.n3312 DVDD.n3311 0.114184
R5651 DVDD.n3299 DVDD.n3259 0.114184
R5652 DVDD.n5760 DVDD.n172 0.114184
R5653 DVDD.n3377 DVDD.n3376 0.114184
R5654 DVDD.n4647 DVDD.n3393 0.114184
R5655 DVDD.n4639 DVDD.n4638 0.114184
R5656 DVDD.n4545 DVDD.n3423 0.114184
R5657 DVDD.n4698 DVDD.n4697 0.110634
R5658 DVDD.n3048 DVDD.n3047 0.110634
R5659 DVDD.n3487 DVDD.n3485 0.110634
R5660 DVDD.n239 DVDD.n238 0.110634
R5661 DVDD.n4511 DVDD.n3429 0.110634
R5662 DVDD.n5135 DVDD.n5134 0.110634
R5663 DVDD.n3192 DVDD.n3191 0.110634
R5664 DVDD.n5364 DVDD.n5363 0.110634
R5665 DVDD.n3355 DVDD.n3354 0.109447
R5666 DVDD.n5759 DVDD.n173 0.109447
R5667 DVDD.n4683 DVDD.n4682 0.109447
R5668 DVDD.n4603 DVDD.n3421 0.109447
R5669 DVDD.n2455 DVDD.n2453 0.10805
R5670 DVDD.n5638 DVDD.n5637 0.10805
R5671 DVDD.n2955 DVDD.n2954 0.10805
R5672 DVDD.n2437 DVDD.n2436 0.10805
R5673 DVDD.n41 DVDD 0.102342
R5674 DVDD DVDD.n6019 0.101194
R5675 DVDD.n2684 DVDD 0.10093
R5676 DVDD.n4078 DVDD 0.10093
R5677 DVDD.n5482 DVDD.n606 0.10085
R5678 DVDD.n5471 DVDD.n626 0.10085
R5679 DVDD.n5705 DVDD.n261 0.10085
R5680 DVDD.n5712 DVDD.n5711 0.10085
R5681 DVDD.n4122 DVDD.n4121 0.0983469
R5682 DVDD.n3762 DVDD.n3761 0.0983469
R5683 DVDD.n2929 DVDD.n526 0.09275
R5684 DVDD.n5562 DVDD.n527 0.09275
R5685 DVDD.n2861 DVDD.n486 0.09275
R5686 DVDD.n2912 DVDD.n2863 0.09275
R5687 DVDD.n4846 DVDD.n4845 0.0881316
R5688 DVDD.n5809 DVDD.n169 0.0881316
R5689 DVDD.n4319 DVDD.n4318 0.0881316
R5690 DVDD.n5983 DVDD.n28 0.0881316
R5691 DVDD.n4786 DVDD.n4785 0.0833947
R5692 DVDD.n5807 DVDD.n5806 0.0833947
R5693 DVDD.n4261 DVDD.n4216 0.0833947
R5694 DVDD.n4562 DVDD.n27 0.0833947
R5695 DVDD.n2569 DVDD.n2568 0.0824403
R5696 DVDD.n5566 DVDD.n524 0.0824403
R5697 DVDD.n2786 DVDD.n524 0.0824403
R5698 DVDD.n2790 DVDD.n2786 0.0824403
R5699 DVDD.n2794 DVDD.n2790 0.0824403
R5700 DVDD.n2798 DVDD.n2794 0.0824403
R5701 DVDD.n2806 DVDD.n2802 0.0824403
R5702 DVDD.n2810 DVDD.n2806 0.0824403
R5703 DVDD.n2814 DVDD.n2810 0.0824403
R5704 DVDD.n2818 DVDD.n2814 0.0824403
R5705 DVDD.n2822 DVDD.n2818 0.0824403
R5706 DVDD.n2826 DVDD.n2822 0.0824403
R5707 DVDD.n2828 DVDD.n2826 0.0824403
R5708 DVDD.n2828 DVDD.n555 0.0824403
R5709 DVDD.n5522 DVDD.n555 0.0824403
R5710 DVDD.n4182 DVDD.n4181 0.0737695
R5711 DVDD.n3800 DVDD.n3508 0.0737695
R5712 DVDD.n2911 DVDD.n2906 0.0718295
R5713 DVDD.n4322 DVDD.n4212 0.0718207
R5714 DVDD.n3704 DVDD.n3699 0.0718204
R5715 DVDD.n4182 DVDD.n16 0.0683695
R5716 DVDD.n3508 DVDD.n3505 0.0683695
R5717 DVDD.n1349 DVDD 0.0638222
R5718 DVDD.n2259 DVDD 0.0638222
R5719 DVDD.n1651 DVDD 0.0638222
R5720 DVDD.n2295 DVDD 0.0638222
R5721 DVDD.n5411 DVDD 0.0638222
R5722 DVDD.n5308 DVDD.n5307 0.0609478
R5723 DVDD DVDD.n1730 0.059934
R5724 DVDD DVDD.n2043 0.059934
R5725 DVDD DVDD.n5650 0.059934
R5726 DVDD DVDD.n1492 0.059934
R5727 DVDD DVDD.n1506 0.059934
R5728 DVDD DVDD.n1520 0.059934
R5729 DVDD DVDD.n1534 0.059934
R5730 DVDD DVDD.n2225 0.059934
R5731 DVDD DVDD.n1550 0.059934
R5732 DVDD DVDD.n1232 0.059934
R5733 DVDD DVDD.n1250 0.059934
R5734 DVDD DVDD.n2446 0.059934
R5735 DVDD DVDD.n1262 0.059934
R5736 DVDD DVDD.n1208 0.059934
R5737 DVDD DVDD.n2524 0.059934
R5738 DVDD DVDD.n2539 0.059934
R5739 DVDD DVDD.n2557 0.059934
R5740 DVDD DVDD.n977 0.059934
R5741 DVDD DVDD.n5627 0.059934
R5742 DVDD DVDD.n1012 0.059934
R5743 DVDD DVDD.n2566 0.059934
R5744 DVDD DVDD.n2571 0.059934
R5745 DVDD DVDD.n2594 0.059934
R5746 DVDD DVDD.n2919 0.059934
R5747 DVDD DVDD.n5564 0.059934
R5748 DVDD DVDD.n2767 0.059934
R5749 DVDD DVDD.n2784 0.059934
R5750 DVDD DVDD.n2788 0.059934
R5751 DVDD DVDD.n2792 0.059934
R5752 DVDD DVDD.n2796 0.059934
R5753 DVDD DVDD.n2800 0.059934
R5754 DVDD DVDD.n2804 0.059934
R5755 DVDD DVDD.n2808 0.059934
R5756 DVDD DVDD.n2812 0.059934
R5757 DVDD DVDD.n2816 0.059934
R5758 DVDD DVDD.n2820 0.059934
R5759 DVDD DVDD.n2824 0.059934
R5760 DVDD DVDD.n2782 0.059934
R5761 DVDD DVDD.n2843 0.059934
R5762 DVDD DVDD.n5520 0.059934
R5763 DVDD.n3831 DVDD.n3830 0.059934
R5764 DVDD.n3845 DVDD.n3538 0.059934
R5765 DVDD.n2906 DVDD.n2864 0.0594957
R5766 DVDD.n3742 DVDD.n3704 0.059485
R5767 DVDD.n4212 DVDD.n3481 0.0594844
R5768 DVDD.n5483 DVDD.n5482 0.05945
R5769 DVDD.n5471 DVDD.n5470 0.05945
R5770 DVDD.n5705 DVDD.n5704 0.05945
R5771 DVDD.n5711 DVDD.n256 0.05945
R5772 DVDD.n1552 DVDD.n1221 0.0577575
R5773 DVDD.n4114 DVDD.n4113 0.0569562
R5774 DVDD.n4109 DVDD.n3557 0.0569562
R5775 DVDD.n4110 DVDD.n3556 0.0569562
R5776 DVDD.n4111 DVDD.n3555 0.0569562
R5777 DVDD.n21 DVDD.n20 0.0569562
R5778 DVDD.n20 DVDD.n19 0.0569562
R5779 DVDD.n19 DVDD.n18 0.0569562
R5780 DVDD.n5985 DVDD.n23 0.0569562
R5781 DVDD.n25 DVDD.n24 0.0569562
R5782 DVDD.n5369 DVDD.n5368 0.0569562
R5783 DVDD.n5371 DVDD.n5370 0.0569562
R5784 DVDD.n5373 DVDD.n5372 0.0569562
R5785 DVDD.n5375 DVDD.n5374 0.0569562
R5786 DVDD.n5377 DVDD.n5376 0.0569562
R5787 DVDD.n5379 DVDD.n5378 0.0569562
R5788 DVDD.n5381 DVDD.n5380 0.0569562
R5789 DVDD.n5383 DVDD.n5382 0.0569562
R5790 DVDD.n5385 DVDD.n5384 0.0569562
R5791 DVDD.n5387 DVDD.n5386 0.0569562
R5792 DVDD.n5390 DVDD.n5389 0.0569562
R5793 DVDD.n5485 DVDD.n5484 0.0569562
R5794 DVDD.n5487 DVDD.n5486 0.0569562
R5795 DVDD.n5489 DVDD.n5488 0.0569562
R5796 DVDD.n5491 DVDD.n5490 0.0569562
R5797 DVDD.n5493 DVDD.n5492 0.0569562
R5798 DVDD.n602 DVDD.n601 0.0569562
R5799 DVDD.n596 DVDD.n595 0.0569562
R5800 DVDD.n595 DVDD.n594 0.0569562
R5801 DVDD.n593 DVDD.n592 0.0569562
R5802 DVDD.n591 DVDD.n590 0.0569562
R5803 DVDD.n589 DVDD.n588 0.0569562
R5804 DVDD.n586 DVDD.n585 0.0569562
R5805 DVDD.n1373 DVDD.n1372 0.0569562
R5806 DVDD.n1376 DVDD.n1375 0.0569562
R5807 DVDD.n1379 DVDD.n1378 0.0569562
R5808 DVDD.n1382 DVDD.n1381 0.0569562
R5809 DVDD.n1385 DVDD.n1384 0.0569562
R5810 DVDD.n2234 DVDD.n2230 0.0569562
R5811 DVDD.n1103 DVDD.n1102 0.0569562
R5812 DVDD.n1105 DVDD.n1104 0.0569562
R5813 DVDD.n1107 DVDD.n1106 0.0569562
R5814 DVDD.n1109 DVDD.n1108 0.0569562
R5815 DVDD.n1111 DVDD.n1110 0.0569562
R5816 DVDD.n1114 DVDD.n1113 0.0569562
R5817 DVDD.n2451 DVDD.n1116 0.0569562
R5818 DVDD.n2454 DVDD.n1098 0.0569562
R5819 DVDD.n1001 DVDD.n989 0.0569562
R5820 DVDD.n1002 DVDD.n991 0.0569562
R5821 DVDD.n1000 DVDD.n986 0.0569562
R5822 DVDD.n999 DVDD.n993 0.0569562
R5823 DVDD.n1003 DVDD.n993 0.0569562
R5824 DVDD.n994 DVDD.n981 0.0569562
R5825 DVDD.n1004 DVDD.n994 0.0569562
R5826 DVDD.n998 DVDD.n996 0.0569562
R5827 DVDD.n1005 DVDD.n996 0.0569562
R5828 DVDD.n2579 DVDD.n2574 0.0569562
R5829 DVDD.n2926 DVDD.n2579 0.0569562
R5830 DVDD.n2925 DVDD.n2581 0.0569562
R5831 DVDD.n2924 DVDD.n2581 0.0569562
R5832 DVDD.n4111 DVDD.n3554 0.0569562
R5833 DVDD.n4110 DVDD.n3555 0.0569562
R5834 DVDD.n4109 DVDD.n3556 0.0569562
R5835 DVDD.n4113 DVDD.n3557 0.0569562
R5836 DVDD.n4114 DVDD.n3551 0.0569562
R5837 DVDD.n5370 DVDD.n5369 0.0569562
R5838 DVDD.n5372 DVDD.n5371 0.0569562
R5839 DVDD.n5374 DVDD.n5373 0.0569562
R5840 DVDD.n5376 DVDD.n5375 0.0569562
R5841 DVDD.n5378 DVDD.n5377 0.0569562
R5842 DVDD.n5380 DVDD.n5379 0.0569562
R5843 DVDD.n5382 DVDD.n5381 0.0569562
R5844 DVDD.n5384 DVDD.n5383 0.0569562
R5845 DVDD.n5386 DVDD.n5385 0.0569562
R5846 DVDD.n5389 DVDD.n5387 0.0569562
R5847 DVDD.n5390 DVDD.n5388 0.0569562
R5848 DVDD.n5486 DVDD.n5485 0.0569562
R5849 DVDD.n5488 DVDD.n5487 0.0569562
R5850 DVDD.n5490 DVDD.n5489 0.0569562
R5851 DVDD.n5492 DVDD.n5491 0.0569562
R5852 DVDD.n5495 DVDD.n602 0.0569562
R5853 DVDD.n601 DVDD.n600 0.0569562
R5854 DVDD.n594 DVDD.n593 0.0569562
R5855 DVDD.n592 DVDD.n591 0.0569562
R5856 DVDD.n590 DVDD.n589 0.0569562
R5857 DVDD.n588 DVDD.n587 0.0569562
R5858 DVDD.n585 DVDD.n584 0.0569562
R5859 DVDD.n1374 DVDD.n1373 0.0569562
R5860 DVDD.n1377 DVDD.n1376 0.0569562
R5861 DVDD.n1380 DVDD.n1379 0.0569562
R5862 DVDD.n1383 DVDD.n1382 0.0569562
R5863 DVDD.n1386 DVDD.n1385 0.0569562
R5864 DVDD.n2235 DVDD.n2234 0.0569562
R5865 DVDD.n1104 DVDD.n1103 0.0569562
R5866 DVDD.n1106 DVDD.n1105 0.0569562
R5867 DVDD.n1108 DVDD.n1107 0.0569562
R5868 DVDD.n1110 DVDD.n1109 0.0569562
R5869 DVDD.n1112 DVDD.n1111 0.0569562
R5870 DVDD.n1115 DVDD.n1114 0.0569562
R5871 DVDD.n1001 DVDD.n990 0.0569562
R5872 DVDD.n1000 DVDD.n985 0.0569562
R5873 DVDD.n2928 DVDD.n2582 0.0569562
R5874 DVDD.n4191 DVDD.n4190 0.0569562
R5875 DVDD.n4190 DVDD.n4189 0.0569562
R5876 DVDD.n4189 DVDD.n4188 0.0569562
R5877 DVDD.n4188 DVDD.n4187 0.0569562
R5878 DVDD.n4542 DVDD.n4541 0.0569562
R5879 DVDD.n4540 DVDD.n4539 0.0569562
R5880 DVDD.n5202 DVDD.n5144 0.0569562
R5881 DVDD.n5203 DVDD.n5145 0.0569562
R5882 DVDD.n5204 DVDD.n5146 0.0569562
R5883 DVDD.n5205 DVDD.n5147 0.0569562
R5884 DVDD.n5206 DVDD.n5148 0.0569562
R5885 DVDD.n5207 DVDD.n5149 0.0569562
R5886 DVDD.n5208 DVDD.n5150 0.0569562
R5887 DVDD.n5209 DVDD.n5151 0.0569562
R5888 DVDD.n5210 DVDD.n5152 0.0569562
R5889 DVDD.n5211 DVDD.n5153 0.0569562
R5890 DVDD.n5214 DVDD.n5213 0.0569562
R5891 DVDD.n633 DVDD.n627 0.0569562
R5892 DVDD.n637 DVDD.n632 0.0569562
R5893 DVDD.n636 DVDD.n631 0.0569562
R5894 DVDD.n635 DVDD.n630 0.0569562
R5895 DVDD.n634 DVDD.n629 0.0569562
R5896 DVDD.n1698 DVDD.n1600 0.0569562
R5897 DVDD.n1699 DVDD.n1601 0.0569562
R5898 DVDD.n1702 DVDD.n1595 0.0569562
R5899 DVDD.n1702 DVDD.n1602 0.0569562
R5900 DVDD.n1703 DVDD.n1603 0.0569562
R5901 DVDD.n1704 DVDD.n1604 0.0569562
R5902 DVDD.n1705 DVDD.n1605 0.0569562
R5903 DVDD.n1707 DVDD.n1607 0.0569562
R5904 DVDD.n369 DVDD.n361 0.0569562
R5905 DVDD.n2069 DVDD.n371 0.0569562
R5906 DVDD.n2071 DVDD.n373 0.0569562
R5907 DVDD.n2073 DVDD.n375 0.0569562
R5908 DVDD.n2075 DVDD.n377 0.0569562
R5909 DVDD.n2077 DVDD.n379 0.0569562
R5910 DVDD.n402 DVDD.n390 0.0569562
R5911 DVDD.n403 DVDD.n391 0.0569562
R5912 DVDD.n404 DVDD.n392 0.0569562
R5913 DVDD.n405 DVDD.n393 0.0569562
R5914 DVDD.n406 DVDD.n394 0.0569562
R5915 DVDD.n408 DVDD.n396 0.0569562
R5916 DVDD.n410 DVDD.n398 0.0569562
R5917 DVDD.n5640 DVDD.n384 0.0569562
R5918 DVDD.n421 DVDD.n412 0.0569562
R5919 DVDD.n438 DVDD.n423 0.0569562
R5920 DVDD.n434 DVDD.n418 0.0569562
R5921 DVDD.n440 DVDD.n416 0.0569562
R5922 DVDD.n440 DVDD.n425 0.0569562
R5923 DVDD.n442 DVDD.n415 0.0569562
R5924 DVDD.n442 DVDD.n426 0.0569562
R5925 DVDD.n5632 DVDD.n414 0.0569562
R5926 DVDD.n5632 DVDD.n427 0.0569562
R5927 DVDD.n2748 DVDD.n2612 0.0569562
R5928 DVDD.n2749 DVDD.n2612 0.0569562
R5929 DVDD.n2613 DVDD.n2606 0.0569562
R5930 DVDD.n2750 DVDD.n2613 0.0569562
R5931 DVDD.n2753 DVDD.n2752 0.0569562
R5932 DVDD.n5203 DVDD.n5144 0.0569562
R5933 DVDD.n5204 DVDD.n5145 0.0569562
R5934 DVDD.n5205 DVDD.n5146 0.0569562
R5935 DVDD.n5206 DVDD.n5147 0.0569562
R5936 DVDD.n5207 DVDD.n5148 0.0569562
R5937 DVDD.n5208 DVDD.n5149 0.0569562
R5938 DVDD.n5209 DVDD.n5150 0.0569562
R5939 DVDD.n5210 DVDD.n5151 0.0569562
R5940 DVDD.n5211 DVDD.n5152 0.0569562
R5941 DVDD.n5213 DVDD.n5153 0.0569562
R5942 DVDD.n5214 DVDD.n5154 0.0569562
R5943 DVDD.n637 DVDD.n633 0.0569562
R5944 DVDD.n636 DVDD.n632 0.0569562
R5945 DVDD.n635 DVDD.n631 0.0569562
R5946 DVDD.n634 DVDD.n630 0.0569562
R5947 DVDD.n1699 DVDD.n1600 0.0569562
R5948 DVDD.n1703 DVDD.n1602 0.0569562
R5949 DVDD.n1704 DVDD.n1603 0.0569562
R5950 DVDD.n1705 DVDD.n1604 0.0569562
R5951 DVDD.n1706 DVDD.n1605 0.0569562
R5952 DVDD.n1710 DVDD.n1607 0.0569562
R5953 DVDD.n2068 DVDD.n369 0.0569562
R5954 DVDD.n2070 DVDD.n371 0.0569562
R5955 DVDD.n2072 DVDD.n373 0.0569562
R5956 DVDD.n2074 DVDD.n375 0.0569562
R5957 DVDD.n2076 DVDD.n377 0.0569562
R5958 DVDD.n380 DVDD.n379 0.0569562
R5959 DVDD.n403 DVDD.n390 0.0569562
R5960 DVDD.n404 DVDD.n391 0.0569562
R5961 DVDD.n405 DVDD.n392 0.0569562
R5962 DVDD.n406 DVDD.n393 0.0569562
R5963 DVDD.n407 DVDD.n394 0.0569562
R5964 DVDD.n409 DVDD.n396 0.0569562
R5965 DVDD.n437 DVDD.n421 0.0569562
R5966 DVDD.n433 DVDD.n418 0.0569562
R5967 DVDD.n3515 DVDD.n3514 0.0569562
R5968 DVDD.n3514 DVDD.n3513 0.0569562
R5969 DVDD.n3513 DVDD.n3512 0.0569562
R5970 DVDD.n3512 DVDD.n3511 0.0569562
R5971 DVDD.n4687 DVDD.n4686 0.0569562
R5972 DVDD.n4689 DVDD.n4688 0.0569562
R5973 DVDD.n747 DVDD.n744 0.0569562
R5974 DVDD.n3028 DVDD.n748 0.0569562
R5975 DVDD.n3029 DVDD.n749 0.0569562
R5976 DVDD.n3030 DVDD.n750 0.0569562
R5977 DVDD.n3031 DVDD.n751 0.0569562
R5978 DVDD.n3032 DVDD.n752 0.0569562
R5979 DVDD.n3033 DVDD.n753 0.0569562
R5980 DVDD.n3034 DVDD.n754 0.0569562
R5981 DVDD.n3035 DVDD.n755 0.0569562
R5982 DVDD.n3036 DVDD.n756 0.0569562
R5983 DVDD.n3039 DVDD.n3038 0.0569562
R5984 DVDD.n268 DVDD.n262 0.0569562
R5985 DVDD.n272 DVDD.n267 0.0569562
R5986 DVDD.n271 DVDD.n266 0.0569562
R5987 DVDD.n270 DVDD.n265 0.0569562
R5988 DVDD.n269 DVDD.n264 0.0569562
R5989 DVDD.n2025 DVDD.n1724 0.0569562
R5990 DVDD.n2026 DVDD.n1725 0.0569562
R5991 DVDD.n2029 DVDD.n1719 0.0569562
R5992 DVDD.n2029 DVDD.n1726 0.0569562
R5993 DVDD.n2030 DVDD.n1727 0.0569562
R5994 DVDD.n2031 DVDD.n1728 0.0569562
R5995 DVDD.n2032 DVDD.n1729 0.0569562
R5996 DVDD.n2036 DVDD.n2035 0.0569562
R5997 DVDD.n908 DVDD.n900 0.0569562
R5998 DVDD.n1437 DVDD.n910 0.0569562
R5999 DVDD.n1439 DVDD.n912 0.0569562
R6000 DVDD.n1441 DVDD.n914 0.0569562
R6001 DVDD.n1443 DVDD.n916 0.0569562
R6002 DVDD.n1445 DVDD.n918 0.0569562
R6003 DVDD.n941 DVDD.n929 0.0569562
R6004 DVDD.n942 DVDD.n930 0.0569562
R6005 DVDD.n943 DVDD.n931 0.0569562
R6006 DVDD.n944 DVDD.n932 0.0569562
R6007 DVDD.n945 DVDD.n933 0.0569562
R6008 DVDD.n947 DVDD.n935 0.0569562
R6009 DVDD.n949 DVDD.n937 0.0569562
R6010 DVDD.n2957 DVDD.n923 0.0569562
R6011 DVDD.n960 DVDD.n951 0.0569562
R6012 DVDD.n974 DVDD.n962 0.0569562
R6013 DVDD.n970 DVDD.n957 0.0569562
R6014 DVDD.n976 DVDD.n955 0.0569562
R6015 DVDD.n976 DVDD.n964 0.0569562
R6016 DVDD.n2947 DVDD.n954 0.0569562
R6017 DVDD.n2947 DVDD.n965 0.0569562
R6018 DVDD.n2950 DVDD.n953 0.0569562
R6019 DVDD.n2951 DVDD.n2950 0.0569562
R6020 DVDD.n482 DVDD.n477 0.0569562
R6021 DVDD.n5610 DVDD.n482 0.0569562
R6022 DVDD.n5609 DVDD.n484 0.0569562
R6023 DVDD.n5611 DVDD.n484 0.0569562
R6024 DVDD.n5614 DVDD.n5613 0.0569562
R6025 DVDD.n3028 DVDD.n747 0.0569562
R6026 DVDD.n3029 DVDD.n748 0.0569562
R6027 DVDD.n3030 DVDD.n749 0.0569562
R6028 DVDD.n3031 DVDD.n750 0.0569562
R6029 DVDD.n3032 DVDD.n751 0.0569562
R6030 DVDD.n3033 DVDD.n752 0.0569562
R6031 DVDD.n3034 DVDD.n753 0.0569562
R6032 DVDD.n3035 DVDD.n754 0.0569562
R6033 DVDD.n3036 DVDD.n755 0.0569562
R6034 DVDD.n3038 DVDD.n756 0.0569562
R6035 DVDD.n3039 DVDD.n757 0.0569562
R6036 DVDD.n272 DVDD.n268 0.0569562
R6037 DVDD.n271 DVDD.n267 0.0569562
R6038 DVDD.n270 DVDD.n266 0.0569562
R6039 DVDD.n269 DVDD.n265 0.0569562
R6040 DVDD.n2026 DVDD.n1724 0.0569562
R6041 DVDD.n2030 DVDD.n1726 0.0569562
R6042 DVDD.n2031 DVDD.n1727 0.0569562
R6043 DVDD.n2032 DVDD.n1728 0.0569562
R6044 DVDD.n2033 DVDD.n1729 0.0569562
R6045 DVDD.n2036 DVDD.n1743 0.0569562
R6046 DVDD.n1436 DVDD.n908 0.0569562
R6047 DVDD.n1438 DVDD.n910 0.0569562
R6048 DVDD.n1440 DVDD.n912 0.0569562
R6049 DVDD.n1442 DVDD.n914 0.0569562
R6050 DVDD.n1444 DVDD.n916 0.0569562
R6051 DVDD.n919 DVDD.n918 0.0569562
R6052 DVDD.n942 DVDD.n929 0.0569562
R6053 DVDD.n943 DVDD.n930 0.0569562
R6054 DVDD.n944 DVDD.n931 0.0569562
R6055 DVDD.n945 DVDD.n932 0.0569562
R6056 DVDD.n946 DVDD.n933 0.0569562
R6057 DVDD.n948 DVDD.n935 0.0569562
R6058 DVDD.n973 DVDD.n960 0.0569562
R6059 DVDD.n969 DVDD.n957 0.0569562
R6060 DVDD.n3755 DVDD.n3754 0.0569562
R6061 DVDD.n3754 DVDD.n3753 0.0569562
R6062 DVDD.n3753 DVDD.n3752 0.0569562
R6063 DVDD.n3752 DVDD.n3751 0.0569562
R6064 DVDD.n3751 DVDD.n3750 0.0569562
R6065 DVDD.n3750 DVDD.n3749 0.0569562
R6066 DVDD.n3749 DVDD.n3748 0.0569562
R6067 DVDD.n3748 DVDD.n3747 0.0569562
R6068 DVDD.n3747 DVDD.n3746 0.0569562
R6069 DVDD.n4213 DVDD.n3507 0.0569562
R6070 DVDD.n4214 DVDD.n3507 0.0569562
R6071 DVDD.n4214 DVDD.n3506 0.0569562
R6072 DVDD.n4323 DVDD.n4209 0.0569562
R6073 DVDD.n4324 DVDD.n4210 0.0569562
R6074 DVDD.n244 DVDD.n241 0.0569562
R6075 DVDD.n774 DVDD.n245 0.0569562
R6076 DVDD.n775 DVDD.n246 0.0569562
R6077 DVDD.n776 DVDD.n247 0.0569562
R6078 DVDD.n777 DVDD.n248 0.0569562
R6079 DVDD.n778 DVDD.n249 0.0569562
R6080 DVDD.n779 DVDD.n250 0.0569562
R6081 DVDD.n780 DVDD.n251 0.0569562
R6082 DVDD.n781 DVDD.n252 0.0569562
R6083 DVDD.n782 DVDD.n253 0.0569562
R6084 DVDD.n783 DVDD.n254 0.0569562
R6085 DVDD.n838 DVDD.n833 0.0569562
R6086 DVDD.n837 DVDD.n832 0.0569562
R6087 DVDD.n836 DVDD.n831 0.0569562
R6088 DVDD.n835 DVDD.n830 0.0569562
R6089 DVDD.n834 DVDD.n829 0.0569562
R6090 DVDD.n888 DVDD.n881 0.0569562
R6091 DVDD.n1788 DVDD.n889 0.0569562
R6092 DVDD.n1791 DVDD.n885 0.0569562
R6093 DVDD.n1791 DVDD.n890 0.0569562
R6094 DVDD.n1792 DVDD.n891 0.0569562
R6095 DVDD.n1793 DVDD.n892 0.0569562
R6096 DVDD.n1794 DVDD.n893 0.0569562
R6097 DVDD.n1796 DVDD.n895 0.0569562
R6098 DVDD.n2206 DVDD.n1399 0.0569562
R6099 DVDD.n2208 DVDD.n1401 0.0569562
R6100 DVDD.n2210 DVDD.n1403 0.0569562
R6101 DVDD.n2212 DVDD.n1405 0.0569562
R6102 DVDD.n2214 DVDD.n1407 0.0569562
R6103 DVDD.n1408 DVDD.n1392 0.0569562
R6104 DVDD.n2427 DVDD.n1130 0.0569562
R6105 DVDD.n2428 DVDD.n1131 0.0569562
R6106 DVDD.n2429 DVDD.n1132 0.0569562
R6107 DVDD.n2430 DVDD.n1133 0.0569562
R6108 DVDD.n2431 DVDD.n1134 0.0569562
R6109 DVDD.n2433 DVDD.n1136 0.0569562
R6110 DVDD.n1137 DVDD.n1122 0.0569562
R6111 DVDD.n2439 DVDD.n1124 0.0569562
R6112 DVDD.n467 DVDD.n455 0.0569562
R6113 DVDD.n468 DVDD.n457 0.0569562
R6114 DVDD.n466 DVDD.n452 0.0569562
R6115 DVDD.n465 DVDD.n459 0.0569562
R6116 DVDD.n469 DVDD.n459 0.0569562
R6117 DVDD.n464 DVDD.n461 0.0569562
R6118 DVDD.n470 DVDD.n461 0.0569562
R6119 DVDD.n462 DVDD.n447 0.0569562
R6120 DVDD.n471 DVDD.n462 0.0569562
R6121 DVDD.n2908 DVDD.n2593 0.0569562
R6122 DVDD.n2909 DVDD.n2593 0.0569562
R6123 DVDD.n2907 DVDD.n2765 0.0569562
R6124 DVDD.n2910 DVDD.n2765 0.0569562
R6125 DVDD.n2913 DVDD.n2588 0.0569562
R6126 DVDD.n774 DVDD.n244 0.0569562
R6127 DVDD.n775 DVDD.n245 0.0569562
R6128 DVDD.n776 DVDD.n246 0.0569562
R6129 DVDD.n777 DVDD.n247 0.0569562
R6130 DVDD.n778 DVDD.n248 0.0569562
R6131 DVDD.n779 DVDD.n249 0.0569562
R6132 DVDD.n780 DVDD.n250 0.0569562
R6133 DVDD.n781 DVDD.n251 0.0569562
R6134 DVDD.n782 DVDD.n252 0.0569562
R6135 DVDD.n783 DVDD.n253 0.0569562
R6136 DVDD.n255 DVDD.n254 0.0569562
R6137 DVDD.n837 DVDD.n833 0.0569562
R6138 DVDD.n836 DVDD.n832 0.0569562
R6139 DVDD.n835 DVDD.n831 0.0569562
R6140 DVDD.n834 DVDD.n830 0.0569562
R6141 DVDD.n1788 DVDD.n888 0.0569562
R6142 DVDD.n1792 DVDD.n890 0.0569562
R6143 DVDD.n1793 DVDD.n891 0.0569562
R6144 DVDD.n1794 DVDD.n892 0.0569562
R6145 DVDD.n1795 DVDD.n893 0.0569562
R6146 DVDD.n1797 DVDD.n895 0.0569562
R6147 DVDD.n2207 DVDD.n1399 0.0569562
R6148 DVDD.n2209 DVDD.n1401 0.0569562
R6149 DVDD.n2211 DVDD.n1403 0.0569562
R6150 DVDD.n2213 DVDD.n1405 0.0569562
R6151 DVDD.n2215 DVDD.n1407 0.0569562
R6152 DVDD.n2217 DVDD.n1408 0.0569562
R6153 DVDD.n2428 DVDD.n1130 0.0569562
R6154 DVDD.n2429 DVDD.n1131 0.0569562
R6155 DVDD.n2430 DVDD.n1132 0.0569562
R6156 DVDD.n2431 DVDD.n1133 0.0569562
R6157 DVDD.n2432 DVDD.n1134 0.0569562
R6158 DVDD.n2434 DVDD.n1136 0.0569562
R6159 DVDD.n467 DVDD.n456 0.0569562
R6160 DVDD.n466 DVDD.n451 0.0569562
R6161 DVDD.n4324 DVDD.n4323 0.0569562
R6162 DVDD.n4688 DVDD.n4687 0.0569562
R6163 DVDD.n4541 DVDD.n4540 0.0569562
R6164 DVDD.n24 DVDD.n23 0.0569562
R6165 DVDD.n3187 DVDD.n3185 0.0563
R6166 DVDD.n3187 DVDD.n3186 0.0563
R6167 DVDD.n3186 DVDD.n3178 0.0563
R6168 DVDD.n3198 DVDD.n3178 0.0563
R6169 DVDD.n3199 DVDD.n3198 0.0563
R6170 DVDD.n3239 DVDD.n3199 0.0563
R6171 DVDD.n3239 DVDD.n3238 0.0563
R6172 DVDD.n3238 DVDD.n3200 0.0563
R6173 DVDD.n3231 DVDD.n3200 0.0563
R6174 DVDD.n3231 DVDD.n170 0.0563
R6175 DVDD.n3213 DVDD.n171 0.0563
R6176 DVDD.n3223 DVDD.n3213 0.0563
R6177 DVDD.n3223 DVDD.n3222 0.0563
R6178 DVDD.n3222 DVDD.n3214 0.0563
R6179 DVDD.n3214 DVDD.n725 0.0563
R6180 DVDD.n5325 DVDD.n725 0.0563
R6181 DVDD.n5326 DVDD.n5325 0.0563
R6182 DVDD.n5327 DVDD.n5326 0.0563
R6183 DVDD.n5327 DVDD.n716 0.0563
R6184 DVDD.n5337 DVDD.n716 0.0563
R6185 DVDD.n5340 DVDD.n5338 0.0563
R6186 DVDD.n5340 DVDD.n5339 0.0563
R6187 DVDD.n5339 DVDD.n707 0.0563
R6188 DVDD.n5351 DVDD.n707 0.0563
R6189 DVDD.n5352 DVDD.n5351 0.0563
R6190 DVDD.n5357 DVDD.n5352 0.0563
R6191 DVDD.n5358 DVDD.n5357 0.0563
R6192 DVDD.n5359 DVDD.n5358 0.0563
R6193 DVDD.n5359 DVDD.n700 0.0563
R6194 DVDD.n5366 DVDD.n700 0.0563
R6195 DVDD.n4537 DVDD.n3428 0.0563
R6196 DVDD.n4503 DVDD.n3428 0.0563
R6197 DVDD.n4515 DVDD.n4503 0.0563
R6198 DVDD.n4517 DVDD.n4515 0.0563
R6199 DVDD.n4517 DVDD.n4516 0.0563
R6200 DVDD.n4516 DVDD.n3149 0.0563
R6201 DVDD.n4871 DVDD.n3149 0.0563
R6202 DVDD.n4873 DVDD.n4871 0.0563
R6203 DVDD.n4873 DVDD.n4872 0.0563
R6204 DVDD.n4872 DVDD.n174 0.0563
R6205 DVDD.n5757 DVDD.n175 0.0563
R6206 DVDD.n3131 DVDD.n175 0.0563
R6207 DVDD.n4896 DVDD.n3131 0.0563
R6208 DVDD.n4897 DVDD.n4896 0.0563
R6209 DVDD.n4897 DVDD.n727 0.0563
R6210 DVDD.n5086 DVDD.n727 0.0563
R6211 DVDD.n5087 DVDD.n5086 0.0563
R6212 DVDD.n5104 DVDD.n5087 0.0563
R6213 DVDD.n5105 DVDD.n5104 0.0563
R6214 DVDD.n5106 DVDD.n5105 0.0563
R6215 DVDD.n5108 DVDD.n5107 0.0563
R6216 DVDD.n5108 DVDD.n5079 0.0563
R6217 DVDD.n5121 DVDD.n5079 0.0563
R6218 DVDD.n5122 DVDD.n5121 0.0563
R6219 DVDD.n5123 DVDD.n5122 0.0563
R6220 DVDD.n5124 DVDD.n5123 0.0563
R6221 DVDD.n5125 DVDD.n5124 0.0563
R6222 DVDD.n5139 DVDD.n5125 0.0563
R6223 DVDD.n5140 DVDD.n5139 0.0563
R6224 DVDD.n5141 DVDD.n5140 0.0563
R6225 DVDD.n4693 DVDD.n4691 0.0563
R6226 DVDD.n4693 DVDD.n4692 0.0563
R6227 DVDD.n4692 DVDD.n3367 0.0563
R6228 DVDD.n4704 DVDD.n3367 0.0563
R6229 DVDD.n4705 DVDD.n4704 0.0563
R6230 DVDD.n4706 DVDD.n4705 0.0563
R6231 DVDD.n4706 DVDD.n3364 0.0563
R6232 DVDD.n4715 DVDD.n3364 0.0563
R6233 DVDD.n4716 DVDD.n4715 0.0563
R6234 DVDD.n4716 DVDD.n3256 0.0563
R6235 DVDD.n4739 DVDD.n3356 0.0563
R6236 DVDD.n4726 DVDD.n3356 0.0563
R6237 DVDD.n4727 DVDD.n4726 0.0563
R6238 DVDD.n4728 DVDD.n4727 0.0563
R6239 DVDD.n4728 DVDD.n3078 0.0563
R6240 DVDD.n3078 DVDD.n3077 0.0563
R6241 DVDD.n3077 DVDD.n3073 0.0563
R6242 DVDD.n3073 DVDD.n3072 0.0563
R6243 DVDD.n3072 DVDD.n3069 0.0563
R6244 DVDD.n3069 DVDD.n3068 0.0563
R6245 DVDD.n3066 DVDD.n3063 0.0563
R6246 DVDD.n3063 DVDD.n3060 0.0563
R6247 DVDD.n3060 DVDD.n3059 0.0563
R6248 DVDD.n3059 DVDD.n3057 0.0563
R6249 DVDD.n3057 DVDD.n3054 0.0563
R6250 DVDD.n3054 DVDD.n3053 0.0563
R6251 DVDD.n3053 DVDD.n735 0.0563
R6252 DVDD.n743 DVDD.n735 0.0563
R6253 DVDD.n3043 DVDD.n743 0.0563
R6254 DVDD.n3043 DVDD.n3042 0.0563
R6255 DVDD.n3503 DVDD.n3484 0.0563
R6256 DVDD.n3492 DVDD.n3484 0.0563
R6257 DVDD.n3496 DVDD.n3492 0.0563
R6258 DVDD.n3496 DVDD.n3495 0.0563
R6259 DVDD.n3495 DVDD.n3247 0.0563
R6260 DVDD.n4857 DVDD.n3247 0.0563
R6261 DVDD.n4857 DVDD.n4856 0.0563
R6262 DVDD.n4856 DVDD.n3248 0.0563
R6263 DVDD.n4849 DVDD.n3248 0.0563
R6264 DVDD.n4849 DVDD.n4848 0.0563
R6265 DVDD.n4811 DVDD.n4787 0.0563
R6266 DVDD.n4800 DVDD.n4787 0.0563
R6267 DVDD.n4803 DVDD.n4800 0.0563
R6268 DVDD.n4803 DVDD.n4802 0.0563
R6269 DVDD.n4802 DVDD.n3128 0.0563
R6270 DVDD.n3128 DVDD.n3127 0.0563
R6271 DVDD.n3127 DVDD.n3081 0.0563
R6272 DVDD.n3120 DVDD.n3081 0.0563
R6273 DVDD.n3120 DVDD.n3119 0.0563
R6274 DVDD.n3119 DVDD.n3118 0.0563
R6275 DVDD.n3110 DVDD.n3088 0.0563
R6276 DVDD.n3110 DVDD.n3109 0.0563
R6277 DVDD.n3109 DVDD.n3108 0.0563
R6278 DVDD.n3108 DVDD.n3098 0.0563
R6279 DVDD.n3098 DVDD.n235 0.0563
R6280 DVDD.n5724 DVDD.n235 0.0563
R6281 DVDD.n5724 DVDD.n5723 0.0563
R6282 DVDD.n5723 DVDD.n236 0.0563
R6283 DVDD.n5716 DVDD.n236 0.0563
R6284 DVDD.n5716 DVDD.n5715 0.0563
R6285 DVDD.n1260 DVDD.n1099 0.05585
R6286 DVDD.n2536 DVDD.n987 0.05585
R6287 DVDD.n400 DVDD.n399 0.05585
R6288 DVDD.n2537 DVDD.n435 0.05585
R6289 DVDD.n939 DVDD.n938 0.05585
R6290 DVDD.n2530 DVDD.n971 0.05585
R6291 DVDD.n1139 DVDD.n1138 0.05585
R6292 DVDD.n2532 DVDD.n453 0.05585
R6293 DVDD.n5984 DVDD.n26 0.0554
R6294 DVDD.n4544 DVDD.n3425 0.0554
R6295 DVDD.n4684 DVDD.n3375 0.0554
R6296 DVDD.n4320 DVDD.n4215 0.0554
R6297 DVDD.n5755 DVDD.n178 0.0538955
R6298 DVDD.n2450 DVDD.n2449 0.05315
R6299 DVDD.n2521 DVDD.n2520 0.05315
R6300 DVDD.n1118 DVDD.n385 0.05315
R6301 DVDD.n2522 DVDD.n419 0.05315
R6302 DVDD.n1120 DVDD.n924 0.05315
R6303 DVDD.n2513 DVDD.n958 0.05315
R6304 DVDD.n2443 DVDD.n2442 0.05315
R6305 DVDD.n2516 DVDD.n2515 0.05315
R6306 DVDD.n2554 DVDD.n2553 0.05225
R6307 DVDD.n2555 DVDD.n417 0.05225
R6308 DVDD.n2548 DVDD.n956 0.05225
R6309 DVDD.n2550 DVDD.n2549 0.05225
R6310 DVDD.n5456 DVDD.n646 0.0515891
R6311 DVDD.n863 DVDD.n850 0.0515891
R6312 DVDD.n4861 DVDD.n3167 0.0515849
R6313 DVDD.n230 DVDD.n215 0.0515849
R6314 DVDD.n230 DVDD.n221 0.0515849
R6315 DVDD.n4861 DVDD.n3163 0.0515849
R6316 DVDD.n5745 DVDD.n191 0.0515835
R6317 DVDD.n5745 DVDD.n196 0.0515835
R6318 DVDD.n4183 DVDD.n22 0.0509
R6319 DVDD.n4208 DVDD.n4207 0.0509
R6320 DVDD.n4862 DVDD.n4861 0.0498479
R6321 DVDD.n4861 DVDD.n3159 0.0498479
R6322 DVDD.n3905 DVDD.n3904 0.049839
R6323 DVDD.n3671 DVDD.n3669 0.049839
R6324 DVDD.n3675 DVDD.n3673 0.049839
R6325 DVDD.n3522 DVDD.n3520 0.049839
R6326 DVDD.n3851 DVDD.n3850 0.049839
R6327 DVDD.n4195 DVDD.n4194 0.049839
R6328 DVDD.n3917 DVDD.n3916 0.049839
R6329 DVDD.n4202 DVDD.n3518 0.049839
R6330 DVDD.n230 DVDD.n225 0.0497891
R6331 DVDD.n230 DVDD.n218 0.0497891
R6332 DVDD.n5455 DVDD.n646 0.0497849
R6333 DVDD.n850 DVDD.n849 0.0497849
R6334 DVDD.n5745 DVDD.n188 0.0497849
R6335 DVDD.n5745 DVDD.n197 0.0497849
R6336 DVDD.n2229 DVDD.n2228 0.04955
R6337 DVDD.n1247 DVDD.n1246 0.04955
R6338 DVDD.n2453 DVDD.n2452 0.04955
R6339 DVDD.n1388 DVDD.n363 0.04955
R6340 DVDD.n1248 DVDD.n386 0.04955
R6341 DVDD.n5637 DVDD.n5636 0.04955
R6342 DVDD.n1390 DVDD.n902 0.04955
R6343 DVDD.n1241 DVDD.n925 0.04955
R6344 DVDD.n2954 DVDD.n2953 0.04955
R6345 DVDD.n2222 DVDD.n2221 0.04955
R6346 DVDD.n1242 DVDD.n1125 0.04955
R6347 DVDD.n2436 DVDD.n2435 0.04955
R6348 DVDD.n4123 DVDD.n4122 0.0491
R6349 DVDD.n4123 DVDD.n3547 0.0491
R6350 DVDD.n4127 DVDD.n3547 0.0491
R6351 DVDD.n4128 DVDD.n4127 0.0491
R6352 DVDD.n4129 DVDD.n4128 0.0491
R6353 DVDD.n4129 DVDD.n3545 0.0491
R6354 DVDD.n4133 DVDD.n3545 0.0491
R6355 DVDD.n4134 DVDD.n4133 0.0491
R6356 DVDD.n4135 DVDD.n4134 0.0491
R6357 DVDD.n4135 DVDD.n3543 0.0491
R6358 DVDD.n4139 DVDD.n3543 0.0491
R6359 DVDD.n4140 DVDD.n4139 0.0491
R6360 DVDD.n4141 DVDD.n4140 0.0491
R6361 DVDD.n4141 DVDD.n3541 0.0491
R6362 DVDD.n4145 DVDD.n3541 0.0491
R6363 DVDD.n4146 DVDD.n4145 0.0491
R6364 DVDD.n4147 DVDD.n4146 0.0491
R6365 DVDD.n4147 DVDD.n3539 0.0491
R6366 DVDD.n4151 DVDD.n3539 0.0491
R6367 DVDD.n4152 DVDD.n4151 0.0491
R6368 DVDD.n4152 DVDD.n3537 0.0491
R6369 DVDD.n4156 DVDD.n3537 0.0491
R6370 DVDD.n4157 DVDD.n4156 0.0491
R6371 DVDD.n4158 DVDD.n4157 0.0491
R6372 DVDD.n4158 DVDD.n3535 0.0491
R6373 DVDD.n4162 DVDD.n3535 0.0491
R6374 DVDD.n4163 DVDD.n4162 0.0491
R6375 DVDD.n4164 DVDD.n4163 0.0491
R6376 DVDD.n4164 DVDD.n3533 0.0491
R6377 DVDD.n4168 DVDD.n3533 0.0491
R6378 DVDD.n4169 DVDD.n4168 0.0491
R6379 DVDD.n4170 DVDD.n4169 0.0491
R6380 DVDD.n4170 DVDD.n3531 0.0491
R6381 DVDD.n4174 DVDD.n3531 0.0491
R6382 DVDD.n4175 DVDD.n4174 0.0491
R6383 DVDD.n4176 DVDD.n4175 0.0491
R6384 DVDD.n4176 DVDD.n3529 0.0491
R6385 DVDD.n4180 DVDD.n3529 0.0491
R6386 DVDD.n4181 DVDD.n4180 0.0491
R6387 DVDD DVDD.n3683 0.0491
R6388 DVDD.n3907 DVDD.n3683 0.0491
R6389 DVDD DVDD.n3680 0.0491
R6390 DVDD.n3910 DVDD.n3680 0.0491
R6391 DVDD.n3674 DVDD 0.0491
R6392 DVDD.n3678 DVDD.n3674 0.0491
R6393 DVDD DVDD.n3524 0.0491
R6394 DVDD.n4198 DVDD.n3524 0.0491
R6395 DVDD.n3858 DVDD.n3857 0.0491
R6396 DVDD.n3874 DVDD.n3873 0.0491
R6397 DVDD.n3880 DVDD.n3879 0.0491
R6398 DVDD.n3880 DVDD.n3854 0.0491
R6399 DVDD.n3884 DVDD.n3854 0.0491
R6400 DVDD.n3885 DVDD.n3884 0.0491
R6401 DVDD.n3886 DVDD.n3885 0.0491
R6402 DVDD.n3886 DVDD.n3852 0.0491
R6403 DVDD.n3891 DVDD.n3852 0.0491
R6404 DVDD.n3932 DVDD.n3931 0.0491
R6405 DVDD.n3954 DVDD.n3661 0.0491
R6406 DVDD.n3948 DVDD.n3947 0.0491
R6407 DVDD.n3947 DVDD.n3946 0.0491
R6408 DVDD.n3946 DVDD.n3664 0.0491
R6409 DVDD.n3942 DVDD.n3664 0.0491
R6410 DVDD.n3942 DVDD.n3941 0.0491
R6411 DVDD.n3941 DVDD.n3940 0.0491
R6412 DVDD.n3940 DVDD.n3919 0.0491
R6413 DVDD.n3762 DVDD.n3696 0.0491
R6414 DVDD.n3766 DVDD.n3696 0.0491
R6415 DVDD.n3767 DVDD.n3766 0.0491
R6416 DVDD.n3768 DVDD.n3767 0.0491
R6417 DVDD.n3768 DVDD.n3694 0.0491
R6418 DVDD.n3772 DVDD.n3694 0.0491
R6419 DVDD.n3773 DVDD.n3772 0.0491
R6420 DVDD.n3774 DVDD.n3773 0.0491
R6421 DVDD.n3774 DVDD.n3692 0.0491
R6422 DVDD.n3778 DVDD.n3692 0.0491
R6423 DVDD.n3779 DVDD.n3778 0.0491
R6424 DVDD.n3780 DVDD.n3779 0.0491
R6425 DVDD.n3780 DVDD.n3690 0.0491
R6426 DVDD.n3784 DVDD.n3690 0.0491
R6427 DVDD.n3785 DVDD.n3784 0.0491
R6428 DVDD.n3786 DVDD.n3785 0.0491
R6429 DVDD.n3786 DVDD.n3688 0.0491
R6430 DVDD.n3790 DVDD.n3688 0.0491
R6431 DVDD.n3791 DVDD.n3790 0.0491
R6432 DVDD.n3828 DVDD.n3791 0.0491
R6433 DVDD.n3828 DVDD.n3827 0.0491
R6434 DVDD.n3827 DVDD.n3826 0.0491
R6435 DVDD.n3826 DVDD.n3792 0.0491
R6436 DVDD.n3822 DVDD.n3792 0.0491
R6437 DVDD.n3822 DVDD.n3821 0.0491
R6438 DVDD.n3821 DVDD.n3820 0.0491
R6439 DVDD.n3820 DVDD.n3794 0.0491
R6440 DVDD.n3816 DVDD.n3794 0.0491
R6441 DVDD.n3816 DVDD.n3815 0.0491
R6442 DVDD.n3815 DVDD.n3814 0.0491
R6443 DVDD.n3814 DVDD.n3796 0.0491
R6444 DVDD.n3810 DVDD.n3796 0.0491
R6445 DVDD.n3810 DVDD.n3809 0.0491
R6446 DVDD.n3809 DVDD.n3808 0.0491
R6447 DVDD.n3808 DVDD.n3798 0.0491
R6448 DVDD.n3804 DVDD.n3798 0.0491
R6449 DVDD.n3804 DVDD.n3803 0.0491
R6450 DVDD.n3803 DVDD.n3802 0.0491
R6451 DVDD.n3802 DVDD.n3800 0.0491
R6452 DVDD.n2295 DVDD 0.0487259
R6453 DVDD DVDD.n1349 0.0487259
R6454 DVDD DVDD.n2259 0.0487259
R6455 DVDD.n1651 DVDD 0.0487259
R6456 DVDD.n5411 DVDD 0.0487259
R6457 DVDD.n2937 DVDD.n980 0.04865
R6458 DVDD.n2938 DVDD.n432 0.04865
R6459 DVDD.n2945 DVDD.n968 0.04865
R6460 DVDD.n2943 DVDD.n450 0.04865
R6461 DVDD.n5499 DVDD.n579 0.04775
R6462 DVDD.n5502 DVDD.n575 0.04775
R6463 DVDD.n5510 DVDD.n564 0.04775
R6464 DVDD.n5513 DVDD.n560 0.04775
R6465 DVDD.n5653 DVDD.n5652 0.047347
R6466 DVDD.n3870 DVDD.n3582 0.04685
R6467 DVDD.n3955 DVDD.n3660 0.04685
R6468 DVDD.n1531 DVDD.n1530 0.04595
R6469 DVDD.n1229 DVDD.n1228 0.04595
R6470 DVDD.n3860 DVDD.n3585 0.04595
R6471 DVDD.n1532 DVDD.n364 0.04595
R6472 DVDD.n1230 DVDD.n387 0.04595
R6473 DVDD.n3928 DVDD.n3657 0.04595
R6474 DVDD.n1525 DVDD.n903 0.04595
R6475 DVDD.n1223 DVDD.n926 0.04595
R6476 DVDD.n1526 DVDD.n1394 0.04595
R6477 DVDD.n1224 DVDD.n1126 0.04595
R6478 DVDD.n984 DVDD.n443 0.04505
R6479 DVDD.n3587 DVDD.n3576 0.04505
R6480 DVDD.n5630 DVDD.n431 0.04505
R6481 DVDD.n3934 DVDD.n3658 0.04505
R6482 DVDD.n967 DVDD.n445 0.04505
R6483 DVDD.n5624 DVDD.n446 0.04505
R6484 DVDD.n3936 DVDD.n3935 0.0449703
R6485 DVDD.n3855 DVDD.n3586 0.0449123
R6486 DVDD.n2604 DVDD.n2577 0.04415
R6487 DVDD.n3876 DVDD.n3580 0.04415
R6488 DVDD.n2756 DVDD.n2605 0.04415
R6489 DVDD.n3950 DVDD.n3653 0.04415
R6490 DVDD.n2761 DVDD.n480 0.04415
R6491 DVDD.n2763 DVDD.n2590 0.04415
R6492 DVDD.n5479 DVDD.n5478 0.0431316
R6493 DVDD.n1517 DVDD.n1516 0.04235
R6494 DVDD.n1518 DVDD.n365 0.04235
R6495 DVDD.n1511 DVDD.n904 0.04235
R6496 DVDD.n1512 DVDD.n1395 0.04235
R6497 DVDD.n997 DVDD.n983 0.04145
R6498 DVDD.n430 DVDD.n428 0.04145
R6499 DVDD.n1008 DVDD.n966 0.04145
R6500 DVDD.n463 DVDD.n449 0.04145
R6501 DVDD.n4845 DVDD.n4786 0.0407632
R6502 DVDD.n5807 DVDD.n169 0.0407632
R6503 DVDD.n4318 DVDD.n4216 0.0407632
R6504 DVDD.n28 DVDD.n27 0.0407632
R6505 DVDD.n2372 DVDD.n1210 0.0406306
R6506 DVDD.n5498 DVDD.n577 0.04055
R6507 DVDD.n2922 DVDD.n2576 0.04055
R6508 DVDD.n576 DVDD.n573 0.04055
R6509 DVDD.n2608 DVDD.n2584 0.04055
R6510 DVDD.n565 DVDD.n562 0.04055
R6511 DVDD.n2586 DVDD.n479 0.04055
R6512 DVDD.n561 DVDD.n558 0.04055
R6513 DVDD.n2916 DVDD.n2587 0.04055
R6514 DVDD.n3868 DVDD.n3579 0.03965
R6515 DVDD.n3920 DVDD.n3649 0.03965
R6516 DVDD.n1713 DVDD.n1712 0.03875
R6517 DVDD.n1503 DVDD.n1502 0.03875
R6518 DVDD.n3862 DVDD.n3577 0.03875
R6519 DVDD.n2046 DVDD.n1593 0.03875
R6520 DVDD.n1504 DVDD.n366 0.03875
R6521 DVDD.n3926 DVDD.n3652 0.03875
R6522 DVDD.n2039 DVDD.n2038 0.03875
R6523 DVDD.n1497 DVDD.n905 0.03875
R6524 DVDD.n2040 DVDD.n883 0.03875
R6525 DVDD.n1498 DVDD.n1396 0.03875
R6526 DVDD.n5280 DVDD.n616 0.037944
R6527 DVDD DVDD.t162 0.0375588
R6528 DVDD DVDD.t156 0.0375588
R6529 DVDD DVDD.t159 0.0375588
R6530 DVDD DVDD.t160 0.0375588
R6531 DVDD.n3879 DVDD.n3581 0.03695
R6532 DVDD.n3948 DVDD.n3655 0.03695
R6533 DVDD.n4846 DVDD.n4842 0.0360263
R6534 DVDD.n5810 DVDD.n5809 0.0360263
R6535 DVDD.n4319 DVDD.n4217 0.0360263
R6536 DVDD.n5983 DVDD.n5982 0.0360263
R6537 DVDD.n1733 DVDD.n1732 0.03515
R6538 DVDD.n1489 DVDD.n1488 0.03515
R6539 DVDD.n1734 DVDD.n1594 0.03515
R6540 DVDD.n1490 DVDD.n367 0.03515
R6541 DVDD.n1741 DVDD.n1718 0.03515
R6542 DVDD.n1483 DVDD.n906 0.03515
R6543 DVDD.n1739 DVDD.n884 0.03515
R6544 DVDD.n1484 DVDD.n1397 0.03515
R6545 DVDD.n5567 DVDD.n5566 0.0349216
R6546 DVDD.n1855 DVDD.n1854 0.0336863
R6547 DVDD.n1777 DVDD.n1775 0.0336863
R6548 DVDD.n1781 DVDD.n1780 0.0336863
R6549 DVDD.n828 DVDD.n787 0.0336863
R6550 DVDD.n3847 DVDD.n3846 0.0336579
R6551 DVDD.n3844 DVDD.n3843 0.0336579
R6552 DVDD.n599 DVDD.n598 0.03335
R6553 DVDD.n1700 DVDD.n1596 0.03335
R6554 DVDD.n2027 DVDD.n1720 0.03335
R6555 DVDD.n1789 DVDD.n886 0.03335
R6556 DVDD.n5520 DVDD.t113 0.03326
R6557 DVDD.n5520 DVDD.t110 0.03326
R6558 DVDD.n1730 DVDD.t153 0.03326
R6559 DVDD.n1730 DVDD.t99 0.03326
R6560 DVDD.n2043 DVDD.t150 0.03326
R6561 DVDD.n2043 DVDD.t106 0.03326
R6562 DVDD.n5650 DVDD.t139 0.03326
R6563 DVDD.n5650 DVDD.t128 0.03326
R6564 DVDD.n1492 DVDD.t89 0.03326
R6565 DVDD.n1492 DVDD.t77 0.03326
R6566 DVDD.n1506 DVDD.t136 0.03326
R6567 DVDD.n1506 DVDD.t92 0.03326
R6568 DVDD.n1520 DVDD.t146 0.03326
R6569 DVDD.n1520 DVDD.t145 0.03326
R6570 DVDD.n1534 DVDD.t135 0.03326
R6571 DVDD.n1534 DVDD.t104 0.03326
R6572 DVDD.n2225 DVDD.t130 0.03326
R6573 DVDD.n2225 DVDD.t147 0.03326
R6574 DVDD.n1550 DVDD.t100 0.03326
R6575 DVDD.n1550 DVDD.t144 0.03326
R6576 DVDD.n1232 DVDD.t112 0.03326
R6577 DVDD.n1232 DVDD.t132 0.03326
R6578 DVDD.n1250 DVDD.t126 0.03326
R6579 DVDD.n1250 DVDD.t78 0.03326
R6580 DVDD.n2446 DVDD.t98 0.03326
R6581 DVDD.n2446 DVDD.t111 0.03326
R6582 DVDD.n1262 DVDD.t76 0.03326
R6583 DVDD.n1262 DVDD.t90 0.03326
R6584 DVDD.n1208 DVDD.t119 0.03326
R6585 DVDD.n1208 DVDD.t151 0.03326
R6586 DVDD.n2524 DVDD.t96 0.03326
R6587 DVDD.n2524 DVDD.t140 0.03326
R6588 DVDD.n2539 DVDD.t109 0.03326
R6589 DVDD.n2539 DVDD.t83 0.03326
R6590 DVDD.n2557 DVDD.t97 0.03326
R6591 DVDD.n2557 DVDD.t107 0.03326
R6592 DVDD.n977 DVDD.t131 0.03326
R6593 DVDD.n977 DVDD.t141 0.03326
R6594 DVDD.n5627 DVDD.t117 0.03326
R6595 DVDD.n5627 DVDD.t118 0.03326
R6596 DVDD.n1012 DVDD.t143 0.03326
R6597 DVDD.n1012 DVDD.t86 0.03326
R6598 DVDD.n2566 DVDD.t142 0.03326
R6599 DVDD.n2566 DVDD.t124 0.03326
R6600 DVDD.n2571 DVDD.t133 0.03326
R6601 DVDD.n2571 DVDD.t85 0.03326
R6602 DVDD.n2594 DVDD.t103 0.03326
R6603 DVDD.n2594 DVDD.t87 0.03326
R6604 DVDD.n2919 DVDD.t80 0.03326
R6605 DVDD.n2919 DVDD.t91 0.03326
R6606 DVDD.n5564 DVDD.t120 0.03326
R6607 DVDD.n5564 DVDD.t95 0.03326
R6608 DVDD.n2767 DVDD.t79 0.03326
R6609 DVDD.n2767 DVDD.t94 0.03326
R6610 DVDD.n2784 DVDD.t122 0.03326
R6611 DVDD.n2784 DVDD.t105 0.03326
R6612 DVDD.n2788 DVDD.t101 0.03326
R6613 DVDD.n2788 DVDD.t102 0.03326
R6614 DVDD.n2792 DVDD.t93 0.03326
R6615 DVDD.n2792 DVDD.t148 0.03326
R6616 DVDD.n2796 DVDD.t82 0.03326
R6617 DVDD.n2796 DVDD.t114 0.03326
R6618 DVDD.n2800 DVDD.t121 0.03326
R6619 DVDD.n2800 DVDD.t152 0.03326
R6620 DVDD.n2804 DVDD.t125 0.03326
R6621 DVDD.n2804 DVDD.t154 0.03326
R6622 DVDD.n2808 DVDD.t116 0.03326
R6623 DVDD.n2808 DVDD.t134 0.03326
R6624 DVDD.n2812 DVDD.t127 0.03326
R6625 DVDD.n2812 DVDD.t149 0.03326
R6626 DVDD.n2816 DVDD.t115 0.03326
R6627 DVDD.n2816 DVDD.t138 0.03326
R6628 DVDD.n2820 DVDD.t84 0.03326
R6629 DVDD.n2820 DVDD.t81 0.03326
R6630 DVDD.n2824 DVDD.t88 0.03326
R6631 DVDD.n2824 DVDD.t123 0.03326
R6632 DVDD.n2782 DVDD.t75 0.03326
R6633 DVDD.n2782 DVDD.t129 0.03326
R6634 DVDD.n2843 DVDD.t137 0.03326
R6635 DVDD.n2843 DVDD.t108 0.03326
R6636 DVDD.n1857 DVDD.n1856 0.0332409
R6637 DVDD.n5029 DVDD.n5013 0.03245
R6638 DVDD.n5029 DVDD.n5011 0.03245
R6639 DVDD.n5034 DVDD.n5011 0.03245
R6640 DVDD.n5664 DVDD.n302 0.03245
R6641 DVDD.n5664 DVDD.n303 0.03245
R6642 DVDD.n5660 DVDD.n303 0.03245
R6643 DVDD.n5751 DVDD.n5750 0.03245
R6644 DVDD.n5750 DVDD.n183 0.03245
R6645 DVDD.n5746 DVDD.n183 0.03245
R6646 DVDD.n5316 DVDD.n200 0.03245
R6647 DVDD.n5316 DVDD.n4906 0.03245
R6648 DVDD.n5312 DVDD.n4906 0.03245
R6649 DVDD.n5304 DVDD.n5303 0.03245
R6650 DVDD.n5303 DVDD.n5300 0.03245
R6651 DVDD.n5300 DVDD.n5299 0.03245
R6652 DVDD.n5291 DVDD.n4927 0.03245
R6653 DVDD.n5291 DVDD.n4928 0.03245
R6654 DVDD.n5287 DVDD.n4928 0.03245
R6655 DVDD.n4532 DVDD.n4531 0.03245
R6656 DVDD.n4531 DVDD.n4528 0.03245
R6657 DVDD.n4528 DVDD.n3171 0.03245
R6658 DVDD.n3170 DVDD.n3144 0.03245
R6659 DVDD.n4879 DVDD.n3144 0.03245
R6660 DVDD.n4879 DVDD.n3142 0.03245
R6661 DVDD.n3866 DVDD.n3583 0.03245
R6662 DVDD.n3922 DVDD.n3659 0.03245
R6663 DVDD.n1371 DVDD.n359 0.03155
R6664 DVDD.n3864 DVDD.n3584 0.03155
R6665 DVDD.n5648 DVDD.n5647 0.03155
R6666 DVDD.n3924 DVDD.n3656 0.03155
R6667 DVDD.n2965 DVDD.n2964 0.03155
R6668 DVDD.n2967 DVDD.n898 0.03155
R6669 DVDD.n1856 DVDD.n1773 0.0309017
R6670 DVDD.n1854 DVDD.n1853 0.0304416
R6671 DVDD.n1849 DVDD.n1777 0.0304416
R6672 DVDD.n1848 DVDD.n1781 0.0304416
R6673 DVDD.n787 DVDD.n786 0.0304416
R6674 DVDD.n4206 DVDD.n4205 0.0296033
R6675 DVDD.n4185 DVDD.n4184 0.0296033
R6676 DVDD.n4116 DVDD.n3551 0.0287281
R6677 DVDD.n3554 DVDD.n3550 0.0287281
R6678 DVDD.n26 DVDD.n18 0.0287281
R6679 DVDD.n5388 DVDD.n606 0.0287281
R6680 DVDD.n5496 DVDD.n5495 0.0287281
R6681 DVDD.n600 DVDD.n579 0.0287281
R6682 DVDD.n1731 DVDD.n587 0.0287281
R6683 DVDD.n1711 DVDD.n584 0.0287281
R6684 DVDD.n583 DVDD.n582 0.0287281
R6685 DVDD.n1487 DVDD.n1374 0.0287281
R6686 DVDD.n1501 DVDD.n1377 0.0287281
R6687 DVDD.n1515 DVDD.n1380 0.0287281
R6688 DVDD.n1529 DVDD.n1383 0.0287281
R6689 DVDD.n1387 DVDD.n1386 0.0287281
R6690 DVDD.n2235 DVDD.n2233 0.0287281
R6691 DVDD.n1227 DVDD.n1101 0.0287281
R6692 DVDD.n1245 DVDD.n1112 0.0287281
R6693 DVDD.n1117 DVDD.n1115 0.0287281
R6694 DVDD.n2519 DVDD.n990 0.0287281
R6695 DVDD.n2553 DVDD.n985 0.0287281
R6696 DVDD.n2926 DVDD.n2577 0.0287281
R6697 DVDD.n2924 DVDD.n2576 0.0287281
R6698 DVDD.n2923 DVDD.n2582 0.0287281
R6699 DVDD.n2929 DVDD.n2928 0.0287281
R6700 DVDD.n5368 DVDD.n5367 0.0287281
R6701 DVDD.n5484 DVDD.n5483 0.0287281
R6702 DVDD.n5494 DVDD.n5493 0.0287281
R6703 DVDD.n597 DVDD.n596 0.0287281
R6704 DVDD.n1732 DVDD.n586 0.0287281
R6705 DVDD.n1712 DVDD.n583 0.0287281
R6706 DVDD.n1372 DVDD.n1371 0.0287281
R6707 DVDD.n1488 DVDD.n1375 0.0287281
R6708 DVDD.n1502 DVDD.n1378 0.0287281
R6709 DVDD.n1516 DVDD.n1381 0.0287281
R6710 DVDD.n1530 DVDD.n1384 0.0287281
R6711 DVDD.n2230 DVDD.n2229 0.0287281
R6712 DVDD.n2231 DVDD.n1101 0.0287281
R6713 DVDD.n1228 DVDD.n1102 0.0287281
R6714 DVDD.n1246 DVDD.n1113 0.0287281
R6715 DVDD.n2451 DVDD.n2450 0.0287281
R6716 DVDD.n1116 DVDD.n1099 0.0287281
R6717 DVDD.n1259 DVDD.n1098 0.0287281
R6718 DVDD.n2455 DVDD.n2454 0.0287281
R6719 DVDD.n2452 DVDD.n989 0.0287281
R6720 DVDD.n2520 DVDD.n991 0.0287281
R6721 DVDD.n1002 DVDD.n987 0.0287281
R6722 DVDD.n2535 DVDD.n986 0.0287281
R6723 DVDD.n999 DVDD.n992 0.0287281
R6724 DVDD.n1003 DVDD.n980 0.0287281
R6725 DVDD.n2936 DVDD.n981 0.0287281
R6726 DVDD.n1004 DVDD.n984 0.0287281
R6727 DVDD.n998 DVDD.n995 0.0287281
R6728 DVDD.n1005 DVDD.n983 0.0287281
R6729 DVDD.n2931 DVDD.n2574 0.0287281
R6730 DVDD.n2925 DVDD.n2580 0.0287281
R6731 DVDD.n4187 DVDD.n3425 0.0287281
R6732 DVDD.n5154 DVDD.n626 0.0287281
R6733 DVDD.n1706 DVDD.n1606 0.0287281
R6734 DVDD.n2047 DVDD.n1710 0.0287281
R6735 DVDD.n1708 DVDD.n360 0.0287281
R6736 DVDD.n2068 DVDD.n370 0.0287281
R6737 DVDD.n2070 DVDD.n372 0.0287281
R6738 DVDD.n2072 DVDD.n374 0.0287281
R6739 DVDD.n2074 DVDD.n376 0.0287281
R6740 DVDD.n2076 DVDD.n378 0.0287281
R6741 DVDD.n5645 DVDD.n380 0.0287281
R6742 DVDD.n389 DVDD.n382 0.0287281
R6743 DVDD.n407 DVDD.n395 0.0287281
R6744 DVDD.n409 DVDD.n397 0.0287281
R6745 DVDD.n437 DVDD.n422 0.0287281
R6746 DVDD.n433 DVDD.n417 0.0287281
R6747 DVDD.n2753 DVDD.n527 0.0287281
R6748 DVDD.n5202 DVDD.n5142 0.0287281
R6749 DVDD.n5470 DVDD.n627 0.0287281
R6750 DVDD.n1597 DVDD.n629 0.0287281
R6751 DVDD.n1698 DVDD.n1598 0.0287281
R6752 DVDD.n1601 DVDD.n575 0.0287281
R6753 DVDD.n1701 DVDD.n1595 0.0287281
R6754 DVDD.n1707 DVDD.n1594 0.0287281
R6755 DVDD.n1708 DVDD.n1593 0.0287281
R6756 DVDD.n5647 DVDD.n361 0.0287281
R6757 DVDD.n2069 DVDD.n367 0.0287281
R6758 DVDD.n2071 DVDD.n366 0.0287281
R6759 DVDD.n2073 DVDD.n365 0.0287281
R6760 DVDD.n2075 DVDD.n364 0.0287281
R6761 DVDD.n2077 DVDD.n363 0.0287281
R6762 DVDD.n5643 DVDD.n382 0.0287281
R6763 DVDD.n402 DVDD.n387 0.0287281
R6764 DVDD.n408 DVDD.n386 0.0287281
R6765 DVDD.n410 DVDD.n385 0.0287281
R6766 DVDD.n400 DVDD.n398 0.0287281
R6767 DVDD.n5641 DVDD.n5640 0.0287281
R6768 DVDD.n5638 DVDD.n384 0.0287281
R6769 DVDD.n5636 DVDD.n412 0.0287281
R6770 DVDD.n438 DVDD.n419 0.0287281
R6771 DVDD.n435 DVDD.n423 0.0287281
R6772 DVDD.n434 DVDD.n424 0.0287281
R6773 DVDD.n439 DVDD.n416 0.0287281
R6774 DVDD.n432 DVDD.n425 0.0287281
R6775 DVDD.n441 DVDD.n415 0.0287281
R6776 DVDD.n431 DVDD.n426 0.0287281
R6777 DVDD.n5631 DVDD.n414 0.0287281
R6778 DVDD.n430 DVDD.n427 0.0287281
R6779 DVDD.n2748 DVDD.n2611 0.0287281
R6780 DVDD.n2749 DVDD.n2605 0.0287281
R6781 DVDD.n2755 DVDD.n2606 0.0287281
R6782 DVDD.n2750 DVDD.n2608 0.0287281
R6783 DVDD.n2752 DVDD.n2614 0.0287281
R6784 DVDD.n3511 DVDD.n3375 0.0287281
R6785 DVDD.n757 DVDD.n261 0.0287281
R6786 DVDD.n2033 DVDD.n1742 0.0287281
R6787 DVDD.n1743 DVDD.n1715 0.0287281
R6788 DVDD.n1716 DVDD.n899 0.0287281
R6789 DVDD.n1436 DVDD.n909 0.0287281
R6790 DVDD.n1438 DVDD.n911 0.0287281
R6791 DVDD.n1440 DVDD.n913 0.0287281
R6792 DVDD.n1442 DVDD.n915 0.0287281
R6793 DVDD.n1444 DVDD.n917 0.0287281
R6794 DVDD.n2962 DVDD.n919 0.0287281
R6795 DVDD.n928 DVDD.n921 0.0287281
R6796 DVDD.n946 DVDD.n934 0.0287281
R6797 DVDD.n948 DVDD.n936 0.0287281
R6798 DVDD.n973 DVDD.n961 0.0287281
R6799 DVDD.n969 DVDD.n956 0.0287281
R6800 DVDD.n5614 DVDD.n486 0.0287281
R6801 DVDD.n3041 DVDD.n744 0.0287281
R6802 DVDD.n5704 DVDD.n262 0.0287281
R6803 DVDD.n1721 DVDD.n264 0.0287281
R6804 DVDD.n2025 DVDD.n1722 0.0287281
R6805 DVDD.n1725 DVDD.n564 0.0287281
R6806 DVDD.n2028 DVDD.n1719 0.0287281
R6807 DVDD.n2035 DVDD.n1718 0.0287281
R6808 DVDD.n2038 DVDD.n1716 0.0287281
R6809 DVDD.n2964 DVDD.n900 0.0287281
R6810 DVDD.n1437 DVDD.n906 0.0287281
R6811 DVDD.n1439 DVDD.n905 0.0287281
R6812 DVDD.n1441 DVDD.n904 0.0287281
R6813 DVDD.n1443 DVDD.n903 0.0287281
R6814 DVDD.n1445 DVDD.n902 0.0287281
R6815 DVDD.n2960 DVDD.n921 0.0287281
R6816 DVDD.n941 DVDD.n926 0.0287281
R6817 DVDD.n947 DVDD.n925 0.0287281
R6818 DVDD.n949 DVDD.n924 0.0287281
R6819 DVDD.n939 DVDD.n937 0.0287281
R6820 DVDD.n2958 DVDD.n2957 0.0287281
R6821 DVDD.n2955 DVDD.n923 0.0287281
R6822 DVDD.n2953 DVDD.n951 0.0287281
R6823 DVDD.n974 DVDD.n958 0.0287281
R6824 DVDD.n971 DVDD.n962 0.0287281
R6825 DVDD.n970 DVDD.n963 0.0287281
R6826 DVDD.n975 DVDD.n955 0.0287281
R6827 DVDD.n968 DVDD.n964 0.0287281
R6828 DVDD.n2946 DVDD.n954 0.0287281
R6829 DVDD.n967 DVDD.n965 0.0287281
R6830 DVDD.n2948 DVDD.n953 0.0287281
R6831 DVDD.n2951 DVDD.n966 0.0287281
R6832 DVDD.n5616 DVDD.n477 0.0287281
R6833 DVDD.n5610 DVDD.n480 0.0287281
R6834 DVDD.n5609 DVDD.n483 0.0287281
R6835 DVDD.n5611 DVDD.n479 0.0287281
R6836 DVDD.n5613 DVDD.n485 0.0287281
R6837 DVDD.n3746 DVDD.n3698 0.0287281
R6838 DVDD.n4215 DVDD.n3506 0.0287281
R6839 DVDD.n5712 DVDD.n255 0.0287281
R6840 DVDD.n1795 DVDD.n894 0.0287281
R6841 DVDD.n1797 DVDD.n896 0.0287281
R6842 DVDD.n2968 DVDD.n897 0.0287281
R6843 DVDD.n2207 DVDD.n1400 0.0287281
R6844 DVDD.n2209 DVDD.n1402 0.0287281
R6845 DVDD.n2211 DVDD.n1404 0.0287281
R6846 DVDD.n2213 DVDD.n1406 0.0287281
R6847 DVDD.n2215 DVDD.n1391 0.0287281
R6848 DVDD.n2219 DVDD.n2217 0.0287281
R6849 DVDD.n2426 DVDD.n1129 0.0287281
R6850 DVDD.n2432 DVDD.n1135 0.0287281
R6851 DVDD.n2434 DVDD.n1121 0.0287281
R6852 DVDD.n2514 DVDD.n456 0.0287281
R6853 DVDD.n2549 DVDD.n451 0.0287281
R6854 DVDD.n2913 DVDD.n2912 0.0287281
R6855 DVDD.n3756 DVDD.n3755 0.0287281
R6856 DVDD.n5714 DVDD.n241 0.0287281
R6857 DVDD.n838 DVDD.n256 0.0287281
R6858 DVDD.n2971 DVDD.n829 0.0287281
R6859 DVDD.n2970 DVDD.n881 0.0287281
R6860 DVDD.n889 DVDD.n560 0.0287281
R6861 DVDD.n1790 DVDD.n885 0.0287281
R6862 DVDD.n1796 DVDD.n884 0.0287281
R6863 DVDD.n897 DVDD.n883 0.0287281
R6864 DVDD.n2206 DVDD.n898 0.0287281
R6865 DVDD.n2208 DVDD.n1397 0.0287281
R6866 DVDD.n2210 DVDD.n1396 0.0287281
R6867 DVDD.n2212 DVDD.n1395 0.0287281
R6868 DVDD.n2214 DVDD.n1394 0.0287281
R6869 DVDD.n2221 DVDD.n1392 0.0287281
R6870 DVDD.n2426 DVDD.n1127 0.0287281
R6871 DVDD.n2427 DVDD.n1126 0.0287281
R6872 DVDD.n2433 DVDD.n1125 0.0287281
R6873 DVDD.n2442 DVDD.n1122 0.0287281
R6874 DVDD.n1139 DVDD.n1137 0.0287281
R6875 DVDD.n2440 DVDD.n2439 0.0287281
R6876 DVDD.n2437 DVDD.n1124 0.0287281
R6877 DVDD.n2435 DVDD.n455 0.0287281
R6878 DVDD.n2515 DVDD.n457 0.0287281
R6879 DVDD.n468 DVDD.n453 0.0287281
R6880 DVDD.n2531 DVDD.n452 0.0287281
R6881 DVDD.n465 DVDD.n458 0.0287281
R6882 DVDD.n469 DVDD.n450 0.0287281
R6883 DVDD.n464 DVDD.n460 0.0287281
R6884 DVDD.n470 DVDD.n446 0.0287281
R6885 DVDD.n5623 DVDD.n447 0.0287281
R6886 DVDD.n471 DVDD.n449 0.0287281
R6887 DVDD.n2908 DVDD.n2592 0.0287281
R6888 DVDD.n2909 DVDD.n2590 0.0287281
R6889 DVDD.n2907 DVDD.n2764 0.0287281
R6890 DVDD.n2910 DVDD.n2587 0.0287281
R6891 DVDD.n2915 DVDD.n2588 0.0287281
R6892 DVDD.n4213 DVDD.n4208 0.0287281
R6893 DVDD.n4210 DVDD.n3504 0.0287281
R6894 DVDD.n4321 DVDD.n4209 0.0287281
R6895 DVDD.n3516 DVDD.n3515 0.0287281
R6896 DVDD.n4690 DVDD.n4689 0.0287281
R6897 DVDD.n4686 DVDD.n4685 0.0287281
R6898 DVDD.n4192 DVDD.n4191 0.0287281
R6899 DVDD.n4539 DVDD.n4538 0.0287281
R6900 DVDD.n4543 DVDD.n4542 0.0287281
R6901 DVDD.n22 DVDD.n21 0.0287281
R6902 DVDD.n3184 DVDD.n25 0.0287281
R6903 DVDD.n5986 DVDD.n5985 0.0287281
R6904 DVDD.n5020 DVDD.n5018 0.0284
R6905 DVDD.n5658 DVDD.n307 0.0284
R6906 DVDD.n4505 DVDD.n4497 0.0284
R6907 DVDD.n4882 DVDD.n3141 0.0284
R6908 DVDD.n5754 DVDD.n5753 0.0284
R6909 DVDD.n5310 DVDD.n4910 0.0284
R6910 DVDD.n5109 DVDD.n4917 0.0284
R6911 DVDD.n5285 DVDD.n4929 0.0284
R6912 DVDD.n5019 DVDD.n5014 0.027725
R6913 DVDD.n4877 DVDD.n3146 0.027725
R6914 DVDD.n5752 DVDD.n181 0.027725
R6915 DVDD.n5286 DVDD.n4931 0.027725
R6916 DVDD.n5659 DVDD.n305 0.027275
R6917 DVDD.n4534 DVDD.n4533 0.027275
R6918 DVDD.n5311 DVDD.n4908 0.027275
R6919 DVDD.n5306 DVDD.n5305 0.027275
R6920 DVDD.n3764 DVDD.n3763 0.026913
R6921 DVDD.n3765 DVDD.n3764 0.026913
R6922 DVDD.n3765 DVDD.n3695 0.026913
R6923 DVDD.n3769 DVDD.n3695 0.026913
R6924 DVDD.n3770 DVDD.n3769 0.026913
R6925 DVDD.n3771 DVDD.n3770 0.026913
R6926 DVDD.n3771 DVDD.n3693 0.026913
R6927 DVDD.n3775 DVDD.n3693 0.026913
R6928 DVDD.n3776 DVDD.n3775 0.026913
R6929 DVDD.n3777 DVDD.n3776 0.026913
R6930 DVDD.n3777 DVDD.n3691 0.026913
R6931 DVDD.n3781 DVDD.n3691 0.026913
R6932 DVDD.n3782 DVDD.n3781 0.026913
R6933 DVDD.n3783 DVDD.n3782 0.026913
R6934 DVDD.n3783 DVDD.n3689 0.026913
R6935 DVDD.n3787 DVDD.n3689 0.026913
R6936 DVDD.n3788 DVDD.n3787 0.026913
R6937 DVDD.n3789 DVDD.n3788 0.026913
R6938 DVDD.n3789 DVDD.n3686 0.026913
R6939 DVDD.n3829 DVDD.n3687 0.026913
R6940 DVDD.n3825 DVDD.n3687 0.026913
R6941 DVDD.n3825 DVDD.n3824 0.026913
R6942 DVDD.n3824 DVDD.n3823 0.026913
R6943 DVDD.n3823 DVDD.n3793 0.026913
R6944 DVDD.n3819 DVDD.n3793 0.026913
R6945 DVDD.n3819 DVDD.n3818 0.026913
R6946 DVDD.n3818 DVDD.n3817 0.026913
R6947 DVDD.n3817 DVDD.n3795 0.026913
R6948 DVDD.n3813 DVDD.n3795 0.026913
R6949 DVDD.n3813 DVDD.n3812 0.026913
R6950 DVDD.n3812 DVDD.n3811 0.026913
R6951 DVDD.n3811 DVDD.n3797 0.026913
R6952 DVDD.n3807 DVDD.n3797 0.026913
R6953 DVDD.n3807 DVDD.n3806 0.026913
R6954 DVDD.n3806 DVDD.n3805 0.026913
R6955 DVDD.n3805 DVDD.n3799 0.026913
R6956 DVDD.n3801 DVDD.n3799 0.026913
R6957 DVDD.n3801 DVDD.n3509 0.026913
R6958 DVDD.n3667 DVDD.n3666 0.026913
R6959 DVDD.n3895 DVDD.n3847 0.026913
R6960 DVDD.n3900 DVDD.n3848 0.026913
R6961 DVDD.n3894 DVDD.n3893 0.026913
R6962 DVDD.n4124 DVDD.n3548 0.026913
R6963 DVDD.n4125 DVDD.n4124 0.026913
R6964 DVDD.n4126 DVDD.n4125 0.026913
R6965 DVDD.n4126 DVDD.n3546 0.026913
R6966 DVDD.n4130 DVDD.n3546 0.026913
R6967 DVDD.n4131 DVDD.n4130 0.026913
R6968 DVDD.n4132 DVDD.n4131 0.026913
R6969 DVDD.n4132 DVDD.n3544 0.026913
R6970 DVDD.n4136 DVDD.n3544 0.026913
R6971 DVDD.n4137 DVDD.n4136 0.026913
R6972 DVDD.n4138 DVDD.n4137 0.026913
R6973 DVDD.n4138 DVDD.n3542 0.026913
R6974 DVDD.n4142 DVDD.n3542 0.026913
R6975 DVDD.n4143 DVDD.n4142 0.026913
R6976 DVDD.n4144 DVDD.n4143 0.026913
R6977 DVDD.n4144 DVDD.n3540 0.026913
R6978 DVDD.n4148 DVDD.n3540 0.026913
R6979 DVDD.n4149 DVDD.n4148 0.026913
R6980 DVDD.n4150 DVDD.n4149 0.026913
R6981 DVDD.n4154 DVDD.n4153 0.026913
R6982 DVDD.n4155 DVDD.n4154 0.026913
R6983 DVDD.n4155 DVDD.n3536 0.026913
R6984 DVDD.n4159 DVDD.n3536 0.026913
R6985 DVDD.n4160 DVDD.n4159 0.026913
R6986 DVDD.n4161 DVDD.n4160 0.026913
R6987 DVDD.n4161 DVDD.n3534 0.026913
R6988 DVDD.n4165 DVDD.n3534 0.026913
R6989 DVDD.n4166 DVDD.n4165 0.026913
R6990 DVDD.n4167 DVDD.n4166 0.026913
R6991 DVDD.n4167 DVDD.n3532 0.026913
R6992 DVDD.n4171 DVDD.n3532 0.026913
R6993 DVDD.n4172 DVDD.n4171 0.026913
R6994 DVDD.n4173 DVDD.n4172 0.026913
R6995 DVDD.n4173 DVDD.n3530 0.026913
R6996 DVDD.n4177 DVDD.n3530 0.026913
R6997 DVDD.n4178 DVDD.n4177 0.026913
R6998 DVDD.n4179 DVDD.n4178 0.026913
R6999 DVDD.n4179 DVDD.n3528 0.026913
R7000 DVDD.n4204 DVDD.n3510 0.026913
R7001 DVDD.n3841 DVDD.n3837 0.026913
R7002 DVDD.n4186 DVDD.n3527 0.026913
R7003 DVDD.n5526 DVDD.n547 0.026913
R7004 DVDD.n551 DVDD.n543 0.026913
R7005 DVDD.n4212 DVDD.n4211 0.0262333
R7006 DVDD.n3704 DVDD.n3702 0.0262332
R7007 DVDD.n2906 DVDD.n2905 0.026229
R7008 DVDD.n230 DVDD.n226 0.0255962
R7009 DVDD.n4861 DVDD.n3153 0.0255962
R7010 DVDD.n5745 DVDD.n187 0.0255952
R7011 DVDD.n804 DVDD.n803 0.0255952
R7012 DVDD.n306 DVDD.n301 0.025475
R7013 DVDD.n4499 DVDD.n4498 0.025475
R7014 DVDD.n4909 DVDD.n4905 0.025475
R7015 DVDD.n4920 DVDD.n4918 0.025475
R7016 DVDD.n571 DVDD.n545 0.0253032
R7017 DVDD.n5527 DVDD.n5526 0.0253032
R7018 DVDD.n3864 DVDD.n3578 0.02525
R7019 DVDD.n3924 DVDD.n3650 0.02525
R7020 DVDD.n3851 DVDD.n3682 0.0251695
R7021 DVDD.n4194 DVDD.n4193 0.0251695
R7022 DVDD.n3892 DVDD.n3850 0.0251695
R7023 DVDD.n4196 DVDD.n4195 0.0251695
R7024 DVDD.n4200 DVDD.n3520 0.0251695
R7025 DVDD DVDD.n3522 0.0251695
R7026 DVDD.n3676 DVDD.n3673 0.0251695
R7027 DVDD.n3675 DVDD 0.0251695
R7028 DVDD.n3912 DVDD.n3669 0.0251695
R7029 DVDD DVDD.n3671 0.0251695
R7030 DVDD.n3904 DVDD.n3668 0.0251695
R7031 DVDD.n3905 DVDD 0.0251695
R7032 DVDD.n3916 DVDD.n3915 0.0251695
R7033 DVDD.n3518 DVDD.n3517 0.0251695
R7034 DVDD.n4203 DVDD.n4202 0.0251695
R7035 DVDD.n3918 DVDD.n3917 0.0251695
R7036 DVDD.n4861 DVDD.n3154 0.0249058
R7037 DVDD.n230 DVDD.n227 0.0247655
R7038 DVDD.n803 DVDD.n801 0.0247646
R7039 DVDD.n5745 DVDD.n186 0.0247619
R7040 DVDD.n3866 DVDD.n3578 0.02435
R7041 DVDD.n3922 DVDD.n3650 0.02435
R7042 DVDD.n5028 DVDD.n5027 0.023675
R7043 DVDD.n4878 DVDD.n3145 0.023675
R7044 DVDD.n4899 DVDD.n182 0.023675
R7045 DVDD.n4930 DVDD.n4926 0.023675
R7046 DVDD.n598 DVDD.n597 0.02345
R7047 DVDD.n1701 DVDD.n1700 0.02345
R7048 DVDD.n2028 DVDD.n2027 0.02345
R7049 DVDD.n1790 DVDD.n1789 0.02345
R7050 DVDD.n4861 DVDD.n3162 0.0229382
R7051 DVDD.n673 DVDD.n672 0.0227712
R7052 DVDD.n230 DVDD.n214 0.0227712
R7053 DVDD.n5745 DVDD.n195 0.0227712
R7054 DVDD.n5017 DVDD.n616 0.0224963
R7055 DVDD.n674 DVDD 0.022387
R7056 DVDD.n5959 DVDD 0.0218158
R7057 DVDD.n5031 DVDD.n5030 0.0218
R7058 DVDD.n5033 DVDD.n5031 0.0218
R7059 DVDD.n5663 DVDD.n304 0.0218
R7060 DVDD.n5663 DVDD.n5662 0.0218
R7061 DVDD.n5749 DVDD.n5748 0.0218
R7062 DVDD.n5748 DVDD.n5747 0.0218
R7063 DVDD.n5315 DVDD.n4907 0.0218
R7064 DVDD.n5315 DVDD.n5314 0.0218
R7065 DVDD.n5302 DVDD.n5301 0.0218
R7066 DVDD.n5301 DVDD.n223 0.0218
R7067 DVDD.n5290 DVDD.n222 0.0218
R7068 DVDD.n5290 DVDD.n5289 0.0218
R7069 DVDD.n4530 DVDD.n4529 0.0218
R7070 DVDD.n4529 DVDD.n3158 0.0218
R7071 DVDD.n3157 DVDD.n3143 0.0218
R7072 DVDD.n4880 DVDD.n3143 0.0218
R7073 DVDD.n1733 DVDD.n1731 0.02165
R7074 DVDD.n1489 DVDD.n1487 0.02165
R7075 DVDD.n1734 DVDD.n1606 0.02165
R7076 DVDD.n1490 DVDD.n370 0.02165
R7077 DVDD.n1742 DVDD.n1741 0.02165
R7078 DVDD.n1483 DVDD.n909 0.02165
R7079 DVDD.n1739 DVDD.n894 0.02165
R7080 DVDD.n1484 DVDD.n1400 0.02165
R7081 DVDD.n5666 DVDD.n5665 0.021425
R7082 DVDD.n4527 DVDD.n4526 0.021425
R7083 DVDD.n5318 DVDD.n5317 0.021425
R7084 DVDD.n5297 DVDD.n4919 0.021425
R7085 DVDD.n4535 DVDD.n4495 0.0213209
R7086 DVDD.n4506 DVDD.n4495 0.0213209
R7087 DVDD.n4506 DVDD.n4501 0.0213209
R7088 DVDD.n4525 DVDD.n4501 0.0213209
R7089 DVDD.n4525 DVDD.n4524 0.0213209
R7090 DVDD.n4524 DVDD.n4523 0.0213209
R7091 DVDD.n4523 DVDD.n3147 0.0213209
R7092 DVDD.n4876 DVDD.n3147 0.0213209
R7093 DVDD.n4876 DVDD.n3140 0.0213209
R7094 DVDD.n4883 DVDD.n3140 0.0213209
R7095 DVDD.n5755 DVDD.n179 0.0213209
R7096 DVDD.n3132 DVDD.n179 0.0213209
R7097 DVDD.n3132 DVDD.n3129 0.0213209
R7098 DVDD.n4902 DVDD.n3129 0.0213209
R7099 DVDD.n5320 DVDD.n4902 0.0213209
R7100 DVDD.n5320 DVDD.n5319 0.0213209
R7101 DVDD.n5319 DVDD.n4904 0.0213209
R7102 DVDD.n4911 DVDD.n4904 0.0213209
R7103 DVDD.n5309 DVDD.n4911 0.0213209
R7104 DVDD.n5309 DVDD.n5308 0.0213209
R7105 DVDD.n5307 DVDD.n4915 0.0213209
R7106 DVDD.n5110 DVDD.n4915 0.0213209
R7107 DVDD.n5110 DVDD.n4921 0.0213209
R7108 DVDD.n5296 DVDD.n4921 0.0213209
R7109 DVDD.n5296 DVDD.n5295 0.0213209
R7110 DVDD.n5295 DVDD.n5294 0.0213209
R7111 DVDD.n5294 DVDD.n4924 0.0213209
R7112 DVDD.n4932 DVDD.n4924 0.0213209
R7113 DVDD.n5284 DVDD.n4932 0.0213209
R7114 DVDD.n5284 DVDD.n5283 0.0213209
R7115 DVDD.n5022 DVDD.n5021 0.0213209
R7116 DVDD.n5026 DVDD.n5025 0.0213209
R7117 DVDD.n5668 DVDD.n5667 0.0213209
R7118 DVDD.n309 DVDD.n308 0.0213209
R7119 DVDD.n5657 DVDD.n5656 0.0213209
R7120 DVDD.n1265 DVDD.n1264 0.021153
R7121 DVDD.n2541 DVDD.n2529 0.021153
R7122 DVDD.n4640 DVDD.n3399 0.0209851
R7123 DVDD.n730 DVDD 0.0209756
R7124 DVDD.n232 DVDD 0.0202739
R7125 DVDD DVDD.n3174 0.0202739
R7126 DVDD.n1212 DVDD.n1119 0.0201455
R7127 DVDD.n2526 DVDD.n1038 0.0201455
R7128 DVDD.n2559 DVDD.n1034 0.0198097
R7129 DVDD.n5024 DVDD.n5015 0.019625
R7130 DVDD.n4522 DVDD.n4521 0.019625
R7131 DVDD.n4901 DVDD.n4900 0.019625
R7132 DVDD.n5293 DVDD.n5292 0.019625
R7133 DVDD.n5808 DVDD.n170 0.0194
R7134 DVDD.n5758 DVDD.n174 0.0194
R7135 DVDD.n4740 DVDD.n3256 0.0194
R7136 DVDD.n4848 DVDD.n4847 0.0194
R7137 DVDD.n1471 DVDD.n1389 0.0188022
R7138 DVDD.n1252 DVDD.n1214 0.0188022
R7139 DVDD.n1210 DVDD.n1042 0.0188022
R7140 DVDD.n2941 DVDD.n978 0.0184664
R7141 DVDD.n5507 DVDD.n324 0.0181306
R7142 DVDD.n1713 DVDD.n1711 0.01805
R7143 DVDD.n1503 DVDD.n1501 0.01805
R7144 DVDD.n3862 DVDD.n3584 0.01805
R7145 DVDD.n2047 DVDD.n2046 0.01805
R7146 DVDD.n1504 DVDD.n372 0.01805
R7147 DVDD.n3926 DVDD.n3656 0.01805
R7148 DVDD.n2039 DVDD.n1715 0.01805
R7149 DVDD.n1497 DVDD.n911 0.01805
R7150 DVDD.n2040 DVDD.n896 0.01805
R7151 DVDD.n1498 DVDD.n1402 0.01805
R7152 DVDD.n1536 DVDD.n1473 0.017459
R7153 DVDD.n1234 DVDD.n1220 0.017459
R7154 DVDD.n5669 DVDD.n298 0.017375
R7155 DVDD.n5035 DVDD.n302 0.017375
R7156 DVDD.n4500 DVDD.n3169 0.017375
R7157 DVDD.n5321 DVDD.n733 0.017375
R7158 DVDD.n5745 DVDD.n200 0.017375
R7159 DVDD.n5298 DVDD.n233 0.017375
R7160 DVDD.n5299 DVDD.n230 0.017375
R7161 DVDD.n4861 DVDD.n3171 0.017375
R7162 DVDD.n3868 DVDD.n3583 0.01715
R7163 DVDD.n3920 DVDD.n3659 0.01715
R7164 DVDD.n1024 DVDD.n444 0.0171231
R7165 DVDD.n2759 DVDD.n2603 0.0167873
R7166 DVDD.n5661 DVDD.n5660 0.0166964
R7167 DVDD.n5013 DVDD.n5012 0.0166964
R7168 DVDD.n5313 DVDD.n5312 0.0166964
R7169 DVDD.n5751 DVDD.n180 0.0166964
R7170 DVDD.n5288 DVDD.n5287 0.0166964
R7171 DVDD.n5304 DVDD.n4916 0.0166964
R7172 DVDD.n4881 DVDD.n3142 0.0166964
R7173 DVDD.n4532 DVDD.n4496 0.0166964
R7174 DVDD.n599 DVDD.n577 0.01625
R7175 DVDD.n2923 DVDD.n2922 0.01625
R7176 DVDD.n1596 DVDD.n573 0.01625
R7177 DVDD.n2614 DVDD.n2584 0.01625
R7178 DVDD.n1720 DVDD.n562 0.01625
R7179 DVDD.n2586 DVDD.n485 0.01625
R7180 DVDD.n886 DVDD.n558 0.01625
R7181 DVDD.n2916 DVDD.n2915 0.01625
R7182 DVDD.n1522 DVDD.n1475 0.0161157
R7183 DVDD.n1019 DVDD.n1014 0.0157799
R7184 DVDD.n5669 DVDD.n297 0.015575
R7185 DVDD.n5035 DVDD.n5034 0.015575
R7186 DVDD.n4520 DVDD.n3169 0.015575
R7187 DVDD.n5321 DVDD.n185 0.015575
R7188 DVDD.n5746 DVDD.n5745 0.015575
R7189 DVDD.n4925 DVDD.n233 0.015575
R7190 DVDD.n4927 DVDD.n230 0.015575
R7191 DVDD.n4861 DVDD.n3170 0.015575
R7192 DVDD.n566 DVDD.n331 0.015444
R7193 DVDD.n2596 DVDD.n2585 0.015444
R7194 DVDD.n2934 DVDD.n997 0.01535
R7195 DVDD.n5634 DVDD.n428 0.01535
R7196 DVDD.n1008 DVDD.n475 0.01535
R7197 DVDD.n5621 DVDD.n463 0.01535
R7198 DVDD.n1714 DVDD.n315 0.0147724
R7199 DVDD.n1508 DVDD.n1477 0.0147724
R7200 DVDD.n3355 DVDD.n3255 0.0147105
R7201 DVDD.n5760 DVDD.n5759 0.0147105
R7202 DVDD.n4683 DVDD.n3377 0.0147105
R7203 DVDD.n3423 DVDD.n3421 0.0147105
R7204 DVDD.n1517 DVDD.n1515 0.01445
R7205 DVDD.n1518 DVDD.n374 0.01445
R7206 DVDD.n1511 DVDD.n913 0.01445
R7207 DVDD.n1512 DVDD.n1404 0.01445
R7208 DVDD.n2685 DVDD.n2684 0.0142903
R7209 DVDD.n4079 DVDD.n4078 0.0142903
R7210 DVDD.n6019 DVDD.n6018 0.0142808
R7211 DVDD.n3895 DVDD.n3685 0.0141679
R7212 DVDD.n3898 DVDD.n3847 0.0141679
R7213 DVDD.n3838 DVDD.n3836 0.0141679
R7214 DVDD.n3835 DVDD.n3832 0.0141679
R7215 DVDD.n3843 DVDD.n3833 0.0141679
R7216 DVDD.n3836 DVDD.n3835 0.0141679
R7217 DVDD.n3843 DVDD.n3832 0.0141679
R7218 DVDD.n3837 DVDD.n3833 0.0141679
R7219 DVDD.n3897 DVDD.n3685 0.0141679
R7220 DVDD.n3898 DVDD.n3848 0.0141679
R7221 DVDD.n5514 DVDD.n559 0.0141679
R7222 DVDD.n5509 DVDD.n563 0.0141679
R7223 DVDD.n569 DVDD.n567 0.0141679
R7224 DVDD.n570 DVDD.n569 0.0141679
R7225 DVDD.n5504 DVDD.n568 0.0141679
R7226 DVDD.n572 DVDD.n568 0.0141679
R7227 DVDD.n5503 DVDD.n574 0.0141679
R7228 DVDD.n5500 DVDD.n578 0.0141679
R7229 DVDD.n5511 DVDD.n563 0.0141679
R7230 DVDD.n5508 DVDD.n567 0.0141679
R7231 DVDD.n5504 DVDD.n571 0.0141679
R7232 DVDD.n5501 DVDD.n574 0.0141679
R7233 DVDD.n578 DVDD.n544 0.0141679
R7234 DVDD.n571 DVDD.n570 0.0141679
R7235 DVDD.n5506 DVDD.n572 0.0141679
R7236 DVDD.n554 DVDD.n547 0.0141679
R7237 DVDD.n551 DVDD.n548 0.0141679
R7238 DVDD.n5524 DVDD.n554 0.0141679
R7239 DVDD.n5526 DVDD.n548 0.0141679
R7240 DVDD.n5512 DVDD.n559 0.0141679
R7241 DVDD.n3830 DVDD.n3686 0.0137065
R7242 DVDD.n3830 DVDD.n3829 0.0137065
R7243 DVDD.n4150 DVDD.n3538 0.0137065
R7244 DVDD.n4153 DVDD.n3538 0.0137065
R7245 DVDD.n1737 DVDD.n317 0.0134291
R7246 DVDD.n1494 DVDD.n1479 0.0134291
R7247 DVDD.n5024 DVDD.n297 0.013325
R7248 DVDD.n4522 DVDD.n4520 0.013325
R7249 DVDD.n4901 DVDD.n185 0.013325
R7250 DVDD.n5293 DVDD.n4925 0.013325
R7251 DVDD.n1785 DVDD.n1781 0.0127609
R7252 DVDD.n1784 DVDD.n1777 0.0127609
R7253 DVDD.n1854 DVDD.n1776 0.0127609
R7254 DVDD.n2977 DVDD.n787 0.0127609
R7255 DVDD.n5505 DVDD.n323 0.0127575
R7256 DVDD.n1856 DVDD.n1774 0.0127528
R7257 DVDD.n2604 DVDD.n2580 0.01265
R7258 DVDD.n3876 DVDD.n3581 0.01265
R7259 DVDD.n2756 DVDD.n2755 0.01265
R7260 DVDD.n3950 DVDD.n3655 0.01265
R7261 DVDD.n2761 DVDD.n483 0.01265
R7262 DVDD.n2764 DVDD.n2763 0.01265
R7263 DVDD.n5515 DVDD.n546 0.01221
R7264 DVDD.n5529 DVDD.n5528 0.01221
R7265 DVDD.n5652 DVDD.n357 0.0120858
R7266 DVDD.n5032 DVDD.n304 0.01175
R7267 DVDD.n4907 DVDD.n184 0.01175
R7268 DVDD.n5729 DVDD.n223 0.01175
R7269 DVDD.n4863 DVDD.n3158 0.01175
R7270 DVDD.n995 DVDD.n443 0.01175
R7271 DVDD.n4036 DVDD.n3587 0.01175
R7272 DVDD.n5631 DVDD.n5630 0.01175
R7273 DVDD.n3934 DVDD.n3651 0.01175
R7274 DVDD.n2948 DVDD.n445 0.01175
R7275 DVDD.n5624 DVDD.n5623 0.01175
R7276 DVDD.n5666 DVDD.n298 0.011525
R7277 DVDD.n4526 DVDD.n4500 0.011525
R7278 DVDD.n5318 DVDD.n733 0.011525
R7279 DVDD.n5298 DVDD.n5297 0.011525
R7280 DVDD.n3616 DVDD.n3606 0.0113864
R7281 DVDD.n3621 DVDD.n3615 0.0113864
R7282 DVDD.n3623 DVDD.n3607 0.0113864
R7283 DVDD.n3620 DVDD.n3614 0.0113864
R7284 DVDD.n3624 DVDD.n3608 0.0113864
R7285 DVDD.n3619 DVDD.n3613 0.0113864
R7286 DVDD.n3625 DVDD.n3609 0.0113864
R7287 DVDD.n3618 DVDD.n3612 0.0113864
R7288 DVDD.n3626 DVDD.n3610 0.0113864
R7289 DVDD.n3617 DVDD.n3611 0.0113864
R7290 DVDD.n4490 DVDD.n4489 0.0113864
R7291 DVDD.n3446 DVDD.n3436 0.0113864
R7292 DVDD.n4486 DVDD.n3443 0.0113864
R7293 DVDD.n3447 DVDD.n3437 0.0113864
R7294 DVDD.n3442 DVDD.n3399 0.0113864
R7295 DVDD.n3444 DVDD.n3439 0.0113864
R7296 DVDD.n4487 DVDD.n3434 0.0113864
R7297 DVDD.n4492 DVDD.n3440 0.0113864
R7298 DVDD.n4494 DVDD.n3431 0.0113864
R7299 DVDD.n5247 DVDD.n4935 0.0113864
R7300 DVDD.n5246 DVDD.n4949 0.0113864
R7301 DVDD.n5268 DVDD.n5249 0.0113864
R7302 DVDD.n5248 DVDD.n4948 0.0113864
R7303 DVDD.n5269 DVDD.n5251 0.0113864
R7304 DVDD.n5250 DVDD.n4947 0.0113864
R7305 DVDD.n5270 DVDD.n5253 0.0113864
R7306 DVDD.n5252 DVDD.n4946 0.0113864
R7307 DVDD.n5271 DVDD.n5255 0.0113864
R7308 DVDD.n5254 DVDD.n4945 0.0113864
R7309 DVDD.n5272 DVDD.n5257 0.0113864
R7310 DVDD.n5256 DVDD.n4944 0.0113864
R7311 DVDD.n5273 DVDD.n5259 0.0113864
R7312 DVDD.n5258 DVDD.n4943 0.0113864
R7313 DVDD.n5274 DVDD.n5261 0.0113864
R7314 DVDD.n5260 DVDD.n4942 0.0113864
R7315 DVDD.n5275 DVDD.n5263 0.0113864
R7316 DVDD.n5262 DVDD.n4941 0.0113864
R7317 DVDD.n5276 DVDD.n5265 0.0113864
R7318 DVDD.n5264 DVDD.n4940 0.0113864
R7319 DVDD.n5277 DVDD.n5267 0.0113864
R7320 DVDD.n5266 DVDD.n4939 0.0113864
R7321 DVDD.n5280 DVDD.n5279 0.0113864
R7322 DVDD.n5021 DVDD.n5016 0.0113864
R7323 DVDD.n5026 DVDD.n5023 0.0113864
R7324 DVDD.n5668 DVDD.n299 0.0113864
R7325 DVDD.n308 DVDD.n300 0.0113864
R7326 DVDD.n5657 DVDD.n310 0.0113864
R7327 DVDD.n328 DVDD.n311 0.0113864
R7328 DVDD.n327 DVDD.n325 0.0113864
R7329 DVDD.n347 DVDD.n330 0.0113864
R7330 DVDD.n329 DVDD.n324 0.0113864
R7331 DVDD.n332 DVDD.n322 0.0113864
R7332 DVDD.n348 DVDD.n335 0.0113864
R7333 DVDD.n334 DVDD.n321 0.0113864
R7334 DVDD.n349 DVDD.n337 0.0113864
R7335 DVDD.n336 DVDD.n320 0.0113864
R7336 DVDD.n350 DVDD.n339 0.0113864
R7337 DVDD.n338 DVDD.n319 0.0113864
R7338 DVDD.n351 DVDD.n341 0.0113864
R7339 DVDD.n340 DVDD.n318 0.0113864
R7340 DVDD.n352 DVDD.n342 0.0113864
R7341 DVDD.n353 DVDD.n344 0.0113864
R7342 DVDD.n343 DVDD.n316 0.0113864
R7343 DVDD.n354 DVDD.n345 0.0113864
R7344 DVDD.n5653 DVDD.n356 0.0113864
R7345 DVDD.n1553 DVDD.n1482 0.0113864
R7346 DVDD.n1547 DVDD.n1480 0.0113864
R7347 DVDD.n1554 DVDD.n1495 0.0113864
R7348 DVDD.n1555 DVDD.n1496 0.0113864
R7349 DVDD.n1546 DVDD.n1478 0.0113864
R7350 DVDD.n1556 DVDD.n1509 0.0113864
R7351 DVDD.n1557 DVDD.n1510 0.0113864
R7352 DVDD.n1545 DVDD.n1476 0.0113864
R7353 DVDD.n1558 DVDD.n1523 0.0113864
R7354 DVDD.n1559 DVDD.n1524 0.0113864
R7355 DVDD.n1544 DVDD.n1474 0.0113864
R7356 DVDD.n1560 DVDD.n1537 0.0113864
R7357 DVDD.n1561 DVDD.n1538 0.0113864
R7358 DVDD.n1543 DVDD.n1472 0.0113864
R7359 DVDD.n1562 DVDD.n1539 0.0113864
R7360 DVDD.n1563 DVDD.n1540 0.0113864
R7361 DVDD.n1542 DVDD.n1470 0.0113864
R7362 DVDD.n2153 DVDD.n1541 0.0113864
R7363 DVDD.n1235 DVDD.n1196 0.0113864
R7364 DVDD.n1236 DVDD.n1197 0.0113864
R7365 DVDD.n1272 DVDD.n1219 0.0113864
R7366 DVDD.n1237 DVDD.n1198 0.0113864
R7367 DVDD.n1271 DVDD.n1218 0.0113864
R7368 DVDD.n1238 DVDD.n1199 0.0113864
R7369 DVDD.n1270 DVDD.n1217 0.0113864
R7370 DVDD.n1239 DVDD.n1200 0.0113864
R7371 DVDD.n1269 DVDD.n1216 0.0113864
R7372 DVDD.n1240 DVDD.n1201 0.0113864
R7373 DVDD.n1268 DVDD.n1215 0.0113864
R7374 DVDD.n1253 DVDD.n1202 0.0113864
R7375 DVDD.n1254 DVDD.n1203 0.0113864
R7376 DVDD.n1267 DVDD.n1213 0.0113864
R7377 DVDD.n1255 DVDD.n1204 0.0113864
R7378 DVDD.n1256 DVDD.n1205 0.0113864
R7379 DVDD.n1266 DVDD.n1265 0.0113864
R7380 DVDD.n1211 DVDD.n1194 0.0113864
R7381 DVDD.n2372 DVDD.n1206 0.0113864
R7382 DVDD.n1041 DVDD.n1040 0.0113864
R7383 DVDD.n2511 DVDD.n1039 0.0113864
R7384 DVDD.n2527 DVDD.n2512 0.0113864
R7385 DVDD.n1037 DVDD.n1036 0.0113864
R7386 DVDD.n2529 DVDD.n1035 0.0113864
R7387 DVDD.n2546 DVDD.n2545 0.0113864
R7388 DVDD.n2547 DVDD.n2544 0.0113864
R7389 DVDD.n2543 DVDD.n1034 0.0113864
R7390 DVDD.n2560 DVDD.n1033 0.0113864
R7391 DVDD.n1032 DVDD.n1031 0.0113864
R7392 DVDD.n1030 DVDD.n978 0.0113864
R7393 DVDD.n1029 DVDD.n1026 0.0113864
R7394 DVDD.n1028 DVDD.n1027 0.0113864
R7395 DVDD.n1025 DVDD.n1024 0.0113864
R7396 DVDD.n2562 DVDD.n1023 0.0113864
R7397 DVDD.n1022 DVDD.n1021 0.0113864
R7398 DVDD.n1020 DVDD.n1019 0.0113864
R7399 DVDD.n517 DVDD.n515 0.0113864
R7400 DVDD.n2598 DVDD.n2597 0.0113864
R7401 DVDD.n2603 DVDD.n514 0.0113864
R7402 DVDD.n519 DVDD.n513 0.0113864
R7403 DVDD.n2600 DVDD.n2599 0.0113864
R7404 DVDD.n2596 DVDD.n512 0.0113864
R7405 DVDD.n521 DVDD.n511 0.0113864
R7406 DVDD.n5567 DVDD.n523 0.0113864
R7407 DVDD.n3617 DVDD.n3610 0.0113864
R7408 DVDD.n3626 DVDD.n3612 0.0113864
R7409 DVDD.n3618 DVDD.n3609 0.0113864
R7410 DVDD.n3625 DVDD.n3613 0.0113864
R7411 DVDD.n3619 DVDD.n3608 0.0113864
R7412 DVDD.n3624 DVDD.n3614 0.0113864
R7413 DVDD.n3620 DVDD.n3607 0.0113864
R7414 DVDD.n3623 DVDD.n3615 0.0113864
R7415 DVDD.n3621 DVDD.n3606 0.0113864
R7416 DVDD.n4000 DVDD.n3616 0.0113864
R7417 DVDD.n5282 DVDD.n4935 0.0113864
R7418 DVDD.n5247 DVDD.n5246 0.0113864
R7419 DVDD.n5268 DVDD.n4949 0.0113864
R7420 DVDD.n5249 DVDD.n5248 0.0113864
R7421 DVDD.n5269 DVDD.n4948 0.0113864
R7422 DVDD.n5251 DVDD.n5250 0.0113864
R7423 DVDD.n5270 DVDD.n4947 0.0113864
R7424 DVDD.n5253 DVDD.n5252 0.0113864
R7425 DVDD.n5271 DVDD.n4946 0.0113864
R7426 DVDD.n5255 DVDD.n5254 0.0113864
R7427 DVDD.n5272 DVDD.n4945 0.0113864
R7428 DVDD.n5257 DVDD.n5256 0.0113864
R7429 DVDD.n5273 DVDD.n4944 0.0113864
R7430 DVDD.n5259 DVDD.n5258 0.0113864
R7431 DVDD.n5274 DVDD.n4943 0.0113864
R7432 DVDD.n5261 DVDD.n5260 0.0113864
R7433 DVDD.n5275 DVDD.n4942 0.0113864
R7434 DVDD.n5263 DVDD.n5262 0.0113864
R7435 DVDD.n5276 DVDD.n4941 0.0113864
R7436 DVDD.n5265 DVDD.n5264 0.0113864
R7437 DVDD.n5277 DVDD.n4940 0.0113864
R7438 DVDD.n5267 DVDD.n5266 0.0113864
R7439 DVDD.n5279 DVDD.n4939 0.0113864
R7440 DVDD.n5017 DVDD.n5016 0.0113864
R7441 DVDD.n5023 DVDD.n5022 0.0113864
R7442 DVDD.n5025 DVDD.n299 0.0113864
R7443 DVDD.n5667 DVDD.n300 0.0113864
R7444 DVDD.n310 DVDD.n309 0.0113864
R7445 DVDD.n5655 DVDD.n311 0.0113864
R7446 DVDD.n328 DVDD.n327 0.0113864
R7447 DVDD.n347 DVDD.n325 0.0113864
R7448 DVDD.n330 DVDD.n329 0.0113864
R7449 DVDD.n333 DVDD.n332 0.0113864
R7450 DVDD.n348 DVDD.n322 0.0113864
R7451 DVDD.n335 DVDD.n334 0.0113864
R7452 DVDD.n349 DVDD.n321 0.0113864
R7453 DVDD.n337 DVDD.n336 0.0113864
R7454 DVDD.n350 DVDD.n320 0.0113864
R7455 DVDD.n339 DVDD.n338 0.0113864
R7456 DVDD.n351 DVDD.n319 0.0113864
R7457 DVDD.n341 DVDD.n340 0.0113864
R7458 DVDD.n352 DVDD.n318 0.0113864
R7459 DVDD.n353 DVDD.n317 0.0113864
R7460 DVDD.n344 DVDD.n343 0.0113864
R7461 DVDD.n354 DVDD.n316 0.0113864
R7462 DVDD.n356 DVDD.n315 0.0113864
R7463 DVDD.n1553 DVDD.n357 0.0113864
R7464 DVDD.n1547 DVDD.n1482 0.0113864
R7465 DVDD.n1554 DVDD.n1480 0.0113864
R7466 DVDD.n1555 DVDD.n1479 0.0113864
R7467 DVDD.n1546 DVDD.n1496 0.0113864
R7468 DVDD.n1556 DVDD.n1478 0.0113864
R7469 DVDD.n1557 DVDD.n1477 0.0113864
R7470 DVDD.n1545 DVDD.n1510 0.0113864
R7471 DVDD.n1558 DVDD.n1476 0.0113864
R7472 DVDD.n1559 DVDD.n1475 0.0113864
R7473 DVDD.n1544 DVDD.n1524 0.0113864
R7474 DVDD.n1560 DVDD.n1474 0.0113864
R7475 DVDD.n1561 DVDD.n1473 0.0113864
R7476 DVDD.n1543 DVDD.n1538 0.0113864
R7477 DVDD.n1562 DVDD.n1472 0.0113864
R7478 DVDD.n1563 DVDD.n1471 0.0113864
R7479 DVDD.n1542 DVDD.n1540 0.0113864
R7480 DVDD.n1541 DVDD.n1470 0.0113864
R7481 DVDD.n1221 DVDD.n1196 0.0113864
R7482 DVDD.n1220 DVDD.n1197 0.0113864
R7483 DVDD.n1272 DVDD.n1236 0.0113864
R7484 DVDD.n1219 DVDD.n1198 0.0113864
R7485 DVDD.n1271 DVDD.n1237 0.0113864
R7486 DVDD.n1218 DVDD.n1199 0.0113864
R7487 DVDD.n1270 DVDD.n1238 0.0113864
R7488 DVDD.n1217 DVDD.n1200 0.0113864
R7489 DVDD.n1269 DVDD.n1239 0.0113864
R7490 DVDD.n1216 DVDD.n1201 0.0113864
R7491 DVDD.n1268 DVDD.n1240 0.0113864
R7492 DVDD.n1215 DVDD.n1202 0.0113864
R7493 DVDD.n1214 DVDD.n1203 0.0113864
R7494 DVDD.n1267 DVDD.n1254 0.0113864
R7495 DVDD.n1213 DVDD.n1204 0.0113864
R7496 DVDD.n1212 DVDD.n1205 0.0113864
R7497 DVDD.n1266 DVDD.n1256 0.0113864
R7498 DVDD.n2370 DVDD.n1194 0.0113864
R7499 DVDD.n1211 DVDD.n1206 0.0113864
R7500 DVDD.n1042 DVDD.n1041 0.0113864
R7501 DVDD.n1040 DVDD.n1039 0.0113864
R7502 DVDD.n2512 DVDD.n2511 0.0113864
R7503 DVDD.n1038 DVDD.n1037 0.0113864
R7504 DVDD.n1036 DVDD.n1035 0.0113864
R7505 DVDD.n2545 DVDD.n2542 0.0113864
R7506 DVDD.n2547 DVDD.n2546 0.0113864
R7507 DVDD.n2544 DVDD.n2543 0.0113864
R7508 DVDD.n2561 DVDD.n2560 0.0113864
R7509 DVDD.n1033 DVDD.n1032 0.0113864
R7510 DVDD.n1031 DVDD.n1030 0.0113864
R7511 DVDD.n1026 DVDD.n979 0.0113864
R7512 DVDD.n1029 DVDD.n1028 0.0113864
R7513 DVDD.n1027 DVDD.n1025 0.0113864
R7514 DVDD.n2563 DVDD.n2562 0.0113864
R7515 DVDD.n1023 DVDD.n1022 0.0113864
R7516 DVDD.n1021 DVDD.n1020 0.0113864
R7517 DVDD.n518 DVDD.n517 0.0113864
R7518 DVDD.n2598 DVDD.n515 0.0113864
R7519 DVDD.n2597 DVDD.n514 0.0113864
R7520 DVDD.n520 DVDD.n519 0.0113864
R7521 DVDD.n2600 DVDD.n513 0.0113864
R7522 DVDD.n2599 DVDD.n512 0.0113864
R7523 DVDD.n522 DVDD.n521 0.0113864
R7524 DVDD.n523 DVDD.n511 0.0113864
R7525 DVDD.n3447 DVDD.n3442 0.0113864
R7526 DVDD.n4486 DVDD.n3437 0.0113864
R7527 DVDD.n3446 DVDD.n3443 0.0113864
R7528 DVDD.n4489 DVDD.n3436 0.0113864
R7529 DVDD.n4490 DVDD.n3435 0.0113864
R7530 DVDD.n4487 DVDD.n3439 0.0113864
R7531 DVDD.n3440 DVDD.n3434 0.0113864
R7532 DVDD.n4492 DVDD.n3431 0.0113864
R7533 DVDD.n3444 DVDD.n3401 0.0113864
R7534 DVDD.n1531 DVDD.n1529 0.01085
R7535 DVDD.n1229 DVDD.n1227 0.01085
R7536 DVDD.n3860 DVDD.n3577 0.01085
R7537 DVDD.n1532 DVDD.n376 0.01085
R7538 DVDD.n1230 DVDD.n389 0.01085
R7539 DVDD.n3928 DVDD.n3652 0.01085
R7540 DVDD.n1525 DVDD.n915 0.01085
R7541 DVDD.n1223 DVDD.n928 0.01085
R7542 DVDD.n1526 DVDD.n1406 0.01085
R7543 DVDD.n1224 DVDD.n1129 0.01085
R7544 DVDD.n5033 DVDD.n5032 0.01055
R7545 DVDD.n5747 DVDD.n184 0.01055
R7546 DVDD.n5729 DVDD.n222 0.01055
R7547 DVDD.n4863 DVDD.n3157 0.01055
R7548 DVDD.n4885 DVDD.n176 0.0104
R7549 DVDD.n4791 DVDD.n3253 0.0104
R7550 DVDD.n4719 DVDD.n3357 0.0104
R7551 DVDD.n4789 DVDD.n4788 0.0104
R7552 DVDD.n4887 DVDD.n4886 0.0104
R7553 DVDD.n4720 DVDD.n3359 0.0104
R7554 DVDD.n3227 DVDD.n3205 0.0104
R7555 DVDD.n3229 DVDD.n3228 0.0104
R7556 DVDD.n3935 DVDD.n3933 0.01022
R7557 DVDD.n3933 DVDD.n3930 0.01022
R7558 DVDD.n3930 DVDD.n3929 0.01022
R7559 DVDD.n3929 DVDD.n3927 0.01022
R7560 DVDD.n3927 DVDD.n3925 0.01022
R7561 DVDD.n3925 DVDD.n3923 0.01022
R7562 DVDD.n3923 DVDD.n3921 0.01022
R7563 DVDD.n3921 DVDD.n3662 0.01022
R7564 DVDD.n3953 DVDD.n3662 0.01022
R7565 DVDD.n3953 DVDD.n3952 0.01022
R7566 DVDD.n3952 DVDD.n3951 0.01022
R7567 DVDD.n3951 DVDD.n3949 0.01022
R7568 DVDD.n3949 DVDD.n3663 0.01022
R7569 DVDD.n3945 DVDD.n3663 0.01022
R7570 DVDD.n3945 DVDD.n3944 0.01022
R7571 DVDD.n3944 DVDD.n3943 0.01022
R7572 DVDD.n3943 DVDD.n3665 0.01022
R7573 DVDD.n3939 DVDD.n3665 0.01022
R7574 DVDD.n3939 DVDD.n3938 0.01022
R7575 DVDD.n3856 DVDD.n3855 0.01022
R7576 DVDD.n3859 DVDD.n3856 0.01022
R7577 DVDD.n3861 DVDD.n3859 0.01022
R7578 DVDD.n3863 DVDD.n3861 0.01022
R7579 DVDD.n3865 DVDD.n3863 0.01022
R7580 DVDD.n3867 DVDD.n3865 0.01022
R7581 DVDD.n3869 DVDD.n3867 0.01022
R7582 DVDD.n3871 DVDD.n3869 0.01022
R7583 DVDD.n3872 DVDD.n3871 0.01022
R7584 DVDD.n3875 DVDD.n3872 0.01022
R7585 DVDD.n3877 DVDD.n3875 0.01022
R7586 DVDD.n3878 DVDD.n3877 0.01022
R7587 DVDD.n3881 DVDD.n3878 0.01022
R7588 DVDD.n3882 DVDD.n3881 0.01022
R7589 DVDD.n3883 DVDD.n3882 0.01022
R7590 DVDD.n3883 DVDD.n3853 0.01022
R7591 DVDD.n3887 DVDD.n3853 0.01022
R7592 DVDD.n3888 DVDD.n3887 0.01022
R7593 DVDD.n3890 DVDD.n3888 0.01022
R7594 DVDD.n3896 DVDD.n3849 0.0100489
R7595 DVDD.n3901 DVDD.n3684 0.0100489
R7596 DVDD.n3906 DVDD.n3903 0.0100489
R7597 DVDD.n3911 DVDD.n3670 0.0100489
R7598 DVDD.n3677 DVDD.n3672 0.0100489
R7599 DVDD.n4199 DVDD.n3521 0.0100489
R7600 DVDD.n3839 DVDD.n3523 0.0100489
R7601 DVDD.n3842 DVDD.n3834 0.0100489
R7602 DVDD.n5525 DVDD.n550 0.0100489
R7603 DVDD.n552 DVDD.n549 0.0100489
R7604 DVDD.n3840 DVDD.n3839 0.0100489
R7605 DVDD.n3840 DVDD.n3834 0.0100489
R7606 DVDD.n3525 DVDD.n3521 0.0100489
R7607 DVDD.n3679 DVDD.n3672 0.0100489
R7608 DVDD.n3681 DVDD.n3670 0.0100489
R7609 DVDD.n3903 DVDD.n3902 0.0100489
R7610 DVDD.n3849 DVDD.n3684 0.0100489
R7611 DVDD.n3899 DVDD.n3896 0.0100489
R7612 DVDD.n5525 DVDD.n552 0.0100489
R7613 DVDD.n5523 DVDD.n550 0.0100489
R7614 DVDD.n4742 DVDD.n4741 0.00997368
R7615 DVDD.n3311 DVDD.n3310 0.00997368
R7616 DVDD.n3302 DVDD.n3259 0.00997368
R7617 DVDD.n5763 DVDD.n172 0.00997368
R7618 DVDD.n4278 DVDD.n3376 0.00997368
R7619 DVDD.n3395 DVDD.n3393 0.00997368
R7620 DVDD.n4639 DVDD.n3402 0.00997368
R7621 DVDD.n4598 DVDD.n4545 0.00997368
R7622 DVDD.n3870 DVDD.n3579 0.00995
R7623 DVDD.n3660 DVDD.n3649 0.00995
R7624 DVDD.n5096 DVDD.n5095 0.00992
R7625 DVDD.n3115 DVDD.n3114 0.00992
R7626 DVDD.n3064 DVDD.n207 0.00992
R7627 DVDD.n3116 DVDD.n3090 0.00992
R7628 DVDD.n5097 DVDD.n5085 0.00992
R7629 DVDD.n5738 DVDD.n208 0.00992
R7630 DVDD.n5334 DVDD.n711 0.00992
R7631 DVDD.n5335 DVDD.n718 0.00992
R7632 DVDD.n2905 DVDD.n2904 0.00962857
R7633 DVDD.n2904 DVDD.n2903 0.00962857
R7634 DVDD.n2903 DVDD.n2865 0.00962857
R7635 DVDD.n2899 DVDD.n2865 0.00962857
R7636 DVDD.n2899 DVDD.n2868 0.00962857
R7637 DVDD.n2895 DVDD.n2868 0.00962857
R7638 DVDD.n2895 DVDD.n2871 0.00962857
R7639 DVDD.n2891 DVDD.n2871 0.00962857
R7640 DVDD.n2891 DVDD.n2873 0.00962857
R7641 DVDD.n2887 DVDD.n2873 0.00962857
R7642 DVDD.n2887 DVDD.n2875 0.00962857
R7643 DVDD.n2883 DVDD.n2875 0.00962857
R7644 DVDD.n2883 DVDD.n2877 0.00962857
R7645 DVDD.n2879 DVDD.n2877 0.00962857
R7646 DVDD.n2879 DVDD.n488 0.00962857
R7647 DVDD.n5607 DVDD.n488 0.00962857
R7648 DVDD.n5607 DVDD.n489 0.00962857
R7649 DVDD.n5603 DVDD.n489 0.00962857
R7650 DVDD.n5603 DVDD.n5602 0.00962857
R7651 DVDD.n5602 DVDD.n492 0.00962857
R7652 DVDD.n5598 DVDD.n492 0.00962857
R7653 DVDD.n5598 DVDD.n494 0.00962857
R7654 DVDD.n5594 DVDD.n494 0.00962857
R7655 DVDD.n5594 DVDD.n497 0.00962857
R7656 DVDD.n5590 DVDD.n497 0.00962857
R7657 DVDD.n5590 DVDD.n499 0.00962857
R7658 DVDD.n5586 DVDD.n499 0.00962857
R7659 DVDD.n5586 DVDD.n501 0.00962857
R7660 DVDD.n5582 DVDD.n501 0.00962857
R7661 DVDD.n5582 DVDD.n503 0.00962857
R7662 DVDD.n5578 DVDD.n503 0.00962857
R7663 DVDD.n5578 DVDD.n505 0.00962857
R7664 DVDD.n5574 DVDD.n505 0.00962857
R7665 DVDD.n5574 DVDD.n507 0.00962857
R7666 DVDD.n5570 DVDD.n507 0.00962857
R7667 DVDD.n5570 DVDD.n509 0.00962857
R7668 DVDD.n2631 DVDD.n509 0.00962857
R7669 DVDD.n2631 DVDD.n2629 0.00962857
R7670 DVDD.n2635 DVDD.n2629 0.00962857
R7671 DVDD.n2635 DVDD.n2627 0.00962857
R7672 DVDD.n2639 DVDD.n2627 0.00962857
R7673 DVDD.n2639 DVDD.n2625 0.00962857
R7674 DVDD.n2643 DVDD.n2625 0.00962857
R7675 DVDD.n2643 DVDD.n2623 0.00962857
R7676 DVDD.n2647 DVDD.n2623 0.00962857
R7677 DVDD.n2647 DVDD.n2621 0.00962857
R7678 DVDD.n2651 DVDD.n2621 0.00962857
R7679 DVDD.n2651 DVDD.n2619 0.00962857
R7680 DVDD.n2655 DVDD.n2619 0.00962857
R7681 DVDD.n2655 DVDD.n2616 0.00962857
R7682 DVDD.n2746 DVDD.n2616 0.00962857
R7683 DVDD.n2746 DVDD.n2617 0.00962857
R7684 DVDD.n2742 DVDD.n2617 0.00962857
R7685 DVDD.n2742 DVDD.n2741 0.00962857
R7686 DVDD.n2741 DVDD.n2659 0.00962857
R7687 DVDD.n2737 DVDD.n2659 0.00962857
R7688 DVDD.n2737 DVDD.n2661 0.00962857
R7689 DVDD.n2733 DVDD.n2661 0.00962857
R7690 DVDD.n2733 DVDD.n2664 0.00962857
R7691 DVDD.n2729 DVDD.n2664 0.00962857
R7692 DVDD.n2729 DVDD.n2666 0.00962857
R7693 DVDD.n2725 DVDD.n2666 0.00962857
R7694 DVDD.n2725 DVDD.n2668 0.00962857
R7695 DVDD.n2721 DVDD.n2668 0.00962857
R7696 DVDD.n2721 DVDD.n2670 0.00962857
R7697 DVDD.n2717 DVDD.n2670 0.00962857
R7698 DVDD.n2717 DVDD.n2714 0.00962857
R7699 DVDD.n2714 DVDD.n2713 0.00962857
R7700 DVDD.n2713 DVDD.n2672 0.00962857
R7701 DVDD.n2709 DVDD.n2672 0.00962857
R7702 DVDD.n2709 DVDD.n2708 0.00962857
R7703 DVDD.n2708 DVDD.n2674 0.00962857
R7704 DVDD.n2704 DVDD.n2674 0.00962857
R7705 DVDD.n2704 DVDD.n2676 0.00962857
R7706 DVDD.n2700 DVDD.n2676 0.00962857
R7707 DVDD.n2700 DVDD.n2679 0.00962857
R7708 DVDD.n2696 DVDD.n2679 0.00962857
R7709 DVDD.n2696 DVDD.n2681 0.00962857
R7710 DVDD.n2692 DVDD.n2681 0.00962857
R7711 DVDD.n2692 DVDD.n2683 0.00962857
R7712 DVDD.n2688 DVDD.n2683 0.00962857
R7713 DVDD.n2902 DVDD.n2591 0.00962857
R7714 DVDD.n2902 DVDD.n2901 0.00962857
R7715 DVDD.n2901 DVDD.n2900 0.00962857
R7716 DVDD.n2900 DVDD.n2867 0.00962857
R7717 DVDD.n2894 DVDD.n2867 0.00962857
R7718 DVDD.n2894 DVDD.n2893 0.00962857
R7719 DVDD.n2893 DVDD.n2892 0.00962857
R7720 DVDD.n2892 DVDD.n2872 0.00962857
R7721 DVDD.n2886 DVDD.n2872 0.00962857
R7722 DVDD.n2886 DVDD.n2885 0.00962857
R7723 DVDD.n2885 DVDD.n2884 0.00962857
R7724 DVDD.n2884 DVDD.n2876 0.00962857
R7725 DVDD.n2878 DVDD.n2876 0.00962857
R7726 DVDD.n2878 DVDD.n487 0.00962857
R7727 DVDD.n5608 DVDD.n487 0.00962857
R7728 DVDD.n5601 DVDD.n481 0.00962857
R7729 DVDD.n5601 DVDD.n5600 0.00962857
R7730 DVDD.n5600 DVDD.n5599 0.00962857
R7731 DVDD.n5599 DVDD.n493 0.00962857
R7732 DVDD.n5593 DVDD.n493 0.00962857
R7733 DVDD.n5593 DVDD.n5592 0.00962857
R7734 DVDD.n5592 DVDD.n5591 0.00962857
R7735 DVDD.n5591 DVDD.n498 0.00962857
R7736 DVDD.n5585 DVDD.n498 0.00962857
R7737 DVDD.n5585 DVDD.n5584 0.00962857
R7738 DVDD.n5584 DVDD.n5583 0.00962857
R7739 DVDD.n5583 DVDD.n502 0.00962857
R7740 DVDD.n5577 DVDD.n502 0.00962857
R7741 DVDD.n5577 DVDD.n5576 0.00962857
R7742 DVDD.n5576 DVDD.n5575 0.00962857
R7743 DVDD.n2630 DVDD.n516 0.00962857
R7744 DVDD.n2630 DVDD.n2628 0.00962857
R7745 DVDD.n2636 DVDD.n2628 0.00962857
R7746 DVDD.n2637 DVDD.n2636 0.00962857
R7747 DVDD.n2638 DVDD.n2637 0.00962857
R7748 DVDD.n2638 DVDD.n2624 0.00962857
R7749 DVDD.n2644 DVDD.n2624 0.00962857
R7750 DVDD.n2645 DVDD.n2644 0.00962857
R7751 DVDD.n2646 DVDD.n2645 0.00962857
R7752 DVDD.n2646 DVDD.n2620 0.00962857
R7753 DVDD.n2652 DVDD.n2620 0.00962857
R7754 DVDD.n2653 DVDD.n2652 0.00962857
R7755 DVDD.n2654 DVDD.n2653 0.00962857
R7756 DVDD.n2654 DVDD.n2615 0.00962857
R7757 DVDD.n2747 DVDD.n2615 0.00962857
R7758 DVDD.n2740 DVDD.n2609 0.00962857
R7759 DVDD.n2740 DVDD.n2739 0.00962857
R7760 DVDD.n2739 DVDD.n2738 0.00962857
R7761 DVDD.n2738 DVDD.n2660 0.00962857
R7762 DVDD.n2732 DVDD.n2660 0.00962857
R7763 DVDD.n2732 DVDD.n2731 0.00962857
R7764 DVDD.n2731 DVDD.n2730 0.00962857
R7765 DVDD.n2730 DVDD.n2665 0.00962857
R7766 DVDD.n2724 DVDD.n2665 0.00962857
R7767 DVDD.n2724 DVDD.n2723 0.00962857
R7768 DVDD.n2723 DVDD.n2722 0.00962857
R7769 DVDD.n2722 DVDD.n2669 0.00962857
R7770 DVDD.n2716 DVDD.n2669 0.00962857
R7771 DVDD.n2716 DVDD.n2715 0.00962857
R7772 DVDD.n2715 DVDD.n2583 0.00962857
R7773 DVDD.n2707 DVDD.n2578 0.00962857
R7774 DVDD.n2707 DVDD.n2706 0.00962857
R7775 DVDD.n2706 DVDD.n2705 0.00962857
R7776 DVDD.n2705 DVDD.n2675 0.00962857
R7777 DVDD.n2699 DVDD.n2675 0.00962857
R7778 DVDD.n2699 DVDD.n2698 0.00962857
R7779 DVDD.n2698 DVDD.n2697 0.00962857
R7780 DVDD.n2697 DVDD.n2680 0.00962857
R7781 DVDD.n2691 DVDD.n2680 0.00962857
R7782 DVDD.n2691 DVDD.n2690 0.00962857
R7783 DVDD.n2690 DVDD.n2689 0.00962857
R7784 DVDD.n3743 DVDD.n3702 0.00962857
R7785 DVDD.n3743 DVDD.n3703 0.00962857
R7786 DVDD.n3739 DVDD.n3703 0.00962857
R7787 DVDD.n3739 DVDD.n3706 0.00962857
R7788 DVDD.n3735 DVDD.n3706 0.00962857
R7789 DVDD.n3735 DVDD.n3708 0.00962857
R7790 DVDD.n3731 DVDD.n3708 0.00962857
R7791 DVDD.n3731 DVDD.n3710 0.00962857
R7792 DVDD.n3727 DVDD.n3710 0.00962857
R7793 DVDD.n3727 DVDD.n3712 0.00962857
R7794 DVDD.n3723 DVDD.n3712 0.00962857
R7795 DVDD.n3723 DVDD.n3714 0.00962857
R7796 DVDD.n3719 DVDD.n3714 0.00962857
R7797 DVDD.n3719 DVDD.n3716 0.00962857
R7798 DVDD.n3716 DVDD.n3647 0.00962857
R7799 DVDD.n3958 DVDD.n3647 0.00962857
R7800 DVDD.n3958 DVDD.n3645 0.00962857
R7801 DVDD.n3962 DVDD.n3645 0.00962857
R7802 DVDD.n3962 DVDD.n3643 0.00962857
R7803 DVDD.n3966 DVDD.n3643 0.00962857
R7804 DVDD.n3966 DVDD.n3641 0.00962857
R7805 DVDD.n3970 DVDD.n3641 0.00962857
R7806 DVDD.n3970 DVDD.n3639 0.00962857
R7807 DVDD.n3974 DVDD.n3639 0.00962857
R7808 DVDD.n3974 DVDD.n3637 0.00962857
R7809 DVDD.n3978 DVDD.n3637 0.00962857
R7810 DVDD.n3978 DVDD.n3635 0.00962857
R7811 DVDD.n3982 DVDD.n3635 0.00962857
R7812 DVDD.n3982 DVDD.n3633 0.00962857
R7813 DVDD.n3986 DVDD.n3633 0.00962857
R7814 DVDD.n3986 DVDD.n3631 0.00962857
R7815 DVDD.n3991 DVDD.n3631 0.00962857
R7816 DVDD.n3991 DVDD.n3628 0.00962857
R7817 DVDD.n3996 DVDD.n3628 0.00962857
R7818 DVDD.n3996 DVDD.n3629 0.00962857
R7819 DVDD.n3629 DVDD.n3604 0.00962857
R7820 DVDD.n4004 DVDD.n3604 0.00962857
R7821 DVDD.n4004 DVDD.n3602 0.00962857
R7822 DVDD.n4008 DVDD.n3602 0.00962857
R7823 DVDD.n4008 DVDD.n3600 0.00962857
R7824 DVDD.n4012 DVDD.n3600 0.00962857
R7825 DVDD.n4012 DVDD.n3598 0.00962857
R7826 DVDD.n4016 DVDD.n3598 0.00962857
R7827 DVDD.n4016 DVDD.n3596 0.00962857
R7828 DVDD.n4020 DVDD.n3596 0.00962857
R7829 DVDD.n4020 DVDD.n3594 0.00962857
R7830 DVDD.n4024 DVDD.n3594 0.00962857
R7831 DVDD.n4024 DVDD.n3592 0.00962857
R7832 DVDD.n4028 DVDD.n3592 0.00962857
R7833 DVDD.n4028 DVDD.n3589 0.00962857
R7834 DVDD.n4033 DVDD.n3589 0.00962857
R7835 DVDD.n4033 DVDD.n3590 0.00962857
R7836 DVDD.n3590 DVDD.n3574 0.00962857
R7837 DVDD.n4040 DVDD.n3574 0.00962857
R7838 DVDD.n4040 DVDD.n3572 0.00962857
R7839 DVDD.n4044 DVDD.n3572 0.00962857
R7840 DVDD.n4044 DVDD.n3570 0.00962857
R7841 DVDD.n4048 DVDD.n3570 0.00962857
R7842 DVDD.n4048 DVDD.n3568 0.00962857
R7843 DVDD.n4052 DVDD.n3568 0.00962857
R7844 DVDD.n4052 DVDD.n3566 0.00962857
R7845 DVDD.n4056 DVDD.n3566 0.00962857
R7846 DVDD.n4056 DVDD.n3564 0.00962857
R7847 DVDD.n4060 DVDD.n3564 0.00962857
R7848 DVDD.n4060 DVDD.n3562 0.00962857
R7849 DVDD.n4064 DVDD.n3562 0.00962857
R7850 DVDD.n4064 DVDD.n3559 0.00962857
R7851 DVDD.n4107 DVDD.n3559 0.00962857
R7852 DVDD.n4107 DVDD.n3560 0.00962857
R7853 DVDD.n4103 DVDD.n3560 0.00962857
R7854 DVDD.n4103 DVDD.n4102 0.00962857
R7855 DVDD.n4102 DVDD.n4068 0.00962857
R7856 DVDD.n4098 DVDD.n4068 0.00962857
R7857 DVDD.n4098 DVDD.n4070 0.00962857
R7858 DVDD.n4094 DVDD.n4070 0.00962857
R7859 DVDD.n4094 DVDD.n4073 0.00962857
R7860 DVDD.n4090 DVDD.n4073 0.00962857
R7861 DVDD.n4090 DVDD.n4075 0.00962857
R7862 DVDD.n4086 DVDD.n4075 0.00962857
R7863 DVDD.n4086 DVDD.n4077 0.00962857
R7864 DVDD.n4082 DVDD.n4077 0.00962857
R7865 DVDD.n3744 DVDD.n3701 0.00962857
R7866 DVDD.n3738 DVDD.n3701 0.00962857
R7867 DVDD.n3738 DVDD.n3737 0.00962857
R7868 DVDD.n3737 DVDD.n3736 0.00962857
R7869 DVDD.n3736 DVDD.n3707 0.00962857
R7870 DVDD.n3730 DVDD.n3707 0.00962857
R7871 DVDD.n3730 DVDD.n3729 0.00962857
R7872 DVDD.n3729 DVDD.n3728 0.00962857
R7873 DVDD.n3728 DVDD.n3711 0.00962857
R7874 DVDD.n3722 DVDD.n3711 0.00962857
R7875 DVDD.n3722 DVDD.n3721 0.00962857
R7876 DVDD.n3721 DVDD.n3720 0.00962857
R7877 DVDD.n3720 DVDD.n3715 0.00962857
R7878 DVDD.n3715 DVDD.n3648 0.00962857
R7879 DVDD.n3957 DVDD.n3648 0.00962857
R7880 DVDD.n3964 DVDD.n3963 0.00962857
R7881 DVDD.n3965 DVDD.n3964 0.00962857
R7882 DVDD.n3965 DVDD.n3640 0.00962857
R7883 DVDD.n3971 DVDD.n3640 0.00962857
R7884 DVDD.n3972 DVDD.n3971 0.00962857
R7885 DVDD.n3973 DVDD.n3972 0.00962857
R7886 DVDD.n3973 DVDD.n3636 0.00962857
R7887 DVDD.n3979 DVDD.n3636 0.00962857
R7888 DVDD.n3980 DVDD.n3979 0.00962857
R7889 DVDD.n3981 DVDD.n3980 0.00962857
R7890 DVDD.n3981 DVDD.n3632 0.00962857
R7891 DVDD.n3987 DVDD.n3632 0.00962857
R7892 DVDD.n3988 DVDD.n3987 0.00962857
R7893 DVDD.n3990 DVDD.n3988 0.00962857
R7894 DVDD.n3990 DVDD.n3989 0.00962857
R7895 DVDD.n4003 DVDD.n4002 0.00962857
R7896 DVDD.n4003 DVDD.n3601 0.00962857
R7897 DVDD.n4009 DVDD.n3601 0.00962857
R7898 DVDD.n4010 DVDD.n4009 0.00962857
R7899 DVDD.n4011 DVDD.n4010 0.00962857
R7900 DVDD.n4011 DVDD.n3597 0.00962857
R7901 DVDD.n4017 DVDD.n3597 0.00962857
R7902 DVDD.n4018 DVDD.n4017 0.00962857
R7903 DVDD.n4019 DVDD.n4018 0.00962857
R7904 DVDD.n4019 DVDD.n3593 0.00962857
R7905 DVDD.n4025 DVDD.n3593 0.00962857
R7906 DVDD.n4026 DVDD.n4025 0.00962857
R7907 DVDD.n4027 DVDD.n4026 0.00962857
R7908 DVDD.n4027 DVDD.n3588 0.00962857
R7909 DVDD.n4034 DVDD.n3588 0.00962857
R7910 DVDD.n4039 DVDD.n4038 0.00962857
R7911 DVDD.n4039 DVDD.n3571 0.00962857
R7912 DVDD.n4045 DVDD.n3571 0.00962857
R7913 DVDD.n4046 DVDD.n4045 0.00962857
R7914 DVDD.n4047 DVDD.n4046 0.00962857
R7915 DVDD.n4047 DVDD.n3567 0.00962857
R7916 DVDD.n4053 DVDD.n3567 0.00962857
R7917 DVDD.n4054 DVDD.n4053 0.00962857
R7918 DVDD.n4055 DVDD.n4054 0.00962857
R7919 DVDD.n4055 DVDD.n3563 0.00962857
R7920 DVDD.n4061 DVDD.n3563 0.00962857
R7921 DVDD.n4062 DVDD.n4061 0.00962857
R7922 DVDD.n4063 DVDD.n4062 0.00962857
R7923 DVDD.n4063 DVDD.n3558 0.00962857
R7924 DVDD.n4108 DVDD.n3558 0.00962857
R7925 DVDD.n4101 DVDD.n3553 0.00962857
R7926 DVDD.n4101 DVDD.n4100 0.00962857
R7927 DVDD.n4100 DVDD.n4099 0.00962857
R7928 DVDD.n4099 DVDD.n4069 0.00962857
R7929 DVDD.n4093 DVDD.n4069 0.00962857
R7930 DVDD.n4093 DVDD.n4092 0.00962857
R7931 DVDD.n4092 DVDD.n4091 0.00962857
R7932 DVDD.n4091 DVDD.n4074 0.00962857
R7933 DVDD.n4085 DVDD.n4074 0.00962857
R7934 DVDD.n4085 DVDD.n4084 0.00962857
R7935 DVDD.n4084 DVDD.n4083 0.00962857
R7936 DVDD.n4327 DVDD.n4326 0.00962857
R7937 DVDD.n4327 DVDD.n3479 0.00962857
R7938 DVDD.n4333 DVDD.n3479 0.00962857
R7939 DVDD.n4334 DVDD.n4333 0.00962857
R7940 DVDD.n4335 DVDD.n4334 0.00962857
R7941 DVDD.n4335 DVDD.n3475 0.00962857
R7942 DVDD.n4341 DVDD.n3475 0.00962857
R7943 DVDD.n4342 DVDD.n4341 0.00962857
R7944 DVDD.n4343 DVDD.n4342 0.00962857
R7945 DVDD.n4343 DVDD.n3471 0.00962857
R7946 DVDD.n4349 DVDD.n3471 0.00962857
R7947 DVDD.n4350 DVDD.n4349 0.00962857
R7948 DVDD.n4352 DVDD.n4350 0.00962857
R7949 DVDD.n4352 DVDD.n4351 0.00962857
R7950 DVDD.n4351 DVDD.n3468 0.00962857
R7951 DVDD.n4360 DVDD.n3464 0.00962857
R7952 DVDD.n4366 DVDD.n3464 0.00962857
R7953 DVDD.n4367 DVDD.n4366 0.00962857
R7954 DVDD.n4368 DVDD.n4367 0.00962857
R7955 DVDD.n4368 DVDD.n3460 0.00962857
R7956 DVDD.n4374 DVDD.n3460 0.00962857
R7957 DVDD.n4375 DVDD.n4374 0.00962857
R7958 DVDD.n4376 DVDD.n4375 0.00962857
R7959 DVDD.n4376 DVDD.n3456 0.00962857
R7960 DVDD.n4382 DVDD.n3456 0.00962857
R7961 DVDD.n4383 DVDD.n4382 0.00962857
R7962 DVDD.n4385 DVDD.n4383 0.00962857
R7963 DVDD.n4385 DVDD.n4384 0.00962857
R7964 DVDD.n4384 DVDD.n3453 0.00962857
R7965 DVDD.n3453 DVDD.n3433 0.00962857
R7966 DVDD.n4485 DVDD.n3448 0.00962857
R7967 DVDD.n4479 DVDD.n3448 0.00962857
R7968 DVDD.n4479 DVDD.n4478 0.00962857
R7969 DVDD.n4478 DVDD.n4477 0.00962857
R7970 DVDD.n4477 DVDD.n4397 0.00962857
R7971 DVDD.n4471 DVDD.n4397 0.00962857
R7972 DVDD.n4471 DVDD.n4470 0.00962857
R7973 DVDD.n4470 DVDD.n4469 0.00962857
R7974 DVDD.n4469 DVDD.n4401 0.00962857
R7975 DVDD.n4463 DVDD.n4401 0.00962857
R7976 DVDD.n4463 DVDD.n4462 0.00962857
R7977 DVDD.n4462 DVDD.n4461 0.00962857
R7978 DVDD.n4461 DVDD.n4405 0.00962857
R7979 DVDD.n4455 DVDD.n4405 0.00962857
R7980 DVDD.n4455 DVDD.n4454 0.00962857
R7981 DVDD.n4447 DVDD.n4412 0.00962857
R7982 DVDD.n4447 DVDD.n4446 0.00962857
R7983 DVDD.n4446 DVDD.n4445 0.00962857
R7984 DVDD.n4445 DVDD.n4413 0.00962857
R7985 DVDD.n4439 DVDD.n4413 0.00962857
R7986 DVDD.n4439 DVDD.n4438 0.00962857
R7987 DVDD.n4438 DVDD.n4437 0.00962857
R7988 DVDD.n4437 DVDD.n4417 0.00962857
R7989 DVDD.n4431 DVDD.n4417 0.00962857
R7990 DVDD.n4431 DVDD.n4430 0.00962857
R7991 DVDD.n4430 DVDD.n4429 0.00962857
R7992 DVDD.n4429 DVDD.n4421 0.00962857
R7993 DVDD.n4423 DVDD.n4421 0.00962857
R7994 DVDD.n4423 DVDD.n15 0.00962857
R7995 DVDD.n5988 DVDD.n15 0.00962857
R7996 DVDD.n5995 DVDD.n5994 0.00962857
R7997 DVDD.n5996 DVDD.n5995 0.00962857
R7998 DVDD.n5996 DVDD.n7 0.00962857
R7999 DVDD.n6002 DVDD.n7 0.00962857
R8000 DVDD.n6003 DVDD.n6002 0.00962857
R8001 DVDD.n6004 DVDD.n6003 0.00962857
R8002 DVDD.n6004 DVDD.n3 0.00962857
R8003 DVDD.n6011 DVDD.n3 0.00962857
R8004 DVDD.n6012 DVDD.n6011 0.00962857
R8005 DVDD.n6013 DVDD.n6012 0.00962857
R8006 DVDD.n6013 DVDD.n0 0.00962857
R8007 DVDD.n4211 DVDD.n3482 0.00962857
R8008 DVDD.n4328 DVDD.n3482 0.00962857
R8009 DVDD.n4328 DVDD.n3480 0.00962857
R8010 DVDD.n4332 DVDD.n3480 0.00962857
R8011 DVDD.n4332 DVDD.n3478 0.00962857
R8012 DVDD.n4336 DVDD.n3478 0.00962857
R8013 DVDD.n4336 DVDD.n3476 0.00962857
R8014 DVDD.n4340 DVDD.n3476 0.00962857
R8015 DVDD.n4340 DVDD.n3474 0.00962857
R8016 DVDD.n4344 DVDD.n3474 0.00962857
R8017 DVDD.n4344 DVDD.n3472 0.00962857
R8018 DVDD.n4348 DVDD.n3472 0.00962857
R8019 DVDD.n4348 DVDD.n3470 0.00962857
R8020 DVDD.n4353 DVDD.n3470 0.00962857
R8021 DVDD.n4353 DVDD.n3467 0.00962857
R8022 DVDD.n4357 DVDD.n3467 0.00962857
R8023 DVDD.n4359 DVDD.n4357 0.00962857
R8024 DVDD.n4361 DVDD.n4359 0.00962857
R8025 DVDD.n4361 DVDD.n3465 0.00962857
R8026 DVDD.n4365 DVDD.n3465 0.00962857
R8027 DVDD.n4365 DVDD.n3463 0.00962857
R8028 DVDD.n4369 DVDD.n3463 0.00962857
R8029 DVDD.n4369 DVDD.n3461 0.00962857
R8030 DVDD.n4373 DVDD.n3461 0.00962857
R8031 DVDD.n4373 DVDD.n3459 0.00962857
R8032 DVDD.n4377 DVDD.n3459 0.00962857
R8033 DVDD.n4377 DVDD.n3457 0.00962857
R8034 DVDD.n4381 DVDD.n3457 0.00962857
R8035 DVDD.n4381 DVDD.n3455 0.00962857
R8036 DVDD.n4386 DVDD.n3455 0.00962857
R8037 DVDD.n4386 DVDD.n3452 0.00962857
R8038 DVDD.n4390 DVDD.n3452 0.00962857
R8039 DVDD.n4391 DVDD.n4390 0.00962857
R8040 DVDD.n4392 DVDD.n4391 0.00962857
R8041 DVDD.n4392 DVDD.n3449 0.00962857
R8042 DVDD.n4484 DVDD.n3449 0.00962857
R8043 DVDD.n4484 DVDD.n3450 0.00962857
R8044 DVDD.n4480 DVDD.n3450 0.00962857
R8045 DVDD.n4480 DVDD.n4396 0.00962857
R8046 DVDD.n4476 DVDD.n4396 0.00962857
R8047 DVDD.n4476 DVDD.n4398 0.00962857
R8048 DVDD.n4472 DVDD.n4398 0.00962857
R8049 DVDD.n4472 DVDD.n4400 0.00962857
R8050 DVDD.n4468 DVDD.n4400 0.00962857
R8051 DVDD.n4468 DVDD.n4402 0.00962857
R8052 DVDD.n4464 DVDD.n4402 0.00962857
R8053 DVDD.n4464 DVDD.n4404 0.00962857
R8054 DVDD.n4460 DVDD.n4404 0.00962857
R8055 DVDD.n4460 DVDD.n4406 0.00962857
R8056 DVDD.n4456 DVDD.n4406 0.00962857
R8057 DVDD.n4456 DVDD.n4453 0.00962857
R8058 DVDD.n4453 DVDD.n4452 0.00962857
R8059 DVDD.n4452 DVDD.n4408 0.00962857
R8060 DVDD.n4448 DVDD.n4408 0.00962857
R8061 DVDD.n4448 DVDD.n4411 0.00962857
R8062 DVDD.n4444 DVDD.n4411 0.00962857
R8063 DVDD.n4444 DVDD.n4414 0.00962857
R8064 DVDD.n4440 DVDD.n4414 0.00962857
R8065 DVDD.n4440 DVDD.n4416 0.00962857
R8066 DVDD.n4436 DVDD.n4416 0.00962857
R8067 DVDD.n4436 DVDD.n4418 0.00962857
R8068 DVDD.n4432 DVDD.n4418 0.00962857
R8069 DVDD.n4432 DVDD.n4420 0.00962857
R8070 DVDD.n4428 DVDD.n4420 0.00962857
R8071 DVDD.n4428 DVDD.n4422 0.00962857
R8072 DVDD.n4424 DVDD.n4422 0.00962857
R8073 DVDD.n4424 DVDD.n14 0.00962857
R8074 DVDD.n5989 DVDD.n14 0.00962857
R8075 DVDD.n5989 DVDD.n12 0.00962857
R8076 DVDD.n5993 DVDD.n12 0.00962857
R8077 DVDD.n5993 DVDD.n10 0.00962857
R8078 DVDD.n5997 DVDD.n10 0.00962857
R8079 DVDD.n5997 DVDD.n8 0.00962857
R8080 DVDD.n6001 DVDD.n8 0.00962857
R8081 DVDD.n6001 DVDD.n6 0.00962857
R8082 DVDD.n6005 DVDD.n6 0.00962857
R8083 DVDD.n6005 DVDD.n4 0.00962857
R8084 DVDD.n6010 DVDD.n4 0.00962857
R8085 DVDD.n6010 DVDD.n2 0.00962857
R8086 DVDD.n6014 DVDD.n2 0.00962857
R8087 DVDD.n6015 DVDD.n6014 0.00962857
R8088 DVDD.n5027 DVDD.n5015 0.009275
R8089 DVDD.n4521 DVDD.n3145 0.009275
R8090 DVDD.n4900 DVDD.n4899 0.009275
R8091 DVDD.n5292 DVDD.n4926 0.009275
R8092 DVDD.n2751 DVDD.n2747 0.00917857
R8093 DVDD.n4035 DVDD.n4034 0.00917857
R8094 DVDD.n4454 DVDD.n3426 0.00917857
R8095 DVDD.n5505 DVDD.n333 0.00906343
R8096 DVDD.n5499 DVDD.n5498 0.00905
R8097 DVDD.n2932 DVDD.n2931 0.00905
R8098 DVDD.n5502 DVDD.n576 0.00905
R8099 DVDD.n2611 DVDD.n2610 0.00905
R8100 DVDD.n5510 DVDD.n565 0.00905
R8101 DVDD.n5617 DVDD.n5616 0.00905
R8102 DVDD.n5513 DVDD.n561 0.00905
R8103 DVDD.n2592 DVDD.n473 0.00905
R8104 DVDD.n5615 DVDD.n481 0.00892143
R8105 DVDD.n3963 DVDD.n3644 0.00892143
R8106 DVDD.n4360 DVDD.n3373 0.00892143
R8107 DVDD.n858 DVDD.n848 0.0084875
R8108 DVDD.n858 DVDD.n857 0.0084875
R8109 DVDD.n857 DVDD.n856 0.0084875
R8110 DVDD.n856 DVDD.n263 0.0084875
R8111 DVDD.n5696 DVDD.n279 0.0084875
R8112 DVDD.n5696 DVDD.n5695 0.0084875
R8113 DVDD.n5695 DVDD.n5694 0.0084875
R8114 DVDD.n5694 DVDD.n280 0.0084875
R8115 DVDD.n5687 DVDD.n5686 0.0084875
R8116 DVDD.n5686 DVDD.n5685 0.0084875
R8117 DVDD.n5685 DVDD.n288 0.0084875
R8118 DVDD.n5679 DVDD.n288 0.0084875
R8119 DVDD.n5679 DVDD.n5678 0.0084875
R8120 DVDD.n5678 DVDD.n5677 0.0084875
R8121 DVDD.n5677 DVDD.n292 0.0084875
R8122 DVDD.n5671 DVDD.n292 0.0084875
R8123 DVDD.n5671 DVDD.n5670 0.0084875
R8124 DVDD.n5038 DVDD.n5037 0.0084875
R8125 DVDD.n5038 DVDD.n5008 0.0084875
R8126 DVDD.n5044 DVDD.n5008 0.0084875
R8127 DVDD.n5045 DVDD.n5044 0.0084875
R8128 DVDD.n5046 DVDD.n5045 0.0084875
R8129 DVDD.n5046 DVDD.n5004 0.0084875
R8130 DVDD.n5052 DVDD.n5004 0.0084875
R8131 DVDD.n5053 DVDD.n5052 0.0084875
R8132 DVDD.n5055 DVDD.n5053 0.0084875
R8133 DVDD.n5055 DVDD.n5054 0.0084875
R8134 DVDD.n5066 DVDD.n5061 0.0084875
R8135 DVDD.n5066 DVDD.n5065 0.0084875
R8136 DVDD.n5065 DVDD.n5064 0.0084875
R8137 DVDD.n5064 DVDD.n628 0.0084875
R8138 DVDD.n5462 DVDD.n644 0.0084875
R8139 DVDD.n5462 DVDD.n5461 0.0084875
R8140 DVDD.n5461 DVDD.n5460 0.0084875
R8141 DVDD.n5452 DVDD.n5451 0.0084875
R8142 DVDD.n5451 DVDD.n5450 0.0084875
R8143 DVDD.n5450 DVDD.n649 0.0084875
R8144 DVDD.n5444 DVDD.n649 0.0084875
R8145 DVDD.n5444 DVDD.n5443 0.0084875
R8146 DVDD.n5443 DVDD.n5442 0.0084875
R8147 DVDD.n5442 DVDD.n653 0.0084875
R8148 DVDD.n5436 DVDD.n653 0.0084875
R8149 DVDD.n695 DVDD.n662 0.0084875
R8150 DVDD.n666 DVDD.n662 0.0084875
R8151 DVDD.n688 DVDD.n666 0.0084875
R8152 DVDD.n688 DVDD.n687 0.0084875
R8153 DVDD.n687 DVDD.n686 0.0084875
R8154 DVDD.n686 DVDD.n667 0.0084875
R8155 DVDD.n680 DVDD.n667 0.0084875
R8156 DVDD.n680 DVDD.n679 0.0084875
R8157 DVDD.n679 DVDD.n678 0.0084875
R8158 DVDD.n5453 DVDD.n648 0.0084875
R8159 DVDD.n5449 DVDD.n648 0.0084875
R8160 DVDD.n5449 DVDD.n650 0.0084875
R8161 DVDD.n5445 DVDD.n650 0.0084875
R8162 DVDD.n5445 DVDD.n652 0.0084875
R8163 DVDD.n5441 DVDD.n652 0.0084875
R8164 DVDD.n5441 DVDD.n654 0.0084875
R8165 DVDD.n5437 DVDD.n654 0.0084875
R8166 DVDD.n5437 DVDD.n5435 0.0084875
R8167 DVDD.n5435 DVDD.n5433 0.0084875
R8168 DVDD.n694 DVDD.n693 0.0084875
R8169 DVDD.n693 DVDD.n663 0.0084875
R8170 DVDD.n689 DVDD.n663 0.0084875
R8171 DVDD.n689 DVDD.n665 0.0084875
R8172 DVDD.n685 DVDD.n665 0.0084875
R8173 DVDD.n685 DVDD.n668 0.0084875
R8174 DVDD.n681 DVDD.n668 0.0084875
R8175 DVDD.n681 DVDD.n670 0.0084875
R8176 DVDD.n677 DVDD.n670 0.0084875
R8177 DVDD.n5039 DVDD.n5036 0.0084875
R8178 DVDD.n5039 DVDD.n5009 0.0084875
R8179 DVDD.n5043 DVDD.n5009 0.0084875
R8180 DVDD.n5043 DVDD.n5007 0.0084875
R8181 DVDD.n5047 DVDD.n5007 0.0084875
R8182 DVDD.n5047 DVDD.n5005 0.0084875
R8183 DVDD.n5051 DVDD.n5005 0.0084875
R8184 DVDD.n5051 DVDD.n5003 0.0084875
R8185 DVDD.n5056 DVDD.n5003 0.0084875
R8186 DVDD.n5056 DVDD.n5000 0.0084875
R8187 DVDD.n5067 DVDD.n5001 0.0084875
R8188 DVDD.n5067 DVDD.n5060 0.0084875
R8189 DVDD.n5063 DVDD.n5060 0.0084875
R8190 DVDD.n5063 DVDD.n639 0.0084875
R8191 DVDD.n5467 DVDD.n639 0.0084875
R8192 DVDD.n5467 DVDD.n640 0.0084875
R8193 DVDD.n5463 DVDD.n640 0.0084875
R8194 DVDD.n5463 DVDD.n643 0.0084875
R8195 DVDD.n5459 DVDD.n643 0.0084875
R8196 DVDD.n860 DVDD.n859 0.0084875
R8197 DVDD.n859 DVDD.n852 0.0084875
R8198 DVDD.n855 DVDD.n852 0.0084875
R8199 DVDD.n855 DVDD.n274 0.0084875
R8200 DVDD.n5701 DVDD.n274 0.0084875
R8201 DVDD.n5701 DVDD.n275 0.0084875
R8202 DVDD.n5697 DVDD.n275 0.0084875
R8203 DVDD.n5697 DVDD.n278 0.0084875
R8204 DVDD.n5693 DVDD.n278 0.0084875
R8205 DVDD.n5693 DVDD.n281 0.0084875
R8206 DVDD.n5688 DVDD.n286 0.0084875
R8207 DVDD.n5684 DVDD.n286 0.0084875
R8208 DVDD.n5684 DVDD.n289 0.0084875
R8209 DVDD.n5680 DVDD.n289 0.0084875
R8210 DVDD.n5680 DVDD.n291 0.0084875
R8211 DVDD.n5676 DVDD.n291 0.0084875
R8212 DVDD.n5676 DVDD.n293 0.0084875
R8213 DVDD.n5672 DVDD.n293 0.0084875
R8214 DVDD.n5672 DVDD.n295 0.0084875
R8215 DVDD.n808 DVDD.n800 0.0084875
R8216 DVDD.n808 DVDD.n798 0.0084875
R8217 DVDD.n812 DVDD.n798 0.0084875
R8218 DVDD.n812 DVDD.n796 0.0084875
R8219 DVDD.n816 DVDD.n796 0.0084875
R8220 DVDD.n816 DVDD.n794 0.0084875
R8221 DVDD.n820 DVDD.n794 0.0084875
R8222 DVDD.n820 DVDD.n792 0.0084875
R8223 DVDD.n825 DVDD.n792 0.0084875
R8224 DVDD.n825 DVDD.n788 0.0084875
R8225 DVDD.n2976 DVDD.n789 0.0084875
R8226 DVDD.n879 DVDD.n789 0.0084875
R8227 DVDD.n879 DVDD.n840 0.0084875
R8228 DVDD.n875 DVDD.n840 0.0084875
R8229 DVDD.n875 DVDD.n843 0.0084875
R8230 DVDD.n871 DVDD.n843 0.0084875
R8231 DVDD.n871 DVDD.n845 0.0084875
R8232 DVDD.n867 DVDD.n845 0.0084875
R8233 DVDD.n867 DVDD.n847 0.0084875
R8234 DVDD.n809 DVDD.n799 0.0084875
R8235 DVDD.n810 DVDD.n809 0.0084875
R8236 DVDD.n811 DVDD.n810 0.0084875
R8237 DVDD.n811 DVDD.n795 0.0084875
R8238 DVDD.n817 DVDD.n795 0.0084875
R8239 DVDD.n818 DVDD.n817 0.0084875
R8240 DVDD.n819 DVDD.n818 0.0084875
R8241 DVDD.n819 DVDD.n791 0.0084875
R8242 DVDD.n826 DVDD.n791 0.0084875
R8243 DVDD.n827 DVDD.n826 0.0084875
R8244 DVDD.n880 DVDD.n839 0.0084875
R8245 DVDD.n874 DVDD.n839 0.0084875
R8246 DVDD.n874 DVDD.n873 0.0084875
R8247 DVDD.n873 DVDD.n872 0.0084875
R8248 DVDD.n872 DVDD.n844 0.0084875
R8249 DVDD.n866 DVDD.n844 0.0084875
R8250 DVDD.n866 DVDD.n865 0.0084875
R8251 DVDD.n1737 DVDD.n342 0.00839179
R8252 DVDD.n1495 DVDD.n1494 0.00839179
R8253 DVDD.n2937 DVDD.n2936 0.00815
R8254 DVDD.n2938 DVDD.n441 0.00815
R8255 DVDD.n2946 DVDD.n2945 0.00815
R8256 DVDD.n2943 DVDD.n460 0.00815
R8257 DVDD.n5469 DVDD.n628 0.00809375
R8258 DVDD.n5569 DVDD.n5568 0.00802143
R8259 DVDD.n2754 DVDD.n2607 0.00802143
R8260 DVDD.n4001 DVDD.n3605 0.00802143
R8261 DVDD.n4037 DVDD.n3575 0.00802143
R8262 DVDD.n4488 DVDD.n3441 0.00802143
R8263 DVDD.n4409 DVDD.n3427 0.00802143
R8264 DVDD.n279 DVDD.n273 0.00786875
R8265 DVDD.n2688 DVDD 0.00782857
R8266 DVDD.n2689 DVDD 0.00782857
R8267 DVDD.n4082 DVDD 0.00782857
R8268 DVDD.n4083 DVDD 0.00782857
R8269 DVDD DVDD.n0 0.00782857
R8270 DVDD.n6015 DVDD 0.00782857
R8271 DVDD.n5612 DVDD.n478 0.00776429
R8272 DVDD.n2595 DVDD.n506 0.00776429
R8273 DVDD.n3956 DVDD.n3654 0.00776429
R8274 DVDD.n3997 DVDD.n3627 0.00776429
R8275 DVDD.n4358 DVDD.n3374 0.00776429
R8276 DVDD.n4493 DVDD.n3438 0.00776429
R8277 DVDD.n2296 DVDD.n2295 0.00772462
R8278 DVDD.n1652 DVDD.n1651 0.00772462
R8279 DVDD.n2259 DVDD.n2258 0.00772462
R8280 DVDD.n1349 DVDD.n1348 0.00772462
R8281 DVDD.n5412 DVDD.n5411 0.00772462
R8282 DVDD.n5321 DVDD.n731 0.00770384
R8283 DVDD.n5745 DVDD.n194 0.00770384
R8284 DVDD.n850 DVDD.n847 0.0077
R8285 DVDD.n865 DVDD.n864 0.0077
R8286 DVDD.n4883 DVDD.n178 0.00755224
R8287 DVDD.n5665 DVDD.n301 0.007475
R8288 DVDD.n4527 DVDD.n4499 0.007475
R8289 DVDD.n5317 DVDD.n4905 0.007475
R8290 DVDD.n4920 DVDD.n4919 0.007475
R8291 DVDD.n5670 DVDD.n5669 0.00725
R8292 DVDD.n5035 DVDD.n295 0.00725
R8293 DVDD.n2228 DVDD.n1387 0.00725
R8294 DVDD.n1247 DVDD.n1245 0.00725
R8295 DVDD.n1388 DVDD.n378 0.00725
R8296 DVDD.n1248 DVDD.n395 0.00725
R8297 DVDD.n1390 DVDD.n917 0.00725
R8298 DVDD.n1241 DVDD.n934 0.00725
R8299 DVDD.n2222 DVDD.n1391 0.00725
R8300 DVDD.n1242 DVDD.n1135 0.00725
R8301 DVDD.n5396 DVDD.n695 0.0071375
R8302 DVDD.n694 DVDD.n656 0.0071375
R8303 DVDD.n4722 DVDD.n4721 0.0071
R8304 DVDD.n4793 DVDD.n4792 0.0071
R8305 DVDD.n4888 DVDD.n3137 0.0071
R8306 DVDD.n3208 DVDD.n3207 0.0071
R8307 DVDD.n5468 DVDD.n638 0.00708125
R8308 DVDD.n1714 DVDD.n345 0.00704851
R8309 DVDD.n1509 DVDD.n1508 0.00704851
R8310 DVDD.n5703 DVDD.n5702 0.00685625
R8311 DVDD.n5460 DVDD.n645 0.0068
R8312 DVDD.n5459 DVDD.n646 0.0068
R8313 DVDD.n5737 DVDD.n5736 0.00678
R8314 DVDD.n3093 DVDD.n3092 0.00678
R8315 DVDD.n5098 DVDD.n5084 0.00678
R8316 DVDD.n5333 DVDD.n710 0.00678
R8317 DVDD.n5061 DVDD.n4997 0.0066875
R8318 DVDD.n5224 DVDD.n5001 0.0066875
R8319 DVDD.n4329 DVDD.n3481 0.00658571
R8320 DVDD.n4330 DVDD.n4329 0.00658571
R8321 DVDD.n4331 DVDD.n4330 0.00658571
R8322 DVDD.n4331 DVDD.n3477 0.00658571
R8323 DVDD.n4337 DVDD.n3477 0.00658571
R8324 DVDD.n4338 DVDD.n4337 0.00658571
R8325 DVDD.n4339 DVDD.n4338 0.00658571
R8326 DVDD.n4339 DVDD.n3473 0.00658571
R8327 DVDD.n4345 DVDD.n3473 0.00658571
R8328 DVDD.n4346 DVDD.n4345 0.00658571
R8329 DVDD.n4347 DVDD.n4346 0.00658571
R8330 DVDD.n4347 DVDD.n3469 0.00658571
R8331 DVDD.n4354 DVDD.n3469 0.00658571
R8332 DVDD.n4355 DVDD.n4354 0.00658571
R8333 DVDD.n4356 DVDD.n4355 0.00658571
R8334 DVDD.n4356 DVDD.n3466 0.00658571
R8335 DVDD.n4362 DVDD.n3466 0.00658571
R8336 DVDD.n4363 DVDD.n4362 0.00658571
R8337 DVDD.n4364 DVDD.n4363 0.00658571
R8338 DVDD.n4364 DVDD.n3462 0.00658571
R8339 DVDD.n4370 DVDD.n3462 0.00658571
R8340 DVDD.n4371 DVDD.n4370 0.00658571
R8341 DVDD.n4372 DVDD.n4371 0.00658571
R8342 DVDD.n4372 DVDD.n3458 0.00658571
R8343 DVDD.n4378 DVDD.n3458 0.00658571
R8344 DVDD.n4379 DVDD.n4378 0.00658571
R8345 DVDD.n4380 DVDD.n4379 0.00658571
R8346 DVDD.n4380 DVDD.n3454 0.00658571
R8347 DVDD.n4387 DVDD.n3454 0.00658571
R8348 DVDD.n4388 DVDD.n4387 0.00658571
R8349 DVDD.n4389 DVDD.n4388 0.00658571
R8350 DVDD.n4389 DVDD.n3451 0.00658571
R8351 DVDD.n4393 DVDD.n3451 0.00658571
R8352 DVDD.n4394 DVDD.n4393 0.00658571
R8353 DVDD.n4483 DVDD.n4394 0.00658571
R8354 DVDD.n4483 DVDD.n4482 0.00658571
R8355 DVDD.n4482 DVDD.n4481 0.00658571
R8356 DVDD.n4481 DVDD.n4395 0.00658571
R8357 DVDD.n4475 DVDD.n4395 0.00658571
R8358 DVDD.n4475 DVDD.n4474 0.00658571
R8359 DVDD.n4474 DVDD.n4473 0.00658571
R8360 DVDD.n4473 DVDD.n4399 0.00658571
R8361 DVDD.n4467 DVDD.n4399 0.00658571
R8362 DVDD.n4467 DVDD.n4466 0.00658571
R8363 DVDD.n4466 DVDD.n4465 0.00658571
R8364 DVDD.n4465 DVDD.n4403 0.00658571
R8365 DVDD.n4459 DVDD.n4403 0.00658571
R8366 DVDD.n4459 DVDD.n4458 0.00658571
R8367 DVDD.n4458 DVDD.n4457 0.00658571
R8368 DVDD.n4457 DVDD.n4407 0.00658571
R8369 DVDD.n4451 DVDD.n4407 0.00658571
R8370 DVDD.n4451 DVDD.n4450 0.00658571
R8371 DVDD.n4450 DVDD.n4449 0.00658571
R8372 DVDD.n4449 DVDD.n4410 0.00658571
R8373 DVDD.n4443 DVDD.n4410 0.00658571
R8374 DVDD.n4443 DVDD.n4442 0.00658571
R8375 DVDD.n4442 DVDD.n4441 0.00658571
R8376 DVDD.n4441 DVDD.n4415 0.00658571
R8377 DVDD.n4435 DVDD.n4415 0.00658571
R8378 DVDD.n4435 DVDD.n4434 0.00658571
R8379 DVDD.n4434 DVDD.n4433 0.00658571
R8380 DVDD.n4433 DVDD.n4419 0.00658571
R8381 DVDD.n4427 DVDD.n4419 0.00658571
R8382 DVDD.n4427 DVDD.n4426 0.00658571
R8383 DVDD.n4426 DVDD.n4425 0.00658571
R8384 DVDD.n4425 DVDD.n13 0.00658571
R8385 DVDD.n5990 DVDD.n13 0.00658571
R8386 DVDD.n5991 DVDD.n5990 0.00658571
R8387 DVDD.n5992 DVDD.n5991 0.00658571
R8388 DVDD.n5992 DVDD.n9 0.00658571
R8389 DVDD.n5998 DVDD.n9 0.00658571
R8390 DVDD.n5999 DVDD.n5998 0.00658571
R8391 DVDD.n6000 DVDD.n5999 0.00658571
R8392 DVDD.n6000 DVDD.n5 0.00658571
R8393 DVDD.n6006 DVDD.n5 0.00658571
R8394 DVDD.n6007 DVDD.n6006 0.00658571
R8395 DVDD.n6009 DVDD.n6007 0.00658571
R8396 DVDD.n6009 DVDD.n6008 0.00658571
R8397 DVDD.n6008 DVDD.n1 0.00658571
R8398 DVDD.n6016 DVDD.n1 0.00658571
R8399 DVDD.n6017 DVDD.n6016 0.00658571
R8400 DVDD.n2866 DVDD.n2864 0.00658571
R8401 DVDD.n2869 DVDD.n2866 0.00658571
R8402 DVDD.n2898 DVDD.n2869 0.00658571
R8403 DVDD.n2898 DVDD.n2897 0.00658571
R8404 DVDD.n2897 DVDD.n2896 0.00658571
R8405 DVDD.n2896 DVDD.n2870 0.00658571
R8406 DVDD.n2890 DVDD.n2870 0.00658571
R8407 DVDD.n2890 DVDD.n2889 0.00658571
R8408 DVDD.n2889 DVDD.n2888 0.00658571
R8409 DVDD.n2888 DVDD.n2874 0.00658571
R8410 DVDD.n2882 DVDD.n2874 0.00658571
R8411 DVDD.n2882 DVDD.n2881 0.00658571
R8412 DVDD.n2881 DVDD.n2880 0.00658571
R8413 DVDD.n2880 DVDD.n490 0.00658571
R8414 DVDD.n5606 DVDD.n490 0.00658571
R8415 DVDD.n5606 DVDD.n5605 0.00658571
R8416 DVDD.n5605 DVDD.n5604 0.00658571
R8417 DVDD.n5604 DVDD.n491 0.00658571
R8418 DVDD.n495 DVDD.n491 0.00658571
R8419 DVDD.n5597 DVDD.n495 0.00658571
R8420 DVDD.n5597 DVDD.n5596 0.00658571
R8421 DVDD.n5596 DVDD.n5595 0.00658571
R8422 DVDD.n5595 DVDD.n496 0.00658571
R8423 DVDD.n5589 DVDD.n496 0.00658571
R8424 DVDD.n5589 DVDD.n5588 0.00658571
R8425 DVDD.n5588 DVDD.n5587 0.00658571
R8426 DVDD.n5587 DVDD.n500 0.00658571
R8427 DVDD.n5581 DVDD.n500 0.00658571
R8428 DVDD.n5581 DVDD.n5580 0.00658571
R8429 DVDD.n5580 DVDD.n5579 0.00658571
R8430 DVDD.n5579 DVDD.n504 0.00658571
R8431 DVDD.n5573 DVDD.n504 0.00658571
R8432 DVDD.n5573 DVDD.n5572 0.00658571
R8433 DVDD.n5572 DVDD.n5571 0.00658571
R8434 DVDD.n5571 DVDD.n508 0.00658571
R8435 DVDD.n2632 DVDD.n508 0.00658571
R8436 DVDD.n2633 DVDD.n2632 0.00658571
R8437 DVDD.n2634 DVDD.n2633 0.00658571
R8438 DVDD.n2634 DVDD.n2626 0.00658571
R8439 DVDD.n2640 DVDD.n2626 0.00658571
R8440 DVDD.n2641 DVDD.n2640 0.00658571
R8441 DVDD.n2642 DVDD.n2641 0.00658571
R8442 DVDD.n2642 DVDD.n2622 0.00658571
R8443 DVDD.n2648 DVDD.n2622 0.00658571
R8444 DVDD.n2649 DVDD.n2648 0.00658571
R8445 DVDD.n2650 DVDD.n2649 0.00658571
R8446 DVDD.n2650 DVDD.n2618 0.00658571
R8447 DVDD.n2656 DVDD.n2618 0.00658571
R8448 DVDD.n2657 DVDD.n2656 0.00658571
R8449 DVDD.n2745 DVDD.n2657 0.00658571
R8450 DVDD.n2745 DVDD.n2744 0.00658571
R8451 DVDD.n2744 DVDD.n2743 0.00658571
R8452 DVDD.n2743 DVDD.n2658 0.00658571
R8453 DVDD.n2662 DVDD.n2658 0.00658571
R8454 DVDD.n2736 DVDD.n2662 0.00658571
R8455 DVDD.n2736 DVDD.n2735 0.00658571
R8456 DVDD.n2735 DVDD.n2734 0.00658571
R8457 DVDD.n2734 DVDD.n2663 0.00658571
R8458 DVDD.n2728 DVDD.n2663 0.00658571
R8459 DVDD.n2728 DVDD.n2727 0.00658571
R8460 DVDD.n2727 DVDD.n2726 0.00658571
R8461 DVDD.n2726 DVDD.n2667 0.00658571
R8462 DVDD.n2720 DVDD.n2667 0.00658571
R8463 DVDD.n2720 DVDD.n2719 0.00658571
R8464 DVDD.n2719 DVDD.n2718 0.00658571
R8465 DVDD.n2718 DVDD.n2671 0.00658571
R8466 DVDD.n2712 DVDD.n2671 0.00658571
R8467 DVDD.n2712 DVDD.n2711 0.00658571
R8468 DVDD.n2711 DVDD.n2710 0.00658571
R8469 DVDD.n2710 DVDD.n2673 0.00658571
R8470 DVDD.n2677 DVDD.n2673 0.00658571
R8471 DVDD.n2703 DVDD.n2677 0.00658571
R8472 DVDD.n2703 DVDD.n2702 0.00658571
R8473 DVDD.n2702 DVDD.n2701 0.00658571
R8474 DVDD.n2701 DVDD.n2678 0.00658571
R8475 DVDD.n2695 DVDD.n2678 0.00658571
R8476 DVDD.n2695 DVDD.n2694 0.00658571
R8477 DVDD.n2694 DVDD.n2693 0.00658571
R8478 DVDD.n2693 DVDD.n2682 0.00658571
R8479 DVDD.n2687 DVDD.n2682 0.00658571
R8480 DVDD.n3742 DVDD.n3741 0.00658571
R8481 DVDD.n3741 DVDD.n3740 0.00658571
R8482 DVDD.n3740 DVDD.n3705 0.00658571
R8483 DVDD.n3734 DVDD.n3705 0.00658571
R8484 DVDD.n3734 DVDD.n3733 0.00658571
R8485 DVDD.n3733 DVDD.n3732 0.00658571
R8486 DVDD.n3732 DVDD.n3709 0.00658571
R8487 DVDD.n3726 DVDD.n3709 0.00658571
R8488 DVDD.n3726 DVDD.n3725 0.00658571
R8489 DVDD.n3725 DVDD.n3724 0.00658571
R8490 DVDD.n3724 DVDD.n3713 0.00658571
R8491 DVDD.n3718 DVDD.n3713 0.00658571
R8492 DVDD.n3718 DVDD.n3717 0.00658571
R8493 DVDD.n3717 DVDD.n3646 0.00658571
R8494 DVDD.n3959 DVDD.n3646 0.00658571
R8495 DVDD.n3960 DVDD.n3959 0.00658571
R8496 DVDD.n3961 DVDD.n3960 0.00658571
R8497 DVDD.n3961 DVDD.n3642 0.00658571
R8498 DVDD.n3967 DVDD.n3642 0.00658571
R8499 DVDD.n3968 DVDD.n3967 0.00658571
R8500 DVDD.n3969 DVDD.n3968 0.00658571
R8501 DVDD.n3969 DVDD.n3638 0.00658571
R8502 DVDD.n3975 DVDD.n3638 0.00658571
R8503 DVDD.n3976 DVDD.n3975 0.00658571
R8504 DVDD.n3977 DVDD.n3976 0.00658571
R8505 DVDD.n3977 DVDD.n3634 0.00658571
R8506 DVDD.n3983 DVDD.n3634 0.00658571
R8507 DVDD.n3984 DVDD.n3983 0.00658571
R8508 DVDD.n3985 DVDD.n3984 0.00658571
R8509 DVDD.n3985 DVDD.n3630 0.00658571
R8510 DVDD.n3992 DVDD.n3630 0.00658571
R8511 DVDD.n3993 DVDD.n3992 0.00658571
R8512 DVDD.n3995 DVDD.n3993 0.00658571
R8513 DVDD.n3995 DVDD.n3994 0.00658571
R8514 DVDD.n3994 DVDD.n3603 0.00658571
R8515 DVDD.n4005 DVDD.n3603 0.00658571
R8516 DVDD.n4006 DVDD.n4005 0.00658571
R8517 DVDD.n4007 DVDD.n4006 0.00658571
R8518 DVDD.n4007 DVDD.n3599 0.00658571
R8519 DVDD.n4013 DVDD.n3599 0.00658571
R8520 DVDD.n4014 DVDD.n4013 0.00658571
R8521 DVDD.n4015 DVDD.n4014 0.00658571
R8522 DVDD.n4015 DVDD.n3595 0.00658571
R8523 DVDD.n4021 DVDD.n3595 0.00658571
R8524 DVDD.n4022 DVDD.n4021 0.00658571
R8525 DVDD.n4023 DVDD.n4022 0.00658571
R8526 DVDD.n4023 DVDD.n3591 0.00658571
R8527 DVDD.n4029 DVDD.n3591 0.00658571
R8528 DVDD.n4030 DVDD.n4029 0.00658571
R8529 DVDD.n4032 DVDD.n4030 0.00658571
R8530 DVDD.n4032 DVDD.n4031 0.00658571
R8531 DVDD.n4031 DVDD.n3573 0.00658571
R8532 DVDD.n4041 DVDD.n3573 0.00658571
R8533 DVDD.n4042 DVDD.n4041 0.00658571
R8534 DVDD.n4043 DVDD.n4042 0.00658571
R8535 DVDD.n4043 DVDD.n3569 0.00658571
R8536 DVDD.n4049 DVDD.n3569 0.00658571
R8537 DVDD.n4050 DVDD.n4049 0.00658571
R8538 DVDD.n4051 DVDD.n4050 0.00658571
R8539 DVDD.n4051 DVDD.n3565 0.00658571
R8540 DVDD.n4057 DVDD.n3565 0.00658571
R8541 DVDD.n4058 DVDD.n4057 0.00658571
R8542 DVDD.n4059 DVDD.n4058 0.00658571
R8543 DVDD.n4059 DVDD.n3561 0.00658571
R8544 DVDD.n4065 DVDD.n3561 0.00658571
R8545 DVDD.n4066 DVDD.n4065 0.00658571
R8546 DVDD.n4106 DVDD.n4066 0.00658571
R8547 DVDD.n4106 DVDD.n4105 0.00658571
R8548 DVDD.n4105 DVDD.n4104 0.00658571
R8549 DVDD.n4104 DVDD.n4067 0.00658571
R8550 DVDD.n4071 DVDD.n4067 0.00658571
R8551 DVDD.n4097 DVDD.n4071 0.00658571
R8552 DVDD.n4097 DVDD.n4096 0.00658571
R8553 DVDD.n4096 DVDD.n4095 0.00658571
R8554 DVDD.n4095 DVDD.n4072 0.00658571
R8555 DVDD.n4089 DVDD.n4072 0.00658571
R8556 DVDD.n4089 DVDD.n4088 0.00658571
R8557 DVDD.n4088 DVDD.n4087 0.00658571
R8558 DVDD.n4087 DVDD.n4076 0.00658571
R8559 DVDD.n4081 DVDD.n4076 0.00658571
R8560 DVDD.n4081 DVDD.n4080 0.00658571
R8561 DVDD.n2172 DVDD.n1452 0.0065
R8562 DVDD.n1586 DVDD.n1062 0.0065
R8563 DVDD.n1855 DVDD.n1775 0.0065
R8564 DVDD.n2172 DVDD.n1176 0.0065
R8565 DVDD.n1776 DVDD.n1774 0.0065
R8566 DVDD.n2393 DVDD.n1172 0.0065
R8567 DVDD.n1784 DVDD.n1776 0.0065
R8568 DVDD.n2393 DVDD.n1173 0.0065
R8569 DVDD.n2132 DVDD.n2057 0.0065
R8570 DVDD.n2016 DVDD.n1173 0.0065
R8571 DVDD.n1785 DVDD.n1784 0.0065
R8572 DVDD.n1670 DVDD.n1328 0.0065
R8573 DVDD.n1328 DVDD.n1321 0.0065
R8574 DVDD.n2132 DVDD.n1065 0.0065
R8575 DVDD.n1065 DVDD.n1060 0.0065
R8576 DVDD.n2314 DVDD.n1321 0.0065
R8577 DVDD.n1857 DVDD.n1855 0.0065
R8578 DVDD.n1906 DVDD.n1176 0.0065
R8579 DVDD.n2279 DVDD.n2278 0.0065
R8580 DVDD.n2492 DVDD.n1062 0.0065
R8581 DVDD.n2493 DVDD.n2492 0.0065
R8582 DVDD.n2277 DVDD.n1325 0.0065
R8583 DVDD.n2278 DVDD.n2277 0.0065
R8584 DVDD.n1780 DVDD.n1775 0.0065
R8585 DVDD.n566 DVDD.n323 0.00637687
R8586 DVDD.n2585 DVDD.n522 0.00637687
R8587 DVDD.n2927 DVDD.n2583 0.00635
R8588 DVDD.n678 DVDD.n671 0.00635
R8589 DVDD.n677 DVDD.n672 0.00635
R8590 DVDD.n4112 DVDD.n4108 0.00635
R8591 DVDD.n5988 DVDD.n5987 0.00635
R8592 DVDD.n5687 DVDD.n287 0.0062375
R8593 DVDD.n5688 DVDD.n285 0.0062375
R8594 DVDD.n2914 DVDD.n2591 0.00609286
R8595 DVDD.n3745 DVDD.n3744 0.00609286
R8596 DVDD.n4326 DVDD.n4325 0.00609286
R8597 DVDD.n2565 DVDD.n1014 0.00604104
R8598 DVDD.n4183 DVDD.n16 0.0059
R8599 DVDD.n4207 DVDD.n3505 0.0059
R8600 DVDD.n731 DVDD 0.00587887
R8601 DVDD DVDD.n194 0.00587887
R8602 DVDD.n5454 DVDD.n647 0.005825
R8603 DVDD.n5448 DVDD.n647 0.005825
R8604 DVDD.n5448 DVDD.n5447 0.005825
R8605 DVDD.n5447 DVDD.n5446 0.005825
R8606 DVDD.n5446 DVDD.n651 0.005825
R8607 DVDD.n5440 DVDD.n651 0.005825
R8608 DVDD.n5440 DVDD.n5439 0.005825
R8609 DVDD.n5439 DVDD.n5438 0.005825
R8610 DVDD.n5438 DVDD.n655 0.005825
R8611 DVDD.n5432 DVDD.n655 0.005825
R8612 DVDD.n692 DVDD.n658 0.005825
R8613 DVDD.n692 DVDD.n691 0.005825
R8614 DVDD.n691 DVDD.n690 0.005825
R8615 DVDD.n690 DVDD.n664 0.005825
R8616 DVDD.n684 DVDD.n664 0.005825
R8617 DVDD.n684 DVDD.n683 0.005825
R8618 DVDD.n683 DVDD.n682 0.005825
R8619 DVDD.n682 DVDD.n669 0.005825
R8620 DVDD.n676 DVDD.n669 0.005825
R8621 DVDD.n5040 DVDD.n5010 0.005825
R8622 DVDD.n5041 DVDD.n5040 0.005825
R8623 DVDD.n5042 DVDD.n5041 0.005825
R8624 DVDD.n5042 DVDD.n5006 0.005825
R8625 DVDD.n5048 DVDD.n5006 0.005825
R8626 DVDD.n5049 DVDD.n5048 0.005825
R8627 DVDD.n5050 DVDD.n5049 0.005825
R8628 DVDD.n5050 DVDD.n5002 0.005825
R8629 DVDD.n5057 DVDD.n5002 0.005825
R8630 DVDD.n5058 DVDD.n5057 0.005825
R8631 DVDD.n5069 DVDD.n5068 0.005825
R8632 DVDD.n5068 DVDD.n5059 0.005825
R8633 DVDD.n5062 DVDD.n5059 0.005825
R8634 DVDD.n5062 DVDD.n641 0.005825
R8635 DVDD.n5466 DVDD.n641 0.005825
R8636 DVDD.n5466 DVDD.n5465 0.005825
R8637 DVDD.n5465 DVDD.n5464 0.005825
R8638 DVDD.n5464 DVDD.n642 0.005825
R8639 DVDD.n5458 DVDD.n642 0.005825
R8640 DVDD.n861 DVDD.n851 0.005825
R8641 DVDD.n853 DVDD.n851 0.005825
R8642 DVDD.n854 DVDD.n853 0.005825
R8643 DVDD.n854 DVDD.n276 0.005825
R8644 DVDD.n5700 DVDD.n276 0.005825
R8645 DVDD.n5700 DVDD.n5699 0.005825
R8646 DVDD.n5699 DVDD.n5698 0.005825
R8647 DVDD.n5698 DVDD.n277 0.005825
R8648 DVDD.n5692 DVDD.n277 0.005825
R8649 DVDD.n5692 DVDD.n5691 0.005825
R8650 DVDD.n5689 DVDD.n284 0.005825
R8651 DVDD.n5683 DVDD.n284 0.005825
R8652 DVDD.n5683 DVDD.n5682 0.005825
R8653 DVDD.n5682 DVDD.n5681 0.005825
R8654 DVDD.n5681 DVDD.n290 0.005825
R8655 DVDD.n5675 DVDD.n290 0.005825
R8656 DVDD.n5675 DVDD.n5674 0.005825
R8657 DVDD.n5674 DVDD.n5673 0.005825
R8658 DVDD.n5673 DVDD.n294 0.005825
R8659 DVDD.n807 DVDD.n806 0.005825
R8660 DVDD.n807 DVDD.n797 0.005825
R8661 DVDD.n813 DVDD.n797 0.005825
R8662 DVDD.n814 DVDD.n813 0.005825
R8663 DVDD.n815 DVDD.n814 0.005825
R8664 DVDD.n815 DVDD.n793 0.005825
R8665 DVDD.n821 DVDD.n793 0.005825
R8666 DVDD.n822 DVDD.n821 0.005825
R8667 DVDD.n824 DVDD.n822 0.005825
R8668 DVDD.n824 DVDD.n823 0.005825
R8669 DVDD.n841 DVDD.n790 0.005825
R8670 DVDD.n878 DVDD.n841 0.005825
R8671 DVDD.n878 DVDD.n877 0.005825
R8672 DVDD.n877 DVDD.n876 0.005825
R8673 DVDD.n876 DVDD.n842 0.005825
R8674 DVDD.n870 DVDD.n842 0.005825
R8675 DVDD.n870 DVDD.n869 0.005825
R8676 DVDD.n869 DVDD.n868 0.005825
R8677 DVDD.n868 DVDD.n846 0.005825
R8678 DVDD.n2977 DVDD.n2976 0.0057875
R8679 DVDD.n2975 DVDD.n828 0.0057875
R8680 DVDD.n1523 DVDD.n1522 0.00570522
R8681 DVDD.n5436 DVDD.n605 0.00561875
R8682 DVDD.n3874 DVDD.n3580 0.00545
R8683 DVDD.n3661 DVDD.n3653 0.00545
R8684 DVDD.n2972 DVDD.n880 0.00539375
R8685 DVDD.n2687 DVDD 0.00538571
R8686 DVDD.n729 DVDD.n184 0.00530256
R8687 DVDD.n862 DVDD.n846 0.0053
R8688 DVDD.n3307 DVDD.n3257 0.00523684
R8689 DVDD.n3305 DVDD.n3303 0.00523684
R8690 DVDD.n4642 DVDD.n3397 0.00523684
R8691 DVDD.n3400 DVDD.n3398 0.00523684
R8692 DVDD.n5028 DVDD.n5014 0.005225
R8693 DVDD.n4878 DVDD.n4877 0.005225
R8694 DVDD.n182 DVDD.n181 0.005225
R8695 DVDD.n4931 DVDD.n4930 0.005225
R8696 DVDD.n2930 DVDD.n2575 0.00519286
R8697 DVDD.n4115 DVDD.n3552 0.00519286
R8698 DVDD.n17 DVDD.n11 0.00519286
R8699 DVDD.n2759 DVDD.n520 0.00503358
R8700 DVDD.n5032 DVDD.n294 0.005
R8701 DVDD.n4193 DVDD.n4192 0.005
R8702 DVDD.n3517 DVDD.n3516 0.005
R8703 DVDD.n2602 DVDD.n2601 0.00498219
R8704 DVDD.n3999 DVDD.n3998 0.00498219
R8705 DVDD.n3999 DVDD.n3622 0.00498219
R8706 DVDD.n2602 DVDD.n510 0.00498219
R8707 DVDD.n4491 DVDD.n3432 0.00498219
R8708 DVDD.n3445 DVDD.n3432 0.00498219
R8709 DVDD.n2911 DVDD.n2589 0.00493571
R8710 DVDD.n2930 DVDD.n2578 0.00493571
R8711 DVDD.n3700 DVDD.n3699 0.00493571
R8712 DVDD.n4115 DVDD.n3553 0.00493571
R8713 DVDD.n4322 DVDD.n3483 0.00493571
R8714 DVDD.n5994 DVDD.n11 0.00493571
R8715 DVDD.n5431 DVDD.n658 0.004925
R8716 DVDD.n1846 DVDD.n1845 0.00476
R8717 DVDD.n1845 DVDD.n1844 0.00476
R8718 DVDD.n1844 DVDD.n1787 0.00476
R8719 DVDD.n1840 DVDD.n1787 0.00476
R8720 DVDD.n1840 DVDD.n1839 0.00476
R8721 DVDD.n1839 DVDD.n1838 0.00476
R8722 DVDD.n1838 DVDD.n1804 0.00476
R8723 DVDD.n1834 DVDD.n1804 0.00476
R8724 DVDD.n1834 DVDD.n1833 0.00476
R8725 DVDD.n1833 DVDD.n1832 0.00476
R8726 DVDD.n1832 DVDD.n1810 0.00476
R8727 DVDD.n1828 DVDD.n1810 0.00476
R8728 DVDD.n1828 DVDD.n1827 0.00476
R8729 DVDD.n1827 DVDD.n1826 0.00476
R8730 DVDD.n1826 DVDD.n1816 0.00476
R8731 DVDD.n1822 DVDD.n1816 0.00476
R8732 DVDD.n1822 DVDD.n1821 0.00476
R8733 DVDD.n1821 DVDD.n1745 0.00476
R8734 DVDD.n2023 DVDD.n1745 0.00476
R8735 DVDD.n2023 DVDD.n2022 0.00476
R8736 DVDD.n2022 DVDD.n2021 0.00476
R8737 DVDD.n2021 DVDD.n1749 0.00476
R8738 DVDD.n2017 DVDD.n1749 0.00476
R8739 DVDD.n2015 DVDD.n1947 0.00476
R8740 DVDD.n2011 DVDD.n1947 0.00476
R8741 DVDD.n2011 DVDD.n2010 0.00476
R8742 DVDD.n2010 DVDD.n2009 0.00476
R8743 DVDD.n2009 DVDD.n1953 0.00476
R8744 DVDD.n2005 DVDD.n1953 0.00476
R8745 DVDD.n2005 DVDD.n2004 0.00476
R8746 DVDD.n2004 DVDD.n2003 0.00476
R8747 DVDD.n2003 DVDD.n2000 0.00476
R8748 DVDD.n2000 DVDD.n1999 0.00476
R8749 DVDD.n1999 DVDD.n1998 0.00476
R8750 DVDD.n1998 DVDD.n1997 0.00476
R8751 DVDD.n1997 DVDD.n1995 0.00476
R8752 DVDD.n1995 DVDD.n1964 0.00476
R8753 DVDD.n1991 DVDD.n1964 0.00476
R8754 DVDD.n1991 DVDD.n1990 0.00476
R8755 DVDD.n1990 DVDD.n1989 0.00476
R8756 DVDD.n1989 DVDD.n1970 0.00476
R8757 DVDD.n1985 DVDD.n1970 0.00476
R8758 DVDD.n1985 DVDD.n1984 0.00476
R8759 DVDD.n1984 DVDD.n1983 0.00476
R8760 DVDD.n1983 DVDD.n1979 0.00476
R8761 DVDD.n1979 DVDD.n1583 0.00476
R8762 DVDD.n2056 DVDD.n1585 0.00476
R8763 DVDD.n2052 DVDD.n1585 0.00476
R8764 DVDD.n2052 DVDD.n2051 0.00476
R8765 DVDD.n2051 DVDD.n2050 0.00476
R8766 DVDD.n2050 DVDD.n1592 0.00476
R8767 DVDD.n1696 DVDD.n1592 0.00476
R8768 DVDD.n1696 DVDD.n1695 0.00476
R8769 DVDD.n1695 DVDD.n1694 0.00476
R8770 DVDD.n1694 DVDD.n1613 0.00476
R8771 DVDD.n1690 DVDD.n1613 0.00476
R8772 DVDD.n1690 DVDD.n1689 0.00476
R8773 DVDD.n1689 DVDD.n1688 0.00476
R8774 DVDD.n1688 DVDD.n1619 0.00476
R8775 DVDD.n1684 DVDD.n1619 0.00476
R8776 DVDD.n1684 DVDD.n1683 0.00476
R8777 DVDD.n1683 DVDD.n1682 0.00476
R8778 DVDD.n1682 DVDD.n1625 0.00476
R8779 DVDD.n1678 DVDD.n1625 0.00476
R8780 DVDD.n1678 DVDD.n1677 0.00476
R8781 DVDD.n1677 DVDD.n1676 0.00476
R8782 DVDD.n1676 DVDD.n1673 0.00476
R8783 DVDD.n1673 DVDD.n1672 0.00476
R8784 DVDD.n1672 DVDD.n1671 0.00476
R8785 DVDD.n1669 DVDD.n1635 0.00476
R8786 DVDD.n1665 DVDD.n1635 0.00476
R8787 DVDD.n1665 DVDD.n1664 0.00476
R8788 DVDD.n1664 DVDD.n1663 0.00476
R8789 DVDD.n1663 DVDD.n1641 0.00476
R8790 DVDD.n1659 DVDD.n1641 0.00476
R8791 DVDD.n1659 DVDD.n1658 0.00476
R8792 DVDD.n1658 DVDD.n1657 0.00476
R8793 DVDD.n1657 DVDD.n1647 0.00476
R8794 DVDD.n1653 DVDD.n1647 0.00476
R8795 DVDD.n1783 DVDD.n1410 0.00476
R8796 DVDD.n2204 DVDD.n1410 0.00476
R8797 DVDD.n2204 DVDD.n2203 0.00476
R8798 DVDD.n2203 DVDD.n2202 0.00476
R8799 DVDD.n2202 DVDD.n1414 0.00476
R8800 DVDD.n2198 DVDD.n1414 0.00476
R8801 DVDD.n2198 DVDD.n2197 0.00476
R8802 DVDD.n2197 DVDD.n2196 0.00476
R8803 DVDD.n2196 DVDD.n1420 0.00476
R8804 DVDD.n2192 DVDD.n1420 0.00476
R8805 DVDD.n2192 DVDD.n2191 0.00476
R8806 DVDD.n2191 DVDD.n2190 0.00476
R8807 DVDD.n2190 DVDD.n1426 0.00476
R8808 DVDD.n2186 DVDD.n1426 0.00476
R8809 DVDD.n2186 DVDD.n2185 0.00476
R8810 DVDD.n2185 DVDD.n2184 0.00476
R8811 DVDD.n2184 DVDD.n2182 0.00476
R8812 DVDD.n2182 DVDD.n2181 0.00476
R8813 DVDD.n2181 DVDD.n2180 0.00476
R8814 DVDD.n2180 DVDD.n1435 0.00476
R8815 DVDD.n2176 DVDD.n1435 0.00476
R8816 DVDD.n2176 DVDD.n2175 0.00476
R8817 DVDD.n2175 DVDD.n2174 0.00476
R8818 DVDD.n2170 DVDD.n2169 0.00476
R8819 DVDD.n2169 DVDD.n2168 0.00476
R8820 DVDD.n2168 DVDD.n1457 0.00476
R8821 DVDD.n2164 DVDD.n1457 0.00476
R8822 DVDD.n2164 DVDD.n2163 0.00476
R8823 DVDD.n2163 DVDD.n2162 0.00476
R8824 DVDD.n2162 DVDD.n1463 0.00476
R8825 DVDD.n2158 DVDD.n1463 0.00476
R8826 DVDD.n2158 DVDD.n2157 0.00476
R8827 DVDD.n2157 DVDD.n2156 0.00476
R8828 DVDD.n2156 DVDD.n1469 0.00476
R8829 DVDD.n2150 DVDD.n1469 0.00476
R8830 DVDD.n2150 DVDD.n2149 0.00476
R8831 DVDD.n2149 DVDD.n1568 0.00476
R8832 DVDD.n2145 DVDD.n1568 0.00476
R8833 DVDD.n2145 DVDD.n2144 0.00476
R8834 DVDD.n2144 DVDD.n2143 0.00476
R8835 DVDD.n2143 DVDD.n1574 0.00476
R8836 DVDD.n2139 DVDD.n1574 0.00476
R8837 DVDD.n2139 DVDD.n2138 0.00476
R8838 DVDD.n2138 DVDD.n2137 0.00476
R8839 DVDD.n2137 DVDD.n1580 0.00476
R8840 DVDD.n2133 DVDD.n1580 0.00476
R8841 DVDD.n2131 DVDD.n2059 0.00476
R8842 DVDD.n2127 DVDD.n2059 0.00476
R8843 DVDD.n2127 DVDD.n2126 0.00476
R8844 DVDD.n2126 DVDD.n2125 0.00476
R8845 DVDD.n2125 DVDD.n2124 0.00476
R8846 DVDD.n2124 DVDD.n2123 0.00476
R8847 DVDD.n2123 DVDD.n2067 0.00476
R8848 DVDD.n2119 DVDD.n2067 0.00476
R8849 DVDD.n2119 DVDD.n2118 0.00476
R8850 DVDD.n2118 DVDD.n2117 0.00476
R8851 DVDD.n2117 DVDD.n2084 0.00476
R8852 DVDD.n2113 DVDD.n2084 0.00476
R8853 DVDD.n2113 DVDD.n2112 0.00476
R8854 DVDD.n2112 DVDD.n2111 0.00476
R8855 DVDD.n2111 DVDD.n2090 0.00476
R8856 DVDD.n2107 DVDD.n2090 0.00476
R8857 DVDD.n2107 DVDD.n2106 0.00476
R8858 DVDD.n2106 DVDD.n2105 0.00476
R8859 DVDD.n2105 DVDD.n2096 0.00476
R8860 DVDD.n2101 DVDD.n2096 0.00476
R8861 DVDD.n2101 DVDD.n1369 0.00476
R8862 DVDD.n2238 DVDD.n1369 0.00476
R8863 DVDD.n2239 DVDD.n2238 0.00476
R8864 DVDD.n2275 DVDD.n2274 0.00476
R8865 DVDD.n2274 DVDD.n2273 0.00476
R8866 DVDD.n2273 DVDD.n2245 0.00476
R8867 DVDD.n2269 DVDD.n2245 0.00476
R8868 DVDD.n2269 DVDD.n2268 0.00476
R8869 DVDD.n2268 DVDD.n2267 0.00476
R8870 DVDD.n2267 DVDD.n2251 0.00476
R8871 DVDD.n2263 DVDD.n2251 0.00476
R8872 DVDD.n2263 DVDD.n2262 0.00476
R8873 DVDD.n2262 DVDD.n2261 0.00476
R8874 DVDD.n1851 DVDD.n1141 0.00476
R8875 DVDD.n2424 DVDD.n1141 0.00476
R8876 DVDD.n2424 DVDD.n2423 0.00476
R8877 DVDD.n2423 DVDD.n2422 0.00476
R8878 DVDD.n2422 DVDD.n1145 0.00476
R8879 DVDD.n2418 DVDD.n1145 0.00476
R8880 DVDD.n2418 DVDD.n2417 0.00476
R8881 DVDD.n2417 DVDD.n2416 0.00476
R8882 DVDD.n2416 DVDD.n1151 0.00476
R8883 DVDD.n2412 DVDD.n1151 0.00476
R8884 DVDD.n2412 DVDD.n2411 0.00476
R8885 DVDD.n2411 DVDD.n2410 0.00476
R8886 DVDD.n2410 DVDD.n1157 0.00476
R8887 DVDD.n2406 DVDD.n1157 0.00476
R8888 DVDD.n2406 DVDD.n2405 0.00476
R8889 DVDD.n2405 DVDD.n2404 0.00476
R8890 DVDD.n2404 DVDD.n2402 0.00476
R8891 DVDD.n2402 DVDD.n2401 0.00476
R8892 DVDD.n2401 DVDD.n2400 0.00476
R8893 DVDD.n2400 DVDD.n2399 0.00476
R8894 DVDD.n2399 DVDD.n1167 0.00476
R8895 DVDD.n2395 DVDD.n1167 0.00476
R8896 DVDD.n2395 DVDD.n2394 0.00476
R8897 DVDD.n2392 DVDD.n1175 0.00476
R8898 DVDD.n2388 DVDD.n1175 0.00476
R8899 DVDD.n2388 DVDD.n2387 0.00476
R8900 DVDD.n2387 DVDD.n2386 0.00476
R8901 DVDD.n2386 DVDD.n1182 0.00476
R8902 DVDD.n2382 DVDD.n1182 0.00476
R8903 DVDD.n2382 DVDD.n2381 0.00476
R8904 DVDD.n2381 DVDD.n2380 0.00476
R8905 DVDD.n2380 DVDD.n1188 0.00476
R8906 DVDD.n2376 DVDD.n1188 0.00476
R8907 DVDD.n2376 DVDD.n2375 0.00476
R8908 DVDD.n2375 DVDD.n1193 0.00476
R8909 DVDD.n2367 DVDD.n1193 0.00476
R8910 DVDD.n2367 DVDD.n2366 0.00476
R8911 DVDD.n2366 DVDD.n2365 0.00476
R8912 DVDD.n2365 DVDD.n1278 0.00476
R8913 DVDD.n2361 DVDD.n1278 0.00476
R8914 DVDD.n2361 DVDD.n2360 0.00476
R8915 DVDD.n2360 DVDD.n2359 0.00476
R8916 DVDD.n2359 DVDD.n1284 0.00476
R8917 DVDD.n2355 DVDD.n1284 0.00476
R8918 DVDD.n2355 DVDD.n2354 0.00476
R8919 DVDD.n2354 DVDD.n2353 0.00476
R8920 DVDD.n2490 DVDD.n2489 0.00476
R8921 DVDD.n2489 DVDD.n2488 0.00476
R8922 DVDD.n2488 DVDD.n2485 0.00476
R8923 DVDD.n2485 DVDD.n2484 0.00476
R8924 DVDD.n2484 DVDD.n2483 0.00476
R8925 DVDD.n2483 DVDD.n2482 0.00476
R8926 DVDD.n2482 DVDD.n2481 0.00476
R8927 DVDD.n2481 DVDD.n1074 0.00476
R8928 DVDD.n2477 DVDD.n1074 0.00476
R8929 DVDD.n2477 DVDD.n2476 0.00476
R8930 DVDD.n2476 DVDD.n2475 0.00476
R8931 DVDD.n2475 DVDD.n1080 0.00476
R8932 DVDD.n2471 DVDD.n1080 0.00476
R8933 DVDD.n2471 DVDD.n2470 0.00476
R8934 DVDD.n2470 DVDD.n2469 0.00476
R8935 DVDD.n2469 DVDD.n1086 0.00476
R8936 DVDD.n2465 DVDD.n1086 0.00476
R8937 DVDD.n2465 DVDD.n2464 0.00476
R8938 DVDD.n2464 DVDD.n2463 0.00476
R8939 DVDD.n2463 DVDD.n1092 0.00476
R8940 DVDD.n2459 DVDD.n1092 0.00476
R8941 DVDD.n2459 DVDD.n2458 0.00476
R8942 DVDD.n2458 DVDD.n1097 0.00476
R8943 DVDD.n1365 DVDD.n1364 0.00476
R8944 DVDD.n1364 DVDD.n1333 0.00476
R8945 DVDD.n1360 DVDD.n1333 0.00476
R8946 DVDD.n1360 DVDD.n1359 0.00476
R8947 DVDD.n1359 DVDD.n1358 0.00476
R8948 DVDD.n1358 DVDD.n1339 0.00476
R8949 DVDD.n1354 DVDD.n1339 0.00476
R8950 DVDD.n1354 DVDD.n1353 0.00476
R8951 DVDD.n1353 DVDD.n1352 0.00476
R8952 DVDD.n1352 DVDD.n1345 0.00476
R8953 DVDD.n1859 DVDD.n1772 0.00476
R8954 DVDD.n1863 DVDD.n1772 0.00476
R8955 DVDD.n1864 DVDD.n1863 0.00476
R8956 DVDD.n1867 DVDD.n1864 0.00476
R8957 DVDD.n1867 DVDD.n1770 0.00476
R8958 DVDD.n1871 DVDD.n1770 0.00476
R8959 DVDD.n1871 DVDD.n1768 0.00476
R8960 DVDD.n1875 DVDD.n1768 0.00476
R8961 DVDD.n1875 DVDD.n1766 0.00476
R8962 DVDD.n1879 DVDD.n1766 0.00476
R8963 DVDD.n1879 DVDD.n1764 0.00476
R8964 DVDD.n1883 DVDD.n1764 0.00476
R8965 DVDD.n1883 DVDD.n1762 0.00476
R8966 DVDD.n1887 DVDD.n1762 0.00476
R8967 DVDD.n1887 DVDD.n1760 0.00476
R8968 DVDD.n1891 DVDD.n1760 0.00476
R8969 DVDD.n1891 DVDD.n1758 0.00476
R8970 DVDD.n1895 DVDD.n1758 0.00476
R8971 DVDD.n1896 DVDD.n1895 0.00476
R8972 DVDD.n1899 DVDD.n1896 0.00476
R8973 DVDD.n1899 DVDD.n1756 0.00476
R8974 DVDD.n1903 DVDD.n1756 0.00476
R8975 DVDD.n1904 DVDD.n1903 0.00476
R8976 DVDD.n1940 DVDD.n1754 0.00476
R8977 DVDD.n1936 DVDD.n1754 0.00476
R8978 DVDD.n1936 DVDD.n1935 0.00476
R8979 DVDD.n1935 DVDD.n1934 0.00476
R8980 DVDD.n1934 DVDD.n1911 0.00476
R8981 DVDD.n1930 DVDD.n1911 0.00476
R8982 DVDD.n1930 DVDD.n1929 0.00476
R8983 DVDD.n1929 DVDD.n1928 0.00476
R8984 DVDD.n1928 DVDD.n1917 0.00476
R8985 DVDD.n1924 DVDD.n1917 0.00476
R8986 DVDD.n1924 DVDD.n1923 0.00476
R8987 DVDD.n1923 DVDD.n1044 0.00476
R8988 DVDD.n2509 DVDD.n1044 0.00476
R8989 DVDD.n2509 DVDD.n2508 0.00476
R8990 DVDD.n2508 DVDD.n2507 0.00476
R8991 DVDD.n2507 DVDD.n1048 0.00476
R8992 DVDD.n2503 DVDD.n1048 0.00476
R8993 DVDD.n2503 DVDD.n2502 0.00476
R8994 DVDD.n2502 DVDD.n2501 0.00476
R8995 DVDD.n2501 DVDD.n1054 0.00476
R8996 DVDD.n2497 DVDD.n1054 0.00476
R8997 DVDD.n2497 DVDD.n2496 0.00476
R8998 DVDD.n2496 DVDD.n2495 0.00476
R8999 DVDD.n2348 DVDD.n2347 0.00476
R9000 DVDD.n2347 DVDD.n1291 0.00476
R9001 DVDD.n2343 DVDD.n1291 0.00476
R9002 DVDD.n2343 DVDD.n2342 0.00476
R9003 DVDD.n2342 DVDD.n2341 0.00476
R9004 DVDD.n2341 DVDD.n2340 0.00476
R9005 DVDD.n2340 DVDD.n2339 0.00476
R9006 DVDD.n2339 DVDD.n1298 0.00476
R9007 DVDD.n2335 DVDD.n1298 0.00476
R9008 DVDD.n2335 DVDD.n2334 0.00476
R9009 DVDD.n2334 DVDD.n2333 0.00476
R9010 DVDD.n2333 DVDD.n1304 0.00476
R9011 DVDD.n2329 DVDD.n1304 0.00476
R9012 DVDD.n2329 DVDD.n2328 0.00476
R9013 DVDD.n2328 DVDD.n2327 0.00476
R9014 DVDD.n2327 DVDD.n1310 0.00476
R9015 DVDD.n2323 DVDD.n1310 0.00476
R9016 DVDD.n2323 DVDD.n2322 0.00476
R9017 DVDD.n2322 DVDD.n2321 0.00476
R9018 DVDD.n2321 DVDD.n1316 0.00476
R9019 DVDD.n2317 DVDD.n1316 0.00476
R9020 DVDD.n2317 DVDD.n2316 0.00476
R9021 DVDD.n2316 DVDD.n2315 0.00476
R9022 DVDD.n2313 DVDD.n1323 0.00476
R9023 DVDD.n2309 DVDD.n1323 0.00476
R9024 DVDD.n2309 DVDD.n2308 0.00476
R9025 DVDD.n2308 DVDD.n2307 0.00476
R9026 DVDD.n2307 DVDD.n2285 0.00476
R9027 DVDD.n2303 DVDD.n2285 0.00476
R9028 DVDD.n2303 DVDD.n2302 0.00476
R9029 DVDD.n2302 DVDD.n2301 0.00476
R9030 DVDD.n2301 DVDD.n2291 0.00476
R9031 DVDD.n2297 DVDD.n2291 0.00476
R9032 DVDD.n1865 DVDD.n454 0.00476
R9033 DVDD.n1866 DVDD.n1865 0.00476
R9034 DVDD.n1866 DVDD.n1769 0.00476
R9035 DVDD.n1872 DVDD.n1769 0.00476
R9036 DVDD.n1873 DVDD.n1872 0.00476
R9037 DVDD.n1874 DVDD.n1873 0.00476
R9038 DVDD.n1874 DVDD.n1765 0.00476
R9039 DVDD.n1880 DVDD.n1765 0.00476
R9040 DVDD.n1881 DVDD.n1880 0.00476
R9041 DVDD.n1882 DVDD.n1881 0.00476
R9042 DVDD.n1882 DVDD.n1761 0.00476
R9043 DVDD.n1888 DVDD.n1761 0.00476
R9044 DVDD.n1889 DVDD.n1888 0.00476
R9045 DVDD.n1890 DVDD.n1889 0.00476
R9046 DVDD.n1890 DVDD.n952 0.00476
R9047 DVDD.n1898 DVDD.n972 0.00476
R9048 DVDD.n1898 DVDD.n1897 0.00476
R9049 DVDD.n1897 DVDD.n1755 0.00476
R9050 DVDD.n1905 DVDD.n1755 0.00476
R9051 DVDD.n1939 DVDD.n1938 0.00476
R9052 DVDD.n1938 DVDD.n1937 0.00476
R9053 DVDD.n1937 DVDD.n1907 0.00476
R9054 DVDD.n1933 DVDD.n1907 0.00476
R9055 DVDD.n1933 DVDD.n1932 0.00476
R9056 DVDD.n1932 DVDD.n1931 0.00476
R9057 DVDD.n1931 DVDD.n1912 0.00476
R9058 DVDD.n1927 DVDD.n1912 0.00476
R9059 DVDD.n1927 DVDD.n1926 0.00476
R9060 DVDD.n1926 DVDD.n1925 0.00476
R9061 DVDD.n2510 DVDD.n1043 0.00476
R9062 DVDD.n2506 DVDD.n1043 0.00476
R9063 DVDD.n2506 DVDD.n2505 0.00476
R9064 DVDD.n2505 DVDD.n2504 0.00476
R9065 DVDD.n2504 DVDD.n1049 0.00476
R9066 DVDD.n2500 DVDD.n1049 0.00476
R9067 DVDD.n2500 DVDD.n2499 0.00476
R9068 DVDD.n2499 DVDD.n2498 0.00476
R9069 DVDD.n2498 DVDD.n1055 0.00476
R9070 DVDD.n2494 DVDD.n1055 0.00476
R9071 DVDD.n2346 DVDD.n1061 0.00476
R9072 DVDD.n2346 DVDD.n2345 0.00476
R9073 DVDD.n2345 DVDD.n2344 0.00476
R9074 DVDD.n2344 DVDD.n413 0.00476
R9075 DVDD.n2338 DVDD.n436 0.00476
R9076 DVDD.n2338 DVDD.n2337 0.00476
R9077 DVDD.n2337 DVDD.n2336 0.00476
R9078 DVDD.n2336 DVDD.n1299 0.00476
R9079 DVDD.n2332 DVDD.n1299 0.00476
R9080 DVDD.n2332 DVDD.n2331 0.00476
R9081 DVDD.n2331 DVDD.n2330 0.00476
R9082 DVDD.n2330 DVDD.n1305 0.00476
R9083 DVDD.n2326 DVDD.n1305 0.00476
R9084 DVDD.n2326 DVDD.n2325 0.00476
R9085 DVDD.n2325 DVDD.n2324 0.00476
R9086 DVDD.n2324 DVDD.n1311 0.00476
R9087 DVDD.n2320 DVDD.n1311 0.00476
R9088 DVDD.n2320 DVDD.n2319 0.00476
R9089 DVDD.n2319 DVDD.n2318 0.00476
R9090 DVDD.n2312 DVDD.n2311 0.00476
R9091 DVDD.n2311 DVDD.n2310 0.00476
R9092 DVDD.n2310 DVDD.n2280 0.00476
R9093 DVDD.n2306 DVDD.n2280 0.00476
R9094 DVDD.n2306 DVDD.n2305 0.00476
R9095 DVDD.n2305 DVDD.n2304 0.00476
R9096 DVDD.n2304 DVDD.n2286 0.00476
R9097 DVDD.n2300 DVDD.n2286 0.00476
R9098 DVDD.n2300 DVDD.n2299 0.00476
R9099 DVDD.n2299 DVDD.n2298 0.00476
R9100 DVDD.n2425 DVDD.n1140 0.00476
R9101 DVDD.n2421 DVDD.n1140 0.00476
R9102 DVDD.n2421 DVDD.n2420 0.00476
R9103 DVDD.n2420 DVDD.n2419 0.00476
R9104 DVDD.n2419 DVDD.n1146 0.00476
R9105 DVDD.n2415 DVDD.n1146 0.00476
R9106 DVDD.n2415 DVDD.n2414 0.00476
R9107 DVDD.n2414 DVDD.n2413 0.00476
R9108 DVDD.n2413 DVDD.n1152 0.00476
R9109 DVDD.n2409 DVDD.n1152 0.00476
R9110 DVDD.n2409 DVDD.n2408 0.00476
R9111 DVDD.n2408 DVDD.n2407 0.00476
R9112 DVDD.n2407 DVDD.n1158 0.00476
R9113 DVDD.n2403 DVDD.n1158 0.00476
R9114 DVDD.n2403 DVDD.n922 0.00476
R9115 DVDD.n2398 DVDD.n940 0.00476
R9116 DVDD.n2398 DVDD.n2397 0.00476
R9117 DVDD.n2397 DVDD.n2396 0.00476
R9118 DVDD.n2396 DVDD.n1168 0.00476
R9119 DVDD.n2391 DVDD.n2390 0.00476
R9120 DVDD.n2390 DVDD.n2389 0.00476
R9121 DVDD.n2389 DVDD.n1177 0.00476
R9122 DVDD.n2385 DVDD.n1177 0.00476
R9123 DVDD.n2385 DVDD.n2384 0.00476
R9124 DVDD.n2384 DVDD.n2383 0.00476
R9125 DVDD.n2383 DVDD.n1183 0.00476
R9126 DVDD.n2379 DVDD.n1183 0.00476
R9127 DVDD.n2379 DVDD.n2378 0.00476
R9128 DVDD.n2378 DVDD.n2377 0.00476
R9129 DVDD.n2368 DVDD.n1273 0.00476
R9130 DVDD.n2364 DVDD.n1273 0.00476
R9131 DVDD.n2364 DVDD.n2363 0.00476
R9132 DVDD.n2363 DVDD.n2362 0.00476
R9133 DVDD.n2362 DVDD.n1279 0.00476
R9134 DVDD.n2358 DVDD.n1279 0.00476
R9135 DVDD.n2358 DVDD.n2357 0.00476
R9136 DVDD.n2357 DVDD.n2356 0.00476
R9137 DVDD.n2356 DVDD.n1285 0.00476
R9138 DVDD.n1285 DVDD.n1063 0.00476
R9139 DVDD.n2491 DVDD.n1064 0.00476
R9140 DVDD.n2487 DVDD.n1064 0.00476
R9141 DVDD.n2487 DVDD.n2486 0.00476
R9142 DVDD.n2486 DVDD.n383 0.00476
R9143 DVDD.n2480 DVDD.n401 0.00476
R9144 DVDD.n2480 DVDD.n2479 0.00476
R9145 DVDD.n2479 DVDD.n2478 0.00476
R9146 DVDD.n2478 DVDD.n1075 0.00476
R9147 DVDD.n2474 DVDD.n1075 0.00476
R9148 DVDD.n2474 DVDD.n2473 0.00476
R9149 DVDD.n2473 DVDD.n2472 0.00476
R9150 DVDD.n2472 DVDD.n1081 0.00476
R9151 DVDD.n2468 DVDD.n1081 0.00476
R9152 DVDD.n2468 DVDD.n2467 0.00476
R9153 DVDD.n2467 DVDD.n2466 0.00476
R9154 DVDD.n2466 DVDD.n1087 0.00476
R9155 DVDD.n2462 DVDD.n1087 0.00476
R9156 DVDD.n2462 DVDD.n2461 0.00476
R9157 DVDD.n2461 DVDD.n2460 0.00476
R9158 DVDD.n1363 DVDD.n1324 0.00476
R9159 DVDD.n1363 DVDD.n1362 0.00476
R9160 DVDD.n1362 DVDD.n1361 0.00476
R9161 DVDD.n1361 DVDD.n1334 0.00476
R9162 DVDD.n1357 DVDD.n1334 0.00476
R9163 DVDD.n1357 DVDD.n1356 0.00476
R9164 DVDD.n1356 DVDD.n1355 0.00476
R9165 DVDD.n1355 DVDD.n1340 0.00476
R9166 DVDD.n1351 DVDD.n1340 0.00476
R9167 DVDD.n1351 DVDD.n1350 0.00476
R9168 DVDD.n2205 DVDD.n1409 0.00476
R9169 DVDD.n2201 DVDD.n1409 0.00476
R9170 DVDD.n2201 DVDD.n2200 0.00476
R9171 DVDD.n2200 DVDD.n2199 0.00476
R9172 DVDD.n2199 DVDD.n1415 0.00476
R9173 DVDD.n2195 DVDD.n1415 0.00476
R9174 DVDD.n2195 DVDD.n2194 0.00476
R9175 DVDD.n2194 DVDD.n2193 0.00476
R9176 DVDD.n2193 DVDD.n1421 0.00476
R9177 DVDD.n2189 DVDD.n1421 0.00476
R9178 DVDD.n2189 DVDD.n2188 0.00476
R9179 DVDD.n2188 DVDD.n2187 0.00476
R9180 DVDD.n2187 DVDD.n1427 0.00476
R9181 DVDD.n2183 DVDD.n1427 0.00476
R9182 DVDD.n2183 DVDD.n901 0.00476
R9183 DVDD.n2179 DVDD.n2178 0.00476
R9184 DVDD.n2178 DVDD.n2177 0.00476
R9185 DVDD.n2177 DVDD.n1447 0.00476
R9186 DVDD.n2173 DVDD.n1447 0.00476
R9187 DVDD.n2171 DVDD.n1453 0.00476
R9188 DVDD.n2167 DVDD.n1453 0.00476
R9189 DVDD.n2167 DVDD.n2166 0.00476
R9190 DVDD.n2166 DVDD.n2165 0.00476
R9191 DVDD.n2165 DVDD.n1458 0.00476
R9192 DVDD.n2161 DVDD.n1458 0.00476
R9193 DVDD.n2161 DVDD.n2160 0.00476
R9194 DVDD.n2160 DVDD.n2159 0.00476
R9195 DVDD.n2159 DVDD.n1464 0.00476
R9196 DVDD.n2155 DVDD.n1464 0.00476
R9197 DVDD.n2148 DVDD.n2147 0.00476
R9198 DVDD.n2147 DVDD.n2146 0.00476
R9199 DVDD.n2146 DVDD.n1569 0.00476
R9200 DVDD.n2142 DVDD.n1569 0.00476
R9201 DVDD.n2142 DVDD.n2141 0.00476
R9202 DVDD.n2141 DVDD.n2140 0.00476
R9203 DVDD.n2140 DVDD.n1575 0.00476
R9204 DVDD.n2136 DVDD.n1575 0.00476
R9205 DVDD.n2136 DVDD.n2135 0.00476
R9206 DVDD.n2135 DVDD.n2134 0.00476
R9207 DVDD.n2130 DVDD.n2129 0.00476
R9208 DVDD.n2129 DVDD.n2128 0.00476
R9209 DVDD.n2128 DVDD.n2060 0.00476
R9210 DVDD.n2060 DVDD.n362 0.00476
R9211 DVDD.n2122 DVDD.n2121 0.00476
R9212 DVDD.n2121 DVDD.n2120 0.00476
R9213 DVDD.n2120 DVDD.n2079 0.00476
R9214 DVDD.n2116 DVDD.n2079 0.00476
R9215 DVDD.n2116 DVDD.n2115 0.00476
R9216 DVDD.n2115 DVDD.n2114 0.00476
R9217 DVDD.n2114 DVDD.n2085 0.00476
R9218 DVDD.n2110 DVDD.n2085 0.00476
R9219 DVDD.n2110 DVDD.n2109 0.00476
R9220 DVDD.n2109 DVDD.n2108 0.00476
R9221 DVDD.n2108 DVDD.n2091 0.00476
R9222 DVDD.n2104 DVDD.n2091 0.00476
R9223 DVDD.n2104 DVDD.n2103 0.00476
R9224 DVDD.n2103 DVDD.n2102 0.00476
R9225 DVDD.n2102 DVDD.n2097 0.00476
R9226 DVDD.n2276 DVDD.n1327 0.00476
R9227 DVDD.n2272 DVDD.n1327 0.00476
R9228 DVDD.n2272 DVDD.n2271 0.00476
R9229 DVDD.n2271 DVDD.n2270 0.00476
R9230 DVDD.n2270 DVDD.n2246 0.00476
R9231 DVDD.n2266 DVDD.n2246 0.00476
R9232 DVDD.n2266 DVDD.n2265 0.00476
R9233 DVDD.n2265 DVDD.n2264 0.00476
R9234 DVDD.n2264 DVDD.n2252 0.00476
R9235 DVDD.n2260 DVDD.n2252 0.00476
R9236 DVDD.n1843 DVDD.n1842 0.00476
R9237 DVDD.n1842 DVDD.n1841 0.00476
R9238 DVDD.n1841 DVDD.n1799 0.00476
R9239 DVDD.n1837 DVDD.n1799 0.00476
R9240 DVDD.n1837 DVDD.n1836 0.00476
R9241 DVDD.n1836 DVDD.n1835 0.00476
R9242 DVDD.n1835 DVDD.n1805 0.00476
R9243 DVDD.n1831 DVDD.n1805 0.00476
R9244 DVDD.n1831 DVDD.n1830 0.00476
R9245 DVDD.n1830 DVDD.n1829 0.00476
R9246 DVDD.n1829 DVDD.n1811 0.00476
R9247 DVDD.n1825 DVDD.n1811 0.00476
R9248 DVDD.n1825 DVDD.n1824 0.00476
R9249 DVDD.n1824 DVDD.n1823 0.00476
R9250 DVDD.n1823 DVDD.n1717 0.00476
R9251 DVDD.n2024 DVDD.n1744 0.00476
R9252 DVDD.n2020 DVDD.n1744 0.00476
R9253 DVDD.n2020 DVDD.n2019 0.00476
R9254 DVDD.n2019 DVDD.n2018 0.00476
R9255 DVDD.n2014 DVDD.n2013 0.00476
R9256 DVDD.n2013 DVDD.n2012 0.00476
R9257 DVDD.n2012 DVDD.n1948 0.00476
R9258 DVDD.n2008 DVDD.n1948 0.00476
R9259 DVDD.n2008 DVDD.n2007 0.00476
R9260 DVDD.n2007 DVDD.n2006 0.00476
R9261 DVDD.n2006 DVDD.n1954 0.00476
R9262 DVDD.n2002 DVDD.n1954 0.00476
R9263 DVDD.n2002 DVDD.n2001 0.00476
R9264 DVDD.n2001 DVDD.n314 0.00476
R9265 DVDD.n1994 DVDD.n1993 0.00476
R9266 DVDD.n1993 DVDD.n1992 0.00476
R9267 DVDD.n1992 DVDD.n1965 0.00476
R9268 DVDD.n1988 DVDD.n1965 0.00476
R9269 DVDD.n1988 DVDD.n1987 0.00476
R9270 DVDD.n1987 DVDD.n1986 0.00476
R9271 DVDD.n1986 DVDD.n1971 0.00476
R9272 DVDD.n1982 DVDD.n1971 0.00476
R9273 DVDD.n1982 DVDD.n1981 0.00476
R9274 DVDD.n1981 DVDD.n1980 0.00476
R9275 DVDD.n2055 DVDD.n2054 0.00476
R9276 DVDD.n2054 DVDD.n2053 0.00476
R9277 DVDD.n2053 DVDD.n1587 0.00476
R9278 DVDD.n2049 DVDD.n1587 0.00476
R9279 DVDD.n1697 DVDD.n1608 0.00476
R9280 DVDD.n1693 DVDD.n1608 0.00476
R9281 DVDD.n1693 DVDD.n1692 0.00476
R9282 DVDD.n1692 DVDD.n1691 0.00476
R9283 DVDD.n1691 DVDD.n1614 0.00476
R9284 DVDD.n1687 DVDD.n1614 0.00476
R9285 DVDD.n1687 DVDD.n1686 0.00476
R9286 DVDD.n1686 DVDD.n1685 0.00476
R9287 DVDD.n1685 DVDD.n1620 0.00476
R9288 DVDD.n1681 DVDD.n1620 0.00476
R9289 DVDD.n1681 DVDD.n1680 0.00476
R9290 DVDD.n1680 DVDD.n1679 0.00476
R9291 DVDD.n1679 DVDD.n1626 0.00476
R9292 DVDD.n1675 DVDD.n1626 0.00476
R9293 DVDD.n1675 DVDD.n1674 0.00476
R9294 DVDD.n1668 DVDD.n1667 0.00476
R9295 DVDD.n1667 DVDD.n1666 0.00476
R9296 DVDD.n1666 DVDD.n1636 0.00476
R9297 DVDD.n1662 DVDD.n1636 0.00476
R9298 DVDD.n1662 DVDD.n1661 0.00476
R9299 DVDD.n1661 DVDD.n1660 0.00476
R9300 DVDD.n1660 DVDD.n1642 0.00476
R9301 DVDD.n1656 DVDD.n1642 0.00476
R9302 DVDD.n1656 DVDD.n1655 0.00476
R9303 DVDD.n1655 DVDD.n1654 0.00476
R9304 DVDD.n2978 DVDD.n785 0.00476
R9305 DVDD.n2982 DVDD.n785 0.00476
R9306 DVDD.n2982 DVDD.n773 0.00476
R9307 DVDD.n2986 DVDD.n773 0.00476
R9308 DVDD.n2986 DVDD.n771 0.00476
R9309 DVDD.n2990 DVDD.n771 0.00476
R9310 DVDD.n2990 DVDD.n769 0.00476
R9311 DVDD.n2994 DVDD.n769 0.00476
R9312 DVDD.n2994 DVDD.n767 0.00476
R9313 DVDD.n2998 DVDD.n767 0.00476
R9314 DVDD.n2998 DVDD.n765 0.00476
R9315 DVDD.n3002 DVDD.n765 0.00476
R9316 DVDD.n3002 DVDD.n763 0.00476
R9317 DVDD.n3007 DVDD.n763 0.00476
R9318 DVDD.n3007 DVDD.n761 0.00476
R9319 DVDD.n3011 DVDD.n761 0.00476
R9320 DVDD.n3012 DVDD.n3011 0.00476
R9321 DVDD.n3012 DVDD.n759 0.00476
R9322 DVDD.n3026 DVDD.n759 0.00476
R9323 DVDD.n3026 DVDD.n3025 0.00476
R9324 DVDD.n3025 DVDD.n3024 0.00476
R9325 DVDD.n3024 DVDD.n3019 0.00476
R9326 DVDD.n3020 DVDD.n3019 0.00476
R9327 DVDD.n4962 DVDD.n4959 0.00476
R9328 DVDD.n4962 DVDD.n4958 0.00476
R9329 DVDD.n4966 DVDD.n4958 0.00476
R9330 DVDD.n4966 DVDD.n4956 0.00476
R9331 DVDD.n4970 DVDD.n4956 0.00476
R9332 DVDD.n4970 DVDD.n4954 0.00476
R9333 DVDD.n4974 DVDD.n4954 0.00476
R9334 DVDD.n4974 DVDD.n4952 0.00476
R9335 DVDD.n4978 DVDD.n4952 0.00476
R9336 DVDD.n4978 DVDD.n4950 0.00476
R9337 DVDD.n5244 DVDD.n4950 0.00476
R9338 DVDD.n5244 DVDD.n5243 0.00476
R9339 DVDD.n5243 DVDD.n5241 0.00476
R9340 DVDD.n5241 DVDD.n4984 0.00476
R9341 DVDD.n5237 DVDD.n4984 0.00476
R9342 DVDD.n5237 DVDD.n5236 0.00476
R9343 DVDD.n5236 DVDD.n5235 0.00476
R9344 DVDD.n5235 DVDD.n4990 0.00476
R9345 DVDD.n5231 DVDD.n4990 0.00476
R9346 DVDD.n5231 DVDD.n5230 0.00476
R9347 DVDD.n5230 DVDD.n5229 0.00476
R9348 DVDD.n5229 DVDD.n4996 0.00476
R9349 DVDD.n5225 DVDD.n4996 0.00476
R9350 DVDD.n5223 DVDD.n5072 0.00476
R9351 DVDD.n5219 DVDD.n5072 0.00476
R9352 DVDD.n5219 DVDD.n5218 0.00476
R9353 DVDD.n5218 DVDD.n5217 0.00476
R9354 DVDD.n5217 DVDD.n5078 0.00476
R9355 DVDD.n5200 DVDD.n5078 0.00476
R9356 DVDD.n5200 DVDD.n5199 0.00476
R9357 DVDD.n5199 DVDD.n5198 0.00476
R9358 DVDD.n5198 DVDD.n5160 0.00476
R9359 DVDD.n5194 DVDD.n5160 0.00476
R9360 DVDD.n5194 DVDD.n5193 0.00476
R9361 DVDD.n5193 DVDD.n5192 0.00476
R9362 DVDD.n5192 DVDD.n5166 0.00476
R9363 DVDD.n5188 DVDD.n5166 0.00476
R9364 DVDD.n5188 DVDD.n5187 0.00476
R9365 DVDD.n5187 DVDD.n5186 0.00476
R9366 DVDD.n5186 DVDD.n5172 0.00476
R9367 DVDD.n5182 DVDD.n5172 0.00476
R9368 DVDD.n5182 DVDD.n5181 0.00476
R9369 DVDD.n5181 DVDD.n5180 0.00476
R9370 DVDD.n5180 DVDD.n697 0.00476
R9371 DVDD.n5393 DVDD.n697 0.00476
R9372 DVDD.n5394 DVDD.n5393 0.00476
R9373 DVDD.n5429 DVDD.n661 0.00476
R9374 DVDD.n5425 DVDD.n661 0.00476
R9375 DVDD.n5425 DVDD.n5424 0.00476
R9376 DVDD.n5424 DVDD.n5423 0.00476
R9377 DVDD.n5423 DVDD.n5401 0.00476
R9378 DVDD.n5419 DVDD.n5401 0.00476
R9379 DVDD.n5419 DVDD.n5418 0.00476
R9380 DVDD.n5418 DVDD.n5417 0.00476
R9381 DVDD.n5417 DVDD.n5407 0.00476
R9382 DVDD.n5413 DVDD.n5407 0.00476
R9383 DVDD.n2984 DVDD.n2983 0.00476
R9384 DVDD.n2985 DVDD.n2984 0.00476
R9385 DVDD.n2985 DVDD.n770 0.00476
R9386 DVDD.n2991 DVDD.n770 0.00476
R9387 DVDD.n2992 DVDD.n2991 0.00476
R9388 DVDD.n2993 DVDD.n2992 0.00476
R9389 DVDD.n2993 DVDD.n766 0.00476
R9390 DVDD.n2999 DVDD.n766 0.00476
R9391 DVDD.n3000 DVDD.n2999 0.00476
R9392 DVDD.n3001 DVDD.n3000 0.00476
R9393 DVDD.n3001 DVDD.n762 0.00476
R9394 DVDD.n3008 DVDD.n762 0.00476
R9395 DVDD.n3009 DVDD.n3008 0.00476
R9396 DVDD.n3010 DVDD.n3009 0.00476
R9397 DVDD.n3010 DVDD.n745 0.00476
R9398 DVDD.n3027 DVDD.n758 0.00476
R9399 DVDD.n3023 DVDD.n758 0.00476
R9400 DVDD.n3023 DVDD.n3022 0.00476
R9401 DVDD.n3022 DVDD.n3021 0.00476
R9402 DVDD.n4961 DVDD.n4960 0.00476
R9403 DVDD.n4961 DVDD.n4957 0.00476
R9404 DVDD.n4967 DVDD.n4957 0.00476
R9405 DVDD.n4968 DVDD.n4967 0.00476
R9406 DVDD.n4969 DVDD.n4968 0.00476
R9407 DVDD.n4969 DVDD.n4953 0.00476
R9408 DVDD.n4975 DVDD.n4953 0.00476
R9409 DVDD.n4976 DVDD.n4975 0.00476
R9410 DVDD.n4977 DVDD.n4976 0.00476
R9411 DVDD.n4977 DVDD.n4938 0.00476
R9412 DVDD.n5240 DVDD.n5239 0.00476
R9413 DVDD.n5239 DVDD.n5238 0.00476
R9414 DVDD.n5238 DVDD.n4985 0.00476
R9415 DVDD.n5234 DVDD.n4985 0.00476
R9416 DVDD.n5234 DVDD.n5233 0.00476
R9417 DVDD.n5233 DVDD.n5232 0.00476
R9418 DVDD.n5232 DVDD.n4991 0.00476
R9419 DVDD.n5228 DVDD.n4991 0.00476
R9420 DVDD.n5228 DVDD.n5227 0.00476
R9421 DVDD.n5227 DVDD.n5226 0.00476
R9422 DVDD.n5222 DVDD.n5221 0.00476
R9423 DVDD.n5221 DVDD.n5220 0.00476
R9424 DVDD.n5220 DVDD.n5073 0.00476
R9425 DVDD.n5216 DVDD.n5073 0.00476
R9426 DVDD.n5201 DVDD.n5155 0.00476
R9427 DVDD.n5197 DVDD.n5155 0.00476
R9428 DVDD.n5197 DVDD.n5196 0.00476
R9429 DVDD.n5196 DVDD.n5195 0.00476
R9430 DVDD.n5195 DVDD.n5161 0.00476
R9431 DVDD.n5191 DVDD.n5161 0.00476
R9432 DVDD.n5191 DVDD.n5190 0.00476
R9433 DVDD.n5190 DVDD.n5189 0.00476
R9434 DVDD.n5189 DVDD.n5167 0.00476
R9435 DVDD.n5185 DVDD.n5167 0.00476
R9436 DVDD.n5185 DVDD.n5184 0.00476
R9437 DVDD.n5184 DVDD.n5183 0.00476
R9438 DVDD.n5183 DVDD.n5173 0.00476
R9439 DVDD.n5179 DVDD.n5173 0.00476
R9440 DVDD.n5179 DVDD.n699 0.00476
R9441 DVDD.n5428 DVDD.n5427 0.00476
R9442 DVDD.n5427 DVDD.n5426 0.00476
R9443 DVDD.n5426 DVDD.n5397 0.00476
R9444 DVDD.n5422 DVDD.n5397 0.00476
R9445 DVDD.n5422 DVDD.n5421 0.00476
R9446 DVDD.n5421 DVDD.n5420 0.00476
R9447 DVDD.n5420 DVDD.n5402 0.00476
R9448 DVDD.n5416 DVDD.n5402 0.00476
R9449 DVDD.n5416 DVDD.n5415 0.00476
R9450 DVDD.n5415 DVDD.n5414 0.00476
R9451 DVDD.n3500 DVDD.n3499 0.00476
R9452 DVDD.n3499 DVDD.n3489 0.00476
R9453 DVDD.n3489 DVDD.n3244 0.00476
R9454 DVDD.n4860 DVDD.n3245 0.00476
R9455 DVDD.n4853 DVDD.n3245 0.00476
R9456 DVDD.n4853 DVDD.n4852 0.00476
R9457 DVDD.n4852 DVDD.n3253 0.00476
R9458 DVDD.n4807 DVDD.n4791 0.00476
R9459 DVDD.n4807 DVDD.n4806 0.00476
R9460 DVDD.n4806 DVDD.n4798 0.00476
R9461 DVDD.n4798 DVDD.n190 0.00476
R9462 DVDD.n3124 DVDD.n189 0.00476
R9463 DVDD.n3124 DVDD.n3123 0.00476
R9464 DVDD.n3123 DVDD.n3086 0.00476
R9465 DVDD.n3115 DVDD.n3086 0.00476
R9466 DVDD.n3114 DVDD.n3113 0.00476
R9467 DVDD.n3113 DVDD.n3095 0.00476
R9468 DVDD.n3105 DVDD.n3095 0.00476
R9469 DVDD.n3105 DVDD.n3104 0.00476
R9470 DVDD.n5727 DVDD.n231 0.00476
R9471 DVDD.n5720 DVDD.n231 0.00476
R9472 DVDD.n5720 DVDD.n5719 0.00476
R9473 DVDD.n4512 DVDD.n4508 0.00476
R9474 DVDD.n4512 DVDD.n4509 0.00476
R9475 DVDD.n4509 DVDD.n3243 0.00476
R9476 DVDD.n4868 DVDD.n3151 0.00476
R9477 DVDD.n4868 DVDD.n3152 0.00476
R9478 DVDD.n3152 DVDD.n3138 0.00476
R9479 DVDD.n4886 DVDD.n3138 0.00476
R9480 DVDD.n4887 DVDD.n3135 0.00476
R9481 DVDD.n4893 DVDD.n3135 0.00476
R9482 DVDD.n4893 DVDD.n3136 0.00476
R9483 DVDD.n3136 DVDD.n199 0.00476
R9484 DVDD.n5090 DVDD.n198 0.00476
R9485 DVDD.n5101 DVDD.n5090 0.00476
R9486 DVDD.n5101 DVDD.n5092 0.00476
R9487 DVDD.n5097 DVDD.n5092 0.00476
R9488 DVDD.n5114 DVDD.n5085 0.00476
R9489 DVDD.n5114 DVDD.n5081 0.00476
R9490 DVDD.n5118 DVDD.n5081 0.00476
R9491 DVDD.n5118 DVDD.n5083 0.00476
R9492 DVDD.n5132 DVDD.n5129 0.00476
R9493 DVDD.n5132 DVDD.n5127 0.00476
R9494 DVDD.n5136 DVDD.n5127 0.00476
R9495 DVDD.n4696 DVDD.n3369 0.00476
R9496 DVDD.n4700 DVDD.n3369 0.00476
R9497 DVDD.n4700 DVDD.n3173 0.00476
R9498 DVDD.n4709 DVDD.n3172 0.00476
R9499 DVDD.n4712 DVDD.n4709 0.00476
R9500 DVDD.n4712 DVDD.n3362 0.00476
R9501 DVDD.n4720 DVDD.n3362 0.00476
R9502 DVDD.n4735 DVDD.n3359 0.00476
R9503 DVDD.n4735 DVDD.n3360 0.00476
R9504 DVDD.n4731 DVDD.n3360 0.00476
R9505 DVDD.n4731 DVDD.n201 0.00476
R9506 DVDD.n5744 DVDD.n203 0.00476
R9507 DVDD.n5740 DVDD.n203 0.00476
R9508 DVDD.n5740 DVDD.n5739 0.00476
R9509 DVDD.n5739 DVDD.n5738 0.00476
R9510 DVDD.n5734 DVDD.n208 0.00476
R9511 DVDD.n5734 DVDD.n5733 0.00476
R9512 DVDD.n5733 DVDD.n5732 0.00476
R9513 DVDD.n5732 DVDD.n213 0.00476
R9514 DVDD.n3050 DVDD.n738 0.00476
R9515 DVDD.n3050 DVDD.n739 0.00476
R9516 DVDD.n3046 DVDD.n739 0.00476
R9517 DVDD.n3190 DVDD.n3180 0.00476
R9518 DVDD.n3194 DVDD.n3180 0.00476
R9519 DVDD.n3194 DVDD.n3175 0.00476
R9520 DVDD.n3242 DVDD.n3176 0.00476
R9521 DVDD.n3235 DVDD.n3176 0.00476
R9522 DVDD.n3235 DVDD.n3234 0.00476
R9523 DVDD.n3234 DVDD.n3205 0.00476
R9524 DVDD.n3227 DVDD.n3226 0.00476
R9525 DVDD.n3226 DVDD.n3210 0.00476
R9526 DVDD.n3219 DVDD.n3210 0.00476
R9527 DVDD.n3219 DVDD.n193 0.00476
R9528 DVDD.n722 DVDD.n192 0.00476
R9529 DVDD.n5330 DVDD.n722 0.00476
R9530 DVDD.n5330 DVDD.n719 0.00476
R9531 DVDD.n5334 DVDD.n719 0.00476
R9532 DVDD.n5343 DVDD.n711 0.00476
R9533 DVDD.n5343 DVDD.n709 0.00476
R9534 DVDD.n5347 DVDD.n709 0.00476
R9535 DVDD.n5348 DVDD.n5347 0.00476
R9536 DVDD.n5353 DVDD.n704 0.00476
R9537 DVDD.n5362 DVDD.n704 0.00476
R9538 DVDD.n5362 DVDD.n702 0.00476
R9539 DVDD.n5458 DVDD.n5457 0.0047
R9540 DVDD.n2563 DVDD.n444 0.00469776
R9541 DVDD.n5070 DVDD.n5069 0.004625
R9542 DVDD.n5434 DVDD.n604 0.00460625
R9543 DVDD.n2975 DVDD.n2974 0.00460625
R9544 DVDD.n5635 DVDD.n413 0.00455
R9545 DVDD.n5642 DVDD.n383 0.00455
R9546 DVDD.n5646 DVDD.n362 0.00455
R9547 DVDD.n2049 DVDD.n2048 0.00455
R9548 DVDD.n5216 DVDD.n5215 0.00455
R9549 DVDD.n2554 DVDD.n992 0.00455
R9550 DVDD.n3857 DVDD.n3576 0.00455
R9551 DVDD.n2555 DVDD.n439 0.00455
R9552 DVDD.n3932 DVDD.n3658 0.00455
R9553 DVDD.n2548 DVDD.n975 0.00455
R9554 DVDD.n2550 DVDD.n458 0.00455
R9555 DVDD.n1945 DVDD.n1944 0.0045
R9556 DVDD.n1976 DVDD.n1289 0.0045
R9557 DVDD.n1853 DVDD.n1849 0.0045
R9558 DVDD.n1944 DVDD.n1943 0.0045
R9559 DVDD.n1853 DVDD.n1773 0.0045
R9560 DVDD.n1943 DVDD.n1942 0.0045
R9561 DVDD.n1367 DVDD.n1330 0.0045
R9562 DVDD.n2351 DVDD.n1289 0.0045
R9563 DVDD.n2351 DVDD.n2350 0.0045
R9564 DVDD.n2241 DVDD.n1329 0.0045
R9565 DVDD.n2241 DVDD.n1367 0.0045
R9566 DVDD.n1849 DVDD.n1848 0.0045
R9567 DVDD.n2949 DVDD.n972 0.00443
R9568 DVDD.n2956 DVDD.n940 0.00443
R9569 DVDD.n2179 DVDD.n1446 0.00443
R9570 DVDD.n2034 DVDD.n2024 0.00443
R9571 DVDD.n3037 DVDD.n3027 0.00443
R9572 DVDD.n676 DVDD.n675 0.0044
R9573 DVDD.n657 DVDD.n604 0.00438125
R9574 DVDD.n2974 DVDD.n2973 0.00438125
R9575 DVDD.n1537 DVDD.n1536 0.00436194
R9576 DVDD.n1235 DVDD.n1234 0.00436194
R9577 DVDD.n5690 DVDD.n5689 0.004325
R9578 DVDD.n2152 DVDD.n1564 0.00422
R9579 DVDD.n5278 DVDD.n4937 0.00422
R9580 DVDD.n4507 DVDD.n4504 0.00422
R9581 DVDD.n4884 DVDD.n3139 0.00422
R9582 DVDD.n5756 DVDD.n177 0.00422
R9583 DVDD.n5103 DVDD.n4912 0.00422
R9584 DVDD.n5112 DVDD.n5111 0.00422
R9585 DVDD.n4934 DVDD.n4933 0.00422
R9586 DVDD.n4694 DVDD.n3372 0.00422
R9587 DVDD.n4718 DVDD.n4717 0.00422
R9588 DVDD.n4738 DVDD.n4737 0.00422
R9589 DVDD.n3071 DVDD.n3070 0.00422
R9590 DVDD.n3062 DVDD.n3061 0.00422
R9591 DVDD.n3044 DVDD.n740 0.00422
R9592 DVDD.n3490 DVDD.n3486 0.00422
R9593 DVDD.n4850 DVDD.n3254 0.00422
R9594 DVDD.n4810 DVDD.n4809 0.00422
R9595 DVDD.n3121 DVDD.n3087 0.00422
R9596 DVDD.n3111 DVDD.n3097 0.00422
R9597 DVDD.n5717 DVDD.n240 0.00422
R9598 DVDD.n3188 DVDD.n3183 0.00422
R9599 DVDD.n3232 DVDD.n3230 0.00422
R9600 DVDD.n3211 DVDD.n3206 0.00422
R9601 DVDD.n5328 DVDD.n724 0.00422
R9602 DVDD.n5341 DVDD.n715 0.00422
R9603 DVDD.n5365 DVDD.n701 0.00422
R9604 DVDD.n4875 DVDD.n4874 0.00413
R9605 DVDD.n3134 DVDD.n3133 0.00413
R9606 DVDD.n5138 DVDD.n5137 0.00413
R9607 DVDD.n4714 DVDD.n3363 0.00413
R9608 DVDD.n4736 DVDD.n3358 0.00413
R9609 DVDD.n3045 DVDD.n742 0.00413
R9610 DVDD.n4851 DVDD.n3249 0.00413
R9611 DVDD.n4808 DVDD.n4790 0.00413
R9612 DVDD.n5718 DVDD.n237 0.00413
R9613 DVDD.n3233 DVDD.n3201 0.00413
R9614 DVDD.n3225 DVDD.n3224 0.00413
R9615 DVDD.n5360 DVDD.n706 0.00413
R9616 DVDD DVDD.n729 0.00408591
R9617 DVDD.n4536 DVDD.n3430 0.00407
R9618 DVDD.n5091 DVDD.n4913 0.00407
R9619 DVDD.n5113 DVDD.n4914 0.00407
R9620 DVDD.n4695 DVDD.n3370 0.00407
R9621 DVDD.n3067 DVDD.n206 0.00407
R9622 DVDD.n3065 DVDD.n210 0.00407
R9623 DVDD.n3502 DVDD.n3501 0.00407
R9624 DVDD.n3117 DVDD.n3089 0.00407
R9625 DVDD.n3112 DVDD.n3096 0.00407
R9626 DVDD.n3189 DVDD.n3181 0.00407
R9627 DVDD.n5336 DVDD.n717 0.00407
R9628 DVDD.n5342 DVDD.n712 0.00407
R9629 DVDD.n1670 DVDD.n1669 0.00404
R9630 DVDD.n2275 DVDD.n1328 0.00404
R9631 DVDD.n1365 DVDD.n1321 0.00404
R9632 DVDD.n2314 DVDD.n2313 0.00404
R9633 DVDD.n2312 DVDD.n2279 0.00404
R9634 DVDD.n2278 DVDD.n1324 0.00404
R9635 DVDD.n2277 DVDD.n2276 0.00404
R9636 DVDD.n1668 DVDD.n1325 0.00404
R9637 DVDD.n5429 DVDD.n656 0.00404
R9638 DVDD.n5428 DVDD.n5396 0.00404
R9639 DVDD.n2914 DVDD.n2589 0.00403571
R9640 DVDD.n3745 DVDD.n3700 0.00403571
R9641 DVDD.n4325 DVDD.n3483 0.00403571
R9642 DVDD.n790 DVDD.n786 0.004025
R9643 DVDD.n2564 DVDD.n1018 0.00401
R9644 DVDD.n5633 DVDD.n420 0.00401
R9645 DVDD.n2369 DVDD.n1222 0.00401
R9646 DVDD.n5639 DVDD.n388 0.00401
R9647 DVDD.n2151 DVDD.n1548 0.00401
R9648 DVDD.n2078 DVDD.n368 0.00401
R9649 DVDD.n1996 DVDD.n312 0.00401
R9650 DVDD.n1709 DVDD.n1599 0.00401
R9651 DVDD.n5242 DVDD.n4936 0.00401
R9652 DVDD.n5212 DVDD.n5143 0.00401
R9653 DVDD.n1653 DVDD 0.00392
R9654 DVDD.n2261 DVDD 0.00392
R9655 DVDD DVDD.n1345 0.00392
R9656 DVDD.n2297 DVDD 0.00392
R9657 DVDD.n2298 DVDD 0.00392
R9658 DVDD.n1350 DVDD 0.00392
R9659 DVDD.n2260 DVDD 0.00392
R9660 DVDD.n1654 DVDD 0.00392
R9661 DVDD.n5413 DVDD 0.00392
R9662 DVDD.n5414 DVDD 0.00392
R9663 DVDD.n2952 DVDD.n959 0.00389
R9664 DVDD.n1922 DVDD.n1016 0.00389
R9665 DVDD.n2959 DVDD.n927 0.00389
R9666 DVDD.n2374 DVDD.n1189 0.00389
R9667 DVDD.n2963 DVDD.n907 0.00389
R9668 DVDD.n2154 DVDD.n1481 0.00389
R9669 DVDD.n2037 DVDD.n1723 0.00389
R9670 DVDD.n5654 DVDD.n326 0.00389
R9671 DVDD.n3040 DVDD.n746 0.00389
R9672 DVDD.n5281 DVDD.n5245 0.00389
R9673 DVDD.n4514 DVDD.n4513 0.00383
R9674 DVDD.n5102 DVDD.n5088 0.00383
R9675 DVDD.n5120 DVDD.n5080 0.00383
R9676 DVDD.n3371 DVDD.n3368 0.00383
R9677 DVDD.n3074 DVDD.n205 0.00383
R9678 DVDD.n3058 DVDD.n211 0.00383
R9679 DVDD.n3498 DVDD.n3497 0.00383
R9680 DVDD.n3122 DVDD.n3082 0.00383
R9681 DVDD.n3107 DVDD.n3099 0.00383
R9682 DVDD.n3182 DVDD.n3179 0.00383
R9683 DVDD.n5329 DVDD.n723 0.00383
R9684 DVDD.n714 DVDD.n713 0.00383
R9685 DVDD.n2057 DVDD.n2056 0.0038
R9686 DVDD.n2132 DVDD.n2131 0.0038
R9687 DVDD.n2490 DVDD.n1065 0.0038
R9688 DVDD.n2348 DVDD.n1060 0.0038
R9689 DVDD.n2493 DVDD.n1061 0.0038
R9690 DVDD.n2492 DVDD.n2491 0.0038
R9691 DVDD.n2130 DVDD.n1062 0.0038
R9692 DVDD.n2055 DVDD.n1586 0.0038
R9693 DVDD.n5224 DVDD.n5223 0.0038
R9694 DVDD.n5222 DVDD.n4997 0.0038
R9695 DVDD.n2927 DVDD.n2575 0.00377857
R9696 DVDD.n4112 DVDD.n3552 0.00377857
R9697 DVDD.n5987 DVDD.n17 0.00377857
R9698 DVDD.n233 DVDD 0.00376574
R9699 DVDD DVDD.n230 0.00376574
R9700 DVDD DVDD.n3169 0.00376574
R9701 DVDD.n4861 DVDD 0.00376574
R9702 DVDD.n5507 DVDD.n331 0.0036903
R9703 DVDD.n2569 DVDD.n518 0.0036903
R9704 DVDD.n5452 DVDD.n645 0.00365
R9705 DVDD.n5453 DVDD.n646 0.00365
R9706 DVDD.n2233 DVDD.n2232 0.00365
R9707 DVDD.n2449 DVDD.n1117 0.00365
R9708 DVDD.n2521 DVDD.n2519 0.00365
R9709 DVDD.n3858 DVDD.n3585 0.00365
R9710 DVDD.n5645 DVDD.n5644 0.00365
R9711 DVDD.n1118 DVDD.n397 0.00365
R9712 DVDD.n2522 DVDD.n422 0.00365
R9713 DVDD.n3931 DVDD.n3657 0.00365
R9714 DVDD.n2962 DVDD.n2961 0.00365
R9715 DVDD.n1120 DVDD.n936 0.00365
R9716 DVDD.n2513 DVDD.n961 0.00365
R9717 DVDD.n2219 DVDD.n2218 0.00365
R9718 DVDD.n2443 DVDD.n1121 0.00365
R9719 DVDD.n2516 DVDD.n2514 0.00365
R9720 DVDD.n2973 DVDD.n2972 0.00359375
R9721 DVDD.n4870 DVDD.n3148 0.00359
R9722 DVDD.n4895 DVDD.n4894 0.00359
R9723 DVDD.n5130 DVDD.n5126 0.00359
R9724 DVDD.n4713 DVDD.n3365 0.00359
R9725 DVDD.n4725 DVDD.n4724 0.00359
R9726 DVDD.n741 DVDD.n737 0.00359
R9727 DVDD.n4855 DVDD.n4854 0.00359
R9728 DVDD.n4805 DVDD.n4804 0.00359
R9729 DVDD.n5722 DVDD.n5721 0.00359
R9730 DVDD.n3237 DVDD.n3236 0.00359
R9731 DVDD.n3221 DVDD.n3212 0.00359
R9732 DVDD.n5361 DVDD.n705 0.00359
R9733 DVDD.n2016 DVDD.n2015 0.00356
R9734 DVDD.n2170 DVDD.n1173 0.00356
R9735 DVDD.n2393 DVDD.n2392 0.00356
R9736 DVDD.n1940 DVDD.n1172 0.00356
R9737 DVDD.n1939 DVDD.n1906 0.00356
R9738 DVDD.n2391 DVDD.n1176 0.00356
R9739 DVDD.n2172 DVDD.n2171 0.00356
R9740 DVDD.n2014 DVDD.n1452 0.00356
R9741 DVDD.n4959 DVDD.n285 0.00356
R9742 DVDD.n4960 DVDD.n287 0.00356
R9743 DVDD.n307 DVDD.n306 0.003425
R9744 DVDD.n4505 DVDD.n4498 0.003425
R9745 DVDD.n4910 DVDD.n4909 0.003425
R9746 DVDD.n5109 DVDD.n4918 0.003425
R9747 DVDD.n5434 DVDD.n605 0.00336875
R9748 DVDD.n2941 DVDD.n979 0.00335448
R9749 DVDD.n1861 DVDD.n1860 0.00334
R9750 DVDD.n1862 DVDD.n1861 0.00334
R9751 DVDD.n1862 DVDD.n1771 0.00334
R9752 DVDD.n1868 DVDD.n1771 0.00334
R9753 DVDD.n1869 DVDD.n1868 0.00334
R9754 DVDD.n1870 DVDD.n1869 0.00334
R9755 DVDD.n1870 DVDD.n1767 0.00334
R9756 DVDD.n1876 DVDD.n1767 0.00334
R9757 DVDD.n1877 DVDD.n1876 0.00334
R9758 DVDD.n1878 DVDD.n1877 0.00334
R9759 DVDD.n1878 DVDD.n1763 0.00334
R9760 DVDD.n1884 DVDD.n1763 0.00334
R9761 DVDD.n1885 DVDD.n1884 0.00334
R9762 DVDD.n1886 DVDD.n1885 0.00334
R9763 DVDD.n1886 DVDD.n1759 0.00334
R9764 DVDD.n1892 DVDD.n1759 0.00334
R9765 DVDD.n1893 DVDD.n1892 0.00334
R9766 DVDD.n1894 DVDD.n1893 0.00334
R9767 DVDD.n1894 DVDD.n1757 0.00334
R9768 DVDD.n1900 DVDD.n1757 0.00334
R9769 DVDD.n1901 DVDD.n1900 0.00334
R9770 DVDD.n1902 DVDD.n1901 0.00334
R9771 DVDD.n1902 DVDD.n1752 0.00334
R9772 DVDD.n1941 DVDD.n1753 0.00334
R9773 DVDD.n1908 DVDD.n1753 0.00334
R9774 DVDD.n1909 DVDD.n1908 0.00334
R9775 DVDD.n1910 DVDD.n1909 0.00334
R9776 DVDD.n1913 DVDD.n1910 0.00334
R9777 DVDD.n1914 DVDD.n1913 0.00334
R9778 DVDD.n1915 DVDD.n1914 0.00334
R9779 DVDD.n1916 DVDD.n1915 0.00334
R9780 DVDD.n1918 DVDD.n1916 0.00334
R9781 DVDD.n1919 DVDD.n1918 0.00334
R9782 DVDD.n1921 DVDD.n1919 0.00334
R9783 DVDD.n1921 DVDD.n1920 0.00334
R9784 DVDD.n1920 DVDD.n1045 0.00334
R9785 DVDD.n1046 DVDD.n1045 0.00334
R9786 DVDD.n1047 DVDD.n1046 0.00334
R9787 DVDD.n1050 DVDD.n1047 0.00334
R9788 DVDD.n1051 DVDD.n1050 0.00334
R9789 DVDD.n1052 DVDD.n1051 0.00334
R9790 DVDD.n1053 DVDD.n1052 0.00334
R9791 DVDD.n1056 DVDD.n1053 0.00334
R9792 DVDD.n1057 DVDD.n1056 0.00334
R9793 DVDD.n1058 DVDD.n1057 0.00334
R9794 DVDD.n1059 DVDD.n1058 0.00334
R9795 DVDD.n2349 DVDD.n1290 0.00334
R9796 DVDD.n1292 DVDD.n1290 0.00334
R9797 DVDD.n1293 DVDD.n1292 0.00334
R9798 DVDD.n1294 DVDD.n1293 0.00334
R9799 DVDD.n1295 DVDD.n1294 0.00334
R9800 DVDD.n1296 DVDD.n1295 0.00334
R9801 DVDD.n1297 DVDD.n1296 0.00334
R9802 DVDD.n1300 DVDD.n1297 0.00334
R9803 DVDD.n1301 DVDD.n1300 0.00334
R9804 DVDD.n1302 DVDD.n1301 0.00334
R9805 DVDD.n1303 DVDD.n1302 0.00334
R9806 DVDD.n1306 DVDD.n1303 0.00334
R9807 DVDD.n1307 DVDD.n1306 0.00334
R9808 DVDD.n1308 DVDD.n1307 0.00334
R9809 DVDD.n1309 DVDD.n1308 0.00334
R9810 DVDD.n1312 DVDD.n1309 0.00334
R9811 DVDD.n1313 DVDD.n1312 0.00334
R9812 DVDD.n1314 DVDD.n1313 0.00334
R9813 DVDD.n1315 DVDD.n1314 0.00334
R9814 DVDD.n1317 DVDD.n1315 0.00334
R9815 DVDD.n1318 DVDD.n1317 0.00334
R9816 DVDD.n1319 DVDD.n1318 0.00334
R9817 DVDD.n1320 DVDD.n1319 0.00334
R9818 DVDD.n2281 DVDD.n1322 0.00334
R9819 DVDD.n2282 DVDD.n2281 0.00334
R9820 DVDD.n2283 DVDD.n2282 0.00334
R9821 DVDD.n2284 DVDD.n2283 0.00334
R9822 DVDD.n2287 DVDD.n2284 0.00334
R9823 DVDD.n2288 DVDD.n2287 0.00334
R9824 DVDD.n2289 DVDD.n2288 0.00334
R9825 DVDD.n2290 DVDD.n2289 0.00334
R9826 DVDD.n2292 DVDD.n2290 0.00334
R9827 DVDD.n2293 DVDD.n2292 0.00334
R9828 DVDD.n1852 DVDD.n1850 0.00334
R9829 DVDD.n1850 DVDD.n1142 0.00334
R9830 DVDD.n1143 DVDD.n1142 0.00334
R9831 DVDD.n1144 DVDD.n1143 0.00334
R9832 DVDD.n1147 DVDD.n1144 0.00334
R9833 DVDD.n1148 DVDD.n1147 0.00334
R9834 DVDD.n1149 DVDD.n1148 0.00334
R9835 DVDD.n1150 DVDD.n1149 0.00334
R9836 DVDD.n1153 DVDD.n1150 0.00334
R9837 DVDD.n1154 DVDD.n1153 0.00334
R9838 DVDD.n1155 DVDD.n1154 0.00334
R9839 DVDD.n1156 DVDD.n1155 0.00334
R9840 DVDD.n1159 DVDD.n1156 0.00334
R9841 DVDD.n1160 DVDD.n1159 0.00334
R9842 DVDD.n1161 DVDD.n1160 0.00334
R9843 DVDD.n1162 DVDD.n1161 0.00334
R9844 DVDD.n1163 DVDD.n1162 0.00334
R9845 DVDD.n1164 DVDD.n1163 0.00334
R9846 DVDD.n1165 DVDD.n1164 0.00334
R9847 DVDD.n1166 DVDD.n1165 0.00334
R9848 DVDD.n1169 DVDD.n1166 0.00334
R9849 DVDD.n1170 DVDD.n1169 0.00334
R9850 DVDD.n1171 DVDD.n1170 0.00334
R9851 DVDD.n1178 DVDD.n1174 0.00334
R9852 DVDD.n1179 DVDD.n1178 0.00334
R9853 DVDD.n1180 DVDD.n1179 0.00334
R9854 DVDD.n1181 DVDD.n1180 0.00334
R9855 DVDD.n1184 DVDD.n1181 0.00334
R9856 DVDD.n1185 DVDD.n1184 0.00334
R9857 DVDD.n1186 DVDD.n1185 0.00334
R9858 DVDD.n1187 DVDD.n1186 0.00334
R9859 DVDD.n1190 DVDD.n1187 0.00334
R9860 DVDD.n1191 DVDD.n1190 0.00334
R9861 DVDD.n1192 DVDD.n1191 0.00334
R9862 DVDD.n1274 DVDD.n1192 0.00334
R9863 DVDD.n1275 DVDD.n1274 0.00334
R9864 DVDD.n1276 DVDD.n1275 0.00334
R9865 DVDD.n1277 DVDD.n1276 0.00334
R9866 DVDD.n1280 DVDD.n1277 0.00334
R9867 DVDD.n1281 DVDD.n1280 0.00334
R9868 DVDD.n1282 DVDD.n1281 0.00334
R9869 DVDD.n1283 DVDD.n1282 0.00334
R9870 DVDD.n1286 DVDD.n1283 0.00334
R9871 DVDD.n1287 DVDD.n1286 0.00334
R9872 DVDD.n1288 DVDD.n1287 0.00334
R9873 DVDD.n2352 DVDD.n1288 0.00334
R9874 DVDD.n1067 DVDD.n1066 0.00334
R9875 DVDD.n1068 DVDD.n1067 0.00334
R9876 DVDD.n1069 DVDD.n1068 0.00334
R9877 DVDD.n1070 DVDD.n1069 0.00334
R9878 DVDD.n1071 DVDD.n1070 0.00334
R9879 DVDD.n1072 DVDD.n1071 0.00334
R9880 DVDD.n1073 DVDD.n1072 0.00334
R9881 DVDD.n1076 DVDD.n1073 0.00334
R9882 DVDD.n1077 DVDD.n1076 0.00334
R9883 DVDD.n1078 DVDD.n1077 0.00334
R9884 DVDD.n1079 DVDD.n1078 0.00334
R9885 DVDD.n1082 DVDD.n1079 0.00334
R9886 DVDD.n1083 DVDD.n1082 0.00334
R9887 DVDD.n1084 DVDD.n1083 0.00334
R9888 DVDD.n1085 DVDD.n1084 0.00334
R9889 DVDD.n1088 DVDD.n1085 0.00334
R9890 DVDD.n1089 DVDD.n1088 0.00334
R9891 DVDD.n1090 DVDD.n1089 0.00334
R9892 DVDD.n1091 DVDD.n1090 0.00334
R9893 DVDD.n1094 DVDD.n1091 0.00334
R9894 DVDD.n1095 DVDD.n1094 0.00334
R9895 DVDD.n1096 DVDD.n1095 0.00334
R9896 DVDD.n1331 DVDD.n1096 0.00334
R9897 DVDD.n1366 DVDD.n1332 0.00334
R9898 DVDD.n1335 DVDD.n1332 0.00334
R9899 DVDD.n1336 DVDD.n1335 0.00334
R9900 DVDD.n1337 DVDD.n1336 0.00334
R9901 DVDD.n1338 DVDD.n1337 0.00334
R9902 DVDD.n1341 DVDD.n1338 0.00334
R9903 DVDD.n1342 DVDD.n1341 0.00334
R9904 DVDD.n1343 DVDD.n1342 0.00334
R9905 DVDD.n1344 DVDD.n1343 0.00334
R9906 DVDD.n1346 DVDD.n1344 0.00334
R9907 DVDD.n1779 DVDD.n1778 0.00334
R9908 DVDD.n1778 DVDD.n1411 0.00334
R9909 DVDD.n1412 DVDD.n1411 0.00334
R9910 DVDD.n1413 DVDD.n1412 0.00334
R9911 DVDD.n1416 DVDD.n1413 0.00334
R9912 DVDD.n1417 DVDD.n1416 0.00334
R9913 DVDD.n1418 DVDD.n1417 0.00334
R9914 DVDD.n1419 DVDD.n1418 0.00334
R9915 DVDD.n1422 DVDD.n1419 0.00334
R9916 DVDD.n1423 DVDD.n1422 0.00334
R9917 DVDD.n1424 DVDD.n1423 0.00334
R9918 DVDD.n1425 DVDD.n1424 0.00334
R9919 DVDD.n1428 DVDD.n1425 0.00334
R9920 DVDD.n1429 DVDD.n1428 0.00334
R9921 DVDD.n1430 DVDD.n1429 0.00334
R9922 DVDD.n1431 DVDD.n1430 0.00334
R9923 DVDD.n1432 DVDD.n1431 0.00334
R9924 DVDD.n1433 DVDD.n1432 0.00334
R9925 DVDD.n1434 DVDD.n1433 0.00334
R9926 DVDD.n1448 DVDD.n1434 0.00334
R9927 DVDD.n1449 DVDD.n1448 0.00334
R9928 DVDD.n1450 DVDD.n1449 0.00334
R9929 DVDD.n1451 DVDD.n1450 0.00334
R9930 DVDD.n1455 DVDD.n1454 0.00334
R9931 DVDD.n1456 DVDD.n1455 0.00334
R9932 DVDD.n1459 DVDD.n1456 0.00334
R9933 DVDD.n1460 DVDD.n1459 0.00334
R9934 DVDD.n1461 DVDD.n1460 0.00334
R9935 DVDD.n1462 DVDD.n1461 0.00334
R9936 DVDD.n1465 DVDD.n1462 0.00334
R9937 DVDD.n1466 DVDD.n1465 0.00334
R9938 DVDD.n1467 DVDD.n1466 0.00334
R9939 DVDD.n1468 DVDD.n1467 0.00334
R9940 DVDD.n1565 DVDD.n1468 0.00334
R9941 DVDD.n1566 DVDD.n1565 0.00334
R9942 DVDD.n1567 DVDD.n1566 0.00334
R9943 DVDD.n1570 DVDD.n1567 0.00334
R9944 DVDD.n1571 DVDD.n1570 0.00334
R9945 DVDD.n1572 DVDD.n1571 0.00334
R9946 DVDD.n1573 DVDD.n1572 0.00334
R9947 DVDD.n1576 DVDD.n1573 0.00334
R9948 DVDD.n1577 DVDD.n1576 0.00334
R9949 DVDD.n1578 DVDD.n1577 0.00334
R9950 DVDD.n1579 DVDD.n1578 0.00334
R9951 DVDD.n1581 DVDD.n1579 0.00334
R9952 DVDD.n1582 DVDD.n1581 0.00334
R9953 DVDD.n2061 DVDD.n2058 0.00334
R9954 DVDD.n2062 DVDD.n2061 0.00334
R9955 DVDD.n2063 DVDD.n2062 0.00334
R9956 DVDD.n2064 DVDD.n2063 0.00334
R9957 DVDD.n2065 DVDD.n2064 0.00334
R9958 DVDD.n2066 DVDD.n2065 0.00334
R9959 DVDD.n2080 DVDD.n2066 0.00334
R9960 DVDD.n2081 DVDD.n2080 0.00334
R9961 DVDD.n2082 DVDD.n2081 0.00334
R9962 DVDD.n2083 DVDD.n2082 0.00334
R9963 DVDD.n2086 DVDD.n2083 0.00334
R9964 DVDD.n2087 DVDD.n2086 0.00334
R9965 DVDD.n2088 DVDD.n2087 0.00334
R9966 DVDD.n2089 DVDD.n2088 0.00334
R9967 DVDD.n2092 DVDD.n2089 0.00334
R9968 DVDD.n2093 DVDD.n2092 0.00334
R9969 DVDD.n2094 DVDD.n2093 0.00334
R9970 DVDD.n2095 DVDD.n2094 0.00334
R9971 DVDD.n2098 DVDD.n2095 0.00334
R9972 DVDD.n2100 DVDD.n2098 0.00334
R9973 DVDD.n2100 DVDD.n2099 0.00334
R9974 DVDD.n2099 DVDD.n1368 0.00334
R9975 DVDD.n2240 DVDD.n1368 0.00334
R9976 DVDD.n2243 DVDD.n2242 0.00334
R9977 DVDD.n2244 DVDD.n2243 0.00334
R9978 DVDD.n2247 DVDD.n2244 0.00334
R9979 DVDD.n2248 DVDD.n2247 0.00334
R9980 DVDD.n2249 DVDD.n2248 0.00334
R9981 DVDD.n2250 DVDD.n2249 0.00334
R9982 DVDD.n2253 DVDD.n2250 0.00334
R9983 DVDD.n2254 DVDD.n2253 0.00334
R9984 DVDD.n2255 DVDD.n2254 0.00334
R9985 DVDD.n2256 DVDD.n2255 0.00334
R9986 DVDD.n2257 DVDD.n2256 0.00334
R9987 DVDD.n1847 DVDD.n1782 0.00334
R9988 DVDD.n1786 DVDD.n1782 0.00334
R9989 DVDD.n1800 DVDD.n1786 0.00334
R9990 DVDD.n1801 DVDD.n1800 0.00334
R9991 DVDD.n1802 DVDD.n1801 0.00334
R9992 DVDD.n1803 DVDD.n1802 0.00334
R9993 DVDD.n1806 DVDD.n1803 0.00334
R9994 DVDD.n1807 DVDD.n1806 0.00334
R9995 DVDD.n1808 DVDD.n1807 0.00334
R9996 DVDD.n1809 DVDD.n1808 0.00334
R9997 DVDD.n1812 DVDD.n1809 0.00334
R9998 DVDD.n1813 DVDD.n1812 0.00334
R9999 DVDD.n1814 DVDD.n1813 0.00334
R10000 DVDD.n1815 DVDD.n1814 0.00334
R10001 DVDD.n1817 DVDD.n1815 0.00334
R10002 DVDD.n1818 DVDD.n1817 0.00334
R10003 DVDD.n1820 DVDD.n1818 0.00334
R10004 DVDD.n1820 DVDD.n1819 0.00334
R10005 DVDD.n1819 DVDD.n1746 0.00334
R10006 DVDD.n1747 DVDD.n1746 0.00334
R10007 DVDD.n1748 DVDD.n1747 0.00334
R10008 DVDD.n1750 DVDD.n1748 0.00334
R10009 DVDD.n1751 DVDD.n1750 0.00334
R10010 DVDD.n1949 DVDD.n1946 0.00334
R10011 DVDD.n1950 DVDD.n1949 0.00334
R10012 DVDD.n1951 DVDD.n1950 0.00334
R10013 DVDD.n1952 DVDD.n1951 0.00334
R10014 DVDD.n1955 DVDD.n1952 0.00334
R10015 DVDD.n1956 DVDD.n1955 0.00334
R10016 DVDD.n1957 DVDD.n1956 0.00334
R10017 DVDD.n1958 DVDD.n1957 0.00334
R10018 DVDD.n1959 DVDD.n1958 0.00334
R10019 DVDD.n1960 DVDD.n1959 0.00334
R10020 DVDD.n1961 DVDD.n1960 0.00334
R10021 DVDD.n1962 DVDD.n1961 0.00334
R10022 DVDD.n1963 DVDD.n1962 0.00334
R10023 DVDD.n1966 DVDD.n1963 0.00334
R10024 DVDD.n1967 DVDD.n1966 0.00334
R10025 DVDD.n1968 DVDD.n1967 0.00334
R10026 DVDD.n1969 DVDD.n1968 0.00334
R10027 DVDD.n1972 DVDD.n1969 0.00334
R10028 DVDD.n1973 DVDD.n1972 0.00334
R10029 DVDD.n1974 DVDD.n1973 0.00334
R10030 DVDD.n1975 DVDD.n1974 0.00334
R10031 DVDD.n1978 DVDD.n1975 0.00334
R10032 DVDD.n1978 DVDD.n1977 0.00334
R10033 DVDD.n1588 DVDD.n1584 0.00334
R10034 DVDD.n1589 DVDD.n1588 0.00334
R10035 DVDD.n1590 DVDD.n1589 0.00334
R10036 DVDD.n1591 DVDD.n1590 0.00334
R10037 DVDD.n1609 DVDD.n1591 0.00334
R10038 DVDD.n1610 DVDD.n1609 0.00334
R10039 DVDD.n1611 DVDD.n1610 0.00334
R10040 DVDD.n1612 DVDD.n1611 0.00334
R10041 DVDD.n1615 DVDD.n1612 0.00334
R10042 DVDD.n1616 DVDD.n1615 0.00334
R10043 DVDD.n1617 DVDD.n1616 0.00334
R10044 DVDD.n1618 DVDD.n1617 0.00334
R10045 DVDD.n1621 DVDD.n1618 0.00334
R10046 DVDD.n1622 DVDD.n1621 0.00334
R10047 DVDD.n1623 DVDD.n1622 0.00334
R10048 DVDD.n1624 DVDD.n1623 0.00334
R10049 DVDD.n1627 DVDD.n1624 0.00334
R10050 DVDD.n1628 DVDD.n1627 0.00334
R10051 DVDD.n1629 DVDD.n1628 0.00334
R10052 DVDD.n1630 DVDD.n1629 0.00334
R10053 DVDD.n1631 DVDD.n1630 0.00334
R10054 DVDD.n1632 DVDD.n1631 0.00334
R10055 DVDD.n1633 DVDD.n1632 0.00334
R10056 DVDD.n1637 DVDD.n1634 0.00334
R10057 DVDD.n1638 DVDD.n1637 0.00334
R10058 DVDD.n1639 DVDD.n1638 0.00334
R10059 DVDD.n1640 DVDD.n1639 0.00334
R10060 DVDD.n1643 DVDD.n1640 0.00334
R10061 DVDD.n1644 DVDD.n1643 0.00334
R10062 DVDD.n1645 DVDD.n1644 0.00334
R10063 DVDD.n1646 DVDD.n1645 0.00334
R10064 DVDD.n1648 DVDD.n1646 0.00334
R10065 DVDD.n1649 DVDD.n1648 0.00334
R10066 DVDD.n2980 DVDD.n2979 0.00334
R10067 DVDD.n2981 DVDD.n2980 0.00334
R10068 DVDD.n2981 DVDD.n772 0.00334
R10069 DVDD.n2987 DVDD.n772 0.00334
R10070 DVDD.n2988 DVDD.n2987 0.00334
R10071 DVDD.n2989 DVDD.n2988 0.00334
R10072 DVDD.n2989 DVDD.n768 0.00334
R10073 DVDD.n2995 DVDD.n768 0.00334
R10074 DVDD.n2996 DVDD.n2995 0.00334
R10075 DVDD.n2997 DVDD.n2996 0.00334
R10076 DVDD.n2997 DVDD.n764 0.00334
R10077 DVDD.n3003 DVDD.n764 0.00334
R10078 DVDD.n3004 DVDD.n3003 0.00334
R10079 DVDD.n3006 DVDD.n3004 0.00334
R10080 DVDD.n3006 DVDD.n3005 0.00334
R10081 DVDD.n3005 DVDD.n760 0.00334
R10082 DVDD.n3013 DVDD.n760 0.00334
R10083 DVDD.n3014 DVDD.n3013 0.00334
R10084 DVDD.n3015 DVDD.n3014 0.00334
R10085 DVDD.n3016 DVDD.n3015 0.00334
R10086 DVDD.n3017 DVDD.n3016 0.00334
R10087 DVDD.n3018 DVDD.n3017 0.00334
R10088 DVDD.n3018 DVDD.n282 0.00334
R10089 DVDD.n4963 DVDD.n283 0.00334
R10090 DVDD.n4964 DVDD.n4963 0.00334
R10091 DVDD.n4965 DVDD.n4964 0.00334
R10092 DVDD.n4965 DVDD.n4955 0.00334
R10093 DVDD.n4971 DVDD.n4955 0.00334
R10094 DVDD.n4972 DVDD.n4971 0.00334
R10095 DVDD.n4973 DVDD.n4972 0.00334
R10096 DVDD.n4973 DVDD.n4951 0.00334
R10097 DVDD.n4979 DVDD.n4951 0.00334
R10098 DVDD.n4980 DVDD.n4979 0.00334
R10099 DVDD.n4981 DVDD.n4980 0.00334
R10100 DVDD.n4982 DVDD.n4981 0.00334
R10101 DVDD.n4983 DVDD.n4982 0.00334
R10102 DVDD.n4986 DVDD.n4983 0.00334
R10103 DVDD.n4987 DVDD.n4986 0.00334
R10104 DVDD.n4988 DVDD.n4987 0.00334
R10105 DVDD.n4989 DVDD.n4988 0.00334
R10106 DVDD.n4992 DVDD.n4989 0.00334
R10107 DVDD.n4993 DVDD.n4992 0.00334
R10108 DVDD.n4994 DVDD.n4993 0.00334
R10109 DVDD.n4995 DVDD.n4994 0.00334
R10110 DVDD.n4998 DVDD.n4995 0.00334
R10111 DVDD.n4999 DVDD.n4998 0.00334
R10112 DVDD.n5074 DVDD.n5071 0.00334
R10113 DVDD.n5075 DVDD.n5074 0.00334
R10114 DVDD.n5076 DVDD.n5075 0.00334
R10115 DVDD.n5077 DVDD.n5076 0.00334
R10116 DVDD.n5156 DVDD.n5077 0.00334
R10117 DVDD.n5157 DVDD.n5156 0.00334
R10118 DVDD.n5158 DVDD.n5157 0.00334
R10119 DVDD.n5159 DVDD.n5158 0.00334
R10120 DVDD.n5162 DVDD.n5159 0.00334
R10121 DVDD.n5163 DVDD.n5162 0.00334
R10122 DVDD.n5164 DVDD.n5163 0.00334
R10123 DVDD.n5165 DVDD.n5164 0.00334
R10124 DVDD.n5168 DVDD.n5165 0.00334
R10125 DVDD.n5169 DVDD.n5168 0.00334
R10126 DVDD.n5170 DVDD.n5169 0.00334
R10127 DVDD.n5171 DVDD.n5170 0.00334
R10128 DVDD.n5174 DVDD.n5171 0.00334
R10129 DVDD.n5175 DVDD.n5174 0.00334
R10130 DVDD.n5176 DVDD.n5175 0.00334
R10131 DVDD.n5178 DVDD.n5176 0.00334
R10132 DVDD.n5178 DVDD.n5177 0.00334
R10133 DVDD.n5177 DVDD.n698 0.00334
R10134 DVDD.n698 DVDD.n659 0.00334
R10135 DVDD.n5430 DVDD.n660 0.00334
R10136 DVDD.n5398 DVDD.n660 0.00334
R10137 DVDD.n5399 DVDD.n5398 0.00334
R10138 DVDD.n5400 DVDD.n5399 0.00334
R10139 DVDD.n5403 DVDD.n5400 0.00334
R10140 DVDD.n5404 DVDD.n5403 0.00334
R10141 DVDD.n5405 DVDD.n5404 0.00334
R10142 DVDD.n5406 DVDD.n5405 0.00334
R10143 DVDD.n5408 DVDD.n5406 0.00334
R10144 DVDD.n5409 DVDD.n5408 0.00334
R10145 DVDD.n4699 DVDD.n4698 0.00334
R10146 DVDD.n4699 DVDD.n3155 0.00334
R10147 DVDD.n4710 DVDD.n3164 0.00334
R10148 DVDD.n4711 DVDD.n4710 0.00334
R10149 DVDD.n4711 DVDD.n3361 0.00334
R10150 DVDD.n4721 DVDD.n3361 0.00334
R10151 DVDD.n4734 DVDD.n4722 0.00334
R10152 DVDD.n4734 DVDD.n4733 0.00334
R10153 DVDD.n4733 DVDD.n4732 0.00334
R10154 DVDD.n4732 DVDD.n4723 0.00334
R10155 DVDD.n5743 DVDD.n5742 0.00334
R10156 DVDD.n5742 DVDD.n5741 0.00334
R10157 DVDD.n5741 DVDD.n204 0.00334
R10158 DVDD.n5737 DVDD.n204 0.00334
R10159 DVDD.n5736 DVDD.n5735 0.00334
R10160 DVDD.n5735 DVDD.n209 0.00334
R10161 DVDD.n5731 DVDD.n209 0.00334
R10162 DVDD.n5731 DVDD.n5730 0.00334
R10163 DVDD.n3049 DVDD.n224 0.00334
R10164 DVDD.n3049 DVDD.n3048 0.00334
R10165 DVDD.n3488 DVDD.n3487 0.00334
R10166 DVDD.n3488 DVDD.n3165 0.00334
R10167 DVDD.n3250 DVDD.n3166 0.00334
R10168 DVDD.n3251 DVDD.n3250 0.00334
R10169 DVDD.n3252 DVDD.n3251 0.00334
R10170 DVDD.n4792 DVDD.n3252 0.00334
R10171 DVDD.n4794 DVDD.n4793 0.00334
R10172 DVDD.n4795 DVDD.n4794 0.00334
R10173 DVDD.n4797 DVDD.n4795 0.00334
R10174 DVDD.n4797 DVDD.n4796 0.00334
R10175 DVDD.n3084 DVDD.n3083 0.00334
R10176 DVDD.n3085 DVDD.n3084 0.00334
R10177 DVDD.n3091 DVDD.n3085 0.00334
R10178 DVDD.n3092 DVDD.n3091 0.00334
R10179 DVDD.n3094 DVDD.n3093 0.00334
R10180 DVDD.n3101 DVDD.n3094 0.00334
R10181 DVDD.n3102 DVDD.n3101 0.00334
R10182 DVDD.n3102 DVDD.n228 0.00334
R10183 DVDD.n5728 DVDD.n229 0.00334
R10184 DVDD.n238 DVDD.n229 0.00334
R10185 DVDD.n4511 DVDD.n4510 0.00334
R10186 DVDD.n4510 DVDD.n3156 0.00334
R10187 DVDD.n4867 DVDD.n4864 0.00334
R10188 DVDD.n4867 DVDD.n4866 0.00334
R10189 DVDD.n4866 DVDD.n4865 0.00334
R10190 DVDD.n4865 DVDD.n3137 0.00334
R10191 DVDD.n4889 DVDD.n4888 0.00334
R10192 DVDD.n4892 DVDD.n4889 0.00334
R10193 DVDD.n4892 DVDD.n4891 0.00334
R10194 DVDD.n4891 DVDD.n4890 0.00334
R10195 DVDD.n5094 DVDD.n5093 0.00334
R10196 DVDD.n5100 DVDD.n5094 0.00334
R10197 DVDD.n5100 DVDD.n5099 0.00334
R10198 DVDD.n5099 DVDD.n5098 0.00334
R10199 DVDD.n5115 DVDD.n5084 0.00334
R10200 DVDD.n5116 DVDD.n5115 0.00334
R10201 DVDD.n5117 DVDD.n5116 0.00334
R10202 DVDD.n5117 DVDD.n219 0.00334
R10203 DVDD.n5133 DVDD.n220 0.00334
R10204 DVDD.n5134 DVDD.n5133 0.00334
R10205 DVDD.n3193 DVDD.n3192 0.00334
R10206 DVDD.n3193 DVDD.n3160 0.00334
R10207 DVDD.n3202 DVDD.n3161 0.00334
R10208 DVDD.n3203 DVDD.n3202 0.00334
R10209 DVDD.n3204 DVDD.n3203 0.00334
R10210 DVDD.n3207 DVDD.n3204 0.00334
R10211 DVDD.n3209 DVDD.n3208 0.00334
R10212 DVDD.n3216 DVDD.n3209 0.00334
R10213 DVDD.n3218 DVDD.n3216 0.00334
R10214 DVDD.n3218 DVDD.n3217 0.00334
R10215 DVDD.n721 DVDD.n720 0.00334
R10216 DVDD.n5331 DVDD.n721 0.00334
R10217 DVDD.n5332 DVDD.n5331 0.00334
R10218 DVDD.n5333 DVDD.n5332 0.00334
R10219 DVDD.n5344 DVDD.n710 0.00334
R10220 DVDD.n5345 DVDD.n5344 0.00334
R10221 DVDD.n5346 DVDD.n5345 0.00334
R10222 DVDD.n5346 DVDD.n217 0.00334
R10223 DVDD.n703 DVDD.n216 0.00334
R10224 DVDD.n5363 DVDD.n703 0.00334
R10225 DVDD.n1846 DVDD.n1785 0.00332
R10226 DVDD.n1784 DVDD.n1783 0.00332
R10227 DVDD.n1851 DVDD.n1776 0.00332
R10228 DVDD.n1859 DVDD.n1774 0.00332
R10229 DVDD.n1858 DVDD.n1857 0.00332
R10230 DVDD.n1855 DVDD.n1123 0.00332
R10231 DVDD.n1775 DVDD.n1393 0.00332
R10232 DVDD.n1780 DVDD.n882 0.00332
R10233 DVDD.n2978 DVDD.n2977 0.00332
R10234 DVDD.n828 DVDD.n242 0.00332
R10235 DVDD.n4519 DVDD.n4502 0.00329
R10236 DVDD.n5089 DVDD.n4903 0.00329
R10237 DVDD.n5119 DVDD.n4922 0.00329
R10238 DVDD.n4703 DVDD.n4701 0.00329
R10239 DVDD.n3076 DVDD.n3075 0.00329
R10240 DVDD.n3056 DVDD.n212 0.00329
R10241 DVDD.n3494 DVDD.n3491 0.00329
R10242 DVDD.n3126 DVDD.n3125 0.00329
R10243 DVDD.n3106 DVDD.n3100 0.00329
R10244 DVDD.n3197 DVDD.n3195 0.00329
R10245 DVDD.n5324 DVDD.n5323 0.00329
R10246 DVDD.n5350 DVDD.n708 0.00329
R10247 DVDD.n2318 DVDD.n1006 0.00323
R10248 DVDD.n2460 DVDD.n1093 0.00323
R10249 DVDD.n2097 DVDD.n1370 0.00323
R10250 DVDD.n1674 DVDD.n580 0.00323
R10251 DVDD.n5391 DVDD.n699 0.00323
R10252 DVDD.n5036 DVDD.n5035 0.0032
R10253 DVDD.n2977 DVDD.n788 0.0032
R10254 DVDD.n828 DVDD.n827 0.0032
R10255 DVDD.n5622 DVDD.n454 0.00311
R10256 DVDD.n2438 DVDD.n2425 0.00311
R10257 DVDD.n2216 DVDD.n2205 0.00311
R10258 DVDD.n1843 DVDD.n1798 0.00311
R10259 DVDD.n2983 DVDD.n784 0.00311
R10260 DVDD.n5719 DVDD.n239 0.00309529
R10261 DVDD.n3500 DVDD.n3485 0.00309529
R10262 DVDD.n3047 DVDD.n3046 0.00309529
R10263 DVDD.n4697 DVDD.n4696 0.00309529
R10264 DVDD.n5136 DVDD.n5135 0.00309529
R10265 DVDD.n4508 DVDD.n3429 0.00309529
R10266 DVDD.n5364 DVDD.n702 0.00309529
R10267 DVDD.n3191 DVDD.n3190 0.00309529
R10268 DVDD.n4869 DVDD.n3150 0.00305
R10269 DVDD.n4898 DVDD.n3130 0.00305
R10270 DVDD.n5131 DVDD.n4923 0.00305
R10271 DVDD.n4708 DVDD.n4707 0.00305
R10272 DVDD.n4730 DVDD.n4729 0.00305
R10273 DVDD.n3052 DVDD.n3051 0.00305
R10274 DVDD.n4858 DVDD.n3246 0.00305
R10275 DVDD.n4801 DVDD.n4799 0.00305
R10276 DVDD.n5725 DVDD.n234 0.00305
R10277 DVDD.n3240 DVDD.n3177 0.00305
R10278 DVDD.n3220 DVDD.n3215 0.00305
R10279 DVDD.n5356 DVDD.n5355 0.00305
R10280 DVDD.n1539 DVDD.n1389 0.00301866
R10281 DVDD.n1253 DVDD.n1252 0.00301866
R10282 DVDD.n3763 DVDD.n3697 0.00294565
R10283 DVDD.n4205 DVDD.n3509 0.00294565
R10284 DVDD.n3549 DVDD.n3548 0.00294565
R10285 DVDD.n4185 DVDD.n3528 0.00294565
R10286 DVDD.n1330 DVDD.n1322 0.00286
R10287 DVDD.n1367 DVDD.n1366 0.00286
R10288 DVDD.n2242 DVDD.n2241 0.00286
R10289 DVDD.n1634 DVDD.n1329 0.00286
R10290 DVDD.n5431 DVDD.n5430 0.00286
R10291 DVDD.n2528 DVDD.n1017 0.00285923
R10292 DVDD.n2373 DVDD.n1195 0.00285923
R10293 DVDD.n355 DVDD.n346 0.00285923
R10294 DVDD.n346 DVDD.n313 0.00285923
R10295 DVDD.n2371 DVDD.n1195 0.00285923
R10296 DVDD.n2528 DVDD.n1015 0.00285923
R10297 DVDD DVDD.n2293 0.00278
R10298 DVDD DVDD.n1346 0.00278
R10299 DVDD DVDD.n1649 0.00278
R10300 DVDD DVDD.n5409 0.00278
R10301 DVDD.n864 DVDD.n848 0.00275
R10302 DVDD.n287 DVDD.n280 0.00275
R10303 DVDD.n860 DVDD.n850 0.00275
R10304 DVDD.n285 DVDD.n281 0.00275
R10305 DVDD.n4518 DVDD.n3169 0.00275
R10306 DVDD.n5321 DVDD.n732 0.00275
R10307 DVDD.n5082 DVDD.n233 0.00275
R10308 DVDD.n4861 DVDD.n3244 0.00275
R10309 DVDD.n5745 DVDD.n189 0.00275
R10310 DVDD.n3104 DVDD.n230 0.00275
R10311 DVDD.n4702 DVDD.n3169 0.00275
R10312 DVDD.n5321 DVDD.n202 0.00275
R10313 DVDD.n3055 DVDD.n233 0.00275
R10314 DVDD.n3493 DVDD.n3169 0.00275
R10315 DVDD.n5321 DVDD.n3080 0.00275
R10316 DVDD.n3103 DVDD.n233 0.00275
R10317 DVDD.n4861 DVDD.n3243 0.00275
R10318 DVDD.n5745 DVDD.n198 0.00275
R10319 DVDD.n5083 DVDD.n230 0.00275
R10320 DVDD.n4861 DVDD.n3173 0.00275
R10321 DVDD.n5745 DVDD.n5744 0.00275
R10322 DVDD.n230 DVDD.n213 0.00275
R10323 DVDD.n4861 DVDD.n3175 0.00275
R10324 DVDD.n5745 DVDD.n192 0.00275
R10325 DVDD.n5348 DVDD.n230 0.00275
R10326 DVDD.n3196 DVDD.n3169 0.00275
R10327 DVDD.n5322 DVDD.n5321 0.00275
R10328 DVDD.n5349 DVDD.n233 0.00275
R10329 DVDD.n3873 DVDD.n3582 0.00275
R10330 DVDD.n3955 DVDD.n3954 0.00275
R10331 DVDD.n2350 DVDD.n2349 0.0027
R10332 DVDD.n2351 DVDD.n1066 0.0027
R10333 DVDD.n2058 DVDD.n1289 0.0027
R10334 DVDD.n1976 DVDD.n1584 0.0027
R10335 DVDD.n5071 DVDD.n5070 0.0027
R10336 DVDD.n1858 DVDD.n472 0.00269
R10337 DVDD.n2935 DVDD.n982 0.00269
R10338 DVDD.n2441 DVDD.n1123 0.00269
R10339 DVDD.n2457 DVDD.n2456 0.00269
R10340 DVDD.n2220 DVDD.n1393 0.00269
R10341 DVDD.n2237 DVDD.n2236 0.00269
R10342 DVDD.n2969 DVDD.n882 0.00269
R10343 DVDD.n5497 DVDD.n581 0.00269
R10344 DVDD.n5713 DVDD.n242 0.00269
R10345 DVDD.n5392 DVDD.n696 0.00269
R10346 DVDD.n5729 DVDD 0.00267716
R10347 DVDD.n4863 DVDD 0.00267716
R10348 DVDD.n5457 DVDD.n5454 0.0026
R10349 DVDD.n472 DVDD.n448 0.00257
R10350 DVDD.n2935 DVDD.n988 0.00257
R10351 DVDD.n2441 DVDD.n1128 0.00257
R10352 DVDD.n2456 DVDD.n1100 0.00257
R10353 DVDD.n2220 DVDD.n1398 0.00257
R10354 DVDD.n2236 DVDD.n1326 0.00257
R10355 DVDD.n2969 DVDD.n887 0.00257
R10356 DVDD.n5497 DVDD.n603 0.00257
R10357 DVDD.n5713 DVDD.n243 0.00257
R10358 DVDD.n5395 DVDD.n696 0.00257
R10359 DVDD.n1942 DVDD.n1941 0.00254
R10360 DVDD.n1943 DVDD.n1174 0.00254
R10361 DVDD.n1944 DVDD.n1454 0.00254
R10362 DVDD.n1946 DVDD.n1945 0.00254
R10363 DVDD.n5690 DVDD.n283 0.00254
R10364 DVDD.n3169 DVDD.n3168 0.00251
R10365 DVDD.n5321 DVDD.n726 0.00251
R10366 DVDD.n5128 DVDD.n233 0.00251
R10367 DVDD.n4861 DVDD.n4860 0.00251
R10368 DVDD.n5745 DVDD.n190 0.00251
R10369 DVDD.n5727 DVDD.n230 0.00251
R10370 DVDD.n3366 DVDD.n3169 0.00251
R10371 DVDD.n5321 DVDD.n734 0.00251
R10372 DVDD.n736 DVDD.n233 0.00251
R10373 DVDD.n4859 DVDD.n3169 0.00251
R10374 DVDD.n5321 DVDD.n3079 0.00251
R10375 DVDD.n5726 DVDD.n233 0.00251
R10376 DVDD.n4861 DVDD.n3151 0.00251
R10377 DVDD.n5745 DVDD.n199 0.00251
R10378 DVDD.n5129 DVDD.n230 0.00251
R10379 DVDD.n4861 DVDD.n3172 0.00251
R10380 DVDD.n5745 DVDD.n201 0.00251
R10381 DVDD.n738 DVDD.n230 0.00251
R10382 DVDD.n4861 DVDD.n3242 0.00251
R10383 DVDD.n5745 DVDD.n193 0.00251
R10384 DVDD.n5353 DVDD.n230 0.00251
R10385 DVDD.n3241 DVDD.n3169 0.00251
R10386 DVDD.n5321 DVDD.n728 0.00251
R10387 DVDD.n5354 DVDD.n233 0.00251
R10388 DVDD.n1860 DVDD.n1773 0.00238
R10389 DVDD.n1853 DVDD.n1852 0.00238
R10390 DVDD.n1849 DVDD.n1779 0.00238
R10391 DVDD.n1848 DVDD.n1847 0.00238
R10392 DVDD.n2979 DVDD.n786 0.00238
R10393 DVDD.n5612 DVDD.n5608 0.00236429
R10394 DVDD.n5575 DVDD.n506 0.00236429
R10395 DVDD.n3957 DVDD.n3956 0.00236429
R10396 DVDD.n3989 DVDD.n3627 0.00236429
R10397 DVDD.n3468 DVDD.n3374 0.00236429
R10398 DVDD.n4493 DVDD.n3433 0.00236429
R10399 DVDD.n2685 DVDD 0.0023
R10400 DVDD.n5054 DVDD.n4997 0.0023
R10401 DVDD.n5224 DVDD.n5000 0.0023
R10402 DVDD.n5032 DVDD.n5010 0.0023
R10403 DVDD.n823 DVDD.n786 0.0023
R10404 DVDD.n803 DVDD.n800 0.0023
R10405 DVDD.n802 DVDD.n799 0.0023
R10406 DVDD.n4079 DVDD 0.0023
R10407 DVDD.n6018 DVDD 0.0023
R10408 DVDD.n3168 DVDD.n3150 0.00221
R10409 DVDD.n4898 DVDD.n726 0.00221
R10410 DVDD.n5128 DVDD.n4923 0.00221
R10411 DVDD.n4707 DVDD.n3366 0.00221
R10412 DVDD.n4729 DVDD.n734 0.00221
R10413 DVDD.n3052 DVDD.n736 0.00221
R10414 DVDD.n4859 DVDD.n4858 0.00221
R10415 DVDD.n4801 DVDD.n3079 0.00221
R10416 DVDD.n5726 DVDD.n5725 0.00221
R10417 DVDD.n3241 DVDD.n3240 0.00221
R10418 DVDD.n3215 DVDD.n728 0.00221
R10419 DVDD.n5356 DVDD.n5354 0.00221
R10420 DVDD.n3842 DVDD.n3435 0.0021791
R10421 DVDD.n5622 DVDD.n448 0.00215
R10422 DVDD.n2438 DVDD.n1128 0.00215
R10423 DVDD.n2216 DVDD.n1398 0.00215
R10424 DVDD.n1798 DVDD.n887 0.00215
R10425 DVDD.n784 DVDD.n243 0.00215
R10426 DVDD.n5703 DVDD.n263 0.00213125
R10427 DVDD.n5568 DVDD.n516 0.00210714
R10428 DVDD.n2754 DVDD.n2609 0.00210714
R10429 DVDD.n4002 DVDD.n4001 0.00210714
R10430 DVDD.n4038 DVDD.n4037 0.00210714
R10431 DVDD.n4488 DVDD.n4485 0.00210714
R10432 DVDD.n4412 DVDD.n3427 0.00210714
R10433 DVDD.n1006 DVDD.n982 0.00203
R10434 DVDD.n2457 DVDD.n1093 0.00203
R10435 DVDD.n2237 DVDD.n1370 0.00203
R10436 DVDD.n581 DVDD.n580 0.00203
R10437 DVDD.n5392 DVDD.n5391 0.00203
R10438 DVDD.n2561 DVDD.n2559 0.00201119
R10439 DVDD.n862 DVDD.n861 0.002
R10440 DVDD.n5691 DVDD.n5690 0.002
R10441 DVDD.n4863 DVDD.n3155 0.002
R10442 DVDD.n5743 DVDD.n184 0.002
R10443 DVDD.n5730 DVDD.n5729 0.002
R10444 DVDD.n4863 DVDD.n3165 0.002
R10445 DVDD.n3083 DVDD.n184 0.002
R10446 DVDD.n5729 DVDD.n228 0.002
R10447 DVDD.n4863 DVDD.n3156 0.002
R10448 DVDD.n5093 DVDD.n184 0.002
R10449 DVDD.n5729 DVDD.n219 0.002
R10450 DVDD.n4863 DVDD.n3160 0.002
R10451 DVDD.n720 DVDD.n184 0.002
R10452 DVDD.n5729 DVDD.n217 0.002
R10453 DVDD.n4519 DVDD.n4518 0.00197
R10454 DVDD.n4903 DVDD.n732 0.00197
R10455 DVDD.n5082 DVDD.n4922 0.00197
R10456 DVDD.n4703 DVDD.n4702 0.00197
R10457 DVDD.n3076 DVDD.n202 0.00197
R10458 DVDD.n3056 DVDD.n3055 0.00197
R10459 DVDD.n3494 DVDD.n3493 0.00197
R10460 DVDD.n3126 DVDD.n3080 0.00197
R10461 DVDD.n3103 DVDD.n3100 0.00197
R10462 DVDD.n3197 DVDD.n3196 0.00197
R10463 DVDD.n5324 DVDD.n5322 0.00197
R10464 DVDD.n5350 DVDD.n5349 0.00197
R10465 DVDD.n5037 DVDD.n296 0.00190625
R10466 DVDD.n644 DVDD.n638 0.00190625
R10467 DVDD.n5396 DVDD.n657 0.00185
R10468 DVDD.n5433 DVDD.n656 0.00185
R10469 DVDD.n4863 DVDD.n3164 0.00184
R10470 DVDD.n4723 DVDD.n184 0.00184
R10471 DVDD.n5729 DVDD.n224 0.00184
R10472 DVDD.n4863 DVDD.n3166 0.00184
R10473 DVDD.n4796 DVDD.n184 0.00184
R10474 DVDD.n5729 DVDD.n5728 0.00184
R10475 DVDD.n4864 DVDD.n4863 0.00184
R10476 DVDD.n4890 DVDD.n184 0.00184
R10477 DVDD.n5729 DVDD.n220 0.00184
R10478 DVDD.n4863 DVDD.n3161 0.00184
R10479 DVDD.n3217 DVDD.n184 0.00184
R10480 DVDD.n5729 DVDD.n216 0.00184
R10481 DVDD.n5669 DVDD.n296 0.00179375
R10482 DVDD DVDD.n2686 0.0017
R10483 DVDD.n2017 DVDD.n2016 0.0017
R10484 DVDD.n2174 DVDD.n1173 0.0017
R10485 DVDD.n2394 DVDD.n2393 0.0017
R10486 DVDD.n1904 DVDD.n1172 0.0017
R10487 DVDD.n1906 DVDD.n1905 0.0017
R10488 DVDD.n1176 DVDD.n1168 0.0017
R10489 DVDD.n2173 DVDD.n2172 0.0017
R10490 DVDD.n2018 DVDD.n1452 0.0017
R10491 DVDD.n5070 DVDD.n5058 0.0017
R10492 DVDD.n806 DVDD.n805 0.0017
R10493 DVDD.n3020 DVDD.n285 0.0017
R10494 DVDD.n3021 DVDD.n287 0.0017
R10495 DVDD.n2153 DVDD.n1552 0.00167537
R10496 DVDD.n1255 DVDD.n1119 0.00167537
R10497 DVDD.n2527 DVDD.n2526 0.00167537
R10498 DVDD.n4870 DVDD.n4869 0.00167
R10499 DVDD.n4895 DVDD.n3130 0.00167
R10500 DVDD.n5131 DVDD.n5130 0.00167
R10501 DVDD.n4708 DVDD.n3365 0.00167
R10502 DVDD.n4730 DVDD.n4725 0.00167
R10503 DVDD.n3051 DVDD.n737 0.00167
R10504 DVDD.n4855 DVDD.n3246 0.00167
R10505 DVDD.n4804 DVDD.n4799 0.00167
R10506 DVDD.n5722 DVDD.n234 0.00167
R10507 DVDD.n3237 DVDD.n3177 0.00167
R10508 DVDD.n3221 DVDD.n3220 0.00167
R10509 DVDD.n5355 DVDD.n705 0.00167
R10510 DVDD DVDD.n671 0.00165261
R10511 DVDD DVDD.n672 0.00165261
R10512 DVDD.n5659 DVDD.n5658 0.001625
R10513 DVDD.n4533 DVDD.n4497 0.001625
R10514 DVDD.n5311 DVDD.n5310 0.001625
R10515 DVDD.n5305 DVDD.n4917 0.001625
R10516 DVDD.n2057 DVDD.n1583 0.00146
R10517 DVDD.n2133 DVDD.n2132 0.00146
R10518 DVDD.n2353 DVDD.n1065 0.00146
R10519 DVDD.n2495 DVDD.n1060 0.00146
R10520 DVDD.n2494 DVDD.n2493 0.00146
R10521 DVDD.n2492 DVDD.n1063 0.00146
R10522 DVDD.n2134 DVDD.n1062 0.00146
R10523 DVDD.n1980 DVDD.n1586 0.00146
R10524 DVDD.n5225 DVDD.n5224 0.00146
R10525 DVDD.n5226 DVDD.n4997 0.00146
R10526 DVDD.n4514 DVDD.n4502 0.00143
R10527 DVDD.n5089 DVDD.n5088 0.00143
R10528 DVDD.n5120 DVDD.n5119 0.00143
R10529 DVDD.n4701 DVDD.n3368 0.00143
R10530 DVDD.n3075 DVDD.n3074 0.00143
R10531 DVDD.n3058 DVDD.n212 0.00143
R10532 DVDD.n3497 DVDD.n3491 0.00143
R10533 DVDD.n3125 DVDD.n3082 0.00143
R10534 DVDD.n3107 DVDD.n3106 0.00143
R10535 DVDD.n3195 DVDD.n3179 0.00143
R10536 DVDD.n5323 DVDD.n723 0.00143
R10537 DVDD.n713 DVDD.n708 0.00143
R10538 DVDD.n5432 DVDD.n5431 0.0014
R10539 DVDD.n5986 DVDD.n5984 0.0014
R10540 DVDD.n4544 DVDD.n4543 0.0014
R10541 DVDD.n4685 DVDD.n4684 0.0014
R10542 DVDD.n4321 DVDD.n4320 0.0014
R10543 DVDD.n2952 DVDD.n952 0.00137
R10544 DVDD.n1925 DVDD.n1016 0.00137
R10545 DVDD.n2959 DVDD.n922 0.00137
R10546 DVDD.n2377 DVDD.n1189 0.00137
R10547 DVDD.n2963 DVDD.n901 0.00137
R10548 DVDD.n2155 DVDD.n2154 0.00137
R10549 DVDD.n2037 DVDD.n1717 0.00137
R10550 DVDD.n5654 DVDD.n314 0.00137
R10551 DVDD.n3040 DVDD.n745 0.00137
R10552 DVDD.n5281 DVDD.n4938 0.00137
R10553 DVDD DVDD.n1652 0.00134
R10554 DVDD.n2258 DVDD 0.00134
R10555 DVDD.n1348 DVDD 0.00134
R10556 DVDD DVDD.n2296 0.00134
R10557 DVDD DVDD.n5412 0.00134
R10558 DVDD.n1942 DVDD.n1752 0.0013
R10559 DVDD.n1943 DVDD.n1171 0.0013
R10560 DVDD.n1944 DVDD.n1451 0.0013
R10561 DVDD.n1945 DVDD.n1751 0.0013
R10562 DVDD.n5690 DVDD.n282 0.0013
R10563 DVDD.n675 DVDD 0.00126841
R10564 DVDD.n2564 DVDD.n2510 0.00125
R10565 DVDD.n5633 DVDD.n436 0.00125
R10566 DVDD.n2369 DVDD.n2368 0.00125
R10567 DVDD.n5639 DVDD.n401 0.00125
R10568 DVDD.n2148 DVDD.n1548 0.00125
R10569 DVDD.n2122 DVDD.n2078 0.00125
R10570 DVDD.n1994 DVDD.n312 0.00125
R10571 DVDD.n1709 DVDD.n1697 0.00125
R10572 DVDD.n5240 DVDD.n4936 0.00125
R10573 DVDD.n5212 DVDD.n5201 0.00125
R10574 DVDD.n1671 DVDD.n1670 0.00122
R10575 DVDD.n2239 DVDD.n1328 0.00122
R10576 DVDD.n1321 DVDD.n1097 0.00122
R10577 DVDD.n2315 DVDD.n2314 0.00122
R10578 DVDD.n2279 DVDD.n988 0.00122
R10579 DVDD.n2278 DVDD.n1100 0.00122
R10580 DVDD.n2277 DVDD.n1326 0.00122
R10581 DVDD.n1325 DVDD.n603 0.00122
R10582 DVDD.n5394 DVDD.n656 0.00122
R10583 DVDD.n5396 DVDD.n5395 0.00122
R10584 DVDD.n5615 DVDD.n478 0.00120714
R10585 DVDD.n2601 DVDD.n2595 0.00120714
R10586 DVDD.n3654 DVDD.n3644 0.00120714
R10587 DVDD.n3998 DVDD.n3997 0.00120714
R10588 DVDD.n4358 DVDD.n3373 0.00120714
R10589 DVDD.n3445 DVDD.n3438 0.00120714
R10590 DVDD.n5096 DVDD.n4913 0.00119
R10591 DVDD.n5095 DVDD.n4914 0.00119
R10592 DVDD.n3067 DVDD.n207 0.00119
R10593 DVDD.n3065 DVDD.n3064 0.00119
R10594 DVDD.n3117 DVDD.n3116 0.00119
R10595 DVDD.n3096 DVDD.n3090 0.00119
R10596 DVDD.n5336 DVDD.n5335 0.00119
R10597 DVDD.n718 DVDD.n712 0.00119
R10598 DVDD.n5020 DVDD.n5019 0.001175
R10599 DVDD.n3146 DVDD.n3141 0.001175
R10600 DVDD.n5753 DVDD.n5752 0.001175
R10601 DVDD.n5286 DVDD.n5285 0.001175
R10602 DVDD.n2350 DVDD.n1059 0.00114
R10603 DVDD.n2352 DVDD.n2351 0.00114
R10604 DVDD.n1582 DVDD.n1289 0.00114
R10605 DVDD.n1977 DVDD.n1976 0.00114
R10606 DVDD.n5070 DVDD.n4999 0.00114
R10607 DVDD.n4875 DVDD.n3148 0.00113
R10608 DVDD.n4894 DVDD.n3133 0.00113
R10609 DVDD.n5138 DVDD.n5126 0.00113
R10610 DVDD.n4714 DVDD.n4713 0.00113
R10611 DVDD.n4724 DVDD.n3358 0.00113
R10612 DVDD.n742 DVDD.n741 0.00113
R10613 DVDD.n4854 DVDD.n3249 0.00113
R10614 DVDD.n4805 DVDD.n4790 0.00113
R10615 DVDD.n5721 DVDD.n237 0.00113
R10616 DVDD.n3236 DVDD.n3201 0.00113
R10617 DVDD.n3224 DVDD.n3212 0.00113
R10618 DVDD.n5361 DVDD.n5360 0.00113
R10619 DVDD.n5702 DVDD.n273 0.00111875
R10620 DVDD.n2294 DVDD 0.00106
R10621 DVDD.n1347 DVDD 0.00106
R10622 DVDD.n1650 DVDD 0.00106
R10623 DVDD.n5410 DVDD 0.00106
R10624 DVDD.n1330 DVDD.n1320 0.00098
R10625 DVDD.n1367 DVDD.n1331 0.00098
R10626 DVDD.n2241 DVDD.n2240 0.00098
R10627 DVDD.n1633 DVDD.n1329 0.00098
R10628 DVDD.n5431 DVDD.n659 0.00098
R10629 DVDD.n5569 DVDD.n510 0.00095
R10630 DVDD.n2751 DVDD.n2607 0.00095
R10631 DVDD.n4885 DVDD.n4884 0.00095
R10632 DVDD.n5756 DVDD.n176 0.00095
R10633 DVDD.n4719 DVDD.n4718 0.00095
R10634 DVDD.n4738 DVDD.n3357 0.00095
R10635 DVDD.n4788 DVDD.n3254 0.00095
R10636 DVDD.n4810 DVDD.n4789 0.00095
R10637 DVDD.n3230 DVDD.n3229 0.00095
R10638 DVDD.n3228 DVDD.n3206 0.00095
R10639 DVDD.n3622 DVDD.n3605 0.00095
R10640 DVDD.n4035 DVDD.n3575 0.00095
R10641 DVDD.n1260 DVDD.n1259 0.00095
R10642 DVDD.n2536 DVDD.n2535 0.00095
R10643 DVDD.n5641 DVDD.n399 0.00095
R10644 DVDD.n2537 DVDD.n424 0.00095
R10645 DVDD.n2958 DVDD.n938 0.00095
R10646 DVDD.n2530 DVDD.n963 0.00095
R10647 DVDD.n2440 DVDD.n1138 0.00095
R10648 DVDD.n2532 DVDD.n2531 0.00095
R10649 DVDD.n4491 DVDD.n3441 0.00095
R10650 DVDD.n4409 DVDD.n3426 0.00095
R10651 DVDD.n5469 DVDD.n5468 0.00089375
R10652 DVDD.n4513 DVDD.n4507 0.00089
R10653 DVDD.n5103 DVDD.n5102 0.00089
R10654 DVDD.n5111 DVDD.n5080 0.00089
R10655 DVDD.n3372 DVDD.n3371 0.00089
R10656 DVDD.n3071 DVDD.n205 0.00089
R10657 DVDD.n3061 DVDD.n211 0.00089
R10658 DVDD.n3498 DVDD.n3490 0.00089
R10659 DVDD.n3122 DVDD.n3121 0.00089
R10660 DVDD.n3099 DVDD.n3097 0.00089
R10661 DVDD.n3183 DVDD.n3182 0.00089
R10662 DVDD.n5329 DVDD.n5328 0.00089
R10663 DVDD.n715 DVDD.n714 0.00089
R10664 DVDD.n4640 DVDD.n3401 0.000835821
R10665 DVDD.n2949 DVDD.n959 0.00083
R10666 DVDD.n1922 DVDD.n1017 0.00083
R10667 DVDD.n2956 DVDD.n927 0.00083
R10668 DVDD.n2374 DVDD.n2373 0.00083
R10669 DVDD.n1446 DVDD.n907 0.00083
R10670 DVDD.n1564 DVDD.n1481 0.00083
R10671 DVDD.n2034 DVDD.n1723 0.00083
R10672 DVDD.n355 DVDD.n326 0.00083
R10673 DVDD.n3037 DVDD.n746 0.00083
R10674 DVDD.n5278 DVDD.n5245 0.00083
R10675 DVDD.n1018 DVDD.n1015 0.00071
R10676 DVDD.n5635 DVDD.n420 0.00071
R10677 DVDD.n2371 DVDD.n1222 0.00071
R10678 DVDD.n5642 DVDD.n388 0.00071
R10679 DVDD.n2152 DVDD.n2151 0.00071
R10680 DVDD.n5646 DVDD.n368 0.00071
R10681 DVDD.n1996 DVDD.n313 0.00071
R10682 DVDD.n2048 DVDD.n1599 0.00071
R10683 DVDD.n5242 DVDD.n4937 0.00071
R10684 DVDD.n5215 DVDD.n5143 0.00071
R10685 DVDD.n6017 DVDD 0.000671429
R10686 DVDD.n2686 DVDD 0.000671429
R10687 DVDD.n4080 DVDD 0.000671429
R10688 DVDD.n2370 DVDD.n1264 0.00066791
R10689 DVDD.n2542 DVDD.n2541 0.00066791
R10690 DVDD.n4504 DVDD.n3430 0.00065
R10691 DVDD.n5091 DVDD.n4912 0.00065
R10692 DVDD.n5113 DVDD.n5112 0.00065
R10693 DVDD.n4695 DVDD.n4694 0.00065
R10694 DVDD.n3070 DVDD.n206 0.00065
R10695 DVDD.n3062 DVDD.n210 0.00065
R10696 DVDD.n3501 DVDD.n3486 0.00065
R10697 DVDD.n3089 DVDD.n3087 0.00065
R10698 DVDD.n3112 DVDD.n3111 0.00065
R10699 DVDD.n3189 DVDD.n3188 0.00065
R10700 DVDD.n724 DVDD.n717 0.00065
R10701 DVDD.n5342 DVDD.n5341 0.00065
R10702 DVDD.n4874 DVDD.n3139 0.00059
R10703 DVDD.n3134 DVDD.n177 0.00059
R10704 DVDD.n5137 DVDD.n4933 0.00059
R10705 DVDD.n4717 DVDD.n3363 0.00059
R10706 DVDD.n4737 DVDD.n4736 0.00059
R10707 DVDD.n3045 DVDD.n3044 0.00059
R10708 DVDD.n4851 DVDD.n4850 0.00059
R10709 DVDD.n4809 DVDD.n4808 0.00059
R10710 DVDD.n5718 DVDD.n5717 0.00059
R10711 DVDD.n3233 DVDD.n3232 0.00059
R10712 DVDD.n3225 DVDD.n3211 0.00059
R10713 DVDD.n706 DVDD.n701 0.00059
R10714 DVDD DVDD.n2294 0.00058
R10715 DVDD.n1347 DVDD 0.00058
R10716 DVDD.n2257 DVDD 0.00058
R10717 DVDD DVDD.n1650 0.00058
R10718 DVDD DVDD.n5410 0.00058
R10719 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n246 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.t71 273.524
R10720 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.t71 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n245 273.524
R10721 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n227 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.t65 273.524
R10722 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.t65 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n226 273.524
R10723 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.t37 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n112 273.524
R10724 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n113 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.t37 273.524
R10725 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n131 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.t19 273.524
R10726 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.t19 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n130 273.524
R10727 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n151 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.t67 273.524
R10728 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.t67 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n150 273.524
R10729 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.t64 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n168 273.524
R10730 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n169 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.t64 273.524
R10731 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.t20 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n189 273.524
R10732 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n190 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.t20 273.524
R10733 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n208 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.t87 273.524
R10734 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.t87 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n207 273.524
R10735 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n226 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.t38 263.844
R10736 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n227 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.t38 263.844
R10737 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n225 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.t56 263.844
R10738 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n228 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.t56 263.844
R10739 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n224 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.t28 263.844
R10740 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n229 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.t28 263.844
R10741 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n223 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.t73 263.844
R10742 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n230 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.t73 263.844
R10743 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n222 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.t23 263.844
R10744 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n231 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.t23 263.844
R10745 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n221 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.t63 263.844
R10746 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n232 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.t63 263.844
R10747 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n220 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.t93 263.844
R10748 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n233 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.t93 263.844
R10749 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n219 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.t49 263.844
R10750 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n234 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.t49 263.844
R10751 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.t91 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n218 263.844
R10752 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n235 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.t91 263.844
R10753 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n254 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.t42 263.844
R10754 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n237 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.t42 263.844
R10755 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n253 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.t81 263.844
R10756 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n238 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.t81 263.844
R10757 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n252 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.t33 263.844
R10758 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n239 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.t33 263.844
R10759 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n251 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.t77 263.844
R10760 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n240 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.t77 263.844
R10761 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n250 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.t48 263.844
R10762 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n241 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.t48 263.844
R10763 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n249 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.t62 263.844
R10764 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n242 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.t62 263.844
R10765 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n248 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.t22 263.844
R10766 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n243 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.t22 263.844
R10767 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n247 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.t55 263.844
R10768 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n244 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.t55 263.844
R10769 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n246 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.t95 263.844
R10770 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n245 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.t95 263.844
R10771 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n130 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.t69 263.844
R10772 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n131 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.t69 263.844
R10773 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n129 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.t30 263.844
R10774 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n132 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.t30 263.844
R10775 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n128 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.t53 263.844
R10776 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n133 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.t53 263.844
R10777 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n127 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.t36 263.844
R10778 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n134 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.t36 263.844
R10779 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n126 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.t59 263.844
R10780 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n135 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.t59 263.844
R10781 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n125 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.t46 263.844
R10782 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n136 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.t46 263.844
R10783 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n124 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.t89 263.844
R10784 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n137 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.t89 263.844
R10785 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n123 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.t31 263.844
R10786 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n138 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.t31 263.844
R10787 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n122 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.t96 263.844
R10788 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n139 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.t96 263.844
R10789 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n104 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.t41 263.844
R10790 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n121 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.t41 263.844
R10791 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n105 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.t26 263.844
R10792 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n120 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.t26 263.844
R10793 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n106 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.t47 263.844
R10794 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n119 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.t47 263.844
R10795 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n107 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.t90 263.844
R10796 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n118 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.t90 263.844
R10797 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n108 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.t61 263.844
R10798 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n117 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.t61 263.844
R10799 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n109 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.t21 263.844
R10800 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n116 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.t21 263.844
R10801 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n110 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.t85 263.844
R10802 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n115 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.t85 263.844
R10803 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n111 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.t27 263.844
R10804 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n114 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.t27 263.844
R10805 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n112 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.t72 263.844
R10806 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n113 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.t72 263.844
R10807 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n169 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.t24 263.844
R10808 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n168 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.t24 263.844
R10809 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n170 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.t78 263.844
R10810 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n167 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.t78 263.844
R10811 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n171 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.t34 263.844
R10812 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n166 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.t34 263.844
R10813 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n172 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.t18 263.844
R10814 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n165 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.t18 263.844
R10815 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n173 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.t39 263.844
R10816 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n164 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.t39 263.844
R10817 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n174 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.t86 263.844
R10818 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n163 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.t86 263.844
R10819 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n175 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.t51 263.844
R10820 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n162 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.t51 263.844
R10821 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n176 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.t94 263.844
R10822 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n161 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.t94 263.844
R10823 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n177 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.t58 263.844
R10824 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n160 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.t58 263.844
R10825 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n159 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.t25 263.844
R10826 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n142 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.t25 263.844
R10827 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n158 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.t68 263.844
R10828 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n143 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.t68 263.844
R10829 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n157 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.t29 263.844
R10830 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n144 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.t29 263.844
R10831 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n156 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.t76 263.844
R10832 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n145 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.t76 263.844
R10833 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n155 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.t84 263.844
R10834 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n146 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.t84 263.844
R10835 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n154 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.t43 263.844
R10836 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n147 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.t43 263.844
R10837 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n153 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.t70 263.844
R10838 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n148 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.t70 263.844
R10839 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n152 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.t52 263.844
R10840 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n149 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.t52 263.844
R10841 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n151 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.t80 263.844
R10842 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n150 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.t80 263.844
R10843 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n207 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.t50 263.844
R10844 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n208 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.t50 263.844
R10845 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n206 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.t17 263.844
R10846 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n209 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.t17 263.844
R10847 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n205 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.t57 263.844
R10848 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n210 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.t57 263.844
R10849 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n204 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.t82 263.844
R10850 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n211 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.t82 263.844
R10851 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n203 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.t74 263.844
R10852 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n212 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.t74 263.844
R10853 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n202 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.t92 263.844
R10854 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n213 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.t92 263.844
R10855 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n201 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.t79 263.844
R10856 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n214 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.t79 263.844
R10857 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n200 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.t35 263.844
R10858 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n215 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.t35 263.844
R10859 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n199 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.t66 263.844
R10860 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n216 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.t66 263.844
R10861 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n181 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.t44 263.844
R10862 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n198 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.t44 263.844
R10863 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n182 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.t75 263.844
R10864 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n197 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.t75 263.844
R10865 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n183 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.t54 263.844
R10866 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n196 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.t54 263.844
R10867 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n184 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.t83 263.844
R10868 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n195 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.t83 263.844
R10869 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n185 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.t40 263.844
R10870 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n194 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.t40 263.844
R10871 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n186 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.t88 263.844
R10872 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n193 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.t88 263.844
R10873 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n187 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.t45 263.844
R10874 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n192 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.t45 263.844
R10875 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n188 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.t32 263.844
R10876 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n191 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.t32 263.844
R10877 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n189 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.t60 263.844
R10878 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n190 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.t60 263.844
R10879 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n228 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n227 9.68093
R10880 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n229 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n228 9.68093
R10881 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n230 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n229 9.68093
R10882 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n231 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n230 9.68093
R10883 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n232 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n231 9.68093
R10884 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n233 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n232 9.68093
R10885 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n234 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n233 9.68093
R10886 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n235 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n234 9.68093
R10887 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n238 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n237 9.68093
R10888 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n239 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n238 9.68093
R10889 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n240 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n239 9.68093
R10890 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n241 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n240 9.68093
R10891 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n242 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n241 9.68093
R10892 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n243 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n242 9.68093
R10893 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n244 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n243 9.68093
R10894 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n245 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n244 9.68093
R10895 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n226 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n225 9.68093
R10896 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n225 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n224 9.68093
R10897 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n224 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n223 9.68093
R10898 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n223 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n222 9.68093
R10899 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n222 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n221 9.68093
R10900 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n221 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n220 9.68093
R10901 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n220 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n219 9.68093
R10902 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n219 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n218 9.68093
R10903 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n254 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n253 9.68093
R10904 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n253 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n252 9.68093
R10905 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n252 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n251 9.68093
R10906 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n251 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n250 9.68093
R10907 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n250 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n249 9.68093
R10908 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n249 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n248 9.68093
R10909 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n248 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n247 9.68093
R10910 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n247 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n246 9.68093
R10911 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n114 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n113 9.68093
R10912 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n115 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n114 9.68093
R10913 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n116 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n115 9.68093
R10914 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n117 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n116 9.68093
R10915 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n118 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n117 9.68093
R10916 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n119 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n118 9.68093
R10917 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n120 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n119 9.68093
R10918 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n121 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n120 9.68093
R10919 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n139 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n138 9.68093
R10920 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n138 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n137 9.68093
R10921 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n137 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n136 9.68093
R10922 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n136 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n135 9.68093
R10923 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n135 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n134 9.68093
R10924 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n134 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n133 9.68093
R10925 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n133 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n132 9.68093
R10926 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n132 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n131 9.68093
R10927 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n112 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n111 9.68093
R10928 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n111 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n110 9.68093
R10929 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n110 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n109 9.68093
R10930 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n109 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n108 9.68093
R10931 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n108 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n107 9.68093
R10932 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n107 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n106 9.68093
R10933 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n106 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n105 9.68093
R10934 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n105 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n104 9.68093
R10935 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n123 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n122 9.68093
R10936 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n124 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n123 9.68093
R10937 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n125 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n124 9.68093
R10938 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n126 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n125 9.68093
R10939 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n127 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n126 9.68093
R10940 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n128 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n127 9.68093
R10941 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n129 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n128 9.68093
R10942 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n130 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n129 9.68093
R10943 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n150 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n149 9.68093
R10944 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n149 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n148 9.68093
R10945 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n148 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n147 9.68093
R10946 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n147 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n146 9.68093
R10947 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n146 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n145 9.68093
R10948 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n145 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n144 9.68093
R10949 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n144 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n143 9.68093
R10950 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n143 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n142 9.68093
R10951 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n161 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n160 9.68093
R10952 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n162 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n161 9.68093
R10953 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n163 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n162 9.68093
R10954 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n164 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n163 9.68093
R10955 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n165 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n164 9.68093
R10956 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n166 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n165 9.68093
R10957 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n167 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n166 9.68093
R10958 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n168 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n167 9.68093
R10959 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n152 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n151 9.68093
R10960 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n153 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n152 9.68093
R10961 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n154 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n153 9.68093
R10962 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n155 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n154 9.68093
R10963 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n156 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n155 9.68093
R10964 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n157 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n156 9.68093
R10965 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n158 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n157 9.68093
R10966 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n159 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n158 9.68093
R10967 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n177 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n176 9.68093
R10968 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n176 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n175 9.68093
R10969 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n175 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n174 9.68093
R10970 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n174 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n173 9.68093
R10971 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n173 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n172 9.68093
R10972 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n172 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n171 9.68093
R10973 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n171 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n170 9.68093
R10974 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n170 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n169 9.68093
R10975 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n191 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n190 9.68093
R10976 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n192 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n191 9.68093
R10977 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n193 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n192 9.68093
R10978 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n194 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n193 9.68093
R10979 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n195 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n194 9.68093
R10980 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n196 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n195 9.68093
R10981 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n197 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n196 9.68093
R10982 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n198 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n197 9.68093
R10983 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n216 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n215 9.68093
R10984 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n215 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n214 9.68093
R10985 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n214 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n213 9.68093
R10986 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n213 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n212 9.68093
R10987 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n212 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n211 9.68093
R10988 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n211 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n210 9.68093
R10989 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n210 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n209 9.68093
R10990 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n209 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n208 9.68093
R10991 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n189 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n188 9.68093
R10992 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n188 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n187 9.68093
R10993 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n187 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n186 9.68093
R10994 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n186 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n185 9.68093
R10995 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n185 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n184 9.68093
R10996 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n184 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n183 9.68093
R10997 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n183 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n182 9.68093
R10998 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n182 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n181 9.68093
R10999 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n200 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n199 9.68093
R11000 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n201 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n200 9.68093
R11001 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n202 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n201 9.68093
R11002 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n203 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n202 9.68093
R11003 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n204 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n203 9.68093
R11004 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n205 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n204 9.68093
R11005 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n206 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n205 9.68093
R11006 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n207 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n206 9.68093
R11007 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n236 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n235 4.84072
R11008 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n237 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n236 4.84072
R11009 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n7 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n218 4.84072
R11010 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n7 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n254 4.84072
R11011 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n140 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n121 4.84072
R11012 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n140 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n139 4.84072
R11013 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n104 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n103 4.84072
R11014 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n122 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n103 4.84072
R11015 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n142 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n141 4.84072
R11016 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n160 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n141 4.84072
R11017 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n178 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n159 4.84072
R11018 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n178 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n177 4.84072
R11019 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n217 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n198 4.84072
R11020 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n217 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n216 4.84072
R11021 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n181 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n180 4.84072
R11022 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n199 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n180 4.84072
R11023 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n85 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n0 5.09602
R11024 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n1 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n62 5.10883
R11025 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n40 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n4 5.09332
R11026 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n7 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n12 4.98233
R11027 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n257 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n84 4.33869
R11028 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n260 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n91 4.14642
R11029 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n257 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n0 4.13574
R11030 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n17 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n15 0.10684
R11031 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n16 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n14 0.226809
R11032 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n13 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n11 0.226809
R11033 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n12 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n10 1.11398
R11034 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n18 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n89 1.11398
R11035 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n19 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n20 0.534346
R11036 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n21 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n22 0.534346
R11037 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n23 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n24 0.534346
R11038 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n25 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n26 0.534346
R11039 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n27 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n28 0.534346
R11040 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n29 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n30 0.534346
R11041 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n31 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n32 0.534346
R11042 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n33 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n34 0.534346
R11043 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n35 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n36 0.534346
R11044 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n37 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n38 0.534346
R11045 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n39 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n40 0.73001
R11046 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n88 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n87 1.11398
R11047 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n43 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n42 0.534346
R11048 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n45 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n41 0.534346
R11049 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n47 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n44 0.534346
R11050 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n49 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n46 0.534346
R11051 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n51 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n48 0.534346
R11052 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n53 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n50 0.534346
R11053 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n55 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n52 0.534346
R11054 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n57 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n54 0.534346
R11055 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n59 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n56 0.534346
R11056 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n61 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n58 0.534346
R11057 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n62 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n60 0.73001
R11058 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n63 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n86 1.11398
R11059 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n64 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n65 0.534346
R11060 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n66 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n67 0.534346
R11061 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n68 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n69 0.534346
R11062 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n70 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n71 0.534346
R11063 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n72 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n73 0.534346
R11064 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n74 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n75 0.534346
R11065 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n76 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n77 0.534346
R11066 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n78 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n79 0.534346
R11067 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n80 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n81 0.534346
R11068 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n82 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n83 0.534346
R11069 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n84 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n85 0.73001
R11070 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.t12 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.t4 1.8765
R11071 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n91 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.t3 1.29859
R11072 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n90 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.t11 1.29859
R11073 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n92 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.t5 1.29859
R11074 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n95 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.t7 1.29859
R11075 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n94 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.t10 1.29859
R11076 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n96 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.t9 1.29859
R11077 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n97 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.t1 1.29859
R11078 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n98 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.t2 1.29859
R11079 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n99 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.t14 1.29859
R11080 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n259 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n102 1.16318
R11081 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n102 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n257 0.97572
R11082 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n93 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n100 0.931354
R11083 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n101 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.t13 0.912457
R11084 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n261 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.t8 0.912457
R11085 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n260 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n259 0.578395
R11086 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n91 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n90 0.578395
R11087 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n90 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n92 0.578395
R11088 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n92 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n93 0.578395
R11089 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n93 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n95 0.578395
R11090 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n95 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n94 0.578395
R11091 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n94 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n96 0.578395
R11092 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n96 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n97 0.578395
R11093 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n97 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n98 0.578395
R11094 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n98 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n99 0.578395
R11095 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n99 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.t12 0.578395
R11096 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n2 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n1 0.620373
R11097 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n5 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n4 0.630944
R11098 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n63 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n60 0.5045
R11099 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n87 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n39 0.5045
R11100 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n18 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n10 0.5045
R11101 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n259 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n101 0.467486
R11102 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n261 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n260 0.467486
R11103 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n102 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n258 0.467055
R11104 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n100 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.t15 0.3645
R11105 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n100 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.t0 0.3645
R11106 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n258 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.t16 0.3281
R11107 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n258 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.t6 0.3281
R11108 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n17 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n7 6.11209
R11109 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n101 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D 0.149031
R11110 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n261 0.149031
R11111 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n11 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n10 0.229028
R11112 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n256 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n103 0.0821327
R11113 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n179 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n178 0.0821327
R11114 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n255 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n180 0.0821327
R11115 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n83 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n85 0.169667
R11116 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n81 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n83 0.192757
R11117 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n79 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n81 0.192757
R11118 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n77 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n79 0.192757
R11119 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n75 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n77 0.192757
R11120 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n75 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n256 0.0723285
R11121 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n73 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n256 0.120928
R11122 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n71 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n73 0.192757
R11123 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n69 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n71 0.192757
R11124 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n67 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n69 0.192757
R11125 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n65 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n67 0.192757
R11126 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n65 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n86 0.145469
R11127 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n2 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n0 0.188574
R11128 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n3 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n2 0.150067
R11129 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n3 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n140 0.191209
R11130 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n86 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n3 5.29016
R11131 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n61 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n62 0.169667
R11132 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n59 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n61 0.192757
R11133 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n57 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n59 0.192757
R11134 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n55 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n57 0.192757
R11135 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n53 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n55 0.192757
R11136 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n179 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n53 0.0723285
R11137 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n51 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n179 0.120928
R11138 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n49 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n51 0.192757
R11139 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n47 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n49 0.192757
R11140 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n45 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n47 0.192757
R11141 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n43 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n45 0.192757
R11142 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n88 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n43 0.145469
R11143 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n5 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n1 0.221781
R11144 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n6 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n5 0.102099
R11145 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n6 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n141 0.168375
R11146 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n88 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n6 5.31608
R11147 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n38 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n40 0.169667
R11148 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n36 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n38 0.192757
R11149 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n34 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n36 0.192757
R11150 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n32 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n34 0.192757
R11151 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n30 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n32 0.192757
R11152 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n30 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n255 0.0723285
R11153 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n28 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n255 0.120928
R11154 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n26 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n28 0.192757
R11155 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n24 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n26 0.192757
R11156 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n22 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n24 0.192757
R11157 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n20 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n22 0.192757
R11158 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n20 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n89 0.145469
R11159 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n8 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n7 1.04643
R11160 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n16 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n13 0.385014
R11161 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n16 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n15 0.24315
R11162 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n84 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n82 0.1949
R11163 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n82 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n80 0.1949
R11164 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n80 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n78 0.1949
R11165 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n78 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n76 0.1949
R11166 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n76 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n74 0.1949
R11167 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n74 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n72 0.1949
R11168 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n72 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n70 0.1949
R11169 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n70 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n68 0.1949
R11170 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n68 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n66 0.1949
R11171 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n66 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n64 0.1949
R11172 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n64 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n63 0.1949
R11173 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n58 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n60 0.1949
R11174 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n56 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n58 0.1949
R11175 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n54 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n56 0.1949
R11176 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n52 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n54 0.1949
R11177 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n50 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n52 0.1949
R11178 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n48 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n50 0.1949
R11179 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n46 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n48 0.1949
R11180 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n44 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n46 0.1949
R11181 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n41 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n44 0.1949
R11182 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n42 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n41 0.1949
R11183 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n87 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n42 0.1949
R11184 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n39 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n37 0.1949
R11185 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n37 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n35 0.1949
R11186 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n35 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n33 0.1949
R11187 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n33 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n31 0.1949
R11188 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n31 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n29 0.1949
R11189 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n29 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n27 0.1949
R11190 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n27 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n25 0.1949
R11191 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n25 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n23 0.1949
R11192 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n23 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n21 0.1949
R11193 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n21 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n19 0.1949
R11194 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n19 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n18 0.1949
R11195 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n14 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n11 0.360357
R11196 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n17 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n14 0.482631
R11197 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n13 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n12 0.337726
R11198 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n236 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n15 0.155273
R11199 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n8 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n4 0.188574
R11200 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n9 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n8 0.150067
R11201 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n9 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n217 0.191209
R11202 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n89 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n9 5.29016
R11203 DVSS.n19912 DVSS.n19911 72044.1
R11204 DVSS.n21442 DVSS.n21441 69584.8
R11205 DVSS.n21442 DVSS.n13369 69568.8
R11206 DVSS.n19912 DVSS.n14849 20790.2
R11207 DVSS.n19911 DVSS.n19910 20768.4
R11208 DVSS.n21441 DVSS.n13370 16041.3
R11209 DVSS.n19907 DVSS.n13369 16041.3
R11210 DVSS.n18159 DVSS.n15142 4180.28
R11211 DVSS.n18160 DVSS.n15143 4158.32
R11212 DVSS.n19911 DVSS.n18529 3646.5
R11213 DVSS.n19913 DVSS.n19912 3646.5
R11214 DVSS.n17484 DVSS.t190 3372.16
R11215 DVSS.n17525 DVSS.t190 3372.16
R11216 DVSS.n18529 DVSS.n15143 3351.4
R11217 DVSS.n19913 DVSS.n15142 3351.4
R11218 DVSS.n19201 DVSS.t187 2629.04
R11219 DVSS.n18161 DVSS.n13368 2402.48
R11220 DVSS.n21443 DVSS.n13368 2401.2
R11221 DVSS.n18161 DVSS.n13367 2400.01
R11222 DVSS.n21443 DVSS.n13367 2398.73
R11223 DVSS.n19906 DVSS.n18998 1820
R11224 DVSS.n14848 DVSS.n13370 1467.09
R11225 DVSS.n19908 DVSS.n19907 1467.09
R11226 DVSS.n14849 DVSS.n14848 1270.34
R11227 DVSS.n19909 DVSS.n19908 1270.34
R11228 DVSS.n19178 DVSS.n18998 1093.94
R11229 DVSS.n19204 DVSS.n19180 867.129
R11230 DVSS.t166 DVSS.n19178 846.384
R11231 DVSS.n16488 DVSS.n15143 551.231
R11232 DVSS.n15584 DVSS.n15142 551.231
R11233 DVSS.t187 DVSS.n19180 425.957
R11234 DVSS.t195 DVSS.t166 337.447
R11235 DVSS.t178 DVSS.t185 337.447
R11236 DVSS.t197 DVSS.t162 337.447
R11237 DVSS.t162 DVSS.t180 337.447
R11238 DVSS.t180 DVSS.t182 337.447
R11239 DVSS.t182 DVSS.t176 337.447
R11240 DVSS.t176 DVSS.t164 337.447
R11241 DVSS.t164 DVSS.t170 337.447
R11242 DVSS.t170 DVSS.t172 337.447
R11243 DVSS.n19203 DVSS.n19202 290.19
R11244 DVSS.n19203 DVSS.n19000 266.233
R11245 DVSS.n19905 DVSS.n19000 233.489
R11246 DVSS.n19202 DVSS.n19177 227.811
R11247 DVSS.n19206 DVSS.n19177 201.056
R11248 DVSS.n19596 DVSS.t120 196.893
R11249 DVSS.n22343 DVSS.t52 196.893
R11250 DVSS.n19179 DVSS.t195 192.234
R11251 DVSS.n20474 DVSS.n14849 177.477
R11252 DVSS.n19909 DVSS.n18997 177.222
R11253 DVSS.n19907 DVSS.n19906 177.022
R11254 DVSS.n19201 DVSS.n13370 177.022
R11255 DVSS.t172 DVSS.n19204 175.638
R11256 DVSS.n19205 DVSS.t197 170.107
R11257 DVSS.t156 DVSS.n19595 168.048
R11258 DVSS.n19595 DVSS.t60 168.048
R11259 DVSS.n22231 DVSS.t66 168.048
R11260 DVSS.n22231 DVSS.t154 168.048
R11261 DVSS.n22342 DVSS.t20 168.048
R11262 DVSS.t64 DVSS.n22342 168.048
R11263 DVSS.n19205 DVSS.t178 167.34
R11264 DVSS.n19905 DVSS.n19001 158.357
R11265 DVSS.t185 DVSS.n19179 145.214
R11266 DVSS.n19176 DVSS.n19001 138.911
R11267 DVSS.n16976 DVSS.n16928 130.275
R11268 DVSS.n17485 DVSS.n16976 130.275
R11269 DVSS.n17483 DVSS.n16925 130.275
R11270 DVSS.n17526 DVSS.n16925 130.275
R11271 DVSS.n17484 DVSS.n17053 123.9
R11272 DVSS.n17525 DVSS.n16929 123.9
R11273 DVSS.n17487 DVSS.n17486 75.1538
R11274 DVSS.n17487 DVSS.n16931 75.1538
R11275 DVSS.n17411 DVSS.n17410 75.1538
R11276 DVSS.n17411 DVSS.n16930 75.1538
R11277 DVSS.n17472 DVSS.n17055 75.1538
R11278 DVSS.n17472 DVSS.n16926 75.1538
R11279 DVSS.t120 DVSS.t50 66.3492
R11280 DVSS.t50 DVSS.t140 66.3492
R11281 DVSS.t140 DVSS.t24 66.3492
R11282 DVSS.t24 DVSS.t152 66.3492
R11283 DVSS.t152 DVSS.t72 66.3492
R11284 DVSS.t72 DVSS.t14 66.3492
R11285 DVSS.t14 DVSS.t100 66.3492
R11286 DVSS.t100 DVSS.t142 66.3492
R11287 DVSS.t142 DVSS.t112 66.3492
R11288 DVSS.t112 DVSS.t2 66.3492
R11289 DVSS.t2 DVSS.t132 66.3492
R11290 DVSS.t132 DVSS.t16 66.3492
R11291 DVSS.t16 DVSS.t102 66.3492
R11292 DVSS.t102 DVSS.t76 66.3492
R11293 DVSS.t76 DVSS.t122 66.3492
R11294 DVSS.t122 DVSS.t88 66.3492
R11295 DVSS.t88 DVSS.t134 66.3492
R11296 DVSS.t134 DVSS.t56 66.3492
R11297 DVSS.t56 DVSS.t156 66.3492
R11298 DVSS.t60 DVSS.t34 66.3492
R11299 DVSS.t34 DVSS.t90 66.3492
R11300 DVSS.t90 DVSS.t54 66.3492
R11301 DVSS.t54 DVSS.t108 66.3492
R11302 DVSS.t108 DVSS.t26 66.3492
R11303 DVSS.t26 DVSS.t42 66.3492
R11304 DVSS.t42 DVSS.t136 66.3492
R11305 DVSS.t136 DVSS.t58 66.3492
R11306 DVSS.t58 DVSS.t144 66.3492
R11307 DVSS.t144 DVSS.t78 66.3492
R11308 DVSS.t78 DVSS.t6 66.3492
R11309 DVSS.t6 DVSS.t92 66.3492
R11310 DVSS.t92 DVSS.t22 66.3492
R11311 DVSS.t22 DVSS.t116 66.3492
R11312 DVSS.t116 DVSS.t158 66.3492
R11313 DVSS.t158 DVSS.t126 66.3492
R11314 DVSS.t126 DVSS.t38 66.3492
R11315 DVSS.t38 DVSS.t146 66.3492
R11316 DVSS.t146 DVSS.t66 66.3492
R11317 DVSS.t154 DVSS.t74 66.3492
R11318 DVSS.t74 DVSS.t130 66.3492
R11319 DVSS.t130 DVSS.t104 66.3492
R11320 DVSS.t104 DVSS.t18 66.3492
R11321 DVSS.t18 DVSS.t114 66.3492
R11322 DVSS.t114 DVSS.t28 66.3492
R11323 DVSS.t28 DVSS.t86 66.3492
R11324 DVSS.t86 DVSS.t44 66.3492
R11325 DVSS.t44 DVSS.t106 66.3492
R11326 DVSS.t106 DVSS.t62 66.3492
R11327 DVSS.t62 DVSS.t124 66.3492
R11328 DVSS.t124 DVSS.t36 66.3492
R11329 DVSS.t36 DVSS.t10 66.3492
R11330 DVSS.t10 DVSS.t46 66.3492
R11331 DVSS.t46 DVSS.t30 66.3492
R11332 DVSS.t30 DVSS.t80 66.3492
R11333 DVSS.t80 DVSS.t160 66.3492
R11334 DVSS.t160 DVSS.t94 66.3492
R11335 DVSS.t94 DVSS.t20 66.3492
R11336 DVSS.t118 DVSS.t64 66.3492
R11337 DVSS.t82 DVSS.t118 66.3492
R11338 DVSS.t138 DVSS.t82 66.3492
R11339 DVSS.t48 DVSS.t138 66.3492
R11340 DVSS.t148 DVSS.t48 66.3492
R11341 DVSS.t68 DVSS.t148 66.3492
R11342 DVSS.t8 DVSS.t68 66.3492
R11343 DVSS.t96 DVSS.t8 66.3492
R11344 DVSS.t12 DVSS.t96 66.3492
R11345 DVSS.t110 DVSS.t12 66.3492
R11346 DVSS.t32 DVSS.t110 66.3492
R11347 DVSS.t128 DVSS.t32 66.3492
R11348 DVSS.t40 DVSS.t128 66.3492
R11349 DVSS.t98 DVSS.t40 66.3492
R11350 DVSS.t70 DVSS.t98 66.3492
R11351 DVSS.t150 DVSS.t70 66.3492
R11352 DVSS.t84 DVSS.t150 66.3492
R11353 DVSS.t4 DVSS.t84 66.3492
R11354 DVSS.t52 DVSS.t4 66.3492
R11355 DVSS.n18995 DVSS.n18994 39.3263
R11356 DVSS.n20616 DVSS.n14705 39.3263
R11357 DVSS.n19206 DVSS.n19176 36.5561
R11358 DVSS.n18994 DVSS.n18642 29.1118
R11359 DVSS.n18988 DVSS.n18642 29.1118
R11360 DVSS.n18988 DVSS.n18650 29.1118
R11361 DVSS.n18899 DVSS.n18650 29.1118
R11362 DVSS.n18899 DVSS.n18887 29.1118
R11363 DVSS.n18905 DVSS.n18887 29.1118
R11364 DVSS.n18905 DVSS.n14542 29.1118
R11365 DVSS.n20693 DVSS.n14542 29.1118
R11366 DVSS.n20693 DVSS.n14543 29.1118
R11367 DVSS.n18946 DVSS.n14543 29.1118
R11368 DVSS.n18959 DVSS.n18946 29.1118
R11369 DVSS.n18959 DVSS.n18938 29.1118
R11370 DVSS.n18965 DVSS.n18938 29.1118
R11371 DVSS.n18965 DVSS.n18930 29.1118
R11372 DVSS.n18971 DVSS.n18930 29.1118
R11373 DVSS.n18971 DVSS.n18919 29.1118
R11374 DVSS.n18980 DVSS.n18919 29.1118
R11375 DVSS.n18980 DVSS.n18920 29.1118
R11376 DVSS.n18920 DVSS.n14571 29.1118
R11377 DVSS.n20684 DVSS.n14571 29.1118
R11378 DVSS.n20684 DVSS.n14572 29.1118
R11379 DVSS.n20678 DVSS.n14572 29.1118
R11380 DVSS.n20678 DVSS.n14581 29.1118
R11381 DVSS.n20103 DVSS.n14581 29.1118
R11382 DVSS.n20121 DVSS.n20103 29.1118
R11383 DVSS.n20121 DVSS.n20095 29.1118
R11384 DVSS.n20127 DVSS.n20095 29.1118
R11385 DVSS.n20127 DVSS.n20087 29.1118
R11386 DVSS.n20133 DVSS.n20087 29.1118
R11387 DVSS.n20133 DVSS.n20079 29.1118
R11388 DVSS.n20139 DVSS.n20079 29.1118
R11389 DVSS.n20139 DVSS.n20072 29.1118
R11390 DVSS.n20145 DVSS.n20072 29.1118
R11391 DVSS.n20145 DVSS.n20064 29.1118
R11392 DVSS.n20151 DVSS.n20064 29.1118
R11393 DVSS.n20151 DVSS.n20035 29.1118
R11394 DVSS.n20162 DVSS.n20035 29.1118
R11395 DVSS.n20162 DVSS.n20030 29.1118
R11396 DVSS.n20169 DVSS.n20030 29.1118
R11397 DVSS.n20169 DVSS.n14606 29.1118
R11398 DVSS.n20669 DVSS.n14606 29.1118
R11399 DVSS.n20669 DVSS.n14607 29.1118
R11400 DVSS.n20663 DVSS.n14607 29.1118
R11401 DVSS.n20663 DVSS.n14613 29.1118
R11402 DVSS.n20657 DVSS.n14613 29.1118
R11403 DVSS.n20657 DVSS.n14618 29.1118
R11404 DVSS.n20651 DVSS.n14618 29.1118
R11405 DVSS.n20651 DVSS.n14627 29.1118
R11406 DVSS.n20270 DVSS.n14627 29.1118
R11407 DVSS.n20270 DVSS.n20256 29.1118
R11408 DVSS.n20276 DVSS.n20256 29.1118
R11409 DVSS.n20276 DVSS.n20248 29.1118
R11410 DVSS.n20282 DVSS.n20248 29.1118
R11411 DVSS.n20282 DVSS.n20240 29.1118
R11412 DVSS.n20288 DVSS.n20240 29.1118
R11413 DVSS.n20288 DVSS.n20229 29.1118
R11414 DVSS.n20296 DVSS.n20229 29.1118
R11415 DVSS.n20296 DVSS.n20230 29.1118
R11416 DVSS.n20230 DVSS.n20203 29.1118
R11417 DVSS.n20308 DVSS.n20203 29.1118
R11418 DVSS.n20308 DVSS.n20198 29.1118
R11419 DVSS.n20313 DVSS.n20198 29.1118
R11420 DVSS.n20313 DVSS.n14655 29.1118
R11421 DVSS.n20643 DVSS.n14655 29.1118
R11422 DVSS.n20643 DVSS.n14656 29.1118
R11423 DVSS.n20636 DVSS.n14656 29.1118
R11424 DVSS.n20636 DVSS.n14665 29.1118
R11425 DVSS.n20629 DVSS.n14665 29.1118
R11426 DVSS.n20629 DVSS.n14671 29.1118
R11427 DVSS.n20386 DVSS.n14671 29.1118
R11428 DVSS.n20404 DVSS.n20386 29.1118
R11429 DVSS.n20404 DVSS.n20378 29.1118
R11430 DVSS.n20410 DVSS.n20378 29.1118
R11431 DVSS.n20410 DVSS.n20370 29.1118
R11432 DVSS.n20420 DVSS.n20370 29.1118
R11433 DVSS.n20420 DVSS.n20361 29.1118
R11434 DVSS.n20426 DVSS.n20361 29.1118
R11435 DVSS.n20426 DVSS.n20349 29.1118
R11436 DVSS.n20435 DVSS.n20349 29.1118
R11437 DVSS.n20435 DVSS.n20343 29.1118
R11438 DVSS.n20443 DVSS.n20343 29.1118
R11439 DVSS.n20443 DVSS.n20336 29.1118
R11440 DVSS.n20454 DVSS.n20336 29.1118
R11441 DVSS.n20454 DVSS.n14697 29.1118
R11442 DVSS.n20622 DVSS.n14697 29.1118
R11443 DVSS.n20622 DVSS.n14698 29.1118
R11444 DVSS.n20616 DVSS.n14698 29.1118
R11445 DVSS.n20474 DVSS.n14705 29.1118
R11446 DVSS.n19910 DVSS.n19909 21.9617
R11447 DVSS.n18160 DVSS.n18159 21.96
R11448 DVSS.n16931 DVSS.n16928 7.68902
R11449 DVSS.n17410 DVSS.n16975 7.68902
R11450 DVSS.n17486 DVSS.n16975 7.68902
R11451 DVSS.n17486 DVSS.n17485 7.68902
R11452 DVSS.n16927 DVSS.n16926 7.68902
R11453 DVSS.n16930 DVSS.n16927 7.68902
R11454 DVSS.n17524 DVSS.n16930 7.68902
R11455 DVSS.n17524 DVSS.n16931 7.68902
R11456 DVSS.n17483 DVSS.n17055 7.68902
R11457 DVSS.n17055 DVSS.n17054 7.68902
R11458 DVSS.n17410 DVSS.n17054 7.68902
R11459 DVSS.n17526 DVSS.n16926 7.68902
R11460 DVSS.n20617 DVSS.n14704 5.28481
R11461 DVSS.n20615 DVSS.n14707 5.28481
R11462 DVSS.n20464 DVSS.n14706 5.28481
R11463 DVSS.n18768 DVSS.n18641 5.2005
R11464 DVSS.n18995 DVSS.n18641 5.2005
R11465 DVSS.n18762 DVSS.n18641 5.2005
R11466 DVSS.n18768 DVSS.n18763 5.2005
R11467 DVSS.n18763 DVSS.n18762 5.2005
R11468 DVSS.n18755 DVSS.n18558 5.2005
R11469 DVSS.n18997 DVSS.n18558 5.2005
R11470 DVSS.n18755 DVSS.n18584 5.2005
R11471 DVSS.n18997 DVSS.n18584 5.2005
R11472 DVSS.n18755 DVSS.n18557 5.2005
R11473 DVSS.n18997 DVSS.n18557 5.2005
R11474 DVSS.n18755 DVSS.n18585 5.2005
R11475 DVSS.n18997 DVSS.n18585 5.2005
R11476 DVSS.n18755 DVSS.n18556 5.2005
R11477 DVSS.n18997 DVSS.n18556 5.2005
R11478 DVSS.n18755 DVSS.n18586 5.2005
R11479 DVSS.n18997 DVSS.n18586 5.2005
R11480 DVSS.n18654 DVSS.n18530 5.2005
R11481 DVSS.n18997 DVSS.n18530 5.2005
R11482 DVSS.n18654 DVSS.n18587 5.2005
R11483 DVSS.n14851 DVSS.n14705 5.2005
R11484 DVSS.n14846 DVSS.n14705 5.2005
R11485 DVSS.n14739 DVSS.n14705 5.2005
R11486 DVSS.n20612 DVSS.n14712 5.2005
R11487 DVSS.n14712 DVSS.n14705 5.2005
R11488 DVSS.n20612 DVSS.n14711 5.2005
R11489 DVSS.n14711 DVSS.n14705 5.2005
R11490 DVSS.n20468 DVSS.n14705 5.2005
R11491 DVSS.n20472 DVSS.n20471 5.2005
R11492 DVSS.n20474 DVSS.n20472 5.2005
R11493 DVSS.n20612 DVSS.n14707 5.2005
R11494 DVSS.n14707 DVSS.n14705 5.2005
R11495 DVSS.n20471 DVSS.n14714 5.2005
R11496 DVSS.n20612 DVSS.n14714 5.2005
R11497 DVSS.n14714 DVSS.n14705 5.2005
R11498 DVSS.n20612 DVSS.n14710 5.2005
R11499 DVSS.n14710 DVSS.n14705 5.2005
R11500 DVSS.n20612 DVSS.n20611 5.2005
R11501 DVSS.n20611 DVSS.n14705 5.2005
R11502 DVSS.n20506 DVSS.n14705 5.2005
R11503 DVSS.n21155 DVSS.n21154 4.7928
R11504 DVSS.n19925 DVSS.n19924 4.60071
R11505 DVSS.n18518 DVSS.n18517 4.60071
R11506 DVSS.n15136 DVSS.n15135 4.60071
R11507 DVSS.n18509 DVSS.n18508 4.60071
R11508 DVSS.n21009 DVSS.n21008 4.60071
R11509 DVSS.n13678 DVSS.n13676 4.5005
R11510 DVSS.n13680 DVSS.n13679 4.5005
R11511 DVSS.n21586 DVSS.n869 4.5005
R11512 DVSS.n21586 DVSS.n21577 4.5005
R11513 DVSS.n21586 DVSS.n21585 4.5005
R11514 DVSS.n21586 DVSS.n1176 4.5005
R11515 DVSS.n1313 DVSS.n623 4.5005
R11516 DVSS.n1332 DVSS.n607 4.5005
R11517 DVSS.n21589 DVSS.n21588 4.5005
R11518 DVSS.n21589 DVSS.n1176 4.5005
R11519 DVSS.n20674 DVSS.n13947 4.5005
R11520 DVSS.n14593 DVSS.n13947 4.5005
R11521 DVSS.n14595 DVSS.n13947 4.5005
R11522 DVSS.n14591 DVSS.n13947 4.5005
R11523 DVSS.n14596 DVSS.n13947 4.5005
R11524 DVSS.n14590 DVSS.n13947 4.5005
R11525 DVSS.n14597 DVSS.n13947 4.5005
R11526 DVSS.n14589 DVSS.n13947 4.5005
R11527 DVSS.n14598 DVSS.n13947 4.5005
R11528 DVSS.n14588 DVSS.n13947 4.5005
R11529 DVSS.n14599 DVSS.n13947 4.5005
R11530 DVSS.n14587 DVSS.n13947 4.5005
R11531 DVSS.n14600 DVSS.n13947 4.5005
R11532 DVSS.n14586 DVSS.n13947 4.5005
R11533 DVSS.n14601 DVSS.n13947 4.5005
R11534 DVSS.n20672 DVSS.n13947 4.5005
R11535 DVSS.n20056 DVSS.n20043 4.5005
R11536 DVSS.n20057 DVSS.n20043 4.5005
R11537 DVSS.n20054 DVSS.n20043 4.5005
R11538 DVSS.n20058 DVSS.n20043 4.5005
R11539 DVSS.n20053 DVSS.n20043 4.5005
R11540 DVSS.n20059 DVSS.n20043 4.5005
R11541 DVSS.n20052 DVSS.n20043 4.5005
R11542 DVSS.n20060 DVSS.n20043 4.5005
R11543 DVSS.n20051 DVSS.n20043 4.5005
R11544 DVSS.n20061 DVSS.n20043 4.5005
R11545 DVSS.n20050 DVSS.n20043 4.5005
R11546 DVSS.n20155 DVSS.n20043 4.5005
R11547 DVSS.n20043 DVSS.n20040 4.5005
R11548 DVSS.n20159 DVSS.n20043 4.5005
R11549 DVSS.n20049 DVSS.n20043 4.5005
R11550 DVSS.n20157 DVSS.n20043 4.5005
R11551 DVSS.n20056 DVSS.n20045 4.5005
R11552 DVSS.n20057 DVSS.n20045 4.5005
R11553 DVSS.n20054 DVSS.n20045 4.5005
R11554 DVSS.n20058 DVSS.n20045 4.5005
R11555 DVSS.n20053 DVSS.n20045 4.5005
R11556 DVSS.n20059 DVSS.n20045 4.5005
R11557 DVSS.n20052 DVSS.n20045 4.5005
R11558 DVSS.n20060 DVSS.n20045 4.5005
R11559 DVSS.n20051 DVSS.n20045 4.5005
R11560 DVSS.n20061 DVSS.n20045 4.5005
R11561 DVSS.n20050 DVSS.n20045 4.5005
R11562 DVSS.n20155 DVSS.n20045 4.5005
R11563 DVSS.n20045 DVSS.n20040 4.5005
R11564 DVSS.n20159 DVSS.n20045 4.5005
R11565 DVSS.n20049 DVSS.n20045 4.5005
R11566 DVSS.n20157 DVSS.n20045 4.5005
R11567 DVSS.n20056 DVSS.n20042 4.5005
R11568 DVSS.n20057 DVSS.n20042 4.5005
R11569 DVSS.n20054 DVSS.n20042 4.5005
R11570 DVSS.n20058 DVSS.n20042 4.5005
R11571 DVSS.n20053 DVSS.n20042 4.5005
R11572 DVSS.n20059 DVSS.n20042 4.5005
R11573 DVSS.n20052 DVSS.n20042 4.5005
R11574 DVSS.n20060 DVSS.n20042 4.5005
R11575 DVSS.n20051 DVSS.n20042 4.5005
R11576 DVSS.n20061 DVSS.n20042 4.5005
R11577 DVSS.n20050 DVSS.n20042 4.5005
R11578 DVSS.n20155 DVSS.n20042 4.5005
R11579 DVSS.n20042 DVSS.n20040 4.5005
R11580 DVSS.n20159 DVSS.n20042 4.5005
R11581 DVSS.n20049 DVSS.n20042 4.5005
R11582 DVSS.n20157 DVSS.n20042 4.5005
R11583 DVSS.n20019 DVSS.n14470 4.5005
R11584 DVSS.n20109 DVSS.n14470 4.5005
R11585 DVSS.n20020 DVSS.n14470 4.5005
R11586 DVSS.n20016 DVSS.n14470 4.5005
R11587 DVSS.n20021 DVSS.n14470 4.5005
R11588 DVSS.n20015 DVSS.n14470 4.5005
R11589 DVSS.n20022 DVSS.n14470 4.5005
R11590 DVSS.n20014 DVSS.n14470 4.5005
R11591 DVSS.n20023 DVSS.n14470 4.5005
R11592 DVSS.n20013 DVSS.n14470 4.5005
R11593 DVSS.n20024 DVSS.n14470 4.5005
R11594 DVSS.n20012 DVSS.n14470 4.5005
R11595 DVSS.n20025 DVSS.n14470 4.5005
R11596 DVSS.n20011 DVSS.n14470 4.5005
R11597 DVSS.n20172 DVSS.n14470 4.5005
R11598 DVSS.n20174 DVSS.n14470 4.5005
R11599 DVSS.n20173 DVSS.n20019 4.5005
R11600 DVSS.n20173 DVSS.n20017 4.5005
R11601 DVSS.n20173 DVSS.n20020 4.5005
R11602 DVSS.n20173 DVSS.n20016 4.5005
R11603 DVSS.n20173 DVSS.n20021 4.5005
R11604 DVSS.n20173 DVSS.n20015 4.5005
R11605 DVSS.n20173 DVSS.n20022 4.5005
R11606 DVSS.n20173 DVSS.n20014 4.5005
R11607 DVSS.n20173 DVSS.n20023 4.5005
R11608 DVSS.n20173 DVSS.n20013 4.5005
R11609 DVSS.n20173 DVSS.n20024 4.5005
R11610 DVSS.n20173 DVSS.n20012 4.5005
R11611 DVSS.n20173 DVSS.n20025 4.5005
R11612 DVSS.n20173 DVSS.n20011 4.5005
R11613 DVSS.n20173 DVSS.n20172 4.5005
R11614 DVSS.n20174 DVSS.n20173 4.5005
R11615 DVSS.n20056 DVSS.n20046 4.5005
R11616 DVSS.n20057 DVSS.n20046 4.5005
R11617 DVSS.n20054 DVSS.n20046 4.5005
R11618 DVSS.n20058 DVSS.n20046 4.5005
R11619 DVSS.n20053 DVSS.n20046 4.5005
R11620 DVSS.n20059 DVSS.n20046 4.5005
R11621 DVSS.n20052 DVSS.n20046 4.5005
R11622 DVSS.n20060 DVSS.n20046 4.5005
R11623 DVSS.n20051 DVSS.n20046 4.5005
R11624 DVSS.n20061 DVSS.n20046 4.5005
R11625 DVSS.n20050 DVSS.n20046 4.5005
R11626 DVSS.n20155 DVSS.n20046 4.5005
R11627 DVSS.n20046 DVSS.n20040 4.5005
R11628 DVSS.n20159 DVSS.n20046 4.5005
R11629 DVSS.n20157 DVSS.n20046 4.5005
R11630 DVSS.n20056 DVSS.n20041 4.5005
R11631 DVSS.n20057 DVSS.n20041 4.5005
R11632 DVSS.n20054 DVSS.n20041 4.5005
R11633 DVSS.n20058 DVSS.n20041 4.5005
R11634 DVSS.n20053 DVSS.n20041 4.5005
R11635 DVSS.n20059 DVSS.n20041 4.5005
R11636 DVSS.n20052 DVSS.n20041 4.5005
R11637 DVSS.n20060 DVSS.n20041 4.5005
R11638 DVSS.n20051 DVSS.n20041 4.5005
R11639 DVSS.n20061 DVSS.n20041 4.5005
R11640 DVSS.n20050 DVSS.n20041 4.5005
R11641 DVSS.n20155 DVSS.n20041 4.5005
R11642 DVSS.n20159 DVSS.n20041 4.5005
R11643 DVSS.n20157 DVSS.n20041 4.5005
R11644 DVSS.n20158 DVSS.n20056 4.5005
R11645 DVSS.n20158 DVSS.n20057 4.5005
R11646 DVSS.n20158 DVSS.n20054 4.5005
R11647 DVSS.n20158 DVSS.n20058 4.5005
R11648 DVSS.n20158 DVSS.n20053 4.5005
R11649 DVSS.n20158 DVSS.n20059 4.5005
R11650 DVSS.n20158 DVSS.n20052 4.5005
R11651 DVSS.n20158 DVSS.n20060 4.5005
R11652 DVSS.n20158 DVSS.n20051 4.5005
R11653 DVSS.n20158 DVSS.n20061 4.5005
R11654 DVSS.n20158 DVSS.n20050 4.5005
R11655 DVSS.n20158 DVSS.n20155 4.5005
R11656 DVSS.n20159 DVSS.n20158 4.5005
R11657 DVSS.n20158 DVSS.n20049 4.5005
R11658 DVSS.n20158 DVSS.n20157 4.5005
R11659 DVSS.n20674 DVSS.n20673 4.5005
R11660 DVSS.n20673 DVSS.n14592 4.5005
R11661 DVSS.n20673 DVSS.n14595 4.5005
R11662 DVSS.n20673 DVSS.n14591 4.5005
R11663 DVSS.n20673 DVSS.n14596 4.5005
R11664 DVSS.n20673 DVSS.n14590 4.5005
R11665 DVSS.n20673 DVSS.n14597 4.5005
R11666 DVSS.n20673 DVSS.n14589 4.5005
R11667 DVSS.n20673 DVSS.n14598 4.5005
R11668 DVSS.n20673 DVSS.n14588 4.5005
R11669 DVSS.n20673 DVSS.n14599 4.5005
R11670 DVSS.n20673 DVSS.n14587 4.5005
R11671 DVSS.n20673 DVSS.n14600 4.5005
R11672 DVSS.n20673 DVSS.n14586 4.5005
R11673 DVSS.n20673 DVSS.n14601 4.5005
R11674 DVSS.n20673 DVSS.n20672 4.5005
R11675 DVSS.n17100 DVSS.n17099 4.5005
R11676 DVSS.n17099 DVSS.n17066 4.5005
R11677 DVSS.n17099 DVSS.n17098 4.5005
R11678 DVSS.n17035 DVSS.n15315 4.5005
R11679 DVSS.n17366 DVSS.n17344 4.5005
R11680 DVSS.n17366 DVSS.n16974 4.5005
R11681 DVSS.n17370 DVSS.n17332 4.5005
R11682 DVSS.n17332 DVSS.n16974 4.5005
R11683 DVSS.n17408 DVSS.n17269 4.5005
R11684 DVSS.n17408 DVSS.n17407 4.5005
R11685 DVSS.n17409 DVSS.n17408 4.5005
R11686 DVSS.n17405 DVSS.n17259 4.5005
R11687 DVSS.n17279 DVSS.n17259 4.5005
R11688 DVSS.n17407 DVSS.n17259 4.5005
R11689 DVSS.n17409 DVSS.n17259 4.5005
R11690 DVSS.n17475 DVSS.n17167 4.5005
R11691 DVSS.n17475 DVSS.n17170 4.5005
R11692 DVSS.n17475 DVSS.n17474 4.5005
R11693 DVSS.n17170 DVSS.n17138 4.5005
R11694 DVSS.n17477 DVSS.n17138 4.5005
R11695 DVSS.n17407 DVSS.n17406 4.5005
R11696 DVSS.n17406 DVSS.n17282 4.5005
R11697 DVSS.n17406 DVSS.n17278 4.5005
R11698 DVSS.n17406 DVSS.n17284 4.5005
R11699 DVSS.n17406 DVSS.n17277 4.5005
R11700 DVSS.n17406 DVSS.n17286 4.5005
R11701 DVSS.n17406 DVSS.n17276 4.5005
R11702 DVSS.n17406 DVSS.n17288 4.5005
R11703 DVSS.n17406 DVSS.n17275 4.5005
R11704 DVSS.n17406 DVSS.n17290 4.5005
R11705 DVSS.n17406 DVSS.n17274 4.5005
R11706 DVSS.n17406 DVSS.n17292 4.5005
R11707 DVSS.n17406 DVSS.n17273 4.5005
R11708 DVSS.n17406 DVSS.n17405 4.5005
R11709 DVSS.n17369 DVSS.n17344 4.5005
R11710 DVSS.n17369 DVSS.n17341 4.5005
R11711 DVSS.n17369 DVSS.n17346 4.5005
R11712 DVSS.n17369 DVSS.n17340 4.5005
R11713 DVSS.n17369 DVSS.n17348 4.5005
R11714 DVSS.n17369 DVSS.n17339 4.5005
R11715 DVSS.n17369 DVSS.n17350 4.5005
R11716 DVSS.n17369 DVSS.n17338 4.5005
R11717 DVSS.n17369 DVSS.n17352 4.5005
R11718 DVSS.n17369 DVSS.n17337 4.5005
R11719 DVSS.n17369 DVSS.n17354 4.5005
R11720 DVSS.n17369 DVSS.n17336 4.5005
R11721 DVSS.n17369 DVSS.n17356 4.5005
R11722 DVSS.n17369 DVSS.n17335 4.5005
R11723 DVSS.n17369 DVSS.n17368 4.5005
R11724 DVSS.n17369 DVSS.n17334 4.5005
R11725 DVSS.n17370 DVSS.n17369 4.5005
R11726 DVSS.n17075 DVSS.n17074 4.5005
R11727 DVSS.n17016 DVSS.n15306 4.5005
R11728 DVSS.n17477 DVSS.n16081 4.5005
R11729 DVSS.n17139 DVSS.n16081 4.5005
R11730 DVSS.n17163 DVSS.n16081 4.5005
R11731 DVSS.n17161 DVSS.n16081 4.5005
R11732 DVSS.n17159 DVSS.n16081 4.5005
R11733 DVSS.n17157 DVSS.n16081 4.5005
R11734 DVSS.n17155 DVSS.n16081 4.5005
R11735 DVSS.n17153 DVSS.n16081 4.5005
R11736 DVSS.n17151 DVSS.n16081 4.5005
R11737 DVSS.n17149 DVSS.n16081 4.5005
R11738 DVSS.n17147 DVSS.n16081 4.5005
R11739 DVSS.n17145 DVSS.n16081 4.5005
R11740 DVSS.n17143 DVSS.n16081 4.5005
R11741 DVSS.n17165 DVSS.n16081 4.5005
R11742 DVSS.n17170 DVSS.n16081 4.5005
R11743 DVSS.n17474 DVSS.n16081 4.5005
R11744 DVSS.n16427 DVSS.n16251 4.5005
R11745 DVSS.n16462 DVSS.n16426 4.5005
R11746 DVSS.n16452 DVSS.n16426 4.5005
R11747 DVSS.n16451 DVSS.n16426 4.5005
R11748 DVSS.n16427 DVSS.n16267 4.5005
R11749 DVSS.n16429 DVSS.n16267 4.5005
R11750 DVSS.n16431 DVSS.n16267 4.5005
R11751 DVSS.n16433 DVSS.n16267 4.5005
R11752 DVSS.n16435 DVSS.n16267 4.5005
R11753 DVSS.n16437 DVSS.n16267 4.5005
R11754 DVSS.n16439 DVSS.n16267 4.5005
R11755 DVSS.n16441 DVSS.n16267 4.5005
R11756 DVSS.n16443 DVSS.n16267 4.5005
R11757 DVSS.n16445 DVSS.n16267 4.5005
R11758 DVSS.n16447 DVSS.n16267 4.5005
R11759 DVSS.n16449 DVSS.n16267 4.5005
R11760 DVSS.n16451 DVSS.n16267 4.5005
R11761 DVSS.n16452 DVSS.n16267 4.5005
R11762 DVSS.n16454 DVSS.n16267 4.5005
R11763 DVSS.n16456 DVSS.n16267 4.5005
R11764 DVSS.n16458 DVSS.n16267 4.5005
R11765 DVSS.n16460 DVSS.n16267 4.5005
R11766 DVSS.n16462 DVSS.n16267 4.5005
R11767 DVSS.n13540 DVSS.n13522 4.5005
R11768 DVSS.n13541 DVSS.n13522 4.5005
R11769 DVSS.n13539 DVSS.n13522 4.5005
R11770 DVSS.n13544 DVSS.n13522 4.5005
R11771 DVSS.n13537 DVSS.n13522 4.5005
R11772 DVSS.n13545 DVSS.n13522 4.5005
R11773 DVSS.n13536 DVSS.n13522 4.5005
R11774 DVSS.n13546 DVSS.n13522 4.5005
R11775 DVSS.n13535 DVSS.n13522 4.5005
R11776 DVSS.n21297 DVSS.n13522 4.5005
R11777 DVSS.n21299 DVSS.n13522 4.5005
R11778 DVSS.n13540 DVSS.n13521 4.5005
R11779 DVSS.n13541 DVSS.n13521 4.5005
R11780 DVSS.n13539 DVSS.n13521 4.5005
R11781 DVSS.n13543 DVSS.n13521 4.5005
R11782 DVSS.n13538 DVSS.n13521 4.5005
R11783 DVSS.n13544 DVSS.n13521 4.5005
R11784 DVSS.n13537 DVSS.n13521 4.5005
R11785 DVSS.n13545 DVSS.n13521 4.5005
R11786 DVSS.n13536 DVSS.n13521 4.5005
R11787 DVSS.n13546 DVSS.n13521 4.5005
R11788 DVSS.n13535 DVSS.n13521 4.5005
R11789 DVSS.n13547 DVSS.n13521 4.5005
R11790 DVSS.n21297 DVSS.n13521 4.5005
R11791 DVSS.n21299 DVSS.n13521 4.5005
R11792 DVSS.n13540 DVSS.n13523 4.5005
R11793 DVSS.n13541 DVSS.n13523 4.5005
R11794 DVSS.n13539 DVSS.n13523 4.5005
R11795 DVSS.n13543 DVSS.n13523 4.5005
R11796 DVSS.n13538 DVSS.n13523 4.5005
R11797 DVSS.n13544 DVSS.n13523 4.5005
R11798 DVSS.n13537 DVSS.n13523 4.5005
R11799 DVSS.n13545 DVSS.n13523 4.5005
R11800 DVSS.n13536 DVSS.n13523 4.5005
R11801 DVSS.n13546 DVSS.n13523 4.5005
R11802 DVSS.n13535 DVSS.n13523 4.5005
R11803 DVSS.n13547 DVSS.n13523 4.5005
R11804 DVSS.n21297 DVSS.n13523 4.5005
R11805 DVSS.n21299 DVSS.n13523 4.5005
R11806 DVSS.n13540 DVSS.n13520 4.5005
R11807 DVSS.n13541 DVSS.n13520 4.5005
R11808 DVSS.n13539 DVSS.n13520 4.5005
R11809 DVSS.n13543 DVSS.n13520 4.5005
R11810 DVSS.n13538 DVSS.n13520 4.5005
R11811 DVSS.n13544 DVSS.n13520 4.5005
R11812 DVSS.n13537 DVSS.n13520 4.5005
R11813 DVSS.n13545 DVSS.n13520 4.5005
R11814 DVSS.n13536 DVSS.n13520 4.5005
R11815 DVSS.n13546 DVSS.n13520 4.5005
R11816 DVSS.n13535 DVSS.n13520 4.5005
R11817 DVSS.n13547 DVSS.n13520 4.5005
R11818 DVSS.n21297 DVSS.n13520 4.5005
R11819 DVSS.n21299 DVSS.n13520 4.5005
R11820 DVSS.n13540 DVSS.n13524 4.5005
R11821 DVSS.n13541 DVSS.n13524 4.5005
R11822 DVSS.n13539 DVSS.n13524 4.5005
R11823 DVSS.n13543 DVSS.n13524 4.5005
R11824 DVSS.n13538 DVSS.n13524 4.5005
R11825 DVSS.n13544 DVSS.n13524 4.5005
R11826 DVSS.n13537 DVSS.n13524 4.5005
R11827 DVSS.n13545 DVSS.n13524 4.5005
R11828 DVSS.n13536 DVSS.n13524 4.5005
R11829 DVSS.n13546 DVSS.n13524 4.5005
R11830 DVSS.n13535 DVSS.n13524 4.5005
R11831 DVSS.n13547 DVSS.n13524 4.5005
R11832 DVSS.n21297 DVSS.n13524 4.5005
R11833 DVSS.n21299 DVSS.n13524 4.5005
R11834 DVSS.n13540 DVSS.n13519 4.5005
R11835 DVSS.n13541 DVSS.n13519 4.5005
R11836 DVSS.n13539 DVSS.n13519 4.5005
R11837 DVSS.n13543 DVSS.n13519 4.5005
R11838 DVSS.n13538 DVSS.n13519 4.5005
R11839 DVSS.n13544 DVSS.n13519 4.5005
R11840 DVSS.n13537 DVSS.n13519 4.5005
R11841 DVSS.n13545 DVSS.n13519 4.5005
R11842 DVSS.n13536 DVSS.n13519 4.5005
R11843 DVSS.n13546 DVSS.n13519 4.5005
R11844 DVSS.n13535 DVSS.n13519 4.5005
R11845 DVSS.n13547 DVSS.n13519 4.5005
R11846 DVSS.n21297 DVSS.n13519 4.5005
R11847 DVSS.n21299 DVSS.n13519 4.5005
R11848 DVSS.n13540 DVSS.n13525 4.5005
R11849 DVSS.n13541 DVSS.n13525 4.5005
R11850 DVSS.n13539 DVSS.n13525 4.5005
R11851 DVSS.n13543 DVSS.n13525 4.5005
R11852 DVSS.n13538 DVSS.n13525 4.5005
R11853 DVSS.n13544 DVSS.n13525 4.5005
R11854 DVSS.n13537 DVSS.n13525 4.5005
R11855 DVSS.n13545 DVSS.n13525 4.5005
R11856 DVSS.n13536 DVSS.n13525 4.5005
R11857 DVSS.n13546 DVSS.n13525 4.5005
R11858 DVSS.n13535 DVSS.n13525 4.5005
R11859 DVSS.n13547 DVSS.n13525 4.5005
R11860 DVSS.n21297 DVSS.n13525 4.5005
R11861 DVSS.n21299 DVSS.n13525 4.5005
R11862 DVSS.n13540 DVSS.n13518 4.5005
R11863 DVSS.n13541 DVSS.n13518 4.5005
R11864 DVSS.n13539 DVSS.n13518 4.5005
R11865 DVSS.n13543 DVSS.n13518 4.5005
R11866 DVSS.n13538 DVSS.n13518 4.5005
R11867 DVSS.n13544 DVSS.n13518 4.5005
R11868 DVSS.n13537 DVSS.n13518 4.5005
R11869 DVSS.n13545 DVSS.n13518 4.5005
R11870 DVSS.n13536 DVSS.n13518 4.5005
R11871 DVSS.n13546 DVSS.n13518 4.5005
R11872 DVSS.n13535 DVSS.n13518 4.5005
R11873 DVSS.n13547 DVSS.n13518 4.5005
R11874 DVSS.n21297 DVSS.n13518 4.5005
R11875 DVSS.n21299 DVSS.n13518 4.5005
R11876 DVSS.n13540 DVSS.n13526 4.5005
R11877 DVSS.n13541 DVSS.n13526 4.5005
R11878 DVSS.n13539 DVSS.n13526 4.5005
R11879 DVSS.n13543 DVSS.n13526 4.5005
R11880 DVSS.n13538 DVSS.n13526 4.5005
R11881 DVSS.n13544 DVSS.n13526 4.5005
R11882 DVSS.n13537 DVSS.n13526 4.5005
R11883 DVSS.n13545 DVSS.n13526 4.5005
R11884 DVSS.n13536 DVSS.n13526 4.5005
R11885 DVSS.n13546 DVSS.n13526 4.5005
R11886 DVSS.n13535 DVSS.n13526 4.5005
R11887 DVSS.n13547 DVSS.n13526 4.5005
R11888 DVSS.n21297 DVSS.n13526 4.5005
R11889 DVSS.n21299 DVSS.n13526 4.5005
R11890 DVSS.n13540 DVSS.n13517 4.5005
R11891 DVSS.n13541 DVSS.n13517 4.5005
R11892 DVSS.n13539 DVSS.n13517 4.5005
R11893 DVSS.n13543 DVSS.n13517 4.5005
R11894 DVSS.n13538 DVSS.n13517 4.5005
R11895 DVSS.n13544 DVSS.n13517 4.5005
R11896 DVSS.n13537 DVSS.n13517 4.5005
R11897 DVSS.n13545 DVSS.n13517 4.5005
R11898 DVSS.n13536 DVSS.n13517 4.5005
R11899 DVSS.n13546 DVSS.n13517 4.5005
R11900 DVSS.n13535 DVSS.n13517 4.5005
R11901 DVSS.n13547 DVSS.n13517 4.5005
R11902 DVSS.n21297 DVSS.n13517 4.5005
R11903 DVSS.n21299 DVSS.n13517 4.5005
R11904 DVSS.n21298 DVSS.n13540 4.5005
R11905 DVSS.n21298 DVSS.n13541 4.5005
R11906 DVSS.n21298 DVSS.n13539 4.5005
R11907 DVSS.n21298 DVSS.n13543 4.5005
R11908 DVSS.n21298 DVSS.n13538 4.5005
R11909 DVSS.n21298 DVSS.n13544 4.5005
R11910 DVSS.n21298 DVSS.n13537 4.5005
R11911 DVSS.n21298 DVSS.n13545 4.5005
R11912 DVSS.n21298 DVSS.n13536 4.5005
R11913 DVSS.n21298 DVSS.n13546 4.5005
R11914 DVSS.n21298 DVSS.n13535 4.5005
R11915 DVSS.n21298 DVSS.n13547 4.5005
R11916 DVSS.n21298 DVSS.n21297 4.5005
R11917 DVSS.n21298 DVSS.n13533 4.5005
R11918 DVSS.n21299 DVSS.n21298 4.5005
R11919 DVSS.n21107 DVSS.n21106 4.5005
R11920 DVSS.n21106 DVSS.n13948 4.5005
R11921 DVSS.n21106 DVSS.n13946 4.5005
R11922 DVSS.n21106 DVSS.n13949 4.5005
R11923 DVSS.n21106 DVSS.n13944 4.5005
R11924 DVSS.n21106 DVSS.n13950 4.5005
R11925 DVSS.n21106 DVSS.n13943 4.5005
R11926 DVSS.n21106 DVSS.n13951 4.5005
R11927 DVSS.n21106 DVSS.n13942 4.5005
R11928 DVSS.n21106 DVSS.n13952 4.5005
R11929 DVSS.n21106 DVSS.n21105 4.5005
R11930 DVSS.n13966 DVSS.n13948 4.5005
R11931 DVSS.n13966 DVSS.n13946 4.5005
R11932 DVSS.n13979 DVSS.n13966 4.5005
R11933 DVSS.n13978 DVSS.n13966 4.5005
R11934 DVSS.n13966 DVSS.n13949 4.5005
R11935 DVSS.n13966 DVSS.n13944 4.5005
R11936 DVSS.n13966 DVSS.n13950 4.5005
R11937 DVSS.n13966 DVSS.n13943 4.5005
R11938 DVSS.n13966 DVSS.n13951 4.5005
R11939 DVSS.n13966 DVSS.n13942 4.5005
R11940 DVSS.n21103 DVSS.n13966 4.5005
R11941 DVSS.n13977 DVSS.n13966 4.5005
R11942 DVSS.n13966 DVSS.n13952 4.5005
R11943 DVSS.n21105 DVSS.n13966 4.5005
R11944 DVSS.n13964 DVSS.n13948 4.5005
R11945 DVSS.n13964 DVSS.n13946 4.5005
R11946 DVSS.n13979 DVSS.n13964 4.5005
R11947 DVSS.n13978 DVSS.n13964 4.5005
R11948 DVSS.n13964 DVSS.n13949 4.5005
R11949 DVSS.n13964 DVSS.n13944 4.5005
R11950 DVSS.n13964 DVSS.n13950 4.5005
R11951 DVSS.n13964 DVSS.n13943 4.5005
R11952 DVSS.n13964 DVSS.n13951 4.5005
R11953 DVSS.n13964 DVSS.n13942 4.5005
R11954 DVSS.n21103 DVSS.n13964 4.5005
R11955 DVSS.n13977 DVSS.n13964 4.5005
R11956 DVSS.n13964 DVSS.n13952 4.5005
R11957 DVSS.n21105 DVSS.n13964 4.5005
R11958 DVSS.n13967 DVSS.n13948 4.5005
R11959 DVSS.n13967 DVSS.n13946 4.5005
R11960 DVSS.n13979 DVSS.n13967 4.5005
R11961 DVSS.n13978 DVSS.n13967 4.5005
R11962 DVSS.n13967 DVSS.n13949 4.5005
R11963 DVSS.n13967 DVSS.n13944 4.5005
R11964 DVSS.n13967 DVSS.n13950 4.5005
R11965 DVSS.n13967 DVSS.n13943 4.5005
R11966 DVSS.n13967 DVSS.n13951 4.5005
R11967 DVSS.n13967 DVSS.n13942 4.5005
R11968 DVSS.n21103 DVSS.n13967 4.5005
R11969 DVSS.n13977 DVSS.n13967 4.5005
R11970 DVSS.n13967 DVSS.n13952 4.5005
R11971 DVSS.n21105 DVSS.n13967 4.5005
R11972 DVSS.n13963 DVSS.n13948 4.5005
R11973 DVSS.n13963 DVSS.n13946 4.5005
R11974 DVSS.n13979 DVSS.n13963 4.5005
R11975 DVSS.n13978 DVSS.n13963 4.5005
R11976 DVSS.n13963 DVSS.n13949 4.5005
R11977 DVSS.n13963 DVSS.n13944 4.5005
R11978 DVSS.n13963 DVSS.n13950 4.5005
R11979 DVSS.n13963 DVSS.n13943 4.5005
R11980 DVSS.n13963 DVSS.n13951 4.5005
R11981 DVSS.n13963 DVSS.n13942 4.5005
R11982 DVSS.n21103 DVSS.n13963 4.5005
R11983 DVSS.n13977 DVSS.n13963 4.5005
R11984 DVSS.n13963 DVSS.n13952 4.5005
R11985 DVSS.n21105 DVSS.n13963 4.5005
R11986 DVSS.n13968 DVSS.n13948 4.5005
R11987 DVSS.n13968 DVSS.n13946 4.5005
R11988 DVSS.n13979 DVSS.n13968 4.5005
R11989 DVSS.n13978 DVSS.n13968 4.5005
R11990 DVSS.n13968 DVSS.n13949 4.5005
R11991 DVSS.n13968 DVSS.n13944 4.5005
R11992 DVSS.n13968 DVSS.n13950 4.5005
R11993 DVSS.n13968 DVSS.n13943 4.5005
R11994 DVSS.n13968 DVSS.n13951 4.5005
R11995 DVSS.n13968 DVSS.n13942 4.5005
R11996 DVSS.n21103 DVSS.n13968 4.5005
R11997 DVSS.n13977 DVSS.n13968 4.5005
R11998 DVSS.n13968 DVSS.n13952 4.5005
R11999 DVSS.n21105 DVSS.n13968 4.5005
R12000 DVSS.n13962 DVSS.n13948 4.5005
R12001 DVSS.n13962 DVSS.n13946 4.5005
R12002 DVSS.n13979 DVSS.n13962 4.5005
R12003 DVSS.n13978 DVSS.n13962 4.5005
R12004 DVSS.n13962 DVSS.n13949 4.5005
R12005 DVSS.n13962 DVSS.n13944 4.5005
R12006 DVSS.n13962 DVSS.n13950 4.5005
R12007 DVSS.n13962 DVSS.n13943 4.5005
R12008 DVSS.n13962 DVSS.n13951 4.5005
R12009 DVSS.n13962 DVSS.n13942 4.5005
R12010 DVSS.n21103 DVSS.n13962 4.5005
R12011 DVSS.n13977 DVSS.n13962 4.5005
R12012 DVSS.n13962 DVSS.n13952 4.5005
R12013 DVSS.n21105 DVSS.n13962 4.5005
R12014 DVSS.n13969 DVSS.n13948 4.5005
R12015 DVSS.n13969 DVSS.n13946 4.5005
R12016 DVSS.n13979 DVSS.n13969 4.5005
R12017 DVSS.n13978 DVSS.n13969 4.5005
R12018 DVSS.n13969 DVSS.n13949 4.5005
R12019 DVSS.n13969 DVSS.n13944 4.5005
R12020 DVSS.n13969 DVSS.n13950 4.5005
R12021 DVSS.n13969 DVSS.n13943 4.5005
R12022 DVSS.n13969 DVSS.n13951 4.5005
R12023 DVSS.n13969 DVSS.n13942 4.5005
R12024 DVSS.n21103 DVSS.n13969 4.5005
R12025 DVSS.n13977 DVSS.n13969 4.5005
R12026 DVSS.n13969 DVSS.n13952 4.5005
R12027 DVSS.n21105 DVSS.n13969 4.5005
R12028 DVSS.n13961 DVSS.n13948 4.5005
R12029 DVSS.n13961 DVSS.n13946 4.5005
R12030 DVSS.n13979 DVSS.n13961 4.5005
R12031 DVSS.n13978 DVSS.n13961 4.5005
R12032 DVSS.n13961 DVSS.n13949 4.5005
R12033 DVSS.n13961 DVSS.n13944 4.5005
R12034 DVSS.n13961 DVSS.n13950 4.5005
R12035 DVSS.n13961 DVSS.n13943 4.5005
R12036 DVSS.n13961 DVSS.n13951 4.5005
R12037 DVSS.n13961 DVSS.n13942 4.5005
R12038 DVSS.n21103 DVSS.n13961 4.5005
R12039 DVSS.n13977 DVSS.n13961 4.5005
R12040 DVSS.n13961 DVSS.n13952 4.5005
R12041 DVSS.n21105 DVSS.n13961 4.5005
R12042 DVSS.n13970 DVSS.n13948 4.5005
R12043 DVSS.n13970 DVSS.n13946 4.5005
R12044 DVSS.n13979 DVSS.n13970 4.5005
R12045 DVSS.n13978 DVSS.n13970 4.5005
R12046 DVSS.n13970 DVSS.n13949 4.5005
R12047 DVSS.n13970 DVSS.n13944 4.5005
R12048 DVSS.n13970 DVSS.n13950 4.5005
R12049 DVSS.n13970 DVSS.n13943 4.5005
R12050 DVSS.n13970 DVSS.n13951 4.5005
R12051 DVSS.n13970 DVSS.n13942 4.5005
R12052 DVSS.n21103 DVSS.n13970 4.5005
R12053 DVSS.n13977 DVSS.n13970 4.5005
R12054 DVSS.n13970 DVSS.n13952 4.5005
R12055 DVSS.n21105 DVSS.n13970 4.5005
R12056 DVSS.n13960 DVSS.n13948 4.5005
R12057 DVSS.n13960 DVSS.n13946 4.5005
R12058 DVSS.n13979 DVSS.n13960 4.5005
R12059 DVSS.n13978 DVSS.n13960 4.5005
R12060 DVSS.n13960 DVSS.n13949 4.5005
R12061 DVSS.n13960 DVSS.n13944 4.5005
R12062 DVSS.n13960 DVSS.n13950 4.5005
R12063 DVSS.n13960 DVSS.n13943 4.5005
R12064 DVSS.n13960 DVSS.n13951 4.5005
R12065 DVSS.n13960 DVSS.n13942 4.5005
R12066 DVSS.n21103 DVSS.n13960 4.5005
R12067 DVSS.n13977 DVSS.n13960 4.5005
R12068 DVSS.n13960 DVSS.n13952 4.5005
R12069 DVSS.n21105 DVSS.n13960 4.5005
R12070 DVSS.n13971 DVSS.n13948 4.5005
R12071 DVSS.n13971 DVSS.n13946 4.5005
R12072 DVSS.n13979 DVSS.n13971 4.5005
R12073 DVSS.n13978 DVSS.n13971 4.5005
R12074 DVSS.n13971 DVSS.n13949 4.5005
R12075 DVSS.n13971 DVSS.n13944 4.5005
R12076 DVSS.n13971 DVSS.n13950 4.5005
R12077 DVSS.n13971 DVSS.n13943 4.5005
R12078 DVSS.n13971 DVSS.n13951 4.5005
R12079 DVSS.n13971 DVSS.n13942 4.5005
R12080 DVSS.n21103 DVSS.n13971 4.5005
R12081 DVSS.n13977 DVSS.n13971 4.5005
R12082 DVSS.n13971 DVSS.n13952 4.5005
R12083 DVSS.n21105 DVSS.n13971 4.5005
R12084 DVSS.n13959 DVSS.n13948 4.5005
R12085 DVSS.n13959 DVSS.n13946 4.5005
R12086 DVSS.n13979 DVSS.n13959 4.5005
R12087 DVSS.n13978 DVSS.n13959 4.5005
R12088 DVSS.n13959 DVSS.n13949 4.5005
R12089 DVSS.n13959 DVSS.n13944 4.5005
R12090 DVSS.n13959 DVSS.n13950 4.5005
R12091 DVSS.n13959 DVSS.n13943 4.5005
R12092 DVSS.n13959 DVSS.n13951 4.5005
R12093 DVSS.n13959 DVSS.n13942 4.5005
R12094 DVSS.n21103 DVSS.n13959 4.5005
R12095 DVSS.n13977 DVSS.n13959 4.5005
R12096 DVSS.n13959 DVSS.n13952 4.5005
R12097 DVSS.n21105 DVSS.n13959 4.5005
R12098 DVSS.n13972 DVSS.n13948 4.5005
R12099 DVSS.n13972 DVSS.n13946 4.5005
R12100 DVSS.n13979 DVSS.n13972 4.5005
R12101 DVSS.n13978 DVSS.n13972 4.5005
R12102 DVSS.n13972 DVSS.n13949 4.5005
R12103 DVSS.n13972 DVSS.n13944 4.5005
R12104 DVSS.n13972 DVSS.n13950 4.5005
R12105 DVSS.n13972 DVSS.n13943 4.5005
R12106 DVSS.n13972 DVSS.n13951 4.5005
R12107 DVSS.n13972 DVSS.n13942 4.5005
R12108 DVSS.n21103 DVSS.n13972 4.5005
R12109 DVSS.n13977 DVSS.n13972 4.5005
R12110 DVSS.n13972 DVSS.n13952 4.5005
R12111 DVSS.n21105 DVSS.n13972 4.5005
R12112 DVSS.n13958 DVSS.n13948 4.5005
R12113 DVSS.n13958 DVSS.n13946 4.5005
R12114 DVSS.n13979 DVSS.n13958 4.5005
R12115 DVSS.n13978 DVSS.n13958 4.5005
R12116 DVSS.n13958 DVSS.n13949 4.5005
R12117 DVSS.n13958 DVSS.n13944 4.5005
R12118 DVSS.n13958 DVSS.n13950 4.5005
R12119 DVSS.n13958 DVSS.n13943 4.5005
R12120 DVSS.n13958 DVSS.n13951 4.5005
R12121 DVSS.n13958 DVSS.n13942 4.5005
R12122 DVSS.n21103 DVSS.n13958 4.5005
R12123 DVSS.n13977 DVSS.n13958 4.5005
R12124 DVSS.n13958 DVSS.n13952 4.5005
R12125 DVSS.n21105 DVSS.n13958 4.5005
R12126 DVSS.n13973 DVSS.n13948 4.5005
R12127 DVSS.n13973 DVSS.n13946 4.5005
R12128 DVSS.n13979 DVSS.n13973 4.5005
R12129 DVSS.n13978 DVSS.n13973 4.5005
R12130 DVSS.n13973 DVSS.n13949 4.5005
R12131 DVSS.n13973 DVSS.n13944 4.5005
R12132 DVSS.n13973 DVSS.n13950 4.5005
R12133 DVSS.n13973 DVSS.n13943 4.5005
R12134 DVSS.n13973 DVSS.n13951 4.5005
R12135 DVSS.n13973 DVSS.n13942 4.5005
R12136 DVSS.n21103 DVSS.n13973 4.5005
R12137 DVSS.n13977 DVSS.n13973 4.5005
R12138 DVSS.n13973 DVSS.n13952 4.5005
R12139 DVSS.n21105 DVSS.n13973 4.5005
R12140 DVSS.n13957 DVSS.n13948 4.5005
R12141 DVSS.n13957 DVSS.n13946 4.5005
R12142 DVSS.n13979 DVSS.n13957 4.5005
R12143 DVSS.n13978 DVSS.n13957 4.5005
R12144 DVSS.n13957 DVSS.n13949 4.5005
R12145 DVSS.n13957 DVSS.n13944 4.5005
R12146 DVSS.n13957 DVSS.n13950 4.5005
R12147 DVSS.n13957 DVSS.n13943 4.5005
R12148 DVSS.n13957 DVSS.n13951 4.5005
R12149 DVSS.n13957 DVSS.n13942 4.5005
R12150 DVSS.n21103 DVSS.n13957 4.5005
R12151 DVSS.n13977 DVSS.n13957 4.5005
R12152 DVSS.n13957 DVSS.n13952 4.5005
R12153 DVSS.n21105 DVSS.n13957 4.5005
R12154 DVSS.n13974 DVSS.n13948 4.5005
R12155 DVSS.n13974 DVSS.n13946 4.5005
R12156 DVSS.n13979 DVSS.n13974 4.5005
R12157 DVSS.n13978 DVSS.n13974 4.5005
R12158 DVSS.n13974 DVSS.n13949 4.5005
R12159 DVSS.n13974 DVSS.n13944 4.5005
R12160 DVSS.n13974 DVSS.n13950 4.5005
R12161 DVSS.n13974 DVSS.n13943 4.5005
R12162 DVSS.n13974 DVSS.n13951 4.5005
R12163 DVSS.n13974 DVSS.n13942 4.5005
R12164 DVSS.n21103 DVSS.n13974 4.5005
R12165 DVSS.n13977 DVSS.n13974 4.5005
R12166 DVSS.n13974 DVSS.n13952 4.5005
R12167 DVSS.n21105 DVSS.n13974 4.5005
R12168 DVSS.n13956 DVSS.n13948 4.5005
R12169 DVSS.n13956 DVSS.n13946 4.5005
R12170 DVSS.n13979 DVSS.n13956 4.5005
R12171 DVSS.n13978 DVSS.n13956 4.5005
R12172 DVSS.n13956 DVSS.n13949 4.5005
R12173 DVSS.n13956 DVSS.n13944 4.5005
R12174 DVSS.n13956 DVSS.n13950 4.5005
R12175 DVSS.n13956 DVSS.n13943 4.5005
R12176 DVSS.n13956 DVSS.n13951 4.5005
R12177 DVSS.n13956 DVSS.n13942 4.5005
R12178 DVSS.n21103 DVSS.n13956 4.5005
R12179 DVSS.n13977 DVSS.n13956 4.5005
R12180 DVSS.n13956 DVSS.n13952 4.5005
R12181 DVSS.n21105 DVSS.n13956 4.5005
R12182 DVSS.n13975 DVSS.n13948 4.5005
R12183 DVSS.n13975 DVSS.n13946 4.5005
R12184 DVSS.n13979 DVSS.n13975 4.5005
R12185 DVSS.n13978 DVSS.n13975 4.5005
R12186 DVSS.n13975 DVSS.n13949 4.5005
R12187 DVSS.n13975 DVSS.n13944 4.5005
R12188 DVSS.n13975 DVSS.n13950 4.5005
R12189 DVSS.n13975 DVSS.n13943 4.5005
R12190 DVSS.n13975 DVSS.n13951 4.5005
R12191 DVSS.n13975 DVSS.n13942 4.5005
R12192 DVSS.n21103 DVSS.n13975 4.5005
R12193 DVSS.n13977 DVSS.n13975 4.5005
R12194 DVSS.n13975 DVSS.n13952 4.5005
R12195 DVSS.n21105 DVSS.n13975 4.5005
R12196 DVSS.n13955 DVSS.n13948 4.5005
R12197 DVSS.n13955 DVSS.n13946 4.5005
R12198 DVSS.n13979 DVSS.n13955 4.5005
R12199 DVSS.n13978 DVSS.n13955 4.5005
R12200 DVSS.n13955 DVSS.n13949 4.5005
R12201 DVSS.n13955 DVSS.n13944 4.5005
R12202 DVSS.n13955 DVSS.n13950 4.5005
R12203 DVSS.n13955 DVSS.n13943 4.5005
R12204 DVSS.n13955 DVSS.n13951 4.5005
R12205 DVSS.n13955 DVSS.n13942 4.5005
R12206 DVSS.n21103 DVSS.n13955 4.5005
R12207 DVSS.n13977 DVSS.n13955 4.5005
R12208 DVSS.n13955 DVSS.n13952 4.5005
R12209 DVSS.n21105 DVSS.n13955 4.5005
R12210 DVSS.n21104 DVSS.n13948 4.5005
R12211 DVSS.n21104 DVSS.n13946 4.5005
R12212 DVSS.n21104 DVSS.n13979 4.5005
R12213 DVSS.n21104 DVSS.n13978 4.5005
R12214 DVSS.n21104 DVSS.n13949 4.5005
R12215 DVSS.n21104 DVSS.n13944 4.5005
R12216 DVSS.n21104 DVSS.n13950 4.5005
R12217 DVSS.n21104 DVSS.n13943 4.5005
R12218 DVSS.n21104 DVSS.n13951 4.5005
R12219 DVSS.n21104 DVSS.n13942 4.5005
R12220 DVSS.n21104 DVSS.n21103 4.5005
R12221 DVSS.n21104 DVSS.n13977 4.5005
R12222 DVSS.n21104 DVSS.n13952 4.5005
R12223 DVSS.n21105 DVSS.n21104 4.5005
R12224 DVSS.n13954 DVSS.n13948 4.5005
R12225 DVSS.n13954 DVSS.n13946 4.5005
R12226 DVSS.n13979 DVSS.n13954 4.5005
R12227 DVSS.n13978 DVSS.n13954 4.5005
R12228 DVSS.n13954 DVSS.n13949 4.5005
R12229 DVSS.n13954 DVSS.n13944 4.5005
R12230 DVSS.n13954 DVSS.n13950 4.5005
R12231 DVSS.n13954 DVSS.n13943 4.5005
R12232 DVSS.n13954 DVSS.n13951 4.5005
R12233 DVSS.n13954 DVSS.n13942 4.5005
R12234 DVSS.n21103 DVSS.n13954 4.5005
R12235 DVSS.n13977 DVSS.n13954 4.5005
R12236 DVSS.n13954 DVSS.n13952 4.5005
R12237 DVSS.n21096 DVSS.n13954 4.5005
R12238 DVSS.n21105 DVSS.n13954 4.5005
R12239 DVSS.n21107 DVSS.n13927 4.5005
R12240 DVSS.n13948 DVSS.n13927 4.5005
R12241 DVSS.n13946 DVSS.n13927 4.5005
R12242 DVSS.n13979 DVSS.n13927 4.5005
R12243 DVSS.n13978 DVSS.n13927 4.5005
R12244 DVSS.n13949 DVSS.n13927 4.5005
R12245 DVSS.n13944 DVSS.n13927 4.5005
R12246 DVSS.n13950 DVSS.n13927 4.5005
R12247 DVSS.n13943 DVSS.n13927 4.5005
R12248 DVSS.n13951 DVSS.n13927 4.5005
R12249 DVSS.n13942 DVSS.n13927 4.5005
R12250 DVSS.n21103 DVSS.n13927 4.5005
R12251 DVSS.n13977 DVSS.n13927 4.5005
R12252 DVSS.n13952 DVSS.n13927 4.5005
R12253 DVSS.n21096 DVSS.n13927 4.5005
R12254 DVSS.n21105 DVSS.n13927 4.5005
R12255 DVSS.n20818 DVSS.n14465 4.5005
R12256 DVSS.n14483 DVSS.n14465 4.5005
R12257 DVSS.n14481 DVSS.n14465 4.5005
R12258 DVSS.n14486 DVSS.n14465 4.5005
R12259 DVSS.n14479 DVSS.n14465 4.5005
R12260 DVSS.n14487 DVSS.n14465 4.5005
R12261 DVSS.n14478 DVSS.n14465 4.5005
R12262 DVSS.n14488 DVSS.n14465 4.5005
R12263 DVSS.n14477 DVSS.n14465 4.5005
R12264 DVSS.n20847 DVSS.n14465 4.5005
R12265 DVSS.n14475 DVSS.n14465 4.5005
R12266 DVSS.n20849 DVSS.n14465 4.5005
R12267 DVSS.n20818 DVSS.n14464 4.5005
R12268 DVSS.n14483 DVSS.n14464 4.5005
R12269 DVSS.n14481 DVSS.n14464 4.5005
R12270 DVSS.n14485 DVSS.n14464 4.5005
R12271 DVSS.n14480 DVSS.n14464 4.5005
R12272 DVSS.n14486 DVSS.n14464 4.5005
R12273 DVSS.n14479 DVSS.n14464 4.5005
R12274 DVSS.n14487 DVSS.n14464 4.5005
R12275 DVSS.n14478 DVSS.n14464 4.5005
R12276 DVSS.n14488 DVSS.n14464 4.5005
R12277 DVSS.n14477 DVSS.n14464 4.5005
R12278 DVSS.n14490 DVSS.n14464 4.5005
R12279 DVSS.n14476 DVSS.n14464 4.5005
R12280 DVSS.n20847 DVSS.n14464 4.5005
R12281 DVSS.n14475 DVSS.n14464 4.5005
R12282 DVSS.n20849 DVSS.n14464 4.5005
R12283 DVSS.n20818 DVSS.n14466 4.5005
R12284 DVSS.n14483 DVSS.n14466 4.5005
R12285 DVSS.n14481 DVSS.n14466 4.5005
R12286 DVSS.n14485 DVSS.n14466 4.5005
R12287 DVSS.n14480 DVSS.n14466 4.5005
R12288 DVSS.n14486 DVSS.n14466 4.5005
R12289 DVSS.n14479 DVSS.n14466 4.5005
R12290 DVSS.n14487 DVSS.n14466 4.5005
R12291 DVSS.n14478 DVSS.n14466 4.5005
R12292 DVSS.n14488 DVSS.n14466 4.5005
R12293 DVSS.n14477 DVSS.n14466 4.5005
R12294 DVSS.n14490 DVSS.n14466 4.5005
R12295 DVSS.n14476 DVSS.n14466 4.5005
R12296 DVSS.n20847 DVSS.n14466 4.5005
R12297 DVSS.n20849 DVSS.n14466 4.5005
R12298 DVSS.n14483 DVSS.n14463 4.5005
R12299 DVSS.n14481 DVSS.n14463 4.5005
R12300 DVSS.n14485 DVSS.n14463 4.5005
R12301 DVSS.n14480 DVSS.n14463 4.5005
R12302 DVSS.n14486 DVSS.n14463 4.5005
R12303 DVSS.n14479 DVSS.n14463 4.5005
R12304 DVSS.n14487 DVSS.n14463 4.5005
R12305 DVSS.n14478 DVSS.n14463 4.5005
R12306 DVSS.n14488 DVSS.n14463 4.5005
R12307 DVSS.n14477 DVSS.n14463 4.5005
R12308 DVSS.n14490 DVSS.n14463 4.5005
R12309 DVSS.n14476 DVSS.n14463 4.5005
R12310 DVSS.n20847 DVSS.n14463 4.5005
R12311 DVSS.n20849 DVSS.n14463 4.5005
R12312 DVSS.n14483 DVSS.n14467 4.5005
R12313 DVSS.n14481 DVSS.n14467 4.5005
R12314 DVSS.n14485 DVSS.n14467 4.5005
R12315 DVSS.n14480 DVSS.n14467 4.5005
R12316 DVSS.n14486 DVSS.n14467 4.5005
R12317 DVSS.n14479 DVSS.n14467 4.5005
R12318 DVSS.n14487 DVSS.n14467 4.5005
R12319 DVSS.n14478 DVSS.n14467 4.5005
R12320 DVSS.n14488 DVSS.n14467 4.5005
R12321 DVSS.n14477 DVSS.n14467 4.5005
R12322 DVSS.n14490 DVSS.n14467 4.5005
R12323 DVSS.n14476 DVSS.n14467 4.5005
R12324 DVSS.n20847 DVSS.n14467 4.5005
R12325 DVSS.n20849 DVSS.n14467 4.5005
R12326 DVSS.n14483 DVSS.n14462 4.5005
R12327 DVSS.n14481 DVSS.n14462 4.5005
R12328 DVSS.n14485 DVSS.n14462 4.5005
R12329 DVSS.n14480 DVSS.n14462 4.5005
R12330 DVSS.n14486 DVSS.n14462 4.5005
R12331 DVSS.n14479 DVSS.n14462 4.5005
R12332 DVSS.n14487 DVSS.n14462 4.5005
R12333 DVSS.n14478 DVSS.n14462 4.5005
R12334 DVSS.n14488 DVSS.n14462 4.5005
R12335 DVSS.n14477 DVSS.n14462 4.5005
R12336 DVSS.n14490 DVSS.n14462 4.5005
R12337 DVSS.n14476 DVSS.n14462 4.5005
R12338 DVSS.n20847 DVSS.n14462 4.5005
R12339 DVSS.n20849 DVSS.n14462 4.5005
R12340 DVSS.n14483 DVSS.n14468 4.5005
R12341 DVSS.n14481 DVSS.n14468 4.5005
R12342 DVSS.n14485 DVSS.n14468 4.5005
R12343 DVSS.n14480 DVSS.n14468 4.5005
R12344 DVSS.n14486 DVSS.n14468 4.5005
R12345 DVSS.n14479 DVSS.n14468 4.5005
R12346 DVSS.n14487 DVSS.n14468 4.5005
R12347 DVSS.n14478 DVSS.n14468 4.5005
R12348 DVSS.n14488 DVSS.n14468 4.5005
R12349 DVSS.n14477 DVSS.n14468 4.5005
R12350 DVSS.n14490 DVSS.n14468 4.5005
R12351 DVSS.n14476 DVSS.n14468 4.5005
R12352 DVSS.n20847 DVSS.n14468 4.5005
R12353 DVSS.n20849 DVSS.n14468 4.5005
R12354 DVSS.n14483 DVSS.n14461 4.5005
R12355 DVSS.n14481 DVSS.n14461 4.5005
R12356 DVSS.n14485 DVSS.n14461 4.5005
R12357 DVSS.n14480 DVSS.n14461 4.5005
R12358 DVSS.n14486 DVSS.n14461 4.5005
R12359 DVSS.n14479 DVSS.n14461 4.5005
R12360 DVSS.n14487 DVSS.n14461 4.5005
R12361 DVSS.n14478 DVSS.n14461 4.5005
R12362 DVSS.n14488 DVSS.n14461 4.5005
R12363 DVSS.n14477 DVSS.n14461 4.5005
R12364 DVSS.n14490 DVSS.n14461 4.5005
R12365 DVSS.n14476 DVSS.n14461 4.5005
R12366 DVSS.n20847 DVSS.n14461 4.5005
R12367 DVSS.n20849 DVSS.n14461 4.5005
R12368 DVSS.n14483 DVSS.n14469 4.5005
R12369 DVSS.n14481 DVSS.n14469 4.5005
R12370 DVSS.n14485 DVSS.n14469 4.5005
R12371 DVSS.n14480 DVSS.n14469 4.5005
R12372 DVSS.n14486 DVSS.n14469 4.5005
R12373 DVSS.n14479 DVSS.n14469 4.5005
R12374 DVSS.n14487 DVSS.n14469 4.5005
R12375 DVSS.n14478 DVSS.n14469 4.5005
R12376 DVSS.n14488 DVSS.n14469 4.5005
R12377 DVSS.n14477 DVSS.n14469 4.5005
R12378 DVSS.n14490 DVSS.n14469 4.5005
R12379 DVSS.n14476 DVSS.n14469 4.5005
R12380 DVSS.n20847 DVSS.n14469 4.5005
R12381 DVSS.n20849 DVSS.n14469 4.5005
R12382 DVSS.n14483 DVSS.n14460 4.5005
R12383 DVSS.n14481 DVSS.n14460 4.5005
R12384 DVSS.n14485 DVSS.n14460 4.5005
R12385 DVSS.n14480 DVSS.n14460 4.5005
R12386 DVSS.n14486 DVSS.n14460 4.5005
R12387 DVSS.n14479 DVSS.n14460 4.5005
R12388 DVSS.n14487 DVSS.n14460 4.5005
R12389 DVSS.n14478 DVSS.n14460 4.5005
R12390 DVSS.n14488 DVSS.n14460 4.5005
R12391 DVSS.n14477 DVSS.n14460 4.5005
R12392 DVSS.n14490 DVSS.n14460 4.5005
R12393 DVSS.n14476 DVSS.n14460 4.5005
R12394 DVSS.n20847 DVSS.n14460 4.5005
R12395 DVSS.n20849 DVSS.n14460 4.5005
R12396 DVSS.n20848 DVSS.n14483 4.5005
R12397 DVSS.n20848 DVSS.n14481 4.5005
R12398 DVSS.n20848 DVSS.n14485 4.5005
R12399 DVSS.n20848 DVSS.n14480 4.5005
R12400 DVSS.n20848 DVSS.n14486 4.5005
R12401 DVSS.n20848 DVSS.n14479 4.5005
R12402 DVSS.n20848 DVSS.n14487 4.5005
R12403 DVSS.n20848 DVSS.n14478 4.5005
R12404 DVSS.n20848 DVSS.n14488 4.5005
R12405 DVSS.n20848 DVSS.n14477 4.5005
R12406 DVSS.n20848 DVSS.n14490 4.5005
R12407 DVSS.n20848 DVSS.n14476 4.5005
R12408 DVSS.n20848 DVSS.n20847 4.5005
R12409 DVSS.n20848 DVSS.n14475 4.5005
R12410 DVSS.n20849 DVSS.n20848 4.5005
R12411 DVSS.n20009 DVSS.n14882 4.5005
R12412 DVSS.n20009 DVSS.n14883 4.5005
R12413 DVSS.n20009 DVSS.n14881 4.5005
R12414 DVSS.n20009 DVSS.n14884 4.5005
R12415 DVSS.n20009 DVSS.n14879 4.5005
R12416 DVSS.n20009 DVSS.n14885 4.5005
R12417 DVSS.n20009 DVSS.n14878 4.5005
R12418 DVSS.n20009 DVSS.n14886 4.5005
R12419 DVSS.n20009 DVSS.n14877 4.5005
R12420 DVSS.n20009 DVSS.n14887 4.5005
R12421 DVSS.n20009 DVSS.n20008 4.5005
R12422 DVSS.n14893 DVSS.n14883 4.5005
R12423 DVSS.n14893 DVSS.n14881 4.5005
R12424 DVSS.n14912 DVSS.n14893 4.5005
R12425 DVSS.n14910 DVSS.n14893 4.5005
R12426 DVSS.n14893 DVSS.n14884 4.5005
R12427 DVSS.n14893 DVSS.n14879 4.5005
R12428 DVSS.n14893 DVSS.n14885 4.5005
R12429 DVSS.n14893 DVSS.n14878 4.5005
R12430 DVSS.n14893 DVSS.n14886 4.5005
R12431 DVSS.n14893 DVSS.n14877 4.5005
R12432 DVSS.n20006 DVSS.n14893 4.5005
R12433 DVSS.n14909 DVSS.n14893 4.5005
R12434 DVSS.n14893 DVSS.n14887 4.5005
R12435 DVSS.n20008 DVSS.n14893 4.5005
R12436 DVSS.n14896 DVSS.n14883 4.5005
R12437 DVSS.n14896 DVSS.n14881 4.5005
R12438 DVSS.n14912 DVSS.n14896 4.5005
R12439 DVSS.n14910 DVSS.n14896 4.5005
R12440 DVSS.n14896 DVSS.n14884 4.5005
R12441 DVSS.n14896 DVSS.n14879 4.5005
R12442 DVSS.n14896 DVSS.n14885 4.5005
R12443 DVSS.n14896 DVSS.n14878 4.5005
R12444 DVSS.n14896 DVSS.n14886 4.5005
R12445 DVSS.n14896 DVSS.n14877 4.5005
R12446 DVSS.n20006 DVSS.n14896 4.5005
R12447 DVSS.n14909 DVSS.n14896 4.5005
R12448 DVSS.n14896 DVSS.n14887 4.5005
R12449 DVSS.n20008 DVSS.n14896 4.5005
R12450 DVSS.n14892 DVSS.n14883 4.5005
R12451 DVSS.n14892 DVSS.n14881 4.5005
R12452 DVSS.n14912 DVSS.n14892 4.5005
R12453 DVSS.n14910 DVSS.n14892 4.5005
R12454 DVSS.n14892 DVSS.n14884 4.5005
R12455 DVSS.n14892 DVSS.n14879 4.5005
R12456 DVSS.n14892 DVSS.n14885 4.5005
R12457 DVSS.n14892 DVSS.n14878 4.5005
R12458 DVSS.n14892 DVSS.n14886 4.5005
R12459 DVSS.n14892 DVSS.n14877 4.5005
R12460 DVSS.n20006 DVSS.n14892 4.5005
R12461 DVSS.n14909 DVSS.n14892 4.5005
R12462 DVSS.n14892 DVSS.n14887 4.5005
R12463 DVSS.n20008 DVSS.n14892 4.5005
R12464 DVSS.n14898 DVSS.n14883 4.5005
R12465 DVSS.n14898 DVSS.n14881 4.5005
R12466 DVSS.n14912 DVSS.n14898 4.5005
R12467 DVSS.n14910 DVSS.n14898 4.5005
R12468 DVSS.n14898 DVSS.n14884 4.5005
R12469 DVSS.n14898 DVSS.n14879 4.5005
R12470 DVSS.n14898 DVSS.n14885 4.5005
R12471 DVSS.n14898 DVSS.n14878 4.5005
R12472 DVSS.n14898 DVSS.n14886 4.5005
R12473 DVSS.n14898 DVSS.n14877 4.5005
R12474 DVSS.n20006 DVSS.n14898 4.5005
R12475 DVSS.n14909 DVSS.n14898 4.5005
R12476 DVSS.n14898 DVSS.n14887 4.5005
R12477 DVSS.n20008 DVSS.n14898 4.5005
R12478 DVSS.n14891 DVSS.n14883 4.5005
R12479 DVSS.n14891 DVSS.n14881 4.5005
R12480 DVSS.n14912 DVSS.n14891 4.5005
R12481 DVSS.n14910 DVSS.n14891 4.5005
R12482 DVSS.n14891 DVSS.n14884 4.5005
R12483 DVSS.n14891 DVSS.n14879 4.5005
R12484 DVSS.n14891 DVSS.n14885 4.5005
R12485 DVSS.n14891 DVSS.n14878 4.5005
R12486 DVSS.n14891 DVSS.n14886 4.5005
R12487 DVSS.n14891 DVSS.n14877 4.5005
R12488 DVSS.n20006 DVSS.n14891 4.5005
R12489 DVSS.n14909 DVSS.n14891 4.5005
R12490 DVSS.n14891 DVSS.n14887 4.5005
R12491 DVSS.n20008 DVSS.n14891 4.5005
R12492 DVSS.n14900 DVSS.n14883 4.5005
R12493 DVSS.n14900 DVSS.n14881 4.5005
R12494 DVSS.n14912 DVSS.n14900 4.5005
R12495 DVSS.n14910 DVSS.n14900 4.5005
R12496 DVSS.n14900 DVSS.n14884 4.5005
R12497 DVSS.n14900 DVSS.n14879 4.5005
R12498 DVSS.n14900 DVSS.n14885 4.5005
R12499 DVSS.n14900 DVSS.n14878 4.5005
R12500 DVSS.n14900 DVSS.n14886 4.5005
R12501 DVSS.n14900 DVSS.n14877 4.5005
R12502 DVSS.n20006 DVSS.n14900 4.5005
R12503 DVSS.n14909 DVSS.n14900 4.5005
R12504 DVSS.n14900 DVSS.n14887 4.5005
R12505 DVSS.n20008 DVSS.n14900 4.5005
R12506 DVSS.n14890 DVSS.n14883 4.5005
R12507 DVSS.n14890 DVSS.n14881 4.5005
R12508 DVSS.n14912 DVSS.n14890 4.5005
R12509 DVSS.n14910 DVSS.n14890 4.5005
R12510 DVSS.n14890 DVSS.n14884 4.5005
R12511 DVSS.n14890 DVSS.n14879 4.5005
R12512 DVSS.n14890 DVSS.n14885 4.5005
R12513 DVSS.n14890 DVSS.n14878 4.5005
R12514 DVSS.n14890 DVSS.n14886 4.5005
R12515 DVSS.n14890 DVSS.n14877 4.5005
R12516 DVSS.n20006 DVSS.n14890 4.5005
R12517 DVSS.n14909 DVSS.n14890 4.5005
R12518 DVSS.n14890 DVSS.n14887 4.5005
R12519 DVSS.n20008 DVSS.n14890 4.5005
R12520 DVSS.n14902 DVSS.n14883 4.5005
R12521 DVSS.n14902 DVSS.n14881 4.5005
R12522 DVSS.n14912 DVSS.n14902 4.5005
R12523 DVSS.n14910 DVSS.n14902 4.5005
R12524 DVSS.n14902 DVSS.n14884 4.5005
R12525 DVSS.n14902 DVSS.n14879 4.5005
R12526 DVSS.n14902 DVSS.n14885 4.5005
R12527 DVSS.n14902 DVSS.n14878 4.5005
R12528 DVSS.n14902 DVSS.n14886 4.5005
R12529 DVSS.n14902 DVSS.n14877 4.5005
R12530 DVSS.n20006 DVSS.n14902 4.5005
R12531 DVSS.n14909 DVSS.n14902 4.5005
R12532 DVSS.n14902 DVSS.n14887 4.5005
R12533 DVSS.n20008 DVSS.n14902 4.5005
R12534 DVSS.n14889 DVSS.n14883 4.5005
R12535 DVSS.n14889 DVSS.n14881 4.5005
R12536 DVSS.n14912 DVSS.n14889 4.5005
R12537 DVSS.n14910 DVSS.n14889 4.5005
R12538 DVSS.n14889 DVSS.n14884 4.5005
R12539 DVSS.n14889 DVSS.n14879 4.5005
R12540 DVSS.n14889 DVSS.n14885 4.5005
R12541 DVSS.n14889 DVSS.n14878 4.5005
R12542 DVSS.n14889 DVSS.n14886 4.5005
R12543 DVSS.n14889 DVSS.n14877 4.5005
R12544 DVSS.n20006 DVSS.n14889 4.5005
R12545 DVSS.n14909 DVSS.n14889 4.5005
R12546 DVSS.n14889 DVSS.n14887 4.5005
R12547 DVSS.n20008 DVSS.n14889 4.5005
R12548 DVSS.n20007 DVSS.n14883 4.5005
R12549 DVSS.n20007 DVSS.n14881 4.5005
R12550 DVSS.n20007 DVSS.n14912 4.5005
R12551 DVSS.n20007 DVSS.n14910 4.5005
R12552 DVSS.n20007 DVSS.n14884 4.5005
R12553 DVSS.n20007 DVSS.n14879 4.5005
R12554 DVSS.n20007 DVSS.n14885 4.5005
R12555 DVSS.n20007 DVSS.n14878 4.5005
R12556 DVSS.n20007 DVSS.n14886 4.5005
R12557 DVSS.n20007 DVSS.n14877 4.5005
R12558 DVSS.n20007 DVSS.n20006 4.5005
R12559 DVSS.n20007 DVSS.n14909 4.5005
R12560 DVSS.n20007 DVSS.n14887 4.5005
R12561 DVSS.n20007 DVSS.n14908 4.5005
R12562 DVSS.n20008 DVSS.n20007 4.5005
R12563 DVSS.n15291 DVSS.n14903 4.5005
R12564 DVSS.n18345 DVSS.n14903 4.5005
R12565 DVSS.n15318 DVSS.n14903 4.5005
R12566 DVSS.n15313 DVSS.n14903 4.5005
R12567 DVSS.n15319 DVSS.n14903 4.5005
R12568 DVSS.n15312 DVSS.n14903 4.5005
R12569 DVSS.n15320 DVSS.n14903 4.5005
R12570 DVSS.n15311 DVSS.n14903 4.5005
R12571 DVSS.n15323 DVSS.n14903 4.5005
R12572 DVSS.n15309 DVSS.n14903 4.5005
R12573 DVSS.n18343 DVSS.n14903 4.5005
R12574 DVSS.n15297 DVSS.n15291 4.5005
R12575 DVSS.n18345 DVSS.n15297 4.5005
R12576 DVSS.n15317 DVSS.n15297 4.5005
R12577 DVSS.n15314 DVSS.n15297 4.5005
R12578 DVSS.n15318 DVSS.n15297 4.5005
R12579 DVSS.n15313 DVSS.n15297 4.5005
R12580 DVSS.n15319 DVSS.n15297 4.5005
R12581 DVSS.n15312 DVSS.n15297 4.5005
R12582 DVSS.n15320 DVSS.n15297 4.5005
R12583 DVSS.n15311 DVSS.n15297 4.5005
R12584 DVSS.n15322 DVSS.n15297 4.5005
R12585 DVSS.n15310 DVSS.n15297 4.5005
R12586 DVSS.n15323 DVSS.n15297 4.5005
R12587 DVSS.n15309 DVSS.n15297 4.5005
R12588 DVSS.n18343 DVSS.n15297 4.5005
R12589 DVSS.n15300 DVSS.n15291 4.5005
R12590 DVSS.n18345 DVSS.n15300 4.5005
R12591 DVSS.n15317 DVSS.n15300 4.5005
R12592 DVSS.n15314 DVSS.n15300 4.5005
R12593 DVSS.n15318 DVSS.n15300 4.5005
R12594 DVSS.n15313 DVSS.n15300 4.5005
R12595 DVSS.n15319 DVSS.n15300 4.5005
R12596 DVSS.n15312 DVSS.n15300 4.5005
R12597 DVSS.n15320 DVSS.n15300 4.5005
R12598 DVSS.n15311 DVSS.n15300 4.5005
R12599 DVSS.n15322 DVSS.n15300 4.5005
R12600 DVSS.n15310 DVSS.n15300 4.5005
R12601 DVSS.n15323 DVSS.n15300 4.5005
R12602 DVSS.n18343 DVSS.n15300 4.5005
R12603 DVSS.n15295 DVSS.n15291 4.5005
R12604 DVSS.n18345 DVSS.n15295 4.5005
R12605 DVSS.n15317 DVSS.n15295 4.5005
R12606 DVSS.n15314 DVSS.n15295 4.5005
R12607 DVSS.n15318 DVSS.n15295 4.5005
R12608 DVSS.n15313 DVSS.n15295 4.5005
R12609 DVSS.n15319 DVSS.n15295 4.5005
R12610 DVSS.n15312 DVSS.n15295 4.5005
R12611 DVSS.n15320 DVSS.n15295 4.5005
R12612 DVSS.n15311 DVSS.n15295 4.5005
R12613 DVSS.n15322 DVSS.n15295 4.5005
R12614 DVSS.n15310 DVSS.n15295 4.5005
R12615 DVSS.n15323 DVSS.n15295 4.5005
R12616 DVSS.n18343 DVSS.n15295 4.5005
R12617 DVSS.n15302 DVSS.n15291 4.5005
R12618 DVSS.n18345 DVSS.n15302 4.5005
R12619 DVSS.n15317 DVSS.n15302 4.5005
R12620 DVSS.n15314 DVSS.n15302 4.5005
R12621 DVSS.n15318 DVSS.n15302 4.5005
R12622 DVSS.n15313 DVSS.n15302 4.5005
R12623 DVSS.n15319 DVSS.n15302 4.5005
R12624 DVSS.n15312 DVSS.n15302 4.5005
R12625 DVSS.n15320 DVSS.n15302 4.5005
R12626 DVSS.n15311 DVSS.n15302 4.5005
R12627 DVSS.n15322 DVSS.n15302 4.5005
R12628 DVSS.n15310 DVSS.n15302 4.5005
R12629 DVSS.n15323 DVSS.n15302 4.5005
R12630 DVSS.n18343 DVSS.n15302 4.5005
R12631 DVSS.n15294 DVSS.n15291 4.5005
R12632 DVSS.n18345 DVSS.n15294 4.5005
R12633 DVSS.n15317 DVSS.n15294 4.5005
R12634 DVSS.n15314 DVSS.n15294 4.5005
R12635 DVSS.n15318 DVSS.n15294 4.5005
R12636 DVSS.n15313 DVSS.n15294 4.5005
R12637 DVSS.n15319 DVSS.n15294 4.5005
R12638 DVSS.n15312 DVSS.n15294 4.5005
R12639 DVSS.n15320 DVSS.n15294 4.5005
R12640 DVSS.n15311 DVSS.n15294 4.5005
R12641 DVSS.n15322 DVSS.n15294 4.5005
R12642 DVSS.n15310 DVSS.n15294 4.5005
R12643 DVSS.n15323 DVSS.n15294 4.5005
R12644 DVSS.n18343 DVSS.n15294 4.5005
R12645 DVSS.n15304 DVSS.n15291 4.5005
R12646 DVSS.n18345 DVSS.n15304 4.5005
R12647 DVSS.n15317 DVSS.n15304 4.5005
R12648 DVSS.n15314 DVSS.n15304 4.5005
R12649 DVSS.n15318 DVSS.n15304 4.5005
R12650 DVSS.n15313 DVSS.n15304 4.5005
R12651 DVSS.n15319 DVSS.n15304 4.5005
R12652 DVSS.n15312 DVSS.n15304 4.5005
R12653 DVSS.n15320 DVSS.n15304 4.5005
R12654 DVSS.n15311 DVSS.n15304 4.5005
R12655 DVSS.n15322 DVSS.n15304 4.5005
R12656 DVSS.n15310 DVSS.n15304 4.5005
R12657 DVSS.n15323 DVSS.n15304 4.5005
R12658 DVSS.n15309 DVSS.n15304 4.5005
R12659 DVSS.n18343 DVSS.n15304 4.5005
R12660 DVSS.n15293 DVSS.n15286 4.5005
R12661 DVSS.n15293 DVSS.n15291 4.5005
R12662 DVSS.n18345 DVSS.n15293 4.5005
R12663 DVSS.n15317 DVSS.n15293 4.5005
R12664 DVSS.n15314 DVSS.n15293 4.5005
R12665 DVSS.n15318 DVSS.n15293 4.5005
R12666 DVSS.n15313 DVSS.n15293 4.5005
R12667 DVSS.n15319 DVSS.n15293 4.5005
R12668 DVSS.n15312 DVSS.n15293 4.5005
R12669 DVSS.n15320 DVSS.n15293 4.5005
R12670 DVSS.n15311 DVSS.n15293 4.5005
R12671 DVSS.n15322 DVSS.n15293 4.5005
R12672 DVSS.n15310 DVSS.n15293 4.5005
R12673 DVSS.n15323 DVSS.n15293 4.5005
R12674 DVSS.n15309 DVSS.n15293 4.5005
R12675 DVSS.n18343 DVSS.n15293 4.5005
R12676 DVSS.n17644 DVSS.n17643 4.5005
R12677 DVSS.n17643 DVSS.n16082 4.5005
R12678 DVSS.n17643 DVSS.n16080 4.5005
R12679 DVSS.n17643 DVSS.n16083 4.5005
R12680 DVSS.n17643 DVSS.n16078 4.5005
R12681 DVSS.n17643 DVSS.n16084 4.5005
R12682 DVSS.n17643 DVSS.n16077 4.5005
R12683 DVSS.n17643 DVSS.n16085 4.5005
R12684 DVSS.n17643 DVSS.n16076 4.5005
R12685 DVSS.n17643 DVSS.n16086 4.5005
R12686 DVSS.n17643 DVSS.n17642 4.5005
R12687 DVSS.n16092 DVSS.n16082 4.5005
R12688 DVSS.n16092 DVSS.n16080 4.5005
R12689 DVSS.n16103 DVSS.n16092 4.5005
R12690 DVSS.n16102 DVSS.n16092 4.5005
R12691 DVSS.n16092 DVSS.n16083 4.5005
R12692 DVSS.n16092 DVSS.n16078 4.5005
R12693 DVSS.n16092 DVSS.n16084 4.5005
R12694 DVSS.n16092 DVSS.n16077 4.5005
R12695 DVSS.n16092 DVSS.n16085 4.5005
R12696 DVSS.n16092 DVSS.n16076 4.5005
R12697 DVSS.n17640 DVSS.n16092 4.5005
R12698 DVSS.n16101 DVSS.n16092 4.5005
R12699 DVSS.n16092 DVSS.n16086 4.5005
R12700 DVSS.n17642 DVSS.n16092 4.5005
R12701 DVSS.n16094 DVSS.n16082 4.5005
R12702 DVSS.n16094 DVSS.n16080 4.5005
R12703 DVSS.n16103 DVSS.n16094 4.5005
R12704 DVSS.n16102 DVSS.n16094 4.5005
R12705 DVSS.n16094 DVSS.n16083 4.5005
R12706 DVSS.n16094 DVSS.n16078 4.5005
R12707 DVSS.n16094 DVSS.n16084 4.5005
R12708 DVSS.n16094 DVSS.n16077 4.5005
R12709 DVSS.n16094 DVSS.n16085 4.5005
R12710 DVSS.n16094 DVSS.n16076 4.5005
R12711 DVSS.n17640 DVSS.n16094 4.5005
R12712 DVSS.n16101 DVSS.n16094 4.5005
R12713 DVSS.n16094 DVSS.n16086 4.5005
R12714 DVSS.n17642 DVSS.n16094 4.5005
R12715 DVSS.n16091 DVSS.n16082 4.5005
R12716 DVSS.n16091 DVSS.n16080 4.5005
R12717 DVSS.n16103 DVSS.n16091 4.5005
R12718 DVSS.n16102 DVSS.n16091 4.5005
R12719 DVSS.n16091 DVSS.n16083 4.5005
R12720 DVSS.n16091 DVSS.n16078 4.5005
R12721 DVSS.n16091 DVSS.n16084 4.5005
R12722 DVSS.n16091 DVSS.n16077 4.5005
R12723 DVSS.n16091 DVSS.n16085 4.5005
R12724 DVSS.n16091 DVSS.n16076 4.5005
R12725 DVSS.n17640 DVSS.n16091 4.5005
R12726 DVSS.n16101 DVSS.n16091 4.5005
R12727 DVSS.n16091 DVSS.n16086 4.5005
R12728 DVSS.n17642 DVSS.n16091 4.5005
R12729 DVSS.n16095 DVSS.n16082 4.5005
R12730 DVSS.n16095 DVSS.n16080 4.5005
R12731 DVSS.n16103 DVSS.n16095 4.5005
R12732 DVSS.n16102 DVSS.n16095 4.5005
R12733 DVSS.n16095 DVSS.n16083 4.5005
R12734 DVSS.n16095 DVSS.n16078 4.5005
R12735 DVSS.n16095 DVSS.n16084 4.5005
R12736 DVSS.n16095 DVSS.n16077 4.5005
R12737 DVSS.n16095 DVSS.n16085 4.5005
R12738 DVSS.n16095 DVSS.n16076 4.5005
R12739 DVSS.n17640 DVSS.n16095 4.5005
R12740 DVSS.n16101 DVSS.n16095 4.5005
R12741 DVSS.n16095 DVSS.n16086 4.5005
R12742 DVSS.n16099 DVSS.n16095 4.5005
R12743 DVSS.n17642 DVSS.n16095 4.5005
R12744 DVSS.n16090 DVSS.n16082 4.5005
R12745 DVSS.n16090 DVSS.n16080 4.5005
R12746 DVSS.n16103 DVSS.n16090 4.5005
R12747 DVSS.n16102 DVSS.n16090 4.5005
R12748 DVSS.n16090 DVSS.n16083 4.5005
R12749 DVSS.n16090 DVSS.n16078 4.5005
R12750 DVSS.n16090 DVSS.n16084 4.5005
R12751 DVSS.n16090 DVSS.n16077 4.5005
R12752 DVSS.n16090 DVSS.n16085 4.5005
R12753 DVSS.n16090 DVSS.n16076 4.5005
R12754 DVSS.n17640 DVSS.n16090 4.5005
R12755 DVSS.n16101 DVSS.n16090 4.5005
R12756 DVSS.n16090 DVSS.n16086 4.5005
R12757 DVSS.n17642 DVSS.n16090 4.5005
R12758 DVSS.n17644 DVSS.n16070 4.5005
R12759 DVSS.n16082 DVSS.n16070 4.5005
R12760 DVSS.n16080 DVSS.n16070 4.5005
R12761 DVSS.n16103 DVSS.n16070 4.5005
R12762 DVSS.n16102 DVSS.n16070 4.5005
R12763 DVSS.n16083 DVSS.n16070 4.5005
R12764 DVSS.n16078 DVSS.n16070 4.5005
R12765 DVSS.n16084 DVSS.n16070 4.5005
R12766 DVSS.n16077 DVSS.n16070 4.5005
R12767 DVSS.n16085 DVSS.n16070 4.5005
R12768 DVSS.n16076 DVSS.n16070 4.5005
R12769 DVSS.n17640 DVSS.n16070 4.5005
R12770 DVSS.n16086 DVSS.n16070 4.5005
R12771 DVSS.n17642 DVSS.n16070 4.5005
R12772 DVSS.n16089 DVSS.n16082 4.5005
R12773 DVSS.n16089 DVSS.n16080 4.5005
R12774 DVSS.n16103 DVSS.n16089 4.5005
R12775 DVSS.n16102 DVSS.n16089 4.5005
R12776 DVSS.n16089 DVSS.n16083 4.5005
R12777 DVSS.n16089 DVSS.n16078 4.5005
R12778 DVSS.n16089 DVSS.n16084 4.5005
R12779 DVSS.n16089 DVSS.n16077 4.5005
R12780 DVSS.n16089 DVSS.n16085 4.5005
R12781 DVSS.n16089 DVSS.n16076 4.5005
R12782 DVSS.n17640 DVSS.n16089 4.5005
R12783 DVSS.n16089 DVSS.n16086 4.5005
R12784 DVSS.n16099 DVSS.n16089 4.5005
R12785 DVSS.n17642 DVSS.n16089 4.5005
R12786 DVSS.n17641 DVSS.n16082 4.5005
R12787 DVSS.n17641 DVSS.n16080 4.5005
R12788 DVSS.n17641 DVSS.n16103 4.5005
R12789 DVSS.n17641 DVSS.n16102 4.5005
R12790 DVSS.n17641 DVSS.n16083 4.5005
R12791 DVSS.n17641 DVSS.n16078 4.5005
R12792 DVSS.n17641 DVSS.n16084 4.5005
R12793 DVSS.n17641 DVSS.n16077 4.5005
R12794 DVSS.n17641 DVSS.n16085 4.5005
R12795 DVSS.n17641 DVSS.n16076 4.5005
R12796 DVSS.n17641 DVSS.n17640 4.5005
R12797 DVSS.n17641 DVSS.n16101 4.5005
R12798 DVSS.n17641 DVSS.n16086 4.5005
R12799 DVSS.n17641 DVSS.n16099 4.5005
R12800 DVSS.n17642 DVSS.n17641 4.5005
R12801 DVSS.n16266 DVSS.n16096 4.5005
R12802 DVSS.n16268 DVSS.n16096 4.5005
R12803 DVSS.n16261 DVSS.n16096 4.5005
R12804 DVSS.n16271 DVSS.n16096 4.5005
R12805 DVSS.n16259 DVSS.n16096 4.5005
R12806 DVSS.n16272 DVSS.n16096 4.5005
R12807 DVSS.n16258 DVSS.n16096 4.5005
R12808 DVSS.n16273 DVSS.n16096 4.5005
R12809 DVSS.n16257 DVSS.n16096 4.5005
R12810 DVSS.n16679 DVSS.n16096 4.5005
R12811 DVSS.n16681 DVSS.n16096 4.5005
R12812 DVSS.n16268 DVSS.n16246 4.5005
R12813 DVSS.n16261 DVSS.n16246 4.5005
R12814 DVSS.n16270 DVSS.n16246 4.5005
R12815 DVSS.n16260 DVSS.n16246 4.5005
R12816 DVSS.n16271 DVSS.n16246 4.5005
R12817 DVSS.n16259 DVSS.n16246 4.5005
R12818 DVSS.n16272 DVSS.n16246 4.5005
R12819 DVSS.n16258 DVSS.n16246 4.5005
R12820 DVSS.n16273 DVSS.n16246 4.5005
R12821 DVSS.n16257 DVSS.n16246 4.5005
R12822 DVSS.n16275 DVSS.n16246 4.5005
R12823 DVSS.n16256 DVSS.n16246 4.5005
R12824 DVSS.n16679 DVSS.n16246 4.5005
R12825 DVSS.n16681 DVSS.n16246 4.5005
R12826 DVSS.n16268 DVSS.n16247 4.5005
R12827 DVSS.n16261 DVSS.n16247 4.5005
R12828 DVSS.n16270 DVSS.n16247 4.5005
R12829 DVSS.n16260 DVSS.n16247 4.5005
R12830 DVSS.n16271 DVSS.n16247 4.5005
R12831 DVSS.n16259 DVSS.n16247 4.5005
R12832 DVSS.n16272 DVSS.n16247 4.5005
R12833 DVSS.n16258 DVSS.n16247 4.5005
R12834 DVSS.n16273 DVSS.n16247 4.5005
R12835 DVSS.n16257 DVSS.n16247 4.5005
R12836 DVSS.n16275 DVSS.n16247 4.5005
R12837 DVSS.n16256 DVSS.n16247 4.5005
R12838 DVSS.n16679 DVSS.n16247 4.5005
R12839 DVSS.n16255 DVSS.n16247 4.5005
R12840 DVSS.n16681 DVSS.n16247 4.5005
R12841 DVSS.n16268 DVSS.n16245 4.5005
R12842 DVSS.n16261 DVSS.n16245 4.5005
R12843 DVSS.n16270 DVSS.n16245 4.5005
R12844 DVSS.n16260 DVSS.n16245 4.5005
R12845 DVSS.n16271 DVSS.n16245 4.5005
R12846 DVSS.n16259 DVSS.n16245 4.5005
R12847 DVSS.n16272 DVSS.n16245 4.5005
R12848 DVSS.n16258 DVSS.n16245 4.5005
R12849 DVSS.n16273 DVSS.n16245 4.5005
R12850 DVSS.n16257 DVSS.n16245 4.5005
R12851 DVSS.n16275 DVSS.n16245 4.5005
R12852 DVSS.n16256 DVSS.n16245 4.5005
R12853 DVSS.n16679 DVSS.n16245 4.5005
R12854 DVSS.n16681 DVSS.n16245 4.5005
R12855 DVSS.n16268 DVSS.n16248 4.5005
R12856 DVSS.n16261 DVSS.n16248 4.5005
R12857 DVSS.n16270 DVSS.n16248 4.5005
R12858 DVSS.n16260 DVSS.n16248 4.5005
R12859 DVSS.n16271 DVSS.n16248 4.5005
R12860 DVSS.n16259 DVSS.n16248 4.5005
R12861 DVSS.n16272 DVSS.n16248 4.5005
R12862 DVSS.n16258 DVSS.n16248 4.5005
R12863 DVSS.n16273 DVSS.n16248 4.5005
R12864 DVSS.n16257 DVSS.n16248 4.5005
R12865 DVSS.n16275 DVSS.n16248 4.5005
R12866 DVSS.n16256 DVSS.n16248 4.5005
R12867 DVSS.n16679 DVSS.n16248 4.5005
R12868 DVSS.n16681 DVSS.n16248 4.5005
R12869 DVSS.n16268 DVSS.n16244 4.5005
R12870 DVSS.n16261 DVSS.n16244 4.5005
R12871 DVSS.n16270 DVSS.n16244 4.5005
R12872 DVSS.n16260 DVSS.n16244 4.5005
R12873 DVSS.n16271 DVSS.n16244 4.5005
R12874 DVSS.n16259 DVSS.n16244 4.5005
R12875 DVSS.n16272 DVSS.n16244 4.5005
R12876 DVSS.n16258 DVSS.n16244 4.5005
R12877 DVSS.n16273 DVSS.n16244 4.5005
R12878 DVSS.n16257 DVSS.n16244 4.5005
R12879 DVSS.n16275 DVSS.n16244 4.5005
R12880 DVSS.n16256 DVSS.n16244 4.5005
R12881 DVSS.n16679 DVSS.n16244 4.5005
R12882 DVSS.n16681 DVSS.n16244 4.5005
R12883 DVSS.n16268 DVSS.n16249 4.5005
R12884 DVSS.n16261 DVSS.n16249 4.5005
R12885 DVSS.n16270 DVSS.n16249 4.5005
R12886 DVSS.n16260 DVSS.n16249 4.5005
R12887 DVSS.n16271 DVSS.n16249 4.5005
R12888 DVSS.n16259 DVSS.n16249 4.5005
R12889 DVSS.n16272 DVSS.n16249 4.5005
R12890 DVSS.n16258 DVSS.n16249 4.5005
R12891 DVSS.n16273 DVSS.n16249 4.5005
R12892 DVSS.n16257 DVSS.n16249 4.5005
R12893 DVSS.n16275 DVSS.n16249 4.5005
R12894 DVSS.n16256 DVSS.n16249 4.5005
R12895 DVSS.n16679 DVSS.n16249 4.5005
R12896 DVSS.n16681 DVSS.n16249 4.5005
R12897 DVSS.n16268 DVSS.n16243 4.5005
R12898 DVSS.n16261 DVSS.n16243 4.5005
R12899 DVSS.n16270 DVSS.n16243 4.5005
R12900 DVSS.n16260 DVSS.n16243 4.5005
R12901 DVSS.n16271 DVSS.n16243 4.5005
R12902 DVSS.n16259 DVSS.n16243 4.5005
R12903 DVSS.n16272 DVSS.n16243 4.5005
R12904 DVSS.n16258 DVSS.n16243 4.5005
R12905 DVSS.n16273 DVSS.n16243 4.5005
R12906 DVSS.n16257 DVSS.n16243 4.5005
R12907 DVSS.n16275 DVSS.n16243 4.5005
R12908 DVSS.n16256 DVSS.n16243 4.5005
R12909 DVSS.n16679 DVSS.n16243 4.5005
R12910 DVSS.n16255 DVSS.n16243 4.5005
R12911 DVSS.n16681 DVSS.n16243 4.5005
R12912 DVSS.n15811 DVSS.n15790 4.5005
R12913 DVSS.n15813 DVSS.n15790 4.5005
R12914 DVSS.n15806 DVSS.n15790 4.5005
R12915 DVSS.n15816 DVSS.n15790 4.5005
R12916 DVSS.n15804 DVSS.n15790 4.5005
R12917 DVSS.n15817 DVSS.n15790 4.5005
R12918 DVSS.n15803 DVSS.n15790 4.5005
R12919 DVSS.n15818 DVSS.n15790 4.5005
R12920 DVSS.n15802 DVSS.n15790 4.5005
R12921 DVSS.n17906 DVSS.n15790 4.5005
R12922 DVSS.n17908 DVSS.n15790 4.5005
R12923 DVSS.n15813 DVSS.n15791 4.5005
R12924 DVSS.n15806 DVSS.n15791 4.5005
R12925 DVSS.n15815 DVSS.n15791 4.5005
R12926 DVSS.n15805 DVSS.n15791 4.5005
R12927 DVSS.n15816 DVSS.n15791 4.5005
R12928 DVSS.n15804 DVSS.n15791 4.5005
R12929 DVSS.n15817 DVSS.n15791 4.5005
R12930 DVSS.n15803 DVSS.n15791 4.5005
R12931 DVSS.n15818 DVSS.n15791 4.5005
R12932 DVSS.n15802 DVSS.n15791 4.5005
R12933 DVSS.n15820 DVSS.n15791 4.5005
R12934 DVSS.n15801 DVSS.n15791 4.5005
R12935 DVSS.n17906 DVSS.n15791 4.5005
R12936 DVSS.n17908 DVSS.n15791 4.5005
R12937 DVSS.n15813 DVSS.n15789 4.5005
R12938 DVSS.n15806 DVSS.n15789 4.5005
R12939 DVSS.n15815 DVSS.n15789 4.5005
R12940 DVSS.n15805 DVSS.n15789 4.5005
R12941 DVSS.n15816 DVSS.n15789 4.5005
R12942 DVSS.n15804 DVSS.n15789 4.5005
R12943 DVSS.n15817 DVSS.n15789 4.5005
R12944 DVSS.n15803 DVSS.n15789 4.5005
R12945 DVSS.n15818 DVSS.n15789 4.5005
R12946 DVSS.n15802 DVSS.n15789 4.5005
R12947 DVSS.n15820 DVSS.n15789 4.5005
R12948 DVSS.n15801 DVSS.n15789 4.5005
R12949 DVSS.n17906 DVSS.n15789 4.5005
R12950 DVSS.n17908 DVSS.n15789 4.5005
R12951 DVSS.n15813 DVSS.n15792 4.5005
R12952 DVSS.n15806 DVSS.n15792 4.5005
R12953 DVSS.n15815 DVSS.n15792 4.5005
R12954 DVSS.n15805 DVSS.n15792 4.5005
R12955 DVSS.n15816 DVSS.n15792 4.5005
R12956 DVSS.n15804 DVSS.n15792 4.5005
R12957 DVSS.n15817 DVSS.n15792 4.5005
R12958 DVSS.n15803 DVSS.n15792 4.5005
R12959 DVSS.n15818 DVSS.n15792 4.5005
R12960 DVSS.n15802 DVSS.n15792 4.5005
R12961 DVSS.n15820 DVSS.n15792 4.5005
R12962 DVSS.n15801 DVSS.n15792 4.5005
R12963 DVSS.n17906 DVSS.n15792 4.5005
R12964 DVSS.n17908 DVSS.n15792 4.5005
R12965 DVSS.n15813 DVSS.n15788 4.5005
R12966 DVSS.n15806 DVSS.n15788 4.5005
R12967 DVSS.n15815 DVSS.n15788 4.5005
R12968 DVSS.n15805 DVSS.n15788 4.5005
R12969 DVSS.n15816 DVSS.n15788 4.5005
R12970 DVSS.n15804 DVSS.n15788 4.5005
R12971 DVSS.n15817 DVSS.n15788 4.5005
R12972 DVSS.n15803 DVSS.n15788 4.5005
R12973 DVSS.n15818 DVSS.n15788 4.5005
R12974 DVSS.n15802 DVSS.n15788 4.5005
R12975 DVSS.n15820 DVSS.n15788 4.5005
R12976 DVSS.n15801 DVSS.n15788 4.5005
R12977 DVSS.n17906 DVSS.n15788 4.5005
R12978 DVSS.n17908 DVSS.n15788 4.5005
R12979 DVSS.n15813 DVSS.n15793 4.5005
R12980 DVSS.n15806 DVSS.n15793 4.5005
R12981 DVSS.n15815 DVSS.n15793 4.5005
R12982 DVSS.n15805 DVSS.n15793 4.5005
R12983 DVSS.n15816 DVSS.n15793 4.5005
R12984 DVSS.n15804 DVSS.n15793 4.5005
R12985 DVSS.n15817 DVSS.n15793 4.5005
R12986 DVSS.n15803 DVSS.n15793 4.5005
R12987 DVSS.n15818 DVSS.n15793 4.5005
R12988 DVSS.n15802 DVSS.n15793 4.5005
R12989 DVSS.n15820 DVSS.n15793 4.5005
R12990 DVSS.n15801 DVSS.n15793 4.5005
R12991 DVSS.n17906 DVSS.n15793 4.5005
R12992 DVSS.n17908 DVSS.n15793 4.5005
R12993 DVSS.n15813 DVSS.n15787 4.5005
R12994 DVSS.n15806 DVSS.n15787 4.5005
R12995 DVSS.n15815 DVSS.n15787 4.5005
R12996 DVSS.n15805 DVSS.n15787 4.5005
R12997 DVSS.n15816 DVSS.n15787 4.5005
R12998 DVSS.n15804 DVSS.n15787 4.5005
R12999 DVSS.n15817 DVSS.n15787 4.5005
R13000 DVSS.n15803 DVSS.n15787 4.5005
R13001 DVSS.n15818 DVSS.n15787 4.5005
R13002 DVSS.n15802 DVSS.n15787 4.5005
R13003 DVSS.n15820 DVSS.n15787 4.5005
R13004 DVSS.n15801 DVSS.n15787 4.5005
R13005 DVSS.n17906 DVSS.n15787 4.5005
R13006 DVSS.n17908 DVSS.n15787 4.5005
R13007 DVSS.n15813 DVSS.n15794 4.5005
R13008 DVSS.n15806 DVSS.n15794 4.5005
R13009 DVSS.n15815 DVSS.n15794 4.5005
R13010 DVSS.n15805 DVSS.n15794 4.5005
R13011 DVSS.n15816 DVSS.n15794 4.5005
R13012 DVSS.n15804 DVSS.n15794 4.5005
R13013 DVSS.n15817 DVSS.n15794 4.5005
R13014 DVSS.n15803 DVSS.n15794 4.5005
R13015 DVSS.n15818 DVSS.n15794 4.5005
R13016 DVSS.n15802 DVSS.n15794 4.5005
R13017 DVSS.n15820 DVSS.n15794 4.5005
R13018 DVSS.n15801 DVSS.n15794 4.5005
R13019 DVSS.n17906 DVSS.n15794 4.5005
R13020 DVSS.n17908 DVSS.n15794 4.5005
R13021 DVSS.n15813 DVSS.n15786 4.5005
R13022 DVSS.n15806 DVSS.n15786 4.5005
R13023 DVSS.n15815 DVSS.n15786 4.5005
R13024 DVSS.n15805 DVSS.n15786 4.5005
R13025 DVSS.n15816 DVSS.n15786 4.5005
R13026 DVSS.n15804 DVSS.n15786 4.5005
R13027 DVSS.n15817 DVSS.n15786 4.5005
R13028 DVSS.n15803 DVSS.n15786 4.5005
R13029 DVSS.n15818 DVSS.n15786 4.5005
R13030 DVSS.n15802 DVSS.n15786 4.5005
R13031 DVSS.n15820 DVSS.n15786 4.5005
R13032 DVSS.n15801 DVSS.n15786 4.5005
R13033 DVSS.n17906 DVSS.n15786 4.5005
R13034 DVSS.n15800 DVSS.n15786 4.5005
R13035 DVSS.n17908 DVSS.n15786 4.5005
R13036 DVSS.n17907 DVSS.n15811 4.5005
R13037 DVSS.n17907 DVSS.n15813 4.5005
R13038 DVSS.n17907 DVSS.n15806 4.5005
R13039 DVSS.n17907 DVSS.n15815 4.5005
R13040 DVSS.n17907 DVSS.n15805 4.5005
R13041 DVSS.n17907 DVSS.n15816 4.5005
R13042 DVSS.n17907 DVSS.n15804 4.5005
R13043 DVSS.n17907 DVSS.n15817 4.5005
R13044 DVSS.n17907 DVSS.n15803 4.5005
R13045 DVSS.n17907 DVSS.n15818 4.5005
R13046 DVSS.n17907 DVSS.n15802 4.5005
R13047 DVSS.n17907 DVSS.n15820 4.5005
R13048 DVSS.n17907 DVSS.n15801 4.5005
R13049 DVSS.n17907 DVSS.n17906 4.5005
R13050 DVSS.n17907 DVSS.n15800 4.5005
R13051 DVSS.n17908 DVSS.n17907 4.5005
R13052 DVSS.n16268 DVSS.n16250 4.5005
R13053 DVSS.n16261 DVSS.n16250 4.5005
R13054 DVSS.n16270 DVSS.n16250 4.5005
R13055 DVSS.n16260 DVSS.n16250 4.5005
R13056 DVSS.n16271 DVSS.n16250 4.5005
R13057 DVSS.n16259 DVSS.n16250 4.5005
R13058 DVSS.n16272 DVSS.n16250 4.5005
R13059 DVSS.n16258 DVSS.n16250 4.5005
R13060 DVSS.n16273 DVSS.n16250 4.5005
R13061 DVSS.n16257 DVSS.n16250 4.5005
R13062 DVSS.n16275 DVSS.n16250 4.5005
R13063 DVSS.n16256 DVSS.n16250 4.5005
R13064 DVSS.n16679 DVSS.n16250 4.5005
R13065 DVSS.n16255 DVSS.n16250 4.5005
R13066 DVSS.n16681 DVSS.n16250 4.5005
R13067 DVSS.n16266 DVSS.n16242 4.5005
R13068 DVSS.n16268 DVSS.n16242 4.5005
R13069 DVSS.n16261 DVSS.n16242 4.5005
R13070 DVSS.n16270 DVSS.n16242 4.5005
R13071 DVSS.n16260 DVSS.n16242 4.5005
R13072 DVSS.n16271 DVSS.n16242 4.5005
R13073 DVSS.n16259 DVSS.n16242 4.5005
R13074 DVSS.n16272 DVSS.n16242 4.5005
R13075 DVSS.n16258 DVSS.n16242 4.5005
R13076 DVSS.n16273 DVSS.n16242 4.5005
R13077 DVSS.n16257 DVSS.n16242 4.5005
R13078 DVSS.n16275 DVSS.n16242 4.5005
R13079 DVSS.n16256 DVSS.n16242 4.5005
R13080 DVSS.n16679 DVSS.n16242 4.5005
R13081 DVSS.n16255 DVSS.n16242 4.5005
R13082 DVSS.n16681 DVSS.n16242 4.5005
R13083 DVSS.n16680 DVSS.n16266 4.5005
R13084 DVSS.n16680 DVSS.n16268 4.5005
R13085 DVSS.n16680 DVSS.n16261 4.5005
R13086 DVSS.n16680 DVSS.n16270 4.5005
R13087 DVSS.n16680 DVSS.n16260 4.5005
R13088 DVSS.n16680 DVSS.n16271 4.5005
R13089 DVSS.n16680 DVSS.n16259 4.5005
R13090 DVSS.n16680 DVSS.n16272 4.5005
R13091 DVSS.n16680 DVSS.n16258 4.5005
R13092 DVSS.n16680 DVSS.n16273 4.5005
R13093 DVSS.n16680 DVSS.n16257 4.5005
R13094 DVSS.n16680 DVSS.n16275 4.5005
R13095 DVSS.n16680 DVSS.n16256 4.5005
R13096 DVSS.n16680 DVSS.n16679 4.5005
R13097 DVSS.n16680 DVSS.n16255 4.5005
R13098 DVSS.n16681 DVSS.n16680 4.5005
R13099 DVSS.n16088 DVSS.n16082 4.5005
R13100 DVSS.n16088 DVSS.n16080 4.5005
R13101 DVSS.n16103 DVSS.n16088 4.5005
R13102 DVSS.n16102 DVSS.n16088 4.5005
R13103 DVSS.n16088 DVSS.n16083 4.5005
R13104 DVSS.n16088 DVSS.n16078 4.5005
R13105 DVSS.n16088 DVSS.n16084 4.5005
R13106 DVSS.n16088 DVSS.n16077 4.5005
R13107 DVSS.n16088 DVSS.n16085 4.5005
R13108 DVSS.n16088 DVSS.n16076 4.5005
R13109 DVSS.n17640 DVSS.n16088 4.5005
R13110 DVSS.n16101 DVSS.n16088 4.5005
R13111 DVSS.n16088 DVSS.n16086 4.5005
R13112 DVSS.n16099 DVSS.n16088 4.5005
R13113 DVSS.n17642 DVSS.n16088 4.5005
R13114 DVSS.n17644 DVSS.n16067 4.5005
R13115 DVSS.n16082 DVSS.n16067 4.5005
R13116 DVSS.n16080 DVSS.n16067 4.5005
R13117 DVSS.n16103 DVSS.n16067 4.5005
R13118 DVSS.n16102 DVSS.n16067 4.5005
R13119 DVSS.n16083 DVSS.n16067 4.5005
R13120 DVSS.n16078 DVSS.n16067 4.5005
R13121 DVSS.n16084 DVSS.n16067 4.5005
R13122 DVSS.n16077 DVSS.n16067 4.5005
R13123 DVSS.n16085 DVSS.n16067 4.5005
R13124 DVSS.n16076 DVSS.n16067 4.5005
R13125 DVSS.n17640 DVSS.n16067 4.5005
R13126 DVSS.n16101 DVSS.n16067 4.5005
R13127 DVSS.n16086 DVSS.n16067 4.5005
R13128 DVSS.n16099 DVSS.n16067 4.5005
R13129 DVSS.n17642 DVSS.n16067 4.5005
R13130 DVSS.n15305 DVSS.n15286 4.5005
R13131 DVSS.n15305 DVSS.n15291 4.5005
R13132 DVSS.n18345 DVSS.n15305 4.5005
R13133 DVSS.n15317 DVSS.n15305 4.5005
R13134 DVSS.n15314 DVSS.n15305 4.5005
R13135 DVSS.n15318 DVSS.n15305 4.5005
R13136 DVSS.n15313 DVSS.n15305 4.5005
R13137 DVSS.n15319 DVSS.n15305 4.5005
R13138 DVSS.n15312 DVSS.n15305 4.5005
R13139 DVSS.n15320 DVSS.n15305 4.5005
R13140 DVSS.n15311 DVSS.n15305 4.5005
R13141 DVSS.n15322 DVSS.n15305 4.5005
R13142 DVSS.n15310 DVSS.n15305 4.5005
R13143 DVSS.n15323 DVSS.n15305 4.5005
R13144 DVSS.n15309 DVSS.n15305 4.5005
R13145 DVSS.n18343 DVSS.n15305 4.5005
R13146 DVSS.n15292 DVSS.n15291 4.5005
R13147 DVSS.n18345 DVSS.n15292 4.5005
R13148 DVSS.n15317 DVSS.n15292 4.5005
R13149 DVSS.n15314 DVSS.n15292 4.5005
R13150 DVSS.n15318 DVSS.n15292 4.5005
R13151 DVSS.n15313 DVSS.n15292 4.5005
R13152 DVSS.n15319 DVSS.n15292 4.5005
R13153 DVSS.n15312 DVSS.n15292 4.5005
R13154 DVSS.n15320 DVSS.n15292 4.5005
R13155 DVSS.n15311 DVSS.n15292 4.5005
R13156 DVSS.n15322 DVSS.n15292 4.5005
R13157 DVSS.n15310 DVSS.n15292 4.5005
R13158 DVSS.n15323 DVSS.n15292 4.5005
R13159 DVSS.n15309 DVSS.n15292 4.5005
R13160 DVSS.n18343 DVSS.n15292 4.5005
R13161 DVSS.n18344 DVSS.n15286 4.5005
R13162 DVSS.n18344 DVSS.n15291 4.5005
R13163 DVSS.n18345 DVSS.n18344 4.5005
R13164 DVSS.n18344 DVSS.n15317 4.5005
R13165 DVSS.n18344 DVSS.n15314 4.5005
R13166 DVSS.n18344 DVSS.n15318 4.5005
R13167 DVSS.n18344 DVSS.n15313 4.5005
R13168 DVSS.n18344 DVSS.n15319 4.5005
R13169 DVSS.n18344 DVSS.n15312 4.5005
R13170 DVSS.n18344 DVSS.n15320 4.5005
R13171 DVSS.n18344 DVSS.n15311 4.5005
R13172 DVSS.n18344 DVSS.n15322 4.5005
R13173 DVSS.n18344 DVSS.n15310 4.5005
R13174 DVSS.n18344 DVSS.n15323 4.5005
R13175 DVSS.n18344 DVSS.n15309 4.5005
R13176 DVSS.n18344 DVSS.n18343 4.5005
R13177 DVSS.n1197 DVSS.n1196 4.5005
R13178 DVSS.n22338 DVSS.n1197 4.5005
R13179 DVSS.n1292 DVSS.n573 4.5005
R13180 DVSS.n1311 DVSS.n562 4.5005
R13181 DVSS.n22340 DVSS.n22339 4.5005
R13182 DVSS.n22339 DVSS.n22338 4.5005
R13183 DVSS.n14631 DVSS.n14630 4.5005
R13184 DVSS.n20648 DVSS.n14631 4.5005
R13185 DVSS.n14641 DVSS.n14631 4.5005
R13186 DVSS.n14640 DVSS.n14631 4.5005
R13187 DVSS.n14642 DVSS.n14631 4.5005
R13188 DVSS.n14639 DVSS.n14631 4.5005
R13189 DVSS.n14643 DVSS.n14631 4.5005
R13190 DVSS.n14638 DVSS.n14631 4.5005
R13191 DVSS.n14644 DVSS.n14631 4.5005
R13192 DVSS.n14637 DVSS.n14631 4.5005
R13193 DVSS.n14645 DVSS.n14631 4.5005
R13194 DVSS.n14636 DVSS.n14631 4.5005
R13195 DVSS.n14646 DVSS.n14631 4.5005
R13196 DVSS.n14635 DVSS.n14631 4.5005
R13197 DVSS.n14647 DVSS.n14631 4.5005
R13198 DVSS.n20646 DVSS.n14631 4.5005
R13199 DVSS.n14625 DVSS.n14074 4.5005
R13200 DVSS.n20221 DVSS.n14074 4.5005
R13201 DVSS.n20219 DVSS.n14074 4.5005
R13202 DVSS.n20222 DVSS.n14074 4.5005
R13203 DVSS.n20218 DVSS.n14074 4.5005
R13204 DVSS.n20223 DVSS.n14074 4.5005
R13205 DVSS.n20217 DVSS.n14074 4.5005
R13206 DVSS.n20224 DVSS.n14074 4.5005
R13207 DVSS.n20216 DVSS.n14074 4.5005
R13208 DVSS.n20298 DVSS.n14074 4.5005
R13209 DVSS.n20215 DVSS.n14074 4.5005
R13210 DVSS.n20208 DVSS.n14074 4.5005
R13211 DVSS.n20305 DVSS.n14074 4.5005
R13212 DVSS.n20302 DVSS.n14074 4.5005
R13213 DVSS.n20300 DVSS.n14074 4.5005
R13214 DVSS.n14660 DVSS.n14074 4.5005
R13215 DVSS.n20211 DVSS.n14625 4.5005
R13216 DVSS.n20221 DVSS.n20211 4.5005
R13217 DVSS.n20219 DVSS.n20211 4.5005
R13218 DVSS.n20222 DVSS.n20211 4.5005
R13219 DVSS.n20218 DVSS.n20211 4.5005
R13220 DVSS.n20223 DVSS.n20211 4.5005
R13221 DVSS.n20217 DVSS.n20211 4.5005
R13222 DVSS.n20224 DVSS.n20211 4.5005
R13223 DVSS.n20216 DVSS.n20211 4.5005
R13224 DVSS.n20298 DVSS.n20211 4.5005
R13225 DVSS.n20215 DVSS.n20211 4.5005
R13226 DVSS.n20211 DVSS.n20208 4.5005
R13227 DVSS.n20305 DVSS.n20211 4.5005
R13228 DVSS.n20302 DVSS.n20211 4.5005
R13229 DVSS.n20300 DVSS.n20211 4.5005
R13230 DVSS.n20211 DVSS.n14660 4.5005
R13231 DVSS.n20209 DVSS.n14625 4.5005
R13232 DVSS.n20221 DVSS.n20209 4.5005
R13233 DVSS.n20219 DVSS.n20209 4.5005
R13234 DVSS.n20222 DVSS.n20209 4.5005
R13235 DVSS.n20218 DVSS.n20209 4.5005
R13236 DVSS.n20223 DVSS.n20209 4.5005
R13237 DVSS.n20217 DVSS.n20209 4.5005
R13238 DVSS.n20224 DVSS.n20209 4.5005
R13239 DVSS.n20216 DVSS.n20209 4.5005
R13240 DVSS.n20298 DVSS.n20209 4.5005
R13241 DVSS.n20215 DVSS.n20209 4.5005
R13242 DVSS.n20209 DVSS.n20208 4.5005
R13243 DVSS.n20305 DVSS.n20209 4.5005
R13244 DVSS.n20302 DVSS.n20209 4.5005
R13245 DVSS.n20300 DVSS.n20209 4.5005
R13246 DVSS.n20209 DVSS.n14660 4.5005
R13247 DVSS.n20185 DVSS.n14425 4.5005
R13248 DVSS.n14873 DVSS.n14425 4.5005
R13249 DVSS.n20186 DVSS.n14425 4.5005
R13250 DVSS.n14872 DVSS.n14425 4.5005
R13251 DVSS.n20187 DVSS.n14425 4.5005
R13252 DVSS.n14871 DVSS.n14425 4.5005
R13253 DVSS.n20188 DVSS.n14425 4.5005
R13254 DVSS.n14870 DVSS.n14425 4.5005
R13255 DVSS.n20189 DVSS.n14425 4.5005
R13256 DVSS.n14869 DVSS.n14425 4.5005
R13257 DVSS.n20190 DVSS.n14425 4.5005
R13258 DVSS.n14868 DVSS.n14425 4.5005
R13259 DVSS.n20191 DVSS.n14425 4.5005
R13260 DVSS.n14867 DVSS.n14425 4.5005
R13261 DVSS.n20192 DVSS.n14425 4.5005
R13262 DVSS.n20317 DVSS.n14425 4.5005
R13263 DVSS.n20316 DVSS.n20185 4.5005
R13264 DVSS.n20316 DVSS.n14873 4.5005
R13265 DVSS.n20316 DVSS.n20186 4.5005
R13266 DVSS.n20316 DVSS.n14872 4.5005
R13267 DVSS.n20316 DVSS.n20187 4.5005
R13268 DVSS.n20316 DVSS.n14871 4.5005
R13269 DVSS.n20316 DVSS.n20188 4.5005
R13270 DVSS.n20316 DVSS.n14870 4.5005
R13271 DVSS.n20316 DVSS.n20189 4.5005
R13272 DVSS.n20316 DVSS.n14869 4.5005
R13273 DVSS.n20316 DVSS.n20190 4.5005
R13274 DVSS.n20316 DVSS.n14868 4.5005
R13275 DVSS.n20316 DVSS.n20191 4.5005
R13276 DVSS.n20316 DVSS.n14867 4.5005
R13277 DVSS.n20316 DVSS.n20192 4.5005
R13278 DVSS.n20316 DVSS.n14866 4.5005
R13279 DVSS.n20316 DVSS.n20315 4.5005
R13280 DVSS.n20317 DVSS.n20316 4.5005
R13281 DVSS.n20212 DVSS.n14625 4.5005
R13282 DVSS.n20221 DVSS.n20212 4.5005
R13283 DVSS.n20219 DVSS.n20212 4.5005
R13284 DVSS.n20222 DVSS.n20212 4.5005
R13285 DVSS.n20218 DVSS.n20212 4.5005
R13286 DVSS.n20223 DVSS.n20212 4.5005
R13287 DVSS.n20217 DVSS.n20212 4.5005
R13288 DVSS.n20224 DVSS.n20212 4.5005
R13289 DVSS.n20216 DVSS.n20212 4.5005
R13290 DVSS.n20298 DVSS.n20212 4.5005
R13291 DVSS.n20215 DVSS.n20212 4.5005
R13292 DVSS.n20212 DVSS.n20208 4.5005
R13293 DVSS.n20305 DVSS.n20212 4.5005
R13294 DVSS.n20302 DVSS.n20212 4.5005
R13295 DVSS.n20212 DVSS.n14660 4.5005
R13296 DVSS.n20303 DVSS.n14625 4.5005
R13297 DVSS.n20303 DVSS.n20221 4.5005
R13298 DVSS.n20303 DVSS.n20219 4.5005
R13299 DVSS.n20303 DVSS.n20222 4.5005
R13300 DVSS.n20303 DVSS.n20218 4.5005
R13301 DVSS.n20303 DVSS.n20223 4.5005
R13302 DVSS.n20303 DVSS.n20217 4.5005
R13303 DVSS.n20303 DVSS.n20224 4.5005
R13304 DVSS.n20303 DVSS.n20216 4.5005
R13305 DVSS.n20303 DVSS.n20298 4.5005
R13306 DVSS.n20303 DVSS.n20215 4.5005
R13307 DVSS.n20303 DVSS.n20208 4.5005
R13308 DVSS.n20303 DVSS.n20302 4.5005
R13309 DVSS.n20303 DVSS.n14660 4.5005
R13310 DVSS.n14625 DVSS.n14044 4.5005
R13311 DVSS.n20221 DVSS.n14044 4.5005
R13312 DVSS.n20219 DVSS.n14044 4.5005
R13313 DVSS.n20222 DVSS.n14044 4.5005
R13314 DVSS.n20218 DVSS.n14044 4.5005
R13315 DVSS.n20223 DVSS.n14044 4.5005
R13316 DVSS.n20217 DVSS.n14044 4.5005
R13317 DVSS.n20224 DVSS.n14044 4.5005
R13318 DVSS.n20216 DVSS.n14044 4.5005
R13319 DVSS.n20298 DVSS.n14044 4.5005
R13320 DVSS.n20215 DVSS.n14044 4.5005
R13321 DVSS.n20208 DVSS.n14044 4.5005
R13322 DVSS.n20302 DVSS.n14044 4.5005
R13323 DVSS.n20300 DVSS.n14044 4.5005
R13324 DVSS.n14660 DVSS.n14044 4.5005
R13325 DVSS.n20647 DVSS.n14630 4.5005
R13326 DVSS.n20648 DVSS.n20647 4.5005
R13327 DVSS.n20647 DVSS.n14641 4.5005
R13328 DVSS.n20647 DVSS.n14640 4.5005
R13329 DVSS.n20647 DVSS.n14642 4.5005
R13330 DVSS.n20647 DVSS.n14639 4.5005
R13331 DVSS.n20647 DVSS.n14643 4.5005
R13332 DVSS.n20647 DVSS.n14638 4.5005
R13333 DVSS.n20647 DVSS.n14644 4.5005
R13334 DVSS.n20647 DVSS.n14637 4.5005
R13335 DVSS.n20647 DVSS.n14645 4.5005
R13336 DVSS.n20647 DVSS.n14636 4.5005
R13337 DVSS.n20647 DVSS.n14646 4.5005
R13338 DVSS.n20647 DVSS.n14635 4.5005
R13339 DVSS.n20647 DVSS.n14647 4.5005
R13340 DVSS.n20647 DVSS.n14634 4.5005
R13341 DVSS.n20647 DVSS.n14649 4.5005
R13342 DVSS.n20647 DVSS.n20646 4.5005
R13343 DVSS.n17077 DVSS.n16827 4.5005
R13344 DVSS.n17014 DVSS.n15387 4.5005
R13345 DVSS.n17492 DVSS.n17491 4.5005
R13346 DVSS.n17493 DVSS.n17492 4.5005
R13347 DVSS.n17489 DVSS.n16940 4.5005
R13348 DVSS.n17493 DVSS.n16940 4.5005
R13349 DVSS.n17416 DVSS.n17234 4.5005
R13350 DVSS.n17416 DVSS.n17415 4.5005
R13351 DVSS.n17417 DVSS.n17416 4.5005
R13352 DVSS.n17413 DVSS.n17224 4.5005
R13353 DVSS.n17244 DVSS.n17224 4.5005
R13354 DVSS.n17415 DVSS.n17224 4.5005
R13355 DVSS.n17417 DVSS.n17224 4.5005
R13356 DVSS.n17468 DVSS.n17467 4.5005
R13357 DVSS.n17468 DVSS.n17196 4.5005
R13358 DVSS.n17469 DVSS.n17468 4.5005
R13359 DVSS.n17196 DVSS.n17173 4.5005
R13360 DVSS.n17471 DVSS.n17173 4.5005
R13361 DVSS.n17415 DVSS.n17414 4.5005
R13362 DVSS.n17414 DVSS.n17247 4.5005
R13363 DVSS.n17414 DVSS.n17243 4.5005
R13364 DVSS.n17414 DVSS.n17249 4.5005
R13365 DVSS.n17414 DVSS.n17242 4.5005
R13366 DVSS.n17414 DVSS.n17251 4.5005
R13367 DVSS.n17414 DVSS.n17241 4.5005
R13368 DVSS.n17414 DVSS.n17253 4.5005
R13369 DVSS.n17414 DVSS.n17240 4.5005
R13370 DVSS.n17414 DVSS.n17255 4.5005
R13371 DVSS.n17414 DVSS.n17239 4.5005
R13372 DVSS.n17414 DVSS.n17257 4.5005
R13373 DVSS.n17414 DVSS.n17238 4.5005
R13374 DVSS.n17414 DVSS.n17413 4.5005
R13375 DVSS.n17491 DVSS.n17490 4.5005
R13376 DVSS.n17490 DVSS.n16959 4.5005
R13377 DVSS.n17490 DVSS.n16961 4.5005
R13378 DVSS.n17490 DVSS.n16958 4.5005
R13379 DVSS.n17490 DVSS.n16963 4.5005
R13380 DVSS.n17490 DVSS.n16957 4.5005
R13381 DVSS.n17490 DVSS.n16965 4.5005
R13382 DVSS.n17490 DVSS.n16956 4.5005
R13383 DVSS.n17490 DVSS.n16967 4.5005
R13384 DVSS.n17490 DVSS.n16955 4.5005
R13385 DVSS.n17490 DVSS.n16969 4.5005
R13386 DVSS.n17490 DVSS.n16954 4.5005
R13387 DVSS.n17490 DVSS.n16971 4.5005
R13388 DVSS.n17490 DVSS.n16953 4.5005
R13389 DVSS.n17490 DVSS.n16973 4.5005
R13390 DVSS.n17490 DVSS.n16952 4.5005
R13391 DVSS.n17490 DVSS.n17489 4.5005
R13392 DVSS.n17096 DVSS.n16843 4.5005
R13393 DVSS.n16995 DVSS.n15373 4.5005
R13394 DVSS.n17471 DVSS.n17470 4.5005
R13395 DVSS.n17470 DVSS.n17182 4.5005
R13396 DVSS.n17470 DVSS.n17184 4.5005
R13397 DVSS.n17470 DVSS.n17181 4.5005
R13398 DVSS.n17470 DVSS.n17186 4.5005
R13399 DVSS.n17470 DVSS.n17180 4.5005
R13400 DVSS.n17470 DVSS.n17188 4.5005
R13401 DVSS.n17470 DVSS.n17179 4.5005
R13402 DVSS.n17470 DVSS.n17190 4.5005
R13403 DVSS.n17470 DVSS.n17178 4.5005
R13404 DVSS.n17470 DVSS.n17192 4.5005
R13405 DVSS.n17470 DVSS.n17177 4.5005
R13406 DVSS.n17470 DVSS.n17194 4.5005
R13407 DVSS.n17470 DVSS.n17176 4.5005
R13408 DVSS.n17470 DVSS.n17196 4.5005
R13409 DVSS.n17470 DVSS.n17469 4.5005
R13410 DVSS.n16200 DVSS.n16176 4.5005
R13411 DVSS.n16192 DVSS.n16176 4.5005
R13412 DVSS.n16195 DVSS.n16176 4.5005
R13413 DVSS.n16222 DVSS.n16220 4.5005
R13414 DVSS.n16223 DVSS.n16195 4.5005
R13415 DVSS.n16223 DVSS.n16194 4.5005
R13416 DVSS.n16223 DVSS.n16197 4.5005
R13417 DVSS.n16223 DVSS.n16193 4.5005
R13418 DVSS.n16223 DVSS.n16199 4.5005
R13419 DVSS.n16223 DVSS.n16192 4.5005
R13420 DVSS.n16223 DVSS.n16200 4.5005
R13421 DVSS.n16223 DVSS.n16191 4.5005
R13422 DVSS.n16223 DVSS.n16202 4.5005
R13423 DVSS.n16223 DVSS.n16190 4.5005
R13424 DVSS.n16223 DVSS.n16204 4.5005
R13425 DVSS.n16223 DVSS.n16189 4.5005
R13426 DVSS.n16223 DVSS.n16206 4.5005
R13427 DVSS.n16223 DVSS.n16188 4.5005
R13428 DVSS.n16223 DVSS.n16208 4.5005
R13429 DVSS.n16223 DVSS.n16187 4.5005
R13430 DVSS.n16223 DVSS.n16210 4.5005
R13431 DVSS.n16223 DVSS.n16186 4.5005
R13432 DVSS.n16223 DVSS.n16222 4.5005
R13433 DVSS.n13488 DVSS.n13472 4.5005
R13434 DVSS.n13489 DVSS.n13472 4.5005
R13435 DVSS.n13487 DVSS.n13472 4.5005
R13436 DVSS.n13492 DVSS.n13472 4.5005
R13437 DVSS.n13485 DVSS.n13472 4.5005
R13438 DVSS.n13493 DVSS.n13472 4.5005
R13439 DVSS.n13484 DVSS.n13472 4.5005
R13440 DVSS.n13494 DVSS.n13472 4.5005
R13441 DVSS.n13483 DVSS.n13472 4.5005
R13442 DVSS.n21338 DVSS.n13472 4.5005
R13443 DVSS.n21340 DVSS.n13472 4.5005
R13444 DVSS.n13488 DVSS.n13470 4.5005
R13445 DVSS.n13489 DVSS.n13470 4.5005
R13446 DVSS.n13487 DVSS.n13470 4.5005
R13447 DVSS.n13491 DVSS.n13470 4.5005
R13448 DVSS.n13486 DVSS.n13470 4.5005
R13449 DVSS.n13492 DVSS.n13470 4.5005
R13450 DVSS.n13485 DVSS.n13470 4.5005
R13451 DVSS.n13493 DVSS.n13470 4.5005
R13452 DVSS.n13484 DVSS.n13470 4.5005
R13453 DVSS.n13494 DVSS.n13470 4.5005
R13454 DVSS.n13483 DVSS.n13470 4.5005
R13455 DVSS.n13495 DVSS.n13470 4.5005
R13456 DVSS.n21338 DVSS.n13470 4.5005
R13457 DVSS.n21340 DVSS.n13470 4.5005
R13458 DVSS.n13488 DVSS.n13474 4.5005
R13459 DVSS.n13489 DVSS.n13474 4.5005
R13460 DVSS.n13487 DVSS.n13474 4.5005
R13461 DVSS.n13491 DVSS.n13474 4.5005
R13462 DVSS.n13486 DVSS.n13474 4.5005
R13463 DVSS.n13492 DVSS.n13474 4.5005
R13464 DVSS.n13485 DVSS.n13474 4.5005
R13465 DVSS.n13493 DVSS.n13474 4.5005
R13466 DVSS.n13484 DVSS.n13474 4.5005
R13467 DVSS.n13494 DVSS.n13474 4.5005
R13468 DVSS.n13483 DVSS.n13474 4.5005
R13469 DVSS.n13495 DVSS.n13474 4.5005
R13470 DVSS.n21338 DVSS.n13474 4.5005
R13471 DVSS.n21340 DVSS.n13474 4.5005
R13472 DVSS.n13488 DVSS.n13469 4.5005
R13473 DVSS.n13489 DVSS.n13469 4.5005
R13474 DVSS.n13487 DVSS.n13469 4.5005
R13475 DVSS.n13491 DVSS.n13469 4.5005
R13476 DVSS.n13486 DVSS.n13469 4.5005
R13477 DVSS.n13492 DVSS.n13469 4.5005
R13478 DVSS.n13485 DVSS.n13469 4.5005
R13479 DVSS.n13493 DVSS.n13469 4.5005
R13480 DVSS.n13484 DVSS.n13469 4.5005
R13481 DVSS.n13494 DVSS.n13469 4.5005
R13482 DVSS.n13483 DVSS.n13469 4.5005
R13483 DVSS.n13495 DVSS.n13469 4.5005
R13484 DVSS.n21338 DVSS.n13469 4.5005
R13485 DVSS.n21340 DVSS.n13469 4.5005
R13486 DVSS.n13488 DVSS.n13476 4.5005
R13487 DVSS.n13489 DVSS.n13476 4.5005
R13488 DVSS.n13487 DVSS.n13476 4.5005
R13489 DVSS.n13491 DVSS.n13476 4.5005
R13490 DVSS.n13486 DVSS.n13476 4.5005
R13491 DVSS.n13492 DVSS.n13476 4.5005
R13492 DVSS.n13485 DVSS.n13476 4.5005
R13493 DVSS.n13493 DVSS.n13476 4.5005
R13494 DVSS.n13484 DVSS.n13476 4.5005
R13495 DVSS.n13494 DVSS.n13476 4.5005
R13496 DVSS.n13483 DVSS.n13476 4.5005
R13497 DVSS.n13495 DVSS.n13476 4.5005
R13498 DVSS.n21338 DVSS.n13476 4.5005
R13499 DVSS.n21340 DVSS.n13476 4.5005
R13500 DVSS.n13488 DVSS.n13468 4.5005
R13501 DVSS.n13489 DVSS.n13468 4.5005
R13502 DVSS.n13487 DVSS.n13468 4.5005
R13503 DVSS.n13491 DVSS.n13468 4.5005
R13504 DVSS.n13486 DVSS.n13468 4.5005
R13505 DVSS.n13492 DVSS.n13468 4.5005
R13506 DVSS.n13485 DVSS.n13468 4.5005
R13507 DVSS.n13493 DVSS.n13468 4.5005
R13508 DVSS.n13484 DVSS.n13468 4.5005
R13509 DVSS.n13494 DVSS.n13468 4.5005
R13510 DVSS.n13483 DVSS.n13468 4.5005
R13511 DVSS.n13495 DVSS.n13468 4.5005
R13512 DVSS.n21338 DVSS.n13468 4.5005
R13513 DVSS.n21340 DVSS.n13468 4.5005
R13514 DVSS.n13488 DVSS.n13478 4.5005
R13515 DVSS.n13489 DVSS.n13478 4.5005
R13516 DVSS.n13487 DVSS.n13478 4.5005
R13517 DVSS.n13491 DVSS.n13478 4.5005
R13518 DVSS.n13486 DVSS.n13478 4.5005
R13519 DVSS.n13492 DVSS.n13478 4.5005
R13520 DVSS.n13485 DVSS.n13478 4.5005
R13521 DVSS.n13493 DVSS.n13478 4.5005
R13522 DVSS.n13484 DVSS.n13478 4.5005
R13523 DVSS.n13494 DVSS.n13478 4.5005
R13524 DVSS.n13483 DVSS.n13478 4.5005
R13525 DVSS.n13495 DVSS.n13478 4.5005
R13526 DVSS.n21338 DVSS.n13478 4.5005
R13527 DVSS.n21340 DVSS.n13478 4.5005
R13528 DVSS.n13488 DVSS.n13467 4.5005
R13529 DVSS.n13489 DVSS.n13467 4.5005
R13530 DVSS.n13487 DVSS.n13467 4.5005
R13531 DVSS.n13491 DVSS.n13467 4.5005
R13532 DVSS.n13486 DVSS.n13467 4.5005
R13533 DVSS.n13492 DVSS.n13467 4.5005
R13534 DVSS.n13485 DVSS.n13467 4.5005
R13535 DVSS.n13493 DVSS.n13467 4.5005
R13536 DVSS.n13484 DVSS.n13467 4.5005
R13537 DVSS.n13494 DVSS.n13467 4.5005
R13538 DVSS.n13483 DVSS.n13467 4.5005
R13539 DVSS.n13495 DVSS.n13467 4.5005
R13540 DVSS.n21338 DVSS.n13467 4.5005
R13541 DVSS.n21340 DVSS.n13467 4.5005
R13542 DVSS.n13488 DVSS.n13480 4.5005
R13543 DVSS.n13489 DVSS.n13480 4.5005
R13544 DVSS.n13487 DVSS.n13480 4.5005
R13545 DVSS.n13491 DVSS.n13480 4.5005
R13546 DVSS.n13486 DVSS.n13480 4.5005
R13547 DVSS.n13492 DVSS.n13480 4.5005
R13548 DVSS.n13485 DVSS.n13480 4.5005
R13549 DVSS.n13493 DVSS.n13480 4.5005
R13550 DVSS.n13484 DVSS.n13480 4.5005
R13551 DVSS.n13494 DVSS.n13480 4.5005
R13552 DVSS.n13483 DVSS.n13480 4.5005
R13553 DVSS.n13495 DVSS.n13480 4.5005
R13554 DVSS.n21338 DVSS.n13480 4.5005
R13555 DVSS.n21340 DVSS.n13480 4.5005
R13556 DVSS.n13488 DVSS.n13466 4.5005
R13557 DVSS.n13489 DVSS.n13466 4.5005
R13558 DVSS.n13487 DVSS.n13466 4.5005
R13559 DVSS.n13491 DVSS.n13466 4.5005
R13560 DVSS.n13486 DVSS.n13466 4.5005
R13561 DVSS.n13492 DVSS.n13466 4.5005
R13562 DVSS.n13485 DVSS.n13466 4.5005
R13563 DVSS.n13493 DVSS.n13466 4.5005
R13564 DVSS.n13484 DVSS.n13466 4.5005
R13565 DVSS.n13494 DVSS.n13466 4.5005
R13566 DVSS.n13483 DVSS.n13466 4.5005
R13567 DVSS.n13495 DVSS.n13466 4.5005
R13568 DVSS.n21338 DVSS.n13466 4.5005
R13569 DVSS.n21340 DVSS.n13466 4.5005
R13570 DVSS.n21339 DVSS.n13488 4.5005
R13571 DVSS.n21339 DVSS.n13489 4.5005
R13572 DVSS.n21339 DVSS.n13487 4.5005
R13573 DVSS.n21339 DVSS.n13491 4.5005
R13574 DVSS.n21339 DVSS.n13486 4.5005
R13575 DVSS.n21339 DVSS.n13492 4.5005
R13576 DVSS.n21339 DVSS.n13485 4.5005
R13577 DVSS.n21339 DVSS.n13493 4.5005
R13578 DVSS.n21339 DVSS.n13484 4.5005
R13579 DVSS.n21339 DVSS.n13494 4.5005
R13580 DVSS.n21339 DVSS.n13483 4.5005
R13581 DVSS.n21339 DVSS.n13495 4.5005
R13582 DVSS.n21339 DVSS.n21338 4.5005
R13583 DVSS.n21339 DVSS.n13465 4.5005
R13584 DVSS.n21340 DVSS.n21339 4.5005
R13585 DVSS.n21076 DVSS.n14031 4.5005
R13586 DVSS.n14075 DVSS.n14031 4.5005
R13587 DVSS.n14073 DVSS.n14031 4.5005
R13588 DVSS.n14078 DVSS.n14031 4.5005
R13589 DVSS.n14071 DVSS.n14031 4.5005
R13590 DVSS.n14079 DVSS.n14031 4.5005
R13591 DVSS.n14070 DVSS.n14031 4.5005
R13592 DVSS.n14080 DVSS.n14031 4.5005
R13593 DVSS.n14069 DVSS.n14031 4.5005
R13594 DVSS.n14083 DVSS.n14031 4.5005
R13595 DVSS.n21074 DVSS.n14031 4.5005
R13596 DVSS.n21076 DVSS.n14033 4.5005
R13597 DVSS.n14075 DVSS.n14033 4.5005
R13598 DVSS.n14073 DVSS.n14033 4.5005
R13599 DVSS.n14077 DVSS.n14033 4.5005
R13600 DVSS.n14072 DVSS.n14033 4.5005
R13601 DVSS.n14078 DVSS.n14033 4.5005
R13602 DVSS.n14071 DVSS.n14033 4.5005
R13603 DVSS.n14079 DVSS.n14033 4.5005
R13604 DVSS.n14070 DVSS.n14033 4.5005
R13605 DVSS.n14080 DVSS.n14033 4.5005
R13606 DVSS.n14069 DVSS.n14033 4.5005
R13607 DVSS.n14082 DVSS.n14033 4.5005
R13608 DVSS.n14083 DVSS.n14033 4.5005
R13609 DVSS.n21074 DVSS.n14033 4.5005
R13610 DVSS.n21076 DVSS.n14030 4.5005
R13611 DVSS.n14075 DVSS.n14030 4.5005
R13612 DVSS.n14073 DVSS.n14030 4.5005
R13613 DVSS.n14077 DVSS.n14030 4.5005
R13614 DVSS.n14072 DVSS.n14030 4.5005
R13615 DVSS.n14078 DVSS.n14030 4.5005
R13616 DVSS.n14071 DVSS.n14030 4.5005
R13617 DVSS.n14079 DVSS.n14030 4.5005
R13618 DVSS.n14070 DVSS.n14030 4.5005
R13619 DVSS.n14080 DVSS.n14030 4.5005
R13620 DVSS.n14069 DVSS.n14030 4.5005
R13621 DVSS.n14082 DVSS.n14030 4.5005
R13622 DVSS.n14083 DVSS.n14030 4.5005
R13623 DVSS.n21074 DVSS.n14030 4.5005
R13624 DVSS.n21076 DVSS.n14034 4.5005
R13625 DVSS.n14075 DVSS.n14034 4.5005
R13626 DVSS.n14073 DVSS.n14034 4.5005
R13627 DVSS.n14077 DVSS.n14034 4.5005
R13628 DVSS.n14072 DVSS.n14034 4.5005
R13629 DVSS.n14078 DVSS.n14034 4.5005
R13630 DVSS.n14071 DVSS.n14034 4.5005
R13631 DVSS.n14079 DVSS.n14034 4.5005
R13632 DVSS.n14070 DVSS.n14034 4.5005
R13633 DVSS.n14080 DVSS.n14034 4.5005
R13634 DVSS.n14069 DVSS.n14034 4.5005
R13635 DVSS.n14082 DVSS.n14034 4.5005
R13636 DVSS.n14083 DVSS.n14034 4.5005
R13637 DVSS.n21074 DVSS.n14034 4.5005
R13638 DVSS.n21076 DVSS.n14029 4.5005
R13639 DVSS.n14075 DVSS.n14029 4.5005
R13640 DVSS.n14073 DVSS.n14029 4.5005
R13641 DVSS.n14077 DVSS.n14029 4.5005
R13642 DVSS.n14072 DVSS.n14029 4.5005
R13643 DVSS.n14078 DVSS.n14029 4.5005
R13644 DVSS.n14071 DVSS.n14029 4.5005
R13645 DVSS.n14079 DVSS.n14029 4.5005
R13646 DVSS.n14070 DVSS.n14029 4.5005
R13647 DVSS.n14080 DVSS.n14029 4.5005
R13648 DVSS.n14069 DVSS.n14029 4.5005
R13649 DVSS.n14082 DVSS.n14029 4.5005
R13650 DVSS.n14083 DVSS.n14029 4.5005
R13651 DVSS.n21074 DVSS.n14029 4.5005
R13652 DVSS.n21076 DVSS.n14035 4.5005
R13653 DVSS.n14075 DVSS.n14035 4.5005
R13654 DVSS.n14073 DVSS.n14035 4.5005
R13655 DVSS.n14077 DVSS.n14035 4.5005
R13656 DVSS.n14072 DVSS.n14035 4.5005
R13657 DVSS.n14078 DVSS.n14035 4.5005
R13658 DVSS.n14071 DVSS.n14035 4.5005
R13659 DVSS.n14079 DVSS.n14035 4.5005
R13660 DVSS.n14070 DVSS.n14035 4.5005
R13661 DVSS.n14080 DVSS.n14035 4.5005
R13662 DVSS.n14069 DVSS.n14035 4.5005
R13663 DVSS.n14082 DVSS.n14035 4.5005
R13664 DVSS.n14083 DVSS.n14035 4.5005
R13665 DVSS.n21074 DVSS.n14035 4.5005
R13666 DVSS.n21076 DVSS.n14028 4.5005
R13667 DVSS.n14075 DVSS.n14028 4.5005
R13668 DVSS.n14073 DVSS.n14028 4.5005
R13669 DVSS.n14077 DVSS.n14028 4.5005
R13670 DVSS.n14072 DVSS.n14028 4.5005
R13671 DVSS.n14078 DVSS.n14028 4.5005
R13672 DVSS.n14071 DVSS.n14028 4.5005
R13673 DVSS.n14079 DVSS.n14028 4.5005
R13674 DVSS.n14070 DVSS.n14028 4.5005
R13675 DVSS.n14080 DVSS.n14028 4.5005
R13676 DVSS.n14069 DVSS.n14028 4.5005
R13677 DVSS.n14082 DVSS.n14028 4.5005
R13678 DVSS.n14083 DVSS.n14028 4.5005
R13679 DVSS.n21074 DVSS.n14028 4.5005
R13680 DVSS.n21076 DVSS.n14036 4.5005
R13681 DVSS.n14075 DVSS.n14036 4.5005
R13682 DVSS.n14073 DVSS.n14036 4.5005
R13683 DVSS.n14077 DVSS.n14036 4.5005
R13684 DVSS.n14072 DVSS.n14036 4.5005
R13685 DVSS.n14078 DVSS.n14036 4.5005
R13686 DVSS.n14071 DVSS.n14036 4.5005
R13687 DVSS.n14079 DVSS.n14036 4.5005
R13688 DVSS.n14070 DVSS.n14036 4.5005
R13689 DVSS.n14080 DVSS.n14036 4.5005
R13690 DVSS.n14069 DVSS.n14036 4.5005
R13691 DVSS.n14082 DVSS.n14036 4.5005
R13692 DVSS.n14083 DVSS.n14036 4.5005
R13693 DVSS.n21074 DVSS.n14036 4.5005
R13694 DVSS.n21076 DVSS.n14027 4.5005
R13695 DVSS.n14075 DVSS.n14027 4.5005
R13696 DVSS.n14073 DVSS.n14027 4.5005
R13697 DVSS.n14077 DVSS.n14027 4.5005
R13698 DVSS.n14072 DVSS.n14027 4.5005
R13699 DVSS.n14078 DVSS.n14027 4.5005
R13700 DVSS.n14071 DVSS.n14027 4.5005
R13701 DVSS.n14079 DVSS.n14027 4.5005
R13702 DVSS.n14070 DVSS.n14027 4.5005
R13703 DVSS.n14080 DVSS.n14027 4.5005
R13704 DVSS.n14069 DVSS.n14027 4.5005
R13705 DVSS.n14082 DVSS.n14027 4.5005
R13706 DVSS.n14083 DVSS.n14027 4.5005
R13707 DVSS.n21074 DVSS.n14027 4.5005
R13708 DVSS.n21076 DVSS.n14037 4.5005
R13709 DVSS.n14075 DVSS.n14037 4.5005
R13710 DVSS.n14073 DVSS.n14037 4.5005
R13711 DVSS.n14077 DVSS.n14037 4.5005
R13712 DVSS.n14072 DVSS.n14037 4.5005
R13713 DVSS.n14078 DVSS.n14037 4.5005
R13714 DVSS.n14071 DVSS.n14037 4.5005
R13715 DVSS.n14079 DVSS.n14037 4.5005
R13716 DVSS.n14070 DVSS.n14037 4.5005
R13717 DVSS.n14080 DVSS.n14037 4.5005
R13718 DVSS.n14069 DVSS.n14037 4.5005
R13719 DVSS.n14082 DVSS.n14037 4.5005
R13720 DVSS.n14083 DVSS.n14037 4.5005
R13721 DVSS.n21074 DVSS.n14037 4.5005
R13722 DVSS.n21076 DVSS.n14026 4.5005
R13723 DVSS.n14075 DVSS.n14026 4.5005
R13724 DVSS.n14073 DVSS.n14026 4.5005
R13725 DVSS.n14077 DVSS.n14026 4.5005
R13726 DVSS.n14072 DVSS.n14026 4.5005
R13727 DVSS.n14078 DVSS.n14026 4.5005
R13728 DVSS.n14071 DVSS.n14026 4.5005
R13729 DVSS.n14079 DVSS.n14026 4.5005
R13730 DVSS.n14070 DVSS.n14026 4.5005
R13731 DVSS.n14080 DVSS.n14026 4.5005
R13732 DVSS.n14069 DVSS.n14026 4.5005
R13733 DVSS.n14082 DVSS.n14026 4.5005
R13734 DVSS.n14083 DVSS.n14026 4.5005
R13735 DVSS.n21074 DVSS.n14026 4.5005
R13736 DVSS.n21076 DVSS.n14038 4.5005
R13737 DVSS.n14075 DVSS.n14038 4.5005
R13738 DVSS.n14073 DVSS.n14038 4.5005
R13739 DVSS.n14077 DVSS.n14038 4.5005
R13740 DVSS.n14072 DVSS.n14038 4.5005
R13741 DVSS.n14078 DVSS.n14038 4.5005
R13742 DVSS.n14071 DVSS.n14038 4.5005
R13743 DVSS.n14079 DVSS.n14038 4.5005
R13744 DVSS.n14070 DVSS.n14038 4.5005
R13745 DVSS.n14080 DVSS.n14038 4.5005
R13746 DVSS.n14069 DVSS.n14038 4.5005
R13747 DVSS.n14082 DVSS.n14038 4.5005
R13748 DVSS.n14083 DVSS.n14038 4.5005
R13749 DVSS.n21074 DVSS.n14038 4.5005
R13750 DVSS.n21076 DVSS.n14025 4.5005
R13751 DVSS.n14075 DVSS.n14025 4.5005
R13752 DVSS.n14073 DVSS.n14025 4.5005
R13753 DVSS.n14077 DVSS.n14025 4.5005
R13754 DVSS.n14072 DVSS.n14025 4.5005
R13755 DVSS.n14078 DVSS.n14025 4.5005
R13756 DVSS.n14071 DVSS.n14025 4.5005
R13757 DVSS.n14079 DVSS.n14025 4.5005
R13758 DVSS.n14070 DVSS.n14025 4.5005
R13759 DVSS.n14080 DVSS.n14025 4.5005
R13760 DVSS.n14069 DVSS.n14025 4.5005
R13761 DVSS.n14082 DVSS.n14025 4.5005
R13762 DVSS.n14083 DVSS.n14025 4.5005
R13763 DVSS.n21074 DVSS.n14025 4.5005
R13764 DVSS.n21076 DVSS.n14039 4.5005
R13765 DVSS.n14075 DVSS.n14039 4.5005
R13766 DVSS.n14073 DVSS.n14039 4.5005
R13767 DVSS.n14077 DVSS.n14039 4.5005
R13768 DVSS.n14072 DVSS.n14039 4.5005
R13769 DVSS.n14078 DVSS.n14039 4.5005
R13770 DVSS.n14071 DVSS.n14039 4.5005
R13771 DVSS.n14079 DVSS.n14039 4.5005
R13772 DVSS.n14070 DVSS.n14039 4.5005
R13773 DVSS.n14080 DVSS.n14039 4.5005
R13774 DVSS.n14069 DVSS.n14039 4.5005
R13775 DVSS.n14082 DVSS.n14039 4.5005
R13776 DVSS.n14083 DVSS.n14039 4.5005
R13777 DVSS.n21074 DVSS.n14039 4.5005
R13778 DVSS.n21076 DVSS.n14024 4.5005
R13779 DVSS.n14075 DVSS.n14024 4.5005
R13780 DVSS.n14073 DVSS.n14024 4.5005
R13781 DVSS.n14077 DVSS.n14024 4.5005
R13782 DVSS.n14072 DVSS.n14024 4.5005
R13783 DVSS.n14078 DVSS.n14024 4.5005
R13784 DVSS.n14071 DVSS.n14024 4.5005
R13785 DVSS.n14079 DVSS.n14024 4.5005
R13786 DVSS.n14070 DVSS.n14024 4.5005
R13787 DVSS.n14080 DVSS.n14024 4.5005
R13788 DVSS.n14069 DVSS.n14024 4.5005
R13789 DVSS.n14082 DVSS.n14024 4.5005
R13790 DVSS.n14083 DVSS.n14024 4.5005
R13791 DVSS.n21074 DVSS.n14024 4.5005
R13792 DVSS.n21076 DVSS.n14040 4.5005
R13793 DVSS.n14075 DVSS.n14040 4.5005
R13794 DVSS.n14073 DVSS.n14040 4.5005
R13795 DVSS.n14077 DVSS.n14040 4.5005
R13796 DVSS.n14072 DVSS.n14040 4.5005
R13797 DVSS.n14078 DVSS.n14040 4.5005
R13798 DVSS.n14071 DVSS.n14040 4.5005
R13799 DVSS.n14079 DVSS.n14040 4.5005
R13800 DVSS.n14070 DVSS.n14040 4.5005
R13801 DVSS.n14080 DVSS.n14040 4.5005
R13802 DVSS.n14069 DVSS.n14040 4.5005
R13803 DVSS.n14082 DVSS.n14040 4.5005
R13804 DVSS.n14083 DVSS.n14040 4.5005
R13805 DVSS.n21074 DVSS.n14040 4.5005
R13806 DVSS.n21076 DVSS.n14023 4.5005
R13807 DVSS.n14075 DVSS.n14023 4.5005
R13808 DVSS.n14073 DVSS.n14023 4.5005
R13809 DVSS.n14077 DVSS.n14023 4.5005
R13810 DVSS.n14072 DVSS.n14023 4.5005
R13811 DVSS.n14078 DVSS.n14023 4.5005
R13812 DVSS.n14071 DVSS.n14023 4.5005
R13813 DVSS.n14079 DVSS.n14023 4.5005
R13814 DVSS.n14070 DVSS.n14023 4.5005
R13815 DVSS.n14080 DVSS.n14023 4.5005
R13816 DVSS.n14069 DVSS.n14023 4.5005
R13817 DVSS.n14082 DVSS.n14023 4.5005
R13818 DVSS.n14083 DVSS.n14023 4.5005
R13819 DVSS.n21074 DVSS.n14023 4.5005
R13820 DVSS.n21076 DVSS.n14041 4.5005
R13821 DVSS.n14075 DVSS.n14041 4.5005
R13822 DVSS.n14073 DVSS.n14041 4.5005
R13823 DVSS.n14077 DVSS.n14041 4.5005
R13824 DVSS.n14072 DVSS.n14041 4.5005
R13825 DVSS.n14078 DVSS.n14041 4.5005
R13826 DVSS.n14071 DVSS.n14041 4.5005
R13827 DVSS.n14079 DVSS.n14041 4.5005
R13828 DVSS.n14070 DVSS.n14041 4.5005
R13829 DVSS.n14080 DVSS.n14041 4.5005
R13830 DVSS.n14069 DVSS.n14041 4.5005
R13831 DVSS.n14082 DVSS.n14041 4.5005
R13832 DVSS.n14083 DVSS.n14041 4.5005
R13833 DVSS.n21074 DVSS.n14041 4.5005
R13834 DVSS.n21076 DVSS.n14022 4.5005
R13835 DVSS.n14075 DVSS.n14022 4.5005
R13836 DVSS.n14073 DVSS.n14022 4.5005
R13837 DVSS.n14077 DVSS.n14022 4.5005
R13838 DVSS.n14072 DVSS.n14022 4.5005
R13839 DVSS.n14078 DVSS.n14022 4.5005
R13840 DVSS.n14071 DVSS.n14022 4.5005
R13841 DVSS.n14079 DVSS.n14022 4.5005
R13842 DVSS.n14070 DVSS.n14022 4.5005
R13843 DVSS.n14080 DVSS.n14022 4.5005
R13844 DVSS.n14069 DVSS.n14022 4.5005
R13845 DVSS.n14082 DVSS.n14022 4.5005
R13846 DVSS.n14083 DVSS.n14022 4.5005
R13847 DVSS.n21074 DVSS.n14022 4.5005
R13848 DVSS.n21076 DVSS.n14042 4.5005
R13849 DVSS.n14075 DVSS.n14042 4.5005
R13850 DVSS.n14073 DVSS.n14042 4.5005
R13851 DVSS.n14077 DVSS.n14042 4.5005
R13852 DVSS.n14072 DVSS.n14042 4.5005
R13853 DVSS.n14078 DVSS.n14042 4.5005
R13854 DVSS.n14071 DVSS.n14042 4.5005
R13855 DVSS.n14079 DVSS.n14042 4.5005
R13856 DVSS.n14070 DVSS.n14042 4.5005
R13857 DVSS.n14080 DVSS.n14042 4.5005
R13858 DVSS.n14069 DVSS.n14042 4.5005
R13859 DVSS.n14082 DVSS.n14042 4.5005
R13860 DVSS.n14083 DVSS.n14042 4.5005
R13861 DVSS.n21074 DVSS.n14042 4.5005
R13862 DVSS.n21076 DVSS.n14021 4.5005
R13863 DVSS.n14075 DVSS.n14021 4.5005
R13864 DVSS.n14073 DVSS.n14021 4.5005
R13865 DVSS.n14077 DVSS.n14021 4.5005
R13866 DVSS.n14072 DVSS.n14021 4.5005
R13867 DVSS.n14078 DVSS.n14021 4.5005
R13868 DVSS.n14071 DVSS.n14021 4.5005
R13869 DVSS.n14079 DVSS.n14021 4.5005
R13870 DVSS.n14070 DVSS.n14021 4.5005
R13871 DVSS.n14080 DVSS.n14021 4.5005
R13872 DVSS.n14069 DVSS.n14021 4.5005
R13873 DVSS.n14082 DVSS.n14021 4.5005
R13874 DVSS.n14083 DVSS.n14021 4.5005
R13875 DVSS.n21074 DVSS.n14021 4.5005
R13876 DVSS.n21076 DVSS.n14043 4.5005
R13877 DVSS.n14075 DVSS.n14043 4.5005
R13878 DVSS.n14073 DVSS.n14043 4.5005
R13879 DVSS.n14077 DVSS.n14043 4.5005
R13880 DVSS.n14072 DVSS.n14043 4.5005
R13881 DVSS.n14078 DVSS.n14043 4.5005
R13882 DVSS.n14071 DVSS.n14043 4.5005
R13883 DVSS.n14079 DVSS.n14043 4.5005
R13884 DVSS.n14070 DVSS.n14043 4.5005
R13885 DVSS.n14080 DVSS.n14043 4.5005
R13886 DVSS.n14069 DVSS.n14043 4.5005
R13887 DVSS.n14082 DVSS.n14043 4.5005
R13888 DVSS.n14083 DVSS.n14043 4.5005
R13889 DVSS.n21074 DVSS.n14043 4.5005
R13890 DVSS.n21076 DVSS.n14020 4.5005
R13891 DVSS.n14075 DVSS.n14020 4.5005
R13892 DVSS.n14073 DVSS.n14020 4.5005
R13893 DVSS.n14077 DVSS.n14020 4.5005
R13894 DVSS.n14072 DVSS.n14020 4.5005
R13895 DVSS.n14078 DVSS.n14020 4.5005
R13896 DVSS.n14071 DVSS.n14020 4.5005
R13897 DVSS.n14079 DVSS.n14020 4.5005
R13898 DVSS.n14070 DVSS.n14020 4.5005
R13899 DVSS.n14080 DVSS.n14020 4.5005
R13900 DVSS.n14069 DVSS.n14020 4.5005
R13901 DVSS.n14082 DVSS.n14020 4.5005
R13902 DVSS.n14083 DVSS.n14020 4.5005
R13903 DVSS.n14056 DVSS.n14020 4.5005
R13904 DVSS.n21074 DVSS.n14020 4.5005
R13905 DVSS.n21076 DVSS.n21075 4.5005
R13906 DVSS.n21075 DVSS.n14075 4.5005
R13907 DVSS.n21075 DVSS.n14073 4.5005
R13908 DVSS.n21075 DVSS.n14077 4.5005
R13909 DVSS.n21075 DVSS.n14072 4.5005
R13910 DVSS.n21075 DVSS.n14078 4.5005
R13911 DVSS.n21075 DVSS.n14071 4.5005
R13912 DVSS.n21075 DVSS.n14079 4.5005
R13913 DVSS.n21075 DVSS.n14070 4.5005
R13914 DVSS.n21075 DVSS.n14080 4.5005
R13915 DVSS.n21075 DVSS.n14069 4.5005
R13916 DVSS.n21075 DVSS.n14082 4.5005
R13917 DVSS.n21075 DVSS.n14068 4.5005
R13918 DVSS.n21075 DVSS.n14083 4.5005
R13919 DVSS.n21075 DVSS.n14056 4.5005
R13920 DVSS.n21075 DVSS.n21074 4.5005
R13921 DVSS.n14432 DVSS.n14416 4.5005
R13922 DVSS.n14433 DVSS.n14416 4.5005
R13923 DVSS.n14431 DVSS.n14416 4.5005
R13924 DVSS.n14436 DVSS.n14416 4.5005
R13925 DVSS.n14429 DVSS.n14416 4.5005
R13926 DVSS.n14437 DVSS.n14416 4.5005
R13927 DVSS.n14428 DVSS.n14416 4.5005
R13928 DVSS.n14438 DVSS.n14416 4.5005
R13929 DVSS.n14427 DVSS.n14416 4.5005
R13930 DVSS.n20888 DVSS.n14416 4.5005
R13931 DVSS.n14416 DVSS.n14410 4.5005
R13932 DVSS.n20890 DVSS.n14416 4.5005
R13933 DVSS.n14432 DVSS.n14415 4.5005
R13934 DVSS.n14433 DVSS.n14415 4.5005
R13935 DVSS.n14431 DVSS.n14415 4.5005
R13936 DVSS.n14435 DVSS.n14415 4.5005
R13937 DVSS.n14430 DVSS.n14415 4.5005
R13938 DVSS.n14436 DVSS.n14415 4.5005
R13939 DVSS.n14429 DVSS.n14415 4.5005
R13940 DVSS.n14437 DVSS.n14415 4.5005
R13941 DVSS.n14428 DVSS.n14415 4.5005
R13942 DVSS.n14438 DVSS.n14415 4.5005
R13943 DVSS.n14427 DVSS.n14415 4.5005
R13944 DVSS.n14439 DVSS.n14415 4.5005
R13945 DVSS.n14444 DVSS.n14415 4.5005
R13946 DVSS.n20888 DVSS.n14415 4.5005
R13947 DVSS.n14415 DVSS.n14410 4.5005
R13948 DVSS.n20890 DVSS.n14415 4.5005
R13949 DVSS.n14432 DVSS.n14418 4.5005
R13950 DVSS.n14433 DVSS.n14418 4.5005
R13951 DVSS.n14431 DVSS.n14418 4.5005
R13952 DVSS.n14435 DVSS.n14418 4.5005
R13953 DVSS.n14430 DVSS.n14418 4.5005
R13954 DVSS.n14436 DVSS.n14418 4.5005
R13955 DVSS.n14429 DVSS.n14418 4.5005
R13956 DVSS.n14437 DVSS.n14418 4.5005
R13957 DVSS.n14428 DVSS.n14418 4.5005
R13958 DVSS.n14438 DVSS.n14418 4.5005
R13959 DVSS.n14427 DVSS.n14418 4.5005
R13960 DVSS.n14439 DVSS.n14418 4.5005
R13961 DVSS.n14444 DVSS.n14418 4.5005
R13962 DVSS.n20888 DVSS.n14418 4.5005
R13963 DVSS.n20890 DVSS.n14418 4.5005
R13964 DVSS.n14432 DVSS.n14414 4.5005
R13965 DVSS.n14433 DVSS.n14414 4.5005
R13966 DVSS.n14431 DVSS.n14414 4.5005
R13967 DVSS.n14435 DVSS.n14414 4.5005
R13968 DVSS.n14430 DVSS.n14414 4.5005
R13969 DVSS.n14436 DVSS.n14414 4.5005
R13970 DVSS.n14429 DVSS.n14414 4.5005
R13971 DVSS.n14437 DVSS.n14414 4.5005
R13972 DVSS.n14428 DVSS.n14414 4.5005
R13973 DVSS.n14438 DVSS.n14414 4.5005
R13974 DVSS.n14427 DVSS.n14414 4.5005
R13975 DVSS.n14439 DVSS.n14414 4.5005
R13976 DVSS.n20888 DVSS.n14414 4.5005
R13977 DVSS.n20890 DVSS.n14414 4.5005
R13978 DVSS.n14432 DVSS.n14420 4.5005
R13979 DVSS.n14433 DVSS.n14420 4.5005
R13980 DVSS.n14431 DVSS.n14420 4.5005
R13981 DVSS.n14435 DVSS.n14420 4.5005
R13982 DVSS.n14430 DVSS.n14420 4.5005
R13983 DVSS.n14436 DVSS.n14420 4.5005
R13984 DVSS.n14429 DVSS.n14420 4.5005
R13985 DVSS.n14437 DVSS.n14420 4.5005
R13986 DVSS.n14428 DVSS.n14420 4.5005
R13987 DVSS.n14438 DVSS.n14420 4.5005
R13988 DVSS.n14427 DVSS.n14420 4.5005
R13989 DVSS.n14439 DVSS.n14420 4.5005
R13990 DVSS.n20888 DVSS.n14420 4.5005
R13991 DVSS.n20890 DVSS.n14420 4.5005
R13992 DVSS.n14432 DVSS.n14413 4.5005
R13993 DVSS.n14433 DVSS.n14413 4.5005
R13994 DVSS.n14431 DVSS.n14413 4.5005
R13995 DVSS.n14435 DVSS.n14413 4.5005
R13996 DVSS.n14430 DVSS.n14413 4.5005
R13997 DVSS.n14436 DVSS.n14413 4.5005
R13998 DVSS.n14429 DVSS.n14413 4.5005
R13999 DVSS.n14437 DVSS.n14413 4.5005
R14000 DVSS.n14428 DVSS.n14413 4.5005
R14001 DVSS.n14438 DVSS.n14413 4.5005
R14002 DVSS.n14427 DVSS.n14413 4.5005
R14003 DVSS.n14439 DVSS.n14413 4.5005
R14004 DVSS.n20888 DVSS.n14413 4.5005
R14005 DVSS.n20890 DVSS.n14413 4.5005
R14006 DVSS.n14432 DVSS.n14422 4.5005
R14007 DVSS.n14433 DVSS.n14422 4.5005
R14008 DVSS.n14431 DVSS.n14422 4.5005
R14009 DVSS.n14435 DVSS.n14422 4.5005
R14010 DVSS.n14430 DVSS.n14422 4.5005
R14011 DVSS.n14436 DVSS.n14422 4.5005
R14012 DVSS.n14429 DVSS.n14422 4.5005
R14013 DVSS.n14437 DVSS.n14422 4.5005
R14014 DVSS.n14428 DVSS.n14422 4.5005
R14015 DVSS.n14438 DVSS.n14422 4.5005
R14016 DVSS.n14427 DVSS.n14422 4.5005
R14017 DVSS.n14439 DVSS.n14422 4.5005
R14018 DVSS.n20888 DVSS.n14422 4.5005
R14019 DVSS.n20890 DVSS.n14422 4.5005
R14020 DVSS.n14432 DVSS.n14412 4.5005
R14021 DVSS.n14433 DVSS.n14412 4.5005
R14022 DVSS.n14431 DVSS.n14412 4.5005
R14023 DVSS.n14435 DVSS.n14412 4.5005
R14024 DVSS.n14430 DVSS.n14412 4.5005
R14025 DVSS.n14436 DVSS.n14412 4.5005
R14026 DVSS.n14429 DVSS.n14412 4.5005
R14027 DVSS.n14437 DVSS.n14412 4.5005
R14028 DVSS.n14428 DVSS.n14412 4.5005
R14029 DVSS.n14438 DVSS.n14412 4.5005
R14030 DVSS.n14427 DVSS.n14412 4.5005
R14031 DVSS.n14439 DVSS.n14412 4.5005
R14032 DVSS.n20888 DVSS.n14412 4.5005
R14033 DVSS.n20890 DVSS.n14412 4.5005
R14034 DVSS.n14432 DVSS.n14424 4.5005
R14035 DVSS.n14433 DVSS.n14424 4.5005
R14036 DVSS.n14431 DVSS.n14424 4.5005
R14037 DVSS.n14435 DVSS.n14424 4.5005
R14038 DVSS.n14430 DVSS.n14424 4.5005
R14039 DVSS.n14436 DVSS.n14424 4.5005
R14040 DVSS.n14429 DVSS.n14424 4.5005
R14041 DVSS.n14437 DVSS.n14424 4.5005
R14042 DVSS.n14428 DVSS.n14424 4.5005
R14043 DVSS.n14438 DVSS.n14424 4.5005
R14044 DVSS.n14427 DVSS.n14424 4.5005
R14045 DVSS.n14439 DVSS.n14424 4.5005
R14046 DVSS.n20888 DVSS.n14424 4.5005
R14047 DVSS.n20890 DVSS.n14424 4.5005
R14048 DVSS.n14432 DVSS.n14411 4.5005
R14049 DVSS.n14433 DVSS.n14411 4.5005
R14050 DVSS.n14431 DVSS.n14411 4.5005
R14051 DVSS.n14435 DVSS.n14411 4.5005
R14052 DVSS.n14430 DVSS.n14411 4.5005
R14053 DVSS.n14436 DVSS.n14411 4.5005
R14054 DVSS.n14429 DVSS.n14411 4.5005
R14055 DVSS.n14437 DVSS.n14411 4.5005
R14056 DVSS.n14428 DVSS.n14411 4.5005
R14057 DVSS.n14438 DVSS.n14411 4.5005
R14058 DVSS.n14427 DVSS.n14411 4.5005
R14059 DVSS.n14439 DVSS.n14411 4.5005
R14060 DVSS.n20888 DVSS.n14411 4.5005
R14061 DVSS.n20890 DVSS.n14411 4.5005
R14062 DVSS.n20889 DVSS.n14432 4.5005
R14063 DVSS.n20889 DVSS.n14433 4.5005
R14064 DVSS.n20889 DVSS.n14431 4.5005
R14065 DVSS.n20889 DVSS.n14435 4.5005
R14066 DVSS.n20889 DVSS.n14430 4.5005
R14067 DVSS.n20889 DVSS.n14436 4.5005
R14068 DVSS.n20889 DVSS.n14429 4.5005
R14069 DVSS.n20889 DVSS.n14437 4.5005
R14070 DVSS.n20889 DVSS.n14428 4.5005
R14071 DVSS.n20889 DVSS.n14438 4.5005
R14072 DVSS.n20889 DVSS.n14427 4.5005
R14073 DVSS.n20889 DVSS.n14439 4.5005
R14074 DVSS.n20889 DVSS.n20888 4.5005
R14075 DVSS.n20889 DVSS.n14410 4.5005
R14076 DVSS.n20890 DVSS.n20889 4.5005
R14077 DVSS.n14927 DVSS.n14864 4.5005
R14078 DVSS.n19983 DVSS.n14864 4.5005
R14079 DVSS.n14950 DVSS.n14864 4.5005
R14080 DVSS.n14953 DVSS.n14864 4.5005
R14081 DVSS.n14948 DVSS.n14864 4.5005
R14082 DVSS.n14954 DVSS.n14864 4.5005
R14083 DVSS.n14947 DVSS.n14864 4.5005
R14084 DVSS.n14955 DVSS.n14864 4.5005
R14085 DVSS.n14946 DVSS.n14864 4.5005
R14086 DVSS.n14957 DVSS.n14864 4.5005
R14087 DVSS.n19981 DVSS.n14864 4.5005
R14088 DVSS.n14932 DVSS.n14927 4.5005
R14089 DVSS.n19983 DVSS.n14932 4.5005
R14090 DVSS.n14950 DVSS.n14932 4.5005
R14091 DVSS.n14952 DVSS.n14932 4.5005
R14092 DVSS.n14949 DVSS.n14932 4.5005
R14093 DVSS.n14953 DVSS.n14932 4.5005
R14094 DVSS.n14948 DVSS.n14932 4.5005
R14095 DVSS.n14954 DVSS.n14932 4.5005
R14096 DVSS.n14947 DVSS.n14932 4.5005
R14097 DVSS.n14955 DVSS.n14932 4.5005
R14098 DVSS.n14946 DVSS.n14932 4.5005
R14099 DVSS.n14956 DVSS.n14932 4.5005
R14100 DVSS.n14957 DVSS.n14932 4.5005
R14101 DVSS.n19981 DVSS.n14932 4.5005
R14102 DVSS.n14934 DVSS.n14927 4.5005
R14103 DVSS.n19983 DVSS.n14934 4.5005
R14104 DVSS.n14950 DVSS.n14934 4.5005
R14105 DVSS.n14952 DVSS.n14934 4.5005
R14106 DVSS.n14949 DVSS.n14934 4.5005
R14107 DVSS.n14953 DVSS.n14934 4.5005
R14108 DVSS.n14948 DVSS.n14934 4.5005
R14109 DVSS.n14954 DVSS.n14934 4.5005
R14110 DVSS.n14947 DVSS.n14934 4.5005
R14111 DVSS.n14955 DVSS.n14934 4.5005
R14112 DVSS.n14946 DVSS.n14934 4.5005
R14113 DVSS.n14956 DVSS.n14934 4.5005
R14114 DVSS.n14957 DVSS.n14934 4.5005
R14115 DVSS.n19981 DVSS.n14934 4.5005
R14116 DVSS.n14931 DVSS.n14927 4.5005
R14117 DVSS.n19983 DVSS.n14931 4.5005
R14118 DVSS.n14950 DVSS.n14931 4.5005
R14119 DVSS.n14952 DVSS.n14931 4.5005
R14120 DVSS.n14949 DVSS.n14931 4.5005
R14121 DVSS.n14953 DVSS.n14931 4.5005
R14122 DVSS.n14948 DVSS.n14931 4.5005
R14123 DVSS.n14954 DVSS.n14931 4.5005
R14124 DVSS.n14947 DVSS.n14931 4.5005
R14125 DVSS.n14955 DVSS.n14931 4.5005
R14126 DVSS.n14946 DVSS.n14931 4.5005
R14127 DVSS.n14956 DVSS.n14931 4.5005
R14128 DVSS.n14957 DVSS.n14931 4.5005
R14129 DVSS.n19981 DVSS.n14931 4.5005
R14130 DVSS.n14935 DVSS.n14927 4.5005
R14131 DVSS.n19983 DVSS.n14935 4.5005
R14132 DVSS.n14950 DVSS.n14935 4.5005
R14133 DVSS.n14952 DVSS.n14935 4.5005
R14134 DVSS.n14949 DVSS.n14935 4.5005
R14135 DVSS.n14953 DVSS.n14935 4.5005
R14136 DVSS.n14948 DVSS.n14935 4.5005
R14137 DVSS.n14954 DVSS.n14935 4.5005
R14138 DVSS.n14947 DVSS.n14935 4.5005
R14139 DVSS.n14955 DVSS.n14935 4.5005
R14140 DVSS.n14946 DVSS.n14935 4.5005
R14141 DVSS.n14956 DVSS.n14935 4.5005
R14142 DVSS.n14957 DVSS.n14935 4.5005
R14143 DVSS.n19981 DVSS.n14935 4.5005
R14144 DVSS.n14930 DVSS.n14927 4.5005
R14145 DVSS.n19983 DVSS.n14930 4.5005
R14146 DVSS.n14950 DVSS.n14930 4.5005
R14147 DVSS.n14952 DVSS.n14930 4.5005
R14148 DVSS.n14949 DVSS.n14930 4.5005
R14149 DVSS.n14953 DVSS.n14930 4.5005
R14150 DVSS.n14948 DVSS.n14930 4.5005
R14151 DVSS.n14954 DVSS.n14930 4.5005
R14152 DVSS.n14947 DVSS.n14930 4.5005
R14153 DVSS.n14955 DVSS.n14930 4.5005
R14154 DVSS.n14946 DVSS.n14930 4.5005
R14155 DVSS.n14956 DVSS.n14930 4.5005
R14156 DVSS.n14957 DVSS.n14930 4.5005
R14157 DVSS.n19981 DVSS.n14930 4.5005
R14158 DVSS.n14936 DVSS.n14927 4.5005
R14159 DVSS.n19983 DVSS.n14936 4.5005
R14160 DVSS.n14950 DVSS.n14936 4.5005
R14161 DVSS.n14952 DVSS.n14936 4.5005
R14162 DVSS.n14949 DVSS.n14936 4.5005
R14163 DVSS.n14953 DVSS.n14936 4.5005
R14164 DVSS.n14948 DVSS.n14936 4.5005
R14165 DVSS.n14954 DVSS.n14936 4.5005
R14166 DVSS.n14947 DVSS.n14936 4.5005
R14167 DVSS.n14955 DVSS.n14936 4.5005
R14168 DVSS.n14946 DVSS.n14936 4.5005
R14169 DVSS.n14956 DVSS.n14936 4.5005
R14170 DVSS.n14957 DVSS.n14936 4.5005
R14171 DVSS.n19981 DVSS.n14936 4.5005
R14172 DVSS.n14929 DVSS.n14927 4.5005
R14173 DVSS.n19983 DVSS.n14929 4.5005
R14174 DVSS.n14950 DVSS.n14929 4.5005
R14175 DVSS.n14952 DVSS.n14929 4.5005
R14176 DVSS.n14949 DVSS.n14929 4.5005
R14177 DVSS.n14953 DVSS.n14929 4.5005
R14178 DVSS.n14948 DVSS.n14929 4.5005
R14179 DVSS.n14954 DVSS.n14929 4.5005
R14180 DVSS.n14947 DVSS.n14929 4.5005
R14181 DVSS.n14955 DVSS.n14929 4.5005
R14182 DVSS.n14946 DVSS.n14929 4.5005
R14183 DVSS.n14956 DVSS.n14929 4.5005
R14184 DVSS.n14957 DVSS.n14929 4.5005
R14185 DVSS.n19981 DVSS.n14929 4.5005
R14186 DVSS.n14937 DVSS.n14927 4.5005
R14187 DVSS.n19983 DVSS.n14937 4.5005
R14188 DVSS.n14950 DVSS.n14937 4.5005
R14189 DVSS.n14952 DVSS.n14937 4.5005
R14190 DVSS.n14949 DVSS.n14937 4.5005
R14191 DVSS.n14953 DVSS.n14937 4.5005
R14192 DVSS.n14948 DVSS.n14937 4.5005
R14193 DVSS.n14954 DVSS.n14937 4.5005
R14194 DVSS.n14947 DVSS.n14937 4.5005
R14195 DVSS.n14955 DVSS.n14937 4.5005
R14196 DVSS.n14946 DVSS.n14937 4.5005
R14197 DVSS.n14956 DVSS.n14937 4.5005
R14198 DVSS.n14957 DVSS.n14937 4.5005
R14199 DVSS.n19981 DVSS.n14937 4.5005
R14200 DVSS.n14928 DVSS.n14927 4.5005
R14201 DVSS.n19983 DVSS.n14928 4.5005
R14202 DVSS.n14950 DVSS.n14928 4.5005
R14203 DVSS.n14952 DVSS.n14928 4.5005
R14204 DVSS.n14949 DVSS.n14928 4.5005
R14205 DVSS.n14953 DVSS.n14928 4.5005
R14206 DVSS.n14948 DVSS.n14928 4.5005
R14207 DVSS.n14954 DVSS.n14928 4.5005
R14208 DVSS.n14947 DVSS.n14928 4.5005
R14209 DVSS.n14955 DVSS.n14928 4.5005
R14210 DVSS.n14946 DVSS.n14928 4.5005
R14211 DVSS.n14956 DVSS.n14928 4.5005
R14212 DVSS.n14957 DVSS.n14928 4.5005
R14213 DVSS.n19981 DVSS.n14928 4.5005
R14214 DVSS.n19982 DVSS.n14927 4.5005
R14215 DVSS.n19983 DVSS.n19982 4.5005
R14216 DVSS.n19982 DVSS.n14950 4.5005
R14217 DVSS.n19982 DVSS.n14952 4.5005
R14218 DVSS.n19982 DVSS.n14949 4.5005
R14219 DVSS.n19982 DVSS.n14953 4.5005
R14220 DVSS.n19982 DVSS.n14948 4.5005
R14221 DVSS.n19982 DVSS.n14954 4.5005
R14222 DVSS.n19982 DVSS.n14947 4.5005
R14223 DVSS.n19982 DVSS.n14955 4.5005
R14224 DVSS.n19982 DVSS.n14946 4.5005
R14225 DVSS.n19982 DVSS.n14956 4.5005
R14226 DVSS.n19982 DVSS.n14957 4.5005
R14227 DVSS.n19982 DVSS.n14944 4.5005
R14228 DVSS.n19982 DVSS.n19981 4.5005
R14229 DVSS.n15362 DVSS.n14938 4.5005
R14230 DVSS.n18327 DVSS.n14938 4.5005
R14231 DVSS.n15386 DVSS.n14938 4.5005
R14232 DVSS.n15390 DVSS.n14938 4.5005
R14233 DVSS.n15384 DVSS.n14938 4.5005
R14234 DVSS.n15391 DVSS.n14938 4.5005
R14235 DVSS.n15383 DVSS.n14938 4.5005
R14236 DVSS.n15392 DVSS.n14938 4.5005
R14237 DVSS.n15382 DVSS.n14938 4.5005
R14238 DVSS.n15395 DVSS.n14938 4.5005
R14239 DVSS.n18325 DVSS.n14938 4.5005
R14240 DVSS.n15367 DVSS.n15362 4.5005
R14241 DVSS.n18327 DVSS.n15367 4.5005
R14242 DVSS.n15386 DVSS.n15367 4.5005
R14243 DVSS.n15389 DVSS.n15367 4.5005
R14244 DVSS.n15385 DVSS.n15367 4.5005
R14245 DVSS.n15390 DVSS.n15367 4.5005
R14246 DVSS.n15384 DVSS.n15367 4.5005
R14247 DVSS.n15391 DVSS.n15367 4.5005
R14248 DVSS.n15383 DVSS.n15367 4.5005
R14249 DVSS.n15392 DVSS.n15367 4.5005
R14250 DVSS.n15382 DVSS.n15367 4.5005
R14251 DVSS.n15394 DVSS.n15367 4.5005
R14252 DVSS.n15381 DVSS.n15367 4.5005
R14253 DVSS.n15395 DVSS.n15367 4.5005
R14254 DVSS.n18325 DVSS.n15367 4.5005
R14255 DVSS.n15369 DVSS.n15362 4.5005
R14256 DVSS.n18327 DVSS.n15369 4.5005
R14257 DVSS.n15386 DVSS.n15369 4.5005
R14258 DVSS.n15389 DVSS.n15369 4.5005
R14259 DVSS.n15385 DVSS.n15369 4.5005
R14260 DVSS.n15390 DVSS.n15369 4.5005
R14261 DVSS.n15384 DVSS.n15369 4.5005
R14262 DVSS.n15391 DVSS.n15369 4.5005
R14263 DVSS.n15383 DVSS.n15369 4.5005
R14264 DVSS.n15392 DVSS.n15369 4.5005
R14265 DVSS.n15382 DVSS.n15369 4.5005
R14266 DVSS.n15394 DVSS.n15369 4.5005
R14267 DVSS.n15395 DVSS.n15369 4.5005
R14268 DVSS.n18325 DVSS.n15369 4.5005
R14269 DVSS.n15366 DVSS.n15362 4.5005
R14270 DVSS.n18327 DVSS.n15366 4.5005
R14271 DVSS.n15386 DVSS.n15366 4.5005
R14272 DVSS.n15389 DVSS.n15366 4.5005
R14273 DVSS.n15385 DVSS.n15366 4.5005
R14274 DVSS.n15390 DVSS.n15366 4.5005
R14275 DVSS.n15384 DVSS.n15366 4.5005
R14276 DVSS.n15391 DVSS.n15366 4.5005
R14277 DVSS.n15383 DVSS.n15366 4.5005
R14278 DVSS.n15392 DVSS.n15366 4.5005
R14279 DVSS.n15382 DVSS.n15366 4.5005
R14280 DVSS.n15394 DVSS.n15366 4.5005
R14281 DVSS.n15395 DVSS.n15366 4.5005
R14282 DVSS.n18325 DVSS.n15366 4.5005
R14283 DVSS.n15370 DVSS.n15362 4.5005
R14284 DVSS.n18327 DVSS.n15370 4.5005
R14285 DVSS.n15386 DVSS.n15370 4.5005
R14286 DVSS.n15389 DVSS.n15370 4.5005
R14287 DVSS.n15385 DVSS.n15370 4.5005
R14288 DVSS.n15390 DVSS.n15370 4.5005
R14289 DVSS.n15384 DVSS.n15370 4.5005
R14290 DVSS.n15391 DVSS.n15370 4.5005
R14291 DVSS.n15383 DVSS.n15370 4.5005
R14292 DVSS.n15392 DVSS.n15370 4.5005
R14293 DVSS.n15382 DVSS.n15370 4.5005
R14294 DVSS.n15394 DVSS.n15370 4.5005
R14295 DVSS.n15395 DVSS.n15370 4.5005
R14296 DVSS.n18325 DVSS.n15370 4.5005
R14297 DVSS.n15365 DVSS.n15362 4.5005
R14298 DVSS.n18327 DVSS.n15365 4.5005
R14299 DVSS.n15386 DVSS.n15365 4.5005
R14300 DVSS.n15389 DVSS.n15365 4.5005
R14301 DVSS.n15385 DVSS.n15365 4.5005
R14302 DVSS.n15390 DVSS.n15365 4.5005
R14303 DVSS.n15384 DVSS.n15365 4.5005
R14304 DVSS.n15391 DVSS.n15365 4.5005
R14305 DVSS.n15383 DVSS.n15365 4.5005
R14306 DVSS.n15392 DVSS.n15365 4.5005
R14307 DVSS.n15382 DVSS.n15365 4.5005
R14308 DVSS.n15394 DVSS.n15365 4.5005
R14309 DVSS.n15395 DVSS.n15365 4.5005
R14310 DVSS.n18325 DVSS.n15365 4.5005
R14311 DVSS.n15371 DVSS.n15362 4.5005
R14312 DVSS.n18327 DVSS.n15371 4.5005
R14313 DVSS.n15386 DVSS.n15371 4.5005
R14314 DVSS.n15389 DVSS.n15371 4.5005
R14315 DVSS.n15385 DVSS.n15371 4.5005
R14316 DVSS.n15390 DVSS.n15371 4.5005
R14317 DVSS.n15384 DVSS.n15371 4.5005
R14318 DVSS.n15391 DVSS.n15371 4.5005
R14319 DVSS.n15383 DVSS.n15371 4.5005
R14320 DVSS.n15392 DVSS.n15371 4.5005
R14321 DVSS.n15382 DVSS.n15371 4.5005
R14322 DVSS.n15394 DVSS.n15371 4.5005
R14323 DVSS.n15395 DVSS.n15371 4.5005
R14324 DVSS.n15377 DVSS.n15371 4.5005
R14325 DVSS.n18325 DVSS.n15371 4.5005
R14326 DVSS.n15364 DVSS.n15362 4.5005
R14327 DVSS.n18327 DVSS.n15364 4.5005
R14328 DVSS.n15386 DVSS.n15364 4.5005
R14329 DVSS.n15389 DVSS.n15364 4.5005
R14330 DVSS.n15385 DVSS.n15364 4.5005
R14331 DVSS.n15390 DVSS.n15364 4.5005
R14332 DVSS.n15384 DVSS.n15364 4.5005
R14333 DVSS.n15391 DVSS.n15364 4.5005
R14334 DVSS.n15383 DVSS.n15364 4.5005
R14335 DVSS.n15392 DVSS.n15364 4.5005
R14336 DVSS.n15382 DVSS.n15364 4.5005
R14337 DVSS.n15394 DVSS.n15364 4.5005
R14338 DVSS.n15381 DVSS.n15364 4.5005
R14339 DVSS.n15395 DVSS.n15364 4.5005
R14340 DVSS.n15377 DVSS.n15364 4.5005
R14341 DVSS.n18325 DVSS.n15364 4.5005
R14342 DVSS.n16148 DVSS.n16141 4.5005
R14343 DVSS.n17617 DVSS.n16148 4.5005
R14344 DVSS.n16842 DVSS.n16148 4.5005
R14345 DVSS.n16846 DVSS.n16148 4.5005
R14346 DVSS.n16840 DVSS.n16148 4.5005
R14347 DVSS.n16847 DVSS.n16148 4.5005
R14348 DVSS.n16839 DVSS.n16148 4.5005
R14349 DVSS.n16848 DVSS.n16148 4.5005
R14350 DVSS.n16838 DVSS.n16148 4.5005
R14351 DVSS.n16851 DVSS.n16148 4.5005
R14352 DVSS.n17615 DVSS.n16148 4.5005
R14353 DVSS.n16146 DVSS.n16141 4.5005
R14354 DVSS.n17617 DVSS.n16146 4.5005
R14355 DVSS.n16842 DVSS.n16146 4.5005
R14356 DVSS.n16845 DVSS.n16146 4.5005
R14357 DVSS.n16841 DVSS.n16146 4.5005
R14358 DVSS.n16846 DVSS.n16146 4.5005
R14359 DVSS.n16840 DVSS.n16146 4.5005
R14360 DVSS.n16847 DVSS.n16146 4.5005
R14361 DVSS.n16839 DVSS.n16146 4.5005
R14362 DVSS.n16848 DVSS.n16146 4.5005
R14363 DVSS.n16838 DVSS.n16146 4.5005
R14364 DVSS.n16850 DVSS.n16146 4.5005
R14365 DVSS.n16851 DVSS.n16146 4.5005
R14366 DVSS.n17615 DVSS.n16146 4.5005
R14367 DVSS.n16149 DVSS.n16141 4.5005
R14368 DVSS.n17617 DVSS.n16149 4.5005
R14369 DVSS.n16842 DVSS.n16149 4.5005
R14370 DVSS.n16845 DVSS.n16149 4.5005
R14371 DVSS.n16841 DVSS.n16149 4.5005
R14372 DVSS.n16846 DVSS.n16149 4.5005
R14373 DVSS.n16840 DVSS.n16149 4.5005
R14374 DVSS.n16847 DVSS.n16149 4.5005
R14375 DVSS.n16839 DVSS.n16149 4.5005
R14376 DVSS.n16848 DVSS.n16149 4.5005
R14377 DVSS.n16838 DVSS.n16149 4.5005
R14378 DVSS.n16850 DVSS.n16149 4.5005
R14379 DVSS.n16851 DVSS.n16149 4.5005
R14380 DVSS.n17615 DVSS.n16149 4.5005
R14381 DVSS.n16145 DVSS.n16141 4.5005
R14382 DVSS.n17617 DVSS.n16145 4.5005
R14383 DVSS.n16842 DVSS.n16145 4.5005
R14384 DVSS.n16845 DVSS.n16145 4.5005
R14385 DVSS.n16841 DVSS.n16145 4.5005
R14386 DVSS.n16846 DVSS.n16145 4.5005
R14387 DVSS.n16840 DVSS.n16145 4.5005
R14388 DVSS.n16847 DVSS.n16145 4.5005
R14389 DVSS.n16839 DVSS.n16145 4.5005
R14390 DVSS.n16848 DVSS.n16145 4.5005
R14391 DVSS.n16838 DVSS.n16145 4.5005
R14392 DVSS.n16850 DVSS.n16145 4.5005
R14393 DVSS.n16851 DVSS.n16145 4.5005
R14394 DVSS.n17615 DVSS.n16145 4.5005
R14395 DVSS.n16150 DVSS.n16141 4.5005
R14396 DVSS.n17617 DVSS.n16150 4.5005
R14397 DVSS.n16842 DVSS.n16150 4.5005
R14398 DVSS.n16845 DVSS.n16150 4.5005
R14399 DVSS.n16841 DVSS.n16150 4.5005
R14400 DVSS.n16846 DVSS.n16150 4.5005
R14401 DVSS.n16840 DVSS.n16150 4.5005
R14402 DVSS.n16847 DVSS.n16150 4.5005
R14403 DVSS.n16839 DVSS.n16150 4.5005
R14404 DVSS.n16848 DVSS.n16150 4.5005
R14405 DVSS.n16838 DVSS.n16150 4.5005
R14406 DVSS.n16850 DVSS.n16150 4.5005
R14407 DVSS.n16851 DVSS.n16150 4.5005
R14408 DVSS.n16832 DVSS.n16150 4.5005
R14409 DVSS.n17615 DVSS.n16150 4.5005
R14410 DVSS.n16144 DVSS.n16141 4.5005
R14411 DVSS.n17617 DVSS.n16144 4.5005
R14412 DVSS.n16842 DVSS.n16144 4.5005
R14413 DVSS.n16845 DVSS.n16144 4.5005
R14414 DVSS.n16841 DVSS.n16144 4.5005
R14415 DVSS.n16846 DVSS.n16144 4.5005
R14416 DVSS.n16840 DVSS.n16144 4.5005
R14417 DVSS.n16847 DVSS.n16144 4.5005
R14418 DVSS.n16839 DVSS.n16144 4.5005
R14419 DVSS.n16848 DVSS.n16144 4.5005
R14420 DVSS.n16838 DVSS.n16144 4.5005
R14421 DVSS.n16850 DVSS.n16144 4.5005
R14422 DVSS.n16851 DVSS.n16144 4.5005
R14423 DVSS.n17615 DVSS.n16144 4.5005
R14424 DVSS.n16151 DVSS.n16141 4.5005
R14425 DVSS.n17617 DVSS.n16151 4.5005
R14426 DVSS.n16842 DVSS.n16151 4.5005
R14427 DVSS.n16845 DVSS.n16151 4.5005
R14428 DVSS.n16841 DVSS.n16151 4.5005
R14429 DVSS.n16846 DVSS.n16151 4.5005
R14430 DVSS.n16840 DVSS.n16151 4.5005
R14431 DVSS.n16847 DVSS.n16151 4.5005
R14432 DVSS.n16839 DVSS.n16151 4.5005
R14433 DVSS.n16848 DVSS.n16151 4.5005
R14434 DVSS.n16838 DVSS.n16151 4.5005
R14435 DVSS.n16850 DVSS.n16151 4.5005
R14436 DVSS.n16851 DVSS.n16151 4.5005
R14437 DVSS.n17615 DVSS.n16151 4.5005
R14438 DVSS.n16143 DVSS.n16141 4.5005
R14439 DVSS.n17617 DVSS.n16143 4.5005
R14440 DVSS.n16842 DVSS.n16143 4.5005
R14441 DVSS.n16845 DVSS.n16143 4.5005
R14442 DVSS.n16841 DVSS.n16143 4.5005
R14443 DVSS.n16846 DVSS.n16143 4.5005
R14444 DVSS.n16840 DVSS.n16143 4.5005
R14445 DVSS.n16847 DVSS.n16143 4.5005
R14446 DVSS.n16839 DVSS.n16143 4.5005
R14447 DVSS.n16848 DVSS.n16143 4.5005
R14448 DVSS.n16838 DVSS.n16143 4.5005
R14449 DVSS.n16850 DVSS.n16143 4.5005
R14450 DVSS.n16851 DVSS.n16143 4.5005
R14451 DVSS.n17615 DVSS.n16143 4.5005
R14452 DVSS.n16826 DVSS.n16141 4.5005
R14453 DVSS.n17617 DVSS.n16826 4.5005
R14454 DVSS.n16842 DVSS.n16826 4.5005
R14455 DVSS.n16845 DVSS.n16826 4.5005
R14456 DVSS.n16841 DVSS.n16826 4.5005
R14457 DVSS.n16846 DVSS.n16826 4.5005
R14458 DVSS.n16840 DVSS.n16826 4.5005
R14459 DVSS.n16847 DVSS.n16826 4.5005
R14460 DVSS.n16839 DVSS.n16826 4.5005
R14461 DVSS.n16848 DVSS.n16826 4.5005
R14462 DVSS.n16838 DVSS.n16826 4.5005
R14463 DVSS.n16850 DVSS.n16826 4.5005
R14464 DVSS.n16837 DVSS.n16826 4.5005
R14465 DVSS.n16851 DVSS.n16826 4.5005
R14466 DVSS.n17615 DVSS.n16826 4.5005
R14467 DVSS.n16825 DVSS.n16159 4.5005
R14468 DVSS.n16825 DVSS.n16160 4.5005
R14469 DVSS.n16825 DVSS.n16158 4.5005
R14470 DVSS.n16825 DVSS.n16161 4.5005
R14471 DVSS.n16825 DVSS.n16156 4.5005
R14472 DVSS.n16825 DVSS.n16162 4.5005
R14473 DVSS.n16825 DVSS.n16155 4.5005
R14474 DVSS.n16825 DVSS.n16163 4.5005
R14475 DVSS.n16825 DVSS.n16154 4.5005
R14476 DVSS.n16825 DVSS.n16164 4.5005
R14477 DVSS.n16825 DVSS.n16824 4.5005
R14478 DVSS.n16170 DVSS.n16159 4.5005
R14479 DVSS.n16170 DVSS.n16160 4.5005
R14480 DVSS.n16170 DVSS.n16158 4.5005
R14481 DVSS.n16224 DVSS.n16170 4.5005
R14482 DVSS.n16185 DVSS.n16170 4.5005
R14483 DVSS.n16170 DVSS.n16161 4.5005
R14484 DVSS.n16170 DVSS.n16156 4.5005
R14485 DVSS.n16170 DVSS.n16162 4.5005
R14486 DVSS.n16170 DVSS.n16155 4.5005
R14487 DVSS.n16170 DVSS.n16163 4.5005
R14488 DVSS.n16170 DVSS.n16154 4.5005
R14489 DVSS.n16822 DVSS.n16170 4.5005
R14490 DVSS.n16170 DVSS.n16164 4.5005
R14491 DVSS.n16824 DVSS.n16170 4.5005
R14492 DVSS.n16172 DVSS.n16159 4.5005
R14493 DVSS.n16172 DVSS.n16160 4.5005
R14494 DVSS.n16172 DVSS.n16158 4.5005
R14495 DVSS.n16224 DVSS.n16172 4.5005
R14496 DVSS.n16185 DVSS.n16172 4.5005
R14497 DVSS.n16172 DVSS.n16161 4.5005
R14498 DVSS.n16172 DVSS.n16156 4.5005
R14499 DVSS.n16172 DVSS.n16162 4.5005
R14500 DVSS.n16172 DVSS.n16155 4.5005
R14501 DVSS.n16172 DVSS.n16163 4.5005
R14502 DVSS.n16172 DVSS.n16154 4.5005
R14503 DVSS.n16822 DVSS.n16172 4.5005
R14504 DVSS.n16172 DVSS.n16164 4.5005
R14505 DVSS.n16179 DVSS.n16172 4.5005
R14506 DVSS.n16824 DVSS.n16172 4.5005
R14507 DVSS.n16169 DVSS.n16159 4.5005
R14508 DVSS.n16169 DVSS.n16160 4.5005
R14509 DVSS.n16169 DVSS.n16158 4.5005
R14510 DVSS.n16224 DVSS.n16169 4.5005
R14511 DVSS.n16185 DVSS.n16169 4.5005
R14512 DVSS.n16169 DVSS.n16161 4.5005
R14513 DVSS.n16169 DVSS.n16156 4.5005
R14514 DVSS.n16169 DVSS.n16162 4.5005
R14515 DVSS.n16169 DVSS.n16155 4.5005
R14516 DVSS.n16169 DVSS.n16163 4.5005
R14517 DVSS.n16169 DVSS.n16154 4.5005
R14518 DVSS.n16822 DVSS.n16169 4.5005
R14519 DVSS.n16169 DVSS.n16164 4.5005
R14520 DVSS.n16824 DVSS.n16169 4.5005
R14521 DVSS.n16173 DVSS.n16159 4.5005
R14522 DVSS.n16173 DVSS.n16160 4.5005
R14523 DVSS.n16173 DVSS.n16158 4.5005
R14524 DVSS.n16224 DVSS.n16173 4.5005
R14525 DVSS.n16185 DVSS.n16173 4.5005
R14526 DVSS.n16173 DVSS.n16161 4.5005
R14527 DVSS.n16173 DVSS.n16156 4.5005
R14528 DVSS.n16173 DVSS.n16162 4.5005
R14529 DVSS.n16173 DVSS.n16155 4.5005
R14530 DVSS.n16173 DVSS.n16163 4.5005
R14531 DVSS.n16173 DVSS.n16154 4.5005
R14532 DVSS.n16822 DVSS.n16173 4.5005
R14533 DVSS.n16173 DVSS.n16164 4.5005
R14534 DVSS.n16824 DVSS.n16173 4.5005
R14535 DVSS.n16168 DVSS.n16159 4.5005
R14536 DVSS.n16168 DVSS.n16160 4.5005
R14537 DVSS.n16168 DVSS.n16158 4.5005
R14538 DVSS.n16224 DVSS.n16168 4.5005
R14539 DVSS.n16185 DVSS.n16168 4.5005
R14540 DVSS.n16168 DVSS.n16161 4.5005
R14541 DVSS.n16168 DVSS.n16156 4.5005
R14542 DVSS.n16168 DVSS.n16162 4.5005
R14543 DVSS.n16168 DVSS.n16155 4.5005
R14544 DVSS.n16168 DVSS.n16163 4.5005
R14545 DVSS.n16168 DVSS.n16154 4.5005
R14546 DVSS.n16822 DVSS.n16168 4.5005
R14547 DVSS.n16168 DVSS.n16164 4.5005
R14548 DVSS.n16824 DVSS.n16168 4.5005
R14549 DVSS.n16174 DVSS.n16159 4.5005
R14550 DVSS.n16174 DVSS.n16160 4.5005
R14551 DVSS.n16174 DVSS.n16158 4.5005
R14552 DVSS.n16224 DVSS.n16174 4.5005
R14553 DVSS.n16185 DVSS.n16174 4.5005
R14554 DVSS.n16174 DVSS.n16161 4.5005
R14555 DVSS.n16174 DVSS.n16156 4.5005
R14556 DVSS.n16174 DVSS.n16162 4.5005
R14557 DVSS.n16174 DVSS.n16155 4.5005
R14558 DVSS.n16174 DVSS.n16163 4.5005
R14559 DVSS.n16174 DVSS.n16154 4.5005
R14560 DVSS.n16822 DVSS.n16174 4.5005
R14561 DVSS.n16174 DVSS.n16164 4.5005
R14562 DVSS.n16824 DVSS.n16174 4.5005
R14563 DVSS.n16167 DVSS.n16159 4.5005
R14564 DVSS.n16167 DVSS.n16160 4.5005
R14565 DVSS.n16167 DVSS.n16158 4.5005
R14566 DVSS.n16224 DVSS.n16167 4.5005
R14567 DVSS.n16185 DVSS.n16167 4.5005
R14568 DVSS.n16167 DVSS.n16161 4.5005
R14569 DVSS.n16167 DVSS.n16156 4.5005
R14570 DVSS.n16167 DVSS.n16162 4.5005
R14571 DVSS.n16167 DVSS.n16155 4.5005
R14572 DVSS.n16167 DVSS.n16163 4.5005
R14573 DVSS.n16167 DVSS.n16154 4.5005
R14574 DVSS.n16822 DVSS.n16167 4.5005
R14575 DVSS.n16167 DVSS.n16164 4.5005
R14576 DVSS.n16179 DVSS.n16167 4.5005
R14577 DVSS.n16824 DVSS.n16167 4.5005
R14578 DVSS.n15762 DVSS.n15743 4.5005
R14579 DVSS.n15763 DVSS.n15743 4.5005
R14580 DVSS.n15761 DVSS.n15743 4.5005
R14581 DVSS.n15766 DVSS.n15743 4.5005
R14582 DVSS.n15759 DVSS.n15743 4.5005
R14583 DVSS.n15767 DVSS.n15743 4.5005
R14584 DVSS.n15758 DVSS.n15743 4.5005
R14585 DVSS.n15768 DVSS.n15743 4.5005
R14586 DVSS.n15757 DVSS.n15743 4.5005
R14587 DVSS.n17947 DVSS.n15743 4.5005
R14588 DVSS.n17949 DVSS.n15743 4.5005
R14589 DVSS.n15762 DVSS.n15745 4.5005
R14590 DVSS.n15763 DVSS.n15745 4.5005
R14591 DVSS.n15761 DVSS.n15745 4.5005
R14592 DVSS.n15765 DVSS.n15745 4.5005
R14593 DVSS.n15760 DVSS.n15745 4.5005
R14594 DVSS.n15766 DVSS.n15745 4.5005
R14595 DVSS.n15759 DVSS.n15745 4.5005
R14596 DVSS.n15767 DVSS.n15745 4.5005
R14597 DVSS.n15758 DVSS.n15745 4.5005
R14598 DVSS.n15768 DVSS.n15745 4.5005
R14599 DVSS.n15757 DVSS.n15745 4.5005
R14600 DVSS.n15770 DVSS.n15745 4.5005
R14601 DVSS.n17947 DVSS.n15745 4.5005
R14602 DVSS.n17949 DVSS.n15745 4.5005
R14603 DVSS.n15762 DVSS.n15742 4.5005
R14604 DVSS.n15763 DVSS.n15742 4.5005
R14605 DVSS.n15761 DVSS.n15742 4.5005
R14606 DVSS.n15765 DVSS.n15742 4.5005
R14607 DVSS.n15760 DVSS.n15742 4.5005
R14608 DVSS.n15766 DVSS.n15742 4.5005
R14609 DVSS.n15759 DVSS.n15742 4.5005
R14610 DVSS.n15767 DVSS.n15742 4.5005
R14611 DVSS.n15758 DVSS.n15742 4.5005
R14612 DVSS.n15768 DVSS.n15742 4.5005
R14613 DVSS.n15757 DVSS.n15742 4.5005
R14614 DVSS.n15770 DVSS.n15742 4.5005
R14615 DVSS.n17947 DVSS.n15742 4.5005
R14616 DVSS.n17949 DVSS.n15742 4.5005
R14617 DVSS.n15762 DVSS.n15747 4.5005
R14618 DVSS.n15763 DVSS.n15747 4.5005
R14619 DVSS.n15761 DVSS.n15747 4.5005
R14620 DVSS.n15765 DVSS.n15747 4.5005
R14621 DVSS.n15760 DVSS.n15747 4.5005
R14622 DVSS.n15766 DVSS.n15747 4.5005
R14623 DVSS.n15759 DVSS.n15747 4.5005
R14624 DVSS.n15767 DVSS.n15747 4.5005
R14625 DVSS.n15758 DVSS.n15747 4.5005
R14626 DVSS.n15768 DVSS.n15747 4.5005
R14627 DVSS.n15757 DVSS.n15747 4.5005
R14628 DVSS.n15770 DVSS.n15747 4.5005
R14629 DVSS.n17947 DVSS.n15747 4.5005
R14630 DVSS.n17949 DVSS.n15747 4.5005
R14631 DVSS.n15762 DVSS.n15741 4.5005
R14632 DVSS.n15763 DVSS.n15741 4.5005
R14633 DVSS.n15761 DVSS.n15741 4.5005
R14634 DVSS.n15765 DVSS.n15741 4.5005
R14635 DVSS.n15760 DVSS.n15741 4.5005
R14636 DVSS.n15766 DVSS.n15741 4.5005
R14637 DVSS.n15759 DVSS.n15741 4.5005
R14638 DVSS.n15767 DVSS.n15741 4.5005
R14639 DVSS.n15758 DVSS.n15741 4.5005
R14640 DVSS.n15768 DVSS.n15741 4.5005
R14641 DVSS.n15757 DVSS.n15741 4.5005
R14642 DVSS.n15770 DVSS.n15741 4.5005
R14643 DVSS.n17947 DVSS.n15741 4.5005
R14644 DVSS.n17949 DVSS.n15741 4.5005
R14645 DVSS.n15762 DVSS.n15749 4.5005
R14646 DVSS.n15763 DVSS.n15749 4.5005
R14647 DVSS.n15761 DVSS.n15749 4.5005
R14648 DVSS.n15765 DVSS.n15749 4.5005
R14649 DVSS.n15760 DVSS.n15749 4.5005
R14650 DVSS.n15766 DVSS.n15749 4.5005
R14651 DVSS.n15759 DVSS.n15749 4.5005
R14652 DVSS.n15767 DVSS.n15749 4.5005
R14653 DVSS.n15758 DVSS.n15749 4.5005
R14654 DVSS.n15768 DVSS.n15749 4.5005
R14655 DVSS.n15757 DVSS.n15749 4.5005
R14656 DVSS.n15770 DVSS.n15749 4.5005
R14657 DVSS.n17947 DVSS.n15749 4.5005
R14658 DVSS.n17949 DVSS.n15749 4.5005
R14659 DVSS.n15762 DVSS.n15740 4.5005
R14660 DVSS.n15763 DVSS.n15740 4.5005
R14661 DVSS.n15761 DVSS.n15740 4.5005
R14662 DVSS.n15765 DVSS.n15740 4.5005
R14663 DVSS.n15760 DVSS.n15740 4.5005
R14664 DVSS.n15766 DVSS.n15740 4.5005
R14665 DVSS.n15759 DVSS.n15740 4.5005
R14666 DVSS.n15767 DVSS.n15740 4.5005
R14667 DVSS.n15758 DVSS.n15740 4.5005
R14668 DVSS.n15768 DVSS.n15740 4.5005
R14669 DVSS.n15757 DVSS.n15740 4.5005
R14670 DVSS.n15770 DVSS.n15740 4.5005
R14671 DVSS.n17947 DVSS.n15740 4.5005
R14672 DVSS.n17949 DVSS.n15740 4.5005
R14673 DVSS.n15762 DVSS.n15751 4.5005
R14674 DVSS.n15763 DVSS.n15751 4.5005
R14675 DVSS.n15761 DVSS.n15751 4.5005
R14676 DVSS.n15765 DVSS.n15751 4.5005
R14677 DVSS.n15760 DVSS.n15751 4.5005
R14678 DVSS.n15766 DVSS.n15751 4.5005
R14679 DVSS.n15759 DVSS.n15751 4.5005
R14680 DVSS.n15767 DVSS.n15751 4.5005
R14681 DVSS.n15758 DVSS.n15751 4.5005
R14682 DVSS.n15768 DVSS.n15751 4.5005
R14683 DVSS.n15757 DVSS.n15751 4.5005
R14684 DVSS.n15770 DVSS.n15751 4.5005
R14685 DVSS.n17947 DVSS.n15751 4.5005
R14686 DVSS.n17949 DVSS.n15751 4.5005
R14687 DVSS.n15762 DVSS.n15739 4.5005
R14688 DVSS.n15763 DVSS.n15739 4.5005
R14689 DVSS.n15761 DVSS.n15739 4.5005
R14690 DVSS.n15765 DVSS.n15739 4.5005
R14691 DVSS.n15760 DVSS.n15739 4.5005
R14692 DVSS.n15766 DVSS.n15739 4.5005
R14693 DVSS.n15759 DVSS.n15739 4.5005
R14694 DVSS.n15767 DVSS.n15739 4.5005
R14695 DVSS.n15758 DVSS.n15739 4.5005
R14696 DVSS.n15768 DVSS.n15739 4.5005
R14697 DVSS.n15757 DVSS.n15739 4.5005
R14698 DVSS.n15770 DVSS.n15739 4.5005
R14699 DVSS.n17947 DVSS.n15739 4.5005
R14700 DVSS.n15739 DVSS.n15738 4.5005
R14701 DVSS.n17949 DVSS.n15739 4.5005
R14702 DVSS.n17948 DVSS.n15762 4.5005
R14703 DVSS.n17948 DVSS.n15763 4.5005
R14704 DVSS.n17948 DVSS.n15761 4.5005
R14705 DVSS.n17948 DVSS.n15765 4.5005
R14706 DVSS.n17948 DVSS.n15760 4.5005
R14707 DVSS.n17948 DVSS.n15766 4.5005
R14708 DVSS.n17948 DVSS.n15759 4.5005
R14709 DVSS.n17948 DVSS.n15767 4.5005
R14710 DVSS.n17948 DVSS.n15758 4.5005
R14711 DVSS.n17948 DVSS.n15768 4.5005
R14712 DVSS.n17948 DVSS.n15757 4.5005
R14713 DVSS.n17948 DVSS.n15770 4.5005
R14714 DVSS.n17948 DVSS.n15756 4.5005
R14715 DVSS.n17948 DVSS.n17947 4.5005
R14716 DVSS.n17948 DVSS.n15738 4.5005
R14717 DVSS.n17949 DVSS.n17948 4.5005
R14718 DVSS.n16175 DVSS.n16159 4.5005
R14719 DVSS.n16175 DVSS.n16160 4.5005
R14720 DVSS.n16175 DVSS.n16158 4.5005
R14721 DVSS.n16224 DVSS.n16175 4.5005
R14722 DVSS.n16185 DVSS.n16175 4.5005
R14723 DVSS.n16175 DVSS.n16161 4.5005
R14724 DVSS.n16175 DVSS.n16156 4.5005
R14725 DVSS.n16175 DVSS.n16162 4.5005
R14726 DVSS.n16175 DVSS.n16155 4.5005
R14727 DVSS.n16175 DVSS.n16163 4.5005
R14728 DVSS.n16175 DVSS.n16154 4.5005
R14729 DVSS.n16822 DVSS.n16175 4.5005
R14730 DVSS.n16175 DVSS.n16164 4.5005
R14731 DVSS.n16179 DVSS.n16175 4.5005
R14732 DVSS.n16824 DVSS.n16175 4.5005
R14733 DVSS.n16166 DVSS.n16159 4.5005
R14734 DVSS.n16166 DVSS.n16160 4.5005
R14735 DVSS.n16166 DVSS.n16158 4.5005
R14736 DVSS.n16224 DVSS.n16166 4.5005
R14737 DVSS.n16185 DVSS.n16166 4.5005
R14738 DVSS.n16166 DVSS.n16161 4.5005
R14739 DVSS.n16166 DVSS.n16156 4.5005
R14740 DVSS.n16166 DVSS.n16162 4.5005
R14741 DVSS.n16166 DVSS.n16155 4.5005
R14742 DVSS.n16166 DVSS.n16163 4.5005
R14743 DVSS.n16166 DVSS.n16154 4.5005
R14744 DVSS.n16822 DVSS.n16166 4.5005
R14745 DVSS.n16184 DVSS.n16166 4.5005
R14746 DVSS.n16166 DVSS.n16164 4.5005
R14747 DVSS.n16179 DVSS.n16166 4.5005
R14748 DVSS.n16824 DVSS.n16166 4.5005
R14749 DVSS.n16823 DVSS.n16159 4.5005
R14750 DVSS.n16823 DVSS.n16160 4.5005
R14751 DVSS.n16823 DVSS.n16158 4.5005
R14752 DVSS.n16823 DVSS.n16224 4.5005
R14753 DVSS.n16823 DVSS.n16185 4.5005
R14754 DVSS.n16823 DVSS.n16161 4.5005
R14755 DVSS.n16823 DVSS.n16156 4.5005
R14756 DVSS.n16823 DVSS.n16162 4.5005
R14757 DVSS.n16823 DVSS.n16155 4.5005
R14758 DVSS.n16823 DVSS.n16163 4.5005
R14759 DVSS.n16823 DVSS.n16154 4.5005
R14760 DVSS.n16823 DVSS.n16822 4.5005
R14761 DVSS.n16823 DVSS.n16184 4.5005
R14762 DVSS.n16823 DVSS.n16164 4.5005
R14763 DVSS.n16823 DVSS.n16179 4.5005
R14764 DVSS.n16824 DVSS.n16823 4.5005
R14765 DVSS.n16142 DVSS.n16141 4.5005
R14766 DVSS.n17617 DVSS.n16142 4.5005
R14767 DVSS.n16842 DVSS.n16142 4.5005
R14768 DVSS.n16845 DVSS.n16142 4.5005
R14769 DVSS.n16841 DVSS.n16142 4.5005
R14770 DVSS.n16846 DVSS.n16142 4.5005
R14771 DVSS.n16840 DVSS.n16142 4.5005
R14772 DVSS.n16847 DVSS.n16142 4.5005
R14773 DVSS.n16839 DVSS.n16142 4.5005
R14774 DVSS.n16848 DVSS.n16142 4.5005
R14775 DVSS.n16838 DVSS.n16142 4.5005
R14776 DVSS.n16850 DVSS.n16142 4.5005
R14777 DVSS.n16851 DVSS.n16142 4.5005
R14778 DVSS.n16832 DVSS.n16142 4.5005
R14779 DVSS.n17615 DVSS.n16142 4.5005
R14780 DVSS.n17616 DVSS.n16141 4.5005
R14781 DVSS.n17617 DVSS.n17616 4.5005
R14782 DVSS.n17616 DVSS.n16842 4.5005
R14783 DVSS.n17616 DVSS.n16845 4.5005
R14784 DVSS.n17616 DVSS.n16841 4.5005
R14785 DVSS.n17616 DVSS.n16846 4.5005
R14786 DVSS.n17616 DVSS.n16840 4.5005
R14787 DVSS.n17616 DVSS.n16847 4.5005
R14788 DVSS.n17616 DVSS.n16839 4.5005
R14789 DVSS.n17616 DVSS.n16848 4.5005
R14790 DVSS.n17616 DVSS.n16838 4.5005
R14791 DVSS.n17616 DVSS.n16850 4.5005
R14792 DVSS.n17616 DVSS.n16837 4.5005
R14793 DVSS.n17616 DVSS.n16851 4.5005
R14794 DVSS.n17616 DVSS.n16832 4.5005
R14795 DVSS.n17616 DVSS.n17615 4.5005
R14796 DVSS.n15372 DVSS.n15362 4.5005
R14797 DVSS.n18327 DVSS.n15372 4.5005
R14798 DVSS.n15386 DVSS.n15372 4.5005
R14799 DVSS.n15389 DVSS.n15372 4.5005
R14800 DVSS.n15385 DVSS.n15372 4.5005
R14801 DVSS.n15390 DVSS.n15372 4.5005
R14802 DVSS.n15384 DVSS.n15372 4.5005
R14803 DVSS.n15391 DVSS.n15372 4.5005
R14804 DVSS.n15383 DVSS.n15372 4.5005
R14805 DVSS.n15392 DVSS.n15372 4.5005
R14806 DVSS.n15382 DVSS.n15372 4.5005
R14807 DVSS.n15394 DVSS.n15372 4.5005
R14808 DVSS.n15381 DVSS.n15372 4.5005
R14809 DVSS.n15395 DVSS.n15372 4.5005
R14810 DVSS.n15377 DVSS.n15372 4.5005
R14811 DVSS.n18325 DVSS.n15372 4.5005
R14812 DVSS.n15363 DVSS.n15362 4.5005
R14813 DVSS.n18327 DVSS.n15363 4.5005
R14814 DVSS.n15386 DVSS.n15363 4.5005
R14815 DVSS.n15389 DVSS.n15363 4.5005
R14816 DVSS.n15385 DVSS.n15363 4.5005
R14817 DVSS.n15390 DVSS.n15363 4.5005
R14818 DVSS.n15384 DVSS.n15363 4.5005
R14819 DVSS.n15391 DVSS.n15363 4.5005
R14820 DVSS.n15383 DVSS.n15363 4.5005
R14821 DVSS.n15392 DVSS.n15363 4.5005
R14822 DVSS.n15382 DVSS.n15363 4.5005
R14823 DVSS.n15394 DVSS.n15363 4.5005
R14824 DVSS.n15395 DVSS.n15363 4.5005
R14825 DVSS.n15377 DVSS.n15363 4.5005
R14826 DVSS.n18325 DVSS.n15363 4.5005
R14827 DVSS.n18326 DVSS.n15362 4.5005
R14828 DVSS.n18327 DVSS.n18326 4.5005
R14829 DVSS.n18326 DVSS.n15386 4.5005
R14830 DVSS.n18326 DVSS.n15389 4.5005
R14831 DVSS.n18326 DVSS.n15385 4.5005
R14832 DVSS.n18326 DVSS.n15390 4.5005
R14833 DVSS.n18326 DVSS.n15384 4.5005
R14834 DVSS.n18326 DVSS.n15391 4.5005
R14835 DVSS.n18326 DVSS.n15383 4.5005
R14836 DVSS.n18326 DVSS.n15392 4.5005
R14837 DVSS.n18326 DVSS.n15382 4.5005
R14838 DVSS.n18326 DVSS.n15394 4.5005
R14839 DVSS.n18326 DVSS.n15381 4.5005
R14840 DVSS.n18326 DVSS.n15395 4.5005
R14841 DVSS.n18326 DVSS.n15377 4.5005
R14842 DVSS.n18326 DVSS.n18325 4.5005
R14843 DVSS.n22460 DVSS.n867 4.5005
R14844 DVSS.n22460 DVSS.n22459 4.5005
R14845 DVSS.n1333 DVSS.n680 4.5005
R14846 DVSS.n1352 DVSS.n669 4.5005
R14847 DVSS.n22458 DVSS.n22457 4.5005
R14848 DVSS.n22459 DVSS.n22458 4.5005
R14849 DVSS.n20688 DVSS.n14557 4.5005
R14850 DVSS.n20688 DVSS.n14556 4.5005
R14851 DVSS.n20688 DVSS.n14558 4.5005
R14852 DVSS.n20688 DVSS.n14555 4.5005
R14853 DVSS.n20688 DVSS.n14559 4.5005
R14854 DVSS.n20689 DVSS.n20688 4.5005
R14855 DVSS.n20688 DVSS.n14562 4.5005
R14856 DVSS.n20688 DVSS.n14554 4.5005
R14857 DVSS.n20688 DVSS.n14563 4.5005
R14858 DVSS.n20688 DVSS.n14553 4.5005
R14859 DVSS.n20688 DVSS.n14564 4.5005
R14860 DVSS.n20688 DVSS.n14552 4.5005
R14861 DVSS.n20688 DVSS.n14565 4.5005
R14862 DVSS.n20688 DVSS.n14551 4.5005
R14863 DVSS.n20688 DVSS.n14566 4.5005
R14864 DVSS.n20688 DVSS.n20687 4.5005
R14865 DVSS.n18985 DVSS.n13879 4.5005
R14866 DVSS.n18882 DVSS.n13879 4.5005
R14867 DVSS.n18881 DVSS.n13879 4.5005
R14868 DVSS.n18908 DVSS.n13879 4.5005
R14869 DVSS.n18880 DVSS.n13879 4.5005
R14870 DVSS.n18910 DVSS.n13879 4.5005
R14871 DVSS.n18879 DVSS.n13879 4.5005
R14872 DVSS.n18911 DVSS.n13879 4.5005
R14873 DVSS.n18878 DVSS.n13879 4.5005
R14874 DVSS.n18912 DVSS.n13879 4.5005
R14875 DVSS.n18877 DVSS.n13879 4.5005
R14876 DVSS.n18913 DVSS.n13879 4.5005
R14877 DVSS.n18876 DVSS.n13879 4.5005
R14878 DVSS.n18983 DVSS.n13879 4.5005
R14879 DVSS.n18915 DVSS.n13879 4.5005
R14880 DVSS.n14576 DVSS.n13879 4.5005
R14881 DVSS.n18985 DVSS.n18873 4.5005
R14882 DVSS.n18882 DVSS.n18873 4.5005
R14883 DVSS.n18881 DVSS.n18873 4.5005
R14884 DVSS.n18908 DVSS.n18873 4.5005
R14885 DVSS.n18880 DVSS.n18873 4.5005
R14886 DVSS.n18910 DVSS.n18873 4.5005
R14887 DVSS.n18879 DVSS.n18873 4.5005
R14888 DVSS.n18911 DVSS.n18873 4.5005
R14889 DVSS.n18878 DVSS.n18873 4.5005
R14890 DVSS.n18912 DVSS.n18873 4.5005
R14891 DVSS.n18877 DVSS.n18873 4.5005
R14892 DVSS.n18913 DVSS.n18873 4.5005
R14893 DVSS.n18876 DVSS.n18873 4.5005
R14894 DVSS.n18983 DVSS.n18873 4.5005
R14895 DVSS.n18915 DVSS.n18873 4.5005
R14896 DVSS.n18873 DVSS.n14576 4.5005
R14897 DVSS.n18985 DVSS.n18871 4.5005
R14898 DVSS.n18882 DVSS.n18871 4.5005
R14899 DVSS.n18881 DVSS.n18871 4.5005
R14900 DVSS.n18908 DVSS.n18871 4.5005
R14901 DVSS.n18880 DVSS.n18871 4.5005
R14902 DVSS.n18910 DVSS.n18871 4.5005
R14903 DVSS.n18879 DVSS.n18871 4.5005
R14904 DVSS.n18911 DVSS.n18871 4.5005
R14905 DVSS.n18878 DVSS.n18871 4.5005
R14906 DVSS.n18912 DVSS.n18871 4.5005
R14907 DVSS.n18877 DVSS.n18871 4.5005
R14908 DVSS.n18913 DVSS.n18871 4.5005
R14909 DVSS.n18876 DVSS.n18871 4.5005
R14910 DVSS.n18983 DVSS.n18871 4.5005
R14911 DVSS.n18915 DVSS.n18871 4.5005
R14912 DVSS.n18871 DVSS.n14576 4.5005
R14913 DVSS.n20699 DVSS.n14526 4.5005
R14914 DVSS.n20699 DVSS.n14525 4.5005
R14915 DVSS.n20699 DVSS.n14527 4.5005
R14916 DVSS.n20699 DVSS.n14524 4.5005
R14917 DVSS.n20699 DVSS.n14528 4.5005
R14918 DVSS.n20699 DVSS.n14523 4.5005
R14919 DVSS.n20699 DVSS.n14529 4.5005
R14920 DVSS.n20699 DVSS.n14521 4.5005
R14921 DVSS.n20699 DVSS.n14530 4.5005
R14922 DVSS.n20699 DVSS.n14520 4.5005
R14923 DVSS.n20699 DVSS.n14531 4.5005
R14924 DVSS.n20699 DVSS.n14519 4.5005
R14925 DVSS.n20699 DVSS.n14532 4.5005
R14926 DVSS.n20699 DVSS.n14518 4.5005
R14927 DVSS.n20699 DVSS.n14533 4.5005
R14928 DVSS.n20699 DVSS.n20698 4.5005
R14929 DVSS.n20697 DVSS.n14526 4.5005
R14930 DVSS.n20697 DVSS.n14525 4.5005
R14931 DVSS.n20697 DVSS.n14527 4.5005
R14932 DVSS.n20697 DVSS.n14524 4.5005
R14933 DVSS.n20697 DVSS.n14528 4.5005
R14934 DVSS.n20697 DVSS.n14537 4.5005
R14935 DVSS.n20697 DVSS.n14529 4.5005
R14936 DVSS.n20697 DVSS.n14521 4.5005
R14937 DVSS.n20697 DVSS.n14530 4.5005
R14938 DVSS.n20697 DVSS.n14520 4.5005
R14939 DVSS.n20697 DVSS.n14531 4.5005
R14940 DVSS.n20697 DVSS.n14519 4.5005
R14941 DVSS.n20697 DVSS.n14532 4.5005
R14942 DVSS.n20697 DVSS.n14518 4.5005
R14943 DVSS.n20697 DVSS.n14533 4.5005
R14944 DVSS.n20698 DVSS.n20697 4.5005
R14945 DVSS.n18985 DVSS.n18984 4.5005
R14946 DVSS.n18984 DVSS.n18882 4.5005
R14947 DVSS.n18984 DVSS.n18881 4.5005
R14948 DVSS.n18984 DVSS.n18908 4.5005
R14949 DVSS.n18984 DVSS.n18880 4.5005
R14950 DVSS.n18984 DVSS.n18910 4.5005
R14951 DVSS.n18984 DVSS.n18879 4.5005
R14952 DVSS.n18984 DVSS.n18911 4.5005
R14953 DVSS.n18984 DVSS.n18878 4.5005
R14954 DVSS.n18984 DVSS.n18912 4.5005
R14955 DVSS.n18984 DVSS.n18877 4.5005
R14956 DVSS.n18984 DVSS.n18913 4.5005
R14957 DVSS.n18984 DVSS.n18876 4.5005
R14958 DVSS.n18984 DVSS.n18983 4.5005
R14959 DVSS.n18984 DVSS.n14576 4.5005
R14960 DVSS.n18985 DVSS.n18870 4.5005
R14961 DVSS.n18882 DVSS.n18870 4.5005
R14962 DVSS.n18881 DVSS.n18870 4.5005
R14963 DVSS.n18908 DVSS.n18870 4.5005
R14964 DVSS.n18880 DVSS.n18870 4.5005
R14965 DVSS.n18910 DVSS.n18870 4.5005
R14966 DVSS.n18879 DVSS.n18870 4.5005
R14967 DVSS.n18911 DVSS.n18870 4.5005
R14968 DVSS.n18878 DVSS.n18870 4.5005
R14969 DVSS.n18912 DVSS.n18870 4.5005
R14970 DVSS.n18877 DVSS.n18870 4.5005
R14971 DVSS.n18913 DVSS.n18870 4.5005
R14972 DVSS.n18983 DVSS.n18870 4.5005
R14973 DVSS.n18870 DVSS.n14576 4.5005
R14974 DVSS.n18985 DVSS.n13849 4.5005
R14975 DVSS.n18882 DVSS.n13849 4.5005
R14976 DVSS.n18881 DVSS.n13849 4.5005
R14977 DVSS.n18908 DVSS.n13849 4.5005
R14978 DVSS.n18880 DVSS.n13849 4.5005
R14979 DVSS.n18910 DVSS.n13849 4.5005
R14980 DVSS.n18879 DVSS.n13849 4.5005
R14981 DVSS.n18911 DVSS.n13849 4.5005
R14982 DVSS.n18878 DVSS.n13849 4.5005
R14983 DVSS.n18912 DVSS.n13849 4.5005
R14984 DVSS.n18877 DVSS.n13849 4.5005
R14985 DVSS.n18913 DVSS.n13849 4.5005
R14986 DVSS.n18983 DVSS.n13849 4.5005
R14987 DVSS.n18915 DVSS.n13849 4.5005
R14988 DVSS.n14576 DVSS.n13849 4.5005
R14989 DVSS.n14556 DVSS.n14548 4.5005
R14990 DVSS.n14558 DVSS.n14548 4.5005
R14991 DVSS.n14555 DVSS.n14548 4.5005
R14992 DVSS.n14559 DVSS.n14548 4.5005
R14993 DVSS.n14560 DVSS.n14548 4.5005
R14994 DVSS.n14562 DVSS.n14548 4.5005
R14995 DVSS.n14554 DVSS.n14548 4.5005
R14996 DVSS.n14563 DVSS.n14548 4.5005
R14997 DVSS.n14553 DVSS.n14548 4.5005
R14998 DVSS.n14564 DVSS.n14548 4.5005
R14999 DVSS.n14552 DVSS.n14548 4.5005
R15000 DVSS.n14565 DVSS.n14548 4.5005
R15001 DVSS.n14551 DVSS.n14548 4.5005
R15002 DVSS.n14566 DVSS.n14548 4.5005
R15003 DVSS.n20687 DVSS.n14548 4.5005
R15004 DVSS.n14557 DVSS.n14548 4.5005
R15005 DVSS.n17056 DVSS.n16005 4.5005
R15006 DVSS.n17115 DVSS.n16005 4.5005
R15007 DVSS.n17101 DVSS.n16005 4.5005
R15008 DVSS.n16977 DVSS.n15273 4.5005
R15009 DVSS.n17312 DVSS.n17310 4.5005
R15010 DVSS.n17379 DVSS.n17312 4.5005
R15011 DVSS.n17319 DVSS.n17312 4.5005
R15012 DVSS.n17371 DVSS.n17312 4.5005
R15013 DVSS.n17372 DVSS.n17310 4.5005
R15014 DVSS.n17372 DVSS.n17371 4.5005
R15015 DVSS.n17401 DVSS.n17383 4.5005
R15016 DVSS.n17403 DVSS.n17383 4.5005
R15017 DVSS.n17403 DVSS.n17309 4.5005
R15018 DVSS.n17403 DVSS.n17384 4.5005
R15019 DVSS.n17403 DVSS.n17402 4.5005
R15020 DVSS.n17404 DVSS.n17403 4.5005
R15021 DVSS.n17383 DVSS.n17302 4.5005
R15022 DVSS.n17309 DVSS.n17302 4.5005
R15023 DVSS.n17391 DVSS.n17302 4.5005
R15024 DVSS.n17393 DVSS.n17302 4.5005
R15025 DVSS.n17402 DVSS.n17302 4.5005
R15026 DVSS.n17404 DVSS.n17302 4.5005
R15027 DVSS.n17301 DVSS.n17118 4.5005
R15028 DVSS.n17119 DVSS.n17118 4.5005
R15029 DVSS.n17480 DVSS.n17119 4.5005
R15030 DVSS.n17299 DVSS.n17119 4.5005
R15031 DVSS.n17135 DVSS.n17119 4.5005
R15032 DVSS.n17478 DVSS.n17119 4.5005
R15033 DVSS.n17301 DVSS.n17135 4.5005
R15034 DVSS.n17402 DVSS.n17401 4.5005
R15035 DVSS.n17401 DVSS.n17396 4.5005
R15036 DVSS.n17401 DVSS.n17390 4.5005
R15037 DVSS.n17401 DVSS.n17398 4.5005
R15038 DVSS.n17401 DVSS.n17389 4.5005
R15039 DVSS.n17401 DVSS.n17400 4.5005
R15040 DVSS.n17401 DVSS.n17388 4.5005
R15041 DVSS.n17378 DVSS.n17319 4.5005
R15042 DVSS.n17378 DVSS.n17317 4.5005
R15043 DVSS.n17378 DVSS.n17321 4.5005
R15044 DVSS.n17378 DVSS.n17316 4.5005
R15045 DVSS.n17378 DVSS.n17323 4.5005
R15046 DVSS.n17378 DVSS.n17315 4.5005
R15047 DVSS.n17378 DVSS.n17325 4.5005
R15048 DVSS.n17378 DVSS.n17314 4.5005
R15049 DVSS.n17378 DVSS.n17375 4.5005
R15050 DVSS.n17378 DVSS.n17313 4.5005
R15051 DVSS.n17378 DVSS.n17377 4.5005
R15052 DVSS.n17379 DVSS.n17378 4.5005
R15053 DVSS.n17378 DVSS.n17310 4.5005
R15054 DVSS.n17056 DVSS.n16021 4.5005
R15055 DVSS.n16977 DVSS.n15267 4.5005
R15056 DVSS.n17050 DVSS.n15267 4.5005
R15057 DVSS.n17036 DVSS.n15267 4.5005
R15058 DVSS.n17479 DVSS.n17118 4.5005
R15059 DVSS.n17480 DVSS.n17479 4.5005
R15060 DVSS.n17479 DVSS.n17127 4.5005
R15061 DVSS.n17479 DVSS.n17125 4.5005
R15062 DVSS.n17479 DVSS.n17129 4.5005
R15063 DVSS.n17479 DVSS.n17124 4.5005
R15064 DVSS.n17479 DVSS.n17131 4.5005
R15065 DVSS.n17479 DVSS.n17123 4.5005
R15066 DVSS.n17479 DVSS.n17133 4.5005
R15067 DVSS.n17479 DVSS.n17122 4.5005
R15068 DVSS.n17479 DVSS.n17135 4.5005
R15069 DVSS.n17479 DVSS.n17478 4.5005
R15070 DVSS.n16471 DVSS.n16360 4.5005
R15071 DVSS.n16365 DVSS.n16360 4.5005
R15072 DVSS.n16470 DVSS.n16365 4.5005
R15073 DVSS.n16470 DVSS.n16367 4.5005
R15074 DVSS.n16470 DVSS.n16364 4.5005
R15075 DVSS.n16470 DVSS.n16369 4.5005
R15076 DVSS.n16470 DVSS.n16363 4.5005
R15077 DVSS.n16470 DVSS.n16371 4.5005
R15078 DVSS.n16470 DVSS.n16362 4.5005
R15079 DVSS.n16470 DVSS.n16469 4.5005
R15080 DVSS.n16470 DVSS.n16361 4.5005
R15081 DVSS.n16471 DVSS.n16470 4.5005
R15082 DVSS.n13601 DVSS.n13576 4.5005
R15083 DVSS.n13587 DVSS.n13576 4.5005
R15084 DVSS.n13602 DVSS.n13576 4.5005
R15085 DVSS.n13586 DVSS.n13576 4.5005
R15086 DVSS.n13603 DVSS.n13576 4.5005
R15087 DVSS.n13585 DVSS.n13576 4.5005
R15088 DVSS.n21252 DVSS.n13576 4.5005
R15089 DVSS.n13584 DVSS.n13576 4.5005
R15090 DVSS.n21255 DVSS.n13576 4.5005
R15091 DVSS.n13576 DVSS.n13570 4.5005
R15092 DVSS.n21257 DVSS.n13576 4.5005
R15093 DVSS.n13587 DVSS.n13575 4.5005
R15094 DVSS.n13602 DVSS.n13575 4.5005
R15095 DVSS.n13586 DVSS.n13575 4.5005
R15096 DVSS.n13603 DVSS.n13575 4.5005
R15097 DVSS.n13585 DVSS.n13575 4.5005
R15098 DVSS.n21252 DVSS.n13575 4.5005
R15099 DVSS.n13584 DVSS.n13575 4.5005
R15100 DVSS.n21255 DVSS.n13575 4.5005
R15101 DVSS.n13575 DVSS.n13570 4.5005
R15102 DVSS.n21257 DVSS.n13575 4.5005
R15103 DVSS.n13591 DVSS.n13577 4.5005
R15104 DVSS.n13587 DVSS.n13577 4.5005
R15105 DVSS.n13602 DVSS.n13577 4.5005
R15106 DVSS.n13586 DVSS.n13577 4.5005
R15107 DVSS.n13603 DVSS.n13577 4.5005
R15108 DVSS.n13585 DVSS.n13577 4.5005
R15109 DVSS.n21252 DVSS.n13577 4.5005
R15110 DVSS.n13584 DVSS.n13577 4.5005
R15111 DVSS.n21255 DVSS.n13577 4.5005
R15112 DVSS.n13577 DVSS.n13570 4.5005
R15113 DVSS.n21257 DVSS.n13577 4.5005
R15114 DVSS.n13591 DVSS.n13574 4.5005
R15115 DVSS.n13587 DVSS.n13574 4.5005
R15116 DVSS.n13602 DVSS.n13574 4.5005
R15117 DVSS.n13586 DVSS.n13574 4.5005
R15118 DVSS.n13603 DVSS.n13574 4.5005
R15119 DVSS.n13585 DVSS.n13574 4.5005
R15120 DVSS.n21252 DVSS.n13574 4.5005
R15121 DVSS.n13584 DVSS.n13574 4.5005
R15122 DVSS.n21255 DVSS.n13574 4.5005
R15123 DVSS.n13574 DVSS.n13570 4.5005
R15124 DVSS.n21257 DVSS.n13574 4.5005
R15125 DVSS.n13587 DVSS.n13578 4.5005
R15126 DVSS.n13602 DVSS.n13578 4.5005
R15127 DVSS.n13586 DVSS.n13578 4.5005
R15128 DVSS.n13603 DVSS.n13578 4.5005
R15129 DVSS.n13585 DVSS.n13578 4.5005
R15130 DVSS.n21252 DVSS.n13578 4.5005
R15131 DVSS.n13584 DVSS.n13578 4.5005
R15132 DVSS.n21255 DVSS.n13578 4.5005
R15133 DVSS.n13578 DVSS.n13570 4.5005
R15134 DVSS.n21257 DVSS.n13578 4.5005
R15135 DVSS.n13587 DVSS.n13573 4.5005
R15136 DVSS.n13602 DVSS.n13573 4.5005
R15137 DVSS.n13586 DVSS.n13573 4.5005
R15138 DVSS.n13603 DVSS.n13573 4.5005
R15139 DVSS.n13585 DVSS.n13573 4.5005
R15140 DVSS.n21252 DVSS.n13573 4.5005
R15141 DVSS.n13584 DVSS.n13573 4.5005
R15142 DVSS.n21255 DVSS.n13573 4.5005
R15143 DVSS.n13573 DVSS.n13570 4.5005
R15144 DVSS.n21257 DVSS.n13573 4.5005
R15145 DVSS.n13587 DVSS.n13579 4.5005
R15146 DVSS.n13602 DVSS.n13579 4.5005
R15147 DVSS.n13586 DVSS.n13579 4.5005
R15148 DVSS.n13603 DVSS.n13579 4.5005
R15149 DVSS.n13585 DVSS.n13579 4.5005
R15150 DVSS.n21252 DVSS.n13579 4.5005
R15151 DVSS.n13584 DVSS.n13579 4.5005
R15152 DVSS.n21255 DVSS.n13579 4.5005
R15153 DVSS.n13579 DVSS.n13570 4.5005
R15154 DVSS.n21257 DVSS.n13579 4.5005
R15155 DVSS.n13587 DVSS.n13572 4.5005
R15156 DVSS.n13602 DVSS.n13572 4.5005
R15157 DVSS.n13586 DVSS.n13572 4.5005
R15158 DVSS.n13603 DVSS.n13572 4.5005
R15159 DVSS.n13585 DVSS.n13572 4.5005
R15160 DVSS.n21252 DVSS.n13572 4.5005
R15161 DVSS.n13584 DVSS.n13572 4.5005
R15162 DVSS.n21257 DVSS.n13572 4.5005
R15163 DVSS.n13591 DVSS.n13580 4.5005
R15164 DVSS.n13587 DVSS.n13580 4.5005
R15165 DVSS.n13602 DVSS.n13580 4.5005
R15166 DVSS.n13586 DVSS.n13580 4.5005
R15167 DVSS.n13603 DVSS.n13580 4.5005
R15168 DVSS.n13585 DVSS.n13580 4.5005
R15169 DVSS.n21252 DVSS.n13580 4.5005
R15170 DVSS.n21255 DVSS.n13580 4.5005
R15171 DVSS.n13580 DVSS.n13570 4.5005
R15172 DVSS.n21257 DVSS.n13580 4.5005
R15173 DVSS.n13593 DVSS.n13571 4.5005
R15174 DVSS.n13594 DVSS.n13571 4.5005
R15175 DVSS.n13592 DVSS.n13571 4.5005
R15176 DVSS.n13595 DVSS.n13571 4.5005
R15177 DVSS.n13591 DVSS.n13571 4.5005
R15178 DVSS.n13602 DVSS.n13571 4.5005
R15179 DVSS.n13586 DVSS.n13571 4.5005
R15180 DVSS.n13603 DVSS.n13571 4.5005
R15181 DVSS.n13585 DVSS.n13571 4.5005
R15182 DVSS.n21252 DVSS.n13571 4.5005
R15183 DVSS.n21255 DVSS.n13571 4.5005
R15184 DVSS.n21257 DVSS.n13571 4.5005
R15185 DVSS.n21256 DVSS.n13593 4.5005
R15186 DVSS.n21256 DVSS.n13594 4.5005
R15187 DVSS.n21256 DVSS.n13592 4.5005
R15188 DVSS.n21256 DVSS.n13595 4.5005
R15189 DVSS.n21256 DVSS.n13591 4.5005
R15190 DVSS.n21256 DVSS.n13601 4.5005
R15191 DVSS.n21256 DVSS.n13587 4.5005
R15192 DVSS.n21256 DVSS.n13602 4.5005
R15193 DVSS.n21256 DVSS.n13586 4.5005
R15194 DVSS.n21256 DVSS.n13603 4.5005
R15195 DVSS.n21256 DVSS.n13585 4.5005
R15196 DVSS.n21256 DVSS.n21252 4.5005
R15197 DVSS.n21256 DVSS.n13584 4.5005
R15198 DVSS.n21256 DVSS.n21255 4.5005
R15199 DVSS.n21257 DVSS.n21256 4.5005
R15200 DVSS.n13836 DVSS.n13824 4.5005
R15201 DVSS.n21116 DVSS.n13836 4.5005
R15202 DVSS.n13878 DVSS.n13836 4.5005
R15203 DVSS.n13880 DVSS.n13836 4.5005
R15204 DVSS.n13877 DVSS.n13836 4.5005
R15205 DVSS.n13883 DVSS.n13836 4.5005
R15206 DVSS.n13875 DVSS.n13836 4.5005
R15207 DVSS.n13884 DVSS.n13836 4.5005
R15208 DVSS.n13874 DVSS.n13836 4.5005
R15209 DVSS.n13885 DVSS.n13836 4.5005
R15210 DVSS.n13873 DVSS.n13836 4.5005
R15211 DVSS.n13887 DVSS.n13836 4.5005
R15212 DVSS.n21114 DVSS.n13836 4.5005
R15213 DVSS.n13838 DVSS.n13824 4.5005
R15214 DVSS.n21116 DVSS.n13838 4.5005
R15215 DVSS.n13878 DVSS.n13838 4.5005
R15216 DVSS.n13880 DVSS.n13838 4.5005
R15217 DVSS.n13877 DVSS.n13838 4.5005
R15218 DVSS.n13882 DVSS.n13838 4.5005
R15219 DVSS.n13876 DVSS.n13838 4.5005
R15220 DVSS.n13883 DVSS.n13838 4.5005
R15221 DVSS.n13875 DVSS.n13838 4.5005
R15222 DVSS.n13884 DVSS.n13838 4.5005
R15223 DVSS.n13874 DVSS.n13838 4.5005
R15224 DVSS.n13885 DVSS.n13838 4.5005
R15225 DVSS.n13887 DVSS.n13838 4.5005
R15226 DVSS.n21114 DVSS.n13838 4.5005
R15227 DVSS.n13835 DVSS.n13824 4.5005
R15228 DVSS.n21116 DVSS.n13835 4.5005
R15229 DVSS.n13878 DVSS.n13835 4.5005
R15230 DVSS.n13880 DVSS.n13835 4.5005
R15231 DVSS.n13877 DVSS.n13835 4.5005
R15232 DVSS.n13882 DVSS.n13835 4.5005
R15233 DVSS.n13876 DVSS.n13835 4.5005
R15234 DVSS.n13883 DVSS.n13835 4.5005
R15235 DVSS.n13875 DVSS.n13835 4.5005
R15236 DVSS.n13884 DVSS.n13835 4.5005
R15237 DVSS.n13874 DVSS.n13835 4.5005
R15238 DVSS.n13885 DVSS.n13835 4.5005
R15239 DVSS.n13887 DVSS.n13835 4.5005
R15240 DVSS.n21114 DVSS.n13835 4.5005
R15241 DVSS.n13839 DVSS.n13824 4.5005
R15242 DVSS.n21116 DVSS.n13839 4.5005
R15243 DVSS.n13878 DVSS.n13839 4.5005
R15244 DVSS.n13880 DVSS.n13839 4.5005
R15245 DVSS.n13877 DVSS.n13839 4.5005
R15246 DVSS.n13882 DVSS.n13839 4.5005
R15247 DVSS.n13876 DVSS.n13839 4.5005
R15248 DVSS.n13883 DVSS.n13839 4.5005
R15249 DVSS.n13875 DVSS.n13839 4.5005
R15250 DVSS.n13884 DVSS.n13839 4.5005
R15251 DVSS.n13874 DVSS.n13839 4.5005
R15252 DVSS.n13885 DVSS.n13839 4.5005
R15253 DVSS.n13887 DVSS.n13839 4.5005
R15254 DVSS.n21114 DVSS.n13839 4.5005
R15255 DVSS.n13834 DVSS.n13824 4.5005
R15256 DVSS.n21116 DVSS.n13834 4.5005
R15257 DVSS.n13878 DVSS.n13834 4.5005
R15258 DVSS.n13880 DVSS.n13834 4.5005
R15259 DVSS.n13877 DVSS.n13834 4.5005
R15260 DVSS.n13882 DVSS.n13834 4.5005
R15261 DVSS.n13876 DVSS.n13834 4.5005
R15262 DVSS.n13883 DVSS.n13834 4.5005
R15263 DVSS.n13875 DVSS.n13834 4.5005
R15264 DVSS.n13884 DVSS.n13834 4.5005
R15265 DVSS.n13874 DVSS.n13834 4.5005
R15266 DVSS.n13885 DVSS.n13834 4.5005
R15267 DVSS.n13887 DVSS.n13834 4.5005
R15268 DVSS.n21114 DVSS.n13834 4.5005
R15269 DVSS.n13840 DVSS.n13824 4.5005
R15270 DVSS.n21116 DVSS.n13840 4.5005
R15271 DVSS.n13878 DVSS.n13840 4.5005
R15272 DVSS.n13880 DVSS.n13840 4.5005
R15273 DVSS.n13877 DVSS.n13840 4.5005
R15274 DVSS.n13882 DVSS.n13840 4.5005
R15275 DVSS.n13876 DVSS.n13840 4.5005
R15276 DVSS.n13883 DVSS.n13840 4.5005
R15277 DVSS.n13875 DVSS.n13840 4.5005
R15278 DVSS.n13884 DVSS.n13840 4.5005
R15279 DVSS.n13874 DVSS.n13840 4.5005
R15280 DVSS.n13885 DVSS.n13840 4.5005
R15281 DVSS.n13887 DVSS.n13840 4.5005
R15282 DVSS.n21114 DVSS.n13840 4.5005
R15283 DVSS.n13833 DVSS.n13824 4.5005
R15284 DVSS.n21116 DVSS.n13833 4.5005
R15285 DVSS.n13878 DVSS.n13833 4.5005
R15286 DVSS.n13880 DVSS.n13833 4.5005
R15287 DVSS.n13877 DVSS.n13833 4.5005
R15288 DVSS.n13882 DVSS.n13833 4.5005
R15289 DVSS.n13876 DVSS.n13833 4.5005
R15290 DVSS.n13883 DVSS.n13833 4.5005
R15291 DVSS.n13875 DVSS.n13833 4.5005
R15292 DVSS.n13884 DVSS.n13833 4.5005
R15293 DVSS.n13874 DVSS.n13833 4.5005
R15294 DVSS.n13885 DVSS.n13833 4.5005
R15295 DVSS.n13887 DVSS.n13833 4.5005
R15296 DVSS.n21114 DVSS.n13833 4.5005
R15297 DVSS.n13841 DVSS.n13824 4.5005
R15298 DVSS.n21116 DVSS.n13841 4.5005
R15299 DVSS.n13878 DVSS.n13841 4.5005
R15300 DVSS.n13880 DVSS.n13841 4.5005
R15301 DVSS.n13877 DVSS.n13841 4.5005
R15302 DVSS.n13882 DVSS.n13841 4.5005
R15303 DVSS.n13876 DVSS.n13841 4.5005
R15304 DVSS.n13883 DVSS.n13841 4.5005
R15305 DVSS.n13875 DVSS.n13841 4.5005
R15306 DVSS.n13884 DVSS.n13841 4.5005
R15307 DVSS.n13874 DVSS.n13841 4.5005
R15308 DVSS.n13885 DVSS.n13841 4.5005
R15309 DVSS.n13887 DVSS.n13841 4.5005
R15310 DVSS.n21114 DVSS.n13841 4.5005
R15311 DVSS.n13832 DVSS.n13824 4.5005
R15312 DVSS.n21116 DVSS.n13832 4.5005
R15313 DVSS.n13878 DVSS.n13832 4.5005
R15314 DVSS.n13880 DVSS.n13832 4.5005
R15315 DVSS.n13877 DVSS.n13832 4.5005
R15316 DVSS.n13882 DVSS.n13832 4.5005
R15317 DVSS.n13876 DVSS.n13832 4.5005
R15318 DVSS.n13883 DVSS.n13832 4.5005
R15319 DVSS.n13875 DVSS.n13832 4.5005
R15320 DVSS.n13884 DVSS.n13832 4.5005
R15321 DVSS.n13874 DVSS.n13832 4.5005
R15322 DVSS.n13885 DVSS.n13832 4.5005
R15323 DVSS.n13887 DVSS.n13832 4.5005
R15324 DVSS.n21114 DVSS.n13832 4.5005
R15325 DVSS.n13842 DVSS.n13824 4.5005
R15326 DVSS.n21116 DVSS.n13842 4.5005
R15327 DVSS.n13878 DVSS.n13842 4.5005
R15328 DVSS.n13880 DVSS.n13842 4.5005
R15329 DVSS.n13877 DVSS.n13842 4.5005
R15330 DVSS.n13882 DVSS.n13842 4.5005
R15331 DVSS.n13876 DVSS.n13842 4.5005
R15332 DVSS.n13883 DVSS.n13842 4.5005
R15333 DVSS.n13875 DVSS.n13842 4.5005
R15334 DVSS.n13884 DVSS.n13842 4.5005
R15335 DVSS.n13874 DVSS.n13842 4.5005
R15336 DVSS.n13885 DVSS.n13842 4.5005
R15337 DVSS.n13887 DVSS.n13842 4.5005
R15338 DVSS.n21114 DVSS.n13842 4.5005
R15339 DVSS.n13831 DVSS.n13824 4.5005
R15340 DVSS.n21116 DVSS.n13831 4.5005
R15341 DVSS.n13878 DVSS.n13831 4.5005
R15342 DVSS.n13880 DVSS.n13831 4.5005
R15343 DVSS.n13877 DVSS.n13831 4.5005
R15344 DVSS.n13882 DVSS.n13831 4.5005
R15345 DVSS.n13876 DVSS.n13831 4.5005
R15346 DVSS.n13883 DVSS.n13831 4.5005
R15347 DVSS.n13875 DVSS.n13831 4.5005
R15348 DVSS.n13884 DVSS.n13831 4.5005
R15349 DVSS.n13874 DVSS.n13831 4.5005
R15350 DVSS.n13885 DVSS.n13831 4.5005
R15351 DVSS.n13887 DVSS.n13831 4.5005
R15352 DVSS.n21114 DVSS.n13831 4.5005
R15353 DVSS.n13843 DVSS.n13824 4.5005
R15354 DVSS.n21116 DVSS.n13843 4.5005
R15355 DVSS.n13878 DVSS.n13843 4.5005
R15356 DVSS.n13880 DVSS.n13843 4.5005
R15357 DVSS.n13877 DVSS.n13843 4.5005
R15358 DVSS.n13882 DVSS.n13843 4.5005
R15359 DVSS.n13876 DVSS.n13843 4.5005
R15360 DVSS.n13883 DVSS.n13843 4.5005
R15361 DVSS.n13875 DVSS.n13843 4.5005
R15362 DVSS.n13884 DVSS.n13843 4.5005
R15363 DVSS.n13874 DVSS.n13843 4.5005
R15364 DVSS.n13885 DVSS.n13843 4.5005
R15365 DVSS.n13887 DVSS.n13843 4.5005
R15366 DVSS.n21114 DVSS.n13843 4.5005
R15367 DVSS.n13830 DVSS.n13824 4.5005
R15368 DVSS.n21116 DVSS.n13830 4.5005
R15369 DVSS.n13878 DVSS.n13830 4.5005
R15370 DVSS.n13880 DVSS.n13830 4.5005
R15371 DVSS.n13877 DVSS.n13830 4.5005
R15372 DVSS.n13882 DVSS.n13830 4.5005
R15373 DVSS.n13876 DVSS.n13830 4.5005
R15374 DVSS.n13883 DVSS.n13830 4.5005
R15375 DVSS.n13875 DVSS.n13830 4.5005
R15376 DVSS.n13884 DVSS.n13830 4.5005
R15377 DVSS.n13874 DVSS.n13830 4.5005
R15378 DVSS.n13885 DVSS.n13830 4.5005
R15379 DVSS.n13887 DVSS.n13830 4.5005
R15380 DVSS.n21114 DVSS.n13830 4.5005
R15381 DVSS.n13844 DVSS.n13824 4.5005
R15382 DVSS.n21116 DVSS.n13844 4.5005
R15383 DVSS.n13878 DVSS.n13844 4.5005
R15384 DVSS.n13880 DVSS.n13844 4.5005
R15385 DVSS.n13877 DVSS.n13844 4.5005
R15386 DVSS.n13882 DVSS.n13844 4.5005
R15387 DVSS.n13876 DVSS.n13844 4.5005
R15388 DVSS.n13883 DVSS.n13844 4.5005
R15389 DVSS.n13875 DVSS.n13844 4.5005
R15390 DVSS.n13884 DVSS.n13844 4.5005
R15391 DVSS.n13874 DVSS.n13844 4.5005
R15392 DVSS.n13885 DVSS.n13844 4.5005
R15393 DVSS.n13887 DVSS.n13844 4.5005
R15394 DVSS.n21114 DVSS.n13844 4.5005
R15395 DVSS.n13829 DVSS.n13824 4.5005
R15396 DVSS.n21116 DVSS.n13829 4.5005
R15397 DVSS.n13878 DVSS.n13829 4.5005
R15398 DVSS.n13880 DVSS.n13829 4.5005
R15399 DVSS.n13877 DVSS.n13829 4.5005
R15400 DVSS.n13882 DVSS.n13829 4.5005
R15401 DVSS.n13876 DVSS.n13829 4.5005
R15402 DVSS.n13883 DVSS.n13829 4.5005
R15403 DVSS.n13875 DVSS.n13829 4.5005
R15404 DVSS.n13884 DVSS.n13829 4.5005
R15405 DVSS.n13874 DVSS.n13829 4.5005
R15406 DVSS.n13885 DVSS.n13829 4.5005
R15407 DVSS.n13887 DVSS.n13829 4.5005
R15408 DVSS.n21114 DVSS.n13829 4.5005
R15409 DVSS.n13845 DVSS.n13824 4.5005
R15410 DVSS.n21116 DVSS.n13845 4.5005
R15411 DVSS.n13878 DVSS.n13845 4.5005
R15412 DVSS.n13880 DVSS.n13845 4.5005
R15413 DVSS.n13877 DVSS.n13845 4.5005
R15414 DVSS.n13882 DVSS.n13845 4.5005
R15415 DVSS.n13876 DVSS.n13845 4.5005
R15416 DVSS.n13883 DVSS.n13845 4.5005
R15417 DVSS.n13875 DVSS.n13845 4.5005
R15418 DVSS.n13884 DVSS.n13845 4.5005
R15419 DVSS.n13874 DVSS.n13845 4.5005
R15420 DVSS.n13885 DVSS.n13845 4.5005
R15421 DVSS.n13887 DVSS.n13845 4.5005
R15422 DVSS.n21114 DVSS.n13845 4.5005
R15423 DVSS.n13828 DVSS.n13824 4.5005
R15424 DVSS.n21116 DVSS.n13828 4.5005
R15425 DVSS.n13878 DVSS.n13828 4.5005
R15426 DVSS.n13880 DVSS.n13828 4.5005
R15427 DVSS.n13877 DVSS.n13828 4.5005
R15428 DVSS.n13882 DVSS.n13828 4.5005
R15429 DVSS.n13876 DVSS.n13828 4.5005
R15430 DVSS.n13883 DVSS.n13828 4.5005
R15431 DVSS.n13875 DVSS.n13828 4.5005
R15432 DVSS.n13884 DVSS.n13828 4.5005
R15433 DVSS.n13874 DVSS.n13828 4.5005
R15434 DVSS.n13885 DVSS.n13828 4.5005
R15435 DVSS.n13887 DVSS.n13828 4.5005
R15436 DVSS.n21114 DVSS.n13828 4.5005
R15437 DVSS.n13846 DVSS.n13824 4.5005
R15438 DVSS.n21116 DVSS.n13846 4.5005
R15439 DVSS.n13878 DVSS.n13846 4.5005
R15440 DVSS.n13880 DVSS.n13846 4.5005
R15441 DVSS.n13877 DVSS.n13846 4.5005
R15442 DVSS.n13882 DVSS.n13846 4.5005
R15443 DVSS.n13876 DVSS.n13846 4.5005
R15444 DVSS.n13883 DVSS.n13846 4.5005
R15445 DVSS.n13875 DVSS.n13846 4.5005
R15446 DVSS.n13884 DVSS.n13846 4.5005
R15447 DVSS.n13874 DVSS.n13846 4.5005
R15448 DVSS.n13885 DVSS.n13846 4.5005
R15449 DVSS.n13887 DVSS.n13846 4.5005
R15450 DVSS.n21114 DVSS.n13846 4.5005
R15451 DVSS.n13827 DVSS.n13824 4.5005
R15452 DVSS.n21116 DVSS.n13827 4.5005
R15453 DVSS.n13878 DVSS.n13827 4.5005
R15454 DVSS.n13880 DVSS.n13827 4.5005
R15455 DVSS.n13877 DVSS.n13827 4.5005
R15456 DVSS.n13882 DVSS.n13827 4.5005
R15457 DVSS.n13876 DVSS.n13827 4.5005
R15458 DVSS.n13883 DVSS.n13827 4.5005
R15459 DVSS.n13875 DVSS.n13827 4.5005
R15460 DVSS.n13884 DVSS.n13827 4.5005
R15461 DVSS.n13874 DVSS.n13827 4.5005
R15462 DVSS.n13885 DVSS.n13827 4.5005
R15463 DVSS.n13887 DVSS.n13827 4.5005
R15464 DVSS.n21114 DVSS.n13827 4.5005
R15465 DVSS.n13847 DVSS.n13824 4.5005
R15466 DVSS.n21116 DVSS.n13847 4.5005
R15467 DVSS.n13878 DVSS.n13847 4.5005
R15468 DVSS.n13880 DVSS.n13847 4.5005
R15469 DVSS.n13877 DVSS.n13847 4.5005
R15470 DVSS.n13882 DVSS.n13847 4.5005
R15471 DVSS.n13876 DVSS.n13847 4.5005
R15472 DVSS.n13883 DVSS.n13847 4.5005
R15473 DVSS.n13875 DVSS.n13847 4.5005
R15474 DVSS.n13884 DVSS.n13847 4.5005
R15475 DVSS.n13874 DVSS.n13847 4.5005
R15476 DVSS.n13885 DVSS.n13847 4.5005
R15477 DVSS.n13887 DVSS.n13847 4.5005
R15478 DVSS.n21114 DVSS.n13847 4.5005
R15479 DVSS.n13826 DVSS.n13824 4.5005
R15480 DVSS.n21116 DVSS.n13826 4.5005
R15481 DVSS.n13878 DVSS.n13826 4.5005
R15482 DVSS.n13880 DVSS.n13826 4.5005
R15483 DVSS.n13877 DVSS.n13826 4.5005
R15484 DVSS.n13882 DVSS.n13826 4.5005
R15485 DVSS.n13876 DVSS.n13826 4.5005
R15486 DVSS.n13883 DVSS.n13826 4.5005
R15487 DVSS.n13875 DVSS.n13826 4.5005
R15488 DVSS.n13884 DVSS.n13826 4.5005
R15489 DVSS.n13874 DVSS.n13826 4.5005
R15490 DVSS.n13885 DVSS.n13826 4.5005
R15491 DVSS.n13887 DVSS.n13826 4.5005
R15492 DVSS.n21114 DVSS.n13826 4.5005
R15493 DVSS.n13848 DVSS.n13824 4.5005
R15494 DVSS.n21116 DVSS.n13848 4.5005
R15495 DVSS.n13878 DVSS.n13848 4.5005
R15496 DVSS.n13880 DVSS.n13848 4.5005
R15497 DVSS.n13877 DVSS.n13848 4.5005
R15498 DVSS.n13882 DVSS.n13848 4.5005
R15499 DVSS.n13876 DVSS.n13848 4.5005
R15500 DVSS.n13883 DVSS.n13848 4.5005
R15501 DVSS.n13875 DVSS.n13848 4.5005
R15502 DVSS.n13884 DVSS.n13848 4.5005
R15503 DVSS.n13874 DVSS.n13848 4.5005
R15504 DVSS.n13885 DVSS.n13848 4.5005
R15505 DVSS.n13887 DVSS.n13848 4.5005
R15506 DVSS.n21114 DVSS.n13848 4.5005
R15507 DVSS.n13825 DVSS.n13824 4.5005
R15508 DVSS.n21116 DVSS.n13825 4.5005
R15509 DVSS.n13878 DVSS.n13825 4.5005
R15510 DVSS.n13880 DVSS.n13825 4.5005
R15511 DVSS.n13877 DVSS.n13825 4.5005
R15512 DVSS.n13882 DVSS.n13825 4.5005
R15513 DVSS.n13876 DVSS.n13825 4.5005
R15514 DVSS.n13883 DVSS.n13825 4.5005
R15515 DVSS.n13875 DVSS.n13825 4.5005
R15516 DVSS.n13884 DVSS.n13825 4.5005
R15517 DVSS.n13874 DVSS.n13825 4.5005
R15518 DVSS.n13885 DVSS.n13825 4.5005
R15519 DVSS.n21114 DVSS.n13825 4.5005
R15520 DVSS.n21115 DVSS.n13824 4.5005
R15521 DVSS.n21116 DVSS.n21115 4.5005
R15522 DVSS.n21115 DVSS.n13878 4.5005
R15523 DVSS.n21115 DVSS.n13880 4.5005
R15524 DVSS.n21115 DVSS.n13877 4.5005
R15525 DVSS.n21115 DVSS.n13882 4.5005
R15526 DVSS.n21115 DVSS.n13876 4.5005
R15527 DVSS.n21115 DVSS.n13883 4.5005
R15528 DVSS.n21115 DVSS.n13875 4.5005
R15529 DVSS.n21115 DVSS.n13884 4.5005
R15530 DVSS.n21115 DVSS.n13874 4.5005
R15531 DVSS.n21115 DVSS.n13885 4.5005
R15532 DVSS.n21115 DVSS.n13873 4.5005
R15533 DVSS.n21115 DVSS.n13887 4.5005
R15534 DVSS.n21115 DVSS.n13861 4.5005
R15535 DVSS.n21115 DVSS.n21114 4.5005
R15536 DVSS.n20711 DVSS.n14512 4.5005
R15537 DVSS.n20712 DVSS.n14512 4.5005
R15538 DVSS.n20710 DVSS.n14512 4.5005
R15539 DVSS.n20713 DVSS.n14512 4.5005
R15540 DVSS.n20709 DVSS.n14512 4.5005
R15541 DVSS.n20716 DVSS.n14512 4.5005
R15542 DVSS.n20707 DVSS.n14512 4.5005
R15543 DVSS.n20717 DVSS.n14512 4.5005
R15544 DVSS.n20706 DVSS.n14512 4.5005
R15545 DVSS.n20718 DVSS.n14512 4.5005
R15546 DVSS.n20722 DVSS.n14512 4.5005
R15547 DVSS.n20805 DVSS.n14512 4.5005
R15548 DVSS.n20711 DVSS.n14511 4.5005
R15549 DVSS.n20712 DVSS.n14511 4.5005
R15550 DVSS.n20710 DVSS.n14511 4.5005
R15551 DVSS.n20713 DVSS.n14511 4.5005
R15552 DVSS.n20709 DVSS.n14511 4.5005
R15553 DVSS.n20715 DVSS.n14511 4.5005
R15554 DVSS.n20708 DVSS.n14511 4.5005
R15555 DVSS.n20716 DVSS.n14511 4.5005
R15556 DVSS.n20707 DVSS.n14511 4.5005
R15557 DVSS.n20717 DVSS.n14511 4.5005
R15558 DVSS.n20706 DVSS.n14511 4.5005
R15559 DVSS.n20718 DVSS.n14511 4.5005
R15560 DVSS.n20722 DVSS.n14511 4.5005
R15561 DVSS.n20803 DVSS.n14511 4.5005
R15562 DVSS.n20704 DVSS.n14511 4.5005
R15563 DVSS.n20805 DVSS.n14511 4.5005
R15564 DVSS.n20711 DVSS.n14513 4.5005
R15565 DVSS.n20712 DVSS.n14513 4.5005
R15566 DVSS.n20710 DVSS.n14513 4.5005
R15567 DVSS.n20713 DVSS.n14513 4.5005
R15568 DVSS.n20709 DVSS.n14513 4.5005
R15569 DVSS.n20715 DVSS.n14513 4.5005
R15570 DVSS.n20708 DVSS.n14513 4.5005
R15571 DVSS.n20716 DVSS.n14513 4.5005
R15572 DVSS.n20707 DVSS.n14513 4.5005
R15573 DVSS.n20717 DVSS.n14513 4.5005
R15574 DVSS.n20706 DVSS.n14513 4.5005
R15575 DVSS.n20718 DVSS.n14513 4.5005
R15576 DVSS.n20722 DVSS.n14513 4.5005
R15577 DVSS.n20803 DVSS.n14513 4.5005
R15578 DVSS.n20805 DVSS.n14513 4.5005
R15579 DVSS.n20711 DVSS.n14510 4.5005
R15580 DVSS.n20712 DVSS.n14510 4.5005
R15581 DVSS.n20710 DVSS.n14510 4.5005
R15582 DVSS.n20713 DVSS.n14510 4.5005
R15583 DVSS.n20709 DVSS.n14510 4.5005
R15584 DVSS.n20715 DVSS.n14510 4.5005
R15585 DVSS.n20708 DVSS.n14510 4.5005
R15586 DVSS.n20716 DVSS.n14510 4.5005
R15587 DVSS.n20707 DVSS.n14510 4.5005
R15588 DVSS.n20717 DVSS.n14510 4.5005
R15589 DVSS.n20706 DVSS.n14510 4.5005
R15590 DVSS.n20718 DVSS.n14510 4.5005
R15591 DVSS.n20803 DVSS.n14510 4.5005
R15592 DVSS.n20805 DVSS.n14510 4.5005
R15593 DVSS.n20711 DVSS.n14514 4.5005
R15594 DVSS.n20712 DVSS.n14514 4.5005
R15595 DVSS.n20710 DVSS.n14514 4.5005
R15596 DVSS.n20713 DVSS.n14514 4.5005
R15597 DVSS.n20709 DVSS.n14514 4.5005
R15598 DVSS.n20715 DVSS.n14514 4.5005
R15599 DVSS.n20708 DVSS.n14514 4.5005
R15600 DVSS.n20716 DVSS.n14514 4.5005
R15601 DVSS.n20707 DVSS.n14514 4.5005
R15602 DVSS.n20717 DVSS.n14514 4.5005
R15603 DVSS.n20706 DVSS.n14514 4.5005
R15604 DVSS.n20718 DVSS.n14514 4.5005
R15605 DVSS.n20803 DVSS.n14514 4.5005
R15606 DVSS.n20805 DVSS.n14514 4.5005
R15607 DVSS.n20711 DVSS.n14509 4.5005
R15608 DVSS.n20712 DVSS.n14509 4.5005
R15609 DVSS.n20710 DVSS.n14509 4.5005
R15610 DVSS.n20713 DVSS.n14509 4.5005
R15611 DVSS.n20709 DVSS.n14509 4.5005
R15612 DVSS.n20715 DVSS.n14509 4.5005
R15613 DVSS.n20708 DVSS.n14509 4.5005
R15614 DVSS.n20716 DVSS.n14509 4.5005
R15615 DVSS.n20707 DVSS.n14509 4.5005
R15616 DVSS.n20717 DVSS.n14509 4.5005
R15617 DVSS.n20706 DVSS.n14509 4.5005
R15618 DVSS.n20718 DVSS.n14509 4.5005
R15619 DVSS.n20803 DVSS.n14509 4.5005
R15620 DVSS.n20805 DVSS.n14509 4.5005
R15621 DVSS.n20711 DVSS.n14515 4.5005
R15622 DVSS.n20712 DVSS.n14515 4.5005
R15623 DVSS.n20710 DVSS.n14515 4.5005
R15624 DVSS.n20713 DVSS.n14515 4.5005
R15625 DVSS.n20709 DVSS.n14515 4.5005
R15626 DVSS.n20715 DVSS.n14515 4.5005
R15627 DVSS.n20708 DVSS.n14515 4.5005
R15628 DVSS.n20716 DVSS.n14515 4.5005
R15629 DVSS.n20707 DVSS.n14515 4.5005
R15630 DVSS.n20717 DVSS.n14515 4.5005
R15631 DVSS.n20706 DVSS.n14515 4.5005
R15632 DVSS.n20718 DVSS.n14515 4.5005
R15633 DVSS.n20803 DVSS.n14515 4.5005
R15634 DVSS.n20805 DVSS.n14515 4.5005
R15635 DVSS.n20711 DVSS.n14508 4.5005
R15636 DVSS.n20712 DVSS.n14508 4.5005
R15637 DVSS.n20710 DVSS.n14508 4.5005
R15638 DVSS.n20713 DVSS.n14508 4.5005
R15639 DVSS.n20709 DVSS.n14508 4.5005
R15640 DVSS.n20715 DVSS.n14508 4.5005
R15641 DVSS.n20708 DVSS.n14508 4.5005
R15642 DVSS.n20716 DVSS.n14508 4.5005
R15643 DVSS.n20707 DVSS.n14508 4.5005
R15644 DVSS.n20717 DVSS.n14508 4.5005
R15645 DVSS.n20706 DVSS.n14508 4.5005
R15646 DVSS.n20718 DVSS.n14508 4.5005
R15647 DVSS.n20803 DVSS.n14508 4.5005
R15648 DVSS.n20805 DVSS.n14508 4.5005
R15649 DVSS.n20711 DVSS.n14516 4.5005
R15650 DVSS.n20712 DVSS.n14516 4.5005
R15651 DVSS.n20710 DVSS.n14516 4.5005
R15652 DVSS.n20713 DVSS.n14516 4.5005
R15653 DVSS.n20709 DVSS.n14516 4.5005
R15654 DVSS.n20715 DVSS.n14516 4.5005
R15655 DVSS.n20708 DVSS.n14516 4.5005
R15656 DVSS.n20716 DVSS.n14516 4.5005
R15657 DVSS.n20707 DVSS.n14516 4.5005
R15658 DVSS.n20717 DVSS.n14516 4.5005
R15659 DVSS.n20706 DVSS.n14516 4.5005
R15660 DVSS.n20718 DVSS.n14516 4.5005
R15661 DVSS.n20803 DVSS.n14516 4.5005
R15662 DVSS.n20805 DVSS.n14516 4.5005
R15663 DVSS.n20711 DVSS.n14507 4.5005
R15664 DVSS.n20712 DVSS.n14507 4.5005
R15665 DVSS.n20710 DVSS.n14507 4.5005
R15666 DVSS.n20713 DVSS.n14507 4.5005
R15667 DVSS.n20709 DVSS.n14507 4.5005
R15668 DVSS.n20715 DVSS.n14507 4.5005
R15669 DVSS.n20708 DVSS.n14507 4.5005
R15670 DVSS.n20716 DVSS.n14507 4.5005
R15671 DVSS.n20707 DVSS.n14507 4.5005
R15672 DVSS.n20717 DVSS.n14507 4.5005
R15673 DVSS.n20706 DVSS.n14507 4.5005
R15674 DVSS.n20718 DVSS.n14507 4.5005
R15675 DVSS.n20803 DVSS.n14507 4.5005
R15676 DVSS.n20805 DVSS.n14507 4.5005
R15677 DVSS.n20804 DVSS.n20711 4.5005
R15678 DVSS.n20804 DVSS.n20712 4.5005
R15679 DVSS.n20804 DVSS.n20710 4.5005
R15680 DVSS.n20804 DVSS.n20713 4.5005
R15681 DVSS.n20804 DVSS.n20709 4.5005
R15682 DVSS.n20804 DVSS.n20715 4.5005
R15683 DVSS.n20804 DVSS.n20708 4.5005
R15684 DVSS.n20804 DVSS.n20716 4.5005
R15685 DVSS.n20804 DVSS.n20707 4.5005
R15686 DVSS.n20804 DVSS.n20717 4.5005
R15687 DVSS.n20804 DVSS.n20706 4.5005
R15688 DVSS.n20804 DVSS.n20718 4.5005
R15689 DVSS.n20804 DVSS.n20803 4.5005
R15690 DVSS.n20804 DVSS.n20704 4.5005
R15691 DVSS.n20805 DVSS.n20804 4.5005
R15692 DVSS.n15223 DVSS.n14536 4.5005
R15693 DVSS.n15228 DVSS.n14536 4.5005
R15694 DVSS.n18474 DVSS.n14536 4.5005
R15695 DVSS.n18387 DVSS.n14536 4.5005
R15696 DVSS.n18386 DVSS.n14536 4.5005
R15697 DVSS.n18390 DVSS.n14536 4.5005
R15698 DVSS.n18384 DVSS.n14536 4.5005
R15699 DVSS.n18391 DVSS.n14536 4.5005
R15700 DVSS.n18383 DVSS.n14536 4.5005
R15701 DVSS.n18392 DVSS.n14536 4.5005
R15702 DVSS.n18432 DVSS.n14536 4.5005
R15703 DVSS.n18433 DVSS.n14536 4.5005
R15704 DVSS.n18472 DVSS.n14536 4.5005
R15705 DVSS.n15233 DVSS.n15223 4.5005
R15706 DVSS.n15233 DVSS.n15228 4.5005
R15707 DVSS.n18474 DVSS.n15233 4.5005
R15708 DVSS.n18387 DVSS.n15233 4.5005
R15709 DVSS.n18386 DVSS.n15233 4.5005
R15710 DVSS.n18389 DVSS.n15233 4.5005
R15711 DVSS.n18385 DVSS.n15233 4.5005
R15712 DVSS.n18390 DVSS.n15233 4.5005
R15713 DVSS.n18384 DVSS.n15233 4.5005
R15714 DVSS.n18391 DVSS.n15233 4.5005
R15715 DVSS.n18383 DVSS.n15233 4.5005
R15716 DVSS.n18392 DVSS.n15233 4.5005
R15717 DVSS.n18433 DVSS.n15233 4.5005
R15718 DVSS.n18472 DVSS.n15233 4.5005
R15719 DVSS.n15235 DVSS.n15223 4.5005
R15720 DVSS.n15235 DVSS.n15228 4.5005
R15721 DVSS.n18474 DVSS.n15235 4.5005
R15722 DVSS.n18387 DVSS.n15235 4.5005
R15723 DVSS.n18386 DVSS.n15235 4.5005
R15724 DVSS.n18389 DVSS.n15235 4.5005
R15725 DVSS.n18385 DVSS.n15235 4.5005
R15726 DVSS.n18390 DVSS.n15235 4.5005
R15727 DVSS.n18384 DVSS.n15235 4.5005
R15728 DVSS.n18391 DVSS.n15235 4.5005
R15729 DVSS.n18383 DVSS.n15235 4.5005
R15730 DVSS.n18392 DVSS.n15235 4.5005
R15731 DVSS.n18433 DVSS.n15235 4.5005
R15732 DVSS.n18472 DVSS.n15235 4.5005
R15733 DVSS.n15232 DVSS.n15223 4.5005
R15734 DVSS.n15232 DVSS.n15228 4.5005
R15735 DVSS.n18474 DVSS.n15232 4.5005
R15736 DVSS.n18387 DVSS.n15232 4.5005
R15737 DVSS.n18386 DVSS.n15232 4.5005
R15738 DVSS.n18389 DVSS.n15232 4.5005
R15739 DVSS.n18385 DVSS.n15232 4.5005
R15740 DVSS.n18390 DVSS.n15232 4.5005
R15741 DVSS.n18384 DVSS.n15232 4.5005
R15742 DVSS.n18391 DVSS.n15232 4.5005
R15743 DVSS.n18383 DVSS.n15232 4.5005
R15744 DVSS.n18392 DVSS.n15232 4.5005
R15745 DVSS.n18433 DVSS.n15232 4.5005
R15746 DVSS.n18472 DVSS.n15232 4.5005
R15747 DVSS.n15236 DVSS.n15223 4.5005
R15748 DVSS.n15236 DVSS.n15228 4.5005
R15749 DVSS.n18474 DVSS.n15236 4.5005
R15750 DVSS.n18387 DVSS.n15236 4.5005
R15751 DVSS.n18386 DVSS.n15236 4.5005
R15752 DVSS.n18389 DVSS.n15236 4.5005
R15753 DVSS.n18385 DVSS.n15236 4.5005
R15754 DVSS.n18390 DVSS.n15236 4.5005
R15755 DVSS.n18384 DVSS.n15236 4.5005
R15756 DVSS.n18391 DVSS.n15236 4.5005
R15757 DVSS.n18383 DVSS.n15236 4.5005
R15758 DVSS.n18392 DVSS.n15236 4.5005
R15759 DVSS.n18433 DVSS.n15236 4.5005
R15760 DVSS.n18472 DVSS.n15236 4.5005
R15761 DVSS.n15231 DVSS.n15223 4.5005
R15762 DVSS.n15231 DVSS.n15228 4.5005
R15763 DVSS.n18474 DVSS.n15231 4.5005
R15764 DVSS.n18387 DVSS.n15231 4.5005
R15765 DVSS.n18386 DVSS.n15231 4.5005
R15766 DVSS.n18389 DVSS.n15231 4.5005
R15767 DVSS.n18385 DVSS.n15231 4.5005
R15768 DVSS.n18390 DVSS.n15231 4.5005
R15769 DVSS.n18384 DVSS.n15231 4.5005
R15770 DVSS.n18391 DVSS.n15231 4.5005
R15771 DVSS.n18383 DVSS.n15231 4.5005
R15772 DVSS.n18392 DVSS.n15231 4.5005
R15773 DVSS.n18433 DVSS.n15231 4.5005
R15774 DVSS.n18472 DVSS.n15231 4.5005
R15775 DVSS.n15237 DVSS.n15223 4.5005
R15776 DVSS.n15237 DVSS.n15228 4.5005
R15777 DVSS.n18474 DVSS.n15237 4.5005
R15778 DVSS.n18387 DVSS.n15237 4.5005
R15779 DVSS.n18386 DVSS.n15237 4.5005
R15780 DVSS.n18389 DVSS.n15237 4.5005
R15781 DVSS.n18385 DVSS.n15237 4.5005
R15782 DVSS.n18390 DVSS.n15237 4.5005
R15783 DVSS.n18384 DVSS.n15237 4.5005
R15784 DVSS.n18391 DVSS.n15237 4.5005
R15785 DVSS.n18383 DVSS.n15237 4.5005
R15786 DVSS.n18392 DVSS.n15237 4.5005
R15787 DVSS.n18433 DVSS.n15237 4.5005
R15788 DVSS.n18472 DVSS.n15237 4.5005
R15789 DVSS.n15230 DVSS.n15223 4.5005
R15790 DVSS.n15230 DVSS.n15228 4.5005
R15791 DVSS.n18474 DVSS.n15230 4.5005
R15792 DVSS.n18387 DVSS.n15230 4.5005
R15793 DVSS.n18386 DVSS.n15230 4.5005
R15794 DVSS.n18389 DVSS.n15230 4.5005
R15795 DVSS.n18385 DVSS.n15230 4.5005
R15796 DVSS.n18390 DVSS.n15230 4.5005
R15797 DVSS.n18384 DVSS.n15230 4.5005
R15798 DVSS.n18391 DVSS.n15230 4.5005
R15799 DVSS.n18383 DVSS.n15230 4.5005
R15800 DVSS.n18392 DVSS.n15230 4.5005
R15801 DVSS.n18433 DVSS.n15230 4.5005
R15802 DVSS.n18472 DVSS.n15230 4.5005
R15803 DVSS.n15238 DVSS.n15223 4.5005
R15804 DVSS.n15238 DVSS.n15228 4.5005
R15805 DVSS.n18474 DVSS.n15238 4.5005
R15806 DVSS.n18387 DVSS.n15238 4.5005
R15807 DVSS.n18386 DVSS.n15238 4.5005
R15808 DVSS.n18389 DVSS.n15238 4.5005
R15809 DVSS.n18385 DVSS.n15238 4.5005
R15810 DVSS.n18390 DVSS.n15238 4.5005
R15811 DVSS.n18384 DVSS.n15238 4.5005
R15812 DVSS.n18391 DVSS.n15238 4.5005
R15813 DVSS.n18383 DVSS.n15238 4.5005
R15814 DVSS.n18392 DVSS.n15238 4.5005
R15815 DVSS.n18433 DVSS.n15238 4.5005
R15816 DVSS.n18472 DVSS.n15238 4.5005
R15817 DVSS.n15229 DVSS.n15223 4.5005
R15818 DVSS.n15229 DVSS.n15228 4.5005
R15819 DVSS.n18474 DVSS.n15229 4.5005
R15820 DVSS.n18387 DVSS.n15229 4.5005
R15821 DVSS.n18386 DVSS.n15229 4.5005
R15822 DVSS.n18389 DVSS.n15229 4.5005
R15823 DVSS.n18385 DVSS.n15229 4.5005
R15824 DVSS.n18390 DVSS.n15229 4.5005
R15825 DVSS.n18384 DVSS.n15229 4.5005
R15826 DVSS.n18391 DVSS.n15229 4.5005
R15827 DVSS.n18383 DVSS.n15229 4.5005
R15828 DVSS.n18392 DVSS.n15229 4.5005
R15829 DVSS.n18433 DVSS.n15229 4.5005
R15830 DVSS.n18472 DVSS.n15229 4.5005
R15831 DVSS.n18473 DVSS.n15223 4.5005
R15832 DVSS.n18473 DVSS.n15228 4.5005
R15833 DVSS.n18474 DVSS.n18473 4.5005
R15834 DVSS.n18473 DVSS.n18387 4.5005
R15835 DVSS.n18473 DVSS.n18386 4.5005
R15836 DVSS.n18473 DVSS.n18389 4.5005
R15837 DVSS.n18473 DVSS.n18385 4.5005
R15838 DVSS.n18473 DVSS.n18390 4.5005
R15839 DVSS.n18473 DVSS.n18384 4.5005
R15840 DVSS.n18473 DVSS.n18391 4.5005
R15841 DVSS.n18473 DVSS.n18383 4.5005
R15842 DVSS.n18473 DVSS.n18392 4.5005
R15843 DVSS.n18473 DVSS.n18472 4.5005
R15844 DVSS.n18381 DVSS.n15246 4.5005
R15845 DVSS.n18381 DVSS.n15247 4.5005
R15846 DVSS.n18381 DVSS.n15245 4.5005
R15847 DVSS.n18381 DVSS.n15248 4.5005
R15848 DVSS.n18381 DVSS.n15244 4.5005
R15849 DVSS.n18381 DVSS.n15249 4.5005
R15850 DVSS.n18381 DVSS.n15242 4.5005
R15851 DVSS.n18381 DVSS.n15250 4.5005
R15852 DVSS.n18381 DVSS.n15241 4.5005
R15853 DVSS.n18381 DVSS.n15251 4.5005
R15854 DVSS.n18381 DVSS.n15240 4.5005
R15855 DVSS.n18381 DVSS.n15252 4.5005
R15856 DVSS.n18381 DVSS.n18380 4.5005
R15857 DVSS.n15258 DVSS.n15246 4.5005
R15858 DVSS.n15258 DVSS.n15247 4.5005
R15859 DVSS.n15258 DVSS.n15245 4.5005
R15860 DVSS.n15258 DVSS.n15248 4.5005
R15861 DVSS.n15258 DVSS.n15244 4.5005
R15862 DVSS.n18378 DVSS.n15258 4.5005
R15863 DVSS.n15272 DVSS.n15258 4.5005
R15864 DVSS.n15258 DVSS.n15249 4.5005
R15865 DVSS.n15258 DVSS.n15242 4.5005
R15866 DVSS.n15258 DVSS.n15250 4.5005
R15867 DVSS.n15258 DVSS.n15241 4.5005
R15868 DVSS.n15258 DVSS.n15251 4.5005
R15869 DVSS.n15258 DVSS.n15240 4.5005
R15870 DVSS.n15258 DVSS.n15252 4.5005
R15871 DVSS.n18380 DVSS.n15258 4.5005
R15872 DVSS.n15261 DVSS.n15246 4.5005
R15873 DVSS.n15261 DVSS.n15247 4.5005
R15874 DVSS.n15261 DVSS.n15245 4.5005
R15875 DVSS.n15261 DVSS.n15248 4.5005
R15876 DVSS.n15261 DVSS.n15244 4.5005
R15877 DVSS.n18378 DVSS.n15261 4.5005
R15878 DVSS.n15272 DVSS.n15261 4.5005
R15879 DVSS.n15261 DVSS.n15249 4.5005
R15880 DVSS.n15261 DVSS.n15242 4.5005
R15881 DVSS.n15261 DVSS.n15250 4.5005
R15882 DVSS.n15261 DVSS.n15241 4.5005
R15883 DVSS.n15261 DVSS.n15251 4.5005
R15884 DVSS.n15261 DVSS.n15252 4.5005
R15885 DVSS.n18380 DVSS.n15261 4.5005
R15886 DVSS.n15257 DVSS.n15246 4.5005
R15887 DVSS.n15257 DVSS.n15247 4.5005
R15888 DVSS.n15257 DVSS.n15245 4.5005
R15889 DVSS.n15257 DVSS.n15248 4.5005
R15890 DVSS.n15257 DVSS.n15244 4.5005
R15891 DVSS.n18378 DVSS.n15257 4.5005
R15892 DVSS.n15272 DVSS.n15257 4.5005
R15893 DVSS.n15257 DVSS.n15249 4.5005
R15894 DVSS.n15257 DVSS.n15242 4.5005
R15895 DVSS.n15257 DVSS.n15250 4.5005
R15896 DVSS.n15257 DVSS.n15241 4.5005
R15897 DVSS.n15257 DVSS.n15251 4.5005
R15898 DVSS.n15257 DVSS.n15252 4.5005
R15899 DVSS.n18380 DVSS.n15257 4.5005
R15900 DVSS.n15263 DVSS.n15246 4.5005
R15901 DVSS.n15263 DVSS.n15247 4.5005
R15902 DVSS.n15263 DVSS.n15245 4.5005
R15903 DVSS.n15263 DVSS.n15248 4.5005
R15904 DVSS.n15263 DVSS.n15244 4.5005
R15905 DVSS.n18378 DVSS.n15263 4.5005
R15906 DVSS.n15272 DVSS.n15263 4.5005
R15907 DVSS.n15263 DVSS.n15249 4.5005
R15908 DVSS.n15263 DVSS.n15242 4.5005
R15909 DVSS.n15263 DVSS.n15250 4.5005
R15910 DVSS.n15263 DVSS.n15241 4.5005
R15911 DVSS.n15263 DVSS.n15251 4.5005
R15912 DVSS.n15263 DVSS.n15252 4.5005
R15913 DVSS.n18380 DVSS.n15263 4.5005
R15914 DVSS.n15256 DVSS.n15246 4.5005
R15915 DVSS.n15256 DVSS.n15247 4.5005
R15916 DVSS.n15256 DVSS.n15245 4.5005
R15917 DVSS.n15256 DVSS.n15248 4.5005
R15918 DVSS.n15256 DVSS.n15244 4.5005
R15919 DVSS.n18378 DVSS.n15256 4.5005
R15920 DVSS.n15272 DVSS.n15256 4.5005
R15921 DVSS.n15256 DVSS.n15249 4.5005
R15922 DVSS.n15256 DVSS.n15242 4.5005
R15923 DVSS.n15256 DVSS.n15250 4.5005
R15924 DVSS.n15256 DVSS.n15241 4.5005
R15925 DVSS.n15256 DVSS.n15251 4.5005
R15926 DVSS.n15256 DVSS.n15252 4.5005
R15927 DVSS.n18380 DVSS.n15256 4.5005
R15928 DVSS.n15265 DVSS.n15246 4.5005
R15929 DVSS.n15265 DVSS.n15247 4.5005
R15930 DVSS.n15265 DVSS.n15245 4.5005
R15931 DVSS.n15265 DVSS.n15248 4.5005
R15932 DVSS.n15265 DVSS.n15244 4.5005
R15933 DVSS.n18378 DVSS.n15265 4.5005
R15934 DVSS.n15272 DVSS.n15265 4.5005
R15935 DVSS.n15265 DVSS.n15249 4.5005
R15936 DVSS.n15265 DVSS.n15242 4.5005
R15937 DVSS.n15265 DVSS.n15250 4.5005
R15938 DVSS.n15265 DVSS.n15241 4.5005
R15939 DVSS.n15265 DVSS.n15251 4.5005
R15940 DVSS.n18380 DVSS.n15265 4.5005
R15941 DVSS.n15255 DVSS.n15246 4.5005
R15942 DVSS.n15255 DVSS.n15247 4.5005
R15943 DVSS.n15255 DVSS.n15245 4.5005
R15944 DVSS.n15255 DVSS.n15248 4.5005
R15945 DVSS.n15255 DVSS.n15244 4.5005
R15946 DVSS.n18378 DVSS.n15255 4.5005
R15947 DVSS.n15272 DVSS.n15255 4.5005
R15948 DVSS.n15255 DVSS.n15249 4.5005
R15949 DVSS.n15255 DVSS.n15242 4.5005
R15950 DVSS.n15255 DVSS.n15250 4.5005
R15951 DVSS.n15255 DVSS.n15241 4.5005
R15952 DVSS.n15255 DVSS.n15251 4.5005
R15953 DVSS.n15255 DVSS.n15240 4.5005
R15954 DVSS.n15255 DVSS.n15252 4.5005
R15955 DVSS.n15271 DVSS.n15255 4.5005
R15956 DVSS.n18380 DVSS.n15255 4.5005
R15957 DVSS.n16000 DVSS.n15993 4.5005
R15958 DVSS.n17655 DVSS.n16000 4.5005
R15959 DVSS.n16020 DVSS.n16000 4.5005
R15960 DVSS.n16022 DVSS.n16000 4.5005
R15961 DVSS.n16019 DVSS.n16000 4.5005
R15962 DVSS.n16025 DVSS.n16000 4.5005
R15963 DVSS.n16017 DVSS.n16000 4.5005
R15964 DVSS.n16026 DVSS.n16000 4.5005
R15965 DVSS.n16016 DVSS.n16000 4.5005
R15966 DVSS.n16027 DVSS.n16000 4.5005
R15967 DVSS.n16015 DVSS.n16000 4.5005
R15968 DVSS.n16029 DVSS.n16000 4.5005
R15969 DVSS.n17653 DVSS.n16000 4.5005
R15970 DVSS.n15998 DVSS.n15993 4.5005
R15971 DVSS.n17655 DVSS.n15998 4.5005
R15972 DVSS.n16020 DVSS.n15998 4.5005
R15973 DVSS.n16022 DVSS.n15998 4.5005
R15974 DVSS.n16019 DVSS.n15998 4.5005
R15975 DVSS.n16024 DVSS.n15998 4.5005
R15976 DVSS.n16018 DVSS.n15998 4.5005
R15977 DVSS.n16025 DVSS.n15998 4.5005
R15978 DVSS.n16017 DVSS.n15998 4.5005
R15979 DVSS.n16026 DVSS.n15998 4.5005
R15980 DVSS.n16016 DVSS.n15998 4.5005
R15981 DVSS.n16027 DVSS.n15998 4.5005
R15982 DVSS.n16029 DVSS.n15998 4.5005
R15983 DVSS.n17653 DVSS.n15998 4.5005
R15984 DVSS.n16001 DVSS.n15993 4.5005
R15985 DVSS.n17655 DVSS.n16001 4.5005
R15986 DVSS.n16020 DVSS.n16001 4.5005
R15987 DVSS.n16022 DVSS.n16001 4.5005
R15988 DVSS.n16019 DVSS.n16001 4.5005
R15989 DVSS.n16024 DVSS.n16001 4.5005
R15990 DVSS.n16018 DVSS.n16001 4.5005
R15991 DVSS.n16025 DVSS.n16001 4.5005
R15992 DVSS.n16017 DVSS.n16001 4.5005
R15993 DVSS.n16026 DVSS.n16001 4.5005
R15994 DVSS.n16016 DVSS.n16001 4.5005
R15995 DVSS.n16027 DVSS.n16001 4.5005
R15996 DVSS.n16029 DVSS.n16001 4.5005
R15997 DVSS.n17653 DVSS.n16001 4.5005
R15998 DVSS.n15997 DVSS.n15993 4.5005
R15999 DVSS.n17655 DVSS.n15997 4.5005
R16000 DVSS.n16020 DVSS.n15997 4.5005
R16001 DVSS.n16022 DVSS.n15997 4.5005
R16002 DVSS.n16019 DVSS.n15997 4.5005
R16003 DVSS.n16024 DVSS.n15997 4.5005
R16004 DVSS.n16018 DVSS.n15997 4.5005
R16005 DVSS.n16025 DVSS.n15997 4.5005
R16006 DVSS.n16017 DVSS.n15997 4.5005
R16007 DVSS.n16026 DVSS.n15997 4.5005
R16008 DVSS.n16016 DVSS.n15997 4.5005
R16009 DVSS.n16027 DVSS.n15997 4.5005
R16010 DVSS.n16029 DVSS.n15997 4.5005
R16011 DVSS.n17653 DVSS.n15997 4.5005
R16012 DVSS.n16002 DVSS.n15993 4.5005
R16013 DVSS.n17655 DVSS.n16002 4.5005
R16014 DVSS.n16020 DVSS.n16002 4.5005
R16015 DVSS.n16022 DVSS.n16002 4.5005
R16016 DVSS.n16019 DVSS.n16002 4.5005
R16017 DVSS.n16024 DVSS.n16002 4.5005
R16018 DVSS.n16018 DVSS.n16002 4.5005
R16019 DVSS.n16025 DVSS.n16002 4.5005
R16020 DVSS.n16017 DVSS.n16002 4.5005
R16021 DVSS.n16026 DVSS.n16002 4.5005
R16022 DVSS.n16016 DVSS.n16002 4.5005
R16023 DVSS.n16027 DVSS.n16002 4.5005
R16024 DVSS.n17653 DVSS.n16002 4.5005
R16025 DVSS.n15996 DVSS.n15993 4.5005
R16026 DVSS.n17655 DVSS.n15996 4.5005
R16027 DVSS.n16020 DVSS.n15996 4.5005
R16028 DVSS.n16022 DVSS.n15996 4.5005
R16029 DVSS.n16019 DVSS.n15996 4.5005
R16030 DVSS.n16024 DVSS.n15996 4.5005
R16031 DVSS.n16018 DVSS.n15996 4.5005
R16032 DVSS.n16025 DVSS.n15996 4.5005
R16033 DVSS.n16017 DVSS.n15996 4.5005
R16034 DVSS.n16026 DVSS.n15996 4.5005
R16035 DVSS.n16016 DVSS.n15996 4.5005
R16036 DVSS.n16027 DVSS.n15996 4.5005
R16037 DVSS.n16029 DVSS.n15996 4.5005
R16038 DVSS.n17653 DVSS.n15996 4.5005
R16039 DVSS.n16003 DVSS.n15993 4.5005
R16040 DVSS.n17655 DVSS.n16003 4.5005
R16041 DVSS.n16020 DVSS.n16003 4.5005
R16042 DVSS.n16022 DVSS.n16003 4.5005
R16043 DVSS.n16019 DVSS.n16003 4.5005
R16044 DVSS.n16024 DVSS.n16003 4.5005
R16045 DVSS.n16018 DVSS.n16003 4.5005
R16046 DVSS.n16025 DVSS.n16003 4.5005
R16047 DVSS.n16017 DVSS.n16003 4.5005
R16048 DVSS.n16026 DVSS.n16003 4.5005
R16049 DVSS.n16016 DVSS.n16003 4.5005
R16050 DVSS.n16027 DVSS.n16003 4.5005
R16051 DVSS.n16029 DVSS.n16003 4.5005
R16052 DVSS.n17653 DVSS.n16003 4.5005
R16053 DVSS.n15995 DVSS.n15993 4.5005
R16054 DVSS.n17655 DVSS.n15995 4.5005
R16055 DVSS.n16020 DVSS.n15995 4.5005
R16056 DVSS.n16022 DVSS.n15995 4.5005
R16057 DVSS.n16019 DVSS.n15995 4.5005
R16058 DVSS.n16024 DVSS.n15995 4.5005
R16059 DVSS.n16018 DVSS.n15995 4.5005
R16060 DVSS.n16025 DVSS.n15995 4.5005
R16061 DVSS.n16017 DVSS.n15995 4.5005
R16062 DVSS.n16026 DVSS.n15995 4.5005
R16063 DVSS.n16016 DVSS.n15995 4.5005
R16064 DVSS.n16027 DVSS.n15995 4.5005
R16065 DVSS.n16029 DVSS.n15995 4.5005
R16066 DVSS.n17653 DVSS.n15995 4.5005
R16067 DVSS.n16004 DVSS.n15993 4.5005
R16068 DVSS.n17655 DVSS.n16004 4.5005
R16069 DVSS.n16020 DVSS.n16004 4.5005
R16070 DVSS.n16022 DVSS.n16004 4.5005
R16071 DVSS.n16019 DVSS.n16004 4.5005
R16072 DVSS.n16024 DVSS.n16004 4.5005
R16073 DVSS.n16018 DVSS.n16004 4.5005
R16074 DVSS.n16025 DVSS.n16004 4.5005
R16075 DVSS.n16017 DVSS.n16004 4.5005
R16076 DVSS.n16026 DVSS.n16004 4.5005
R16077 DVSS.n16016 DVSS.n16004 4.5005
R16078 DVSS.n16027 DVSS.n16004 4.5005
R16079 DVSS.n16015 DVSS.n16004 4.5005
R16080 DVSS.n16029 DVSS.n16004 4.5005
R16081 DVSS.n17653 DVSS.n16004 4.5005
R16082 DVSS.n16312 DVSS.n16299 4.5005
R16083 DVSS.n16314 DVSS.n16299 4.5005
R16084 DVSS.n16311 DVSS.n16299 4.5005
R16085 DVSS.n16315 DVSS.n16299 4.5005
R16086 DVSS.n16310 DVSS.n16299 4.5005
R16087 DVSS.n16318 DVSS.n16299 4.5005
R16088 DVSS.n16308 DVSS.n16299 4.5005
R16089 DVSS.n16319 DVSS.n16299 4.5005
R16090 DVSS.n16307 DVSS.n16299 4.5005
R16091 DVSS.n16634 DVSS.n16299 4.5005
R16092 DVSS.n16306 DVSS.n16299 4.5005
R16093 DVSS.n16637 DVSS.n16299 4.5005
R16094 DVSS.n16639 DVSS.n16299 4.5005
R16095 DVSS.n16312 DVSS.n16297 4.5005
R16096 DVSS.n16314 DVSS.n16297 4.5005
R16097 DVSS.n16311 DVSS.n16297 4.5005
R16098 DVSS.n16315 DVSS.n16297 4.5005
R16099 DVSS.n16310 DVSS.n16297 4.5005
R16100 DVSS.n16317 DVSS.n16297 4.5005
R16101 DVSS.n16309 DVSS.n16297 4.5005
R16102 DVSS.n16318 DVSS.n16297 4.5005
R16103 DVSS.n16308 DVSS.n16297 4.5005
R16104 DVSS.n16319 DVSS.n16297 4.5005
R16105 DVSS.n16307 DVSS.n16297 4.5005
R16106 DVSS.n16634 DVSS.n16297 4.5005
R16107 DVSS.n16637 DVSS.n16297 4.5005
R16108 DVSS.n16639 DVSS.n16297 4.5005
R16109 DVSS.n16312 DVSS.n16300 4.5005
R16110 DVSS.n16314 DVSS.n16300 4.5005
R16111 DVSS.n16311 DVSS.n16300 4.5005
R16112 DVSS.n16315 DVSS.n16300 4.5005
R16113 DVSS.n16310 DVSS.n16300 4.5005
R16114 DVSS.n16317 DVSS.n16300 4.5005
R16115 DVSS.n16309 DVSS.n16300 4.5005
R16116 DVSS.n16318 DVSS.n16300 4.5005
R16117 DVSS.n16308 DVSS.n16300 4.5005
R16118 DVSS.n16319 DVSS.n16300 4.5005
R16119 DVSS.n16307 DVSS.n16300 4.5005
R16120 DVSS.n16634 DVSS.n16300 4.5005
R16121 DVSS.n16639 DVSS.n16300 4.5005
R16122 DVSS.n16308 DVSS.n16296 4.5005
R16123 DVSS.n16319 DVSS.n16296 4.5005
R16124 DVSS.n16307 DVSS.n16296 4.5005
R16125 DVSS.n16634 DVSS.n16296 4.5005
R16126 DVSS.n16306 DVSS.n16296 4.5005
R16127 DVSS.n16637 DVSS.n16296 4.5005
R16128 DVSS.n16296 DVSS.n16292 4.5005
R16129 DVSS.n16639 DVSS.n16296 4.5005
R16130 DVSS.n16308 DVSS.n16301 4.5005
R16131 DVSS.n16319 DVSS.n16301 4.5005
R16132 DVSS.n16307 DVSS.n16301 4.5005
R16133 DVSS.n16634 DVSS.n16301 4.5005
R16134 DVSS.n16306 DVSS.n16301 4.5005
R16135 DVSS.n16637 DVSS.n16301 4.5005
R16136 DVSS.n16301 DVSS.n16292 4.5005
R16137 DVSS.n16639 DVSS.n16301 4.5005
R16138 DVSS.n16308 DVSS.n16295 4.5005
R16139 DVSS.n16319 DVSS.n16295 4.5005
R16140 DVSS.n16307 DVSS.n16295 4.5005
R16141 DVSS.n16634 DVSS.n16295 4.5005
R16142 DVSS.n16306 DVSS.n16295 4.5005
R16143 DVSS.n16637 DVSS.n16295 4.5005
R16144 DVSS.n16295 DVSS.n16292 4.5005
R16145 DVSS.n16639 DVSS.n16295 4.5005
R16146 DVSS.n16312 DVSS.n16302 4.5005
R16147 DVSS.n16314 DVSS.n16302 4.5005
R16148 DVSS.n16311 DVSS.n16302 4.5005
R16149 DVSS.n16315 DVSS.n16302 4.5005
R16150 DVSS.n16310 DVSS.n16302 4.5005
R16151 DVSS.n16317 DVSS.n16302 4.5005
R16152 DVSS.n16309 DVSS.n16302 4.5005
R16153 DVSS.n16318 DVSS.n16302 4.5005
R16154 DVSS.n16308 DVSS.n16302 4.5005
R16155 DVSS.n16319 DVSS.n16302 4.5005
R16156 DVSS.n16307 DVSS.n16302 4.5005
R16157 DVSS.n16634 DVSS.n16302 4.5005
R16158 DVSS.n16306 DVSS.n16302 4.5005
R16159 DVSS.n16637 DVSS.n16302 4.5005
R16160 DVSS.n16302 DVSS.n16292 4.5005
R16161 DVSS.n16639 DVSS.n16302 4.5005
R16162 DVSS.n16312 DVSS.n16294 4.5005
R16163 DVSS.n16314 DVSS.n16294 4.5005
R16164 DVSS.n16311 DVSS.n16294 4.5005
R16165 DVSS.n16315 DVSS.n16294 4.5005
R16166 DVSS.n16310 DVSS.n16294 4.5005
R16167 DVSS.n16317 DVSS.n16294 4.5005
R16168 DVSS.n16309 DVSS.n16294 4.5005
R16169 DVSS.n16318 DVSS.n16294 4.5005
R16170 DVSS.n16308 DVSS.n16294 4.5005
R16171 DVSS.n16319 DVSS.n16294 4.5005
R16172 DVSS.n16307 DVSS.n16294 4.5005
R16173 DVSS.n16634 DVSS.n16294 4.5005
R16174 DVSS.n16306 DVSS.n16294 4.5005
R16175 DVSS.n16637 DVSS.n16294 4.5005
R16176 DVSS.n16294 DVSS.n16292 4.5005
R16177 DVSS.n16639 DVSS.n16294 4.5005
R16178 DVSS.n16312 DVSS.n16303 4.5005
R16179 DVSS.n16314 DVSS.n16303 4.5005
R16180 DVSS.n16311 DVSS.n16303 4.5005
R16181 DVSS.n16315 DVSS.n16303 4.5005
R16182 DVSS.n16310 DVSS.n16303 4.5005
R16183 DVSS.n16317 DVSS.n16303 4.5005
R16184 DVSS.n16309 DVSS.n16303 4.5005
R16185 DVSS.n16318 DVSS.n16303 4.5005
R16186 DVSS.n16308 DVSS.n16303 4.5005
R16187 DVSS.n16319 DVSS.n16303 4.5005
R16188 DVSS.n16307 DVSS.n16303 4.5005
R16189 DVSS.n16634 DVSS.n16303 4.5005
R16190 DVSS.n16306 DVSS.n16303 4.5005
R16191 DVSS.n16637 DVSS.n16303 4.5005
R16192 DVSS.n16303 DVSS.n16292 4.5005
R16193 DVSS.n16639 DVSS.n16303 4.5005
R16194 DVSS.n16312 DVSS.n16293 4.5005
R16195 DVSS.n16314 DVSS.n16293 4.5005
R16196 DVSS.n16311 DVSS.n16293 4.5005
R16197 DVSS.n16315 DVSS.n16293 4.5005
R16198 DVSS.n16310 DVSS.n16293 4.5005
R16199 DVSS.n16317 DVSS.n16293 4.5005
R16200 DVSS.n16309 DVSS.n16293 4.5005
R16201 DVSS.n16318 DVSS.n16293 4.5005
R16202 DVSS.n16308 DVSS.n16293 4.5005
R16203 DVSS.n16319 DVSS.n16293 4.5005
R16204 DVSS.n16307 DVSS.n16293 4.5005
R16205 DVSS.n16634 DVSS.n16293 4.5005
R16206 DVSS.n16306 DVSS.n16293 4.5005
R16207 DVSS.n16637 DVSS.n16293 4.5005
R16208 DVSS.n16293 DVSS.n16292 4.5005
R16209 DVSS.n16639 DVSS.n16293 4.5005
R16210 DVSS.n16638 DVSS.n16312 4.5005
R16211 DVSS.n16638 DVSS.n16314 4.5005
R16212 DVSS.n16638 DVSS.n16311 4.5005
R16213 DVSS.n16638 DVSS.n16315 4.5005
R16214 DVSS.n16638 DVSS.n16310 4.5005
R16215 DVSS.n16638 DVSS.n16317 4.5005
R16216 DVSS.n16638 DVSS.n16309 4.5005
R16217 DVSS.n16638 DVSS.n16318 4.5005
R16218 DVSS.n16638 DVSS.n16308 4.5005
R16219 DVSS.n16638 DVSS.n16319 4.5005
R16220 DVSS.n16638 DVSS.n16307 4.5005
R16221 DVSS.n16638 DVSS.n16634 4.5005
R16222 DVSS.n16638 DVSS.n16306 4.5005
R16223 DVSS.n16638 DVSS.n16637 4.5005
R16224 DVSS.n16638 DVSS.n16292 4.5005
R16225 DVSS.n16639 DVSS.n16638 4.5005
R16226 DVSS.n15856 DVSS.n15841 4.5005
R16227 DVSS.n15858 DVSS.n15841 4.5005
R16228 DVSS.n15855 DVSS.n15841 4.5005
R16229 DVSS.n15859 DVSS.n15841 4.5005
R16230 DVSS.n15854 DVSS.n15841 4.5005
R16231 DVSS.n15862 DVSS.n15841 4.5005
R16232 DVSS.n15852 DVSS.n15841 4.5005
R16233 DVSS.n15863 DVSS.n15841 4.5005
R16234 DVSS.n15851 DVSS.n15841 4.5005
R16235 DVSS.n17860 DVSS.n15841 4.5005
R16236 DVSS.n15850 DVSS.n15841 4.5005
R16237 DVSS.n17865 DVSS.n15841 4.5005
R16238 DVSS.n15856 DVSS.n15842 4.5005
R16239 DVSS.n15858 DVSS.n15842 4.5005
R16240 DVSS.n15855 DVSS.n15842 4.5005
R16241 DVSS.n15859 DVSS.n15842 4.5005
R16242 DVSS.n15854 DVSS.n15842 4.5005
R16243 DVSS.n15861 DVSS.n15842 4.5005
R16244 DVSS.n15853 DVSS.n15842 4.5005
R16245 DVSS.n15862 DVSS.n15842 4.5005
R16246 DVSS.n15852 DVSS.n15842 4.5005
R16247 DVSS.n15863 DVSS.n15842 4.5005
R16248 DVSS.n15851 DVSS.n15842 4.5005
R16249 DVSS.n17860 DVSS.n15842 4.5005
R16250 DVSS.n15850 DVSS.n15842 4.5005
R16251 DVSS.n17863 DVSS.n15842 4.5005
R16252 DVSS.n15842 DVSS.n15836 4.5005
R16253 DVSS.n17865 DVSS.n15842 4.5005
R16254 DVSS.n15856 DVSS.n15840 4.5005
R16255 DVSS.n15858 DVSS.n15840 4.5005
R16256 DVSS.n15855 DVSS.n15840 4.5005
R16257 DVSS.n15859 DVSS.n15840 4.5005
R16258 DVSS.n15854 DVSS.n15840 4.5005
R16259 DVSS.n15861 DVSS.n15840 4.5005
R16260 DVSS.n15853 DVSS.n15840 4.5005
R16261 DVSS.n15862 DVSS.n15840 4.5005
R16262 DVSS.n15852 DVSS.n15840 4.5005
R16263 DVSS.n15863 DVSS.n15840 4.5005
R16264 DVSS.n15851 DVSS.n15840 4.5005
R16265 DVSS.n17860 DVSS.n15840 4.5005
R16266 DVSS.n15850 DVSS.n15840 4.5005
R16267 DVSS.n17863 DVSS.n15840 4.5005
R16268 DVSS.n15840 DVSS.n15836 4.5005
R16269 DVSS.n17865 DVSS.n15840 4.5005
R16270 DVSS.n15856 DVSS.n15843 4.5005
R16271 DVSS.n15858 DVSS.n15843 4.5005
R16272 DVSS.n15855 DVSS.n15843 4.5005
R16273 DVSS.n15859 DVSS.n15843 4.5005
R16274 DVSS.n15854 DVSS.n15843 4.5005
R16275 DVSS.n15861 DVSS.n15843 4.5005
R16276 DVSS.n15853 DVSS.n15843 4.5005
R16277 DVSS.n15862 DVSS.n15843 4.5005
R16278 DVSS.n15852 DVSS.n15843 4.5005
R16279 DVSS.n15863 DVSS.n15843 4.5005
R16280 DVSS.n15851 DVSS.n15843 4.5005
R16281 DVSS.n17860 DVSS.n15843 4.5005
R16282 DVSS.n15850 DVSS.n15843 4.5005
R16283 DVSS.n17863 DVSS.n15843 4.5005
R16284 DVSS.n15843 DVSS.n15836 4.5005
R16285 DVSS.n17865 DVSS.n15843 4.5005
R16286 DVSS.n15856 DVSS.n15839 4.5005
R16287 DVSS.n15858 DVSS.n15839 4.5005
R16288 DVSS.n15855 DVSS.n15839 4.5005
R16289 DVSS.n15859 DVSS.n15839 4.5005
R16290 DVSS.n15854 DVSS.n15839 4.5005
R16291 DVSS.n15861 DVSS.n15839 4.5005
R16292 DVSS.n15853 DVSS.n15839 4.5005
R16293 DVSS.n15862 DVSS.n15839 4.5005
R16294 DVSS.n15852 DVSS.n15839 4.5005
R16295 DVSS.n15863 DVSS.n15839 4.5005
R16296 DVSS.n15851 DVSS.n15839 4.5005
R16297 DVSS.n17860 DVSS.n15839 4.5005
R16298 DVSS.n15850 DVSS.n15839 4.5005
R16299 DVSS.n17863 DVSS.n15839 4.5005
R16300 DVSS.n15839 DVSS.n15836 4.5005
R16301 DVSS.n17865 DVSS.n15839 4.5005
R16302 DVSS.n15856 DVSS.n15845 4.5005
R16303 DVSS.n15858 DVSS.n15845 4.5005
R16304 DVSS.n15855 DVSS.n15845 4.5005
R16305 DVSS.n15859 DVSS.n15845 4.5005
R16306 DVSS.n15854 DVSS.n15845 4.5005
R16307 DVSS.n15861 DVSS.n15845 4.5005
R16308 DVSS.n15853 DVSS.n15845 4.5005
R16309 DVSS.n15862 DVSS.n15845 4.5005
R16310 DVSS.n15852 DVSS.n15845 4.5005
R16311 DVSS.n15863 DVSS.n15845 4.5005
R16312 DVSS.n15851 DVSS.n15845 4.5005
R16313 DVSS.n17860 DVSS.n15845 4.5005
R16314 DVSS.n15850 DVSS.n15845 4.5005
R16315 DVSS.n17863 DVSS.n15845 4.5005
R16316 DVSS.n17865 DVSS.n15845 4.5005
R16317 DVSS.n15856 DVSS.n15838 4.5005
R16318 DVSS.n15858 DVSS.n15838 4.5005
R16319 DVSS.n15855 DVSS.n15838 4.5005
R16320 DVSS.n15859 DVSS.n15838 4.5005
R16321 DVSS.n15854 DVSS.n15838 4.5005
R16322 DVSS.n15861 DVSS.n15838 4.5005
R16323 DVSS.n15853 DVSS.n15838 4.5005
R16324 DVSS.n15862 DVSS.n15838 4.5005
R16325 DVSS.n15852 DVSS.n15838 4.5005
R16326 DVSS.n15863 DVSS.n15838 4.5005
R16327 DVSS.n15851 DVSS.n15838 4.5005
R16328 DVSS.n17860 DVSS.n15838 4.5005
R16329 DVSS.n17863 DVSS.n15838 4.5005
R16330 DVSS.n17865 DVSS.n15838 4.5005
R16331 DVSS.n15856 DVSS.n15847 4.5005
R16332 DVSS.n15858 DVSS.n15847 4.5005
R16333 DVSS.n15855 DVSS.n15847 4.5005
R16334 DVSS.n15859 DVSS.n15847 4.5005
R16335 DVSS.n15854 DVSS.n15847 4.5005
R16336 DVSS.n15861 DVSS.n15847 4.5005
R16337 DVSS.n15853 DVSS.n15847 4.5005
R16338 DVSS.n15862 DVSS.n15847 4.5005
R16339 DVSS.n15852 DVSS.n15847 4.5005
R16340 DVSS.n15863 DVSS.n15847 4.5005
R16341 DVSS.n15851 DVSS.n15847 4.5005
R16342 DVSS.n17860 DVSS.n15847 4.5005
R16343 DVSS.n17863 DVSS.n15847 4.5005
R16344 DVSS.n17865 DVSS.n15847 4.5005
R16345 DVSS.n15856 DVSS.n15837 4.5005
R16346 DVSS.n15858 DVSS.n15837 4.5005
R16347 DVSS.n15855 DVSS.n15837 4.5005
R16348 DVSS.n15859 DVSS.n15837 4.5005
R16349 DVSS.n15854 DVSS.n15837 4.5005
R16350 DVSS.n15861 DVSS.n15837 4.5005
R16351 DVSS.n15853 DVSS.n15837 4.5005
R16352 DVSS.n15862 DVSS.n15837 4.5005
R16353 DVSS.n15852 DVSS.n15837 4.5005
R16354 DVSS.n15863 DVSS.n15837 4.5005
R16355 DVSS.n15851 DVSS.n15837 4.5005
R16356 DVSS.n17860 DVSS.n15837 4.5005
R16357 DVSS.n15850 DVSS.n15837 4.5005
R16358 DVSS.n17863 DVSS.n15837 4.5005
R16359 DVSS.n17865 DVSS.n15837 4.5005
R16360 DVSS.n17864 DVSS.n15856 4.5005
R16361 DVSS.n17864 DVSS.n15858 4.5005
R16362 DVSS.n17864 DVSS.n15855 4.5005
R16363 DVSS.n17864 DVSS.n15859 4.5005
R16364 DVSS.n17864 DVSS.n15854 4.5005
R16365 DVSS.n17864 DVSS.n15861 4.5005
R16366 DVSS.n17864 DVSS.n15853 4.5005
R16367 DVSS.n17864 DVSS.n15862 4.5005
R16368 DVSS.n17864 DVSS.n15852 4.5005
R16369 DVSS.n17864 DVSS.n15863 4.5005
R16370 DVSS.n17864 DVSS.n15851 4.5005
R16371 DVSS.n17864 DVSS.n17860 4.5005
R16372 DVSS.n17864 DVSS.n15850 4.5005
R16373 DVSS.n17864 DVSS.n17863 4.5005
R16374 DVSS.n17864 DVSS.n15836 4.5005
R16375 DVSS.n17865 DVSS.n17864 4.5005
R16376 DVSS.n16318 DVSS.n16295 4.5005
R16377 DVSS.n16309 DVSS.n16295 4.5005
R16378 DVSS.n16317 DVSS.n16295 4.5005
R16379 DVSS.n16310 DVSS.n16295 4.5005
R16380 DVSS.n16315 DVSS.n16295 4.5005
R16381 DVSS.n16311 DVSS.n16295 4.5005
R16382 DVSS.n16314 DVSS.n16295 4.5005
R16383 DVSS.n16312 DVSS.n16295 4.5005
R16384 DVSS.n16318 DVSS.n16301 4.5005
R16385 DVSS.n16309 DVSS.n16301 4.5005
R16386 DVSS.n16317 DVSS.n16301 4.5005
R16387 DVSS.n16310 DVSS.n16301 4.5005
R16388 DVSS.n16315 DVSS.n16301 4.5005
R16389 DVSS.n16311 DVSS.n16301 4.5005
R16390 DVSS.n16314 DVSS.n16301 4.5005
R16391 DVSS.n16312 DVSS.n16301 4.5005
R16392 DVSS.n16318 DVSS.n16296 4.5005
R16393 DVSS.n16309 DVSS.n16296 4.5005
R16394 DVSS.n16317 DVSS.n16296 4.5005
R16395 DVSS.n16310 DVSS.n16296 4.5005
R16396 DVSS.n16315 DVSS.n16296 4.5005
R16397 DVSS.n16311 DVSS.n16296 4.5005
R16398 DVSS.n16314 DVSS.n16296 4.5005
R16399 DVSS.n16312 DVSS.n16296 4.5005
R16400 DVSS.n15994 DVSS.n15993 4.5005
R16401 DVSS.n17655 DVSS.n15994 4.5005
R16402 DVSS.n16020 DVSS.n15994 4.5005
R16403 DVSS.n16022 DVSS.n15994 4.5005
R16404 DVSS.n16019 DVSS.n15994 4.5005
R16405 DVSS.n16024 DVSS.n15994 4.5005
R16406 DVSS.n16018 DVSS.n15994 4.5005
R16407 DVSS.n16025 DVSS.n15994 4.5005
R16408 DVSS.n16017 DVSS.n15994 4.5005
R16409 DVSS.n16026 DVSS.n15994 4.5005
R16410 DVSS.n16016 DVSS.n15994 4.5005
R16411 DVSS.n16027 DVSS.n15994 4.5005
R16412 DVSS.n16029 DVSS.n15994 4.5005
R16413 DVSS.n16010 DVSS.n15994 4.5005
R16414 DVSS.n17653 DVSS.n15994 4.5005
R16415 DVSS.n17654 DVSS.n15993 4.5005
R16416 DVSS.n17655 DVSS.n17654 4.5005
R16417 DVSS.n17654 DVSS.n16020 4.5005
R16418 DVSS.n17654 DVSS.n16022 4.5005
R16419 DVSS.n17654 DVSS.n16019 4.5005
R16420 DVSS.n17654 DVSS.n16024 4.5005
R16421 DVSS.n17654 DVSS.n16018 4.5005
R16422 DVSS.n17654 DVSS.n16025 4.5005
R16423 DVSS.n17654 DVSS.n16017 4.5005
R16424 DVSS.n17654 DVSS.n16026 4.5005
R16425 DVSS.n17654 DVSS.n16016 4.5005
R16426 DVSS.n17654 DVSS.n16027 4.5005
R16427 DVSS.n17654 DVSS.n16015 4.5005
R16428 DVSS.n17654 DVSS.n16029 4.5005
R16429 DVSS.n17654 DVSS.n16010 4.5005
R16430 DVSS.n17654 DVSS.n17653 4.5005
R16431 DVSS.n15266 DVSS.n15246 4.5005
R16432 DVSS.n15266 DVSS.n15247 4.5005
R16433 DVSS.n15266 DVSS.n15245 4.5005
R16434 DVSS.n15266 DVSS.n15248 4.5005
R16435 DVSS.n15266 DVSS.n15244 4.5005
R16436 DVSS.n18378 DVSS.n15266 4.5005
R16437 DVSS.n15272 DVSS.n15266 4.5005
R16438 DVSS.n15266 DVSS.n15249 4.5005
R16439 DVSS.n15266 DVSS.n15242 4.5005
R16440 DVSS.n15266 DVSS.n15250 4.5005
R16441 DVSS.n15266 DVSS.n15241 4.5005
R16442 DVSS.n15266 DVSS.n15251 4.5005
R16443 DVSS.n15266 DVSS.n15240 4.5005
R16444 DVSS.n15266 DVSS.n15252 4.5005
R16445 DVSS.n15271 DVSS.n15266 4.5005
R16446 DVSS.n18380 DVSS.n15266 4.5005
R16447 DVSS.n15254 DVSS.n15246 4.5005
R16448 DVSS.n15254 DVSS.n15247 4.5005
R16449 DVSS.n15254 DVSS.n15245 4.5005
R16450 DVSS.n15254 DVSS.n15248 4.5005
R16451 DVSS.n15254 DVSS.n15244 4.5005
R16452 DVSS.n18378 DVSS.n15254 4.5005
R16453 DVSS.n15272 DVSS.n15254 4.5005
R16454 DVSS.n15254 DVSS.n15249 4.5005
R16455 DVSS.n15254 DVSS.n15242 4.5005
R16456 DVSS.n15254 DVSS.n15250 4.5005
R16457 DVSS.n15254 DVSS.n15241 4.5005
R16458 DVSS.n15254 DVSS.n15251 4.5005
R16459 DVSS.n15254 DVSS.n15252 4.5005
R16460 DVSS.n15271 DVSS.n15254 4.5005
R16461 DVSS.n18380 DVSS.n15254 4.5005
R16462 DVSS.n18379 DVSS.n15246 4.5005
R16463 DVSS.n18379 DVSS.n15247 4.5005
R16464 DVSS.n18379 DVSS.n15245 4.5005
R16465 DVSS.n18379 DVSS.n15248 4.5005
R16466 DVSS.n18379 DVSS.n15244 4.5005
R16467 DVSS.n18379 DVSS.n18378 4.5005
R16468 DVSS.n18379 DVSS.n15272 4.5005
R16469 DVSS.n18379 DVSS.n15249 4.5005
R16470 DVSS.n18379 DVSS.n15242 4.5005
R16471 DVSS.n18379 DVSS.n15250 4.5005
R16472 DVSS.n18379 DVSS.n15241 4.5005
R16473 DVSS.n18379 DVSS.n15251 4.5005
R16474 DVSS.n18379 DVSS.n15240 4.5005
R16475 DVSS.n18379 DVSS.n15252 4.5005
R16476 DVSS.n18379 DVSS.n15271 4.5005
R16477 DVSS.n18380 DVSS.n18379 4.5005
R16478 DVSS.n13595 DVSS.n13580 4.5005
R16479 DVSS.n13592 DVSS.n13580 4.5005
R16480 DVSS.n13594 DVSS.n13580 4.5005
R16481 DVSS.n13593 DVSS.n13580 4.5005
R16482 DVSS.n13595 DVSS.n13572 4.5005
R16483 DVSS.n13592 DVSS.n13572 4.5005
R16484 DVSS.n13594 DVSS.n13572 4.5005
R16485 DVSS.n13593 DVSS.n13572 4.5005
R16486 DVSS.n13595 DVSS.n13579 4.5005
R16487 DVSS.n13592 DVSS.n13579 4.5005
R16488 DVSS.n13594 DVSS.n13579 4.5005
R16489 DVSS.n13593 DVSS.n13579 4.5005
R16490 DVSS.n13595 DVSS.n13573 4.5005
R16491 DVSS.n13592 DVSS.n13573 4.5005
R16492 DVSS.n13594 DVSS.n13573 4.5005
R16493 DVSS.n13593 DVSS.n13573 4.5005
R16494 DVSS.n13595 DVSS.n13578 4.5005
R16495 DVSS.n13592 DVSS.n13578 4.5005
R16496 DVSS.n13594 DVSS.n13578 4.5005
R16497 DVSS.n13593 DVSS.n13578 4.5005
R16498 DVSS.n13595 DVSS.n13574 4.5005
R16499 DVSS.n13592 DVSS.n13574 4.5005
R16500 DVSS.n13594 DVSS.n13574 4.5005
R16501 DVSS.n13593 DVSS.n13574 4.5005
R16502 DVSS.n13595 DVSS.n13577 4.5005
R16503 DVSS.n13592 DVSS.n13577 4.5005
R16504 DVSS.n13594 DVSS.n13577 4.5005
R16505 DVSS.n13593 DVSS.n13577 4.5005
R16506 DVSS.n13595 DVSS.n13575 4.5005
R16507 DVSS.n13592 DVSS.n13575 4.5005
R16508 DVSS.n13594 DVSS.n13575 4.5005
R16509 DVSS.n13593 DVSS.n13575 4.5005
R16510 DVSS.n13595 DVSS.n13576 4.5005
R16511 DVSS.n13592 DVSS.n13576 4.5005
R16512 DVSS.n13594 DVSS.n13576 4.5005
R16513 DVSS.n13593 DVSS.n13576 4.5005
R16514 DVSS.n19592 DVSS.n19591 4.5005
R16515 DVSS.n19593 DVSS.n19592 4.5005
R16516 DVSS.n19089 DVSS.n19088 4.5005
R16517 DVSS.n19849 DVSS.n19089 4.5005
R16518 DVSS.n19513 DVSS.n19512 4.5005
R16519 DVSS.n19512 DVSS.n19504 4.5005
R16520 DVSS.n19502 DVSS.n19065 4.5005
R16521 DVSS.n19593 DVSS.n19065 4.5005
R16522 DVSS.n19850 DVSS.n19078 4.5005
R16523 DVSS.n19850 DVSS.n19849 4.5005
R16524 DVSS.n16549 DVSS.n16548 4.5005
R16525 DVSS.n16548 DVSS.n16472 4.5005
R16526 DVSS.n16550 DVSS.n16472 4.5005
R16527 DVSS.n16550 DVSS.n16473 4.5005
R16528 DVSS.n16550 DVSS.n16358 4.5005
R16529 DVSS.n16550 DVSS.n16474 4.5005
R16530 DVSS.n16550 DVSS.n16357 4.5005
R16531 DVSS.n16550 DVSS.n16475 4.5005
R16532 DVSS.n16550 DVSS.n16356 4.5005
R16533 DVSS.n16550 DVSS.n16476 4.5005
R16534 DVSS.n16550 DVSS.n16355 4.5005
R16535 DVSS.n16550 DVSS.n16477 4.5005
R16536 DVSS.n16550 DVSS.n16354 4.5005
R16537 DVSS.n16550 DVSS.n16549 4.5005
R16538 DVSS.n13642 DVSS.n13624 4.5005
R16539 DVSS.n13640 DVSS.n13624 4.5005
R16540 DVSS.n13645 DVSS.n13624 4.5005
R16541 DVSS.n13639 DVSS.n13624 4.5005
R16542 DVSS.n13646 DVSS.n13624 4.5005
R16543 DVSS.n13638 DVSS.n13624 4.5005
R16544 DVSS.n13647 DVSS.n13624 4.5005
R16545 DVSS.n21205 DVSS.n13624 4.5005
R16546 DVSS.n21213 DVSS.n13624 4.5005
R16547 DVSS.n21215 DVSS.n13624 4.5005
R16548 DVSS.n13642 DVSS.n13623 4.5005
R16549 DVSS.n13641 DVSS.n13623 4.5005
R16550 DVSS.n13644 DVSS.n13623 4.5005
R16551 DVSS.n13640 DVSS.n13623 4.5005
R16552 DVSS.n13645 DVSS.n13623 4.5005
R16553 DVSS.n13639 DVSS.n13623 4.5005
R16554 DVSS.n13646 DVSS.n13623 4.5005
R16555 DVSS.n13638 DVSS.n13623 4.5005
R16556 DVSS.n13647 DVSS.n13623 4.5005
R16557 DVSS.n13637 DVSS.n13623 4.5005
R16558 DVSS.n13649 DVSS.n13623 4.5005
R16559 DVSS.n21213 DVSS.n13623 4.5005
R16560 DVSS.n21215 DVSS.n13623 4.5005
R16561 DVSS.n13642 DVSS.n13625 4.5005
R16562 DVSS.n13641 DVSS.n13625 4.5005
R16563 DVSS.n13644 DVSS.n13625 4.5005
R16564 DVSS.n13640 DVSS.n13625 4.5005
R16565 DVSS.n13645 DVSS.n13625 4.5005
R16566 DVSS.n13639 DVSS.n13625 4.5005
R16567 DVSS.n13646 DVSS.n13625 4.5005
R16568 DVSS.n13638 DVSS.n13625 4.5005
R16569 DVSS.n13647 DVSS.n13625 4.5005
R16570 DVSS.n13637 DVSS.n13625 4.5005
R16571 DVSS.n13649 DVSS.n13625 4.5005
R16572 DVSS.n21213 DVSS.n13625 4.5005
R16573 DVSS.n21215 DVSS.n13625 4.5005
R16574 DVSS.n13642 DVSS.n13622 4.5005
R16575 DVSS.n13641 DVSS.n13622 4.5005
R16576 DVSS.n13644 DVSS.n13622 4.5005
R16577 DVSS.n13640 DVSS.n13622 4.5005
R16578 DVSS.n13645 DVSS.n13622 4.5005
R16579 DVSS.n13639 DVSS.n13622 4.5005
R16580 DVSS.n13646 DVSS.n13622 4.5005
R16581 DVSS.n13638 DVSS.n13622 4.5005
R16582 DVSS.n13647 DVSS.n13622 4.5005
R16583 DVSS.n13637 DVSS.n13622 4.5005
R16584 DVSS.n13649 DVSS.n13622 4.5005
R16585 DVSS.n21213 DVSS.n13622 4.5005
R16586 DVSS.n21215 DVSS.n13622 4.5005
R16587 DVSS.n13642 DVSS.n13626 4.5005
R16588 DVSS.n13641 DVSS.n13626 4.5005
R16589 DVSS.n13644 DVSS.n13626 4.5005
R16590 DVSS.n13640 DVSS.n13626 4.5005
R16591 DVSS.n13645 DVSS.n13626 4.5005
R16592 DVSS.n13639 DVSS.n13626 4.5005
R16593 DVSS.n13646 DVSS.n13626 4.5005
R16594 DVSS.n13638 DVSS.n13626 4.5005
R16595 DVSS.n13647 DVSS.n13626 4.5005
R16596 DVSS.n13637 DVSS.n13626 4.5005
R16597 DVSS.n13649 DVSS.n13626 4.5005
R16598 DVSS.n21213 DVSS.n13626 4.5005
R16599 DVSS.n21215 DVSS.n13626 4.5005
R16600 DVSS.n13642 DVSS.n13621 4.5005
R16601 DVSS.n13641 DVSS.n13621 4.5005
R16602 DVSS.n13644 DVSS.n13621 4.5005
R16603 DVSS.n13640 DVSS.n13621 4.5005
R16604 DVSS.n13645 DVSS.n13621 4.5005
R16605 DVSS.n13639 DVSS.n13621 4.5005
R16606 DVSS.n13646 DVSS.n13621 4.5005
R16607 DVSS.n13638 DVSS.n13621 4.5005
R16608 DVSS.n13647 DVSS.n13621 4.5005
R16609 DVSS.n13637 DVSS.n13621 4.5005
R16610 DVSS.n13649 DVSS.n13621 4.5005
R16611 DVSS.n21213 DVSS.n13621 4.5005
R16612 DVSS.n21215 DVSS.n13621 4.5005
R16613 DVSS.n13642 DVSS.n13627 4.5005
R16614 DVSS.n13641 DVSS.n13627 4.5005
R16615 DVSS.n13644 DVSS.n13627 4.5005
R16616 DVSS.n13640 DVSS.n13627 4.5005
R16617 DVSS.n13645 DVSS.n13627 4.5005
R16618 DVSS.n13639 DVSS.n13627 4.5005
R16619 DVSS.n13646 DVSS.n13627 4.5005
R16620 DVSS.n13638 DVSS.n13627 4.5005
R16621 DVSS.n13647 DVSS.n13627 4.5005
R16622 DVSS.n13637 DVSS.n13627 4.5005
R16623 DVSS.n13649 DVSS.n13627 4.5005
R16624 DVSS.n21213 DVSS.n13627 4.5005
R16625 DVSS.n21215 DVSS.n13627 4.5005
R16626 DVSS.n13642 DVSS.n13620 4.5005
R16627 DVSS.n13641 DVSS.n13620 4.5005
R16628 DVSS.n13644 DVSS.n13620 4.5005
R16629 DVSS.n13640 DVSS.n13620 4.5005
R16630 DVSS.n13645 DVSS.n13620 4.5005
R16631 DVSS.n13639 DVSS.n13620 4.5005
R16632 DVSS.n13646 DVSS.n13620 4.5005
R16633 DVSS.n13638 DVSS.n13620 4.5005
R16634 DVSS.n13647 DVSS.n13620 4.5005
R16635 DVSS.n13637 DVSS.n13620 4.5005
R16636 DVSS.n13649 DVSS.n13620 4.5005
R16637 DVSS.n21213 DVSS.n13620 4.5005
R16638 DVSS.n21215 DVSS.n13620 4.5005
R16639 DVSS.n13642 DVSS.n13628 4.5005
R16640 DVSS.n13641 DVSS.n13628 4.5005
R16641 DVSS.n13644 DVSS.n13628 4.5005
R16642 DVSS.n13640 DVSS.n13628 4.5005
R16643 DVSS.n13645 DVSS.n13628 4.5005
R16644 DVSS.n13639 DVSS.n13628 4.5005
R16645 DVSS.n13646 DVSS.n13628 4.5005
R16646 DVSS.n13638 DVSS.n13628 4.5005
R16647 DVSS.n13647 DVSS.n13628 4.5005
R16648 DVSS.n13637 DVSS.n13628 4.5005
R16649 DVSS.n13649 DVSS.n13628 4.5005
R16650 DVSS.n21213 DVSS.n13628 4.5005
R16651 DVSS.n21215 DVSS.n13628 4.5005
R16652 DVSS.n13642 DVSS.n13619 4.5005
R16653 DVSS.n13641 DVSS.n13619 4.5005
R16654 DVSS.n13644 DVSS.n13619 4.5005
R16655 DVSS.n13640 DVSS.n13619 4.5005
R16656 DVSS.n13645 DVSS.n13619 4.5005
R16657 DVSS.n13639 DVSS.n13619 4.5005
R16658 DVSS.n13646 DVSS.n13619 4.5005
R16659 DVSS.n13638 DVSS.n13619 4.5005
R16660 DVSS.n13647 DVSS.n13619 4.5005
R16661 DVSS.n13637 DVSS.n13619 4.5005
R16662 DVSS.n13649 DVSS.n13619 4.5005
R16663 DVSS.n21213 DVSS.n13619 4.5005
R16664 DVSS.n21215 DVSS.n13619 4.5005
R16665 DVSS.n21214 DVSS.n13642 4.5005
R16666 DVSS.n21214 DVSS.n13641 4.5005
R16667 DVSS.n21214 DVSS.n13644 4.5005
R16668 DVSS.n21214 DVSS.n13640 4.5005
R16669 DVSS.n21214 DVSS.n13645 4.5005
R16670 DVSS.n21214 DVSS.n13639 4.5005
R16671 DVSS.n21214 DVSS.n13646 4.5005
R16672 DVSS.n21214 DVSS.n13638 4.5005
R16673 DVSS.n21214 DVSS.n13647 4.5005
R16674 DVSS.n21214 DVSS.n13637 4.5005
R16675 DVSS.n21214 DVSS.n13649 4.5005
R16676 DVSS.n21214 DVSS.n21213 4.5005
R16677 DVSS.n21214 DVSS.n13635 4.5005
R16678 DVSS.n21215 DVSS.n21214 4.5005
R16679 DVSS.n13736 DVSS.n13629 4.5005
R16680 DVSS.n13734 DVSS.n13629 4.5005
R16681 DVSS.n13739 DVSS.n13629 4.5005
R16682 DVSS.n13733 DVSS.n13629 4.5005
R16683 DVSS.n13740 DVSS.n13629 4.5005
R16684 DVSS.n13732 DVSS.n13629 4.5005
R16685 DVSS.n13741 DVSS.n13629 4.5005
R16686 DVSS.n13730 DVSS.n13629 4.5005
R16687 DVSS.n13744 DVSS.n13629 4.5005
R16688 DVSS.n21142 DVSS.n13629 4.5005
R16689 DVSS.n13759 DVSS.n13736 4.5005
R16690 DVSS.n13759 DVSS.n13735 4.5005
R16691 DVSS.n13759 DVSS.n13738 4.5005
R16692 DVSS.n13759 DVSS.n13734 4.5005
R16693 DVSS.n13759 DVSS.n13739 4.5005
R16694 DVSS.n13759 DVSS.n13733 4.5005
R16695 DVSS.n13759 DVSS.n13740 4.5005
R16696 DVSS.n13759 DVSS.n13732 4.5005
R16697 DVSS.n13759 DVSS.n13741 4.5005
R16698 DVSS.n13759 DVSS.n13731 4.5005
R16699 DVSS.n13759 DVSS.n13743 4.5005
R16700 DVSS.n13759 DVSS.n13744 4.5005
R16701 DVSS.n21142 DVSS.n13759 4.5005
R16702 DVSS.n13756 DVSS.n13736 4.5005
R16703 DVSS.n13756 DVSS.n13735 4.5005
R16704 DVSS.n13756 DVSS.n13738 4.5005
R16705 DVSS.n13756 DVSS.n13734 4.5005
R16706 DVSS.n13756 DVSS.n13739 4.5005
R16707 DVSS.n13756 DVSS.n13733 4.5005
R16708 DVSS.n13756 DVSS.n13740 4.5005
R16709 DVSS.n13756 DVSS.n13732 4.5005
R16710 DVSS.n13756 DVSS.n13741 4.5005
R16711 DVSS.n13756 DVSS.n13731 4.5005
R16712 DVSS.n13756 DVSS.n13743 4.5005
R16713 DVSS.n13756 DVSS.n13744 4.5005
R16714 DVSS.n21142 DVSS.n13756 4.5005
R16715 DVSS.n13761 DVSS.n13736 4.5005
R16716 DVSS.n13761 DVSS.n13735 4.5005
R16717 DVSS.n13761 DVSS.n13738 4.5005
R16718 DVSS.n13761 DVSS.n13734 4.5005
R16719 DVSS.n13761 DVSS.n13739 4.5005
R16720 DVSS.n13761 DVSS.n13733 4.5005
R16721 DVSS.n13761 DVSS.n13740 4.5005
R16722 DVSS.n13761 DVSS.n13732 4.5005
R16723 DVSS.n13761 DVSS.n13741 4.5005
R16724 DVSS.n13761 DVSS.n13731 4.5005
R16725 DVSS.n13761 DVSS.n13743 4.5005
R16726 DVSS.n13761 DVSS.n13744 4.5005
R16727 DVSS.n21142 DVSS.n13761 4.5005
R16728 DVSS.n13755 DVSS.n13736 4.5005
R16729 DVSS.n13755 DVSS.n13735 4.5005
R16730 DVSS.n13755 DVSS.n13738 4.5005
R16731 DVSS.n13755 DVSS.n13734 4.5005
R16732 DVSS.n13755 DVSS.n13739 4.5005
R16733 DVSS.n13755 DVSS.n13733 4.5005
R16734 DVSS.n13755 DVSS.n13740 4.5005
R16735 DVSS.n13755 DVSS.n13732 4.5005
R16736 DVSS.n13755 DVSS.n13741 4.5005
R16737 DVSS.n13755 DVSS.n13731 4.5005
R16738 DVSS.n13755 DVSS.n13743 4.5005
R16739 DVSS.n13755 DVSS.n13744 4.5005
R16740 DVSS.n21142 DVSS.n13755 4.5005
R16741 DVSS.n13763 DVSS.n13736 4.5005
R16742 DVSS.n13763 DVSS.n13735 4.5005
R16743 DVSS.n13763 DVSS.n13738 4.5005
R16744 DVSS.n13763 DVSS.n13734 4.5005
R16745 DVSS.n13763 DVSS.n13739 4.5005
R16746 DVSS.n13763 DVSS.n13733 4.5005
R16747 DVSS.n13763 DVSS.n13740 4.5005
R16748 DVSS.n13763 DVSS.n13732 4.5005
R16749 DVSS.n13763 DVSS.n13741 4.5005
R16750 DVSS.n13763 DVSS.n13731 4.5005
R16751 DVSS.n13763 DVSS.n13743 4.5005
R16752 DVSS.n13763 DVSS.n13744 4.5005
R16753 DVSS.n21142 DVSS.n13763 4.5005
R16754 DVSS.n13754 DVSS.n13736 4.5005
R16755 DVSS.n13754 DVSS.n13735 4.5005
R16756 DVSS.n13754 DVSS.n13738 4.5005
R16757 DVSS.n13754 DVSS.n13734 4.5005
R16758 DVSS.n13754 DVSS.n13739 4.5005
R16759 DVSS.n13754 DVSS.n13733 4.5005
R16760 DVSS.n13754 DVSS.n13740 4.5005
R16761 DVSS.n13754 DVSS.n13732 4.5005
R16762 DVSS.n13754 DVSS.n13741 4.5005
R16763 DVSS.n13754 DVSS.n13731 4.5005
R16764 DVSS.n13754 DVSS.n13743 4.5005
R16765 DVSS.n13754 DVSS.n13744 4.5005
R16766 DVSS.n21142 DVSS.n13754 4.5005
R16767 DVSS.n13765 DVSS.n13736 4.5005
R16768 DVSS.n13765 DVSS.n13735 4.5005
R16769 DVSS.n13765 DVSS.n13738 4.5005
R16770 DVSS.n13765 DVSS.n13734 4.5005
R16771 DVSS.n13765 DVSS.n13739 4.5005
R16772 DVSS.n13765 DVSS.n13733 4.5005
R16773 DVSS.n13765 DVSS.n13740 4.5005
R16774 DVSS.n13765 DVSS.n13732 4.5005
R16775 DVSS.n13765 DVSS.n13741 4.5005
R16776 DVSS.n13765 DVSS.n13731 4.5005
R16777 DVSS.n13765 DVSS.n13743 4.5005
R16778 DVSS.n13765 DVSS.n13744 4.5005
R16779 DVSS.n21142 DVSS.n13765 4.5005
R16780 DVSS.n13753 DVSS.n13736 4.5005
R16781 DVSS.n13753 DVSS.n13735 4.5005
R16782 DVSS.n13753 DVSS.n13738 4.5005
R16783 DVSS.n13753 DVSS.n13734 4.5005
R16784 DVSS.n13753 DVSS.n13739 4.5005
R16785 DVSS.n13753 DVSS.n13733 4.5005
R16786 DVSS.n13753 DVSS.n13740 4.5005
R16787 DVSS.n13753 DVSS.n13732 4.5005
R16788 DVSS.n13753 DVSS.n13741 4.5005
R16789 DVSS.n13753 DVSS.n13731 4.5005
R16790 DVSS.n13753 DVSS.n13743 4.5005
R16791 DVSS.n13753 DVSS.n13744 4.5005
R16792 DVSS.n21142 DVSS.n13753 4.5005
R16793 DVSS.n13767 DVSS.n13736 4.5005
R16794 DVSS.n13767 DVSS.n13735 4.5005
R16795 DVSS.n13767 DVSS.n13738 4.5005
R16796 DVSS.n13767 DVSS.n13734 4.5005
R16797 DVSS.n13767 DVSS.n13739 4.5005
R16798 DVSS.n13767 DVSS.n13733 4.5005
R16799 DVSS.n13767 DVSS.n13740 4.5005
R16800 DVSS.n13767 DVSS.n13732 4.5005
R16801 DVSS.n13767 DVSS.n13741 4.5005
R16802 DVSS.n13767 DVSS.n13731 4.5005
R16803 DVSS.n13767 DVSS.n13743 4.5005
R16804 DVSS.n13767 DVSS.n13744 4.5005
R16805 DVSS.n21142 DVSS.n13767 4.5005
R16806 DVSS.n13752 DVSS.n13736 4.5005
R16807 DVSS.n13752 DVSS.n13735 4.5005
R16808 DVSS.n13752 DVSS.n13738 4.5005
R16809 DVSS.n13752 DVSS.n13734 4.5005
R16810 DVSS.n13752 DVSS.n13739 4.5005
R16811 DVSS.n13752 DVSS.n13733 4.5005
R16812 DVSS.n13752 DVSS.n13740 4.5005
R16813 DVSS.n13752 DVSS.n13732 4.5005
R16814 DVSS.n13752 DVSS.n13741 4.5005
R16815 DVSS.n13752 DVSS.n13731 4.5005
R16816 DVSS.n13752 DVSS.n13743 4.5005
R16817 DVSS.n13752 DVSS.n13744 4.5005
R16818 DVSS.n21142 DVSS.n13752 4.5005
R16819 DVSS.n13769 DVSS.n13736 4.5005
R16820 DVSS.n13769 DVSS.n13735 4.5005
R16821 DVSS.n13769 DVSS.n13738 4.5005
R16822 DVSS.n13769 DVSS.n13734 4.5005
R16823 DVSS.n13769 DVSS.n13739 4.5005
R16824 DVSS.n13769 DVSS.n13733 4.5005
R16825 DVSS.n13769 DVSS.n13740 4.5005
R16826 DVSS.n13769 DVSS.n13732 4.5005
R16827 DVSS.n13769 DVSS.n13741 4.5005
R16828 DVSS.n13769 DVSS.n13731 4.5005
R16829 DVSS.n13769 DVSS.n13743 4.5005
R16830 DVSS.n13769 DVSS.n13744 4.5005
R16831 DVSS.n21142 DVSS.n13769 4.5005
R16832 DVSS.n13751 DVSS.n13736 4.5005
R16833 DVSS.n13751 DVSS.n13735 4.5005
R16834 DVSS.n13751 DVSS.n13738 4.5005
R16835 DVSS.n13751 DVSS.n13734 4.5005
R16836 DVSS.n13751 DVSS.n13739 4.5005
R16837 DVSS.n13751 DVSS.n13733 4.5005
R16838 DVSS.n13751 DVSS.n13740 4.5005
R16839 DVSS.n13751 DVSS.n13732 4.5005
R16840 DVSS.n13751 DVSS.n13741 4.5005
R16841 DVSS.n13751 DVSS.n13731 4.5005
R16842 DVSS.n13751 DVSS.n13743 4.5005
R16843 DVSS.n13751 DVSS.n13744 4.5005
R16844 DVSS.n21142 DVSS.n13751 4.5005
R16845 DVSS.n13771 DVSS.n13736 4.5005
R16846 DVSS.n13771 DVSS.n13735 4.5005
R16847 DVSS.n13771 DVSS.n13738 4.5005
R16848 DVSS.n13771 DVSS.n13734 4.5005
R16849 DVSS.n13771 DVSS.n13739 4.5005
R16850 DVSS.n13771 DVSS.n13733 4.5005
R16851 DVSS.n13771 DVSS.n13740 4.5005
R16852 DVSS.n13771 DVSS.n13732 4.5005
R16853 DVSS.n13771 DVSS.n13741 4.5005
R16854 DVSS.n13771 DVSS.n13731 4.5005
R16855 DVSS.n13771 DVSS.n13743 4.5005
R16856 DVSS.n13771 DVSS.n13744 4.5005
R16857 DVSS.n21142 DVSS.n13771 4.5005
R16858 DVSS.n13750 DVSS.n13736 4.5005
R16859 DVSS.n13750 DVSS.n13735 4.5005
R16860 DVSS.n13750 DVSS.n13738 4.5005
R16861 DVSS.n13750 DVSS.n13734 4.5005
R16862 DVSS.n13750 DVSS.n13739 4.5005
R16863 DVSS.n13750 DVSS.n13733 4.5005
R16864 DVSS.n13750 DVSS.n13740 4.5005
R16865 DVSS.n13750 DVSS.n13732 4.5005
R16866 DVSS.n13750 DVSS.n13741 4.5005
R16867 DVSS.n13750 DVSS.n13731 4.5005
R16868 DVSS.n13750 DVSS.n13743 4.5005
R16869 DVSS.n13750 DVSS.n13744 4.5005
R16870 DVSS.n21142 DVSS.n13750 4.5005
R16871 DVSS.n13773 DVSS.n13736 4.5005
R16872 DVSS.n13773 DVSS.n13735 4.5005
R16873 DVSS.n13773 DVSS.n13738 4.5005
R16874 DVSS.n13773 DVSS.n13734 4.5005
R16875 DVSS.n13773 DVSS.n13739 4.5005
R16876 DVSS.n13773 DVSS.n13733 4.5005
R16877 DVSS.n13773 DVSS.n13740 4.5005
R16878 DVSS.n13773 DVSS.n13732 4.5005
R16879 DVSS.n13773 DVSS.n13741 4.5005
R16880 DVSS.n13773 DVSS.n13731 4.5005
R16881 DVSS.n13773 DVSS.n13743 4.5005
R16882 DVSS.n13773 DVSS.n13744 4.5005
R16883 DVSS.n21142 DVSS.n13773 4.5005
R16884 DVSS.n13749 DVSS.n13736 4.5005
R16885 DVSS.n13749 DVSS.n13735 4.5005
R16886 DVSS.n13749 DVSS.n13738 4.5005
R16887 DVSS.n13749 DVSS.n13734 4.5005
R16888 DVSS.n13749 DVSS.n13739 4.5005
R16889 DVSS.n13749 DVSS.n13733 4.5005
R16890 DVSS.n13749 DVSS.n13740 4.5005
R16891 DVSS.n13749 DVSS.n13732 4.5005
R16892 DVSS.n13749 DVSS.n13741 4.5005
R16893 DVSS.n13749 DVSS.n13731 4.5005
R16894 DVSS.n13749 DVSS.n13743 4.5005
R16895 DVSS.n13749 DVSS.n13744 4.5005
R16896 DVSS.n21142 DVSS.n13749 4.5005
R16897 DVSS.n13775 DVSS.n13736 4.5005
R16898 DVSS.n13775 DVSS.n13735 4.5005
R16899 DVSS.n13775 DVSS.n13738 4.5005
R16900 DVSS.n13775 DVSS.n13734 4.5005
R16901 DVSS.n13775 DVSS.n13739 4.5005
R16902 DVSS.n13775 DVSS.n13733 4.5005
R16903 DVSS.n13775 DVSS.n13740 4.5005
R16904 DVSS.n13775 DVSS.n13732 4.5005
R16905 DVSS.n13775 DVSS.n13741 4.5005
R16906 DVSS.n13775 DVSS.n13731 4.5005
R16907 DVSS.n13775 DVSS.n13743 4.5005
R16908 DVSS.n13775 DVSS.n13744 4.5005
R16909 DVSS.n21142 DVSS.n13775 4.5005
R16910 DVSS.n13748 DVSS.n13736 4.5005
R16911 DVSS.n13748 DVSS.n13735 4.5005
R16912 DVSS.n13748 DVSS.n13738 4.5005
R16913 DVSS.n13748 DVSS.n13734 4.5005
R16914 DVSS.n13748 DVSS.n13739 4.5005
R16915 DVSS.n13748 DVSS.n13733 4.5005
R16916 DVSS.n13748 DVSS.n13740 4.5005
R16917 DVSS.n13748 DVSS.n13732 4.5005
R16918 DVSS.n13748 DVSS.n13741 4.5005
R16919 DVSS.n13748 DVSS.n13731 4.5005
R16920 DVSS.n13748 DVSS.n13743 4.5005
R16921 DVSS.n13748 DVSS.n13744 4.5005
R16922 DVSS.n21142 DVSS.n13748 4.5005
R16923 DVSS.n13777 DVSS.n13736 4.5005
R16924 DVSS.n13777 DVSS.n13735 4.5005
R16925 DVSS.n13777 DVSS.n13738 4.5005
R16926 DVSS.n13777 DVSS.n13734 4.5005
R16927 DVSS.n13777 DVSS.n13739 4.5005
R16928 DVSS.n13777 DVSS.n13733 4.5005
R16929 DVSS.n13777 DVSS.n13740 4.5005
R16930 DVSS.n13777 DVSS.n13732 4.5005
R16931 DVSS.n13777 DVSS.n13741 4.5005
R16932 DVSS.n13777 DVSS.n13731 4.5005
R16933 DVSS.n13777 DVSS.n13743 4.5005
R16934 DVSS.n13777 DVSS.n13744 4.5005
R16935 DVSS.n21142 DVSS.n13777 4.5005
R16936 DVSS.n13747 DVSS.n13736 4.5005
R16937 DVSS.n13747 DVSS.n13735 4.5005
R16938 DVSS.n13747 DVSS.n13738 4.5005
R16939 DVSS.n13747 DVSS.n13734 4.5005
R16940 DVSS.n13747 DVSS.n13739 4.5005
R16941 DVSS.n13747 DVSS.n13733 4.5005
R16942 DVSS.n13747 DVSS.n13740 4.5005
R16943 DVSS.n13747 DVSS.n13732 4.5005
R16944 DVSS.n13747 DVSS.n13741 4.5005
R16945 DVSS.n13747 DVSS.n13731 4.5005
R16946 DVSS.n13747 DVSS.n13743 4.5005
R16947 DVSS.n13747 DVSS.n13744 4.5005
R16948 DVSS.n21142 DVSS.n13747 4.5005
R16949 DVSS.n21141 DVSS.n13736 4.5005
R16950 DVSS.n21141 DVSS.n13735 4.5005
R16951 DVSS.n21141 DVSS.n13738 4.5005
R16952 DVSS.n21141 DVSS.n13734 4.5005
R16953 DVSS.n21141 DVSS.n13739 4.5005
R16954 DVSS.n21141 DVSS.n13733 4.5005
R16955 DVSS.n21141 DVSS.n13740 4.5005
R16956 DVSS.n21141 DVSS.n13732 4.5005
R16957 DVSS.n21141 DVSS.n13741 4.5005
R16958 DVSS.n21141 DVSS.n13731 4.5005
R16959 DVSS.n21141 DVSS.n13743 4.5005
R16960 DVSS.n21141 DVSS.n13744 4.5005
R16961 DVSS.n21142 DVSS.n21141 4.5005
R16962 DVSS.n13746 DVSS.n13736 4.5005
R16963 DVSS.n13746 DVSS.n13735 4.5005
R16964 DVSS.n13746 DVSS.n13738 4.5005
R16965 DVSS.n13746 DVSS.n13734 4.5005
R16966 DVSS.n13746 DVSS.n13739 4.5005
R16967 DVSS.n13746 DVSS.n13733 4.5005
R16968 DVSS.n13746 DVSS.n13740 4.5005
R16969 DVSS.n13746 DVSS.n13732 4.5005
R16970 DVSS.n13746 DVSS.n13741 4.5005
R16971 DVSS.n13746 DVSS.n13731 4.5005
R16972 DVSS.n13746 DVSS.n13743 4.5005
R16973 DVSS.n13746 DVSS.n13744 4.5005
R16974 DVSS.n21142 DVSS.n13746 4.5005
R16975 DVSS.n21143 DVSS.n13736 4.5005
R16976 DVSS.n21143 DVSS.n13735 4.5005
R16977 DVSS.n21143 DVSS.n13738 4.5005
R16978 DVSS.n21143 DVSS.n13734 4.5005
R16979 DVSS.n21143 DVSS.n13739 4.5005
R16980 DVSS.n21143 DVSS.n13733 4.5005
R16981 DVSS.n21143 DVSS.n13740 4.5005
R16982 DVSS.n21143 DVSS.n13732 4.5005
R16983 DVSS.n21143 DVSS.n13741 4.5005
R16984 DVSS.n21143 DVSS.n13731 4.5005
R16985 DVSS.n21143 DVSS.n13743 4.5005
R16986 DVSS.n21143 DVSS.n13730 4.5005
R16987 DVSS.n21143 DVSS.n13744 4.5005
R16988 DVSS.n21143 DVSS.n21142 4.5005
R16989 DVSS.n21144 DVSS.n13691 4.5005
R16990 DVSS.n21144 DVSS.n13712 4.5005
R16991 DVSS.n21144 DVSS.n13715 4.5005
R16992 DVSS.n21144 DVSS.n13711 4.5005
R16993 DVSS.n21144 DVSS.n13716 4.5005
R16994 DVSS.n21144 DVSS.n13710 4.5005
R16995 DVSS.n21144 DVSS.n13717 4.5005
R16996 DVSS.n21144 DVSS.n13727 4.5005
R16997 DVSS.n21144 DVSS.n13719 4.5005
R16998 DVSS.n21145 DVSS.n21144 4.5005
R16999 DVSS.n13696 DVSS.n13691 4.5005
R17000 DVSS.n21147 DVSS.n13696 4.5005
R17001 DVSS.n13714 DVSS.n13696 4.5005
R17002 DVSS.n13712 DVSS.n13696 4.5005
R17003 DVSS.n13715 DVSS.n13696 4.5005
R17004 DVSS.n13711 DVSS.n13696 4.5005
R17005 DVSS.n13716 DVSS.n13696 4.5005
R17006 DVSS.n13710 DVSS.n13696 4.5005
R17007 DVSS.n13717 DVSS.n13696 4.5005
R17008 DVSS.n13709 DVSS.n13696 4.5005
R17009 DVSS.n13718 DVSS.n13696 4.5005
R17010 DVSS.n13719 DVSS.n13696 4.5005
R17011 DVSS.n21145 DVSS.n13696 4.5005
R17012 DVSS.n13698 DVSS.n13691 4.5005
R17013 DVSS.n21147 DVSS.n13698 4.5005
R17014 DVSS.n13714 DVSS.n13698 4.5005
R17015 DVSS.n13712 DVSS.n13698 4.5005
R17016 DVSS.n13715 DVSS.n13698 4.5005
R17017 DVSS.n13711 DVSS.n13698 4.5005
R17018 DVSS.n13716 DVSS.n13698 4.5005
R17019 DVSS.n13710 DVSS.n13698 4.5005
R17020 DVSS.n13717 DVSS.n13698 4.5005
R17021 DVSS.n13709 DVSS.n13698 4.5005
R17022 DVSS.n13718 DVSS.n13698 4.5005
R17023 DVSS.n13719 DVSS.n13698 4.5005
R17024 DVSS.n21145 DVSS.n13698 4.5005
R17025 DVSS.n13695 DVSS.n13691 4.5005
R17026 DVSS.n21147 DVSS.n13695 4.5005
R17027 DVSS.n13714 DVSS.n13695 4.5005
R17028 DVSS.n13712 DVSS.n13695 4.5005
R17029 DVSS.n13715 DVSS.n13695 4.5005
R17030 DVSS.n13711 DVSS.n13695 4.5005
R17031 DVSS.n13716 DVSS.n13695 4.5005
R17032 DVSS.n13710 DVSS.n13695 4.5005
R17033 DVSS.n13717 DVSS.n13695 4.5005
R17034 DVSS.n13709 DVSS.n13695 4.5005
R17035 DVSS.n13718 DVSS.n13695 4.5005
R17036 DVSS.n13719 DVSS.n13695 4.5005
R17037 DVSS.n21145 DVSS.n13695 4.5005
R17038 DVSS.n13699 DVSS.n13691 4.5005
R17039 DVSS.n21147 DVSS.n13699 4.5005
R17040 DVSS.n13714 DVSS.n13699 4.5005
R17041 DVSS.n13712 DVSS.n13699 4.5005
R17042 DVSS.n13715 DVSS.n13699 4.5005
R17043 DVSS.n13711 DVSS.n13699 4.5005
R17044 DVSS.n13716 DVSS.n13699 4.5005
R17045 DVSS.n13710 DVSS.n13699 4.5005
R17046 DVSS.n13717 DVSS.n13699 4.5005
R17047 DVSS.n13709 DVSS.n13699 4.5005
R17048 DVSS.n13718 DVSS.n13699 4.5005
R17049 DVSS.n13719 DVSS.n13699 4.5005
R17050 DVSS.n21145 DVSS.n13699 4.5005
R17051 DVSS.n13694 DVSS.n13691 4.5005
R17052 DVSS.n21147 DVSS.n13694 4.5005
R17053 DVSS.n13714 DVSS.n13694 4.5005
R17054 DVSS.n13712 DVSS.n13694 4.5005
R17055 DVSS.n13715 DVSS.n13694 4.5005
R17056 DVSS.n13711 DVSS.n13694 4.5005
R17057 DVSS.n13716 DVSS.n13694 4.5005
R17058 DVSS.n13710 DVSS.n13694 4.5005
R17059 DVSS.n13717 DVSS.n13694 4.5005
R17060 DVSS.n13709 DVSS.n13694 4.5005
R17061 DVSS.n13718 DVSS.n13694 4.5005
R17062 DVSS.n13719 DVSS.n13694 4.5005
R17063 DVSS.n21145 DVSS.n13694 4.5005
R17064 DVSS.n13700 DVSS.n13691 4.5005
R17065 DVSS.n21147 DVSS.n13700 4.5005
R17066 DVSS.n13714 DVSS.n13700 4.5005
R17067 DVSS.n13712 DVSS.n13700 4.5005
R17068 DVSS.n13715 DVSS.n13700 4.5005
R17069 DVSS.n13711 DVSS.n13700 4.5005
R17070 DVSS.n13716 DVSS.n13700 4.5005
R17071 DVSS.n13710 DVSS.n13700 4.5005
R17072 DVSS.n13717 DVSS.n13700 4.5005
R17073 DVSS.n13709 DVSS.n13700 4.5005
R17074 DVSS.n13718 DVSS.n13700 4.5005
R17075 DVSS.n13719 DVSS.n13700 4.5005
R17076 DVSS.n21145 DVSS.n13700 4.5005
R17077 DVSS.n13693 DVSS.n13691 4.5005
R17078 DVSS.n21147 DVSS.n13693 4.5005
R17079 DVSS.n13714 DVSS.n13693 4.5005
R17080 DVSS.n13712 DVSS.n13693 4.5005
R17081 DVSS.n13715 DVSS.n13693 4.5005
R17082 DVSS.n13711 DVSS.n13693 4.5005
R17083 DVSS.n13716 DVSS.n13693 4.5005
R17084 DVSS.n13710 DVSS.n13693 4.5005
R17085 DVSS.n13717 DVSS.n13693 4.5005
R17086 DVSS.n13709 DVSS.n13693 4.5005
R17087 DVSS.n13718 DVSS.n13693 4.5005
R17088 DVSS.n13719 DVSS.n13693 4.5005
R17089 DVSS.n21145 DVSS.n13693 4.5005
R17090 DVSS.n13701 DVSS.n13691 4.5005
R17091 DVSS.n21147 DVSS.n13701 4.5005
R17092 DVSS.n13714 DVSS.n13701 4.5005
R17093 DVSS.n13712 DVSS.n13701 4.5005
R17094 DVSS.n13715 DVSS.n13701 4.5005
R17095 DVSS.n13711 DVSS.n13701 4.5005
R17096 DVSS.n13716 DVSS.n13701 4.5005
R17097 DVSS.n13710 DVSS.n13701 4.5005
R17098 DVSS.n13717 DVSS.n13701 4.5005
R17099 DVSS.n13709 DVSS.n13701 4.5005
R17100 DVSS.n13718 DVSS.n13701 4.5005
R17101 DVSS.n13719 DVSS.n13701 4.5005
R17102 DVSS.n21145 DVSS.n13701 4.5005
R17103 DVSS.n13692 DVSS.n13691 4.5005
R17104 DVSS.n21147 DVSS.n13692 4.5005
R17105 DVSS.n13714 DVSS.n13692 4.5005
R17106 DVSS.n13712 DVSS.n13692 4.5005
R17107 DVSS.n13715 DVSS.n13692 4.5005
R17108 DVSS.n13711 DVSS.n13692 4.5005
R17109 DVSS.n13716 DVSS.n13692 4.5005
R17110 DVSS.n13710 DVSS.n13692 4.5005
R17111 DVSS.n13717 DVSS.n13692 4.5005
R17112 DVSS.n13709 DVSS.n13692 4.5005
R17113 DVSS.n13718 DVSS.n13692 4.5005
R17114 DVSS.n13719 DVSS.n13692 4.5005
R17115 DVSS.n21145 DVSS.n13692 4.5005
R17116 DVSS.n21146 DVSS.n13691 4.5005
R17117 DVSS.n21147 DVSS.n21146 4.5005
R17118 DVSS.n21146 DVSS.n13714 4.5005
R17119 DVSS.n21146 DVSS.n13712 4.5005
R17120 DVSS.n21146 DVSS.n13715 4.5005
R17121 DVSS.n21146 DVSS.n13711 4.5005
R17122 DVSS.n21146 DVSS.n13716 4.5005
R17123 DVSS.n21146 DVSS.n13710 4.5005
R17124 DVSS.n21146 DVSS.n13717 4.5005
R17125 DVSS.n21146 DVSS.n13709 4.5005
R17126 DVSS.n21146 DVSS.n13718 4.5005
R17127 DVSS.n21146 DVSS.n13719 4.5005
R17128 DVSS.n21146 DVSS.n13707 4.5005
R17129 DVSS.n21146 DVSS.n21145 4.5005
R17130 DVSS.n15153 DVSS.n13702 4.5005
R17131 DVSS.n15175 DVSS.n13702 4.5005
R17132 DVSS.n15178 DVSS.n13702 4.5005
R17133 DVSS.n15174 DVSS.n13702 4.5005
R17134 DVSS.n15179 DVSS.n13702 4.5005
R17135 DVSS.n15173 DVSS.n13702 4.5005
R17136 DVSS.n15180 DVSS.n13702 4.5005
R17137 DVSS.n15214 DVSS.n13702 4.5005
R17138 DVSS.n15183 DVSS.n13702 4.5005
R17139 DVSS.n18490 DVSS.n13702 4.5005
R17140 DVSS.n15158 DVSS.n15153 4.5005
R17141 DVSS.n18492 DVSS.n15158 4.5005
R17142 DVSS.n15177 DVSS.n15158 4.5005
R17143 DVSS.n15175 DVSS.n15158 4.5005
R17144 DVSS.n15178 DVSS.n15158 4.5005
R17145 DVSS.n15174 DVSS.n15158 4.5005
R17146 DVSS.n15179 DVSS.n15158 4.5005
R17147 DVSS.n15173 DVSS.n15158 4.5005
R17148 DVSS.n15180 DVSS.n15158 4.5005
R17149 DVSS.n15172 DVSS.n15158 4.5005
R17150 DVSS.n15182 DVSS.n15158 4.5005
R17151 DVSS.n15183 DVSS.n15158 4.5005
R17152 DVSS.n18490 DVSS.n15158 4.5005
R17153 DVSS.n15160 DVSS.n15153 4.5005
R17154 DVSS.n18492 DVSS.n15160 4.5005
R17155 DVSS.n15177 DVSS.n15160 4.5005
R17156 DVSS.n15175 DVSS.n15160 4.5005
R17157 DVSS.n15178 DVSS.n15160 4.5005
R17158 DVSS.n15174 DVSS.n15160 4.5005
R17159 DVSS.n15179 DVSS.n15160 4.5005
R17160 DVSS.n15173 DVSS.n15160 4.5005
R17161 DVSS.n15180 DVSS.n15160 4.5005
R17162 DVSS.n15172 DVSS.n15160 4.5005
R17163 DVSS.n15182 DVSS.n15160 4.5005
R17164 DVSS.n15183 DVSS.n15160 4.5005
R17165 DVSS.n18490 DVSS.n15160 4.5005
R17166 DVSS.n15157 DVSS.n15153 4.5005
R17167 DVSS.n18492 DVSS.n15157 4.5005
R17168 DVSS.n15177 DVSS.n15157 4.5005
R17169 DVSS.n15175 DVSS.n15157 4.5005
R17170 DVSS.n15178 DVSS.n15157 4.5005
R17171 DVSS.n15174 DVSS.n15157 4.5005
R17172 DVSS.n15179 DVSS.n15157 4.5005
R17173 DVSS.n15173 DVSS.n15157 4.5005
R17174 DVSS.n15180 DVSS.n15157 4.5005
R17175 DVSS.n15172 DVSS.n15157 4.5005
R17176 DVSS.n15182 DVSS.n15157 4.5005
R17177 DVSS.n15183 DVSS.n15157 4.5005
R17178 DVSS.n18490 DVSS.n15157 4.5005
R17179 DVSS.n15161 DVSS.n15153 4.5005
R17180 DVSS.n18492 DVSS.n15161 4.5005
R17181 DVSS.n15177 DVSS.n15161 4.5005
R17182 DVSS.n15175 DVSS.n15161 4.5005
R17183 DVSS.n15178 DVSS.n15161 4.5005
R17184 DVSS.n15174 DVSS.n15161 4.5005
R17185 DVSS.n15179 DVSS.n15161 4.5005
R17186 DVSS.n15173 DVSS.n15161 4.5005
R17187 DVSS.n15180 DVSS.n15161 4.5005
R17188 DVSS.n15172 DVSS.n15161 4.5005
R17189 DVSS.n15182 DVSS.n15161 4.5005
R17190 DVSS.n15183 DVSS.n15161 4.5005
R17191 DVSS.n18490 DVSS.n15161 4.5005
R17192 DVSS.n15156 DVSS.n15153 4.5005
R17193 DVSS.n18492 DVSS.n15156 4.5005
R17194 DVSS.n15177 DVSS.n15156 4.5005
R17195 DVSS.n15175 DVSS.n15156 4.5005
R17196 DVSS.n15178 DVSS.n15156 4.5005
R17197 DVSS.n15174 DVSS.n15156 4.5005
R17198 DVSS.n15179 DVSS.n15156 4.5005
R17199 DVSS.n15173 DVSS.n15156 4.5005
R17200 DVSS.n15180 DVSS.n15156 4.5005
R17201 DVSS.n15172 DVSS.n15156 4.5005
R17202 DVSS.n15182 DVSS.n15156 4.5005
R17203 DVSS.n15183 DVSS.n15156 4.5005
R17204 DVSS.n18490 DVSS.n15156 4.5005
R17205 DVSS.n15162 DVSS.n15153 4.5005
R17206 DVSS.n18492 DVSS.n15162 4.5005
R17207 DVSS.n15177 DVSS.n15162 4.5005
R17208 DVSS.n15175 DVSS.n15162 4.5005
R17209 DVSS.n15178 DVSS.n15162 4.5005
R17210 DVSS.n15174 DVSS.n15162 4.5005
R17211 DVSS.n15179 DVSS.n15162 4.5005
R17212 DVSS.n15173 DVSS.n15162 4.5005
R17213 DVSS.n15180 DVSS.n15162 4.5005
R17214 DVSS.n15172 DVSS.n15162 4.5005
R17215 DVSS.n15182 DVSS.n15162 4.5005
R17216 DVSS.n15183 DVSS.n15162 4.5005
R17217 DVSS.n18490 DVSS.n15162 4.5005
R17218 DVSS.n15155 DVSS.n15153 4.5005
R17219 DVSS.n18492 DVSS.n15155 4.5005
R17220 DVSS.n15177 DVSS.n15155 4.5005
R17221 DVSS.n15175 DVSS.n15155 4.5005
R17222 DVSS.n15178 DVSS.n15155 4.5005
R17223 DVSS.n15174 DVSS.n15155 4.5005
R17224 DVSS.n15179 DVSS.n15155 4.5005
R17225 DVSS.n15173 DVSS.n15155 4.5005
R17226 DVSS.n15180 DVSS.n15155 4.5005
R17227 DVSS.n15172 DVSS.n15155 4.5005
R17228 DVSS.n15182 DVSS.n15155 4.5005
R17229 DVSS.n15183 DVSS.n15155 4.5005
R17230 DVSS.n18490 DVSS.n15155 4.5005
R17231 DVSS.n15163 DVSS.n15153 4.5005
R17232 DVSS.n18492 DVSS.n15163 4.5005
R17233 DVSS.n15177 DVSS.n15163 4.5005
R17234 DVSS.n15175 DVSS.n15163 4.5005
R17235 DVSS.n15178 DVSS.n15163 4.5005
R17236 DVSS.n15174 DVSS.n15163 4.5005
R17237 DVSS.n15179 DVSS.n15163 4.5005
R17238 DVSS.n15173 DVSS.n15163 4.5005
R17239 DVSS.n15180 DVSS.n15163 4.5005
R17240 DVSS.n15172 DVSS.n15163 4.5005
R17241 DVSS.n15182 DVSS.n15163 4.5005
R17242 DVSS.n15183 DVSS.n15163 4.5005
R17243 DVSS.n18490 DVSS.n15163 4.5005
R17244 DVSS.n15154 DVSS.n15153 4.5005
R17245 DVSS.n18492 DVSS.n15154 4.5005
R17246 DVSS.n15177 DVSS.n15154 4.5005
R17247 DVSS.n15175 DVSS.n15154 4.5005
R17248 DVSS.n15178 DVSS.n15154 4.5005
R17249 DVSS.n15174 DVSS.n15154 4.5005
R17250 DVSS.n15179 DVSS.n15154 4.5005
R17251 DVSS.n15173 DVSS.n15154 4.5005
R17252 DVSS.n15180 DVSS.n15154 4.5005
R17253 DVSS.n15172 DVSS.n15154 4.5005
R17254 DVSS.n15182 DVSS.n15154 4.5005
R17255 DVSS.n15183 DVSS.n15154 4.5005
R17256 DVSS.n18490 DVSS.n15154 4.5005
R17257 DVSS.n18491 DVSS.n15153 4.5005
R17258 DVSS.n18492 DVSS.n18491 4.5005
R17259 DVSS.n18491 DVSS.n15177 4.5005
R17260 DVSS.n18491 DVSS.n15175 4.5005
R17261 DVSS.n18491 DVSS.n15178 4.5005
R17262 DVSS.n18491 DVSS.n15174 4.5005
R17263 DVSS.n18491 DVSS.n15179 4.5005
R17264 DVSS.n18491 DVSS.n15173 4.5005
R17265 DVSS.n18491 DVSS.n15180 4.5005
R17266 DVSS.n18491 DVSS.n15172 4.5005
R17267 DVSS.n18491 DVSS.n15182 4.5005
R17268 DVSS.n18491 DVSS.n15183 4.5005
R17269 DVSS.n18491 DVSS.n15170 4.5005
R17270 DVSS.n18491 DVSS.n18490 4.5005
R17271 DVSS.n17682 DVSS.n15164 4.5005
R17272 DVSS.n17680 DVSS.n15164 4.5005
R17273 DVSS.n17685 DVSS.n15164 4.5005
R17274 DVSS.n17679 DVSS.n15164 4.5005
R17275 DVSS.n17686 DVSS.n15164 4.5005
R17276 DVSS.n17678 DVSS.n15164 4.5005
R17277 DVSS.n17687 DVSS.n15164 4.5005
R17278 DVSS.n17771 DVSS.n15164 4.5005
R17279 DVSS.n17690 DVSS.n15164 4.5005
R17280 DVSS.n17774 DVSS.n15164 4.5005
R17281 DVSS.n17697 DVSS.n17682 4.5005
R17282 DVSS.n17697 DVSS.n17681 4.5005
R17283 DVSS.n17697 DVSS.n17684 4.5005
R17284 DVSS.n17697 DVSS.n17680 4.5005
R17285 DVSS.n17697 DVSS.n17685 4.5005
R17286 DVSS.n17697 DVSS.n17679 4.5005
R17287 DVSS.n17697 DVSS.n17686 4.5005
R17288 DVSS.n17697 DVSS.n17678 4.5005
R17289 DVSS.n17697 DVSS.n17687 4.5005
R17290 DVSS.n17697 DVSS.n17677 4.5005
R17291 DVSS.n17697 DVSS.n17689 4.5005
R17292 DVSS.n17697 DVSS.n17690 4.5005
R17293 DVSS.n17774 DVSS.n17697 4.5005
R17294 DVSS.n17700 DVSS.n17682 4.5005
R17295 DVSS.n17700 DVSS.n17681 4.5005
R17296 DVSS.n17700 DVSS.n17684 4.5005
R17297 DVSS.n17700 DVSS.n17680 4.5005
R17298 DVSS.n17700 DVSS.n17685 4.5005
R17299 DVSS.n17700 DVSS.n17679 4.5005
R17300 DVSS.n17700 DVSS.n17686 4.5005
R17301 DVSS.n17700 DVSS.n17678 4.5005
R17302 DVSS.n17700 DVSS.n17687 4.5005
R17303 DVSS.n17700 DVSS.n17677 4.5005
R17304 DVSS.n17700 DVSS.n17689 4.5005
R17305 DVSS.n17700 DVSS.n17690 4.5005
R17306 DVSS.n17774 DVSS.n17700 4.5005
R17307 DVSS.n17695 DVSS.n17682 4.5005
R17308 DVSS.n17695 DVSS.n17681 4.5005
R17309 DVSS.n17695 DVSS.n17684 4.5005
R17310 DVSS.n17695 DVSS.n17680 4.5005
R17311 DVSS.n17695 DVSS.n17685 4.5005
R17312 DVSS.n17695 DVSS.n17679 4.5005
R17313 DVSS.n17695 DVSS.n17686 4.5005
R17314 DVSS.n17695 DVSS.n17678 4.5005
R17315 DVSS.n17695 DVSS.n17687 4.5005
R17316 DVSS.n17695 DVSS.n17677 4.5005
R17317 DVSS.n17695 DVSS.n17689 4.5005
R17318 DVSS.n17695 DVSS.n17690 4.5005
R17319 DVSS.n17774 DVSS.n17695 4.5005
R17320 DVSS.n17702 DVSS.n17682 4.5005
R17321 DVSS.n17702 DVSS.n17681 4.5005
R17322 DVSS.n17702 DVSS.n17684 4.5005
R17323 DVSS.n17702 DVSS.n17680 4.5005
R17324 DVSS.n17702 DVSS.n17685 4.5005
R17325 DVSS.n17702 DVSS.n17679 4.5005
R17326 DVSS.n17702 DVSS.n17686 4.5005
R17327 DVSS.n17702 DVSS.n17678 4.5005
R17328 DVSS.n17702 DVSS.n17687 4.5005
R17329 DVSS.n17702 DVSS.n17677 4.5005
R17330 DVSS.n17702 DVSS.n17689 4.5005
R17331 DVSS.n17702 DVSS.n17690 4.5005
R17332 DVSS.n17774 DVSS.n17702 4.5005
R17333 DVSS.n17694 DVSS.n17682 4.5005
R17334 DVSS.n17694 DVSS.n17681 4.5005
R17335 DVSS.n17694 DVSS.n17684 4.5005
R17336 DVSS.n17694 DVSS.n17680 4.5005
R17337 DVSS.n17694 DVSS.n17685 4.5005
R17338 DVSS.n17694 DVSS.n17679 4.5005
R17339 DVSS.n17694 DVSS.n17686 4.5005
R17340 DVSS.n17694 DVSS.n17678 4.5005
R17341 DVSS.n17694 DVSS.n17687 4.5005
R17342 DVSS.n17694 DVSS.n17677 4.5005
R17343 DVSS.n17694 DVSS.n17689 4.5005
R17344 DVSS.n17694 DVSS.n17690 4.5005
R17345 DVSS.n17774 DVSS.n17694 4.5005
R17346 DVSS.n17704 DVSS.n17682 4.5005
R17347 DVSS.n17704 DVSS.n17681 4.5005
R17348 DVSS.n17704 DVSS.n17684 4.5005
R17349 DVSS.n17704 DVSS.n17680 4.5005
R17350 DVSS.n17704 DVSS.n17685 4.5005
R17351 DVSS.n17704 DVSS.n17679 4.5005
R17352 DVSS.n17704 DVSS.n17686 4.5005
R17353 DVSS.n17704 DVSS.n17678 4.5005
R17354 DVSS.n17704 DVSS.n17687 4.5005
R17355 DVSS.n17704 DVSS.n17677 4.5005
R17356 DVSS.n17704 DVSS.n17689 4.5005
R17357 DVSS.n17704 DVSS.n17690 4.5005
R17358 DVSS.n17774 DVSS.n17704 4.5005
R17359 DVSS.n17693 DVSS.n17682 4.5005
R17360 DVSS.n17693 DVSS.n17681 4.5005
R17361 DVSS.n17693 DVSS.n17684 4.5005
R17362 DVSS.n17693 DVSS.n17680 4.5005
R17363 DVSS.n17693 DVSS.n17685 4.5005
R17364 DVSS.n17693 DVSS.n17679 4.5005
R17365 DVSS.n17693 DVSS.n17686 4.5005
R17366 DVSS.n17693 DVSS.n17678 4.5005
R17367 DVSS.n17693 DVSS.n17687 4.5005
R17368 DVSS.n17693 DVSS.n17677 4.5005
R17369 DVSS.n17693 DVSS.n17689 4.5005
R17370 DVSS.n17693 DVSS.n17690 4.5005
R17371 DVSS.n17774 DVSS.n17693 4.5005
R17372 DVSS.n17773 DVSS.n17682 4.5005
R17373 DVSS.n17773 DVSS.n17681 4.5005
R17374 DVSS.n17773 DVSS.n17684 4.5005
R17375 DVSS.n17773 DVSS.n17680 4.5005
R17376 DVSS.n17773 DVSS.n17685 4.5005
R17377 DVSS.n17773 DVSS.n17679 4.5005
R17378 DVSS.n17773 DVSS.n17686 4.5005
R17379 DVSS.n17773 DVSS.n17678 4.5005
R17380 DVSS.n17773 DVSS.n17687 4.5005
R17381 DVSS.n17773 DVSS.n17677 4.5005
R17382 DVSS.n17773 DVSS.n17689 4.5005
R17383 DVSS.n17773 DVSS.n17690 4.5005
R17384 DVSS.n17774 DVSS.n17773 4.5005
R17385 DVSS.n17692 DVSS.n17682 4.5005
R17386 DVSS.n17692 DVSS.n17681 4.5005
R17387 DVSS.n17692 DVSS.n17684 4.5005
R17388 DVSS.n17692 DVSS.n17680 4.5005
R17389 DVSS.n17692 DVSS.n17685 4.5005
R17390 DVSS.n17692 DVSS.n17679 4.5005
R17391 DVSS.n17692 DVSS.n17686 4.5005
R17392 DVSS.n17692 DVSS.n17678 4.5005
R17393 DVSS.n17692 DVSS.n17687 4.5005
R17394 DVSS.n17692 DVSS.n17677 4.5005
R17395 DVSS.n17692 DVSS.n17689 4.5005
R17396 DVSS.n17692 DVSS.n17690 4.5005
R17397 DVSS.n17774 DVSS.n17692 4.5005
R17398 DVSS.n17775 DVSS.n17682 4.5005
R17399 DVSS.n17775 DVSS.n17681 4.5005
R17400 DVSS.n17775 DVSS.n17684 4.5005
R17401 DVSS.n17775 DVSS.n17680 4.5005
R17402 DVSS.n17775 DVSS.n17685 4.5005
R17403 DVSS.n17775 DVSS.n17679 4.5005
R17404 DVSS.n17775 DVSS.n17686 4.5005
R17405 DVSS.n17775 DVSS.n17678 4.5005
R17406 DVSS.n17775 DVSS.n17687 4.5005
R17407 DVSS.n17775 DVSS.n17677 4.5005
R17408 DVSS.n17775 DVSS.n17689 4.5005
R17409 DVSS.n17775 DVSS.n17690 4.5005
R17410 DVSS.n17775 DVSS.n17675 4.5005
R17411 DVSS.n17775 DVSS.n17774 4.5005
R17412 DVSS.n17776 DVSS.n15926 4.5005
R17413 DVSS.n17776 DVSS.n15947 4.5005
R17414 DVSS.n17776 DVSS.n15950 4.5005
R17415 DVSS.n17776 DVSS.n15946 4.5005
R17416 DVSS.n17776 DVSS.n15951 4.5005
R17417 DVSS.n17776 DVSS.n15945 4.5005
R17418 DVSS.n17776 DVSS.n15952 4.5005
R17419 DVSS.n17776 DVSS.n17673 4.5005
R17420 DVSS.n17776 DVSS.n15954 4.5005
R17421 DVSS.n17777 DVSS.n17776 4.5005
R17422 DVSS.n15931 DVSS.n15926 4.5005
R17423 DVSS.n17779 DVSS.n15931 4.5005
R17424 DVSS.n15949 DVSS.n15931 4.5005
R17425 DVSS.n15947 DVSS.n15931 4.5005
R17426 DVSS.n15950 DVSS.n15931 4.5005
R17427 DVSS.n15946 DVSS.n15931 4.5005
R17428 DVSS.n15951 DVSS.n15931 4.5005
R17429 DVSS.n15945 DVSS.n15931 4.5005
R17430 DVSS.n15952 DVSS.n15931 4.5005
R17431 DVSS.n15944 DVSS.n15931 4.5005
R17432 DVSS.n15953 DVSS.n15931 4.5005
R17433 DVSS.n15954 DVSS.n15931 4.5005
R17434 DVSS.n17777 DVSS.n15931 4.5005
R17435 DVSS.n15933 DVSS.n15926 4.5005
R17436 DVSS.n17779 DVSS.n15933 4.5005
R17437 DVSS.n15949 DVSS.n15933 4.5005
R17438 DVSS.n15947 DVSS.n15933 4.5005
R17439 DVSS.n15950 DVSS.n15933 4.5005
R17440 DVSS.n15946 DVSS.n15933 4.5005
R17441 DVSS.n15951 DVSS.n15933 4.5005
R17442 DVSS.n15945 DVSS.n15933 4.5005
R17443 DVSS.n15952 DVSS.n15933 4.5005
R17444 DVSS.n15944 DVSS.n15933 4.5005
R17445 DVSS.n15953 DVSS.n15933 4.5005
R17446 DVSS.n15954 DVSS.n15933 4.5005
R17447 DVSS.n17777 DVSS.n15933 4.5005
R17448 DVSS.n15930 DVSS.n15926 4.5005
R17449 DVSS.n17779 DVSS.n15930 4.5005
R17450 DVSS.n15949 DVSS.n15930 4.5005
R17451 DVSS.n15947 DVSS.n15930 4.5005
R17452 DVSS.n15950 DVSS.n15930 4.5005
R17453 DVSS.n15946 DVSS.n15930 4.5005
R17454 DVSS.n15951 DVSS.n15930 4.5005
R17455 DVSS.n15945 DVSS.n15930 4.5005
R17456 DVSS.n15952 DVSS.n15930 4.5005
R17457 DVSS.n15944 DVSS.n15930 4.5005
R17458 DVSS.n15953 DVSS.n15930 4.5005
R17459 DVSS.n15954 DVSS.n15930 4.5005
R17460 DVSS.n17777 DVSS.n15930 4.5005
R17461 DVSS.n15934 DVSS.n15926 4.5005
R17462 DVSS.n17779 DVSS.n15934 4.5005
R17463 DVSS.n15949 DVSS.n15934 4.5005
R17464 DVSS.n15947 DVSS.n15934 4.5005
R17465 DVSS.n15950 DVSS.n15934 4.5005
R17466 DVSS.n15946 DVSS.n15934 4.5005
R17467 DVSS.n15951 DVSS.n15934 4.5005
R17468 DVSS.n15945 DVSS.n15934 4.5005
R17469 DVSS.n15952 DVSS.n15934 4.5005
R17470 DVSS.n15944 DVSS.n15934 4.5005
R17471 DVSS.n15953 DVSS.n15934 4.5005
R17472 DVSS.n15954 DVSS.n15934 4.5005
R17473 DVSS.n17777 DVSS.n15934 4.5005
R17474 DVSS.n15929 DVSS.n15926 4.5005
R17475 DVSS.n17779 DVSS.n15929 4.5005
R17476 DVSS.n15949 DVSS.n15929 4.5005
R17477 DVSS.n15947 DVSS.n15929 4.5005
R17478 DVSS.n15950 DVSS.n15929 4.5005
R17479 DVSS.n15946 DVSS.n15929 4.5005
R17480 DVSS.n15951 DVSS.n15929 4.5005
R17481 DVSS.n15945 DVSS.n15929 4.5005
R17482 DVSS.n15952 DVSS.n15929 4.5005
R17483 DVSS.n15944 DVSS.n15929 4.5005
R17484 DVSS.n15953 DVSS.n15929 4.5005
R17485 DVSS.n15954 DVSS.n15929 4.5005
R17486 DVSS.n17777 DVSS.n15929 4.5005
R17487 DVSS.n15935 DVSS.n15926 4.5005
R17488 DVSS.n17779 DVSS.n15935 4.5005
R17489 DVSS.n15949 DVSS.n15935 4.5005
R17490 DVSS.n15947 DVSS.n15935 4.5005
R17491 DVSS.n15950 DVSS.n15935 4.5005
R17492 DVSS.n15946 DVSS.n15935 4.5005
R17493 DVSS.n15951 DVSS.n15935 4.5005
R17494 DVSS.n15945 DVSS.n15935 4.5005
R17495 DVSS.n15952 DVSS.n15935 4.5005
R17496 DVSS.n15944 DVSS.n15935 4.5005
R17497 DVSS.n15953 DVSS.n15935 4.5005
R17498 DVSS.n15954 DVSS.n15935 4.5005
R17499 DVSS.n17777 DVSS.n15935 4.5005
R17500 DVSS.n15928 DVSS.n15926 4.5005
R17501 DVSS.n17779 DVSS.n15928 4.5005
R17502 DVSS.n15949 DVSS.n15928 4.5005
R17503 DVSS.n15947 DVSS.n15928 4.5005
R17504 DVSS.n15950 DVSS.n15928 4.5005
R17505 DVSS.n15946 DVSS.n15928 4.5005
R17506 DVSS.n15951 DVSS.n15928 4.5005
R17507 DVSS.n15945 DVSS.n15928 4.5005
R17508 DVSS.n15952 DVSS.n15928 4.5005
R17509 DVSS.n15944 DVSS.n15928 4.5005
R17510 DVSS.n15953 DVSS.n15928 4.5005
R17511 DVSS.n15954 DVSS.n15928 4.5005
R17512 DVSS.n17777 DVSS.n15928 4.5005
R17513 DVSS.n15936 DVSS.n15926 4.5005
R17514 DVSS.n17779 DVSS.n15936 4.5005
R17515 DVSS.n15949 DVSS.n15936 4.5005
R17516 DVSS.n15947 DVSS.n15936 4.5005
R17517 DVSS.n15950 DVSS.n15936 4.5005
R17518 DVSS.n15946 DVSS.n15936 4.5005
R17519 DVSS.n15951 DVSS.n15936 4.5005
R17520 DVSS.n15945 DVSS.n15936 4.5005
R17521 DVSS.n15952 DVSS.n15936 4.5005
R17522 DVSS.n15944 DVSS.n15936 4.5005
R17523 DVSS.n15953 DVSS.n15936 4.5005
R17524 DVSS.n15954 DVSS.n15936 4.5005
R17525 DVSS.n17777 DVSS.n15936 4.5005
R17526 DVSS.n15927 DVSS.n15926 4.5005
R17527 DVSS.n17779 DVSS.n15927 4.5005
R17528 DVSS.n15949 DVSS.n15927 4.5005
R17529 DVSS.n15947 DVSS.n15927 4.5005
R17530 DVSS.n15950 DVSS.n15927 4.5005
R17531 DVSS.n15946 DVSS.n15927 4.5005
R17532 DVSS.n15951 DVSS.n15927 4.5005
R17533 DVSS.n15945 DVSS.n15927 4.5005
R17534 DVSS.n15952 DVSS.n15927 4.5005
R17535 DVSS.n15944 DVSS.n15927 4.5005
R17536 DVSS.n15953 DVSS.n15927 4.5005
R17537 DVSS.n15954 DVSS.n15927 4.5005
R17538 DVSS.n17777 DVSS.n15927 4.5005
R17539 DVSS.n17778 DVSS.n15926 4.5005
R17540 DVSS.n17779 DVSS.n17778 4.5005
R17541 DVSS.n17778 DVSS.n15949 4.5005
R17542 DVSS.n17778 DVSS.n15947 4.5005
R17543 DVSS.n17778 DVSS.n15950 4.5005
R17544 DVSS.n17778 DVSS.n15946 4.5005
R17545 DVSS.n17778 DVSS.n15951 4.5005
R17546 DVSS.n17778 DVSS.n15945 4.5005
R17547 DVSS.n17778 DVSS.n15952 4.5005
R17548 DVSS.n17778 DVSS.n15944 4.5005
R17549 DVSS.n17778 DVSS.n15953 4.5005
R17550 DVSS.n17778 DVSS.n15954 4.5005
R17551 DVSS.n17778 DVSS.n15942 4.5005
R17552 DVSS.n17778 DVSS.n17777 4.5005
R17553 DVSS.n16551 DVSS.n15937 4.5005
R17554 DVSS.n16352 DVSS.n15937 4.5005
R17555 DVSS.n16554 DVSS.n15937 4.5005
R17556 DVSS.n16351 DVSS.n15937 4.5005
R17557 DVSS.n16555 DVSS.n15937 4.5005
R17558 DVSS.n16350 DVSS.n15937 4.5005
R17559 DVSS.n16556 DVSS.n15937 4.5005
R17560 DVSS.n16348 DVSS.n15937 4.5005
R17561 DVSS.n16595 DVSS.n15937 4.5005
R17562 DVSS.n16597 DVSS.n15937 4.5005
R17563 DVSS.n16551 DVSS.n16339 4.5005
R17564 DVSS.n16353 DVSS.n16339 4.5005
R17565 DVSS.n16553 DVSS.n16339 4.5005
R17566 DVSS.n16352 DVSS.n16339 4.5005
R17567 DVSS.n16554 DVSS.n16339 4.5005
R17568 DVSS.n16351 DVSS.n16339 4.5005
R17569 DVSS.n16555 DVSS.n16339 4.5005
R17570 DVSS.n16350 DVSS.n16339 4.5005
R17571 DVSS.n16556 DVSS.n16339 4.5005
R17572 DVSS.n16349 DVSS.n16339 4.5005
R17573 DVSS.n16558 DVSS.n16339 4.5005
R17574 DVSS.n16595 DVSS.n16339 4.5005
R17575 DVSS.n16597 DVSS.n16339 4.5005
R17576 DVSS.n16551 DVSS.n16340 4.5005
R17577 DVSS.n16353 DVSS.n16340 4.5005
R17578 DVSS.n16553 DVSS.n16340 4.5005
R17579 DVSS.n16352 DVSS.n16340 4.5005
R17580 DVSS.n16554 DVSS.n16340 4.5005
R17581 DVSS.n16351 DVSS.n16340 4.5005
R17582 DVSS.n16555 DVSS.n16340 4.5005
R17583 DVSS.n16350 DVSS.n16340 4.5005
R17584 DVSS.n16556 DVSS.n16340 4.5005
R17585 DVSS.n16349 DVSS.n16340 4.5005
R17586 DVSS.n16558 DVSS.n16340 4.5005
R17587 DVSS.n16595 DVSS.n16340 4.5005
R17588 DVSS.n16346 DVSS.n16340 4.5005
R17589 DVSS.n16597 DVSS.n16340 4.5005
R17590 DVSS.n16551 DVSS.n16338 4.5005
R17591 DVSS.n16353 DVSS.n16338 4.5005
R17592 DVSS.n16553 DVSS.n16338 4.5005
R17593 DVSS.n16352 DVSS.n16338 4.5005
R17594 DVSS.n16554 DVSS.n16338 4.5005
R17595 DVSS.n16351 DVSS.n16338 4.5005
R17596 DVSS.n16555 DVSS.n16338 4.5005
R17597 DVSS.n16350 DVSS.n16338 4.5005
R17598 DVSS.n16556 DVSS.n16338 4.5005
R17599 DVSS.n16349 DVSS.n16338 4.5005
R17600 DVSS.n16558 DVSS.n16338 4.5005
R17601 DVSS.n16348 DVSS.n16338 4.5005
R17602 DVSS.n16595 DVSS.n16338 4.5005
R17603 DVSS.n16346 DVSS.n16338 4.5005
R17604 DVSS.n16597 DVSS.n16338 4.5005
R17605 DVSS.n16551 DVSS.n16341 4.5005
R17606 DVSS.n16353 DVSS.n16341 4.5005
R17607 DVSS.n16553 DVSS.n16341 4.5005
R17608 DVSS.n16352 DVSS.n16341 4.5005
R17609 DVSS.n16554 DVSS.n16341 4.5005
R17610 DVSS.n16351 DVSS.n16341 4.5005
R17611 DVSS.n16555 DVSS.n16341 4.5005
R17612 DVSS.n16350 DVSS.n16341 4.5005
R17613 DVSS.n16556 DVSS.n16341 4.5005
R17614 DVSS.n16349 DVSS.n16341 4.5005
R17615 DVSS.n16558 DVSS.n16341 4.5005
R17616 DVSS.n16348 DVSS.n16341 4.5005
R17617 DVSS.n16595 DVSS.n16341 4.5005
R17618 DVSS.n16346 DVSS.n16341 4.5005
R17619 DVSS.n16597 DVSS.n16341 4.5005
R17620 DVSS.n16551 DVSS.n16337 4.5005
R17621 DVSS.n16353 DVSS.n16337 4.5005
R17622 DVSS.n16553 DVSS.n16337 4.5005
R17623 DVSS.n16352 DVSS.n16337 4.5005
R17624 DVSS.n16554 DVSS.n16337 4.5005
R17625 DVSS.n16351 DVSS.n16337 4.5005
R17626 DVSS.n16555 DVSS.n16337 4.5005
R17627 DVSS.n16350 DVSS.n16337 4.5005
R17628 DVSS.n16556 DVSS.n16337 4.5005
R17629 DVSS.n16349 DVSS.n16337 4.5005
R17630 DVSS.n16558 DVSS.n16337 4.5005
R17631 DVSS.n16348 DVSS.n16337 4.5005
R17632 DVSS.n16595 DVSS.n16337 4.5005
R17633 DVSS.n16346 DVSS.n16337 4.5005
R17634 DVSS.n16597 DVSS.n16337 4.5005
R17635 DVSS.n16551 DVSS.n16342 4.5005
R17636 DVSS.n16353 DVSS.n16342 4.5005
R17637 DVSS.n16553 DVSS.n16342 4.5005
R17638 DVSS.n16352 DVSS.n16342 4.5005
R17639 DVSS.n16554 DVSS.n16342 4.5005
R17640 DVSS.n16351 DVSS.n16342 4.5005
R17641 DVSS.n16555 DVSS.n16342 4.5005
R17642 DVSS.n16350 DVSS.n16342 4.5005
R17643 DVSS.n16556 DVSS.n16342 4.5005
R17644 DVSS.n16349 DVSS.n16342 4.5005
R17645 DVSS.n16558 DVSS.n16342 4.5005
R17646 DVSS.n16348 DVSS.n16342 4.5005
R17647 DVSS.n16595 DVSS.n16342 4.5005
R17648 DVSS.n16346 DVSS.n16342 4.5005
R17649 DVSS.n16597 DVSS.n16342 4.5005
R17650 DVSS.n16551 DVSS.n16336 4.5005
R17651 DVSS.n16353 DVSS.n16336 4.5005
R17652 DVSS.n16553 DVSS.n16336 4.5005
R17653 DVSS.n16352 DVSS.n16336 4.5005
R17654 DVSS.n16554 DVSS.n16336 4.5005
R17655 DVSS.n16351 DVSS.n16336 4.5005
R17656 DVSS.n16555 DVSS.n16336 4.5005
R17657 DVSS.n16350 DVSS.n16336 4.5005
R17658 DVSS.n16556 DVSS.n16336 4.5005
R17659 DVSS.n16349 DVSS.n16336 4.5005
R17660 DVSS.n16558 DVSS.n16336 4.5005
R17661 DVSS.n16348 DVSS.n16336 4.5005
R17662 DVSS.n16595 DVSS.n16336 4.5005
R17663 DVSS.n16346 DVSS.n16336 4.5005
R17664 DVSS.n16597 DVSS.n16336 4.5005
R17665 DVSS.n15900 DVSS.n15883 4.5005
R17666 DVSS.n15897 DVSS.n15883 4.5005
R17667 DVSS.n15903 DVSS.n15883 4.5005
R17668 DVSS.n15896 DVSS.n15883 4.5005
R17669 DVSS.n15904 DVSS.n15883 4.5005
R17670 DVSS.n15895 DVSS.n15883 4.5005
R17671 DVSS.n15905 DVSS.n15883 4.5005
R17672 DVSS.n15893 DVSS.n15883 4.5005
R17673 DVSS.n17821 DVSS.n15883 4.5005
R17674 DVSS.n15891 DVSS.n15883 4.5005
R17675 DVSS.n17823 DVSS.n15883 4.5005
R17676 DVSS.n15900 DVSS.n15884 4.5005
R17677 DVSS.n15898 DVSS.n15884 4.5005
R17678 DVSS.n15902 DVSS.n15884 4.5005
R17679 DVSS.n15897 DVSS.n15884 4.5005
R17680 DVSS.n15903 DVSS.n15884 4.5005
R17681 DVSS.n15896 DVSS.n15884 4.5005
R17682 DVSS.n15904 DVSS.n15884 4.5005
R17683 DVSS.n15895 DVSS.n15884 4.5005
R17684 DVSS.n15905 DVSS.n15884 4.5005
R17685 DVSS.n15894 DVSS.n15884 4.5005
R17686 DVSS.n15907 DVSS.n15884 4.5005
R17687 DVSS.n15893 DVSS.n15884 4.5005
R17688 DVSS.n17821 DVSS.n15884 4.5005
R17689 DVSS.n15891 DVSS.n15884 4.5005
R17690 DVSS.n17823 DVSS.n15884 4.5005
R17691 DVSS.n15900 DVSS.n15882 4.5005
R17692 DVSS.n15898 DVSS.n15882 4.5005
R17693 DVSS.n15902 DVSS.n15882 4.5005
R17694 DVSS.n15897 DVSS.n15882 4.5005
R17695 DVSS.n15903 DVSS.n15882 4.5005
R17696 DVSS.n15896 DVSS.n15882 4.5005
R17697 DVSS.n15904 DVSS.n15882 4.5005
R17698 DVSS.n15895 DVSS.n15882 4.5005
R17699 DVSS.n15905 DVSS.n15882 4.5005
R17700 DVSS.n15894 DVSS.n15882 4.5005
R17701 DVSS.n15907 DVSS.n15882 4.5005
R17702 DVSS.n15893 DVSS.n15882 4.5005
R17703 DVSS.n17821 DVSS.n15882 4.5005
R17704 DVSS.n15891 DVSS.n15882 4.5005
R17705 DVSS.n17823 DVSS.n15882 4.5005
R17706 DVSS.n15900 DVSS.n15885 4.5005
R17707 DVSS.n15898 DVSS.n15885 4.5005
R17708 DVSS.n15902 DVSS.n15885 4.5005
R17709 DVSS.n15897 DVSS.n15885 4.5005
R17710 DVSS.n15903 DVSS.n15885 4.5005
R17711 DVSS.n15896 DVSS.n15885 4.5005
R17712 DVSS.n15904 DVSS.n15885 4.5005
R17713 DVSS.n15895 DVSS.n15885 4.5005
R17714 DVSS.n15905 DVSS.n15885 4.5005
R17715 DVSS.n15894 DVSS.n15885 4.5005
R17716 DVSS.n15907 DVSS.n15885 4.5005
R17717 DVSS.n15893 DVSS.n15885 4.5005
R17718 DVSS.n17821 DVSS.n15885 4.5005
R17719 DVSS.n15891 DVSS.n15885 4.5005
R17720 DVSS.n17823 DVSS.n15885 4.5005
R17721 DVSS.n15900 DVSS.n15881 4.5005
R17722 DVSS.n15898 DVSS.n15881 4.5005
R17723 DVSS.n15902 DVSS.n15881 4.5005
R17724 DVSS.n15897 DVSS.n15881 4.5005
R17725 DVSS.n15903 DVSS.n15881 4.5005
R17726 DVSS.n15896 DVSS.n15881 4.5005
R17727 DVSS.n15904 DVSS.n15881 4.5005
R17728 DVSS.n15895 DVSS.n15881 4.5005
R17729 DVSS.n15905 DVSS.n15881 4.5005
R17730 DVSS.n15894 DVSS.n15881 4.5005
R17731 DVSS.n15907 DVSS.n15881 4.5005
R17732 DVSS.n15893 DVSS.n15881 4.5005
R17733 DVSS.n17821 DVSS.n15881 4.5005
R17734 DVSS.n15891 DVSS.n15881 4.5005
R17735 DVSS.n17823 DVSS.n15881 4.5005
R17736 DVSS.n15900 DVSS.n15886 4.5005
R17737 DVSS.n15898 DVSS.n15886 4.5005
R17738 DVSS.n15902 DVSS.n15886 4.5005
R17739 DVSS.n15897 DVSS.n15886 4.5005
R17740 DVSS.n15903 DVSS.n15886 4.5005
R17741 DVSS.n15896 DVSS.n15886 4.5005
R17742 DVSS.n15904 DVSS.n15886 4.5005
R17743 DVSS.n15895 DVSS.n15886 4.5005
R17744 DVSS.n15905 DVSS.n15886 4.5005
R17745 DVSS.n15894 DVSS.n15886 4.5005
R17746 DVSS.n15907 DVSS.n15886 4.5005
R17747 DVSS.n15893 DVSS.n15886 4.5005
R17748 DVSS.n17821 DVSS.n15886 4.5005
R17749 DVSS.n17823 DVSS.n15886 4.5005
R17750 DVSS.n15900 DVSS.n15880 4.5005
R17751 DVSS.n15898 DVSS.n15880 4.5005
R17752 DVSS.n15902 DVSS.n15880 4.5005
R17753 DVSS.n15897 DVSS.n15880 4.5005
R17754 DVSS.n15903 DVSS.n15880 4.5005
R17755 DVSS.n15896 DVSS.n15880 4.5005
R17756 DVSS.n15904 DVSS.n15880 4.5005
R17757 DVSS.n15895 DVSS.n15880 4.5005
R17758 DVSS.n15905 DVSS.n15880 4.5005
R17759 DVSS.n15894 DVSS.n15880 4.5005
R17760 DVSS.n15907 DVSS.n15880 4.5005
R17761 DVSS.n17821 DVSS.n15880 4.5005
R17762 DVSS.n17823 DVSS.n15880 4.5005
R17763 DVSS.n15900 DVSS.n15887 4.5005
R17764 DVSS.n15898 DVSS.n15887 4.5005
R17765 DVSS.n15902 DVSS.n15887 4.5005
R17766 DVSS.n15897 DVSS.n15887 4.5005
R17767 DVSS.n15903 DVSS.n15887 4.5005
R17768 DVSS.n15896 DVSS.n15887 4.5005
R17769 DVSS.n15904 DVSS.n15887 4.5005
R17770 DVSS.n15895 DVSS.n15887 4.5005
R17771 DVSS.n15905 DVSS.n15887 4.5005
R17772 DVSS.n15894 DVSS.n15887 4.5005
R17773 DVSS.n15907 DVSS.n15887 4.5005
R17774 DVSS.n17821 DVSS.n15887 4.5005
R17775 DVSS.n17823 DVSS.n15887 4.5005
R17776 DVSS.n15900 DVSS.n15879 4.5005
R17777 DVSS.n15898 DVSS.n15879 4.5005
R17778 DVSS.n15902 DVSS.n15879 4.5005
R17779 DVSS.n15897 DVSS.n15879 4.5005
R17780 DVSS.n15903 DVSS.n15879 4.5005
R17781 DVSS.n15896 DVSS.n15879 4.5005
R17782 DVSS.n15904 DVSS.n15879 4.5005
R17783 DVSS.n15895 DVSS.n15879 4.5005
R17784 DVSS.n15905 DVSS.n15879 4.5005
R17785 DVSS.n15894 DVSS.n15879 4.5005
R17786 DVSS.n15907 DVSS.n15879 4.5005
R17787 DVSS.n15893 DVSS.n15879 4.5005
R17788 DVSS.n17821 DVSS.n15879 4.5005
R17789 DVSS.n17823 DVSS.n15879 4.5005
R17790 DVSS.n17822 DVSS.n15900 4.5005
R17791 DVSS.n17822 DVSS.n15898 4.5005
R17792 DVSS.n17822 DVSS.n15902 4.5005
R17793 DVSS.n17822 DVSS.n15897 4.5005
R17794 DVSS.n17822 DVSS.n15903 4.5005
R17795 DVSS.n17822 DVSS.n15896 4.5005
R17796 DVSS.n17822 DVSS.n15904 4.5005
R17797 DVSS.n17822 DVSS.n15895 4.5005
R17798 DVSS.n17822 DVSS.n15905 4.5005
R17799 DVSS.n17822 DVSS.n15894 4.5005
R17800 DVSS.n17822 DVSS.n15907 4.5005
R17801 DVSS.n17822 DVSS.n15893 4.5005
R17802 DVSS.n17822 DVSS.n17821 4.5005
R17803 DVSS.n17822 DVSS.n15891 4.5005
R17804 DVSS.n17823 DVSS.n17822 4.5005
R17805 DVSS.n16551 DVSS.n16343 4.5005
R17806 DVSS.n16353 DVSS.n16343 4.5005
R17807 DVSS.n16553 DVSS.n16343 4.5005
R17808 DVSS.n16352 DVSS.n16343 4.5005
R17809 DVSS.n16554 DVSS.n16343 4.5005
R17810 DVSS.n16351 DVSS.n16343 4.5005
R17811 DVSS.n16555 DVSS.n16343 4.5005
R17812 DVSS.n16350 DVSS.n16343 4.5005
R17813 DVSS.n16556 DVSS.n16343 4.5005
R17814 DVSS.n16349 DVSS.n16343 4.5005
R17815 DVSS.n16558 DVSS.n16343 4.5005
R17816 DVSS.n16348 DVSS.n16343 4.5005
R17817 DVSS.n16595 DVSS.n16343 4.5005
R17818 DVSS.n16346 DVSS.n16343 4.5005
R17819 DVSS.n16597 DVSS.n16343 4.5005
R17820 DVSS.n16551 DVSS.n16335 4.5005
R17821 DVSS.n16353 DVSS.n16335 4.5005
R17822 DVSS.n16553 DVSS.n16335 4.5005
R17823 DVSS.n16352 DVSS.n16335 4.5005
R17824 DVSS.n16554 DVSS.n16335 4.5005
R17825 DVSS.n16351 DVSS.n16335 4.5005
R17826 DVSS.n16555 DVSS.n16335 4.5005
R17827 DVSS.n16350 DVSS.n16335 4.5005
R17828 DVSS.n16556 DVSS.n16335 4.5005
R17829 DVSS.n16349 DVSS.n16335 4.5005
R17830 DVSS.n16558 DVSS.n16335 4.5005
R17831 DVSS.n16348 DVSS.n16335 4.5005
R17832 DVSS.n16595 DVSS.n16335 4.5005
R17833 DVSS.n16346 DVSS.n16335 4.5005
R17834 DVSS.n16597 DVSS.n16335 4.5005
R17835 DVSS.n16596 DVSS.n16551 4.5005
R17836 DVSS.n16596 DVSS.n16353 4.5005
R17837 DVSS.n16596 DVSS.n16553 4.5005
R17838 DVSS.n16596 DVSS.n16352 4.5005
R17839 DVSS.n16596 DVSS.n16554 4.5005
R17840 DVSS.n16596 DVSS.n16351 4.5005
R17841 DVSS.n16596 DVSS.n16555 4.5005
R17842 DVSS.n16596 DVSS.n16350 4.5005
R17843 DVSS.n16596 DVSS.n16556 4.5005
R17844 DVSS.n16596 DVSS.n16349 4.5005
R17845 DVSS.n16596 DVSS.n16558 4.5005
R17846 DVSS.n16596 DVSS.n16348 4.5005
R17847 DVSS.n16596 DVSS.n16595 4.5005
R17848 DVSS.n16596 DVSS.n16346 4.5005
R17849 DVSS.n16597 DVSS.n16596 4.5005
R17850 DVSS.n19312 DVSS.n19311 4.5005
R17851 DVSS.n19313 DVSS.n19312 4.5005
R17852 DVSS.n19314 DVSS.n19313 4.5005
R17853 DVSS.n19899 DVSS.n19898 4.5005
R17854 DVSS.n19900 DVSS.n19899 4.5005
R17855 DVSS.n19247 DVSS.n19041 4.5005
R17856 DVSS.n19250 DVSS.n19041 4.5005
R17857 DVSS.n19621 DVSS.n19159 4.5005
R17858 DVSS.n19624 DVSS.n19159 4.5005
R17859 DVSS.n19029 DVSS.n19012 4.5005
R17860 DVSS.n19898 DVSS.n19029 4.5005
R17861 DVSS.n19900 DVSS.n19029 4.5005
R17862 DVSS.n19171 DVSS.n19030 4.5005
R17863 DVSS.n19247 DVSS.n19171 4.5005
R17864 DVSS.n19250 DVSS.n19171 4.5005
R17865 DVSS.n19598 DVSS.n19157 4.5005
R17866 DVSS.n19621 DVSS.n19157 4.5005
R17867 DVSS.n19624 DVSS.n19157 4.5005
R17868 DVSS.n19901 DVSS.n19012 4.5005
R17869 DVSS.n19901 DVSS.n19011 4.5005
R17870 DVSS.n19901 DVSS.n19013 4.5005
R17871 DVSS.n19901 DVSS.n19010 4.5005
R17872 DVSS.n19901 DVSS.n19014 4.5005
R17873 DVSS.n19901 DVSS.n19009 4.5005
R17874 DVSS.n19901 DVSS.n19015 4.5005
R17875 DVSS.n19901 DVSS.n19008 4.5005
R17876 DVSS.n19901 DVSS.n19016 4.5005
R17877 DVSS.n19901 DVSS.n19007 4.5005
R17878 DVSS.n19901 DVSS.n19017 4.5005
R17879 DVSS.n19901 DVSS.n19006 4.5005
R17880 DVSS.n19901 DVSS.n19018 4.5005
R17881 DVSS.n19901 DVSS.n19005 4.5005
R17882 DVSS.n19901 DVSS.n19019 4.5005
R17883 DVSS.n19901 DVSS.n19900 4.5005
R17884 DVSS.n19249 DVSS.n19030 4.5005
R17885 DVSS.n19249 DVSS.n19224 4.5005
R17886 DVSS.n19249 DVSS.n19227 4.5005
R17887 DVSS.n19249 DVSS.n19222 4.5005
R17888 DVSS.n19249 DVSS.n19230 4.5005
R17889 DVSS.n19249 DVSS.n19221 4.5005
R17890 DVSS.n19249 DVSS.n19233 4.5005
R17891 DVSS.n19249 DVSS.n19220 4.5005
R17892 DVSS.n19249 DVSS.n19236 4.5005
R17893 DVSS.n19249 DVSS.n19219 4.5005
R17894 DVSS.n19249 DVSS.n19239 4.5005
R17895 DVSS.n19249 DVSS.n19218 4.5005
R17896 DVSS.n19249 DVSS.n19242 4.5005
R17897 DVSS.n19249 DVSS.n19217 4.5005
R17898 DVSS.n19249 DVSS.n19244 4.5005
R17899 DVSS.n19250 DVSS.n19249 4.5005
R17900 DVSS.n19623 DVSS.n19598 4.5005
R17901 DVSS.n19623 DVSS.n19168 4.5005
R17902 DVSS.n19623 DVSS.n19601 4.5005
R17903 DVSS.n19623 DVSS.n19167 4.5005
R17904 DVSS.n19623 DVSS.n19604 4.5005
R17905 DVSS.n19623 DVSS.n19166 4.5005
R17906 DVSS.n19623 DVSS.n19607 4.5005
R17907 DVSS.n19623 DVSS.n19165 4.5005
R17908 DVSS.n19623 DVSS.n19610 4.5005
R17909 DVSS.n19623 DVSS.n19164 4.5005
R17910 DVSS.n19623 DVSS.n19613 4.5005
R17911 DVSS.n19623 DVSS.n19163 4.5005
R17912 DVSS.n19623 DVSS.n19616 4.5005
R17913 DVSS.n19623 DVSS.n19162 4.5005
R17914 DVSS.n19623 DVSS.n19618 4.5005
R17915 DVSS.n19624 DVSS.n19623 4.5005
R17916 DVSS.n22433 DVSS.n22432 4.5005
R17917 DVSS.n22430 DVSS.n1012 4.5005
R17918 DVSS.n22431 DVSS.n22430 4.5005
R17919 DVSS.n22431 DVSS.n22429 4.5005
R17920 DVSS.n22432 DVSS.n22431 4.5005
R17921 DVSS.n22383 DVSS.n22382 4.5005
R17922 DVSS.n22384 DVSS.n22383 4.5005
R17923 DVSS.n22369 DVSS.n22368 4.5005
R17924 DVSS.n22370 DVSS.n22369 4.5005
R17925 DVSS.n13086 DVSS.n12961 4.5005
R17926 DVSS.n13089 DVSS.n12961 4.5005
R17927 DVSS.n22386 DVSS.n1015 4.5005
R17928 DVSS.n22384 DVSS.n1015 4.5005
R17929 DVSS.n22371 DVSS.n1043 4.5005
R17930 DVSS.n22371 DVSS.n22370 4.5005
R17931 DVSS.n12959 DVSS.n1175 4.5005
R17932 DVSS.n13089 DVSS.n12959 4.5005
R17933 DVSS.n22386 DVSS.n22385 4.5005
R17934 DVSS.n22385 DVSS.n1025 4.5005
R17935 DVSS.n22385 DVSS.n1028 4.5005
R17936 DVSS.n22385 DVSS.n1024 4.5005
R17937 DVSS.n22385 DVSS.n1030 4.5005
R17938 DVSS.n22385 DVSS.n1023 4.5005
R17939 DVSS.n22385 DVSS.n1032 4.5005
R17940 DVSS.n22385 DVSS.n1022 4.5005
R17941 DVSS.n22385 DVSS.n1034 4.5005
R17942 DVSS.n22385 DVSS.n1021 4.5005
R17943 DVSS.n22385 DVSS.n1036 4.5005
R17944 DVSS.n22385 DVSS.n1020 4.5005
R17945 DVSS.n22385 DVSS.n1038 4.5005
R17946 DVSS.n22385 DVSS.n1019 4.5005
R17947 DVSS.n22385 DVSS.n1040 4.5005
R17948 DVSS.n22385 DVSS.n1018 4.5005
R17949 DVSS.n22385 DVSS.n22384 4.5005
R17950 DVSS.n1153 DVSS.n1043 4.5005
R17951 DVSS.n22365 DVSS.n1153 4.5005
R17952 DVSS.n22363 DVSS.n1153 4.5005
R17953 DVSS.n22362 DVSS.n1153 4.5005
R17954 DVSS.n22360 DVSS.n1153 4.5005
R17955 DVSS.n22359 DVSS.n1153 4.5005
R17956 DVSS.n22357 DVSS.n1153 4.5005
R17957 DVSS.n22356 DVSS.n1153 4.5005
R17958 DVSS.n22354 DVSS.n1153 4.5005
R17959 DVSS.n22353 DVSS.n1153 4.5005
R17960 DVSS.n22351 DVSS.n1153 4.5005
R17961 DVSS.n22350 DVSS.n1153 4.5005
R17962 DVSS.n22348 DVSS.n1153 4.5005
R17963 DVSS.n22347 DVSS.n1153 4.5005
R17964 DVSS.n22345 DVSS.n1153 4.5005
R17965 DVSS.n22344 DVSS.n1153 4.5005
R17966 DVSS.n22370 DVSS.n1153 4.5005
R17967 DVSS.n13088 DVSS.n1175 4.5005
R17968 DVSS.n13088 DVSS.n12971 4.5005
R17969 DVSS.n13088 DVSS.n13066 4.5005
R17970 DVSS.n13088 DVSS.n12969 4.5005
R17971 DVSS.n13088 DVSS.n13069 4.5005
R17972 DVSS.n13088 DVSS.n12968 4.5005
R17973 DVSS.n13088 DVSS.n13072 4.5005
R17974 DVSS.n13088 DVSS.n12967 4.5005
R17975 DVSS.n13088 DVSS.n13075 4.5005
R17976 DVSS.n13088 DVSS.n12966 4.5005
R17977 DVSS.n13088 DVSS.n13078 4.5005
R17978 DVSS.n13088 DVSS.n12965 4.5005
R17979 DVSS.n13088 DVSS.n13081 4.5005
R17980 DVSS.n13088 DVSS.n12964 4.5005
R17981 DVSS.n13088 DVSS.n13084 4.5005
R17982 DVSS.n13088 DVSS.n12963 4.5005
R17983 DVSS.n13089 DVSS.n13088 4.5005
R17984 DVSS.n13093 DVSS.n12957 4.5005
R17985 DVSS.n13094 DVSS.n13093 4.5005
R17986 DVSS.n12955 DVSS.n369 4.5005
R17987 DVSS.n12953 DVSS.n369 4.5005
R17988 DVSS.n12951 DVSS.n369 4.5005
R17989 DVSS.n12949 DVSS.n369 4.5005
R17990 DVSS.n12947 DVSS.n369 4.5005
R17991 DVSS.n12945 DVSS.n369 4.5005
R17992 DVSS.n12943 DVSS.n369 4.5005
R17993 DVSS.n12941 DVSS.n369 4.5005
R17994 DVSS.n12939 DVSS.n369 4.5005
R17995 DVSS.n12937 DVSS.n369 4.5005
R17996 DVSS.n12935 DVSS.n369 4.5005
R17997 DVSS.n12933 DVSS.n369 4.5005
R17998 DVSS.n12931 DVSS.n369 4.5005
R17999 DVSS.n12929 DVSS.n369 4.5005
R18000 DVSS.n12927 DVSS.n369 4.5005
R18001 DVSS.n12925 DVSS.n369 4.5005
R18002 DVSS.n13094 DVSS.n369 4.5005
R18003 DVSS.n19649 DVSS.n19146 4.5005
R18004 DVSS.n19652 DVSS.n19146 4.5005
R18005 DVSS.n19626 DVSS.n19142 4.5005
R18006 DVSS.n19649 DVSS.n19142 4.5005
R18007 DVSS.n19652 DVSS.n19142 4.5005
R18008 DVSS.n19651 DVSS.n19626 4.5005
R18009 DVSS.n19651 DVSS.n19155 4.5005
R18010 DVSS.n19651 DVSS.n19629 4.5005
R18011 DVSS.n19651 DVSS.n19154 4.5005
R18012 DVSS.n19651 DVSS.n19632 4.5005
R18013 DVSS.n19651 DVSS.n19153 4.5005
R18014 DVSS.n19651 DVSS.n19635 4.5005
R18015 DVSS.n19651 DVSS.n19152 4.5005
R18016 DVSS.n19651 DVSS.n19638 4.5005
R18017 DVSS.n19651 DVSS.n19151 4.5005
R18018 DVSS.n19651 DVSS.n19641 4.5005
R18019 DVSS.n19651 DVSS.n19150 4.5005
R18020 DVSS.n19651 DVSS.n19644 4.5005
R18021 DVSS.n19651 DVSS.n19149 4.5005
R18022 DVSS.n19651 DVSS.n19646 4.5005
R18023 DVSS.n19652 DVSS.n19651 4.5005
R18024 DVSS.n1218 DVSS.n1217 4.5005
R18025 DVSS.n22335 DVSS.n1218 4.5005
R18026 DVSS.n1271 DVSS.n523 4.5005
R18027 DVSS.n19109 DVSS.n19108 4.5005
R18028 DVSS.n19846 DVSS.n19109 4.5005
R18029 DVSS.n19848 DVSS.n19847 4.5005
R18030 DVSS.n19847 DVSS.n19846 4.5005
R18031 DVSS.n1291 DVSS.n507 4.5005
R18032 DVSS.n22337 DVSS.n22336 4.5005
R18033 DVSS.n22336 DVSS.n22335 4.5005
R18034 DVSS.n20632 DVSS.n14668 4.5005
R18035 DVSS.n14669 DVSS.n14668 4.5005
R18036 DVSS.n20397 DVSS.n14668 4.5005
R18037 DVSS.n20399 DVSS.n14668 4.5005
R18038 DVSS.n20401 DVSS.n14668 4.5005
R18039 DVSS.n20376 DVSS.n14668 4.5005
R18040 DVSS.n20413 DVSS.n14668 4.5005
R18041 DVSS.n20415 DVSS.n14668 4.5005
R18042 DVSS.n20417 DVSS.n14668 4.5005
R18043 DVSS.n20359 DVSS.n14668 4.5005
R18044 DVSS.n20429 DVSS.n14668 4.5005
R18045 DVSS.n20431 DVSS.n14668 4.5005
R18046 DVSS.n20341 DVSS.n14668 4.5005
R18047 DVSS.n20446 DVSS.n14668 4.5005
R18048 DVSS.n20448 DVSS.n14668 4.5005
R18049 DVSS.n14702 DVSS.n14668 4.5005
R18050 DVSS.n20627 DVSS.n14180 4.5005
R18051 DVSS.n14686 DVSS.n14180 4.5005
R18052 DVSS.n14685 DVSS.n14180 4.5005
R18053 DVSS.n14687 DVSS.n14180 4.5005
R18054 DVSS.n14684 DVSS.n14180 4.5005
R18055 DVSS.n14688 DVSS.n14180 4.5005
R18056 DVSS.n14683 DVSS.n14180 4.5005
R18057 DVSS.n14689 DVSS.n14180 4.5005
R18058 DVSS.n14682 DVSS.n14180 4.5005
R18059 DVSS.n14690 DVSS.n14180 4.5005
R18060 DVSS.n14681 DVSS.n14180 4.5005
R18061 DVSS.n14691 DVSS.n14180 4.5005
R18062 DVSS.n14680 DVSS.n14180 4.5005
R18063 DVSS.n14692 DVSS.n14180 4.5005
R18064 DVSS.n20337 DVSS.n14180 4.5005
R18065 DVSS.n20625 DVSS.n14180 4.5005
R18066 DVSS.n20627 DVSS.n14677 4.5005
R18067 DVSS.n14686 DVSS.n14677 4.5005
R18068 DVSS.n14685 DVSS.n14677 4.5005
R18069 DVSS.n14687 DVSS.n14677 4.5005
R18070 DVSS.n14684 DVSS.n14677 4.5005
R18071 DVSS.n14688 DVSS.n14677 4.5005
R18072 DVSS.n14683 DVSS.n14677 4.5005
R18073 DVSS.n14689 DVSS.n14677 4.5005
R18074 DVSS.n14682 DVSS.n14677 4.5005
R18075 DVSS.n14690 DVSS.n14677 4.5005
R18076 DVSS.n14681 DVSS.n14677 4.5005
R18077 DVSS.n14691 DVSS.n14677 4.5005
R18078 DVSS.n14680 DVSS.n14677 4.5005
R18079 DVSS.n14692 DVSS.n14677 4.5005
R18080 DVSS.n20337 DVSS.n14677 4.5005
R18081 DVSS.n20625 DVSS.n14677 4.5005
R18082 DVSS.n20627 DVSS.n14675 4.5005
R18083 DVSS.n14686 DVSS.n14675 4.5005
R18084 DVSS.n14685 DVSS.n14675 4.5005
R18085 DVSS.n14687 DVSS.n14675 4.5005
R18086 DVSS.n14684 DVSS.n14675 4.5005
R18087 DVSS.n14688 DVSS.n14675 4.5005
R18088 DVSS.n14683 DVSS.n14675 4.5005
R18089 DVSS.n14689 DVSS.n14675 4.5005
R18090 DVSS.n14682 DVSS.n14675 4.5005
R18091 DVSS.n14690 DVSS.n14675 4.5005
R18092 DVSS.n14681 DVSS.n14675 4.5005
R18093 DVSS.n14691 DVSS.n14675 4.5005
R18094 DVSS.n14680 DVSS.n14675 4.5005
R18095 DVSS.n14692 DVSS.n14675 4.5005
R18096 DVSS.n20337 DVSS.n14675 4.5005
R18097 DVSS.n20625 DVSS.n14675 4.5005
R18098 DVSS.n20325 DVSS.n14376 4.5005
R18099 DVSS.n14862 DVSS.n14376 4.5005
R18100 DVSS.n20326 DVSS.n14376 4.5005
R18101 DVSS.n14861 DVSS.n14376 4.5005
R18102 DVSS.n20327 DVSS.n14376 4.5005
R18103 DVSS.n14860 DVSS.n14376 4.5005
R18104 DVSS.n20328 DVSS.n14376 4.5005
R18105 DVSS.n14859 DVSS.n14376 4.5005
R18106 DVSS.n20329 DVSS.n14376 4.5005
R18107 DVSS.n14858 DVSS.n14376 4.5005
R18108 DVSS.n20330 DVSS.n14376 4.5005
R18109 DVSS.n20362 DVSS.n14376 4.5005
R18110 DVSS.n20331 DVSS.n14376 4.5005
R18111 DVSS.n14855 DVSS.n14376 4.5005
R18112 DVSS.n20457 DVSS.n14376 4.5005
R18113 DVSS.n20459 DVSS.n14376 4.5005
R18114 DVSS.n20458 DVSS.n20325 4.5005
R18115 DVSS.n20458 DVSS.n14862 4.5005
R18116 DVSS.n20458 DVSS.n20326 4.5005
R18117 DVSS.n20458 DVSS.n14861 4.5005
R18118 DVSS.n20458 DVSS.n20327 4.5005
R18119 DVSS.n20458 DVSS.n14860 4.5005
R18120 DVSS.n20458 DVSS.n20328 4.5005
R18121 DVSS.n20458 DVSS.n14859 4.5005
R18122 DVSS.n20458 DVSS.n20329 4.5005
R18123 DVSS.n20458 DVSS.n14858 4.5005
R18124 DVSS.n20458 DVSS.n20330 4.5005
R18125 DVSS.n20458 DVSS.n14856 4.5005
R18126 DVSS.n20458 DVSS.n20331 4.5005
R18127 DVSS.n20458 DVSS.n14855 4.5005
R18128 DVSS.n20458 DVSS.n20457 4.5005
R18129 DVSS.n20459 DVSS.n20458 4.5005
R18130 DVSS.n20627 DVSS.n20626 4.5005
R18131 DVSS.n20626 DVSS.n14686 4.5005
R18132 DVSS.n20626 DVSS.n14685 4.5005
R18133 DVSS.n20626 DVSS.n14687 4.5005
R18134 DVSS.n20626 DVSS.n14684 4.5005
R18135 DVSS.n20626 DVSS.n14688 4.5005
R18136 DVSS.n20626 DVSS.n14683 4.5005
R18137 DVSS.n20626 DVSS.n14689 4.5005
R18138 DVSS.n20626 DVSS.n14682 4.5005
R18139 DVSS.n20626 DVSS.n14690 4.5005
R18140 DVSS.n20626 DVSS.n14681 4.5005
R18141 DVSS.n20626 DVSS.n14691 4.5005
R18142 DVSS.n20626 DVSS.n14680 4.5005
R18143 DVSS.n20626 DVSS.n14692 4.5005
R18144 DVSS.n20626 DVSS.n20625 4.5005
R18145 DVSS.n20627 DVSS.n14674 4.5005
R18146 DVSS.n14686 DVSS.n14674 4.5005
R18147 DVSS.n14685 DVSS.n14674 4.5005
R18148 DVSS.n14687 DVSS.n14674 4.5005
R18149 DVSS.n14684 DVSS.n14674 4.5005
R18150 DVSS.n14688 DVSS.n14674 4.5005
R18151 DVSS.n14683 DVSS.n14674 4.5005
R18152 DVSS.n14689 DVSS.n14674 4.5005
R18153 DVSS.n14682 DVSS.n14674 4.5005
R18154 DVSS.n14690 DVSS.n14674 4.5005
R18155 DVSS.n14681 DVSS.n14674 4.5005
R18156 DVSS.n14691 DVSS.n14674 4.5005
R18157 DVSS.n14692 DVSS.n14674 4.5005
R18158 DVSS.n20625 DVSS.n14674 4.5005
R18159 DVSS.n20627 DVSS.n14150 4.5005
R18160 DVSS.n14686 DVSS.n14150 4.5005
R18161 DVSS.n14685 DVSS.n14150 4.5005
R18162 DVSS.n14687 DVSS.n14150 4.5005
R18163 DVSS.n14684 DVSS.n14150 4.5005
R18164 DVSS.n14688 DVSS.n14150 4.5005
R18165 DVSS.n14683 DVSS.n14150 4.5005
R18166 DVSS.n14689 DVSS.n14150 4.5005
R18167 DVSS.n14682 DVSS.n14150 4.5005
R18168 DVSS.n14690 DVSS.n14150 4.5005
R18169 DVSS.n14681 DVSS.n14150 4.5005
R18170 DVSS.n14691 DVSS.n14150 4.5005
R18171 DVSS.n14692 DVSS.n14150 4.5005
R18172 DVSS.n20337 DVSS.n14150 4.5005
R18173 DVSS.n20625 DVSS.n14150 4.5005
R18174 DVSS.n20632 DVSS.n13430 4.5005
R18175 DVSS.n14669 DVSS.n13430 4.5005
R18176 DVSS.n20397 DVSS.n13430 4.5005
R18177 DVSS.n20399 DVSS.n13430 4.5005
R18178 DVSS.n20401 DVSS.n13430 4.5005
R18179 DVSS.n20376 DVSS.n13430 4.5005
R18180 DVSS.n20413 DVSS.n13430 4.5005
R18181 DVSS.n20415 DVSS.n13430 4.5005
R18182 DVSS.n20417 DVSS.n13430 4.5005
R18183 DVSS.n20359 DVSS.n13430 4.5005
R18184 DVSS.n20429 DVSS.n13430 4.5005
R18185 DVSS.n20357 DVSS.n13430 4.5005
R18186 DVSS.n20341 DVSS.n13430 4.5005
R18187 DVSS.n20446 DVSS.n13430 4.5005
R18188 DVSS.n20448 DVSS.n13430 4.5005
R18189 DVSS.n14702 DVSS.n13430 4.5005
R18190 DVSS.n17456 DVSS.n17433 4.5005
R18191 DVSS.n17530 DVSS.n16920 4.5005
R18192 DVSS.n17529 DVSS.n16900 4.5005
R18193 DVSS.n16978 DVSS.n15452 4.5005
R18194 DVSS.n16980 DVSS.n15452 4.5005
R18195 DVSS.n16994 DVSS.n15452 4.5005
R18196 DVSS.n17494 DVSS.n16936 4.5005
R18197 DVSS.n17502 DVSS.n16938 4.5005
R18198 DVSS.n17424 DVSS.n17209 4.5005
R18199 DVSS.n17423 DVSS.n17418 4.5005
R18200 DVSS.n17423 DVSS.n17420 4.5005
R18201 DVSS.n17425 DVSS.n17206 4.5005
R18202 DVSS.n17433 DVSS.n17426 4.5005
R18203 DVSS.n17452 DVSS.n17451 4.5005
R18204 DVSS.n17455 DVSS.n17452 4.5005
R18205 DVSS.n17452 DVSS.n17433 4.5005
R18206 DVSS.n17457 DVSS.n17426 4.5005
R18207 DVSS.n17425 DVSS.n17424 4.5005
R18208 DVSS.n17424 DVSS.n17423 4.5005
R18209 DVSS.n17421 DVSS.n17209 4.5005
R18210 DVSS.n17420 DVSS.n17209 4.5005
R18211 DVSS.n17212 DVSS.n17209 4.5005
R18212 DVSS.n17211 DVSS.n17209 4.5005
R18213 DVSS.n17215 DVSS.n17209 4.5005
R18214 DVSS.n17214 DVSS.n17209 4.5005
R18215 DVSS.n17218 DVSS.n17209 4.5005
R18216 DVSS.n17217 DVSS.n17209 4.5005
R18217 DVSS.n17221 DVSS.n17209 4.5005
R18218 DVSS.n17220 DVSS.n17209 4.5005
R18219 DVSS.n17418 DVSS.n17209 4.5005
R18220 DVSS.n17521 DVSS.n16938 4.5005
R18221 DVSS.n17521 DVSS.n16936 4.5005
R18222 DVSS.n17520 DVSS.n17504 4.5005
R18223 DVSS.n17520 DVSS.n17499 4.5005
R18224 DVSS.n17520 DVSS.n17507 4.5005
R18225 DVSS.n17520 DVSS.n17498 4.5005
R18226 DVSS.n17520 DVSS.n17510 4.5005
R18227 DVSS.n17520 DVSS.n17497 4.5005
R18228 DVSS.n17520 DVSS.n17513 4.5005
R18229 DVSS.n17520 DVSS.n17496 4.5005
R18230 DVSS.n17520 DVSS.n17516 4.5005
R18231 DVSS.n17520 DVSS.n17495 4.5005
R18232 DVSS.n17520 DVSS.n17519 4.5005
R18233 DVSS.n17520 DVSS.n17494 4.5005
R18234 DVSS.n17521 DVSS.n17520 4.5005
R18235 DVSS.n17530 DVSS.n16909 4.5005
R18236 DVSS.n16978 DVSS.n15443 4.5005
R18237 DVSS.n17530 DVSS.n17529 4.5005
R18238 DVSS.n17457 DVSS.n17456 4.5005
R18239 DVSS.n17456 DVSS.n17432 4.5005
R18240 DVSS.n17456 DVSS.n17436 4.5005
R18241 DVSS.n17456 DVSS.n17431 4.5005
R18242 DVSS.n17456 DVSS.n17438 4.5005
R18243 DVSS.n17456 DVSS.n17430 4.5005
R18244 DVSS.n17456 DVSS.n17440 4.5005
R18245 DVSS.n17456 DVSS.n17429 4.5005
R18246 DVSS.n17456 DVSS.n17442 4.5005
R18247 DVSS.n17456 DVSS.n17428 4.5005
R18248 DVSS.n17456 DVSS.n17455 4.5005
R18249 DVSS.n18087 DVSS.n15629 4.5005
R18250 DVSS.n18089 DVSS.n15629 4.5005
R18251 DVSS.n18089 DVSS.n18088 4.5005
R18252 DVSS.n18088 DVSS.n15637 4.5005
R18253 DVSS.n18088 DVSS.n15634 4.5005
R18254 DVSS.n18088 DVSS.n15639 4.5005
R18255 DVSS.n18088 DVSS.n15633 4.5005
R18256 DVSS.n18088 DVSS.n15641 4.5005
R18257 DVSS.n18088 DVSS.n15632 4.5005
R18258 DVSS.n18088 DVSS.n15643 4.5005
R18259 DVSS.n18088 DVSS.n15631 4.5005
R18260 DVSS.n18088 DVSS.n18087 4.5005
R18261 DVSS.n21382 DVSS.n13425 4.5005
R18262 DVSS.n13425 DVSS.n13419 4.5005
R18263 DVSS.n21384 DVSS.n13425 4.5005
R18264 DVSS.n13424 DVSS.n13419 4.5005
R18265 DVSS.n21384 DVSS.n13424 4.5005
R18266 DVSS.n13436 DVSS.n13426 4.5005
R18267 DVSS.n13426 DVSS.n13419 4.5005
R18268 DVSS.n21384 DVSS.n13426 4.5005
R18269 DVSS.n13436 DVSS.n13423 4.5005
R18270 DVSS.n13423 DVSS.n13419 4.5005
R18271 DVSS.n21384 DVSS.n13423 4.5005
R18272 DVSS.n13427 DVSS.n13419 4.5005
R18273 DVSS.n21384 DVSS.n13427 4.5005
R18274 DVSS.n13422 DVSS.n13419 4.5005
R18275 DVSS.n21384 DVSS.n13422 4.5005
R18276 DVSS.n13428 DVSS.n13419 4.5005
R18277 DVSS.n21384 DVSS.n13428 4.5005
R18278 DVSS.n13421 DVSS.n13419 4.5005
R18279 DVSS.n21384 DVSS.n13421 4.5005
R18280 DVSS.n13429 DVSS.n13419 4.5005
R18281 DVSS.n21384 DVSS.n13429 4.5005
R18282 DVSS.n13442 DVSS.n13420 4.5005
R18283 DVSS.n13445 DVSS.n13420 4.5005
R18284 DVSS.n13440 DVSS.n13420 4.5005
R18285 DVSS.n13446 DVSS.n13420 4.5005
R18286 DVSS.n13439 DVSS.n13420 4.5005
R18287 DVSS.n13447 DVSS.n13420 4.5005
R18288 DVSS.n13438 DVSS.n13420 4.5005
R18289 DVSS.n13450 DVSS.n13420 4.5005
R18290 DVSS.n21382 DVSS.n13420 4.5005
R18291 DVSS.n21384 DVSS.n13420 4.5005
R18292 DVSS.n21383 DVSS.n13442 4.5005
R18293 DVSS.n21383 DVSS.n13444 4.5005
R18294 DVSS.n21383 DVSS.n13441 4.5005
R18295 DVSS.n21383 DVSS.n13445 4.5005
R18296 DVSS.n21383 DVSS.n13440 4.5005
R18297 DVSS.n21383 DVSS.n13446 4.5005
R18298 DVSS.n21383 DVSS.n13439 4.5005
R18299 DVSS.n21383 DVSS.n13447 4.5005
R18300 DVSS.n21383 DVSS.n13438 4.5005
R18301 DVSS.n21383 DVSS.n13449 4.5005
R18302 DVSS.n21383 DVSS.n13437 4.5005
R18303 DVSS.n21383 DVSS.n13450 4.5005
R18304 DVSS.n21383 DVSS.n13436 4.5005
R18305 DVSS.n21383 DVSS.n21382 4.5005
R18306 DVSS.n21384 DVSS.n21383 4.5005
R18307 DVSS.n21067 DVSS.n14137 4.5005
R18308 DVSS.n14183 DVSS.n14137 4.5005
R18309 DVSS.n14178 DVSS.n14137 4.5005
R18310 DVSS.n14184 DVSS.n14137 4.5005
R18311 DVSS.n14177 DVSS.n14137 4.5005
R18312 DVSS.n14185 DVSS.n14137 4.5005
R18313 DVSS.n14176 DVSS.n14137 4.5005
R18314 DVSS.n14188 DVSS.n14137 4.5005
R18315 DVSS.n14174 DVSS.n14137 4.5005
R18316 DVSS.n14189 DVSS.n14137 4.5005
R18317 DVSS.n21065 DVSS.n14137 4.5005
R18318 DVSS.n21067 DVSS.n14139 4.5005
R18319 DVSS.n14182 DVSS.n14139 4.5005
R18320 DVSS.n14179 DVSS.n14139 4.5005
R18321 DVSS.n14183 DVSS.n14139 4.5005
R18322 DVSS.n14178 DVSS.n14139 4.5005
R18323 DVSS.n14184 DVSS.n14139 4.5005
R18324 DVSS.n14177 DVSS.n14139 4.5005
R18325 DVSS.n14185 DVSS.n14139 4.5005
R18326 DVSS.n14176 DVSS.n14139 4.5005
R18327 DVSS.n14187 DVSS.n14139 4.5005
R18328 DVSS.n14175 DVSS.n14139 4.5005
R18329 DVSS.n14188 DVSS.n14139 4.5005
R18330 DVSS.n14189 DVSS.n14139 4.5005
R18331 DVSS.n21065 DVSS.n14139 4.5005
R18332 DVSS.n21067 DVSS.n14136 4.5005
R18333 DVSS.n14182 DVSS.n14136 4.5005
R18334 DVSS.n14179 DVSS.n14136 4.5005
R18335 DVSS.n14183 DVSS.n14136 4.5005
R18336 DVSS.n14178 DVSS.n14136 4.5005
R18337 DVSS.n14184 DVSS.n14136 4.5005
R18338 DVSS.n14177 DVSS.n14136 4.5005
R18339 DVSS.n14185 DVSS.n14136 4.5005
R18340 DVSS.n14176 DVSS.n14136 4.5005
R18341 DVSS.n14187 DVSS.n14136 4.5005
R18342 DVSS.n14175 DVSS.n14136 4.5005
R18343 DVSS.n14188 DVSS.n14136 4.5005
R18344 DVSS.n14189 DVSS.n14136 4.5005
R18345 DVSS.n21065 DVSS.n14136 4.5005
R18346 DVSS.n21067 DVSS.n14140 4.5005
R18347 DVSS.n14182 DVSS.n14140 4.5005
R18348 DVSS.n14179 DVSS.n14140 4.5005
R18349 DVSS.n14183 DVSS.n14140 4.5005
R18350 DVSS.n14178 DVSS.n14140 4.5005
R18351 DVSS.n14184 DVSS.n14140 4.5005
R18352 DVSS.n14177 DVSS.n14140 4.5005
R18353 DVSS.n14185 DVSS.n14140 4.5005
R18354 DVSS.n14176 DVSS.n14140 4.5005
R18355 DVSS.n14187 DVSS.n14140 4.5005
R18356 DVSS.n14175 DVSS.n14140 4.5005
R18357 DVSS.n14188 DVSS.n14140 4.5005
R18358 DVSS.n14189 DVSS.n14140 4.5005
R18359 DVSS.n21065 DVSS.n14140 4.5005
R18360 DVSS.n21067 DVSS.n14135 4.5005
R18361 DVSS.n14182 DVSS.n14135 4.5005
R18362 DVSS.n14179 DVSS.n14135 4.5005
R18363 DVSS.n14183 DVSS.n14135 4.5005
R18364 DVSS.n14178 DVSS.n14135 4.5005
R18365 DVSS.n14184 DVSS.n14135 4.5005
R18366 DVSS.n14177 DVSS.n14135 4.5005
R18367 DVSS.n14185 DVSS.n14135 4.5005
R18368 DVSS.n14176 DVSS.n14135 4.5005
R18369 DVSS.n14187 DVSS.n14135 4.5005
R18370 DVSS.n14175 DVSS.n14135 4.5005
R18371 DVSS.n14188 DVSS.n14135 4.5005
R18372 DVSS.n14189 DVSS.n14135 4.5005
R18373 DVSS.n21065 DVSS.n14135 4.5005
R18374 DVSS.n21067 DVSS.n14141 4.5005
R18375 DVSS.n14182 DVSS.n14141 4.5005
R18376 DVSS.n14179 DVSS.n14141 4.5005
R18377 DVSS.n14183 DVSS.n14141 4.5005
R18378 DVSS.n14178 DVSS.n14141 4.5005
R18379 DVSS.n14184 DVSS.n14141 4.5005
R18380 DVSS.n14177 DVSS.n14141 4.5005
R18381 DVSS.n14185 DVSS.n14141 4.5005
R18382 DVSS.n14176 DVSS.n14141 4.5005
R18383 DVSS.n14187 DVSS.n14141 4.5005
R18384 DVSS.n14175 DVSS.n14141 4.5005
R18385 DVSS.n14188 DVSS.n14141 4.5005
R18386 DVSS.n14189 DVSS.n14141 4.5005
R18387 DVSS.n21065 DVSS.n14141 4.5005
R18388 DVSS.n21067 DVSS.n14134 4.5005
R18389 DVSS.n14182 DVSS.n14134 4.5005
R18390 DVSS.n14179 DVSS.n14134 4.5005
R18391 DVSS.n14183 DVSS.n14134 4.5005
R18392 DVSS.n14178 DVSS.n14134 4.5005
R18393 DVSS.n14184 DVSS.n14134 4.5005
R18394 DVSS.n14177 DVSS.n14134 4.5005
R18395 DVSS.n14185 DVSS.n14134 4.5005
R18396 DVSS.n14176 DVSS.n14134 4.5005
R18397 DVSS.n14187 DVSS.n14134 4.5005
R18398 DVSS.n14175 DVSS.n14134 4.5005
R18399 DVSS.n14188 DVSS.n14134 4.5005
R18400 DVSS.n14189 DVSS.n14134 4.5005
R18401 DVSS.n21065 DVSS.n14134 4.5005
R18402 DVSS.n21067 DVSS.n14142 4.5005
R18403 DVSS.n14182 DVSS.n14142 4.5005
R18404 DVSS.n14179 DVSS.n14142 4.5005
R18405 DVSS.n14183 DVSS.n14142 4.5005
R18406 DVSS.n14178 DVSS.n14142 4.5005
R18407 DVSS.n14184 DVSS.n14142 4.5005
R18408 DVSS.n14177 DVSS.n14142 4.5005
R18409 DVSS.n14185 DVSS.n14142 4.5005
R18410 DVSS.n14176 DVSS.n14142 4.5005
R18411 DVSS.n14187 DVSS.n14142 4.5005
R18412 DVSS.n14175 DVSS.n14142 4.5005
R18413 DVSS.n14188 DVSS.n14142 4.5005
R18414 DVSS.n14189 DVSS.n14142 4.5005
R18415 DVSS.n21065 DVSS.n14142 4.5005
R18416 DVSS.n21067 DVSS.n14133 4.5005
R18417 DVSS.n14182 DVSS.n14133 4.5005
R18418 DVSS.n14179 DVSS.n14133 4.5005
R18419 DVSS.n14183 DVSS.n14133 4.5005
R18420 DVSS.n14178 DVSS.n14133 4.5005
R18421 DVSS.n14184 DVSS.n14133 4.5005
R18422 DVSS.n14177 DVSS.n14133 4.5005
R18423 DVSS.n14185 DVSS.n14133 4.5005
R18424 DVSS.n14176 DVSS.n14133 4.5005
R18425 DVSS.n14187 DVSS.n14133 4.5005
R18426 DVSS.n14175 DVSS.n14133 4.5005
R18427 DVSS.n14188 DVSS.n14133 4.5005
R18428 DVSS.n14189 DVSS.n14133 4.5005
R18429 DVSS.n21065 DVSS.n14133 4.5005
R18430 DVSS.n21067 DVSS.n14143 4.5005
R18431 DVSS.n14182 DVSS.n14143 4.5005
R18432 DVSS.n14179 DVSS.n14143 4.5005
R18433 DVSS.n14183 DVSS.n14143 4.5005
R18434 DVSS.n14178 DVSS.n14143 4.5005
R18435 DVSS.n14184 DVSS.n14143 4.5005
R18436 DVSS.n14177 DVSS.n14143 4.5005
R18437 DVSS.n14185 DVSS.n14143 4.5005
R18438 DVSS.n14176 DVSS.n14143 4.5005
R18439 DVSS.n14187 DVSS.n14143 4.5005
R18440 DVSS.n14175 DVSS.n14143 4.5005
R18441 DVSS.n14188 DVSS.n14143 4.5005
R18442 DVSS.n14189 DVSS.n14143 4.5005
R18443 DVSS.n21065 DVSS.n14143 4.5005
R18444 DVSS.n21067 DVSS.n14132 4.5005
R18445 DVSS.n14182 DVSS.n14132 4.5005
R18446 DVSS.n14179 DVSS.n14132 4.5005
R18447 DVSS.n14183 DVSS.n14132 4.5005
R18448 DVSS.n14178 DVSS.n14132 4.5005
R18449 DVSS.n14184 DVSS.n14132 4.5005
R18450 DVSS.n14177 DVSS.n14132 4.5005
R18451 DVSS.n14185 DVSS.n14132 4.5005
R18452 DVSS.n14176 DVSS.n14132 4.5005
R18453 DVSS.n14187 DVSS.n14132 4.5005
R18454 DVSS.n14175 DVSS.n14132 4.5005
R18455 DVSS.n14188 DVSS.n14132 4.5005
R18456 DVSS.n14189 DVSS.n14132 4.5005
R18457 DVSS.n21065 DVSS.n14132 4.5005
R18458 DVSS.n21067 DVSS.n14144 4.5005
R18459 DVSS.n14182 DVSS.n14144 4.5005
R18460 DVSS.n14179 DVSS.n14144 4.5005
R18461 DVSS.n14183 DVSS.n14144 4.5005
R18462 DVSS.n14178 DVSS.n14144 4.5005
R18463 DVSS.n14184 DVSS.n14144 4.5005
R18464 DVSS.n14177 DVSS.n14144 4.5005
R18465 DVSS.n14185 DVSS.n14144 4.5005
R18466 DVSS.n14176 DVSS.n14144 4.5005
R18467 DVSS.n14187 DVSS.n14144 4.5005
R18468 DVSS.n14175 DVSS.n14144 4.5005
R18469 DVSS.n14188 DVSS.n14144 4.5005
R18470 DVSS.n14189 DVSS.n14144 4.5005
R18471 DVSS.n21065 DVSS.n14144 4.5005
R18472 DVSS.n21067 DVSS.n14131 4.5005
R18473 DVSS.n14182 DVSS.n14131 4.5005
R18474 DVSS.n14179 DVSS.n14131 4.5005
R18475 DVSS.n14183 DVSS.n14131 4.5005
R18476 DVSS.n14178 DVSS.n14131 4.5005
R18477 DVSS.n14184 DVSS.n14131 4.5005
R18478 DVSS.n14177 DVSS.n14131 4.5005
R18479 DVSS.n14185 DVSS.n14131 4.5005
R18480 DVSS.n14176 DVSS.n14131 4.5005
R18481 DVSS.n14187 DVSS.n14131 4.5005
R18482 DVSS.n14175 DVSS.n14131 4.5005
R18483 DVSS.n14188 DVSS.n14131 4.5005
R18484 DVSS.n14189 DVSS.n14131 4.5005
R18485 DVSS.n21065 DVSS.n14131 4.5005
R18486 DVSS.n21067 DVSS.n14145 4.5005
R18487 DVSS.n14182 DVSS.n14145 4.5005
R18488 DVSS.n14179 DVSS.n14145 4.5005
R18489 DVSS.n14183 DVSS.n14145 4.5005
R18490 DVSS.n14178 DVSS.n14145 4.5005
R18491 DVSS.n14184 DVSS.n14145 4.5005
R18492 DVSS.n14177 DVSS.n14145 4.5005
R18493 DVSS.n14185 DVSS.n14145 4.5005
R18494 DVSS.n14176 DVSS.n14145 4.5005
R18495 DVSS.n14187 DVSS.n14145 4.5005
R18496 DVSS.n14175 DVSS.n14145 4.5005
R18497 DVSS.n14188 DVSS.n14145 4.5005
R18498 DVSS.n14189 DVSS.n14145 4.5005
R18499 DVSS.n21065 DVSS.n14145 4.5005
R18500 DVSS.n21067 DVSS.n14130 4.5005
R18501 DVSS.n14182 DVSS.n14130 4.5005
R18502 DVSS.n14179 DVSS.n14130 4.5005
R18503 DVSS.n14183 DVSS.n14130 4.5005
R18504 DVSS.n14178 DVSS.n14130 4.5005
R18505 DVSS.n14184 DVSS.n14130 4.5005
R18506 DVSS.n14177 DVSS.n14130 4.5005
R18507 DVSS.n14185 DVSS.n14130 4.5005
R18508 DVSS.n14176 DVSS.n14130 4.5005
R18509 DVSS.n14187 DVSS.n14130 4.5005
R18510 DVSS.n14175 DVSS.n14130 4.5005
R18511 DVSS.n14188 DVSS.n14130 4.5005
R18512 DVSS.n14189 DVSS.n14130 4.5005
R18513 DVSS.n21065 DVSS.n14130 4.5005
R18514 DVSS.n21067 DVSS.n14146 4.5005
R18515 DVSS.n14182 DVSS.n14146 4.5005
R18516 DVSS.n14179 DVSS.n14146 4.5005
R18517 DVSS.n14183 DVSS.n14146 4.5005
R18518 DVSS.n14178 DVSS.n14146 4.5005
R18519 DVSS.n14184 DVSS.n14146 4.5005
R18520 DVSS.n14177 DVSS.n14146 4.5005
R18521 DVSS.n14185 DVSS.n14146 4.5005
R18522 DVSS.n14176 DVSS.n14146 4.5005
R18523 DVSS.n14187 DVSS.n14146 4.5005
R18524 DVSS.n14175 DVSS.n14146 4.5005
R18525 DVSS.n14188 DVSS.n14146 4.5005
R18526 DVSS.n14189 DVSS.n14146 4.5005
R18527 DVSS.n21065 DVSS.n14146 4.5005
R18528 DVSS.n21067 DVSS.n14129 4.5005
R18529 DVSS.n14182 DVSS.n14129 4.5005
R18530 DVSS.n14179 DVSS.n14129 4.5005
R18531 DVSS.n14183 DVSS.n14129 4.5005
R18532 DVSS.n14178 DVSS.n14129 4.5005
R18533 DVSS.n14184 DVSS.n14129 4.5005
R18534 DVSS.n14177 DVSS.n14129 4.5005
R18535 DVSS.n14185 DVSS.n14129 4.5005
R18536 DVSS.n14176 DVSS.n14129 4.5005
R18537 DVSS.n14187 DVSS.n14129 4.5005
R18538 DVSS.n14175 DVSS.n14129 4.5005
R18539 DVSS.n14188 DVSS.n14129 4.5005
R18540 DVSS.n14189 DVSS.n14129 4.5005
R18541 DVSS.n21065 DVSS.n14129 4.5005
R18542 DVSS.n21067 DVSS.n14147 4.5005
R18543 DVSS.n14182 DVSS.n14147 4.5005
R18544 DVSS.n14179 DVSS.n14147 4.5005
R18545 DVSS.n14183 DVSS.n14147 4.5005
R18546 DVSS.n14178 DVSS.n14147 4.5005
R18547 DVSS.n14184 DVSS.n14147 4.5005
R18548 DVSS.n14177 DVSS.n14147 4.5005
R18549 DVSS.n14185 DVSS.n14147 4.5005
R18550 DVSS.n14176 DVSS.n14147 4.5005
R18551 DVSS.n14187 DVSS.n14147 4.5005
R18552 DVSS.n14175 DVSS.n14147 4.5005
R18553 DVSS.n14188 DVSS.n14147 4.5005
R18554 DVSS.n14189 DVSS.n14147 4.5005
R18555 DVSS.n21065 DVSS.n14147 4.5005
R18556 DVSS.n21067 DVSS.n14128 4.5005
R18557 DVSS.n14182 DVSS.n14128 4.5005
R18558 DVSS.n14179 DVSS.n14128 4.5005
R18559 DVSS.n14183 DVSS.n14128 4.5005
R18560 DVSS.n14178 DVSS.n14128 4.5005
R18561 DVSS.n14184 DVSS.n14128 4.5005
R18562 DVSS.n14177 DVSS.n14128 4.5005
R18563 DVSS.n14185 DVSS.n14128 4.5005
R18564 DVSS.n14176 DVSS.n14128 4.5005
R18565 DVSS.n14187 DVSS.n14128 4.5005
R18566 DVSS.n14175 DVSS.n14128 4.5005
R18567 DVSS.n14188 DVSS.n14128 4.5005
R18568 DVSS.n14189 DVSS.n14128 4.5005
R18569 DVSS.n21065 DVSS.n14128 4.5005
R18570 DVSS.n21067 DVSS.n14148 4.5005
R18571 DVSS.n14182 DVSS.n14148 4.5005
R18572 DVSS.n14179 DVSS.n14148 4.5005
R18573 DVSS.n14183 DVSS.n14148 4.5005
R18574 DVSS.n14178 DVSS.n14148 4.5005
R18575 DVSS.n14184 DVSS.n14148 4.5005
R18576 DVSS.n14177 DVSS.n14148 4.5005
R18577 DVSS.n14185 DVSS.n14148 4.5005
R18578 DVSS.n14176 DVSS.n14148 4.5005
R18579 DVSS.n14187 DVSS.n14148 4.5005
R18580 DVSS.n14175 DVSS.n14148 4.5005
R18581 DVSS.n14188 DVSS.n14148 4.5005
R18582 DVSS.n14189 DVSS.n14148 4.5005
R18583 DVSS.n21065 DVSS.n14148 4.5005
R18584 DVSS.n21067 DVSS.n14127 4.5005
R18585 DVSS.n14182 DVSS.n14127 4.5005
R18586 DVSS.n14179 DVSS.n14127 4.5005
R18587 DVSS.n14183 DVSS.n14127 4.5005
R18588 DVSS.n14178 DVSS.n14127 4.5005
R18589 DVSS.n14184 DVSS.n14127 4.5005
R18590 DVSS.n14177 DVSS.n14127 4.5005
R18591 DVSS.n14185 DVSS.n14127 4.5005
R18592 DVSS.n14176 DVSS.n14127 4.5005
R18593 DVSS.n14187 DVSS.n14127 4.5005
R18594 DVSS.n14175 DVSS.n14127 4.5005
R18595 DVSS.n14188 DVSS.n14127 4.5005
R18596 DVSS.n14189 DVSS.n14127 4.5005
R18597 DVSS.n21065 DVSS.n14127 4.5005
R18598 DVSS.n21067 DVSS.n14149 4.5005
R18599 DVSS.n14182 DVSS.n14149 4.5005
R18600 DVSS.n14179 DVSS.n14149 4.5005
R18601 DVSS.n14183 DVSS.n14149 4.5005
R18602 DVSS.n14178 DVSS.n14149 4.5005
R18603 DVSS.n14184 DVSS.n14149 4.5005
R18604 DVSS.n14177 DVSS.n14149 4.5005
R18605 DVSS.n14185 DVSS.n14149 4.5005
R18606 DVSS.n14176 DVSS.n14149 4.5005
R18607 DVSS.n14187 DVSS.n14149 4.5005
R18608 DVSS.n14175 DVSS.n14149 4.5005
R18609 DVSS.n14188 DVSS.n14149 4.5005
R18610 DVSS.n14189 DVSS.n14149 4.5005
R18611 DVSS.n21065 DVSS.n14149 4.5005
R18612 DVSS.n21067 DVSS.n14126 4.5005
R18613 DVSS.n14182 DVSS.n14126 4.5005
R18614 DVSS.n14179 DVSS.n14126 4.5005
R18615 DVSS.n14183 DVSS.n14126 4.5005
R18616 DVSS.n14178 DVSS.n14126 4.5005
R18617 DVSS.n14184 DVSS.n14126 4.5005
R18618 DVSS.n14177 DVSS.n14126 4.5005
R18619 DVSS.n14185 DVSS.n14126 4.5005
R18620 DVSS.n14176 DVSS.n14126 4.5005
R18621 DVSS.n14187 DVSS.n14126 4.5005
R18622 DVSS.n14175 DVSS.n14126 4.5005
R18623 DVSS.n14188 DVSS.n14126 4.5005
R18624 DVSS.n14189 DVSS.n14126 4.5005
R18625 DVSS.n14162 DVSS.n14126 4.5005
R18626 DVSS.n21065 DVSS.n14126 4.5005
R18627 DVSS.n21067 DVSS.n21066 4.5005
R18628 DVSS.n21066 DVSS.n14182 4.5005
R18629 DVSS.n21066 DVSS.n14179 4.5005
R18630 DVSS.n21066 DVSS.n14183 4.5005
R18631 DVSS.n21066 DVSS.n14178 4.5005
R18632 DVSS.n21066 DVSS.n14184 4.5005
R18633 DVSS.n21066 DVSS.n14177 4.5005
R18634 DVSS.n21066 DVSS.n14185 4.5005
R18635 DVSS.n21066 DVSS.n14176 4.5005
R18636 DVSS.n21066 DVSS.n14187 4.5005
R18637 DVSS.n21066 DVSS.n14175 4.5005
R18638 DVSS.n21066 DVSS.n14188 4.5005
R18639 DVSS.n21066 DVSS.n14174 4.5005
R18640 DVSS.n21066 DVSS.n14189 4.5005
R18641 DVSS.n21066 DVSS.n14162 4.5005
R18642 DVSS.n21066 DVSS.n21065 4.5005
R18643 DVSS.n14383 DVSS.n14367 4.5005
R18644 DVSS.n14386 DVSS.n14367 4.5005
R18645 DVSS.n14381 DVSS.n14367 4.5005
R18646 DVSS.n14387 DVSS.n14367 4.5005
R18647 DVSS.n14380 DVSS.n14367 4.5005
R18648 DVSS.n14388 DVSS.n14367 4.5005
R18649 DVSS.n14379 DVSS.n14367 4.5005
R18650 DVSS.n14391 DVSS.n14367 4.5005
R18651 DVSS.n14395 DVSS.n14367 4.5005
R18652 DVSS.n20928 DVSS.n14367 4.5005
R18653 DVSS.n14367 DVSS.n14361 4.5005
R18654 DVSS.n20930 DVSS.n14367 4.5005
R18655 DVSS.n14383 DVSS.n14366 4.5005
R18656 DVSS.n14385 DVSS.n14366 4.5005
R18657 DVSS.n14382 DVSS.n14366 4.5005
R18658 DVSS.n14386 DVSS.n14366 4.5005
R18659 DVSS.n14381 DVSS.n14366 4.5005
R18660 DVSS.n14387 DVSS.n14366 4.5005
R18661 DVSS.n14380 DVSS.n14366 4.5005
R18662 DVSS.n14388 DVSS.n14366 4.5005
R18663 DVSS.n14379 DVSS.n14366 4.5005
R18664 DVSS.n14390 DVSS.n14366 4.5005
R18665 DVSS.n14378 DVSS.n14366 4.5005
R18666 DVSS.n14391 DVSS.n14366 4.5005
R18667 DVSS.n14395 DVSS.n14366 4.5005
R18668 DVSS.n20928 DVSS.n14366 4.5005
R18669 DVSS.n14366 DVSS.n14361 4.5005
R18670 DVSS.n20930 DVSS.n14366 4.5005
R18671 DVSS.n14383 DVSS.n14369 4.5005
R18672 DVSS.n14385 DVSS.n14369 4.5005
R18673 DVSS.n14382 DVSS.n14369 4.5005
R18674 DVSS.n14386 DVSS.n14369 4.5005
R18675 DVSS.n14381 DVSS.n14369 4.5005
R18676 DVSS.n14387 DVSS.n14369 4.5005
R18677 DVSS.n14380 DVSS.n14369 4.5005
R18678 DVSS.n14388 DVSS.n14369 4.5005
R18679 DVSS.n14379 DVSS.n14369 4.5005
R18680 DVSS.n14390 DVSS.n14369 4.5005
R18681 DVSS.n14378 DVSS.n14369 4.5005
R18682 DVSS.n14391 DVSS.n14369 4.5005
R18683 DVSS.n14395 DVSS.n14369 4.5005
R18684 DVSS.n20928 DVSS.n14369 4.5005
R18685 DVSS.n20930 DVSS.n14369 4.5005
R18686 DVSS.n14383 DVSS.n14365 4.5005
R18687 DVSS.n14385 DVSS.n14365 4.5005
R18688 DVSS.n14382 DVSS.n14365 4.5005
R18689 DVSS.n14386 DVSS.n14365 4.5005
R18690 DVSS.n14381 DVSS.n14365 4.5005
R18691 DVSS.n14387 DVSS.n14365 4.5005
R18692 DVSS.n14380 DVSS.n14365 4.5005
R18693 DVSS.n14388 DVSS.n14365 4.5005
R18694 DVSS.n14379 DVSS.n14365 4.5005
R18695 DVSS.n14390 DVSS.n14365 4.5005
R18696 DVSS.n14378 DVSS.n14365 4.5005
R18697 DVSS.n14391 DVSS.n14365 4.5005
R18698 DVSS.n20928 DVSS.n14365 4.5005
R18699 DVSS.n20930 DVSS.n14365 4.5005
R18700 DVSS.n14383 DVSS.n14371 4.5005
R18701 DVSS.n14385 DVSS.n14371 4.5005
R18702 DVSS.n14382 DVSS.n14371 4.5005
R18703 DVSS.n14386 DVSS.n14371 4.5005
R18704 DVSS.n14381 DVSS.n14371 4.5005
R18705 DVSS.n14387 DVSS.n14371 4.5005
R18706 DVSS.n14380 DVSS.n14371 4.5005
R18707 DVSS.n14388 DVSS.n14371 4.5005
R18708 DVSS.n14379 DVSS.n14371 4.5005
R18709 DVSS.n14390 DVSS.n14371 4.5005
R18710 DVSS.n14378 DVSS.n14371 4.5005
R18711 DVSS.n14391 DVSS.n14371 4.5005
R18712 DVSS.n20928 DVSS.n14371 4.5005
R18713 DVSS.n20930 DVSS.n14371 4.5005
R18714 DVSS.n14383 DVSS.n14364 4.5005
R18715 DVSS.n14385 DVSS.n14364 4.5005
R18716 DVSS.n14382 DVSS.n14364 4.5005
R18717 DVSS.n14386 DVSS.n14364 4.5005
R18718 DVSS.n14381 DVSS.n14364 4.5005
R18719 DVSS.n14387 DVSS.n14364 4.5005
R18720 DVSS.n14380 DVSS.n14364 4.5005
R18721 DVSS.n14388 DVSS.n14364 4.5005
R18722 DVSS.n14379 DVSS.n14364 4.5005
R18723 DVSS.n14390 DVSS.n14364 4.5005
R18724 DVSS.n14378 DVSS.n14364 4.5005
R18725 DVSS.n14391 DVSS.n14364 4.5005
R18726 DVSS.n20928 DVSS.n14364 4.5005
R18727 DVSS.n20930 DVSS.n14364 4.5005
R18728 DVSS.n14383 DVSS.n14373 4.5005
R18729 DVSS.n14385 DVSS.n14373 4.5005
R18730 DVSS.n14382 DVSS.n14373 4.5005
R18731 DVSS.n14386 DVSS.n14373 4.5005
R18732 DVSS.n14381 DVSS.n14373 4.5005
R18733 DVSS.n14387 DVSS.n14373 4.5005
R18734 DVSS.n14380 DVSS.n14373 4.5005
R18735 DVSS.n14388 DVSS.n14373 4.5005
R18736 DVSS.n14379 DVSS.n14373 4.5005
R18737 DVSS.n14390 DVSS.n14373 4.5005
R18738 DVSS.n14378 DVSS.n14373 4.5005
R18739 DVSS.n14391 DVSS.n14373 4.5005
R18740 DVSS.n20928 DVSS.n14373 4.5005
R18741 DVSS.n20930 DVSS.n14373 4.5005
R18742 DVSS.n14383 DVSS.n14363 4.5005
R18743 DVSS.n14385 DVSS.n14363 4.5005
R18744 DVSS.n14382 DVSS.n14363 4.5005
R18745 DVSS.n14386 DVSS.n14363 4.5005
R18746 DVSS.n14381 DVSS.n14363 4.5005
R18747 DVSS.n14387 DVSS.n14363 4.5005
R18748 DVSS.n14380 DVSS.n14363 4.5005
R18749 DVSS.n14388 DVSS.n14363 4.5005
R18750 DVSS.n14379 DVSS.n14363 4.5005
R18751 DVSS.n14390 DVSS.n14363 4.5005
R18752 DVSS.n14378 DVSS.n14363 4.5005
R18753 DVSS.n14391 DVSS.n14363 4.5005
R18754 DVSS.n20928 DVSS.n14363 4.5005
R18755 DVSS.n20930 DVSS.n14363 4.5005
R18756 DVSS.n14383 DVSS.n14375 4.5005
R18757 DVSS.n14385 DVSS.n14375 4.5005
R18758 DVSS.n14382 DVSS.n14375 4.5005
R18759 DVSS.n14386 DVSS.n14375 4.5005
R18760 DVSS.n14381 DVSS.n14375 4.5005
R18761 DVSS.n14387 DVSS.n14375 4.5005
R18762 DVSS.n14380 DVSS.n14375 4.5005
R18763 DVSS.n14388 DVSS.n14375 4.5005
R18764 DVSS.n14379 DVSS.n14375 4.5005
R18765 DVSS.n14390 DVSS.n14375 4.5005
R18766 DVSS.n14378 DVSS.n14375 4.5005
R18767 DVSS.n14391 DVSS.n14375 4.5005
R18768 DVSS.n20928 DVSS.n14375 4.5005
R18769 DVSS.n20930 DVSS.n14375 4.5005
R18770 DVSS.n14383 DVSS.n14362 4.5005
R18771 DVSS.n14385 DVSS.n14362 4.5005
R18772 DVSS.n14382 DVSS.n14362 4.5005
R18773 DVSS.n14386 DVSS.n14362 4.5005
R18774 DVSS.n14381 DVSS.n14362 4.5005
R18775 DVSS.n14387 DVSS.n14362 4.5005
R18776 DVSS.n14380 DVSS.n14362 4.5005
R18777 DVSS.n14388 DVSS.n14362 4.5005
R18778 DVSS.n14379 DVSS.n14362 4.5005
R18779 DVSS.n14390 DVSS.n14362 4.5005
R18780 DVSS.n14378 DVSS.n14362 4.5005
R18781 DVSS.n14391 DVSS.n14362 4.5005
R18782 DVSS.n20928 DVSS.n14362 4.5005
R18783 DVSS.n20930 DVSS.n14362 4.5005
R18784 DVSS.n20929 DVSS.n14383 4.5005
R18785 DVSS.n20929 DVSS.n14385 4.5005
R18786 DVSS.n20929 DVSS.n14382 4.5005
R18787 DVSS.n20929 DVSS.n14386 4.5005
R18788 DVSS.n20929 DVSS.n14381 4.5005
R18789 DVSS.n20929 DVSS.n14387 4.5005
R18790 DVSS.n20929 DVSS.n14380 4.5005
R18791 DVSS.n20929 DVSS.n14388 4.5005
R18792 DVSS.n20929 DVSS.n14379 4.5005
R18793 DVSS.n20929 DVSS.n14390 4.5005
R18794 DVSS.n20929 DVSS.n14378 4.5005
R18795 DVSS.n20929 DVSS.n14391 4.5005
R18796 DVSS.n20929 DVSS.n20928 4.5005
R18797 DVSS.n20929 DVSS.n14361 4.5005
R18798 DVSS.n20930 DVSS.n20929 4.5005
R18799 DVSS.n19972 DVSS.n14853 4.5005
R18800 DVSS.n15026 DVSS.n14853 4.5005
R18801 DVSS.n15022 DVSS.n14853 4.5005
R18802 DVSS.n15027 DVSS.n14853 4.5005
R18803 DVSS.n15021 DVSS.n14853 4.5005
R18804 DVSS.n15028 DVSS.n14853 4.5005
R18805 DVSS.n15020 DVSS.n14853 4.5005
R18806 DVSS.n15031 DVSS.n14853 4.5005
R18807 DVSS.n15071 DVSS.n14853 4.5005
R18808 DVSS.n15032 DVSS.n14853 4.5005
R18809 DVSS.n19970 DVSS.n14853 4.5005
R18810 DVSS.n19972 DVSS.n15005 4.5005
R18811 DVSS.n15025 DVSS.n15005 4.5005
R18812 DVSS.n15023 DVSS.n15005 4.5005
R18813 DVSS.n15026 DVSS.n15005 4.5005
R18814 DVSS.n15022 DVSS.n15005 4.5005
R18815 DVSS.n15027 DVSS.n15005 4.5005
R18816 DVSS.n15021 DVSS.n15005 4.5005
R18817 DVSS.n15028 DVSS.n15005 4.5005
R18818 DVSS.n15020 DVSS.n15005 4.5005
R18819 DVSS.n15030 DVSS.n15005 4.5005
R18820 DVSS.n15019 DVSS.n15005 4.5005
R18821 DVSS.n15031 DVSS.n15005 4.5005
R18822 DVSS.n15032 DVSS.n15005 4.5005
R18823 DVSS.n19970 DVSS.n15005 4.5005
R18824 DVSS.n19972 DVSS.n15007 4.5005
R18825 DVSS.n15025 DVSS.n15007 4.5005
R18826 DVSS.n15023 DVSS.n15007 4.5005
R18827 DVSS.n15026 DVSS.n15007 4.5005
R18828 DVSS.n15022 DVSS.n15007 4.5005
R18829 DVSS.n15027 DVSS.n15007 4.5005
R18830 DVSS.n15021 DVSS.n15007 4.5005
R18831 DVSS.n15028 DVSS.n15007 4.5005
R18832 DVSS.n15020 DVSS.n15007 4.5005
R18833 DVSS.n15030 DVSS.n15007 4.5005
R18834 DVSS.n15019 DVSS.n15007 4.5005
R18835 DVSS.n15031 DVSS.n15007 4.5005
R18836 DVSS.n15032 DVSS.n15007 4.5005
R18837 DVSS.n19970 DVSS.n15007 4.5005
R18838 DVSS.n19972 DVSS.n15004 4.5005
R18839 DVSS.n15025 DVSS.n15004 4.5005
R18840 DVSS.n15023 DVSS.n15004 4.5005
R18841 DVSS.n15026 DVSS.n15004 4.5005
R18842 DVSS.n15022 DVSS.n15004 4.5005
R18843 DVSS.n15027 DVSS.n15004 4.5005
R18844 DVSS.n15021 DVSS.n15004 4.5005
R18845 DVSS.n15028 DVSS.n15004 4.5005
R18846 DVSS.n15020 DVSS.n15004 4.5005
R18847 DVSS.n15030 DVSS.n15004 4.5005
R18848 DVSS.n15019 DVSS.n15004 4.5005
R18849 DVSS.n15031 DVSS.n15004 4.5005
R18850 DVSS.n15032 DVSS.n15004 4.5005
R18851 DVSS.n19970 DVSS.n15004 4.5005
R18852 DVSS.n19972 DVSS.n15008 4.5005
R18853 DVSS.n15025 DVSS.n15008 4.5005
R18854 DVSS.n15023 DVSS.n15008 4.5005
R18855 DVSS.n15026 DVSS.n15008 4.5005
R18856 DVSS.n15022 DVSS.n15008 4.5005
R18857 DVSS.n15027 DVSS.n15008 4.5005
R18858 DVSS.n15021 DVSS.n15008 4.5005
R18859 DVSS.n15028 DVSS.n15008 4.5005
R18860 DVSS.n15020 DVSS.n15008 4.5005
R18861 DVSS.n15030 DVSS.n15008 4.5005
R18862 DVSS.n15019 DVSS.n15008 4.5005
R18863 DVSS.n15031 DVSS.n15008 4.5005
R18864 DVSS.n15032 DVSS.n15008 4.5005
R18865 DVSS.n19970 DVSS.n15008 4.5005
R18866 DVSS.n19972 DVSS.n15003 4.5005
R18867 DVSS.n15025 DVSS.n15003 4.5005
R18868 DVSS.n15023 DVSS.n15003 4.5005
R18869 DVSS.n15026 DVSS.n15003 4.5005
R18870 DVSS.n15022 DVSS.n15003 4.5005
R18871 DVSS.n15027 DVSS.n15003 4.5005
R18872 DVSS.n15021 DVSS.n15003 4.5005
R18873 DVSS.n15028 DVSS.n15003 4.5005
R18874 DVSS.n15020 DVSS.n15003 4.5005
R18875 DVSS.n15030 DVSS.n15003 4.5005
R18876 DVSS.n15019 DVSS.n15003 4.5005
R18877 DVSS.n15031 DVSS.n15003 4.5005
R18878 DVSS.n15032 DVSS.n15003 4.5005
R18879 DVSS.n19970 DVSS.n15003 4.5005
R18880 DVSS.n19972 DVSS.n15009 4.5005
R18881 DVSS.n15025 DVSS.n15009 4.5005
R18882 DVSS.n15023 DVSS.n15009 4.5005
R18883 DVSS.n15026 DVSS.n15009 4.5005
R18884 DVSS.n15022 DVSS.n15009 4.5005
R18885 DVSS.n15027 DVSS.n15009 4.5005
R18886 DVSS.n15021 DVSS.n15009 4.5005
R18887 DVSS.n15028 DVSS.n15009 4.5005
R18888 DVSS.n15020 DVSS.n15009 4.5005
R18889 DVSS.n15030 DVSS.n15009 4.5005
R18890 DVSS.n15019 DVSS.n15009 4.5005
R18891 DVSS.n15031 DVSS.n15009 4.5005
R18892 DVSS.n15032 DVSS.n15009 4.5005
R18893 DVSS.n19970 DVSS.n15009 4.5005
R18894 DVSS.n19972 DVSS.n15002 4.5005
R18895 DVSS.n15025 DVSS.n15002 4.5005
R18896 DVSS.n15023 DVSS.n15002 4.5005
R18897 DVSS.n15026 DVSS.n15002 4.5005
R18898 DVSS.n15022 DVSS.n15002 4.5005
R18899 DVSS.n15027 DVSS.n15002 4.5005
R18900 DVSS.n15021 DVSS.n15002 4.5005
R18901 DVSS.n15028 DVSS.n15002 4.5005
R18902 DVSS.n15020 DVSS.n15002 4.5005
R18903 DVSS.n15030 DVSS.n15002 4.5005
R18904 DVSS.n15019 DVSS.n15002 4.5005
R18905 DVSS.n15031 DVSS.n15002 4.5005
R18906 DVSS.n15032 DVSS.n15002 4.5005
R18907 DVSS.n19970 DVSS.n15002 4.5005
R18908 DVSS.n19972 DVSS.n15010 4.5005
R18909 DVSS.n15025 DVSS.n15010 4.5005
R18910 DVSS.n15023 DVSS.n15010 4.5005
R18911 DVSS.n15026 DVSS.n15010 4.5005
R18912 DVSS.n15022 DVSS.n15010 4.5005
R18913 DVSS.n15027 DVSS.n15010 4.5005
R18914 DVSS.n15021 DVSS.n15010 4.5005
R18915 DVSS.n15028 DVSS.n15010 4.5005
R18916 DVSS.n15020 DVSS.n15010 4.5005
R18917 DVSS.n15030 DVSS.n15010 4.5005
R18918 DVSS.n15019 DVSS.n15010 4.5005
R18919 DVSS.n15031 DVSS.n15010 4.5005
R18920 DVSS.n15032 DVSS.n15010 4.5005
R18921 DVSS.n19970 DVSS.n15010 4.5005
R18922 DVSS.n19972 DVSS.n15001 4.5005
R18923 DVSS.n15025 DVSS.n15001 4.5005
R18924 DVSS.n15023 DVSS.n15001 4.5005
R18925 DVSS.n15026 DVSS.n15001 4.5005
R18926 DVSS.n15022 DVSS.n15001 4.5005
R18927 DVSS.n15027 DVSS.n15001 4.5005
R18928 DVSS.n15021 DVSS.n15001 4.5005
R18929 DVSS.n15028 DVSS.n15001 4.5005
R18930 DVSS.n15020 DVSS.n15001 4.5005
R18931 DVSS.n15030 DVSS.n15001 4.5005
R18932 DVSS.n15019 DVSS.n15001 4.5005
R18933 DVSS.n15031 DVSS.n15001 4.5005
R18934 DVSS.n15032 DVSS.n15001 4.5005
R18935 DVSS.n19970 DVSS.n15001 4.5005
R18936 DVSS.n19972 DVSS.n19971 4.5005
R18937 DVSS.n19971 DVSS.n15025 4.5005
R18938 DVSS.n19971 DVSS.n15023 4.5005
R18939 DVSS.n19971 DVSS.n15026 4.5005
R18940 DVSS.n19971 DVSS.n15022 4.5005
R18941 DVSS.n19971 DVSS.n15027 4.5005
R18942 DVSS.n19971 DVSS.n15021 4.5005
R18943 DVSS.n19971 DVSS.n15028 4.5005
R18944 DVSS.n19971 DVSS.n15020 4.5005
R18945 DVSS.n19971 DVSS.n15030 4.5005
R18946 DVSS.n19971 DVSS.n15019 4.5005
R18947 DVSS.n19971 DVSS.n15031 4.5005
R18948 DVSS.n19971 DVSS.n15032 4.5005
R18949 DVSS.n19971 DVSS.n15017 4.5005
R18950 DVSS.n19971 DVSS.n19970 4.5005
R18951 DVSS.n18316 DVSS.n15011 4.5005
R18952 DVSS.n15445 DVSS.n15011 4.5005
R18953 DVSS.n15465 DVSS.n15011 4.5005
R18954 DVSS.n15446 DVSS.n15011 4.5005
R18955 DVSS.n15464 DVSS.n15011 4.5005
R18956 DVSS.n15447 DVSS.n15011 4.5005
R18957 DVSS.n15463 DVSS.n15011 4.5005
R18958 DVSS.n15449 DVSS.n15011 4.5005
R18959 DVSS.n15460 DVSS.n15011 4.5005
R18960 DVSS.n15451 DVSS.n15011 4.5005
R18961 DVSS.n15450 DVSS.n15011 4.5005
R18962 DVSS.n18316 DVSS.n15437 4.5005
R18963 DVSS.n15444 DVSS.n15437 4.5005
R18964 DVSS.n18314 DVSS.n15437 4.5005
R18965 DVSS.n15445 DVSS.n15437 4.5005
R18966 DVSS.n15465 DVSS.n15437 4.5005
R18967 DVSS.n15446 DVSS.n15437 4.5005
R18968 DVSS.n15464 DVSS.n15437 4.5005
R18969 DVSS.n15447 DVSS.n15437 4.5005
R18970 DVSS.n15463 DVSS.n15437 4.5005
R18971 DVSS.n15448 DVSS.n15437 4.5005
R18972 DVSS.n15462 DVSS.n15437 4.5005
R18973 DVSS.n15449 DVSS.n15437 4.5005
R18974 DVSS.n15460 DVSS.n15437 4.5005
R18975 DVSS.n15451 DVSS.n15437 4.5005
R18976 DVSS.n15450 DVSS.n15437 4.5005
R18977 DVSS.n18315 DVSS.n15451 4.5005
R18978 DVSS.n18315 DVSS.n15456 4.5005
R18979 DVSS.n18315 DVSS.n15450 4.5005
R18980 DVSS.n15451 DVSS.n15433 4.5005
R18981 DVSS.n15456 DVSS.n15433 4.5005
R18982 DVSS.n15450 DVSS.n15433 4.5005
R18983 DVSS.n18316 DVSS.n15439 4.5005
R18984 DVSS.n15444 DVSS.n15439 4.5005
R18985 DVSS.n18314 DVSS.n15439 4.5005
R18986 DVSS.n15445 DVSS.n15439 4.5005
R18987 DVSS.n15465 DVSS.n15439 4.5005
R18988 DVSS.n15446 DVSS.n15439 4.5005
R18989 DVSS.n15464 DVSS.n15439 4.5005
R18990 DVSS.n15447 DVSS.n15439 4.5005
R18991 DVSS.n15463 DVSS.n15439 4.5005
R18992 DVSS.n15448 DVSS.n15439 4.5005
R18993 DVSS.n15462 DVSS.n15439 4.5005
R18994 DVSS.n15449 DVSS.n15439 4.5005
R18995 DVSS.n15451 DVSS.n15439 4.5005
R18996 DVSS.n15450 DVSS.n15439 4.5005
R18997 DVSS.n18316 DVSS.n15436 4.5005
R18998 DVSS.n15444 DVSS.n15436 4.5005
R18999 DVSS.n18314 DVSS.n15436 4.5005
R19000 DVSS.n15445 DVSS.n15436 4.5005
R19001 DVSS.n15465 DVSS.n15436 4.5005
R19002 DVSS.n15446 DVSS.n15436 4.5005
R19003 DVSS.n15464 DVSS.n15436 4.5005
R19004 DVSS.n15447 DVSS.n15436 4.5005
R19005 DVSS.n15463 DVSS.n15436 4.5005
R19006 DVSS.n15448 DVSS.n15436 4.5005
R19007 DVSS.n15462 DVSS.n15436 4.5005
R19008 DVSS.n15449 DVSS.n15436 4.5005
R19009 DVSS.n15451 DVSS.n15436 4.5005
R19010 DVSS.n15450 DVSS.n15436 4.5005
R19011 DVSS.n18316 DVSS.n15440 4.5005
R19012 DVSS.n15444 DVSS.n15440 4.5005
R19013 DVSS.n18314 DVSS.n15440 4.5005
R19014 DVSS.n15445 DVSS.n15440 4.5005
R19015 DVSS.n15465 DVSS.n15440 4.5005
R19016 DVSS.n15446 DVSS.n15440 4.5005
R19017 DVSS.n15464 DVSS.n15440 4.5005
R19018 DVSS.n15447 DVSS.n15440 4.5005
R19019 DVSS.n15463 DVSS.n15440 4.5005
R19020 DVSS.n15448 DVSS.n15440 4.5005
R19021 DVSS.n15462 DVSS.n15440 4.5005
R19022 DVSS.n15449 DVSS.n15440 4.5005
R19023 DVSS.n15451 DVSS.n15440 4.5005
R19024 DVSS.n15450 DVSS.n15440 4.5005
R19025 DVSS.n18316 DVSS.n15435 4.5005
R19026 DVSS.n15444 DVSS.n15435 4.5005
R19027 DVSS.n18314 DVSS.n15435 4.5005
R19028 DVSS.n15445 DVSS.n15435 4.5005
R19029 DVSS.n15465 DVSS.n15435 4.5005
R19030 DVSS.n15446 DVSS.n15435 4.5005
R19031 DVSS.n15464 DVSS.n15435 4.5005
R19032 DVSS.n15447 DVSS.n15435 4.5005
R19033 DVSS.n15463 DVSS.n15435 4.5005
R19034 DVSS.n15448 DVSS.n15435 4.5005
R19035 DVSS.n15462 DVSS.n15435 4.5005
R19036 DVSS.n15449 DVSS.n15435 4.5005
R19037 DVSS.n15451 DVSS.n15435 4.5005
R19038 DVSS.n15450 DVSS.n15435 4.5005
R19039 DVSS.n18316 DVSS.n15441 4.5005
R19040 DVSS.n15444 DVSS.n15441 4.5005
R19041 DVSS.n18314 DVSS.n15441 4.5005
R19042 DVSS.n15445 DVSS.n15441 4.5005
R19043 DVSS.n15465 DVSS.n15441 4.5005
R19044 DVSS.n15446 DVSS.n15441 4.5005
R19045 DVSS.n15464 DVSS.n15441 4.5005
R19046 DVSS.n15447 DVSS.n15441 4.5005
R19047 DVSS.n15463 DVSS.n15441 4.5005
R19048 DVSS.n15448 DVSS.n15441 4.5005
R19049 DVSS.n15462 DVSS.n15441 4.5005
R19050 DVSS.n15449 DVSS.n15441 4.5005
R19051 DVSS.n15451 DVSS.n15441 4.5005
R19052 DVSS.n15456 DVSS.n15441 4.5005
R19053 DVSS.n15450 DVSS.n15441 4.5005
R19054 DVSS.n18316 DVSS.n15434 4.5005
R19055 DVSS.n15444 DVSS.n15434 4.5005
R19056 DVSS.n18314 DVSS.n15434 4.5005
R19057 DVSS.n15445 DVSS.n15434 4.5005
R19058 DVSS.n15465 DVSS.n15434 4.5005
R19059 DVSS.n15446 DVSS.n15434 4.5005
R19060 DVSS.n15464 DVSS.n15434 4.5005
R19061 DVSS.n15447 DVSS.n15434 4.5005
R19062 DVSS.n15463 DVSS.n15434 4.5005
R19063 DVSS.n15448 DVSS.n15434 4.5005
R19064 DVSS.n15462 DVSS.n15434 4.5005
R19065 DVSS.n15449 DVSS.n15434 4.5005
R19066 DVSS.n15460 DVSS.n15434 4.5005
R19067 DVSS.n15451 DVSS.n15434 4.5005
R19068 DVSS.n15456 DVSS.n15434 4.5005
R19069 DVSS.n15450 DVSS.n15434 4.5005
R19070 DVSS.n15451 DVSS.n15442 4.5005
R19071 DVSS.n15456 DVSS.n15442 4.5005
R19072 DVSS.n15450 DVSS.n15442 4.5005
R19073 DVSS.n17606 DVSS.n16895 4.5005
R19074 DVSS.n16902 DVSS.n16895 4.5005
R19075 DVSS.n17545 DVSS.n16895 4.5005
R19076 DVSS.n16903 DVSS.n16895 4.5005
R19077 DVSS.n17544 DVSS.n16895 4.5005
R19078 DVSS.n16904 DVSS.n16895 4.5005
R19079 DVSS.n17543 DVSS.n16895 4.5005
R19080 DVSS.n16906 DVSS.n16895 4.5005
R19081 DVSS.n17540 DVSS.n16895 4.5005
R19082 DVSS.n16908 DVSS.n16895 4.5005
R19083 DVSS.n16907 DVSS.n16895 4.5005
R19084 DVSS.n17606 DVSS.n16893 4.5005
R19085 DVSS.n16901 DVSS.n16893 4.5005
R19086 DVSS.n17604 DVSS.n16893 4.5005
R19087 DVSS.n16902 DVSS.n16893 4.5005
R19088 DVSS.n17545 DVSS.n16893 4.5005
R19089 DVSS.n16903 DVSS.n16893 4.5005
R19090 DVSS.n17544 DVSS.n16893 4.5005
R19091 DVSS.n16904 DVSS.n16893 4.5005
R19092 DVSS.n17543 DVSS.n16893 4.5005
R19093 DVSS.n16905 DVSS.n16893 4.5005
R19094 DVSS.n17542 DVSS.n16893 4.5005
R19095 DVSS.n16906 DVSS.n16893 4.5005
R19096 DVSS.n16908 DVSS.n16893 4.5005
R19097 DVSS.n16907 DVSS.n16893 4.5005
R19098 DVSS.n17606 DVSS.n16896 4.5005
R19099 DVSS.n16901 DVSS.n16896 4.5005
R19100 DVSS.n17604 DVSS.n16896 4.5005
R19101 DVSS.n16902 DVSS.n16896 4.5005
R19102 DVSS.n17545 DVSS.n16896 4.5005
R19103 DVSS.n16903 DVSS.n16896 4.5005
R19104 DVSS.n17544 DVSS.n16896 4.5005
R19105 DVSS.n16904 DVSS.n16896 4.5005
R19106 DVSS.n17543 DVSS.n16896 4.5005
R19107 DVSS.n16905 DVSS.n16896 4.5005
R19108 DVSS.n17542 DVSS.n16896 4.5005
R19109 DVSS.n16906 DVSS.n16896 4.5005
R19110 DVSS.n16908 DVSS.n16896 4.5005
R19111 DVSS.n16907 DVSS.n16896 4.5005
R19112 DVSS.n17606 DVSS.n16892 4.5005
R19113 DVSS.n16901 DVSS.n16892 4.5005
R19114 DVSS.n17604 DVSS.n16892 4.5005
R19115 DVSS.n16902 DVSS.n16892 4.5005
R19116 DVSS.n17545 DVSS.n16892 4.5005
R19117 DVSS.n16903 DVSS.n16892 4.5005
R19118 DVSS.n17544 DVSS.n16892 4.5005
R19119 DVSS.n16904 DVSS.n16892 4.5005
R19120 DVSS.n17543 DVSS.n16892 4.5005
R19121 DVSS.n16905 DVSS.n16892 4.5005
R19122 DVSS.n17542 DVSS.n16892 4.5005
R19123 DVSS.n16906 DVSS.n16892 4.5005
R19124 DVSS.n16908 DVSS.n16892 4.5005
R19125 DVSS.n16907 DVSS.n16892 4.5005
R19126 DVSS.n17606 DVSS.n16897 4.5005
R19127 DVSS.n16901 DVSS.n16897 4.5005
R19128 DVSS.n17604 DVSS.n16897 4.5005
R19129 DVSS.n16902 DVSS.n16897 4.5005
R19130 DVSS.n17545 DVSS.n16897 4.5005
R19131 DVSS.n16903 DVSS.n16897 4.5005
R19132 DVSS.n17544 DVSS.n16897 4.5005
R19133 DVSS.n16904 DVSS.n16897 4.5005
R19134 DVSS.n17543 DVSS.n16897 4.5005
R19135 DVSS.n16905 DVSS.n16897 4.5005
R19136 DVSS.n17542 DVSS.n16897 4.5005
R19137 DVSS.n16906 DVSS.n16897 4.5005
R19138 DVSS.n16908 DVSS.n16897 4.5005
R19139 DVSS.n17535 DVSS.n16897 4.5005
R19140 DVSS.n16907 DVSS.n16897 4.5005
R19141 DVSS.n17605 DVSS.n16908 4.5005
R19142 DVSS.n17605 DVSS.n17535 4.5005
R19143 DVSS.n17605 DVSS.n16907 4.5005
R19144 DVSS.n16908 DVSS.n16889 4.5005
R19145 DVSS.n17535 DVSS.n16889 4.5005
R19146 DVSS.n16907 DVSS.n16889 4.5005
R19147 DVSS.n17606 DVSS.n16891 4.5005
R19148 DVSS.n16901 DVSS.n16891 4.5005
R19149 DVSS.n17604 DVSS.n16891 4.5005
R19150 DVSS.n16902 DVSS.n16891 4.5005
R19151 DVSS.n17545 DVSS.n16891 4.5005
R19152 DVSS.n16903 DVSS.n16891 4.5005
R19153 DVSS.n17544 DVSS.n16891 4.5005
R19154 DVSS.n16904 DVSS.n16891 4.5005
R19155 DVSS.n17543 DVSS.n16891 4.5005
R19156 DVSS.n16905 DVSS.n16891 4.5005
R19157 DVSS.n17542 DVSS.n16891 4.5005
R19158 DVSS.n16906 DVSS.n16891 4.5005
R19159 DVSS.n16908 DVSS.n16891 4.5005
R19160 DVSS.n16907 DVSS.n16891 4.5005
R19161 DVSS.n17606 DVSS.n16898 4.5005
R19162 DVSS.n16901 DVSS.n16898 4.5005
R19163 DVSS.n17604 DVSS.n16898 4.5005
R19164 DVSS.n16902 DVSS.n16898 4.5005
R19165 DVSS.n17545 DVSS.n16898 4.5005
R19166 DVSS.n16903 DVSS.n16898 4.5005
R19167 DVSS.n17544 DVSS.n16898 4.5005
R19168 DVSS.n16904 DVSS.n16898 4.5005
R19169 DVSS.n17543 DVSS.n16898 4.5005
R19170 DVSS.n16905 DVSS.n16898 4.5005
R19171 DVSS.n17542 DVSS.n16898 4.5005
R19172 DVSS.n16906 DVSS.n16898 4.5005
R19173 DVSS.n16908 DVSS.n16898 4.5005
R19174 DVSS.n16907 DVSS.n16898 4.5005
R19175 DVSS.n17606 DVSS.n16890 4.5005
R19176 DVSS.n16901 DVSS.n16890 4.5005
R19177 DVSS.n17604 DVSS.n16890 4.5005
R19178 DVSS.n16902 DVSS.n16890 4.5005
R19179 DVSS.n17545 DVSS.n16890 4.5005
R19180 DVSS.n16903 DVSS.n16890 4.5005
R19181 DVSS.n17544 DVSS.n16890 4.5005
R19182 DVSS.n16904 DVSS.n16890 4.5005
R19183 DVSS.n17543 DVSS.n16890 4.5005
R19184 DVSS.n16905 DVSS.n16890 4.5005
R19185 DVSS.n17542 DVSS.n16890 4.5005
R19186 DVSS.n16906 DVSS.n16890 4.5005
R19187 DVSS.n16908 DVSS.n16890 4.5005
R19188 DVSS.n16907 DVSS.n16890 4.5005
R19189 DVSS.n17606 DVSS.n16899 4.5005
R19190 DVSS.n16901 DVSS.n16899 4.5005
R19191 DVSS.n17604 DVSS.n16899 4.5005
R19192 DVSS.n16902 DVSS.n16899 4.5005
R19193 DVSS.n17545 DVSS.n16899 4.5005
R19194 DVSS.n16903 DVSS.n16899 4.5005
R19195 DVSS.n17544 DVSS.n16899 4.5005
R19196 DVSS.n16904 DVSS.n16899 4.5005
R19197 DVSS.n17543 DVSS.n16899 4.5005
R19198 DVSS.n16905 DVSS.n16899 4.5005
R19199 DVSS.n17542 DVSS.n16899 4.5005
R19200 DVSS.n16906 DVSS.n16899 4.5005
R19201 DVSS.n17540 DVSS.n16899 4.5005
R19202 DVSS.n16908 DVSS.n16899 4.5005
R19203 DVSS.n16907 DVSS.n16899 4.5005
R19204 DVSS.n15677 DVSS.n15660 4.5005
R19205 DVSS.n15677 DVSS.n15662 4.5005
R19206 DVSS.n15677 DVSS.n15658 4.5005
R19207 DVSS.n15677 DVSS.n15663 4.5005
R19208 DVSS.n15677 DVSS.n15657 4.5005
R19209 DVSS.n15677 DVSS.n15664 4.5005
R19210 DVSS.n15677 DVSS.n15656 4.5005
R19211 DVSS.n15677 DVSS.n15666 4.5005
R19212 DVSS.n15677 DVSS.n15654 4.5005
R19213 DVSS.n15677 DVSS.n15667 4.5005
R19214 DVSS.n18079 DVSS.n15677 4.5005
R19215 DVSS.n15672 DVSS.n15660 4.5005
R19216 DVSS.n15672 DVSS.n15661 4.5005
R19217 DVSS.n15672 DVSS.n15659 4.5005
R19218 DVSS.n15672 DVSS.n15662 4.5005
R19219 DVSS.n15672 DVSS.n15658 4.5005
R19220 DVSS.n15672 DVSS.n15663 4.5005
R19221 DVSS.n15672 DVSS.n15657 4.5005
R19222 DVSS.n15672 DVSS.n15664 4.5005
R19223 DVSS.n15672 DVSS.n15656 4.5005
R19224 DVSS.n15672 DVSS.n15665 4.5005
R19225 DVSS.n15672 DVSS.n15655 4.5005
R19226 DVSS.n15672 DVSS.n15666 4.5005
R19227 DVSS.n15672 DVSS.n15667 4.5005
R19228 DVSS.n18079 DVSS.n15672 4.5005
R19229 DVSS.n15660 DVSS.n15635 4.5005
R19230 DVSS.n15661 DVSS.n15635 4.5005
R19231 DVSS.n15659 DVSS.n15635 4.5005
R19232 DVSS.n15662 DVSS.n15635 4.5005
R19233 DVSS.n15658 DVSS.n15635 4.5005
R19234 DVSS.n15663 DVSS.n15635 4.5005
R19235 DVSS.n15657 DVSS.n15635 4.5005
R19236 DVSS.n15664 DVSS.n15635 4.5005
R19237 DVSS.n15656 DVSS.n15635 4.5005
R19238 DVSS.n15665 DVSS.n15635 4.5005
R19239 DVSS.n15655 DVSS.n15635 4.5005
R19240 DVSS.n15666 DVSS.n15635 4.5005
R19241 DVSS.n15667 DVSS.n15635 4.5005
R19242 DVSS.n15653 DVSS.n15635 4.5005
R19243 DVSS.n18079 DVSS.n15635 4.5005
R19244 DVSS.n18080 DVSS.n15660 4.5005
R19245 DVSS.n18080 DVSS.n15661 4.5005
R19246 DVSS.n18080 DVSS.n15659 4.5005
R19247 DVSS.n18080 DVSS.n15662 4.5005
R19248 DVSS.n18080 DVSS.n15658 4.5005
R19249 DVSS.n18080 DVSS.n15663 4.5005
R19250 DVSS.n18080 DVSS.n15657 4.5005
R19251 DVSS.n18080 DVSS.n15664 4.5005
R19252 DVSS.n18080 DVSS.n15656 4.5005
R19253 DVSS.n18080 DVSS.n15665 4.5005
R19254 DVSS.n18080 DVSS.n15655 4.5005
R19255 DVSS.n18080 DVSS.n15666 4.5005
R19256 DVSS.n18080 DVSS.n15654 4.5005
R19257 DVSS.n18080 DVSS.n15667 4.5005
R19258 DVSS.n18080 DVSS.n15653 4.5005
R19259 DVSS.n18080 DVSS.n18079 4.5005
R19260 DVSS.n15678 DVSS.n15660 4.5005
R19261 DVSS.n15678 DVSS.n15661 4.5005
R19262 DVSS.n15678 DVSS.n15659 4.5005
R19263 DVSS.n15678 DVSS.n15662 4.5005
R19264 DVSS.n15678 DVSS.n15658 4.5005
R19265 DVSS.n15678 DVSS.n15663 4.5005
R19266 DVSS.n15678 DVSS.n15657 4.5005
R19267 DVSS.n15678 DVSS.n15664 4.5005
R19268 DVSS.n15678 DVSS.n15656 4.5005
R19269 DVSS.n15678 DVSS.n15665 4.5005
R19270 DVSS.n15678 DVSS.n15655 4.5005
R19271 DVSS.n15678 DVSS.n15666 4.5005
R19272 DVSS.n15678 DVSS.n15654 4.5005
R19273 DVSS.n15678 DVSS.n15667 4.5005
R19274 DVSS.n15678 DVSS.n15653 4.5005
R19275 DVSS.n18079 DVSS.n15678 4.5005
R19276 DVSS.n15670 DVSS.n15660 4.5005
R19277 DVSS.n15670 DVSS.n15661 4.5005
R19278 DVSS.n15670 DVSS.n15659 4.5005
R19279 DVSS.n15670 DVSS.n15662 4.5005
R19280 DVSS.n15670 DVSS.n15658 4.5005
R19281 DVSS.n15670 DVSS.n15663 4.5005
R19282 DVSS.n15670 DVSS.n15657 4.5005
R19283 DVSS.n15670 DVSS.n15664 4.5005
R19284 DVSS.n15670 DVSS.n15656 4.5005
R19285 DVSS.n15670 DVSS.n15665 4.5005
R19286 DVSS.n15670 DVSS.n15655 4.5005
R19287 DVSS.n15670 DVSS.n15666 4.5005
R19288 DVSS.n15670 DVSS.n15654 4.5005
R19289 DVSS.n15670 DVSS.n15667 4.5005
R19290 DVSS.n15670 DVSS.n15653 4.5005
R19291 DVSS.n18079 DVSS.n15670 4.5005
R19292 DVSS.n18078 DVSS.n15660 4.5005
R19293 DVSS.n18078 DVSS.n15661 4.5005
R19294 DVSS.n18078 DVSS.n15659 4.5005
R19295 DVSS.n18078 DVSS.n15662 4.5005
R19296 DVSS.n18078 DVSS.n15658 4.5005
R19297 DVSS.n18078 DVSS.n15663 4.5005
R19298 DVSS.n18078 DVSS.n15657 4.5005
R19299 DVSS.n18078 DVSS.n15664 4.5005
R19300 DVSS.n18078 DVSS.n15656 4.5005
R19301 DVSS.n18078 DVSS.n15665 4.5005
R19302 DVSS.n18078 DVSS.n15655 4.5005
R19303 DVSS.n18078 DVSS.n15666 4.5005
R19304 DVSS.n18078 DVSS.n15654 4.5005
R19305 DVSS.n18078 DVSS.n15667 4.5005
R19306 DVSS.n18078 DVSS.n15653 4.5005
R19307 DVSS.n18079 DVSS.n18078 4.5005
R19308 DVSS.n15669 DVSS.n15660 4.5005
R19309 DVSS.n15669 DVSS.n15661 4.5005
R19310 DVSS.n15669 DVSS.n15659 4.5005
R19311 DVSS.n15669 DVSS.n15662 4.5005
R19312 DVSS.n15669 DVSS.n15658 4.5005
R19313 DVSS.n15669 DVSS.n15663 4.5005
R19314 DVSS.n15669 DVSS.n15657 4.5005
R19315 DVSS.n15669 DVSS.n15664 4.5005
R19316 DVSS.n15669 DVSS.n15656 4.5005
R19317 DVSS.n15669 DVSS.n15665 4.5005
R19318 DVSS.n15669 DVSS.n15655 4.5005
R19319 DVSS.n15669 DVSS.n15666 4.5005
R19320 DVSS.n15669 DVSS.n15654 4.5005
R19321 DVSS.n15669 DVSS.n15667 4.5005
R19322 DVSS.n15669 DVSS.n15653 4.5005
R19323 DVSS.n18079 DVSS.n15669 4.5005
R19324 DVSS.n18047 DVSS.n15697 4.5005
R19325 DVSS.n18047 DVSS.n15698 4.5005
R19326 DVSS.n18047 DVSS.n15695 4.5005
R19327 DVSS.n18047 DVSS.n15699 4.5005
R19328 DVSS.n18047 DVSS.n15694 4.5005
R19329 DVSS.n18047 DVSS.n15700 4.5005
R19330 DVSS.n18047 DVSS.n15693 4.5005
R19331 DVSS.n18047 DVSS.n15701 4.5005
R19332 DVSS.n18047 DVSS.n15691 4.5005
R19333 DVSS.n18047 DVSS.n15702 4.5005
R19334 DVSS.n18047 DVSS.n15690 4.5005
R19335 DVSS.n18047 DVSS.n18046 4.5005
R19336 DVSS.n15709 DVSS.n15697 4.5005
R19337 DVSS.n15725 DVSS.n15709 4.5005
R19338 DVSS.n15724 DVSS.n15709 4.5005
R19339 DVSS.n15709 DVSS.n15698 4.5005
R19340 DVSS.n15709 DVSS.n15695 4.5005
R19341 DVSS.n15709 DVSS.n15699 4.5005
R19342 DVSS.n15709 DVSS.n15694 4.5005
R19343 DVSS.n15709 DVSS.n15700 4.5005
R19344 DVSS.n15709 DVSS.n15693 4.5005
R19345 DVSS.n18044 DVSS.n15709 4.5005
R19346 DVSS.n15723 DVSS.n15709 4.5005
R19347 DVSS.n15709 DVSS.n15701 4.5005
R19348 DVSS.n15709 DVSS.n15691 4.5005
R19349 DVSS.n15709 DVSS.n15702 4.5005
R19350 DVSS.n15709 DVSS.n15690 4.5005
R19351 DVSS.n18046 DVSS.n15709 4.5005
R19352 DVSS.n15707 DVSS.n15697 4.5005
R19353 DVSS.n15725 DVSS.n15707 4.5005
R19354 DVSS.n15724 DVSS.n15707 4.5005
R19355 DVSS.n15707 DVSS.n15698 4.5005
R19356 DVSS.n15707 DVSS.n15695 4.5005
R19357 DVSS.n15707 DVSS.n15699 4.5005
R19358 DVSS.n15707 DVSS.n15694 4.5005
R19359 DVSS.n15707 DVSS.n15700 4.5005
R19360 DVSS.n15707 DVSS.n15693 4.5005
R19361 DVSS.n18044 DVSS.n15707 4.5005
R19362 DVSS.n15723 DVSS.n15707 4.5005
R19363 DVSS.n15707 DVSS.n15701 4.5005
R19364 DVSS.n15707 DVSS.n15691 4.5005
R19365 DVSS.n15707 DVSS.n15702 4.5005
R19366 DVSS.n15707 DVSS.n15690 4.5005
R19367 DVSS.n18046 DVSS.n15707 4.5005
R19368 DVSS.n15710 DVSS.n15697 4.5005
R19369 DVSS.n15725 DVSS.n15710 4.5005
R19370 DVSS.n15724 DVSS.n15710 4.5005
R19371 DVSS.n15710 DVSS.n15698 4.5005
R19372 DVSS.n15710 DVSS.n15695 4.5005
R19373 DVSS.n15710 DVSS.n15699 4.5005
R19374 DVSS.n15710 DVSS.n15694 4.5005
R19375 DVSS.n15710 DVSS.n15700 4.5005
R19376 DVSS.n15710 DVSS.n15693 4.5005
R19377 DVSS.n18044 DVSS.n15710 4.5005
R19378 DVSS.n15723 DVSS.n15710 4.5005
R19379 DVSS.n15710 DVSS.n15701 4.5005
R19380 DVSS.n15710 DVSS.n15691 4.5005
R19381 DVSS.n15710 DVSS.n15702 4.5005
R19382 DVSS.n15710 DVSS.n15690 4.5005
R19383 DVSS.n18046 DVSS.n15710 4.5005
R19384 DVSS.n15706 DVSS.n15697 4.5005
R19385 DVSS.n15725 DVSS.n15706 4.5005
R19386 DVSS.n15724 DVSS.n15706 4.5005
R19387 DVSS.n15706 DVSS.n15698 4.5005
R19388 DVSS.n15706 DVSS.n15695 4.5005
R19389 DVSS.n15706 DVSS.n15699 4.5005
R19390 DVSS.n15706 DVSS.n15694 4.5005
R19391 DVSS.n15706 DVSS.n15700 4.5005
R19392 DVSS.n15706 DVSS.n15693 4.5005
R19393 DVSS.n18044 DVSS.n15706 4.5005
R19394 DVSS.n15723 DVSS.n15706 4.5005
R19395 DVSS.n15706 DVSS.n15701 4.5005
R19396 DVSS.n15706 DVSS.n15691 4.5005
R19397 DVSS.n15706 DVSS.n15702 4.5005
R19398 DVSS.n15706 DVSS.n15690 4.5005
R19399 DVSS.n18046 DVSS.n15706 4.5005
R19400 DVSS.n15719 DVSS.n15697 4.5005
R19401 DVSS.n15725 DVSS.n15719 4.5005
R19402 DVSS.n15724 DVSS.n15719 4.5005
R19403 DVSS.n15719 DVSS.n15698 4.5005
R19404 DVSS.n15719 DVSS.n15695 4.5005
R19405 DVSS.n15719 DVSS.n15699 4.5005
R19406 DVSS.n15719 DVSS.n15694 4.5005
R19407 DVSS.n15719 DVSS.n15700 4.5005
R19408 DVSS.n15719 DVSS.n15693 4.5005
R19409 DVSS.n18044 DVSS.n15719 4.5005
R19410 DVSS.n15723 DVSS.n15719 4.5005
R19411 DVSS.n15719 DVSS.n15701 4.5005
R19412 DVSS.n15719 DVSS.n15691 4.5005
R19413 DVSS.n15719 DVSS.n15702 4.5005
R19414 DVSS.n18046 DVSS.n15719 4.5005
R19415 DVSS.n15705 DVSS.n15697 4.5005
R19416 DVSS.n15725 DVSS.n15705 4.5005
R19417 DVSS.n15724 DVSS.n15705 4.5005
R19418 DVSS.n15705 DVSS.n15698 4.5005
R19419 DVSS.n15705 DVSS.n15695 4.5005
R19420 DVSS.n15705 DVSS.n15699 4.5005
R19421 DVSS.n15705 DVSS.n15694 4.5005
R19422 DVSS.n15705 DVSS.n15700 4.5005
R19423 DVSS.n15705 DVSS.n15693 4.5005
R19424 DVSS.n18044 DVSS.n15705 4.5005
R19425 DVSS.n15723 DVSS.n15705 4.5005
R19426 DVSS.n15705 DVSS.n15701 4.5005
R19427 DVSS.n15705 DVSS.n15702 4.5005
R19428 DVSS.n18046 DVSS.n15705 4.5005
R19429 DVSS.n15722 DVSS.n15697 4.5005
R19430 DVSS.n15725 DVSS.n15722 4.5005
R19431 DVSS.n15724 DVSS.n15722 4.5005
R19432 DVSS.n15722 DVSS.n15698 4.5005
R19433 DVSS.n15722 DVSS.n15695 4.5005
R19434 DVSS.n15722 DVSS.n15699 4.5005
R19435 DVSS.n15722 DVSS.n15694 4.5005
R19436 DVSS.n15722 DVSS.n15700 4.5005
R19437 DVSS.n15722 DVSS.n15693 4.5005
R19438 DVSS.n18044 DVSS.n15722 4.5005
R19439 DVSS.n15723 DVSS.n15722 4.5005
R19440 DVSS.n15722 DVSS.n15701 4.5005
R19441 DVSS.n15722 DVSS.n15702 4.5005
R19442 DVSS.n18046 DVSS.n15722 4.5005
R19443 DVSS.n15704 DVSS.n15697 4.5005
R19444 DVSS.n15725 DVSS.n15704 4.5005
R19445 DVSS.n15724 DVSS.n15704 4.5005
R19446 DVSS.n15704 DVSS.n15698 4.5005
R19447 DVSS.n15704 DVSS.n15695 4.5005
R19448 DVSS.n15704 DVSS.n15699 4.5005
R19449 DVSS.n15704 DVSS.n15694 4.5005
R19450 DVSS.n15704 DVSS.n15700 4.5005
R19451 DVSS.n15704 DVSS.n15693 4.5005
R19452 DVSS.n18044 DVSS.n15704 4.5005
R19453 DVSS.n15723 DVSS.n15704 4.5005
R19454 DVSS.n15704 DVSS.n15701 4.5005
R19455 DVSS.n15704 DVSS.n15691 4.5005
R19456 DVSS.n15704 DVSS.n15702 4.5005
R19457 DVSS.n18046 DVSS.n15704 4.5005
R19458 DVSS.n18045 DVSS.n15697 4.5005
R19459 DVSS.n18045 DVSS.n15725 4.5005
R19460 DVSS.n18045 DVSS.n15724 4.5005
R19461 DVSS.n18045 DVSS.n15698 4.5005
R19462 DVSS.n18045 DVSS.n15695 4.5005
R19463 DVSS.n18045 DVSS.n15699 4.5005
R19464 DVSS.n18045 DVSS.n15694 4.5005
R19465 DVSS.n18045 DVSS.n15700 4.5005
R19466 DVSS.n18045 DVSS.n15693 4.5005
R19467 DVSS.n18045 DVSS.n18044 4.5005
R19468 DVSS.n18045 DVSS.n15723 4.5005
R19469 DVSS.n18045 DVSS.n15701 4.5005
R19470 DVSS.n18045 DVSS.n15691 4.5005
R19471 DVSS.n18045 DVSS.n15702 4.5005
R19472 DVSS.n18045 DVSS.n15690 4.5005
R19473 DVSS.n18046 DVSS.n18045 4.5005
R19474 DVSS.n15660 DVSS.n15646 4.5005
R19475 DVSS.n15661 DVSS.n15646 4.5005
R19476 DVSS.n15659 DVSS.n15646 4.5005
R19477 DVSS.n15662 DVSS.n15646 4.5005
R19478 DVSS.n15658 DVSS.n15646 4.5005
R19479 DVSS.n15663 DVSS.n15646 4.5005
R19480 DVSS.n15657 DVSS.n15646 4.5005
R19481 DVSS.n15664 DVSS.n15646 4.5005
R19482 DVSS.n15656 DVSS.n15646 4.5005
R19483 DVSS.n15665 DVSS.n15646 4.5005
R19484 DVSS.n15655 DVSS.n15646 4.5005
R19485 DVSS.n15666 DVSS.n15646 4.5005
R19486 DVSS.n15654 DVSS.n15646 4.5005
R19487 DVSS.n15667 DVSS.n15646 4.5005
R19488 DVSS.n15653 DVSS.n15646 4.5005
R19489 DVSS.n18079 DVSS.n15646 4.5005
R19490 DVSS.n15660 DVSS.n15650 4.5005
R19491 DVSS.n15661 DVSS.n15650 4.5005
R19492 DVSS.n15659 DVSS.n15650 4.5005
R19493 DVSS.n15662 DVSS.n15650 4.5005
R19494 DVSS.n15658 DVSS.n15650 4.5005
R19495 DVSS.n15663 DVSS.n15650 4.5005
R19496 DVSS.n15657 DVSS.n15650 4.5005
R19497 DVSS.n15664 DVSS.n15650 4.5005
R19498 DVSS.n15656 DVSS.n15650 4.5005
R19499 DVSS.n15665 DVSS.n15650 4.5005
R19500 DVSS.n15655 DVSS.n15650 4.5005
R19501 DVSS.n15666 DVSS.n15650 4.5005
R19502 DVSS.n15654 DVSS.n15650 4.5005
R19503 DVSS.n15667 DVSS.n15650 4.5005
R19504 DVSS.n15653 DVSS.n15650 4.5005
R19505 DVSS.n18079 DVSS.n15650 4.5005
R19506 DVSS.n15660 DVSS.n15630 4.5005
R19507 DVSS.n15661 DVSS.n15630 4.5005
R19508 DVSS.n15659 DVSS.n15630 4.5005
R19509 DVSS.n15662 DVSS.n15630 4.5005
R19510 DVSS.n15658 DVSS.n15630 4.5005
R19511 DVSS.n15663 DVSS.n15630 4.5005
R19512 DVSS.n15657 DVSS.n15630 4.5005
R19513 DVSS.n15664 DVSS.n15630 4.5005
R19514 DVSS.n15656 DVSS.n15630 4.5005
R19515 DVSS.n15665 DVSS.n15630 4.5005
R19516 DVSS.n15655 DVSS.n15630 4.5005
R19517 DVSS.n15666 DVSS.n15630 4.5005
R19518 DVSS.n15654 DVSS.n15630 4.5005
R19519 DVSS.n15667 DVSS.n15630 4.5005
R19520 DVSS.n15653 DVSS.n15630 4.5005
R19521 DVSS.n18079 DVSS.n15630 4.5005
R19522 DVSS.n16906 DVSS.n16889 4.5005
R19523 DVSS.n17542 DVSS.n16889 4.5005
R19524 DVSS.n16905 DVSS.n16889 4.5005
R19525 DVSS.n17543 DVSS.n16889 4.5005
R19526 DVSS.n16904 DVSS.n16889 4.5005
R19527 DVSS.n17544 DVSS.n16889 4.5005
R19528 DVSS.n16903 DVSS.n16889 4.5005
R19529 DVSS.n17545 DVSS.n16889 4.5005
R19530 DVSS.n16902 DVSS.n16889 4.5005
R19531 DVSS.n17604 DVSS.n16889 4.5005
R19532 DVSS.n16901 DVSS.n16889 4.5005
R19533 DVSS.n17606 DVSS.n16889 4.5005
R19534 DVSS.n17605 DVSS.n17540 4.5005
R19535 DVSS.n17605 DVSS.n16906 4.5005
R19536 DVSS.n17605 DVSS.n17542 4.5005
R19537 DVSS.n17605 DVSS.n16905 4.5005
R19538 DVSS.n17605 DVSS.n17543 4.5005
R19539 DVSS.n17605 DVSS.n16904 4.5005
R19540 DVSS.n17605 DVSS.n17544 4.5005
R19541 DVSS.n17605 DVSS.n16903 4.5005
R19542 DVSS.n17605 DVSS.n17545 4.5005
R19543 DVSS.n17605 DVSS.n16902 4.5005
R19544 DVSS.n17605 DVSS.n17604 4.5005
R19545 DVSS.n17605 DVSS.n16901 4.5005
R19546 DVSS.n17606 DVSS.n17605 4.5005
R19547 DVSS.n15460 DVSS.n15442 4.5005
R19548 DVSS.n15449 DVSS.n15442 4.5005
R19549 DVSS.n15462 DVSS.n15442 4.5005
R19550 DVSS.n15448 DVSS.n15442 4.5005
R19551 DVSS.n15463 DVSS.n15442 4.5005
R19552 DVSS.n15447 DVSS.n15442 4.5005
R19553 DVSS.n15464 DVSS.n15442 4.5005
R19554 DVSS.n15446 DVSS.n15442 4.5005
R19555 DVSS.n15465 DVSS.n15442 4.5005
R19556 DVSS.n15445 DVSS.n15442 4.5005
R19557 DVSS.n18314 DVSS.n15442 4.5005
R19558 DVSS.n15444 DVSS.n15442 4.5005
R19559 DVSS.n18316 DVSS.n15442 4.5005
R19560 DVSS.n15449 DVSS.n15433 4.5005
R19561 DVSS.n15462 DVSS.n15433 4.5005
R19562 DVSS.n15448 DVSS.n15433 4.5005
R19563 DVSS.n15463 DVSS.n15433 4.5005
R19564 DVSS.n15447 DVSS.n15433 4.5005
R19565 DVSS.n15464 DVSS.n15433 4.5005
R19566 DVSS.n15446 DVSS.n15433 4.5005
R19567 DVSS.n15465 DVSS.n15433 4.5005
R19568 DVSS.n15445 DVSS.n15433 4.5005
R19569 DVSS.n18314 DVSS.n15433 4.5005
R19570 DVSS.n15444 DVSS.n15433 4.5005
R19571 DVSS.n18316 DVSS.n15433 4.5005
R19572 DVSS.n18315 DVSS.n15460 4.5005
R19573 DVSS.n18315 DVSS.n15449 4.5005
R19574 DVSS.n18315 DVSS.n15462 4.5005
R19575 DVSS.n18315 DVSS.n15448 4.5005
R19576 DVSS.n18315 DVSS.n15463 4.5005
R19577 DVSS.n18315 DVSS.n15447 4.5005
R19578 DVSS.n18315 DVSS.n15464 4.5005
R19579 DVSS.n18315 DVSS.n15446 4.5005
R19580 DVSS.n18315 DVSS.n15465 4.5005
R19581 DVSS.n18315 DVSS.n15445 4.5005
R19582 DVSS.n18315 DVSS.n18314 4.5005
R19583 DVSS.n18315 DVSS.n15444 4.5005
R19584 DVSS.n18316 DVSS.n18315 4.5005
R19585 DVSS.n13450 DVSS.n13429 4.5005
R19586 DVSS.n13437 DVSS.n13429 4.5005
R19587 DVSS.n13449 DVSS.n13429 4.5005
R19588 DVSS.n13438 DVSS.n13429 4.5005
R19589 DVSS.n13447 DVSS.n13429 4.5005
R19590 DVSS.n13439 DVSS.n13429 4.5005
R19591 DVSS.n13446 DVSS.n13429 4.5005
R19592 DVSS.n13440 DVSS.n13429 4.5005
R19593 DVSS.n13445 DVSS.n13429 4.5005
R19594 DVSS.n13441 DVSS.n13429 4.5005
R19595 DVSS.n13444 DVSS.n13429 4.5005
R19596 DVSS.n13442 DVSS.n13429 4.5005
R19597 DVSS.n13450 DVSS.n13421 4.5005
R19598 DVSS.n13437 DVSS.n13421 4.5005
R19599 DVSS.n13449 DVSS.n13421 4.5005
R19600 DVSS.n13438 DVSS.n13421 4.5005
R19601 DVSS.n13447 DVSS.n13421 4.5005
R19602 DVSS.n13439 DVSS.n13421 4.5005
R19603 DVSS.n13446 DVSS.n13421 4.5005
R19604 DVSS.n13440 DVSS.n13421 4.5005
R19605 DVSS.n13445 DVSS.n13421 4.5005
R19606 DVSS.n13441 DVSS.n13421 4.5005
R19607 DVSS.n13444 DVSS.n13421 4.5005
R19608 DVSS.n13442 DVSS.n13421 4.5005
R19609 DVSS.n13450 DVSS.n13428 4.5005
R19610 DVSS.n13437 DVSS.n13428 4.5005
R19611 DVSS.n13449 DVSS.n13428 4.5005
R19612 DVSS.n13438 DVSS.n13428 4.5005
R19613 DVSS.n13447 DVSS.n13428 4.5005
R19614 DVSS.n13439 DVSS.n13428 4.5005
R19615 DVSS.n13446 DVSS.n13428 4.5005
R19616 DVSS.n13440 DVSS.n13428 4.5005
R19617 DVSS.n13445 DVSS.n13428 4.5005
R19618 DVSS.n13441 DVSS.n13428 4.5005
R19619 DVSS.n13444 DVSS.n13428 4.5005
R19620 DVSS.n13442 DVSS.n13428 4.5005
R19621 DVSS.n13450 DVSS.n13422 4.5005
R19622 DVSS.n13437 DVSS.n13422 4.5005
R19623 DVSS.n13449 DVSS.n13422 4.5005
R19624 DVSS.n13438 DVSS.n13422 4.5005
R19625 DVSS.n13447 DVSS.n13422 4.5005
R19626 DVSS.n13439 DVSS.n13422 4.5005
R19627 DVSS.n13446 DVSS.n13422 4.5005
R19628 DVSS.n13440 DVSS.n13422 4.5005
R19629 DVSS.n13445 DVSS.n13422 4.5005
R19630 DVSS.n13441 DVSS.n13422 4.5005
R19631 DVSS.n13444 DVSS.n13422 4.5005
R19632 DVSS.n13442 DVSS.n13422 4.5005
R19633 DVSS.n13450 DVSS.n13427 4.5005
R19634 DVSS.n13437 DVSS.n13427 4.5005
R19635 DVSS.n13449 DVSS.n13427 4.5005
R19636 DVSS.n13438 DVSS.n13427 4.5005
R19637 DVSS.n13447 DVSS.n13427 4.5005
R19638 DVSS.n13439 DVSS.n13427 4.5005
R19639 DVSS.n13446 DVSS.n13427 4.5005
R19640 DVSS.n13440 DVSS.n13427 4.5005
R19641 DVSS.n13445 DVSS.n13427 4.5005
R19642 DVSS.n13441 DVSS.n13427 4.5005
R19643 DVSS.n13444 DVSS.n13427 4.5005
R19644 DVSS.n13442 DVSS.n13427 4.5005
R19645 DVSS.n13450 DVSS.n13423 4.5005
R19646 DVSS.n13437 DVSS.n13423 4.5005
R19647 DVSS.n13449 DVSS.n13423 4.5005
R19648 DVSS.n13438 DVSS.n13423 4.5005
R19649 DVSS.n13447 DVSS.n13423 4.5005
R19650 DVSS.n13439 DVSS.n13423 4.5005
R19651 DVSS.n13446 DVSS.n13423 4.5005
R19652 DVSS.n13440 DVSS.n13423 4.5005
R19653 DVSS.n13445 DVSS.n13423 4.5005
R19654 DVSS.n13441 DVSS.n13423 4.5005
R19655 DVSS.n13444 DVSS.n13423 4.5005
R19656 DVSS.n13442 DVSS.n13423 4.5005
R19657 DVSS.n13450 DVSS.n13426 4.5005
R19658 DVSS.n13437 DVSS.n13426 4.5005
R19659 DVSS.n13449 DVSS.n13426 4.5005
R19660 DVSS.n13438 DVSS.n13426 4.5005
R19661 DVSS.n13447 DVSS.n13426 4.5005
R19662 DVSS.n13439 DVSS.n13426 4.5005
R19663 DVSS.n13446 DVSS.n13426 4.5005
R19664 DVSS.n13440 DVSS.n13426 4.5005
R19665 DVSS.n13445 DVSS.n13426 4.5005
R19666 DVSS.n13441 DVSS.n13426 4.5005
R19667 DVSS.n13444 DVSS.n13426 4.5005
R19668 DVSS.n13442 DVSS.n13426 4.5005
R19669 DVSS.n13450 DVSS.n13424 4.5005
R19670 DVSS.n13437 DVSS.n13424 4.5005
R19671 DVSS.n13449 DVSS.n13424 4.5005
R19672 DVSS.n13438 DVSS.n13424 4.5005
R19673 DVSS.n13447 DVSS.n13424 4.5005
R19674 DVSS.n13439 DVSS.n13424 4.5005
R19675 DVSS.n13446 DVSS.n13424 4.5005
R19676 DVSS.n13440 DVSS.n13424 4.5005
R19677 DVSS.n13445 DVSS.n13424 4.5005
R19678 DVSS.n13441 DVSS.n13424 4.5005
R19679 DVSS.n13444 DVSS.n13424 4.5005
R19680 DVSS.n13442 DVSS.n13424 4.5005
R19681 DVSS.n13450 DVSS.n13425 4.5005
R19682 DVSS.n13437 DVSS.n13425 4.5005
R19683 DVSS.n13449 DVSS.n13425 4.5005
R19684 DVSS.n13438 DVSS.n13425 4.5005
R19685 DVSS.n13447 DVSS.n13425 4.5005
R19686 DVSS.n13439 DVSS.n13425 4.5005
R19687 DVSS.n13446 DVSS.n13425 4.5005
R19688 DVSS.n13440 DVSS.n13425 4.5005
R19689 DVSS.n13445 DVSS.n13425 4.5005
R19690 DVSS.n13441 DVSS.n13425 4.5005
R19691 DVSS.n13444 DVSS.n13425 4.5005
R19692 DVSS.n13442 DVSS.n13425 4.5005
R19693 DVSS.n6655 DVSS.n6654 4.5005
R19694 DVSS.n6655 DVSS.n6652 4.5005
R19695 DVSS.n6655 DVSS.n6602 4.5005
R19696 DVSS.n6655 DVSS.n6259 4.5005
R19697 DVSS.n12745 DVSS.n12359 4.5005
R19698 DVSS.n12745 DVSS.n12506 4.5005
R19699 DVSS.n12745 DVSS.n12360 4.5005
R19700 DVSS.n12745 DVSS.n12553 4.5005
R19701 DVSS.n6654 DVSS.n6309 4.5005
R19702 DVSS.n6602 DVSS.n6309 4.5005
R19703 DVSS.n6656 DVSS.n6309 4.5005
R19704 DVSS.n12743 DVSS.n12359 4.5005
R19705 DVSS.n12743 DVSS.n12506 4.5005
R19706 DVSS.n12743 DVSS.n12360 4.5005
R19707 DVSS.n12411 DVSS.n12359 4.5005
R19708 DVSS.n12411 DVSS.n12360 4.5005
R19709 DVSS.n12768 DVSS.n12411 4.5005
R19710 DVSS.n12409 DVSS.n12359 4.5005
R19711 DVSS.n12409 DVSS.n12360 4.5005
R19712 DVSS.n12768 DVSS.n12409 4.5005
R19713 DVSS.n12412 DVSS.n12359 4.5005
R19714 DVSS.n12412 DVSS.n12360 4.5005
R19715 DVSS.n12768 DVSS.n12412 4.5005
R19716 DVSS.n12408 DVSS.n12359 4.5005
R19717 DVSS.n12408 DVSS.n12360 4.5005
R19718 DVSS.n12768 DVSS.n12408 4.5005
R19719 DVSS.n12413 DVSS.n12359 4.5005
R19720 DVSS.n12413 DVSS.n12360 4.5005
R19721 DVSS.n12768 DVSS.n12413 4.5005
R19722 DVSS.n12407 DVSS.n12359 4.5005
R19723 DVSS.n12407 DVSS.n12360 4.5005
R19724 DVSS.n12768 DVSS.n12407 4.5005
R19725 DVSS.n12414 DVSS.n12359 4.5005
R19726 DVSS.n12414 DVSS.n12360 4.5005
R19727 DVSS.n12768 DVSS.n12414 4.5005
R19728 DVSS.n12406 DVSS.n12359 4.5005
R19729 DVSS.n12406 DVSS.n12360 4.5005
R19730 DVSS.n12768 DVSS.n12406 4.5005
R19731 DVSS.n12415 DVSS.n12359 4.5005
R19732 DVSS.n12415 DVSS.n12360 4.5005
R19733 DVSS.n12768 DVSS.n12415 4.5005
R19734 DVSS.n12405 DVSS.n12359 4.5005
R19735 DVSS.n12405 DVSS.n12360 4.5005
R19736 DVSS.n12768 DVSS.n12405 4.5005
R19737 DVSS.n12416 DVSS.n12359 4.5005
R19738 DVSS.n12416 DVSS.n12360 4.5005
R19739 DVSS.n12768 DVSS.n12416 4.5005
R19740 DVSS.n12404 DVSS.n12359 4.5005
R19741 DVSS.n12404 DVSS.n12360 4.5005
R19742 DVSS.n12768 DVSS.n12404 4.5005
R19743 DVSS.n12417 DVSS.n12359 4.5005
R19744 DVSS.n12417 DVSS.n12360 4.5005
R19745 DVSS.n12768 DVSS.n12417 4.5005
R19746 DVSS.n12403 DVSS.n12359 4.5005
R19747 DVSS.n12403 DVSS.n12360 4.5005
R19748 DVSS.n12768 DVSS.n12403 4.5005
R19749 DVSS.n12418 DVSS.n12359 4.5005
R19750 DVSS.n12418 DVSS.n12360 4.5005
R19751 DVSS.n12768 DVSS.n12418 4.5005
R19752 DVSS.n12402 DVSS.n12359 4.5005
R19753 DVSS.n12402 DVSS.n12360 4.5005
R19754 DVSS.n12768 DVSS.n12402 4.5005
R19755 DVSS.n12419 DVSS.n12359 4.5005
R19756 DVSS.n12419 DVSS.n12360 4.5005
R19757 DVSS.n12768 DVSS.n12419 4.5005
R19758 DVSS.n12401 DVSS.n12359 4.5005
R19759 DVSS.n12401 DVSS.n12360 4.5005
R19760 DVSS.n12768 DVSS.n12401 4.5005
R19761 DVSS.n12420 DVSS.n12359 4.5005
R19762 DVSS.n12420 DVSS.n12360 4.5005
R19763 DVSS.n12768 DVSS.n12420 4.5005
R19764 DVSS.n12400 DVSS.n12359 4.5005
R19765 DVSS.n12400 DVSS.n12360 4.5005
R19766 DVSS.n12768 DVSS.n12400 4.5005
R19767 DVSS.n12421 DVSS.n12359 4.5005
R19768 DVSS.n12421 DVSS.n12360 4.5005
R19769 DVSS.n12768 DVSS.n12421 4.5005
R19770 DVSS.n12399 DVSS.n12359 4.5005
R19771 DVSS.n12399 DVSS.n12360 4.5005
R19772 DVSS.n12768 DVSS.n12399 4.5005
R19773 DVSS.n12422 DVSS.n12359 4.5005
R19774 DVSS.n12422 DVSS.n12360 4.5005
R19775 DVSS.n12768 DVSS.n12422 4.5005
R19776 DVSS.n12398 DVSS.n12359 4.5005
R19777 DVSS.n12398 DVSS.n12360 4.5005
R19778 DVSS.n12768 DVSS.n12398 4.5005
R19779 DVSS.n12423 DVSS.n12359 4.5005
R19780 DVSS.n12423 DVSS.n12360 4.5005
R19781 DVSS.n12768 DVSS.n12423 4.5005
R19782 DVSS.n12397 DVSS.n12359 4.5005
R19783 DVSS.n12397 DVSS.n12360 4.5005
R19784 DVSS.n12768 DVSS.n12397 4.5005
R19785 DVSS.n12424 DVSS.n12359 4.5005
R19786 DVSS.n12424 DVSS.n12360 4.5005
R19787 DVSS.n12768 DVSS.n12424 4.5005
R19788 DVSS.n12396 DVSS.n12359 4.5005
R19789 DVSS.n12396 DVSS.n12360 4.5005
R19790 DVSS.n12768 DVSS.n12396 4.5005
R19791 DVSS.n12425 DVSS.n12359 4.5005
R19792 DVSS.n12425 DVSS.n12360 4.5005
R19793 DVSS.n12768 DVSS.n12425 4.5005
R19794 DVSS.n12395 DVSS.n12359 4.5005
R19795 DVSS.n12395 DVSS.n12360 4.5005
R19796 DVSS.n12768 DVSS.n12395 4.5005
R19797 DVSS.n12426 DVSS.n12359 4.5005
R19798 DVSS.n12426 DVSS.n12360 4.5005
R19799 DVSS.n12768 DVSS.n12426 4.5005
R19800 DVSS.n12394 DVSS.n12359 4.5005
R19801 DVSS.n12394 DVSS.n12360 4.5005
R19802 DVSS.n12768 DVSS.n12394 4.5005
R19803 DVSS.n12427 DVSS.n12359 4.5005
R19804 DVSS.n12427 DVSS.n12360 4.5005
R19805 DVSS.n12768 DVSS.n12427 4.5005
R19806 DVSS.n12393 DVSS.n12359 4.5005
R19807 DVSS.n12393 DVSS.n12360 4.5005
R19808 DVSS.n12768 DVSS.n12393 4.5005
R19809 DVSS.n12428 DVSS.n12359 4.5005
R19810 DVSS.n12428 DVSS.n12360 4.5005
R19811 DVSS.n12768 DVSS.n12428 4.5005
R19812 DVSS.n12392 DVSS.n12359 4.5005
R19813 DVSS.n12392 DVSS.n12360 4.5005
R19814 DVSS.n12768 DVSS.n12392 4.5005
R19815 DVSS.n12429 DVSS.n12359 4.5005
R19816 DVSS.n12429 DVSS.n12360 4.5005
R19817 DVSS.n12768 DVSS.n12429 4.5005
R19818 DVSS.n12391 DVSS.n12359 4.5005
R19819 DVSS.n12391 DVSS.n12360 4.5005
R19820 DVSS.n12768 DVSS.n12391 4.5005
R19821 DVSS.n12430 DVSS.n12359 4.5005
R19822 DVSS.n12430 DVSS.n12360 4.5005
R19823 DVSS.n12768 DVSS.n12430 4.5005
R19824 DVSS.n12390 DVSS.n12359 4.5005
R19825 DVSS.n12390 DVSS.n12360 4.5005
R19826 DVSS.n12768 DVSS.n12390 4.5005
R19827 DVSS.n12431 DVSS.n12359 4.5005
R19828 DVSS.n12431 DVSS.n12360 4.5005
R19829 DVSS.n12768 DVSS.n12431 4.5005
R19830 DVSS.n12389 DVSS.n12359 4.5005
R19831 DVSS.n12389 DVSS.n12360 4.5005
R19832 DVSS.n12768 DVSS.n12389 4.5005
R19833 DVSS.n12432 DVSS.n12359 4.5005
R19834 DVSS.n12432 DVSS.n12360 4.5005
R19835 DVSS.n12768 DVSS.n12432 4.5005
R19836 DVSS.n12388 DVSS.n12359 4.5005
R19837 DVSS.n12388 DVSS.n12360 4.5005
R19838 DVSS.n12768 DVSS.n12388 4.5005
R19839 DVSS.n12433 DVSS.n12359 4.5005
R19840 DVSS.n12433 DVSS.n12360 4.5005
R19841 DVSS.n12768 DVSS.n12433 4.5005
R19842 DVSS.n12387 DVSS.n12359 4.5005
R19843 DVSS.n12387 DVSS.n12360 4.5005
R19844 DVSS.n12768 DVSS.n12387 4.5005
R19845 DVSS.n12434 DVSS.n12359 4.5005
R19846 DVSS.n12434 DVSS.n12360 4.5005
R19847 DVSS.n12768 DVSS.n12434 4.5005
R19848 DVSS.n12386 DVSS.n12359 4.5005
R19849 DVSS.n12386 DVSS.n12360 4.5005
R19850 DVSS.n12768 DVSS.n12386 4.5005
R19851 DVSS.n12435 DVSS.n12359 4.5005
R19852 DVSS.n12435 DVSS.n12360 4.5005
R19853 DVSS.n12768 DVSS.n12435 4.5005
R19854 DVSS.n12385 DVSS.n12359 4.5005
R19855 DVSS.n12385 DVSS.n12360 4.5005
R19856 DVSS.n12768 DVSS.n12385 4.5005
R19857 DVSS.n12436 DVSS.n12359 4.5005
R19858 DVSS.n12436 DVSS.n12360 4.5005
R19859 DVSS.n12768 DVSS.n12436 4.5005
R19860 DVSS.n12384 DVSS.n12359 4.5005
R19861 DVSS.n12384 DVSS.n12360 4.5005
R19862 DVSS.n12768 DVSS.n12384 4.5005
R19863 DVSS.n12437 DVSS.n12359 4.5005
R19864 DVSS.n12437 DVSS.n12360 4.5005
R19865 DVSS.n12768 DVSS.n12437 4.5005
R19866 DVSS.n12383 DVSS.n12359 4.5005
R19867 DVSS.n12383 DVSS.n12360 4.5005
R19868 DVSS.n12768 DVSS.n12383 4.5005
R19869 DVSS.n12438 DVSS.n12359 4.5005
R19870 DVSS.n12438 DVSS.n12360 4.5005
R19871 DVSS.n12768 DVSS.n12438 4.5005
R19872 DVSS.n12382 DVSS.n12359 4.5005
R19873 DVSS.n12382 DVSS.n12360 4.5005
R19874 DVSS.n12768 DVSS.n12382 4.5005
R19875 DVSS.n12439 DVSS.n12359 4.5005
R19876 DVSS.n12439 DVSS.n12360 4.5005
R19877 DVSS.n12768 DVSS.n12439 4.5005
R19878 DVSS.n12381 DVSS.n12359 4.5005
R19879 DVSS.n12381 DVSS.n12360 4.5005
R19880 DVSS.n12768 DVSS.n12381 4.5005
R19881 DVSS.n12440 DVSS.n12359 4.5005
R19882 DVSS.n12440 DVSS.n12360 4.5005
R19883 DVSS.n12768 DVSS.n12440 4.5005
R19884 DVSS.n12380 DVSS.n12359 4.5005
R19885 DVSS.n12380 DVSS.n12360 4.5005
R19886 DVSS.n12768 DVSS.n12380 4.5005
R19887 DVSS.n12441 DVSS.n12359 4.5005
R19888 DVSS.n12441 DVSS.n12360 4.5005
R19889 DVSS.n12768 DVSS.n12441 4.5005
R19890 DVSS.n12379 DVSS.n12359 4.5005
R19891 DVSS.n12379 DVSS.n12360 4.5005
R19892 DVSS.n12768 DVSS.n12379 4.5005
R19893 DVSS.n12442 DVSS.n12359 4.5005
R19894 DVSS.n12442 DVSS.n12360 4.5005
R19895 DVSS.n12768 DVSS.n12442 4.5005
R19896 DVSS.n12378 DVSS.n12359 4.5005
R19897 DVSS.n12378 DVSS.n12360 4.5005
R19898 DVSS.n12768 DVSS.n12378 4.5005
R19899 DVSS.n12443 DVSS.n12359 4.5005
R19900 DVSS.n12443 DVSS.n12360 4.5005
R19901 DVSS.n12768 DVSS.n12443 4.5005
R19902 DVSS.n12377 DVSS.n12359 4.5005
R19903 DVSS.n12377 DVSS.n12360 4.5005
R19904 DVSS.n12768 DVSS.n12377 4.5005
R19905 DVSS.n12444 DVSS.n12359 4.5005
R19906 DVSS.n12444 DVSS.n12360 4.5005
R19907 DVSS.n12768 DVSS.n12444 4.5005
R19908 DVSS.n12376 DVSS.n12359 4.5005
R19909 DVSS.n12376 DVSS.n12360 4.5005
R19910 DVSS.n12768 DVSS.n12376 4.5005
R19911 DVSS.n12445 DVSS.n12359 4.5005
R19912 DVSS.n12445 DVSS.n12360 4.5005
R19913 DVSS.n12768 DVSS.n12445 4.5005
R19914 DVSS.n12375 DVSS.n12359 4.5005
R19915 DVSS.n12375 DVSS.n12360 4.5005
R19916 DVSS.n12768 DVSS.n12375 4.5005
R19917 DVSS.n12446 DVSS.n12359 4.5005
R19918 DVSS.n12446 DVSS.n12360 4.5005
R19919 DVSS.n12768 DVSS.n12446 4.5005
R19920 DVSS.n12374 DVSS.n12359 4.5005
R19921 DVSS.n12374 DVSS.n12360 4.5005
R19922 DVSS.n12768 DVSS.n12374 4.5005
R19923 DVSS.n12447 DVSS.n12359 4.5005
R19924 DVSS.n12447 DVSS.n12360 4.5005
R19925 DVSS.n12768 DVSS.n12447 4.5005
R19926 DVSS.n12373 DVSS.n12359 4.5005
R19927 DVSS.n12373 DVSS.n12360 4.5005
R19928 DVSS.n12768 DVSS.n12373 4.5005
R19929 DVSS.n12448 DVSS.n12359 4.5005
R19930 DVSS.n12448 DVSS.n12360 4.5005
R19931 DVSS.n12768 DVSS.n12448 4.5005
R19932 DVSS.n12372 DVSS.n12359 4.5005
R19933 DVSS.n12372 DVSS.n12360 4.5005
R19934 DVSS.n12768 DVSS.n12372 4.5005
R19935 DVSS.n12449 DVSS.n12359 4.5005
R19936 DVSS.n12449 DVSS.n12360 4.5005
R19937 DVSS.n12768 DVSS.n12449 4.5005
R19938 DVSS.n12371 DVSS.n12359 4.5005
R19939 DVSS.n12371 DVSS.n12360 4.5005
R19940 DVSS.n12768 DVSS.n12371 4.5005
R19941 DVSS.n12450 DVSS.n12359 4.5005
R19942 DVSS.n12450 DVSS.n12360 4.5005
R19943 DVSS.n12768 DVSS.n12450 4.5005
R19944 DVSS.n12370 DVSS.n12359 4.5005
R19945 DVSS.n12370 DVSS.n12360 4.5005
R19946 DVSS.n12768 DVSS.n12370 4.5005
R19947 DVSS.n12451 DVSS.n12359 4.5005
R19948 DVSS.n12451 DVSS.n12360 4.5005
R19949 DVSS.n12768 DVSS.n12451 4.5005
R19950 DVSS.n12369 DVSS.n12359 4.5005
R19951 DVSS.n12369 DVSS.n12360 4.5005
R19952 DVSS.n12768 DVSS.n12369 4.5005
R19953 DVSS.n12452 DVSS.n12359 4.5005
R19954 DVSS.n12452 DVSS.n12360 4.5005
R19955 DVSS.n12768 DVSS.n12452 4.5005
R19956 DVSS.n12368 DVSS.n12359 4.5005
R19957 DVSS.n12368 DVSS.n12360 4.5005
R19958 DVSS.n12768 DVSS.n12368 4.5005
R19959 DVSS.n12453 DVSS.n12359 4.5005
R19960 DVSS.n12453 DVSS.n12360 4.5005
R19961 DVSS.n12768 DVSS.n12453 4.5005
R19962 DVSS.n12367 DVSS.n12359 4.5005
R19963 DVSS.n12367 DVSS.n12360 4.5005
R19964 DVSS.n12768 DVSS.n12367 4.5005
R19965 DVSS.n12454 DVSS.n12359 4.5005
R19966 DVSS.n12454 DVSS.n12360 4.5005
R19967 DVSS.n12768 DVSS.n12454 4.5005
R19968 DVSS.n12366 DVSS.n12359 4.5005
R19969 DVSS.n12366 DVSS.n12360 4.5005
R19970 DVSS.n12768 DVSS.n12366 4.5005
R19971 DVSS.n12455 DVSS.n12359 4.5005
R19972 DVSS.n12455 DVSS.n12360 4.5005
R19973 DVSS.n12768 DVSS.n12455 4.5005
R19974 DVSS.n12365 DVSS.n12359 4.5005
R19975 DVSS.n12365 DVSS.n12360 4.5005
R19976 DVSS.n12768 DVSS.n12365 4.5005
R19977 DVSS.n12456 DVSS.n12359 4.5005
R19978 DVSS.n12456 DVSS.n12360 4.5005
R19979 DVSS.n12768 DVSS.n12456 4.5005
R19980 DVSS.n12364 DVSS.n12359 4.5005
R19981 DVSS.n12364 DVSS.n12360 4.5005
R19982 DVSS.n12768 DVSS.n12364 4.5005
R19983 DVSS.n12457 DVSS.n12359 4.5005
R19984 DVSS.n12457 DVSS.n12360 4.5005
R19985 DVSS.n12768 DVSS.n12457 4.5005
R19986 DVSS.n12363 DVSS.n12359 4.5005
R19987 DVSS.n12363 DVSS.n12360 4.5005
R19988 DVSS.n12768 DVSS.n12363 4.5005
R19989 DVSS.n12769 DVSS.n12359 4.5005
R19990 DVSS.n12769 DVSS.n12360 4.5005
R19991 DVSS.n12769 DVSS.n12768 4.5005
R19992 DVSS.n12362 DVSS.n12359 4.5005
R19993 DVSS.n12362 DVSS.n12360 4.5005
R19994 DVSS.n12553 DVSS.n12362 4.5005
R19995 DVSS.n12768 DVSS.n12362 4.5005
R19996 DVSS.n6257 DVSS.n6248 4.5005
R19997 DVSS.n6258 DVSS.n6248 4.5005
R19998 DVSS.n6256 DVSS.n6248 4.5005
R19999 DVSS.n6661 DVSS.n6248 4.5005
R20000 DVSS.n6248 DVSS.n6237 4.5005
R20001 DVSS.n12756 DVSS.n12354 4.5005
R20002 DVSS.n12758 DVSS.n12354 4.5005
R20003 DVSS.n12361 DVSS.n12354 4.5005
R20004 DVSS.n6659 DVSS.n6257 4.5005
R20005 DVSS.n6659 DVSS.n6258 4.5005
R20006 DVSS.n6659 DVSS.n6256 4.5005
R20007 DVSS.n6661 DVSS.n6659 4.5005
R20008 DVSS.n6659 DVSS.n6237 4.5005
R20009 DVSS.n12760 DVSS.n12752 4.5005
R20010 DVSS.n12757 DVSS.n12752 4.5005
R20011 DVSS.n12756 DVSS.n12752 4.5005
R20012 DVSS.n12758 DVSS.n12752 4.5005
R20013 DVSS.n12752 DVSS.n12361 4.5005
R20014 DVSS.n6662 DVSS.n6257 4.5005
R20015 DVSS.n6662 DVSS.n6258 4.5005
R20016 DVSS.n6662 DVSS.n6256 4.5005
R20017 DVSS.n6662 DVSS.n6661 4.5005
R20018 DVSS.n6662 DVSS.n6237 4.5005
R20019 DVSS.n12760 DVSS.n12749 4.5005
R20020 DVSS.n12757 DVSS.n12749 4.5005
R20021 DVSS.n12756 DVSS.n12749 4.5005
R20022 DVSS.n12758 DVSS.n12749 4.5005
R20023 DVSS.n12749 DVSS.n12361 4.5005
R20024 DVSS.n6660 DVSS.n6257 4.5005
R20025 DVSS.n6660 DVSS.n6258 4.5005
R20026 DVSS.n6660 DVSS.n6256 4.5005
R20027 DVSS.n6661 DVSS.n6660 4.5005
R20028 DVSS.n6660 DVSS.n6237 4.5005
R20029 DVSS.n12760 DVSS.n12759 4.5005
R20030 DVSS.n12759 DVSS.n12757 4.5005
R20031 DVSS.n12759 DVSS.n12756 4.5005
R20032 DVSS.n12759 DVSS.n12758 4.5005
R20033 DVSS.n12759 DVSS.n12361 4.5005
R20034 DVSS.n11980 DVSS.n11688 4.5005
R20035 DVSS.n11980 DVSS.n11979 4.5005
R20036 DVSS.n13324 DVSS.n13323 4.5005
R20037 DVSS.n13323 DVSS.n13322 4.5005
R20038 DVSS.n13338 DVSS.n13337 4.5005
R20039 DVSS.n13337 DVSS.n13336 4.5005
R20040 DVSS.n11102 DVSS.n10766 4.5005
R20041 DVSS.n10894 DVSS.n10766 4.5005
R20042 DVSS.n10754 DVSS.n1565 4.5005
R20043 DVSS.n10754 DVSS.n10753 4.5005
R20044 DVSS.n1959 DVSS.n1620 4.5005
R20045 DVSS.n1712 DVSS.n1620 4.5005
R20046 DVSS.n10475 DVSS.n2009 4.5005
R20047 DVSS.n10475 DVSS.n10474 4.5005
R20048 DVSS.n10166 DVSS.n2069 4.5005
R20049 DVSS.n10166 DVSS.n10165 4.5005
R20050 DVSS.n10141 DVSS.n2412 4.5005
R20051 DVSS.n10141 DVSS.n10140 4.5005
R20052 DVSS.n9860 DVSS.n2720 4.5005
R20053 DVSS.n10107 DVSS.n2720 4.5005
R20054 DVSS.n9757 DVSS.n2728 4.5005
R20055 DVSS.n9510 DVSS.n2728 4.5005
R20056 DVSS.n9455 DVSS.n2829 4.5005
R20057 DVSS.n9455 DVSS.n9454 4.5005
R20058 DVSS.n9185 DVSS.n9184 4.5005
R20059 DVSS.n9184 DVSS.n9183 4.5005
R20060 DVSS.n8967 DVSS.n3052 4.5005
R20061 DVSS.n8720 DVSS.n3052 4.5005
R20062 DVSS.n3153 DVSS.n3059 4.5005
R20063 DVSS.n3400 DVSS.n3059 4.5005
R20064 DVSS.n8602 DVSS.n8601 4.5005
R20065 DVSS.n8601 DVSS.n8600 4.5005
R20066 DVSS.n8588 DVSS.n3797 4.5005
R20067 DVSS.n8588 DVSS.n8587 4.5005
R20068 DVSS.n8318 DVSS.n8317 4.5005
R20069 DVSS.n8317 DVSS.n8316 4.5005
R20070 DVSS.n4109 DVSS.n4022 4.5005
R20071 DVSS.n4356 DVSS.n4022 4.5005
R20072 DVSS.n8088 DVSS.n4362 4.5005
R20073 DVSS.n7841 DVSS.n4362 4.5005
R20074 DVSS.n4805 DVSS.n4471 4.5005
R20075 DVSS.n4597 DVSS.n4471 4.5005
R20076 DVSS.n7793 DVSS.n4811 4.5005
R20077 DVSS.n7546 DVSS.n4811 4.5005
R20078 DVSS.n7442 DVSS.n4825 4.5005
R20079 DVSS.n7234 DVSS.n4825 4.5005
R20080 DVSS.n7102 DVSS.n4882 4.5005
R20081 DVSS.n7102 DVSS.n7101 4.5005
R20082 DVSS.n5272 DVSS.n5184 4.5005
R20083 DVSS.n5519 DVSS.n5184 4.5005
R20084 DVSS.n7059 DVSS.n5573 4.5005
R20085 DVSS.n7059 DVSS.n7058 4.5005
R20086 DVSS.n6656 DVSS.n6308 4.5005
R20087 DVSS.n6308 DVSS.n6259 4.5005
R20088 DVSS.n6602 DVSS.n6308 4.5005
R20089 DVSS.n6654 DVSS.n6308 4.5005
R20090 DVSS.n6656 DVSS.n6311 4.5005
R20091 DVSS.n6602 DVSS.n6311 4.5005
R20092 DVSS.n6654 DVSS.n6311 4.5005
R20093 DVSS.n6656 DVSS.n6307 4.5005
R20094 DVSS.n6602 DVSS.n6307 4.5005
R20095 DVSS.n6654 DVSS.n6307 4.5005
R20096 DVSS.n6656 DVSS.n6313 4.5005
R20097 DVSS.n6602 DVSS.n6313 4.5005
R20098 DVSS.n6654 DVSS.n6313 4.5005
R20099 DVSS.n6656 DVSS.n6306 4.5005
R20100 DVSS.n6602 DVSS.n6306 4.5005
R20101 DVSS.n6654 DVSS.n6306 4.5005
R20102 DVSS.n6656 DVSS.n6315 4.5005
R20103 DVSS.n6602 DVSS.n6315 4.5005
R20104 DVSS.n6654 DVSS.n6315 4.5005
R20105 DVSS.n6656 DVSS.n6305 4.5005
R20106 DVSS.n6602 DVSS.n6305 4.5005
R20107 DVSS.n6654 DVSS.n6305 4.5005
R20108 DVSS.n6656 DVSS.n6317 4.5005
R20109 DVSS.n6602 DVSS.n6317 4.5005
R20110 DVSS.n6654 DVSS.n6317 4.5005
R20111 DVSS.n6656 DVSS.n6304 4.5005
R20112 DVSS.n6602 DVSS.n6304 4.5005
R20113 DVSS.n6654 DVSS.n6304 4.5005
R20114 DVSS.n6656 DVSS.n6319 4.5005
R20115 DVSS.n6602 DVSS.n6319 4.5005
R20116 DVSS.n6654 DVSS.n6319 4.5005
R20117 DVSS.n6656 DVSS.n6303 4.5005
R20118 DVSS.n6602 DVSS.n6303 4.5005
R20119 DVSS.n6654 DVSS.n6303 4.5005
R20120 DVSS.n6656 DVSS.n6321 4.5005
R20121 DVSS.n6602 DVSS.n6321 4.5005
R20122 DVSS.n6654 DVSS.n6321 4.5005
R20123 DVSS.n6656 DVSS.n6302 4.5005
R20124 DVSS.n6602 DVSS.n6302 4.5005
R20125 DVSS.n6654 DVSS.n6302 4.5005
R20126 DVSS.n6656 DVSS.n6323 4.5005
R20127 DVSS.n6602 DVSS.n6323 4.5005
R20128 DVSS.n6654 DVSS.n6323 4.5005
R20129 DVSS.n6656 DVSS.n6301 4.5005
R20130 DVSS.n6602 DVSS.n6301 4.5005
R20131 DVSS.n6654 DVSS.n6301 4.5005
R20132 DVSS.n6656 DVSS.n6325 4.5005
R20133 DVSS.n6602 DVSS.n6325 4.5005
R20134 DVSS.n6654 DVSS.n6325 4.5005
R20135 DVSS.n6656 DVSS.n6300 4.5005
R20136 DVSS.n6602 DVSS.n6300 4.5005
R20137 DVSS.n6654 DVSS.n6300 4.5005
R20138 DVSS.n6656 DVSS.n6327 4.5005
R20139 DVSS.n6602 DVSS.n6327 4.5005
R20140 DVSS.n6654 DVSS.n6327 4.5005
R20141 DVSS.n6656 DVSS.n6299 4.5005
R20142 DVSS.n6602 DVSS.n6299 4.5005
R20143 DVSS.n6654 DVSS.n6299 4.5005
R20144 DVSS.n6656 DVSS.n6329 4.5005
R20145 DVSS.n6602 DVSS.n6329 4.5005
R20146 DVSS.n6654 DVSS.n6329 4.5005
R20147 DVSS.n6656 DVSS.n6298 4.5005
R20148 DVSS.n6602 DVSS.n6298 4.5005
R20149 DVSS.n6654 DVSS.n6298 4.5005
R20150 DVSS.n6656 DVSS.n6331 4.5005
R20151 DVSS.n6602 DVSS.n6331 4.5005
R20152 DVSS.n6654 DVSS.n6331 4.5005
R20153 DVSS.n6656 DVSS.n6297 4.5005
R20154 DVSS.n6602 DVSS.n6297 4.5005
R20155 DVSS.n6654 DVSS.n6297 4.5005
R20156 DVSS.n6656 DVSS.n6333 4.5005
R20157 DVSS.n6602 DVSS.n6333 4.5005
R20158 DVSS.n6654 DVSS.n6333 4.5005
R20159 DVSS.n6656 DVSS.n6296 4.5005
R20160 DVSS.n6602 DVSS.n6296 4.5005
R20161 DVSS.n6654 DVSS.n6296 4.5005
R20162 DVSS.n6656 DVSS.n6335 4.5005
R20163 DVSS.n6602 DVSS.n6335 4.5005
R20164 DVSS.n6654 DVSS.n6335 4.5005
R20165 DVSS.n6656 DVSS.n6295 4.5005
R20166 DVSS.n6602 DVSS.n6295 4.5005
R20167 DVSS.n6654 DVSS.n6295 4.5005
R20168 DVSS.n6656 DVSS.n6337 4.5005
R20169 DVSS.n6602 DVSS.n6337 4.5005
R20170 DVSS.n6654 DVSS.n6337 4.5005
R20171 DVSS.n6656 DVSS.n6294 4.5005
R20172 DVSS.n6602 DVSS.n6294 4.5005
R20173 DVSS.n6654 DVSS.n6294 4.5005
R20174 DVSS.n6656 DVSS.n6339 4.5005
R20175 DVSS.n6602 DVSS.n6339 4.5005
R20176 DVSS.n6654 DVSS.n6339 4.5005
R20177 DVSS.n6656 DVSS.n6293 4.5005
R20178 DVSS.n6602 DVSS.n6293 4.5005
R20179 DVSS.n6654 DVSS.n6293 4.5005
R20180 DVSS.n6656 DVSS.n6341 4.5005
R20181 DVSS.n6602 DVSS.n6341 4.5005
R20182 DVSS.n6654 DVSS.n6341 4.5005
R20183 DVSS.n6656 DVSS.n6292 4.5005
R20184 DVSS.n6602 DVSS.n6292 4.5005
R20185 DVSS.n6654 DVSS.n6292 4.5005
R20186 DVSS.n6656 DVSS.n6343 4.5005
R20187 DVSS.n6602 DVSS.n6343 4.5005
R20188 DVSS.n6654 DVSS.n6343 4.5005
R20189 DVSS.n6656 DVSS.n6291 4.5005
R20190 DVSS.n6602 DVSS.n6291 4.5005
R20191 DVSS.n6654 DVSS.n6291 4.5005
R20192 DVSS.n6656 DVSS.n6345 4.5005
R20193 DVSS.n6602 DVSS.n6345 4.5005
R20194 DVSS.n6654 DVSS.n6345 4.5005
R20195 DVSS.n6656 DVSS.n6290 4.5005
R20196 DVSS.n6602 DVSS.n6290 4.5005
R20197 DVSS.n6654 DVSS.n6290 4.5005
R20198 DVSS.n6656 DVSS.n6347 4.5005
R20199 DVSS.n6602 DVSS.n6347 4.5005
R20200 DVSS.n6654 DVSS.n6347 4.5005
R20201 DVSS.n6656 DVSS.n6289 4.5005
R20202 DVSS.n6602 DVSS.n6289 4.5005
R20203 DVSS.n6654 DVSS.n6289 4.5005
R20204 DVSS.n6656 DVSS.n6349 4.5005
R20205 DVSS.n6602 DVSS.n6349 4.5005
R20206 DVSS.n6654 DVSS.n6349 4.5005
R20207 DVSS.n6656 DVSS.n6288 4.5005
R20208 DVSS.n6602 DVSS.n6288 4.5005
R20209 DVSS.n6654 DVSS.n6288 4.5005
R20210 DVSS.n6656 DVSS.n6351 4.5005
R20211 DVSS.n6602 DVSS.n6351 4.5005
R20212 DVSS.n6654 DVSS.n6351 4.5005
R20213 DVSS.n6656 DVSS.n6287 4.5005
R20214 DVSS.n6602 DVSS.n6287 4.5005
R20215 DVSS.n6654 DVSS.n6287 4.5005
R20216 DVSS.n6656 DVSS.n6353 4.5005
R20217 DVSS.n6602 DVSS.n6353 4.5005
R20218 DVSS.n6654 DVSS.n6353 4.5005
R20219 DVSS.n6656 DVSS.n6286 4.5005
R20220 DVSS.n6602 DVSS.n6286 4.5005
R20221 DVSS.n6654 DVSS.n6286 4.5005
R20222 DVSS.n6656 DVSS.n6355 4.5005
R20223 DVSS.n6602 DVSS.n6355 4.5005
R20224 DVSS.n6654 DVSS.n6355 4.5005
R20225 DVSS.n6656 DVSS.n6285 4.5005
R20226 DVSS.n6602 DVSS.n6285 4.5005
R20227 DVSS.n6654 DVSS.n6285 4.5005
R20228 DVSS.n6656 DVSS.n6357 4.5005
R20229 DVSS.n6602 DVSS.n6357 4.5005
R20230 DVSS.n6654 DVSS.n6357 4.5005
R20231 DVSS.n6656 DVSS.n6284 4.5005
R20232 DVSS.n6602 DVSS.n6284 4.5005
R20233 DVSS.n6654 DVSS.n6284 4.5005
R20234 DVSS.n6656 DVSS.n6359 4.5005
R20235 DVSS.n6602 DVSS.n6359 4.5005
R20236 DVSS.n6654 DVSS.n6359 4.5005
R20237 DVSS.n6656 DVSS.n6283 4.5005
R20238 DVSS.n6602 DVSS.n6283 4.5005
R20239 DVSS.n6654 DVSS.n6283 4.5005
R20240 DVSS.n6656 DVSS.n6361 4.5005
R20241 DVSS.n6602 DVSS.n6361 4.5005
R20242 DVSS.n6654 DVSS.n6361 4.5005
R20243 DVSS.n6656 DVSS.n6282 4.5005
R20244 DVSS.n6602 DVSS.n6282 4.5005
R20245 DVSS.n6654 DVSS.n6282 4.5005
R20246 DVSS.n6656 DVSS.n6363 4.5005
R20247 DVSS.n6602 DVSS.n6363 4.5005
R20248 DVSS.n6654 DVSS.n6363 4.5005
R20249 DVSS.n6656 DVSS.n6281 4.5005
R20250 DVSS.n6602 DVSS.n6281 4.5005
R20251 DVSS.n6654 DVSS.n6281 4.5005
R20252 DVSS.n6656 DVSS.n6365 4.5005
R20253 DVSS.n6602 DVSS.n6365 4.5005
R20254 DVSS.n6654 DVSS.n6365 4.5005
R20255 DVSS.n6656 DVSS.n6280 4.5005
R20256 DVSS.n6602 DVSS.n6280 4.5005
R20257 DVSS.n6654 DVSS.n6280 4.5005
R20258 DVSS.n6656 DVSS.n6367 4.5005
R20259 DVSS.n6602 DVSS.n6367 4.5005
R20260 DVSS.n6654 DVSS.n6367 4.5005
R20261 DVSS.n6656 DVSS.n6279 4.5005
R20262 DVSS.n6602 DVSS.n6279 4.5005
R20263 DVSS.n6654 DVSS.n6279 4.5005
R20264 DVSS.n6656 DVSS.n6369 4.5005
R20265 DVSS.n6602 DVSS.n6369 4.5005
R20266 DVSS.n6654 DVSS.n6369 4.5005
R20267 DVSS.n6656 DVSS.n6278 4.5005
R20268 DVSS.n6602 DVSS.n6278 4.5005
R20269 DVSS.n6654 DVSS.n6278 4.5005
R20270 DVSS.n6656 DVSS.n6371 4.5005
R20271 DVSS.n6602 DVSS.n6371 4.5005
R20272 DVSS.n6654 DVSS.n6371 4.5005
R20273 DVSS.n6656 DVSS.n6277 4.5005
R20274 DVSS.n6602 DVSS.n6277 4.5005
R20275 DVSS.n6654 DVSS.n6277 4.5005
R20276 DVSS.n6656 DVSS.n6373 4.5005
R20277 DVSS.n6602 DVSS.n6373 4.5005
R20278 DVSS.n6654 DVSS.n6373 4.5005
R20279 DVSS.n6656 DVSS.n6276 4.5005
R20280 DVSS.n6602 DVSS.n6276 4.5005
R20281 DVSS.n6654 DVSS.n6276 4.5005
R20282 DVSS.n6656 DVSS.n6375 4.5005
R20283 DVSS.n6602 DVSS.n6375 4.5005
R20284 DVSS.n6654 DVSS.n6375 4.5005
R20285 DVSS.n6656 DVSS.n6275 4.5005
R20286 DVSS.n6602 DVSS.n6275 4.5005
R20287 DVSS.n6654 DVSS.n6275 4.5005
R20288 DVSS.n6656 DVSS.n6377 4.5005
R20289 DVSS.n6602 DVSS.n6377 4.5005
R20290 DVSS.n6654 DVSS.n6377 4.5005
R20291 DVSS.n6656 DVSS.n6274 4.5005
R20292 DVSS.n6602 DVSS.n6274 4.5005
R20293 DVSS.n6654 DVSS.n6274 4.5005
R20294 DVSS.n6656 DVSS.n6379 4.5005
R20295 DVSS.n6602 DVSS.n6379 4.5005
R20296 DVSS.n6654 DVSS.n6379 4.5005
R20297 DVSS.n6656 DVSS.n6273 4.5005
R20298 DVSS.n6602 DVSS.n6273 4.5005
R20299 DVSS.n6654 DVSS.n6273 4.5005
R20300 DVSS.n6656 DVSS.n6381 4.5005
R20301 DVSS.n6602 DVSS.n6381 4.5005
R20302 DVSS.n6654 DVSS.n6381 4.5005
R20303 DVSS.n6656 DVSS.n6272 4.5005
R20304 DVSS.n6602 DVSS.n6272 4.5005
R20305 DVSS.n6654 DVSS.n6272 4.5005
R20306 DVSS.n6656 DVSS.n6383 4.5005
R20307 DVSS.n6602 DVSS.n6383 4.5005
R20308 DVSS.n6654 DVSS.n6383 4.5005
R20309 DVSS.n6656 DVSS.n6271 4.5005
R20310 DVSS.n6602 DVSS.n6271 4.5005
R20311 DVSS.n6654 DVSS.n6271 4.5005
R20312 DVSS.n6656 DVSS.n6385 4.5005
R20313 DVSS.n6602 DVSS.n6385 4.5005
R20314 DVSS.n6654 DVSS.n6385 4.5005
R20315 DVSS.n6656 DVSS.n6270 4.5005
R20316 DVSS.n6602 DVSS.n6270 4.5005
R20317 DVSS.n6654 DVSS.n6270 4.5005
R20318 DVSS.n6656 DVSS.n6387 4.5005
R20319 DVSS.n6602 DVSS.n6387 4.5005
R20320 DVSS.n6654 DVSS.n6387 4.5005
R20321 DVSS.n6656 DVSS.n6269 4.5005
R20322 DVSS.n6602 DVSS.n6269 4.5005
R20323 DVSS.n6654 DVSS.n6269 4.5005
R20324 DVSS.n6656 DVSS.n6389 4.5005
R20325 DVSS.n6602 DVSS.n6389 4.5005
R20326 DVSS.n6654 DVSS.n6389 4.5005
R20327 DVSS.n6656 DVSS.n6268 4.5005
R20328 DVSS.n6602 DVSS.n6268 4.5005
R20329 DVSS.n6654 DVSS.n6268 4.5005
R20330 DVSS.n6656 DVSS.n6391 4.5005
R20331 DVSS.n6602 DVSS.n6391 4.5005
R20332 DVSS.n6654 DVSS.n6391 4.5005
R20333 DVSS.n6656 DVSS.n6267 4.5005
R20334 DVSS.n6602 DVSS.n6267 4.5005
R20335 DVSS.n6654 DVSS.n6267 4.5005
R20336 DVSS.n6656 DVSS.n6393 4.5005
R20337 DVSS.n6602 DVSS.n6393 4.5005
R20338 DVSS.n6654 DVSS.n6393 4.5005
R20339 DVSS.n6656 DVSS.n6266 4.5005
R20340 DVSS.n6602 DVSS.n6266 4.5005
R20341 DVSS.n6654 DVSS.n6266 4.5005
R20342 DVSS.n6656 DVSS.n6395 4.5005
R20343 DVSS.n6602 DVSS.n6395 4.5005
R20344 DVSS.n6654 DVSS.n6395 4.5005
R20345 DVSS.n6656 DVSS.n6265 4.5005
R20346 DVSS.n6602 DVSS.n6265 4.5005
R20347 DVSS.n6654 DVSS.n6265 4.5005
R20348 DVSS.n6656 DVSS.n6397 4.5005
R20349 DVSS.n6602 DVSS.n6397 4.5005
R20350 DVSS.n6654 DVSS.n6397 4.5005
R20351 DVSS.n6656 DVSS.n6264 4.5005
R20352 DVSS.n6602 DVSS.n6264 4.5005
R20353 DVSS.n6654 DVSS.n6264 4.5005
R20354 DVSS.n6656 DVSS.n6399 4.5005
R20355 DVSS.n6602 DVSS.n6399 4.5005
R20356 DVSS.n6654 DVSS.n6399 4.5005
R20357 DVSS.n6656 DVSS.n6263 4.5005
R20358 DVSS.n6602 DVSS.n6263 4.5005
R20359 DVSS.n6654 DVSS.n6263 4.5005
R20360 DVSS.n6656 DVSS.n6401 4.5005
R20361 DVSS.n6602 DVSS.n6401 4.5005
R20362 DVSS.n6654 DVSS.n6401 4.5005
R20363 DVSS.n6656 DVSS.n6262 4.5005
R20364 DVSS.n6602 DVSS.n6262 4.5005
R20365 DVSS.n6654 DVSS.n6262 4.5005
R20366 DVSS.n6656 DVSS.n6403 4.5005
R20367 DVSS.n6602 DVSS.n6403 4.5005
R20368 DVSS.n6654 DVSS.n6403 4.5005
R20369 DVSS.n6656 DVSS.n6261 4.5005
R20370 DVSS.n6602 DVSS.n6261 4.5005
R20371 DVSS.n6654 DVSS.n6261 4.5005
R20372 DVSS.n6656 DVSS.n6601 4.5005
R20373 DVSS.n6602 DVSS.n6601 4.5005
R20374 DVSS.n6654 DVSS.n6601 4.5005
R20375 DVSS.n6656 DVSS.n6260 4.5005
R20376 DVSS.n6260 DVSS.n6259 4.5005
R20377 DVSS.n6602 DVSS.n6260 4.5005
R20378 DVSS.n6654 DVSS.n6260 4.5005
R20379 DVSS.n12768 DVSS.n12767 4.5005
R20380 DVSS.n12767 DVSS.n12553 4.5005
R20381 DVSS.n12767 DVSS.n12360 4.5005
R20382 DVSS.n12767 DVSS.n12506 4.5005
R20383 DVSS.n12767 DVSS.n12359 4.5005
R20384 DVSS.n6656 DVSS.n6655 4.5005
R20385 DVSS.n6777 DVSS.n5878 4.5005
R20386 DVSS.n7025 DVSS.n5878 4.5005
R20387 DVSS.n12336 DVSS.n12044 4.5005
R20388 DVSS.n12336 DVSS.n12335 4.5005
R20389 DVSS.n5938 DVSS.n5888 4.5005
R20390 DVSS.n5983 DVSS.n5888 4.5005
R20391 DVSS.n12351 DVSS.n12345 4.5005
R20392 DVSS.n13103 DVSS.n12345 4.5005
R20393 DVSS.n13105 DVSS.n12345 4.5005
R20394 DVSS.n6666 DVSS.n6244 4.5005
R20395 DVSS.n6252 DVSS.n6244 4.5005
R20396 DVSS.n6664 DVSS.n6244 4.5005
R20397 DVSS.n12352 DVSS.n12349 4.5005
R20398 DVSS.n12775 DVSS.n12349 4.5005
R20399 DVSS.n12351 DVSS.n12349 4.5005
R20400 DVSS.n13103 DVSS.n12349 4.5005
R20401 DVSS.n13105 DVSS.n12349 4.5005
R20402 DVSS.n6663 DVSS.n6246 4.5005
R20403 DVSS.n6663 DVSS.n6252 4.5005
R20404 DVSS.n6664 DVSS.n6663 4.5005
R20405 DVSS.n12352 DVSS.n12344 4.5005
R20406 DVSS.n12775 DVSS.n12344 4.5005
R20407 DVSS.n12351 DVSS.n12344 4.5005
R20408 DVSS.n13103 DVSS.n12344 4.5005
R20409 DVSS.n13105 DVSS.n12344 4.5005
R20410 DVSS.n6666 DVSS.n6243 4.5005
R20411 DVSS.n6250 DVSS.n6243 4.5005
R20412 DVSS.n6246 DVSS.n6243 4.5005
R20413 DVSS.n6252 DVSS.n6243 4.5005
R20414 DVSS.n6664 DVSS.n6243 4.5005
R20415 DVSS.n13104 DVSS.n12352 4.5005
R20416 DVSS.n13104 DVSS.n12775 4.5005
R20417 DVSS.n13104 DVSS.n12351 4.5005
R20418 DVSS.n13104 DVSS.n13103 4.5005
R20419 DVSS.n13105 DVSS.n13104 4.5005
R20420 DVSS.n6666 DVSS.n6665 4.5005
R20421 DVSS.n6665 DVSS.n6250 4.5005
R20422 DVSS.n6665 DVSS.n6246 4.5005
R20423 DVSS.n6665 DVSS.n6252 4.5005
R20424 DVSS.n6665 DVSS.n6664 4.5005
R20425 DVSS.n19653 DVSS.n19138 4.5005
R20426 DVSS.n19656 DVSS.n19138 4.5005
R20427 DVSS.n19654 DVSS.n19653 4.5005
R20428 DVSS.n18113 DVSS.n18112 4.5005
R20429 DVSS.n18112 DVSS.n15622 4.5005
R20430 DVSS.n18114 DVSS.n15622 4.5005
R20431 DVSS.n18114 DVSS.n15623 4.5005
R20432 DVSS.n18114 DVSS.n15621 4.5005
R20433 DVSS.n18114 DVSS.n15624 4.5005
R20434 DVSS.n18114 DVSS.n15620 4.5005
R20435 DVSS.n18114 DVSS.n15625 4.5005
R20436 DVSS.n18114 DVSS.n15619 4.5005
R20437 DVSS.n18114 DVSS.n15626 4.5005
R20438 DVSS.n18114 DVSS.n15618 4.5005
R20439 DVSS.n18114 DVSS.n15627 4.5005
R20440 DVSS.n18114 DVSS.n15617 4.5005
R20441 DVSS.n18114 DVSS.n18113 4.5005
R20442 DVSS.n18151 DVSS.n15569 4.5005
R20443 DVSS.n15569 DVSS.n15549 4.5005
R20444 DVSS.n15569 DVSS.n15556 4.5005
R20445 DVSS.n15569 DVSS.n15554 4.5005
R20446 DVSS.n15569 DVSS.n15557 4.5005
R20447 DVSS.n15569 DVSS.n15553 4.5005
R20448 DVSS.n15569 DVSS.n15558 4.5005
R20449 DVSS.n15569 DVSS.n15560 4.5005
R20450 DVSS.n15569 DVSS.n15561 4.5005
R20451 DVSS.n18151 DVSS.n15573 4.5005
R20452 DVSS.n15573 DVSS.n15548 4.5005
R20453 DVSS.n15573 DVSS.n15562 4.5005
R20454 DVSS.n15573 DVSS.n15549 4.5005
R20455 DVSS.n15573 DVSS.n15556 4.5005
R20456 DVSS.n15573 DVSS.n15554 4.5005
R20457 DVSS.n15573 DVSS.n15557 4.5005
R20458 DVSS.n15573 DVSS.n15553 4.5005
R20459 DVSS.n15573 DVSS.n15558 4.5005
R20460 DVSS.n15573 DVSS.n15552 4.5005
R20461 DVSS.n15573 DVSS.n15559 4.5005
R20462 DVSS.n15573 DVSS.n15560 4.5005
R20463 DVSS.n15573 DVSS.n15561 4.5005
R20464 DVSS.n18151 DVSS.n15547 4.5005
R20465 DVSS.n15548 DVSS.n15547 4.5005
R20466 DVSS.n15562 DVSS.n15547 4.5005
R20467 DVSS.n15549 DVSS.n15547 4.5005
R20468 DVSS.n15556 DVSS.n15547 4.5005
R20469 DVSS.n15554 DVSS.n15547 4.5005
R20470 DVSS.n15557 DVSS.n15547 4.5005
R20471 DVSS.n15553 DVSS.n15547 4.5005
R20472 DVSS.n15558 DVSS.n15547 4.5005
R20473 DVSS.n15552 DVSS.n15547 4.5005
R20474 DVSS.n15559 DVSS.n15547 4.5005
R20475 DVSS.n15551 DVSS.n15547 4.5005
R20476 DVSS.n15560 DVSS.n15547 4.5005
R20477 DVSS.n15561 DVSS.n15547 4.5005
R20478 DVSS.n18152 DVSS.n15556 4.5005
R20479 DVSS.n18152 DVSS.n15554 4.5005
R20480 DVSS.n18152 DVSS.n15557 4.5005
R20481 DVSS.n18152 DVSS.n15553 4.5005
R20482 DVSS.n18152 DVSS.n15558 4.5005
R20483 DVSS.n18152 DVSS.n15552 4.5005
R20484 DVSS.n18152 DVSS.n15559 4.5005
R20485 DVSS.n18152 DVSS.n15551 4.5005
R20486 DVSS.n18152 DVSS.n15560 4.5005
R20487 DVSS.n18152 DVSS.n15550 4.5005
R20488 DVSS.n18152 DVSS.n15561 4.5005
R20489 DVSS.n18152 DVSS.n15549 4.5005
R20490 DVSS.n18152 DVSS.n15562 4.5005
R20491 DVSS.n18152 DVSS.n15548 4.5005
R20492 DVSS.n18152 DVSS.n18151 4.5005
R20493 DVSS.n15566 DVSS.n15556 4.5005
R20494 DVSS.n15566 DVSS.n15554 4.5005
R20495 DVSS.n15566 DVSS.n15557 4.5005
R20496 DVSS.n15566 DVSS.n15553 4.5005
R20497 DVSS.n15566 DVSS.n15558 4.5005
R20498 DVSS.n15566 DVSS.n15552 4.5005
R20499 DVSS.n15566 DVSS.n15559 4.5005
R20500 DVSS.n15566 DVSS.n15551 4.5005
R20501 DVSS.n15566 DVSS.n15560 4.5005
R20502 DVSS.n15566 DVSS.n15550 4.5005
R20503 DVSS.n15566 DVSS.n15561 4.5005
R20504 DVSS.n15566 DVSS.n15549 4.5005
R20505 DVSS.n15566 DVSS.n15562 4.5005
R20506 DVSS.n15566 DVSS.n15548 4.5005
R20507 DVSS.n18151 DVSS.n15566 4.5005
R20508 DVSS.n15574 DVSS.n15556 4.5005
R20509 DVSS.n15574 DVSS.n15554 4.5005
R20510 DVSS.n15574 DVSS.n15557 4.5005
R20511 DVSS.n15574 DVSS.n15553 4.5005
R20512 DVSS.n15574 DVSS.n15558 4.5005
R20513 DVSS.n15574 DVSS.n15552 4.5005
R20514 DVSS.n15574 DVSS.n15559 4.5005
R20515 DVSS.n15574 DVSS.n15551 4.5005
R20516 DVSS.n15574 DVSS.n15560 4.5005
R20517 DVSS.n15574 DVSS.n15550 4.5005
R20518 DVSS.n15574 DVSS.n15561 4.5005
R20519 DVSS.n15574 DVSS.n15549 4.5005
R20520 DVSS.n15574 DVSS.n15562 4.5005
R20521 DVSS.n15574 DVSS.n15548 4.5005
R20522 DVSS.n18151 DVSS.n15574 4.5005
R20523 DVSS.n15565 DVSS.n15556 4.5005
R20524 DVSS.n15565 DVSS.n15554 4.5005
R20525 DVSS.n15565 DVSS.n15557 4.5005
R20526 DVSS.n15565 DVSS.n15553 4.5005
R20527 DVSS.n15565 DVSS.n15558 4.5005
R20528 DVSS.n15565 DVSS.n15552 4.5005
R20529 DVSS.n15565 DVSS.n15559 4.5005
R20530 DVSS.n15565 DVSS.n15551 4.5005
R20531 DVSS.n15565 DVSS.n15560 4.5005
R20532 DVSS.n15565 DVSS.n15550 4.5005
R20533 DVSS.n15565 DVSS.n15561 4.5005
R20534 DVSS.n15565 DVSS.n15549 4.5005
R20535 DVSS.n15565 DVSS.n15562 4.5005
R20536 DVSS.n15565 DVSS.n15548 4.5005
R20537 DVSS.n18151 DVSS.n15565 4.5005
R20538 DVSS.n18148 DVSS.n15556 4.5005
R20539 DVSS.n18148 DVSS.n15554 4.5005
R20540 DVSS.n18148 DVSS.n15557 4.5005
R20541 DVSS.n18148 DVSS.n15553 4.5005
R20542 DVSS.n18148 DVSS.n15558 4.5005
R20543 DVSS.n18148 DVSS.n15552 4.5005
R20544 DVSS.n18148 DVSS.n15559 4.5005
R20545 DVSS.n18148 DVSS.n15551 4.5005
R20546 DVSS.n18148 DVSS.n15560 4.5005
R20547 DVSS.n18148 DVSS.n15550 4.5005
R20548 DVSS.n18148 DVSS.n15561 4.5005
R20549 DVSS.n18148 DVSS.n15549 4.5005
R20550 DVSS.n18148 DVSS.n15562 4.5005
R20551 DVSS.n18148 DVSS.n15548 4.5005
R20552 DVSS.n18151 DVSS.n18148 4.5005
R20553 DVSS.n15599 DVSS.n15589 4.5005
R20554 DVSS.n15597 DVSS.n15589 4.5005
R20555 DVSS.n15600 DVSS.n15589 4.5005
R20556 DVSS.n15596 DVSS.n15589 4.5005
R20557 DVSS.n15601 DVSS.n15589 4.5005
R20558 DVSS.n15594 DVSS.n15589 4.5005
R20559 DVSS.n15604 DVSS.n15589 4.5005
R20560 DVSS.n15593 DVSS.n15589 4.5005
R20561 DVSS.n15605 DVSS.n15589 4.5005
R20562 DVSS.n15592 DVSS.n15589 4.5005
R20563 DVSS.n18119 DVSS.n15589 4.5005
R20564 DVSS.n18120 DVSS.n15599 4.5005
R20565 DVSS.n18120 DVSS.n15597 4.5005
R20566 DVSS.n18120 DVSS.n15600 4.5005
R20567 DVSS.n18120 DVSS.n15596 4.5005
R20568 DVSS.n18120 DVSS.n15601 4.5005
R20569 DVSS.n18120 DVSS.n15595 4.5005
R20570 DVSS.n18120 DVSS.n15603 4.5005
R20571 DVSS.n18120 DVSS.n15594 4.5005
R20572 DVSS.n18120 DVSS.n15604 4.5005
R20573 DVSS.n18120 DVSS.n15593 4.5005
R20574 DVSS.n18120 DVSS.n15605 4.5005
R20575 DVSS.n18120 DVSS.n15592 4.5005
R20576 DVSS.n18120 DVSS.n15607 4.5005
R20577 DVSS.n18120 DVSS.n15591 4.5005
R20578 DVSS.n18120 DVSS.n18119 4.5005
R20579 DVSS.n15614 DVSS.n15599 4.5005
R20580 DVSS.n15614 DVSS.n15597 4.5005
R20581 DVSS.n15614 DVSS.n15600 4.5005
R20582 DVSS.n15614 DVSS.n15596 4.5005
R20583 DVSS.n15614 DVSS.n15601 4.5005
R20584 DVSS.n15614 DVSS.n15595 4.5005
R20585 DVSS.n15614 DVSS.n15603 4.5005
R20586 DVSS.n15614 DVSS.n15594 4.5005
R20587 DVSS.n15614 DVSS.n15604 4.5005
R20588 DVSS.n15614 DVSS.n15593 4.5005
R20589 DVSS.n15614 DVSS.n15605 4.5005
R20590 DVSS.n15614 DVSS.n15592 4.5005
R20591 DVSS.n15614 DVSS.n15607 4.5005
R20592 DVSS.n15614 DVSS.n15591 4.5005
R20593 DVSS.n18119 DVSS.n15614 4.5005
R20594 DVSS.n15612 DVSS.n15599 4.5005
R20595 DVSS.n15612 DVSS.n15597 4.5005
R20596 DVSS.n15612 DVSS.n15600 4.5005
R20597 DVSS.n15612 DVSS.n15596 4.5005
R20598 DVSS.n15612 DVSS.n15601 4.5005
R20599 DVSS.n15612 DVSS.n15595 4.5005
R20600 DVSS.n15612 DVSS.n15603 4.5005
R20601 DVSS.n15612 DVSS.n15594 4.5005
R20602 DVSS.n15612 DVSS.n15604 4.5005
R20603 DVSS.n15612 DVSS.n15593 4.5005
R20604 DVSS.n15612 DVSS.n15605 4.5005
R20605 DVSS.n15612 DVSS.n15592 4.5005
R20606 DVSS.n15612 DVSS.n15607 4.5005
R20607 DVSS.n15612 DVSS.n15591 4.5005
R20608 DVSS.n18119 DVSS.n15612 4.5005
R20609 DVSS.n15615 DVSS.n15599 4.5005
R20610 DVSS.n15615 DVSS.n15597 4.5005
R20611 DVSS.n15615 DVSS.n15600 4.5005
R20612 DVSS.n15615 DVSS.n15596 4.5005
R20613 DVSS.n15615 DVSS.n15601 4.5005
R20614 DVSS.n15615 DVSS.n15595 4.5005
R20615 DVSS.n15615 DVSS.n15603 4.5005
R20616 DVSS.n15615 DVSS.n15594 4.5005
R20617 DVSS.n15615 DVSS.n15604 4.5005
R20618 DVSS.n15615 DVSS.n15593 4.5005
R20619 DVSS.n15615 DVSS.n15605 4.5005
R20620 DVSS.n15615 DVSS.n15592 4.5005
R20621 DVSS.n15615 DVSS.n15607 4.5005
R20622 DVSS.n15615 DVSS.n15591 4.5005
R20623 DVSS.n18119 DVSS.n15615 4.5005
R20624 DVSS.n15611 DVSS.n15599 4.5005
R20625 DVSS.n15611 DVSS.n15597 4.5005
R20626 DVSS.n15611 DVSS.n15600 4.5005
R20627 DVSS.n15611 DVSS.n15596 4.5005
R20628 DVSS.n15611 DVSS.n15601 4.5005
R20629 DVSS.n15611 DVSS.n15595 4.5005
R20630 DVSS.n15611 DVSS.n15603 4.5005
R20631 DVSS.n15611 DVSS.n15594 4.5005
R20632 DVSS.n15611 DVSS.n15604 4.5005
R20633 DVSS.n15611 DVSS.n15593 4.5005
R20634 DVSS.n15611 DVSS.n15605 4.5005
R20635 DVSS.n15611 DVSS.n15592 4.5005
R20636 DVSS.n15611 DVSS.n15607 4.5005
R20637 DVSS.n15611 DVSS.n15591 4.5005
R20638 DVSS.n18119 DVSS.n15611 4.5005
R20639 DVSS.n15616 DVSS.n15599 4.5005
R20640 DVSS.n15616 DVSS.n15597 4.5005
R20641 DVSS.n15616 DVSS.n15600 4.5005
R20642 DVSS.n15616 DVSS.n15596 4.5005
R20643 DVSS.n15616 DVSS.n15601 4.5005
R20644 DVSS.n15616 DVSS.n15595 4.5005
R20645 DVSS.n15616 DVSS.n15603 4.5005
R20646 DVSS.n15616 DVSS.n15594 4.5005
R20647 DVSS.n15616 DVSS.n15604 4.5005
R20648 DVSS.n15616 DVSS.n15593 4.5005
R20649 DVSS.n15616 DVSS.n15605 4.5005
R20650 DVSS.n15616 DVSS.n15592 4.5005
R20651 DVSS.n15616 DVSS.n15607 4.5005
R20652 DVSS.n15616 DVSS.n15591 4.5005
R20653 DVSS.n18119 DVSS.n15616 4.5005
R20654 DVSS.n15610 DVSS.n15599 4.5005
R20655 DVSS.n15610 DVSS.n15597 4.5005
R20656 DVSS.n15610 DVSS.n15600 4.5005
R20657 DVSS.n15610 DVSS.n15596 4.5005
R20658 DVSS.n15610 DVSS.n15601 4.5005
R20659 DVSS.n15610 DVSS.n15595 4.5005
R20660 DVSS.n15610 DVSS.n15603 4.5005
R20661 DVSS.n15610 DVSS.n15594 4.5005
R20662 DVSS.n15610 DVSS.n15604 4.5005
R20663 DVSS.n15610 DVSS.n15593 4.5005
R20664 DVSS.n15610 DVSS.n15605 4.5005
R20665 DVSS.n15610 DVSS.n15592 4.5005
R20666 DVSS.n15610 DVSS.n15607 4.5005
R20667 DVSS.n15610 DVSS.n15591 4.5005
R20668 DVSS.n18119 DVSS.n15610 4.5005
R20669 DVSS.n18119 DVSS.n18116 4.5005
R20670 DVSS.n18116 DVSS.n15591 4.5005
R20671 DVSS.n18116 DVSS.n15607 4.5005
R20672 DVSS.n18116 DVSS.n15592 4.5005
R20673 DVSS.n18116 DVSS.n15599 4.5005
R20674 DVSS.n18116 DVSS.n15597 4.5005
R20675 DVSS.n18116 DVSS.n15600 4.5005
R20676 DVSS.n18116 DVSS.n15596 4.5005
R20677 DVSS.n18116 DVSS.n15601 4.5005
R20678 DVSS.n18116 DVSS.n15595 4.5005
R20679 DVSS.n18116 DVSS.n15603 4.5005
R20680 DVSS.n18116 DVSS.n15594 4.5005
R20681 DVSS.n18116 DVSS.n15604 4.5005
R20682 DVSS.n18116 DVSS.n15605 4.5005
R20683 DVSS.n18119 DVSS.n15609 4.5005
R20684 DVSS.n15609 DVSS.n15591 4.5005
R20685 DVSS.n15609 DVSS.n15607 4.5005
R20686 DVSS.n15609 DVSS.n15592 4.5005
R20687 DVSS.n15609 DVSS.n15599 4.5005
R20688 DVSS.n15609 DVSS.n15597 4.5005
R20689 DVSS.n15609 DVSS.n15600 4.5005
R20690 DVSS.n15609 DVSS.n15596 4.5005
R20691 DVSS.n15609 DVSS.n15601 4.5005
R20692 DVSS.n15609 DVSS.n15595 4.5005
R20693 DVSS.n15609 DVSS.n15603 4.5005
R20694 DVSS.n15609 DVSS.n15604 4.5005
R20695 DVSS.n15609 DVSS.n15605 4.5005
R20696 DVSS.n18119 DVSS.n18118 4.5005
R20697 DVSS.n18118 DVSS.n15591 4.5005
R20698 DVSS.n18118 DVSS.n15607 4.5005
R20699 DVSS.n18118 DVSS.n15592 4.5005
R20700 DVSS.n18118 DVSS.n15599 4.5005
R20701 DVSS.n18118 DVSS.n15597 4.5005
R20702 DVSS.n18118 DVSS.n15600 4.5005
R20703 DVSS.n18118 DVSS.n15596 4.5005
R20704 DVSS.n18118 DVSS.n15601 4.5005
R20705 DVSS.n18118 DVSS.n15595 4.5005
R20706 DVSS.n18118 DVSS.n15603 4.5005
R20707 DVSS.n18118 DVSS.n15604 4.5005
R20708 DVSS.n18118 DVSS.n15593 4.5005
R20709 DVSS.n18118 DVSS.n15605 4.5005
R20710 DVSS.n15515 DVSS.n15498 4.5005
R20711 DVSS.n15515 DVSS.n15496 4.5005
R20712 DVSS.n15515 DVSS.n15500 4.5005
R20713 DVSS.n15515 DVSS.n15495 4.5005
R20714 DVSS.n15515 DVSS.n15501 4.5005
R20715 DVSS.n15515 DVSS.n15494 4.5005
R20716 DVSS.n15515 DVSS.n15502 4.5005
R20717 DVSS.n18201 DVSS.n15515 4.5005
R20718 DVSS.n15515 DVSS.n15504 4.5005
R20719 DVSS.n18205 DVSS.n15515 4.5005
R20720 DVSS.n15510 DVSS.n15498 4.5005
R20721 DVSS.n15510 DVSS.n15497 4.5005
R20722 DVSS.n15510 DVSS.n15499 4.5005
R20723 DVSS.n15510 DVSS.n15496 4.5005
R20724 DVSS.n15510 DVSS.n15500 4.5005
R20725 DVSS.n15510 DVSS.n15495 4.5005
R20726 DVSS.n15510 DVSS.n15501 4.5005
R20727 DVSS.n15510 DVSS.n15494 4.5005
R20728 DVSS.n15510 DVSS.n15502 4.5005
R20729 DVSS.n15510 DVSS.n15493 4.5005
R20730 DVSS.n15510 DVSS.n15503 4.5005
R20731 DVSS.n15510 DVSS.n15504 4.5005
R20732 DVSS.n18205 DVSS.n15510 4.5005
R20733 DVSS.n15517 DVSS.n15498 4.5005
R20734 DVSS.n15517 DVSS.n15497 4.5005
R20735 DVSS.n15517 DVSS.n15499 4.5005
R20736 DVSS.n15517 DVSS.n15496 4.5005
R20737 DVSS.n15517 DVSS.n15500 4.5005
R20738 DVSS.n15517 DVSS.n15495 4.5005
R20739 DVSS.n15517 DVSS.n15501 4.5005
R20740 DVSS.n15517 DVSS.n15494 4.5005
R20741 DVSS.n15517 DVSS.n15502 4.5005
R20742 DVSS.n15517 DVSS.n15493 4.5005
R20743 DVSS.n15517 DVSS.n15503 4.5005
R20744 DVSS.n15517 DVSS.n15504 4.5005
R20745 DVSS.n18205 DVSS.n15517 4.5005
R20746 DVSS.n15509 DVSS.n15498 4.5005
R20747 DVSS.n15509 DVSS.n15497 4.5005
R20748 DVSS.n15509 DVSS.n15499 4.5005
R20749 DVSS.n15509 DVSS.n15496 4.5005
R20750 DVSS.n15509 DVSS.n15500 4.5005
R20751 DVSS.n15509 DVSS.n15495 4.5005
R20752 DVSS.n15509 DVSS.n15501 4.5005
R20753 DVSS.n15509 DVSS.n15494 4.5005
R20754 DVSS.n15509 DVSS.n15502 4.5005
R20755 DVSS.n15509 DVSS.n15493 4.5005
R20756 DVSS.n15509 DVSS.n15503 4.5005
R20757 DVSS.n15509 DVSS.n15504 4.5005
R20758 DVSS.n18205 DVSS.n15509 4.5005
R20759 DVSS.n15519 DVSS.n15498 4.5005
R20760 DVSS.n15519 DVSS.n15497 4.5005
R20761 DVSS.n15519 DVSS.n15499 4.5005
R20762 DVSS.n15519 DVSS.n15496 4.5005
R20763 DVSS.n15519 DVSS.n15500 4.5005
R20764 DVSS.n15519 DVSS.n15495 4.5005
R20765 DVSS.n15519 DVSS.n15501 4.5005
R20766 DVSS.n15519 DVSS.n15494 4.5005
R20767 DVSS.n15519 DVSS.n15502 4.5005
R20768 DVSS.n15519 DVSS.n15493 4.5005
R20769 DVSS.n15519 DVSS.n15503 4.5005
R20770 DVSS.n15519 DVSS.n15504 4.5005
R20771 DVSS.n18205 DVSS.n15519 4.5005
R20772 DVSS.n15508 DVSS.n15498 4.5005
R20773 DVSS.n15508 DVSS.n15497 4.5005
R20774 DVSS.n15508 DVSS.n15499 4.5005
R20775 DVSS.n15508 DVSS.n15496 4.5005
R20776 DVSS.n15508 DVSS.n15500 4.5005
R20777 DVSS.n15508 DVSS.n15495 4.5005
R20778 DVSS.n15508 DVSS.n15501 4.5005
R20779 DVSS.n15508 DVSS.n15494 4.5005
R20780 DVSS.n15508 DVSS.n15502 4.5005
R20781 DVSS.n15508 DVSS.n15493 4.5005
R20782 DVSS.n15508 DVSS.n15503 4.5005
R20783 DVSS.n15508 DVSS.n15504 4.5005
R20784 DVSS.n18205 DVSS.n15508 4.5005
R20785 DVSS.n15521 DVSS.n15498 4.5005
R20786 DVSS.n15521 DVSS.n15497 4.5005
R20787 DVSS.n15521 DVSS.n15499 4.5005
R20788 DVSS.n15521 DVSS.n15496 4.5005
R20789 DVSS.n15521 DVSS.n15500 4.5005
R20790 DVSS.n15521 DVSS.n15495 4.5005
R20791 DVSS.n15521 DVSS.n15501 4.5005
R20792 DVSS.n15521 DVSS.n15494 4.5005
R20793 DVSS.n15521 DVSS.n15502 4.5005
R20794 DVSS.n15521 DVSS.n15493 4.5005
R20795 DVSS.n15521 DVSS.n15503 4.5005
R20796 DVSS.n15521 DVSS.n15504 4.5005
R20797 DVSS.n18205 DVSS.n15521 4.5005
R20798 DVSS.n15507 DVSS.n15498 4.5005
R20799 DVSS.n15507 DVSS.n15497 4.5005
R20800 DVSS.n15507 DVSS.n15499 4.5005
R20801 DVSS.n15507 DVSS.n15496 4.5005
R20802 DVSS.n15507 DVSS.n15500 4.5005
R20803 DVSS.n15507 DVSS.n15495 4.5005
R20804 DVSS.n15507 DVSS.n15501 4.5005
R20805 DVSS.n15507 DVSS.n15494 4.5005
R20806 DVSS.n15507 DVSS.n15502 4.5005
R20807 DVSS.n15507 DVSS.n15493 4.5005
R20808 DVSS.n15507 DVSS.n15503 4.5005
R20809 DVSS.n15507 DVSS.n15504 4.5005
R20810 DVSS.n18205 DVSS.n15507 4.5005
R20811 DVSS.n18204 DVSS.n15498 4.5005
R20812 DVSS.n18204 DVSS.n15497 4.5005
R20813 DVSS.n18204 DVSS.n15499 4.5005
R20814 DVSS.n18204 DVSS.n15496 4.5005
R20815 DVSS.n18204 DVSS.n15500 4.5005
R20816 DVSS.n18204 DVSS.n15495 4.5005
R20817 DVSS.n18204 DVSS.n15501 4.5005
R20818 DVSS.n18204 DVSS.n15494 4.5005
R20819 DVSS.n18204 DVSS.n15502 4.5005
R20820 DVSS.n18204 DVSS.n15493 4.5005
R20821 DVSS.n18204 DVSS.n15503 4.5005
R20822 DVSS.n18204 DVSS.n15504 4.5005
R20823 DVSS.n18205 DVSS.n18204 4.5005
R20824 DVSS.n15506 DVSS.n15498 4.5005
R20825 DVSS.n15506 DVSS.n15497 4.5005
R20826 DVSS.n15506 DVSS.n15499 4.5005
R20827 DVSS.n15506 DVSS.n15496 4.5005
R20828 DVSS.n15506 DVSS.n15500 4.5005
R20829 DVSS.n15506 DVSS.n15495 4.5005
R20830 DVSS.n15506 DVSS.n15501 4.5005
R20831 DVSS.n15506 DVSS.n15494 4.5005
R20832 DVSS.n15506 DVSS.n15502 4.5005
R20833 DVSS.n15506 DVSS.n15493 4.5005
R20834 DVSS.n15506 DVSS.n15503 4.5005
R20835 DVSS.n15506 DVSS.n15504 4.5005
R20836 DVSS.n18205 DVSS.n15506 4.5005
R20837 DVSS.n18206 DVSS.n15498 4.5005
R20838 DVSS.n18206 DVSS.n15497 4.5005
R20839 DVSS.n18206 DVSS.n15499 4.5005
R20840 DVSS.n18206 DVSS.n15496 4.5005
R20841 DVSS.n18206 DVSS.n15500 4.5005
R20842 DVSS.n18206 DVSS.n15495 4.5005
R20843 DVSS.n18206 DVSS.n15501 4.5005
R20844 DVSS.n18206 DVSS.n15494 4.5005
R20845 DVSS.n18206 DVSS.n15502 4.5005
R20846 DVSS.n18206 DVSS.n15493 4.5005
R20847 DVSS.n18206 DVSS.n15503 4.5005
R20848 DVSS.n18206 DVSS.n15504 4.5005
R20849 DVSS.n18206 DVSS.n15492 4.5005
R20850 DVSS.n18206 DVSS.n18205 4.5005
R20851 DVSS.n18224 DVSS.n18207 4.5005
R20852 DVSS.n18222 DVSS.n18207 4.5005
R20853 DVSS.n18227 DVSS.n18207 4.5005
R20854 DVSS.n18221 DVSS.n18207 4.5005
R20855 DVSS.n18228 DVSS.n18207 4.5005
R20856 DVSS.n18220 DVSS.n18207 4.5005
R20857 DVSS.n18229 DVSS.n18207 4.5005
R20858 DVSS.n18237 DVSS.n18207 4.5005
R20859 DVSS.n18274 DVSS.n18207 4.5005
R20860 DVSS.n18276 DVSS.n18207 4.5005
R20861 DVSS.n18224 DVSS.n15489 4.5005
R20862 DVSS.n18223 DVSS.n15489 4.5005
R20863 DVSS.n18226 DVSS.n15489 4.5005
R20864 DVSS.n18222 DVSS.n15489 4.5005
R20865 DVSS.n18227 DVSS.n15489 4.5005
R20866 DVSS.n18221 DVSS.n15489 4.5005
R20867 DVSS.n18228 DVSS.n15489 4.5005
R20868 DVSS.n18220 DVSS.n15489 4.5005
R20869 DVSS.n18229 DVSS.n15489 4.5005
R20870 DVSS.n18219 DVSS.n15489 4.5005
R20871 DVSS.n18231 DVSS.n15489 4.5005
R20872 DVSS.n18274 DVSS.n15489 4.5005
R20873 DVSS.n18276 DVSS.n15489 4.5005
R20874 DVSS.n18224 DVSS.n18208 4.5005
R20875 DVSS.n18223 DVSS.n18208 4.5005
R20876 DVSS.n18226 DVSS.n18208 4.5005
R20877 DVSS.n18222 DVSS.n18208 4.5005
R20878 DVSS.n18227 DVSS.n18208 4.5005
R20879 DVSS.n18221 DVSS.n18208 4.5005
R20880 DVSS.n18228 DVSS.n18208 4.5005
R20881 DVSS.n18220 DVSS.n18208 4.5005
R20882 DVSS.n18229 DVSS.n18208 4.5005
R20883 DVSS.n18219 DVSS.n18208 4.5005
R20884 DVSS.n18231 DVSS.n18208 4.5005
R20885 DVSS.n18274 DVSS.n18208 4.5005
R20886 DVSS.n18276 DVSS.n18208 4.5005
R20887 DVSS.n18224 DVSS.n15488 4.5005
R20888 DVSS.n18223 DVSS.n15488 4.5005
R20889 DVSS.n18226 DVSS.n15488 4.5005
R20890 DVSS.n18222 DVSS.n15488 4.5005
R20891 DVSS.n18227 DVSS.n15488 4.5005
R20892 DVSS.n18221 DVSS.n15488 4.5005
R20893 DVSS.n18228 DVSS.n15488 4.5005
R20894 DVSS.n18220 DVSS.n15488 4.5005
R20895 DVSS.n18229 DVSS.n15488 4.5005
R20896 DVSS.n18219 DVSS.n15488 4.5005
R20897 DVSS.n18231 DVSS.n15488 4.5005
R20898 DVSS.n18274 DVSS.n15488 4.5005
R20899 DVSS.n18276 DVSS.n15488 4.5005
R20900 DVSS.n18224 DVSS.n18209 4.5005
R20901 DVSS.n18223 DVSS.n18209 4.5005
R20902 DVSS.n18226 DVSS.n18209 4.5005
R20903 DVSS.n18222 DVSS.n18209 4.5005
R20904 DVSS.n18227 DVSS.n18209 4.5005
R20905 DVSS.n18221 DVSS.n18209 4.5005
R20906 DVSS.n18228 DVSS.n18209 4.5005
R20907 DVSS.n18220 DVSS.n18209 4.5005
R20908 DVSS.n18229 DVSS.n18209 4.5005
R20909 DVSS.n18219 DVSS.n18209 4.5005
R20910 DVSS.n18231 DVSS.n18209 4.5005
R20911 DVSS.n18274 DVSS.n18209 4.5005
R20912 DVSS.n18276 DVSS.n18209 4.5005
R20913 DVSS.n18224 DVSS.n15487 4.5005
R20914 DVSS.n18223 DVSS.n15487 4.5005
R20915 DVSS.n18226 DVSS.n15487 4.5005
R20916 DVSS.n18222 DVSS.n15487 4.5005
R20917 DVSS.n18227 DVSS.n15487 4.5005
R20918 DVSS.n18221 DVSS.n15487 4.5005
R20919 DVSS.n18228 DVSS.n15487 4.5005
R20920 DVSS.n18220 DVSS.n15487 4.5005
R20921 DVSS.n18229 DVSS.n15487 4.5005
R20922 DVSS.n18219 DVSS.n15487 4.5005
R20923 DVSS.n18231 DVSS.n15487 4.5005
R20924 DVSS.n18274 DVSS.n15487 4.5005
R20925 DVSS.n18276 DVSS.n15487 4.5005
R20926 DVSS.n18224 DVSS.n18210 4.5005
R20927 DVSS.n18223 DVSS.n18210 4.5005
R20928 DVSS.n18226 DVSS.n18210 4.5005
R20929 DVSS.n18222 DVSS.n18210 4.5005
R20930 DVSS.n18227 DVSS.n18210 4.5005
R20931 DVSS.n18221 DVSS.n18210 4.5005
R20932 DVSS.n18228 DVSS.n18210 4.5005
R20933 DVSS.n18220 DVSS.n18210 4.5005
R20934 DVSS.n18229 DVSS.n18210 4.5005
R20935 DVSS.n18219 DVSS.n18210 4.5005
R20936 DVSS.n18231 DVSS.n18210 4.5005
R20937 DVSS.n18274 DVSS.n18210 4.5005
R20938 DVSS.n18276 DVSS.n18210 4.5005
R20939 DVSS.n18224 DVSS.n15486 4.5005
R20940 DVSS.n18223 DVSS.n15486 4.5005
R20941 DVSS.n18226 DVSS.n15486 4.5005
R20942 DVSS.n18222 DVSS.n15486 4.5005
R20943 DVSS.n18227 DVSS.n15486 4.5005
R20944 DVSS.n18221 DVSS.n15486 4.5005
R20945 DVSS.n18228 DVSS.n15486 4.5005
R20946 DVSS.n18220 DVSS.n15486 4.5005
R20947 DVSS.n18229 DVSS.n15486 4.5005
R20948 DVSS.n18219 DVSS.n15486 4.5005
R20949 DVSS.n18231 DVSS.n15486 4.5005
R20950 DVSS.n18274 DVSS.n15486 4.5005
R20951 DVSS.n18276 DVSS.n15486 4.5005
R20952 DVSS.n18224 DVSS.n18211 4.5005
R20953 DVSS.n18223 DVSS.n18211 4.5005
R20954 DVSS.n18226 DVSS.n18211 4.5005
R20955 DVSS.n18222 DVSS.n18211 4.5005
R20956 DVSS.n18227 DVSS.n18211 4.5005
R20957 DVSS.n18221 DVSS.n18211 4.5005
R20958 DVSS.n18228 DVSS.n18211 4.5005
R20959 DVSS.n18220 DVSS.n18211 4.5005
R20960 DVSS.n18229 DVSS.n18211 4.5005
R20961 DVSS.n18219 DVSS.n18211 4.5005
R20962 DVSS.n18231 DVSS.n18211 4.5005
R20963 DVSS.n18274 DVSS.n18211 4.5005
R20964 DVSS.n18276 DVSS.n18211 4.5005
R20965 DVSS.n18224 DVSS.n15485 4.5005
R20966 DVSS.n18223 DVSS.n15485 4.5005
R20967 DVSS.n18226 DVSS.n15485 4.5005
R20968 DVSS.n18222 DVSS.n15485 4.5005
R20969 DVSS.n18227 DVSS.n15485 4.5005
R20970 DVSS.n18221 DVSS.n15485 4.5005
R20971 DVSS.n18228 DVSS.n15485 4.5005
R20972 DVSS.n18220 DVSS.n15485 4.5005
R20973 DVSS.n18229 DVSS.n15485 4.5005
R20974 DVSS.n18219 DVSS.n15485 4.5005
R20975 DVSS.n18231 DVSS.n15485 4.5005
R20976 DVSS.n18274 DVSS.n15485 4.5005
R20977 DVSS.n18276 DVSS.n15485 4.5005
R20978 DVSS.n18275 DVSS.n18224 4.5005
R20979 DVSS.n18275 DVSS.n18223 4.5005
R20980 DVSS.n18275 DVSS.n18226 4.5005
R20981 DVSS.n18275 DVSS.n18222 4.5005
R20982 DVSS.n18275 DVSS.n18227 4.5005
R20983 DVSS.n18275 DVSS.n18221 4.5005
R20984 DVSS.n18275 DVSS.n18228 4.5005
R20985 DVSS.n18275 DVSS.n18220 4.5005
R20986 DVSS.n18275 DVSS.n18229 4.5005
R20987 DVSS.n18275 DVSS.n18219 4.5005
R20988 DVSS.n18275 DVSS.n18231 4.5005
R20989 DVSS.n18275 DVSS.n18274 4.5005
R20990 DVSS.n18275 DVSS.n18218 4.5005
R20991 DVSS.n18276 DVSS.n18275 4.5005
R20992 DVSS.n15108 DVSS.n15093 4.5005
R20993 DVSS.n15106 DVSS.n15093 4.5005
R20994 DVSS.n15111 DVSS.n15093 4.5005
R20995 DVSS.n15105 DVSS.n15093 4.5005
R20996 DVSS.n15112 DVSS.n15093 4.5005
R20997 DVSS.n15104 DVSS.n15093 4.5005
R20998 DVSS.n15113 DVSS.n15093 4.5005
R20999 DVSS.n15118 DVSS.n15093 4.5005
R21000 DVSS.n19954 DVSS.n15093 4.5005
R21001 DVSS.n15093 DVSS.n15080 4.5005
R21002 DVSS.n15108 DVSS.n15090 4.5005
R21003 DVSS.n15107 DVSS.n15090 4.5005
R21004 DVSS.n15110 DVSS.n15090 4.5005
R21005 DVSS.n15106 DVSS.n15090 4.5005
R21006 DVSS.n15111 DVSS.n15090 4.5005
R21007 DVSS.n15105 DVSS.n15090 4.5005
R21008 DVSS.n15112 DVSS.n15090 4.5005
R21009 DVSS.n15104 DVSS.n15090 4.5005
R21010 DVSS.n15113 DVSS.n15090 4.5005
R21011 DVSS.n15103 DVSS.n15090 4.5005
R21012 DVSS.n19952 DVSS.n15090 4.5005
R21013 DVSS.n19954 DVSS.n15090 4.5005
R21014 DVSS.n15090 DVSS.n15080 4.5005
R21015 DVSS.n15108 DVSS.n15095 4.5005
R21016 DVSS.n15107 DVSS.n15095 4.5005
R21017 DVSS.n15110 DVSS.n15095 4.5005
R21018 DVSS.n15106 DVSS.n15095 4.5005
R21019 DVSS.n15111 DVSS.n15095 4.5005
R21020 DVSS.n15105 DVSS.n15095 4.5005
R21021 DVSS.n15112 DVSS.n15095 4.5005
R21022 DVSS.n15104 DVSS.n15095 4.5005
R21023 DVSS.n15113 DVSS.n15095 4.5005
R21024 DVSS.n15103 DVSS.n15095 4.5005
R21025 DVSS.n19952 DVSS.n15095 4.5005
R21026 DVSS.n19954 DVSS.n15095 4.5005
R21027 DVSS.n15095 DVSS.n15080 4.5005
R21028 DVSS.n15108 DVSS.n15089 4.5005
R21029 DVSS.n15107 DVSS.n15089 4.5005
R21030 DVSS.n15110 DVSS.n15089 4.5005
R21031 DVSS.n15106 DVSS.n15089 4.5005
R21032 DVSS.n15111 DVSS.n15089 4.5005
R21033 DVSS.n15105 DVSS.n15089 4.5005
R21034 DVSS.n15112 DVSS.n15089 4.5005
R21035 DVSS.n15104 DVSS.n15089 4.5005
R21036 DVSS.n15113 DVSS.n15089 4.5005
R21037 DVSS.n15103 DVSS.n15089 4.5005
R21038 DVSS.n19952 DVSS.n15089 4.5005
R21039 DVSS.n19954 DVSS.n15089 4.5005
R21040 DVSS.n15089 DVSS.n15080 4.5005
R21041 DVSS.n15108 DVSS.n15097 4.5005
R21042 DVSS.n15107 DVSS.n15097 4.5005
R21043 DVSS.n15110 DVSS.n15097 4.5005
R21044 DVSS.n15106 DVSS.n15097 4.5005
R21045 DVSS.n15111 DVSS.n15097 4.5005
R21046 DVSS.n15105 DVSS.n15097 4.5005
R21047 DVSS.n15112 DVSS.n15097 4.5005
R21048 DVSS.n15104 DVSS.n15097 4.5005
R21049 DVSS.n15113 DVSS.n15097 4.5005
R21050 DVSS.n15103 DVSS.n15097 4.5005
R21051 DVSS.n19952 DVSS.n15097 4.5005
R21052 DVSS.n19954 DVSS.n15097 4.5005
R21053 DVSS.n15097 DVSS.n15080 4.5005
R21054 DVSS.n15108 DVSS.n15088 4.5005
R21055 DVSS.n15107 DVSS.n15088 4.5005
R21056 DVSS.n15110 DVSS.n15088 4.5005
R21057 DVSS.n15106 DVSS.n15088 4.5005
R21058 DVSS.n15111 DVSS.n15088 4.5005
R21059 DVSS.n15105 DVSS.n15088 4.5005
R21060 DVSS.n15112 DVSS.n15088 4.5005
R21061 DVSS.n15104 DVSS.n15088 4.5005
R21062 DVSS.n15113 DVSS.n15088 4.5005
R21063 DVSS.n15103 DVSS.n15088 4.5005
R21064 DVSS.n19952 DVSS.n15088 4.5005
R21065 DVSS.n19954 DVSS.n15088 4.5005
R21066 DVSS.n15088 DVSS.n15080 4.5005
R21067 DVSS.n15108 DVSS.n15099 4.5005
R21068 DVSS.n15107 DVSS.n15099 4.5005
R21069 DVSS.n15110 DVSS.n15099 4.5005
R21070 DVSS.n15106 DVSS.n15099 4.5005
R21071 DVSS.n15111 DVSS.n15099 4.5005
R21072 DVSS.n15105 DVSS.n15099 4.5005
R21073 DVSS.n15112 DVSS.n15099 4.5005
R21074 DVSS.n15104 DVSS.n15099 4.5005
R21075 DVSS.n15113 DVSS.n15099 4.5005
R21076 DVSS.n15103 DVSS.n15099 4.5005
R21077 DVSS.n19952 DVSS.n15099 4.5005
R21078 DVSS.n19954 DVSS.n15099 4.5005
R21079 DVSS.n15099 DVSS.n15080 4.5005
R21080 DVSS.n15108 DVSS.n15087 4.5005
R21081 DVSS.n15107 DVSS.n15087 4.5005
R21082 DVSS.n15110 DVSS.n15087 4.5005
R21083 DVSS.n15106 DVSS.n15087 4.5005
R21084 DVSS.n15111 DVSS.n15087 4.5005
R21085 DVSS.n15105 DVSS.n15087 4.5005
R21086 DVSS.n15112 DVSS.n15087 4.5005
R21087 DVSS.n15104 DVSS.n15087 4.5005
R21088 DVSS.n15113 DVSS.n15087 4.5005
R21089 DVSS.n15103 DVSS.n15087 4.5005
R21090 DVSS.n19952 DVSS.n15087 4.5005
R21091 DVSS.n19954 DVSS.n15087 4.5005
R21092 DVSS.n15087 DVSS.n15080 4.5005
R21093 DVSS.n15108 DVSS.n15101 4.5005
R21094 DVSS.n15107 DVSS.n15101 4.5005
R21095 DVSS.n15110 DVSS.n15101 4.5005
R21096 DVSS.n15106 DVSS.n15101 4.5005
R21097 DVSS.n15111 DVSS.n15101 4.5005
R21098 DVSS.n15105 DVSS.n15101 4.5005
R21099 DVSS.n15112 DVSS.n15101 4.5005
R21100 DVSS.n15104 DVSS.n15101 4.5005
R21101 DVSS.n15113 DVSS.n15101 4.5005
R21102 DVSS.n15103 DVSS.n15101 4.5005
R21103 DVSS.n19952 DVSS.n15101 4.5005
R21104 DVSS.n19954 DVSS.n15101 4.5005
R21105 DVSS.n15101 DVSS.n15080 4.5005
R21106 DVSS.n15108 DVSS.n15086 4.5005
R21107 DVSS.n15107 DVSS.n15086 4.5005
R21108 DVSS.n15110 DVSS.n15086 4.5005
R21109 DVSS.n15106 DVSS.n15086 4.5005
R21110 DVSS.n15111 DVSS.n15086 4.5005
R21111 DVSS.n15105 DVSS.n15086 4.5005
R21112 DVSS.n15112 DVSS.n15086 4.5005
R21113 DVSS.n15104 DVSS.n15086 4.5005
R21114 DVSS.n15113 DVSS.n15086 4.5005
R21115 DVSS.n15103 DVSS.n15086 4.5005
R21116 DVSS.n19952 DVSS.n15086 4.5005
R21117 DVSS.n19954 DVSS.n15086 4.5005
R21118 DVSS.n15086 DVSS.n15080 4.5005
R21119 DVSS.n19953 DVSS.n15108 4.5005
R21120 DVSS.n19953 DVSS.n15107 4.5005
R21121 DVSS.n19953 DVSS.n15110 4.5005
R21122 DVSS.n19953 DVSS.n15106 4.5005
R21123 DVSS.n19953 DVSS.n15111 4.5005
R21124 DVSS.n19953 DVSS.n15105 4.5005
R21125 DVSS.n19953 DVSS.n15112 4.5005
R21126 DVSS.n19953 DVSS.n15104 4.5005
R21127 DVSS.n19953 DVSS.n15113 4.5005
R21128 DVSS.n19953 DVSS.n15103 4.5005
R21129 DVSS.n19953 DVSS.n19952 4.5005
R21130 DVSS.n19954 DVSS.n19953 4.5005
R21131 DVSS.n19953 DVSS.n15085 4.5005
R21132 DVSS.n19953 DVSS.n15080 4.5005
R21133 DVSS.n20978 DVSS.n14326 4.5005
R21134 DVSS.n14341 DVSS.n14326 4.5005
R21135 DVSS.n14345 DVSS.n14326 4.5005
R21136 DVSS.n14340 DVSS.n14326 4.5005
R21137 DVSS.n14346 DVSS.n14326 4.5005
R21138 DVSS.n14339 DVSS.n14326 4.5005
R21139 DVSS.n14347 DVSS.n14326 4.5005
R21140 DVSS.n20968 DVSS.n14326 4.5005
R21141 DVSS.n14350 DVSS.n14326 4.5005
R21142 DVSS.n20976 DVSS.n14326 4.5005
R21143 DVSS.n20978 DVSS.n14325 4.5005
R21144 DVSS.n14325 DVSS.n14320 4.5005
R21145 DVSS.n14344 DVSS.n14325 4.5005
R21146 DVSS.n14341 DVSS.n14325 4.5005
R21147 DVSS.n14345 DVSS.n14325 4.5005
R21148 DVSS.n14340 DVSS.n14325 4.5005
R21149 DVSS.n14346 DVSS.n14325 4.5005
R21150 DVSS.n14339 DVSS.n14325 4.5005
R21151 DVSS.n14347 DVSS.n14325 4.5005
R21152 DVSS.n14338 DVSS.n14325 4.5005
R21153 DVSS.n14349 DVSS.n14325 4.5005
R21154 DVSS.n14350 DVSS.n14325 4.5005
R21155 DVSS.n20976 DVSS.n14325 4.5005
R21156 DVSS.n20978 DVSS.n14327 4.5005
R21157 DVSS.n14327 DVSS.n14320 4.5005
R21158 DVSS.n14344 DVSS.n14327 4.5005
R21159 DVSS.n14341 DVSS.n14327 4.5005
R21160 DVSS.n14345 DVSS.n14327 4.5005
R21161 DVSS.n14340 DVSS.n14327 4.5005
R21162 DVSS.n14346 DVSS.n14327 4.5005
R21163 DVSS.n14339 DVSS.n14327 4.5005
R21164 DVSS.n14347 DVSS.n14327 4.5005
R21165 DVSS.n14338 DVSS.n14327 4.5005
R21166 DVSS.n14349 DVSS.n14327 4.5005
R21167 DVSS.n14350 DVSS.n14327 4.5005
R21168 DVSS.n20976 DVSS.n14327 4.5005
R21169 DVSS.n20978 DVSS.n14324 4.5005
R21170 DVSS.n14324 DVSS.n14320 4.5005
R21171 DVSS.n14344 DVSS.n14324 4.5005
R21172 DVSS.n14341 DVSS.n14324 4.5005
R21173 DVSS.n14345 DVSS.n14324 4.5005
R21174 DVSS.n14340 DVSS.n14324 4.5005
R21175 DVSS.n14346 DVSS.n14324 4.5005
R21176 DVSS.n14339 DVSS.n14324 4.5005
R21177 DVSS.n14347 DVSS.n14324 4.5005
R21178 DVSS.n14338 DVSS.n14324 4.5005
R21179 DVSS.n14349 DVSS.n14324 4.5005
R21180 DVSS.n14350 DVSS.n14324 4.5005
R21181 DVSS.n20976 DVSS.n14324 4.5005
R21182 DVSS.n20978 DVSS.n14328 4.5005
R21183 DVSS.n14328 DVSS.n14320 4.5005
R21184 DVSS.n14344 DVSS.n14328 4.5005
R21185 DVSS.n14341 DVSS.n14328 4.5005
R21186 DVSS.n14345 DVSS.n14328 4.5005
R21187 DVSS.n14340 DVSS.n14328 4.5005
R21188 DVSS.n14346 DVSS.n14328 4.5005
R21189 DVSS.n14339 DVSS.n14328 4.5005
R21190 DVSS.n14347 DVSS.n14328 4.5005
R21191 DVSS.n14338 DVSS.n14328 4.5005
R21192 DVSS.n14349 DVSS.n14328 4.5005
R21193 DVSS.n14350 DVSS.n14328 4.5005
R21194 DVSS.n20976 DVSS.n14328 4.5005
R21195 DVSS.n20978 DVSS.n14323 4.5005
R21196 DVSS.n14323 DVSS.n14320 4.5005
R21197 DVSS.n14344 DVSS.n14323 4.5005
R21198 DVSS.n14341 DVSS.n14323 4.5005
R21199 DVSS.n14345 DVSS.n14323 4.5005
R21200 DVSS.n14340 DVSS.n14323 4.5005
R21201 DVSS.n14346 DVSS.n14323 4.5005
R21202 DVSS.n14339 DVSS.n14323 4.5005
R21203 DVSS.n14347 DVSS.n14323 4.5005
R21204 DVSS.n14338 DVSS.n14323 4.5005
R21205 DVSS.n14349 DVSS.n14323 4.5005
R21206 DVSS.n14350 DVSS.n14323 4.5005
R21207 DVSS.n20976 DVSS.n14323 4.5005
R21208 DVSS.n20978 DVSS.n14329 4.5005
R21209 DVSS.n14329 DVSS.n14320 4.5005
R21210 DVSS.n14344 DVSS.n14329 4.5005
R21211 DVSS.n14341 DVSS.n14329 4.5005
R21212 DVSS.n14345 DVSS.n14329 4.5005
R21213 DVSS.n14340 DVSS.n14329 4.5005
R21214 DVSS.n14346 DVSS.n14329 4.5005
R21215 DVSS.n14339 DVSS.n14329 4.5005
R21216 DVSS.n14347 DVSS.n14329 4.5005
R21217 DVSS.n14338 DVSS.n14329 4.5005
R21218 DVSS.n14349 DVSS.n14329 4.5005
R21219 DVSS.n14350 DVSS.n14329 4.5005
R21220 DVSS.n20976 DVSS.n14329 4.5005
R21221 DVSS.n20978 DVSS.n14322 4.5005
R21222 DVSS.n14322 DVSS.n14320 4.5005
R21223 DVSS.n14344 DVSS.n14322 4.5005
R21224 DVSS.n14341 DVSS.n14322 4.5005
R21225 DVSS.n14345 DVSS.n14322 4.5005
R21226 DVSS.n14340 DVSS.n14322 4.5005
R21227 DVSS.n14346 DVSS.n14322 4.5005
R21228 DVSS.n14339 DVSS.n14322 4.5005
R21229 DVSS.n14347 DVSS.n14322 4.5005
R21230 DVSS.n14338 DVSS.n14322 4.5005
R21231 DVSS.n14349 DVSS.n14322 4.5005
R21232 DVSS.n14350 DVSS.n14322 4.5005
R21233 DVSS.n20976 DVSS.n14322 4.5005
R21234 DVSS.n20978 DVSS.n14330 4.5005
R21235 DVSS.n14330 DVSS.n14320 4.5005
R21236 DVSS.n14344 DVSS.n14330 4.5005
R21237 DVSS.n14341 DVSS.n14330 4.5005
R21238 DVSS.n14345 DVSS.n14330 4.5005
R21239 DVSS.n14340 DVSS.n14330 4.5005
R21240 DVSS.n14346 DVSS.n14330 4.5005
R21241 DVSS.n14339 DVSS.n14330 4.5005
R21242 DVSS.n14347 DVSS.n14330 4.5005
R21243 DVSS.n14338 DVSS.n14330 4.5005
R21244 DVSS.n14349 DVSS.n14330 4.5005
R21245 DVSS.n14350 DVSS.n14330 4.5005
R21246 DVSS.n20976 DVSS.n14330 4.5005
R21247 DVSS.n20978 DVSS.n14321 4.5005
R21248 DVSS.n14321 DVSS.n14320 4.5005
R21249 DVSS.n14344 DVSS.n14321 4.5005
R21250 DVSS.n14341 DVSS.n14321 4.5005
R21251 DVSS.n14345 DVSS.n14321 4.5005
R21252 DVSS.n14340 DVSS.n14321 4.5005
R21253 DVSS.n14346 DVSS.n14321 4.5005
R21254 DVSS.n14339 DVSS.n14321 4.5005
R21255 DVSS.n14347 DVSS.n14321 4.5005
R21256 DVSS.n14338 DVSS.n14321 4.5005
R21257 DVSS.n14349 DVSS.n14321 4.5005
R21258 DVSS.n14350 DVSS.n14321 4.5005
R21259 DVSS.n20976 DVSS.n14321 4.5005
R21260 DVSS.n20978 DVSS.n20977 4.5005
R21261 DVSS.n20977 DVSS.n14320 4.5005
R21262 DVSS.n20977 DVSS.n14344 4.5005
R21263 DVSS.n20977 DVSS.n14341 4.5005
R21264 DVSS.n20977 DVSS.n14345 4.5005
R21265 DVSS.n20977 DVSS.n14340 4.5005
R21266 DVSS.n20977 DVSS.n14346 4.5005
R21267 DVSS.n20977 DVSS.n14339 4.5005
R21268 DVSS.n20977 DVSS.n14347 4.5005
R21269 DVSS.n20977 DVSS.n14338 4.5005
R21270 DVSS.n20977 DVSS.n14349 4.5005
R21271 DVSS.n20977 DVSS.n14350 4.5005
R21272 DVSS.n20977 DVSS.n14337 4.5005
R21273 DVSS.n20977 DVSS.n20976 4.5005
R21274 DVSS.n14276 DVSS.n14258 4.5005
R21275 DVSS.n14276 DVSS.n14256 4.5005
R21276 DVSS.n14276 DVSS.n14260 4.5005
R21277 DVSS.n14276 DVSS.n14255 4.5005
R21278 DVSS.n14276 DVSS.n14261 4.5005
R21279 DVSS.n14276 DVSS.n14254 4.5005
R21280 DVSS.n14276 DVSS.n14262 4.5005
R21281 DVSS.n21047 DVSS.n14276 4.5005
R21282 DVSS.n21051 DVSS.n14276 4.5005
R21283 DVSS.n14276 DVSS.n14234 4.5005
R21284 DVSS.n14278 DVSS.n14258 4.5005
R21285 DVSS.n14278 DVSS.n14257 4.5005
R21286 DVSS.n14278 DVSS.n14259 4.5005
R21287 DVSS.n14278 DVSS.n14256 4.5005
R21288 DVSS.n14278 DVSS.n14260 4.5005
R21289 DVSS.n14278 DVSS.n14255 4.5005
R21290 DVSS.n14278 DVSS.n14261 4.5005
R21291 DVSS.n14278 DVSS.n14254 4.5005
R21292 DVSS.n14278 DVSS.n14262 4.5005
R21293 DVSS.n14278 DVSS.n14253 4.5005
R21294 DVSS.n14278 DVSS.n14263 4.5005
R21295 DVSS.n21051 DVSS.n14278 4.5005
R21296 DVSS.n14278 DVSS.n14234 4.5005
R21297 DVSS.n14273 DVSS.n14258 4.5005
R21298 DVSS.n14273 DVSS.n14257 4.5005
R21299 DVSS.n14273 DVSS.n14259 4.5005
R21300 DVSS.n14273 DVSS.n14256 4.5005
R21301 DVSS.n14273 DVSS.n14260 4.5005
R21302 DVSS.n14273 DVSS.n14255 4.5005
R21303 DVSS.n14273 DVSS.n14261 4.5005
R21304 DVSS.n14273 DVSS.n14254 4.5005
R21305 DVSS.n14273 DVSS.n14262 4.5005
R21306 DVSS.n14273 DVSS.n14253 4.5005
R21307 DVSS.n14273 DVSS.n14263 4.5005
R21308 DVSS.n21051 DVSS.n14273 4.5005
R21309 DVSS.n14273 DVSS.n14234 4.5005
R21310 DVSS.n14279 DVSS.n14258 4.5005
R21311 DVSS.n14279 DVSS.n14257 4.5005
R21312 DVSS.n14279 DVSS.n14259 4.5005
R21313 DVSS.n14279 DVSS.n14256 4.5005
R21314 DVSS.n14279 DVSS.n14260 4.5005
R21315 DVSS.n14279 DVSS.n14255 4.5005
R21316 DVSS.n14279 DVSS.n14261 4.5005
R21317 DVSS.n14279 DVSS.n14254 4.5005
R21318 DVSS.n14279 DVSS.n14262 4.5005
R21319 DVSS.n14279 DVSS.n14253 4.5005
R21320 DVSS.n14279 DVSS.n14263 4.5005
R21321 DVSS.n21051 DVSS.n14279 4.5005
R21322 DVSS.n14279 DVSS.n14234 4.5005
R21323 DVSS.n14272 DVSS.n14258 4.5005
R21324 DVSS.n14272 DVSS.n14257 4.5005
R21325 DVSS.n14272 DVSS.n14259 4.5005
R21326 DVSS.n14272 DVSS.n14256 4.5005
R21327 DVSS.n14272 DVSS.n14260 4.5005
R21328 DVSS.n14272 DVSS.n14255 4.5005
R21329 DVSS.n14272 DVSS.n14261 4.5005
R21330 DVSS.n14272 DVSS.n14254 4.5005
R21331 DVSS.n14272 DVSS.n14262 4.5005
R21332 DVSS.n14272 DVSS.n14253 4.5005
R21333 DVSS.n14272 DVSS.n14263 4.5005
R21334 DVSS.n21051 DVSS.n14272 4.5005
R21335 DVSS.n14272 DVSS.n14234 4.5005
R21336 DVSS.n14280 DVSS.n14258 4.5005
R21337 DVSS.n14280 DVSS.n14257 4.5005
R21338 DVSS.n14280 DVSS.n14259 4.5005
R21339 DVSS.n14280 DVSS.n14256 4.5005
R21340 DVSS.n14280 DVSS.n14260 4.5005
R21341 DVSS.n14280 DVSS.n14255 4.5005
R21342 DVSS.n14280 DVSS.n14261 4.5005
R21343 DVSS.n14280 DVSS.n14254 4.5005
R21344 DVSS.n14280 DVSS.n14262 4.5005
R21345 DVSS.n14280 DVSS.n14253 4.5005
R21346 DVSS.n14280 DVSS.n14263 4.5005
R21347 DVSS.n21051 DVSS.n14280 4.5005
R21348 DVSS.n14280 DVSS.n14234 4.5005
R21349 DVSS.n14271 DVSS.n14258 4.5005
R21350 DVSS.n14271 DVSS.n14257 4.5005
R21351 DVSS.n14271 DVSS.n14259 4.5005
R21352 DVSS.n14271 DVSS.n14256 4.5005
R21353 DVSS.n14271 DVSS.n14260 4.5005
R21354 DVSS.n14271 DVSS.n14255 4.5005
R21355 DVSS.n14271 DVSS.n14261 4.5005
R21356 DVSS.n14271 DVSS.n14254 4.5005
R21357 DVSS.n14271 DVSS.n14262 4.5005
R21358 DVSS.n14271 DVSS.n14253 4.5005
R21359 DVSS.n14271 DVSS.n14263 4.5005
R21360 DVSS.n21051 DVSS.n14271 4.5005
R21361 DVSS.n14271 DVSS.n14234 4.5005
R21362 DVSS.n14281 DVSS.n14258 4.5005
R21363 DVSS.n14281 DVSS.n14257 4.5005
R21364 DVSS.n14281 DVSS.n14259 4.5005
R21365 DVSS.n14281 DVSS.n14256 4.5005
R21366 DVSS.n14281 DVSS.n14260 4.5005
R21367 DVSS.n14281 DVSS.n14255 4.5005
R21368 DVSS.n14281 DVSS.n14261 4.5005
R21369 DVSS.n14281 DVSS.n14254 4.5005
R21370 DVSS.n14281 DVSS.n14262 4.5005
R21371 DVSS.n14281 DVSS.n14253 4.5005
R21372 DVSS.n14281 DVSS.n14263 4.5005
R21373 DVSS.n21051 DVSS.n14281 4.5005
R21374 DVSS.n14281 DVSS.n14234 4.5005
R21375 DVSS.n14270 DVSS.n14258 4.5005
R21376 DVSS.n14270 DVSS.n14257 4.5005
R21377 DVSS.n14270 DVSS.n14259 4.5005
R21378 DVSS.n14270 DVSS.n14256 4.5005
R21379 DVSS.n14270 DVSS.n14260 4.5005
R21380 DVSS.n14270 DVSS.n14255 4.5005
R21381 DVSS.n14270 DVSS.n14261 4.5005
R21382 DVSS.n14270 DVSS.n14254 4.5005
R21383 DVSS.n14270 DVSS.n14262 4.5005
R21384 DVSS.n14270 DVSS.n14253 4.5005
R21385 DVSS.n14270 DVSS.n14263 4.5005
R21386 DVSS.n21051 DVSS.n14270 4.5005
R21387 DVSS.n14270 DVSS.n14234 4.5005
R21388 DVSS.n14282 DVSS.n14258 4.5005
R21389 DVSS.n14282 DVSS.n14257 4.5005
R21390 DVSS.n14282 DVSS.n14259 4.5005
R21391 DVSS.n14282 DVSS.n14256 4.5005
R21392 DVSS.n14282 DVSS.n14260 4.5005
R21393 DVSS.n14282 DVSS.n14255 4.5005
R21394 DVSS.n14282 DVSS.n14261 4.5005
R21395 DVSS.n14282 DVSS.n14254 4.5005
R21396 DVSS.n14282 DVSS.n14262 4.5005
R21397 DVSS.n14282 DVSS.n14253 4.5005
R21398 DVSS.n14282 DVSS.n14263 4.5005
R21399 DVSS.n21051 DVSS.n14282 4.5005
R21400 DVSS.n14282 DVSS.n14234 4.5005
R21401 DVSS.n14269 DVSS.n14258 4.5005
R21402 DVSS.n14269 DVSS.n14257 4.5005
R21403 DVSS.n14269 DVSS.n14259 4.5005
R21404 DVSS.n14269 DVSS.n14256 4.5005
R21405 DVSS.n14269 DVSS.n14260 4.5005
R21406 DVSS.n14269 DVSS.n14255 4.5005
R21407 DVSS.n14269 DVSS.n14261 4.5005
R21408 DVSS.n14269 DVSS.n14254 4.5005
R21409 DVSS.n14269 DVSS.n14262 4.5005
R21410 DVSS.n14269 DVSS.n14253 4.5005
R21411 DVSS.n14269 DVSS.n14263 4.5005
R21412 DVSS.n21051 DVSS.n14269 4.5005
R21413 DVSS.n14269 DVSS.n14234 4.5005
R21414 DVSS.n14283 DVSS.n14258 4.5005
R21415 DVSS.n14283 DVSS.n14257 4.5005
R21416 DVSS.n14283 DVSS.n14259 4.5005
R21417 DVSS.n14283 DVSS.n14256 4.5005
R21418 DVSS.n14283 DVSS.n14260 4.5005
R21419 DVSS.n14283 DVSS.n14255 4.5005
R21420 DVSS.n14283 DVSS.n14261 4.5005
R21421 DVSS.n14283 DVSS.n14254 4.5005
R21422 DVSS.n14283 DVSS.n14262 4.5005
R21423 DVSS.n14283 DVSS.n14253 4.5005
R21424 DVSS.n14283 DVSS.n14263 4.5005
R21425 DVSS.n21051 DVSS.n14283 4.5005
R21426 DVSS.n14283 DVSS.n14234 4.5005
R21427 DVSS.n14268 DVSS.n14258 4.5005
R21428 DVSS.n14268 DVSS.n14257 4.5005
R21429 DVSS.n14268 DVSS.n14259 4.5005
R21430 DVSS.n14268 DVSS.n14256 4.5005
R21431 DVSS.n14268 DVSS.n14260 4.5005
R21432 DVSS.n14268 DVSS.n14255 4.5005
R21433 DVSS.n14268 DVSS.n14261 4.5005
R21434 DVSS.n14268 DVSS.n14254 4.5005
R21435 DVSS.n14268 DVSS.n14262 4.5005
R21436 DVSS.n14268 DVSS.n14253 4.5005
R21437 DVSS.n14268 DVSS.n14263 4.5005
R21438 DVSS.n21051 DVSS.n14268 4.5005
R21439 DVSS.n14268 DVSS.n14234 4.5005
R21440 DVSS.n14284 DVSS.n14258 4.5005
R21441 DVSS.n14284 DVSS.n14257 4.5005
R21442 DVSS.n14284 DVSS.n14259 4.5005
R21443 DVSS.n14284 DVSS.n14256 4.5005
R21444 DVSS.n14284 DVSS.n14260 4.5005
R21445 DVSS.n14284 DVSS.n14255 4.5005
R21446 DVSS.n14284 DVSS.n14261 4.5005
R21447 DVSS.n14284 DVSS.n14254 4.5005
R21448 DVSS.n14284 DVSS.n14262 4.5005
R21449 DVSS.n14284 DVSS.n14253 4.5005
R21450 DVSS.n14284 DVSS.n14263 4.5005
R21451 DVSS.n21051 DVSS.n14284 4.5005
R21452 DVSS.n14284 DVSS.n14234 4.5005
R21453 DVSS.n14267 DVSS.n14258 4.5005
R21454 DVSS.n14267 DVSS.n14257 4.5005
R21455 DVSS.n14267 DVSS.n14259 4.5005
R21456 DVSS.n14267 DVSS.n14256 4.5005
R21457 DVSS.n14267 DVSS.n14260 4.5005
R21458 DVSS.n14267 DVSS.n14255 4.5005
R21459 DVSS.n14267 DVSS.n14261 4.5005
R21460 DVSS.n14267 DVSS.n14254 4.5005
R21461 DVSS.n14267 DVSS.n14262 4.5005
R21462 DVSS.n14267 DVSS.n14253 4.5005
R21463 DVSS.n14267 DVSS.n14263 4.5005
R21464 DVSS.n21051 DVSS.n14267 4.5005
R21465 DVSS.n14267 DVSS.n14234 4.5005
R21466 DVSS.n14285 DVSS.n14258 4.5005
R21467 DVSS.n14285 DVSS.n14257 4.5005
R21468 DVSS.n14285 DVSS.n14259 4.5005
R21469 DVSS.n14285 DVSS.n14256 4.5005
R21470 DVSS.n14285 DVSS.n14260 4.5005
R21471 DVSS.n14285 DVSS.n14255 4.5005
R21472 DVSS.n14285 DVSS.n14261 4.5005
R21473 DVSS.n14285 DVSS.n14254 4.5005
R21474 DVSS.n14285 DVSS.n14262 4.5005
R21475 DVSS.n14285 DVSS.n14253 4.5005
R21476 DVSS.n14285 DVSS.n14263 4.5005
R21477 DVSS.n21051 DVSS.n14285 4.5005
R21478 DVSS.n14285 DVSS.n14234 4.5005
R21479 DVSS.n14266 DVSS.n14258 4.5005
R21480 DVSS.n14266 DVSS.n14257 4.5005
R21481 DVSS.n14266 DVSS.n14259 4.5005
R21482 DVSS.n14266 DVSS.n14256 4.5005
R21483 DVSS.n14266 DVSS.n14260 4.5005
R21484 DVSS.n14266 DVSS.n14255 4.5005
R21485 DVSS.n14266 DVSS.n14261 4.5005
R21486 DVSS.n14266 DVSS.n14254 4.5005
R21487 DVSS.n14266 DVSS.n14262 4.5005
R21488 DVSS.n14266 DVSS.n14253 4.5005
R21489 DVSS.n14266 DVSS.n14263 4.5005
R21490 DVSS.n21051 DVSS.n14266 4.5005
R21491 DVSS.n14266 DVSS.n14234 4.5005
R21492 DVSS.n14286 DVSS.n14258 4.5005
R21493 DVSS.n14286 DVSS.n14257 4.5005
R21494 DVSS.n14286 DVSS.n14259 4.5005
R21495 DVSS.n14286 DVSS.n14256 4.5005
R21496 DVSS.n14286 DVSS.n14260 4.5005
R21497 DVSS.n14286 DVSS.n14255 4.5005
R21498 DVSS.n14286 DVSS.n14261 4.5005
R21499 DVSS.n14286 DVSS.n14254 4.5005
R21500 DVSS.n14286 DVSS.n14262 4.5005
R21501 DVSS.n14286 DVSS.n14253 4.5005
R21502 DVSS.n14286 DVSS.n14263 4.5005
R21503 DVSS.n21051 DVSS.n14286 4.5005
R21504 DVSS.n14286 DVSS.n14234 4.5005
R21505 DVSS.n14265 DVSS.n14258 4.5005
R21506 DVSS.n14265 DVSS.n14257 4.5005
R21507 DVSS.n14265 DVSS.n14259 4.5005
R21508 DVSS.n14265 DVSS.n14256 4.5005
R21509 DVSS.n14265 DVSS.n14260 4.5005
R21510 DVSS.n14265 DVSS.n14255 4.5005
R21511 DVSS.n14265 DVSS.n14261 4.5005
R21512 DVSS.n14265 DVSS.n14254 4.5005
R21513 DVSS.n14265 DVSS.n14262 4.5005
R21514 DVSS.n14265 DVSS.n14253 4.5005
R21515 DVSS.n14265 DVSS.n14263 4.5005
R21516 DVSS.n21051 DVSS.n14265 4.5005
R21517 DVSS.n14265 DVSS.n14234 4.5005
R21518 DVSS.n21049 DVSS.n14258 4.5005
R21519 DVSS.n21049 DVSS.n14257 4.5005
R21520 DVSS.n21049 DVSS.n14259 4.5005
R21521 DVSS.n21049 DVSS.n14256 4.5005
R21522 DVSS.n21049 DVSS.n14260 4.5005
R21523 DVSS.n21049 DVSS.n14255 4.5005
R21524 DVSS.n21049 DVSS.n14261 4.5005
R21525 DVSS.n21049 DVSS.n14254 4.5005
R21526 DVSS.n21049 DVSS.n14262 4.5005
R21527 DVSS.n21049 DVSS.n14253 4.5005
R21528 DVSS.n21049 DVSS.n14263 4.5005
R21529 DVSS.n21051 DVSS.n21049 4.5005
R21530 DVSS.n21049 DVSS.n14234 4.5005
R21531 DVSS.n14264 DVSS.n14258 4.5005
R21532 DVSS.n14264 DVSS.n14257 4.5005
R21533 DVSS.n14264 DVSS.n14259 4.5005
R21534 DVSS.n14264 DVSS.n14256 4.5005
R21535 DVSS.n14264 DVSS.n14260 4.5005
R21536 DVSS.n14264 DVSS.n14255 4.5005
R21537 DVSS.n14264 DVSS.n14261 4.5005
R21538 DVSS.n14264 DVSS.n14254 4.5005
R21539 DVSS.n14264 DVSS.n14262 4.5005
R21540 DVSS.n14264 DVSS.n14253 4.5005
R21541 DVSS.n14264 DVSS.n14263 4.5005
R21542 DVSS.n21051 DVSS.n14264 4.5005
R21543 DVSS.n14264 DVSS.n14234 4.5005
R21544 DVSS.n21050 DVSS.n14258 4.5005
R21545 DVSS.n21050 DVSS.n14257 4.5005
R21546 DVSS.n21050 DVSS.n14259 4.5005
R21547 DVSS.n21050 DVSS.n14256 4.5005
R21548 DVSS.n21050 DVSS.n14260 4.5005
R21549 DVSS.n21050 DVSS.n14255 4.5005
R21550 DVSS.n21050 DVSS.n14261 4.5005
R21551 DVSS.n21050 DVSS.n14254 4.5005
R21552 DVSS.n21050 DVSS.n14262 4.5005
R21553 DVSS.n21050 DVSS.n14253 4.5005
R21554 DVSS.n21050 DVSS.n14263 4.5005
R21555 DVSS.n21051 DVSS.n21050 4.5005
R21556 DVSS.n21050 DVSS.n14234 4.5005
R21557 DVSS.n21052 DVSS.n14258 4.5005
R21558 DVSS.n21052 DVSS.n14257 4.5005
R21559 DVSS.n21052 DVSS.n14259 4.5005
R21560 DVSS.n21052 DVSS.n14256 4.5005
R21561 DVSS.n21052 DVSS.n14260 4.5005
R21562 DVSS.n21052 DVSS.n14255 4.5005
R21563 DVSS.n21052 DVSS.n14261 4.5005
R21564 DVSS.n21052 DVSS.n14254 4.5005
R21565 DVSS.n21052 DVSS.n14262 4.5005
R21566 DVSS.n21052 DVSS.n14253 4.5005
R21567 DVSS.n21052 DVSS.n14263 4.5005
R21568 DVSS.n21052 DVSS.n21051 4.5005
R21569 DVSS.n21052 DVSS.n14234 4.5005
R21570 DVSS.n14258 DVSS.n14251 4.5005
R21571 DVSS.n14257 DVSS.n14251 4.5005
R21572 DVSS.n14259 DVSS.n14251 4.5005
R21573 DVSS.n14256 DVSS.n14251 4.5005
R21574 DVSS.n14260 DVSS.n14251 4.5005
R21575 DVSS.n14255 DVSS.n14251 4.5005
R21576 DVSS.n14261 DVSS.n14251 4.5005
R21577 DVSS.n14254 DVSS.n14251 4.5005
R21578 DVSS.n14262 DVSS.n14251 4.5005
R21579 DVSS.n14253 DVSS.n14251 4.5005
R21580 DVSS.n14263 DVSS.n14251 4.5005
R21581 DVSS.n21047 DVSS.n14251 4.5005
R21582 DVSS.n21051 DVSS.n14251 4.5005
R21583 DVSS.n14251 DVSS.n14234 4.5005
R21584 DVSS.n21432 DVSS.n13383 4.5005
R21585 DVSS.n13398 DVSS.n13383 4.5005
R21586 DVSS.n13403 DVSS.n13383 4.5005
R21587 DVSS.n13397 DVSS.n13383 4.5005
R21588 DVSS.n13404 DVSS.n13383 4.5005
R21589 DVSS.n13396 DVSS.n13383 4.5005
R21590 DVSS.n13405 DVSS.n13383 4.5005
R21591 DVSS.n21422 DVSS.n13383 4.5005
R21592 DVSS.n13408 DVSS.n13383 4.5005
R21593 DVSS.n21430 DVSS.n13383 4.5005
R21594 DVSS.n21432 DVSS.n13382 4.5005
R21595 DVSS.n13382 DVSS.n13377 4.5005
R21596 DVSS.n13402 DVSS.n13382 4.5005
R21597 DVSS.n13398 DVSS.n13382 4.5005
R21598 DVSS.n13403 DVSS.n13382 4.5005
R21599 DVSS.n13397 DVSS.n13382 4.5005
R21600 DVSS.n13404 DVSS.n13382 4.5005
R21601 DVSS.n13396 DVSS.n13382 4.5005
R21602 DVSS.n13405 DVSS.n13382 4.5005
R21603 DVSS.n13395 DVSS.n13382 4.5005
R21604 DVSS.n13407 DVSS.n13382 4.5005
R21605 DVSS.n13408 DVSS.n13382 4.5005
R21606 DVSS.n21430 DVSS.n13382 4.5005
R21607 DVSS.n21432 DVSS.n13384 4.5005
R21608 DVSS.n13384 DVSS.n13377 4.5005
R21609 DVSS.n13402 DVSS.n13384 4.5005
R21610 DVSS.n13398 DVSS.n13384 4.5005
R21611 DVSS.n13403 DVSS.n13384 4.5005
R21612 DVSS.n13397 DVSS.n13384 4.5005
R21613 DVSS.n13404 DVSS.n13384 4.5005
R21614 DVSS.n13396 DVSS.n13384 4.5005
R21615 DVSS.n13405 DVSS.n13384 4.5005
R21616 DVSS.n13395 DVSS.n13384 4.5005
R21617 DVSS.n13407 DVSS.n13384 4.5005
R21618 DVSS.n13408 DVSS.n13384 4.5005
R21619 DVSS.n21430 DVSS.n13384 4.5005
R21620 DVSS.n21432 DVSS.n13381 4.5005
R21621 DVSS.n13381 DVSS.n13377 4.5005
R21622 DVSS.n13402 DVSS.n13381 4.5005
R21623 DVSS.n13398 DVSS.n13381 4.5005
R21624 DVSS.n13403 DVSS.n13381 4.5005
R21625 DVSS.n13397 DVSS.n13381 4.5005
R21626 DVSS.n13404 DVSS.n13381 4.5005
R21627 DVSS.n13396 DVSS.n13381 4.5005
R21628 DVSS.n13405 DVSS.n13381 4.5005
R21629 DVSS.n13395 DVSS.n13381 4.5005
R21630 DVSS.n13407 DVSS.n13381 4.5005
R21631 DVSS.n13408 DVSS.n13381 4.5005
R21632 DVSS.n21430 DVSS.n13381 4.5005
R21633 DVSS.n21432 DVSS.n13385 4.5005
R21634 DVSS.n13385 DVSS.n13377 4.5005
R21635 DVSS.n13402 DVSS.n13385 4.5005
R21636 DVSS.n13398 DVSS.n13385 4.5005
R21637 DVSS.n13403 DVSS.n13385 4.5005
R21638 DVSS.n13397 DVSS.n13385 4.5005
R21639 DVSS.n13404 DVSS.n13385 4.5005
R21640 DVSS.n13396 DVSS.n13385 4.5005
R21641 DVSS.n13405 DVSS.n13385 4.5005
R21642 DVSS.n13395 DVSS.n13385 4.5005
R21643 DVSS.n13407 DVSS.n13385 4.5005
R21644 DVSS.n13408 DVSS.n13385 4.5005
R21645 DVSS.n21430 DVSS.n13385 4.5005
R21646 DVSS.n21432 DVSS.n13380 4.5005
R21647 DVSS.n13380 DVSS.n13377 4.5005
R21648 DVSS.n13402 DVSS.n13380 4.5005
R21649 DVSS.n13398 DVSS.n13380 4.5005
R21650 DVSS.n13403 DVSS.n13380 4.5005
R21651 DVSS.n13397 DVSS.n13380 4.5005
R21652 DVSS.n13404 DVSS.n13380 4.5005
R21653 DVSS.n13396 DVSS.n13380 4.5005
R21654 DVSS.n13405 DVSS.n13380 4.5005
R21655 DVSS.n13395 DVSS.n13380 4.5005
R21656 DVSS.n13407 DVSS.n13380 4.5005
R21657 DVSS.n13408 DVSS.n13380 4.5005
R21658 DVSS.n21430 DVSS.n13380 4.5005
R21659 DVSS.n21432 DVSS.n13386 4.5005
R21660 DVSS.n13386 DVSS.n13377 4.5005
R21661 DVSS.n13402 DVSS.n13386 4.5005
R21662 DVSS.n13398 DVSS.n13386 4.5005
R21663 DVSS.n13403 DVSS.n13386 4.5005
R21664 DVSS.n13397 DVSS.n13386 4.5005
R21665 DVSS.n13404 DVSS.n13386 4.5005
R21666 DVSS.n13396 DVSS.n13386 4.5005
R21667 DVSS.n13405 DVSS.n13386 4.5005
R21668 DVSS.n13395 DVSS.n13386 4.5005
R21669 DVSS.n13407 DVSS.n13386 4.5005
R21670 DVSS.n13408 DVSS.n13386 4.5005
R21671 DVSS.n21430 DVSS.n13386 4.5005
R21672 DVSS.n21432 DVSS.n13379 4.5005
R21673 DVSS.n13379 DVSS.n13377 4.5005
R21674 DVSS.n13402 DVSS.n13379 4.5005
R21675 DVSS.n13398 DVSS.n13379 4.5005
R21676 DVSS.n13403 DVSS.n13379 4.5005
R21677 DVSS.n13397 DVSS.n13379 4.5005
R21678 DVSS.n13404 DVSS.n13379 4.5005
R21679 DVSS.n13396 DVSS.n13379 4.5005
R21680 DVSS.n13405 DVSS.n13379 4.5005
R21681 DVSS.n13395 DVSS.n13379 4.5005
R21682 DVSS.n13407 DVSS.n13379 4.5005
R21683 DVSS.n13408 DVSS.n13379 4.5005
R21684 DVSS.n21430 DVSS.n13379 4.5005
R21685 DVSS.n21432 DVSS.n13387 4.5005
R21686 DVSS.n13387 DVSS.n13377 4.5005
R21687 DVSS.n13402 DVSS.n13387 4.5005
R21688 DVSS.n13398 DVSS.n13387 4.5005
R21689 DVSS.n13403 DVSS.n13387 4.5005
R21690 DVSS.n13397 DVSS.n13387 4.5005
R21691 DVSS.n13404 DVSS.n13387 4.5005
R21692 DVSS.n13396 DVSS.n13387 4.5005
R21693 DVSS.n13405 DVSS.n13387 4.5005
R21694 DVSS.n13395 DVSS.n13387 4.5005
R21695 DVSS.n13407 DVSS.n13387 4.5005
R21696 DVSS.n13408 DVSS.n13387 4.5005
R21697 DVSS.n21430 DVSS.n13387 4.5005
R21698 DVSS.n21432 DVSS.n13378 4.5005
R21699 DVSS.n13378 DVSS.n13377 4.5005
R21700 DVSS.n13402 DVSS.n13378 4.5005
R21701 DVSS.n13398 DVSS.n13378 4.5005
R21702 DVSS.n13403 DVSS.n13378 4.5005
R21703 DVSS.n13397 DVSS.n13378 4.5005
R21704 DVSS.n13404 DVSS.n13378 4.5005
R21705 DVSS.n13396 DVSS.n13378 4.5005
R21706 DVSS.n13405 DVSS.n13378 4.5005
R21707 DVSS.n13395 DVSS.n13378 4.5005
R21708 DVSS.n13407 DVSS.n13378 4.5005
R21709 DVSS.n13408 DVSS.n13378 4.5005
R21710 DVSS.n21430 DVSS.n13378 4.5005
R21711 DVSS.n21432 DVSS.n21431 4.5005
R21712 DVSS.n21431 DVSS.n13377 4.5005
R21713 DVSS.n21431 DVSS.n13402 4.5005
R21714 DVSS.n21431 DVSS.n13398 4.5005
R21715 DVSS.n21431 DVSS.n13403 4.5005
R21716 DVSS.n21431 DVSS.n13397 4.5005
R21717 DVSS.n21431 DVSS.n13404 4.5005
R21718 DVSS.n21431 DVSS.n13396 4.5005
R21719 DVSS.n21431 DVSS.n13405 4.5005
R21720 DVSS.n21431 DVSS.n13395 4.5005
R21721 DVSS.n21431 DVSS.n13407 4.5005
R21722 DVSS.n21431 DVSS.n13408 4.5005
R21723 DVSS.n21431 DVSS.n13394 4.5005
R21724 DVSS.n21431 DVSS.n21430 4.5005
R21725 DVSS.n15564 DVSS.n15561 4.5005
R21726 DVSS.n15564 DVSS.n15550 4.5005
R21727 DVSS.n15564 DVSS.n15560 4.5005
R21728 DVSS.n15564 DVSS.n15551 4.5005
R21729 DVSS.n15564 DVSS.n15559 4.5005
R21730 DVSS.n15564 DVSS.n15552 4.5005
R21731 DVSS.n15564 DVSS.n15558 4.5005
R21732 DVSS.n15564 DVSS.n15553 4.5005
R21733 DVSS.n15564 DVSS.n15557 4.5005
R21734 DVSS.n15564 DVSS.n15554 4.5005
R21735 DVSS.n15564 DVSS.n15556 4.5005
R21736 DVSS.n15564 DVSS.n15549 4.5005
R21737 DVSS.n15564 DVSS.n15562 4.5005
R21738 DVSS.n15564 DVSS.n15548 4.5005
R21739 DVSS.n18151 DVSS.n15564 4.5005
R21740 DVSS.n18151 DVSS.n18150 4.5005
R21741 DVSS.n18150 DVSS.n15561 4.5005
R21742 DVSS.n18150 DVSS.n15560 4.5005
R21743 DVSS.n18150 DVSS.n15551 4.5005
R21744 DVSS.n18150 DVSS.n15559 4.5005
R21745 DVSS.n18150 DVSS.n15552 4.5005
R21746 DVSS.n18150 DVSS.n15558 4.5005
R21747 DVSS.n18150 DVSS.n15553 4.5005
R21748 DVSS.n18150 DVSS.n15557 4.5005
R21749 DVSS.n18150 DVSS.n15554 4.5005
R21750 DVSS.n18150 DVSS.n15556 4.5005
R21751 DVSS.n18150 DVSS.n15549 4.5005
R21752 DVSS.n18150 DVSS.n15562 4.5005
R21753 DVSS.n18150 DVSS.n15548 4.5005
R21754 DVSS.n22879 DVSS.n464 4.5005
R21755 DVSS.n470 DVSS.n464 4.5005
R21756 DVSS.n22874 DVSS.n464 4.5005
R21757 DVSS.n471 DVSS.n464 4.5005
R21758 DVSS.n482 DVSS.n464 4.5005
R21759 DVSS.n472 DVSS.n464 4.5005
R21760 DVSS.n481 DVSS.n464 4.5005
R21761 DVSS.n474 DVSS.n464 4.5005
R21762 DVSS.n478 DVSS.n464 4.5005
R21763 DVSS.n477 DVSS.n464 4.5005
R21764 DVSS.n475 DVSS.n464 4.5005
R21765 DVSS.n22879 DVSS.n463 4.5005
R21766 DVSS.n463 DVSS.n458 4.5005
R21767 DVSS.n22877 DVSS.n463 4.5005
R21768 DVSS.n470 DVSS.n463 4.5005
R21769 DVSS.n22874 DVSS.n463 4.5005
R21770 DVSS.n471 DVSS.n463 4.5005
R21771 DVSS.n482 DVSS.n463 4.5005
R21772 DVSS.n472 DVSS.n463 4.5005
R21773 DVSS.n481 DVSS.n463 4.5005
R21774 DVSS.n473 DVSS.n463 4.5005
R21775 DVSS.n480 DVSS.n463 4.5005
R21776 DVSS.n474 DVSS.n463 4.5005
R21777 DVSS.n478 DVSS.n463 4.5005
R21778 DVSS.n477 DVSS.n463 4.5005
R21779 DVSS.n475 DVSS.n463 4.5005
R21780 DVSS.n477 DVSS.n465 4.5005
R21781 DVSS.n475 DVSS.n465 4.5005
R21782 DVSS.n478 DVSS.n465 4.5005
R21783 DVSS.n474 DVSS.n465 4.5005
R21784 DVSS.n480 DVSS.n465 4.5005
R21785 DVSS.n473 DVSS.n465 4.5005
R21786 DVSS.n481 DVSS.n465 4.5005
R21787 DVSS.n472 DVSS.n465 4.5005
R21788 DVSS.n482 DVSS.n465 4.5005
R21789 DVSS.n471 DVSS.n465 4.5005
R21790 DVSS.n22874 DVSS.n465 4.5005
R21791 DVSS.n470 DVSS.n465 4.5005
R21792 DVSS.n22877 DVSS.n465 4.5005
R21793 DVSS.n465 DVSS.n458 4.5005
R21794 DVSS.n22879 DVSS.n465 4.5005
R21795 DVSS.n477 DVSS.n462 4.5005
R21796 DVSS.n475 DVSS.n462 4.5005
R21797 DVSS.n478 DVSS.n462 4.5005
R21798 DVSS.n474 DVSS.n462 4.5005
R21799 DVSS.n480 DVSS.n462 4.5005
R21800 DVSS.n473 DVSS.n462 4.5005
R21801 DVSS.n481 DVSS.n462 4.5005
R21802 DVSS.n472 DVSS.n462 4.5005
R21803 DVSS.n482 DVSS.n462 4.5005
R21804 DVSS.n471 DVSS.n462 4.5005
R21805 DVSS.n22874 DVSS.n462 4.5005
R21806 DVSS.n470 DVSS.n462 4.5005
R21807 DVSS.n22877 DVSS.n462 4.5005
R21808 DVSS.n462 DVSS.n458 4.5005
R21809 DVSS.n22879 DVSS.n462 4.5005
R21810 DVSS.n477 DVSS.n466 4.5005
R21811 DVSS.n475 DVSS.n466 4.5005
R21812 DVSS.n478 DVSS.n466 4.5005
R21813 DVSS.n474 DVSS.n466 4.5005
R21814 DVSS.n480 DVSS.n466 4.5005
R21815 DVSS.n473 DVSS.n466 4.5005
R21816 DVSS.n481 DVSS.n466 4.5005
R21817 DVSS.n472 DVSS.n466 4.5005
R21818 DVSS.n482 DVSS.n466 4.5005
R21819 DVSS.n471 DVSS.n466 4.5005
R21820 DVSS.n22874 DVSS.n466 4.5005
R21821 DVSS.n470 DVSS.n466 4.5005
R21822 DVSS.n22877 DVSS.n466 4.5005
R21823 DVSS.n466 DVSS.n458 4.5005
R21824 DVSS.n22879 DVSS.n466 4.5005
R21825 DVSS.n477 DVSS.n461 4.5005
R21826 DVSS.n475 DVSS.n461 4.5005
R21827 DVSS.n478 DVSS.n461 4.5005
R21828 DVSS.n474 DVSS.n461 4.5005
R21829 DVSS.n480 DVSS.n461 4.5005
R21830 DVSS.n473 DVSS.n461 4.5005
R21831 DVSS.n481 DVSS.n461 4.5005
R21832 DVSS.n472 DVSS.n461 4.5005
R21833 DVSS.n482 DVSS.n461 4.5005
R21834 DVSS.n471 DVSS.n461 4.5005
R21835 DVSS.n22874 DVSS.n461 4.5005
R21836 DVSS.n470 DVSS.n461 4.5005
R21837 DVSS.n22877 DVSS.n461 4.5005
R21838 DVSS.n461 DVSS.n458 4.5005
R21839 DVSS.n22879 DVSS.n461 4.5005
R21840 DVSS.n22879 DVSS.n467 4.5005
R21841 DVSS.n467 DVSS.n458 4.5005
R21842 DVSS.n22877 DVSS.n467 4.5005
R21843 DVSS.n470 DVSS.n467 4.5005
R21844 DVSS.n22874 DVSS.n467 4.5005
R21845 DVSS.n471 DVSS.n467 4.5005
R21846 DVSS.n482 DVSS.n467 4.5005
R21847 DVSS.n472 DVSS.n467 4.5005
R21848 DVSS.n481 DVSS.n467 4.5005
R21849 DVSS.n473 DVSS.n467 4.5005
R21850 DVSS.n480 DVSS.n467 4.5005
R21851 DVSS.n474 DVSS.n467 4.5005
R21852 DVSS.n478 DVSS.n467 4.5005
R21853 DVSS.n477 DVSS.n467 4.5005
R21854 DVSS.n475 DVSS.n467 4.5005
R21855 DVSS.n22879 DVSS.n460 4.5005
R21856 DVSS.n460 DVSS.n458 4.5005
R21857 DVSS.n22877 DVSS.n460 4.5005
R21858 DVSS.n470 DVSS.n460 4.5005
R21859 DVSS.n22874 DVSS.n460 4.5005
R21860 DVSS.n471 DVSS.n460 4.5005
R21861 DVSS.n482 DVSS.n460 4.5005
R21862 DVSS.n472 DVSS.n460 4.5005
R21863 DVSS.n481 DVSS.n460 4.5005
R21864 DVSS.n473 DVSS.n460 4.5005
R21865 DVSS.n480 DVSS.n460 4.5005
R21866 DVSS.n474 DVSS.n460 4.5005
R21867 DVSS.n478 DVSS.n460 4.5005
R21868 DVSS.n477 DVSS.n460 4.5005
R21869 DVSS.n475 DVSS.n460 4.5005
R21870 DVSS.n22879 DVSS.n468 4.5005
R21871 DVSS.n468 DVSS.n458 4.5005
R21872 DVSS.n22877 DVSS.n468 4.5005
R21873 DVSS.n470 DVSS.n468 4.5005
R21874 DVSS.n22874 DVSS.n468 4.5005
R21875 DVSS.n471 DVSS.n468 4.5005
R21876 DVSS.n482 DVSS.n468 4.5005
R21877 DVSS.n472 DVSS.n468 4.5005
R21878 DVSS.n481 DVSS.n468 4.5005
R21879 DVSS.n473 DVSS.n468 4.5005
R21880 DVSS.n480 DVSS.n468 4.5005
R21881 DVSS.n474 DVSS.n468 4.5005
R21882 DVSS.n478 DVSS.n468 4.5005
R21883 DVSS.n477 DVSS.n468 4.5005
R21884 DVSS.n475 DVSS.n468 4.5005
R21885 DVSS.n477 DVSS.n459 4.5005
R21886 DVSS.n475 DVSS.n459 4.5005
R21887 DVSS.n478 DVSS.n459 4.5005
R21888 DVSS.n474 DVSS.n459 4.5005
R21889 DVSS.n480 DVSS.n459 4.5005
R21890 DVSS.n473 DVSS.n459 4.5005
R21891 DVSS.n481 DVSS.n459 4.5005
R21892 DVSS.n472 DVSS.n459 4.5005
R21893 DVSS.n482 DVSS.n459 4.5005
R21894 DVSS.n471 DVSS.n459 4.5005
R21895 DVSS.n22874 DVSS.n459 4.5005
R21896 DVSS.n470 DVSS.n459 4.5005
R21897 DVSS.n22877 DVSS.n459 4.5005
R21898 DVSS.n459 DVSS.n458 4.5005
R21899 DVSS.n22879 DVSS.n459 4.5005
R21900 DVSS.n22878 DVSS.n477 4.5005
R21901 DVSS.n22878 DVSS.n475 4.5005
R21902 DVSS.n22878 DVSS.n478 4.5005
R21903 DVSS.n22878 DVSS.n474 4.5005
R21904 DVSS.n22878 DVSS.n480 4.5005
R21905 DVSS.n22878 DVSS.n473 4.5005
R21906 DVSS.n22878 DVSS.n481 4.5005
R21907 DVSS.n22878 DVSS.n472 4.5005
R21908 DVSS.n22878 DVSS.n482 4.5005
R21909 DVSS.n22878 DVSS.n471 4.5005
R21910 DVSS.n22878 DVSS.n22874 4.5005
R21911 DVSS.n22878 DVSS.n470 4.5005
R21912 DVSS.n22878 DVSS.n22877 4.5005
R21913 DVSS.n22878 DVSS.n458 4.5005
R21914 DVSS.n22879 DVSS.n22878 4.5005
R21915 DVSS.n22671 DVSS.n707 4.5005
R21916 DVSS.n714 DVSS.n707 4.5005
R21917 DVSS.n726 DVSS.n707 4.5005
R21918 DVSS.n715 DVSS.n707 4.5005
R21919 DVSS.n725 DVSS.n707 4.5005
R21920 DVSS.n716 DVSS.n707 4.5005
R21921 DVSS.n724 DVSS.n707 4.5005
R21922 DVSS.n718 DVSS.n707 4.5005
R21923 DVSS.n721 DVSS.n707 4.5005
R21924 DVSS.n720 DVSS.n707 4.5005
R21925 DVSS.n22673 DVSS.n707 4.5005
R21926 DVSS.n22671 DVSS.n706 4.5005
R21927 DVSS.n713 DVSS.n706 4.5005
R21928 DVSS.n728 DVSS.n706 4.5005
R21929 DVSS.n714 DVSS.n706 4.5005
R21930 DVSS.n726 DVSS.n706 4.5005
R21931 DVSS.n715 DVSS.n706 4.5005
R21932 DVSS.n725 DVSS.n706 4.5005
R21933 DVSS.n716 DVSS.n706 4.5005
R21934 DVSS.n724 DVSS.n706 4.5005
R21935 DVSS.n717 DVSS.n706 4.5005
R21936 DVSS.n723 DVSS.n706 4.5005
R21937 DVSS.n718 DVSS.n706 4.5005
R21938 DVSS.n721 DVSS.n706 4.5005
R21939 DVSS.n720 DVSS.n706 4.5005
R21940 DVSS.n22673 DVSS.n706 4.5005
R21941 DVSS.n720 DVSS.n708 4.5005
R21942 DVSS.n22673 DVSS.n708 4.5005
R21943 DVSS.n720 DVSS.n705 4.5005
R21944 DVSS.n22673 DVSS.n705 4.5005
R21945 DVSS.n720 DVSS.n709 4.5005
R21946 DVSS.n22673 DVSS.n709 4.5005
R21947 DVSS.n22671 DVSS.n704 4.5005
R21948 DVSS.n713 DVSS.n704 4.5005
R21949 DVSS.n728 DVSS.n704 4.5005
R21950 DVSS.n714 DVSS.n704 4.5005
R21951 DVSS.n726 DVSS.n704 4.5005
R21952 DVSS.n715 DVSS.n704 4.5005
R21953 DVSS.n725 DVSS.n704 4.5005
R21954 DVSS.n716 DVSS.n704 4.5005
R21955 DVSS.n724 DVSS.n704 4.5005
R21956 DVSS.n717 DVSS.n704 4.5005
R21957 DVSS.n723 DVSS.n704 4.5005
R21958 DVSS.n718 DVSS.n704 4.5005
R21959 DVSS.n721 DVSS.n704 4.5005
R21960 DVSS.n720 DVSS.n704 4.5005
R21961 DVSS.n22673 DVSS.n704 4.5005
R21962 DVSS.n22671 DVSS.n710 4.5005
R21963 DVSS.n713 DVSS.n710 4.5005
R21964 DVSS.n728 DVSS.n710 4.5005
R21965 DVSS.n714 DVSS.n710 4.5005
R21966 DVSS.n726 DVSS.n710 4.5005
R21967 DVSS.n715 DVSS.n710 4.5005
R21968 DVSS.n725 DVSS.n710 4.5005
R21969 DVSS.n716 DVSS.n710 4.5005
R21970 DVSS.n724 DVSS.n710 4.5005
R21971 DVSS.n717 DVSS.n710 4.5005
R21972 DVSS.n723 DVSS.n710 4.5005
R21973 DVSS.n718 DVSS.n710 4.5005
R21974 DVSS.n721 DVSS.n710 4.5005
R21975 DVSS.n720 DVSS.n710 4.5005
R21976 DVSS.n22673 DVSS.n710 4.5005
R21977 DVSS.n22671 DVSS.n703 4.5005
R21978 DVSS.n713 DVSS.n703 4.5005
R21979 DVSS.n728 DVSS.n703 4.5005
R21980 DVSS.n714 DVSS.n703 4.5005
R21981 DVSS.n726 DVSS.n703 4.5005
R21982 DVSS.n715 DVSS.n703 4.5005
R21983 DVSS.n725 DVSS.n703 4.5005
R21984 DVSS.n716 DVSS.n703 4.5005
R21985 DVSS.n724 DVSS.n703 4.5005
R21986 DVSS.n717 DVSS.n703 4.5005
R21987 DVSS.n723 DVSS.n703 4.5005
R21988 DVSS.n718 DVSS.n703 4.5005
R21989 DVSS.n721 DVSS.n703 4.5005
R21990 DVSS.n720 DVSS.n703 4.5005
R21991 DVSS.n22673 DVSS.n703 4.5005
R21992 DVSS.n22671 DVSS.n711 4.5005
R21993 DVSS.n713 DVSS.n711 4.5005
R21994 DVSS.n728 DVSS.n711 4.5005
R21995 DVSS.n714 DVSS.n711 4.5005
R21996 DVSS.n726 DVSS.n711 4.5005
R21997 DVSS.n715 DVSS.n711 4.5005
R21998 DVSS.n725 DVSS.n711 4.5005
R21999 DVSS.n716 DVSS.n711 4.5005
R22000 DVSS.n724 DVSS.n711 4.5005
R22001 DVSS.n717 DVSS.n711 4.5005
R22002 DVSS.n723 DVSS.n711 4.5005
R22003 DVSS.n718 DVSS.n711 4.5005
R22004 DVSS.n721 DVSS.n711 4.5005
R22005 DVSS.n720 DVSS.n711 4.5005
R22006 DVSS.n22673 DVSS.n711 4.5005
R22007 DVSS.n720 DVSS.n702 4.5005
R22008 DVSS.n22673 DVSS.n702 4.5005
R22009 DVSS.n22672 DVSS.n720 4.5005
R22010 DVSS.n22673 DVSS.n22672 4.5005
R22011 DVSS.n22672 DVSS.n721 4.5005
R22012 DVSS.n22672 DVSS.n718 4.5005
R22013 DVSS.n22672 DVSS.n723 4.5005
R22014 DVSS.n22672 DVSS.n717 4.5005
R22015 DVSS.n22672 DVSS.n724 4.5005
R22016 DVSS.n22672 DVSS.n716 4.5005
R22017 DVSS.n22672 DVSS.n725 4.5005
R22018 DVSS.n22672 DVSS.n715 4.5005
R22019 DVSS.n22672 DVSS.n726 4.5005
R22020 DVSS.n22672 DVSS.n714 4.5005
R22021 DVSS.n22672 DVSS.n728 4.5005
R22022 DVSS.n22672 DVSS.n713 4.5005
R22023 DVSS.n22672 DVSS.n22671 4.5005
R22024 DVSS.n721 DVSS.n702 4.5005
R22025 DVSS.n718 DVSS.n702 4.5005
R22026 DVSS.n723 DVSS.n702 4.5005
R22027 DVSS.n717 DVSS.n702 4.5005
R22028 DVSS.n724 DVSS.n702 4.5005
R22029 DVSS.n716 DVSS.n702 4.5005
R22030 DVSS.n725 DVSS.n702 4.5005
R22031 DVSS.n715 DVSS.n702 4.5005
R22032 DVSS.n726 DVSS.n702 4.5005
R22033 DVSS.n714 DVSS.n702 4.5005
R22034 DVSS.n728 DVSS.n702 4.5005
R22035 DVSS.n713 DVSS.n702 4.5005
R22036 DVSS.n22671 DVSS.n702 4.5005
R22037 DVSS.n721 DVSS.n709 4.5005
R22038 DVSS.n718 DVSS.n709 4.5005
R22039 DVSS.n723 DVSS.n709 4.5005
R22040 DVSS.n717 DVSS.n709 4.5005
R22041 DVSS.n724 DVSS.n709 4.5005
R22042 DVSS.n716 DVSS.n709 4.5005
R22043 DVSS.n725 DVSS.n709 4.5005
R22044 DVSS.n715 DVSS.n709 4.5005
R22045 DVSS.n726 DVSS.n709 4.5005
R22046 DVSS.n714 DVSS.n709 4.5005
R22047 DVSS.n728 DVSS.n709 4.5005
R22048 DVSS.n713 DVSS.n709 4.5005
R22049 DVSS.n22671 DVSS.n709 4.5005
R22050 DVSS.n721 DVSS.n705 4.5005
R22051 DVSS.n718 DVSS.n705 4.5005
R22052 DVSS.n723 DVSS.n705 4.5005
R22053 DVSS.n717 DVSS.n705 4.5005
R22054 DVSS.n724 DVSS.n705 4.5005
R22055 DVSS.n716 DVSS.n705 4.5005
R22056 DVSS.n725 DVSS.n705 4.5005
R22057 DVSS.n715 DVSS.n705 4.5005
R22058 DVSS.n726 DVSS.n705 4.5005
R22059 DVSS.n714 DVSS.n705 4.5005
R22060 DVSS.n728 DVSS.n705 4.5005
R22061 DVSS.n713 DVSS.n705 4.5005
R22062 DVSS.n22671 DVSS.n705 4.5005
R22063 DVSS.n721 DVSS.n708 4.5005
R22064 DVSS.n718 DVSS.n708 4.5005
R22065 DVSS.n723 DVSS.n708 4.5005
R22066 DVSS.n717 DVSS.n708 4.5005
R22067 DVSS.n724 DVSS.n708 4.5005
R22068 DVSS.n716 DVSS.n708 4.5005
R22069 DVSS.n725 DVSS.n708 4.5005
R22070 DVSS.n715 DVSS.n708 4.5005
R22071 DVSS.n726 DVSS.n708 4.5005
R22072 DVSS.n714 DVSS.n708 4.5005
R22073 DVSS.n728 DVSS.n708 4.5005
R22074 DVSS.n713 DVSS.n708 4.5005
R22075 DVSS.n22671 DVSS.n708 4.5005
R22076 DVSS.n679 DVSS.n655 4.5005
R22077 DVSS.n681 DVSS.n655 4.5005
R22078 DVSS.n678 DVSS.n655 4.5005
R22079 DVSS.n682 DVSS.n655 4.5005
R22080 DVSS.n677 DVSS.n655 4.5005
R22081 DVSS.n685 DVSS.n655 4.5005
R22082 DVSS.n675 DVSS.n655 4.5005
R22083 DVSS.n686 DVSS.n655 4.5005
R22084 DVSS.n674 DVSS.n655 4.5005
R22085 DVSS.n22710 DVSS.n655 4.5005
R22086 DVSS.n673 DVSS.n655 4.5005
R22087 DVSS.n22713 DVSS.n655 4.5005
R22088 DVSS.n22715 DVSS.n655 4.5005
R22089 DVSS.n679 DVSS.n653 4.5005
R22090 DVSS.n681 DVSS.n653 4.5005
R22091 DVSS.n678 DVSS.n653 4.5005
R22092 DVSS.n682 DVSS.n653 4.5005
R22093 DVSS.n677 DVSS.n653 4.5005
R22094 DVSS.n684 DVSS.n653 4.5005
R22095 DVSS.n676 DVSS.n653 4.5005
R22096 DVSS.n685 DVSS.n653 4.5005
R22097 DVSS.n675 DVSS.n653 4.5005
R22098 DVSS.n686 DVSS.n653 4.5005
R22099 DVSS.n674 DVSS.n653 4.5005
R22100 DVSS.n22710 DVSS.n653 4.5005
R22101 DVSS.n22713 DVSS.n653 4.5005
R22102 DVSS.n22715 DVSS.n653 4.5005
R22103 DVSS.n679 DVSS.n657 4.5005
R22104 DVSS.n681 DVSS.n657 4.5005
R22105 DVSS.n678 DVSS.n657 4.5005
R22106 DVSS.n682 DVSS.n657 4.5005
R22107 DVSS.n677 DVSS.n657 4.5005
R22108 DVSS.n684 DVSS.n657 4.5005
R22109 DVSS.n676 DVSS.n657 4.5005
R22110 DVSS.n685 DVSS.n657 4.5005
R22111 DVSS.n675 DVSS.n657 4.5005
R22112 DVSS.n686 DVSS.n657 4.5005
R22113 DVSS.n674 DVSS.n657 4.5005
R22114 DVSS.n22710 DVSS.n657 4.5005
R22115 DVSS.n22713 DVSS.n657 4.5005
R22116 DVSS.n22715 DVSS.n657 4.5005
R22117 DVSS.n679 DVSS.n652 4.5005
R22118 DVSS.n681 DVSS.n652 4.5005
R22119 DVSS.n678 DVSS.n652 4.5005
R22120 DVSS.n682 DVSS.n652 4.5005
R22121 DVSS.n677 DVSS.n652 4.5005
R22122 DVSS.n684 DVSS.n652 4.5005
R22123 DVSS.n676 DVSS.n652 4.5005
R22124 DVSS.n685 DVSS.n652 4.5005
R22125 DVSS.n675 DVSS.n652 4.5005
R22126 DVSS.n686 DVSS.n652 4.5005
R22127 DVSS.n674 DVSS.n652 4.5005
R22128 DVSS.n22710 DVSS.n652 4.5005
R22129 DVSS.n673 DVSS.n652 4.5005
R22130 DVSS.n22713 DVSS.n652 4.5005
R22131 DVSS.n22715 DVSS.n652 4.5005
R22132 DVSS.n679 DVSS.n665 4.5005
R22133 DVSS.n681 DVSS.n665 4.5005
R22134 DVSS.n678 DVSS.n665 4.5005
R22135 DVSS.n682 DVSS.n665 4.5005
R22136 DVSS.n677 DVSS.n665 4.5005
R22137 DVSS.n684 DVSS.n665 4.5005
R22138 DVSS.n676 DVSS.n665 4.5005
R22139 DVSS.n685 DVSS.n665 4.5005
R22140 DVSS.n675 DVSS.n665 4.5005
R22141 DVSS.n686 DVSS.n665 4.5005
R22142 DVSS.n674 DVSS.n665 4.5005
R22143 DVSS.n22710 DVSS.n665 4.5005
R22144 DVSS.n673 DVSS.n665 4.5005
R22145 DVSS.n22713 DVSS.n665 4.5005
R22146 DVSS.n22715 DVSS.n665 4.5005
R22147 DVSS.n679 DVSS.n651 4.5005
R22148 DVSS.n681 DVSS.n651 4.5005
R22149 DVSS.n678 DVSS.n651 4.5005
R22150 DVSS.n682 DVSS.n651 4.5005
R22151 DVSS.n677 DVSS.n651 4.5005
R22152 DVSS.n684 DVSS.n651 4.5005
R22153 DVSS.n676 DVSS.n651 4.5005
R22154 DVSS.n685 DVSS.n651 4.5005
R22155 DVSS.n675 DVSS.n651 4.5005
R22156 DVSS.n686 DVSS.n651 4.5005
R22157 DVSS.n674 DVSS.n651 4.5005
R22158 DVSS.n22710 DVSS.n651 4.5005
R22159 DVSS.n22713 DVSS.n651 4.5005
R22160 DVSS.n22715 DVSS.n651 4.5005
R22161 DVSS.n679 DVSS.n666 4.5005
R22162 DVSS.n681 DVSS.n666 4.5005
R22163 DVSS.n678 DVSS.n666 4.5005
R22164 DVSS.n682 DVSS.n666 4.5005
R22165 DVSS.n677 DVSS.n666 4.5005
R22166 DVSS.n684 DVSS.n666 4.5005
R22167 DVSS.n676 DVSS.n666 4.5005
R22168 DVSS.n685 DVSS.n666 4.5005
R22169 DVSS.n675 DVSS.n666 4.5005
R22170 DVSS.n686 DVSS.n666 4.5005
R22171 DVSS.n674 DVSS.n666 4.5005
R22172 DVSS.n22710 DVSS.n666 4.5005
R22173 DVSS.n22715 DVSS.n666 4.5005
R22174 DVSS.n679 DVSS.n650 4.5005
R22175 DVSS.n681 DVSS.n650 4.5005
R22176 DVSS.n678 DVSS.n650 4.5005
R22177 DVSS.n682 DVSS.n650 4.5005
R22178 DVSS.n677 DVSS.n650 4.5005
R22179 DVSS.n684 DVSS.n650 4.5005
R22180 DVSS.n676 DVSS.n650 4.5005
R22181 DVSS.n685 DVSS.n650 4.5005
R22182 DVSS.n675 DVSS.n650 4.5005
R22183 DVSS.n686 DVSS.n650 4.5005
R22184 DVSS.n674 DVSS.n650 4.5005
R22185 DVSS.n22710 DVSS.n650 4.5005
R22186 DVSS.n22713 DVSS.n650 4.5005
R22187 DVSS.n22715 DVSS.n650 4.5005
R22188 DVSS.n679 DVSS.n668 4.5005
R22189 DVSS.n681 DVSS.n668 4.5005
R22190 DVSS.n678 DVSS.n668 4.5005
R22191 DVSS.n682 DVSS.n668 4.5005
R22192 DVSS.n677 DVSS.n668 4.5005
R22193 DVSS.n684 DVSS.n668 4.5005
R22194 DVSS.n676 DVSS.n668 4.5005
R22195 DVSS.n685 DVSS.n668 4.5005
R22196 DVSS.n675 DVSS.n668 4.5005
R22197 DVSS.n686 DVSS.n668 4.5005
R22198 DVSS.n674 DVSS.n668 4.5005
R22199 DVSS.n22710 DVSS.n668 4.5005
R22200 DVSS.n673 DVSS.n668 4.5005
R22201 DVSS.n22713 DVSS.n668 4.5005
R22202 DVSS.n22715 DVSS.n668 4.5005
R22203 DVSS.n679 DVSS.n649 4.5005
R22204 DVSS.n681 DVSS.n649 4.5005
R22205 DVSS.n678 DVSS.n649 4.5005
R22206 DVSS.n682 DVSS.n649 4.5005
R22207 DVSS.n677 DVSS.n649 4.5005
R22208 DVSS.n684 DVSS.n649 4.5005
R22209 DVSS.n676 DVSS.n649 4.5005
R22210 DVSS.n685 DVSS.n649 4.5005
R22211 DVSS.n675 DVSS.n649 4.5005
R22212 DVSS.n686 DVSS.n649 4.5005
R22213 DVSS.n674 DVSS.n649 4.5005
R22214 DVSS.n22710 DVSS.n649 4.5005
R22215 DVSS.n22713 DVSS.n649 4.5005
R22216 DVSS.n649 DVSS.n648 4.5005
R22217 DVSS.n22715 DVSS.n649 4.5005
R22218 DVSS.n22714 DVSS.n679 4.5005
R22219 DVSS.n22714 DVSS.n681 4.5005
R22220 DVSS.n22714 DVSS.n678 4.5005
R22221 DVSS.n22714 DVSS.n682 4.5005
R22222 DVSS.n22714 DVSS.n677 4.5005
R22223 DVSS.n22714 DVSS.n684 4.5005
R22224 DVSS.n22714 DVSS.n676 4.5005
R22225 DVSS.n22714 DVSS.n685 4.5005
R22226 DVSS.n22714 DVSS.n675 4.5005
R22227 DVSS.n22714 DVSS.n686 4.5005
R22228 DVSS.n22714 DVSS.n674 4.5005
R22229 DVSS.n22714 DVSS.n22710 4.5005
R22230 DVSS.n22714 DVSS.n673 4.5005
R22231 DVSS.n22714 DVSS.n22713 4.5005
R22232 DVSS.n22714 DVSS.n648 4.5005
R22233 DVSS.n22715 DVSS.n22714 4.5005
R22234 DVSS.n622 DVSS.n602 4.5005
R22235 DVSS.n624 DVSS.n602 4.5005
R22236 DVSS.n621 DVSS.n602 4.5005
R22237 DVSS.n627 DVSS.n602 4.5005
R22238 DVSS.n619 DVSS.n602 4.5005
R22239 DVSS.n628 DVSS.n602 4.5005
R22240 DVSS.n618 DVSS.n602 4.5005
R22241 DVSS.n629 DVSS.n602 4.5005
R22242 DVSS.n617 DVSS.n602 4.5005
R22243 DVSS.n22755 DVSS.n602 4.5005
R22244 DVSS.n22757 DVSS.n602 4.5005
R22245 DVSS.n622 DVSS.n601 4.5005
R22246 DVSS.n624 DVSS.n601 4.5005
R22247 DVSS.n621 DVSS.n601 4.5005
R22248 DVSS.n626 DVSS.n601 4.5005
R22249 DVSS.n620 DVSS.n601 4.5005
R22250 DVSS.n627 DVSS.n601 4.5005
R22251 DVSS.n619 DVSS.n601 4.5005
R22252 DVSS.n628 DVSS.n601 4.5005
R22253 DVSS.n618 DVSS.n601 4.5005
R22254 DVSS.n629 DVSS.n601 4.5005
R22255 DVSS.n617 DVSS.n601 4.5005
R22256 DVSS.n631 DVSS.n601 4.5005
R22257 DVSS.n22755 DVSS.n601 4.5005
R22258 DVSS.n22757 DVSS.n601 4.5005
R22259 DVSS.n622 DVSS.n603 4.5005
R22260 DVSS.n624 DVSS.n603 4.5005
R22261 DVSS.n621 DVSS.n603 4.5005
R22262 DVSS.n626 DVSS.n603 4.5005
R22263 DVSS.n620 DVSS.n603 4.5005
R22264 DVSS.n627 DVSS.n603 4.5005
R22265 DVSS.n619 DVSS.n603 4.5005
R22266 DVSS.n628 DVSS.n603 4.5005
R22267 DVSS.n618 DVSS.n603 4.5005
R22268 DVSS.n629 DVSS.n603 4.5005
R22269 DVSS.n617 DVSS.n603 4.5005
R22270 DVSS.n631 DVSS.n603 4.5005
R22271 DVSS.n22755 DVSS.n603 4.5005
R22272 DVSS.n22757 DVSS.n603 4.5005
R22273 DVSS.n622 DVSS.n600 4.5005
R22274 DVSS.n624 DVSS.n600 4.5005
R22275 DVSS.n621 DVSS.n600 4.5005
R22276 DVSS.n626 DVSS.n600 4.5005
R22277 DVSS.n620 DVSS.n600 4.5005
R22278 DVSS.n627 DVSS.n600 4.5005
R22279 DVSS.n619 DVSS.n600 4.5005
R22280 DVSS.n628 DVSS.n600 4.5005
R22281 DVSS.n618 DVSS.n600 4.5005
R22282 DVSS.n629 DVSS.n600 4.5005
R22283 DVSS.n617 DVSS.n600 4.5005
R22284 DVSS.n631 DVSS.n600 4.5005
R22285 DVSS.n616 DVSS.n600 4.5005
R22286 DVSS.n22755 DVSS.n600 4.5005
R22287 DVSS.n22757 DVSS.n600 4.5005
R22288 DVSS.n622 DVSS.n604 4.5005
R22289 DVSS.n624 DVSS.n604 4.5005
R22290 DVSS.n621 DVSS.n604 4.5005
R22291 DVSS.n626 DVSS.n604 4.5005
R22292 DVSS.n620 DVSS.n604 4.5005
R22293 DVSS.n627 DVSS.n604 4.5005
R22294 DVSS.n619 DVSS.n604 4.5005
R22295 DVSS.n628 DVSS.n604 4.5005
R22296 DVSS.n618 DVSS.n604 4.5005
R22297 DVSS.n629 DVSS.n604 4.5005
R22298 DVSS.n617 DVSS.n604 4.5005
R22299 DVSS.n631 DVSS.n604 4.5005
R22300 DVSS.n616 DVSS.n604 4.5005
R22301 DVSS.n22755 DVSS.n604 4.5005
R22302 DVSS.n22757 DVSS.n604 4.5005
R22303 DVSS.n622 DVSS.n599 4.5005
R22304 DVSS.n624 DVSS.n599 4.5005
R22305 DVSS.n621 DVSS.n599 4.5005
R22306 DVSS.n626 DVSS.n599 4.5005
R22307 DVSS.n620 DVSS.n599 4.5005
R22308 DVSS.n627 DVSS.n599 4.5005
R22309 DVSS.n619 DVSS.n599 4.5005
R22310 DVSS.n628 DVSS.n599 4.5005
R22311 DVSS.n618 DVSS.n599 4.5005
R22312 DVSS.n629 DVSS.n599 4.5005
R22313 DVSS.n617 DVSS.n599 4.5005
R22314 DVSS.n631 DVSS.n599 4.5005
R22315 DVSS.n22755 DVSS.n599 4.5005
R22316 DVSS.n22757 DVSS.n599 4.5005
R22317 DVSS.n622 DVSS.n605 4.5005
R22318 DVSS.n624 DVSS.n605 4.5005
R22319 DVSS.n621 DVSS.n605 4.5005
R22320 DVSS.n626 DVSS.n605 4.5005
R22321 DVSS.n620 DVSS.n605 4.5005
R22322 DVSS.n627 DVSS.n605 4.5005
R22323 DVSS.n619 DVSS.n605 4.5005
R22324 DVSS.n628 DVSS.n605 4.5005
R22325 DVSS.n618 DVSS.n605 4.5005
R22326 DVSS.n629 DVSS.n605 4.5005
R22327 DVSS.n617 DVSS.n605 4.5005
R22328 DVSS.n631 DVSS.n605 4.5005
R22329 DVSS.n22755 DVSS.n605 4.5005
R22330 DVSS.n612 DVSS.n605 4.5005
R22331 DVSS.n22757 DVSS.n605 4.5005
R22332 DVSS.n622 DVSS.n598 4.5005
R22333 DVSS.n624 DVSS.n598 4.5005
R22334 DVSS.n621 DVSS.n598 4.5005
R22335 DVSS.n626 DVSS.n598 4.5005
R22336 DVSS.n620 DVSS.n598 4.5005
R22337 DVSS.n627 DVSS.n598 4.5005
R22338 DVSS.n619 DVSS.n598 4.5005
R22339 DVSS.n628 DVSS.n598 4.5005
R22340 DVSS.n618 DVSS.n598 4.5005
R22341 DVSS.n629 DVSS.n598 4.5005
R22342 DVSS.n617 DVSS.n598 4.5005
R22343 DVSS.n631 DVSS.n598 4.5005
R22344 DVSS.n22755 DVSS.n598 4.5005
R22345 DVSS.n22757 DVSS.n598 4.5005
R22346 DVSS.n622 DVSS.n606 4.5005
R22347 DVSS.n624 DVSS.n606 4.5005
R22348 DVSS.n621 DVSS.n606 4.5005
R22349 DVSS.n626 DVSS.n606 4.5005
R22350 DVSS.n620 DVSS.n606 4.5005
R22351 DVSS.n627 DVSS.n606 4.5005
R22352 DVSS.n619 DVSS.n606 4.5005
R22353 DVSS.n628 DVSS.n606 4.5005
R22354 DVSS.n618 DVSS.n606 4.5005
R22355 DVSS.n629 DVSS.n606 4.5005
R22356 DVSS.n617 DVSS.n606 4.5005
R22357 DVSS.n631 DVSS.n606 4.5005
R22358 DVSS.n616 DVSS.n606 4.5005
R22359 DVSS.n22755 DVSS.n606 4.5005
R22360 DVSS.n22757 DVSS.n606 4.5005
R22361 DVSS.n622 DVSS.n597 4.5005
R22362 DVSS.n624 DVSS.n597 4.5005
R22363 DVSS.n621 DVSS.n597 4.5005
R22364 DVSS.n626 DVSS.n597 4.5005
R22365 DVSS.n620 DVSS.n597 4.5005
R22366 DVSS.n627 DVSS.n597 4.5005
R22367 DVSS.n619 DVSS.n597 4.5005
R22368 DVSS.n628 DVSS.n597 4.5005
R22369 DVSS.n618 DVSS.n597 4.5005
R22370 DVSS.n629 DVSS.n597 4.5005
R22371 DVSS.n617 DVSS.n597 4.5005
R22372 DVSS.n631 DVSS.n597 4.5005
R22373 DVSS.n22755 DVSS.n597 4.5005
R22374 DVSS.n612 DVSS.n597 4.5005
R22375 DVSS.n22757 DVSS.n597 4.5005
R22376 DVSS.n22756 DVSS.n622 4.5005
R22377 DVSS.n22756 DVSS.n624 4.5005
R22378 DVSS.n22756 DVSS.n621 4.5005
R22379 DVSS.n22756 DVSS.n626 4.5005
R22380 DVSS.n22756 DVSS.n620 4.5005
R22381 DVSS.n22756 DVSS.n627 4.5005
R22382 DVSS.n22756 DVSS.n619 4.5005
R22383 DVSS.n22756 DVSS.n628 4.5005
R22384 DVSS.n22756 DVSS.n618 4.5005
R22385 DVSS.n22756 DVSS.n629 4.5005
R22386 DVSS.n22756 DVSS.n617 4.5005
R22387 DVSS.n22756 DVSS.n631 4.5005
R22388 DVSS.n22756 DVSS.n616 4.5005
R22389 DVSS.n22756 DVSS.n22755 4.5005
R22390 DVSS.n22756 DVSS.n612 4.5005
R22391 DVSS.n22757 DVSS.n22756 4.5005
R22392 DVSS.n572 DVSS.n554 4.5005
R22393 DVSS.n574 DVSS.n554 4.5005
R22394 DVSS.n571 DVSS.n554 4.5005
R22395 DVSS.n577 DVSS.n554 4.5005
R22396 DVSS.n569 DVSS.n554 4.5005
R22397 DVSS.n578 DVSS.n554 4.5005
R22398 DVSS.n568 DVSS.n554 4.5005
R22399 DVSS.n579 DVSS.n554 4.5005
R22400 DVSS.n567 DVSS.n554 4.5005
R22401 DVSS.n22796 DVSS.n554 4.5005
R22402 DVSS.n22798 DVSS.n554 4.5005
R22403 DVSS.n572 DVSS.n552 4.5005
R22404 DVSS.n574 DVSS.n552 4.5005
R22405 DVSS.n571 DVSS.n552 4.5005
R22406 DVSS.n576 DVSS.n552 4.5005
R22407 DVSS.n570 DVSS.n552 4.5005
R22408 DVSS.n577 DVSS.n552 4.5005
R22409 DVSS.n569 DVSS.n552 4.5005
R22410 DVSS.n578 DVSS.n552 4.5005
R22411 DVSS.n568 DVSS.n552 4.5005
R22412 DVSS.n579 DVSS.n552 4.5005
R22413 DVSS.n567 DVSS.n552 4.5005
R22414 DVSS.n581 DVSS.n552 4.5005
R22415 DVSS.n22796 DVSS.n552 4.5005
R22416 DVSS.n22798 DVSS.n552 4.5005
R22417 DVSS.n572 DVSS.n556 4.5005
R22418 DVSS.n574 DVSS.n556 4.5005
R22419 DVSS.n571 DVSS.n556 4.5005
R22420 DVSS.n576 DVSS.n556 4.5005
R22421 DVSS.n570 DVSS.n556 4.5005
R22422 DVSS.n577 DVSS.n556 4.5005
R22423 DVSS.n569 DVSS.n556 4.5005
R22424 DVSS.n578 DVSS.n556 4.5005
R22425 DVSS.n568 DVSS.n556 4.5005
R22426 DVSS.n579 DVSS.n556 4.5005
R22427 DVSS.n567 DVSS.n556 4.5005
R22428 DVSS.n581 DVSS.n556 4.5005
R22429 DVSS.n22796 DVSS.n556 4.5005
R22430 DVSS.n22798 DVSS.n556 4.5005
R22431 DVSS.n572 DVSS.n551 4.5005
R22432 DVSS.n574 DVSS.n551 4.5005
R22433 DVSS.n571 DVSS.n551 4.5005
R22434 DVSS.n576 DVSS.n551 4.5005
R22435 DVSS.n570 DVSS.n551 4.5005
R22436 DVSS.n577 DVSS.n551 4.5005
R22437 DVSS.n569 DVSS.n551 4.5005
R22438 DVSS.n578 DVSS.n551 4.5005
R22439 DVSS.n568 DVSS.n551 4.5005
R22440 DVSS.n579 DVSS.n551 4.5005
R22441 DVSS.n567 DVSS.n551 4.5005
R22442 DVSS.n581 DVSS.n551 4.5005
R22443 DVSS.n566 DVSS.n551 4.5005
R22444 DVSS.n22796 DVSS.n551 4.5005
R22445 DVSS.n22798 DVSS.n551 4.5005
R22446 DVSS.n572 DVSS.n558 4.5005
R22447 DVSS.n574 DVSS.n558 4.5005
R22448 DVSS.n571 DVSS.n558 4.5005
R22449 DVSS.n576 DVSS.n558 4.5005
R22450 DVSS.n570 DVSS.n558 4.5005
R22451 DVSS.n577 DVSS.n558 4.5005
R22452 DVSS.n569 DVSS.n558 4.5005
R22453 DVSS.n578 DVSS.n558 4.5005
R22454 DVSS.n568 DVSS.n558 4.5005
R22455 DVSS.n579 DVSS.n558 4.5005
R22456 DVSS.n567 DVSS.n558 4.5005
R22457 DVSS.n581 DVSS.n558 4.5005
R22458 DVSS.n566 DVSS.n558 4.5005
R22459 DVSS.n22796 DVSS.n558 4.5005
R22460 DVSS.n22798 DVSS.n558 4.5005
R22461 DVSS.n572 DVSS.n550 4.5005
R22462 DVSS.n574 DVSS.n550 4.5005
R22463 DVSS.n571 DVSS.n550 4.5005
R22464 DVSS.n576 DVSS.n550 4.5005
R22465 DVSS.n570 DVSS.n550 4.5005
R22466 DVSS.n577 DVSS.n550 4.5005
R22467 DVSS.n569 DVSS.n550 4.5005
R22468 DVSS.n578 DVSS.n550 4.5005
R22469 DVSS.n568 DVSS.n550 4.5005
R22470 DVSS.n579 DVSS.n550 4.5005
R22471 DVSS.n567 DVSS.n550 4.5005
R22472 DVSS.n581 DVSS.n550 4.5005
R22473 DVSS.n22796 DVSS.n550 4.5005
R22474 DVSS.n22798 DVSS.n550 4.5005
R22475 DVSS.n572 DVSS.n559 4.5005
R22476 DVSS.n574 DVSS.n559 4.5005
R22477 DVSS.n571 DVSS.n559 4.5005
R22478 DVSS.n576 DVSS.n559 4.5005
R22479 DVSS.n570 DVSS.n559 4.5005
R22480 DVSS.n577 DVSS.n559 4.5005
R22481 DVSS.n569 DVSS.n559 4.5005
R22482 DVSS.n578 DVSS.n559 4.5005
R22483 DVSS.n568 DVSS.n559 4.5005
R22484 DVSS.n579 DVSS.n559 4.5005
R22485 DVSS.n567 DVSS.n559 4.5005
R22486 DVSS.n581 DVSS.n559 4.5005
R22487 DVSS.n22796 DVSS.n559 4.5005
R22488 DVSS.n559 DVSS.n547 4.5005
R22489 DVSS.n22798 DVSS.n559 4.5005
R22490 DVSS.n572 DVSS.n549 4.5005
R22491 DVSS.n574 DVSS.n549 4.5005
R22492 DVSS.n571 DVSS.n549 4.5005
R22493 DVSS.n576 DVSS.n549 4.5005
R22494 DVSS.n570 DVSS.n549 4.5005
R22495 DVSS.n577 DVSS.n549 4.5005
R22496 DVSS.n569 DVSS.n549 4.5005
R22497 DVSS.n578 DVSS.n549 4.5005
R22498 DVSS.n568 DVSS.n549 4.5005
R22499 DVSS.n579 DVSS.n549 4.5005
R22500 DVSS.n567 DVSS.n549 4.5005
R22501 DVSS.n581 DVSS.n549 4.5005
R22502 DVSS.n22796 DVSS.n549 4.5005
R22503 DVSS.n22798 DVSS.n549 4.5005
R22504 DVSS.n572 DVSS.n561 4.5005
R22505 DVSS.n574 DVSS.n561 4.5005
R22506 DVSS.n571 DVSS.n561 4.5005
R22507 DVSS.n576 DVSS.n561 4.5005
R22508 DVSS.n570 DVSS.n561 4.5005
R22509 DVSS.n577 DVSS.n561 4.5005
R22510 DVSS.n569 DVSS.n561 4.5005
R22511 DVSS.n578 DVSS.n561 4.5005
R22512 DVSS.n568 DVSS.n561 4.5005
R22513 DVSS.n579 DVSS.n561 4.5005
R22514 DVSS.n567 DVSS.n561 4.5005
R22515 DVSS.n581 DVSS.n561 4.5005
R22516 DVSS.n566 DVSS.n561 4.5005
R22517 DVSS.n22796 DVSS.n561 4.5005
R22518 DVSS.n22798 DVSS.n561 4.5005
R22519 DVSS.n572 DVSS.n548 4.5005
R22520 DVSS.n574 DVSS.n548 4.5005
R22521 DVSS.n571 DVSS.n548 4.5005
R22522 DVSS.n576 DVSS.n548 4.5005
R22523 DVSS.n570 DVSS.n548 4.5005
R22524 DVSS.n577 DVSS.n548 4.5005
R22525 DVSS.n569 DVSS.n548 4.5005
R22526 DVSS.n578 DVSS.n548 4.5005
R22527 DVSS.n568 DVSS.n548 4.5005
R22528 DVSS.n579 DVSS.n548 4.5005
R22529 DVSS.n567 DVSS.n548 4.5005
R22530 DVSS.n581 DVSS.n548 4.5005
R22531 DVSS.n22796 DVSS.n548 4.5005
R22532 DVSS.n548 DVSS.n547 4.5005
R22533 DVSS.n22798 DVSS.n548 4.5005
R22534 DVSS.n22797 DVSS.n572 4.5005
R22535 DVSS.n22797 DVSS.n574 4.5005
R22536 DVSS.n22797 DVSS.n571 4.5005
R22537 DVSS.n22797 DVSS.n576 4.5005
R22538 DVSS.n22797 DVSS.n570 4.5005
R22539 DVSS.n22797 DVSS.n577 4.5005
R22540 DVSS.n22797 DVSS.n569 4.5005
R22541 DVSS.n22797 DVSS.n578 4.5005
R22542 DVSS.n22797 DVSS.n568 4.5005
R22543 DVSS.n22797 DVSS.n579 4.5005
R22544 DVSS.n22797 DVSS.n567 4.5005
R22545 DVSS.n22797 DVSS.n581 4.5005
R22546 DVSS.n22797 DVSS.n566 4.5005
R22547 DVSS.n22797 DVSS.n22796 4.5005
R22548 DVSS.n22797 DVSS.n547 4.5005
R22549 DVSS.n22798 DVSS.n22797 4.5005
R22550 DVSS.n522 DVSS.n502 4.5005
R22551 DVSS.n526 DVSS.n502 4.5005
R22552 DVSS.n520 DVSS.n502 4.5005
R22553 DVSS.n527 DVSS.n502 4.5005
R22554 DVSS.n519 DVSS.n502 4.5005
R22555 DVSS.n528 DVSS.n502 4.5005
R22556 DVSS.n518 DVSS.n502 4.5005
R22557 DVSS.n531 DVSS.n502 4.5005
R22558 DVSS.n516 DVSS.n502 4.5005
R22559 DVSS.n22837 DVSS.n502 4.5005
R22560 DVSS.n22839 DVSS.n502 4.5005
R22561 DVSS.n522 DVSS.n501 4.5005
R22562 DVSS.n525 DVSS.n501 4.5005
R22563 DVSS.n521 DVSS.n501 4.5005
R22564 DVSS.n526 DVSS.n501 4.5005
R22565 DVSS.n520 DVSS.n501 4.5005
R22566 DVSS.n527 DVSS.n501 4.5005
R22567 DVSS.n519 DVSS.n501 4.5005
R22568 DVSS.n528 DVSS.n501 4.5005
R22569 DVSS.n518 DVSS.n501 4.5005
R22570 DVSS.n530 DVSS.n501 4.5005
R22571 DVSS.n517 DVSS.n501 4.5005
R22572 DVSS.n531 DVSS.n501 4.5005
R22573 DVSS.n22837 DVSS.n501 4.5005
R22574 DVSS.n22839 DVSS.n501 4.5005
R22575 DVSS.n522 DVSS.n503 4.5005
R22576 DVSS.n525 DVSS.n503 4.5005
R22577 DVSS.n521 DVSS.n503 4.5005
R22578 DVSS.n526 DVSS.n503 4.5005
R22579 DVSS.n520 DVSS.n503 4.5005
R22580 DVSS.n527 DVSS.n503 4.5005
R22581 DVSS.n519 DVSS.n503 4.5005
R22582 DVSS.n528 DVSS.n503 4.5005
R22583 DVSS.n518 DVSS.n503 4.5005
R22584 DVSS.n530 DVSS.n503 4.5005
R22585 DVSS.n517 DVSS.n503 4.5005
R22586 DVSS.n531 DVSS.n503 4.5005
R22587 DVSS.n22837 DVSS.n503 4.5005
R22588 DVSS.n22839 DVSS.n503 4.5005
R22589 DVSS.n522 DVSS.n500 4.5005
R22590 DVSS.n525 DVSS.n500 4.5005
R22591 DVSS.n521 DVSS.n500 4.5005
R22592 DVSS.n526 DVSS.n500 4.5005
R22593 DVSS.n520 DVSS.n500 4.5005
R22594 DVSS.n527 DVSS.n500 4.5005
R22595 DVSS.n519 DVSS.n500 4.5005
R22596 DVSS.n528 DVSS.n500 4.5005
R22597 DVSS.n518 DVSS.n500 4.5005
R22598 DVSS.n530 DVSS.n500 4.5005
R22599 DVSS.n517 DVSS.n500 4.5005
R22600 DVSS.n531 DVSS.n500 4.5005
R22601 DVSS.n516 DVSS.n500 4.5005
R22602 DVSS.n22837 DVSS.n500 4.5005
R22603 DVSS.n22839 DVSS.n500 4.5005
R22604 DVSS.n522 DVSS.n504 4.5005
R22605 DVSS.n525 DVSS.n504 4.5005
R22606 DVSS.n521 DVSS.n504 4.5005
R22607 DVSS.n526 DVSS.n504 4.5005
R22608 DVSS.n520 DVSS.n504 4.5005
R22609 DVSS.n527 DVSS.n504 4.5005
R22610 DVSS.n519 DVSS.n504 4.5005
R22611 DVSS.n528 DVSS.n504 4.5005
R22612 DVSS.n518 DVSS.n504 4.5005
R22613 DVSS.n530 DVSS.n504 4.5005
R22614 DVSS.n517 DVSS.n504 4.5005
R22615 DVSS.n531 DVSS.n504 4.5005
R22616 DVSS.n516 DVSS.n504 4.5005
R22617 DVSS.n22837 DVSS.n504 4.5005
R22618 DVSS.n22839 DVSS.n504 4.5005
R22619 DVSS.n522 DVSS.n499 4.5005
R22620 DVSS.n525 DVSS.n499 4.5005
R22621 DVSS.n521 DVSS.n499 4.5005
R22622 DVSS.n526 DVSS.n499 4.5005
R22623 DVSS.n520 DVSS.n499 4.5005
R22624 DVSS.n527 DVSS.n499 4.5005
R22625 DVSS.n519 DVSS.n499 4.5005
R22626 DVSS.n528 DVSS.n499 4.5005
R22627 DVSS.n518 DVSS.n499 4.5005
R22628 DVSS.n530 DVSS.n499 4.5005
R22629 DVSS.n517 DVSS.n499 4.5005
R22630 DVSS.n531 DVSS.n499 4.5005
R22631 DVSS.n22837 DVSS.n499 4.5005
R22632 DVSS.n22839 DVSS.n499 4.5005
R22633 DVSS.n522 DVSS.n505 4.5005
R22634 DVSS.n525 DVSS.n505 4.5005
R22635 DVSS.n521 DVSS.n505 4.5005
R22636 DVSS.n526 DVSS.n505 4.5005
R22637 DVSS.n520 DVSS.n505 4.5005
R22638 DVSS.n527 DVSS.n505 4.5005
R22639 DVSS.n519 DVSS.n505 4.5005
R22640 DVSS.n528 DVSS.n505 4.5005
R22641 DVSS.n518 DVSS.n505 4.5005
R22642 DVSS.n530 DVSS.n505 4.5005
R22643 DVSS.n517 DVSS.n505 4.5005
R22644 DVSS.n531 DVSS.n505 4.5005
R22645 DVSS.n22837 DVSS.n505 4.5005
R22646 DVSS.n512 DVSS.n505 4.5005
R22647 DVSS.n22839 DVSS.n505 4.5005
R22648 DVSS.n522 DVSS.n498 4.5005
R22649 DVSS.n525 DVSS.n498 4.5005
R22650 DVSS.n521 DVSS.n498 4.5005
R22651 DVSS.n526 DVSS.n498 4.5005
R22652 DVSS.n520 DVSS.n498 4.5005
R22653 DVSS.n527 DVSS.n498 4.5005
R22654 DVSS.n519 DVSS.n498 4.5005
R22655 DVSS.n528 DVSS.n498 4.5005
R22656 DVSS.n518 DVSS.n498 4.5005
R22657 DVSS.n530 DVSS.n498 4.5005
R22658 DVSS.n517 DVSS.n498 4.5005
R22659 DVSS.n531 DVSS.n498 4.5005
R22660 DVSS.n22837 DVSS.n498 4.5005
R22661 DVSS.n22839 DVSS.n498 4.5005
R22662 DVSS.n522 DVSS.n506 4.5005
R22663 DVSS.n525 DVSS.n506 4.5005
R22664 DVSS.n521 DVSS.n506 4.5005
R22665 DVSS.n526 DVSS.n506 4.5005
R22666 DVSS.n520 DVSS.n506 4.5005
R22667 DVSS.n527 DVSS.n506 4.5005
R22668 DVSS.n519 DVSS.n506 4.5005
R22669 DVSS.n528 DVSS.n506 4.5005
R22670 DVSS.n518 DVSS.n506 4.5005
R22671 DVSS.n530 DVSS.n506 4.5005
R22672 DVSS.n517 DVSS.n506 4.5005
R22673 DVSS.n531 DVSS.n506 4.5005
R22674 DVSS.n516 DVSS.n506 4.5005
R22675 DVSS.n22837 DVSS.n506 4.5005
R22676 DVSS.n22839 DVSS.n506 4.5005
R22677 DVSS.n522 DVSS.n497 4.5005
R22678 DVSS.n525 DVSS.n497 4.5005
R22679 DVSS.n521 DVSS.n497 4.5005
R22680 DVSS.n526 DVSS.n497 4.5005
R22681 DVSS.n520 DVSS.n497 4.5005
R22682 DVSS.n527 DVSS.n497 4.5005
R22683 DVSS.n519 DVSS.n497 4.5005
R22684 DVSS.n528 DVSS.n497 4.5005
R22685 DVSS.n518 DVSS.n497 4.5005
R22686 DVSS.n530 DVSS.n497 4.5005
R22687 DVSS.n517 DVSS.n497 4.5005
R22688 DVSS.n531 DVSS.n497 4.5005
R22689 DVSS.n22837 DVSS.n497 4.5005
R22690 DVSS.n512 DVSS.n497 4.5005
R22691 DVSS.n22839 DVSS.n497 4.5005
R22692 DVSS.n22838 DVSS.n522 4.5005
R22693 DVSS.n22838 DVSS.n525 4.5005
R22694 DVSS.n22838 DVSS.n521 4.5005
R22695 DVSS.n22838 DVSS.n526 4.5005
R22696 DVSS.n22838 DVSS.n520 4.5005
R22697 DVSS.n22838 DVSS.n527 4.5005
R22698 DVSS.n22838 DVSS.n519 4.5005
R22699 DVSS.n22838 DVSS.n528 4.5005
R22700 DVSS.n22838 DVSS.n518 4.5005
R22701 DVSS.n22838 DVSS.n530 4.5005
R22702 DVSS.n22838 DVSS.n517 4.5005
R22703 DVSS.n22838 DVSS.n531 4.5005
R22704 DVSS.n22838 DVSS.n516 4.5005
R22705 DVSS.n22838 DVSS.n22837 4.5005
R22706 DVSS.n22838 DVSS.n512 4.5005
R22707 DVSS.n22839 DVSS.n22838 4.5005
R22708 DVSS.n21461 DVSS.n21460 4.5005
R22709 DVSS.n21459 DVSS.n21452 4.5005
R22710 DVSS.n21457 DVSS.n21456 4.5005
R22711 DVSS.n21455 DVSS.n21454 4.5005
R22712 DVSS.n21453 DVSS.n757 4.5005
R22713 DVSS.n22572 DVSS.n756 4.5005
R22714 DVSS.n22574 DVSS.n22573 4.5005
R22715 DVSS.n22575 DVSS.n755 4.5005
R22716 DVSS.n22577 DVSS.n22576 4.5005
R22717 DVSS.n22578 DVSS.n754 4.5005
R22718 DVSS.n22580 DVSS.n22579 4.5005
R22719 DVSS.n22582 DVSS.n753 4.5005
R22720 DVSS.n22584 DVSS.n22583 4.5005
R22721 DVSS.n22588 DVSS.n22587 4.5005
R22722 DVSS.n22589 DVSS.n750 4.5005
R22723 DVSS.n22592 DVSS.n22591 4.5005
R22724 DVSS.n22593 DVSS.n749 4.5005
R22725 DVSS.n22595 DVSS.n22594 4.5005
R22726 DVSS.n22596 DVSS.n748 4.5005
R22727 DVSS.n22598 DVSS.n22597 4.5005
R22728 DVSS.n22599 DVSS.n747 4.5005
R22729 DVSS.n22601 DVSS.n22600 4.5005
R22730 DVSS.n22602 DVSS.n746 4.5005
R22731 DVSS.n22604 DVSS.n22603 4.5005
R22732 DVSS.n22606 DVSS.n22605 4.5005
R22733 DVSS.n22608 DVSS.n22607 4.5005
R22734 DVSS.n22610 DVSS.n22609 4.5005
R22735 DVSS.n22611 DVSS.n742 4.5005
R22736 DVSS.n22613 DVSS.n22612 4.5005
R22737 DVSS.n22614 DVSS.n741 4.5005
R22738 DVSS.n22616 DVSS.n22615 4.5005
R22739 DVSS.n22617 DVSS.n740 4.5005
R22740 DVSS.n22619 DVSS.n22618 4.5005
R22741 DVSS.n22620 DVSS.n739 4.5005
R22742 DVSS.n22622 DVSS.n22621 4.5005
R22743 DVSS.n22624 DVSS.n738 4.5005
R22744 DVSS.n22626 DVSS.n22625 4.5005
R22745 DVSS.n22630 DVSS.n736 4.5005
R22746 DVSS.n22632 DVSS.n22631 4.5005
R22747 DVSS.n22634 DVSS.n22633 4.5005
R22748 DVSS.n22635 DVSS.n733 4.5005
R22749 DVSS.n21177 DVSS.n13660 4.5005
R22750 DVSS.n21179 DVSS.n21178 4.5005
R22751 DVSS.n13661 DVSS.n13659 4.5005
R22752 DVSS.n13667 DVSS.n13666 4.5005
R22753 DVSS.n21160 DVSS.n21159 4.5005
R22754 DVSS.n21158 DVSS.n13683 4.5005
R22755 DVSS.n18507 DVSS.n18506 4.5005
R22756 DVSS.n18508 DVSS.n18505 4.5005
R22757 DVSS.n18519 DVSS.n18518 4.5005
R22758 DVSS.n18520 DVSS.n15148 4.5005
R22759 DVSS.n18522 DVSS.n18521 4.5005
R22760 DVSS.n18523 DVSS.n15147 4.5005
R22761 DVSS.n18525 DVSS.n18524 4.5005
R22762 DVSS.n17787 DVSS.n15921 4.5005
R22763 DVSS.n17789 DVSS.n17788 4.5005
R22764 DVSS.n18170 DVSS.n18169 4.5005
R22765 DVSS.n18171 DVSS.n15532 4.5005
R22766 DVSS.n19918 DVSS.n19917 4.5005
R22767 DVSS.n19919 DVSS.n15139 4.5005
R22768 DVSS.n19921 DVSS.n19920 4.5005
R22769 DVSS.n19922 DVSS.n15138 4.5005
R22770 DVSS.n19924 DVSS.n19923 4.5005
R22771 DVSS.n15135 DVSS.n15134 4.5005
R22772 DVSS.n15133 DVSS.n15127 4.5005
R22773 DVSS.n15131 DVSS.n15130 4.5005
R22774 DVSS.n15129 DVSS.n15128 4.5005
R22775 DVSS.n14315 DVSS.n14314 4.5005
R22776 DVSS.n14313 DVSS.n14312 4.5005
R22777 DVSS.n20990 DVSS.n20989 4.5005
R22778 DVSS.n20991 DVSS.n14311 4.5005
R22779 DVSS.n20993 DVSS.n20992 4.5005
R22780 DVSS.n20994 DVSS.n14309 4.5005
R22781 DVSS.n21024 DVSS.n21023 4.5005
R22782 DVSS.n21022 DVSS.n14310 4.5005
R22783 DVSS.n21021 DVSS.n21020 4.5005
R22784 DVSS.n21019 DVSS.n20995 4.5005
R22785 DVSS.n21018 DVSS.n21017 4.5005
R22786 DVSS.n21016 DVSS.n20996 4.5005
R22787 DVSS.n21011 DVSS.n20997 4.5005
R22788 DVSS.n21012 DVSS.n20998 4.5005
R22789 DVSS.n21008 DVSS.n21007 4.5005
R22790 DVSS.n21006 DVSS.n21000 4.5005
R22791 DVSS.n21004 DVSS.n21003 4.5005
R22792 DVSS.n21002 DVSS.n21001 4.5005
R22793 DVSS.n13372 DVSS.n13371 4.5005
R22794 DVSS.n22886 DVSS.n452 4.5005
R22795 DVSS.n22888 DVSS.n22887 4.5005
R22796 DVSS.n22890 DVSS.n451 4.5005
R22797 DVSS.n22892 DVSS.n22891 4.5005
R22798 DVSS.n22896 DVSS.n22895 4.5005
R22799 DVSS.n22897 DVSS.n448 4.5005
R22800 DVSS.n22900 DVSS.n22899 4.5005
R22801 DVSS.n22901 DVSS.n447 4.5005
R22802 DVSS.n22903 DVSS.n22902 4.5005
R22803 DVSS.n22904 DVSS.n446 4.5005
R22804 DVSS.n22906 DVSS.n22905 4.5005
R22805 DVSS.n22907 DVSS.n445 4.5005
R22806 DVSS.n22909 DVSS.n22908 4.5005
R22807 DVSS.n22910 DVSS.n444 4.5005
R22808 DVSS.n22912 DVSS.n22911 4.5005
R22809 DVSS.n22914 DVSS.n22913 4.5005
R22810 DVSS.n22916 DVSS.n22915 4.5005
R22811 DVSS.n22918 DVSS.n22917 4.5005
R22812 DVSS.n22919 DVSS.n440 4.5005
R22813 DVSS.n22921 DVSS.n22920 4.5005
R22814 DVSS.n22922 DVSS.n439 4.5005
R22815 DVSS.n22924 DVSS.n22923 4.5005
R22816 DVSS.n22925 DVSS.n438 4.5005
R22817 DVSS.n22927 DVSS.n22926 4.5005
R22818 DVSS.n22928 DVSS.n437 4.5005
R22819 DVSS.n22930 DVSS.n22929 4.5005
R22820 DVSS.n22932 DVSS.n436 4.5005
R22821 DVSS.n22934 DVSS.n22933 4.5005
R22822 DVSS.n22938 DVSS.n22937 4.5005
R22823 DVSS.n22939 DVSS.n433 4.5005
R22824 DVSS.n22942 DVSS.n22941 4.5005
R22825 DVSS.n22943 DVSS.n432 4.5005
R22826 DVSS.n22945 DVSS.n22944 4.5005
R22827 DVSS.n22946 DVSS.n431 4.5005
R22828 DVSS.n22948 DVSS.n22947 4.5005
R22829 DVSS.n22949 DVSS.n430 4.5005
R22830 DVSS.n22952 DVSS.n22951 4.5005
R22831 DVSS.n22953 DVSS.n429 4.5005
R22832 DVSS.n22955 DVSS.n22954 4.5005
R22833 DVSS.n22957 DVSS.n22956 4.5005
R22834 DVSS.n22958 DVSS.n427 4.5005
R22835 DVSS.n426 DVSS.n425 4.5005
R22836 DVSS.n22965 DVSS.n22964 4.5005
R22837 DVSS.n22966 DVSS.n424 4.5005
R22838 DVSS.n22968 DVSS.n22967 4.5005
R22839 DVSS.n22969 DVSS.n422 4.5005
R22840 DVSS.n21471 DVSS.n1500 4.5005
R22841 DVSS.n21470 DVSS.n21469 4.5005
R22842 DVSS.n21468 DVSS.n21448 4.5005
R22843 DVSS.n21467 DVSS.n21466 4.5005
R22844 DVSS.n21450 DVSS.n21449 4.5005
R22845 DVSS.n12808 DVSS.n12785 4.5005
R22846 DVSS.n12808 DVSS.n12782 4.5005
R22847 DVSS.n12808 DVSS.n12787 4.5005
R22848 DVSS.n12808 DVSS.n12781 4.5005
R22849 DVSS.n12808 DVSS.n12789 4.5005
R22850 DVSS.n12808 DVSS.n12780 4.5005
R22851 DVSS.n12808 DVSS.n12790 4.5005
R22852 DVSS.n12808 DVSS.n12778 4.5005
R22853 DVSS.n12808 DVSS.n12793 4.5005
R22854 DVSS.n12808 DVSS.n12777 4.5005
R22855 DVSS.n13099 DVSS.n12808 4.5005
R22856 DVSS.n12809 DVSS.n12785 4.5005
R22857 DVSS.n12809 DVSS.n12783 4.5005
R22858 DVSS.n12809 DVSS.n12786 4.5005
R22859 DVSS.n12809 DVSS.n12782 4.5005
R22860 DVSS.n12809 DVSS.n12787 4.5005
R22861 DVSS.n12809 DVSS.n12781 4.5005
R22862 DVSS.n12809 DVSS.n12789 4.5005
R22863 DVSS.n12809 DVSS.n12780 4.5005
R22864 DVSS.n12809 DVSS.n12790 4.5005
R22865 DVSS.n12809 DVSS.n12779 4.5005
R22866 DVSS.n12809 DVSS.n12792 4.5005
R22867 DVSS.n12809 DVSS.n12778 4.5005
R22868 DVSS.n12809 DVSS.n12793 4.5005
R22869 DVSS.n12809 DVSS.n12777 4.5005
R22870 DVSS.n13099 DVSS.n12809 4.5005
R22871 DVSS.n12805 DVSS.n12785 4.5005
R22872 DVSS.n12805 DVSS.n12783 4.5005
R22873 DVSS.n12805 DVSS.n12786 4.5005
R22874 DVSS.n12805 DVSS.n12782 4.5005
R22875 DVSS.n12805 DVSS.n12787 4.5005
R22876 DVSS.n12805 DVSS.n12781 4.5005
R22877 DVSS.n12805 DVSS.n12789 4.5005
R22878 DVSS.n12805 DVSS.n12780 4.5005
R22879 DVSS.n12805 DVSS.n12790 4.5005
R22880 DVSS.n12805 DVSS.n12779 4.5005
R22881 DVSS.n12805 DVSS.n12792 4.5005
R22882 DVSS.n12805 DVSS.n12778 4.5005
R22883 DVSS.n12805 DVSS.n12793 4.5005
R22884 DVSS.n12805 DVSS.n12777 4.5005
R22885 DVSS.n13099 DVSS.n12805 4.5005
R22886 DVSS.n12810 DVSS.n12785 4.5005
R22887 DVSS.n12810 DVSS.n12783 4.5005
R22888 DVSS.n12810 DVSS.n12786 4.5005
R22889 DVSS.n12810 DVSS.n12782 4.5005
R22890 DVSS.n12810 DVSS.n12787 4.5005
R22891 DVSS.n12810 DVSS.n12781 4.5005
R22892 DVSS.n12810 DVSS.n12789 4.5005
R22893 DVSS.n12810 DVSS.n12780 4.5005
R22894 DVSS.n12810 DVSS.n12790 4.5005
R22895 DVSS.n12810 DVSS.n12779 4.5005
R22896 DVSS.n12810 DVSS.n12792 4.5005
R22897 DVSS.n12810 DVSS.n12778 4.5005
R22898 DVSS.n12810 DVSS.n12793 4.5005
R22899 DVSS.n12810 DVSS.n12777 4.5005
R22900 DVSS.n13099 DVSS.n12810 4.5005
R22901 DVSS.n12804 DVSS.n12777 4.5005
R22902 DVSS.n13099 DVSS.n12804 4.5005
R22903 DVSS.n12804 DVSS.n12793 4.5005
R22904 DVSS.n12804 DVSS.n12778 4.5005
R22905 DVSS.n12804 DVSS.n12792 4.5005
R22906 DVSS.n12804 DVSS.n12779 4.5005
R22907 DVSS.n12804 DVSS.n12790 4.5005
R22908 DVSS.n12804 DVSS.n12780 4.5005
R22909 DVSS.n12804 DVSS.n12789 4.5005
R22910 DVSS.n12804 DVSS.n12781 4.5005
R22911 DVSS.n12804 DVSS.n12787 4.5005
R22912 DVSS.n12804 DVSS.n12782 4.5005
R22913 DVSS.n12804 DVSS.n12786 4.5005
R22914 DVSS.n12804 DVSS.n12783 4.5005
R22915 DVSS.n12804 DVSS.n12785 4.5005
R22916 DVSS.n12811 DVSS.n12777 4.5005
R22917 DVSS.n13099 DVSS.n12811 4.5005
R22918 DVSS.n12811 DVSS.n12793 4.5005
R22919 DVSS.n12811 DVSS.n12778 4.5005
R22920 DVSS.n12811 DVSS.n12792 4.5005
R22921 DVSS.n12811 DVSS.n12779 4.5005
R22922 DVSS.n12811 DVSS.n12790 4.5005
R22923 DVSS.n12811 DVSS.n12780 4.5005
R22924 DVSS.n12811 DVSS.n12789 4.5005
R22925 DVSS.n12811 DVSS.n12781 4.5005
R22926 DVSS.n12811 DVSS.n12787 4.5005
R22927 DVSS.n12811 DVSS.n12782 4.5005
R22928 DVSS.n12811 DVSS.n12786 4.5005
R22929 DVSS.n12811 DVSS.n12783 4.5005
R22930 DVSS.n12811 DVSS.n12785 4.5005
R22931 DVSS.n12803 DVSS.n12777 4.5005
R22932 DVSS.n13099 DVSS.n12803 4.5005
R22933 DVSS.n12803 DVSS.n12793 4.5005
R22934 DVSS.n12803 DVSS.n12778 4.5005
R22935 DVSS.n12803 DVSS.n12792 4.5005
R22936 DVSS.n12803 DVSS.n12779 4.5005
R22937 DVSS.n12803 DVSS.n12790 4.5005
R22938 DVSS.n12803 DVSS.n12780 4.5005
R22939 DVSS.n12803 DVSS.n12789 4.5005
R22940 DVSS.n12803 DVSS.n12781 4.5005
R22941 DVSS.n12803 DVSS.n12787 4.5005
R22942 DVSS.n12803 DVSS.n12782 4.5005
R22943 DVSS.n12803 DVSS.n12786 4.5005
R22944 DVSS.n12803 DVSS.n12783 4.5005
R22945 DVSS.n12803 DVSS.n12785 4.5005
R22946 DVSS.n12812 DVSS.n12785 4.5005
R22947 DVSS.n12812 DVSS.n12783 4.5005
R22948 DVSS.n12812 DVSS.n12786 4.5005
R22949 DVSS.n12812 DVSS.n12782 4.5005
R22950 DVSS.n12812 DVSS.n12787 4.5005
R22951 DVSS.n12812 DVSS.n12781 4.5005
R22952 DVSS.n12812 DVSS.n12789 4.5005
R22953 DVSS.n12812 DVSS.n12780 4.5005
R22954 DVSS.n12812 DVSS.n12790 4.5005
R22955 DVSS.n12812 DVSS.n12779 4.5005
R22956 DVSS.n12812 DVSS.n12792 4.5005
R22957 DVSS.n12812 DVSS.n12778 4.5005
R22958 DVSS.n12812 DVSS.n12793 4.5005
R22959 DVSS.n12812 DVSS.n12777 4.5005
R22960 DVSS.n13099 DVSS.n12812 4.5005
R22961 DVSS.n12802 DVSS.n12785 4.5005
R22962 DVSS.n12802 DVSS.n12783 4.5005
R22963 DVSS.n12802 DVSS.n12786 4.5005
R22964 DVSS.n12802 DVSS.n12782 4.5005
R22965 DVSS.n12802 DVSS.n12787 4.5005
R22966 DVSS.n12802 DVSS.n12781 4.5005
R22967 DVSS.n12802 DVSS.n12789 4.5005
R22968 DVSS.n12802 DVSS.n12780 4.5005
R22969 DVSS.n12802 DVSS.n12790 4.5005
R22970 DVSS.n12802 DVSS.n12779 4.5005
R22971 DVSS.n12802 DVSS.n12792 4.5005
R22972 DVSS.n12802 DVSS.n12778 4.5005
R22973 DVSS.n12802 DVSS.n12793 4.5005
R22974 DVSS.n12802 DVSS.n12777 4.5005
R22975 DVSS.n13099 DVSS.n12802 4.5005
R22976 DVSS.n12813 DVSS.n12785 4.5005
R22977 DVSS.n12813 DVSS.n12783 4.5005
R22978 DVSS.n12813 DVSS.n12786 4.5005
R22979 DVSS.n12813 DVSS.n12782 4.5005
R22980 DVSS.n12813 DVSS.n12787 4.5005
R22981 DVSS.n12813 DVSS.n12781 4.5005
R22982 DVSS.n12813 DVSS.n12789 4.5005
R22983 DVSS.n12813 DVSS.n12780 4.5005
R22984 DVSS.n12813 DVSS.n12790 4.5005
R22985 DVSS.n12813 DVSS.n12779 4.5005
R22986 DVSS.n12813 DVSS.n12792 4.5005
R22987 DVSS.n12813 DVSS.n12778 4.5005
R22988 DVSS.n12813 DVSS.n12793 4.5005
R22989 DVSS.n12813 DVSS.n12777 4.5005
R22990 DVSS.n13099 DVSS.n12813 4.5005
R22991 DVSS.n12801 DVSS.n12777 4.5005
R22992 DVSS.n13099 DVSS.n12801 4.5005
R22993 DVSS.n12801 DVSS.n12793 4.5005
R22994 DVSS.n12801 DVSS.n12778 4.5005
R22995 DVSS.n12801 DVSS.n12792 4.5005
R22996 DVSS.n12801 DVSS.n12779 4.5005
R22997 DVSS.n12801 DVSS.n12790 4.5005
R22998 DVSS.n12801 DVSS.n12780 4.5005
R22999 DVSS.n12801 DVSS.n12789 4.5005
R23000 DVSS.n12801 DVSS.n12781 4.5005
R23001 DVSS.n12801 DVSS.n12787 4.5005
R23002 DVSS.n12801 DVSS.n12782 4.5005
R23003 DVSS.n12801 DVSS.n12786 4.5005
R23004 DVSS.n12801 DVSS.n12783 4.5005
R23005 DVSS.n12801 DVSS.n12785 4.5005
R23006 DVSS.n12814 DVSS.n12777 4.5005
R23007 DVSS.n13099 DVSS.n12814 4.5005
R23008 DVSS.n12814 DVSS.n12793 4.5005
R23009 DVSS.n12814 DVSS.n12778 4.5005
R23010 DVSS.n12814 DVSS.n12792 4.5005
R23011 DVSS.n12814 DVSS.n12779 4.5005
R23012 DVSS.n12814 DVSS.n12790 4.5005
R23013 DVSS.n12814 DVSS.n12780 4.5005
R23014 DVSS.n12814 DVSS.n12789 4.5005
R23015 DVSS.n12814 DVSS.n12781 4.5005
R23016 DVSS.n12814 DVSS.n12787 4.5005
R23017 DVSS.n12814 DVSS.n12782 4.5005
R23018 DVSS.n12814 DVSS.n12786 4.5005
R23019 DVSS.n12814 DVSS.n12783 4.5005
R23020 DVSS.n12814 DVSS.n12785 4.5005
R23021 DVSS.n12800 DVSS.n12777 4.5005
R23022 DVSS.n13099 DVSS.n12800 4.5005
R23023 DVSS.n12800 DVSS.n12793 4.5005
R23024 DVSS.n12800 DVSS.n12778 4.5005
R23025 DVSS.n12800 DVSS.n12792 4.5005
R23026 DVSS.n12800 DVSS.n12779 4.5005
R23027 DVSS.n12800 DVSS.n12790 4.5005
R23028 DVSS.n12800 DVSS.n12780 4.5005
R23029 DVSS.n12800 DVSS.n12789 4.5005
R23030 DVSS.n12800 DVSS.n12781 4.5005
R23031 DVSS.n12800 DVSS.n12787 4.5005
R23032 DVSS.n12800 DVSS.n12782 4.5005
R23033 DVSS.n12800 DVSS.n12786 4.5005
R23034 DVSS.n12800 DVSS.n12783 4.5005
R23035 DVSS.n12800 DVSS.n12785 4.5005
R23036 DVSS.n12815 DVSS.n12777 4.5005
R23037 DVSS.n13099 DVSS.n12815 4.5005
R23038 DVSS.n12815 DVSS.n12793 4.5005
R23039 DVSS.n12815 DVSS.n12778 4.5005
R23040 DVSS.n12815 DVSS.n12792 4.5005
R23041 DVSS.n12815 DVSS.n12779 4.5005
R23042 DVSS.n12815 DVSS.n12790 4.5005
R23043 DVSS.n12815 DVSS.n12780 4.5005
R23044 DVSS.n12815 DVSS.n12789 4.5005
R23045 DVSS.n12815 DVSS.n12781 4.5005
R23046 DVSS.n12815 DVSS.n12787 4.5005
R23047 DVSS.n12815 DVSS.n12782 4.5005
R23048 DVSS.n12815 DVSS.n12786 4.5005
R23049 DVSS.n12815 DVSS.n12783 4.5005
R23050 DVSS.n12815 DVSS.n12785 4.5005
R23051 DVSS.n12799 DVSS.n12785 4.5005
R23052 DVSS.n12799 DVSS.n12783 4.5005
R23053 DVSS.n12799 DVSS.n12786 4.5005
R23054 DVSS.n12799 DVSS.n12782 4.5005
R23055 DVSS.n12799 DVSS.n12787 4.5005
R23056 DVSS.n12799 DVSS.n12781 4.5005
R23057 DVSS.n12799 DVSS.n12789 4.5005
R23058 DVSS.n12799 DVSS.n12780 4.5005
R23059 DVSS.n12799 DVSS.n12790 4.5005
R23060 DVSS.n12799 DVSS.n12779 4.5005
R23061 DVSS.n12799 DVSS.n12792 4.5005
R23062 DVSS.n12799 DVSS.n12778 4.5005
R23063 DVSS.n12799 DVSS.n12793 4.5005
R23064 DVSS.n12799 DVSS.n12777 4.5005
R23065 DVSS.n13099 DVSS.n12799 4.5005
R23066 DVSS.n12816 DVSS.n12785 4.5005
R23067 DVSS.n12816 DVSS.n12783 4.5005
R23068 DVSS.n12816 DVSS.n12786 4.5005
R23069 DVSS.n12816 DVSS.n12782 4.5005
R23070 DVSS.n12816 DVSS.n12787 4.5005
R23071 DVSS.n12816 DVSS.n12781 4.5005
R23072 DVSS.n12816 DVSS.n12789 4.5005
R23073 DVSS.n12816 DVSS.n12780 4.5005
R23074 DVSS.n12816 DVSS.n12790 4.5005
R23075 DVSS.n12816 DVSS.n12779 4.5005
R23076 DVSS.n12816 DVSS.n12792 4.5005
R23077 DVSS.n12816 DVSS.n12778 4.5005
R23078 DVSS.n12816 DVSS.n12793 4.5005
R23079 DVSS.n12816 DVSS.n12777 4.5005
R23080 DVSS.n13099 DVSS.n12816 4.5005
R23081 DVSS.n12798 DVSS.n12785 4.5005
R23082 DVSS.n12798 DVSS.n12783 4.5005
R23083 DVSS.n12798 DVSS.n12786 4.5005
R23084 DVSS.n12798 DVSS.n12782 4.5005
R23085 DVSS.n12798 DVSS.n12787 4.5005
R23086 DVSS.n12798 DVSS.n12781 4.5005
R23087 DVSS.n12798 DVSS.n12789 4.5005
R23088 DVSS.n12798 DVSS.n12780 4.5005
R23089 DVSS.n12798 DVSS.n12790 4.5005
R23090 DVSS.n12798 DVSS.n12779 4.5005
R23091 DVSS.n12798 DVSS.n12792 4.5005
R23092 DVSS.n12798 DVSS.n12778 4.5005
R23093 DVSS.n12798 DVSS.n12793 4.5005
R23094 DVSS.n12798 DVSS.n12777 4.5005
R23095 DVSS.n13099 DVSS.n12798 4.5005
R23096 DVSS.n12817 DVSS.n12777 4.5005
R23097 DVSS.n13099 DVSS.n12817 4.5005
R23098 DVSS.n12817 DVSS.n12793 4.5005
R23099 DVSS.n12817 DVSS.n12778 4.5005
R23100 DVSS.n12817 DVSS.n12792 4.5005
R23101 DVSS.n12817 DVSS.n12779 4.5005
R23102 DVSS.n12817 DVSS.n12790 4.5005
R23103 DVSS.n12817 DVSS.n12780 4.5005
R23104 DVSS.n12817 DVSS.n12789 4.5005
R23105 DVSS.n12817 DVSS.n12781 4.5005
R23106 DVSS.n12817 DVSS.n12787 4.5005
R23107 DVSS.n12817 DVSS.n12782 4.5005
R23108 DVSS.n12817 DVSS.n12786 4.5005
R23109 DVSS.n12817 DVSS.n12783 4.5005
R23110 DVSS.n12817 DVSS.n12785 4.5005
R23111 DVSS.n12797 DVSS.n12777 4.5005
R23112 DVSS.n13099 DVSS.n12797 4.5005
R23113 DVSS.n12797 DVSS.n12793 4.5005
R23114 DVSS.n12797 DVSS.n12778 4.5005
R23115 DVSS.n12797 DVSS.n12792 4.5005
R23116 DVSS.n12797 DVSS.n12779 4.5005
R23117 DVSS.n12797 DVSS.n12790 4.5005
R23118 DVSS.n12797 DVSS.n12780 4.5005
R23119 DVSS.n12797 DVSS.n12789 4.5005
R23120 DVSS.n12797 DVSS.n12781 4.5005
R23121 DVSS.n12797 DVSS.n12787 4.5005
R23122 DVSS.n12797 DVSS.n12782 4.5005
R23123 DVSS.n12797 DVSS.n12786 4.5005
R23124 DVSS.n12797 DVSS.n12783 4.5005
R23125 DVSS.n12797 DVSS.n12785 4.5005
R23126 DVSS.n12818 DVSS.n12777 4.5005
R23127 DVSS.n13099 DVSS.n12818 4.5005
R23128 DVSS.n12818 DVSS.n12793 4.5005
R23129 DVSS.n12818 DVSS.n12778 4.5005
R23130 DVSS.n12818 DVSS.n12792 4.5005
R23131 DVSS.n12818 DVSS.n12779 4.5005
R23132 DVSS.n12818 DVSS.n12790 4.5005
R23133 DVSS.n12818 DVSS.n12780 4.5005
R23134 DVSS.n12818 DVSS.n12789 4.5005
R23135 DVSS.n12818 DVSS.n12781 4.5005
R23136 DVSS.n12818 DVSS.n12787 4.5005
R23137 DVSS.n12818 DVSS.n12782 4.5005
R23138 DVSS.n12818 DVSS.n12786 4.5005
R23139 DVSS.n12818 DVSS.n12783 4.5005
R23140 DVSS.n12818 DVSS.n12785 4.5005
R23141 DVSS.n12796 DVSS.n12785 4.5005
R23142 DVSS.n12796 DVSS.n12783 4.5005
R23143 DVSS.n12796 DVSS.n12786 4.5005
R23144 DVSS.n12796 DVSS.n12782 4.5005
R23145 DVSS.n12796 DVSS.n12787 4.5005
R23146 DVSS.n12796 DVSS.n12781 4.5005
R23147 DVSS.n12796 DVSS.n12789 4.5005
R23148 DVSS.n12796 DVSS.n12780 4.5005
R23149 DVSS.n12796 DVSS.n12790 4.5005
R23150 DVSS.n12796 DVSS.n12779 4.5005
R23151 DVSS.n12796 DVSS.n12792 4.5005
R23152 DVSS.n12796 DVSS.n12778 4.5005
R23153 DVSS.n12796 DVSS.n12793 4.5005
R23154 DVSS.n12796 DVSS.n12777 4.5005
R23155 DVSS.n13099 DVSS.n12796 4.5005
R23156 DVSS.n13098 DVSS.n12785 4.5005
R23157 DVSS.n13098 DVSS.n12783 4.5005
R23158 DVSS.n13098 DVSS.n12786 4.5005
R23159 DVSS.n13098 DVSS.n12782 4.5005
R23160 DVSS.n13098 DVSS.n12787 4.5005
R23161 DVSS.n13098 DVSS.n12781 4.5005
R23162 DVSS.n13098 DVSS.n12789 4.5005
R23163 DVSS.n13098 DVSS.n12780 4.5005
R23164 DVSS.n13098 DVSS.n12790 4.5005
R23165 DVSS.n13098 DVSS.n12779 4.5005
R23166 DVSS.n13098 DVSS.n12792 4.5005
R23167 DVSS.n13098 DVSS.n12778 4.5005
R23168 DVSS.n13098 DVSS.n12793 4.5005
R23169 DVSS.n13098 DVSS.n12777 4.5005
R23170 DVSS.n13099 DVSS.n13098 4.5005
R23171 DVSS.n12795 DVSS.n12785 4.5005
R23172 DVSS.n12795 DVSS.n12783 4.5005
R23173 DVSS.n12795 DVSS.n12786 4.5005
R23174 DVSS.n12795 DVSS.n12782 4.5005
R23175 DVSS.n12795 DVSS.n12787 4.5005
R23176 DVSS.n12795 DVSS.n12781 4.5005
R23177 DVSS.n12795 DVSS.n12789 4.5005
R23178 DVSS.n12795 DVSS.n12780 4.5005
R23179 DVSS.n12795 DVSS.n12790 4.5005
R23180 DVSS.n12795 DVSS.n12779 4.5005
R23181 DVSS.n12795 DVSS.n12792 4.5005
R23182 DVSS.n12795 DVSS.n12778 4.5005
R23183 DVSS.n12795 DVSS.n12793 4.5005
R23184 DVSS.n12795 DVSS.n12777 4.5005
R23185 DVSS.n13099 DVSS.n12795 4.5005
R23186 DVSS.n13100 DVSS.n12785 4.5005
R23187 DVSS.n13100 DVSS.n12783 4.5005
R23188 DVSS.n13100 DVSS.n12786 4.5005
R23189 DVSS.n13100 DVSS.n12782 4.5005
R23190 DVSS.n13100 DVSS.n12787 4.5005
R23191 DVSS.n13100 DVSS.n12781 4.5005
R23192 DVSS.n13100 DVSS.n12789 4.5005
R23193 DVSS.n13100 DVSS.n12780 4.5005
R23194 DVSS.n13100 DVSS.n12790 4.5005
R23195 DVSS.n13100 DVSS.n12779 4.5005
R23196 DVSS.n13100 DVSS.n12792 4.5005
R23197 DVSS.n13100 DVSS.n12778 4.5005
R23198 DVSS.n13100 DVSS.n12793 4.5005
R23199 DVSS.n13100 DVSS.n12777 4.5005
R23200 DVSS.n13100 DVSS.n13099 4.5005
R23201 DVSS.n22435 DVSS.n1000 4.5005
R23202 DVSS.n1000 DVSS.n973 4.5005
R23203 DVSS.n1000 DVSS.n985 4.5005
R23204 DVSS.n1000 DVSS.n974 4.5005
R23205 DVSS.n1000 DVSS.n984 4.5005
R23206 DVSS.n1000 DVSS.n975 4.5005
R23207 DVSS.n1000 DVSS.n983 4.5005
R23208 DVSS.n1000 DVSS.n977 4.5005
R23209 DVSS.n1000 DVSS.n981 4.5005
R23210 DVSS.n1000 DVSS.n980 4.5005
R23211 DVSS.n1000 DVSS.n978 4.5005
R23212 DVSS.n22434 DVSS.n980 4.5005
R23213 DVSS.n22434 DVSS.n978 4.5005
R23214 DVSS.n988 DVSS.n980 4.5005
R23215 DVSS.n988 DVSS.n978 4.5005
R23216 DVSS.n1011 DVSS.n980 4.5005
R23217 DVSS.n1011 DVSS.n978 4.5005
R23218 DVSS.n22435 DVSS.n1002 4.5005
R23219 DVSS.n1002 DVSS.n972 4.5005
R23220 DVSS.n1002 DVSS.n986 4.5005
R23221 DVSS.n1002 DVSS.n973 4.5005
R23222 DVSS.n1002 DVSS.n985 4.5005
R23223 DVSS.n1002 DVSS.n974 4.5005
R23224 DVSS.n1002 DVSS.n984 4.5005
R23225 DVSS.n1002 DVSS.n975 4.5005
R23226 DVSS.n1002 DVSS.n983 4.5005
R23227 DVSS.n1002 DVSS.n976 4.5005
R23228 DVSS.n1002 DVSS.n982 4.5005
R23229 DVSS.n1002 DVSS.n977 4.5005
R23230 DVSS.n1002 DVSS.n981 4.5005
R23231 DVSS.n1002 DVSS.n980 4.5005
R23232 DVSS.n1002 DVSS.n978 4.5005
R23233 DVSS.n22435 DVSS.n997 4.5005
R23234 DVSS.n997 DVSS.n972 4.5005
R23235 DVSS.n997 DVSS.n986 4.5005
R23236 DVSS.n997 DVSS.n973 4.5005
R23237 DVSS.n997 DVSS.n985 4.5005
R23238 DVSS.n997 DVSS.n974 4.5005
R23239 DVSS.n997 DVSS.n984 4.5005
R23240 DVSS.n997 DVSS.n975 4.5005
R23241 DVSS.n997 DVSS.n983 4.5005
R23242 DVSS.n997 DVSS.n976 4.5005
R23243 DVSS.n997 DVSS.n982 4.5005
R23244 DVSS.n997 DVSS.n977 4.5005
R23245 DVSS.n997 DVSS.n981 4.5005
R23246 DVSS.n997 DVSS.n980 4.5005
R23247 DVSS.n997 DVSS.n978 4.5005
R23248 DVSS.n22435 DVSS.n1003 4.5005
R23249 DVSS.n1003 DVSS.n972 4.5005
R23250 DVSS.n1003 DVSS.n986 4.5005
R23251 DVSS.n1003 DVSS.n973 4.5005
R23252 DVSS.n1003 DVSS.n985 4.5005
R23253 DVSS.n1003 DVSS.n974 4.5005
R23254 DVSS.n1003 DVSS.n984 4.5005
R23255 DVSS.n1003 DVSS.n975 4.5005
R23256 DVSS.n1003 DVSS.n983 4.5005
R23257 DVSS.n1003 DVSS.n976 4.5005
R23258 DVSS.n1003 DVSS.n982 4.5005
R23259 DVSS.n1003 DVSS.n977 4.5005
R23260 DVSS.n1003 DVSS.n981 4.5005
R23261 DVSS.n1003 DVSS.n980 4.5005
R23262 DVSS.n1003 DVSS.n978 4.5005
R23263 DVSS.n989 DVSS.n980 4.5005
R23264 DVSS.n989 DVSS.n978 4.5005
R23265 DVSS.n1010 DVSS.n980 4.5005
R23266 DVSS.n1010 DVSS.n978 4.5005
R23267 DVSS.n990 DVSS.n980 4.5005
R23268 DVSS.n990 DVSS.n978 4.5005
R23269 DVSS.n22435 DVSS.n996 4.5005
R23270 DVSS.n996 DVSS.n972 4.5005
R23271 DVSS.n996 DVSS.n986 4.5005
R23272 DVSS.n996 DVSS.n973 4.5005
R23273 DVSS.n996 DVSS.n985 4.5005
R23274 DVSS.n996 DVSS.n974 4.5005
R23275 DVSS.n996 DVSS.n984 4.5005
R23276 DVSS.n996 DVSS.n975 4.5005
R23277 DVSS.n996 DVSS.n983 4.5005
R23278 DVSS.n996 DVSS.n976 4.5005
R23279 DVSS.n996 DVSS.n982 4.5005
R23280 DVSS.n996 DVSS.n977 4.5005
R23281 DVSS.n996 DVSS.n981 4.5005
R23282 DVSS.n996 DVSS.n980 4.5005
R23283 DVSS.n996 DVSS.n978 4.5005
R23284 DVSS.n22435 DVSS.n1004 4.5005
R23285 DVSS.n1004 DVSS.n972 4.5005
R23286 DVSS.n1004 DVSS.n986 4.5005
R23287 DVSS.n1004 DVSS.n973 4.5005
R23288 DVSS.n1004 DVSS.n985 4.5005
R23289 DVSS.n1004 DVSS.n974 4.5005
R23290 DVSS.n1004 DVSS.n984 4.5005
R23291 DVSS.n1004 DVSS.n975 4.5005
R23292 DVSS.n1004 DVSS.n983 4.5005
R23293 DVSS.n1004 DVSS.n976 4.5005
R23294 DVSS.n1004 DVSS.n982 4.5005
R23295 DVSS.n1004 DVSS.n977 4.5005
R23296 DVSS.n1004 DVSS.n981 4.5005
R23297 DVSS.n1004 DVSS.n980 4.5005
R23298 DVSS.n1004 DVSS.n978 4.5005
R23299 DVSS.n22435 DVSS.n995 4.5005
R23300 DVSS.n995 DVSS.n972 4.5005
R23301 DVSS.n995 DVSS.n986 4.5005
R23302 DVSS.n995 DVSS.n973 4.5005
R23303 DVSS.n995 DVSS.n985 4.5005
R23304 DVSS.n995 DVSS.n974 4.5005
R23305 DVSS.n995 DVSS.n984 4.5005
R23306 DVSS.n995 DVSS.n975 4.5005
R23307 DVSS.n995 DVSS.n983 4.5005
R23308 DVSS.n995 DVSS.n976 4.5005
R23309 DVSS.n995 DVSS.n982 4.5005
R23310 DVSS.n995 DVSS.n977 4.5005
R23311 DVSS.n995 DVSS.n981 4.5005
R23312 DVSS.n995 DVSS.n980 4.5005
R23313 DVSS.n995 DVSS.n978 4.5005
R23314 DVSS.n22435 DVSS.n1005 4.5005
R23315 DVSS.n1005 DVSS.n972 4.5005
R23316 DVSS.n1005 DVSS.n986 4.5005
R23317 DVSS.n1005 DVSS.n973 4.5005
R23318 DVSS.n1005 DVSS.n985 4.5005
R23319 DVSS.n1005 DVSS.n974 4.5005
R23320 DVSS.n1005 DVSS.n984 4.5005
R23321 DVSS.n1005 DVSS.n975 4.5005
R23322 DVSS.n1005 DVSS.n983 4.5005
R23323 DVSS.n1005 DVSS.n976 4.5005
R23324 DVSS.n1005 DVSS.n982 4.5005
R23325 DVSS.n1005 DVSS.n977 4.5005
R23326 DVSS.n1005 DVSS.n981 4.5005
R23327 DVSS.n1005 DVSS.n980 4.5005
R23328 DVSS.n1005 DVSS.n978 4.5005
R23329 DVSS.n1009 DVSS.n980 4.5005
R23330 DVSS.n1009 DVSS.n978 4.5005
R23331 DVSS.n991 DVSS.n980 4.5005
R23332 DVSS.n991 DVSS.n978 4.5005
R23333 DVSS.n1008 DVSS.n980 4.5005
R23334 DVSS.n1008 DVSS.n978 4.5005
R23335 DVSS.n22435 DVSS.n994 4.5005
R23336 DVSS.n994 DVSS.n972 4.5005
R23337 DVSS.n994 DVSS.n986 4.5005
R23338 DVSS.n994 DVSS.n973 4.5005
R23339 DVSS.n994 DVSS.n985 4.5005
R23340 DVSS.n994 DVSS.n974 4.5005
R23341 DVSS.n994 DVSS.n984 4.5005
R23342 DVSS.n994 DVSS.n975 4.5005
R23343 DVSS.n994 DVSS.n983 4.5005
R23344 DVSS.n994 DVSS.n976 4.5005
R23345 DVSS.n994 DVSS.n982 4.5005
R23346 DVSS.n994 DVSS.n977 4.5005
R23347 DVSS.n994 DVSS.n981 4.5005
R23348 DVSS.n994 DVSS.n980 4.5005
R23349 DVSS.n994 DVSS.n978 4.5005
R23350 DVSS.n22435 DVSS.n1006 4.5005
R23351 DVSS.n1006 DVSS.n972 4.5005
R23352 DVSS.n1006 DVSS.n986 4.5005
R23353 DVSS.n1006 DVSS.n973 4.5005
R23354 DVSS.n1006 DVSS.n985 4.5005
R23355 DVSS.n1006 DVSS.n974 4.5005
R23356 DVSS.n1006 DVSS.n984 4.5005
R23357 DVSS.n1006 DVSS.n975 4.5005
R23358 DVSS.n1006 DVSS.n983 4.5005
R23359 DVSS.n1006 DVSS.n976 4.5005
R23360 DVSS.n1006 DVSS.n982 4.5005
R23361 DVSS.n1006 DVSS.n977 4.5005
R23362 DVSS.n1006 DVSS.n981 4.5005
R23363 DVSS.n1006 DVSS.n980 4.5005
R23364 DVSS.n1006 DVSS.n978 4.5005
R23365 DVSS.n22435 DVSS.n993 4.5005
R23366 DVSS.n993 DVSS.n972 4.5005
R23367 DVSS.n993 DVSS.n986 4.5005
R23368 DVSS.n993 DVSS.n973 4.5005
R23369 DVSS.n993 DVSS.n985 4.5005
R23370 DVSS.n993 DVSS.n974 4.5005
R23371 DVSS.n993 DVSS.n984 4.5005
R23372 DVSS.n993 DVSS.n975 4.5005
R23373 DVSS.n993 DVSS.n983 4.5005
R23374 DVSS.n993 DVSS.n976 4.5005
R23375 DVSS.n993 DVSS.n982 4.5005
R23376 DVSS.n993 DVSS.n977 4.5005
R23377 DVSS.n993 DVSS.n981 4.5005
R23378 DVSS.n993 DVSS.n980 4.5005
R23379 DVSS.n993 DVSS.n978 4.5005
R23380 DVSS.n22435 DVSS.n1007 4.5005
R23381 DVSS.n1007 DVSS.n972 4.5005
R23382 DVSS.n1007 DVSS.n986 4.5005
R23383 DVSS.n1007 DVSS.n973 4.5005
R23384 DVSS.n1007 DVSS.n985 4.5005
R23385 DVSS.n1007 DVSS.n974 4.5005
R23386 DVSS.n1007 DVSS.n984 4.5005
R23387 DVSS.n1007 DVSS.n975 4.5005
R23388 DVSS.n1007 DVSS.n983 4.5005
R23389 DVSS.n1007 DVSS.n976 4.5005
R23390 DVSS.n1007 DVSS.n982 4.5005
R23391 DVSS.n1007 DVSS.n977 4.5005
R23392 DVSS.n1007 DVSS.n981 4.5005
R23393 DVSS.n1007 DVSS.n980 4.5005
R23394 DVSS.n1007 DVSS.n978 4.5005
R23395 DVSS.n992 DVSS.n980 4.5005
R23396 DVSS.n992 DVSS.n978 4.5005
R23397 DVSS.n22436 DVSS.n980 4.5005
R23398 DVSS.n22436 DVSS.n978 4.5005
R23399 DVSS.n980 DVSS.n970 4.5005
R23400 DVSS.n978 DVSS.n970 4.5005
R23401 DVSS.n981 DVSS.n970 4.5005
R23402 DVSS.n977 DVSS.n970 4.5005
R23403 DVSS.n982 DVSS.n970 4.5005
R23404 DVSS.n976 DVSS.n970 4.5005
R23405 DVSS.n983 DVSS.n970 4.5005
R23406 DVSS.n975 DVSS.n970 4.5005
R23407 DVSS.n984 DVSS.n970 4.5005
R23408 DVSS.n974 DVSS.n970 4.5005
R23409 DVSS.n985 DVSS.n970 4.5005
R23410 DVSS.n973 DVSS.n970 4.5005
R23411 DVSS.n986 DVSS.n970 4.5005
R23412 DVSS.n972 DVSS.n970 4.5005
R23413 DVSS.n22435 DVSS.n970 4.5005
R23414 DVSS.n22436 DVSS.n981 4.5005
R23415 DVSS.n22436 DVSS.n977 4.5005
R23416 DVSS.n22436 DVSS.n982 4.5005
R23417 DVSS.n22436 DVSS.n976 4.5005
R23418 DVSS.n22436 DVSS.n983 4.5005
R23419 DVSS.n22436 DVSS.n975 4.5005
R23420 DVSS.n22436 DVSS.n984 4.5005
R23421 DVSS.n22436 DVSS.n974 4.5005
R23422 DVSS.n22436 DVSS.n985 4.5005
R23423 DVSS.n22436 DVSS.n973 4.5005
R23424 DVSS.n22436 DVSS.n986 4.5005
R23425 DVSS.n22436 DVSS.n972 4.5005
R23426 DVSS.n22436 DVSS.n22435 4.5005
R23427 DVSS.n992 DVSS.n981 4.5005
R23428 DVSS.n992 DVSS.n977 4.5005
R23429 DVSS.n992 DVSS.n982 4.5005
R23430 DVSS.n992 DVSS.n976 4.5005
R23431 DVSS.n992 DVSS.n983 4.5005
R23432 DVSS.n992 DVSS.n975 4.5005
R23433 DVSS.n992 DVSS.n984 4.5005
R23434 DVSS.n992 DVSS.n974 4.5005
R23435 DVSS.n992 DVSS.n985 4.5005
R23436 DVSS.n992 DVSS.n973 4.5005
R23437 DVSS.n992 DVSS.n986 4.5005
R23438 DVSS.n992 DVSS.n972 4.5005
R23439 DVSS.n22435 DVSS.n992 4.5005
R23440 DVSS.n1008 DVSS.n981 4.5005
R23441 DVSS.n1008 DVSS.n977 4.5005
R23442 DVSS.n1008 DVSS.n982 4.5005
R23443 DVSS.n1008 DVSS.n976 4.5005
R23444 DVSS.n1008 DVSS.n983 4.5005
R23445 DVSS.n1008 DVSS.n975 4.5005
R23446 DVSS.n1008 DVSS.n984 4.5005
R23447 DVSS.n1008 DVSS.n974 4.5005
R23448 DVSS.n1008 DVSS.n985 4.5005
R23449 DVSS.n1008 DVSS.n973 4.5005
R23450 DVSS.n1008 DVSS.n986 4.5005
R23451 DVSS.n1008 DVSS.n972 4.5005
R23452 DVSS.n22435 DVSS.n1008 4.5005
R23453 DVSS.n991 DVSS.n981 4.5005
R23454 DVSS.n991 DVSS.n977 4.5005
R23455 DVSS.n991 DVSS.n982 4.5005
R23456 DVSS.n991 DVSS.n976 4.5005
R23457 DVSS.n991 DVSS.n983 4.5005
R23458 DVSS.n991 DVSS.n975 4.5005
R23459 DVSS.n991 DVSS.n984 4.5005
R23460 DVSS.n991 DVSS.n974 4.5005
R23461 DVSS.n991 DVSS.n985 4.5005
R23462 DVSS.n991 DVSS.n973 4.5005
R23463 DVSS.n991 DVSS.n986 4.5005
R23464 DVSS.n991 DVSS.n972 4.5005
R23465 DVSS.n22435 DVSS.n991 4.5005
R23466 DVSS.n1009 DVSS.n981 4.5005
R23467 DVSS.n1009 DVSS.n977 4.5005
R23468 DVSS.n1009 DVSS.n982 4.5005
R23469 DVSS.n1009 DVSS.n976 4.5005
R23470 DVSS.n1009 DVSS.n983 4.5005
R23471 DVSS.n1009 DVSS.n975 4.5005
R23472 DVSS.n1009 DVSS.n984 4.5005
R23473 DVSS.n1009 DVSS.n974 4.5005
R23474 DVSS.n1009 DVSS.n985 4.5005
R23475 DVSS.n1009 DVSS.n973 4.5005
R23476 DVSS.n1009 DVSS.n986 4.5005
R23477 DVSS.n1009 DVSS.n972 4.5005
R23478 DVSS.n22435 DVSS.n1009 4.5005
R23479 DVSS.n990 DVSS.n981 4.5005
R23480 DVSS.n990 DVSS.n977 4.5005
R23481 DVSS.n990 DVSS.n982 4.5005
R23482 DVSS.n990 DVSS.n976 4.5005
R23483 DVSS.n990 DVSS.n983 4.5005
R23484 DVSS.n990 DVSS.n975 4.5005
R23485 DVSS.n990 DVSS.n984 4.5005
R23486 DVSS.n990 DVSS.n974 4.5005
R23487 DVSS.n990 DVSS.n985 4.5005
R23488 DVSS.n990 DVSS.n973 4.5005
R23489 DVSS.n990 DVSS.n986 4.5005
R23490 DVSS.n990 DVSS.n972 4.5005
R23491 DVSS.n22435 DVSS.n990 4.5005
R23492 DVSS.n1010 DVSS.n981 4.5005
R23493 DVSS.n1010 DVSS.n977 4.5005
R23494 DVSS.n1010 DVSS.n982 4.5005
R23495 DVSS.n1010 DVSS.n976 4.5005
R23496 DVSS.n1010 DVSS.n983 4.5005
R23497 DVSS.n1010 DVSS.n975 4.5005
R23498 DVSS.n1010 DVSS.n984 4.5005
R23499 DVSS.n1010 DVSS.n974 4.5005
R23500 DVSS.n1010 DVSS.n985 4.5005
R23501 DVSS.n1010 DVSS.n973 4.5005
R23502 DVSS.n1010 DVSS.n986 4.5005
R23503 DVSS.n1010 DVSS.n972 4.5005
R23504 DVSS.n22435 DVSS.n1010 4.5005
R23505 DVSS.n989 DVSS.n981 4.5005
R23506 DVSS.n989 DVSS.n977 4.5005
R23507 DVSS.n989 DVSS.n982 4.5005
R23508 DVSS.n989 DVSS.n976 4.5005
R23509 DVSS.n989 DVSS.n983 4.5005
R23510 DVSS.n989 DVSS.n975 4.5005
R23511 DVSS.n989 DVSS.n984 4.5005
R23512 DVSS.n989 DVSS.n974 4.5005
R23513 DVSS.n989 DVSS.n985 4.5005
R23514 DVSS.n989 DVSS.n973 4.5005
R23515 DVSS.n989 DVSS.n986 4.5005
R23516 DVSS.n989 DVSS.n972 4.5005
R23517 DVSS.n22435 DVSS.n989 4.5005
R23518 DVSS.n1011 DVSS.n981 4.5005
R23519 DVSS.n1011 DVSS.n977 4.5005
R23520 DVSS.n1011 DVSS.n982 4.5005
R23521 DVSS.n1011 DVSS.n976 4.5005
R23522 DVSS.n1011 DVSS.n983 4.5005
R23523 DVSS.n1011 DVSS.n975 4.5005
R23524 DVSS.n1011 DVSS.n984 4.5005
R23525 DVSS.n1011 DVSS.n974 4.5005
R23526 DVSS.n1011 DVSS.n985 4.5005
R23527 DVSS.n1011 DVSS.n973 4.5005
R23528 DVSS.n1011 DVSS.n986 4.5005
R23529 DVSS.n1011 DVSS.n972 4.5005
R23530 DVSS.n22435 DVSS.n1011 4.5005
R23531 DVSS.n988 DVSS.n981 4.5005
R23532 DVSS.n988 DVSS.n977 4.5005
R23533 DVSS.n988 DVSS.n982 4.5005
R23534 DVSS.n988 DVSS.n976 4.5005
R23535 DVSS.n988 DVSS.n983 4.5005
R23536 DVSS.n988 DVSS.n975 4.5005
R23537 DVSS.n988 DVSS.n984 4.5005
R23538 DVSS.n988 DVSS.n974 4.5005
R23539 DVSS.n988 DVSS.n985 4.5005
R23540 DVSS.n988 DVSS.n973 4.5005
R23541 DVSS.n988 DVSS.n986 4.5005
R23542 DVSS.n988 DVSS.n972 4.5005
R23543 DVSS.n22435 DVSS.n988 4.5005
R23544 DVSS.n22434 DVSS.n981 4.5005
R23545 DVSS.n22434 DVSS.n977 4.5005
R23546 DVSS.n22434 DVSS.n982 4.5005
R23547 DVSS.n22434 DVSS.n976 4.5005
R23548 DVSS.n22434 DVSS.n983 4.5005
R23549 DVSS.n22434 DVSS.n975 4.5005
R23550 DVSS.n22434 DVSS.n984 4.5005
R23551 DVSS.n22434 DVSS.n974 4.5005
R23552 DVSS.n22434 DVSS.n985 4.5005
R23553 DVSS.n22434 DVSS.n973 4.5005
R23554 DVSS.n22434 DVSS.n986 4.5005
R23555 DVSS.n22434 DVSS.n972 4.5005
R23556 DVSS.n22435 DVSS.n22434 4.5005
R23557 DVSS.n1082 DVSS.n1059 4.5005
R23558 DVSS.n1082 DVSS.n1060 4.5005
R23559 DVSS.n1082 DVSS.n1058 4.5005
R23560 DVSS.n1082 DVSS.n1061 4.5005
R23561 DVSS.n1082 DVSS.n1057 4.5005
R23562 DVSS.n1082 DVSS.n1063 4.5005
R23563 DVSS.n1082 DVSS.n1055 4.5005
R23564 DVSS.n1082 DVSS.n1064 4.5005
R23565 DVSS.n1082 DVSS.n1054 4.5005
R23566 DVSS.n1082 DVSS.n1065 4.5005
R23567 DVSS.n1082 DVSS.n1053 4.5005
R23568 DVSS.n1082 DVSS.n1066 4.5005
R23569 DVSS.n22379 DVSS.n1082 4.5005
R23570 DVSS.n22380 DVSS.n1059 4.5005
R23571 DVSS.n22380 DVSS.n1060 4.5005
R23572 DVSS.n22380 DVSS.n1058 4.5005
R23573 DVSS.n22380 DVSS.n1061 4.5005
R23574 DVSS.n22380 DVSS.n1057 4.5005
R23575 DVSS.n22380 DVSS.n1062 4.5005
R23576 DVSS.n22380 DVSS.n1056 4.5005
R23577 DVSS.n22380 DVSS.n1063 4.5005
R23578 DVSS.n22380 DVSS.n1055 4.5005
R23579 DVSS.n22380 DVSS.n1064 4.5005
R23580 DVSS.n22380 DVSS.n1054 4.5005
R23581 DVSS.n22380 DVSS.n1065 4.5005
R23582 DVSS.n22380 DVSS.n1053 4.5005
R23583 DVSS.n22380 DVSS.n1066 4.5005
R23584 DVSS.n22380 DVSS.n22379 4.5005
R23585 DVSS.n1080 DVSS.n1059 4.5005
R23586 DVSS.n1080 DVSS.n1060 4.5005
R23587 DVSS.n1080 DVSS.n1058 4.5005
R23588 DVSS.n1080 DVSS.n1061 4.5005
R23589 DVSS.n1080 DVSS.n1057 4.5005
R23590 DVSS.n1080 DVSS.n1062 4.5005
R23591 DVSS.n1080 DVSS.n1056 4.5005
R23592 DVSS.n1080 DVSS.n1063 4.5005
R23593 DVSS.n1080 DVSS.n1055 4.5005
R23594 DVSS.n1080 DVSS.n1064 4.5005
R23595 DVSS.n1080 DVSS.n1054 4.5005
R23596 DVSS.n1080 DVSS.n1065 4.5005
R23597 DVSS.n1080 DVSS.n1066 4.5005
R23598 DVSS.n22379 DVSS.n1080 4.5005
R23599 DVSS.n1085 DVSS.n1059 4.5005
R23600 DVSS.n1085 DVSS.n1060 4.5005
R23601 DVSS.n1085 DVSS.n1058 4.5005
R23602 DVSS.n1085 DVSS.n1061 4.5005
R23603 DVSS.n1085 DVSS.n1057 4.5005
R23604 DVSS.n1085 DVSS.n1062 4.5005
R23605 DVSS.n1085 DVSS.n1056 4.5005
R23606 DVSS.n1085 DVSS.n1063 4.5005
R23607 DVSS.n1085 DVSS.n1055 4.5005
R23608 DVSS.n1085 DVSS.n1064 4.5005
R23609 DVSS.n1085 DVSS.n1054 4.5005
R23610 DVSS.n1085 DVSS.n1065 4.5005
R23611 DVSS.n1085 DVSS.n1066 4.5005
R23612 DVSS.n22379 DVSS.n1085 4.5005
R23613 DVSS.n1078 DVSS.n1059 4.5005
R23614 DVSS.n1078 DVSS.n1060 4.5005
R23615 DVSS.n1078 DVSS.n1058 4.5005
R23616 DVSS.n1078 DVSS.n1061 4.5005
R23617 DVSS.n1078 DVSS.n1057 4.5005
R23618 DVSS.n1078 DVSS.n1062 4.5005
R23619 DVSS.n1078 DVSS.n1056 4.5005
R23620 DVSS.n1078 DVSS.n1063 4.5005
R23621 DVSS.n1078 DVSS.n1055 4.5005
R23622 DVSS.n1078 DVSS.n1064 4.5005
R23623 DVSS.n1078 DVSS.n1054 4.5005
R23624 DVSS.n1078 DVSS.n1065 4.5005
R23625 DVSS.n22379 DVSS.n1078 4.5005
R23626 DVSS.n1086 DVSS.n1059 4.5005
R23627 DVSS.n1086 DVSS.n1060 4.5005
R23628 DVSS.n1086 DVSS.n1058 4.5005
R23629 DVSS.n1086 DVSS.n1061 4.5005
R23630 DVSS.n1086 DVSS.n1057 4.5005
R23631 DVSS.n1086 DVSS.n1062 4.5005
R23632 DVSS.n1086 DVSS.n1056 4.5005
R23633 DVSS.n1086 DVSS.n1063 4.5005
R23634 DVSS.n1086 DVSS.n1055 4.5005
R23635 DVSS.n1086 DVSS.n1064 4.5005
R23636 DVSS.n1086 DVSS.n1054 4.5005
R23637 DVSS.n1086 DVSS.n1065 4.5005
R23638 DVSS.n1086 DVSS.n1066 4.5005
R23639 DVSS.n22379 DVSS.n1086 4.5005
R23640 DVSS.n1077 DVSS.n1059 4.5005
R23641 DVSS.n1077 DVSS.n1060 4.5005
R23642 DVSS.n1077 DVSS.n1058 4.5005
R23643 DVSS.n1077 DVSS.n1061 4.5005
R23644 DVSS.n1077 DVSS.n1057 4.5005
R23645 DVSS.n1077 DVSS.n1062 4.5005
R23646 DVSS.n1077 DVSS.n1056 4.5005
R23647 DVSS.n1077 DVSS.n1063 4.5005
R23648 DVSS.n1077 DVSS.n1055 4.5005
R23649 DVSS.n1077 DVSS.n1064 4.5005
R23650 DVSS.n1077 DVSS.n1054 4.5005
R23651 DVSS.n1077 DVSS.n1065 4.5005
R23652 DVSS.n1077 DVSS.n1066 4.5005
R23653 DVSS.n22379 DVSS.n1077 4.5005
R23654 DVSS.n1088 DVSS.n1059 4.5005
R23655 DVSS.n1088 DVSS.n1060 4.5005
R23656 DVSS.n1088 DVSS.n1058 4.5005
R23657 DVSS.n1088 DVSS.n1061 4.5005
R23658 DVSS.n1088 DVSS.n1057 4.5005
R23659 DVSS.n1088 DVSS.n1062 4.5005
R23660 DVSS.n1088 DVSS.n1056 4.5005
R23661 DVSS.n1088 DVSS.n1063 4.5005
R23662 DVSS.n1088 DVSS.n1055 4.5005
R23663 DVSS.n1088 DVSS.n1064 4.5005
R23664 DVSS.n1088 DVSS.n1054 4.5005
R23665 DVSS.n1088 DVSS.n1065 4.5005
R23666 DVSS.n1088 DVSS.n1066 4.5005
R23667 DVSS.n1106 DVSS.n1088 4.5005
R23668 DVSS.n22379 DVSS.n1088 4.5005
R23669 DVSS.n1076 DVSS.n1059 4.5005
R23670 DVSS.n1076 DVSS.n1060 4.5005
R23671 DVSS.n1076 DVSS.n1058 4.5005
R23672 DVSS.n1076 DVSS.n1061 4.5005
R23673 DVSS.n1076 DVSS.n1057 4.5005
R23674 DVSS.n1076 DVSS.n1062 4.5005
R23675 DVSS.n1076 DVSS.n1056 4.5005
R23676 DVSS.n1076 DVSS.n1063 4.5005
R23677 DVSS.n1076 DVSS.n1055 4.5005
R23678 DVSS.n1076 DVSS.n1064 4.5005
R23679 DVSS.n1076 DVSS.n1054 4.5005
R23680 DVSS.n1076 DVSS.n1065 4.5005
R23681 DVSS.n1076 DVSS.n1066 4.5005
R23682 DVSS.n22379 DVSS.n1076 4.5005
R23683 DVSS.n1090 DVSS.n1059 4.5005
R23684 DVSS.n1090 DVSS.n1060 4.5005
R23685 DVSS.n1090 DVSS.n1058 4.5005
R23686 DVSS.n1090 DVSS.n1061 4.5005
R23687 DVSS.n1090 DVSS.n1057 4.5005
R23688 DVSS.n1090 DVSS.n1062 4.5005
R23689 DVSS.n1090 DVSS.n1056 4.5005
R23690 DVSS.n1090 DVSS.n1063 4.5005
R23691 DVSS.n1090 DVSS.n1055 4.5005
R23692 DVSS.n1090 DVSS.n1064 4.5005
R23693 DVSS.n1090 DVSS.n1054 4.5005
R23694 DVSS.n1090 DVSS.n1065 4.5005
R23695 DVSS.n1090 DVSS.n1066 4.5005
R23696 DVSS.n22379 DVSS.n1090 4.5005
R23697 DVSS.n1074 DVSS.n1059 4.5005
R23698 DVSS.n1074 DVSS.n1060 4.5005
R23699 DVSS.n1074 DVSS.n1058 4.5005
R23700 DVSS.n1074 DVSS.n1061 4.5005
R23701 DVSS.n1074 DVSS.n1057 4.5005
R23702 DVSS.n1074 DVSS.n1062 4.5005
R23703 DVSS.n1074 DVSS.n1056 4.5005
R23704 DVSS.n1074 DVSS.n1063 4.5005
R23705 DVSS.n1074 DVSS.n1055 4.5005
R23706 DVSS.n1074 DVSS.n1064 4.5005
R23707 DVSS.n1074 DVSS.n1054 4.5005
R23708 DVSS.n1074 DVSS.n1065 4.5005
R23709 DVSS.n1074 DVSS.n1066 4.5005
R23710 DVSS.n1106 DVSS.n1074 4.5005
R23711 DVSS.n22379 DVSS.n1074 4.5005
R23712 DVSS.n1091 DVSS.n1059 4.5005
R23713 DVSS.n1091 DVSS.n1060 4.5005
R23714 DVSS.n1091 DVSS.n1058 4.5005
R23715 DVSS.n1091 DVSS.n1061 4.5005
R23716 DVSS.n1091 DVSS.n1057 4.5005
R23717 DVSS.n1091 DVSS.n1062 4.5005
R23718 DVSS.n1091 DVSS.n1056 4.5005
R23719 DVSS.n1091 DVSS.n1063 4.5005
R23720 DVSS.n1091 DVSS.n1055 4.5005
R23721 DVSS.n1091 DVSS.n1064 4.5005
R23722 DVSS.n1091 DVSS.n1054 4.5005
R23723 DVSS.n1091 DVSS.n1065 4.5005
R23724 DVSS.n1091 DVSS.n1066 4.5005
R23725 DVSS.n22379 DVSS.n1091 4.5005
R23726 DVSS.n1073 DVSS.n1059 4.5005
R23727 DVSS.n1073 DVSS.n1060 4.5005
R23728 DVSS.n1073 DVSS.n1058 4.5005
R23729 DVSS.n1073 DVSS.n1061 4.5005
R23730 DVSS.n1073 DVSS.n1057 4.5005
R23731 DVSS.n1073 DVSS.n1062 4.5005
R23732 DVSS.n1073 DVSS.n1056 4.5005
R23733 DVSS.n1073 DVSS.n1063 4.5005
R23734 DVSS.n1073 DVSS.n1055 4.5005
R23735 DVSS.n1073 DVSS.n1064 4.5005
R23736 DVSS.n1073 DVSS.n1054 4.5005
R23737 DVSS.n1073 DVSS.n1065 4.5005
R23738 DVSS.n1073 DVSS.n1066 4.5005
R23739 DVSS.n22379 DVSS.n1073 4.5005
R23740 DVSS.n1093 DVSS.n1059 4.5005
R23741 DVSS.n1093 DVSS.n1060 4.5005
R23742 DVSS.n1093 DVSS.n1058 4.5005
R23743 DVSS.n1093 DVSS.n1061 4.5005
R23744 DVSS.n1093 DVSS.n1057 4.5005
R23745 DVSS.n1093 DVSS.n1062 4.5005
R23746 DVSS.n1093 DVSS.n1056 4.5005
R23747 DVSS.n1093 DVSS.n1063 4.5005
R23748 DVSS.n1093 DVSS.n1055 4.5005
R23749 DVSS.n1093 DVSS.n1064 4.5005
R23750 DVSS.n1093 DVSS.n1054 4.5005
R23751 DVSS.n1093 DVSS.n1065 4.5005
R23752 DVSS.n1093 DVSS.n1066 4.5005
R23753 DVSS.n1106 DVSS.n1093 4.5005
R23754 DVSS.n22379 DVSS.n1093 4.5005
R23755 DVSS.n1072 DVSS.n1059 4.5005
R23756 DVSS.n1072 DVSS.n1060 4.5005
R23757 DVSS.n1072 DVSS.n1058 4.5005
R23758 DVSS.n1072 DVSS.n1061 4.5005
R23759 DVSS.n1072 DVSS.n1057 4.5005
R23760 DVSS.n1072 DVSS.n1062 4.5005
R23761 DVSS.n1072 DVSS.n1056 4.5005
R23762 DVSS.n1072 DVSS.n1063 4.5005
R23763 DVSS.n1072 DVSS.n1055 4.5005
R23764 DVSS.n1072 DVSS.n1064 4.5005
R23765 DVSS.n1072 DVSS.n1054 4.5005
R23766 DVSS.n1072 DVSS.n1065 4.5005
R23767 DVSS.n1072 DVSS.n1066 4.5005
R23768 DVSS.n22379 DVSS.n1072 4.5005
R23769 DVSS.n1095 DVSS.n1059 4.5005
R23770 DVSS.n1095 DVSS.n1060 4.5005
R23771 DVSS.n1095 DVSS.n1058 4.5005
R23772 DVSS.n1095 DVSS.n1061 4.5005
R23773 DVSS.n1095 DVSS.n1057 4.5005
R23774 DVSS.n1095 DVSS.n1062 4.5005
R23775 DVSS.n1095 DVSS.n1056 4.5005
R23776 DVSS.n1095 DVSS.n1063 4.5005
R23777 DVSS.n1095 DVSS.n1055 4.5005
R23778 DVSS.n1095 DVSS.n1064 4.5005
R23779 DVSS.n1095 DVSS.n1054 4.5005
R23780 DVSS.n1095 DVSS.n1065 4.5005
R23781 DVSS.n1095 DVSS.n1066 4.5005
R23782 DVSS.n22379 DVSS.n1095 4.5005
R23783 DVSS.n1070 DVSS.n1059 4.5005
R23784 DVSS.n1070 DVSS.n1060 4.5005
R23785 DVSS.n1070 DVSS.n1058 4.5005
R23786 DVSS.n1070 DVSS.n1061 4.5005
R23787 DVSS.n1070 DVSS.n1057 4.5005
R23788 DVSS.n1070 DVSS.n1062 4.5005
R23789 DVSS.n1070 DVSS.n1056 4.5005
R23790 DVSS.n1070 DVSS.n1063 4.5005
R23791 DVSS.n1070 DVSS.n1055 4.5005
R23792 DVSS.n1070 DVSS.n1064 4.5005
R23793 DVSS.n1070 DVSS.n1054 4.5005
R23794 DVSS.n1070 DVSS.n1065 4.5005
R23795 DVSS.n1070 DVSS.n1066 4.5005
R23796 DVSS.n1106 DVSS.n1070 4.5005
R23797 DVSS.n22379 DVSS.n1070 4.5005
R23798 DVSS.n1096 DVSS.n1059 4.5005
R23799 DVSS.n1096 DVSS.n1060 4.5005
R23800 DVSS.n1096 DVSS.n1058 4.5005
R23801 DVSS.n1096 DVSS.n1061 4.5005
R23802 DVSS.n1096 DVSS.n1057 4.5005
R23803 DVSS.n1096 DVSS.n1062 4.5005
R23804 DVSS.n1096 DVSS.n1056 4.5005
R23805 DVSS.n1096 DVSS.n1063 4.5005
R23806 DVSS.n1096 DVSS.n1055 4.5005
R23807 DVSS.n1096 DVSS.n1064 4.5005
R23808 DVSS.n1096 DVSS.n1054 4.5005
R23809 DVSS.n1096 DVSS.n1065 4.5005
R23810 DVSS.n1096 DVSS.n1053 4.5005
R23811 DVSS.n1096 DVSS.n1066 4.5005
R23812 DVSS.n1106 DVSS.n1096 4.5005
R23813 DVSS.n22379 DVSS.n1096 4.5005
R23814 DVSS.n1069 DVSS.n1059 4.5005
R23815 DVSS.n1069 DVSS.n1060 4.5005
R23816 DVSS.n1069 DVSS.n1058 4.5005
R23817 DVSS.n1069 DVSS.n1061 4.5005
R23818 DVSS.n1069 DVSS.n1057 4.5005
R23819 DVSS.n1069 DVSS.n1062 4.5005
R23820 DVSS.n1069 DVSS.n1056 4.5005
R23821 DVSS.n1069 DVSS.n1063 4.5005
R23822 DVSS.n1069 DVSS.n1055 4.5005
R23823 DVSS.n1069 DVSS.n1064 4.5005
R23824 DVSS.n1069 DVSS.n1054 4.5005
R23825 DVSS.n1069 DVSS.n1065 4.5005
R23826 DVSS.n1069 DVSS.n1066 4.5005
R23827 DVSS.n1106 DVSS.n1069 4.5005
R23828 DVSS.n22379 DVSS.n1069 4.5005
R23829 DVSS.n1098 DVSS.n1059 4.5005
R23830 DVSS.n1098 DVSS.n1060 4.5005
R23831 DVSS.n1098 DVSS.n1058 4.5005
R23832 DVSS.n1098 DVSS.n1061 4.5005
R23833 DVSS.n1098 DVSS.n1057 4.5005
R23834 DVSS.n1098 DVSS.n1062 4.5005
R23835 DVSS.n1098 DVSS.n1056 4.5005
R23836 DVSS.n1098 DVSS.n1063 4.5005
R23837 DVSS.n1098 DVSS.n1055 4.5005
R23838 DVSS.n1098 DVSS.n1064 4.5005
R23839 DVSS.n1098 DVSS.n1054 4.5005
R23840 DVSS.n1098 DVSS.n1065 4.5005
R23841 DVSS.n1098 DVSS.n1066 4.5005
R23842 DVSS.n1106 DVSS.n1098 4.5005
R23843 DVSS.n22379 DVSS.n1098 4.5005
R23844 DVSS.n1068 DVSS.n1059 4.5005
R23845 DVSS.n1068 DVSS.n1060 4.5005
R23846 DVSS.n1068 DVSS.n1058 4.5005
R23847 DVSS.n1068 DVSS.n1061 4.5005
R23848 DVSS.n1068 DVSS.n1057 4.5005
R23849 DVSS.n1068 DVSS.n1062 4.5005
R23850 DVSS.n1068 DVSS.n1056 4.5005
R23851 DVSS.n1068 DVSS.n1063 4.5005
R23852 DVSS.n1068 DVSS.n1055 4.5005
R23853 DVSS.n1068 DVSS.n1064 4.5005
R23854 DVSS.n1068 DVSS.n1054 4.5005
R23855 DVSS.n1068 DVSS.n1065 4.5005
R23856 DVSS.n1068 DVSS.n1066 4.5005
R23857 DVSS.n1106 DVSS.n1068 4.5005
R23858 DVSS.n22379 DVSS.n1068 4.5005
R23859 DVSS.n22378 DVSS.n1059 4.5005
R23860 DVSS.n22378 DVSS.n1060 4.5005
R23861 DVSS.n22378 DVSS.n1058 4.5005
R23862 DVSS.n22378 DVSS.n1061 4.5005
R23863 DVSS.n22378 DVSS.n1057 4.5005
R23864 DVSS.n22378 DVSS.n1062 4.5005
R23865 DVSS.n22378 DVSS.n1056 4.5005
R23866 DVSS.n22378 DVSS.n1063 4.5005
R23867 DVSS.n22378 DVSS.n1055 4.5005
R23868 DVSS.n22378 DVSS.n1064 4.5005
R23869 DVSS.n22378 DVSS.n1054 4.5005
R23870 DVSS.n22378 DVSS.n1065 4.5005
R23871 DVSS.n22378 DVSS.n1066 4.5005
R23872 DVSS.n22378 DVSS.n1106 4.5005
R23873 DVSS.n22379 DVSS.n22378 4.5005
R23874 DVSS.n1059 DVSS.n1017 4.5005
R23875 DVSS.n1060 DVSS.n1017 4.5005
R23876 DVSS.n1058 DVSS.n1017 4.5005
R23877 DVSS.n1061 DVSS.n1017 4.5005
R23878 DVSS.n1057 DVSS.n1017 4.5005
R23879 DVSS.n1062 DVSS.n1017 4.5005
R23880 DVSS.n1056 DVSS.n1017 4.5005
R23881 DVSS.n1063 DVSS.n1017 4.5005
R23882 DVSS.n1055 DVSS.n1017 4.5005
R23883 DVSS.n1064 DVSS.n1017 4.5005
R23884 DVSS.n1054 DVSS.n1017 4.5005
R23885 DVSS.n1065 DVSS.n1017 4.5005
R23886 DVSS.n1066 DVSS.n1017 4.5005
R23887 DVSS.n1106 DVSS.n1017 4.5005
R23888 DVSS.n22379 DVSS.n1017 4.5005
R23889 DVSS.n1059 DVSS.n1026 4.5005
R23890 DVSS.n1060 DVSS.n1026 4.5005
R23891 DVSS.n1058 DVSS.n1026 4.5005
R23892 DVSS.n1061 DVSS.n1026 4.5005
R23893 DVSS.n1057 DVSS.n1026 4.5005
R23894 DVSS.n1062 DVSS.n1026 4.5005
R23895 DVSS.n1056 DVSS.n1026 4.5005
R23896 DVSS.n1063 DVSS.n1026 4.5005
R23897 DVSS.n1055 DVSS.n1026 4.5005
R23898 DVSS.n1064 DVSS.n1026 4.5005
R23899 DVSS.n1054 DVSS.n1026 4.5005
R23900 DVSS.n1065 DVSS.n1026 4.5005
R23901 DVSS.n1053 DVSS.n1026 4.5005
R23902 DVSS.n1066 DVSS.n1026 4.5005
R23903 DVSS.n1106 DVSS.n1026 4.5005
R23904 DVSS.n22379 DVSS.n1026 4.5005
R23905 DVSS.n1136 DVSS.n1115 4.5005
R23906 DVSS.n1136 DVSS.n1116 4.5005
R23907 DVSS.n1136 DVSS.n1114 4.5005
R23908 DVSS.n1136 DVSS.n1118 4.5005
R23909 DVSS.n1136 DVSS.n1112 4.5005
R23910 DVSS.n1136 DVSS.n1119 4.5005
R23911 DVSS.n1136 DVSS.n1111 4.5005
R23912 DVSS.n1136 DVSS.n1121 4.5005
R23913 DVSS.n1136 DVSS.n1110 4.5005
R23914 DVSS.n1136 DVSS.n1124 4.5005
R23915 DVSS.n22373 DVSS.n1136 4.5005
R23916 DVSS.n1138 DVSS.n1115 4.5005
R23917 DVSS.n1138 DVSS.n1116 4.5005
R23918 DVSS.n1138 DVSS.n1114 4.5005
R23919 DVSS.n1138 DVSS.n1117 4.5005
R23920 DVSS.n1138 DVSS.n1113 4.5005
R23921 DVSS.n1138 DVSS.n1118 4.5005
R23922 DVSS.n1138 DVSS.n1112 4.5005
R23923 DVSS.n1138 DVSS.n1119 4.5005
R23924 DVSS.n1138 DVSS.n1111 4.5005
R23925 DVSS.n1138 DVSS.n1121 4.5005
R23926 DVSS.n1138 DVSS.n1110 4.5005
R23927 DVSS.n1138 DVSS.n1122 4.5005
R23928 DVSS.n1164 DVSS.n1138 4.5005
R23929 DVSS.n1138 DVSS.n1124 4.5005
R23930 DVSS.n22373 DVSS.n1138 4.5005
R23931 DVSS.n1134 DVSS.n1115 4.5005
R23932 DVSS.n1134 DVSS.n1116 4.5005
R23933 DVSS.n1134 DVSS.n1114 4.5005
R23934 DVSS.n1134 DVSS.n1117 4.5005
R23935 DVSS.n1134 DVSS.n1113 4.5005
R23936 DVSS.n1134 DVSS.n1118 4.5005
R23937 DVSS.n1134 DVSS.n1112 4.5005
R23938 DVSS.n1134 DVSS.n1119 4.5005
R23939 DVSS.n1134 DVSS.n1111 4.5005
R23940 DVSS.n1134 DVSS.n1121 4.5005
R23941 DVSS.n1134 DVSS.n1110 4.5005
R23942 DVSS.n1134 DVSS.n1122 4.5005
R23943 DVSS.n1134 DVSS.n1124 4.5005
R23944 DVSS.n22373 DVSS.n1134 4.5005
R23945 DVSS.n1140 DVSS.n1115 4.5005
R23946 DVSS.n1140 DVSS.n1116 4.5005
R23947 DVSS.n1140 DVSS.n1114 4.5005
R23948 DVSS.n1140 DVSS.n1117 4.5005
R23949 DVSS.n1140 DVSS.n1113 4.5005
R23950 DVSS.n1140 DVSS.n1118 4.5005
R23951 DVSS.n1140 DVSS.n1112 4.5005
R23952 DVSS.n1140 DVSS.n1119 4.5005
R23953 DVSS.n1140 DVSS.n1111 4.5005
R23954 DVSS.n1140 DVSS.n1121 4.5005
R23955 DVSS.n1140 DVSS.n1110 4.5005
R23956 DVSS.n1140 DVSS.n1122 4.5005
R23957 DVSS.n1140 DVSS.n1124 4.5005
R23958 DVSS.n22373 DVSS.n1140 4.5005
R23959 DVSS.n22374 DVSS.n1115 4.5005
R23960 DVSS.n22374 DVSS.n1116 4.5005
R23961 DVSS.n22374 DVSS.n1114 4.5005
R23962 DVSS.n22374 DVSS.n1117 4.5005
R23963 DVSS.n22374 DVSS.n1113 4.5005
R23964 DVSS.n22374 DVSS.n1118 4.5005
R23965 DVSS.n22374 DVSS.n1112 4.5005
R23966 DVSS.n22374 DVSS.n1119 4.5005
R23967 DVSS.n22374 DVSS.n1111 4.5005
R23968 DVSS.n22374 DVSS.n1121 4.5005
R23969 DVSS.n22374 DVSS.n1110 4.5005
R23970 DVSS.n22374 DVSS.n1122 4.5005
R23971 DVSS.n22374 DVSS.n1124 4.5005
R23972 DVSS.n22374 DVSS.n1108 4.5005
R23973 DVSS.n22374 DVSS.n22373 4.5005
R23974 DVSS.n1142 DVSS.n1115 4.5005
R23975 DVSS.n1142 DVSS.n1116 4.5005
R23976 DVSS.n1142 DVSS.n1114 4.5005
R23977 DVSS.n1142 DVSS.n1117 4.5005
R23978 DVSS.n1142 DVSS.n1113 4.5005
R23979 DVSS.n1142 DVSS.n1118 4.5005
R23980 DVSS.n1142 DVSS.n1112 4.5005
R23981 DVSS.n1142 DVSS.n1119 4.5005
R23982 DVSS.n1142 DVSS.n1111 4.5005
R23983 DVSS.n1142 DVSS.n1121 4.5005
R23984 DVSS.n1142 DVSS.n1110 4.5005
R23985 DVSS.n1142 DVSS.n1122 4.5005
R23986 DVSS.n1142 DVSS.n1124 4.5005
R23987 DVSS.n22373 DVSS.n1142 4.5005
R23988 DVSS.n1133 DVSS.n1115 4.5005
R23989 DVSS.n1133 DVSS.n1116 4.5005
R23990 DVSS.n1133 DVSS.n1114 4.5005
R23991 DVSS.n1133 DVSS.n1117 4.5005
R23992 DVSS.n1133 DVSS.n1113 4.5005
R23993 DVSS.n1133 DVSS.n1118 4.5005
R23994 DVSS.n1133 DVSS.n1112 4.5005
R23995 DVSS.n1133 DVSS.n1119 4.5005
R23996 DVSS.n1133 DVSS.n1111 4.5005
R23997 DVSS.n1133 DVSS.n1121 4.5005
R23998 DVSS.n1133 DVSS.n1110 4.5005
R23999 DVSS.n1133 DVSS.n1122 4.5005
R24000 DVSS.n1133 DVSS.n1124 4.5005
R24001 DVSS.n22373 DVSS.n1133 4.5005
R24002 DVSS.n1143 DVSS.n1115 4.5005
R24003 DVSS.n1143 DVSS.n1116 4.5005
R24004 DVSS.n1143 DVSS.n1114 4.5005
R24005 DVSS.n1143 DVSS.n1117 4.5005
R24006 DVSS.n1143 DVSS.n1113 4.5005
R24007 DVSS.n1143 DVSS.n1118 4.5005
R24008 DVSS.n1143 DVSS.n1112 4.5005
R24009 DVSS.n1143 DVSS.n1119 4.5005
R24010 DVSS.n1143 DVSS.n1111 4.5005
R24011 DVSS.n1143 DVSS.n1121 4.5005
R24012 DVSS.n1143 DVSS.n1110 4.5005
R24013 DVSS.n1143 DVSS.n1122 4.5005
R24014 DVSS.n1143 DVSS.n1124 4.5005
R24015 DVSS.n1143 DVSS.n1108 4.5005
R24016 DVSS.n22373 DVSS.n1143 4.5005
R24017 DVSS.n1132 DVSS.n1115 4.5005
R24018 DVSS.n1132 DVSS.n1116 4.5005
R24019 DVSS.n1132 DVSS.n1114 4.5005
R24020 DVSS.n1132 DVSS.n1117 4.5005
R24021 DVSS.n1132 DVSS.n1113 4.5005
R24022 DVSS.n1132 DVSS.n1118 4.5005
R24023 DVSS.n1132 DVSS.n1112 4.5005
R24024 DVSS.n1132 DVSS.n1119 4.5005
R24025 DVSS.n1132 DVSS.n1111 4.5005
R24026 DVSS.n1132 DVSS.n1121 4.5005
R24027 DVSS.n1132 DVSS.n1110 4.5005
R24028 DVSS.n1132 DVSS.n1122 4.5005
R24029 DVSS.n1132 DVSS.n1124 4.5005
R24030 DVSS.n22373 DVSS.n1132 4.5005
R24031 DVSS.n1145 DVSS.n1115 4.5005
R24032 DVSS.n1145 DVSS.n1116 4.5005
R24033 DVSS.n1145 DVSS.n1114 4.5005
R24034 DVSS.n1145 DVSS.n1117 4.5005
R24035 DVSS.n1145 DVSS.n1113 4.5005
R24036 DVSS.n1145 DVSS.n1118 4.5005
R24037 DVSS.n1145 DVSS.n1112 4.5005
R24038 DVSS.n1145 DVSS.n1119 4.5005
R24039 DVSS.n1145 DVSS.n1111 4.5005
R24040 DVSS.n1145 DVSS.n1121 4.5005
R24041 DVSS.n1145 DVSS.n1110 4.5005
R24042 DVSS.n1145 DVSS.n1122 4.5005
R24043 DVSS.n1145 DVSS.n1124 4.5005
R24044 DVSS.n22373 DVSS.n1145 4.5005
R24045 DVSS.n1131 DVSS.n1115 4.5005
R24046 DVSS.n1131 DVSS.n1116 4.5005
R24047 DVSS.n1131 DVSS.n1114 4.5005
R24048 DVSS.n1131 DVSS.n1117 4.5005
R24049 DVSS.n1131 DVSS.n1113 4.5005
R24050 DVSS.n1131 DVSS.n1118 4.5005
R24051 DVSS.n1131 DVSS.n1112 4.5005
R24052 DVSS.n1131 DVSS.n1119 4.5005
R24053 DVSS.n1131 DVSS.n1111 4.5005
R24054 DVSS.n1131 DVSS.n1121 4.5005
R24055 DVSS.n1131 DVSS.n1110 4.5005
R24056 DVSS.n1131 DVSS.n1122 4.5005
R24057 DVSS.n1131 DVSS.n1124 4.5005
R24058 DVSS.n1131 DVSS.n1108 4.5005
R24059 DVSS.n22373 DVSS.n1131 4.5005
R24060 DVSS.n1147 DVSS.n1115 4.5005
R24061 DVSS.n1147 DVSS.n1116 4.5005
R24062 DVSS.n1147 DVSS.n1114 4.5005
R24063 DVSS.n1147 DVSS.n1117 4.5005
R24064 DVSS.n1147 DVSS.n1113 4.5005
R24065 DVSS.n1147 DVSS.n1118 4.5005
R24066 DVSS.n1147 DVSS.n1112 4.5005
R24067 DVSS.n1147 DVSS.n1119 4.5005
R24068 DVSS.n1147 DVSS.n1111 4.5005
R24069 DVSS.n1147 DVSS.n1121 4.5005
R24070 DVSS.n1147 DVSS.n1110 4.5005
R24071 DVSS.n1147 DVSS.n1122 4.5005
R24072 DVSS.n1147 DVSS.n1124 4.5005
R24073 DVSS.n22373 DVSS.n1147 4.5005
R24074 DVSS.n1130 DVSS.n1115 4.5005
R24075 DVSS.n1130 DVSS.n1116 4.5005
R24076 DVSS.n1130 DVSS.n1114 4.5005
R24077 DVSS.n1130 DVSS.n1117 4.5005
R24078 DVSS.n1130 DVSS.n1113 4.5005
R24079 DVSS.n1130 DVSS.n1118 4.5005
R24080 DVSS.n1130 DVSS.n1112 4.5005
R24081 DVSS.n1130 DVSS.n1119 4.5005
R24082 DVSS.n1130 DVSS.n1111 4.5005
R24083 DVSS.n1130 DVSS.n1121 4.5005
R24084 DVSS.n1130 DVSS.n1110 4.5005
R24085 DVSS.n1130 DVSS.n1122 4.5005
R24086 DVSS.n1130 DVSS.n1124 4.5005
R24087 DVSS.n22373 DVSS.n1130 4.5005
R24088 DVSS.n1148 DVSS.n1115 4.5005
R24089 DVSS.n1148 DVSS.n1116 4.5005
R24090 DVSS.n1148 DVSS.n1114 4.5005
R24091 DVSS.n1148 DVSS.n1117 4.5005
R24092 DVSS.n1148 DVSS.n1113 4.5005
R24093 DVSS.n1148 DVSS.n1118 4.5005
R24094 DVSS.n1148 DVSS.n1112 4.5005
R24095 DVSS.n1148 DVSS.n1119 4.5005
R24096 DVSS.n1148 DVSS.n1111 4.5005
R24097 DVSS.n1148 DVSS.n1121 4.5005
R24098 DVSS.n1148 DVSS.n1110 4.5005
R24099 DVSS.n1148 DVSS.n1122 4.5005
R24100 DVSS.n1148 DVSS.n1124 4.5005
R24101 DVSS.n1148 DVSS.n1108 4.5005
R24102 DVSS.n22373 DVSS.n1148 4.5005
R24103 DVSS.n1129 DVSS.n1115 4.5005
R24104 DVSS.n1129 DVSS.n1116 4.5005
R24105 DVSS.n1129 DVSS.n1114 4.5005
R24106 DVSS.n1129 DVSS.n1117 4.5005
R24107 DVSS.n1129 DVSS.n1113 4.5005
R24108 DVSS.n1129 DVSS.n1118 4.5005
R24109 DVSS.n1129 DVSS.n1112 4.5005
R24110 DVSS.n1129 DVSS.n1119 4.5005
R24111 DVSS.n1129 DVSS.n1111 4.5005
R24112 DVSS.n1129 DVSS.n1121 4.5005
R24113 DVSS.n1129 DVSS.n1110 4.5005
R24114 DVSS.n1129 DVSS.n1122 4.5005
R24115 DVSS.n1129 DVSS.n1124 4.5005
R24116 DVSS.n22373 DVSS.n1129 4.5005
R24117 DVSS.n1150 DVSS.n1115 4.5005
R24118 DVSS.n1150 DVSS.n1116 4.5005
R24119 DVSS.n1150 DVSS.n1114 4.5005
R24120 DVSS.n1150 DVSS.n1117 4.5005
R24121 DVSS.n1150 DVSS.n1113 4.5005
R24122 DVSS.n1150 DVSS.n1118 4.5005
R24123 DVSS.n1150 DVSS.n1112 4.5005
R24124 DVSS.n1150 DVSS.n1119 4.5005
R24125 DVSS.n1150 DVSS.n1111 4.5005
R24126 DVSS.n1150 DVSS.n1121 4.5005
R24127 DVSS.n1150 DVSS.n1110 4.5005
R24128 DVSS.n1150 DVSS.n1122 4.5005
R24129 DVSS.n1150 DVSS.n1124 4.5005
R24130 DVSS.n22373 DVSS.n1150 4.5005
R24131 DVSS.n1128 DVSS.n1115 4.5005
R24132 DVSS.n1128 DVSS.n1116 4.5005
R24133 DVSS.n1128 DVSS.n1114 4.5005
R24134 DVSS.n1128 DVSS.n1117 4.5005
R24135 DVSS.n1128 DVSS.n1113 4.5005
R24136 DVSS.n1128 DVSS.n1118 4.5005
R24137 DVSS.n1128 DVSS.n1112 4.5005
R24138 DVSS.n1128 DVSS.n1119 4.5005
R24139 DVSS.n1128 DVSS.n1111 4.5005
R24140 DVSS.n1128 DVSS.n1121 4.5005
R24141 DVSS.n1128 DVSS.n1110 4.5005
R24142 DVSS.n1128 DVSS.n1122 4.5005
R24143 DVSS.n1128 DVSS.n1124 4.5005
R24144 DVSS.n1128 DVSS.n1108 4.5005
R24145 DVSS.n22373 DVSS.n1128 4.5005
R24146 DVSS.n1151 DVSS.n1115 4.5005
R24147 DVSS.n1151 DVSS.n1116 4.5005
R24148 DVSS.n1151 DVSS.n1114 4.5005
R24149 DVSS.n1151 DVSS.n1117 4.5005
R24150 DVSS.n1151 DVSS.n1113 4.5005
R24151 DVSS.n1151 DVSS.n1118 4.5005
R24152 DVSS.n1151 DVSS.n1112 4.5005
R24153 DVSS.n1151 DVSS.n1119 4.5005
R24154 DVSS.n1151 DVSS.n1111 4.5005
R24155 DVSS.n1151 DVSS.n1121 4.5005
R24156 DVSS.n1151 DVSS.n1110 4.5005
R24157 DVSS.n1151 DVSS.n1122 4.5005
R24158 DVSS.n1164 DVSS.n1151 4.5005
R24159 DVSS.n1151 DVSS.n1124 4.5005
R24160 DVSS.n1151 DVSS.n1108 4.5005
R24161 DVSS.n22373 DVSS.n1151 4.5005
R24162 DVSS.n1127 DVSS.n1115 4.5005
R24163 DVSS.n1127 DVSS.n1116 4.5005
R24164 DVSS.n1127 DVSS.n1114 4.5005
R24165 DVSS.n1127 DVSS.n1117 4.5005
R24166 DVSS.n1127 DVSS.n1113 4.5005
R24167 DVSS.n1127 DVSS.n1118 4.5005
R24168 DVSS.n1127 DVSS.n1112 4.5005
R24169 DVSS.n1127 DVSS.n1119 4.5005
R24170 DVSS.n1127 DVSS.n1111 4.5005
R24171 DVSS.n1127 DVSS.n1121 4.5005
R24172 DVSS.n1127 DVSS.n1110 4.5005
R24173 DVSS.n1127 DVSS.n1122 4.5005
R24174 DVSS.n1127 DVSS.n1124 4.5005
R24175 DVSS.n1127 DVSS.n1108 4.5005
R24176 DVSS.n22373 DVSS.n1127 4.5005
R24177 DVSS.n1152 DVSS.n1115 4.5005
R24178 DVSS.n1152 DVSS.n1116 4.5005
R24179 DVSS.n1152 DVSS.n1114 4.5005
R24180 DVSS.n1152 DVSS.n1117 4.5005
R24181 DVSS.n1152 DVSS.n1113 4.5005
R24182 DVSS.n1152 DVSS.n1118 4.5005
R24183 DVSS.n1152 DVSS.n1112 4.5005
R24184 DVSS.n1152 DVSS.n1119 4.5005
R24185 DVSS.n1152 DVSS.n1111 4.5005
R24186 DVSS.n1152 DVSS.n1121 4.5005
R24187 DVSS.n1152 DVSS.n1110 4.5005
R24188 DVSS.n1152 DVSS.n1122 4.5005
R24189 DVSS.n1152 DVSS.n1124 4.5005
R24190 DVSS.n1152 DVSS.n1108 4.5005
R24191 DVSS.n22373 DVSS.n1152 4.5005
R24192 DVSS.n1126 DVSS.n1115 4.5005
R24193 DVSS.n1126 DVSS.n1116 4.5005
R24194 DVSS.n1126 DVSS.n1114 4.5005
R24195 DVSS.n1126 DVSS.n1117 4.5005
R24196 DVSS.n1126 DVSS.n1113 4.5005
R24197 DVSS.n1126 DVSS.n1118 4.5005
R24198 DVSS.n1126 DVSS.n1112 4.5005
R24199 DVSS.n1126 DVSS.n1119 4.5005
R24200 DVSS.n1126 DVSS.n1111 4.5005
R24201 DVSS.n1126 DVSS.n1121 4.5005
R24202 DVSS.n1126 DVSS.n1110 4.5005
R24203 DVSS.n1126 DVSS.n1122 4.5005
R24204 DVSS.n1126 DVSS.n1124 4.5005
R24205 DVSS.n1126 DVSS.n1108 4.5005
R24206 DVSS.n22373 DVSS.n1126 4.5005
R24207 DVSS.n1115 DVSS.n1107 4.5005
R24208 DVSS.n1116 DVSS.n1107 4.5005
R24209 DVSS.n1114 DVSS.n1107 4.5005
R24210 DVSS.n1117 DVSS.n1107 4.5005
R24211 DVSS.n1113 DVSS.n1107 4.5005
R24212 DVSS.n1118 DVSS.n1107 4.5005
R24213 DVSS.n1112 DVSS.n1107 4.5005
R24214 DVSS.n1119 DVSS.n1107 4.5005
R24215 DVSS.n1111 DVSS.n1107 4.5005
R24216 DVSS.n1121 DVSS.n1107 4.5005
R24217 DVSS.n1110 DVSS.n1107 4.5005
R24218 DVSS.n1122 DVSS.n1107 4.5005
R24219 DVSS.n1124 DVSS.n1107 4.5005
R24220 DVSS.n1108 DVSS.n1107 4.5005
R24221 DVSS.n22373 DVSS.n1107 4.5005
R24222 DVSS.n1125 DVSS.n1115 4.5005
R24223 DVSS.n1125 DVSS.n1116 4.5005
R24224 DVSS.n1125 DVSS.n1114 4.5005
R24225 DVSS.n1125 DVSS.n1117 4.5005
R24226 DVSS.n1125 DVSS.n1113 4.5005
R24227 DVSS.n1125 DVSS.n1118 4.5005
R24228 DVSS.n1125 DVSS.n1112 4.5005
R24229 DVSS.n1125 DVSS.n1119 4.5005
R24230 DVSS.n1125 DVSS.n1111 4.5005
R24231 DVSS.n1125 DVSS.n1121 4.5005
R24232 DVSS.n1125 DVSS.n1110 4.5005
R24233 DVSS.n1125 DVSS.n1122 4.5005
R24234 DVSS.n1125 DVSS.n1124 4.5005
R24235 DVSS.n1125 DVSS.n1108 4.5005
R24236 DVSS.n22373 DVSS.n1125 4.5005
R24237 DVSS.n22372 DVSS.n1115 4.5005
R24238 DVSS.n22372 DVSS.n1116 4.5005
R24239 DVSS.n22372 DVSS.n1114 4.5005
R24240 DVSS.n22372 DVSS.n1117 4.5005
R24241 DVSS.n22372 DVSS.n1113 4.5005
R24242 DVSS.n22372 DVSS.n1118 4.5005
R24243 DVSS.n22372 DVSS.n1112 4.5005
R24244 DVSS.n22372 DVSS.n1119 4.5005
R24245 DVSS.n22372 DVSS.n1111 4.5005
R24246 DVSS.n22372 DVSS.n1121 4.5005
R24247 DVSS.n22372 DVSS.n1110 4.5005
R24248 DVSS.n22372 DVSS.n1122 4.5005
R24249 DVSS.n22372 DVSS.n1164 4.5005
R24250 DVSS.n22372 DVSS.n1124 4.5005
R24251 DVSS.n22372 DVSS.n1108 4.5005
R24252 DVSS.n22373 DVSS.n22372 4.5005
R24253 DVSS.n13006 DVSS.n12979 4.5005
R24254 DVSS.n13006 DVSS.n12981 4.5005
R24255 DVSS.n13006 DVSS.n12978 4.5005
R24256 DVSS.n13006 DVSS.n12984 4.5005
R24257 DVSS.n13006 DVSS.n12976 4.5005
R24258 DVSS.n13006 DVSS.n12985 4.5005
R24259 DVSS.n13006 DVSS.n12975 4.5005
R24260 DVSS.n13006 DVSS.n12987 4.5005
R24261 DVSS.n13006 DVSS.n12974 4.5005
R24262 DVSS.n13006 DVSS.n12989 4.5005
R24263 DVSS.n13062 DVSS.n13006 4.5005
R24264 DVSS.n13008 DVSS.n12979 4.5005
R24265 DVSS.n13008 DVSS.n12981 4.5005
R24266 DVSS.n13008 DVSS.n12978 4.5005
R24267 DVSS.n13008 DVSS.n12982 4.5005
R24268 DVSS.n13008 DVSS.n12977 4.5005
R24269 DVSS.n13008 DVSS.n12984 4.5005
R24270 DVSS.n13008 DVSS.n12976 4.5005
R24271 DVSS.n13008 DVSS.n12985 4.5005
R24272 DVSS.n13008 DVSS.n12975 4.5005
R24273 DVSS.n13008 DVSS.n12987 4.5005
R24274 DVSS.n13008 DVSS.n12974 4.5005
R24275 DVSS.n13008 DVSS.n12988 4.5005
R24276 DVSS.n13008 DVSS.n12973 4.5005
R24277 DVSS.n13008 DVSS.n12989 4.5005
R24278 DVSS.n13062 DVSS.n13008 4.5005
R24279 DVSS.n13003 DVSS.n12979 4.5005
R24280 DVSS.n13003 DVSS.n12981 4.5005
R24281 DVSS.n13003 DVSS.n12978 4.5005
R24282 DVSS.n13003 DVSS.n12982 4.5005
R24283 DVSS.n13003 DVSS.n12977 4.5005
R24284 DVSS.n13003 DVSS.n12984 4.5005
R24285 DVSS.n13003 DVSS.n12976 4.5005
R24286 DVSS.n13003 DVSS.n12985 4.5005
R24287 DVSS.n13003 DVSS.n12975 4.5005
R24288 DVSS.n13003 DVSS.n12987 4.5005
R24289 DVSS.n13003 DVSS.n12974 4.5005
R24290 DVSS.n13003 DVSS.n12988 4.5005
R24291 DVSS.n13003 DVSS.n12989 4.5005
R24292 DVSS.n13062 DVSS.n13003 4.5005
R24293 DVSS.n13011 DVSS.n12979 4.5005
R24294 DVSS.n13011 DVSS.n12981 4.5005
R24295 DVSS.n13011 DVSS.n12978 4.5005
R24296 DVSS.n13011 DVSS.n12982 4.5005
R24297 DVSS.n13011 DVSS.n12977 4.5005
R24298 DVSS.n13011 DVSS.n12984 4.5005
R24299 DVSS.n13011 DVSS.n12976 4.5005
R24300 DVSS.n13011 DVSS.n12985 4.5005
R24301 DVSS.n13011 DVSS.n12975 4.5005
R24302 DVSS.n13011 DVSS.n12987 4.5005
R24303 DVSS.n13011 DVSS.n12974 4.5005
R24304 DVSS.n13011 DVSS.n12988 4.5005
R24305 DVSS.n13011 DVSS.n12989 4.5005
R24306 DVSS.n13062 DVSS.n13011 4.5005
R24307 DVSS.n13001 DVSS.n12979 4.5005
R24308 DVSS.n13001 DVSS.n12981 4.5005
R24309 DVSS.n13001 DVSS.n12978 4.5005
R24310 DVSS.n13001 DVSS.n12982 4.5005
R24311 DVSS.n13001 DVSS.n12977 4.5005
R24312 DVSS.n13001 DVSS.n12984 4.5005
R24313 DVSS.n13001 DVSS.n12976 4.5005
R24314 DVSS.n13001 DVSS.n12985 4.5005
R24315 DVSS.n13001 DVSS.n12975 4.5005
R24316 DVSS.n13001 DVSS.n12987 4.5005
R24317 DVSS.n13001 DVSS.n12974 4.5005
R24318 DVSS.n13001 DVSS.n12988 4.5005
R24319 DVSS.n13001 DVSS.n12989 4.5005
R24320 DVSS.n13001 DVSS.n12972 4.5005
R24321 DVSS.n13062 DVSS.n13001 4.5005
R24322 DVSS.n13013 DVSS.n12979 4.5005
R24323 DVSS.n13013 DVSS.n12981 4.5005
R24324 DVSS.n13013 DVSS.n12978 4.5005
R24325 DVSS.n13013 DVSS.n12982 4.5005
R24326 DVSS.n13013 DVSS.n12977 4.5005
R24327 DVSS.n13013 DVSS.n12984 4.5005
R24328 DVSS.n13013 DVSS.n12976 4.5005
R24329 DVSS.n13013 DVSS.n12985 4.5005
R24330 DVSS.n13013 DVSS.n12975 4.5005
R24331 DVSS.n13013 DVSS.n12987 4.5005
R24332 DVSS.n13013 DVSS.n12974 4.5005
R24333 DVSS.n13013 DVSS.n12988 4.5005
R24334 DVSS.n13013 DVSS.n12989 4.5005
R24335 DVSS.n13062 DVSS.n13013 4.5005
R24336 DVSS.n13000 DVSS.n12979 4.5005
R24337 DVSS.n13000 DVSS.n12981 4.5005
R24338 DVSS.n13000 DVSS.n12978 4.5005
R24339 DVSS.n13000 DVSS.n12982 4.5005
R24340 DVSS.n13000 DVSS.n12977 4.5005
R24341 DVSS.n13000 DVSS.n12984 4.5005
R24342 DVSS.n13000 DVSS.n12976 4.5005
R24343 DVSS.n13000 DVSS.n12985 4.5005
R24344 DVSS.n13000 DVSS.n12975 4.5005
R24345 DVSS.n13000 DVSS.n12987 4.5005
R24346 DVSS.n13000 DVSS.n12974 4.5005
R24347 DVSS.n13000 DVSS.n12988 4.5005
R24348 DVSS.n13000 DVSS.n12989 4.5005
R24349 DVSS.n13062 DVSS.n13000 4.5005
R24350 DVSS.n13022 DVSS.n12979 4.5005
R24351 DVSS.n13022 DVSS.n12981 4.5005
R24352 DVSS.n13022 DVSS.n12978 4.5005
R24353 DVSS.n13022 DVSS.n12982 4.5005
R24354 DVSS.n13022 DVSS.n12977 4.5005
R24355 DVSS.n13022 DVSS.n12984 4.5005
R24356 DVSS.n13022 DVSS.n12976 4.5005
R24357 DVSS.n13022 DVSS.n12985 4.5005
R24358 DVSS.n13022 DVSS.n12975 4.5005
R24359 DVSS.n13022 DVSS.n12987 4.5005
R24360 DVSS.n13022 DVSS.n12974 4.5005
R24361 DVSS.n13022 DVSS.n12988 4.5005
R24362 DVSS.n13022 DVSS.n12989 4.5005
R24363 DVSS.n13022 DVSS.n12972 4.5005
R24364 DVSS.n13062 DVSS.n13022 4.5005
R24365 DVSS.n12999 DVSS.n12979 4.5005
R24366 DVSS.n12999 DVSS.n12981 4.5005
R24367 DVSS.n12999 DVSS.n12978 4.5005
R24368 DVSS.n12999 DVSS.n12982 4.5005
R24369 DVSS.n12999 DVSS.n12977 4.5005
R24370 DVSS.n12999 DVSS.n12984 4.5005
R24371 DVSS.n12999 DVSS.n12976 4.5005
R24372 DVSS.n12999 DVSS.n12985 4.5005
R24373 DVSS.n12999 DVSS.n12975 4.5005
R24374 DVSS.n12999 DVSS.n12987 4.5005
R24375 DVSS.n12999 DVSS.n12974 4.5005
R24376 DVSS.n12999 DVSS.n12988 4.5005
R24377 DVSS.n12999 DVSS.n12989 4.5005
R24378 DVSS.n13062 DVSS.n12999 4.5005
R24379 DVSS.n13025 DVSS.n12979 4.5005
R24380 DVSS.n13025 DVSS.n12981 4.5005
R24381 DVSS.n13025 DVSS.n12978 4.5005
R24382 DVSS.n13025 DVSS.n12982 4.5005
R24383 DVSS.n13025 DVSS.n12977 4.5005
R24384 DVSS.n13025 DVSS.n12984 4.5005
R24385 DVSS.n13025 DVSS.n12976 4.5005
R24386 DVSS.n13025 DVSS.n12985 4.5005
R24387 DVSS.n13025 DVSS.n12975 4.5005
R24388 DVSS.n13025 DVSS.n12987 4.5005
R24389 DVSS.n13025 DVSS.n12974 4.5005
R24390 DVSS.n13025 DVSS.n12988 4.5005
R24391 DVSS.n13025 DVSS.n12989 4.5005
R24392 DVSS.n13062 DVSS.n13025 4.5005
R24393 DVSS.n12997 DVSS.n12979 4.5005
R24394 DVSS.n12997 DVSS.n12981 4.5005
R24395 DVSS.n12997 DVSS.n12978 4.5005
R24396 DVSS.n12997 DVSS.n12982 4.5005
R24397 DVSS.n12997 DVSS.n12977 4.5005
R24398 DVSS.n12997 DVSS.n12984 4.5005
R24399 DVSS.n12997 DVSS.n12976 4.5005
R24400 DVSS.n12997 DVSS.n12985 4.5005
R24401 DVSS.n12997 DVSS.n12975 4.5005
R24402 DVSS.n12997 DVSS.n12987 4.5005
R24403 DVSS.n12997 DVSS.n12974 4.5005
R24404 DVSS.n12997 DVSS.n12988 4.5005
R24405 DVSS.n12997 DVSS.n12989 4.5005
R24406 DVSS.n12997 DVSS.n12972 4.5005
R24407 DVSS.n13062 DVSS.n12997 4.5005
R24408 DVSS.n13027 DVSS.n12979 4.5005
R24409 DVSS.n13027 DVSS.n12981 4.5005
R24410 DVSS.n13027 DVSS.n12978 4.5005
R24411 DVSS.n13027 DVSS.n12982 4.5005
R24412 DVSS.n13027 DVSS.n12977 4.5005
R24413 DVSS.n13027 DVSS.n12984 4.5005
R24414 DVSS.n13027 DVSS.n12976 4.5005
R24415 DVSS.n13027 DVSS.n12985 4.5005
R24416 DVSS.n13027 DVSS.n12975 4.5005
R24417 DVSS.n13027 DVSS.n12987 4.5005
R24418 DVSS.n13027 DVSS.n12974 4.5005
R24419 DVSS.n13027 DVSS.n12988 4.5005
R24420 DVSS.n13027 DVSS.n12989 4.5005
R24421 DVSS.n13062 DVSS.n13027 4.5005
R24422 DVSS.n12996 DVSS.n12979 4.5005
R24423 DVSS.n12996 DVSS.n12981 4.5005
R24424 DVSS.n12996 DVSS.n12978 4.5005
R24425 DVSS.n12996 DVSS.n12982 4.5005
R24426 DVSS.n12996 DVSS.n12977 4.5005
R24427 DVSS.n12996 DVSS.n12984 4.5005
R24428 DVSS.n12996 DVSS.n12976 4.5005
R24429 DVSS.n12996 DVSS.n12985 4.5005
R24430 DVSS.n12996 DVSS.n12975 4.5005
R24431 DVSS.n12996 DVSS.n12987 4.5005
R24432 DVSS.n12996 DVSS.n12974 4.5005
R24433 DVSS.n12996 DVSS.n12988 4.5005
R24434 DVSS.n12996 DVSS.n12989 4.5005
R24435 DVSS.n13062 DVSS.n12996 4.5005
R24436 DVSS.n13036 DVSS.n12979 4.5005
R24437 DVSS.n13036 DVSS.n12981 4.5005
R24438 DVSS.n13036 DVSS.n12978 4.5005
R24439 DVSS.n13036 DVSS.n12982 4.5005
R24440 DVSS.n13036 DVSS.n12977 4.5005
R24441 DVSS.n13036 DVSS.n12984 4.5005
R24442 DVSS.n13036 DVSS.n12976 4.5005
R24443 DVSS.n13036 DVSS.n12985 4.5005
R24444 DVSS.n13036 DVSS.n12975 4.5005
R24445 DVSS.n13036 DVSS.n12987 4.5005
R24446 DVSS.n13036 DVSS.n12974 4.5005
R24447 DVSS.n13036 DVSS.n12988 4.5005
R24448 DVSS.n13036 DVSS.n12989 4.5005
R24449 DVSS.n13036 DVSS.n12972 4.5005
R24450 DVSS.n13062 DVSS.n13036 4.5005
R24451 DVSS.n12995 DVSS.n12979 4.5005
R24452 DVSS.n12995 DVSS.n12981 4.5005
R24453 DVSS.n12995 DVSS.n12978 4.5005
R24454 DVSS.n12995 DVSS.n12982 4.5005
R24455 DVSS.n12995 DVSS.n12977 4.5005
R24456 DVSS.n12995 DVSS.n12984 4.5005
R24457 DVSS.n12995 DVSS.n12976 4.5005
R24458 DVSS.n12995 DVSS.n12985 4.5005
R24459 DVSS.n12995 DVSS.n12975 4.5005
R24460 DVSS.n12995 DVSS.n12987 4.5005
R24461 DVSS.n12995 DVSS.n12974 4.5005
R24462 DVSS.n12995 DVSS.n12988 4.5005
R24463 DVSS.n12995 DVSS.n12989 4.5005
R24464 DVSS.n13062 DVSS.n12995 4.5005
R24465 DVSS.n13039 DVSS.n12979 4.5005
R24466 DVSS.n13039 DVSS.n12981 4.5005
R24467 DVSS.n13039 DVSS.n12978 4.5005
R24468 DVSS.n13039 DVSS.n12982 4.5005
R24469 DVSS.n13039 DVSS.n12977 4.5005
R24470 DVSS.n13039 DVSS.n12984 4.5005
R24471 DVSS.n13039 DVSS.n12976 4.5005
R24472 DVSS.n13039 DVSS.n12985 4.5005
R24473 DVSS.n13039 DVSS.n12975 4.5005
R24474 DVSS.n13039 DVSS.n12987 4.5005
R24475 DVSS.n13039 DVSS.n12974 4.5005
R24476 DVSS.n13039 DVSS.n12988 4.5005
R24477 DVSS.n13039 DVSS.n12989 4.5005
R24478 DVSS.n13062 DVSS.n13039 4.5005
R24479 DVSS.n12993 DVSS.n12979 4.5005
R24480 DVSS.n12993 DVSS.n12981 4.5005
R24481 DVSS.n12993 DVSS.n12978 4.5005
R24482 DVSS.n12993 DVSS.n12982 4.5005
R24483 DVSS.n12993 DVSS.n12977 4.5005
R24484 DVSS.n12993 DVSS.n12984 4.5005
R24485 DVSS.n12993 DVSS.n12976 4.5005
R24486 DVSS.n12993 DVSS.n12985 4.5005
R24487 DVSS.n12993 DVSS.n12975 4.5005
R24488 DVSS.n12993 DVSS.n12987 4.5005
R24489 DVSS.n12993 DVSS.n12974 4.5005
R24490 DVSS.n12993 DVSS.n12988 4.5005
R24491 DVSS.n12993 DVSS.n12989 4.5005
R24492 DVSS.n12993 DVSS.n12972 4.5005
R24493 DVSS.n13062 DVSS.n12993 4.5005
R24494 DVSS.n13047 DVSS.n12979 4.5005
R24495 DVSS.n13047 DVSS.n12981 4.5005
R24496 DVSS.n13047 DVSS.n12978 4.5005
R24497 DVSS.n13047 DVSS.n12982 4.5005
R24498 DVSS.n13047 DVSS.n12977 4.5005
R24499 DVSS.n13047 DVSS.n12984 4.5005
R24500 DVSS.n13047 DVSS.n12976 4.5005
R24501 DVSS.n13047 DVSS.n12985 4.5005
R24502 DVSS.n13047 DVSS.n12975 4.5005
R24503 DVSS.n13047 DVSS.n12987 4.5005
R24504 DVSS.n13047 DVSS.n12974 4.5005
R24505 DVSS.n13047 DVSS.n12988 4.5005
R24506 DVSS.n13047 DVSS.n12973 4.5005
R24507 DVSS.n13047 DVSS.n12989 4.5005
R24508 DVSS.n13047 DVSS.n12972 4.5005
R24509 DVSS.n13062 DVSS.n13047 4.5005
R24510 DVSS.n12992 DVSS.n12979 4.5005
R24511 DVSS.n12992 DVSS.n12981 4.5005
R24512 DVSS.n12992 DVSS.n12978 4.5005
R24513 DVSS.n12992 DVSS.n12982 4.5005
R24514 DVSS.n12992 DVSS.n12977 4.5005
R24515 DVSS.n12992 DVSS.n12984 4.5005
R24516 DVSS.n12992 DVSS.n12976 4.5005
R24517 DVSS.n12992 DVSS.n12985 4.5005
R24518 DVSS.n12992 DVSS.n12975 4.5005
R24519 DVSS.n12992 DVSS.n12987 4.5005
R24520 DVSS.n12992 DVSS.n12974 4.5005
R24521 DVSS.n12992 DVSS.n12988 4.5005
R24522 DVSS.n12992 DVSS.n12989 4.5005
R24523 DVSS.n12992 DVSS.n12972 4.5005
R24524 DVSS.n13062 DVSS.n12992 4.5005
R24525 DVSS.n13056 DVSS.n12979 4.5005
R24526 DVSS.n13056 DVSS.n12981 4.5005
R24527 DVSS.n13056 DVSS.n12978 4.5005
R24528 DVSS.n13056 DVSS.n12982 4.5005
R24529 DVSS.n13056 DVSS.n12977 4.5005
R24530 DVSS.n13056 DVSS.n12984 4.5005
R24531 DVSS.n13056 DVSS.n12976 4.5005
R24532 DVSS.n13056 DVSS.n12985 4.5005
R24533 DVSS.n13056 DVSS.n12975 4.5005
R24534 DVSS.n13056 DVSS.n12987 4.5005
R24535 DVSS.n13056 DVSS.n12974 4.5005
R24536 DVSS.n13056 DVSS.n12988 4.5005
R24537 DVSS.n13056 DVSS.n12989 4.5005
R24538 DVSS.n13056 DVSS.n12972 4.5005
R24539 DVSS.n13062 DVSS.n13056 4.5005
R24540 DVSS.n12991 DVSS.n12979 4.5005
R24541 DVSS.n12991 DVSS.n12981 4.5005
R24542 DVSS.n12991 DVSS.n12978 4.5005
R24543 DVSS.n12991 DVSS.n12982 4.5005
R24544 DVSS.n12991 DVSS.n12977 4.5005
R24545 DVSS.n12991 DVSS.n12984 4.5005
R24546 DVSS.n12991 DVSS.n12976 4.5005
R24547 DVSS.n12991 DVSS.n12985 4.5005
R24548 DVSS.n12991 DVSS.n12975 4.5005
R24549 DVSS.n12991 DVSS.n12987 4.5005
R24550 DVSS.n12991 DVSS.n12974 4.5005
R24551 DVSS.n12991 DVSS.n12988 4.5005
R24552 DVSS.n12991 DVSS.n12989 4.5005
R24553 DVSS.n12991 DVSS.n12972 4.5005
R24554 DVSS.n13062 DVSS.n12991 4.5005
R24555 DVSS.n13061 DVSS.n12979 4.5005
R24556 DVSS.n13061 DVSS.n12981 4.5005
R24557 DVSS.n13061 DVSS.n12978 4.5005
R24558 DVSS.n13061 DVSS.n12982 4.5005
R24559 DVSS.n13061 DVSS.n12977 4.5005
R24560 DVSS.n13061 DVSS.n12984 4.5005
R24561 DVSS.n13061 DVSS.n12976 4.5005
R24562 DVSS.n13061 DVSS.n12985 4.5005
R24563 DVSS.n13061 DVSS.n12975 4.5005
R24564 DVSS.n13061 DVSS.n12987 4.5005
R24565 DVSS.n13061 DVSS.n12974 4.5005
R24566 DVSS.n13061 DVSS.n12988 4.5005
R24567 DVSS.n13061 DVSS.n12989 4.5005
R24568 DVSS.n13061 DVSS.n12972 4.5005
R24569 DVSS.n13062 DVSS.n13061 4.5005
R24570 DVSS.n12979 DVSS.n12962 4.5005
R24571 DVSS.n12981 DVSS.n12962 4.5005
R24572 DVSS.n12978 DVSS.n12962 4.5005
R24573 DVSS.n12982 DVSS.n12962 4.5005
R24574 DVSS.n12977 DVSS.n12962 4.5005
R24575 DVSS.n12984 DVSS.n12962 4.5005
R24576 DVSS.n12976 DVSS.n12962 4.5005
R24577 DVSS.n12985 DVSS.n12962 4.5005
R24578 DVSS.n12975 DVSS.n12962 4.5005
R24579 DVSS.n12987 DVSS.n12962 4.5005
R24580 DVSS.n12974 DVSS.n12962 4.5005
R24581 DVSS.n12988 DVSS.n12962 4.5005
R24582 DVSS.n12989 DVSS.n12962 4.5005
R24583 DVSS.n12972 DVSS.n12962 4.5005
R24584 DVSS.n13062 DVSS.n12962 4.5005
R24585 DVSS.n13063 DVSS.n12979 4.5005
R24586 DVSS.n13063 DVSS.n12981 4.5005
R24587 DVSS.n13063 DVSS.n12978 4.5005
R24588 DVSS.n13063 DVSS.n12982 4.5005
R24589 DVSS.n13063 DVSS.n12977 4.5005
R24590 DVSS.n13063 DVSS.n12984 4.5005
R24591 DVSS.n13063 DVSS.n12976 4.5005
R24592 DVSS.n13063 DVSS.n12985 4.5005
R24593 DVSS.n13063 DVSS.n12975 4.5005
R24594 DVSS.n13063 DVSS.n12987 4.5005
R24595 DVSS.n13063 DVSS.n12974 4.5005
R24596 DVSS.n13063 DVSS.n12988 4.5005
R24597 DVSS.n13063 DVSS.n12973 4.5005
R24598 DVSS.n13063 DVSS.n12989 4.5005
R24599 DVSS.n13063 DVSS.n12972 4.5005
R24600 DVSS.n13063 DVSS.n13062 4.5005
R24601 DVSS.n383 DVSS.n349 4.5005
R24602 DVSS.n387 DVSS.n349 4.5005
R24603 DVSS.n380 DVSS.n349 4.5005
R24604 DVSS.n389 DVSS.n349 4.5005
R24605 DVSS.n379 DVSS.n349 4.5005
R24606 DVSS.n390 DVSS.n349 4.5005
R24607 DVSS.n378 DVSS.n349 4.5005
R24608 DVSS.n394 DVSS.n349 4.5005
R24609 DVSS.n349 DVSS.n334 4.5005
R24610 DVSS.n23004 DVSS.n349 4.5005
R24611 DVSS.n23002 DVSS.n349 4.5005
R24612 DVSS.n383 DVSS.n351 4.5005
R24613 DVSS.n386 DVSS.n351 4.5005
R24614 DVSS.n381 DVSS.n351 4.5005
R24615 DVSS.n387 DVSS.n351 4.5005
R24616 DVSS.n380 DVSS.n351 4.5005
R24617 DVSS.n389 DVSS.n351 4.5005
R24618 DVSS.n379 DVSS.n351 4.5005
R24619 DVSS.n390 DVSS.n351 4.5005
R24620 DVSS.n378 DVSS.n351 4.5005
R24621 DVSS.n393 DVSS.n351 4.5005
R24622 DVSS.n377 DVSS.n351 4.5005
R24623 DVSS.n394 DVSS.n351 4.5005
R24624 DVSS.n351 DVSS.n334 4.5005
R24625 DVSS.n23004 DVSS.n351 4.5005
R24626 DVSS.n23002 DVSS.n351 4.5005
R24627 DVSS.n383 DVSS.n348 4.5005
R24628 DVSS.n386 DVSS.n348 4.5005
R24629 DVSS.n381 DVSS.n348 4.5005
R24630 DVSS.n387 DVSS.n348 4.5005
R24631 DVSS.n380 DVSS.n348 4.5005
R24632 DVSS.n389 DVSS.n348 4.5005
R24633 DVSS.n379 DVSS.n348 4.5005
R24634 DVSS.n390 DVSS.n348 4.5005
R24635 DVSS.n378 DVSS.n348 4.5005
R24636 DVSS.n393 DVSS.n348 4.5005
R24637 DVSS.n377 DVSS.n348 4.5005
R24638 DVSS.n394 DVSS.n348 4.5005
R24639 DVSS.n23004 DVSS.n348 4.5005
R24640 DVSS.n23002 DVSS.n348 4.5005
R24641 DVSS.n383 DVSS.n353 4.5005
R24642 DVSS.n386 DVSS.n353 4.5005
R24643 DVSS.n381 DVSS.n353 4.5005
R24644 DVSS.n387 DVSS.n353 4.5005
R24645 DVSS.n380 DVSS.n353 4.5005
R24646 DVSS.n389 DVSS.n353 4.5005
R24647 DVSS.n379 DVSS.n353 4.5005
R24648 DVSS.n390 DVSS.n353 4.5005
R24649 DVSS.n378 DVSS.n353 4.5005
R24650 DVSS.n393 DVSS.n353 4.5005
R24651 DVSS.n377 DVSS.n353 4.5005
R24652 DVSS.n394 DVSS.n353 4.5005
R24653 DVSS.n23004 DVSS.n353 4.5005
R24654 DVSS.n23002 DVSS.n353 4.5005
R24655 DVSS.n383 DVSS.n346 4.5005
R24656 DVSS.n386 DVSS.n346 4.5005
R24657 DVSS.n381 DVSS.n346 4.5005
R24658 DVSS.n387 DVSS.n346 4.5005
R24659 DVSS.n380 DVSS.n346 4.5005
R24660 DVSS.n389 DVSS.n346 4.5005
R24661 DVSS.n379 DVSS.n346 4.5005
R24662 DVSS.n390 DVSS.n346 4.5005
R24663 DVSS.n378 DVSS.n346 4.5005
R24664 DVSS.n393 DVSS.n346 4.5005
R24665 DVSS.n377 DVSS.n346 4.5005
R24666 DVSS.n394 DVSS.n346 4.5005
R24667 DVSS.n23004 DVSS.n346 4.5005
R24668 DVSS.n376 DVSS.n346 4.5005
R24669 DVSS.n23002 DVSS.n346 4.5005
R24670 DVSS.n383 DVSS.n354 4.5005
R24671 DVSS.n386 DVSS.n354 4.5005
R24672 DVSS.n381 DVSS.n354 4.5005
R24673 DVSS.n387 DVSS.n354 4.5005
R24674 DVSS.n380 DVSS.n354 4.5005
R24675 DVSS.n389 DVSS.n354 4.5005
R24676 DVSS.n379 DVSS.n354 4.5005
R24677 DVSS.n390 DVSS.n354 4.5005
R24678 DVSS.n378 DVSS.n354 4.5005
R24679 DVSS.n393 DVSS.n354 4.5005
R24680 DVSS.n377 DVSS.n354 4.5005
R24681 DVSS.n394 DVSS.n354 4.5005
R24682 DVSS.n23004 DVSS.n354 4.5005
R24683 DVSS.n23002 DVSS.n354 4.5005
R24684 DVSS.n383 DVSS.n345 4.5005
R24685 DVSS.n386 DVSS.n345 4.5005
R24686 DVSS.n381 DVSS.n345 4.5005
R24687 DVSS.n387 DVSS.n345 4.5005
R24688 DVSS.n380 DVSS.n345 4.5005
R24689 DVSS.n389 DVSS.n345 4.5005
R24690 DVSS.n379 DVSS.n345 4.5005
R24691 DVSS.n390 DVSS.n345 4.5005
R24692 DVSS.n378 DVSS.n345 4.5005
R24693 DVSS.n393 DVSS.n345 4.5005
R24694 DVSS.n377 DVSS.n345 4.5005
R24695 DVSS.n394 DVSS.n345 4.5005
R24696 DVSS.n23004 DVSS.n345 4.5005
R24697 DVSS.n23002 DVSS.n345 4.5005
R24698 DVSS.n383 DVSS.n356 4.5005
R24699 DVSS.n386 DVSS.n356 4.5005
R24700 DVSS.n381 DVSS.n356 4.5005
R24701 DVSS.n387 DVSS.n356 4.5005
R24702 DVSS.n380 DVSS.n356 4.5005
R24703 DVSS.n389 DVSS.n356 4.5005
R24704 DVSS.n379 DVSS.n356 4.5005
R24705 DVSS.n390 DVSS.n356 4.5005
R24706 DVSS.n378 DVSS.n356 4.5005
R24707 DVSS.n393 DVSS.n356 4.5005
R24708 DVSS.n377 DVSS.n356 4.5005
R24709 DVSS.n394 DVSS.n356 4.5005
R24710 DVSS.n23004 DVSS.n356 4.5005
R24711 DVSS.n376 DVSS.n356 4.5005
R24712 DVSS.n23002 DVSS.n356 4.5005
R24713 DVSS.n383 DVSS.n344 4.5005
R24714 DVSS.n386 DVSS.n344 4.5005
R24715 DVSS.n381 DVSS.n344 4.5005
R24716 DVSS.n387 DVSS.n344 4.5005
R24717 DVSS.n380 DVSS.n344 4.5005
R24718 DVSS.n389 DVSS.n344 4.5005
R24719 DVSS.n379 DVSS.n344 4.5005
R24720 DVSS.n390 DVSS.n344 4.5005
R24721 DVSS.n378 DVSS.n344 4.5005
R24722 DVSS.n393 DVSS.n344 4.5005
R24723 DVSS.n377 DVSS.n344 4.5005
R24724 DVSS.n394 DVSS.n344 4.5005
R24725 DVSS.n23004 DVSS.n344 4.5005
R24726 DVSS.n23002 DVSS.n344 4.5005
R24727 DVSS.n383 DVSS.n358 4.5005
R24728 DVSS.n386 DVSS.n358 4.5005
R24729 DVSS.n381 DVSS.n358 4.5005
R24730 DVSS.n387 DVSS.n358 4.5005
R24731 DVSS.n380 DVSS.n358 4.5005
R24732 DVSS.n389 DVSS.n358 4.5005
R24733 DVSS.n379 DVSS.n358 4.5005
R24734 DVSS.n390 DVSS.n358 4.5005
R24735 DVSS.n378 DVSS.n358 4.5005
R24736 DVSS.n393 DVSS.n358 4.5005
R24737 DVSS.n377 DVSS.n358 4.5005
R24738 DVSS.n394 DVSS.n358 4.5005
R24739 DVSS.n23004 DVSS.n358 4.5005
R24740 DVSS.n23002 DVSS.n358 4.5005
R24741 DVSS.n383 DVSS.n342 4.5005
R24742 DVSS.n386 DVSS.n342 4.5005
R24743 DVSS.n381 DVSS.n342 4.5005
R24744 DVSS.n387 DVSS.n342 4.5005
R24745 DVSS.n380 DVSS.n342 4.5005
R24746 DVSS.n389 DVSS.n342 4.5005
R24747 DVSS.n379 DVSS.n342 4.5005
R24748 DVSS.n390 DVSS.n342 4.5005
R24749 DVSS.n378 DVSS.n342 4.5005
R24750 DVSS.n393 DVSS.n342 4.5005
R24751 DVSS.n377 DVSS.n342 4.5005
R24752 DVSS.n394 DVSS.n342 4.5005
R24753 DVSS.n23004 DVSS.n342 4.5005
R24754 DVSS.n376 DVSS.n342 4.5005
R24755 DVSS.n23002 DVSS.n342 4.5005
R24756 DVSS.n383 DVSS.n359 4.5005
R24757 DVSS.n386 DVSS.n359 4.5005
R24758 DVSS.n381 DVSS.n359 4.5005
R24759 DVSS.n387 DVSS.n359 4.5005
R24760 DVSS.n380 DVSS.n359 4.5005
R24761 DVSS.n389 DVSS.n359 4.5005
R24762 DVSS.n379 DVSS.n359 4.5005
R24763 DVSS.n390 DVSS.n359 4.5005
R24764 DVSS.n378 DVSS.n359 4.5005
R24765 DVSS.n393 DVSS.n359 4.5005
R24766 DVSS.n377 DVSS.n359 4.5005
R24767 DVSS.n394 DVSS.n359 4.5005
R24768 DVSS.n23004 DVSS.n359 4.5005
R24769 DVSS.n23002 DVSS.n359 4.5005
R24770 DVSS.n383 DVSS.n341 4.5005
R24771 DVSS.n386 DVSS.n341 4.5005
R24772 DVSS.n381 DVSS.n341 4.5005
R24773 DVSS.n387 DVSS.n341 4.5005
R24774 DVSS.n380 DVSS.n341 4.5005
R24775 DVSS.n389 DVSS.n341 4.5005
R24776 DVSS.n379 DVSS.n341 4.5005
R24777 DVSS.n390 DVSS.n341 4.5005
R24778 DVSS.n378 DVSS.n341 4.5005
R24779 DVSS.n393 DVSS.n341 4.5005
R24780 DVSS.n377 DVSS.n341 4.5005
R24781 DVSS.n394 DVSS.n341 4.5005
R24782 DVSS.n23004 DVSS.n341 4.5005
R24783 DVSS.n23002 DVSS.n341 4.5005
R24784 DVSS.n383 DVSS.n361 4.5005
R24785 DVSS.n386 DVSS.n361 4.5005
R24786 DVSS.n381 DVSS.n361 4.5005
R24787 DVSS.n387 DVSS.n361 4.5005
R24788 DVSS.n380 DVSS.n361 4.5005
R24789 DVSS.n389 DVSS.n361 4.5005
R24790 DVSS.n379 DVSS.n361 4.5005
R24791 DVSS.n390 DVSS.n361 4.5005
R24792 DVSS.n378 DVSS.n361 4.5005
R24793 DVSS.n393 DVSS.n361 4.5005
R24794 DVSS.n377 DVSS.n361 4.5005
R24795 DVSS.n394 DVSS.n361 4.5005
R24796 DVSS.n23004 DVSS.n361 4.5005
R24797 DVSS.n376 DVSS.n361 4.5005
R24798 DVSS.n23002 DVSS.n361 4.5005
R24799 DVSS.n383 DVSS.n340 4.5005
R24800 DVSS.n386 DVSS.n340 4.5005
R24801 DVSS.n381 DVSS.n340 4.5005
R24802 DVSS.n387 DVSS.n340 4.5005
R24803 DVSS.n380 DVSS.n340 4.5005
R24804 DVSS.n389 DVSS.n340 4.5005
R24805 DVSS.n379 DVSS.n340 4.5005
R24806 DVSS.n390 DVSS.n340 4.5005
R24807 DVSS.n378 DVSS.n340 4.5005
R24808 DVSS.n393 DVSS.n340 4.5005
R24809 DVSS.n377 DVSS.n340 4.5005
R24810 DVSS.n394 DVSS.n340 4.5005
R24811 DVSS.n23004 DVSS.n340 4.5005
R24812 DVSS.n23002 DVSS.n340 4.5005
R24813 DVSS.n383 DVSS.n363 4.5005
R24814 DVSS.n386 DVSS.n363 4.5005
R24815 DVSS.n381 DVSS.n363 4.5005
R24816 DVSS.n387 DVSS.n363 4.5005
R24817 DVSS.n380 DVSS.n363 4.5005
R24818 DVSS.n389 DVSS.n363 4.5005
R24819 DVSS.n379 DVSS.n363 4.5005
R24820 DVSS.n390 DVSS.n363 4.5005
R24821 DVSS.n378 DVSS.n363 4.5005
R24822 DVSS.n393 DVSS.n363 4.5005
R24823 DVSS.n377 DVSS.n363 4.5005
R24824 DVSS.n394 DVSS.n363 4.5005
R24825 DVSS.n23004 DVSS.n363 4.5005
R24826 DVSS.n23002 DVSS.n363 4.5005
R24827 DVSS.n383 DVSS.n338 4.5005
R24828 DVSS.n386 DVSS.n338 4.5005
R24829 DVSS.n381 DVSS.n338 4.5005
R24830 DVSS.n387 DVSS.n338 4.5005
R24831 DVSS.n380 DVSS.n338 4.5005
R24832 DVSS.n389 DVSS.n338 4.5005
R24833 DVSS.n379 DVSS.n338 4.5005
R24834 DVSS.n390 DVSS.n338 4.5005
R24835 DVSS.n378 DVSS.n338 4.5005
R24836 DVSS.n393 DVSS.n338 4.5005
R24837 DVSS.n377 DVSS.n338 4.5005
R24838 DVSS.n394 DVSS.n338 4.5005
R24839 DVSS.n23004 DVSS.n338 4.5005
R24840 DVSS.n376 DVSS.n338 4.5005
R24841 DVSS.n23002 DVSS.n338 4.5005
R24842 DVSS.n383 DVSS.n364 4.5005
R24843 DVSS.n386 DVSS.n364 4.5005
R24844 DVSS.n381 DVSS.n364 4.5005
R24845 DVSS.n387 DVSS.n364 4.5005
R24846 DVSS.n380 DVSS.n364 4.5005
R24847 DVSS.n389 DVSS.n364 4.5005
R24848 DVSS.n379 DVSS.n364 4.5005
R24849 DVSS.n390 DVSS.n364 4.5005
R24850 DVSS.n378 DVSS.n364 4.5005
R24851 DVSS.n393 DVSS.n364 4.5005
R24852 DVSS.n377 DVSS.n364 4.5005
R24853 DVSS.n394 DVSS.n364 4.5005
R24854 DVSS.n364 DVSS.n334 4.5005
R24855 DVSS.n23004 DVSS.n364 4.5005
R24856 DVSS.n376 DVSS.n364 4.5005
R24857 DVSS.n23002 DVSS.n364 4.5005
R24858 DVSS.n383 DVSS.n337 4.5005
R24859 DVSS.n386 DVSS.n337 4.5005
R24860 DVSS.n381 DVSS.n337 4.5005
R24861 DVSS.n387 DVSS.n337 4.5005
R24862 DVSS.n380 DVSS.n337 4.5005
R24863 DVSS.n389 DVSS.n337 4.5005
R24864 DVSS.n379 DVSS.n337 4.5005
R24865 DVSS.n390 DVSS.n337 4.5005
R24866 DVSS.n378 DVSS.n337 4.5005
R24867 DVSS.n393 DVSS.n337 4.5005
R24868 DVSS.n377 DVSS.n337 4.5005
R24869 DVSS.n394 DVSS.n337 4.5005
R24870 DVSS.n23004 DVSS.n337 4.5005
R24871 DVSS.n376 DVSS.n337 4.5005
R24872 DVSS.n23002 DVSS.n337 4.5005
R24873 DVSS.n383 DVSS.n366 4.5005
R24874 DVSS.n386 DVSS.n366 4.5005
R24875 DVSS.n381 DVSS.n366 4.5005
R24876 DVSS.n387 DVSS.n366 4.5005
R24877 DVSS.n380 DVSS.n366 4.5005
R24878 DVSS.n389 DVSS.n366 4.5005
R24879 DVSS.n379 DVSS.n366 4.5005
R24880 DVSS.n390 DVSS.n366 4.5005
R24881 DVSS.n378 DVSS.n366 4.5005
R24882 DVSS.n393 DVSS.n366 4.5005
R24883 DVSS.n377 DVSS.n366 4.5005
R24884 DVSS.n394 DVSS.n366 4.5005
R24885 DVSS.n23004 DVSS.n366 4.5005
R24886 DVSS.n376 DVSS.n366 4.5005
R24887 DVSS.n23002 DVSS.n366 4.5005
R24888 DVSS.n383 DVSS.n336 4.5005
R24889 DVSS.n386 DVSS.n336 4.5005
R24890 DVSS.n381 DVSS.n336 4.5005
R24891 DVSS.n387 DVSS.n336 4.5005
R24892 DVSS.n380 DVSS.n336 4.5005
R24893 DVSS.n389 DVSS.n336 4.5005
R24894 DVSS.n379 DVSS.n336 4.5005
R24895 DVSS.n390 DVSS.n336 4.5005
R24896 DVSS.n378 DVSS.n336 4.5005
R24897 DVSS.n393 DVSS.n336 4.5005
R24898 DVSS.n377 DVSS.n336 4.5005
R24899 DVSS.n394 DVSS.n336 4.5005
R24900 DVSS.n23004 DVSS.n336 4.5005
R24901 DVSS.n376 DVSS.n336 4.5005
R24902 DVSS.n23002 DVSS.n336 4.5005
R24903 DVSS.n383 DVSS.n368 4.5005
R24904 DVSS.n386 DVSS.n368 4.5005
R24905 DVSS.n381 DVSS.n368 4.5005
R24906 DVSS.n387 DVSS.n368 4.5005
R24907 DVSS.n380 DVSS.n368 4.5005
R24908 DVSS.n389 DVSS.n368 4.5005
R24909 DVSS.n379 DVSS.n368 4.5005
R24910 DVSS.n390 DVSS.n368 4.5005
R24911 DVSS.n378 DVSS.n368 4.5005
R24912 DVSS.n393 DVSS.n368 4.5005
R24913 DVSS.n377 DVSS.n368 4.5005
R24914 DVSS.n394 DVSS.n368 4.5005
R24915 DVSS.n23004 DVSS.n368 4.5005
R24916 DVSS.n376 DVSS.n368 4.5005
R24917 DVSS.n23002 DVSS.n368 4.5005
R24918 DVSS.n383 DVSS.n335 4.5005
R24919 DVSS.n386 DVSS.n335 4.5005
R24920 DVSS.n381 DVSS.n335 4.5005
R24921 DVSS.n387 DVSS.n335 4.5005
R24922 DVSS.n380 DVSS.n335 4.5005
R24923 DVSS.n389 DVSS.n335 4.5005
R24924 DVSS.n379 DVSS.n335 4.5005
R24925 DVSS.n390 DVSS.n335 4.5005
R24926 DVSS.n378 DVSS.n335 4.5005
R24927 DVSS.n393 DVSS.n335 4.5005
R24928 DVSS.n377 DVSS.n335 4.5005
R24929 DVSS.n394 DVSS.n335 4.5005
R24930 DVSS.n23004 DVSS.n335 4.5005
R24931 DVSS.n376 DVSS.n335 4.5005
R24932 DVSS.n23002 DVSS.n335 4.5005
R24933 DVSS.n23003 DVSS.n383 4.5005
R24934 DVSS.n23003 DVSS.n386 4.5005
R24935 DVSS.n23003 DVSS.n381 4.5005
R24936 DVSS.n23003 DVSS.n387 4.5005
R24937 DVSS.n23003 DVSS.n380 4.5005
R24938 DVSS.n23003 DVSS.n389 4.5005
R24939 DVSS.n23003 DVSS.n379 4.5005
R24940 DVSS.n23003 DVSS.n390 4.5005
R24941 DVSS.n23003 DVSS.n378 4.5005
R24942 DVSS.n23003 DVSS.n393 4.5005
R24943 DVSS.n23003 DVSS.n377 4.5005
R24944 DVSS.n23003 DVSS.n394 4.5005
R24945 DVSS.n23003 DVSS.n334 4.5005
R24946 DVSS.n23004 DVSS.n23003 4.5005
R24947 DVSS.n23003 DVSS.n376 4.5005
R24948 DVSS.n23003 DVSS.n23002 4.5005
R24949 DVSS.n23221 DVSS.n16 4.5005
R24950 DVSS.n30 DVSS.n16 4.5005
R24951 DVSS.n23217 DVSS.n16 4.5005
R24952 DVSS.n31 DVSS.n16 4.5005
R24953 DVSS.n42 DVSS.n16 4.5005
R24954 DVSS.n32 DVSS.n16 4.5005
R24955 DVSS.n41 DVSS.n16 4.5005
R24956 DVSS.n34 DVSS.n16 4.5005
R24957 DVSS.n38 DVSS.n16 4.5005
R24958 DVSS.n37 DVSS.n16 4.5005
R24959 DVSS.n35 DVSS.n16 4.5005
R24960 DVSS.n37 DVSS.n17 4.5005
R24961 DVSS.n35 DVSS.n17 4.5005
R24962 DVSS.n38 DVSS.n17 4.5005
R24963 DVSS.n34 DVSS.n17 4.5005
R24964 DVSS.n40 DVSS.n17 4.5005
R24965 DVSS.n33 DVSS.n17 4.5005
R24966 DVSS.n41 DVSS.n17 4.5005
R24967 DVSS.n32 DVSS.n17 4.5005
R24968 DVSS.n42 DVSS.n17 4.5005
R24969 DVSS.n31 DVSS.n17 4.5005
R24970 DVSS.n23217 DVSS.n17 4.5005
R24971 DVSS.n30 DVSS.n17 4.5005
R24972 DVSS.n23219 DVSS.n17 4.5005
R24973 DVSS.n29 DVSS.n17 4.5005
R24974 DVSS.n23221 DVSS.n17 4.5005
R24975 DVSS.n37 DVSS.n15 4.5005
R24976 DVSS.n35 DVSS.n15 4.5005
R24977 DVSS.n38 DVSS.n15 4.5005
R24978 DVSS.n34 DVSS.n15 4.5005
R24979 DVSS.n40 DVSS.n15 4.5005
R24980 DVSS.n33 DVSS.n15 4.5005
R24981 DVSS.n41 DVSS.n15 4.5005
R24982 DVSS.n32 DVSS.n15 4.5005
R24983 DVSS.n42 DVSS.n15 4.5005
R24984 DVSS.n31 DVSS.n15 4.5005
R24985 DVSS.n23217 DVSS.n15 4.5005
R24986 DVSS.n30 DVSS.n15 4.5005
R24987 DVSS.n23219 DVSS.n15 4.5005
R24988 DVSS.n29 DVSS.n15 4.5005
R24989 DVSS.n23221 DVSS.n15 4.5005
R24990 DVSS.n37 DVSS.n18 4.5005
R24991 DVSS.n35 DVSS.n18 4.5005
R24992 DVSS.n38 DVSS.n18 4.5005
R24993 DVSS.n34 DVSS.n18 4.5005
R24994 DVSS.n40 DVSS.n18 4.5005
R24995 DVSS.n33 DVSS.n18 4.5005
R24996 DVSS.n41 DVSS.n18 4.5005
R24997 DVSS.n32 DVSS.n18 4.5005
R24998 DVSS.n42 DVSS.n18 4.5005
R24999 DVSS.n31 DVSS.n18 4.5005
R25000 DVSS.n23217 DVSS.n18 4.5005
R25001 DVSS.n30 DVSS.n18 4.5005
R25002 DVSS.n23219 DVSS.n18 4.5005
R25003 DVSS.n29 DVSS.n18 4.5005
R25004 DVSS.n23221 DVSS.n18 4.5005
R25005 DVSS.n23221 DVSS.n14 4.5005
R25006 DVSS.n29 DVSS.n14 4.5005
R25007 DVSS.n23219 DVSS.n14 4.5005
R25008 DVSS.n30 DVSS.n14 4.5005
R25009 DVSS.n23217 DVSS.n14 4.5005
R25010 DVSS.n31 DVSS.n14 4.5005
R25011 DVSS.n42 DVSS.n14 4.5005
R25012 DVSS.n32 DVSS.n14 4.5005
R25013 DVSS.n41 DVSS.n14 4.5005
R25014 DVSS.n33 DVSS.n14 4.5005
R25015 DVSS.n40 DVSS.n14 4.5005
R25016 DVSS.n34 DVSS.n14 4.5005
R25017 DVSS.n38 DVSS.n14 4.5005
R25018 DVSS.n37 DVSS.n14 4.5005
R25019 DVSS.n35 DVSS.n14 4.5005
R25020 DVSS.n23221 DVSS.n19 4.5005
R25021 DVSS.n29 DVSS.n19 4.5005
R25022 DVSS.n23219 DVSS.n19 4.5005
R25023 DVSS.n30 DVSS.n19 4.5005
R25024 DVSS.n23217 DVSS.n19 4.5005
R25025 DVSS.n31 DVSS.n19 4.5005
R25026 DVSS.n42 DVSS.n19 4.5005
R25027 DVSS.n32 DVSS.n19 4.5005
R25028 DVSS.n41 DVSS.n19 4.5005
R25029 DVSS.n33 DVSS.n19 4.5005
R25030 DVSS.n40 DVSS.n19 4.5005
R25031 DVSS.n34 DVSS.n19 4.5005
R25032 DVSS.n38 DVSS.n19 4.5005
R25033 DVSS.n37 DVSS.n19 4.5005
R25034 DVSS.n35 DVSS.n19 4.5005
R25035 DVSS.n23221 DVSS.n13 4.5005
R25036 DVSS.n29 DVSS.n13 4.5005
R25037 DVSS.n23219 DVSS.n13 4.5005
R25038 DVSS.n30 DVSS.n13 4.5005
R25039 DVSS.n23217 DVSS.n13 4.5005
R25040 DVSS.n31 DVSS.n13 4.5005
R25041 DVSS.n42 DVSS.n13 4.5005
R25042 DVSS.n32 DVSS.n13 4.5005
R25043 DVSS.n41 DVSS.n13 4.5005
R25044 DVSS.n33 DVSS.n13 4.5005
R25045 DVSS.n40 DVSS.n13 4.5005
R25046 DVSS.n34 DVSS.n13 4.5005
R25047 DVSS.n38 DVSS.n13 4.5005
R25048 DVSS.n37 DVSS.n13 4.5005
R25049 DVSS.n35 DVSS.n13 4.5005
R25050 DVSS.n23221 DVSS.n20 4.5005
R25051 DVSS.n29 DVSS.n20 4.5005
R25052 DVSS.n23219 DVSS.n20 4.5005
R25053 DVSS.n30 DVSS.n20 4.5005
R25054 DVSS.n23217 DVSS.n20 4.5005
R25055 DVSS.n31 DVSS.n20 4.5005
R25056 DVSS.n42 DVSS.n20 4.5005
R25057 DVSS.n32 DVSS.n20 4.5005
R25058 DVSS.n41 DVSS.n20 4.5005
R25059 DVSS.n33 DVSS.n20 4.5005
R25060 DVSS.n40 DVSS.n20 4.5005
R25061 DVSS.n34 DVSS.n20 4.5005
R25062 DVSS.n38 DVSS.n20 4.5005
R25063 DVSS.n37 DVSS.n20 4.5005
R25064 DVSS.n35 DVSS.n20 4.5005
R25065 DVSS.n37 DVSS.n12 4.5005
R25066 DVSS.n35 DVSS.n12 4.5005
R25067 DVSS.n38 DVSS.n12 4.5005
R25068 DVSS.n34 DVSS.n12 4.5005
R25069 DVSS.n40 DVSS.n12 4.5005
R25070 DVSS.n33 DVSS.n12 4.5005
R25071 DVSS.n41 DVSS.n12 4.5005
R25072 DVSS.n32 DVSS.n12 4.5005
R25073 DVSS.n42 DVSS.n12 4.5005
R25074 DVSS.n31 DVSS.n12 4.5005
R25075 DVSS.n23217 DVSS.n12 4.5005
R25076 DVSS.n30 DVSS.n12 4.5005
R25077 DVSS.n23219 DVSS.n12 4.5005
R25078 DVSS.n29 DVSS.n12 4.5005
R25079 DVSS.n23221 DVSS.n12 4.5005
R25080 DVSS.n37 DVSS.n21 4.5005
R25081 DVSS.n35 DVSS.n21 4.5005
R25082 DVSS.n38 DVSS.n21 4.5005
R25083 DVSS.n34 DVSS.n21 4.5005
R25084 DVSS.n40 DVSS.n21 4.5005
R25085 DVSS.n33 DVSS.n21 4.5005
R25086 DVSS.n41 DVSS.n21 4.5005
R25087 DVSS.n32 DVSS.n21 4.5005
R25088 DVSS.n42 DVSS.n21 4.5005
R25089 DVSS.n31 DVSS.n21 4.5005
R25090 DVSS.n23217 DVSS.n21 4.5005
R25091 DVSS.n30 DVSS.n21 4.5005
R25092 DVSS.n23219 DVSS.n21 4.5005
R25093 DVSS.n29 DVSS.n21 4.5005
R25094 DVSS.n23221 DVSS.n21 4.5005
R25095 DVSS.n37 DVSS.n11 4.5005
R25096 DVSS.n35 DVSS.n11 4.5005
R25097 DVSS.n38 DVSS.n11 4.5005
R25098 DVSS.n34 DVSS.n11 4.5005
R25099 DVSS.n40 DVSS.n11 4.5005
R25100 DVSS.n33 DVSS.n11 4.5005
R25101 DVSS.n41 DVSS.n11 4.5005
R25102 DVSS.n32 DVSS.n11 4.5005
R25103 DVSS.n42 DVSS.n11 4.5005
R25104 DVSS.n31 DVSS.n11 4.5005
R25105 DVSS.n23217 DVSS.n11 4.5005
R25106 DVSS.n30 DVSS.n11 4.5005
R25107 DVSS.n23219 DVSS.n11 4.5005
R25108 DVSS.n29 DVSS.n11 4.5005
R25109 DVSS.n23221 DVSS.n11 4.5005
R25110 DVSS.n23221 DVSS.n22 4.5005
R25111 DVSS.n29 DVSS.n22 4.5005
R25112 DVSS.n23219 DVSS.n22 4.5005
R25113 DVSS.n30 DVSS.n22 4.5005
R25114 DVSS.n23217 DVSS.n22 4.5005
R25115 DVSS.n31 DVSS.n22 4.5005
R25116 DVSS.n42 DVSS.n22 4.5005
R25117 DVSS.n32 DVSS.n22 4.5005
R25118 DVSS.n41 DVSS.n22 4.5005
R25119 DVSS.n33 DVSS.n22 4.5005
R25120 DVSS.n40 DVSS.n22 4.5005
R25121 DVSS.n34 DVSS.n22 4.5005
R25122 DVSS.n38 DVSS.n22 4.5005
R25123 DVSS.n37 DVSS.n22 4.5005
R25124 DVSS.n35 DVSS.n22 4.5005
R25125 DVSS.n23221 DVSS.n10 4.5005
R25126 DVSS.n29 DVSS.n10 4.5005
R25127 DVSS.n23219 DVSS.n10 4.5005
R25128 DVSS.n30 DVSS.n10 4.5005
R25129 DVSS.n23217 DVSS.n10 4.5005
R25130 DVSS.n31 DVSS.n10 4.5005
R25131 DVSS.n42 DVSS.n10 4.5005
R25132 DVSS.n32 DVSS.n10 4.5005
R25133 DVSS.n41 DVSS.n10 4.5005
R25134 DVSS.n33 DVSS.n10 4.5005
R25135 DVSS.n40 DVSS.n10 4.5005
R25136 DVSS.n34 DVSS.n10 4.5005
R25137 DVSS.n38 DVSS.n10 4.5005
R25138 DVSS.n37 DVSS.n10 4.5005
R25139 DVSS.n35 DVSS.n10 4.5005
R25140 DVSS.n23221 DVSS.n23 4.5005
R25141 DVSS.n29 DVSS.n23 4.5005
R25142 DVSS.n23219 DVSS.n23 4.5005
R25143 DVSS.n30 DVSS.n23 4.5005
R25144 DVSS.n23217 DVSS.n23 4.5005
R25145 DVSS.n31 DVSS.n23 4.5005
R25146 DVSS.n42 DVSS.n23 4.5005
R25147 DVSS.n32 DVSS.n23 4.5005
R25148 DVSS.n41 DVSS.n23 4.5005
R25149 DVSS.n33 DVSS.n23 4.5005
R25150 DVSS.n40 DVSS.n23 4.5005
R25151 DVSS.n34 DVSS.n23 4.5005
R25152 DVSS.n38 DVSS.n23 4.5005
R25153 DVSS.n37 DVSS.n23 4.5005
R25154 DVSS.n35 DVSS.n23 4.5005
R25155 DVSS.n23221 DVSS.n9 4.5005
R25156 DVSS.n29 DVSS.n9 4.5005
R25157 DVSS.n23219 DVSS.n9 4.5005
R25158 DVSS.n30 DVSS.n9 4.5005
R25159 DVSS.n23217 DVSS.n9 4.5005
R25160 DVSS.n31 DVSS.n9 4.5005
R25161 DVSS.n42 DVSS.n9 4.5005
R25162 DVSS.n32 DVSS.n9 4.5005
R25163 DVSS.n41 DVSS.n9 4.5005
R25164 DVSS.n33 DVSS.n9 4.5005
R25165 DVSS.n40 DVSS.n9 4.5005
R25166 DVSS.n34 DVSS.n9 4.5005
R25167 DVSS.n38 DVSS.n9 4.5005
R25168 DVSS.n37 DVSS.n9 4.5005
R25169 DVSS.n35 DVSS.n9 4.5005
R25170 DVSS.n37 DVSS.n24 4.5005
R25171 DVSS.n35 DVSS.n24 4.5005
R25172 DVSS.n38 DVSS.n24 4.5005
R25173 DVSS.n34 DVSS.n24 4.5005
R25174 DVSS.n40 DVSS.n24 4.5005
R25175 DVSS.n33 DVSS.n24 4.5005
R25176 DVSS.n41 DVSS.n24 4.5005
R25177 DVSS.n32 DVSS.n24 4.5005
R25178 DVSS.n42 DVSS.n24 4.5005
R25179 DVSS.n31 DVSS.n24 4.5005
R25180 DVSS.n23217 DVSS.n24 4.5005
R25181 DVSS.n30 DVSS.n24 4.5005
R25182 DVSS.n23219 DVSS.n24 4.5005
R25183 DVSS.n29 DVSS.n24 4.5005
R25184 DVSS.n23221 DVSS.n24 4.5005
R25185 DVSS.n37 DVSS.n8 4.5005
R25186 DVSS.n35 DVSS.n8 4.5005
R25187 DVSS.n38 DVSS.n8 4.5005
R25188 DVSS.n34 DVSS.n8 4.5005
R25189 DVSS.n40 DVSS.n8 4.5005
R25190 DVSS.n33 DVSS.n8 4.5005
R25191 DVSS.n41 DVSS.n8 4.5005
R25192 DVSS.n32 DVSS.n8 4.5005
R25193 DVSS.n42 DVSS.n8 4.5005
R25194 DVSS.n31 DVSS.n8 4.5005
R25195 DVSS.n23217 DVSS.n8 4.5005
R25196 DVSS.n30 DVSS.n8 4.5005
R25197 DVSS.n23219 DVSS.n8 4.5005
R25198 DVSS.n29 DVSS.n8 4.5005
R25199 DVSS.n23221 DVSS.n8 4.5005
R25200 DVSS.n37 DVSS.n25 4.5005
R25201 DVSS.n35 DVSS.n25 4.5005
R25202 DVSS.n38 DVSS.n25 4.5005
R25203 DVSS.n34 DVSS.n25 4.5005
R25204 DVSS.n40 DVSS.n25 4.5005
R25205 DVSS.n33 DVSS.n25 4.5005
R25206 DVSS.n41 DVSS.n25 4.5005
R25207 DVSS.n32 DVSS.n25 4.5005
R25208 DVSS.n42 DVSS.n25 4.5005
R25209 DVSS.n31 DVSS.n25 4.5005
R25210 DVSS.n23217 DVSS.n25 4.5005
R25211 DVSS.n30 DVSS.n25 4.5005
R25212 DVSS.n23219 DVSS.n25 4.5005
R25213 DVSS.n29 DVSS.n25 4.5005
R25214 DVSS.n23221 DVSS.n25 4.5005
R25215 DVSS.n23221 DVSS.n7 4.5005
R25216 DVSS.n29 DVSS.n7 4.5005
R25217 DVSS.n23219 DVSS.n7 4.5005
R25218 DVSS.n30 DVSS.n7 4.5005
R25219 DVSS.n23217 DVSS.n7 4.5005
R25220 DVSS.n31 DVSS.n7 4.5005
R25221 DVSS.n42 DVSS.n7 4.5005
R25222 DVSS.n32 DVSS.n7 4.5005
R25223 DVSS.n41 DVSS.n7 4.5005
R25224 DVSS.n33 DVSS.n7 4.5005
R25225 DVSS.n40 DVSS.n7 4.5005
R25226 DVSS.n34 DVSS.n7 4.5005
R25227 DVSS.n38 DVSS.n7 4.5005
R25228 DVSS.n37 DVSS.n7 4.5005
R25229 DVSS.n35 DVSS.n7 4.5005
R25230 DVSS.n23221 DVSS.n26 4.5005
R25231 DVSS.n29 DVSS.n26 4.5005
R25232 DVSS.n23219 DVSS.n26 4.5005
R25233 DVSS.n30 DVSS.n26 4.5005
R25234 DVSS.n23217 DVSS.n26 4.5005
R25235 DVSS.n31 DVSS.n26 4.5005
R25236 DVSS.n42 DVSS.n26 4.5005
R25237 DVSS.n32 DVSS.n26 4.5005
R25238 DVSS.n41 DVSS.n26 4.5005
R25239 DVSS.n33 DVSS.n26 4.5005
R25240 DVSS.n40 DVSS.n26 4.5005
R25241 DVSS.n34 DVSS.n26 4.5005
R25242 DVSS.n38 DVSS.n26 4.5005
R25243 DVSS.n37 DVSS.n26 4.5005
R25244 DVSS.n35 DVSS.n26 4.5005
R25245 DVSS.n23221 DVSS.n6 4.5005
R25246 DVSS.n29 DVSS.n6 4.5005
R25247 DVSS.n23219 DVSS.n6 4.5005
R25248 DVSS.n30 DVSS.n6 4.5005
R25249 DVSS.n23217 DVSS.n6 4.5005
R25250 DVSS.n31 DVSS.n6 4.5005
R25251 DVSS.n42 DVSS.n6 4.5005
R25252 DVSS.n32 DVSS.n6 4.5005
R25253 DVSS.n41 DVSS.n6 4.5005
R25254 DVSS.n33 DVSS.n6 4.5005
R25255 DVSS.n40 DVSS.n6 4.5005
R25256 DVSS.n34 DVSS.n6 4.5005
R25257 DVSS.n38 DVSS.n6 4.5005
R25258 DVSS.n37 DVSS.n6 4.5005
R25259 DVSS.n35 DVSS.n6 4.5005
R25260 DVSS.n37 DVSS.n27 4.5005
R25261 DVSS.n35 DVSS.n27 4.5005
R25262 DVSS.n38 DVSS.n27 4.5005
R25263 DVSS.n34 DVSS.n27 4.5005
R25264 DVSS.n40 DVSS.n27 4.5005
R25265 DVSS.n33 DVSS.n27 4.5005
R25266 DVSS.n41 DVSS.n27 4.5005
R25267 DVSS.n32 DVSS.n27 4.5005
R25268 DVSS.n42 DVSS.n27 4.5005
R25269 DVSS.n31 DVSS.n27 4.5005
R25270 DVSS.n23217 DVSS.n27 4.5005
R25271 DVSS.n30 DVSS.n27 4.5005
R25272 DVSS.n23219 DVSS.n27 4.5005
R25273 DVSS.n29 DVSS.n27 4.5005
R25274 DVSS.n23221 DVSS.n27 4.5005
R25275 DVSS.n37 DVSS.n5 4.5005
R25276 DVSS.n35 DVSS.n5 4.5005
R25277 DVSS.n38 DVSS.n5 4.5005
R25278 DVSS.n34 DVSS.n5 4.5005
R25279 DVSS.n40 DVSS.n5 4.5005
R25280 DVSS.n33 DVSS.n5 4.5005
R25281 DVSS.n41 DVSS.n5 4.5005
R25282 DVSS.n32 DVSS.n5 4.5005
R25283 DVSS.n42 DVSS.n5 4.5005
R25284 DVSS.n31 DVSS.n5 4.5005
R25285 DVSS.n23217 DVSS.n5 4.5005
R25286 DVSS.n30 DVSS.n5 4.5005
R25287 DVSS.n23219 DVSS.n5 4.5005
R25288 DVSS.n29 DVSS.n5 4.5005
R25289 DVSS.n23221 DVSS.n5 4.5005
R25290 DVSS.n23220 DVSS.n37 4.5005
R25291 DVSS.n23220 DVSS.n35 4.5005
R25292 DVSS.n23220 DVSS.n38 4.5005
R25293 DVSS.n23220 DVSS.n34 4.5005
R25294 DVSS.n23220 DVSS.n40 4.5005
R25295 DVSS.n23220 DVSS.n33 4.5005
R25296 DVSS.n23220 DVSS.n41 4.5005
R25297 DVSS.n23220 DVSS.n32 4.5005
R25298 DVSS.n23220 DVSS.n42 4.5005
R25299 DVSS.n23220 DVSS.n31 4.5005
R25300 DVSS.n23220 DVSS.n23217 4.5005
R25301 DVSS.n23220 DVSS.n30 4.5005
R25302 DVSS.n23220 DVSS.n23219 4.5005
R25303 DVSS.n23220 DVSS.n29 4.5005
R25304 DVSS.n23221 DVSS.n23220 4.5005
R25305 DVSS.n22452 DVSS.n913 4.5005
R25306 DVSS.n913 DVSS.n883 4.5005
R25307 DVSS.n913 DVSS.n898 4.5005
R25308 DVSS.n913 DVSS.n884 4.5005
R25309 DVSS.n913 DVSS.n896 4.5005
R25310 DVSS.n913 DVSS.n885 4.5005
R25311 DVSS.n913 DVSS.n895 4.5005
R25312 DVSS.n913 DVSS.n887 4.5005
R25313 DVSS.n913 DVSS.n892 4.5005
R25314 DVSS.n913 DVSS.n891 4.5005
R25315 DVSS.n913 DVSS.n888 4.5005
R25316 DVSS.n22452 DVSS.n914 4.5005
R25317 DVSS.n914 DVSS.n882 4.5005
R25318 DVSS.n914 DVSS.n899 4.5005
R25319 DVSS.n914 DVSS.n883 4.5005
R25320 DVSS.n914 DVSS.n898 4.5005
R25321 DVSS.n914 DVSS.n884 4.5005
R25322 DVSS.n914 DVSS.n896 4.5005
R25323 DVSS.n914 DVSS.n885 4.5005
R25324 DVSS.n914 DVSS.n895 4.5005
R25325 DVSS.n914 DVSS.n886 4.5005
R25326 DVSS.n914 DVSS.n893 4.5005
R25327 DVSS.n914 DVSS.n887 4.5005
R25328 DVSS.n914 DVSS.n892 4.5005
R25329 DVSS.n914 DVSS.n891 4.5005
R25330 DVSS.n914 DVSS.n888 4.5005
R25331 DVSS.n22452 DVSS.n910 4.5005
R25332 DVSS.n910 DVSS.n882 4.5005
R25333 DVSS.n910 DVSS.n899 4.5005
R25334 DVSS.n910 DVSS.n883 4.5005
R25335 DVSS.n910 DVSS.n898 4.5005
R25336 DVSS.n910 DVSS.n884 4.5005
R25337 DVSS.n910 DVSS.n896 4.5005
R25338 DVSS.n910 DVSS.n885 4.5005
R25339 DVSS.n910 DVSS.n895 4.5005
R25340 DVSS.n910 DVSS.n886 4.5005
R25341 DVSS.n910 DVSS.n893 4.5005
R25342 DVSS.n910 DVSS.n887 4.5005
R25343 DVSS.n910 DVSS.n892 4.5005
R25344 DVSS.n910 DVSS.n891 4.5005
R25345 DVSS.n910 DVSS.n888 4.5005
R25346 DVSS.n22451 DVSS.n891 4.5005
R25347 DVSS.n22451 DVSS.n888 4.5005
R25348 DVSS.n900 DVSS.n891 4.5005
R25349 DVSS.n900 DVSS.n888 4.5005
R25350 DVSS.n923 DVSS.n891 4.5005
R25351 DVSS.n923 DVSS.n888 4.5005
R25352 DVSS.n22452 DVSS.n915 4.5005
R25353 DVSS.n915 DVSS.n882 4.5005
R25354 DVSS.n915 DVSS.n899 4.5005
R25355 DVSS.n915 DVSS.n883 4.5005
R25356 DVSS.n915 DVSS.n898 4.5005
R25357 DVSS.n915 DVSS.n884 4.5005
R25358 DVSS.n915 DVSS.n896 4.5005
R25359 DVSS.n915 DVSS.n885 4.5005
R25360 DVSS.n915 DVSS.n895 4.5005
R25361 DVSS.n915 DVSS.n886 4.5005
R25362 DVSS.n915 DVSS.n893 4.5005
R25363 DVSS.n915 DVSS.n887 4.5005
R25364 DVSS.n915 DVSS.n892 4.5005
R25365 DVSS.n915 DVSS.n891 4.5005
R25366 DVSS.n915 DVSS.n888 4.5005
R25367 DVSS.n22452 DVSS.n909 4.5005
R25368 DVSS.n909 DVSS.n882 4.5005
R25369 DVSS.n909 DVSS.n899 4.5005
R25370 DVSS.n909 DVSS.n883 4.5005
R25371 DVSS.n909 DVSS.n898 4.5005
R25372 DVSS.n909 DVSS.n884 4.5005
R25373 DVSS.n909 DVSS.n896 4.5005
R25374 DVSS.n909 DVSS.n885 4.5005
R25375 DVSS.n909 DVSS.n895 4.5005
R25376 DVSS.n909 DVSS.n886 4.5005
R25377 DVSS.n909 DVSS.n893 4.5005
R25378 DVSS.n909 DVSS.n887 4.5005
R25379 DVSS.n909 DVSS.n892 4.5005
R25380 DVSS.n909 DVSS.n891 4.5005
R25381 DVSS.n909 DVSS.n888 4.5005
R25382 DVSS.n22452 DVSS.n916 4.5005
R25383 DVSS.n916 DVSS.n882 4.5005
R25384 DVSS.n916 DVSS.n899 4.5005
R25385 DVSS.n916 DVSS.n883 4.5005
R25386 DVSS.n916 DVSS.n898 4.5005
R25387 DVSS.n916 DVSS.n884 4.5005
R25388 DVSS.n916 DVSS.n896 4.5005
R25389 DVSS.n916 DVSS.n885 4.5005
R25390 DVSS.n916 DVSS.n895 4.5005
R25391 DVSS.n916 DVSS.n886 4.5005
R25392 DVSS.n916 DVSS.n893 4.5005
R25393 DVSS.n916 DVSS.n887 4.5005
R25394 DVSS.n916 DVSS.n892 4.5005
R25395 DVSS.n916 DVSS.n891 4.5005
R25396 DVSS.n916 DVSS.n888 4.5005
R25397 DVSS.n22452 DVSS.n908 4.5005
R25398 DVSS.n908 DVSS.n882 4.5005
R25399 DVSS.n908 DVSS.n899 4.5005
R25400 DVSS.n908 DVSS.n883 4.5005
R25401 DVSS.n908 DVSS.n898 4.5005
R25402 DVSS.n908 DVSS.n884 4.5005
R25403 DVSS.n908 DVSS.n896 4.5005
R25404 DVSS.n908 DVSS.n885 4.5005
R25405 DVSS.n908 DVSS.n895 4.5005
R25406 DVSS.n908 DVSS.n886 4.5005
R25407 DVSS.n908 DVSS.n893 4.5005
R25408 DVSS.n908 DVSS.n887 4.5005
R25409 DVSS.n908 DVSS.n892 4.5005
R25410 DVSS.n908 DVSS.n891 4.5005
R25411 DVSS.n908 DVSS.n888 4.5005
R25412 DVSS.n901 DVSS.n891 4.5005
R25413 DVSS.n901 DVSS.n888 4.5005
R25414 DVSS.n922 DVSS.n891 4.5005
R25415 DVSS.n922 DVSS.n888 4.5005
R25416 DVSS.n902 DVSS.n891 4.5005
R25417 DVSS.n902 DVSS.n888 4.5005
R25418 DVSS.n22452 DVSS.n917 4.5005
R25419 DVSS.n917 DVSS.n882 4.5005
R25420 DVSS.n917 DVSS.n899 4.5005
R25421 DVSS.n917 DVSS.n883 4.5005
R25422 DVSS.n917 DVSS.n898 4.5005
R25423 DVSS.n917 DVSS.n884 4.5005
R25424 DVSS.n917 DVSS.n896 4.5005
R25425 DVSS.n917 DVSS.n885 4.5005
R25426 DVSS.n917 DVSS.n895 4.5005
R25427 DVSS.n917 DVSS.n886 4.5005
R25428 DVSS.n917 DVSS.n893 4.5005
R25429 DVSS.n917 DVSS.n887 4.5005
R25430 DVSS.n917 DVSS.n892 4.5005
R25431 DVSS.n917 DVSS.n891 4.5005
R25432 DVSS.n917 DVSS.n888 4.5005
R25433 DVSS.n22452 DVSS.n907 4.5005
R25434 DVSS.n907 DVSS.n882 4.5005
R25435 DVSS.n907 DVSS.n899 4.5005
R25436 DVSS.n907 DVSS.n883 4.5005
R25437 DVSS.n907 DVSS.n898 4.5005
R25438 DVSS.n907 DVSS.n884 4.5005
R25439 DVSS.n907 DVSS.n896 4.5005
R25440 DVSS.n907 DVSS.n885 4.5005
R25441 DVSS.n907 DVSS.n895 4.5005
R25442 DVSS.n907 DVSS.n886 4.5005
R25443 DVSS.n907 DVSS.n893 4.5005
R25444 DVSS.n907 DVSS.n887 4.5005
R25445 DVSS.n907 DVSS.n892 4.5005
R25446 DVSS.n907 DVSS.n891 4.5005
R25447 DVSS.n907 DVSS.n888 4.5005
R25448 DVSS.n22452 DVSS.n918 4.5005
R25449 DVSS.n918 DVSS.n882 4.5005
R25450 DVSS.n918 DVSS.n899 4.5005
R25451 DVSS.n918 DVSS.n883 4.5005
R25452 DVSS.n918 DVSS.n898 4.5005
R25453 DVSS.n918 DVSS.n884 4.5005
R25454 DVSS.n918 DVSS.n896 4.5005
R25455 DVSS.n918 DVSS.n885 4.5005
R25456 DVSS.n918 DVSS.n895 4.5005
R25457 DVSS.n918 DVSS.n886 4.5005
R25458 DVSS.n918 DVSS.n893 4.5005
R25459 DVSS.n918 DVSS.n887 4.5005
R25460 DVSS.n918 DVSS.n892 4.5005
R25461 DVSS.n918 DVSS.n891 4.5005
R25462 DVSS.n918 DVSS.n888 4.5005
R25463 DVSS.n921 DVSS.n891 4.5005
R25464 DVSS.n921 DVSS.n888 4.5005
R25465 DVSS.n903 DVSS.n891 4.5005
R25466 DVSS.n903 DVSS.n888 4.5005
R25467 DVSS.n920 DVSS.n891 4.5005
R25468 DVSS.n920 DVSS.n888 4.5005
R25469 DVSS.n904 DVSS.n891 4.5005
R25470 DVSS.n904 DVSS.n888 4.5005
R25471 DVSS.n22452 DVSS.n906 4.5005
R25472 DVSS.n906 DVSS.n882 4.5005
R25473 DVSS.n906 DVSS.n899 4.5005
R25474 DVSS.n906 DVSS.n883 4.5005
R25475 DVSS.n906 DVSS.n898 4.5005
R25476 DVSS.n906 DVSS.n884 4.5005
R25477 DVSS.n906 DVSS.n896 4.5005
R25478 DVSS.n906 DVSS.n885 4.5005
R25479 DVSS.n906 DVSS.n895 4.5005
R25480 DVSS.n906 DVSS.n886 4.5005
R25481 DVSS.n906 DVSS.n893 4.5005
R25482 DVSS.n906 DVSS.n887 4.5005
R25483 DVSS.n906 DVSS.n892 4.5005
R25484 DVSS.n906 DVSS.n891 4.5005
R25485 DVSS.n906 DVSS.n888 4.5005
R25486 DVSS.n22452 DVSS.n919 4.5005
R25487 DVSS.n919 DVSS.n882 4.5005
R25488 DVSS.n919 DVSS.n899 4.5005
R25489 DVSS.n919 DVSS.n883 4.5005
R25490 DVSS.n919 DVSS.n898 4.5005
R25491 DVSS.n919 DVSS.n884 4.5005
R25492 DVSS.n919 DVSS.n896 4.5005
R25493 DVSS.n919 DVSS.n885 4.5005
R25494 DVSS.n919 DVSS.n895 4.5005
R25495 DVSS.n919 DVSS.n886 4.5005
R25496 DVSS.n919 DVSS.n893 4.5005
R25497 DVSS.n919 DVSS.n887 4.5005
R25498 DVSS.n919 DVSS.n892 4.5005
R25499 DVSS.n919 DVSS.n891 4.5005
R25500 DVSS.n919 DVSS.n888 4.5005
R25501 DVSS.n22452 DVSS.n905 4.5005
R25502 DVSS.n905 DVSS.n882 4.5005
R25503 DVSS.n905 DVSS.n899 4.5005
R25504 DVSS.n905 DVSS.n883 4.5005
R25505 DVSS.n905 DVSS.n898 4.5005
R25506 DVSS.n905 DVSS.n884 4.5005
R25507 DVSS.n905 DVSS.n896 4.5005
R25508 DVSS.n905 DVSS.n885 4.5005
R25509 DVSS.n905 DVSS.n895 4.5005
R25510 DVSS.n905 DVSS.n886 4.5005
R25511 DVSS.n905 DVSS.n893 4.5005
R25512 DVSS.n905 DVSS.n887 4.5005
R25513 DVSS.n905 DVSS.n892 4.5005
R25514 DVSS.n905 DVSS.n891 4.5005
R25515 DVSS.n905 DVSS.n888 4.5005
R25516 DVSS.n22453 DVSS.n891 4.5005
R25517 DVSS.n22453 DVSS.n888 4.5005
R25518 DVSS.n22453 DVSS.n892 4.5005
R25519 DVSS.n22453 DVSS.n887 4.5005
R25520 DVSS.n22453 DVSS.n893 4.5005
R25521 DVSS.n22453 DVSS.n886 4.5005
R25522 DVSS.n22453 DVSS.n895 4.5005
R25523 DVSS.n22453 DVSS.n885 4.5005
R25524 DVSS.n22453 DVSS.n896 4.5005
R25525 DVSS.n22453 DVSS.n884 4.5005
R25526 DVSS.n22453 DVSS.n898 4.5005
R25527 DVSS.n22453 DVSS.n883 4.5005
R25528 DVSS.n22453 DVSS.n899 4.5005
R25529 DVSS.n22453 DVSS.n882 4.5005
R25530 DVSS.n22453 DVSS.n22452 4.5005
R25531 DVSS.n904 DVSS.n892 4.5005
R25532 DVSS.n904 DVSS.n887 4.5005
R25533 DVSS.n904 DVSS.n893 4.5005
R25534 DVSS.n904 DVSS.n886 4.5005
R25535 DVSS.n904 DVSS.n895 4.5005
R25536 DVSS.n904 DVSS.n885 4.5005
R25537 DVSS.n904 DVSS.n896 4.5005
R25538 DVSS.n904 DVSS.n884 4.5005
R25539 DVSS.n904 DVSS.n898 4.5005
R25540 DVSS.n904 DVSS.n883 4.5005
R25541 DVSS.n904 DVSS.n899 4.5005
R25542 DVSS.n904 DVSS.n882 4.5005
R25543 DVSS.n22452 DVSS.n904 4.5005
R25544 DVSS.n920 DVSS.n892 4.5005
R25545 DVSS.n920 DVSS.n887 4.5005
R25546 DVSS.n920 DVSS.n893 4.5005
R25547 DVSS.n920 DVSS.n886 4.5005
R25548 DVSS.n920 DVSS.n895 4.5005
R25549 DVSS.n920 DVSS.n885 4.5005
R25550 DVSS.n920 DVSS.n896 4.5005
R25551 DVSS.n920 DVSS.n884 4.5005
R25552 DVSS.n920 DVSS.n898 4.5005
R25553 DVSS.n920 DVSS.n883 4.5005
R25554 DVSS.n920 DVSS.n899 4.5005
R25555 DVSS.n920 DVSS.n882 4.5005
R25556 DVSS.n22452 DVSS.n920 4.5005
R25557 DVSS.n903 DVSS.n892 4.5005
R25558 DVSS.n903 DVSS.n887 4.5005
R25559 DVSS.n903 DVSS.n893 4.5005
R25560 DVSS.n903 DVSS.n886 4.5005
R25561 DVSS.n903 DVSS.n895 4.5005
R25562 DVSS.n903 DVSS.n885 4.5005
R25563 DVSS.n903 DVSS.n896 4.5005
R25564 DVSS.n903 DVSS.n884 4.5005
R25565 DVSS.n903 DVSS.n898 4.5005
R25566 DVSS.n903 DVSS.n883 4.5005
R25567 DVSS.n903 DVSS.n899 4.5005
R25568 DVSS.n903 DVSS.n882 4.5005
R25569 DVSS.n22452 DVSS.n903 4.5005
R25570 DVSS.n921 DVSS.n892 4.5005
R25571 DVSS.n921 DVSS.n887 4.5005
R25572 DVSS.n921 DVSS.n893 4.5005
R25573 DVSS.n921 DVSS.n886 4.5005
R25574 DVSS.n921 DVSS.n895 4.5005
R25575 DVSS.n921 DVSS.n885 4.5005
R25576 DVSS.n921 DVSS.n896 4.5005
R25577 DVSS.n921 DVSS.n884 4.5005
R25578 DVSS.n921 DVSS.n898 4.5005
R25579 DVSS.n921 DVSS.n883 4.5005
R25580 DVSS.n921 DVSS.n899 4.5005
R25581 DVSS.n921 DVSS.n882 4.5005
R25582 DVSS.n22452 DVSS.n921 4.5005
R25583 DVSS.n902 DVSS.n892 4.5005
R25584 DVSS.n902 DVSS.n887 4.5005
R25585 DVSS.n902 DVSS.n893 4.5005
R25586 DVSS.n902 DVSS.n886 4.5005
R25587 DVSS.n902 DVSS.n895 4.5005
R25588 DVSS.n902 DVSS.n885 4.5005
R25589 DVSS.n902 DVSS.n896 4.5005
R25590 DVSS.n902 DVSS.n884 4.5005
R25591 DVSS.n902 DVSS.n898 4.5005
R25592 DVSS.n902 DVSS.n883 4.5005
R25593 DVSS.n902 DVSS.n899 4.5005
R25594 DVSS.n902 DVSS.n882 4.5005
R25595 DVSS.n22452 DVSS.n902 4.5005
R25596 DVSS.n922 DVSS.n892 4.5005
R25597 DVSS.n922 DVSS.n887 4.5005
R25598 DVSS.n922 DVSS.n893 4.5005
R25599 DVSS.n922 DVSS.n886 4.5005
R25600 DVSS.n922 DVSS.n895 4.5005
R25601 DVSS.n922 DVSS.n885 4.5005
R25602 DVSS.n922 DVSS.n896 4.5005
R25603 DVSS.n922 DVSS.n884 4.5005
R25604 DVSS.n922 DVSS.n898 4.5005
R25605 DVSS.n922 DVSS.n883 4.5005
R25606 DVSS.n922 DVSS.n899 4.5005
R25607 DVSS.n922 DVSS.n882 4.5005
R25608 DVSS.n22452 DVSS.n922 4.5005
R25609 DVSS.n901 DVSS.n892 4.5005
R25610 DVSS.n901 DVSS.n887 4.5005
R25611 DVSS.n901 DVSS.n893 4.5005
R25612 DVSS.n901 DVSS.n886 4.5005
R25613 DVSS.n901 DVSS.n895 4.5005
R25614 DVSS.n901 DVSS.n885 4.5005
R25615 DVSS.n901 DVSS.n896 4.5005
R25616 DVSS.n901 DVSS.n884 4.5005
R25617 DVSS.n901 DVSS.n898 4.5005
R25618 DVSS.n901 DVSS.n883 4.5005
R25619 DVSS.n901 DVSS.n899 4.5005
R25620 DVSS.n901 DVSS.n882 4.5005
R25621 DVSS.n22452 DVSS.n901 4.5005
R25622 DVSS.n923 DVSS.n892 4.5005
R25623 DVSS.n923 DVSS.n887 4.5005
R25624 DVSS.n923 DVSS.n893 4.5005
R25625 DVSS.n923 DVSS.n886 4.5005
R25626 DVSS.n923 DVSS.n895 4.5005
R25627 DVSS.n923 DVSS.n885 4.5005
R25628 DVSS.n923 DVSS.n896 4.5005
R25629 DVSS.n923 DVSS.n884 4.5005
R25630 DVSS.n923 DVSS.n898 4.5005
R25631 DVSS.n923 DVSS.n883 4.5005
R25632 DVSS.n923 DVSS.n899 4.5005
R25633 DVSS.n923 DVSS.n882 4.5005
R25634 DVSS.n22452 DVSS.n923 4.5005
R25635 DVSS.n900 DVSS.n892 4.5005
R25636 DVSS.n900 DVSS.n887 4.5005
R25637 DVSS.n900 DVSS.n893 4.5005
R25638 DVSS.n900 DVSS.n886 4.5005
R25639 DVSS.n900 DVSS.n895 4.5005
R25640 DVSS.n900 DVSS.n885 4.5005
R25641 DVSS.n900 DVSS.n896 4.5005
R25642 DVSS.n900 DVSS.n884 4.5005
R25643 DVSS.n900 DVSS.n898 4.5005
R25644 DVSS.n900 DVSS.n883 4.5005
R25645 DVSS.n900 DVSS.n899 4.5005
R25646 DVSS.n900 DVSS.n882 4.5005
R25647 DVSS.n22452 DVSS.n900 4.5005
R25648 DVSS.n22451 DVSS.n892 4.5005
R25649 DVSS.n22451 DVSS.n887 4.5005
R25650 DVSS.n22451 DVSS.n893 4.5005
R25651 DVSS.n22451 DVSS.n886 4.5005
R25652 DVSS.n22451 DVSS.n895 4.5005
R25653 DVSS.n22451 DVSS.n885 4.5005
R25654 DVSS.n22451 DVSS.n896 4.5005
R25655 DVSS.n22451 DVSS.n884 4.5005
R25656 DVSS.n22451 DVSS.n898 4.5005
R25657 DVSS.n22451 DVSS.n883 4.5005
R25658 DVSS.n22451 DVSS.n899 4.5005
R25659 DVSS.n22451 DVSS.n882 4.5005
R25660 DVSS.n22452 DVSS.n22451 4.5005
R25661 DVSS.n22478 DVSS.n813 4.5005
R25662 DVSS.n22483 DVSS.n813 4.5005
R25663 DVSS.n22477 DVSS.n813 4.5005
R25664 DVSS.n22485 DVSS.n813 4.5005
R25665 DVSS.n22476 DVSS.n813 4.5005
R25666 DVSS.n22489 DVSS.n813 4.5005
R25667 DVSS.n22474 DVSS.n813 4.5005
R25668 DVSS.n22490 DVSS.n813 4.5005
R25669 DVSS.n22473 DVSS.n813 4.5005
R25670 DVSS.n22500 DVSS.n813 4.5005
R25671 DVSS.n22498 DVSS.n813 4.5005
R25672 DVSS.n22504 DVSS.n813 4.5005
R25673 DVSS.n22478 DVSS.n814 4.5005
R25674 DVSS.n22483 DVSS.n814 4.5005
R25675 DVSS.n22477 DVSS.n814 4.5005
R25676 DVSS.n22485 DVSS.n814 4.5005
R25677 DVSS.n22476 DVSS.n814 4.5005
R25678 DVSS.n22487 DVSS.n814 4.5005
R25679 DVSS.n22475 DVSS.n814 4.5005
R25680 DVSS.n22489 DVSS.n814 4.5005
R25681 DVSS.n22474 DVSS.n814 4.5005
R25682 DVSS.n22490 DVSS.n814 4.5005
R25683 DVSS.n22473 DVSS.n814 4.5005
R25684 DVSS.n22500 DVSS.n814 4.5005
R25685 DVSS.n22502 DVSS.n814 4.5005
R25686 DVSS.n22504 DVSS.n814 4.5005
R25687 DVSS.n22478 DVSS.n812 4.5005
R25688 DVSS.n22483 DVSS.n812 4.5005
R25689 DVSS.n22477 DVSS.n812 4.5005
R25690 DVSS.n22485 DVSS.n812 4.5005
R25691 DVSS.n22476 DVSS.n812 4.5005
R25692 DVSS.n22487 DVSS.n812 4.5005
R25693 DVSS.n22475 DVSS.n812 4.5005
R25694 DVSS.n22489 DVSS.n812 4.5005
R25695 DVSS.n22474 DVSS.n812 4.5005
R25696 DVSS.n22490 DVSS.n812 4.5005
R25697 DVSS.n22473 DVSS.n812 4.5005
R25698 DVSS.n22500 DVSS.n812 4.5005
R25699 DVSS.n22502 DVSS.n812 4.5005
R25700 DVSS.n22504 DVSS.n812 4.5005
R25701 DVSS.n22478 DVSS.n822 4.5005
R25702 DVSS.n22483 DVSS.n822 4.5005
R25703 DVSS.n22477 DVSS.n822 4.5005
R25704 DVSS.n22485 DVSS.n822 4.5005
R25705 DVSS.n22476 DVSS.n822 4.5005
R25706 DVSS.n22487 DVSS.n822 4.5005
R25707 DVSS.n22475 DVSS.n822 4.5005
R25708 DVSS.n22489 DVSS.n822 4.5005
R25709 DVSS.n22474 DVSS.n822 4.5005
R25710 DVSS.n22490 DVSS.n822 4.5005
R25711 DVSS.n22473 DVSS.n822 4.5005
R25712 DVSS.n22500 DVSS.n822 4.5005
R25713 DVSS.n22502 DVSS.n822 4.5005
R25714 DVSS.n22472 DVSS.n822 4.5005
R25715 DVSS.n22504 DVSS.n822 4.5005
R25716 DVSS.n22478 DVSS.n811 4.5005
R25717 DVSS.n22483 DVSS.n811 4.5005
R25718 DVSS.n22477 DVSS.n811 4.5005
R25719 DVSS.n22485 DVSS.n811 4.5005
R25720 DVSS.n22476 DVSS.n811 4.5005
R25721 DVSS.n22487 DVSS.n811 4.5005
R25722 DVSS.n22475 DVSS.n811 4.5005
R25723 DVSS.n22489 DVSS.n811 4.5005
R25724 DVSS.n22474 DVSS.n811 4.5005
R25725 DVSS.n22490 DVSS.n811 4.5005
R25726 DVSS.n22473 DVSS.n811 4.5005
R25727 DVSS.n22500 DVSS.n811 4.5005
R25728 DVSS.n22502 DVSS.n811 4.5005
R25729 DVSS.n22504 DVSS.n811 4.5005
R25730 DVSS.n22478 DVSS.n823 4.5005
R25731 DVSS.n22483 DVSS.n823 4.5005
R25732 DVSS.n22477 DVSS.n823 4.5005
R25733 DVSS.n22485 DVSS.n823 4.5005
R25734 DVSS.n22476 DVSS.n823 4.5005
R25735 DVSS.n22487 DVSS.n823 4.5005
R25736 DVSS.n22475 DVSS.n823 4.5005
R25737 DVSS.n22489 DVSS.n823 4.5005
R25738 DVSS.n22474 DVSS.n823 4.5005
R25739 DVSS.n22490 DVSS.n823 4.5005
R25740 DVSS.n22473 DVSS.n823 4.5005
R25741 DVSS.n22500 DVSS.n823 4.5005
R25742 DVSS.n22502 DVSS.n823 4.5005
R25743 DVSS.n22504 DVSS.n823 4.5005
R25744 DVSS.n22478 DVSS.n810 4.5005
R25745 DVSS.n22483 DVSS.n810 4.5005
R25746 DVSS.n22477 DVSS.n810 4.5005
R25747 DVSS.n22485 DVSS.n810 4.5005
R25748 DVSS.n22476 DVSS.n810 4.5005
R25749 DVSS.n22487 DVSS.n810 4.5005
R25750 DVSS.n22475 DVSS.n810 4.5005
R25751 DVSS.n22489 DVSS.n810 4.5005
R25752 DVSS.n22474 DVSS.n810 4.5005
R25753 DVSS.n22490 DVSS.n810 4.5005
R25754 DVSS.n22473 DVSS.n810 4.5005
R25755 DVSS.n22500 DVSS.n810 4.5005
R25756 DVSS.n22502 DVSS.n810 4.5005
R25757 DVSS.n22472 DVSS.n810 4.5005
R25758 DVSS.n22504 DVSS.n810 4.5005
R25759 DVSS.n22478 DVSS.n831 4.5005
R25760 DVSS.n22483 DVSS.n831 4.5005
R25761 DVSS.n22477 DVSS.n831 4.5005
R25762 DVSS.n22485 DVSS.n831 4.5005
R25763 DVSS.n22476 DVSS.n831 4.5005
R25764 DVSS.n22487 DVSS.n831 4.5005
R25765 DVSS.n22475 DVSS.n831 4.5005
R25766 DVSS.n22489 DVSS.n831 4.5005
R25767 DVSS.n22474 DVSS.n831 4.5005
R25768 DVSS.n22490 DVSS.n831 4.5005
R25769 DVSS.n22473 DVSS.n831 4.5005
R25770 DVSS.n22500 DVSS.n831 4.5005
R25771 DVSS.n22498 DVSS.n831 4.5005
R25772 DVSS.n22502 DVSS.n831 4.5005
R25773 DVSS.n22504 DVSS.n831 4.5005
R25774 DVSS.n22478 DVSS.n809 4.5005
R25775 DVSS.n22483 DVSS.n809 4.5005
R25776 DVSS.n22477 DVSS.n809 4.5005
R25777 DVSS.n22485 DVSS.n809 4.5005
R25778 DVSS.n22476 DVSS.n809 4.5005
R25779 DVSS.n22487 DVSS.n809 4.5005
R25780 DVSS.n22475 DVSS.n809 4.5005
R25781 DVSS.n22489 DVSS.n809 4.5005
R25782 DVSS.n22474 DVSS.n809 4.5005
R25783 DVSS.n22490 DVSS.n809 4.5005
R25784 DVSS.n22473 DVSS.n809 4.5005
R25785 DVSS.n22500 DVSS.n809 4.5005
R25786 DVSS.n22502 DVSS.n809 4.5005
R25787 DVSS.n22504 DVSS.n809 4.5005
R25788 DVSS.n22478 DVSS.n832 4.5005
R25789 DVSS.n22483 DVSS.n832 4.5005
R25790 DVSS.n22477 DVSS.n832 4.5005
R25791 DVSS.n22485 DVSS.n832 4.5005
R25792 DVSS.n22476 DVSS.n832 4.5005
R25793 DVSS.n22487 DVSS.n832 4.5005
R25794 DVSS.n22475 DVSS.n832 4.5005
R25795 DVSS.n22489 DVSS.n832 4.5005
R25796 DVSS.n22474 DVSS.n832 4.5005
R25797 DVSS.n22490 DVSS.n832 4.5005
R25798 DVSS.n22473 DVSS.n832 4.5005
R25799 DVSS.n22500 DVSS.n832 4.5005
R25800 DVSS.n22502 DVSS.n832 4.5005
R25801 DVSS.n22504 DVSS.n832 4.5005
R25802 DVSS.n22478 DVSS.n808 4.5005
R25803 DVSS.n22483 DVSS.n808 4.5005
R25804 DVSS.n22477 DVSS.n808 4.5005
R25805 DVSS.n22485 DVSS.n808 4.5005
R25806 DVSS.n22476 DVSS.n808 4.5005
R25807 DVSS.n22487 DVSS.n808 4.5005
R25808 DVSS.n22475 DVSS.n808 4.5005
R25809 DVSS.n22489 DVSS.n808 4.5005
R25810 DVSS.n22474 DVSS.n808 4.5005
R25811 DVSS.n22490 DVSS.n808 4.5005
R25812 DVSS.n22473 DVSS.n808 4.5005
R25813 DVSS.n22500 DVSS.n808 4.5005
R25814 DVSS.n22498 DVSS.n808 4.5005
R25815 DVSS.n22502 DVSS.n808 4.5005
R25816 DVSS.n22504 DVSS.n808 4.5005
R25817 DVSS.n22478 DVSS.n840 4.5005
R25818 DVSS.n22483 DVSS.n840 4.5005
R25819 DVSS.n22477 DVSS.n840 4.5005
R25820 DVSS.n22485 DVSS.n840 4.5005
R25821 DVSS.n22476 DVSS.n840 4.5005
R25822 DVSS.n22487 DVSS.n840 4.5005
R25823 DVSS.n22475 DVSS.n840 4.5005
R25824 DVSS.n22489 DVSS.n840 4.5005
R25825 DVSS.n22474 DVSS.n840 4.5005
R25826 DVSS.n22490 DVSS.n840 4.5005
R25827 DVSS.n22473 DVSS.n840 4.5005
R25828 DVSS.n22500 DVSS.n840 4.5005
R25829 DVSS.n22498 DVSS.n840 4.5005
R25830 DVSS.n22502 DVSS.n840 4.5005
R25831 DVSS.n22504 DVSS.n840 4.5005
R25832 DVSS.n22478 DVSS.n807 4.5005
R25833 DVSS.n22483 DVSS.n807 4.5005
R25834 DVSS.n22477 DVSS.n807 4.5005
R25835 DVSS.n22485 DVSS.n807 4.5005
R25836 DVSS.n22476 DVSS.n807 4.5005
R25837 DVSS.n22487 DVSS.n807 4.5005
R25838 DVSS.n22475 DVSS.n807 4.5005
R25839 DVSS.n22489 DVSS.n807 4.5005
R25840 DVSS.n22474 DVSS.n807 4.5005
R25841 DVSS.n22490 DVSS.n807 4.5005
R25842 DVSS.n22473 DVSS.n807 4.5005
R25843 DVSS.n22500 DVSS.n807 4.5005
R25844 DVSS.n22502 DVSS.n807 4.5005
R25845 DVSS.n22504 DVSS.n807 4.5005
R25846 DVSS.n22478 DVSS.n841 4.5005
R25847 DVSS.n22483 DVSS.n841 4.5005
R25848 DVSS.n22477 DVSS.n841 4.5005
R25849 DVSS.n22485 DVSS.n841 4.5005
R25850 DVSS.n22476 DVSS.n841 4.5005
R25851 DVSS.n22487 DVSS.n841 4.5005
R25852 DVSS.n22475 DVSS.n841 4.5005
R25853 DVSS.n22489 DVSS.n841 4.5005
R25854 DVSS.n22474 DVSS.n841 4.5005
R25855 DVSS.n22490 DVSS.n841 4.5005
R25856 DVSS.n22473 DVSS.n841 4.5005
R25857 DVSS.n22500 DVSS.n841 4.5005
R25858 DVSS.n22502 DVSS.n841 4.5005
R25859 DVSS.n22504 DVSS.n841 4.5005
R25860 DVSS.n22478 DVSS.n806 4.5005
R25861 DVSS.n22483 DVSS.n806 4.5005
R25862 DVSS.n22477 DVSS.n806 4.5005
R25863 DVSS.n22485 DVSS.n806 4.5005
R25864 DVSS.n22476 DVSS.n806 4.5005
R25865 DVSS.n22487 DVSS.n806 4.5005
R25866 DVSS.n22475 DVSS.n806 4.5005
R25867 DVSS.n22489 DVSS.n806 4.5005
R25868 DVSS.n22474 DVSS.n806 4.5005
R25869 DVSS.n22490 DVSS.n806 4.5005
R25870 DVSS.n22473 DVSS.n806 4.5005
R25871 DVSS.n22500 DVSS.n806 4.5005
R25872 DVSS.n22498 DVSS.n806 4.5005
R25873 DVSS.n22502 DVSS.n806 4.5005
R25874 DVSS.n22504 DVSS.n806 4.5005
R25875 DVSS.n22478 DVSS.n849 4.5005
R25876 DVSS.n22483 DVSS.n849 4.5005
R25877 DVSS.n22477 DVSS.n849 4.5005
R25878 DVSS.n22485 DVSS.n849 4.5005
R25879 DVSS.n22476 DVSS.n849 4.5005
R25880 DVSS.n22487 DVSS.n849 4.5005
R25881 DVSS.n22475 DVSS.n849 4.5005
R25882 DVSS.n22489 DVSS.n849 4.5005
R25883 DVSS.n22474 DVSS.n849 4.5005
R25884 DVSS.n22490 DVSS.n849 4.5005
R25885 DVSS.n22473 DVSS.n849 4.5005
R25886 DVSS.n22500 DVSS.n849 4.5005
R25887 DVSS.n22498 DVSS.n849 4.5005
R25888 DVSS.n22502 DVSS.n849 4.5005
R25889 DVSS.n22504 DVSS.n849 4.5005
R25890 DVSS.n22478 DVSS.n805 4.5005
R25891 DVSS.n22483 DVSS.n805 4.5005
R25892 DVSS.n22477 DVSS.n805 4.5005
R25893 DVSS.n22485 DVSS.n805 4.5005
R25894 DVSS.n22476 DVSS.n805 4.5005
R25895 DVSS.n22487 DVSS.n805 4.5005
R25896 DVSS.n22475 DVSS.n805 4.5005
R25897 DVSS.n22489 DVSS.n805 4.5005
R25898 DVSS.n22474 DVSS.n805 4.5005
R25899 DVSS.n22490 DVSS.n805 4.5005
R25900 DVSS.n22473 DVSS.n805 4.5005
R25901 DVSS.n22500 DVSS.n805 4.5005
R25902 DVSS.n22502 DVSS.n805 4.5005
R25903 DVSS.n22504 DVSS.n805 4.5005
R25904 DVSS.n22478 DVSS.n850 4.5005
R25905 DVSS.n22483 DVSS.n850 4.5005
R25906 DVSS.n22477 DVSS.n850 4.5005
R25907 DVSS.n22485 DVSS.n850 4.5005
R25908 DVSS.n22476 DVSS.n850 4.5005
R25909 DVSS.n22487 DVSS.n850 4.5005
R25910 DVSS.n22475 DVSS.n850 4.5005
R25911 DVSS.n22489 DVSS.n850 4.5005
R25912 DVSS.n22474 DVSS.n850 4.5005
R25913 DVSS.n22490 DVSS.n850 4.5005
R25914 DVSS.n22473 DVSS.n850 4.5005
R25915 DVSS.n22500 DVSS.n850 4.5005
R25916 DVSS.n22502 DVSS.n850 4.5005
R25917 DVSS.n22504 DVSS.n850 4.5005
R25918 DVSS.n22478 DVSS.n804 4.5005
R25919 DVSS.n22483 DVSS.n804 4.5005
R25920 DVSS.n22477 DVSS.n804 4.5005
R25921 DVSS.n22485 DVSS.n804 4.5005
R25922 DVSS.n22476 DVSS.n804 4.5005
R25923 DVSS.n22487 DVSS.n804 4.5005
R25924 DVSS.n22475 DVSS.n804 4.5005
R25925 DVSS.n22489 DVSS.n804 4.5005
R25926 DVSS.n22474 DVSS.n804 4.5005
R25927 DVSS.n22490 DVSS.n804 4.5005
R25928 DVSS.n22473 DVSS.n804 4.5005
R25929 DVSS.n22500 DVSS.n804 4.5005
R25930 DVSS.n22498 DVSS.n804 4.5005
R25931 DVSS.n22502 DVSS.n804 4.5005
R25932 DVSS.n22504 DVSS.n804 4.5005
R25933 DVSS.n22478 DVSS.n857 4.5005
R25934 DVSS.n22483 DVSS.n857 4.5005
R25935 DVSS.n22477 DVSS.n857 4.5005
R25936 DVSS.n22485 DVSS.n857 4.5005
R25937 DVSS.n22476 DVSS.n857 4.5005
R25938 DVSS.n22487 DVSS.n857 4.5005
R25939 DVSS.n22475 DVSS.n857 4.5005
R25940 DVSS.n22489 DVSS.n857 4.5005
R25941 DVSS.n22474 DVSS.n857 4.5005
R25942 DVSS.n22490 DVSS.n857 4.5005
R25943 DVSS.n22473 DVSS.n857 4.5005
R25944 DVSS.n22500 DVSS.n857 4.5005
R25945 DVSS.n22498 DVSS.n857 4.5005
R25946 DVSS.n22502 DVSS.n857 4.5005
R25947 DVSS.n22504 DVSS.n857 4.5005
R25948 DVSS.n22478 DVSS.n803 4.5005
R25949 DVSS.n22483 DVSS.n803 4.5005
R25950 DVSS.n22477 DVSS.n803 4.5005
R25951 DVSS.n22485 DVSS.n803 4.5005
R25952 DVSS.n22476 DVSS.n803 4.5005
R25953 DVSS.n22487 DVSS.n803 4.5005
R25954 DVSS.n22475 DVSS.n803 4.5005
R25955 DVSS.n22489 DVSS.n803 4.5005
R25956 DVSS.n22474 DVSS.n803 4.5005
R25957 DVSS.n22490 DVSS.n803 4.5005
R25958 DVSS.n22473 DVSS.n803 4.5005
R25959 DVSS.n22500 DVSS.n803 4.5005
R25960 DVSS.n22502 DVSS.n803 4.5005
R25961 DVSS.n22504 DVSS.n803 4.5005
R25962 DVSS.n22478 DVSS.n22461 4.5005
R25963 DVSS.n22483 DVSS.n22461 4.5005
R25964 DVSS.n22477 DVSS.n22461 4.5005
R25965 DVSS.n22485 DVSS.n22461 4.5005
R25966 DVSS.n22476 DVSS.n22461 4.5005
R25967 DVSS.n22487 DVSS.n22461 4.5005
R25968 DVSS.n22475 DVSS.n22461 4.5005
R25969 DVSS.n22489 DVSS.n22461 4.5005
R25970 DVSS.n22474 DVSS.n22461 4.5005
R25971 DVSS.n22490 DVSS.n22461 4.5005
R25972 DVSS.n22473 DVSS.n22461 4.5005
R25973 DVSS.n22500 DVSS.n22461 4.5005
R25974 DVSS.n22502 DVSS.n22461 4.5005
R25975 DVSS.n22472 DVSS.n22461 4.5005
R25976 DVSS.n22504 DVSS.n22461 4.5005
R25977 DVSS.n22478 DVSS.n802 4.5005
R25978 DVSS.n22483 DVSS.n802 4.5005
R25979 DVSS.n22477 DVSS.n802 4.5005
R25980 DVSS.n22485 DVSS.n802 4.5005
R25981 DVSS.n22476 DVSS.n802 4.5005
R25982 DVSS.n22487 DVSS.n802 4.5005
R25983 DVSS.n22475 DVSS.n802 4.5005
R25984 DVSS.n22489 DVSS.n802 4.5005
R25985 DVSS.n22474 DVSS.n802 4.5005
R25986 DVSS.n22490 DVSS.n802 4.5005
R25987 DVSS.n22473 DVSS.n802 4.5005
R25988 DVSS.n22500 DVSS.n802 4.5005
R25989 DVSS.n22502 DVSS.n802 4.5005
R25990 DVSS.n22472 DVSS.n802 4.5005
R25991 DVSS.n22504 DVSS.n802 4.5005
R25992 DVSS.n22503 DVSS.n22478 4.5005
R25993 DVSS.n22503 DVSS.n22483 4.5005
R25994 DVSS.n22503 DVSS.n22477 4.5005
R25995 DVSS.n22503 DVSS.n22485 4.5005
R25996 DVSS.n22503 DVSS.n22476 4.5005
R25997 DVSS.n22503 DVSS.n22487 4.5005
R25998 DVSS.n22503 DVSS.n22475 4.5005
R25999 DVSS.n22503 DVSS.n22489 4.5005
R26000 DVSS.n22503 DVSS.n22474 4.5005
R26001 DVSS.n22503 DVSS.n22490 4.5005
R26002 DVSS.n22503 DVSS.n22473 4.5005
R26003 DVSS.n22503 DVSS.n22500 4.5005
R26004 DVSS.n22503 DVSS.n22502 4.5005
R26005 DVSS.n22503 DVSS.n22472 4.5005
R26006 DVSS.n22504 DVSS.n22503 4.5005
R26007 DVSS.n245 DVSS.n217 4.5005
R26008 DVSS.n247 DVSS.n217 4.5005
R26009 DVSS.n244 DVSS.n217 4.5005
R26010 DVSS.n250 DVSS.n217 4.5005
R26011 DVSS.n242 DVSS.n217 4.5005
R26012 DVSS.n251 DVSS.n217 4.5005
R26013 DVSS.n241 DVSS.n217 4.5005
R26014 DVSS.n252 DVSS.n217 4.5005
R26015 DVSS.n240 DVSS.n217 4.5005
R26016 DVSS.n23093 DVSS.n217 4.5005
R26017 DVSS.n239 DVSS.n217 4.5005
R26018 DVSS.n23095 DVSS.n217 4.5005
R26019 DVSS.n245 DVSS.n218 4.5005
R26020 DVSS.n247 DVSS.n218 4.5005
R26021 DVSS.n244 DVSS.n218 4.5005
R26022 DVSS.n249 DVSS.n218 4.5005
R26023 DVSS.n243 DVSS.n218 4.5005
R26024 DVSS.n250 DVSS.n218 4.5005
R26025 DVSS.n242 DVSS.n218 4.5005
R26026 DVSS.n251 DVSS.n218 4.5005
R26027 DVSS.n241 DVSS.n218 4.5005
R26028 DVSS.n252 DVSS.n218 4.5005
R26029 DVSS.n240 DVSS.n218 4.5005
R26030 DVSS.n253 DVSS.n218 4.5005
R26031 DVSS.n23093 DVSS.n218 4.5005
R26032 DVSS.n23095 DVSS.n218 4.5005
R26033 DVSS.n245 DVSS.n216 4.5005
R26034 DVSS.n247 DVSS.n216 4.5005
R26035 DVSS.n244 DVSS.n216 4.5005
R26036 DVSS.n249 DVSS.n216 4.5005
R26037 DVSS.n243 DVSS.n216 4.5005
R26038 DVSS.n250 DVSS.n216 4.5005
R26039 DVSS.n242 DVSS.n216 4.5005
R26040 DVSS.n251 DVSS.n216 4.5005
R26041 DVSS.n241 DVSS.n216 4.5005
R26042 DVSS.n252 DVSS.n216 4.5005
R26043 DVSS.n240 DVSS.n216 4.5005
R26044 DVSS.n253 DVSS.n216 4.5005
R26045 DVSS.n23093 DVSS.n216 4.5005
R26046 DVSS.n23095 DVSS.n216 4.5005
R26047 DVSS.n245 DVSS.n219 4.5005
R26048 DVSS.n247 DVSS.n219 4.5005
R26049 DVSS.n244 DVSS.n219 4.5005
R26050 DVSS.n249 DVSS.n219 4.5005
R26051 DVSS.n243 DVSS.n219 4.5005
R26052 DVSS.n250 DVSS.n219 4.5005
R26053 DVSS.n242 DVSS.n219 4.5005
R26054 DVSS.n251 DVSS.n219 4.5005
R26055 DVSS.n241 DVSS.n219 4.5005
R26056 DVSS.n252 DVSS.n219 4.5005
R26057 DVSS.n240 DVSS.n219 4.5005
R26058 DVSS.n253 DVSS.n219 4.5005
R26059 DVSS.n23093 DVSS.n219 4.5005
R26060 DVSS.n239 DVSS.n219 4.5005
R26061 DVSS.n23095 DVSS.n219 4.5005
R26062 DVSS.n245 DVSS.n215 4.5005
R26063 DVSS.n247 DVSS.n215 4.5005
R26064 DVSS.n244 DVSS.n215 4.5005
R26065 DVSS.n249 DVSS.n215 4.5005
R26066 DVSS.n243 DVSS.n215 4.5005
R26067 DVSS.n250 DVSS.n215 4.5005
R26068 DVSS.n242 DVSS.n215 4.5005
R26069 DVSS.n251 DVSS.n215 4.5005
R26070 DVSS.n241 DVSS.n215 4.5005
R26071 DVSS.n252 DVSS.n215 4.5005
R26072 DVSS.n240 DVSS.n215 4.5005
R26073 DVSS.n253 DVSS.n215 4.5005
R26074 DVSS.n23093 DVSS.n215 4.5005
R26075 DVSS.n23095 DVSS.n215 4.5005
R26076 DVSS.n245 DVSS.n220 4.5005
R26077 DVSS.n247 DVSS.n220 4.5005
R26078 DVSS.n244 DVSS.n220 4.5005
R26079 DVSS.n249 DVSS.n220 4.5005
R26080 DVSS.n243 DVSS.n220 4.5005
R26081 DVSS.n250 DVSS.n220 4.5005
R26082 DVSS.n242 DVSS.n220 4.5005
R26083 DVSS.n251 DVSS.n220 4.5005
R26084 DVSS.n241 DVSS.n220 4.5005
R26085 DVSS.n252 DVSS.n220 4.5005
R26086 DVSS.n240 DVSS.n220 4.5005
R26087 DVSS.n253 DVSS.n220 4.5005
R26088 DVSS.n23093 DVSS.n220 4.5005
R26089 DVSS.n23095 DVSS.n220 4.5005
R26090 DVSS.n245 DVSS.n214 4.5005
R26091 DVSS.n247 DVSS.n214 4.5005
R26092 DVSS.n244 DVSS.n214 4.5005
R26093 DVSS.n249 DVSS.n214 4.5005
R26094 DVSS.n243 DVSS.n214 4.5005
R26095 DVSS.n250 DVSS.n214 4.5005
R26096 DVSS.n242 DVSS.n214 4.5005
R26097 DVSS.n251 DVSS.n214 4.5005
R26098 DVSS.n241 DVSS.n214 4.5005
R26099 DVSS.n252 DVSS.n214 4.5005
R26100 DVSS.n240 DVSS.n214 4.5005
R26101 DVSS.n253 DVSS.n214 4.5005
R26102 DVSS.n23093 DVSS.n214 4.5005
R26103 DVSS.n239 DVSS.n214 4.5005
R26104 DVSS.n23095 DVSS.n214 4.5005
R26105 DVSS.n245 DVSS.n221 4.5005
R26106 DVSS.n247 DVSS.n221 4.5005
R26107 DVSS.n244 DVSS.n221 4.5005
R26108 DVSS.n249 DVSS.n221 4.5005
R26109 DVSS.n243 DVSS.n221 4.5005
R26110 DVSS.n250 DVSS.n221 4.5005
R26111 DVSS.n242 DVSS.n221 4.5005
R26112 DVSS.n251 DVSS.n221 4.5005
R26113 DVSS.n241 DVSS.n221 4.5005
R26114 DVSS.n252 DVSS.n221 4.5005
R26115 DVSS.n240 DVSS.n221 4.5005
R26116 DVSS.n253 DVSS.n221 4.5005
R26117 DVSS.n262 DVSS.n221 4.5005
R26118 DVSS.n23093 DVSS.n221 4.5005
R26119 DVSS.n23095 DVSS.n221 4.5005
R26120 DVSS.n245 DVSS.n213 4.5005
R26121 DVSS.n247 DVSS.n213 4.5005
R26122 DVSS.n244 DVSS.n213 4.5005
R26123 DVSS.n249 DVSS.n213 4.5005
R26124 DVSS.n243 DVSS.n213 4.5005
R26125 DVSS.n250 DVSS.n213 4.5005
R26126 DVSS.n242 DVSS.n213 4.5005
R26127 DVSS.n251 DVSS.n213 4.5005
R26128 DVSS.n241 DVSS.n213 4.5005
R26129 DVSS.n252 DVSS.n213 4.5005
R26130 DVSS.n240 DVSS.n213 4.5005
R26131 DVSS.n253 DVSS.n213 4.5005
R26132 DVSS.n23093 DVSS.n213 4.5005
R26133 DVSS.n23095 DVSS.n213 4.5005
R26134 DVSS.n245 DVSS.n222 4.5005
R26135 DVSS.n247 DVSS.n222 4.5005
R26136 DVSS.n244 DVSS.n222 4.5005
R26137 DVSS.n249 DVSS.n222 4.5005
R26138 DVSS.n243 DVSS.n222 4.5005
R26139 DVSS.n250 DVSS.n222 4.5005
R26140 DVSS.n242 DVSS.n222 4.5005
R26141 DVSS.n251 DVSS.n222 4.5005
R26142 DVSS.n241 DVSS.n222 4.5005
R26143 DVSS.n252 DVSS.n222 4.5005
R26144 DVSS.n240 DVSS.n222 4.5005
R26145 DVSS.n253 DVSS.n222 4.5005
R26146 DVSS.n23093 DVSS.n222 4.5005
R26147 DVSS.n23095 DVSS.n222 4.5005
R26148 DVSS.n245 DVSS.n212 4.5005
R26149 DVSS.n247 DVSS.n212 4.5005
R26150 DVSS.n244 DVSS.n212 4.5005
R26151 DVSS.n249 DVSS.n212 4.5005
R26152 DVSS.n243 DVSS.n212 4.5005
R26153 DVSS.n250 DVSS.n212 4.5005
R26154 DVSS.n242 DVSS.n212 4.5005
R26155 DVSS.n251 DVSS.n212 4.5005
R26156 DVSS.n241 DVSS.n212 4.5005
R26157 DVSS.n252 DVSS.n212 4.5005
R26158 DVSS.n240 DVSS.n212 4.5005
R26159 DVSS.n253 DVSS.n212 4.5005
R26160 DVSS.n262 DVSS.n212 4.5005
R26161 DVSS.n23093 DVSS.n212 4.5005
R26162 DVSS.n23095 DVSS.n212 4.5005
R26163 DVSS.n245 DVSS.n223 4.5005
R26164 DVSS.n247 DVSS.n223 4.5005
R26165 DVSS.n244 DVSS.n223 4.5005
R26166 DVSS.n249 DVSS.n223 4.5005
R26167 DVSS.n243 DVSS.n223 4.5005
R26168 DVSS.n250 DVSS.n223 4.5005
R26169 DVSS.n242 DVSS.n223 4.5005
R26170 DVSS.n251 DVSS.n223 4.5005
R26171 DVSS.n241 DVSS.n223 4.5005
R26172 DVSS.n252 DVSS.n223 4.5005
R26173 DVSS.n240 DVSS.n223 4.5005
R26174 DVSS.n253 DVSS.n223 4.5005
R26175 DVSS.n262 DVSS.n223 4.5005
R26176 DVSS.n23093 DVSS.n223 4.5005
R26177 DVSS.n23095 DVSS.n223 4.5005
R26178 DVSS.n245 DVSS.n211 4.5005
R26179 DVSS.n247 DVSS.n211 4.5005
R26180 DVSS.n244 DVSS.n211 4.5005
R26181 DVSS.n249 DVSS.n211 4.5005
R26182 DVSS.n243 DVSS.n211 4.5005
R26183 DVSS.n250 DVSS.n211 4.5005
R26184 DVSS.n242 DVSS.n211 4.5005
R26185 DVSS.n251 DVSS.n211 4.5005
R26186 DVSS.n241 DVSS.n211 4.5005
R26187 DVSS.n252 DVSS.n211 4.5005
R26188 DVSS.n240 DVSS.n211 4.5005
R26189 DVSS.n253 DVSS.n211 4.5005
R26190 DVSS.n23093 DVSS.n211 4.5005
R26191 DVSS.n23095 DVSS.n211 4.5005
R26192 DVSS.n245 DVSS.n224 4.5005
R26193 DVSS.n247 DVSS.n224 4.5005
R26194 DVSS.n244 DVSS.n224 4.5005
R26195 DVSS.n249 DVSS.n224 4.5005
R26196 DVSS.n243 DVSS.n224 4.5005
R26197 DVSS.n250 DVSS.n224 4.5005
R26198 DVSS.n242 DVSS.n224 4.5005
R26199 DVSS.n251 DVSS.n224 4.5005
R26200 DVSS.n241 DVSS.n224 4.5005
R26201 DVSS.n252 DVSS.n224 4.5005
R26202 DVSS.n240 DVSS.n224 4.5005
R26203 DVSS.n253 DVSS.n224 4.5005
R26204 DVSS.n23093 DVSS.n224 4.5005
R26205 DVSS.n23095 DVSS.n224 4.5005
R26206 DVSS.n245 DVSS.n210 4.5005
R26207 DVSS.n247 DVSS.n210 4.5005
R26208 DVSS.n244 DVSS.n210 4.5005
R26209 DVSS.n249 DVSS.n210 4.5005
R26210 DVSS.n243 DVSS.n210 4.5005
R26211 DVSS.n250 DVSS.n210 4.5005
R26212 DVSS.n242 DVSS.n210 4.5005
R26213 DVSS.n251 DVSS.n210 4.5005
R26214 DVSS.n241 DVSS.n210 4.5005
R26215 DVSS.n252 DVSS.n210 4.5005
R26216 DVSS.n240 DVSS.n210 4.5005
R26217 DVSS.n253 DVSS.n210 4.5005
R26218 DVSS.n262 DVSS.n210 4.5005
R26219 DVSS.n23093 DVSS.n210 4.5005
R26220 DVSS.n23095 DVSS.n210 4.5005
R26221 DVSS.n245 DVSS.n225 4.5005
R26222 DVSS.n247 DVSS.n225 4.5005
R26223 DVSS.n244 DVSS.n225 4.5005
R26224 DVSS.n249 DVSS.n225 4.5005
R26225 DVSS.n243 DVSS.n225 4.5005
R26226 DVSS.n250 DVSS.n225 4.5005
R26227 DVSS.n242 DVSS.n225 4.5005
R26228 DVSS.n251 DVSS.n225 4.5005
R26229 DVSS.n241 DVSS.n225 4.5005
R26230 DVSS.n252 DVSS.n225 4.5005
R26231 DVSS.n240 DVSS.n225 4.5005
R26232 DVSS.n253 DVSS.n225 4.5005
R26233 DVSS.n262 DVSS.n225 4.5005
R26234 DVSS.n23093 DVSS.n225 4.5005
R26235 DVSS.n23095 DVSS.n225 4.5005
R26236 DVSS.n245 DVSS.n209 4.5005
R26237 DVSS.n247 DVSS.n209 4.5005
R26238 DVSS.n244 DVSS.n209 4.5005
R26239 DVSS.n249 DVSS.n209 4.5005
R26240 DVSS.n243 DVSS.n209 4.5005
R26241 DVSS.n250 DVSS.n209 4.5005
R26242 DVSS.n242 DVSS.n209 4.5005
R26243 DVSS.n251 DVSS.n209 4.5005
R26244 DVSS.n241 DVSS.n209 4.5005
R26245 DVSS.n252 DVSS.n209 4.5005
R26246 DVSS.n240 DVSS.n209 4.5005
R26247 DVSS.n253 DVSS.n209 4.5005
R26248 DVSS.n23093 DVSS.n209 4.5005
R26249 DVSS.n23095 DVSS.n209 4.5005
R26250 DVSS.n245 DVSS.n226 4.5005
R26251 DVSS.n247 DVSS.n226 4.5005
R26252 DVSS.n244 DVSS.n226 4.5005
R26253 DVSS.n249 DVSS.n226 4.5005
R26254 DVSS.n243 DVSS.n226 4.5005
R26255 DVSS.n250 DVSS.n226 4.5005
R26256 DVSS.n242 DVSS.n226 4.5005
R26257 DVSS.n251 DVSS.n226 4.5005
R26258 DVSS.n241 DVSS.n226 4.5005
R26259 DVSS.n252 DVSS.n226 4.5005
R26260 DVSS.n240 DVSS.n226 4.5005
R26261 DVSS.n253 DVSS.n226 4.5005
R26262 DVSS.n23093 DVSS.n226 4.5005
R26263 DVSS.n23095 DVSS.n226 4.5005
R26264 DVSS.n245 DVSS.n208 4.5005
R26265 DVSS.n247 DVSS.n208 4.5005
R26266 DVSS.n244 DVSS.n208 4.5005
R26267 DVSS.n249 DVSS.n208 4.5005
R26268 DVSS.n243 DVSS.n208 4.5005
R26269 DVSS.n250 DVSS.n208 4.5005
R26270 DVSS.n242 DVSS.n208 4.5005
R26271 DVSS.n251 DVSS.n208 4.5005
R26272 DVSS.n241 DVSS.n208 4.5005
R26273 DVSS.n252 DVSS.n208 4.5005
R26274 DVSS.n240 DVSS.n208 4.5005
R26275 DVSS.n253 DVSS.n208 4.5005
R26276 DVSS.n262 DVSS.n208 4.5005
R26277 DVSS.n23093 DVSS.n208 4.5005
R26278 DVSS.n23095 DVSS.n208 4.5005
R26279 DVSS.n245 DVSS.n227 4.5005
R26280 DVSS.n247 DVSS.n227 4.5005
R26281 DVSS.n244 DVSS.n227 4.5005
R26282 DVSS.n249 DVSS.n227 4.5005
R26283 DVSS.n243 DVSS.n227 4.5005
R26284 DVSS.n250 DVSS.n227 4.5005
R26285 DVSS.n242 DVSS.n227 4.5005
R26286 DVSS.n251 DVSS.n227 4.5005
R26287 DVSS.n241 DVSS.n227 4.5005
R26288 DVSS.n252 DVSS.n227 4.5005
R26289 DVSS.n240 DVSS.n227 4.5005
R26290 DVSS.n253 DVSS.n227 4.5005
R26291 DVSS.n262 DVSS.n227 4.5005
R26292 DVSS.n23093 DVSS.n227 4.5005
R26293 DVSS.n23095 DVSS.n227 4.5005
R26294 DVSS.n245 DVSS.n207 4.5005
R26295 DVSS.n247 DVSS.n207 4.5005
R26296 DVSS.n244 DVSS.n207 4.5005
R26297 DVSS.n249 DVSS.n207 4.5005
R26298 DVSS.n243 DVSS.n207 4.5005
R26299 DVSS.n250 DVSS.n207 4.5005
R26300 DVSS.n242 DVSS.n207 4.5005
R26301 DVSS.n251 DVSS.n207 4.5005
R26302 DVSS.n241 DVSS.n207 4.5005
R26303 DVSS.n252 DVSS.n207 4.5005
R26304 DVSS.n240 DVSS.n207 4.5005
R26305 DVSS.n253 DVSS.n207 4.5005
R26306 DVSS.n23093 DVSS.n207 4.5005
R26307 DVSS.n23095 DVSS.n207 4.5005
R26308 DVSS.n245 DVSS.n228 4.5005
R26309 DVSS.n247 DVSS.n228 4.5005
R26310 DVSS.n244 DVSS.n228 4.5005
R26311 DVSS.n249 DVSS.n228 4.5005
R26312 DVSS.n243 DVSS.n228 4.5005
R26313 DVSS.n250 DVSS.n228 4.5005
R26314 DVSS.n242 DVSS.n228 4.5005
R26315 DVSS.n251 DVSS.n228 4.5005
R26316 DVSS.n241 DVSS.n228 4.5005
R26317 DVSS.n252 DVSS.n228 4.5005
R26318 DVSS.n240 DVSS.n228 4.5005
R26319 DVSS.n253 DVSS.n228 4.5005
R26320 DVSS.n23093 DVSS.n228 4.5005
R26321 DVSS.n239 DVSS.n228 4.5005
R26322 DVSS.n23095 DVSS.n228 4.5005
R26323 DVSS.n245 DVSS.n206 4.5005
R26324 DVSS.n247 DVSS.n206 4.5005
R26325 DVSS.n244 DVSS.n206 4.5005
R26326 DVSS.n249 DVSS.n206 4.5005
R26327 DVSS.n243 DVSS.n206 4.5005
R26328 DVSS.n250 DVSS.n206 4.5005
R26329 DVSS.n242 DVSS.n206 4.5005
R26330 DVSS.n251 DVSS.n206 4.5005
R26331 DVSS.n241 DVSS.n206 4.5005
R26332 DVSS.n252 DVSS.n206 4.5005
R26333 DVSS.n240 DVSS.n206 4.5005
R26334 DVSS.n253 DVSS.n206 4.5005
R26335 DVSS.n23093 DVSS.n206 4.5005
R26336 DVSS.n239 DVSS.n206 4.5005
R26337 DVSS.n23095 DVSS.n206 4.5005
R26338 DVSS.n23094 DVSS.n245 4.5005
R26339 DVSS.n23094 DVSS.n247 4.5005
R26340 DVSS.n23094 DVSS.n244 4.5005
R26341 DVSS.n23094 DVSS.n249 4.5005
R26342 DVSS.n23094 DVSS.n243 4.5005
R26343 DVSS.n23094 DVSS.n250 4.5005
R26344 DVSS.n23094 DVSS.n242 4.5005
R26345 DVSS.n23094 DVSS.n251 4.5005
R26346 DVSS.n23094 DVSS.n241 4.5005
R26347 DVSS.n23094 DVSS.n252 4.5005
R26348 DVSS.n23094 DVSS.n240 4.5005
R26349 DVSS.n23094 DVSS.n253 4.5005
R26350 DVSS.n23094 DVSS.n23093 4.5005
R26351 DVSS.n23094 DVSS.n239 4.5005
R26352 DVSS.n23095 DVSS.n23094 4.5005
R26353 DVSS.n165 DVSS.n137 4.5005
R26354 DVSS.n167 DVSS.n137 4.5005
R26355 DVSS.n164 DVSS.n137 4.5005
R26356 DVSS.n170 DVSS.n137 4.5005
R26357 DVSS.n162 DVSS.n137 4.5005
R26358 DVSS.n171 DVSS.n137 4.5005
R26359 DVSS.n161 DVSS.n137 4.5005
R26360 DVSS.n172 DVSS.n137 4.5005
R26361 DVSS.n160 DVSS.n137 4.5005
R26362 DVSS.n23136 DVSS.n137 4.5005
R26363 DVSS.n159 DVSS.n137 4.5005
R26364 DVSS.n23138 DVSS.n137 4.5005
R26365 DVSS.n165 DVSS.n138 4.5005
R26366 DVSS.n167 DVSS.n138 4.5005
R26367 DVSS.n164 DVSS.n138 4.5005
R26368 DVSS.n169 DVSS.n138 4.5005
R26369 DVSS.n163 DVSS.n138 4.5005
R26370 DVSS.n170 DVSS.n138 4.5005
R26371 DVSS.n162 DVSS.n138 4.5005
R26372 DVSS.n171 DVSS.n138 4.5005
R26373 DVSS.n161 DVSS.n138 4.5005
R26374 DVSS.n172 DVSS.n138 4.5005
R26375 DVSS.n160 DVSS.n138 4.5005
R26376 DVSS.n173 DVSS.n138 4.5005
R26377 DVSS.n23136 DVSS.n138 4.5005
R26378 DVSS.n23138 DVSS.n138 4.5005
R26379 DVSS.n165 DVSS.n136 4.5005
R26380 DVSS.n167 DVSS.n136 4.5005
R26381 DVSS.n164 DVSS.n136 4.5005
R26382 DVSS.n169 DVSS.n136 4.5005
R26383 DVSS.n163 DVSS.n136 4.5005
R26384 DVSS.n170 DVSS.n136 4.5005
R26385 DVSS.n162 DVSS.n136 4.5005
R26386 DVSS.n171 DVSS.n136 4.5005
R26387 DVSS.n161 DVSS.n136 4.5005
R26388 DVSS.n172 DVSS.n136 4.5005
R26389 DVSS.n160 DVSS.n136 4.5005
R26390 DVSS.n173 DVSS.n136 4.5005
R26391 DVSS.n23136 DVSS.n136 4.5005
R26392 DVSS.n23138 DVSS.n136 4.5005
R26393 DVSS.n165 DVSS.n139 4.5005
R26394 DVSS.n167 DVSS.n139 4.5005
R26395 DVSS.n164 DVSS.n139 4.5005
R26396 DVSS.n169 DVSS.n139 4.5005
R26397 DVSS.n163 DVSS.n139 4.5005
R26398 DVSS.n170 DVSS.n139 4.5005
R26399 DVSS.n162 DVSS.n139 4.5005
R26400 DVSS.n171 DVSS.n139 4.5005
R26401 DVSS.n161 DVSS.n139 4.5005
R26402 DVSS.n172 DVSS.n139 4.5005
R26403 DVSS.n160 DVSS.n139 4.5005
R26404 DVSS.n173 DVSS.n139 4.5005
R26405 DVSS.n23136 DVSS.n139 4.5005
R26406 DVSS.n159 DVSS.n139 4.5005
R26407 DVSS.n23138 DVSS.n139 4.5005
R26408 DVSS.n165 DVSS.n135 4.5005
R26409 DVSS.n167 DVSS.n135 4.5005
R26410 DVSS.n164 DVSS.n135 4.5005
R26411 DVSS.n169 DVSS.n135 4.5005
R26412 DVSS.n163 DVSS.n135 4.5005
R26413 DVSS.n170 DVSS.n135 4.5005
R26414 DVSS.n162 DVSS.n135 4.5005
R26415 DVSS.n171 DVSS.n135 4.5005
R26416 DVSS.n161 DVSS.n135 4.5005
R26417 DVSS.n172 DVSS.n135 4.5005
R26418 DVSS.n160 DVSS.n135 4.5005
R26419 DVSS.n173 DVSS.n135 4.5005
R26420 DVSS.n23136 DVSS.n135 4.5005
R26421 DVSS.n23138 DVSS.n135 4.5005
R26422 DVSS.n165 DVSS.n140 4.5005
R26423 DVSS.n167 DVSS.n140 4.5005
R26424 DVSS.n164 DVSS.n140 4.5005
R26425 DVSS.n169 DVSS.n140 4.5005
R26426 DVSS.n163 DVSS.n140 4.5005
R26427 DVSS.n170 DVSS.n140 4.5005
R26428 DVSS.n162 DVSS.n140 4.5005
R26429 DVSS.n171 DVSS.n140 4.5005
R26430 DVSS.n161 DVSS.n140 4.5005
R26431 DVSS.n172 DVSS.n140 4.5005
R26432 DVSS.n160 DVSS.n140 4.5005
R26433 DVSS.n173 DVSS.n140 4.5005
R26434 DVSS.n23136 DVSS.n140 4.5005
R26435 DVSS.n23138 DVSS.n140 4.5005
R26436 DVSS.n165 DVSS.n134 4.5005
R26437 DVSS.n167 DVSS.n134 4.5005
R26438 DVSS.n164 DVSS.n134 4.5005
R26439 DVSS.n169 DVSS.n134 4.5005
R26440 DVSS.n163 DVSS.n134 4.5005
R26441 DVSS.n170 DVSS.n134 4.5005
R26442 DVSS.n162 DVSS.n134 4.5005
R26443 DVSS.n171 DVSS.n134 4.5005
R26444 DVSS.n161 DVSS.n134 4.5005
R26445 DVSS.n172 DVSS.n134 4.5005
R26446 DVSS.n160 DVSS.n134 4.5005
R26447 DVSS.n173 DVSS.n134 4.5005
R26448 DVSS.n23136 DVSS.n134 4.5005
R26449 DVSS.n159 DVSS.n134 4.5005
R26450 DVSS.n23138 DVSS.n134 4.5005
R26451 DVSS.n165 DVSS.n141 4.5005
R26452 DVSS.n167 DVSS.n141 4.5005
R26453 DVSS.n164 DVSS.n141 4.5005
R26454 DVSS.n169 DVSS.n141 4.5005
R26455 DVSS.n163 DVSS.n141 4.5005
R26456 DVSS.n170 DVSS.n141 4.5005
R26457 DVSS.n162 DVSS.n141 4.5005
R26458 DVSS.n171 DVSS.n141 4.5005
R26459 DVSS.n161 DVSS.n141 4.5005
R26460 DVSS.n172 DVSS.n141 4.5005
R26461 DVSS.n160 DVSS.n141 4.5005
R26462 DVSS.n173 DVSS.n141 4.5005
R26463 DVSS.n182 DVSS.n141 4.5005
R26464 DVSS.n23136 DVSS.n141 4.5005
R26465 DVSS.n23138 DVSS.n141 4.5005
R26466 DVSS.n165 DVSS.n133 4.5005
R26467 DVSS.n167 DVSS.n133 4.5005
R26468 DVSS.n164 DVSS.n133 4.5005
R26469 DVSS.n169 DVSS.n133 4.5005
R26470 DVSS.n163 DVSS.n133 4.5005
R26471 DVSS.n170 DVSS.n133 4.5005
R26472 DVSS.n162 DVSS.n133 4.5005
R26473 DVSS.n171 DVSS.n133 4.5005
R26474 DVSS.n161 DVSS.n133 4.5005
R26475 DVSS.n172 DVSS.n133 4.5005
R26476 DVSS.n160 DVSS.n133 4.5005
R26477 DVSS.n173 DVSS.n133 4.5005
R26478 DVSS.n23136 DVSS.n133 4.5005
R26479 DVSS.n23138 DVSS.n133 4.5005
R26480 DVSS.n165 DVSS.n142 4.5005
R26481 DVSS.n167 DVSS.n142 4.5005
R26482 DVSS.n164 DVSS.n142 4.5005
R26483 DVSS.n169 DVSS.n142 4.5005
R26484 DVSS.n163 DVSS.n142 4.5005
R26485 DVSS.n170 DVSS.n142 4.5005
R26486 DVSS.n162 DVSS.n142 4.5005
R26487 DVSS.n171 DVSS.n142 4.5005
R26488 DVSS.n161 DVSS.n142 4.5005
R26489 DVSS.n172 DVSS.n142 4.5005
R26490 DVSS.n160 DVSS.n142 4.5005
R26491 DVSS.n173 DVSS.n142 4.5005
R26492 DVSS.n23136 DVSS.n142 4.5005
R26493 DVSS.n23138 DVSS.n142 4.5005
R26494 DVSS.n165 DVSS.n132 4.5005
R26495 DVSS.n167 DVSS.n132 4.5005
R26496 DVSS.n164 DVSS.n132 4.5005
R26497 DVSS.n169 DVSS.n132 4.5005
R26498 DVSS.n163 DVSS.n132 4.5005
R26499 DVSS.n170 DVSS.n132 4.5005
R26500 DVSS.n162 DVSS.n132 4.5005
R26501 DVSS.n171 DVSS.n132 4.5005
R26502 DVSS.n161 DVSS.n132 4.5005
R26503 DVSS.n172 DVSS.n132 4.5005
R26504 DVSS.n160 DVSS.n132 4.5005
R26505 DVSS.n173 DVSS.n132 4.5005
R26506 DVSS.n182 DVSS.n132 4.5005
R26507 DVSS.n23136 DVSS.n132 4.5005
R26508 DVSS.n23138 DVSS.n132 4.5005
R26509 DVSS.n165 DVSS.n143 4.5005
R26510 DVSS.n167 DVSS.n143 4.5005
R26511 DVSS.n164 DVSS.n143 4.5005
R26512 DVSS.n169 DVSS.n143 4.5005
R26513 DVSS.n163 DVSS.n143 4.5005
R26514 DVSS.n170 DVSS.n143 4.5005
R26515 DVSS.n162 DVSS.n143 4.5005
R26516 DVSS.n171 DVSS.n143 4.5005
R26517 DVSS.n161 DVSS.n143 4.5005
R26518 DVSS.n172 DVSS.n143 4.5005
R26519 DVSS.n160 DVSS.n143 4.5005
R26520 DVSS.n173 DVSS.n143 4.5005
R26521 DVSS.n182 DVSS.n143 4.5005
R26522 DVSS.n23136 DVSS.n143 4.5005
R26523 DVSS.n23138 DVSS.n143 4.5005
R26524 DVSS.n165 DVSS.n131 4.5005
R26525 DVSS.n167 DVSS.n131 4.5005
R26526 DVSS.n164 DVSS.n131 4.5005
R26527 DVSS.n169 DVSS.n131 4.5005
R26528 DVSS.n163 DVSS.n131 4.5005
R26529 DVSS.n170 DVSS.n131 4.5005
R26530 DVSS.n162 DVSS.n131 4.5005
R26531 DVSS.n171 DVSS.n131 4.5005
R26532 DVSS.n161 DVSS.n131 4.5005
R26533 DVSS.n172 DVSS.n131 4.5005
R26534 DVSS.n160 DVSS.n131 4.5005
R26535 DVSS.n173 DVSS.n131 4.5005
R26536 DVSS.n23136 DVSS.n131 4.5005
R26537 DVSS.n23138 DVSS.n131 4.5005
R26538 DVSS.n165 DVSS.n144 4.5005
R26539 DVSS.n167 DVSS.n144 4.5005
R26540 DVSS.n164 DVSS.n144 4.5005
R26541 DVSS.n169 DVSS.n144 4.5005
R26542 DVSS.n163 DVSS.n144 4.5005
R26543 DVSS.n170 DVSS.n144 4.5005
R26544 DVSS.n162 DVSS.n144 4.5005
R26545 DVSS.n171 DVSS.n144 4.5005
R26546 DVSS.n161 DVSS.n144 4.5005
R26547 DVSS.n172 DVSS.n144 4.5005
R26548 DVSS.n160 DVSS.n144 4.5005
R26549 DVSS.n173 DVSS.n144 4.5005
R26550 DVSS.n23136 DVSS.n144 4.5005
R26551 DVSS.n23138 DVSS.n144 4.5005
R26552 DVSS.n165 DVSS.n130 4.5005
R26553 DVSS.n167 DVSS.n130 4.5005
R26554 DVSS.n164 DVSS.n130 4.5005
R26555 DVSS.n169 DVSS.n130 4.5005
R26556 DVSS.n163 DVSS.n130 4.5005
R26557 DVSS.n170 DVSS.n130 4.5005
R26558 DVSS.n162 DVSS.n130 4.5005
R26559 DVSS.n171 DVSS.n130 4.5005
R26560 DVSS.n161 DVSS.n130 4.5005
R26561 DVSS.n172 DVSS.n130 4.5005
R26562 DVSS.n160 DVSS.n130 4.5005
R26563 DVSS.n173 DVSS.n130 4.5005
R26564 DVSS.n182 DVSS.n130 4.5005
R26565 DVSS.n23136 DVSS.n130 4.5005
R26566 DVSS.n23138 DVSS.n130 4.5005
R26567 DVSS.n165 DVSS.n145 4.5005
R26568 DVSS.n167 DVSS.n145 4.5005
R26569 DVSS.n164 DVSS.n145 4.5005
R26570 DVSS.n169 DVSS.n145 4.5005
R26571 DVSS.n163 DVSS.n145 4.5005
R26572 DVSS.n170 DVSS.n145 4.5005
R26573 DVSS.n162 DVSS.n145 4.5005
R26574 DVSS.n171 DVSS.n145 4.5005
R26575 DVSS.n161 DVSS.n145 4.5005
R26576 DVSS.n172 DVSS.n145 4.5005
R26577 DVSS.n160 DVSS.n145 4.5005
R26578 DVSS.n173 DVSS.n145 4.5005
R26579 DVSS.n182 DVSS.n145 4.5005
R26580 DVSS.n23136 DVSS.n145 4.5005
R26581 DVSS.n23138 DVSS.n145 4.5005
R26582 DVSS.n165 DVSS.n129 4.5005
R26583 DVSS.n167 DVSS.n129 4.5005
R26584 DVSS.n164 DVSS.n129 4.5005
R26585 DVSS.n169 DVSS.n129 4.5005
R26586 DVSS.n163 DVSS.n129 4.5005
R26587 DVSS.n170 DVSS.n129 4.5005
R26588 DVSS.n162 DVSS.n129 4.5005
R26589 DVSS.n171 DVSS.n129 4.5005
R26590 DVSS.n161 DVSS.n129 4.5005
R26591 DVSS.n172 DVSS.n129 4.5005
R26592 DVSS.n160 DVSS.n129 4.5005
R26593 DVSS.n173 DVSS.n129 4.5005
R26594 DVSS.n23136 DVSS.n129 4.5005
R26595 DVSS.n23138 DVSS.n129 4.5005
R26596 DVSS.n165 DVSS.n146 4.5005
R26597 DVSS.n167 DVSS.n146 4.5005
R26598 DVSS.n164 DVSS.n146 4.5005
R26599 DVSS.n169 DVSS.n146 4.5005
R26600 DVSS.n163 DVSS.n146 4.5005
R26601 DVSS.n170 DVSS.n146 4.5005
R26602 DVSS.n162 DVSS.n146 4.5005
R26603 DVSS.n171 DVSS.n146 4.5005
R26604 DVSS.n161 DVSS.n146 4.5005
R26605 DVSS.n172 DVSS.n146 4.5005
R26606 DVSS.n160 DVSS.n146 4.5005
R26607 DVSS.n173 DVSS.n146 4.5005
R26608 DVSS.n23136 DVSS.n146 4.5005
R26609 DVSS.n23138 DVSS.n146 4.5005
R26610 DVSS.n165 DVSS.n128 4.5005
R26611 DVSS.n167 DVSS.n128 4.5005
R26612 DVSS.n164 DVSS.n128 4.5005
R26613 DVSS.n169 DVSS.n128 4.5005
R26614 DVSS.n163 DVSS.n128 4.5005
R26615 DVSS.n170 DVSS.n128 4.5005
R26616 DVSS.n162 DVSS.n128 4.5005
R26617 DVSS.n171 DVSS.n128 4.5005
R26618 DVSS.n161 DVSS.n128 4.5005
R26619 DVSS.n172 DVSS.n128 4.5005
R26620 DVSS.n160 DVSS.n128 4.5005
R26621 DVSS.n173 DVSS.n128 4.5005
R26622 DVSS.n182 DVSS.n128 4.5005
R26623 DVSS.n23136 DVSS.n128 4.5005
R26624 DVSS.n23138 DVSS.n128 4.5005
R26625 DVSS.n165 DVSS.n147 4.5005
R26626 DVSS.n167 DVSS.n147 4.5005
R26627 DVSS.n164 DVSS.n147 4.5005
R26628 DVSS.n169 DVSS.n147 4.5005
R26629 DVSS.n163 DVSS.n147 4.5005
R26630 DVSS.n170 DVSS.n147 4.5005
R26631 DVSS.n162 DVSS.n147 4.5005
R26632 DVSS.n171 DVSS.n147 4.5005
R26633 DVSS.n161 DVSS.n147 4.5005
R26634 DVSS.n172 DVSS.n147 4.5005
R26635 DVSS.n160 DVSS.n147 4.5005
R26636 DVSS.n173 DVSS.n147 4.5005
R26637 DVSS.n182 DVSS.n147 4.5005
R26638 DVSS.n23136 DVSS.n147 4.5005
R26639 DVSS.n23138 DVSS.n147 4.5005
R26640 DVSS.n165 DVSS.n127 4.5005
R26641 DVSS.n167 DVSS.n127 4.5005
R26642 DVSS.n164 DVSS.n127 4.5005
R26643 DVSS.n169 DVSS.n127 4.5005
R26644 DVSS.n163 DVSS.n127 4.5005
R26645 DVSS.n170 DVSS.n127 4.5005
R26646 DVSS.n162 DVSS.n127 4.5005
R26647 DVSS.n171 DVSS.n127 4.5005
R26648 DVSS.n161 DVSS.n127 4.5005
R26649 DVSS.n172 DVSS.n127 4.5005
R26650 DVSS.n160 DVSS.n127 4.5005
R26651 DVSS.n173 DVSS.n127 4.5005
R26652 DVSS.n23136 DVSS.n127 4.5005
R26653 DVSS.n23138 DVSS.n127 4.5005
R26654 DVSS.n165 DVSS.n148 4.5005
R26655 DVSS.n167 DVSS.n148 4.5005
R26656 DVSS.n164 DVSS.n148 4.5005
R26657 DVSS.n169 DVSS.n148 4.5005
R26658 DVSS.n163 DVSS.n148 4.5005
R26659 DVSS.n170 DVSS.n148 4.5005
R26660 DVSS.n162 DVSS.n148 4.5005
R26661 DVSS.n171 DVSS.n148 4.5005
R26662 DVSS.n161 DVSS.n148 4.5005
R26663 DVSS.n172 DVSS.n148 4.5005
R26664 DVSS.n160 DVSS.n148 4.5005
R26665 DVSS.n173 DVSS.n148 4.5005
R26666 DVSS.n23136 DVSS.n148 4.5005
R26667 DVSS.n159 DVSS.n148 4.5005
R26668 DVSS.n23138 DVSS.n148 4.5005
R26669 DVSS.n165 DVSS.n126 4.5005
R26670 DVSS.n167 DVSS.n126 4.5005
R26671 DVSS.n164 DVSS.n126 4.5005
R26672 DVSS.n169 DVSS.n126 4.5005
R26673 DVSS.n163 DVSS.n126 4.5005
R26674 DVSS.n170 DVSS.n126 4.5005
R26675 DVSS.n162 DVSS.n126 4.5005
R26676 DVSS.n171 DVSS.n126 4.5005
R26677 DVSS.n161 DVSS.n126 4.5005
R26678 DVSS.n172 DVSS.n126 4.5005
R26679 DVSS.n160 DVSS.n126 4.5005
R26680 DVSS.n173 DVSS.n126 4.5005
R26681 DVSS.n23136 DVSS.n126 4.5005
R26682 DVSS.n159 DVSS.n126 4.5005
R26683 DVSS.n23138 DVSS.n126 4.5005
R26684 DVSS.n23137 DVSS.n165 4.5005
R26685 DVSS.n23137 DVSS.n167 4.5005
R26686 DVSS.n23137 DVSS.n164 4.5005
R26687 DVSS.n23137 DVSS.n169 4.5005
R26688 DVSS.n23137 DVSS.n163 4.5005
R26689 DVSS.n23137 DVSS.n170 4.5005
R26690 DVSS.n23137 DVSS.n162 4.5005
R26691 DVSS.n23137 DVSS.n171 4.5005
R26692 DVSS.n23137 DVSS.n161 4.5005
R26693 DVSS.n23137 DVSS.n172 4.5005
R26694 DVSS.n23137 DVSS.n160 4.5005
R26695 DVSS.n23137 DVSS.n173 4.5005
R26696 DVSS.n23137 DVSS.n23136 4.5005
R26697 DVSS.n23137 DVSS.n159 4.5005
R26698 DVSS.n23138 DVSS.n23137 4.5005
R26699 DVSS.n100 DVSS.n72 4.5005
R26700 DVSS.n104 DVSS.n72 4.5005
R26701 DVSS.n98 DVSS.n72 4.5005
R26702 DVSS.n105 DVSS.n72 4.5005
R26703 DVSS.n97 DVSS.n72 4.5005
R26704 DVSS.n106 DVSS.n72 4.5005
R26705 DVSS.n96 DVSS.n72 4.5005
R26706 DVSS.n109 DVSS.n72 4.5005
R26707 DVSS.n23172 DVSS.n72 4.5005
R26708 DVSS.n23180 DVSS.n72 4.5005
R26709 DVSS.n94 DVSS.n72 4.5005
R26710 DVSS.n23182 DVSS.n72 4.5005
R26711 DVSS.n100 DVSS.n73 4.5005
R26712 DVSS.n103 DVSS.n73 4.5005
R26713 DVSS.n99 DVSS.n73 4.5005
R26714 DVSS.n104 DVSS.n73 4.5005
R26715 DVSS.n98 DVSS.n73 4.5005
R26716 DVSS.n105 DVSS.n73 4.5005
R26717 DVSS.n97 DVSS.n73 4.5005
R26718 DVSS.n106 DVSS.n73 4.5005
R26719 DVSS.n96 DVSS.n73 4.5005
R26720 DVSS.n108 DVSS.n73 4.5005
R26721 DVSS.n95 DVSS.n73 4.5005
R26722 DVSS.n109 DVSS.n73 4.5005
R26723 DVSS.n23180 DVSS.n73 4.5005
R26724 DVSS.n23182 DVSS.n73 4.5005
R26725 DVSS.n100 DVSS.n71 4.5005
R26726 DVSS.n103 DVSS.n71 4.5005
R26727 DVSS.n99 DVSS.n71 4.5005
R26728 DVSS.n104 DVSS.n71 4.5005
R26729 DVSS.n98 DVSS.n71 4.5005
R26730 DVSS.n105 DVSS.n71 4.5005
R26731 DVSS.n97 DVSS.n71 4.5005
R26732 DVSS.n106 DVSS.n71 4.5005
R26733 DVSS.n96 DVSS.n71 4.5005
R26734 DVSS.n108 DVSS.n71 4.5005
R26735 DVSS.n95 DVSS.n71 4.5005
R26736 DVSS.n109 DVSS.n71 4.5005
R26737 DVSS.n23180 DVSS.n71 4.5005
R26738 DVSS.n23182 DVSS.n71 4.5005
R26739 DVSS.n100 DVSS.n74 4.5005
R26740 DVSS.n103 DVSS.n74 4.5005
R26741 DVSS.n99 DVSS.n74 4.5005
R26742 DVSS.n104 DVSS.n74 4.5005
R26743 DVSS.n98 DVSS.n74 4.5005
R26744 DVSS.n105 DVSS.n74 4.5005
R26745 DVSS.n97 DVSS.n74 4.5005
R26746 DVSS.n106 DVSS.n74 4.5005
R26747 DVSS.n96 DVSS.n74 4.5005
R26748 DVSS.n108 DVSS.n74 4.5005
R26749 DVSS.n95 DVSS.n74 4.5005
R26750 DVSS.n109 DVSS.n74 4.5005
R26751 DVSS.n23180 DVSS.n74 4.5005
R26752 DVSS.n94 DVSS.n74 4.5005
R26753 DVSS.n23182 DVSS.n74 4.5005
R26754 DVSS.n100 DVSS.n70 4.5005
R26755 DVSS.n103 DVSS.n70 4.5005
R26756 DVSS.n99 DVSS.n70 4.5005
R26757 DVSS.n104 DVSS.n70 4.5005
R26758 DVSS.n98 DVSS.n70 4.5005
R26759 DVSS.n105 DVSS.n70 4.5005
R26760 DVSS.n97 DVSS.n70 4.5005
R26761 DVSS.n106 DVSS.n70 4.5005
R26762 DVSS.n96 DVSS.n70 4.5005
R26763 DVSS.n108 DVSS.n70 4.5005
R26764 DVSS.n95 DVSS.n70 4.5005
R26765 DVSS.n109 DVSS.n70 4.5005
R26766 DVSS.n23180 DVSS.n70 4.5005
R26767 DVSS.n23182 DVSS.n70 4.5005
R26768 DVSS.n100 DVSS.n75 4.5005
R26769 DVSS.n103 DVSS.n75 4.5005
R26770 DVSS.n99 DVSS.n75 4.5005
R26771 DVSS.n104 DVSS.n75 4.5005
R26772 DVSS.n98 DVSS.n75 4.5005
R26773 DVSS.n105 DVSS.n75 4.5005
R26774 DVSS.n97 DVSS.n75 4.5005
R26775 DVSS.n106 DVSS.n75 4.5005
R26776 DVSS.n96 DVSS.n75 4.5005
R26777 DVSS.n108 DVSS.n75 4.5005
R26778 DVSS.n95 DVSS.n75 4.5005
R26779 DVSS.n109 DVSS.n75 4.5005
R26780 DVSS.n23180 DVSS.n75 4.5005
R26781 DVSS.n23182 DVSS.n75 4.5005
R26782 DVSS.n100 DVSS.n69 4.5005
R26783 DVSS.n103 DVSS.n69 4.5005
R26784 DVSS.n99 DVSS.n69 4.5005
R26785 DVSS.n104 DVSS.n69 4.5005
R26786 DVSS.n98 DVSS.n69 4.5005
R26787 DVSS.n105 DVSS.n69 4.5005
R26788 DVSS.n97 DVSS.n69 4.5005
R26789 DVSS.n106 DVSS.n69 4.5005
R26790 DVSS.n96 DVSS.n69 4.5005
R26791 DVSS.n108 DVSS.n69 4.5005
R26792 DVSS.n95 DVSS.n69 4.5005
R26793 DVSS.n109 DVSS.n69 4.5005
R26794 DVSS.n23180 DVSS.n69 4.5005
R26795 DVSS.n94 DVSS.n69 4.5005
R26796 DVSS.n23182 DVSS.n69 4.5005
R26797 DVSS.n100 DVSS.n76 4.5005
R26798 DVSS.n103 DVSS.n76 4.5005
R26799 DVSS.n99 DVSS.n76 4.5005
R26800 DVSS.n104 DVSS.n76 4.5005
R26801 DVSS.n98 DVSS.n76 4.5005
R26802 DVSS.n105 DVSS.n76 4.5005
R26803 DVSS.n97 DVSS.n76 4.5005
R26804 DVSS.n106 DVSS.n76 4.5005
R26805 DVSS.n96 DVSS.n76 4.5005
R26806 DVSS.n108 DVSS.n76 4.5005
R26807 DVSS.n95 DVSS.n76 4.5005
R26808 DVSS.n109 DVSS.n76 4.5005
R26809 DVSS.n23172 DVSS.n76 4.5005
R26810 DVSS.n23180 DVSS.n76 4.5005
R26811 DVSS.n23182 DVSS.n76 4.5005
R26812 DVSS.n100 DVSS.n68 4.5005
R26813 DVSS.n103 DVSS.n68 4.5005
R26814 DVSS.n99 DVSS.n68 4.5005
R26815 DVSS.n104 DVSS.n68 4.5005
R26816 DVSS.n98 DVSS.n68 4.5005
R26817 DVSS.n105 DVSS.n68 4.5005
R26818 DVSS.n97 DVSS.n68 4.5005
R26819 DVSS.n106 DVSS.n68 4.5005
R26820 DVSS.n96 DVSS.n68 4.5005
R26821 DVSS.n108 DVSS.n68 4.5005
R26822 DVSS.n95 DVSS.n68 4.5005
R26823 DVSS.n109 DVSS.n68 4.5005
R26824 DVSS.n23180 DVSS.n68 4.5005
R26825 DVSS.n23182 DVSS.n68 4.5005
R26826 DVSS.n100 DVSS.n77 4.5005
R26827 DVSS.n103 DVSS.n77 4.5005
R26828 DVSS.n99 DVSS.n77 4.5005
R26829 DVSS.n104 DVSS.n77 4.5005
R26830 DVSS.n98 DVSS.n77 4.5005
R26831 DVSS.n105 DVSS.n77 4.5005
R26832 DVSS.n97 DVSS.n77 4.5005
R26833 DVSS.n106 DVSS.n77 4.5005
R26834 DVSS.n96 DVSS.n77 4.5005
R26835 DVSS.n108 DVSS.n77 4.5005
R26836 DVSS.n95 DVSS.n77 4.5005
R26837 DVSS.n109 DVSS.n77 4.5005
R26838 DVSS.n23180 DVSS.n77 4.5005
R26839 DVSS.n23182 DVSS.n77 4.5005
R26840 DVSS.n100 DVSS.n67 4.5005
R26841 DVSS.n103 DVSS.n67 4.5005
R26842 DVSS.n99 DVSS.n67 4.5005
R26843 DVSS.n104 DVSS.n67 4.5005
R26844 DVSS.n98 DVSS.n67 4.5005
R26845 DVSS.n105 DVSS.n67 4.5005
R26846 DVSS.n97 DVSS.n67 4.5005
R26847 DVSS.n106 DVSS.n67 4.5005
R26848 DVSS.n96 DVSS.n67 4.5005
R26849 DVSS.n108 DVSS.n67 4.5005
R26850 DVSS.n95 DVSS.n67 4.5005
R26851 DVSS.n109 DVSS.n67 4.5005
R26852 DVSS.n23172 DVSS.n67 4.5005
R26853 DVSS.n23180 DVSS.n67 4.5005
R26854 DVSS.n23182 DVSS.n67 4.5005
R26855 DVSS.n100 DVSS.n78 4.5005
R26856 DVSS.n103 DVSS.n78 4.5005
R26857 DVSS.n99 DVSS.n78 4.5005
R26858 DVSS.n104 DVSS.n78 4.5005
R26859 DVSS.n98 DVSS.n78 4.5005
R26860 DVSS.n105 DVSS.n78 4.5005
R26861 DVSS.n97 DVSS.n78 4.5005
R26862 DVSS.n106 DVSS.n78 4.5005
R26863 DVSS.n96 DVSS.n78 4.5005
R26864 DVSS.n108 DVSS.n78 4.5005
R26865 DVSS.n95 DVSS.n78 4.5005
R26866 DVSS.n109 DVSS.n78 4.5005
R26867 DVSS.n23172 DVSS.n78 4.5005
R26868 DVSS.n23180 DVSS.n78 4.5005
R26869 DVSS.n23182 DVSS.n78 4.5005
R26870 DVSS.n100 DVSS.n66 4.5005
R26871 DVSS.n103 DVSS.n66 4.5005
R26872 DVSS.n99 DVSS.n66 4.5005
R26873 DVSS.n104 DVSS.n66 4.5005
R26874 DVSS.n98 DVSS.n66 4.5005
R26875 DVSS.n105 DVSS.n66 4.5005
R26876 DVSS.n97 DVSS.n66 4.5005
R26877 DVSS.n106 DVSS.n66 4.5005
R26878 DVSS.n96 DVSS.n66 4.5005
R26879 DVSS.n108 DVSS.n66 4.5005
R26880 DVSS.n95 DVSS.n66 4.5005
R26881 DVSS.n109 DVSS.n66 4.5005
R26882 DVSS.n23180 DVSS.n66 4.5005
R26883 DVSS.n23182 DVSS.n66 4.5005
R26884 DVSS.n100 DVSS.n79 4.5005
R26885 DVSS.n103 DVSS.n79 4.5005
R26886 DVSS.n99 DVSS.n79 4.5005
R26887 DVSS.n104 DVSS.n79 4.5005
R26888 DVSS.n98 DVSS.n79 4.5005
R26889 DVSS.n105 DVSS.n79 4.5005
R26890 DVSS.n97 DVSS.n79 4.5005
R26891 DVSS.n106 DVSS.n79 4.5005
R26892 DVSS.n96 DVSS.n79 4.5005
R26893 DVSS.n108 DVSS.n79 4.5005
R26894 DVSS.n95 DVSS.n79 4.5005
R26895 DVSS.n109 DVSS.n79 4.5005
R26896 DVSS.n23180 DVSS.n79 4.5005
R26897 DVSS.n23182 DVSS.n79 4.5005
R26898 DVSS.n100 DVSS.n65 4.5005
R26899 DVSS.n103 DVSS.n65 4.5005
R26900 DVSS.n99 DVSS.n65 4.5005
R26901 DVSS.n104 DVSS.n65 4.5005
R26902 DVSS.n98 DVSS.n65 4.5005
R26903 DVSS.n105 DVSS.n65 4.5005
R26904 DVSS.n97 DVSS.n65 4.5005
R26905 DVSS.n106 DVSS.n65 4.5005
R26906 DVSS.n96 DVSS.n65 4.5005
R26907 DVSS.n108 DVSS.n65 4.5005
R26908 DVSS.n95 DVSS.n65 4.5005
R26909 DVSS.n109 DVSS.n65 4.5005
R26910 DVSS.n23172 DVSS.n65 4.5005
R26911 DVSS.n23180 DVSS.n65 4.5005
R26912 DVSS.n23182 DVSS.n65 4.5005
R26913 DVSS.n100 DVSS.n80 4.5005
R26914 DVSS.n103 DVSS.n80 4.5005
R26915 DVSS.n99 DVSS.n80 4.5005
R26916 DVSS.n104 DVSS.n80 4.5005
R26917 DVSS.n98 DVSS.n80 4.5005
R26918 DVSS.n105 DVSS.n80 4.5005
R26919 DVSS.n97 DVSS.n80 4.5005
R26920 DVSS.n106 DVSS.n80 4.5005
R26921 DVSS.n96 DVSS.n80 4.5005
R26922 DVSS.n108 DVSS.n80 4.5005
R26923 DVSS.n95 DVSS.n80 4.5005
R26924 DVSS.n109 DVSS.n80 4.5005
R26925 DVSS.n23172 DVSS.n80 4.5005
R26926 DVSS.n23180 DVSS.n80 4.5005
R26927 DVSS.n23182 DVSS.n80 4.5005
R26928 DVSS.n100 DVSS.n64 4.5005
R26929 DVSS.n103 DVSS.n64 4.5005
R26930 DVSS.n99 DVSS.n64 4.5005
R26931 DVSS.n104 DVSS.n64 4.5005
R26932 DVSS.n98 DVSS.n64 4.5005
R26933 DVSS.n105 DVSS.n64 4.5005
R26934 DVSS.n97 DVSS.n64 4.5005
R26935 DVSS.n106 DVSS.n64 4.5005
R26936 DVSS.n96 DVSS.n64 4.5005
R26937 DVSS.n108 DVSS.n64 4.5005
R26938 DVSS.n95 DVSS.n64 4.5005
R26939 DVSS.n109 DVSS.n64 4.5005
R26940 DVSS.n23180 DVSS.n64 4.5005
R26941 DVSS.n23182 DVSS.n64 4.5005
R26942 DVSS.n100 DVSS.n81 4.5005
R26943 DVSS.n103 DVSS.n81 4.5005
R26944 DVSS.n99 DVSS.n81 4.5005
R26945 DVSS.n104 DVSS.n81 4.5005
R26946 DVSS.n98 DVSS.n81 4.5005
R26947 DVSS.n105 DVSS.n81 4.5005
R26948 DVSS.n97 DVSS.n81 4.5005
R26949 DVSS.n106 DVSS.n81 4.5005
R26950 DVSS.n96 DVSS.n81 4.5005
R26951 DVSS.n108 DVSS.n81 4.5005
R26952 DVSS.n95 DVSS.n81 4.5005
R26953 DVSS.n109 DVSS.n81 4.5005
R26954 DVSS.n23180 DVSS.n81 4.5005
R26955 DVSS.n23182 DVSS.n81 4.5005
R26956 DVSS.n100 DVSS.n63 4.5005
R26957 DVSS.n103 DVSS.n63 4.5005
R26958 DVSS.n99 DVSS.n63 4.5005
R26959 DVSS.n104 DVSS.n63 4.5005
R26960 DVSS.n98 DVSS.n63 4.5005
R26961 DVSS.n105 DVSS.n63 4.5005
R26962 DVSS.n97 DVSS.n63 4.5005
R26963 DVSS.n106 DVSS.n63 4.5005
R26964 DVSS.n96 DVSS.n63 4.5005
R26965 DVSS.n108 DVSS.n63 4.5005
R26966 DVSS.n95 DVSS.n63 4.5005
R26967 DVSS.n109 DVSS.n63 4.5005
R26968 DVSS.n23172 DVSS.n63 4.5005
R26969 DVSS.n23180 DVSS.n63 4.5005
R26970 DVSS.n23182 DVSS.n63 4.5005
R26971 DVSS.n100 DVSS.n82 4.5005
R26972 DVSS.n103 DVSS.n82 4.5005
R26973 DVSS.n99 DVSS.n82 4.5005
R26974 DVSS.n104 DVSS.n82 4.5005
R26975 DVSS.n98 DVSS.n82 4.5005
R26976 DVSS.n105 DVSS.n82 4.5005
R26977 DVSS.n97 DVSS.n82 4.5005
R26978 DVSS.n106 DVSS.n82 4.5005
R26979 DVSS.n96 DVSS.n82 4.5005
R26980 DVSS.n108 DVSS.n82 4.5005
R26981 DVSS.n95 DVSS.n82 4.5005
R26982 DVSS.n109 DVSS.n82 4.5005
R26983 DVSS.n23172 DVSS.n82 4.5005
R26984 DVSS.n23180 DVSS.n82 4.5005
R26985 DVSS.n23182 DVSS.n82 4.5005
R26986 DVSS.n100 DVSS.n62 4.5005
R26987 DVSS.n103 DVSS.n62 4.5005
R26988 DVSS.n99 DVSS.n62 4.5005
R26989 DVSS.n104 DVSS.n62 4.5005
R26990 DVSS.n98 DVSS.n62 4.5005
R26991 DVSS.n105 DVSS.n62 4.5005
R26992 DVSS.n97 DVSS.n62 4.5005
R26993 DVSS.n106 DVSS.n62 4.5005
R26994 DVSS.n96 DVSS.n62 4.5005
R26995 DVSS.n108 DVSS.n62 4.5005
R26996 DVSS.n95 DVSS.n62 4.5005
R26997 DVSS.n109 DVSS.n62 4.5005
R26998 DVSS.n23180 DVSS.n62 4.5005
R26999 DVSS.n23182 DVSS.n62 4.5005
R27000 DVSS.n100 DVSS.n83 4.5005
R27001 DVSS.n103 DVSS.n83 4.5005
R27002 DVSS.n99 DVSS.n83 4.5005
R27003 DVSS.n104 DVSS.n83 4.5005
R27004 DVSS.n98 DVSS.n83 4.5005
R27005 DVSS.n105 DVSS.n83 4.5005
R27006 DVSS.n97 DVSS.n83 4.5005
R27007 DVSS.n106 DVSS.n83 4.5005
R27008 DVSS.n96 DVSS.n83 4.5005
R27009 DVSS.n108 DVSS.n83 4.5005
R27010 DVSS.n95 DVSS.n83 4.5005
R27011 DVSS.n109 DVSS.n83 4.5005
R27012 DVSS.n23180 DVSS.n83 4.5005
R27013 DVSS.n94 DVSS.n83 4.5005
R27014 DVSS.n23182 DVSS.n83 4.5005
R27015 DVSS.n100 DVSS.n61 4.5005
R27016 DVSS.n103 DVSS.n61 4.5005
R27017 DVSS.n99 DVSS.n61 4.5005
R27018 DVSS.n104 DVSS.n61 4.5005
R27019 DVSS.n98 DVSS.n61 4.5005
R27020 DVSS.n105 DVSS.n61 4.5005
R27021 DVSS.n97 DVSS.n61 4.5005
R27022 DVSS.n106 DVSS.n61 4.5005
R27023 DVSS.n96 DVSS.n61 4.5005
R27024 DVSS.n108 DVSS.n61 4.5005
R27025 DVSS.n95 DVSS.n61 4.5005
R27026 DVSS.n109 DVSS.n61 4.5005
R27027 DVSS.n23180 DVSS.n61 4.5005
R27028 DVSS.n94 DVSS.n61 4.5005
R27029 DVSS.n23182 DVSS.n61 4.5005
R27030 DVSS.n23181 DVSS.n100 4.5005
R27031 DVSS.n23181 DVSS.n103 4.5005
R27032 DVSS.n23181 DVSS.n99 4.5005
R27033 DVSS.n23181 DVSS.n104 4.5005
R27034 DVSS.n23181 DVSS.n98 4.5005
R27035 DVSS.n23181 DVSS.n105 4.5005
R27036 DVSS.n23181 DVSS.n97 4.5005
R27037 DVSS.n23181 DVSS.n106 4.5005
R27038 DVSS.n23181 DVSS.n96 4.5005
R27039 DVSS.n23181 DVSS.n108 4.5005
R27040 DVSS.n23181 DVSS.n95 4.5005
R27041 DVSS.n23181 DVSS.n109 4.5005
R27042 DVSS.n23181 DVSS.n23180 4.5005
R27043 DVSS.n23181 DVSS.n94 4.5005
R27044 DVSS.n23182 DVSS.n23181 4.5005
R27045 DVSS.n1251 DVSS.n1224 4.5005
R27046 DVSS.n22325 DVSS.n1251 4.5005
R27047 DVSS.n1251 DVSS.n1237 4.5005
R27048 DVSS.n1251 DVSS.n1225 4.5005
R27049 DVSS.n1251 DVSS.n1235 4.5005
R27050 DVSS.n1251 DVSS.n1227 4.5005
R27051 DVSS.n1251 DVSS.n1234 4.5005
R27052 DVSS.n1251 DVSS.n1228 4.5005
R27053 DVSS.n1251 DVSS.n1233 4.5005
R27054 DVSS.n1251 DVSS.n1229 4.5005
R27055 DVSS.n1251 DVSS.n1231 4.5005
R27056 DVSS.n1253 DVSS.n1224 4.5005
R27057 DVSS.n22325 DVSS.n1253 4.5005
R27058 DVSS.n1253 DVSS.n1237 4.5005
R27059 DVSS.n1253 DVSS.n1225 4.5005
R27060 DVSS.n1253 DVSS.n1236 4.5005
R27061 DVSS.n1253 DVSS.n1226 4.5005
R27062 DVSS.n1253 DVSS.n1235 4.5005
R27063 DVSS.n1253 DVSS.n1227 4.5005
R27064 DVSS.n1253 DVSS.n1234 4.5005
R27065 DVSS.n1253 DVSS.n1228 4.5005
R27066 DVSS.n1253 DVSS.n1233 4.5005
R27067 DVSS.n1253 DVSS.n1229 4.5005
R27068 DVSS.n1253 DVSS.n1232 4.5005
R27069 DVSS.n1253 DVSS.n1230 4.5005
R27070 DVSS.n1253 DVSS.n1231 4.5005
R27071 DVSS.n1248 DVSS.n1231 4.5005
R27072 DVSS.n1248 DVSS.n1230 4.5005
R27073 DVSS.n1248 DVSS.n1232 4.5005
R27074 DVSS.n1248 DVSS.n1229 4.5005
R27075 DVSS.n1248 DVSS.n1233 4.5005
R27076 DVSS.n1248 DVSS.n1228 4.5005
R27077 DVSS.n1248 DVSS.n1234 4.5005
R27078 DVSS.n1248 DVSS.n1227 4.5005
R27079 DVSS.n1248 DVSS.n1235 4.5005
R27080 DVSS.n1248 DVSS.n1226 4.5005
R27081 DVSS.n1248 DVSS.n1236 4.5005
R27082 DVSS.n1248 DVSS.n1225 4.5005
R27083 DVSS.n1248 DVSS.n1237 4.5005
R27084 DVSS.n1248 DVSS.n1224 4.5005
R27085 DVSS.n22325 DVSS.n1248 4.5005
R27086 DVSS.n1254 DVSS.n1231 4.5005
R27087 DVSS.n1254 DVSS.n1230 4.5005
R27088 DVSS.n1254 DVSS.n1232 4.5005
R27089 DVSS.n1254 DVSS.n1229 4.5005
R27090 DVSS.n1254 DVSS.n1233 4.5005
R27091 DVSS.n1254 DVSS.n1228 4.5005
R27092 DVSS.n1254 DVSS.n1234 4.5005
R27093 DVSS.n1254 DVSS.n1227 4.5005
R27094 DVSS.n1254 DVSS.n1235 4.5005
R27095 DVSS.n1254 DVSS.n1226 4.5005
R27096 DVSS.n1254 DVSS.n1236 4.5005
R27097 DVSS.n1254 DVSS.n1225 4.5005
R27098 DVSS.n1254 DVSS.n1237 4.5005
R27099 DVSS.n1254 DVSS.n1224 4.5005
R27100 DVSS.n22325 DVSS.n1254 4.5005
R27101 DVSS.n1247 DVSS.n1231 4.5005
R27102 DVSS.n1247 DVSS.n1230 4.5005
R27103 DVSS.n1247 DVSS.n1232 4.5005
R27104 DVSS.n1247 DVSS.n1229 4.5005
R27105 DVSS.n1247 DVSS.n1233 4.5005
R27106 DVSS.n1247 DVSS.n1228 4.5005
R27107 DVSS.n1247 DVSS.n1234 4.5005
R27108 DVSS.n1247 DVSS.n1227 4.5005
R27109 DVSS.n1247 DVSS.n1235 4.5005
R27110 DVSS.n1247 DVSS.n1226 4.5005
R27111 DVSS.n1247 DVSS.n1236 4.5005
R27112 DVSS.n1247 DVSS.n1225 4.5005
R27113 DVSS.n1247 DVSS.n1237 4.5005
R27114 DVSS.n1247 DVSS.n1224 4.5005
R27115 DVSS.n22325 DVSS.n1247 4.5005
R27116 DVSS.n1255 DVSS.n1224 4.5005
R27117 DVSS.n22325 DVSS.n1255 4.5005
R27118 DVSS.n1255 DVSS.n1237 4.5005
R27119 DVSS.n1255 DVSS.n1225 4.5005
R27120 DVSS.n1255 DVSS.n1236 4.5005
R27121 DVSS.n1255 DVSS.n1226 4.5005
R27122 DVSS.n1255 DVSS.n1235 4.5005
R27123 DVSS.n1255 DVSS.n1227 4.5005
R27124 DVSS.n1255 DVSS.n1234 4.5005
R27125 DVSS.n1255 DVSS.n1228 4.5005
R27126 DVSS.n1255 DVSS.n1233 4.5005
R27127 DVSS.n1255 DVSS.n1229 4.5005
R27128 DVSS.n1255 DVSS.n1232 4.5005
R27129 DVSS.n1255 DVSS.n1230 4.5005
R27130 DVSS.n1255 DVSS.n1231 4.5005
R27131 DVSS.n1246 DVSS.n1224 4.5005
R27132 DVSS.n22325 DVSS.n1246 4.5005
R27133 DVSS.n1246 DVSS.n1237 4.5005
R27134 DVSS.n1246 DVSS.n1225 4.5005
R27135 DVSS.n1246 DVSS.n1236 4.5005
R27136 DVSS.n1246 DVSS.n1226 4.5005
R27137 DVSS.n1246 DVSS.n1235 4.5005
R27138 DVSS.n1246 DVSS.n1227 4.5005
R27139 DVSS.n1246 DVSS.n1234 4.5005
R27140 DVSS.n1246 DVSS.n1228 4.5005
R27141 DVSS.n1246 DVSS.n1233 4.5005
R27142 DVSS.n1246 DVSS.n1229 4.5005
R27143 DVSS.n1246 DVSS.n1232 4.5005
R27144 DVSS.n1246 DVSS.n1230 4.5005
R27145 DVSS.n1246 DVSS.n1231 4.5005
R27146 DVSS.n1256 DVSS.n1224 4.5005
R27147 DVSS.n22325 DVSS.n1256 4.5005
R27148 DVSS.n1256 DVSS.n1237 4.5005
R27149 DVSS.n1256 DVSS.n1225 4.5005
R27150 DVSS.n1256 DVSS.n1236 4.5005
R27151 DVSS.n1256 DVSS.n1226 4.5005
R27152 DVSS.n1256 DVSS.n1235 4.5005
R27153 DVSS.n1256 DVSS.n1227 4.5005
R27154 DVSS.n1256 DVSS.n1234 4.5005
R27155 DVSS.n1256 DVSS.n1228 4.5005
R27156 DVSS.n1256 DVSS.n1233 4.5005
R27157 DVSS.n1256 DVSS.n1229 4.5005
R27158 DVSS.n1256 DVSS.n1232 4.5005
R27159 DVSS.n1256 DVSS.n1230 4.5005
R27160 DVSS.n1256 DVSS.n1231 4.5005
R27161 DVSS.n1245 DVSS.n1224 4.5005
R27162 DVSS.n22325 DVSS.n1245 4.5005
R27163 DVSS.n1245 DVSS.n1237 4.5005
R27164 DVSS.n1245 DVSS.n1225 4.5005
R27165 DVSS.n1245 DVSS.n1236 4.5005
R27166 DVSS.n1245 DVSS.n1226 4.5005
R27167 DVSS.n1245 DVSS.n1235 4.5005
R27168 DVSS.n1245 DVSS.n1227 4.5005
R27169 DVSS.n1245 DVSS.n1234 4.5005
R27170 DVSS.n1245 DVSS.n1228 4.5005
R27171 DVSS.n1245 DVSS.n1233 4.5005
R27172 DVSS.n1245 DVSS.n1229 4.5005
R27173 DVSS.n1245 DVSS.n1232 4.5005
R27174 DVSS.n1245 DVSS.n1230 4.5005
R27175 DVSS.n1245 DVSS.n1231 4.5005
R27176 DVSS.n1257 DVSS.n1231 4.5005
R27177 DVSS.n1257 DVSS.n1230 4.5005
R27178 DVSS.n1257 DVSS.n1232 4.5005
R27179 DVSS.n1257 DVSS.n1229 4.5005
R27180 DVSS.n1257 DVSS.n1233 4.5005
R27181 DVSS.n1257 DVSS.n1228 4.5005
R27182 DVSS.n1257 DVSS.n1234 4.5005
R27183 DVSS.n1257 DVSS.n1227 4.5005
R27184 DVSS.n1257 DVSS.n1235 4.5005
R27185 DVSS.n1257 DVSS.n1226 4.5005
R27186 DVSS.n1257 DVSS.n1236 4.5005
R27187 DVSS.n1257 DVSS.n1225 4.5005
R27188 DVSS.n1257 DVSS.n1237 4.5005
R27189 DVSS.n1257 DVSS.n1224 4.5005
R27190 DVSS.n22325 DVSS.n1257 4.5005
R27191 DVSS.n1244 DVSS.n1231 4.5005
R27192 DVSS.n1244 DVSS.n1230 4.5005
R27193 DVSS.n1244 DVSS.n1232 4.5005
R27194 DVSS.n1244 DVSS.n1229 4.5005
R27195 DVSS.n1244 DVSS.n1233 4.5005
R27196 DVSS.n1244 DVSS.n1228 4.5005
R27197 DVSS.n1244 DVSS.n1234 4.5005
R27198 DVSS.n1244 DVSS.n1227 4.5005
R27199 DVSS.n1244 DVSS.n1235 4.5005
R27200 DVSS.n1244 DVSS.n1226 4.5005
R27201 DVSS.n1244 DVSS.n1236 4.5005
R27202 DVSS.n1244 DVSS.n1225 4.5005
R27203 DVSS.n1244 DVSS.n1237 4.5005
R27204 DVSS.n1244 DVSS.n1224 4.5005
R27205 DVSS.n22325 DVSS.n1244 4.5005
R27206 DVSS.n1258 DVSS.n1231 4.5005
R27207 DVSS.n1258 DVSS.n1230 4.5005
R27208 DVSS.n1258 DVSS.n1232 4.5005
R27209 DVSS.n1258 DVSS.n1229 4.5005
R27210 DVSS.n1258 DVSS.n1233 4.5005
R27211 DVSS.n1258 DVSS.n1228 4.5005
R27212 DVSS.n1258 DVSS.n1234 4.5005
R27213 DVSS.n1258 DVSS.n1227 4.5005
R27214 DVSS.n1258 DVSS.n1235 4.5005
R27215 DVSS.n1258 DVSS.n1226 4.5005
R27216 DVSS.n1258 DVSS.n1236 4.5005
R27217 DVSS.n1258 DVSS.n1225 4.5005
R27218 DVSS.n1258 DVSS.n1237 4.5005
R27219 DVSS.n1258 DVSS.n1224 4.5005
R27220 DVSS.n22325 DVSS.n1258 4.5005
R27221 DVSS.n1243 DVSS.n1224 4.5005
R27222 DVSS.n22325 DVSS.n1243 4.5005
R27223 DVSS.n1243 DVSS.n1237 4.5005
R27224 DVSS.n1243 DVSS.n1225 4.5005
R27225 DVSS.n1243 DVSS.n1236 4.5005
R27226 DVSS.n1243 DVSS.n1226 4.5005
R27227 DVSS.n1243 DVSS.n1235 4.5005
R27228 DVSS.n1243 DVSS.n1227 4.5005
R27229 DVSS.n1243 DVSS.n1234 4.5005
R27230 DVSS.n1243 DVSS.n1228 4.5005
R27231 DVSS.n1243 DVSS.n1233 4.5005
R27232 DVSS.n1243 DVSS.n1229 4.5005
R27233 DVSS.n1243 DVSS.n1232 4.5005
R27234 DVSS.n1243 DVSS.n1230 4.5005
R27235 DVSS.n1243 DVSS.n1231 4.5005
R27236 DVSS.n1259 DVSS.n1224 4.5005
R27237 DVSS.n22325 DVSS.n1259 4.5005
R27238 DVSS.n1259 DVSS.n1237 4.5005
R27239 DVSS.n1259 DVSS.n1225 4.5005
R27240 DVSS.n1259 DVSS.n1236 4.5005
R27241 DVSS.n1259 DVSS.n1226 4.5005
R27242 DVSS.n1259 DVSS.n1235 4.5005
R27243 DVSS.n1259 DVSS.n1227 4.5005
R27244 DVSS.n1259 DVSS.n1234 4.5005
R27245 DVSS.n1259 DVSS.n1228 4.5005
R27246 DVSS.n1259 DVSS.n1233 4.5005
R27247 DVSS.n1259 DVSS.n1229 4.5005
R27248 DVSS.n1259 DVSS.n1232 4.5005
R27249 DVSS.n1259 DVSS.n1230 4.5005
R27250 DVSS.n1259 DVSS.n1231 4.5005
R27251 DVSS.n1242 DVSS.n1224 4.5005
R27252 DVSS.n22325 DVSS.n1242 4.5005
R27253 DVSS.n1242 DVSS.n1237 4.5005
R27254 DVSS.n1242 DVSS.n1225 4.5005
R27255 DVSS.n1242 DVSS.n1236 4.5005
R27256 DVSS.n1242 DVSS.n1226 4.5005
R27257 DVSS.n1242 DVSS.n1235 4.5005
R27258 DVSS.n1242 DVSS.n1227 4.5005
R27259 DVSS.n1242 DVSS.n1234 4.5005
R27260 DVSS.n1242 DVSS.n1228 4.5005
R27261 DVSS.n1242 DVSS.n1233 4.5005
R27262 DVSS.n1242 DVSS.n1229 4.5005
R27263 DVSS.n1242 DVSS.n1232 4.5005
R27264 DVSS.n1242 DVSS.n1230 4.5005
R27265 DVSS.n1242 DVSS.n1231 4.5005
R27266 DVSS.n1260 DVSS.n1231 4.5005
R27267 DVSS.n1260 DVSS.n1230 4.5005
R27268 DVSS.n1260 DVSS.n1232 4.5005
R27269 DVSS.n1260 DVSS.n1229 4.5005
R27270 DVSS.n1260 DVSS.n1233 4.5005
R27271 DVSS.n1260 DVSS.n1228 4.5005
R27272 DVSS.n1260 DVSS.n1234 4.5005
R27273 DVSS.n1260 DVSS.n1227 4.5005
R27274 DVSS.n1260 DVSS.n1235 4.5005
R27275 DVSS.n1260 DVSS.n1226 4.5005
R27276 DVSS.n1260 DVSS.n1236 4.5005
R27277 DVSS.n1260 DVSS.n1225 4.5005
R27278 DVSS.n1260 DVSS.n1237 4.5005
R27279 DVSS.n1260 DVSS.n1224 4.5005
R27280 DVSS.n22325 DVSS.n1260 4.5005
R27281 DVSS.n1241 DVSS.n1231 4.5005
R27282 DVSS.n1241 DVSS.n1230 4.5005
R27283 DVSS.n1241 DVSS.n1232 4.5005
R27284 DVSS.n1241 DVSS.n1229 4.5005
R27285 DVSS.n1241 DVSS.n1233 4.5005
R27286 DVSS.n1241 DVSS.n1228 4.5005
R27287 DVSS.n1241 DVSS.n1234 4.5005
R27288 DVSS.n1241 DVSS.n1227 4.5005
R27289 DVSS.n1241 DVSS.n1235 4.5005
R27290 DVSS.n1241 DVSS.n1226 4.5005
R27291 DVSS.n1241 DVSS.n1236 4.5005
R27292 DVSS.n1241 DVSS.n1225 4.5005
R27293 DVSS.n1241 DVSS.n1237 4.5005
R27294 DVSS.n1241 DVSS.n1224 4.5005
R27295 DVSS.n22325 DVSS.n1241 4.5005
R27296 DVSS.n1261 DVSS.n1231 4.5005
R27297 DVSS.n1261 DVSS.n1230 4.5005
R27298 DVSS.n1261 DVSS.n1232 4.5005
R27299 DVSS.n1261 DVSS.n1229 4.5005
R27300 DVSS.n1261 DVSS.n1233 4.5005
R27301 DVSS.n1261 DVSS.n1228 4.5005
R27302 DVSS.n1261 DVSS.n1234 4.5005
R27303 DVSS.n1261 DVSS.n1227 4.5005
R27304 DVSS.n1261 DVSS.n1235 4.5005
R27305 DVSS.n1261 DVSS.n1226 4.5005
R27306 DVSS.n1261 DVSS.n1236 4.5005
R27307 DVSS.n1261 DVSS.n1225 4.5005
R27308 DVSS.n1261 DVSS.n1237 4.5005
R27309 DVSS.n1261 DVSS.n1224 4.5005
R27310 DVSS.n22325 DVSS.n1261 4.5005
R27311 DVSS.n1240 DVSS.n1231 4.5005
R27312 DVSS.n1240 DVSS.n1230 4.5005
R27313 DVSS.n1240 DVSS.n1232 4.5005
R27314 DVSS.n1240 DVSS.n1229 4.5005
R27315 DVSS.n1240 DVSS.n1233 4.5005
R27316 DVSS.n1240 DVSS.n1228 4.5005
R27317 DVSS.n1240 DVSS.n1234 4.5005
R27318 DVSS.n1240 DVSS.n1227 4.5005
R27319 DVSS.n1240 DVSS.n1235 4.5005
R27320 DVSS.n1240 DVSS.n1226 4.5005
R27321 DVSS.n1240 DVSS.n1236 4.5005
R27322 DVSS.n1240 DVSS.n1225 4.5005
R27323 DVSS.n1240 DVSS.n1237 4.5005
R27324 DVSS.n1240 DVSS.n1224 4.5005
R27325 DVSS.n22325 DVSS.n1240 4.5005
R27326 DVSS.n1262 DVSS.n1224 4.5005
R27327 DVSS.n22325 DVSS.n1262 4.5005
R27328 DVSS.n1262 DVSS.n1237 4.5005
R27329 DVSS.n1262 DVSS.n1225 4.5005
R27330 DVSS.n1262 DVSS.n1236 4.5005
R27331 DVSS.n1262 DVSS.n1226 4.5005
R27332 DVSS.n1262 DVSS.n1235 4.5005
R27333 DVSS.n1262 DVSS.n1227 4.5005
R27334 DVSS.n1262 DVSS.n1234 4.5005
R27335 DVSS.n1262 DVSS.n1228 4.5005
R27336 DVSS.n1262 DVSS.n1233 4.5005
R27337 DVSS.n1262 DVSS.n1229 4.5005
R27338 DVSS.n1262 DVSS.n1232 4.5005
R27339 DVSS.n1262 DVSS.n1230 4.5005
R27340 DVSS.n1262 DVSS.n1231 4.5005
R27341 DVSS.n1239 DVSS.n1224 4.5005
R27342 DVSS.n22325 DVSS.n1239 4.5005
R27343 DVSS.n1239 DVSS.n1237 4.5005
R27344 DVSS.n1239 DVSS.n1225 4.5005
R27345 DVSS.n1239 DVSS.n1236 4.5005
R27346 DVSS.n1239 DVSS.n1226 4.5005
R27347 DVSS.n1239 DVSS.n1235 4.5005
R27348 DVSS.n1239 DVSS.n1227 4.5005
R27349 DVSS.n1239 DVSS.n1234 4.5005
R27350 DVSS.n1239 DVSS.n1228 4.5005
R27351 DVSS.n1239 DVSS.n1233 4.5005
R27352 DVSS.n1239 DVSS.n1229 4.5005
R27353 DVSS.n1239 DVSS.n1232 4.5005
R27354 DVSS.n1239 DVSS.n1230 4.5005
R27355 DVSS.n1239 DVSS.n1231 4.5005
R27356 DVSS.n22324 DVSS.n1224 4.5005
R27357 DVSS.n22325 DVSS.n22324 4.5005
R27358 DVSS.n22324 DVSS.n1237 4.5005
R27359 DVSS.n22324 DVSS.n1225 4.5005
R27360 DVSS.n22324 DVSS.n1236 4.5005
R27361 DVSS.n22324 DVSS.n1226 4.5005
R27362 DVSS.n22324 DVSS.n1235 4.5005
R27363 DVSS.n22324 DVSS.n1227 4.5005
R27364 DVSS.n22324 DVSS.n1234 4.5005
R27365 DVSS.n22324 DVSS.n1228 4.5005
R27366 DVSS.n22324 DVSS.n1233 4.5005
R27367 DVSS.n22324 DVSS.n1229 4.5005
R27368 DVSS.n22324 DVSS.n1232 4.5005
R27369 DVSS.n22324 DVSS.n1230 4.5005
R27370 DVSS.n22324 DVSS.n1231 4.5005
R27371 DVSS.n22326 DVSS.n1231 4.5005
R27372 DVSS.n22326 DVSS.n1230 4.5005
R27373 DVSS.n22326 DVSS.n1232 4.5005
R27374 DVSS.n22326 DVSS.n1229 4.5005
R27375 DVSS.n22326 DVSS.n1233 4.5005
R27376 DVSS.n22326 DVSS.n1228 4.5005
R27377 DVSS.n22326 DVSS.n1234 4.5005
R27378 DVSS.n22326 DVSS.n1227 4.5005
R27379 DVSS.n22326 DVSS.n1235 4.5005
R27380 DVSS.n22326 DVSS.n1226 4.5005
R27381 DVSS.n22326 DVSS.n1236 4.5005
R27382 DVSS.n22326 DVSS.n1225 4.5005
R27383 DVSS.n22326 DVSS.n1237 4.5005
R27384 DVSS.n22326 DVSS.n1224 4.5005
R27385 DVSS.n22326 DVSS.n22325 4.5005
R27386 DVSS.n1231 DVSS.n1221 4.5005
R27387 DVSS.n1230 DVSS.n1221 4.5005
R27388 DVSS.n1232 DVSS.n1221 4.5005
R27389 DVSS.n1229 DVSS.n1221 4.5005
R27390 DVSS.n1233 DVSS.n1221 4.5005
R27391 DVSS.n1228 DVSS.n1221 4.5005
R27392 DVSS.n1234 DVSS.n1221 4.5005
R27393 DVSS.n1227 DVSS.n1221 4.5005
R27394 DVSS.n1235 DVSS.n1221 4.5005
R27395 DVSS.n1226 DVSS.n1221 4.5005
R27396 DVSS.n1236 DVSS.n1221 4.5005
R27397 DVSS.n1225 DVSS.n1221 4.5005
R27398 DVSS.n1237 DVSS.n1221 4.5005
R27399 DVSS.n1224 DVSS.n1221 4.5005
R27400 DVSS.n22325 DVSS.n1221 4.5005
R27401 DVSS.n1392 DVSS.n1363 4.5005
R27402 DVSS.n22184 DVSS.n1392 4.5005
R27403 DVSS.n22120 DVSS.n1363 4.5005
R27404 DVSS.n22184 DVSS.n22120 4.5005
R27405 DVSS.n1391 DVSS.n1371 4.5005
R27406 DVSS.n1391 DVSS.n1368 4.5005
R27407 DVSS.n1391 DVSS.n1373 4.5005
R27408 DVSS.n1391 DVSS.n1367 4.5005
R27409 DVSS.n1391 DVSS.n1374 4.5005
R27410 DVSS.n1391 DVSS.n1366 4.5005
R27411 DVSS.n1391 DVSS.n1375 4.5005
R27412 DVSS.n1391 DVSS.n1364 4.5005
R27413 DVSS.n1391 DVSS.n1377 4.5005
R27414 DVSS.n1391 DVSS.n1363 4.5005
R27415 DVSS.n22184 DVSS.n1391 4.5005
R27416 DVSS.n22121 DVSS.n1371 4.5005
R27417 DVSS.n22121 DVSS.n1369 4.5005
R27418 DVSS.n22121 DVSS.n1372 4.5005
R27419 DVSS.n22121 DVSS.n1368 4.5005
R27420 DVSS.n22121 DVSS.n1373 4.5005
R27421 DVSS.n22121 DVSS.n1367 4.5005
R27422 DVSS.n22121 DVSS.n1374 4.5005
R27423 DVSS.n22121 DVSS.n1366 4.5005
R27424 DVSS.n22121 DVSS.n1375 4.5005
R27425 DVSS.n22121 DVSS.n1365 4.5005
R27426 DVSS.n22121 DVSS.n1376 4.5005
R27427 DVSS.n22121 DVSS.n1364 4.5005
R27428 DVSS.n22121 DVSS.n1377 4.5005
R27429 DVSS.n22121 DVSS.n1363 4.5005
R27430 DVSS.n22184 DVSS.n22121 4.5005
R27431 DVSS.n1388 DVSS.n1371 4.5005
R27432 DVSS.n1388 DVSS.n1369 4.5005
R27433 DVSS.n1388 DVSS.n1372 4.5005
R27434 DVSS.n1388 DVSS.n1368 4.5005
R27435 DVSS.n1388 DVSS.n1373 4.5005
R27436 DVSS.n1388 DVSS.n1367 4.5005
R27437 DVSS.n1388 DVSS.n1374 4.5005
R27438 DVSS.n1388 DVSS.n1366 4.5005
R27439 DVSS.n1388 DVSS.n1375 4.5005
R27440 DVSS.n1388 DVSS.n1365 4.5005
R27441 DVSS.n1388 DVSS.n1376 4.5005
R27442 DVSS.n1388 DVSS.n1364 4.5005
R27443 DVSS.n1388 DVSS.n1377 4.5005
R27444 DVSS.n1388 DVSS.n1363 4.5005
R27445 DVSS.n22184 DVSS.n1388 4.5005
R27446 DVSS.n22122 DVSS.n1363 4.5005
R27447 DVSS.n22184 DVSS.n22122 4.5005
R27448 DVSS.n1387 DVSS.n1363 4.5005
R27449 DVSS.n22184 DVSS.n1387 4.5005
R27450 DVSS.n22123 DVSS.n1363 4.5005
R27451 DVSS.n22184 DVSS.n22123 4.5005
R27452 DVSS.n1386 DVSS.n1363 4.5005
R27453 DVSS.n22184 DVSS.n1386 4.5005
R27454 DVSS.n22124 DVSS.n1371 4.5005
R27455 DVSS.n22124 DVSS.n1369 4.5005
R27456 DVSS.n22124 DVSS.n1372 4.5005
R27457 DVSS.n22124 DVSS.n1368 4.5005
R27458 DVSS.n22124 DVSS.n1373 4.5005
R27459 DVSS.n22124 DVSS.n1367 4.5005
R27460 DVSS.n22124 DVSS.n1374 4.5005
R27461 DVSS.n22124 DVSS.n1366 4.5005
R27462 DVSS.n22124 DVSS.n1375 4.5005
R27463 DVSS.n22124 DVSS.n1365 4.5005
R27464 DVSS.n22124 DVSS.n1376 4.5005
R27465 DVSS.n22124 DVSS.n1364 4.5005
R27466 DVSS.n22124 DVSS.n1377 4.5005
R27467 DVSS.n22124 DVSS.n1363 4.5005
R27468 DVSS.n22184 DVSS.n22124 4.5005
R27469 DVSS.n1385 DVSS.n1371 4.5005
R27470 DVSS.n1385 DVSS.n1369 4.5005
R27471 DVSS.n1385 DVSS.n1372 4.5005
R27472 DVSS.n1385 DVSS.n1368 4.5005
R27473 DVSS.n1385 DVSS.n1373 4.5005
R27474 DVSS.n1385 DVSS.n1367 4.5005
R27475 DVSS.n1385 DVSS.n1374 4.5005
R27476 DVSS.n1385 DVSS.n1366 4.5005
R27477 DVSS.n1385 DVSS.n1375 4.5005
R27478 DVSS.n1385 DVSS.n1365 4.5005
R27479 DVSS.n1385 DVSS.n1376 4.5005
R27480 DVSS.n1385 DVSS.n1364 4.5005
R27481 DVSS.n1385 DVSS.n1377 4.5005
R27482 DVSS.n1385 DVSS.n1363 4.5005
R27483 DVSS.n22184 DVSS.n1385 4.5005
R27484 DVSS.n22125 DVSS.n1371 4.5005
R27485 DVSS.n22125 DVSS.n1369 4.5005
R27486 DVSS.n22125 DVSS.n1372 4.5005
R27487 DVSS.n22125 DVSS.n1368 4.5005
R27488 DVSS.n22125 DVSS.n1373 4.5005
R27489 DVSS.n22125 DVSS.n1367 4.5005
R27490 DVSS.n22125 DVSS.n1374 4.5005
R27491 DVSS.n22125 DVSS.n1366 4.5005
R27492 DVSS.n22125 DVSS.n1375 4.5005
R27493 DVSS.n22125 DVSS.n1365 4.5005
R27494 DVSS.n22125 DVSS.n1376 4.5005
R27495 DVSS.n22125 DVSS.n1364 4.5005
R27496 DVSS.n22125 DVSS.n1377 4.5005
R27497 DVSS.n22125 DVSS.n1363 4.5005
R27498 DVSS.n22184 DVSS.n22125 4.5005
R27499 DVSS.n1384 DVSS.n1363 4.5005
R27500 DVSS.n22184 DVSS.n1384 4.5005
R27501 DVSS.n22126 DVSS.n1363 4.5005
R27502 DVSS.n22184 DVSS.n22126 4.5005
R27503 DVSS.n1383 DVSS.n1363 4.5005
R27504 DVSS.n22184 DVSS.n1383 4.5005
R27505 DVSS.n22127 DVSS.n1371 4.5005
R27506 DVSS.n22127 DVSS.n1369 4.5005
R27507 DVSS.n22127 DVSS.n1372 4.5005
R27508 DVSS.n22127 DVSS.n1368 4.5005
R27509 DVSS.n22127 DVSS.n1373 4.5005
R27510 DVSS.n22127 DVSS.n1367 4.5005
R27511 DVSS.n22127 DVSS.n1374 4.5005
R27512 DVSS.n22127 DVSS.n1366 4.5005
R27513 DVSS.n22127 DVSS.n1375 4.5005
R27514 DVSS.n22127 DVSS.n1365 4.5005
R27515 DVSS.n22127 DVSS.n1376 4.5005
R27516 DVSS.n22127 DVSS.n1364 4.5005
R27517 DVSS.n22127 DVSS.n1377 4.5005
R27518 DVSS.n22127 DVSS.n1363 4.5005
R27519 DVSS.n22184 DVSS.n22127 4.5005
R27520 DVSS.n1382 DVSS.n1371 4.5005
R27521 DVSS.n1382 DVSS.n1369 4.5005
R27522 DVSS.n1382 DVSS.n1372 4.5005
R27523 DVSS.n1382 DVSS.n1368 4.5005
R27524 DVSS.n1382 DVSS.n1373 4.5005
R27525 DVSS.n1382 DVSS.n1367 4.5005
R27526 DVSS.n1382 DVSS.n1374 4.5005
R27527 DVSS.n1382 DVSS.n1366 4.5005
R27528 DVSS.n1382 DVSS.n1375 4.5005
R27529 DVSS.n1382 DVSS.n1365 4.5005
R27530 DVSS.n1382 DVSS.n1376 4.5005
R27531 DVSS.n1382 DVSS.n1364 4.5005
R27532 DVSS.n1382 DVSS.n1377 4.5005
R27533 DVSS.n1382 DVSS.n1363 4.5005
R27534 DVSS.n22184 DVSS.n1382 4.5005
R27535 DVSS.n22128 DVSS.n1371 4.5005
R27536 DVSS.n22128 DVSS.n1369 4.5005
R27537 DVSS.n22128 DVSS.n1372 4.5005
R27538 DVSS.n22128 DVSS.n1368 4.5005
R27539 DVSS.n22128 DVSS.n1373 4.5005
R27540 DVSS.n22128 DVSS.n1367 4.5005
R27541 DVSS.n22128 DVSS.n1374 4.5005
R27542 DVSS.n22128 DVSS.n1366 4.5005
R27543 DVSS.n22128 DVSS.n1375 4.5005
R27544 DVSS.n22128 DVSS.n1365 4.5005
R27545 DVSS.n22128 DVSS.n1376 4.5005
R27546 DVSS.n22128 DVSS.n1364 4.5005
R27547 DVSS.n22128 DVSS.n1377 4.5005
R27548 DVSS.n22128 DVSS.n1363 4.5005
R27549 DVSS.n22184 DVSS.n22128 4.5005
R27550 DVSS.n1381 DVSS.n1371 4.5005
R27551 DVSS.n1381 DVSS.n1369 4.5005
R27552 DVSS.n1381 DVSS.n1372 4.5005
R27553 DVSS.n1381 DVSS.n1368 4.5005
R27554 DVSS.n1381 DVSS.n1373 4.5005
R27555 DVSS.n1381 DVSS.n1367 4.5005
R27556 DVSS.n1381 DVSS.n1374 4.5005
R27557 DVSS.n1381 DVSS.n1366 4.5005
R27558 DVSS.n1381 DVSS.n1375 4.5005
R27559 DVSS.n1381 DVSS.n1365 4.5005
R27560 DVSS.n1381 DVSS.n1376 4.5005
R27561 DVSS.n1381 DVSS.n1364 4.5005
R27562 DVSS.n1381 DVSS.n1377 4.5005
R27563 DVSS.n1381 DVSS.n1363 4.5005
R27564 DVSS.n22184 DVSS.n1381 4.5005
R27565 DVSS.n22129 DVSS.n1363 4.5005
R27566 DVSS.n22184 DVSS.n22129 4.5005
R27567 DVSS.n1380 DVSS.n1363 4.5005
R27568 DVSS.n22184 DVSS.n1380 4.5005
R27569 DVSS.n22183 DVSS.n1363 4.5005
R27570 DVSS.n22184 DVSS.n22183 4.5005
R27571 DVSS.n1379 DVSS.n1371 4.5005
R27572 DVSS.n1379 DVSS.n1369 4.5005
R27573 DVSS.n1379 DVSS.n1372 4.5005
R27574 DVSS.n1379 DVSS.n1368 4.5005
R27575 DVSS.n1379 DVSS.n1373 4.5005
R27576 DVSS.n1379 DVSS.n1367 4.5005
R27577 DVSS.n1379 DVSS.n1374 4.5005
R27578 DVSS.n1379 DVSS.n1366 4.5005
R27579 DVSS.n1379 DVSS.n1375 4.5005
R27580 DVSS.n1379 DVSS.n1365 4.5005
R27581 DVSS.n1379 DVSS.n1376 4.5005
R27582 DVSS.n1379 DVSS.n1364 4.5005
R27583 DVSS.n1379 DVSS.n1377 4.5005
R27584 DVSS.n1379 DVSS.n1363 4.5005
R27585 DVSS.n22184 DVSS.n1379 4.5005
R27586 DVSS.n22185 DVSS.n1371 4.5005
R27587 DVSS.n22185 DVSS.n1369 4.5005
R27588 DVSS.n22185 DVSS.n1372 4.5005
R27589 DVSS.n22185 DVSS.n1368 4.5005
R27590 DVSS.n22185 DVSS.n1373 4.5005
R27591 DVSS.n22185 DVSS.n1367 4.5005
R27592 DVSS.n22185 DVSS.n1374 4.5005
R27593 DVSS.n22185 DVSS.n1366 4.5005
R27594 DVSS.n22185 DVSS.n1375 4.5005
R27595 DVSS.n22185 DVSS.n1365 4.5005
R27596 DVSS.n22185 DVSS.n1376 4.5005
R27597 DVSS.n22185 DVSS.n1364 4.5005
R27598 DVSS.n22185 DVSS.n1377 4.5005
R27599 DVSS.n22185 DVSS.n1363 4.5005
R27600 DVSS.n22185 DVSS.n22184 4.5005
R27601 DVSS.n22183 DVSS.n1377 4.5005
R27602 DVSS.n22183 DVSS.n1364 4.5005
R27603 DVSS.n22183 DVSS.n1376 4.5005
R27604 DVSS.n22183 DVSS.n1365 4.5005
R27605 DVSS.n22183 DVSS.n1375 4.5005
R27606 DVSS.n22183 DVSS.n1366 4.5005
R27607 DVSS.n22183 DVSS.n1374 4.5005
R27608 DVSS.n22183 DVSS.n1367 4.5005
R27609 DVSS.n22183 DVSS.n1373 4.5005
R27610 DVSS.n22183 DVSS.n1368 4.5005
R27611 DVSS.n22183 DVSS.n1372 4.5005
R27612 DVSS.n22183 DVSS.n1369 4.5005
R27613 DVSS.n22183 DVSS.n1371 4.5005
R27614 DVSS.n1380 DVSS.n1377 4.5005
R27615 DVSS.n1380 DVSS.n1364 4.5005
R27616 DVSS.n1380 DVSS.n1376 4.5005
R27617 DVSS.n1380 DVSS.n1365 4.5005
R27618 DVSS.n1380 DVSS.n1375 4.5005
R27619 DVSS.n1380 DVSS.n1366 4.5005
R27620 DVSS.n1380 DVSS.n1374 4.5005
R27621 DVSS.n1380 DVSS.n1367 4.5005
R27622 DVSS.n1380 DVSS.n1373 4.5005
R27623 DVSS.n1380 DVSS.n1368 4.5005
R27624 DVSS.n1380 DVSS.n1372 4.5005
R27625 DVSS.n1380 DVSS.n1369 4.5005
R27626 DVSS.n1380 DVSS.n1371 4.5005
R27627 DVSS.n22129 DVSS.n1377 4.5005
R27628 DVSS.n22129 DVSS.n1364 4.5005
R27629 DVSS.n22129 DVSS.n1376 4.5005
R27630 DVSS.n22129 DVSS.n1365 4.5005
R27631 DVSS.n22129 DVSS.n1375 4.5005
R27632 DVSS.n22129 DVSS.n1366 4.5005
R27633 DVSS.n22129 DVSS.n1374 4.5005
R27634 DVSS.n22129 DVSS.n1367 4.5005
R27635 DVSS.n22129 DVSS.n1373 4.5005
R27636 DVSS.n22129 DVSS.n1368 4.5005
R27637 DVSS.n22129 DVSS.n1372 4.5005
R27638 DVSS.n22129 DVSS.n1369 4.5005
R27639 DVSS.n22129 DVSS.n1371 4.5005
R27640 DVSS.n1383 DVSS.n1377 4.5005
R27641 DVSS.n1383 DVSS.n1364 4.5005
R27642 DVSS.n1383 DVSS.n1376 4.5005
R27643 DVSS.n1383 DVSS.n1365 4.5005
R27644 DVSS.n1383 DVSS.n1375 4.5005
R27645 DVSS.n1383 DVSS.n1366 4.5005
R27646 DVSS.n1383 DVSS.n1374 4.5005
R27647 DVSS.n1383 DVSS.n1367 4.5005
R27648 DVSS.n1383 DVSS.n1373 4.5005
R27649 DVSS.n1383 DVSS.n1368 4.5005
R27650 DVSS.n1383 DVSS.n1372 4.5005
R27651 DVSS.n1383 DVSS.n1369 4.5005
R27652 DVSS.n1383 DVSS.n1371 4.5005
R27653 DVSS.n22126 DVSS.n1377 4.5005
R27654 DVSS.n22126 DVSS.n1364 4.5005
R27655 DVSS.n22126 DVSS.n1376 4.5005
R27656 DVSS.n22126 DVSS.n1365 4.5005
R27657 DVSS.n22126 DVSS.n1375 4.5005
R27658 DVSS.n22126 DVSS.n1366 4.5005
R27659 DVSS.n22126 DVSS.n1374 4.5005
R27660 DVSS.n22126 DVSS.n1367 4.5005
R27661 DVSS.n22126 DVSS.n1373 4.5005
R27662 DVSS.n22126 DVSS.n1368 4.5005
R27663 DVSS.n22126 DVSS.n1372 4.5005
R27664 DVSS.n22126 DVSS.n1369 4.5005
R27665 DVSS.n22126 DVSS.n1371 4.5005
R27666 DVSS.n1384 DVSS.n1377 4.5005
R27667 DVSS.n1384 DVSS.n1364 4.5005
R27668 DVSS.n1384 DVSS.n1376 4.5005
R27669 DVSS.n1384 DVSS.n1365 4.5005
R27670 DVSS.n1384 DVSS.n1375 4.5005
R27671 DVSS.n1384 DVSS.n1366 4.5005
R27672 DVSS.n1384 DVSS.n1374 4.5005
R27673 DVSS.n1384 DVSS.n1367 4.5005
R27674 DVSS.n1384 DVSS.n1373 4.5005
R27675 DVSS.n1384 DVSS.n1368 4.5005
R27676 DVSS.n1384 DVSS.n1372 4.5005
R27677 DVSS.n1384 DVSS.n1369 4.5005
R27678 DVSS.n1384 DVSS.n1371 4.5005
R27679 DVSS.n1386 DVSS.n1377 4.5005
R27680 DVSS.n1386 DVSS.n1364 4.5005
R27681 DVSS.n1386 DVSS.n1376 4.5005
R27682 DVSS.n1386 DVSS.n1365 4.5005
R27683 DVSS.n1386 DVSS.n1375 4.5005
R27684 DVSS.n1386 DVSS.n1366 4.5005
R27685 DVSS.n1386 DVSS.n1374 4.5005
R27686 DVSS.n1386 DVSS.n1367 4.5005
R27687 DVSS.n1386 DVSS.n1373 4.5005
R27688 DVSS.n1386 DVSS.n1368 4.5005
R27689 DVSS.n1386 DVSS.n1372 4.5005
R27690 DVSS.n1386 DVSS.n1369 4.5005
R27691 DVSS.n1386 DVSS.n1371 4.5005
R27692 DVSS.n22123 DVSS.n1377 4.5005
R27693 DVSS.n22123 DVSS.n1364 4.5005
R27694 DVSS.n22123 DVSS.n1376 4.5005
R27695 DVSS.n22123 DVSS.n1365 4.5005
R27696 DVSS.n22123 DVSS.n1375 4.5005
R27697 DVSS.n22123 DVSS.n1366 4.5005
R27698 DVSS.n22123 DVSS.n1374 4.5005
R27699 DVSS.n22123 DVSS.n1367 4.5005
R27700 DVSS.n22123 DVSS.n1373 4.5005
R27701 DVSS.n22123 DVSS.n1368 4.5005
R27702 DVSS.n22123 DVSS.n1372 4.5005
R27703 DVSS.n22123 DVSS.n1369 4.5005
R27704 DVSS.n22123 DVSS.n1371 4.5005
R27705 DVSS.n1387 DVSS.n1377 4.5005
R27706 DVSS.n1387 DVSS.n1364 4.5005
R27707 DVSS.n1387 DVSS.n1376 4.5005
R27708 DVSS.n1387 DVSS.n1365 4.5005
R27709 DVSS.n1387 DVSS.n1375 4.5005
R27710 DVSS.n1387 DVSS.n1366 4.5005
R27711 DVSS.n1387 DVSS.n1374 4.5005
R27712 DVSS.n1387 DVSS.n1367 4.5005
R27713 DVSS.n1387 DVSS.n1373 4.5005
R27714 DVSS.n1387 DVSS.n1368 4.5005
R27715 DVSS.n1387 DVSS.n1372 4.5005
R27716 DVSS.n1387 DVSS.n1369 4.5005
R27717 DVSS.n1387 DVSS.n1371 4.5005
R27718 DVSS.n22122 DVSS.n1377 4.5005
R27719 DVSS.n22122 DVSS.n1364 4.5005
R27720 DVSS.n22122 DVSS.n1376 4.5005
R27721 DVSS.n22122 DVSS.n1365 4.5005
R27722 DVSS.n22122 DVSS.n1375 4.5005
R27723 DVSS.n22122 DVSS.n1366 4.5005
R27724 DVSS.n22122 DVSS.n1374 4.5005
R27725 DVSS.n22122 DVSS.n1367 4.5005
R27726 DVSS.n22122 DVSS.n1373 4.5005
R27727 DVSS.n22122 DVSS.n1368 4.5005
R27728 DVSS.n22122 DVSS.n1372 4.5005
R27729 DVSS.n22122 DVSS.n1369 4.5005
R27730 DVSS.n22122 DVSS.n1371 4.5005
R27731 DVSS.n22120 DVSS.n1377 4.5005
R27732 DVSS.n22120 DVSS.n1364 4.5005
R27733 DVSS.n22120 DVSS.n1376 4.5005
R27734 DVSS.n22120 DVSS.n1365 4.5005
R27735 DVSS.n22120 DVSS.n1375 4.5005
R27736 DVSS.n22120 DVSS.n1366 4.5005
R27737 DVSS.n22120 DVSS.n1374 4.5005
R27738 DVSS.n22120 DVSS.n1367 4.5005
R27739 DVSS.n22120 DVSS.n1373 4.5005
R27740 DVSS.n22120 DVSS.n1368 4.5005
R27741 DVSS.n22120 DVSS.n1372 4.5005
R27742 DVSS.n22120 DVSS.n1369 4.5005
R27743 DVSS.n22120 DVSS.n1371 4.5005
R27744 DVSS.n1392 DVSS.n1377 4.5005
R27745 DVSS.n1392 DVSS.n1364 4.5005
R27746 DVSS.n1392 DVSS.n1376 4.5005
R27747 DVSS.n1392 DVSS.n1365 4.5005
R27748 DVSS.n1392 DVSS.n1375 4.5005
R27749 DVSS.n1392 DVSS.n1366 4.5005
R27750 DVSS.n1392 DVSS.n1374 4.5005
R27751 DVSS.n1392 DVSS.n1367 4.5005
R27752 DVSS.n1392 DVSS.n1373 4.5005
R27753 DVSS.n1392 DVSS.n1368 4.5005
R27754 DVSS.n1392 DVSS.n1372 4.5005
R27755 DVSS.n1392 DVSS.n1369 4.5005
R27756 DVSS.n1392 DVSS.n1371 4.5005
R27757 DVSS.n21858 DVSS.n870 4.5005
R27758 DVSS.n21860 DVSS.n870 4.5005
R27759 DVSS.n21857 DVSS.n870 4.5005
R27760 DVSS.n21861 DVSS.n870 4.5005
R27761 DVSS.n21856 DVSS.n870 4.5005
R27762 DVSS.n21865 DVSS.n870 4.5005
R27763 DVSS.n21854 DVSS.n870 4.5005
R27764 DVSS.n21867 DVSS.n870 4.5005
R27765 DVSS.n21853 DVSS.n870 4.5005
R27766 DVSS.n21868 DVSS.n870 4.5005
R27767 DVSS.n21852 DVSS.n870 4.5005
R27768 DVSS.n21869 DVSS.n870 4.5005
R27769 DVSS.n21944 DVSS.n870 4.5005
R27770 DVSS.n21882 DVSS.n21858 4.5005
R27771 DVSS.n21882 DVSS.n21860 4.5005
R27772 DVSS.n21882 DVSS.n21857 4.5005
R27773 DVSS.n21882 DVSS.n21861 4.5005
R27774 DVSS.n21882 DVSS.n21856 4.5005
R27775 DVSS.n21882 DVSS.n21864 4.5005
R27776 DVSS.n21882 DVSS.n21855 4.5005
R27777 DVSS.n21882 DVSS.n21865 4.5005
R27778 DVSS.n21882 DVSS.n21854 4.5005
R27779 DVSS.n21882 DVSS.n21867 4.5005
R27780 DVSS.n21882 DVSS.n21853 4.5005
R27781 DVSS.n21882 DVSS.n21868 4.5005
R27782 DVSS.n21882 DVSS.n21869 4.5005
R27783 DVSS.n21944 DVSS.n21882 4.5005
R27784 DVSS.n21880 DVSS.n21858 4.5005
R27785 DVSS.n21880 DVSS.n21860 4.5005
R27786 DVSS.n21880 DVSS.n21857 4.5005
R27787 DVSS.n21880 DVSS.n21861 4.5005
R27788 DVSS.n21880 DVSS.n21856 4.5005
R27789 DVSS.n21880 DVSS.n21864 4.5005
R27790 DVSS.n21880 DVSS.n21855 4.5005
R27791 DVSS.n21880 DVSS.n21865 4.5005
R27792 DVSS.n21880 DVSS.n21854 4.5005
R27793 DVSS.n21880 DVSS.n21867 4.5005
R27794 DVSS.n21880 DVSS.n21853 4.5005
R27795 DVSS.n21880 DVSS.n21868 4.5005
R27796 DVSS.n21944 DVSS.n21880 4.5005
R27797 DVSS.n21889 DVSS.n21858 4.5005
R27798 DVSS.n21889 DVSS.n21860 4.5005
R27799 DVSS.n21889 DVSS.n21857 4.5005
R27800 DVSS.n21889 DVSS.n21861 4.5005
R27801 DVSS.n21889 DVSS.n21856 4.5005
R27802 DVSS.n21889 DVSS.n21864 4.5005
R27803 DVSS.n21889 DVSS.n21855 4.5005
R27804 DVSS.n21889 DVSS.n21865 4.5005
R27805 DVSS.n21889 DVSS.n21854 4.5005
R27806 DVSS.n21889 DVSS.n21867 4.5005
R27807 DVSS.n21889 DVSS.n21853 4.5005
R27808 DVSS.n21889 DVSS.n21868 4.5005
R27809 DVSS.n21889 DVSS.n21852 4.5005
R27810 DVSS.n21889 DVSS.n21869 4.5005
R27811 DVSS.n21944 DVSS.n21889 4.5005
R27812 DVSS.n21879 DVSS.n21858 4.5005
R27813 DVSS.n21879 DVSS.n21860 4.5005
R27814 DVSS.n21879 DVSS.n21857 4.5005
R27815 DVSS.n21879 DVSS.n21861 4.5005
R27816 DVSS.n21879 DVSS.n21856 4.5005
R27817 DVSS.n21879 DVSS.n21864 4.5005
R27818 DVSS.n21879 DVSS.n21855 4.5005
R27819 DVSS.n21879 DVSS.n21865 4.5005
R27820 DVSS.n21879 DVSS.n21854 4.5005
R27821 DVSS.n21879 DVSS.n21867 4.5005
R27822 DVSS.n21879 DVSS.n21853 4.5005
R27823 DVSS.n21879 DVSS.n21868 4.5005
R27824 DVSS.n21879 DVSS.n21869 4.5005
R27825 DVSS.n21944 DVSS.n21879 4.5005
R27826 DVSS.n21891 DVSS.n21858 4.5005
R27827 DVSS.n21891 DVSS.n21860 4.5005
R27828 DVSS.n21891 DVSS.n21857 4.5005
R27829 DVSS.n21891 DVSS.n21861 4.5005
R27830 DVSS.n21891 DVSS.n21856 4.5005
R27831 DVSS.n21891 DVSS.n21864 4.5005
R27832 DVSS.n21891 DVSS.n21855 4.5005
R27833 DVSS.n21891 DVSS.n21865 4.5005
R27834 DVSS.n21891 DVSS.n21854 4.5005
R27835 DVSS.n21891 DVSS.n21867 4.5005
R27836 DVSS.n21891 DVSS.n21853 4.5005
R27837 DVSS.n21891 DVSS.n21868 4.5005
R27838 DVSS.n21891 DVSS.n21869 4.5005
R27839 DVSS.n21944 DVSS.n21891 4.5005
R27840 DVSS.n21878 DVSS.n21858 4.5005
R27841 DVSS.n21878 DVSS.n21860 4.5005
R27842 DVSS.n21878 DVSS.n21857 4.5005
R27843 DVSS.n21878 DVSS.n21861 4.5005
R27844 DVSS.n21878 DVSS.n21856 4.5005
R27845 DVSS.n21878 DVSS.n21864 4.5005
R27846 DVSS.n21878 DVSS.n21855 4.5005
R27847 DVSS.n21878 DVSS.n21865 4.5005
R27848 DVSS.n21878 DVSS.n21854 4.5005
R27849 DVSS.n21878 DVSS.n21867 4.5005
R27850 DVSS.n21878 DVSS.n21853 4.5005
R27851 DVSS.n21878 DVSS.n21868 4.5005
R27852 DVSS.n21878 DVSS.n21852 4.5005
R27853 DVSS.n21878 DVSS.n21869 4.5005
R27854 DVSS.n21944 DVSS.n21878 4.5005
R27855 DVSS.n21899 DVSS.n21858 4.5005
R27856 DVSS.n21899 DVSS.n21860 4.5005
R27857 DVSS.n21899 DVSS.n21857 4.5005
R27858 DVSS.n21899 DVSS.n21861 4.5005
R27859 DVSS.n21899 DVSS.n21856 4.5005
R27860 DVSS.n21899 DVSS.n21864 4.5005
R27861 DVSS.n21899 DVSS.n21855 4.5005
R27862 DVSS.n21899 DVSS.n21865 4.5005
R27863 DVSS.n21899 DVSS.n21854 4.5005
R27864 DVSS.n21899 DVSS.n21867 4.5005
R27865 DVSS.n21899 DVSS.n21853 4.5005
R27866 DVSS.n21899 DVSS.n21868 4.5005
R27867 DVSS.n21899 DVSS.n21852 4.5005
R27868 DVSS.n21899 DVSS.n21869 4.5005
R27869 DVSS.n21944 DVSS.n21899 4.5005
R27870 DVSS.n21877 DVSS.n21858 4.5005
R27871 DVSS.n21877 DVSS.n21860 4.5005
R27872 DVSS.n21877 DVSS.n21857 4.5005
R27873 DVSS.n21877 DVSS.n21861 4.5005
R27874 DVSS.n21877 DVSS.n21856 4.5005
R27875 DVSS.n21877 DVSS.n21864 4.5005
R27876 DVSS.n21877 DVSS.n21855 4.5005
R27877 DVSS.n21877 DVSS.n21865 4.5005
R27878 DVSS.n21877 DVSS.n21854 4.5005
R27879 DVSS.n21877 DVSS.n21867 4.5005
R27880 DVSS.n21877 DVSS.n21853 4.5005
R27881 DVSS.n21877 DVSS.n21868 4.5005
R27882 DVSS.n21877 DVSS.n21869 4.5005
R27883 DVSS.n21944 DVSS.n21877 4.5005
R27884 DVSS.n21901 DVSS.n21858 4.5005
R27885 DVSS.n21901 DVSS.n21860 4.5005
R27886 DVSS.n21901 DVSS.n21857 4.5005
R27887 DVSS.n21901 DVSS.n21861 4.5005
R27888 DVSS.n21901 DVSS.n21856 4.5005
R27889 DVSS.n21901 DVSS.n21864 4.5005
R27890 DVSS.n21901 DVSS.n21855 4.5005
R27891 DVSS.n21901 DVSS.n21865 4.5005
R27892 DVSS.n21901 DVSS.n21854 4.5005
R27893 DVSS.n21901 DVSS.n21867 4.5005
R27894 DVSS.n21901 DVSS.n21853 4.5005
R27895 DVSS.n21901 DVSS.n21868 4.5005
R27896 DVSS.n21901 DVSS.n21869 4.5005
R27897 DVSS.n21944 DVSS.n21901 4.5005
R27898 DVSS.n21876 DVSS.n21858 4.5005
R27899 DVSS.n21876 DVSS.n21860 4.5005
R27900 DVSS.n21876 DVSS.n21857 4.5005
R27901 DVSS.n21876 DVSS.n21861 4.5005
R27902 DVSS.n21876 DVSS.n21856 4.5005
R27903 DVSS.n21876 DVSS.n21864 4.5005
R27904 DVSS.n21876 DVSS.n21855 4.5005
R27905 DVSS.n21876 DVSS.n21865 4.5005
R27906 DVSS.n21876 DVSS.n21854 4.5005
R27907 DVSS.n21876 DVSS.n21867 4.5005
R27908 DVSS.n21876 DVSS.n21853 4.5005
R27909 DVSS.n21876 DVSS.n21868 4.5005
R27910 DVSS.n21876 DVSS.n21852 4.5005
R27911 DVSS.n21876 DVSS.n21869 4.5005
R27912 DVSS.n21944 DVSS.n21876 4.5005
R27913 DVSS.n21909 DVSS.n21858 4.5005
R27914 DVSS.n21909 DVSS.n21860 4.5005
R27915 DVSS.n21909 DVSS.n21857 4.5005
R27916 DVSS.n21909 DVSS.n21861 4.5005
R27917 DVSS.n21909 DVSS.n21856 4.5005
R27918 DVSS.n21909 DVSS.n21864 4.5005
R27919 DVSS.n21909 DVSS.n21855 4.5005
R27920 DVSS.n21909 DVSS.n21865 4.5005
R27921 DVSS.n21909 DVSS.n21854 4.5005
R27922 DVSS.n21909 DVSS.n21867 4.5005
R27923 DVSS.n21909 DVSS.n21853 4.5005
R27924 DVSS.n21909 DVSS.n21868 4.5005
R27925 DVSS.n21909 DVSS.n21852 4.5005
R27926 DVSS.n21909 DVSS.n21869 4.5005
R27927 DVSS.n21944 DVSS.n21909 4.5005
R27928 DVSS.n21875 DVSS.n21858 4.5005
R27929 DVSS.n21875 DVSS.n21860 4.5005
R27930 DVSS.n21875 DVSS.n21857 4.5005
R27931 DVSS.n21875 DVSS.n21861 4.5005
R27932 DVSS.n21875 DVSS.n21856 4.5005
R27933 DVSS.n21875 DVSS.n21864 4.5005
R27934 DVSS.n21875 DVSS.n21855 4.5005
R27935 DVSS.n21875 DVSS.n21865 4.5005
R27936 DVSS.n21875 DVSS.n21854 4.5005
R27937 DVSS.n21875 DVSS.n21867 4.5005
R27938 DVSS.n21875 DVSS.n21853 4.5005
R27939 DVSS.n21875 DVSS.n21868 4.5005
R27940 DVSS.n21875 DVSS.n21869 4.5005
R27941 DVSS.n21944 DVSS.n21875 4.5005
R27942 DVSS.n21911 DVSS.n21858 4.5005
R27943 DVSS.n21911 DVSS.n21860 4.5005
R27944 DVSS.n21911 DVSS.n21857 4.5005
R27945 DVSS.n21911 DVSS.n21861 4.5005
R27946 DVSS.n21911 DVSS.n21856 4.5005
R27947 DVSS.n21911 DVSS.n21864 4.5005
R27948 DVSS.n21911 DVSS.n21855 4.5005
R27949 DVSS.n21911 DVSS.n21865 4.5005
R27950 DVSS.n21911 DVSS.n21854 4.5005
R27951 DVSS.n21911 DVSS.n21867 4.5005
R27952 DVSS.n21911 DVSS.n21853 4.5005
R27953 DVSS.n21911 DVSS.n21868 4.5005
R27954 DVSS.n21911 DVSS.n21869 4.5005
R27955 DVSS.n21944 DVSS.n21911 4.5005
R27956 DVSS.n21874 DVSS.n21858 4.5005
R27957 DVSS.n21874 DVSS.n21860 4.5005
R27958 DVSS.n21874 DVSS.n21857 4.5005
R27959 DVSS.n21874 DVSS.n21861 4.5005
R27960 DVSS.n21874 DVSS.n21856 4.5005
R27961 DVSS.n21874 DVSS.n21864 4.5005
R27962 DVSS.n21874 DVSS.n21855 4.5005
R27963 DVSS.n21874 DVSS.n21865 4.5005
R27964 DVSS.n21874 DVSS.n21854 4.5005
R27965 DVSS.n21874 DVSS.n21867 4.5005
R27966 DVSS.n21874 DVSS.n21853 4.5005
R27967 DVSS.n21874 DVSS.n21868 4.5005
R27968 DVSS.n21874 DVSS.n21852 4.5005
R27969 DVSS.n21874 DVSS.n21869 4.5005
R27970 DVSS.n21944 DVSS.n21874 4.5005
R27971 DVSS.n21919 DVSS.n21858 4.5005
R27972 DVSS.n21919 DVSS.n21860 4.5005
R27973 DVSS.n21919 DVSS.n21857 4.5005
R27974 DVSS.n21919 DVSS.n21861 4.5005
R27975 DVSS.n21919 DVSS.n21856 4.5005
R27976 DVSS.n21919 DVSS.n21864 4.5005
R27977 DVSS.n21919 DVSS.n21855 4.5005
R27978 DVSS.n21919 DVSS.n21865 4.5005
R27979 DVSS.n21919 DVSS.n21854 4.5005
R27980 DVSS.n21919 DVSS.n21867 4.5005
R27981 DVSS.n21919 DVSS.n21853 4.5005
R27982 DVSS.n21919 DVSS.n21868 4.5005
R27983 DVSS.n21919 DVSS.n21852 4.5005
R27984 DVSS.n21919 DVSS.n21869 4.5005
R27985 DVSS.n21944 DVSS.n21919 4.5005
R27986 DVSS.n21873 DVSS.n21858 4.5005
R27987 DVSS.n21873 DVSS.n21860 4.5005
R27988 DVSS.n21873 DVSS.n21857 4.5005
R27989 DVSS.n21873 DVSS.n21861 4.5005
R27990 DVSS.n21873 DVSS.n21856 4.5005
R27991 DVSS.n21873 DVSS.n21864 4.5005
R27992 DVSS.n21873 DVSS.n21855 4.5005
R27993 DVSS.n21873 DVSS.n21865 4.5005
R27994 DVSS.n21873 DVSS.n21854 4.5005
R27995 DVSS.n21873 DVSS.n21867 4.5005
R27996 DVSS.n21873 DVSS.n21853 4.5005
R27997 DVSS.n21873 DVSS.n21868 4.5005
R27998 DVSS.n21873 DVSS.n21869 4.5005
R27999 DVSS.n21944 DVSS.n21873 4.5005
R28000 DVSS.n21921 DVSS.n21858 4.5005
R28001 DVSS.n21921 DVSS.n21860 4.5005
R28002 DVSS.n21921 DVSS.n21857 4.5005
R28003 DVSS.n21921 DVSS.n21861 4.5005
R28004 DVSS.n21921 DVSS.n21856 4.5005
R28005 DVSS.n21921 DVSS.n21864 4.5005
R28006 DVSS.n21921 DVSS.n21855 4.5005
R28007 DVSS.n21921 DVSS.n21865 4.5005
R28008 DVSS.n21921 DVSS.n21854 4.5005
R28009 DVSS.n21921 DVSS.n21867 4.5005
R28010 DVSS.n21921 DVSS.n21853 4.5005
R28011 DVSS.n21921 DVSS.n21868 4.5005
R28012 DVSS.n21921 DVSS.n21869 4.5005
R28013 DVSS.n21944 DVSS.n21921 4.5005
R28014 DVSS.n21872 DVSS.n21858 4.5005
R28015 DVSS.n21872 DVSS.n21860 4.5005
R28016 DVSS.n21872 DVSS.n21857 4.5005
R28017 DVSS.n21872 DVSS.n21861 4.5005
R28018 DVSS.n21872 DVSS.n21856 4.5005
R28019 DVSS.n21872 DVSS.n21864 4.5005
R28020 DVSS.n21872 DVSS.n21855 4.5005
R28021 DVSS.n21872 DVSS.n21865 4.5005
R28022 DVSS.n21872 DVSS.n21854 4.5005
R28023 DVSS.n21872 DVSS.n21867 4.5005
R28024 DVSS.n21872 DVSS.n21853 4.5005
R28025 DVSS.n21872 DVSS.n21868 4.5005
R28026 DVSS.n21872 DVSS.n21852 4.5005
R28027 DVSS.n21872 DVSS.n21869 4.5005
R28028 DVSS.n21944 DVSS.n21872 4.5005
R28029 DVSS.n21941 DVSS.n21858 4.5005
R28030 DVSS.n21941 DVSS.n21860 4.5005
R28031 DVSS.n21941 DVSS.n21857 4.5005
R28032 DVSS.n21941 DVSS.n21861 4.5005
R28033 DVSS.n21941 DVSS.n21856 4.5005
R28034 DVSS.n21941 DVSS.n21864 4.5005
R28035 DVSS.n21941 DVSS.n21855 4.5005
R28036 DVSS.n21941 DVSS.n21865 4.5005
R28037 DVSS.n21941 DVSS.n21854 4.5005
R28038 DVSS.n21941 DVSS.n21867 4.5005
R28039 DVSS.n21941 DVSS.n21853 4.5005
R28040 DVSS.n21941 DVSS.n21868 4.5005
R28041 DVSS.n21941 DVSS.n21852 4.5005
R28042 DVSS.n21941 DVSS.n21869 4.5005
R28043 DVSS.n21944 DVSS.n21941 4.5005
R28044 DVSS.n21871 DVSS.n21858 4.5005
R28045 DVSS.n21871 DVSS.n21860 4.5005
R28046 DVSS.n21871 DVSS.n21857 4.5005
R28047 DVSS.n21871 DVSS.n21861 4.5005
R28048 DVSS.n21871 DVSS.n21856 4.5005
R28049 DVSS.n21871 DVSS.n21864 4.5005
R28050 DVSS.n21871 DVSS.n21855 4.5005
R28051 DVSS.n21871 DVSS.n21865 4.5005
R28052 DVSS.n21871 DVSS.n21854 4.5005
R28053 DVSS.n21871 DVSS.n21867 4.5005
R28054 DVSS.n21871 DVSS.n21853 4.5005
R28055 DVSS.n21871 DVSS.n21868 4.5005
R28056 DVSS.n21871 DVSS.n21869 4.5005
R28057 DVSS.n21944 DVSS.n21871 4.5005
R28058 DVSS.n21943 DVSS.n21858 4.5005
R28059 DVSS.n21943 DVSS.n21860 4.5005
R28060 DVSS.n21943 DVSS.n21857 4.5005
R28061 DVSS.n21943 DVSS.n21861 4.5005
R28062 DVSS.n21943 DVSS.n21856 4.5005
R28063 DVSS.n21943 DVSS.n21864 4.5005
R28064 DVSS.n21943 DVSS.n21855 4.5005
R28065 DVSS.n21943 DVSS.n21865 4.5005
R28066 DVSS.n21943 DVSS.n21854 4.5005
R28067 DVSS.n21943 DVSS.n21867 4.5005
R28068 DVSS.n21943 DVSS.n21853 4.5005
R28069 DVSS.n21943 DVSS.n21868 4.5005
R28070 DVSS.n21943 DVSS.n21869 4.5005
R28071 DVSS.n21944 DVSS.n21943 4.5005
R28072 DVSS.n21945 DVSS.n21858 4.5005
R28073 DVSS.n21945 DVSS.n21860 4.5005
R28074 DVSS.n21945 DVSS.n21857 4.5005
R28075 DVSS.n21945 DVSS.n21861 4.5005
R28076 DVSS.n21945 DVSS.n21856 4.5005
R28077 DVSS.n21945 DVSS.n21864 4.5005
R28078 DVSS.n21945 DVSS.n21855 4.5005
R28079 DVSS.n21945 DVSS.n21865 4.5005
R28080 DVSS.n21945 DVSS.n21854 4.5005
R28081 DVSS.n21945 DVSS.n21867 4.5005
R28082 DVSS.n21945 DVSS.n21853 4.5005
R28083 DVSS.n21945 DVSS.n21868 4.5005
R28084 DVSS.n21945 DVSS.n21852 4.5005
R28085 DVSS.n21945 DVSS.n21869 4.5005
R28086 DVSS.n21945 DVSS.n21944 4.5005
R28087 DVSS.n21858 DVSS.n21850 4.5005
R28088 DVSS.n21860 DVSS.n21850 4.5005
R28089 DVSS.n21857 DVSS.n21850 4.5005
R28090 DVSS.n21861 DVSS.n21850 4.5005
R28091 DVSS.n21856 DVSS.n21850 4.5005
R28092 DVSS.n21864 DVSS.n21850 4.5005
R28093 DVSS.n21855 DVSS.n21850 4.5005
R28094 DVSS.n21865 DVSS.n21850 4.5005
R28095 DVSS.n21854 DVSS.n21850 4.5005
R28096 DVSS.n21867 DVSS.n21850 4.5005
R28097 DVSS.n21853 DVSS.n21850 4.5005
R28098 DVSS.n21868 DVSS.n21850 4.5005
R28099 DVSS.n21852 DVSS.n21850 4.5005
R28100 DVSS.n21869 DVSS.n21850 4.5005
R28101 DVSS.n21932 DVSS.n21850 4.5005
R28102 DVSS.n21944 DVSS.n21850 4.5005
R28103 DVSS.n21628 DVSS.n21590 4.5005
R28104 DVSS.n21630 DVSS.n21590 4.5005
R28105 DVSS.n21626 DVSS.n21590 4.5005
R28106 DVSS.n22075 DVSS.n21590 4.5005
R28107 DVSS.n21625 DVSS.n21590 4.5005
R28108 DVSS.n21633 DVSS.n21590 4.5005
R28109 DVSS.n21624 DVSS.n21590 4.5005
R28110 DVSS.n21634 DVSS.n21590 4.5005
R28111 DVSS.n21623 DVSS.n21590 4.5005
R28112 DVSS.n21637 DVSS.n21590 4.5005
R28113 DVSS.n22073 DVSS.n21590 4.5005
R28114 DVSS.n21628 DVSS.n21592 4.5005
R28115 DVSS.n21630 DVSS.n21592 4.5005
R28116 DVSS.n21626 DVSS.n21592 4.5005
R28117 DVSS.n21632 DVSS.n21592 4.5005
R28118 DVSS.n21592 DVSS.n1463 4.5005
R28119 DVSS.n22075 DVSS.n21592 4.5005
R28120 DVSS.n21625 DVSS.n21592 4.5005
R28121 DVSS.n21633 DVSS.n21592 4.5005
R28122 DVSS.n21624 DVSS.n21592 4.5005
R28123 DVSS.n21634 DVSS.n21592 4.5005
R28124 DVSS.n21623 DVSS.n21592 4.5005
R28125 DVSS.n21636 DVSS.n21592 4.5005
R28126 DVSS.n21637 DVSS.n21592 4.5005
R28127 DVSS.n22073 DVSS.n21592 4.5005
R28128 DVSS.n21628 DVSS.n21567 4.5005
R28129 DVSS.n21630 DVSS.n21567 4.5005
R28130 DVSS.n21626 DVSS.n21567 4.5005
R28131 DVSS.n21632 DVSS.n21567 4.5005
R28132 DVSS.n21567 DVSS.n1463 4.5005
R28133 DVSS.n22075 DVSS.n21567 4.5005
R28134 DVSS.n21625 DVSS.n21567 4.5005
R28135 DVSS.n21633 DVSS.n21567 4.5005
R28136 DVSS.n21624 DVSS.n21567 4.5005
R28137 DVSS.n21634 DVSS.n21567 4.5005
R28138 DVSS.n21623 DVSS.n21567 4.5005
R28139 DVSS.n21636 DVSS.n21567 4.5005
R28140 DVSS.n21637 DVSS.n21567 4.5005
R28141 DVSS.n21615 DVSS.n21567 4.5005
R28142 DVSS.n22073 DVSS.n21567 4.5005
R28143 DVSS.n21628 DVSS.n21593 4.5005
R28144 DVSS.n21630 DVSS.n21593 4.5005
R28145 DVSS.n21626 DVSS.n21593 4.5005
R28146 DVSS.n21632 DVSS.n21593 4.5005
R28147 DVSS.n21593 DVSS.n1463 4.5005
R28148 DVSS.n22075 DVSS.n21593 4.5005
R28149 DVSS.n21625 DVSS.n21593 4.5005
R28150 DVSS.n21633 DVSS.n21593 4.5005
R28151 DVSS.n21624 DVSS.n21593 4.5005
R28152 DVSS.n21634 DVSS.n21593 4.5005
R28153 DVSS.n21623 DVSS.n21593 4.5005
R28154 DVSS.n21636 DVSS.n21593 4.5005
R28155 DVSS.n21622 DVSS.n21593 4.5005
R28156 DVSS.n21637 DVSS.n21593 4.5005
R28157 DVSS.n22073 DVSS.n21593 4.5005
R28158 DVSS.n21628 DVSS.n21566 4.5005
R28159 DVSS.n21630 DVSS.n21566 4.5005
R28160 DVSS.n21626 DVSS.n21566 4.5005
R28161 DVSS.n21632 DVSS.n21566 4.5005
R28162 DVSS.n21566 DVSS.n1463 4.5005
R28163 DVSS.n22075 DVSS.n21566 4.5005
R28164 DVSS.n21625 DVSS.n21566 4.5005
R28165 DVSS.n21633 DVSS.n21566 4.5005
R28166 DVSS.n21624 DVSS.n21566 4.5005
R28167 DVSS.n21634 DVSS.n21566 4.5005
R28168 DVSS.n21623 DVSS.n21566 4.5005
R28169 DVSS.n21636 DVSS.n21566 4.5005
R28170 DVSS.n21637 DVSS.n21566 4.5005
R28171 DVSS.n22073 DVSS.n21566 4.5005
R28172 DVSS.n21628 DVSS.n21594 4.5005
R28173 DVSS.n21630 DVSS.n21594 4.5005
R28174 DVSS.n21626 DVSS.n21594 4.5005
R28175 DVSS.n21632 DVSS.n21594 4.5005
R28176 DVSS.n21594 DVSS.n1463 4.5005
R28177 DVSS.n22075 DVSS.n21594 4.5005
R28178 DVSS.n21625 DVSS.n21594 4.5005
R28179 DVSS.n21633 DVSS.n21594 4.5005
R28180 DVSS.n21624 DVSS.n21594 4.5005
R28181 DVSS.n21634 DVSS.n21594 4.5005
R28182 DVSS.n21623 DVSS.n21594 4.5005
R28183 DVSS.n21636 DVSS.n21594 4.5005
R28184 DVSS.n21637 DVSS.n21594 4.5005
R28185 DVSS.n22073 DVSS.n21594 4.5005
R28186 DVSS.n21628 DVSS.n21565 4.5005
R28187 DVSS.n21630 DVSS.n21565 4.5005
R28188 DVSS.n21626 DVSS.n21565 4.5005
R28189 DVSS.n21632 DVSS.n21565 4.5005
R28190 DVSS.n21565 DVSS.n1463 4.5005
R28191 DVSS.n22075 DVSS.n21565 4.5005
R28192 DVSS.n21625 DVSS.n21565 4.5005
R28193 DVSS.n21633 DVSS.n21565 4.5005
R28194 DVSS.n21624 DVSS.n21565 4.5005
R28195 DVSS.n21634 DVSS.n21565 4.5005
R28196 DVSS.n21623 DVSS.n21565 4.5005
R28197 DVSS.n21636 DVSS.n21565 4.5005
R28198 DVSS.n21622 DVSS.n21565 4.5005
R28199 DVSS.n21637 DVSS.n21565 4.5005
R28200 DVSS.n22073 DVSS.n21565 4.5005
R28201 DVSS.n21628 DVSS.n21595 4.5005
R28202 DVSS.n21630 DVSS.n21595 4.5005
R28203 DVSS.n21626 DVSS.n21595 4.5005
R28204 DVSS.n21632 DVSS.n21595 4.5005
R28205 DVSS.n21595 DVSS.n1463 4.5005
R28206 DVSS.n22075 DVSS.n21595 4.5005
R28207 DVSS.n21625 DVSS.n21595 4.5005
R28208 DVSS.n21633 DVSS.n21595 4.5005
R28209 DVSS.n21624 DVSS.n21595 4.5005
R28210 DVSS.n21634 DVSS.n21595 4.5005
R28211 DVSS.n21623 DVSS.n21595 4.5005
R28212 DVSS.n21636 DVSS.n21595 4.5005
R28213 DVSS.n21622 DVSS.n21595 4.5005
R28214 DVSS.n21637 DVSS.n21595 4.5005
R28215 DVSS.n22073 DVSS.n21595 4.5005
R28216 DVSS.n21628 DVSS.n21564 4.5005
R28217 DVSS.n21630 DVSS.n21564 4.5005
R28218 DVSS.n21626 DVSS.n21564 4.5005
R28219 DVSS.n21632 DVSS.n21564 4.5005
R28220 DVSS.n21564 DVSS.n1463 4.5005
R28221 DVSS.n22075 DVSS.n21564 4.5005
R28222 DVSS.n21625 DVSS.n21564 4.5005
R28223 DVSS.n21633 DVSS.n21564 4.5005
R28224 DVSS.n21624 DVSS.n21564 4.5005
R28225 DVSS.n21634 DVSS.n21564 4.5005
R28226 DVSS.n21623 DVSS.n21564 4.5005
R28227 DVSS.n21636 DVSS.n21564 4.5005
R28228 DVSS.n21637 DVSS.n21564 4.5005
R28229 DVSS.n22073 DVSS.n21564 4.5005
R28230 DVSS.n21628 DVSS.n21596 4.5005
R28231 DVSS.n21630 DVSS.n21596 4.5005
R28232 DVSS.n21626 DVSS.n21596 4.5005
R28233 DVSS.n21632 DVSS.n21596 4.5005
R28234 DVSS.n21596 DVSS.n1463 4.5005
R28235 DVSS.n22075 DVSS.n21596 4.5005
R28236 DVSS.n21625 DVSS.n21596 4.5005
R28237 DVSS.n21633 DVSS.n21596 4.5005
R28238 DVSS.n21624 DVSS.n21596 4.5005
R28239 DVSS.n21634 DVSS.n21596 4.5005
R28240 DVSS.n21623 DVSS.n21596 4.5005
R28241 DVSS.n21636 DVSS.n21596 4.5005
R28242 DVSS.n21637 DVSS.n21596 4.5005
R28243 DVSS.n22073 DVSS.n21596 4.5005
R28244 DVSS.n21628 DVSS.n21563 4.5005
R28245 DVSS.n21630 DVSS.n21563 4.5005
R28246 DVSS.n21626 DVSS.n21563 4.5005
R28247 DVSS.n21632 DVSS.n21563 4.5005
R28248 DVSS.n21563 DVSS.n1463 4.5005
R28249 DVSS.n22075 DVSS.n21563 4.5005
R28250 DVSS.n21625 DVSS.n21563 4.5005
R28251 DVSS.n21633 DVSS.n21563 4.5005
R28252 DVSS.n21624 DVSS.n21563 4.5005
R28253 DVSS.n21634 DVSS.n21563 4.5005
R28254 DVSS.n21623 DVSS.n21563 4.5005
R28255 DVSS.n21636 DVSS.n21563 4.5005
R28256 DVSS.n21622 DVSS.n21563 4.5005
R28257 DVSS.n21637 DVSS.n21563 4.5005
R28258 DVSS.n22073 DVSS.n21563 4.5005
R28259 DVSS.n21628 DVSS.n21597 4.5005
R28260 DVSS.n21630 DVSS.n21597 4.5005
R28261 DVSS.n21626 DVSS.n21597 4.5005
R28262 DVSS.n21632 DVSS.n21597 4.5005
R28263 DVSS.n21597 DVSS.n1463 4.5005
R28264 DVSS.n22075 DVSS.n21597 4.5005
R28265 DVSS.n21625 DVSS.n21597 4.5005
R28266 DVSS.n21633 DVSS.n21597 4.5005
R28267 DVSS.n21624 DVSS.n21597 4.5005
R28268 DVSS.n21634 DVSS.n21597 4.5005
R28269 DVSS.n21623 DVSS.n21597 4.5005
R28270 DVSS.n21636 DVSS.n21597 4.5005
R28271 DVSS.n21622 DVSS.n21597 4.5005
R28272 DVSS.n21637 DVSS.n21597 4.5005
R28273 DVSS.n22073 DVSS.n21597 4.5005
R28274 DVSS.n21628 DVSS.n21562 4.5005
R28275 DVSS.n21630 DVSS.n21562 4.5005
R28276 DVSS.n21626 DVSS.n21562 4.5005
R28277 DVSS.n21632 DVSS.n21562 4.5005
R28278 DVSS.n21562 DVSS.n1463 4.5005
R28279 DVSS.n22075 DVSS.n21562 4.5005
R28280 DVSS.n21625 DVSS.n21562 4.5005
R28281 DVSS.n21633 DVSS.n21562 4.5005
R28282 DVSS.n21624 DVSS.n21562 4.5005
R28283 DVSS.n21634 DVSS.n21562 4.5005
R28284 DVSS.n21623 DVSS.n21562 4.5005
R28285 DVSS.n21636 DVSS.n21562 4.5005
R28286 DVSS.n21637 DVSS.n21562 4.5005
R28287 DVSS.n22073 DVSS.n21562 4.5005
R28288 DVSS.n21628 DVSS.n21598 4.5005
R28289 DVSS.n21630 DVSS.n21598 4.5005
R28290 DVSS.n21626 DVSS.n21598 4.5005
R28291 DVSS.n21632 DVSS.n21598 4.5005
R28292 DVSS.n21598 DVSS.n1463 4.5005
R28293 DVSS.n22075 DVSS.n21598 4.5005
R28294 DVSS.n21625 DVSS.n21598 4.5005
R28295 DVSS.n21633 DVSS.n21598 4.5005
R28296 DVSS.n21624 DVSS.n21598 4.5005
R28297 DVSS.n21634 DVSS.n21598 4.5005
R28298 DVSS.n21623 DVSS.n21598 4.5005
R28299 DVSS.n21636 DVSS.n21598 4.5005
R28300 DVSS.n21637 DVSS.n21598 4.5005
R28301 DVSS.n22073 DVSS.n21598 4.5005
R28302 DVSS.n21628 DVSS.n21561 4.5005
R28303 DVSS.n21630 DVSS.n21561 4.5005
R28304 DVSS.n21626 DVSS.n21561 4.5005
R28305 DVSS.n21632 DVSS.n21561 4.5005
R28306 DVSS.n21561 DVSS.n1463 4.5005
R28307 DVSS.n22075 DVSS.n21561 4.5005
R28308 DVSS.n21625 DVSS.n21561 4.5005
R28309 DVSS.n21633 DVSS.n21561 4.5005
R28310 DVSS.n21624 DVSS.n21561 4.5005
R28311 DVSS.n21634 DVSS.n21561 4.5005
R28312 DVSS.n21623 DVSS.n21561 4.5005
R28313 DVSS.n21636 DVSS.n21561 4.5005
R28314 DVSS.n21622 DVSS.n21561 4.5005
R28315 DVSS.n21637 DVSS.n21561 4.5005
R28316 DVSS.n22073 DVSS.n21561 4.5005
R28317 DVSS.n21628 DVSS.n21599 4.5005
R28318 DVSS.n21630 DVSS.n21599 4.5005
R28319 DVSS.n21626 DVSS.n21599 4.5005
R28320 DVSS.n21632 DVSS.n21599 4.5005
R28321 DVSS.n21599 DVSS.n1463 4.5005
R28322 DVSS.n22075 DVSS.n21599 4.5005
R28323 DVSS.n21625 DVSS.n21599 4.5005
R28324 DVSS.n21633 DVSS.n21599 4.5005
R28325 DVSS.n21624 DVSS.n21599 4.5005
R28326 DVSS.n21634 DVSS.n21599 4.5005
R28327 DVSS.n21623 DVSS.n21599 4.5005
R28328 DVSS.n21636 DVSS.n21599 4.5005
R28329 DVSS.n21622 DVSS.n21599 4.5005
R28330 DVSS.n21637 DVSS.n21599 4.5005
R28331 DVSS.n22073 DVSS.n21599 4.5005
R28332 DVSS.n21628 DVSS.n21560 4.5005
R28333 DVSS.n21630 DVSS.n21560 4.5005
R28334 DVSS.n21626 DVSS.n21560 4.5005
R28335 DVSS.n21632 DVSS.n21560 4.5005
R28336 DVSS.n21560 DVSS.n1463 4.5005
R28337 DVSS.n22075 DVSS.n21560 4.5005
R28338 DVSS.n21625 DVSS.n21560 4.5005
R28339 DVSS.n21633 DVSS.n21560 4.5005
R28340 DVSS.n21624 DVSS.n21560 4.5005
R28341 DVSS.n21634 DVSS.n21560 4.5005
R28342 DVSS.n21623 DVSS.n21560 4.5005
R28343 DVSS.n21636 DVSS.n21560 4.5005
R28344 DVSS.n21637 DVSS.n21560 4.5005
R28345 DVSS.n22073 DVSS.n21560 4.5005
R28346 DVSS.n21628 DVSS.n21600 4.5005
R28347 DVSS.n21630 DVSS.n21600 4.5005
R28348 DVSS.n21626 DVSS.n21600 4.5005
R28349 DVSS.n21632 DVSS.n21600 4.5005
R28350 DVSS.n21600 DVSS.n1463 4.5005
R28351 DVSS.n22075 DVSS.n21600 4.5005
R28352 DVSS.n21625 DVSS.n21600 4.5005
R28353 DVSS.n21633 DVSS.n21600 4.5005
R28354 DVSS.n21624 DVSS.n21600 4.5005
R28355 DVSS.n21634 DVSS.n21600 4.5005
R28356 DVSS.n21623 DVSS.n21600 4.5005
R28357 DVSS.n21636 DVSS.n21600 4.5005
R28358 DVSS.n21637 DVSS.n21600 4.5005
R28359 DVSS.n22073 DVSS.n21600 4.5005
R28360 DVSS.n21628 DVSS.n21559 4.5005
R28361 DVSS.n21630 DVSS.n21559 4.5005
R28362 DVSS.n21626 DVSS.n21559 4.5005
R28363 DVSS.n21632 DVSS.n21559 4.5005
R28364 DVSS.n21559 DVSS.n1463 4.5005
R28365 DVSS.n22075 DVSS.n21559 4.5005
R28366 DVSS.n21625 DVSS.n21559 4.5005
R28367 DVSS.n21633 DVSS.n21559 4.5005
R28368 DVSS.n21624 DVSS.n21559 4.5005
R28369 DVSS.n21634 DVSS.n21559 4.5005
R28370 DVSS.n21623 DVSS.n21559 4.5005
R28371 DVSS.n21636 DVSS.n21559 4.5005
R28372 DVSS.n21622 DVSS.n21559 4.5005
R28373 DVSS.n21637 DVSS.n21559 4.5005
R28374 DVSS.n22073 DVSS.n21559 4.5005
R28375 DVSS.n21628 DVSS.n21601 4.5005
R28376 DVSS.n21630 DVSS.n21601 4.5005
R28377 DVSS.n21626 DVSS.n21601 4.5005
R28378 DVSS.n21632 DVSS.n21601 4.5005
R28379 DVSS.n21601 DVSS.n1463 4.5005
R28380 DVSS.n22075 DVSS.n21601 4.5005
R28381 DVSS.n21625 DVSS.n21601 4.5005
R28382 DVSS.n21633 DVSS.n21601 4.5005
R28383 DVSS.n21624 DVSS.n21601 4.5005
R28384 DVSS.n21634 DVSS.n21601 4.5005
R28385 DVSS.n21623 DVSS.n21601 4.5005
R28386 DVSS.n21636 DVSS.n21601 4.5005
R28387 DVSS.n21622 DVSS.n21601 4.5005
R28388 DVSS.n21637 DVSS.n21601 4.5005
R28389 DVSS.n22073 DVSS.n21601 4.5005
R28390 DVSS.n21628 DVSS.n21558 4.5005
R28391 DVSS.n21630 DVSS.n21558 4.5005
R28392 DVSS.n21626 DVSS.n21558 4.5005
R28393 DVSS.n21632 DVSS.n21558 4.5005
R28394 DVSS.n21558 DVSS.n1463 4.5005
R28395 DVSS.n22075 DVSS.n21558 4.5005
R28396 DVSS.n21625 DVSS.n21558 4.5005
R28397 DVSS.n21633 DVSS.n21558 4.5005
R28398 DVSS.n21624 DVSS.n21558 4.5005
R28399 DVSS.n21634 DVSS.n21558 4.5005
R28400 DVSS.n21623 DVSS.n21558 4.5005
R28401 DVSS.n21636 DVSS.n21558 4.5005
R28402 DVSS.n21637 DVSS.n21558 4.5005
R28403 DVSS.n22073 DVSS.n21558 4.5005
R28404 DVSS.n21628 DVSS.n21602 4.5005
R28405 DVSS.n21630 DVSS.n21602 4.5005
R28406 DVSS.n21626 DVSS.n21602 4.5005
R28407 DVSS.n21632 DVSS.n21602 4.5005
R28408 DVSS.n21602 DVSS.n1463 4.5005
R28409 DVSS.n22075 DVSS.n21602 4.5005
R28410 DVSS.n21625 DVSS.n21602 4.5005
R28411 DVSS.n21633 DVSS.n21602 4.5005
R28412 DVSS.n21624 DVSS.n21602 4.5005
R28413 DVSS.n21634 DVSS.n21602 4.5005
R28414 DVSS.n21623 DVSS.n21602 4.5005
R28415 DVSS.n21636 DVSS.n21602 4.5005
R28416 DVSS.n21637 DVSS.n21602 4.5005
R28417 DVSS.n22073 DVSS.n21602 4.5005
R28418 DVSS.n21628 DVSS.n21557 4.5005
R28419 DVSS.n21630 DVSS.n21557 4.5005
R28420 DVSS.n21626 DVSS.n21557 4.5005
R28421 DVSS.n21632 DVSS.n21557 4.5005
R28422 DVSS.n21557 DVSS.n1463 4.5005
R28423 DVSS.n22075 DVSS.n21557 4.5005
R28424 DVSS.n21625 DVSS.n21557 4.5005
R28425 DVSS.n21633 DVSS.n21557 4.5005
R28426 DVSS.n21624 DVSS.n21557 4.5005
R28427 DVSS.n21634 DVSS.n21557 4.5005
R28428 DVSS.n21623 DVSS.n21557 4.5005
R28429 DVSS.n21636 DVSS.n21557 4.5005
R28430 DVSS.n21622 DVSS.n21557 4.5005
R28431 DVSS.n21637 DVSS.n21557 4.5005
R28432 DVSS.n22073 DVSS.n21557 4.5005
R28433 DVSS.n22074 DVSS.n21628 4.5005
R28434 DVSS.n22074 DVSS.n21630 4.5005
R28435 DVSS.n22074 DVSS.n21626 4.5005
R28436 DVSS.n22074 DVSS.n21632 4.5005
R28437 DVSS.n22074 DVSS.n1463 4.5005
R28438 DVSS.n22075 DVSS.n22074 4.5005
R28439 DVSS.n22074 DVSS.n21625 4.5005
R28440 DVSS.n22074 DVSS.n21633 4.5005
R28441 DVSS.n22074 DVSS.n21624 4.5005
R28442 DVSS.n22074 DVSS.n21634 4.5005
R28443 DVSS.n22074 DVSS.n21623 4.5005
R28444 DVSS.n22074 DVSS.n21636 4.5005
R28445 DVSS.n22074 DVSS.n21622 4.5005
R28446 DVSS.n22074 DVSS.n21637 4.5005
R28447 DVSS.n22074 DVSS.n21615 4.5005
R28448 DVSS.n22074 DVSS.n22073 4.5005
R28449 DVSS.n21732 DVSS.n1178 4.5005
R28450 DVSS.n21734 DVSS.n1178 4.5005
R28451 DVSS.n21730 DVSS.n1178 4.5005
R28452 DVSS.n21738 DVSS.n1178 4.5005
R28453 DVSS.n21728 DVSS.n1178 4.5005
R28454 DVSS.n21739 DVSS.n1178 4.5005
R28455 DVSS.n21727 DVSS.n1178 4.5005
R28456 DVSS.n21682 DVSS.n1178 4.5005
R28457 DVSS.n22047 DVSS.n1178 4.5005
R28458 DVSS.n21742 DVSS.n1178 4.5005
R28459 DVSS.n22045 DVSS.n1178 4.5005
R28460 DVSS.n21732 DVSS.n21695 4.5005
R28461 DVSS.n21734 DVSS.n21695 4.5005
R28462 DVSS.n21730 DVSS.n21695 4.5005
R28463 DVSS.n21736 DVSS.n21695 4.5005
R28464 DVSS.n21729 DVSS.n21695 4.5005
R28465 DVSS.n21738 DVSS.n21695 4.5005
R28466 DVSS.n21728 DVSS.n21695 4.5005
R28467 DVSS.n21739 DVSS.n21695 4.5005
R28468 DVSS.n21727 DVSS.n21695 4.5005
R28469 DVSS.n21695 DVSS.n21682 4.5005
R28470 DVSS.n22047 DVSS.n21695 4.5005
R28471 DVSS.n21741 DVSS.n21695 4.5005
R28472 DVSS.n21742 DVSS.n21695 4.5005
R28473 DVSS.n22045 DVSS.n21695 4.5005
R28474 DVSS.n21732 DVSS.n21693 4.5005
R28475 DVSS.n21734 DVSS.n21693 4.5005
R28476 DVSS.n21730 DVSS.n21693 4.5005
R28477 DVSS.n21736 DVSS.n21693 4.5005
R28478 DVSS.n21729 DVSS.n21693 4.5005
R28479 DVSS.n21738 DVSS.n21693 4.5005
R28480 DVSS.n21728 DVSS.n21693 4.5005
R28481 DVSS.n21739 DVSS.n21693 4.5005
R28482 DVSS.n21727 DVSS.n21693 4.5005
R28483 DVSS.n21693 DVSS.n21682 4.5005
R28484 DVSS.n22047 DVSS.n21693 4.5005
R28485 DVSS.n21741 DVSS.n21693 4.5005
R28486 DVSS.n21742 DVSS.n21693 4.5005
R28487 DVSS.n21718 DVSS.n21693 4.5005
R28488 DVSS.n22045 DVSS.n21693 4.5005
R28489 DVSS.n21732 DVSS.n21696 4.5005
R28490 DVSS.n21734 DVSS.n21696 4.5005
R28491 DVSS.n21730 DVSS.n21696 4.5005
R28492 DVSS.n21736 DVSS.n21696 4.5005
R28493 DVSS.n21729 DVSS.n21696 4.5005
R28494 DVSS.n21738 DVSS.n21696 4.5005
R28495 DVSS.n21728 DVSS.n21696 4.5005
R28496 DVSS.n21739 DVSS.n21696 4.5005
R28497 DVSS.n21727 DVSS.n21696 4.5005
R28498 DVSS.n21696 DVSS.n21682 4.5005
R28499 DVSS.n22047 DVSS.n21696 4.5005
R28500 DVSS.n21741 DVSS.n21696 4.5005
R28501 DVSS.n21725 DVSS.n21696 4.5005
R28502 DVSS.n21742 DVSS.n21696 4.5005
R28503 DVSS.n22045 DVSS.n21696 4.5005
R28504 DVSS.n21732 DVSS.n21692 4.5005
R28505 DVSS.n21734 DVSS.n21692 4.5005
R28506 DVSS.n21730 DVSS.n21692 4.5005
R28507 DVSS.n21736 DVSS.n21692 4.5005
R28508 DVSS.n21729 DVSS.n21692 4.5005
R28509 DVSS.n21738 DVSS.n21692 4.5005
R28510 DVSS.n21728 DVSS.n21692 4.5005
R28511 DVSS.n21739 DVSS.n21692 4.5005
R28512 DVSS.n21727 DVSS.n21692 4.5005
R28513 DVSS.n21692 DVSS.n21682 4.5005
R28514 DVSS.n22047 DVSS.n21692 4.5005
R28515 DVSS.n21741 DVSS.n21692 4.5005
R28516 DVSS.n21742 DVSS.n21692 4.5005
R28517 DVSS.n22045 DVSS.n21692 4.5005
R28518 DVSS.n21732 DVSS.n21697 4.5005
R28519 DVSS.n21734 DVSS.n21697 4.5005
R28520 DVSS.n21730 DVSS.n21697 4.5005
R28521 DVSS.n21736 DVSS.n21697 4.5005
R28522 DVSS.n21729 DVSS.n21697 4.5005
R28523 DVSS.n21738 DVSS.n21697 4.5005
R28524 DVSS.n21728 DVSS.n21697 4.5005
R28525 DVSS.n21739 DVSS.n21697 4.5005
R28526 DVSS.n21727 DVSS.n21697 4.5005
R28527 DVSS.n21697 DVSS.n21682 4.5005
R28528 DVSS.n22047 DVSS.n21697 4.5005
R28529 DVSS.n21741 DVSS.n21697 4.5005
R28530 DVSS.n21742 DVSS.n21697 4.5005
R28531 DVSS.n22045 DVSS.n21697 4.5005
R28532 DVSS.n21732 DVSS.n21691 4.5005
R28533 DVSS.n21734 DVSS.n21691 4.5005
R28534 DVSS.n21730 DVSS.n21691 4.5005
R28535 DVSS.n21736 DVSS.n21691 4.5005
R28536 DVSS.n21729 DVSS.n21691 4.5005
R28537 DVSS.n21738 DVSS.n21691 4.5005
R28538 DVSS.n21728 DVSS.n21691 4.5005
R28539 DVSS.n21739 DVSS.n21691 4.5005
R28540 DVSS.n21727 DVSS.n21691 4.5005
R28541 DVSS.n21691 DVSS.n21682 4.5005
R28542 DVSS.n22047 DVSS.n21691 4.5005
R28543 DVSS.n21741 DVSS.n21691 4.5005
R28544 DVSS.n21725 DVSS.n21691 4.5005
R28545 DVSS.n21742 DVSS.n21691 4.5005
R28546 DVSS.n22045 DVSS.n21691 4.5005
R28547 DVSS.n21732 DVSS.n21698 4.5005
R28548 DVSS.n21734 DVSS.n21698 4.5005
R28549 DVSS.n21730 DVSS.n21698 4.5005
R28550 DVSS.n21736 DVSS.n21698 4.5005
R28551 DVSS.n21729 DVSS.n21698 4.5005
R28552 DVSS.n21738 DVSS.n21698 4.5005
R28553 DVSS.n21728 DVSS.n21698 4.5005
R28554 DVSS.n21739 DVSS.n21698 4.5005
R28555 DVSS.n21727 DVSS.n21698 4.5005
R28556 DVSS.n21698 DVSS.n21682 4.5005
R28557 DVSS.n22047 DVSS.n21698 4.5005
R28558 DVSS.n21741 DVSS.n21698 4.5005
R28559 DVSS.n21725 DVSS.n21698 4.5005
R28560 DVSS.n21742 DVSS.n21698 4.5005
R28561 DVSS.n22045 DVSS.n21698 4.5005
R28562 DVSS.n21732 DVSS.n21690 4.5005
R28563 DVSS.n21734 DVSS.n21690 4.5005
R28564 DVSS.n21730 DVSS.n21690 4.5005
R28565 DVSS.n21736 DVSS.n21690 4.5005
R28566 DVSS.n21729 DVSS.n21690 4.5005
R28567 DVSS.n21738 DVSS.n21690 4.5005
R28568 DVSS.n21728 DVSS.n21690 4.5005
R28569 DVSS.n21739 DVSS.n21690 4.5005
R28570 DVSS.n21727 DVSS.n21690 4.5005
R28571 DVSS.n21690 DVSS.n21682 4.5005
R28572 DVSS.n22047 DVSS.n21690 4.5005
R28573 DVSS.n21741 DVSS.n21690 4.5005
R28574 DVSS.n21742 DVSS.n21690 4.5005
R28575 DVSS.n22045 DVSS.n21690 4.5005
R28576 DVSS.n21732 DVSS.n21699 4.5005
R28577 DVSS.n21734 DVSS.n21699 4.5005
R28578 DVSS.n21730 DVSS.n21699 4.5005
R28579 DVSS.n21736 DVSS.n21699 4.5005
R28580 DVSS.n21729 DVSS.n21699 4.5005
R28581 DVSS.n21738 DVSS.n21699 4.5005
R28582 DVSS.n21728 DVSS.n21699 4.5005
R28583 DVSS.n21739 DVSS.n21699 4.5005
R28584 DVSS.n21727 DVSS.n21699 4.5005
R28585 DVSS.n21699 DVSS.n21682 4.5005
R28586 DVSS.n22047 DVSS.n21699 4.5005
R28587 DVSS.n21741 DVSS.n21699 4.5005
R28588 DVSS.n21742 DVSS.n21699 4.5005
R28589 DVSS.n22045 DVSS.n21699 4.5005
R28590 DVSS.n21732 DVSS.n21689 4.5005
R28591 DVSS.n21734 DVSS.n21689 4.5005
R28592 DVSS.n21730 DVSS.n21689 4.5005
R28593 DVSS.n21736 DVSS.n21689 4.5005
R28594 DVSS.n21729 DVSS.n21689 4.5005
R28595 DVSS.n21738 DVSS.n21689 4.5005
R28596 DVSS.n21728 DVSS.n21689 4.5005
R28597 DVSS.n21739 DVSS.n21689 4.5005
R28598 DVSS.n21727 DVSS.n21689 4.5005
R28599 DVSS.n21689 DVSS.n21682 4.5005
R28600 DVSS.n22047 DVSS.n21689 4.5005
R28601 DVSS.n21741 DVSS.n21689 4.5005
R28602 DVSS.n21725 DVSS.n21689 4.5005
R28603 DVSS.n21742 DVSS.n21689 4.5005
R28604 DVSS.n22045 DVSS.n21689 4.5005
R28605 DVSS.n21732 DVSS.n21700 4.5005
R28606 DVSS.n21734 DVSS.n21700 4.5005
R28607 DVSS.n21730 DVSS.n21700 4.5005
R28608 DVSS.n21736 DVSS.n21700 4.5005
R28609 DVSS.n21729 DVSS.n21700 4.5005
R28610 DVSS.n21738 DVSS.n21700 4.5005
R28611 DVSS.n21728 DVSS.n21700 4.5005
R28612 DVSS.n21739 DVSS.n21700 4.5005
R28613 DVSS.n21727 DVSS.n21700 4.5005
R28614 DVSS.n21700 DVSS.n21682 4.5005
R28615 DVSS.n22047 DVSS.n21700 4.5005
R28616 DVSS.n21741 DVSS.n21700 4.5005
R28617 DVSS.n21725 DVSS.n21700 4.5005
R28618 DVSS.n21742 DVSS.n21700 4.5005
R28619 DVSS.n22045 DVSS.n21700 4.5005
R28620 DVSS.n21732 DVSS.n21688 4.5005
R28621 DVSS.n21734 DVSS.n21688 4.5005
R28622 DVSS.n21730 DVSS.n21688 4.5005
R28623 DVSS.n21736 DVSS.n21688 4.5005
R28624 DVSS.n21729 DVSS.n21688 4.5005
R28625 DVSS.n21738 DVSS.n21688 4.5005
R28626 DVSS.n21728 DVSS.n21688 4.5005
R28627 DVSS.n21739 DVSS.n21688 4.5005
R28628 DVSS.n21727 DVSS.n21688 4.5005
R28629 DVSS.n21688 DVSS.n21682 4.5005
R28630 DVSS.n22047 DVSS.n21688 4.5005
R28631 DVSS.n21741 DVSS.n21688 4.5005
R28632 DVSS.n21742 DVSS.n21688 4.5005
R28633 DVSS.n22045 DVSS.n21688 4.5005
R28634 DVSS.n21732 DVSS.n21701 4.5005
R28635 DVSS.n21734 DVSS.n21701 4.5005
R28636 DVSS.n21730 DVSS.n21701 4.5005
R28637 DVSS.n21736 DVSS.n21701 4.5005
R28638 DVSS.n21729 DVSS.n21701 4.5005
R28639 DVSS.n21738 DVSS.n21701 4.5005
R28640 DVSS.n21728 DVSS.n21701 4.5005
R28641 DVSS.n21739 DVSS.n21701 4.5005
R28642 DVSS.n21727 DVSS.n21701 4.5005
R28643 DVSS.n21701 DVSS.n21682 4.5005
R28644 DVSS.n22047 DVSS.n21701 4.5005
R28645 DVSS.n21741 DVSS.n21701 4.5005
R28646 DVSS.n21742 DVSS.n21701 4.5005
R28647 DVSS.n22045 DVSS.n21701 4.5005
R28648 DVSS.n21732 DVSS.n21687 4.5005
R28649 DVSS.n21734 DVSS.n21687 4.5005
R28650 DVSS.n21730 DVSS.n21687 4.5005
R28651 DVSS.n21736 DVSS.n21687 4.5005
R28652 DVSS.n21729 DVSS.n21687 4.5005
R28653 DVSS.n21738 DVSS.n21687 4.5005
R28654 DVSS.n21728 DVSS.n21687 4.5005
R28655 DVSS.n21739 DVSS.n21687 4.5005
R28656 DVSS.n21727 DVSS.n21687 4.5005
R28657 DVSS.n21687 DVSS.n21682 4.5005
R28658 DVSS.n22047 DVSS.n21687 4.5005
R28659 DVSS.n21741 DVSS.n21687 4.5005
R28660 DVSS.n21725 DVSS.n21687 4.5005
R28661 DVSS.n21742 DVSS.n21687 4.5005
R28662 DVSS.n22045 DVSS.n21687 4.5005
R28663 DVSS.n21732 DVSS.n21702 4.5005
R28664 DVSS.n21734 DVSS.n21702 4.5005
R28665 DVSS.n21730 DVSS.n21702 4.5005
R28666 DVSS.n21736 DVSS.n21702 4.5005
R28667 DVSS.n21729 DVSS.n21702 4.5005
R28668 DVSS.n21738 DVSS.n21702 4.5005
R28669 DVSS.n21728 DVSS.n21702 4.5005
R28670 DVSS.n21739 DVSS.n21702 4.5005
R28671 DVSS.n21727 DVSS.n21702 4.5005
R28672 DVSS.n21702 DVSS.n21682 4.5005
R28673 DVSS.n22047 DVSS.n21702 4.5005
R28674 DVSS.n21741 DVSS.n21702 4.5005
R28675 DVSS.n21725 DVSS.n21702 4.5005
R28676 DVSS.n21742 DVSS.n21702 4.5005
R28677 DVSS.n22045 DVSS.n21702 4.5005
R28678 DVSS.n21732 DVSS.n21686 4.5005
R28679 DVSS.n21734 DVSS.n21686 4.5005
R28680 DVSS.n21730 DVSS.n21686 4.5005
R28681 DVSS.n21736 DVSS.n21686 4.5005
R28682 DVSS.n21729 DVSS.n21686 4.5005
R28683 DVSS.n21738 DVSS.n21686 4.5005
R28684 DVSS.n21728 DVSS.n21686 4.5005
R28685 DVSS.n21739 DVSS.n21686 4.5005
R28686 DVSS.n21727 DVSS.n21686 4.5005
R28687 DVSS.n21686 DVSS.n21682 4.5005
R28688 DVSS.n22047 DVSS.n21686 4.5005
R28689 DVSS.n21741 DVSS.n21686 4.5005
R28690 DVSS.n21742 DVSS.n21686 4.5005
R28691 DVSS.n22045 DVSS.n21686 4.5005
R28692 DVSS.n21732 DVSS.n21703 4.5005
R28693 DVSS.n21734 DVSS.n21703 4.5005
R28694 DVSS.n21730 DVSS.n21703 4.5005
R28695 DVSS.n21736 DVSS.n21703 4.5005
R28696 DVSS.n21729 DVSS.n21703 4.5005
R28697 DVSS.n21738 DVSS.n21703 4.5005
R28698 DVSS.n21728 DVSS.n21703 4.5005
R28699 DVSS.n21739 DVSS.n21703 4.5005
R28700 DVSS.n21727 DVSS.n21703 4.5005
R28701 DVSS.n21703 DVSS.n21682 4.5005
R28702 DVSS.n22047 DVSS.n21703 4.5005
R28703 DVSS.n21741 DVSS.n21703 4.5005
R28704 DVSS.n21742 DVSS.n21703 4.5005
R28705 DVSS.n22045 DVSS.n21703 4.5005
R28706 DVSS.n21732 DVSS.n21685 4.5005
R28707 DVSS.n21734 DVSS.n21685 4.5005
R28708 DVSS.n21730 DVSS.n21685 4.5005
R28709 DVSS.n21736 DVSS.n21685 4.5005
R28710 DVSS.n21729 DVSS.n21685 4.5005
R28711 DVSS.n21738 DVSS.n21685 4.5005
R28712 DVSS.n21728 DVSS.n21685 4.5005
R28713 DVSS.n21739 DVSS.n21685 4.5005
R28714 DVSS.n21727 DVSS.n21685 4.5005
R28715 DVSS.n21685 DVSS.n21682 4.5005
R28716 DVSS.n22047 DVSS.n21685 4.5005
R28717 DVSS.n21741 DVSS.n21685 4.5005
R28718 DVSS.n21725 DVSS.n21685 4.5005
R28719 DVSS.n21742 DVSS.n21685 4.5005
R28720 DVSS.n22045 DVSS.n21685 4.5005
R28721 DVSS.n21732 DVSS.n21704 4.5005
R28722 DVSS.n21734 DVSS.n21704 4.5005
R28723 DVSS.n21730 DVSS.n21704 4.5005
R28724 DVSS.n21736 DVSS.n21704 4.5005
R28725 DVSS.n21729 DVSS.n21704 4.5005
R28726 DVSS.n21738 DVSS.n21704 4.5005
R28727 DVSS.n21728 DVSS.n21704 4.5005
R28728 DVSS.n21739 DVSS.n21704 4.5005
R28729 DVSS.n21727 DVSS.n21704 4.5005
R28730 DVSS.n21704 DVSS.n21682 4.5005
R28731 DVSS.n22047 DVSS.n21704 4.5005
R28732 DVSS.n21741 DVSS.n21704 4.5005
R28733 DVSS.n21725 DVSS.n21704 4.5005
R28734 DVSS.n21742 DVSS.n21704 4.5005
R28735 DVSS.n22045 DVSS.n21704 4.5005
R28736 DVSS.n21732 DVSS.n21684 4.5005
R28737 DVSS.n21734 DVSS.n21684 4.5005
R28738 DVSS.n21730 DVSS.n21684 4.5005
R28739 DVSS.n21736 DVSS.n21684 4.5005
R28740 DVSS.n21729 DVSS.n21684 4.5005
R28741 DVSS.n21738 DVSS.n21684 4.5005
R28742 DVSS.n21728 DVSS.n21684 4.5005
R28743 DVSS.n21739 DVSS.n21684 4.5005
R28744 DVSS.n21727 DVSS.n21684 4.5005
R28745 DVSS.n21684 DVSS.n21682 4.5005
R28746 DVSS.n22047 DVSS.n21684 4.5005
R28747 DVSS.n21741 DVSS.n21684 4.5005
R28748 DVSS.n21742 DVSS.n21684 4.5005
R28749 DVSS.n22045 DVSS.n21684 4.5005
R28750 DVSS.n21732 DVSS.n21705 4.5005
R28751 DVSS.n21734 DVSS.n21705 4.5005
R28752 DVSS.n21730 DVSS.n21705 4.5005
R28753 DVSS.n21736 DVSS.n21705 4.5005
R28754 DVSS.n21729 DVSS.n21705 4.5005
R28755 DVSS.n21738 DVSS.n21705 4.5005
R28756 DVSS.n21728 DVSS.n21705 4.5005
R28757 DVSS.n21739 DVSS.n21705 4.5005
R28758 DVSS.n21727 DVSS.n21705 4.5005
R28759 DVSS.n21705 DVSS.n21682 4.5005
R28760 DVSS.n22047 DVSS.n21705 4.5005
R28761 DVSS.n21741 DVSS.n21705 4.5005
R28762 DVSS.n21742 DVSS.n21705 4.5005
R28763 DVSS.n22045 DVSS.n21705 4.5005
R28764 DVSS.n21732 DVSS.n21683 4.5005
R28765 DVSS.n21734 DVSS.n21683 4.5005
R28766 DVSS.n21730 DVSS.n21683 4.5005
R28767 DVSS.n21736 DVSS.n21683 4.5005
R28768 DVSS.n21729 DVSS.n21683 4.5005
R28769 DVSS.n21738 DVSS.n21683 4.5005
R28770 DVSS.n21728 DVSS.n21683 4.5005
R28771 DVSS.n21739 DVSS.n21683 4.5005
R28772 DVSS.n21727 DVSS.n21683 4.5005
R28773 DVSS.n21683 DVSS.n21682 4.5005
R28774 DVSS.n22047 DVSS.n21683 4.5005
R28775 DVSS.n21741 DVSS.n21683 4.5005
R28776 DVSS.n21725 DVSS.n21683 4.5005
R28777 DVSS.n21742 DVSS.n21683 4.5005
R28778 DVSS.n22045 DVSS.n21683 4.5005
R28779 DVSS.n22046 DVSS.n21732 4.5005
R28780 DVSS.n22046 DVSS.n21734 4.5005
R28781 DVSS.n22046 DVSS.n21730 4.5005
R28782 DVSS.n22046 DVSS.n21736 4.5005
R28783 DVSS.n22046 DVSS.n21729 4.5005
R28784 DVSS.n22046 DVSS.n21738 4.5005
R28785 DVSS.n22046 DVSS.n21728 4.5005
R28786 DVSS.n22046 DVSS.n21739 4.5005
R28787 DVSS.n22046 DVSS.n21727 4.5005
R28788 DVSS.n22046 DVSS.n21682 4.5005
R28789 DVSS.n22047 DVSS.n22046 4.5005
R28790 DVSS.n22046 DVSS.n21741 4.5005
R28791 DVSS.n22046 DVSS.n21725 4.5005
R28792 DVSS.n22046 DVSS.n21742 4.5005
R28793 DVSS.n22046 DVSS.n21718 4.5005
R28794 DVSS.n22046 DVSS.n22045 4.5005
R28795 DVSS.n21824 DVSS.n1199 4.5005
R28796 DVSS.n21954 DVSS.n1199 4.5005
R28797 DVSS.n21822 DVSS.n1199 4.5005
R28798 DVSS.n21955 DVSS.n1199 4.5005
R28799 DVSS.n21821 DVSS.n1199 4.5005
R28800 DVSS.n21957 DVSS.n1199 4.5005
R28801 DVSS.n21820 DVSS.n1199 4.5005
R28802 DVSS.n21961 DVSS.n1199 4.5005
R28803 DVSS.n21818 DVSS.n1199 4.5005
R28804 DVSS.n21962 DVSS.n1199 4.5005
R28805 DVSS.n21964 DVSS.n1199 4.5005
R28806 DVSS.n21824 DVSS.n21788 4.5005
R28807 DVSS.n21952 DVSS.n21788 4.5005
R28808 DVSS.n21823 DVSS.n21788 4.5005
R28809 DVSS.n21954 DVSS.n21788 4.5005
R28810 DVSS.n21822 DVSS.n21788 4.5005
R28811 DVSS.n21955 DVSS.n21788 4.5005
R28812 DVSS.n21821 DVSS.n21788 4.5005
R28813 DVSS.n21957 DVSS.n21788 4.5005
R28814 DVSS.n21820 DVSS.n21788 4.5005
R28815 DVSS.n21959 DVSS.n21788 4.5005
R28816 DVSS.n21819 DVSS.n21788 4.5005
R28817 DVSS.n21961 DVSS.n21788 4.5005
R28818 DVSS.n21962 DVSS.n21788 4.5005
R28819 DVSS.n21964 DVSS.n21788 4.5005
R28820 DVSS.n21824 DVSS.n21787 4.5005
R28821 DVSS.n21952 DVSS.n21787 4.5005
R28822 DVSS.n21823 DVSS.n21787 4.5005
R28823 DVSS.n21954 DVSS.n21787 4.5005
R28824 DVSS.n21822 DVSS.n21787 4.5005
R28825 DVSS.n21955 DVSS.n21787 4.5005
R28826 DVSS.n21821 DVSS.n21787 4.5005
R28827 DVSS.n21957 DVSS.n21787 4.5005
R28828 DVSS.n21820 DVSS.n21787 4.5005
R28829 DVSS.n21959 DVSS.n21787 4.5005
R28830 DVSS.n21819 DVSS.n21787 4.5005
R28831 DVSS.n21961 DVSS.n21787 4.5005
R28832 DVSS.n21962 DVSS.n21787 4.5005
R28833 DVSS.n21811 DVSS.n21787 4.5005
R28834 DVSS.n21964 DVSS.n21787 4.5005
R28835 DVSS.n21824 DVSS.n21789 4.5005
R28836 DVSS.n21952 DVSS.n21789 4.5005
R28837 DVSS.n21823 DVSS.n21789 4.5005
R28838 DVSS.n21954 DVSS.n21789 4.5005
R28839 DVSS.n21822 DVSS.n21789 4.5005
R28840 DVSS.n21955 DVSS.n21789 4.5005
R28841 DVSS.n21821 DVSS.n21789 4.5005
R28842 DVSS.n21957 DVSS.n21789 4.5005
R28843 DVSS.n21820 DVSS.n21789 4.5005
R28844 DVSS.n21959 DVSS.n21789 4.5005
R28845 DVSS.n21819 DVSS.n21789 4.5005
R28846 DVSS.n21961 DVSS.n21789 4.5005
R28847 DVSS.n21818 DVSS.n21789 4.5005
R28848 DVSS.n21962 DVSS.n21789 4.5005
R28849 DVSS.n21964 DVSS.n21789 4.5005
R28850 DVSS.n21824 DVSS.n21786 4.5005
R28851 DVSS.n21952 DVSS.n21786 4.5005
R28852 DVSS.n21823 DVSS.n21786 4.5005
R28853 DVSS.n21954 DVSS.n21786 4.5005
R28854 DVSS.n21822 DVSS.n21786 4.5005
R28855 DVSS.n21955 DVSS.n21786 4.5005
R28856 DVSS.n21821 DVSS.n21786 4.5005
R28857 DVSS.n21957 DVSS.n21786 4.5005
R28858 DVSS.n21820 DVSS.n21786 4.5005
R28859 DVSS.n21959 DVSS.n21786 4.5005
R28860 DVSS.n21819 DVSS.n21786 4.5005
R28861 DVSS.n21961 DVSS.n21786 4.5005
R28862 DVSS.n21962 DVSS.n21786 4.5005
R28863 DVSS.n21964 DVSS.n21786 4.5005
R28864 DVSS.n21824 DVSS.n21790 4.5005
R28865 DVSS.n21952 DVSS.n21790 4.5005
R28866 DVSS.n21823 DVSS.n21790 4.5005
R28867 DVSS.n21954 DVSS.n21790 4.5005
R28868 DVSS.n21822 DVSS.n21790 4.5005
R28869 DVSS.n21955 DVSS.n21790 4.5005
R28870 DVSS.n21821 DVSS.n21790 4.5005
R28871 DVSS.n21957 DVSS.n21790 4.5005
R28872 DVSS.n21820 DVSS.n21790 4.5005
R28873 DVSS.n21959 DVSS.n21790 4.5005
R28874 DVSS.n21819 DVSS.n21790 4.5005
R28875 DVSS.n21961 DVSS.n21790 4.5005
R28876 DVSS.n21962 DVSS.n21790 4.5005
R28877 DVSS.n21964 DVSS.n21790 4.5005
R28878 DVSS.n21824 DVSS.n21785 4.5005
R28879 DVSS.n21952 DVSS.n21785 4.5005
R28880 DVSS.n21823 DVSS.n21785 4.5005
R28881 DVSS.n21954 DVSS.n21785 4.5005
R28882 DVSS.n21822 DVSS.n21785 4.5005
R28883 DVSS.n21955 DVSS.n21785 4.5005
R28884 DVSS.n21821 DVSS.n21785 4.5005
R28885 DVSS.n21957 DVSS.n21785 4.5005
R28886 DVSS.n21820 DVSS.n21785 4.5005
R28887 DVSS.n21959 DVSS.n21785 4.5005
R28888 DVSS.n21819 DVSS.n21785 4.5005
R28889 DVSS.n21961 DVSS.n21785 4.5005
R28890 DVSS.n21818 DVSS.n21785 4.5005
R28891 DVSS.n21962 DVSS.n21785 4.5005
R28892 DVSS.n21964 DVSS.n21785 4.5005
R28893 DVSS.n21824 DVSS.n21791 4.5005
R28894 DVSS.n21952 DVSS.n21791 4.5005
R28895 DVSS.n21823 DVSS.n21791 4.5005
R28896 DVSS.n21954 DVSS.n21791 4.5005
R28897 DVSS.n21822 DVSS.n21791 4.5005
R28898 DVSS.n21955 DVSS.n21791 4.5005
R28899 DVSS.n21821 DVSS.n21791 4.5005
R28900 DVSS.n21957 DVSS.n21791 4.5005
R28901 DVSS.n21820 DVSS.n21791 4.5005
R28902 DVSS.n21959 DVSS.n21791 4.5005
R28903 DVSS.n21819 DVSS.n21791 4.5005
R28904 DVSS.n21961 DVSS.n21791 4.5005
R28905 DVSS.n21818 DVSS.n21791 4.5005
R28906 DVSS.n21962 DVSS.n21791 4.5005
R28907 DVSS.n21964 DVSS.n21791 4.5005
R28908 DVSS.n21824 DVSS.n21784 4.5005
R28909 DVSS.n21952 DVSS.n21784 4.5005
R28910 DVSS.n21823 DVSS.n21784 4.5005
R28911 DVSS.n21954 DVSS.n21784 4.5005
R28912 DVSS.n21822 DVSS.n21784 4.5005
R28913 DVSS.n21955 DVSS.n21784 4.5005
R28914 DVSS.n21821 DVSS.n21784 4.5005
R28915 DVSS.n21957 DVSS.n21784 4.5005
R28916 DVSS.n21820 DVSS.n21784 4.5005
R28917 DVSS.n21959 DVSS.n21784 4.5005
R28918 DVSS.n21819 DVSS.n21784 4.5005
R28919 DVSS.n21961 DVSS.n21784 4.5005
R28920 DVSS.n21962 DVSS.n21784 4.5005
R28921 DVSS.n21964 DVSS.n21784 4.5005
R28922 DVSS.n21824 DVSS.n21792 4.5005
R28923 DVSS.n21952 DVSS.n21792 4.5005
R28924 DVSS.n21823 DVSS.n21792 4.5005
R28925 DVSS.n21954 DVSS.n21792 4.5005
R28926 DVSS.n21822 DVSS.n21792 4.5005
R28927 DVSS.n21955 DVSS.n21792 4.5005
R28928 DVSS.n21821 DVSS.n21792 4.5005
R28929 DVSS.n21957 DVSS.n21792 4.5005
R28930 DVSS.n21820 DVSS.n21792 4.5005
R28931 DVSS.n21959 DVSS.n21792 4.5005
R28932 DVSS.n21819 DVSS.n21792 4.5005
R28933 DVSS.n21961 DVSS.n21792 4.5005
R28934 DVSS.n21962 DVSS.n21792 4.5005
R28935 DVSS.n21964 DVSS.n21792 4.5005
R28936 DVSS.n21824 DVSS.n21783 4.5005
R28937 DVSS.n21952 DVSS.n21783 4.5005
R28938 DVSS.n21823 DVSS.n21783 4.5005
R28939 DVSS.n21954 DVSS.n21783 4.5005
R28940 DVSS.n21822 DVSS.n21783 4.5005
R28941 DVSS.n21955 DVSS.n21783 4.5005
R28942 DVSS.n21821 DVSS.n21783 4.5005
R28943 DVSS.n21957 DVSS.n21783 4.5005
R28944 DVSS.n21820 DVSS.n21783 4.5005
R28945 DVSS.n21959 DVSS.n21783 4.5005
R28946 DVSS.n21819 DVSS.n21783 4.5005
R28947 DVSS.n21961 DVSS.n21783 4.5005
R28948 DVSS.n21818 DVSS.n21783 4.5005
R28949 DVSS.n21962 DVSS.n21783 4.5005
R28950 DVSS.n21964 DVSS.n21783 4.5005
R28951 DVSS.n21824 DVSS.n21793 4.5005
R28952 DVSS.n21952 DVSS.n21793 4.5005
R28953 DVSS.n21823 DVSS.n21793 4.5005
R28954 DVSS.n21954 DVSS.n21793 4.5005
R28955 DVSS.n21822 DVSS.n21793 4.5005
R28956 DVSS.n21955 DVSS.n21793 4.5005
R28957 DVSS.n21821 DVSS.n21793 4.5005
R28958 DVSS.n21957 DVSS.n21793 4.5005
R28959 DVSS.n21820 DVSS.n21793 4.5005
R28960 DVSS.n21959 DVSS.n21793 4.5005
R28961 DVSS.n21819 DVSS.n21793 4.5005
R28962 DVSS.n21961 DVSS.n21793 4.5005
R28963 DVSS.n21818 DVSS.n21793 4.5005
R28964 DVSS.n21962 DVSS.n21793 4.5005
R28965 DVSS.n21964 DVSS.n21793 4.5005
R28966 DVSS.n21824 DVSS.n21782 4.5005
R28967 DVSS.n21952 DVSS.n21782 4.5005
R28968 DVSS.n21823 DVSS.n21782 4.5005
R28969 DVSS.n21954 DVSS.n21782 4.5005
R28970 DVSS.n21822 DVSS.n21782 4.5005
R28971 DVSS.n21955 DVSS.n21782 4.5005
R28972 DVSS.n21821 DVSS.n21782 4.5005
R28973 DVSS.n21957 DVSS.n21782 4.5005
R28974 DVSS.n21820 DVSS.n21782 4.5005
R28975 DVSS.n21959 DVSS.n21782 4.5005
R28976 DVSS.n21819 DVSS.n21782 4.5005
R28977 DVSS.n21961 DVSS.n21782 4.5005
R28978 DVSS.n21962 DVSS.n21782 4.5005
R28979 DVSS.n21964 DVSS.n21782 4.5005
R28980 DVSS.n21824 DVSS.n21794 4.5005
R28981 DVSS.n21952 DVSS.n21794 4.5005
R28982 DVSS.n21823 DVSS.n21794 4.5005
R28983 DVSS.n21954 DVSS.n21794 4.5005
R28984 DVSS.n21822 DVSS.n21794 4.5005
R28985 DVSS.n21955 DVSS.n21794 4.5005
R28986 DVSS.n21821 DVSS.n21794 4.5005
R28987 DVSS.n21957 DVSS.n21794 4.5005
R28988 DVSS.n21820 DVSS.n21794 4.5005
R28989 DVSS.n21959 DVSS.n21794 4.5005
R28990 DVSS.n21819 DVSS.n21794 4.5005
R28991 DVSS.n21961 DVSS.n21794 4.5005
R28992 DVSS.n21962 DVSS.n21794 4.5005
R28993 DVSS.n21964 DVSS.n21794 4.5005
R28994 DVSS.n21824 DVSS.n21781 4.5005
R28995 DVSS.n21952 DVSS.n21781 4.5005
R28996 DVSS.n21823 DVSS.n21781 4.5005
R28997 DVSS.n21954 DVSS.n21781 4.5005
R28998 DVSS.n21822 DVSS.n21781 4.5005
R28999 DVSS.n21955 DVSS.n21781 4.5005
R29000 DVSS.n21821 DVSS.n21781 4.5005
R29001 DVSS.n21957 DVSS.n21781 4.5005
R29002 DVSS.n21820 DVSS.n21781 4.5005
R29003 DVSS.n21959 DVSS.n21781 4.5005
R29004 DVSS.n21819 DVSS.n21781 4.5005
R29005 DVSS.n21961 DVSS.n21781 4.5005
R29006 DVSS.n21818 DVSS.n21781 4.5005
R29007 DVSS.n21962 DVSS.n21781 4.5005
R29008 DVSS.n21964 DVSS.n21781 4.5005
R29009 DVSS.n21824 DVSS.n21795 4.5005
R29010 DVSS.n21952 DVSS.n21795 4.5005
R29011 DVSS.n21823 DVSS.n21795 4.5005
R29012 DVSS.n21954 DVSS.n21795 4.5005
R29013 DVSS.n21822 DVSS.n21795 4.5005
R29014 DVSS.n21955 DVSS.n21795 4.5005
R29015 DVSS.n21821 DVSS.n21795 4.5005
R29016 DVSS.n21957 DVSS.n21795 4.5005
R29017 DVSS.n21820 DVSS.n21795 4.5005
R29018 DVSS.n21959 DVSS.n21795 4.5005
R29019 DVSS.n21819 DVSS.n21795 4.5005
R29020 DVSS.n21961 DVSS.n21795 4.5005
R29021 DVSS.n21818 DVSS.n21795 4.5005
R29022 DVSS.n21962 DVSS.n21795 4.5005
R29023 DVSS.n21964 DVSS.n21795 4.5005
R29024 DVSS.n21824 DVSS.n21780 4.5005
R29025 DVSS.n21952 DVSS.n21780 4.5005
R29026 DVSS.n21823 DVSS.n21780 4.5005
R29027 DVSS.n21954 DVSS.n21780 4.5005
R29028 DVSS.n21822 DVSS.n21780 4.5005
R29029 DVSS.n21955 DVSS.n21780 4.5005
R29030 DVSS.n21821 DVSS.n21780 4.5005
R29031 DVSS.n21957 DVSS.n21780 4.5005
R29032 DVSS.n21820 DVSS.n21780 4.5005
R29033 DVSS.n21959 DVSS.n21780 4.5005
R29034 DVSS.n21819 DVSS.n21780 4.5005
R29035 DVSS.n21961 DVSS.n21780 4.5005
R29036 DVSS.n21962 DVSS.n21780 4.5005
R29037 DVSS.n21964 DVSS.n21780 4.5005
R29038 DVSS.n21824 DVSS.n21796 4.5005
R29039 DVSS.n21952 DVSS.n21796 4.5005
R29040 DVSS.n21823 DVSS.n21796 4.5005
R29041 DVSS.n21954 DVSS.n21796 4.5005
R29042 DVSS.n21822 DVSS.n21796 4.5005
R29043 DVSS.n21955 DVSS.n21796 4.5005
R29044 DVSS.n21821 DVSS.n21796 4.5005
R29045 DVSS.n21957 DVSS.n21796 4.5005
R29046 DVSS.n21820 DVSS.n21796 4.5005
R29047 DVSS.n21959 DVSS.n21796 4.5005
R29048 DVSS.n21819 DVSS.n21796 4.5005
R29049 DVSS.n21961 DVSS.n21796 4.5005
R29050 DVSS.n21962 DVSS.n21796 4.5005
R29051 DVSS.n21964 DVSS.n21796 4.5005
R29052 DVSS.n21824 DVSS.n21779 4.5005
R29053 DVSS.n21952 DVSS.n21779 4.5005
R29054 DVSS.n21823 DVSS.n21779 4.5005
R29055 DVSS.n21954 DVSS.n21779 4.5005
R29056 DVSS.n21822 DVSS.n21779 4.5005
R29057 DVSS.n21955 DVSS.n21779 4.5005
R29058 DVSS.n21821 DVSS.n21779 4.5005
R29059 DVSS.n21957 DVSS.n21779 4.5005
R29060 DVSS.n21820 DVSS.n21779 4.5005
R29061 DVSS.n21959 DVSS.n21779 4.5005
R29062 DVSS.n21819 DVSS.n21779 4.5005
R29063 DVSS.n21961 DVSS.n21779 4.5005
R29064 DVSS.n21818 DVSS.n21779 4.5005
R29065 DVSS.n21962 DVSS.n21779 4.5005
R29066 DVSS.n21964 DVSS.n21779 4.5005
R29067 DVSS.n21824 DVSS.n21797 4.5005
R29068 DVSS.n21952 DVSS.n21797 4.5005
R29069 DVSS.n21823 DVSS.n21797 4.5005
R29070 DVSS.n21954 DVSS.n21797 4.5005
R29071 DVSS.n21822 DVSS.n21797 4.5005
R29072 DVSS.n21955 DVSS.n21797 4.5005
R29073 DVSS.n21821 DVSS.n21797 4.5005
R29074 DVSS.n21957 DVSS.n21797 4.5005
R29075 DVSS.n21820 DVSS.n21797 4.5005
R29076 DVSS.n21959 DVSS.n21797 4.5005
R29077 DVSS.n21819 DVSS.n21797 4.5005
R29078 DVSS.n21961 DVSS.n21797 4.5005
R29079 DVSS.n21818 DVSS.n21797 4.5005
R29080 DVSS.n21962 DVSS.n21797 4.5005
R29081 DVSS.n21964 DVSS.n21797 4.5005
R29082 DVSS.n21824 DVSS.n21778 4.5005
R29083 DVSS.n21952 DVSS.n21778 4.5005
R29084 DVSS.n21823 DVSS.n21778 4.5005
R29085 DVSS.n21954 DVSS.n21778 4.5005
R29086 DVSS.n21822 DVSS.n21778 4.5005
R29087 DVSS.n21955 DVSS.n21778 4.5005
R29088 DVSS.n21821 DVSS.n21778 4.5005
R29089 DVSS.n21957 DVSS.n21778 4.5005
R29090 DVSS.n21820 DVSS.n21778 4.5005
R29091 DVSS.n21959 DVSS.n21778 4.5005
R29092 DVSS.n21819 DVSS.n21778 4.5005
R29093 DVSS.n21961 DVSS.n21778 4.5005
R29094 DVSS.n21962 DVSS.n21778 4.5005
R29095 DVSS.n21964 DVSS.n21778 4.5005
R29096 DVSS.n21824 DVSS.n21798 4.5005
R29097 DVSS.n21952 DVSS.n21798 4.5005
R29098 DVSS.n21823 DVSS.n21798 4.5005
R29099 DVSS.n21954 DVSS.n21798 4.5005
R29100 DVSS.n21822 DVSS.n21798 4.5005
R29101 DVSS.n21955 DVSS.n21798 4.5005
R29102 DVSS.n21821 DVSS.n21798 4.5005
R29103 DVSS.n21957 DVSS.n21798 4.5005
R29104 DVSS.n21820 DVSS.n21798 4.5005
R29105 DVSS.n21959 DVSS.n21798 4.5005
R29106 DVSS.n21819 DVSS.n21798 4.5005
R29107 DVSS.n21961 DVSS.n21798 4.5005
R29108 DVSS.n21962 DVSS.n21798 4.5005
R29109 DVSS.n21964 DVSS.n21798 4.5005
R29110 DVSS.n21824 DVSS.n21777 4.5005
R29111 DVSS.n21952 DVSS.n21777 4.5005
R29112 DVSS.n21823 DVSS.n21777 4.5005
R29113 DVSS.n21954 DVSS.n21777 4.5005
R29114 DVSS.n21822 DVSS.n21777 4.5005
R29115 DVSS.n21955 DVSS.n21777 4.5005
R29116 DVSS.n21821 DVSS.n21777 4.5005
R29117 DVSS.n21957 DVSS.n21777 4.5005
R29118 DVSS.n21820 DVSS.n21777 4.5005
R29119 DVSS.n21959 DVSS.n21777 4.5005
R29120 DVSS.n21819 DVSS.n21777 4.5005
R29121 DVSS.n21961 DVSS.n21777 4.5005
R29122 DVSS.n21818 DVSS.n21777 4.5005
R29123 DVSS.n21962 DVSS.n21777 4.5005
R29124 DVSS.n21964 DVSS.n21777 4.5005
R29125 DVSS.n21963 DVSS.n21824 4.5005
R29126 DVSS.n21963 DVSS.n21952 4.5005
R29127 DVSS.n21963 DVSS.n21823 4.5005
R29128 DVSS.n21963 DVSS.n21954 4.5005
R29129 DVSS.n21963 DVSS.n21822 4.5005
R29130 DVSS.n21963 DVSS.n21955 4.5005
R29131 DVSS.n21963 DVSS.n21821 4.5005
R29132 DVSS.n21963 DVSS.n21957 4.5005
R29133 DVSS.n21963 DVSS.n21820 4.5005
R29134 DVSS.n21963 DVSS.n21959 4.5005
R29135 DVSS.n21963 DVSS.n21819 4.5005
R29136 DVSS.n21963 DVSS.n21961 4.5005
R29137 DVSS.n21963 DVSS.n21818 4.5005
R29138 DVSS.n21963 DVSS.n21962 4.5005
R29139 DVSS.n21963 DVSS.n21811 4.5005
R29140 DVSS.n21964 DVSS.n21963 4.5005
R29141 DVSS.n18993 DVSS.n18645 3.91226
R29142 DVSS.n18989 DVSS.n18645 3.91226
R29143 DVSS.n18989 DVSS.n18649 3.91226
R29144 DVSS.n18900 DVSS.n18649 3.91226
R29145 DVSS.n18902 DVSS.n18900 3.91226
R29146 DVSS.n18904 DVSS.n18902 3.91226
R29147 DVSS.n18904 DVSS.n14545 3.91226
R29148 DVSS.n20692 DVSS.n14545 3.91226
R29149 DVSS.n20692 DVSS.n14546 3.91226
R29150 DVSS.n18944 DVSS.n14546 3.91226
R29151 DVSS.n18960 DVSS.n18944 3.91226
R29152 DVSS.n18962 DVSS.n18960 3.91226
R29153 DVSS.n18964 DVSS.n18962 3.91226
R29154 DVSS.n18964 DVSS.n18928 3.91226
R29155 DVSS.n18972 DVSS.n18928 3.91226
R29156 DVSS.n18974 DVSS.n18972 3.91226
R29157 DVSS.n18979 DVSS.n18974 3.91226
R29158 DVSS.n18979 DVSS.n18977 3.91226
R29159 DVSS.n18977 DVSS.n14569 3.91226
R29160 DVSS.n20685 DVSS.n14569 3.91226
R29161 DVSS.n20685 DVSS.n14570 3.91226
R29162 DVSS.n20677 DVSS.n14570 3.91226
R29163 DVSS.n20677 DVSS.n14583 3.91226
R29164 DVSS.n20100 DVSS.n14583 3.91226
R29165 DVSS.n20122 DVSS.n20100 3.91226
R29166 DVSS.n20124 DVSS.n20122 3.91226
R29167 DVSS.n20126 DVSS.n20124 3.91226
R29168 DVSS.n20126 DVSS.n20085 3.91226
R29169 DVSS.n20134 DVSS.n20085 3.91226
R29170 DVSS.n20136 DVSS.n20134 3.91226
R29171 DVSS.n20138 DVSS.n20136 3.91226
R29172 DVSS.n20138 DVSS.n20070 3.91226
R29173 DVSS.n20146 DVSS.n20070 3.91226
R29174 DVSS.n20148 DVSS.n20146 3.91226
R29175 DVSS.n20150 DVSS.n20148 3.91226
R29176 DVSS.n20150 DVSS.n20033 3.91226
R29177 DVSS.n20163 DVSS.n20033 3.91226
R29178 DVSS.n20165 DVSS.n20163 3.91226
R29179 DVSS.n20168 DVSS.n20165 3.91226
R29180 DVSS.n20168 DVSS.n14604 3.91226
R29181 DVSS.n20670 DVSS.n14604 3.91226
R29182 DVSS.n20670 DVSS.n14605 3.91226
R29183 DVSS.n20662 DVSS.n14605 3.91226
R29184 DVSS.n20662 DVSS.n14615 3.91226
R29185 DVSS.n20658 DVSS.n14615 3.91226
R29186 DVSS.n20658 DVSS.n14617 3.91226
R29187 DVSS.n20650 DVSS.n14617 3.91226
R29188 DVSS.n20650 DVSS.n14629 3.91226
R29189 DVSS.n20269 DVSS.n14629 3.91226
R29190 DVSS.n20269 DVSS.n20254 3.91226
R29191 DVSS.n20277 DVSS.n20254 3.91226
R29192 DVSS.n20279 DVSS.n20277 3.91226
R29193 DVSS.n20281 DVSS.n20279 3.91226
R29194 DVSS.n20281 DVSS.n20238 3.91226
R29195 DVSS.n20289 DVSS.n20238 3.91226
R29196 DVSS.n20291 DVSS.n20289 3.91226
R29197 DVSS.n20295 DVSS.n20291 3.91226
R29198 DVSS.n20295 DVSS.n20293 3.91226
R29199 DVSS.n20293 DVSS.n20201 3.91226
R29200 DVSS.n20309 DVSS.n20201 3.91226
R29201 DVSS.n20311 DVSS.n20309 3.91226
R29202 DVSS.n20312 DVSS.n20311 3.91226
R29203 DVSS.n20312 DVSS.n14653 3.91226
R29204 DVSS.n20644 DVSS.n14653 3.91226
R29205 DVSS.n20644 DVSS.n14654 3.91226
R29206 DVSS.n20635 DVSS.n14654 3.91226
R29207 DVSS.n20635 DVSS.n14667 3.91226
R29208 DVSS.n20630 DVSS.n14667 3.91226
R29209 DVSS.n20630 DVSS.n14670 3.91226
R29210 DVSS.n20395 DVSS.n14670 3.91226
R29211 DVSS.n20403 DVSS.n20395 3.91226
R29212 DVSS.n20403 DVSS.n20377 3.91226
R29213 DVSS.n20411 DVSS.n20377 3.91226
R29214 DVSS.n20411 DVSS.n20375 3.91226
R29215 DVSS.n20419 DVSS.n20375 3.91226
R29216 DVSS.n20419 DVSS.n20360 3.91226
R29217 DVSS.n20427 DVSS.n20360 3.91226
R29218 DVSS.n20427 DVSS.n20355 3.91226
R29219 DVSS.n20434 DVSS.n20355 3.91226
R29220 DVSS.n20434 DVSS.n20342 3.91226
R29221 DVSS.n20444 DVSS.n20342 3.91226
R29222 DVSS.n20444 DVSS.n20340 3.91226
R29223 DVSS.n20453 DVSS.n20340 3.91226
R29224 DVSS.n20453 DVSS.n14700 3.91226
R29225 DVSS.n20621 DVSS.n14700 3.91226
R29226 DVSS.n20621 DVSS.n14701 3.91226
R29227 DVSS.n20617 DVSS.n14701 3.91226
R29228 DVSS.n18652 DVSS.n18644 3.91226
R29229 DVSS.n18987 DVSS.n18652 3.91226
R29230 DVSS.n18987 DVSS.n18653 3.91226
R29231 DVSS.n18898 DVSS.n18653 3.91226
R29232 DVSS.n18898 DVSS.n18885 3.91226
R29233 DVSS.n18906 DVSS.n18885 3.91226
R29234 DVSS.n18906 DVSS.n18886 3.91226
R29235 DVSS.n18886 DVSS.n14544 3.91226
R29236 DVSS.n18954 DVSS.n14544 3.91226
R29237 DVSS.n18956 DVSS.n18954 3.91226
R29238 DVSS.n18958 DVSS.n18956 3.91226
R29239 DVSS.n18958 DVSS.n18936 3.91226
R29240 DVSS.n18966 DVSS.n18936 3.91226
R29241 DVSS.n18968 DVSS.n18966 3.91226
R29242 DVSS.n18970 DVSS.n18968 3.91226
R29243 DVSS.n18970 DVSS.n18916 3.91226
R29244 DVSS.n18981 DVSS.n18916 3.91226
R29245 DVSS.n18981 DVSS.n18918 3.91226
R29246 DVSS.n18918 DVSS.n14574 3.91226
R29247 DVSS.n20683 DVSS.n14574 3.91226
R29248 DVSS.n20683 DVSS.n14575 3.91226
R29249 DVSS.n20679 DVSS.n14575 3.91226
R29250 DVSS.n20679 DVSS.n14580 3.91226
R29251 DVSS.n20118 DVSS.n14580 3.91226
R29252 DVSS.n20120 DVSS.n20118 3.91226
R29253 DVSS.n20120 DVSS.n20093 3.91226
R29254 DVSS.n20128 DVSS.n20093 3.91226
R29255 DVSS.n20130 DVSS.n20128 3.91226
R29256 DVSS.n20132 DVSS.n20130 3.91226
R29257 DVSS.n20132 DVSS.n20077 3.91226
R29258 DVSS.n20140 DVSS.n20077 3.91226
R29259 DVSS.n20142 DVSS.n20140 3.91226
R29260 DVSS.n20144 DVSS.n20142 3.91226
R29261 DVSS.n20144 DVSS.n20063 3.91226
R29262 DVSS.n20152 DVSS.n20063 3.91226
R29263 DVSS.n20152 DVSS.n20038 3.91226
R29264 DVSS.n20161 DVSS.n20038 3.91226
R29265 DVSS.n20161 DVSS.n20039 3.91226
R29266 DVSS.n20039 DVSS.n20031 3.91226
R29267 DVSS.n20031 DVSS.n14609 3.91226
R29268 DVSS.n20668 DVSS.n14609 3.91226
R29269 DVSS.n20668 DVSS.n14610 3.91226
R29270 DVSS.n20664 DVSS.n14610 3.91226
R29271 DVSS.n20664 DVSS.n14612 3.91226
R29272 DVSS.n20656 DVSS.n14612 3.91226
R29273 DVSS.n20656 DVSS.n14620 3.91226
R29274 DVSS.n20652 DVSS.n14620 3.91226
R29275 DVSS.n20652 DVSS.n14626 3.91226
R29276 DVSS.n20271 DVSS.n14626 3.91226
R29277 DVSS.n20273 DVSS.n20271 3.91226
R29278 DVSS.n20275 DVSS.n20273 3.91226
R29279 DVSS.n20275 DVSS.n20246 3.91226
R29280 DVSS.n20283 DVSS.n20246 3.91226
R29281 DVSS.n20285 DVSS.n20283 3.91226
R29282 DVSS.n20287 DVSS.n20285 3.91226
R29283 DVSS.n20287 DVSS.n20227 3.91226
R29284 DVSS.n20297 DVSS.n20227 3.91226
R29285 DVSS.n20297 DVSS.n20228 3.91226
R29286 DVSS.n20228 DVSS.n20206 3.91226
R29287 DVSS.n20307 DVSS.n20206 3.91226
R29288 DVSS.n20307 DVSS.n20207 3.91226
R29289 DVSS.n20207 DVSS.n20199 3.91226
R29290 DVSS.n20199 DVSS.n14658 3.91226
R29291 DVSS.n20642 DVSS.n14658 3.91226
R29292 DVSS.n20642 DVSS.n14659 3.91226
R29293 DVSS.n20637 DVSS.n14659 3.91226
R29294 DVSS.n20637 DVSS.n14664 3.91226
R29295 DVSS.n20628 DVSS.n14664 3.91226
R29296 DVSS.n20628 DVSS.n14673 3.91226
R29297 DVSS.n20384 DVSS.n14673 3.91226
R29298 DVSS.n20405 DVSS.n20384 3.91226
R29299 DVSS.n20407 DVSS.n20405 3.91226
R29300 DVSS.n20409 DVSS.n20407 3.91226
R29301 DVSS.n20409 DVSS.n20368 3.91226
R29302 DVSS.n20421 DVSS.n20368 3.91226
R29303 DVSS.n20423 DVSS.n20421 3.91226
R29304 DVSS.n20425 DVSS.n20423 3.91226
R29305 DVSS.n20425 DVSS.n20347 3.91226
R29306 DVSS.n20436 DVSS.n20347 3.91226
R29307 DVSS.n20437 DVSS.n20436 3.91226
R29308 DVSS.n20442 DVSS.n20437 3.91226
R29309 DVSS.n20442 DVSS.n20439 3.91226
R29310 DVSS.n20439 DVSS.n20339 3.91226
R29311 DVSS.n20339 DVSS.n14695 3.91226
R29312 DVSS.n20623 DVSS.n14695 3.91226
R29313 DVSS.n20623 DVSS.n14696 3.91226
R29314 DVSS.n20615 DVSS.n14696 3.91226
R29315 DVSS.n18765 DVSS.n18643 3.91226
R29316 DVSS.n18765 DVSS.n18651 3.91226
R29317 DVSS.n18892 DVSS.n18651 3.91226
R29318 DVSS.n18896 DVSS.n18892 3.91226
R29319 DVSS.n18896 DVSS.n18894 3.91226
R29320 DVSS.n18894 DVSS.n18889 3.91226
R29321 DVSS.n18889 DVSS.n14539 3.91226
R29322 DVSS.n20694 DVSS.n14539 3.91226
R29323 DVSS.n20694 DVSS.n14541 3.91226
R29324 DVSS.n18948 DVSS.n14541 3.91226
R29325 DVSS.n18952 DVSS.n18948 3.91226
R29326 DVSS.n18952 DVSS.n18950 3.91226
R29327 DVSS.n18950 DVSS.n18942 3.91226
R29328 DVSS.n18942 DVSS.n18940 3.91226
R29329 DVSS.n18940 DVSS.n18934 3.91226
R29330 DVSS.n18934 DVSS.n18932 3.91226
R29331 DVSS.n18932 DVSS.n18926 3.91226
R29332 DVSS.n18926 DVSS.n18924 3.91226
R29333 DVSS.n18924 DVSS.n18921 3.91226
R29334 DVSS.n18921 DVSS.n14573 3.91226
R29335 DVSS.n20104 DVSS.n14573 3.91226
R29336 DVSS.n20104 DVSS.n14582 3.91226
R29337 DVSS.n20108 DVSS.n14582 3.91226
R29338 DVSS.n20111 DVSS.n20108 3.91226
R29339 DVSS.n20116 DVSS.n20111 3.91226
R29340 DVSS.n20116 DVSS.n20113 3.91226
R29341 DVSS.n20113 DVSS.n20099 3.91226
R29342 DVSS.n20099 DVSS.n20097 3.91226
R29343 DVSS.n20097 DVSS.n20091 3.91226
R29344 DVSS.n20091 DVSS.n20089 3.91226
R29345 DVSS.n20089 DVSS.n20083 3.91226
R29346 DVSS.n20083 DVSS.n20081 3.91226
R29347 DVSS.n20081 DVSS.n20076 3.91226
R29348 DVSS.n20076 DVSS.n20074 3.91226
R29349 DVSS.n20074 DVSS.n20068 3.91226
R29350 DVSS.n20068 DVSS.n20066 3.91226
R29351 DVSS.n20066 DVSS.n20037 3.91226
R29352 DVSS.n20037 DVSS.n20028 3.91226
R29353 DVSS.n20170 DVSS.n20028 3.91226
R29354 DVSS.n20170 DVSS.n20029 3.91226
R29355 DVSS.n20029 DVSS.n14608 3.91226
R29356 DVSS.n20176 DVSS.n14608 3.91226
R29357 DVSS.n20176 DVSS.n14614 3.91226
R29358 DVSS.n20179 DVSS.n14614 3.91226
R29359 DVSS.n20179 DVSS.n14619 3.91226
R29360 DVSS.n20182 DVSS.n14619 3.91226
R29361 DVSS.n20182 DVSS.n14628 3.91226
R29362 DVSS.n20263 DVSS.n14628 3.91226
R29363 DVSS.n20267 DVSS.n20263 3.91226
R29364 DVSS.n20267 DVSS.n20265 3.91226
R29365 DVSS.n20265 DVSS.n20260 3.91226
R29366 DVSS.n20260 DVSS.n20258 3.91226
R29367 DVSS.n20258 DVSS.n20252 3.91226
R29368 DVSS.n20252 DVSS.n20250 3.91226
R29369 DVSS.n20250 DVSS.n20244 3.91226
R29370 DVSS.n20244 DVSS.n20242 3.91226
R29371 DVSS.n20242 DVSS.n20236 3.91226
R29372 DVSS.n20236 DVSS.n20234 3.91226
R29373 DVSS.n20234 DVSS.n20232 3.91226
R29374 DVSS.n20232 DVSS.n20205 3.91226
R29375 DVSS.n20205 DVSS.n20196 3.91226
R29376 DVSS.n20314 DVSS.n20196 3.91226
R29377 DVSS.n20314 DVSS.n20197 3.91226
R29378 DVSS.n20197 DVSS.n14657 3.91226
R29379 DVSS.n20319 DVSS.n14657 3.91226
R29380 DVSS.n20319 DVSS.n14666 3.91226
R29381 DVSS.n20322 DVSS.n14666 3.91226
R29382 DVSS.n20322 DVSS.n14672 3.91226
R29383 DVSS.n20388 DVSS.n14672 3.91226
R29384 DVSS.n20390 DVSS.n20388 3.91226
R29385 DVSS.n20394 DVSS.n20390 3.91226
R29386 DVSS.n20394 DVSS.n20392 3.91226
R29387 DVSS.n20392 DVSS.n20382 3.91226
R29388 DVSS.n20382 DVSS.n20380 3.91226
R29389 DVSS.n20380 DVSS.n20374 3.91226
R29390 DVSS.n20374 DVSS.n20372 3.91226
R29391 DVSS.n20372 DVSS.n20366 3.91226
R29392 DVSS.n20366 DVSS.n20364 3.91226
R29393 DVSS.n20364 DVSS.n20354 3.91226
R29394 DVSS.n20354 DVSS.n20351 3.91226
R29395 DVSS.n20351 DVSS.n20345 3.91226
R29396 DVSS.n20345 DVSS.n20334 3.91226
R29397 DVSS.n20455 DVSS.n20334 3.91226
R29398 DVSS.n20455 DVSS.n20335 3.91226
R29399 DVSS.n20335 DVSS.n14699 3.91226
R29400 DVSS.n20461 DVSS.n14699 3.91226
R29401 DVSS.n20461 DVSS.n14706 3.91226
R29402 DVSS.n18996 DVSS.n18995 3.83228
R29403 DVSS.n18997 DVSS.n18996 3.83228
R29404 DVSS.n20507 DVSS.n20506 3.39586
R29405 DVSS.n20508 DVSS.n20507 3.39586
R29406 DVSS.n14847 DVSS.n14846 3.12476
R29407 DVSS.n14851 DVSS.n14847 3.12476
R29408 DVSS.n19926 DVSS.n15136 2.66791
R29409 DVSS.n20504 DVSS.n20503 2.62838
R29410 DVSS.n20467 DVSS.n20466 2.62838
R29411 DVSS.n20466 DVSS.n14851 2.62235
R29412 DVSS.n20511 DVSS.n20508 2.61801
R29413 DVSS.n20506 DVSS.n20503 2.61724
R29414 DVSS.n18771 DVSS.n18770 2.6005
R29415 DVSS.n18773 DVSS.n18772 2.6005
R29416 DVSS.n18775 DVSS.n18774 2.6005
R29417 DVSS.n18777 DVSS.n18776 2.6005
R29418 DVSS.n18779 DVSS.n18778 2.6005
R29419 DVSS.n18781 DVSS.n18780 2.6005
R29420 DVSS.n18783 DVSS.n18782 2.6005
R29421 DVSS.n18785 DVSS.n18784 2.6005
R29422 DVSS.n18787 DVSS.n18786 2.6005
R29423 DVSS.n18789 DVSS.n18788 2.6005
R29424 DVSS.n18791 DVSS.n18790 2.6005
R29425 DVSS.n18793 DVSS.n18792 2.6005
R29426 DVSS.n18795 DVSS.n18794 2.6005
R29427 DVSS.n18797 DVSS.n18796 2.6005
R29428 DVSS.n18799 DVSS.n18798 2.6005
R29429 DVSS.n18801 DVSS.n18800 2.6005
R29430 DVSS.n18803 DVSS.n18802 2.6005
R29431 DVSS.n18805 DVSS.n18804 2.6005
R29432 DVSS.n18807 DVSS.n18806 2.6005
R29433 DVSS.n18809 DVSS.n18808 2.6005
R29434 DVSS.n18811 DVSS.n18810 2.6005
R29435 DVSS.n18813 DVSS.n18812 2.6005
R29436 DVSS.n18815 DVSS.n18814 2.6005
R29437 DVSS.n18817 DVSS.n18816 2.6005
R29438 DVSS.n18819 DVSS.n18818 2.6005
R29439 DVSS.n18822 DVSS.n18821 2.6005
R29440 DVSS.n18824 DVSS.n18823 2.6005
R29441 DVSS.n18826 DVSS.n18825 2.6005
R29442 DVSS.n18828 DVSS.n18827 2.6005
R29443 DVSS.n18830 DVSS.n18829 2.6005
R29444 DVSS.n18832 DVSS.n18831 2.6005
R29445 DVSS.n18834 DVSS.n18833 2.6005
R29446 DVSS.n18836 DVSS.n18835 2.6005
R29447 DVSS.n18838 DVSS.n18837 2.6005
R29448 DVSS.n18840 DVSS.n18839 2.6005
R29449 DVSS.n18842 DVSS.n18841 2.6005
R29450 DVSS.n18844 DVSS.n18843 2.6005
R29451 DVSS.n18846 DVSS.n18845 2.6005
R29452 DVSS.n18848 DVSS.n18847 2.6005
R29453 DVSS.n18850 DVSS.n18849 2.6005
R29454 DVSS.n18852 DVSS.n18851 2.6005
R29455 DVSS.n18854 DVSS.n18853 2.6005
R29456 DVSS.n18856 DVSS.n18855 2.6005
R29457 DVSS.n18858 DVSS.n18857 2.6005
R29458 DVSS.n18860 DVSS.n18859 2.6005
R29459 DVSS.n18862 DVSS.n18861 2.6005
R29460 DVSS.n18864 DVSS.n18863 2.6005
R29461 DVSS.n18866 DVSS.n18865 2.6005
R29462 DVSS.n18754 DVSS.n18753 2.6005
R29463 DVSS.n18752 DVSS.n18751 2.6005
R29464 DVSS.n18750 DVSS.n18749 2.6005
R29465 DVSS.n18748 DVSS.n18747 2.6005
R29466 DVSS.n18746 DVSS.n18745 2.6005
R29467 DVSS.n18744 DVSS.n18743 2.6005
R29468 DVSS.n18742 DVSS.n18741 2.6005
R29469 DVSS.n18740 DVSS.n18739 2.6005
R29470 DVSS.n18738 DVSS.n18737 2.6005
R29471 DVSS.n18736 DVSS.n18735 2.6005
R29472 DVSS.n18734 DVSS.n18733 2.6005
R29473 DVSS.n18732 DVSS.n18731 2.6005
R29474 DVSS.n18730 DVSS.n18729 2.6005
R29475 DVSS.n18728 DVSS.n18727 2.6005
R29476 DVSS.n18726 DVSS.n18725 2.6005
R29477 DVSS.n18724 DVSS.n18723 2.6005
R29478 DVSS.n18722 DVSS.n18721 2.6005
R29479 DVSS.n18720 DVSS.n18719 2.6005
R29480 DVSS.n18718 DVSS.n18717 2.6005
R29481 DVSS.n18716 DVSS.n18715 2.6005
R29482 DVSS.n18714 DVSS.n18713 2.6005
R29483 DVSS.n18712 DVSS.n18711 2.6005
R29484 DVSS.n18710 DVSS.n18709 2.6005
R29485 DVSS.n18707 DVSS.n18706 2.6005
R29486 DVSS.n18705 DVSS.n18704 2.6005
R29487 DVSS.n18703 DVSS.n18702 2.6005
R29488 DVSS.n18701 DVSS.n18700 2.6005
R29489 DVSS.n18699 DVSS.n18698 2.6005
R29490 DVSS.n18697 DVSS.n18696 2.6005
R29491 DVSS.n18695 DVSS.n18694 2.6005
R29492 DVSS.n18693 DVSS.n18692 2.6005
R29493 DVSS.n18691 DVSS.n18690 2.6005
R29494 DVSS.n18689 DVSS.n18688 2.6005
R29495 DVSS.n18687 DVSS.n18686 2.6005
R29496 DVSS.n18685 DVSS.n18684 2.6005
R29497 DVSS.n18683 DVSS.n18682 2.6005
R29498 DVSS.n18681 DVSS.n18680 2.6005
R29499 DVSS.n18679 DVSS.n18678 2.6005
R29500 DVSS.n18677 DVSS.n18676 2.6005
R29501 DVSS.n18675 DVSS.n18674 2.6005
R29502 DVSS.n18673 DVSS.n18672 2.6005
R29503 DVSS.n18671 DVSS.n18670 2.6005
R29504 DVSS.n18669 DVSS.n18668 2.6005
R29505 DVSS.n18667 DVSS.n18666 2.6005
R29506 DVSS.n18665 DVSS.n18664 2.6005
R29507 DVSS.n18663 DVSS.n18662 2.6005
R29508 DVSS.n18661 DVSS.n18660 2.6005
R29509 DVSS.n18659 DVSS.n18658 2.6005
R29510 DVSS.n18657 DVSS.n18656 2.6005
R29511 DVSS.n20474 DVSS.n20467 2.6005
R29512 DVSS.n20465 DVSS.n20464 2.6005
R29513 DVSS.n20464 DVSS.n14705 2.6005
R29514 DVSS.n20463 DVSS.n14706 2.6005
R29515 DVSS.n20616 DVSS.n14706 2.6005
R29516 DVSS.n20462 DVSS.n20461 2.6005
R29517 DVSS.n20461 DVSS.n14698 2.6005
R29518 DVSS.n20460 DVSS.n14699 2.6005
R29519 DVSS.n20622 DVSS.n14699 2.6005
R29520 DVSS.n20335 DVSS.n14852 2.6005
R29521 DVSS.n20335 DVSS.n14697 2.6005
R29522 DVSS.n20456 DVSS.n20455 2.6005
R29523 DVSS.n20455 DVSS.n20454 2.6005
R29524 DVSS.n20334 DVSS.n20332 2.6005
R29525 DVSS.n20336 DVSS.n20334 2.6005
R29526 DVSS.n20345 DVSS.n20344 2.6005
R29527 DVSS.n20443 DVSS.n20345 2.6005
R29528 DVSS.n20351 DVSS.n20350 2.6005
R29529 DVSS.n20351 DVSS.n20343 2.6005
R29530 DVSS.n20354 DVSS.n20353 2.6005
R29531 DVSS.n20435 DVSS.n20354 2.6005
R29532 DVSS.n20364 DVSS.n20363 2.6005
R29533 DVSS.n20364 DVSS.n20349 2.6005
R29534 DVSS.n20366 DVSS.n20365 2.6005
R29535 DVSS.n20426 DVSS.n20366 2.6005
R29536 DVSS.n20372 DVSS.n20371 2.6005
R29537 DVSS.n20372 DVSS.n20361 2.6005
R29538 DVSS.n20374 DVSS.n20373 2.6005
R29539 DVSS.n20420 DVSS.n20374 2.6005
R29540 DVSS.n20380 DVSS.n20379 2.6005
R29541 DVSS.n20380 DVSS.n20370 2.6005
R29542 DVSS.n20382 DVSS.n20381 2.6005
R29543 DVSS.n20410 DVSS.n20382 2.6005
R29544 DVSS.n20392 DVSS.n20391 2.6005
R29545 DVSS.n20392 DVSS.n20378 2.6005
R29546 DVSS.n20394 DVSS.n20393 2.6005
R29547 DVSS.n20404 DVSS.n20394 2.6005
R29548 DVSS.n20390 DVSS.n20389 2.6005
R29549 DVSS.n20390 DVSS.n20386 2.6005
R29550 DVSS.n20388 DVSS.n20387 2.6005
R29551 DVSS.n20388 DVSS.n14671 2.6005
R29552 DVSS.n20324 DVSS.n14672 2.6005
R29553 DVSS.n20629 DVSS.n14672 2.6005
R29554 DVSS.n20323 DVSS.n20322 2.6005
R29555 DVSS.n20322 DVSS.n14665 2.6005
R29556 DVSS.n20321 DVSS.n14666 2.6005
R29557 DVSS.n20636 DVSS.n14666 2.6005
R29558 DVSS.n20320 DVSS.n20319 2.6005
R29559 DVSS.n20319 DVSS.n14656 2.6005
R29560 DVSS.n20318 DVSS.n14657 2.6005
R29561 DVSS.n20643 DVSS.n14657 2.6005
R29562 DVSS.n20197 DVSS.n14863 2.6005
R29563 DVSS.n20197 DVSS.n14655 2.6005
R29564 DVSS.n20315 DVSS.n20314 2.6005
R29565 DVSS.n20314 DVSS.n20313 2.6005
R29566 DVSS.n20196 DVSS.n20195 2.6005
R29567 DVSS.n20198 DVSS.n20196 2.6005
R29568 DVSS.n20205 DVSS.n20204 2.6005
R29569 DVSS.n20308 DVSS.n20205 2.6005
R29570 DVSS.n20232 DVSS.n20231 2.6005
R29571 DVSS.n20232 DVSS.n20203 2.6005
R29572 DVSS.n20234 DVSS.n20233 2.6005
R29573 DVSS.n20234 DVSS.n20230 2.6005
R29574 DVSS.n20236 DVSS.n20235 2.6005
R29575 DVSS.n20296 DVSS.n20236 2.6005
R29576 DVSS.n20242 DVSS.n20241 2.6005
R29577 DVSS.n20242 DVSS.n20229 2.6005
R29578 DVSS.n20244 DVSS.n20243 2.6005
R29579 DVSS.n20288 DVSS.n20244 2.6005
R29580 DVSS.n20250 DVSS.n20249 2.6005
R29581 DVSS.n20250 DVSS.n20240 2.6005
R29582 DVSS.n20252 DVSS.n20251 2.6005
R29583 DVSS.n20282 DVSS.n20252 2.6005
R29584 DVSS.n20258 DVSS.n20257 2.6005
R29585 DVSS.n20258 DVSS.n20248 2.6005
R29586 DVSS.n20260 DVSS.n20259 2.6005
R29587 DVSS.n20276 DVSS.n20260 2.6005
R29588 DVSS.n20265 DVSS.n20264 2.6005
R29589 DVSS.n20265 DVSS.n20256 2.6005
R29590 DVSS.n20267 DVSS.n20266 2.6005
R29591 DVSS.n20270 DVSS.n20267 2.6005
R29592 DVSS.n20263 DVSS.n20262 2.6005
R29593 DVSS.n20263 DVSS.n14627 2.6005
R29594 DVSS.n20184 DVSS.n14628 2.6005
R29595 DVSS.n20651 DVSS.n14628 2.6005
R29596 DVSS.n20183 DVSS.n20182 2.6005
R29597 DVSS.n20182 DVSS.n14618 2.6005
R29598 DVSS.n20181 DVSS.n14619 2.6005
R29599 DVSS.n20657 DVSS.n14619 2.6005
R29600 DVSS.n20180 DVSS.n20179 2.6005
R29601 DVSS.n20179 DVSS.n14613 2.6005
R29602 DVSS.n20178 DVSS.n14614 2.6005
R29603 DVSS.n20663 DVSS.n14614 2.6005
R29604 DVSS.n20177 DVSS.n20176 2.6005
R29605 DVSS.n20176 DVSS.n14607 2.6005
R29606 DVSS.n20175 DVSS.n14608 2.6005
R29607 DVSS.n20669 DVSS.n14608 2.6005
R29608 DVSS.n20029 DVSS.n14874 2.6005
R29609 DVSS.n20029 DVSS.n14606 2.6005
R29610 DVSS.n20171 DVSS.n20170 2.6005
R29611 DVSS.n20170 DVSS.n20169 2.6005
R29612 DVSS.n20028 DVSS.n20026 2.6005
R29613 DVSS.n20030 DVSS.n20028 2.6005
R29614 DVSS.n20037 DVSS.n20036 2.6005
R29615 DVSS.n20162 DVSS.n20037 2.6005
R29616 DVSS.n20066 DVSS.n20065 2.6005
R29617 DVSS.n20066 DVSS.n20035 2.6005
R29618 DVSS.n20068 DVSS.n20067 2.6005
R29619 DVSS.n20151 DVSS.n20068 2.6005
R29620 DVSS.n20074 DVSS.n20073 2.6005
R29621 DVSS.n20074 DVSS.n20064 2.6005
R29622 DVSS.n20076 DVSS.n20075 2.6005
R29623 DVSS.n20145 DVSS.n20076 2.6005
R29624 DVSS.n20081 DVSS.n20080 2.6005
R29625 DVSS.n20081 DVSS.n20072 2.6005
R29626 DVSS.n20083 DVSS.n20082 2.6005
R29627 DVSS.n20139 DVSS.n20083 2.6005
R29628 DVSS.n20089 DVSS.n20088 2.6005
R29629 DVSS.n20089 DVSS.n20079 2.6005
R29630 DVSS.n20091 DVSS.n20090 2.6005
R29631 DVSS.n20133 DVSS.n20091 2.6005
R29632 DVSS.n20097 DVSS.n20096 2.6005
R29633 DVSS.n20097 DVSS.n20087 2.6005
R29634 DVSS.n20099 DVSS.n20098 2.6005
R29635 DVSS.n20127 DVSS.n20099 2.6005
R29636 DVSS.n20113 DVSS.n20112 2.6005
R29637 DVSS.n20113 DVSS.n20095 2.6005
R29638 DVSS.n20116 DVSS.n20115 2.6005
R29639 DVSS.n20121 DVSS.n20116 2.6005
R29640 DVSS.n20111 DVSS.n20110 2.6005
R29641 DVSS.n20111 DVSS.n20103 2.6005
R29642 DVSS.n20108 DVSS.n20107 2.6005
R29643 DVSS.n20108 DVSS.n14581 2.6005
R29644 DVSS.n20106 DVSS.n14582 2.6005
R29645 DVSS.n20678 DVSS.n14582 2.6005
R29646 DVSS.n20105 DVSS.n20104 2.6005
R29647 DVSS.n20104 DVSS.n14572 2.6005
R29648 DVSS.n14573 DVSS.n14535 2.6005
R29649 DVSS.n20684 DVSS.n14573 2.6005
R29650 DVSS.n18921 DVSS.n14534 2.6005
R29651 DVSS.n18921 DVSS.n14571 2.6005
R29652 DVSS.n18924 DVSS.n18923 2.6005
R29653 DVSS.n18924 DVSS.n18920 2.6005
R29654 DVSS.n18926 DVSS.n18925 2.6005
R29655 DVSS.n18980 DVSS.n18926 2.6005
R29656 DVSS.n18932 DVSS.n18931 2.6005
R29657 DVSS.n18932 DVSS.n18919 2.6005
R29658 DVSS.n18934 DVSS.n18933 2.6005
R29659 DVSS.n18971 DVSS.n18934 2.6005
R29660 DVSS.n18940 DVSS.n18939 2.6005
R29661 DVSS.n18940 DVSS.n18930 2.6005
R29662 DVSS.n18942 DVSS.n18941 2.6005
R29663 DVSS.n18965 DVSS.n18942 2.6005
R29664 DVSS.n18950 DVSS.n18949 2.6005
R29665 DVSS.n18950 DVSS.n18938 2.6005
R29666 DVSS.n18952 DVSS.n18951 2.6005
R29667 DVSS.n18959 DVSS.n18952 2.6005
R29668 DVSS.n18948 DVSS.n18947 2.6005
R29669 DVSS.n18948 DVSS.n18946 2.6005
R29670 DVSS.n14541 DVSS.n14540 2.6005
R29671 DVSS.n14543 DVSS.n14541 2.6005
R29672 DVSS.n20695 DVSS.n20694 2.6005
R29673 DVSS.n20694 DVSS.n20693 2.6005
R29674 DVSS.n14539 DVSS.n14538 2.6005
R29675 DVSS.n14542 DVSS.n14539 2.6005
R29676 DVSS.n18889 DVSS.n18888 2.6005
R29677 DVSS.n18905 DVSS.n18889 2.6005
R29678 DVSS.n18894 DVSS.n18893 2.6005
R29679 DVSS.n18894 DVSS.n18887 2.6005
R29680 DVSS.n18896 DVSS.n18895 2.6005
R29681 DVSS.n18899 DVSS.n18896 2.6005
R29682 DVSS.n18892 DVSS.n18891 2.6005
R29683 DVSS.n18892 DVSS.n18650 2.6005
R29684 DVSS.n18764 DVSS.n18651 2.6005
R29685 DVSS.n18988 DVSS.n18651 2.6005
R29686 DVSS.n18766 DVSS.n18765 2.6005
R29687 DVSS.n18765 DVSS.n18642 2.6005
R29688 DVSS.n18767 DVSS.n18643 2.6005
R29689 DVSS.n18994 DVSS.n18643 2.6005
R29690 DVSS.n14844 DVSS.n14843 2.6005
R29691 DVSS.n14841 DVSS.n14840 2.6005
R29692 DVSS.n14839 DVSS.n14838 2.6005
R29693 DVSS.n14836 DVSS.n14835 2.6005
R29694 DVSS.n14834 DVSS.n14833 2.6005
R29695 DVSS.n14831 DVSS.n14830 2.6005
R29696 DVSS.n14829 DVSS.n14828 2.6005
R29697 DVSS.n14826 DVSS.n14825 2.6005
R29698 DVSS.n14824 DVSS.n14823 2.6005
R29699 DVSS.n14821 DVSS.n14820 2.6005
R29700 DVSS.n14819 DVSS.n14818 2.6005
R29701 DVSS.n14816 DVSS.n14815 2.6005
R29702 DVSS.n14814 DVSS.n14813 2.6005
R29703 DVSS.n14811 DVSS.n14810 2.6005
R29704 DVSS.n14809 DVSS.n14808 2.6005
R29705 DVSS.n14806 DVSS.n14805 2.6005
R29706 DVSS.n14804 DVSS.n14803 2.6005
R29707 DVSS.n14801 DVSS.n14800 2.6005
R29708 DVSS.n14799 DVSS.n14798 2.6005
R29709 DVSS.n14796 DVSS.n14795 2.6005
R29710 DVSS.n14794 DVSS.n14793 2.6005
R29711 DVSS.n14791 DVSS.n14790 2.6005
R29712 DVSS.n14789 DVSS.n14788 2.6005
R29713 DVSS.n14786 DVSS.n14785 2.6005
R29714 DVSS.n14784 DVSS.n14783 2.6005
R29715 DVSS.n14781 DVSS.n14780 2.6005
R29716 DVSS.n14779 DVSS.n14778 2.6005
R29717 DVSS.n14776 DVSS.n14775 2.6005
R29718 DVSS.n14774 DVSS.n14773 2.6005
R29719 DVSS.n14771 DVSS.n14770 2.6005
R29720 DVSS.n14769 DVSS.n14768 2.6005
R29721 DVSS.n14766 DVSS.n14765 2.6005
R29722 DVSS.n14764 DVSS.n14763 2.6005
R29723 DVSS.n14761 DVSS.n14760 2.6005
R29724 DVSS.n14759 DVSS.n14758 2.6005
R29725 DVSS.n14756 DVSS.n14755 2.6005
R29726 DVSS.n14754 DVSS.n14753 2.6005
R29727 DVSS.n14751 DVSS.n14750 2.6005
R29728 DVSS.n14749 DVSS.n14748 2.6005
R29729 DVSS.n14746 DVSS.n14745 2.6005
R29730 DVSS.n14744 DVSS.n14743 2.6005
R29731 DVSS.n14741 DVSS.n14708 2.6005
R29732 DVSS.n20615 DVSS.n20614 2.6005
R29733 DVSS.n20616 DVSS.n20615 2.6005
R29734 DVSS.n14696 DVSS.n14694 2.6005
R29735 DVSS.n14698 DVSS.n14696 2.6005
R29736 DVSS.n20624 DVSS.n20623 2.6005
R29737 DVSS.n20623 DVSS.n20622 2.6005
R29738 DVSS.n14695 DVSS.n14693 2.6005
R29739 DVSS.n14697 DVSS.n14695 2.6005
R29740 DVSS.n20339 DVSS.n20338 2.6005
R29741 DVSS.n20454 DVSS.n20339 2.6005
R29742 DVSS.n20439 DVSS.n20438 2.6005
R29743 DVSS.n20439 DVSS.n20336 2.6005
R29744 DVSS.n20442 DVSS.n20441 2.6005
R29745 DVSS.n20443 DVSS.n20442 2.6005
R29746 DVSS.n20440 DVSS.n20437 2.6005
R29747 DVSS.n20437 DVSS.n20343 2.6005
R29748 DVSS.n20436 DVSS.n20348 2.6005
R29749 DVSS.n20436 DVSS.n20435 2.6005
R29750 DVSS.n20347 DVSS.n20346 2.6005
R29751 DVSS.n20349 DVSS.n20347 2.6005
R29752 DVSS.n20425 DVSS.n20424 2.6005
R29753 DVSS.n20426 DVSS.n20425 2.6005
R29754 DVSS.n20423 DVSS.n20422 2.6005
R29755 DVSS.n20423 DVSS.n20361 2.6005
R29756 DVSS.n20421 DVSS.n20369 2.6005
R29757 DVSS.n20421 DVSS.n20420 2.6005
R29758 DVSS.n20368 DVSS.n20367 2.6005
R29759 DVSS.n20370 DVSS.n20368 2.6005
R29760 DVSS.n20409 DVSS.n20408 2.6005
R29761 DVSS.n20410 DVSS.n20409 2.6005
R29762 DVSS.n20407 DVSS.n20406 2.6005
R29763 DVSS.n20407 DVSS.n20378 2.6005
R29764 DVSS.n20405 DVSS.n20385 2.6005
R29765 DVSS.n20405 DVSS.n20404 2.6005
R29766 DVSS.n20384 DVSS.n20383 2.6005
R29767 DVSS.n20386 DVSS.n20384 2.6005
R29768 DVSS.n14676 DVSS.n14673 2.6005
R29769 DVSS.n14673 DVSS.n14671 2.6005
R29770 DVSS.n20628 DVSS.n20627 2.6005
R29771 DVSS.n20629 DVSS.n20628 2.6005
R29772 DVSS.n14664 DVSS.n14663 2.6005
R29773 DVSS.n14665 DVSS.n14664 2.6005
R29774 DVSS.n20638 DVSS.n20637 2.6005
R29775 DVSS.n20637 DVSS.n20636 2.6005
R29776 DVSS.n20639 DVSS.n14659 2.6005
R29777 DVSS.n14659 DVSS.n14656 2.6005
R29778 DVSS.n20642 DVSS.n20641 2.6005
R29779 DVSS.n20643 DVSS.n20642 2.6005
R29780 DVSS.n20299 DVSS.n14658 2.6005
R29781 DVSS.n14658 DVSS.n14655 2.6005
R29782 DVSS.n20301 DVSS.n20199 2.6005
R29783 DVSS.n20313 DVSS.n20199 2.6005
R29784 DVSS.n20210 DVSS.n20207 2.6005
R29785 DVSS.n20207 DVSS.n20198 2.6005
R29786 DVSS.n20307 DVSS.n20306 2.6005
R29787 DVSS.n20308 DVSS.n20307 2.6005
R29788 DVSS.n20214 DVSS.n20206 2.6005
R29789 DVSS.n20206 DVSS.n20203 2.6005
R29790 DVSS.n20228 DVSS.n20226 2.6005
R29791 DVSS.n20230 DVSS.n20228 2.6005
R29792 DVSS.n20298 DVSS.n20297 2.6005
R29793 DVSS.n20297 DVSS.n20296 2.6005
R29794 DVSS.n20227 DVSS.n20225 2.6005
R29795 DVSS.n20229 DVSS.n20227 2.6005
R29796 DVSS.n20287 DVSS.n20286 2.6005
R29797 DVSS.n20288 DVSS.n20287 2.6005
R29798 DVSS.n20285 DVSS.n20284 2.6005
R29799 DVSS.n20285 DVSS.n20240 2.6005
R29800 DVSS.n20283 DVSS.n20247 2.6005
R29801 DVSS.n20283 DVSS.n20282 2.6005
R29802 DVSS.n20246 DVSS.n20245 2.6005
R29803 DVSS.n20248 DVSS.n20246 2.6005
R29804 DVSS.n20275 DVSS.n20274 2.6005
R29805 DVSS.n20276 DVSS.n20275 2.6005
R29806 DVSS.n20273 DVSS.n20272 2.6005
R29807 DVSS.n20273 DVSS.n20256 2.6005
R29808 DVSS.n20271 DVSS.n20261 2.6005
R29809 DVSS.n20271 DVSS.n20270 2.6005
R29810 DVSS.n20220 DVSS.n14626 2.6005
R29811 DVSS.n14627 DVSS.n14626 2.6005
R29812 DVSS.n20653 DVSS.n20652 2.6005
R29813 DVSS.n20652 DVSS.n20651 2.6005
R29814 DVSS.n20654 DVSS.n14620 2.6005
R29815 DVSS.n14620 DVSS.n14618 2.6005
R29816 DVSS.n20656 DVSS.n20655 2.6005
R29817 DVSS.n20657 DVSS.n20656 2.6005
R29818 DVSS.n14624 DVSS.n14612 2.6005
R29819 DVSS.n14613 DVSS.n14612 2.6005
R29820 DVSS.n20665 DVSS.n20664 2.6005
R29821 DVSS.n20664 DVSS.n20663 2.6005
R29822 DVSS.n20666 DVSS.n14610 2.6005
R29823 DVSS.n14610 DVSS.n14607 2.6005
R29824 DVSS.n20668 DVSS.n20667 2.6005
R29825 DVSS.n20669 DVSS.n20668 2.6005
R29826 DVSS.n14611 DVSS.n14609 2.6005
R29827 DVSS.n14609 DVSS.n14606 2.6005
R29828 DVSS.n20156 DVSS.n20031 2.6005
R29829 DVSS.n20169 DVSS.n20031 2.6005
R29830 DVSS.n20044 DVSS.n20039 2.6005
R29831 DVSS.n20039 DVSS.n20030 2.6005
R29832 DVSS.n20161 DVSS.n20160 2.6005
R29833 DVSS.n20162 DVSS.n20161 2.6005
R29834 DVSS.n20154 DVSS.n20038 2.6005
R29835 DVSS.n20038 DVSS.n20035 2.6005
R29836 DVSS.n20153 DVSS.n20152 2.6005
R29837 DVSS.n20152 DVSS.n20151 2.6005
R29838 DVSS.n20063 DVSS.n20062 2.6005
R29839 DVSS.n20064 DVSS.n20063 2.6005
R29840 DVSS.n20144 DVSS.n20143 2.6005
R29841 DVSS.n20145 DVSS.n20144 2.6005
R29842 DVSS.n20142 DVSS.n20141 2.6005
R29843 DVSS.n20142 DVSS.n20072 2.6005
R29844 DVSS.n20140 DVSS.n20078 2.6005
R29845 DVSS.n20140 DVSS.n20139 2.6005
R29846 DVSS.n20077 DVSS.n20052 2.6005
R29847 DVSS.n20079 DVSS.n20077 2.6005
R29848 DVSS.n20132 DVSS.n20131 2.6005
R29849 DVSS.n20133 DVSS.n20132 2.6005
R29850 DVSS.n20130 DVSS.n20129 2.6005
R29851 DVSS.n20130 DVSS.n20087 2.6005
R29852 DVSS.n20128 DVSS.n20094 2.6005
R29853 DVSS.n20128 DVSS.n20127 2.6005
R29854 DVSS.n20093 DVSS.n20092 2.6005
R29855 DVSS.n20095 DVSS.n20093 2.6005
R29856 DVSS.n20120 DVSS.n20119 2.6005
R29857 DVSS.n20121 DVSS.n20120 2.6005
R29858 DVSS.n20118 DVSS.n20117 2.6005
R29859 DVSS.n20118 DVSS.n20103 2.6005
R29860 DVSS.n20055 DVSS.n14580 2.6005
R29861 DVSS.n14581 DVSS.n14580 2.6005
R29862 DVSS.n20680 DVSS.n20679 2.6005
R29863 DVSS.n20679 DVSS.n20678 2.6005
R29864 DVSS.n20681 DVSS.n14575 2.6005
R29865 DVSS.n14575 DVSS.n14572 2.6005
R29866 DVSS.n20683 DVSS.n20682 2.6005
R29867 DVSS.n20684 DVSS.n20683 2.6005
R29868 DVSS.n14576 DVSS.n14574 2.6005
R29869 DVSS.n14574 DVSS.n14571 2.6005
R29870 DVSS.n18918 DVSS.n18917 2.6005
R29871 DVSS.n18920 DVSS.n18918 2.6005
R29872 DVSS.n18982 DVSS.n18981 2.6005
R29873 DVSS.n18981 DVSS.n18980 2.6005
R29874 DVSS.n18916 DVSS.n18914 2.6005
R29875 DVSS.n18919 DVSS.n18916 2.6005
R29876 DVSS.n18970 DVSS.n18969 2.6005
R29877 DVSS.n18971 DVSS.n18970 2.6005
R29878 DVSS.n18968 DVSS.n18967 2.6005
R29879 DVSS.n18968 DVSS.n18930 2.6005
R29880 DVSS.n18966 DVSS.n18937 2.6005
R29881 DVSS.n18966 DVSS.n18965 2.6005
R29882 DVSS.n18936 DVSS.n18935 2.6005
R29883 DVSS.n18938 DVSS.n18936 2.6005
R29884 DVSS.n18958 DVSS.n18957 2.6005
R29885 DVSS.n18959 DVSS.n18958 2.6005
R29886 DVSS.n18956 DVSS.n18955 2.6005
R29887 DVSS.n18956 DVSS.n18946 2.6005
R29888 DVSS.n18954 DVSS.n18953 2.6005
R29889 DVSS.n18954 DVSS.n14543 2.6005
R29890 DVSS.n18909 DVSS.n14544 2.6005
R29891 DVSS.n20693 DVSS.n14544 2.6005
R29892 DVSS.n18886 DVSS.n18884 2.6005
R29893 DVSS.n18886 DVSS.n14542 2.6005
R29894 DVSS.n18907 DVSS.n18906 2.6005
R29895 DVSS.n18906 DVSS.n18905 2.6005
R29896 DVSS.n18885 DVSS.n18883 2.6005
R29897 DVSS.n18887 DVSS.n18885 2.6005
R29898 DVSS.n18898 DVSS.n18897 2.6005
R29899 DVSS.n18899 DVSS.n18898 2.6005
R29900 DVSS.n18872 DVSS.n18653 2.6005
R29901 DVSS.n18653 DVSS.n18650 2.6005
R29902 DVSS.n18987 DVSS.n18986 2.6005
R29903 DVSS.n18988 DVSS.n18987 2.6005
R29904 DVSS.n18869 DVSS.n18652 2.6005
R29905 DVSS.n18652 DVSS.n18642 2.6005
R29906 DVSS.n18868 DVSS.n18644 2.6005
R29907 DVSS.n18994 DVSS.n18644 2.6005
R29908 DVSS.n20609 DVSS.n14709 2.6005
R29909 DVSS.n20607 DVSS.n20606 2.6005
R29910 DVSS.n20605 DVSS.n20604 2.6005
R29911 DVSS.n20602 DVSS.n20476 2.6005
R29912 DVSS.n20600 DVSS.n20599 2.6005
R29913 DVSS.n20598 DVSS.n20597 2.6005
R29914 DVSS.n20595 DVSS.n20478 2.6005
R29915 DVSS.n20593 DVSS.n20592 2.6005
R29916 DVSS.n20591 DVSS.n20590 2.6005
R29917 DVSS.n20588 DVSS.n20480 2.6005
R29918 DVSS.n20586 DVSS.n20585 2.6005
R29919 DVSS.n20584 DVSS.n20583 2.6005
R29920 DVSS.n20581 DVSS.n20482 2.6005
R29921 DVSS.n20579 DVSS.n20578 2.6005
R29922 DVSS.n20577 DVSS.n20576 2.6005
R29923 DVSS.n20574 DVSS.n20484 2.6005
R29924 DVSS.n20572 DVSS.n20571 2.6005
R29925 DVSS.n20570 DVSS.n20569 2.6005
R29926 DVSS.n20567 DVSS.n20486 2.6005
R29927 DVSS.n20565 DVSS.n20564 2.6005
R29928 DVSS.n20563 DVSS.n20562 2.6005
R29929 DVSS.n20560 DVSS.n20559 2.6005
R29930 DVSS.n20558 DVSS.n20557 2.6005
R29931 DVSS.n20555 DVSS.n20554 2.6005
R29932 DVSS.n20553 DVSS.n20552 2.6005
R29933 DVSS.n20550 DVSS.n20491 2.6005
R29934 DVSS.n20548 DVSS.n20547 2.6005
R29935 DVSS.n20546 DVSS.n20545 2.6005
R29936 DVSS.n20543 DVSS.n20493 2.6005
R29937 DVSS.n20541 DVSS.n20540 2.6005
R29938 DVSS.n20539 DVSS.n20538 2.6005
R29939 DVSS.n20536 DVSS.n20495 2.6005
R29940 DVSS.n20534 DVSS.n20533 2.6005
R29941 DVSS.n20532 DVSS.n20531 2.6005
R29942 DVSS.n20529 DVSS.n20497 2.6005
R29943 DVSS.n20527 DVSS.n20526 2.6005
R29944 DVSS.n20525 DVSS.n20524 2.6005
R29945 DVSS.n20522 DVSS.n20499 2.6005
R29946 DVSS.n20520 DVSS.n20519 2.6005
R29947 DVSS.n20518 DVSS.n20517 2.6005
R29948 DVSS.n20515 DVSS.n20501 2.6005
R29949 DVSS.n20513 DVSS.n20512 2.6005
R29950 DVSS.n20511 DVSS.n20510 2.6005
R29951 DVSS.n20504 DVSS.n20474 2.6005
R29952 DVSS.n14704 DVSS.n14703 2.6005
R29953 DVSS.n14705 DVSS.n14704 2.6005
R29954 DVSS.n20618 DVSS.n20617 2.6005
R29955 DVSS.n20617 DVSS.n20616 2.6005
R29956 DVSS.n20619 DVSS.n14701 2.6005
R29957 DVSS.n14701 DVSS.n14698 2.6005
R29958 DVSS.n20621 DVSS.n20620 2.6005
R29959 DVSS.n20622 DVSS.n20621 2.6005
R29960 DVSS.n20449 DVSS.n14700 2.6005
R29961 DVSS.n14700 DVSS.n14697 2.6005
R29962 DVSS.n20453 DVSS.n20452 2.6005
R29963 DVSS.n20454 DVSS.n20453 2.6005
R29964 DVSS.n20447 DVSS.n20340 2.6005
R29965 DVSS.n20340 DVSS.n20336 2.6005
R29966 DVSS.n20445 DVSS.n20444 2.6005
R29967 DVSS.n20444 DVSS.n20443 2.6005
R29968 DVSS.n20356 DVSS.n20342 2.6005
R29969 DVSS.n20343 DVSS.n20342 2.6005
R29970 DVSS.n20434 DVSS.n20433 2.6005
R29971 DVSS.n20435 DVSS.n20434 2.6005
R29972 DVSS.n20430 DVSS.n20355 2.6005
R29973 DVSS.n20355 DVSS.n20349 2.6005
R29974 DVSS.n20428 DVSS.n20427 2.6005
R29975 DVSS.n20427 DVSS.n20426 2.6005
R29976 DVSS.n20416 DVSS.n20360 2.6005
R29977 DVSS.n20361 DVSS.n20360 2.6005
R29978 DVSS.n20419 DVSS.n20418 2.6005
R29979 DVSS.n20420 DVSS.n20419 2.6005
R29980 DVSS.n20414 DVSS.n20375 2.6005
R29981 DVSS.n20375 DVSS.n20370 2.6005
R29982 DVSS.n20412 DVSS.n20411 2.6005
R29983 DVSS.n20411 DVSS.n20410 2.6005
R29984 DVSS.n20400 DVSS.n20377 2.6005
R29985 DVSS.n20378 DVSS.n20377 2.6005
R29986 DVSS.n20403 DVSS.n20402 2.6005
R29987 DVSS.n20404 DVSS.n20403 2.6005
R29988 DVSS.n20398 DVSS.n20395 2.6005
R29989 DVSS.n20395 DVSS.n20386 2.6005
R29990 DVSS.n20396 DVSS.n14670 2.6005
R29991 DVSS.n14671 DVSS.n14670 2.6005
R29992 DVSS.n20631 DVSS.n20630 2.6005
R29993 DVSS.n20630 DVSS.n20629 2.6005
R29994 DVSS.n20633 DVSS.n14667 2.6005
R29995 DVSS.n14667 DVSS.n14665 2.6005
R29996 DVSS.n20635 DVSS.n20634 2.6005
R29997 DVSS.n20636 DVSS.n20635 2.6005
R29998 DVSS.n14654 DVSS.n14652 2.6005
R29999 DVSS.n14656 DVSS.n14654 2.6005
R30000 DVSS.n20645 DVSS.n20644 2.6005
R30001 DVSS.n20644 DVSS.n20643 2.6005
R30002 DVSS.n14653 DVSS.n14651 2.6005
R30003 DVSS.n14655 DVSS.n14653 2.6005
R30004 DVSS.n20312 DVSS.n14649 2.6005
R30005 DVSS.n20313 DVSS.n20312 2.6005
R30006 DVSS.n20311 DVSS.n20310 2.6005
R30007 DVSS.n20311 DVSS.n20198 2.6005
R30008 DVSS.n20309 DVSS.n20202 2.6005
R30009 DVSS.n20309 DVSS.n20308 2.6005
R30010 DVSS.n20201 DVSS.n20200 2.6005
R30011 DVSS.n20203 DVSS.n20201 2.6005
R30012 DVSS.n20293 DVSS.n20292 2.6005
R30013 DVSS.n20293 DVSS.n20230 2.6005
R30014 DVSS.n20295 DVSS.n20294 2.6005
R30015 DVSS.n20296 DVSS.n20295 2.6005
R30016 DVSS.n20291 DVSS.n20290 2.6005
R30017 DVSS.n20291 DVSS.n20229 2.6005
R30018 DVSS.n20289 DVSS.n20239 2.6005
R30019 DVSS.n20289 DVSS.n20288 2.6005
R30020 DVSS.n20238 DVSS.n20237 2.6005
R30021 DVSS.n20240 DVSS.n20238 2.6005
R30022 DVSS.n20281 DVSS.n20280 2.6005
R30023 DVSS.n20282 DVSS.n20281 2.6005
R30024 DVSS.n20279 DVSS.n20278 2.6005
R30025 DVSS.n20279 DVSS.n20248 2.6005
R30026 DVSS.n20277 DVSS.n20255 2.6005
R30027 DVSS.n20277 DVSS.n20276 2.6005
R30028 DVSS.n20254 DVSS.n20253 2.6005
R30029 DVSS.n20256 DVSS.n20254 2.6005
R30030 DVSS.n20269 DVSS.n20268 2.6005
R30031 DVSS.n20270 DVSS.n20269 2.6005
R30032 DVSS.n14632 DVSS.n14629 2.6005
R30033 DVSS.n14629 DVSS.n14627 2.6005
R30034 DVSS.n20650 DVSS.n20649 2.6005
R30035 DVSS.n20651 DVSS.n20650 2.6005
R30036 DVSS.n14617 DVSS.n14616 2.6005
R30037 DVSS.n14618 DVSS.n14617 2.6005
R30038 DVSS.n20659 DVSS.n20658 2.6005
R30039 DVSS.n20658 DVSS.n20657 2.6005
R30040 DVSS.n20660 DVSS.n14615 2.6005
R30041 DVSS.n14615 DVSS.n14613 2.6005
R30042 DVSS.n20662 DVSS.n20661 2.6005
R30043 DVSS.n20663 DVSS.n20662 2.6005
R30044 DVSS.n14605 DVSS.n14603 2.6005
R30045 DVSS.n14607 DVSS.n14605 2.6005
R30046 DVSS.n20671 DVSS.n20670 2.6005
R30047 DVSS.n20670 DVSS.n20669 2.6005
R30048 DVSS.n14604 DVSS.n14602 2.6005
R30049 DVSS.n14606 DVSS.n14604 2.6005
R30050 DVSS.n20168 DVSS.n20167 2.6005
R30051 DVSS.n20169 DVSS.n20168 2.6005
R30052 DVSS.n20165 DVSS.n20164 2.6005
R30053 DVSS.n20165 DVSS.n20030 2.6005
R30054 DVSS.n20163 DVSS.n20034 2.6005
R30055 DVSS.n20163 DVSS.n20162 2.6005
R30056 DVSS.n20033 DVSS.n20032 2.6005
R30057 DVSS.n20035 DVSS.n20033 2.6005
R30058 DVSS.n20150 DVSS.n20149 2.6005
R30059 DVSS.n20151 DVSS.n20150 2.6005
R30060 DVSS.n20148 DVSS.n20147 2.6005
R30061 DVSS.n20148 DVSS.n20064 2.6005
R30062 DVSS.n20146 DVSS.n20071 2.6005
R30063 DVSS.n20146 DVSS.n20145 2.6005
R30064 DVSS.n20070 DVSS.n20069 2.6005
R30065 DVSS.n20072 DVSS.n20070 2.6005
R30066 DVSS.n20138 DVSS.n20137 2.6005
R30067 DVSS.n20139 DVSS.n20138 2.6005
R30068 DVSS.n20136 DVSS.n20135 2.6005
R30069 DVSS.n20136 DVSS.n20079 2.6005
R30070 DVSS.n20134 DVSS.n20086 2.6005
R30071 DVSS.n20134 DVSS.n20133 2.6005
R30072 DVSS.n20085 DVSS.n20084 2.6005
R30073 DVSS.n20087 DVSS.n20085 2.6005
R30074 DVSS.n20126 DVSS.n20125 2.6005
R30075 DVSS.n20127 DVSS.n20126 2.6005
R30076 DVSS.n20124 DVSS.n20123 2.6005
R30077 DVSS.n20124 DVSS.n20095 2.6005
R30078 DVSS.n20122 DVSS.n20102 2.6005
R30079 DVSS.n20122 DVSS.n20121 2.6005
R30080 DVSS.n20100 DVSS.n14584 2.6005
R30081 DVSS.n20103 DVSS.n20100 2.6005
R30082 DVSS.n20675 DVSS.n14583 2.6005
R30083 DVSS.n14583 DVSS.n14581 2.6005
R30084 DVSS.n20677 DVSS.n20676 2.6005
R30085 DVSS.n20678 DVSS.n20677 2.6005
R30086 DVSS.n14570 DVSS.n14568 2.6005
R30087 DVSS.n14572 DVSS.n14570 2.6005
R30088 DVSS.n20686 DVSS.n20685 2.6005
R30089 DVSS.n20685 DVSS.n20684 2.6005
R30090 DVSS.n14569 DVSS.n14567 2.6005
R30091 DVSS.n14571 DVSS.n14569 2.6005
R30092 DVSS.n18977 DVSS.n18976 2.6005
R30093 DVSS.n18977 DVSS.n18920 2.6005
R30094 DVSS.n18979 DVSS.n18978 2.6005
R30095 DVSS.n18980 DVSS.n18979 2.6005
R30096 DVSS.n18974 DVSS.n18973 2.6005
R30097 DVSS.n18974 DVSS.n18919 2.6005
R30098 DVSS.n18972 DVSS.n18929 2.6005
R30099 DVSS.n18972 DVSS.n18971 2.6005
R30100 DVSS.n18928 DVSS.n18927 2.6005
R30101 DVSS.n18930 DVSS.n18928 2.6005
R30102 DVSS.n18964 DVSS.n18963 2.6005
R30103 DVSS.n18965 DVSS.n18964 2.6005
R30104 DVSS.n18962 DVSS.n18961 2.6005
R30105 DVSS.n18962 DVSS.n18938 2.6005
R30106 DVSS.n18960 DVSS.n18945 2.6005
R30107 DVSS.n18960 DVSS.n18959 2.6005
R30108 DVSS.n18944 DVSS.n18943 2.6005
R30109 DVSS.n18946 DVSS.n18944 2.6005
R30110 DVSS.n14561 DVSS.n14546 2.6005
R30111 DVSS.n14546 DVSS.n14543 2.6005
R30112 DVSS.n20692 DVSS.n20691 2.6005
R30113 DVSS.n20693 DVSS.n20692 2.6005
R30114 DVSS.n14549 DVSS.n14545 2.6005
R30115 DVSS.n14545 DVSS.n14542 2.6005
R30116 DVSS.n18904 DVSS.n18903 2.6005
R30117 DVSS.n18905 DVSS.n18904 2.6005
R30118 DVSS.n18902 DVSS.n18901 2.6005
R30119 DVSS.n18902 DVSS.n18887 2.6005
R30120 DVSS.n18900 DVSS.n18890 2.6005
R30121 DVSS.n18900 DVSS.n18899 2.6005
R30122 DVSS.n18649 DVSS.n18648 2.6005
R30123 DVSS.n18650 DVSS.n18649 2.6005
R30124 DVSS.n18990 DVSS.n18989 2.6005
R30125 DVSS.n18989 DVSS.n18988 2.6005
R30126 DVSS.n18991 DVSS.n18645 2.6005
R30127 DVSS.n18645 DVSS.n18642 2.6005
R30128 DVSS.n18993 DVSS.n18992 2.6005
R30129 DVSS.n18994 DVSS.n18993 2.6005
R30130 DVSS.n18757 DVSS.n18756 2.5974
R30131 DVSS.n20468 DVSS.n14713 2.5974
R30132 DVSS.n22895 DVSS.n22894 2.37282
R30133 DVSS.n22935 DVSS.n22934 2.37282
R30134 DVSS.n22893 DVSS.n22892 2.37282
R30135 DVSS.n22628 DVSS.n736 2.37282
R30136 DVSS.n22627 DVSS.n22626 2.37282
R30137 DVSS.n22587 DVSS.n22586 2.37282
R30138 DVSS.n20506 DVSS.n20505 2.36815
R30139 DVSS.n14851 DVSS.n14850 2.36815
R30140 DVSS.n16493 DVSS.n16492 2.266
R30141 DVSS.n18156 DVSS.n18155 2.26273
R30142 DVSS.n12750 DVSS.n12354 2.25086
R30143 DVSS.n7053 DVSS.n5576 2.2505
R30144 DVSS.n7055 DVSS.n7054 2.2505
R30145 DVSS.n5863 DVSS.n5578 2.2505
R30146 DVSS.n5862 DVSS.n5861 2.2505
R30147 DVSS.n5857 DVSS.n5579 2.2505
R30148 DVSS.n5853 DVSS.n5852 2.2505
R30149 DVSS.n5851 DVSS.n5580 2.2505
R30150 DVSS.n5850 DVSS.n5849 2.2505
R30151 DVSS.n5845 DVSS.n5581 2.2505
R30152 DVSS.n5841 DVSS.n5840 2.2505
R30153 DVSS.n5839 DVSS.n5582 2.2505
R30154 DVSS.n5838 DVSS.n5837 2.2505
R30155 DVSS.n5833 DVSS.n5583 2.2505
R30156 DVSS.n5829 DVSS.n5828 2.2505
R30157 DVSS.n5827 DVSS.n5584 2.2505
R30158 DVSS.n5826 DVSS.n5825 2.2505
R30159 DVSS.n5821 DVSS.n5585 2.2505
R30160 DVSS.n5817 DVSS.n5816 2.2505
R30161 DVSS.n5815 DVSS.n5586 2.2505
R30162 DVSS.n5814 DVSS.n5813 2.2505
R30163 DVSS.n5809 DVSS.n5587 2.2505
R30164 DVSS.n5805 DVSS.n5804 2.2505
R30165 DVSS.n5803 DVSS.n5588 2.2505
R30166 DVSS.n5802 DVSS.n5801 2.2505
R30167 DVSS.n5797 DVSS.n5589 2.2505
R30168 DVSS.n5793 DVSS.n5792 2.2505
R30169 DVSS.n5791 DVSS.n5590 2.2505
R30170 DVSS.n5790 DVSS.n5789 2.2505
R30171 DVSS.n5785 DVSS.n5591 2.2505
R30172 DVSS.n5781 DVSS.n5780 2.2505
R30173 DVSS.n5779 DVSS.n5592 2.2505
R30174 DVSS.n5778 DVSS.n5777 2.2505
R30175 DVSS.n5773 DVSS.n5593 2.2505
R30176 DVSS.n5769 DVSS.n5768 2.2505
R30177 DVSS.n5767 DVSS.n5594 2.2505
R30178 DVSS.n5766 DVSS.n5765 2.2505
R30179 DVSS.n5761 DVSS.n5595 2.2505
R30180 DVSS.n5757 DVSS.n5756 2.2505
R30181 DVSS.n5755 DVSS.n5596 2.2505
R30182 DVSS.n5754 DVSS.n5753 2.2505
R30183 DVSS.n5749 DVSS.n5597 2.2505
R30184 DVSS.n5745 DVSS.n5744 2.2505
R30185 DVSS.n5743 DVSS.n5598 2.2505
R30186 DVSS.n5742 DVSS.n5741 2.2505
R30187 DVSS.n5737 DVSS.n5599 2.2505
R30188 DVSS.n5733 DVSS.n5732 2.2505
R30189 DVSS.n5731 DVSS.n5600 2.2505
R30190 DVSS.n5730 DVSS.n5729 2.2505
R30191 DVSS.n5725 DVSS.n5601 2.2505
R30192 DVSS.n5721 DVSS.n5720 2.2505
R30193 DVSS.n5719 DVSS.n5602 2.2505
R30194 DVSS.n5718 DVSS.n5717 2.2505
R30195 DVSS.n5713 DVSS.n5603 2.2505
R30196 DVSS.n5709 DVSS.n5708 2.2505
R30197 DVSS.n5707 DVSS.n5604 2.2505
R30198 DVSS.n5706 DVSS.n5705 2.2505
R30199 DVSS.n5701 DVSS.n5605 2.2505
R30200 DVSS.n5697 DVSS.n5696 2.2505
R30201 DVSS.n5695 DVSS.n5606 2.2505
R30202 DVSS.n5694 DVSS.n5693 2.2505
R30203 DVSS.n5689 DVSS.n5607 2.2505
R30204 DVSS.n5685 DVSS.n5684 2.2505
R30205 DVSS.n5683 DVSS.n5608 2.2505
R30206 DVSS.n5682 DVSS.n5681 2.2505
R30207 DVSS.n5677 DVSS.n5609 2.2505
R30208 DVSS.n5673 DVSS.n5672 2.2505
R30209 DVSS.n5671 DVSS.n5610 2.2505
R30210 DVSS.n5670 DVSS.n5669 2.2505
R30211 DVSS.n5665 DVSS.n5611 2.2505
R30212 DVSS.n5661 DVSS.n5660 2.2505
R30213 DVSS.n5659 DVSS.n5612 2.2505
R30214 DVSS.n5658 DVSS.n5657 2.2505
R30215 DVSS.n5653 DVSS.n5613 2.2505
R30216 DVSS.n5649 DVSS.n5648 2.2505
R30217 DVSS.n5647 DVSS.n5614 2.2505
R30218 DVSS.n5646 DVSS.n5645 2.2505
R30219 DVSS.n5641 DVSS.n5615 2.2505
R30220 DVSS.n5637 DVSS.n5636 2.2505
R30221 DVSS.n5635 DVSS.n5616 2.2505
R30222 DVSS.n5634 DVSS.n5633 2.2505
R30223 DVSS.n5629 DVSS.n5617 2.2505
R30224 DVSS.n5625 DVSS.n5624 2.2505
R30225 DVSS.n5623 DVSS.n5620 2.2505
R30226 DVSS.n5622 DVSS.n5621 2.2505
R30227 DVSS.n5621 DVSS.n5573 2.2505
R30228 DVSS.n5620 DVSS.n5619 2.2505
R30229 DVSS.n5626 DVSS.n5625 2.2505
R30230 DVSS.n5629 DVSS.n5628 2.2505
R30231 DVSS.n5633 DVSS.n5632 2.2505
R30232 DVSS.n5630 DVSS.n5616 2.2505
R30233 DVSS.n5638 DVSS.n5637 2.2505
R30234 DVSS.n5641 DVSS.n5640 2.2505
R30235 DVSS.n5645 DVSS.n5644 2.2505
R30236 DVSS.n5642 DVSS.n5614 2.2505
R30237 DVSS.n5650 DVSS.n5649 2.2505
R30238 DVSS.n5653 DVSS.n5652 2.2505
R30239 DVSS.n5657 DVSS.n5656 2.2505
R30240 DVSS.n5654 DVSS.n5612 2.2505
R30241 DVSS.n5662 DVSS.n5661 2.2505
R30242 DVSS.n5665 DVSS.n5664 2.2505
R30243 DVSS.n5669 DVSS.n5668 2.2505
R30244 DVSS.n5666 DVSS.n5610 2.2505
R30245 DVSS.n5674 DVSS.n5673 2.2505
R30246 DVSS.n5677 DVSS.n5676 2.2505
R30247 DVSS.n5681 DVSS.n5680 2.2505
R30248 DVSS.n5678 DVSS.n5608 2.2505
R30249 DVSS.n5686 DVSS.n5685 2.2505
R30250 DVSS.n5689 DVSS.n5688 2.2505
R30251 DVSS.n5693 DVSS.n5692 2.2505
R30252 DVSS.n5690 DVSS.n5606 2.2505
R30253 DVSS.n5698 DVSS.n5697 2.2505
R30254 DVSS.n5701 DVSS.n5700 2.2505
R30255 DVSS.n5705 DVSS.n5704 2.2505
R30256 DVSS.n5702 DVSS.n5604 2.2505
R30257 DVSS.n5710 DVSS.n5709 2.2505
R30258 DVSS.n5713 DVSS.n5712 2.2505
R30259 DVSS.n5717 DVSS.n5716 2.2505
R30260 DVSS.n5714 DVSS.n5602 2.2505
R30261 DVSS.n5722 DVSS.n5721 2.2505
R30262 DVSS.n5725 DVSS.n5724 2.2505
R30263 DVSS.n5729 DVSS.n5728 2.2505
R30264 DVSS.n5726 DVSS.n5600 2.2505
R30265 DVSS.n5734 DVSS.n5733 2.2505
R30266 DVSS.n5737 DVSS.n5736 2.2505
R30267 DVSS.n5741 DVSS.n5740 2.2505
R30268 DVSS.n5738 DVSS.n5598 2.2505
R30269 DVSS.n5746 DVSS.n5745 2.2505
R30270 DVSS.n5749 DVSS.n5748 2.2505
R30271 DVSS.n5753 DVSS.n5752 2.2505
R30272 DVSS.n5750 DVSS.n5596 2.2505
R30273 DVSS.n5758 DVSS.n5757 2.2505
R30274 DVSS.n5761 DVSS.n5760 2.2505
R30275 DVSS.n5765 DVSS.n5764 2.2505
R30276 DVSS.n5762 DVSS.n5594 2.2505
R30277 DVSS.n5770 DVSS.n5769 2.2505
R30278 DVSS.n5773 DVSS.n5772 2.2505
R30279 DVSS.n5777 DVSS.n5776 2.2505
R30280 DVSS.n5774 DVSS.n5592 2.2505
R30281 DVSS.n5782 DVSS.n5781 2.2505
R30282 DVSS.n5785 DVSS.n5784 2.2505
R30283 DVSS.n5789 DVSS.n5788 2.2505
R30284 DVSS.n5786 DVSS.n5590 2.2505
R30285 DVSS.n5794 DVSS.n5793 2.2505
R30286 DVSS.n5797 DVSS.n5796 2.2505
R30287 DVSS.n5801 DVSS.n5800 2.2505
R30288 DVSS.n5798 DVSS.n5588 2.2505
R30289 DVSS.n5806 DVSS.n5805 2.2505
R30290 DVSS.n5809 DVSS.n5808 2.2505
R30291 DVSS.n5813 DVSS.n5812 2.2505
R30292 DVSS.n5810 DVSS.n5586 2.2505
R30293 DVSS.n5818 DVSS.n5817 2.2505
R30294 DVSS.n5821 DVSS.n5820 2.2505
R30295 DVSS.n5825 DVSS.n5824 2.2505
R30296 DVSS.n5822 DVSS.n5584 2.2505
R30297 DVSS.n5830 DVSS.n5829 2.2505
R30298 DVSS.n5833 DVSS.n5832 2.2505
R30299 DVSS.n5837 DVSS.n5836 2.2505
R30300 DVSS.n5834 DVSS.n5582 2.2505
R30301 DVSS.n5842 DVSS.n5841 2.2505
R30302 DVSS.n5845 DVSS.n5844 2.2505
R30303 DVSS.n5849 DVSS.n5848 2.2505
R30304 DVSS.n5846 DVSS.n5580 2.2505
R30305 DVSS.n5854 DVSS.n5853 2.2505
R30306 DVSS.n5857 DVSS.n5856 2.2505
R30307 DVSS.n5861 DVSS.n5860 2.2505
R30308 DVSS.n5858 DVSS.n5578 2.2505
R30309 DVSS.n7056 DVSS.n7055 2.2505
R30310 DVSS.n7058 DVSS.n5576 2.2505
R30311 DVSS.n5521 DVSS.n5520 2.2505
R30312 DVSS.n5188 DVSS.n5187 2.2505
R30313 DVSS.n5510 DVSS.n5189 2.2505
R30314 DVSS.n5512 DVSS.n5511 2.2505
R30315 DVSS.n5509 DVSS.n5191 2.2505
R30316 DVSS.n5508 DVSS.n5507 2.2505
R30317 DVSS.n5193 DVSS.n5192 2.2505
R30318 DVSS.n5499 DVSS.n5498 2.2505
R30319 DVSS.n5497 DVSS.n5195 2.2505
R30320 DVSS.n5496 DVSS.n5495 2.2505
R30321 DVSS.n5197 DVSS.n5196 2.2505
R30322 DVSS.n5487 DVSS.n5486 2.2505
R30323 DVSS.n5485 DVSS.n5199 2.2505
R30324 DVSS.n5484 DVSS.n5483 2.2505
R30325 DVSS.n5201 DVSS.n5200 2.2505
R30326 DVSS.n5475 DVSS.n5474 2.2505
R30327 DVSS.n5473 DVSS.n5203 2.2505
R30328 DVSS.n5472 DVSS.n5471 2.2505
R30329 DVSS.n5205 DVSS.n5204 2.2505
R30330 DVSS.n5463 DVSS.n5462 2.2505
R30331 DVSS.n5461 DVSS.n5207 2.2505
R30332 DVSS.n5460 DVSS.n5459 2.2505
R30333 DVSS.n5209 DVSS.n5208 2.2505
R30334 DVSS.n5451 DVSS.n5450 2.2505
R30335 DVSS.n5449 DVSS.n5211 2.2505
R30336 DVSS.n5448 DVSS.n5447 2.2505
R30337 DVSS.n5213 DVSS.n5212 2.2505
R30338 DVSS.n5439 DVSS.n5438 2.2505
R30339 DVSS.n5437 DVSS.n5215 2.2505
R30340 DVSS.n5436 DVSS.n5435 2.2505
R30341 DVSS.n5217 DVSS.n5216 2.2505
R30342 DVSS.n5427 DVSS.n5426 2.2505
R30343 DVSS.n5425 DVSS.n5219 2.2505
R30344 DVSS.n5424 DVSS.n5423 2.2505
R30345 DVSS.n5221 DVSS.n5220 2.2505
R30346 DVSS.n5415 DVSS.n5414 2.2505
R30347 DVSS.n5413 DVSS.n5223 2.2505
R30348 DVSS.n5412 DVSS.n5411 2.2505
R30349 DVSS.n5225 DVSS.n5224 2.2505
R30350 DVSS.n5403 DVSS.n5402 2.2505
R30351 DVSS.n5401 DVSS.n5227 2.2505
R30352 DVSS.n5400 DVSS.n5399 2.2505
R30353 DVSS.n5229 DVSS.n5228 2.2505
R30354 DVSS.n5391 DVSS.n5390 2.2505
R30355 DVSS.n5389 DVSS.n5231 2.2505
R30356 DVSS.n5388 DVSS.n5387 2.2505
R30357 DVSS.n5233 DVSS.n5232 2.2505
R30358 DVSS.n5379 DVSS.n5378 2.2505
R30359 DVSS.n5377 DVSS.n5235 2.2505
R30360 DVSS.n5376 DVSS.n5375 2.2505
R30361 DVSS.n5237 DVSS.n5236 2.2505
R30362 DVSS.n5367 DVSS.n5366 2.2505
R30363 DVSS.n5365 DVSS.n5239 2.2505
R30364 DVSS.n5364 DVSS.n5363 2.2505
R30365 DVSS.n5241 DVSS.n5240 2.2505
R30366 DVSS.n5355 DVSS.n5354 2.2505
R30367 DVSS.n5353 DVSS.n5243 2.2505
R30368 DVSS.n5352 DVSS.n5351 2.2505
R30369 DVSS.n5245 DVSS.n5244 2.2505
R30370 DVSS.n5343 DVSS.n5342 2.2505
R30371 DVSS.n5341 DVSS.n5247 2.2505
R30372 DVSS.n5340 DVSS.n5339 2.2505
R30373 DVSS.n5249 DVSS.n5248 2.2505
R30374 DVSS.n5331 DVSS.n5330 2.2505
R30375 DVSS.n5329 DVSS.n5251 2.2505
R30376 DVSS.n5328 DVSS.n5327 2.2505
R30377 DVSS.n5253 DVSS.n5252 2.2505
R30378 DVSS.n5319 DVSS.n5318 2.2505
R30379 DVSS.n5317 DVSS.n5255 2.2505
R30380 DVSS.n5316 DVSS.n5315 2.2505
R30381 DVSS.n5257 DVSS.n5256 2.2505
R30382 DVSS.n5307 DVSS.n5306 2.2505
R30383 DVSS.n5305 DVSS.n5259 2.2505
R30384 DVSS.n5304 DVSS.n5303 2.2505
R30385 DVSS.n5261 DVSS.n5260 2.2505
R30386 DVSS.n5295 DVSS.n5294 2.2505
R30387 DVSS.n5293 DVSS.n5263 2.2505
R30388 DVSS.n5292 DVSS.n5291 2.2505
R30389 DVSS.n5265 DVSS.n5264 2.2505
R30390 DVSS.n5283 DVSS.n5282 2.2505
R30391 DVSS.n5281 DVSS.n5267 2.2505
R30392 DVSS.n5280 DVSS.n5279 2.2505
R30393 DVSS.n5269 DVSS.n5268 2.2505
R30394 DVSS.n5271 DVSS.n5270 2.2505
R30395 DVSS.n5272 DVSS.n5271 2.2505
R30396 DVSS.n5274 DVSS.n5269 2.2505
R30397 DVSS.n5279 DVSS.n5278 2.2505
R30398 DVSS.n5276 DVSS.n5267 2.2505
R30399 DVSS.n5284 DVSS.n5283 2.2505
R30400 DVSS.n5286 DVSS.n5265 2.2505
R30401 DVSS.n5291 DVSS.n5290 2.2505
R30402 DVSS.n5288 DVSS.n5263 2.2505
R30403 DVSS.n5296 DVSS.n5295 2.2505
R30404 DVSS.n5298 DVSS.n5261 2.2505
R30405 DVSS.n5303 DVSS.n5302 2.2505
R30406 DVSS.n5300 DVSS.n5259 2.2505
R30407 DVSS.n5308 DVSS.n5307 2.2505
R30408 DVSS.n5310 DVSS.n5257 2.2505
R30409 DVSS.n5315 DVSS.n5314 2.2505
R30410 DVSS.n5312 DVSS.n5255 2.2505
R30411 DVSS.n5320 DVSS.n5319 2.2505
R30412 DVSS.n5322 DVSS.n5253 2.2505
R30413 DVSS.n5327 DVSS.n5326 2.2505
R30414 DVSS.n5324 DVSS.n5251 2.2505
R30415 DVSS.n5332 DVSS.n5331 2.2505
R30416 DVSS.n5334 DVSS.n5249 2.2505
R30417 DVSS.n5339 DVSS.n5338 2.2505
R30418 DVSS.n5336 DVSS.n5247 2.2505
R30419 DVSS.n5344 DVSS.n5343 2.2505
R30420 DVSS.n5346 DVSS.n5245 2.2505
R30421 DVSS.n5351 DVSS.n5350 2.2505
R30422 DVSS.n5348 DVSS.n5243 2.2505
R30423 DVSS.n5356 DVSS.n5355 2.2505
R30424 DVSS.n5358 DVSS.n5241 2.2505
R30425 DVSS.n5363 DVSS.n5362 2.2505
R30426 DVSS.n5360 DVSS.n5239 2.2505
R30427 DVSS.n5368 DVSS.n5367 2.2505
R30428 DVSS.n5370 DVSS.n5237 2.2505
R30429 DVSS.n5375 DVSS.n5374 2.2505
R30430 DVSS.n5372 DVSS.n5235 2.2505
R30431 DVSS.n5380 DVSS.n5379 2.2505
R30432 DVSS.n5382 DVSS.n5233 2.2505
R30433 DVSS.n5387 DVSS.n5386 2.2505
R30434 DVSS.n5384 DVSS.n5231 2.2505
R30435 DVSS.n5392 DVSS.n5391 2.2505
R30436 DVSS.n5394 DVSS.n5229 2.2505
R30437 DVSS.n5399 DVSS.n5398 2.2505
R30438 DVSS.n5396 DVSS.n5227 2.2505
R30439 DVSS.n5404 DVSS.n5403 2.2505
R30440 DVSS.n5406 DVSS.n5225 2.2505
R30441 DVSS.n5411 DVSS.n5410 2.2505
R30442 DVSS.n5408 DVSS.n5223 2.2505
R30443 DVSS.n5416 DVSS.n5415 2.2505
R30444 DVSS.n5418 DVSS.n5221 2.2505
R30445 DVSS.n5423 DVSS.n5422 2.2505
R30446 DVSS.n5420 DVSS.n5219 2.2505
R30447 DVSS.n5428 DVSS.n5427 2.2505
R30448 DVSS.n5430 DVSS.n5217 2.2505
R30449 DVSS.n5435 DVSS.n5434 2.2505
R30450 DVSS.n5432 DVSS.n5215 2.2505
R30451 DVSS.n5440 DVSS.n5439 2.2505
R30452 DVSS.n5442 DVSS.n5213 2.2505
R30453 DVSS.n5447 DVSS.n5446 2.2505
R30454 DVSS.n5444 DVSS.n5211 2.2505
R30455 DVSS.n5452 DVSS.n5451 2.2505
R30456 DVSS.n5454 DVSS.n5209 2.2505
R30457 DVSS.n5459 DVSS.n5458 2.2505
R30458 DVSS.n5456 DVSS.n5207 2.2505
R30459 DVSS.n5464 DVSS.n5463 2.2505
R30460 DVSS.n5466 DVSS.n5205 2.2505
R30461 DVSS.n5471 DVSS.n5470 2.2505
R30462 DVSS.n5468 DVSS.n5203 2.2505
R30463 DVSS.n5476 DVSS.n5475 2.2505
R30464 DVSS.n5478 DVSS.n5201 2.2505
R30465 DVSS.n5483 DVSS.n5482 2.2505
R30466 DVSS.n5480 DVSS.n5199 2.2505
R30467 DVSS.n5488 DVSS.n5487 2.2505
R30468 DVSS.n5490 DVSS.n5197 2.2505
R30469 DVSS.n5495 DVSS.n5494 2.2505
R30470 DVSS.n5492 DVSS.n5195 2.2505
R30471 DVSS.n5500 DVSS.n5499 2.2505
R30472 DVSS.n5502 DVSS.n5193 2.2505
R30473 DVSS.n5507 DVSS.n5506 2.2505
R30474 DVSS.n5504 DVSS.n5191 2.2505
R30475 DVSS.n5513 DVSS.n5512 2.2505
R30476 DVSS.n5515 DVSS.n5189 2.2505
R30477 DVSS.n5517 DVSS.n5188 2.2505
R30478 DVSS.n5520 DVSS.n5519 2.2505
R30479 DVSS.n7096 DVSS.n4884 2.2505
R30480 DVSS.n7098 DVSS.n7097 2.2505
R30481 DVSS.n5172 DVSS.n4887 2.2505
R30482 DVSS.n5171 DVSS.n5170 2.2505
R30483 DVSS.n5166 DVSS.n4888 2.2505
R30484 DVSS.n5162 DVSS.n5161 2.2505
R30485 DVSS.n5160 DVSS.n4889 2.2505
R30486 DVSS.n5159 DVSS.n5158 2.2505
R30487 DVSS.n5154 DVSS.n4890 2.2505
R30488 DVSS.n5150 DVSS.n5149 2.2505
R30489 DVSS.n5148 DVSS.n4891 2.2505
R30490 DVSS.n5147 DVSS.n5146 2.2505
R30491 DVSS.n5142 DVSS.n4892 2.2505
R30492 DVSS.n5138 DVSS.n5137 2.2505
R30493 DVSS.n5136 DVSS.n4893 2.2505
R30494 DVSS.n5135 DVSS.n5134 2.2505
R30495 DVSS.n5130 DVSS.n4894 2.2505
R30496 DVSS.n5126 DVSS.n5125 2.2505
R30497 DVSS.n5124 DVSS.n4895 2.2505
R30498 DVSS.n5123 DVSS.n5122 2.2505
R30499 DVSS.n5118 DVSS.n4896 2.2505
R30500 DVSS.n5114 DVSS.n5113 2.2505
R30501 DVSS.n5112 DVSS.n4897 2.2505
R30502 DVSS.n5111 DVSS.n5110 2.2505
R30503 DVSS.n5106 DVSS.n4898 2.2505
R30504 DVSS.n5102 DVSS.n5101 2.2505
R30505 DVSS.n5100 DVSS.n4899 2.2505
R30506 DVSS.n5099 DVSS.n5098 2.2505
R30507 DVSS.n5094 DVSS.n4900 2.2505
R30508 DVSS.n5090 DVSS.n5089 2.2505
R30509 DVSS.n5088 DVSS.n4901 2.2505
R30510 DVSS.n5087 DVSS.n5086 2.2505
R30511 DVSS.n5082 DVSS.n4902 2.2505
R30512 DVSS.n5078 DVSS.n5077 2.2505
R30513 DVSS.n5076 DVSS.n4903 2.2505
R30514 DVSS.n5075 DVSS.n5074 2.2505
R30515 DVSS.n5070 DVSS.n4904 2.2505
R30516 DVSS.n5066 DVSS.n5065 2.2505
R30517 DVSS.n5064 DVSS.n4905 2.2505
R30518 DVSS.n5063 DVSS.n5062 2.2505
R30519 DVSS.n5058 DVSS.n4906 2.2505
R30520 DVSS.n5054 DVSS.n5053 2.2505
R30521 DVSS.n5052 DVSS.n4907 2.2505
R30522 DVSS.n5051 DVSS.n5050 2.2505
R30523 DVSS.n5046 DVSS.n4908 2.2505
R30524 DVSS.n5042 DVSS.n5041 2.2505
R30525 DVSS.n5040 DVSS.n4909 2.2505
R30526 DVSS.n5039 DVSS.n5038 2.2505
R30527 DVSS.n5034 DVSS.n4910 2.2505
R30528 DVSS.n5030 DVSS.n5029 2.2505
R30529 DVSS.n5028 DVSS.n4911 2.2505
R30530 DVSS.n5027 DVSS.n5026 2.2505
R30531 DVSS.n5022 DVSS.n4912 2.2505
R30532 DVSS.n5018 DVSS.n5017 2.2505
R30533 DVSS.n5016 DVSS.n4913 2.2505
R30534 DVSS.n5015 DVSS.n5014 2.2505
R30535 DVSS.n5010 DVSS.n4914 2.2505
R30536 DVSS.n5006 DVSS.n5005 2.2505
R30537 DVSS.n5004 DVSS.n4915 2.2505
R30538 DVSS.n5003 DVSS.n5002 2.2505
R30539 DVSS.n4998 DVSS.n4916 2.2505
R30540 DVSS.n4994 DVSS.n4993 2.2505
R30541 DVSS.n4992 DVSS.n4917 2.2505
R30542 DVSS.n4991 DVSS.n4990 2.2505
R30543 DVSS.n4986 DVSS.n4918 2.2505
R30544 DVSS.n4982 DVSS.n4981 2.2505
R30545 DVSS.n4980 DVSS.n4919 2.2505
R30546 DVSS.n4979 DVSS.n4978 2.2505
R30547 DVSS.n4974 DVSS.n4920 2.2505
R30548 DVSS.n4970 DVSS.n4969 2.2505
R30549 DVSS.n4968 DVSS.n4921 2.2505
R30550 DVSS.n4967 DVSS.n4966 2.2505
R30551 DVSS.n4962 DVSS.n4922 2.2505
R30552 DVSS.n4958 DVSS.n4957 2.2505
R30553 DVSS.n4956 DVSS.n4923 2.2505
R30554 DVSS.n4955 DVSS.n4954 2.2505
R30555 DVSS.n4950 DVSS.n4924 2.2505
R30556 DVSS.n4946 DVSS.n4945 2.2505
R30557 DVSS.n4944 DVSS.n4925 2.2505
R30558 DVSS.n4943 DVSS.n4942 2.2505
R30559 DVSS.n4938 DVSS.n4926 2.2505
R30560 DVSS.n4934 DVSS.n4933 2.2505
R30561 DVSS.n4932 DVSS.n4929 2.2505
R30562 DVSS.n4931 DVSS.n4930 2.2505
R30563 DVSS.n4930 DVSS.n4882 2.2505
R30564 DVSS.n4929 DVSS.n4928 2.2505
R30565 DVSS.n4935 DVSS.n4934 2.2505
R30566 DVSS.n4938 DVSS.n4937 2.2505
R30567 DVSS.n4942 DVSS.n4941 2.2505
R30568 DVSS.n4939 DVSS.n4925 2.2505
R30569 DVSS.n4947 DVSS.n4946 2.2505
R30570 DVSS.n4950 DVSS.n4949 2.2505
R30571 DVSS.n4954 DVSS.n4953 2.2505
R30572 DVSS.n4951 DVSS.n4923 2.2505
R30573 DVSS.n4959 DVSS.n4958 2.2505
R30574 DVSS.n4962 DVSS.n4961 2.2505
R30575 DVSS.n4966 DVSS.n4965 2.2505
R30576 DVSS.n4963 DVSS.n4921 2.2505
R30577 DVSS.n4971 DVSS.n4970 2.2505
R30578 DVSS.n4974 DVSS.n4973 2.2505
R30579 DVSS.n4978 DVSS.n4977 2.2505
R30580 DVSS.n4975 DVSS.n4919 2.2505
R30581 DVSS.n4983 DVSS.n4982 2.2505
R30582 DVSS.n4986 DVSS.n4985 2.2505
R30583 DVSS.n4990 DVSS.n4989 2.2505
R30584 DVSS.n4987 DVSS.n4917 2.2505
R30585 DVSS.n4995 DVSS.n4994 2.2505
R30586 DVSS.n4998 DVSS.n4997 2.2505
R30587 DVSS.n5002 DVSS.n5001 2.2505
R30588 DVSS.n4999 DVSS.n4915 2.2505
R30589 DVSS.n5007 DVSS.n5006 2.2505
R30590 DVSS.n5010 DVSS.n5009 2.2505
R30591 DVSS.n5014 DVSS.n5013 2.2505
R30592 DVSS.n5011 DVSS.n4913 2.2505
R30593 DVSS.n5019 DVSS.n5018 2.2505
R30594 DVSS.n5022 DVSS.n5021 2.2505
R30595 DVSS.n5026 DVSS.n5025 2.2505
R30596 DVSS.n5023 DVSS.n4911 2.2505
R30597 DVSS.n5031 DVSS.n5030 2.2505
R30598 DVSS.n5034 DVSS.n5033 2.2505
R30599 DVSS.n5038 DVSS.n5037 2.2505
R30600 DVSS.n5035 DVSS.n4909 2.2505
R30601 DVSS.n5043 DVSS.n5042 2.2505
R30602 DVSS.n5046 DVSS.n5045 2.2505
R30603 DVSS.n5050 DVSS.n5049 2.2505
R30604 DVSS.n5047 DVSS.n4907 2.2505
R30605 DVSS.n5055 DVSS.n5054 2.2505
R30606 DVSS.n5058 DVSS.n5057 2.2505
R30607 DVSS.n5062 DVSS.n5061 2.2505
R30608 DVSS.n5059 DVSS.n4905 2.2505
R30609 DVSS.n5067 DVSS.n5066 2.2505
R30610 DVSS.n5070 DVSS.n5069 2.2505
R30611 DVSS.n5074 DVSS.n5073 2.2505
R30612 DVSS.n5071 DVSS.n4903 2.2505
R30613 DVSS.n5079 DVSS.n5078 2.2505
R30614 DVSS.n5082 DVSS.n5081 2.2505
R30615 DVSS.n5086 DVSS.n5085 2.2505
R30616 DVSS.n5083 DVSS.n4901 2.2505
R30617 DVSS.n5091 DVSS.n5090 2.2505
R30618 DVSS.n5094 DVSS.n5093 2.2505
R30619 DVSS.n5098 DVSS.n5097 2.2505
R30620 DVSS.n5095 DVSS.n4899 2.2505
R30621 DVSS.n5103 DVSS.n5102 2.2505
R30622 DVSS.n5106 DVSS.n5105 2.2505
R30623 DVSS.n5110 DVSS.n5109 2.2505
R30624 DVSS.n5107 DVSS.n4897 2.2505
R30625 DVSS.n5115 DVSS.n5114 2.2505
R30626 DVSS.n5118 DVSS.n5117 2.2505
R30627 DVSS.n5122 DVSS.n5121 2.2505
R30628 DVSS.n5119 DVSS.n4895 2.2505
R30629 DVSS.n5127 DVSS.n5126 2.2505
R30630 DVSS.n5130 DVSS.n5129 2.2505
R30631 DVSS.n5134 DVSS.n5133 2.2505
R30632 DVSS.n5131 DVSS.n4893 2.2505
R30633 DVSS.n5139 DVSS.n5138 2.2505
R30634 DVSS.n5142 DVSS.n5141 2.2505
R30635 DVSS.n5146 DVSS.n5145 2.2505
R30636 DVSS.n5143 DVSS.n4891 2.2505
R30637 DVSS.n5151 DVSS.n5150 2.2505
R30638 DVSS.n5154 DVSS.n5153 2.2505
R30639 DVSS.n5158 DVSS.n5157 2.2505
R30640 DVSS.n5155 DVSS.n4889 2.2505
R30641 DVSS.n5163 DVSS.n5162 2.2505
R30642 DVSS.n5166 DVSS.n5165 2.2505
R30643 DVSS.n5170 DVSS.n5169 2.2505
R30644 DVSS.n5167 DVSS.n4887 2.2505
R30645 DVSS.n7099 DVSS.n7098 2.2505
R30646 DVSS.n7101 DVSS.n4884 2.2505
R30647 DVSS.n7235 DVSS.n4828 2.2505
R30648 DVSS.n7237 DVSS.n7236 2.2505
R30649 DVSS.n7230 DVSS.n7229 2.2505
R30650 DVSS.n7244 DVSS.n7243 2.2505
R30651 DVSS.n7245 DVSS.n7228 2.2505
R30652 DVSS.n7247 DVSS.n7246 2.2505
R30653 DVSS.n7224 DVSS.n7223 2.2505
R30654 DVSS.n7254 DVSS.n7253 2.2505
R30655 DVSS.n7255 DVSS.n7222 2.2505
R30656 DVSS.n7257 DVSS.n7256 2.2505
R30657 DVSS.n7218 DVSS.n7217 2.2505
R30658 DVSS.n7264 DVSS.n7263 2.2505
R30659 DVSS.n7265 DVSS.n7216 2.2505
R30660 DVSS.n7267 DVSS.n7266 2.2505
R30661 DVSS.n7212 DVSS.n7211 2.2505
R30662 DVSS.n7274 DVSS.n7273 2.2505
R30663 DVSS.n7275 DVSS.n7210 2.2505
R30664 DVSS.n7277 DVSS.n7276 2.2505
R30665 DVSS.n7206 DVSS.n7205 2.2505
R30666 DVSS.n7284 DVSS.n7283 2.2505
R30667 DVSS.n7285 DVSS.n7204 2.2505
R30668 DVSS.n7287 DVSS.n7286 2.2505
R30669 DVSS.n7200 DVSS.n7199 2.2505
R30670 DVSS.n7294 DVSS.n7293 2.2505
R30671 DVSS.n7295 DVSS.n7198 2.2505
R30672 DVSS.n7297 DVSS.n7296 2.2505
R30673 DVSS.n7194 DVSS.n7193 2.2505
R30674 DVSS.n7304 DVSS.n7303 2.2505
R30675 DVSS.n7305 DVSS.n7192 2.2505
R30676 DVSS.n7307 DVSS.n7306 2.2505
R30677 DVSS.n7188 DVSS.n7187 2.2505
R30678 DVSS.n7314 DVSS.n7313 2.2505
R30679 DVSS.n7315 DVSS.n7186 2.2505
R30680 DVSS.n7317 DVSS.n7316 2.2505
R30681 DVSS.n7182 DVSS.n7181 2.2505
R30682 DVSS.n7324 DVSS.n7323 2.2505
R30683 DVSS.n7325 DVSS.n7180 2.2505
R30684 DVSS.n7327 DVSS.n7326 2.2505
R30685 DVSS.n7176 DVSS.n7175 2.2505
R30686 DVSS.n7334 DVSS.n7333 2.2505
R30687 DVSS.n7335 DVSS.n7174 2.2505
R30688 DVSS.n7337 DVSS.n7336 2.2505
R30689 DVSS.n7170 DVSS.n7169 2.2505
R30690 DVSS.n7344 DVSS.n7343 2.2505
R30691 DVSS.n7345 DVSS.n7168 2.2505
R30692 DVSS.n7347 DVSS.n7346 2.2505
R30693 DVSS.n7164 DVSS.n7163 2.2505
R30694 DVSS.n7354 DVSS.n7353 2.2505
R30695 DVSS.n7355 DVSS.n7162 2.2505
R30696 DVSS.n7357 DVSS.n7356 2.2505
R30697 DVSS.n7158 DVSS.n7157 2.2505
R30698 DVSS.n7364 DVSS.n7363 2.2505
R30699 DVSS.n7365 DVSS.n7156 2.2505
R30700 DVSS.n7367 DVSS.n7366 2.2505
R30701 DVSS.n7152 DVSS.n7151 2.2505
R30702 DVSS.n7374 DVSS.n7373 2.2505
R30703 DVSS.n7375 DVSS.n7150 2.2505
R30704 DVSS.n7377 DVSS.n7376 2.2505
R30705 DVSS.n7146 DVSS.n7145 2.2505
R30706 DVSS.n7384 DVSS.n7383 2.2505
R30707 DVSS.n7385 DVSS.n7144 2.2505
R30708 DVSS.n7387 DVSS.n7386 2.2505
R30709 DVSS.n7140 DVSS.n7139 2.2505
R30710 DVSS.n7394 DVSS.n7393 2.2505
R30711 DVSS.n7395 DVSS.n7138 2.2505
R30712 DVSS.n7397 DVSS.n7396 2.2505
R30713 DVSS.n7134 DVSS.n7133 2.2505
R30714 DVSS.n7404 DVSS.n7403 2.2505
R30715 DVSS.n7405 DVSS.n7132 2.2505
R30716 DVSS.n7407 DVSS.n7406 2.2505
R30717 DVSS.n7128 DVSS.n7127 2.2505
R30718 DVSS.n7414 DVSS.n7413 2.2505
R30719 DVSS.n7415 DVSS.n7126 2.2505
R30720 DVSS.n7417 DVSS.n7416 2.2505
R30721 DVSS.n7122 DVSS.n7121 2.2505
R30722 DVSS.n7424 DVSS.n7423 2.2505
R30723 DVSS.n7425 DVSS.n7120 2.2505
R30724 DVSS.n7427 DVSS.n7426 2.2505
R30725 DVSS.n7116 DVSS.n7115 2.2505
R30726 DVSS.n7434 DVSS.n7433 2.2505
R30727 DVSS.n7435 DVSS.n7114 2.2505
R30728 DVSS.n7437 DVSS.n7436 2.2505
R30729 DVSS.n7112 DVSS.n7111 2.2505
R30730 DVSS.n7444 DVSS.n7443 2.2505
R30731 DVSS.n7443 DVSS.n7442 2.2505
R30732 DVSS.n7440 DVSS.n7112 2.2505
R30733 DVSS.n7438 DVSS.n7437 2.2505
R30734 DVSS.n7117 DVSS.n7114 2.2505
R30735 DVSS.n7433 DVSS.n7432 2.2505
R30736 DVSS.n7430 DVSS.n7116 2.2505
R30737 DVSS.n7428 DVSS.n7427 2.2505
R30738 DVSS.n7123 DVSS.n7120 2.2505
R30739 DVSS.n7423 DVSS.n7422 2.2505
R30740 DVSS.n7420 DVSS.n7122 2.2505
R30741 DVSS.n7418 DVSS.n7417 2.2505
R30742 DVSS.n7129 DVSS.n7126 2.2505
R30743 DVSS.n7413 DVSS.n7412 2.2505
R30744 DVSS.n7410 DVSS.n7128 2.2505
R30745 DVSS.n7408 DVSS.n7407 2.2505
R30746 DVSS.n7135 DVSS.n7132 2.2505
R30747 DVSS.n7403 DVSS.n7402 2.2505
R30748 DVSS.n7400 DVSS.n7134 2.2505
R30749 DVSS.n7398 DVSS.n7397 2.2505
R30750 DVSS.n7141 DVSS.n7138 2.2505
R30751 DVSS.n7393 DVSS.n7392 2.2505
R30752 DVSS.n7390 DVSS.n7140 2.2505
R30753 DVSS.n7388 DVSS.n7387 2.2505
R30754 DVSS.n7147 DVSS.n7144 2.2505
R30755 DVSS.n7383 DVSS.n7382 2.2505
R30756 DVSS.n7380 DVSS.n7146 2.2505
R30757 DVSS.n7378 DVSS.n7377 2.2505
R30758 DVSS.n7153 DVSS.n7150 2.2505
R30759 DVSS.n7373 DVSS.n7372 2.2505
R30760 DVSS.n7370 DVSS.n7152 2.2505
R30761 DVSS.n7368 DVSS.n7367 2.2505
R30762 DVSS.n7159 DVSS.n7156 2.2505
R30763 DVSS.n7363 DVSS.n7362 2.2505
R30764 DVSS.n7360 DVSS.n7158 2.2505
R30765 DVSS.n7358 DVSS.n7357 2.2505
R30766 DVSS.n7165 DVSS.n7162 2.2505
R30767 DVSS.n7353 DVSS.n7352 2.2505
R30768 DVSS.n7350 DVSS.n7164 2.2505
R30769 DVSS.n7348 DVSS.n7347 2.2505
R30770 DVSS.n7171 DVSS.n7168 2.2505
R30771 DVSS.n7343 DVSS.n7342 2.2505
R30772 DVSS.n7340 DVSS.n7170 2.2505
R30773 DVSS.n7338 DVSS.n7337 2.2505
R30774 DVSS.n7177 DVSS.n7174 2.2505
R30775 DVSS.n7333 DVSS.n7332 2.2505
R30776 DVSS.n7330 DVSS.n7176 2.2505
R30777 DVSS.n7328 DVSS.n7327 2.2505
R30778 DVSS.n7183 DVSS.n7180 2.2505
R30779 DVSS.n7323 DVSS.n7322 2.2505
R30780 DVSS.n7320 DVSS.n7182 2.2505
R30781 DVSS.n7318 DVSS.n7317 2.2505
R30782 DVSS.n7189 DVSS.n7186 2.2505
R30783 DVSS.n7313 DVSS.n7312 2.2505
R30784 DVSS.n7310 DVSS.n7188 2.2505
R30785 DVSS.n7308 DVSS.n7307 2.2505
R30786 DVSS.n7195 DVSS.n7192 2.2505
R30787 DVSS.n7303 DVSS.n7302 2.2505
R30788 DVSS.n7300 DVSS.n7194 2.2505
R30789 DVSS.n7298 DVSS.n7297 2.2505
R30790 DVSS.n7201 DVSS.n7198 2.2505
R30791 DVSS.n7293 DVSS.n7292 2.2505
R30792 DVSS.n7290 DVSS.n7200 2.2505
R30793 DVSS.n7288 DVSS.n7287 2.2505
R30794 DVSS.n7207 DVSS.n7204 2.2505
R30795 DVSS.n7283 DVSS.n7282 2.2505
R30796 DVSS.n7280 DVSS.n7206 2.2505
R30797 DVSS.n7278 DVSS.n7277 2.2505
R30798 DVSS.n7213 DVSS.n7210 2.2505
R30799 DVSS.n7273 DVSS.n7272 2.2505
R30800 DVSS.n7270 DVSS.n7212 2.2505
R30801 DVSS.n7268 DVSS.n7267 2.2505
R30802 DVSS.n7219 DVSS.n7216 2.2505
R30803 DVSS.n7263 DVSS.n7262 2.2505
R30804 DVSS.n7260 DVSS.n7218 2.2505
R30805 DVSS.n7258 DVSS.n7257 2.2505
R30806 DVSS.n7225 DVSS.n7222 2.2505
R30807 DVSS.n7253 DVSS.n7252 2.2505
R30808 DVSS.n7250 DVSS.n7224 2.2505
R30809 DVSS.n7248 DVSS.n7247 2.2505
R30810 DVSS.n7231 DVSS.n7228 2.2505
R30811 DVSS.n7243 DVSS.n7242 2.2505
R30812 DVSS.n7240 DVSS.n7230 2.2505
R30813 DVSS.n7238 DVSS.n7237 2.2505
R30814 DVSS.n7235 DVSS.n7234 2.2505
R30815 DVSS.n7547 DVSS.n4814 2.2505
R30816 DVSS.n7549 DVSS.n7548 2.2505
R30817 DVSS.n7554 DVSS.n7550 2.2505
R30818 DVSS.n7555 DVSS.n7545 2.2505
R30819 DVSS.n7560 DVSS.n7559 2.2505
R30820 DVSS.n7561 DVSS.n7544 2.2505
R30821 DVSS.n7566 DVSS.n7562 2.2505
R30822 DVSS.n7567 DVSS.n7543 2.2505
R30823 DVSS.n7572 DVSS.n7571 2.2505
R30824 DVSS.n7573 DVSS.n7542 2.2505
R30825 DVSS.n7578 DVSS.n7574 2.2505
R30826 DVSS.n7579 DVSS.n7541 2.2505
R30827 DVSS.n7584 DVSS.n7583 2.2505
R30828 DVSS.n7585 DVSS.n7540 2.2505
R30829 DVSS.n7590 DVSS.n7586 2.2505
R30830 DVSS.n7591 DVSS.n7539 2.2505
R30831 DVSS.n7596 DVSS.n7595 2.2505
R30832 DVSS.n7597 DVSS.n7538 2.2505
R30833 DVSS.n7602 DVSS.n7598 2.2505
R30834 DVSS.n7603 DVSS.n7537 2.2505
R30835 DVSS.n7608 DVSS.n7607 2.2505
R30836 DVSS.n7609 DVSS.n7536 2.2505
R30837 DVSS.n7614 DVSS.n7610 2.2505
R30838 DVSS.n7615 DVSS.n7535 2.2505
R30839 DVSS.n7620 DVSS.n7619 2.2505
R30840 DVSS.n7621 DVSS.n7534 2.2505
R30841 DVSS.n7626 DVSS.n7622 2.2505
R30842 DVSS.n7627 DVSS.n7533 2.2505
R30843 DVSS.n7632 DVSS.n7631 2.2505
R30844 DVSS.n7633 DVSS.n7532 2.2505
R30845 DVSS.n7638 DVSS.n7634 2.2505
R30846 DVSS.n7639 DVSS.n7531 2.2505
R30847 DVSS.n7644 DVSS.n7643 2.2505
R30848 DVSS.n7645 DVSS.n7530 2.2505
R30849 DVSS.n7650 DVSS.n7646 2.2505
R30850 DVSS.n7651 DVSS.n7529 2.2505
R30851 DVSS.n7656 DVSS.n7655 2.2505
R30852 DVSS.n7657 DVSS.n7528 2.2505
R30853 DVSS.n7662 DVSS.n7658 2.2505
R30854 DVSS.n7663 DVSS.n7527 2.2505
R30855 DVSS.n7668 DVSS.n7667 2.2505
R30856 DVSS.n7669 DVSS.n7526 2.2505
R30857 DVSS.n7674 DVSS.n7670 2.2505
R30858 DVSS.n7675 DVSS.n7525 2.2505
R30859 DVSS.n7680 DVSS.n7679 2.2505
R30860 DVSS.n7681 DVSS.n7524 2.2505
R30861 DVSS.n7686 DVSS.n7682 2.2505
R30862 DVSS.n7687 DVSS.n7523 2.2505
R30863 DVSS.n7692 DVSS.n7691 2.2505
R30864 DVSS.n7693 DVSS.n7522 2.2505
R30865 DVSS.n7698 DVSS.n7694 2.2505
R30866 DVSS.n7699 DVSS.n7521 2.2505
R30867 DVSS.n7704 DVSS.n7703 2.2505
R30868 DVSS.n7705 DVSS.n7520 2.2505
R30869 DVSS.n7710 DVSS.n7706 2.2505
R30870 DVSS.n7711 DVSS.n7519 2.2505
R30871 DVSS.n7716 DVSS.n7715 2.2505
R30872 DVSS.n7717 DVSS.n7518 2.2505
R30873 DVSS.n7722 DVSS.n7718 2.2505
R30874 DVSS.n7723 DVSS.n7517 2.2505
R30875 DVSS.n7728 DVSS.n7727 2.2505
R30876 DVSS.n7729 DVSS.n7516 2.2505
R30877 DVSS.n7734 DVSS.n7730 2.2505
R30878 DVSS.n7735 DVSS.n7515 2.2505
R30879 DVSS.n7740 DVSS.n7739 2.2505
R30880 DVSS.n7741 DVSS.n7514 2.2505
R30881 DVSS.n7746 DVSS.n7742 2.2505
R30882 DVSS.n7747 DVSS.n7513 2.2505
R30883 DVSS.n7752 DVSS.n7751 2.2505
R30884 DVSS.n7753 DVSS.n7512 2.2505
R30885 DVSS.n7758 DVSS.n7754 2.2505
R30886 DVSS.n7759 DVSS.n7511 2.2505
R30887 DVSS.n7764 DVSS.n7763 2.2505
R30888 DVSS.n7765 DVSS.n7510 2.2505
R30889 DVSS.n7770 DVSS.n7766 2.2505
R30890 DVSS.n7771 DVSS.n7509 2.2505
R30891 DVSS.n7776 DVSS.n7775 2.2505
R30892 DVSS.n7777 DVSS.n7508 2.2505
R30893 DVSS.n7782 DVSS.n7778 2.2505
R30894 DVSS.n7783 DVSS.n7507 2.2505
R30895 DVSS.n7788 DVSS.n7787 2.2505
R30896 DVSS.n7789 DVSS.n7506 2.2505
R30897 DVSS.n7791 DVSS.n7790 2.2505
R30898 DVSS.n7792 DVSS.n4821 2.2505
R30899 DVSS.n7793 DVSS.n7792 2.2505
R30900 DVSS.n7791 DVSS.n7503 2.2505
R30901 DVSS.n7506 DVSS.n7505 2.2505
R30902 DVSS.n7787 DVSS.n7786 2.2505
R30903 DVSS.n7784 DVSS.n7783 2.2505
R30904 DVSS.n7782 DVSS.n7781 2.2505
R30905 DVSS.n7779 DVSS.n7508 2.2505
R30906 DVSS.n7775 DVSS.n7774 2.2505
R30907 DVSS.n7772 DVSS.n7771 2.2505
R30908 DVSS.n7770 DVSS.n7769 2.2505
R30909 DVSS.n7767 DVSS.n7510 2.2505
R30910 DVSS.n7763 DVSS.n7762 2.2505
R30911 DVSS.n7760 DVSS.n7759 2.2505
R30912 DVSS.n7758 DVSS.n7757 2.2505
R30913 DVSS.n7755 DVSS.n7512 2.2505
R30914 DVSS.n7751 DVSS.n7750 2.2505
R30915 DVSS.n7748 DVSS.n7747 2.2505
R30916 DVSS.n7746 DVSS.n7745 2.2505
R30917 DVSS.n7743 DVSS.n7514 2.2505
R30918 DVSS.n7739 DVSS.n7738 2.2505
R30919 DVSS.n7736 DVSS.n7735 2.2505
R30920 DVSS.n7734 DVSS.n7733 2.2505
R30921 DVSS.n7731 DVSS.n7516 2.2505
R30922 DVSS.n7727 DVSS.n7726 2.2505
R30923 DVSS.n7724 DVSS.n7723 2.2505
R30924 DVSS.n7722 DVSS.n7721 2.2505
R30925 DVSS.n7719 DVSS.n7518 2.2505
R30926 DVSS.n7715 DVSS.n7714 2.2505
R30927 DVSS.n7712 DVSS.n7711 2.2505
R30928 DVSS.n7710 DVSS.n7709 2.2505
R30929 DVSS.n7707 DVSS.n7520 2.2505
R30930 DVSS.n7703 DVSS.n7702 2.2505
R30931 DVSS.n7700 DVSS.n7699 2.2505
R30932 DVSS.n7698 DVSS.n7697 2.2505
R30933 DVSS.n7695 DVSS.n7522 2.2505
R30934 DVSS.n7691 DVSS.n7690 2.2505
R30935 DVSS.n7688 DVSS.n7687 2.2505
R30936 DVSS.n7686 DVSS.n7685 2.2505
R30937 DVSS.n7683 DVSS.n7524 2.2505
R30938 DVSS.n7679 DVSS.n7678 2.2505
R30939 DVSS.n7676 DVSS.n7675 2.2505
R30940 DVSS.n7674 DVSS.n7673 2.2505
R30941 DVSS.n7671 DVSS.n7526 2.2505
R30942 DVSS.n7667 DVSS.n7666 2.2505
R30943 DVSS.n7664 DVSS.n7663 2.2505
R30944 DVSS.n7662 DVSS.n7661 2.2505
R30945 DVSS.n7659 DVSS.n7528 2.2505
R30946 DVSS.n7655 DVSS.n7654 2.2505
R30947 DVSS.n7652 DVSS.n7651 2.2505
R30948 DVSS.n7650 DVSS.n7649 2.2505
R30949 DVSS.n7647 DVSS.n7530 2.2505
R30950 DVSS.n7643 DVSS.n7642 2.2505
R30951 DVSS.n7640 DVSS.n7639 2.2505
R30952 DVSS.n7638 DVSS.n7637 2.2505
R30953 DVSS.n7635 DVSS.n7532 2.2505
R30954 DVSS.n7631 DVSS.n7630 2.2505
R30955 DVSS.n7628 DVSS.n7627 2.2505
R30956 DVSS.n7626 DVSS.n7625 2.2505
R30957 DVSS.n7623 DVSS.n7534 2.2505
R30958 DVSS.n7619 DVSS.n7618 2.2505
R30959 DVSS.n7616 DVSS.n7615 2.2505
R30960 DVSS.n7614 DVSS.n7613 2.2505
R30961 DVSS.n7611 DVSS.n7536 2.2505
R30962 DVSS.n7607 DVSS.n7606 2.2505
R30963 DVSS.n7604 DVSS.n7603 2.2505
R30964 DVSS.n7602 DVSS.n7601 2.2505
R30965 DVSS.n7599 DVSS.n7538 2.2505
R30966 DVSS.n7595 DVSS.n7594 2.2505
R30967 DVSS.n7592 DVSS.n7591 2.2505
R30968 DVSS.n7590 DVSS.n7589 2.2505
R30969 DVSS.n7587 DVSS.n7540 2.2505
R30970 DVSS.n7583 DVSS.n7582 2.2505
R30971 DVSS.n7580 DVSS.n7579 2.2505
R30972 DVSS.n7578 DVSS.n7577 2.2505
R30973 DVSS.n7575 DVSS.n7542 2.2505
R30974 DVSS.n7571 DVSS.n7570 2.2505
R30975 DVSS.n7568 DVSS.n7567 2.2505
R30976 DVSS.n7566 DVSS.n7565 2.2505
R30977 DVSS.n7563 DVSS.n7544 2.2505
R30978 DVSS.n7559 DVSS.n7558 2.2505
R30979 DVSS.n7556 DVSS.n7555 2.2505
R30980 DVSS.n7554 DVSS.n7553 2.2505
R30981 DVSS.n7551 DVSS.n7548 2.2505
R30982 DVSS.n7547 DVSS.n7546 2.2505
R30983 DVSS.n4598 DVSS.n4462 2.2505
R30984 DVSS.n4600 DVSS.n4599 2.2505
R30985 DVSS.n4593 DVSS.n4592 2.2505
R30986 DVSS.n4607 DVSS.n4606 2.2505
R30987 DVSS.n4608 DVSS.n4591 2.2505
R30988 DVSS.n4610 DVSS.n4609 2.2505
R30989 DVSS.n4587 DVSS.n4586 2.2505
R30990 DVSS.n4617 DVSS.n4616 2.2505
R30991 DVSS.n4618 DVSS.n4585 2.2505
R30992 DVSS.n4620 DVSS.n4619 2.2505
R30993 DVSS.n4581 DVSS.n4580 2.2505
R30994 DVSS.n4627 DVSS.n4626 2.2505
R30995 DVSS.n4628 DVSS.n4579 2.2505
R30996 DVSS.n4630 DVSS.n4629 2.2505
R30997 DVSS.n4575 DVSS.n4574 2.2505
R30998 DVSS.n4637 DVSS.n4636 2.2505
R30999 DVSS.n4638 DVSS.n4573 2.2505
R31000 DVSS.n4640 DVSS.n4639 2.2505
R31001 DVSS.n4569 DVSS.n4568 2.2505
R31002 DVSS.n4647 DVSS.n4646 2.2505
R31003 DVSS.n4648 DVSS.n4567 2.2505
R31004 DVSS.n4650 DVSS.n4649 2.2505
R31005 DVSS.n4563 DVSS.n4562 2.2505
R31006 DVSS.n4657 DVSS.n4656 2.2505
R31007 DVSS.n4658 DVSS.n4561 2.2505
R31008 DVSS.n4660 DVSS.n4659 2.2505
R31009 DVSS.n4557 DVSS.n4556 2.2505
R31010 DVSS.n4667 DVSS.n4666 2.2505
R31011 DVSS.n4668 DVSS.n4555 2.2505
R31012 DVSS.n4670 DVSS.n4669 2.2505
R31013 DVSS.n4551 DVSS.n4550 2.2505
R31014 DVSS.n4677 DVSS.n4676 2.2505
R31015 DVSS.n4678 DVSS.n4549 2.2505
R31016 DVSS.n4680 DVSS.n4679 2.2505
R31017 DVSS.n4545 DVSS.n4544 2.2505
R31018 DVSS.n4687 DVSS.n4686 2.2505
R31019 DVSS.n4688 DVSS.n4543 2.2505
R31020 DVSS.n4690 DVSS.n4689 2.2505
R31021 DVSS.n4539 DVSS.n4538 2.2505
R31022 DVSS.n4697 DVSS.n4696 2.2505
R31023 DVSS.n4698 DVSS.n4537 2.2505
R31024 DVSS.n4700 DVSS.n4699 2.2505
R31025 DVSS.n4533 DVSS.n4532 2.2505
R31026 DVSS.n4707 DVSS.n4706 2.2505
R31027 DVSS.n4708 DVSS.n4531 2.2505
R31028 DVSS.n4710 DVSS.n4709 2.2505
R31029 DVSS.n4527 DVSS.n4526 2.2505
R31030 DVSS.n4717 DVSS.n4716 2.2505
R31031 DVSS.n4718 DVSS.n4525 2.2505
R31032 DVSS.n4720 DVSS.n4719 2.2505
R31033 DVSS.n4521 DVSS.n4520 2.2505
R31034 DVSS.n4727 DVSS.n4726 2.2505
R31035 DVSS.n4728 DVSS.n4519 2.2505
R31036 DVSS.n4730 DVSS.n4729 2.2505
R31037 DVSS.n4515 DVSS.n4514 2.2505
R31038 DVSS.n4737 DVSS.n4736 2.2505
R31039 DVSS.n4738 DVSS.n4513 2.2505
R31040 DVSS.n4740 DVSS.n4739 2.2505
R31041 DVSS.n4509 DVSS.n4508 2.2505
R31042 DVSS.n4747 DVSS.n4746 2.2505
R31043 DVSS.n4748 DVSS.n4507 2.2505
R31044 DVSS.n4750 DVSS.n4749 2.2505
R31045 DVSS.n4503 DVSS.n4502 2.2505
R31046 DVSS.n4757 DVSS.n4756 2.2505
R31047 DVSS.n4758 DVSS.n4501 2.2505
R31048 DVSS.n4760 DVSS.n4759 2.2505
R31049 DVSS.n4497 DVSS.n4496 2.2505
R31050 DVSS.n4767 DVSS.n4766 2.2505
R31051 DVSS.n4768 DVSS.n4495 2.2505
R31052 DVSS.n4770 DVSS.n4769 2.2505
R31053 DVSS.n4491 DVSS.n4490 2.2505
R31054 DVSS.n4777 DVSS.n4776 2.2505
R31055 DVSS.n4778 DVSS.n4489 2.2505
R31056 DVSS.n4780 DVSS.n4779 2.2505
R31057 DVSS.n4485 DVSS.n4484 2.2505
R31058 DVSS.n4787 DVSS.n4786 2.2505
R31059 DVSS.n4788 DVSS.n4483 2.2505
R31060 DVSS.n4790 DVSS.n4789 2.2505
R31061 DVSS.n4479 DVSS.n4478 2.2505
R31062 DVSS.n4797 DVSS.n4796 2.2505
R31063 DVSS.n4798 DVSS.n4477 2.2505
R31064 DVSS.n4800 DVSS.n4799 2.2505
R31065 DVSS.n4475 DVSS.n4474 2.2505
R31066 DVSS.n4807 DVSS.n4806 2.2505
R31067 DVSS.n4806 DVSS.n4805 2.2505
R31068 DVSS.n4803 DVSS.n4475 2.2505
R31069 DVSS.n4801 DVSS.n4800 2.2505
R31070 DVSS.n4480 DVSS.n4477 2.2505
R31071 DVSS.n4796 DVSS.n4795 2.2505
R31072 DVSS.n4793 DVSS.n4479 2.2505
R31073 DVSS.n4791 DVSS.n4790 2.2505
R31074 DVSS.n4486 DVSS.n4483 2.2505
R31075 DVSS.n4786 DVSS.n4785 2.2505
R31076 DVSS.n4783 DVSS.n4485 2.2505
R31077 DVSS.n4781 DVSS.n4780 2.2505
R31078 DVSS.n4492 DVSS.n4489 2.2505
R31079 DVSS.n4776 DVSS.n4775 2.2505
R31080 DVSS.n4773 DVSS.n4491 2.2505
R31081 DVSS.n4771 DVSS.n4770 2.2505
R31082 DVSS.n4498 DVSS.n4495 2.2505
R31083 DVSS.n4766 DVSS.n4765 2.2505
R31084 DVSS.n4763 DVSS.n4497 2.2505
R31085 DVSS.n4761 DVSS.n4760 2.2505
R31086 DVSS.n4504 DVSS.n4501 2.2505
R31087 DVSS.n4756 DVSS.n4755 2.2505
R31088 DVSS.n4753 DVSS.n4503 2.2505
R31089 DVSS.n4751 DVSS.n4750 2.2505
R31090 DVSS.n4510 DVSS.n4507 2.2505
R31091 DVSS.n4746 DVSS.n4745 2.2505
R31092 DVSS.n4743 DVSS.n4509 2.2505
R31093 DVSS.n4741 DVSS.n4740 2.2505
R31094 DVSS.n4516 DVSS.n4513 2.2505
R31095 DVSS.n4736 DVSS.n4735 2.2505
R31096 DVSS.n4733 DVSS.n4515 2.2505
R31097 DVSS.n4731 DVSS.n4730 2.2505
R31098 DVSS.n4522 DVSS.n4519 2.2505
R31099 DVSS.n4726 DVSS.n4725 2.2505
R31100 DVSS.n4723 DVSS.n4521 2.2505
R31101 DVSS.n4721 DVSS.n4720 2.2505
R31102 DVSS.n4528 DVSS.n4525 2.2505
R31103 DVSS.n4716 DVSS.n4715 2.2505
R31104 DVSS.n4713 DVSS.n4527 2.2505
R31105 DVSS.n4711 DVSS.n4710 2.2505
R31106 DVSS.n4534 DVSS.n4531 2.2505
R31107 DVSS.n4706 DVSS.n4705 2.2505
R31108 DVSS.n4703 DVSS.n4533 2.2505
R31109 DVSS.n4701 DVSS.n4700 2.2505
R31110 DVSS.n4540 DVSS.n4537 2.2505
R31111 DVSS.n4696 DVSS.n4695 2.2505
R31112 DVSS.n4693 DVSS.n4539 2.2505
R31113 DVSS.n4691 DVSS.n4690 2.2505
R31114 DVSS.n4546 DVSS.n4543 2.2505
R31115 DVSS.n4686 DVSS.n4685 2.2505
R31116 DVSS.n4683 DVSS.n4545 2.2505
R31117 DVSS.n4681 DVSS.n4680 2.2505
R31118 DVSS.n4552 DVSS.n4549 2.2505
R31119 DVSS.n4676 DVSS.n4675 2.2505
R31120 DVSS.n4673 DVSS.n4551 2.2505
R31121 DVSS.n4671 DVSS.n4670 2.2505
R31122 DVSS.n4558 DVSS.n4555 2.2505
R31123 DVSS.n4666 DVSS.n4665 2.2505
R31124 DVSS.n4663 DVSS.n4557 2.2505
R31125 DVSS.n4661 DVSS.n4660 2.2505
R31126 DVSS.n4564 DVSS.n4561 2.2505
R31127 DVSS.n4656 DVSS.n4655 2.2505
R31128 DVSS.n4653 DVSS.n4563 2.2505
R31129 DVSS.n4651 DVSS.n4650 2.2505
R31130 DVSS.n4570 DVSS.n4567 2.2505
R31131 DVSS.n4646 DVSS.n4645 2.2505
R31132 DVSS.n4643 DVSS.n4569 2.2505
R31133 DVSS.n4641 DVSS.n4640 2.2505
R31134 DVSS.n4576 DVSS.n4573 2.2505
R31135 DVSS.n4636 DVSS.n4635 2.2505
R31136 DVSS.n4633 DVSS.n4575 2.2505
R31137 DVSS.n4631 DVSS.n4630 2.2505
R31138 DVSS.n4582 DVSS.n4579 2.2505
R31139 DVSS.n4626 DVSS.n4625 2.2505
R31140 DVSS.n4623 DVSS.n4581 2.2505
R31141 DVSS.n4621 DVSS.n4620 2.2505
R31142 DVSS.n4588 DVSS.n4585 2.2505
R31143 DVSS.n4616 DVSS.n4615 2.2505
R31144 DVSS.n4613 DVSS.n4587 2.2505
R31145 DVSS.n4611 DVSS.n4610 2.2505
R31146 DVSS.n4594 DVSS.n4591 2.2505
R31147 DVSS.n4606 DVSS.n4605 2.2505
R31148 DVSS.n4603 DVSS.n4593 2.2505
R31149 DVSS.n4601 DVSS.n4600 2.2505
R31150 DVSS.n4598 DVSS.n4597 2.2505
R31151 DVSS.n7843 DVSS.n7842 2.2505
R31152 DVSS.n7844 DVSS.n4457 2.2505
R31153 DVSS.n7849 DVSS.n7845 2.2505
R31154 DVSS.n7850 DVSS.n4456 2.2505
R31155 DVSS.n7855 DVSS.n7854 2.2505
R31156 DVSS.n7856 DVSS.n4455 2.2505
R31157 DVSS.n7861 DVSS.n7857 2.2505
R31158 DVSS.n7862 DVSS.n4454 2.2505
R31159 DVSS.n7867 DVSS.n7866 2.2505
R31160 DVSS.n7868 DVSS.n4453 2.2505
R31161 DVSS.n7873 DVSS.n7869 2.2505
R31162 DVSS.n7874 DVSS.n4452 2.2505
R31163 DVSS.n7879 DVSS.n7878 2.2505
R31164 DVSS.n7880 DVSS.n4451 2.2505
R31165 DVSS.n7885 DVSS.n7881 2.2505
R31166 DVSS.n7886 DVSS.n4450 2.2505
R31167 DVSS.n7891 DVSS.n7890 2.2505
R31168 DVSS.n7892 DVSS.n4449 2.2505
R31169 DVSS.n7897 DVSS.n7893 2.2505
R31170 DVSS.n7898 DVSS.n4448 2.2505
R31171 DVSS.n7903 DVSS.n7902 2.2505
R31172 DVSS.n7904 DVSS.n4447 2.2505
R31173 DVSS.n7909 DVSS.n7905 2.2505
R31174 DVSS.n7910 DVSS.n4446 2.2505
R31175 DVSS.n7915 DVSS.n7914 2.2505
R31176 DVSS.n7916 DVSS.n4445 2.2505
R31177 DVSS.n7921 DVSS.n7917 2.2505
R31178 DVSS.n7922 DVSS.n4444 2.2505
R31179 DVSS.n7927 DVSS.n7926 2.2505
R31180 DVSS.n7928 DVSS.n4443 2.2505
R31181 DVSS.n7933 DVSS.n7929 2.2505
R31182 DVSS.n7934 DVSS.n4442 2.2505
R31183 DVSS.n7939 DVSS.n7938 2.2505
R31184 DVSS.n7940 DVSS.n4441 2.2505
R31185 DVSS.n7945 DVSS.n7941 2.2505
R31186 DVSS.n7946 DVSS.n4440 2.2505
R31187 DVSS.n7951 DVSS.n7950 2.2505
R31188 DVSS.n7952 DVSS.n4439 2.2505
R31189 DVSS.n7957 DVSS.n7953 2.2505
R31190 DVSS.n7958 DVSS.n4438 2.2505
R31191 DVSS.n7963 DVSS.n7962 2.2505
R31192 DVSS.n7964 DVSS.n4437 2.2505
R31193 DVSS.n7969 DVSS.n7965 2.2505
R31194 DVSS.n7970 DVSS.n4436 2.2505
R31195 DVSS.n7975 DVSS.n7974 2.2505
R31196 DVSS.n7976 DVSS.n4435 2.2505
R31197 DVSS.n7981 DVSS.n7977 2.2505
R31198 DVSS.n7982 DVSS.n4434 2.2505
R31199 DVSS.n7987 DVSS.n7986 2.2505
R31200 DVSS.n7988 DVSS.n4433 2.2505
R31201 DVSS.n7993 DVSS.n7989 2.2505
R31202 DVSS.n7994 DVSS.n4432 2.2505
R31203 DVSS.n7999 DVSS.n7998 2.2505
R31204 DVSS.n8000 DVSS.n4431 2.2505
R31205 DVSS.n8005 DVSS.n8001 2.2505
R31206 DVSS.n8006 DVSS.n4430 2.2505
R31207 DVSS.n8011 DVSS.n8010 2.2505
R31208 DVSS.n8012 DVSS.n4429 2.2505
R31209 DVSS.n8017 DVSS.n8013 2.2505
R31210 DVSS.n8018 DVSS.n4428 2.2505
R31211 DVSS.n8023 DVSS.n8022 2.2505
R31212 DVSS.n8024 DVSS.n4427 2.2505
R31213 DVSS.n8029 DVSS.n8025 2.2505
R31214 DVSS.n8030 DVSS.n4426 2.2505
R31215 DVSS.n8035 DVSS.n8034 2.2505
R31216 DVSS.n8036 DVSS.n4425 2.2505
R31217 DVSS.n8041 DVSS.n8037 2.2505
R31218 DVSS.n8042 DVSS.n4424 2.2505
R31219 DVSS.n8047 DVSS.n8046 2.2505
R31220 DVSS.n8048 DVSS.n4423 2.2505
R31221 DVSS.n8053 DVSS.n8049 2.2505
R31222 DVSS.n8054 DVSS.n4422 2.2505
R31223 DVSS.n8059 DVSS.n8058 2.2505
R31224 DVSS.n8060 DVSS.n4421 2.2505
R31225 DVSS.n8065 DVSS.n8061 2.2505
R31226 DVSS.n8066 DVSS.n4420 2.2505
R31227 DVSS.n8071 DVSS.n8070 2.2505
R31228 DVSS.n8072 DVSS.n4419 2.2505
R31229 DVSS.n8077 DVSS.n8073 2.2505
R31230 DVSS.n8078 DVSS.n4418 2.2505
R31231 DVSS.n8083 DVSS.n8082 2.2505
R31232 DVSS.n8084 DVSS.n4417 2.2505
R31233 DVSS.n8086 DVSS.n8085 2.2505
R31234 DVSS.n8087 DVSS.n4365 2.2505
R31235 DVSS.n8088 DVSS.n8087 2.2505
R31236 DVSS.n8086 DVSS.n4414 2.2505
R31237 DVSS.n4417 DVSS.n4416 2.2505
R31238 DVSS.n8082 DVSS.n8081 2.2505
R31239 DVSS.n8079 DVSS.n8078 2.2505
R31240 DVSS.n8077 DVSS.n8076 2.2505
R31241 DVSS.n8074 DVSS.n4419 2.2505
R31242 DVSS.n8070 DVSS.n8069 2.2505
R31243 DVSS.n8067 DVSS.n8066 2.2505
R31244 DVSS.n8065 DVSS.n8064 2.2505
R31245 DVSS.n8062 DVSS.n4421 2.2505
R31246 DVSS.n8058 DVSS.n8057 2.2505
R31247 DVSS.n8055 DVSS.n8054 2.2505
R31248 DVSS.n8053 DVSS.n8052 2.2505
R31249 DVSS.n8050 DVSS.n4423 2.2505
R31250 DVSS.n8046 DVSS.n8045 2.2505
R31251 DVSS.n8043 DVSS.n8042 2.2505
R31252 DVSS.n8041 DVSS.n8040 2.2505
R31253 DVSS.n8038 DVSS.n4425 2.2505
R31254 DVSS.n8034 DVSS.n8033 2.2505
R31255 DVSS.n8031 DVSS.n8030 2.2505
R31256 DVSS.n8029 DVSS.n8028 2.2505
R31257 DVSS.n8026 DVSS.n4427 2.2505
R31258 DVSS.n8022 DVSS.n8021 2.2505
R31259 DVSS.n8019 DVSS.n8018 2.2505
R31260 DVSS.n8017 DVSS.n8016 2.2505
R31261 DVSS.n8014 DVSS.n4429 2.2505
R31262 DVSS.n8010 DVSS.n8009 2.2505
R31263 DVSS.n8007 DVSS.n8006 2.2505
R31264 DVSS.n8005 DVSS.n8004 2.2505
R31265 DVSS.n8002 DVSS.n4431 2.2505
R31266 DVSS.n7998 DVSS.n7997 2.2505
R31267 DVSS.n7995 DVSS.n7994 2.2505
R31268 DVSS.n7993 DVSS.n7992 2.2505
R31269 DVSS.n7990 DVSS.n4433 2.2505
R31270 DVSS.n7986 DVSS.n7985 2.2505
R31271 DVSS.n7983 DVSS.n7982 2.2505
R31272 DVSS.n7981 DVSS.n7980 2.2505
R31273 DVSS.n7978 DVSS.n4435 2.2505
R31274 DVSS.n7974 DVSS.n7973 2.2505
R31275 DVSS.n7971 DVSS.n7970 2.2505
R31276 DVSS.n7969 DVSS.n7968 2.2505
R31277 DVSS.n7966 DVSS.n4437 2.2505
R31278 DVSS.n7962 DVSS.n7961 2.2505
R31279 DVSS.n7959 DVSS.n7958 2.2505
R31280 DVSS.n7957 DVSS.n7956 2.2505
R31281 DVSS.n7954 DVSS.n4439 2.2505
R31282 DVSS.n7950 DVSS.n7949 2.2505
R31283 DVSS.n7947 DVSS.n7946 2.2505
R31284 DVSS.n7945 DVSS.n7944 2.2505
R31285 DVSS.n7942 DVSS.n4441 2.2505
R31286 DVSS.n7938 DVSS.n7937 2.2505
R31287 DVSS.n7935 DVSS.n7934 2.2505
R31288 DVSS.n7933 DVSS.n7932 2.2505
R31289 DVSS.n7930 DVSS.n4443 2.2505
R31290 DVSS.n7926 DVSS.n7925 2.2505
R31291 DVSS.n7923 DVSS.n7922 2.2505
R31292 DVSS.n7921 DVSS.n7920 2.2505
R31293 DVSS.n7918 DVSS.n4445 2.2505
R31294 DVSS.n7914 DVSS.n7913 2.2505
R31295 DVSS.n7911 DVSS.n7910 2.2505
R31296 DVSS.n7909 DVSS.n7908 2.2505
R31297 DVSS.n7906 DVSS.n4447 2.2505
R31298 DVSS.n7902 DVSS.n7901 2.2505
R31299 DVSS.n7899 DVSS.n7898 2.2505
R31300 DVSS.n7897 DVSS.n7896 2.2505
R31301 DVSS.n7894 DVSS.n4449 2.2505
R31302 DVSS.n7890 DVSS.n7889 2.2505
R31303 DVSS.n7887 DVSS.n7886 2.2505
R31304 DVSS.n7885 DVSS.n7884 2.2505
R31305 DVSS.n7882 DVSS.n4451 2.2505
R31306 DVSS.n7878 DVSS.n7877 2.2505
R31307 DVSS.n7875 DVSS.n7874 2.2505
R31308 DVSS.n7873 DVSS.n7872 2.2505
R31309 DVSS.n7870 DVSS.n4453 2.2505
R31310 DVSS.n7866 DVSS.n7865 2.2505
R31311 DVSS.n7863 DVSS.n7862 2.2505
R31312 DVSS.n7861 DVSS.n7860 2.2505
R31313 DVSS.n7858 DVSS.n4455 2.2505
R31314 DVSS.n7854 DVSS.n7853 2.2505
R31315 DVSS.n7851 DVSS.n7850 2.2505
R31316 DVSS.n7849 DVSS.n7848 2.2505
R31317 DVSS.n7846 DVSS.n4457 2.2505
R31318 DVSS.n7842 DVSS.n7841 2.2505
R31319 DVSS.n4358 DVSS.n4357 2.2505
R31320 DVSS.n4026 DVSS.n4025 2.2505
R31321 DVSS.n4347 DVSS.n4027 2.2505
R31322 DVSS.n4349 DVSS.n4348 2.2505
R31323 DVSS.n4346 DVSS.n4029 2.2505
R31324 DVSS.n4345 DVSS.n4344 2.2505
R31325 DVSS.n4031 DVSS.n4030 2.2505
R31326 DVSS.n4336 DVSS.n4335 2.2505
R31327 DVSS.n4334 DVSS.n4033 2.2505
R31328 DVSS.n4333 DVSS.n4332 2.2505
R31329 DVSS.n4035 DVSS.n4034 2.2505
R31330 DVSS.n4324 DVSS.n4323 2.2505
R31331 DVSS.n4322 DVSS.n4037 2.2505
R31332 DVSS.n4321 DVSS.n4320 2.2505
R31333 DVSS.n4039 DVSS.n4038 2.2505
R31334 DVSS.n4312 DVSS.n4311 2.2505
R31335 DVSS.n4310 DVSS.n4041 2.2505
R31336 DVSS.n4309 DVSS.n4308 2.2505
R31337 DVSS.n4043 DVSS.n4042 2.2505
R31338 DVSS.n4300 DVSS.n4299 2.2505
R31339 DVSS.n4298 DVSS.n4045 2.2505
R31340 DVSS.n4297 DVSS.n4296 2.2505
R31341 DVSS.n4047 DVSS.n4046 2.2505
R31342 DVSS.n4288 DVSS.n4287 2.2505
R31343 DVSS.n4286 DVSS.n4049 2.2505
R31344 DVSS.n4285 DVSS.n4284 2.2505
R31345 DVSS.n4051 DVSS.n4050 2.2505
R31346 DVSS.n4276 DVSS.n4275 2.2505
R31347 DVSS.n4274 DVSS.n4053 2.2505
R31348 DVSS.n4273 DVSS.n4272 2.2505
R31349 DVSS.n4055 DVSS.n4054 2.2505
R31350 DVSS.n4264 DVSS.n4263 2.2505
R31351 DVSS.n4262 DVSS.n4057 2.2505
R31352 DVSS.n4261 DVSS.n4260 2.2505
R31353 DVSS.n4059 DVSS.n4058 2.2505
R31354 DVSS.n4252 DVSS.n4251 2.2505
R31355 DVSS.n4250 DVSS.n4061 2.2505
R31356 DVSS.n4249 DVSS.n4248 2.2505
R31357 DVSS.n4063 DVSS.n4062 2.2505
R31358 DVSS.n4240 DVSS.n4239 2.2505
R31359 DVSS.n4238 DVSS.n4065 2.2505
R31360 DVSS.n4237 DVSS.n4236 2.2505
R31361 DVSS.n4067 DVSS.n4066 2.2505
R31362 DVSS.n4228 DVSS.n4227 2.2505
R31363 DVSS.n4226 DVSS.n4069 2.2505
R31364 DVSS.n4225 DVSS.n4224 2.2505
R31365 DVSS.n4071 DVSS.n4070 2.2505
R31366 DVSS.n4216 DVSS.n4215 2.2505
R31367 DVSS.n4214 DVSS.n4073 2.2505
R31368 DVSS.n4213 DVSS.n4212 2.2505
R31369 DVSS.n4075 DVSS.n4074 2.2505
R31370 DVSS.n4204 DVSS.n4203 2.2505
R31371 DVSS.n4202 DVSS.n4077 2.2505
R31372 DVSS.n4201 DVSS.n4200 2.2505
R31373 DVSS.n4079 DVSS.n4078 2.2505
R31374 DVSS.n4192 DVSS.n4191 2.2505
R31375 DVSS.n4190 DVSS.n4081 2.2505
R31376 DVSS.n4189 DVSS.n4188 2.2505
R31377 DVSS.n4083 DVSS.n4082 2.2505
R31378 DVSS.n4180 DVSS.n4179 2.2505
R31379 DVSS.n4178 DVSS.n4085 2.2505
R31380 DVSS.n4177 DVSS.n4176 2.2505
R31381 DVSS.n4087 DVSS.n4086 2.2505
R31382 DVSS.n4168 DVSS.n4167 2.2505
R31383 DVSS.n4166 DVSS.n4089 2.2505
R31384 DVSS.n4165 DVSS.n4164 2.2505
R31385 DVSS.n4091 DVSS.n4090 2.2505
R31386 DVSS.n4156 DVSS.n4155 2.2505
R31387 DVSS.n4154 DVSS.n4093 2.2505
R31388 DVSS.n4153 DVSS.n4152 2.2505
R31389 DVSS.n4095 DVSS.n4094 2.2505
R31390 DVSS.n4144 DVSS.n4143 2.2505
R31391 DVSS.n4142 DVSS.n4097 2.2505
R31392 DVSS.n4141 DVSS.n4140 2.2505
R31393 DVSS.n4099 DVSS.n4098 2.2505
R31394 DVSS.n4132 DVSS.n4131 2.2505
R31395 DVSS.n4130 DVSS.n4101 2.2505
R31396 DVSS.n4129 DVSS.n4128 2.2505
R31397 DVSS.n4103 DVSS.n4102 2.2505
R31398 DVSS.n4120 DVSS.n4119 2.2505
R31399 DVSS.n4118 DVSS.n4105 2.2505
R31400 DVSS.n4117 DVSS.n4116 2.2505
R31401 DVSS.n4107 DVSS.n4106 2.2505
R31402 DVSS.n4108 DVSS.n4017 2.2505
R31403 DVSS.n4109 DVSS.n4108 2.2505
R31404 DVSS.n4111 DVSS.n4107 2.2505
R31405 DVSS.n4116 DVSS.n4115 2.2505
R31406 DVSS.n4113 DVSS.n4105 2.2505
R31407 DVSS.n4121 DVSS.n4120 2.2505
R31408 DVSS.n4123 DVSS.n4103 2.2505
R31409 DVSS.n4128 DVSS.n4127 2.2505
R31410 DVSS.n4125 DVSS.n4101 2.2505
R31411 DVSS.n4133 DVSS.n4132 2.2505
R31412 DVSS.n4135 DVSS.n4099 2.2505
R31413 DVSS.n4140 DVSS.n4139 2.2505
R31414 DVSS.n4137 DVSS.n4097 2.2505
R31415 DVSS.n4145 DVSS.n4144 2.2505
R31416 DVSS.n4147 DVSS.n4095 2.2505
R31417 DVSS.n4152 DVSS.n4151 2.2505
R31418 DVSS.n4149 DVSS.n4093 2.2505
R31419 DVSS.n4157 DVSS.n4156 2.2505
R31420 DVSS.n4159 DVSS.n4091 2.2505
R31421 DVSS.n4164 DVSS.n4163 2.2505
R31422 DVSS.n4161 DVSS.n4089 2.2505
R31423 DVSS.n4169 DVSS.n4168 2.2505
R31424 DVSS.n4171 DVSS.n4087 2.2505
R31425 DVSS.n4176 DVSS.n4175 2.2505
R31426 DVSS.n4173 DVSS.n4085 2.2505
R31427 DVSS.n4181 DVSS.n4180 2.2505
R31428 DVSS.n4183 DVSS.n4083 2.2505
R31429 DVSS.n4188 DVSS.n4187 2.2505
R31430 DVSS.n4185 DVSS.n4081 2.2505
R31431 DVSS.n4193 DVSS.n4192 2.2505
R31432 DVSS.n4195 DVSS.n4079 2.2505
R31433 DVSS.n4200 DVSS.n4199 2.2505
R31434 DVSS.n4197 DVSS.n4077 2.2505
R31435 DVSS.n4205 DVSS.n4204 2.2505
R31436 DVSS.n4207 DVSS.n4075 2.2505
R31437 DVSS.n4212 DVSS.n4211 2.2505
R31438 DVSS.n4209 DVSS.n4073 2.2505
R31439 DVSS.n4217 DVSS.n4216 2.2505
R31440 DVSS.n4219 DVSS.n4071 2.2505
R31441 DVSS.n4224 DVSS.n4223 2.2505
R31442 DVSS.n4221 DVSS.n4069 2.2505
R31443 DVSS.n4229 DVSS.n4228 2.2505
R31444 DVSS.n4231 DVSS.n4067 2.2505
R31445 DVSS.n4236 DVSS.n4235 2.2505
R31446 DVSS.n4233 DVSS.n4065 2.2505
R31447 DVSS.n4241 DVSS.n4240 2.2505
R31448 DVSS.n4243 DVSS.n4063 2.2505
R31449 DVSS.n4248 DVSS.n4247 2.2505
R31450 DVSS.n4245 DVSS.n4061 2.2505
R31451 DVSS.n4253 DVSS.n4252 2.2505
R31452 DVSS.n4255 DVSS.n4059 2.2505
R31453 DVSS.n4260 DVSS.n4259 2.2505
R31454 DVSS.n4257 DVSS.n4057 2.2505
R31455 DVSS.n4265 DVSS.n4264 2.2505
R31456 DVSS.n4267 DVSS.n4055 2.2505
R31457 DVSS.n4272 DVSS.n4271 2.2505
R31458 DVSS.n4269 DVSS.n4053 2.2505
R31459 DVSS.n4277 DVSS.n4276 2.2505
R31460 DVSS.n4279 DVSS.n4051 2.2505
R31461 DVSS.n4284 DVSS.n4283 2.2505
R31462 DVSS.n4281 DVSS.n4049 2.2505
R31463 DVSS.n4289 DVSS.n4288 2.2505
R31464 DVSS.n4291 DVSS.n4047 2.2505
R31465 DVSS.n4296 DVSS.n4295 2.2505
R31466 DVSS.n4293 DVSS.n4045 2.2505
R31467 DVSS.n4301 DVSS.n4300 2.2505
R31468 DVSS.n4303 DVSS.n4043 2.2505
R31469 DVSS.n4308 DVSS.n4307 2.2505
R31470 DVSS.n4305 DVSS.n4041 2.2505
R31471 DVSS.n4313 DVSS.n4312 2.2505
R31472 DVSS.n4315 DVSS.n4039 2.2505
R31473 DVSS.n4320 DVSS.n4319 2.2505
R31474 DVSS.n4317 DVSS.n4037 2.2505
R31475 DVSS.n4325 DVSS.n4324 2.2505
R31476 DVSS.n4327 DVSS.n4035 2.2505
R31477 DVSS.n4332 DVSS.n4331 2.2505
R31478 DVSS.n4329 DVSS.n4033 2.2505
R31479 DVSS.n4337 DVSS.n4336 2.2505
R31480 DVSS.n4339 DVSS.n4031 2.2505
R31481 DVSS.n4344 DVSS.n4343 2.2505
R31482 DVSS.n4341 DVSS.n4029 2.2505
R31483 DVSS.n4350 DVSS.n4349 2.2505
R31484 DVSS.n4352 DVSS.n4027 2.2505
R31485 DVSS.n4354 DVSS.n4026 2.2505
R31486 DVSS.n4357 DVSS.n4356 2.2505
R31487 DVSS.n8315 DVSS.n3852 2.2505
R31488 DVSS.n8314 DVSS.n8312 2.2505
R31489 DVSS.n8311 DVSS.n3948 2.2505
R31490 DVSS.n8310 DVSS.n8309 2.2505
R31491 DVSS.n8307 DVSS.n3949 2.2505
R31492 DVSS.n8305 DVSS.n8303 2.2505
R31493 DVSS.n8302 DVSS.n3951 2.2505
R31494 DVSS.n8301 DVSS.n8300 2.2505
R31495 DVSS.n8298 DVSS.n3952 2.2505
R31496 DVSS.n8296 DVSS.n8294 2.2505
R31497 DVSS.n8293 DVSS.n3954 2.2505
R31498 DVSS.n8292 DVSS.n8291 2.2505
R31499 DVSS.n8289 DVSS.n3955 2.2505
R31500 DVSS.n8287 DVSS.n8285 2.2505
R31501 DVSS.n8284 DVSS.n3957 2.2505
R31502 DVSS.n8283 DVSS.n8282 2.2505
R31503 DVSS.n8280 DVSS.n3958 2.2505
R31504 DVSS.n8278 DVSS.n8276 2.2505
R31505 DVSS.n8275 DVSS.n3960 2.2505
R31506 DVSS.n8274 DVSS.n8273 2.2505
R31507 DVSS.n8271 DVSS.n3961 2.2505
R31508 DVSS.n8269 DVSS.n8267 2.2505
R31509 DVSS.n8266 DVSS.n3963 2.2505
R31510 DVSS.n8265 DVSS.n8264 2.2505
R31511 DVSS.n8262 DVSS.n3964 2.2505
R31512 DVSS.n8260 DVSS.n8258 2.2505
R31513 DVSS.n8257 DVSS.n3966 2.2505
R31514 DVSS.n8256 DVSS.n8255 2.2505
R31515 DVSS.n8253 DVSS.n3967 2.2505
R31516 DVSS.n8251 DVSS.n8249 2.2505
R31517 DVSS.n8248 DVSS.n3969 2.2505
R31518 DVSS.n8247 DVSS.n8246 2.2505
R31519 DVSS.n8244 DVSS.n3970 2.2505
R31520 DVSS.n8242 DVSS.n8240 2.2505
R31521 DVSS.n8239 DVSS.n3972 2.2505
R31522 DVSS.n8238 DVSS.n8237 2.2505
R31523 DVSS.n8235 DVSS.n3973 2.2505
R31524 DVSS.n8233 DVSS.n8231 2.2505
R31525 DVSS.n8230 DVSS.n3975 2.2505
R31526 DVSS.n8229 DVSS.n8228 2.2505
R31527 DVSS.n8226 DVSS.n3976 2.2505
R31528 DVSS.n8224 DVSS.n8222 2.2505
R31529 DVSS.n8221 DVSS.n3978 2.2505
R31530 DVSS.n8220 DVSS.n8219 2.2505
R31531 DVSS.n8217 DVSS.n3979 2.2505
R31532 DVSS.n8215 DVSS.n8213 2.2505
R31533 DVSS.n8212 DVSS.n3981 2.2505
R31534 DVSS.n8211 DVSS.n8210 2.2505
R31535 DVSS.n8208 DVSS.n3982 2.2505
R31536 DVSS.n8206 DVSS.n8204 2.2505
R31537 DVSS.n8203 DVSS.n3984 2.2505
R31538 DVSS.n8202 DVSS.n8201 2.2505
R31539 DVSS.n8199 DVSS.n3985 2.2505
R31540 DVSS.n8197 DVSS.n8195 2.2505
R31541 DVSS.n8194 DVSS.n3987 2.2505
R31542 DVSS.n8193 DVSS.n8192 2.2505
R31543 DVSS.n8190 DVSS.n3988 2.2505
R31544 DVSS.n8188 DVSS.n8186 2.2505
R31545 DVSS.n8185 DVSS.n3990 2.2505
R31546 DVSS.n8184 DVSS.n8183 2.2505
R31547 DVSS.n8181 DVSS.n3991 2.2505
R31548 DVSS.n8179 DVSS.n8177 2.2505
R31549 DVSS.n8176 DVSS.n3993 2.2505
R31550 DVSS.n8175 DVSS.n8174 2.2505
R31551 DVSS.n8172 DVSS.n3994 2.2505
R31552 DVSS.n8170 DVSS.n8168 2.2505
R31553 DVSS.n8167 DVSS.n3996 2.2505
R31554 DVSS.n8166 DVSS.n8165 2.2505
R31555 DVSS.n8163 DVSS.n3997 2.2505
R31556 DVSS.n8161 DVSS.n8159 2.2505
R31557 DVSS.n8158 DVSS.n3999 2.2505
R31558 DVSS.n8157 DVSS.n8156 2.2505
R31559 DVSS.n8154 DVSS.n4000 2.2505
R31560 DVSS.n8152 DVSS.n8150 2.2505
R31561 DVSS.n8149 DVSS.n4002 2.2505
R31562 DVSS.n8148 DVSS.n8147 2.2505
R31563 DVSS.n8145 DVSS.n4003 2.2505
R31564 DVSS.n8143 DVSS.n8141 2.2505
R31565 DVSS.n8140 DVSS.n4005 2.2505
R31566 DVSS.n8139 DVSS.n8138 2.2505
R31567 DVSS.n8136 DVSS.n4006 2.2505
R31568 DVSS.n8134 DVSS.n8132 2.2505
R31569 DVSS.n8131 DVSS.n4007 2.2505
R31570 DVSS.n8130 DVSS.n3903 2.2505
R31571 DVSS.n8318 DVSS.n3903 2.2505
R31572 DVSS.n4007 DVSS.n3901 2.2505
R31573 DVSS.n8134 DVSS.n8133 2.2505
R31574 DVSS.n8136 DVSS.n8135 2.2505
R31575 DVSS.n8138 DVSS.n8137 2.2505
R31576 DVSS.n4005 DVSS.n4004 2.2505
R31577 DVSS.n8143 DVSS.n8142 2.2505
R31578 DVSS.n8145 DVSS.n8144 2.2505
R31579 DVSS.n8147 DVSS.n8146 2.2505
R31580 DVSS.n4002 DVSS.n4001 2.2505
R31581 DVSS.n8152 DVSS.n8151 2.2505
R31582 DVSS.n8154 DVSS.n8153 2.2505
R31583 DVSS.n8156 DVSS.n8155 2.2505
R31584 DVSS.n3999 DVSS.n3998 2.2505
R31585 DVSS.n8161 DVSS.n8160 2.2505
R31586 DVSS.n8163 DVSS.n8162 2.2505
R31587 DVSS.n8165 DVSS.n8164 2.2505
R31588 DVSS.n3996 DVSS.n3995 2.2505
R31589 DVSS.n8170 DVSS.n8169 2.2505
R31590 DVSS.n8172 DVSS.n8171 2.2505
R31591 DVSS.n8174 DVSS.n8173 2.2505
R31592 DVSS.n3993 DVSS.n3992 2.2505
R31593 DVSS.n8179 DVSS.n8178 2.2505
R31594 DVSS.n8181 DVSS.n8180 2.2505
R31595 DVSS.n8183 DVSS.n8182 2.2505
R31596 DVSS.n3990 DVSS.n3989 2.2505
R31597 DVSS.n8188 DVSS.n8187 2.2505
R31598 DVSS.n8190 DVSS.n8189 2.2505
R31599 DVSS.n8192 DVSS.n8191 2.2505
R31600 DVSS.n3987 DVSS.n3986 2.2505
R31601 DVSS.n8197 DVSS.n8196 2.2505
R31602 DVSS.n8199 DVSS.n8198 2.2505
R31603 DVSS.n8201 DVSS.n8200 2.2505
R31604 DVSS.n3984 DVSS.n3983 2.2505
R31605 DVSS.n8206 DVSS.n8205 2.2505
R31606 DVSS.n8208 DVSS.n8207 2.2505
R31607 DVSS.n8210 DVSS.n8209 2.2505
R31608 DVSS.n3981 DVSS.n3980 2.2505
R31609 DVSS.n8215 DVSS.n8214 2.2505
R31610 DVSS.n8217 DVSS.n8216 2.2505
R31611 DVSS.n8219 DVSS.n8218 2.2505
R31612 DVSS.n3978 DVSS.n3977 2.2505
R31613 DVSS.n8224 DVSS.n8223 2.2505
R31614 DVSS.n8226 DVSS.n8225 2.2505
R31615 DVSS.n8228 DVSS.n8227 2.2505
R31616 DVSS.n3975 DVSS.n3974 2.2505
R31617 DVSS.n8233 DVSS.n8232 2.2505
R31618 DVSS.n8235 DVSS.n8234 2.2505
R31619 DVSS.n8237 DVSS.n8236 2.2505
R31620 DVSS.n3972 DVSS.n3971 2.2505
R31621 DVSS.n8242 DVSS.n8241 2.2505
R31622 DVSS.n8244 DVSS.n8243 2.2505
R31623 DVSS.n8246 DVSS.n8245 2.2505
R31624 DVSS.n3969 DVSS.n3968 2.2505
R31625 DVSS.n8251 DVSS.n8250 2.2505
R31626 DVSS.n8253 DVSS.n8252 2.2505
R31627 DVSS.n8255 DVSS.n8254 2.2505
R31628 DVSS.n3966 DVSS.n3965 2.2505
R31629 DVSS.n8260 DVSS.n8259 2.2505
R31630 DVSS.n8262 DVSS.n8261 2.2505
R31631 DVSS.n8264 DVSS.n8263 2.2505
R31632 DVSS.n3963 DVSS.n3962 2.2505
R31633 DVSS.n8269 DVSS.n8268 2.2505
R31634 DVSS.n8271 DVSS.n8270 2.2505
R31635 DVSS.n8273 DVSS.n8272 2.2505
R31636 DVSS.n3960 DVSS.n3959 2.2505
R31637 DVSS.n8278 DVSS.n8277 2.2505
R31638 DVSS.n8280 DVSS.n8279 2.2505
R31639 DVSS.n8282 DVSS.n8281 2.2505
R31640 DVSS.n3957 DVSS.n3956 2.2505
R31641 DVSS.n8287 DVSS.n8286 2.2505
R31642 DVSS.n8289 DVSS.n8288 2.2505
R31643 DVSS.n8291 DVSS.n8290 2.2505
R31644 DVSS.n3954 DVSS.n3953 2.2505
R31645 DVSS.n8296 DVSS.n8295 2.2505
R31646 DVSS.n8298 DVSS.n8297 2.2505
R31647 DVSS.n8300 DVSS.n8299 2.2505
R31648 DVSS.n3951 DVSS.n3950 2.2505
R31649 DVSS.n8305 DVSS.n8304 2.2505
R31650 DVSS.n8307 DVSS.n8306 2.2505
R31651 DVSS.n8309 DVSS.n8308 2.2505
R31652 DVSS.n3948 DVSS.n3947 2.2505
R31653 DVSS.n8314 DVSS.n8313 2.2505
R31654 DVSS.n8316 DVSS.n8315 2.2505
R31655 DVSS.n8582 DVSS.n3798 2.2505
R31656 DVSS.n8584 DVSS.n8583 2.2505
R31657 DVSS.n8581 DVSS.n3800 2.2505
R31658 DVSS.n8580 DVSS.n8579 2.2505
R31659 DVSS.n8575 DVSS.n3801 2.2505
R31660 DVSS.n8571 DVSS.n8570 2.2505
R31661 DVSS.n8569 DVSS.n3802 2.2505
R31662 DVSS.n8568 DVSS.n8567 2.2505
R31663 DVSS.n8563 DVSS.n3803 2.2505
R31664 DVSS.n8559 DVSS.n8558 2.2505
R31665 DVSS.n8557 DVSS.n3804 2.2505
R31666 DVSS.n8556 DVSS.n8555 2.2505
R31667 DVSS.n8551 DVSS.n3805 2.2505
R31668 DVSS.n8547 DVSS.n8546 2.2505
R31669 DVSS.n8545 DVSS.n3806 2.2505
R31670 DVSS.n8544 DVSS.n8543 2.2505
R31671 DVSS.n8539 DVSS.n3807 2.2505
R31672 DVSS.n8535 DVSS.n8534 2.2505
R31673 DVSS.n8533 DVSS.n3808 2.2505
R31674 DVSS.n8532 DVSS.n8531 2.2505
R31675 DVSS.n8527 DVSS.n3809 2.2505
R31676 DVSS.n8523 DVSS.n8522 2.2505
R31677 DVSS.n8521 DVSS.n3810 2.2505
R31678 DVSS.n8520 DVSS.n8519 2.2505
R31679 DVSS.n8515 DVSS.n3811 2.2505
R31680 DVSS.n8511 DVSS.n8510 2.2505
R31681 DVSS.n8509 DVSS.n3812 2.2505
R31682 DVSS.n8508 DVSS.n8507 2.2505
R31683 DVSS.n8503 DVSS.n3813 2.2505
R31684 DVSS.n8499 DVSS.n8498 2.2505
R31685 DVSS.n8497 DVSS.n3814 2.2505
R31686 DVSS.n8496 DVSS.n8495 2.2505
R31687 DVSS.n8491 DVSS.n3815 2.2505
R31688 DVSS.n8487 DVSS.n8486 2.2505
R31689 DVSS.n8485 DVSS.n3816 2.2505
R31690 DVSS.n8484 DVSS.n8483 2.2505
R31691 DVSS.n8479 DVSS.n3817 2.2505
R31692 DVSS.n8475 DVSS.n8474 2.2505
R31693 DVSS.n8473 DVSS.n3818 2.2505
R31694 DVSS.n8472 DVSS.n8471 2.2505
R31695 DVSS.n8467 DVSS.n3819 2.2505
R31696 DVSS.n8463 DVSS.n8462 2.2505
R31697 DVSS.n8461 DVSS.n3820 2.2505
R31698 DVSS.n8460 DVSS.n8459 2.2505
R31699 DVSS.n8455 DVSS.n3821 2.2505
R31700 DVSS.n8451 DVSS.n8450 2.2505
R31701 DVSS.n8449 DVSS.n3822 2.2505
R31702 DVSS.n8448 DVSS.n8447 2.2505
R31703 DVSS.n8443 DVSS.n3823 2.2505
R31704 DVSS.n8439 DVSS.n8438 2.2505
R31705 DVSS.n8437 DVSS.n3824 2.2505
R31706 DVSS.n8436 DVSS.n8435 2.2505
R31707 DVSS.n8431 DVSS.n3825 2.2505
R31708 DVSS.n8427 DVSS.n8426 2.2505
R31709 DVSS.n8425 DVSS.n3826 2.2505
R31710 DVSS.n8424 DVSS.n8423 2.2505
R31711 DVSS.n8419 DVSS.n3827 2.2505
R31712 DVSS.n8415 DVSS.n8414 2.2505
R31713 DVSS.n8413 DVSS.n3828 2.2505
R31714 DVSS.n8412 DVSS.n8411 2.2505
R31715 DVSS.n8407 DVSS.n3829 2.2505
R31716 DVSS.n8403 DVSS.n8402 2.2505
R31717 DVSS.n8401 DVSS.n3830 2.2505
R31718 DVSS.n8400 DVSS.n8399 2.2505
R31719 DVSS.n8395 DVSS.n3831 2.2505
R31720 DVSS.n8391 DVSS.n8390 2.2505
R31721 DVSS.n8389 DVSS.n3832 2.2505
R31722 DVSS.n8388 DVSS.n8387 2.2505
R31723 DVSS.n8383 DVSS.n3833 2.2505
R31724 DVSS.n8379 DVSS.n8378 2.2505
R31725 DVSS.n8377 DVSS.n3834 2.2505
R31726 DVSS.n8376 DVSS.n8375 2.2505
R31727 DVSS.n8371 DVSS.n3835 2.2505
R31728 DVSS.n8367 DVSS.n8366 2.2505
R31729 DVSS.n8365 DVSS.n3836 2.2505
R31730 DVSS.n8364 DVSS.n8363 2.2505
R31731 DVSS.n8359 DVSS.n3837 2.2505
R31732 DVSS.n8355 DVSS.n8354 2.2505
R31733 DVSS.n8353 DVSS.n3838 2.2505
R31734 DVSS.n8352 DVSS.n8351 2.2505
R31735 DVSS.n8347 DVSS.n3839 2.2505
R31736 DVSS.n8343 DVSS.n8342 2.2505
R31737 DVSS.n8341 DVSS.n3842 2.2505
R31738 DVSS.n8340 DVSS.n8339 2.2505
R31739 DVSS.n8339 DVSS.n3797 2.2505
R31740 DVSS.n3842 DVSS.n3841 2.2505
R31741 DVSS.n8344 DVSS.n8343 2.2505
R31742 DVSS.n8347 DVSS.n8346 2.2505
R31743 DVSS.n8351 DVSS.n8350 2.2505
R31744 DVSS.n8348 DVSS.n3838 2.2505
R31745 DVSS.n8356 DVSS.n8355 2.2505
R31746 DVSS.n8359 DVSS.n8358 2.2505
R31747 DVSS.n8363 DVSS.n8362 2.2505
R31748 DVSS.n8360 DVSS.n3836 2.2505
R31749 DVSS.n8368 DVSS.n8367 2.2505
R31750 DVSS.n8371 DVSS.n8370 2.2505
R31751 DVSS.n8375 DVSS.n8374 2.2505
R31752 DVSS.n8372 DVSS.n3834 2.2505
R31753 DVSS.n8380 DVSS.n8379 2.2505
R31754 DVSS.n8383 DVSS.n8382 2.2505
R31755 DVSS.n8387 DVSS.n8386 2.2505
R31756 DVSS.n8384 DVSS.n3832 2.2505
R31757 DVSS.n8392 DVSS.n8391 2.2505
R31758 DVSS.n8395 DVSS.n8394 2.2505
R31759 DVSS.n8399 DVSS.n8398 2.2505
R31760 DVSS.n8396 DVSS.n3830 2.2505
R31761 DVSS.n8404 DVSS.n8403 2.2505
R31762 DVSS.n8407 DVSS.n8406 2.2505
R31763 DVSS.n8411 DVSS.n8410 2.2505
R31764 DVSS.n8408 DVSS.n3828 2.2505
R31765 DVSS.n8416 DVSS.n8415 2.2505
R31766 DVSS.n8419 DVSS.n8418 2.2505
R31767 DVSS.n8423 DVSS.n8422 2.2505
R31768 DVSS.n8420 DVSS.n3826 2.2505
R31769 DVSS.n8428 DVSS.n8427 2.2505
R31770 DVSS.n8431 DVSS.n8430 2.2505
R31771 DVSS.n8435 DVSS.n8434 2.2505
R31772 DVSS.n8432 DVSS.n3824 2.2505
R31773 DVSS.n8440 DVSS.n8439 2.2505
R31774 DVSS.n8443 DVSS.n8442 2.2505
R31775 DVSS.n8447 DVSS.n8446 2.2505
R31776 DVSS.n8444 DVSS.n3822 2.2505
R31777 DVSS.n8452 DVSS.n8451 2.2505
R31778 DVSS.n8455 DVSS.n8454 2.2505
R31779 DVSS.n8459 DVSS.n8458 2.2505
R31780 DVSS.n8456 DVSS.n3820 2.2505
R31781 DVSS.n8464 DVSS.n8463 2.2505
R31782 DVSS.n8467 DVSS.n8466 2.2505
R31783 DVSS.n8471 DVSS.n8470 2.2505
R31784 DVSS.n8468 DVSS.n3818 2.2505
R31785 DVSS.n8476 DVSS.n8475 2.2505
R31786 DVSS.n8479 DVSS.n8478 2.2505
R31787 DVSS.n8483 DVSS.n8482 2.2505
R31788 DVSS.n8480 DVSS.n3816 2.2505
R31789 DVSS.n8488 DVSS.n8487 2.2505
R31790 DVSS.n8491 DVSS.n8490 2.2505
R31791 DVSS.n8495 DVSS.n8494 2.2505
R31792 DVSS.n8492 DVSS.n3814 2.2505
R31793 DVSS.n8500 DVSS.n8499 2.2505
R31794 DVSS.n8503 DVSS.n8502 2.2505
R31795 DVSS.n8507 DVSS.n8506 2.2505
R31796 DVSS.n8504 DVSS.n3812 2.2505
R31797 DVSS.n8512 DVSS.n8511 2.2505
R31798 DVSS.n8515 DVSS.n8514 2.2505
R31799 DVSS.n8519 DVSS.n8518 2.2505
R31800 DVSS.n8516 DVSS.n3810 2.2505
R31801 DVSS.n8524 DVSS.n8523 2.2505
R31802 DVSS.n8527 DVSS.n8526 2.2505
R31803 DVSS.n8531 DVSS.n8530 2.2505
R31804 DVSS.n8528 DVSS.n3808 2.2505
R31805 DVSS.n8536 DVSS.n8535 2.2505
R31806 DVSS.n8539 DVSS.n8538 2.2505
R31807 DVSS.n8543 DVSS.n8542 2.2505
R31808 DVSS.n8540 DVSS.n3806 2.2505
R31809 DVSS.n8548 DVSS.n8547 2.2505
R31810 DVSS.n8551 DVSS.n8550 2.2505
R31811 DVSS.n8555 DVSS.n8554 2.2505
R31812 DVSS.n8552 DVSS.n3804 2.2505
R31813 DVSS.n8560 DVSS.n8559 2.2505
R31814 DVSS.n8563 DVSS.n8562 2.2505
R31815 DVSS.n8567 DVSS.n8566 2.2505
R31816 DVSS.n8564 DVSS.n3802 2.2505
R31817 DVSS.n8572 DVSS.n8571 2.2505
R31818 DVSS.n8575 DVSS.n8574 2.2505
R31819 DVSS.n8579 DVSS.n8578 2.2505
R31820 DVSS.n8576 DVSS.n3800 2.2505
R31821 DVSS.n8585 DVSS.n8584 2.2505
R31822 DVSS.n8587 DVSS.n3798 2.2505
R31823 DVSS.n8599 DVSS.n3748 2.2505
R31824 DVSS.n3747 DVSS.n3504 2.2505
R31825 DVSS.n3746 DVSS.n3745 2.2505
R31826 DVSS.n3743 DVSS.n3505 2.2505
R31827 DVSS.n3741 DVSS.n3739 2.2505
R31828 DVSS.n3738 DVSS.n3507 2.2505
R31829 DVSS.n3737 DVSS.n3736 2.2505
R31830 DVSS.n3734 DVSS.n3508 2.2505
R31831 DVSS.n3732 DVSS.n3730 2.2505
R31832 DVSS.n3729 DVSS.n3510 2.2505
R31833 DVSS.n3728 DVSS.n3727 2.2505
R31834 DVSS.n3725 DVSS.n3511 2.2505
R31835 DVSS.n3723 DVSS.n3721 2.2505
R31836 DVSS.n3720 DVSS.n3513 2.2505
R31837 DVSS.n3719 DVSS.n3718 2.2505
R31838 DVSS.n3716 DVSS.n3514 2.2505
R31839 DVSS.n3714 DVSS.n3712 2.2505
R31840 DVSS.n3711 DVSS.n3516 2.2505
R31841 DVSS.n3710 DVSS.n3709 2.2505
R31842 DVSS.n3707 DVSS.n3517 2.2505
R31843 DVSS.n3705 DVSS.n3703 2.2505
R31844 DVSS.n3702 DVSS.n3519 2.2505
R31845 DVSS.n3701 DVSS.n3700 2.2505
R31846 DVSS.n3698 DVSS.n3520 2.2505
R31847 DVSS.n3696 DVSS.n3694 2.2505
R31848 DVSS.n3693 DVSS.n3522 2.2505
R31849 DVSS.n3692 DVSS.n3691 2.2505
R31850 DVSS.n3689 DVSS.n3523 2.2505
R31851 DVSS.n3687 DVSS.n3685 2.2505
R31852 DVSS.n3684 DVSS.n3525 2.2505
R31853 DVSS.n3683 DVSS.n3682 2.2505
R31854 DVSS.n3680 DVSS.n3526 2.2505
R31855 DVSS.n3678 DVSS.n3676 2.2505
R31856 DVSS.n3675 DVSS.n3528 2.2505
R31857 DVSS.n3674 DVSS.n3673 2.2505
R31858 DVSS.n3671 DVSS.n3529 2.2505
R31859 DVSS.n3669 DVSS.n3667 2.2505
R31860 DVSS.n3666 DVSS.n3531 2.2505
R31861 DVSS.n3665 DVSS.n3664 2.2505
R31862 DVSS.n3662 DVSS.n3532 2.2505
R31863 DVSS.n3660 DVSS.n3658 2.2505
R31864 DVSS.n3657 DVSS.n3534 2.2505
R31865 DVSS.n3656 DVSS.n3655 2.2505
R31866 DVSS.n3653 DVSS.n3535 2.2505
R31867 DVSS.n3651 DVSS.n3649 2.2505
R31868 DVSS.n3648 DVSS.n3537 2.2505
R31869 DVSS.n3647 DVSS.n3646 2.2505
R31870 DVSS.n3644 DVSS.n3538 2.2505
R31871 DVSS.n3642 DVSS.n3640 2.2505
R31872 DVSS.n3639 DVSS.n3540 2.2505
R31873 DVSS.n3638 DVSS.n3637 2.2505
R31874 DVSS.n3635 DVSS.n3541 2.2505
R31875 DVSS.n3633 DVSS.n3631 2.2505
R31876 DVSS.n3630 DVSS.n3543 2.2505
R31877 DVSS.n3629 DVSS.n3628 2.2505
R31878 DVSS.n3626 DVSS.n3544 2.2505
R31879 DVSS.n3624 DVSS.n3622 2.2505
R31880 DVSS.n3621 DVSS.n3546 2.2505
R31881 DVSS.n3620 DVSS.n3619 2.2505
R31882 DVSS.n3617 DVSS.n3547 2.2505
R31883 DVSS.n3615 DVSS.n3613 2.2505
R31884 DVSS.n3612 DVSS.n3549 2.2505
R31885 DVSS.n3611 DVSS.n3610 2.2505
R31886 DVSS.n3608 DVSS.n3550 2.2505
R31887 DVSS.n3606 DVSS.n3604 2.2505
R31888 DVSS.n3603 DVSS.n3552 2.2505
R31889 DVSS.n3602 DVSS.n3601 2.2505
R31890 DVSS.n3599 DVSS.n3553 2.2505
R31891 DVSS.n3597 DVSS.n3595 2.2505
R31892 DVSS.n3594 DVSS.n3555 2.2505
R31893 DVSS.n3593 DVSS.n3592 2.2505
R31894 DVSS.n3590 DVSS.n3556 2.2505
R31895 DVSS.n3588 DVSS.n3586 2.2505
R31896 DVSS.n3585 DVSS.n3558 2.2505
R31897 DVSS.n3584 DVSS.n3583 2.2505
R31898 DVSS.n3581 DVSS.n3559 2.2505
R31899 DVSS.n3579 DVSS.n3577 2.2505
R31900 DVSS.n3576 DVSS.n3561 2.2505
R31901 DVSS.n3575 DVSS.n3574 2.2505
R31902 DVSS.n3572 DVSS.n3562 2.2505
R31903 DVSS.n3570 DVSS.n3568 2.2505
R31904 DVSS.n3567 DVSS.n3564 2.2505
R31905 DVSS.n3566 DVSS.n3565 2.2505
R31906 DVSS.n3459 DVSS.n3409 2.2505
R31907 DVSS.n8602 DVSS.n3459 2.2505
R31908 DVSS.n3565 DVSS.n3458 2.2505
R31909 DVSS.n3564 DVSS.n3563 2.2505
R31910 DVSS.n3570 DVSS.n3569 2.2505
R31911 DVSS.n3572 DVSS.n3571 2.2505
R31912 DVSS.n3574 DVSS.n3573 2.2505
R31913 DVSS.n3561 DVSS.n3560 2.2505
R31914 DVSS.n3579 DVSS.n3578 2.2505
R31915 DVSS.n3581 DVSS.n3580 2.2505
R31916 DVSS.n3583 DVSS.n3582 2.2505
R31917 DVSS.n3558 DVSS.n3557 2.2505
R31918 DVSS.n3588 DVSS.n3587 2.2505
R31919 DVSS.n3590 DVSS.n3589 2.2505
R31920 DVSS.n3592 DVSS.n3591 2.2505
R31921 DVSS.n3555 DVSS.n3554 2.2505
R31922 DVSS.n3597 DVSS.n3596 2.2505
R31923 DVSS.n3599 DVSS.n3598 2.2505
R31924 DVSS.n3601 DVSS.n3600 2.2505
R31925 DVSS.n3552 DVSS.n3551 2.2505
R31926 DVSS.n3606 DVSS.n3605 2.2505
R31927 DVSS.n3608 DVSS.n3607 2.2505
R31928 DVSS.n3610 DVSS.n3609 2.2505
R31929 DVSS.n3549 DVSS.n3548 2.2505
R31930 DVSS.n3615 DVSS.n3614 2.2505
R31931 DVSS.n3617 DVSS.n3616 2.2505
R31932 DVSS.n3619 DVSS.n3618 2.2505
R31933 DVSS.n3546 DVSS.n3545 2.2505
R31934 DVSS.n3624 DVSS.n3623 2.2505
R31935 DVSS.n3626 DVSS.n3625 2.2505
R31936 DVSS.n3628 DVSS.n3627 2.2505
R31937 DVSS.n3543 DVSS.n3542 2.2505
R31938 DVSS.n3633 DVSS.n3632 2.2505
R31939 DVSS.n3635 DVSS.n3634 2.2505
R31940 DVSS.n3637 DVSS.n3636 2.2505
R31941 DVSS.n3540 DVSS.n3539 2.2505
R31942 DVSS.n3642 DVSS.n3641 2.2505
R31943 DVSS.n3644 DVSS.n3643 2.2505
R31944 DVSS.n3646 DVSS.n3645 2.2505
R31945 DVSS.n3537 DVSS.n3536 2.2505
R31946 DVSS.n3651 DVSS.n3650 2.2505
R31947 DVSS.n3653 DVSS.n3652 2.2505
R31948 DVSS.n3655 DVSS.n3654 2.2505
R31949 DVSS.n3534 DVSS.n3533 2.2505
R31950 DVSS.n3660 DVSS.n3659 2.2505
R31951 DVSS.n3662 DVSS.n3661 2.2505
R31952 DVSS.n3664 DVSS.n3663 2.2505
R31953 DVSS.n3531 DVSS.n3530 2.2505
R31954 DVSS.n3669 DVSS.n3668 2.2505
R31955 DVSS.n3671 DVSS.n3670 2.2505
R31956 DVSS.n3673 DVSS.n3672 2.2505
R31957 DVSS.n3528 DVSS.n3527 2.2505
R31958 DVSS.n3678 DVSS.n3677 2.2505
R31959 DVSS.n3680 DVSS.n3679 2.2505
R31960 DVSS.n3682 DVSS.n3681 2.2505
R31961 DVSS.n3525 DVSS.n3524 2.2505
R31962 DVSS.n3687 DVSS.n3686 2.2505
R31963 DVSS.n3689 DVSS.n3688 2.2505
R31964 DVSS.n3691 DVSS.n3690 2.2505
R31965 DVSS.n3522 DVSS.n3521 2.2505
R31966 DVSS.n3696 DVSS.n3695 2.2505
R31967 DVSS.n3698 DVSS.n3697 2.2505
R31968 DVSS.n3700 DVSS.n3699 2.2505
R31969 DVSS.n3519 DVSS.n3518 2.2505
R31970 DVSS.n3705 DVSS.n3704 2.2505
R31971 DVSS.n3707 DVSS.n3706 2.2505
R31972 DVSS.n3709 DVSS.n3708 2.2505
R31973 DVSS.n3516 DVSS.n3515 2.2505
R31974 DVSS.n3714 DVSS.n3713 2.2505
R31975 DVSS.n3716 DVSS.n3715 2.2505
R31976 DVSS.n3718 DVSS.n3717 2.2505
R31977 DVSS.n3513 DVSS.n3512 2.2505
R31978 DVSS.n3723 DVSS.n3722 2.2505
R31979 DVSS.n3725 DVSS.n3724 2.2505
R31980 DVSS.n3727 DVSS.n3726 2.2505
R31981 DVSS.n3510 DVSS.n3509 2.2505
R31982 DVSS.n3732 DVSS.n3731 2.2505
R31983 DVSS.n3734 DVSS.n3733 2.2505
R31984 DVSS.n3736 DVSS.n3735 2.2505
R31985 DVSS.n3507 DVSS.n3506 2.2505
R31986 DVSS.n3741 DVSS.n3740 2.2505
R31987 DVSS.n3743 DVSS.n3742 2.2505
R31988 DVSS.n3745 DVSS.n3744 2.2505
R31989 DVSS.n3504 DVSS.n3503 2.2505
R31990 DVSS.n8600 DVSS.n8599 2.2505
R31991 DVSS.n3402 DVSS.n3401 2.2505
R31992 DVSS.n3070 DVSS.n3069 2.2505
R31993 DVSS.n3391 DVSS.n3071 2.2505
R31994 DVSS.n3393 DVSS.n3392 2.2505
R31995 DVSS.n3390 DVSS.n3073 2.2505
R31996 DVSS.n3389 DVSS.n3388 2.2505
R31997 DVSS.n3075 DVSS.n3074 2.2505
R31998 DVSS.n3380 DVSS.n3379 2.2505
R31999 DVSS.n3378 DVSS.n3077 2.2505
R32000 DVSS.n3377 DVSS.n3376 2.2505
R32001 DVSS.n3079 DVSS.n3078 2.2505
R32002 DVSS.n3368 DVSS.n3367 2.2505
R32003 DVSS.n3366 DVSS.n3081 2.2505
R32004 DVSS.n3365 DVSS.n3364 2.2505
R32005 DVSS.n3083 DVSS.n3082 2.2505
R32006 DVSS.n3356 DVSS.n3355 2.2505
R32007 DVSS.n3354 DVSS.n3085 2.2505
R32008 DVSS.n3353 DVSS.n3352 2.2505
R32009 DVSS.n3087 DVSS.n3086 2.2505
R32010 DVSS.n3344 DVSS.n3343 2.2505
R32011 DVSS.n3342 DVSS.n3089 2.2505
R32012 DVSS.n3341 DVSS.n3340 2.2505
R32013 DVSS.n3091 DVSS.n3090 2.2505
R32014 DVSS.n3332 DVSS.n3331 2.2505
R32015 DVSS.n3330 DVSS.n3093 2.2505
R32016 DVSS.n3329 DVSS.n3328 2.2505
R32017 DVSS.n3095 DVSS.n3094 2.2505
R32018 DVSS.n3320 DVSS.n3319 2.2505
R32019 DVSS.n3318 DVSS.n3097 2.2505
R32020 DVSS.n3317 DVSS.n3316 2.2505
R32021 DVSS.n3099 DVSS.n3098 2.2505
R32022 DVSS.n3308 DVSS.n3307 2.2505
R32023 DVSS.n3306 DVSS.n3101 2.2505
R32024 DVSS.n3305 DVSS.n3304 2.2505
R32025 DVSS.n3103 DVSS.n3102 2.2505
R32026 DVSS.n3296 DVSS.n3295 2.2505
R32027 DVSS.n3294 DVSS.n3105 2.2505
R32028 DVSS.n3293 DVSS.n3292 2.2505
R32029 DVSS.n3107 DVSS.n3106 2.2505
R32030 DVSS.n3284 DVSS.n3283 2.2505
R32031 DVSS.n3282 DVSS.n3109 2.2505
R32032 DVSS.n3281 DVSS.n3280 2.2505
R32033 DVSS.n3111 DVSS.n3110 2.2505
R32034 DVSS.n3272 DVSS.n3271 2.2505
R32035 DVSS.n3270 DVSS.n3113 2.2505
R32036 DVSS.n3269 DVSS.n3268 2.2505
R32037 DVSS.n3115 DVSS.n3114 2.2505
R32038 DVSS.n3260 DVSS.n3259 2.2505
R32039 DVSS.n3258 DVSS.n3117 2.2505
R32040 DVSS.n3257 DVSS.n3256 2.2505
R32041 DVSS.n3119 DVSS.n3118 2.2505
R32042 DVSS.n3248 DVSS.n3247 2.2505
R32043 DVSS.n3246 DVSS.n3121 2.2505
R32044 DVSS.n3245 DVSS.n3244 2.2505
R32045 DVSS.n3123 DVSS.n3122 2.2505
R32046 DVSS.n3236 DVSS.n3235 2.2505
R32047 DVSS.n3234 DVSS.n3125 2.2505
R32048 DVSS.n3233 DVSS.n3232 2.2505
R32049 DVSS.n3127 DVSS.n3126 2.2505
R32050 DVSS.n3224 DVSS.n3223 2.2505
R32051 DVSS.n3222 DVSS.n3129 2.2505
R32052 DVSS.n3221 DVSS.n3220 2.2505
R32053 DVSS.n3131 DVSS.n3130 2.2505
R32054 DVSS.n3212 DVSS.n3211 2.2505
R32055 DVSS.n3210 DVSS.n3133 2.2505
R32056 DVSS.n3209 DVSS.n3208 2.2505
R32057 DVSS.n3135 DVSS.n3134 2.2505
R32058 DVSS.n3200 DVSS.n3199 2.2505
R32059 DVSS.n3198 DVSS.n3137 2.2505
R32060 DVSS.n3197 DVSS.n3196 2.2505
R32061 DVSS.n3139 DVSS.n3138 2.2505
R32062 DVSS.n3188 DVSS.n3187 2.2505
R32063 DVSS.n3186 DVSS.n3141 2.2505
R32064 DVSS.n3185 DVSS.n3184 2.2505
R32065 DVSS.n3143 DVSS.n3142 2.2505
R32066 DVSS.n3176 DVSS.n3175 2.2505
R32067 DVSS.n3174 DVSS.n3145 2.2505
R32068 DVSS.n3173 DVSS.n3172 2.2505
R32069 DVSS.n3147 DVSS.n3146 2.2505
R32070 DVSS.n3164 DVSS.n3163 2.2505
R32071 DVSS.n3162 DVSS.n3149 2.2505
R32072 DVSS.n3161 DVSS.n3160 2.2505
R32073 DVSS.n3151 DVSS.n3150 2.2505
R32074 DVSS.n3152 DVSS.n3062 2.2505
R32075 DVSS.n3153 DVSS.n3152 2.2505
R32076 DVSS.n3155 DVSS.n3151 2.2505
R32077 DVSS.n3160 DVSS.n3159 2.2505
R32078 DVSS.n3157 DVSS.n3149 2.2505
R32079 DVSS.n3165 DVSS.n3164 2.2505
R32080 DVSS.n3167 DVSS.n3147 2.2505
R32081 DVSS.n3172 DVSS.n3171 2.2505
R32082 DVSS.n3169 DVSS.n3145 2.2505
R32083 DVSS.n3177 DVSS.n3176 2.2505
R32084 DVSS.n3179 DVSS.n3143 2.2505
R32085 DVSS.n3184 DVSS.n3183 2.2505
R32086 DVSS.n3181 DVSS.n3141 2.2505
R32087 DVSS.n3189 DVSS.n3188 2.2505
R32088 DVSS.n3191 DVSS.n3139 2.2505
R32089 DVSS.n3196 DVSS.n3195 2.2505
R32090 DVSS.n3193 DVSS.n3137 2.2505
R32091 DVSS.n3201 DVSS.n3200 2.2505
R32092 DVSS.n3203 DVSS.n3135 2.2505
R32093 DVSS.n3208 DVSS.n3207 2.2505
R32094 DVSS.n3205 DVSS.n3133 2.2505
R32095 DVSS.n3213 DVSS.n3212 2.2505
R32096 DVSS.n3215 DVSS.n3131 2.2505
R32097 DVSS.n3220 DVSS.n3219 2.2505
R32098 DVSS.n3217 DVSS.n3129 2.2505
R32099 DVSS.n3225 DVSS.n3224 2.2505
R32100 DVSS.n3227 DVSS.n3127 2.2505
R32101 DVSS.n3232 DVSS.n3231 2.2505
R32102 DVSS.n3229 DVSS.n3125 2.2505
R32103 DVSS.n3237 DVSS.n3236 2.2505
R32104 DVSS.n3239 DVSS.n3123 2.2505
R32105 DVSS.n3244 DVSS.n3243 2.2505
R32106 DVSS.n3241 DVSS.n3121 2.2505
R32107 DVSS.n3249 DVSS.n3248 2.2505
R32108 DVSS.n3251 DVSS.n3119 2.2505
R32109 DVSS.n3256 DVSS.n3255 2.2505
R32110 DVSS.n3253 DVSS.n3117 2.2505
R32111 DVSS.n3261 DVSS.n3260 2.2505
R32112 DVSS.n3263 DVSS.n3115 2.2505
R32113 DVSS.n3268 DVSS.n3267 2.2505
R32114 DVSS.n3265 DVSS.n3113 2.2505
R32115 DVSS.n3273 DVSS.n3272 2.2505
R32116 DVSS.n3275 DVSS.n3111 2.2505
R32117 DVSS.n3280 DVSS.n3279 2.2505
R32118 DVSS.n3277 DVSS.n3109 2.2505
R32119 DVSS.n3285 DVSS.n3284 2.2505
R32120 DVSS.n3287 DVSS.n3107 2.2505
R32121 DVSS.n3292 DVSS.n3291 2.2505
R32122 DVSS.n3289 DVSS.n3105 2.2505
R32123 DVSS.n3297 DVSS.n3296 2.2505
R32124 DVSS.n3299 DVSS.n3103 2.2505
R32125 DVSS.n3304 DVSS.n3303 2.2505
R32126 DVSS.n3301 DVSS.n3101 2.2505
R32127 DVSS.n3309 DVSS.n3308 2.2505
R32128 DVSS.n3311 DVSS.n3099 2.2505
R32129 DVSS.n3316 DVSS.n3315 2.2505
R32130 DVSS.n3313 DVSS.n3097 2.2505
R32131 DVSS.n3321 DVSS.n3320 2.2505
R32132 DVSS.n3323 DVSS.n3095 2.2505
R32133 DVSS.n3328 DVSS.n3327 2.2505
R32134 DVSS.n3325 DVSS.n3093 2.2505
R32135 DVSS.n3333 DVSS.n3332 2.2505
R32136 DVSS.n3335 DVSS.n3091 2.2505
R32137 DVSS.n3340 DVSS.n3339 2.2505
R32138 DVSS.n3337 DVSS.n3089 2.2505
R32139 DVSS.n3345 DVSS.n3344 2.2505
R32140 DVSS.n3347 DVSS.n3087 2.2505
R32141 DVSS.n3352 DVSS.n3351 2.2505
R32142 DVSS.n3349 DVSS.n3085 2.2505
R32143 DVSS.n3357 DVSS.n3356 2.2505
R32144 DVSS.n3359 DVSS.n3083 2.2505
R32145 DVSS.n3364 DVSS.n3363 2.2505
R32146 DVSS.n3361 DVSS.n3081 2.2505
R32147 DVSS.n3369 DVSS.n3368 2.2505
R32148 DVSS.n3371 DVSS.n3079 2.2505
R32149 DVSS.n3376 DVSS.n3375 2.2505
R32150 DVSS.n3373 DVSS.n3077 2.2505
R32151 DVSS.n3381 DVSS.n3380 2.2505
R32152 DVSS.n3383 DVSS.n3075 2.2505
R32153 DVSS.n3388 DVSS.n3387 2.2505
R32154 DVSS.n3385 DVSS.n3073 2.2505
R32155 DVSS.n3394 DVSS.n3393 2.2505
R32156 DVSS.n3396 DVSS.n3071 2.2505
R32157 DVSS.n3398 DVSS.n3070 2.2505
R32158 DVSS.n3401 DVSS.n3400 2.2505
R32159 DVSS.n8721 DVSS.n3055 2.2505
R32160 DVSS.n8723 DVSS.n8722 2.2505
R32161 DVSS.n8728 DVSS.n8724 2.2505
R32162 DVSS.n8729 DVSS.n8719 2.2505
R32163 DVSS.n8734 DVSS.n8733 2.2505
R32164 DVSS.n8735 DVSS.n8718 2.2505
R32165 DVSS.n8740 DVSS.n8736 2.2505
R32166 DVSS.n8741 DVSS.n8717 2.2505
R32167 DVSS.n8746 DVSS.n8745 2.2505
R32168 DVSS.n8747 DVSS.n8716 2.2505
R32169 DVSS.n8752 DVSS.n8748 2.2505
R32170 DVSS.n8753 DVSS.n8715 2.2505
R32171 DVSS.n8758 DVSS.n8757 2.2505
R32172 DVSS.n8759 DVSS.n8714 2.2505
R32173 DVSS.n8764 DVSS.n8760 2.2505
R32174 DVSS.n8765 DVSS.n8713 2.2505
R32175 DVSS.n8770 DVSS.n8769 2.2505
R32176 DVSS.n8771 DVSS.n8712 2.2505
R32177 DVSS.n8776 DVSS.n8772 2.2505
R32178 DVSS.n8777 DVSS.n8711 2.2505
R32179 DVSS.n8782 DVSS.n8781 2.2505
R32180 DVSS.n8783 DVSS.n8710 2.2505
R32181 DVSS.n8788 DVSS.n8784 2.2505
R32182 DVSS.n8789 DVSS.n8709 2.2505
R32183 DVSS.n8794 DVSS.n8793 2.2505
R32184 DVSS.n8795 DVSS.n8708 2.2505
R32185 DVSS.n8800 DVSS.n8796 2.2505
R32186 DVSS.n8801 DVSS.n8707 2.2505
R32187 DVSS.n8806 DVSS.n8805 2.2505
R32188 DVSS.n8807 DVSS.n8706 2.2505
R32189 DVSS.n8812 DVSS.n8808 2.2505
R32190 DVSS.n8813 DVSS.n8705 2.2505
R32191 DVSS.n8818 DVSS.n8817 2.2505
R32192 DVSS.n8819 DVSS.n8704 2.2505
R32193 DVSS.n8824 DVSS.n8820 2.2505
R32194 DVSS.n8825 DVSS.n8703 2.2505
R32195 DVSS.n8830 DVSS.n8829 2.2505
R32196 DVSS.n8831 DVSS.n8702 2.2505
R32197 DVSS.n8836 DVSS.n8832 2.2505
R32198 DVSS.n8837 DVSS.n8701 2.2505
R32199 DVSS.n8842 DVSS.n8841 2.2505
R32200 DVSS.n8843 DVSS.n8700 2.2505
R32201 DVSS.n8848 DVSS.n8844 2.2505
R32202 DVSS.n8849 DVSS.n8699 2.2505
R32203 DVSS.n8854 DVSS.n8853 2.2505
R32204 DVSS.n8855 DVSS.n8698 2.2505
R32205 DVSS.n8860 DVSS.n8856 2.2505
R32206 DVSS.n8861 DVSS.n8697 2.2505
R32207 DVSS.n8866 DVSS.n8865 2.2505
R32208 DVSS.n8867 DVSS.n8696 2.2505
R32209 DVSS.n8872 DVSS.n8868 2.2505
R32210 DVSS.n8873 DVSS.n8695 2.2505
R32211 DVSS.n8878 DVSS.n8877 2.2505
R32212 DVSS.n8879 DVSS.n8694 2.2505
R32213 DVSS.n8884 DVSS.n8880 2.2505
R32214 DVSS.n8885 DVSS.n8693 2.2505
R32215 DVSS.n8890 DVSS.n8889 2.2505
R32216 DVSS.n8891 DVSS.n8692 2.2505
R32217 DVSS.n8896 DVSS.n8892 2.2505
R32218 DVSS.n8897 DVSS.n8691 2.2505
R32219 DVSS.n8902 DVSS.n8901 2.2505
R32220 DVSS.n8903 DVSS.n8690 2.2505
R32221 DVSS.n8908 DVSS.n8904 2.2505
R32222 DVSS.n8909 DVSS.n8689 2.2505
R32223 DVSS.n8914 DVSS.n8913 2.2505
R32224 DVSS.n8915 DVSS.n8688 2.2505
R32225 DVSS.n8920 DVSS.n8916 2.2505
R32226 DVSS.n8921 DVSS.n8687 2.2505
R32227 DVSS.n8926 DVSS.n8925 2.2505
R32228 DVSS.n8927 DVSS.n8686 2.2505
R32229 DVSS.n8932 DVSS.n8928 2.2505
R32230 DVSS.n8933 DVSS.n8685 2.2505
R32231 DVSS.n8938 DVSS.n8937 2.2505
R32232 DVSS.n8939 DVSS.n8684 2.2505
R32233 DVSS.n8944 DVSS.n8940 2.2505
R32234 DVSS.n8945 DVSS.n8683 2.2505
R32235 DVSS.n8950 DVSS.n8949 2.2505
R32236 DVSS.n8951 DVSS.n8682 2.2505
R32237 DVSS.n8956 DVSS.n8952 2.2505
R32238 DVSS.n8957 DVSS.n8681 2.2505
R32239 DVSS.n8962 DVSS.n8961 2.2505
R32240 DVSS.n8963 DVSS.n8680 2.2505
R32241 DVSS.n8965 DVSS.n8964 2.2505
R32242 DVSS.n8966 DVSS.n3048 2.2505
R32243 DVSS.n8967 DVSS.n8966 2.2505
R32244 DVSS.n8965 DVSS.n8677 2.2505
R32245 DVSS.n8680 DVSS.n8679 2.2505
R32246 DVSS.n8961 DVSS.n8960 2.2505
R32247 DVSS.n8958 DVSS.n8957 2.2505
R32248 DVSS.n8956 DVSS.n8955 2.2505
R32249 DVSS.n8953 DVSS.n8682 2.2505
R32250 DVSS.n8949 DVSS.n8948 2.2505
R32251 DVSS.n8946 DVSS.n8945 2.2505
R32252 DVSS.n8944 DVSS.n8943 2.2505
R32253 DVSS.n8941 DVSS.n8684 2.2505
R32254 DVSS.n8937 DVSS.n8936 2.2505
R32255 DVSS.n8934 DVSS.n8933 2.2505
R32256 DVSS.n8932 DVSS.n8931 2.2505
R32257 DVSS.n8929 DVSS.n8686 2.2505
R32258 DVSS.n8925 DVSS.n8924 2.2505
R32259 DVSS.n8922 DVSS.n8921 2.2505
R32260 DVSS.n8920 DVSS.n8919 2.2505
R32261 DVSS.n8917 DVSS.n8688 2.2505
R32262 DVSS.n8913 DVSS.n8912 2.2505
R32263 DVSS.n8910 DVSS.n8909 2.2505
R32264 DVSS.n8908 DVSS.n8907 2.2505
R32265 DVSS.n8905 DVSS.n8690 2.2505
R32266 DVSS.n8901 DVSS.n8900 2.2505
R32267 DVSS.n8898 DVSS.n8897 2.2505
R32268 DVSS.n8896 DVSS.n8895 2.2505
R32269 DVSS.n8893 DVSS.n8692 2.2505
R32270 DVSS.n8889 DVSS.n8888 2.2505
R32271 DVSS.n8886 DVSS.n8885 2.2505
R32272 DVSS.n8884 DVSS.n8883 2.2505
R32273 DVSS.n8881 DVSS.n8694 2.2505
R32274 DVSS.n8877 DVSS.n8876 2.2505
R32275 DVSS.n8874 DVSS.n8873 2.2505
R32276 DVSS.n8872 DVSS.n8871 2.2505
R32277 DVSS.n8869 DVSS.n8696 2.2505
R32278 DVSS.n8865 DVSS.n8864 2.2505
R32279 DVSS.n8862 DVSS.n8861 2.2505
R32280 DVSS.n8860 DVSS.n8859 2.2505
R32281 DVSS.n8857 DVSS.n8698 2.2505
R32282 DVSS.n8853 DVSS.n8852 2.2505
R32283 DVSS.n8850 DVSS.n8849 2.2505
R32284 DVSS.n8848 DVSS.n8847 2.2505
R32285 DVSS.n8845 DVSS.n8700 2.2505
R32286 DVSS.n8841 DVSS.n8840 2.2505
R32287 DVSS.n8838 DVSS.n8837 2.2505
R32288 DVSS.n8836 DVSS.n8835 2.2505
R32289 DVSS.n8833 DVSS.n8702 2.2505
R32290 DVSS.n8829 DVSS.n8828 2.2505
R32291 DVSS.n8826 DVSS.n8825 2.2505
R32292 DVSS.n8824 DVSS.n8823 2.2505
R32293 DVSS.n8821 DVSS.n8704 2.2505
R32294 DVSS.n8817 DVSS.n8816 2.2505
R32295 DVSS.n8814 DVSS.n8813 2.2505
R32296 DVSS.n8812 DVSS.n8811 2.2505
R32297 DVSS.n8809 DVSS.n8706 2.2505
R32298 DVSS.n8805 DVSS.n8804 2.2505
R32299 DVSS.n8802 DVSS.n8801 2.2505
R32300 DVSS.n8800 DVSS.n8799 2.2505
R32301 DVSS.n8797 DVSS.n8708 2.2505
R32302 DVSS.n8793 DVSS.n8792 2.2505
R32303 DVSS.n8790 DVSS.n8789 2.2505
R32304 DVSS.n8788 DVSS.n8787 2.2505
R32305 DVSS.n8785 DVSS.n8710 2.2505
R32306 DVSS.n8781 DVSS.n8780 2.2505
R32307 DVSS.n8778 DVSS.n8777 2.2505
R32308 DVSS.n8776 DVSS.n8775 2.2505
R32309 DVSS.n8773 DVSS.n8712 2.2505
R32310 DVSS.n8769 DVSS.n8768 2.2505
R32311 DVSS.n8766 DVSS.n8765 2.2505
R32312 DVSS.n8764 DVSS.n8763 2.2505
R32313 DVSS.n8761 DVSS.n8714 2.2505
R32314 DVSS.n8757 DVSS.n8756 2.2505
R32315 DVSS.n8754 DVSS.n8753 2.2505
R32316 DVSS.n8752 DVSS.n8751 2.2505
R32317 DVSS.n8749 DVSS.n8716 2.2505
R32318 DVSS.n8745 DVSS.n8744 2.2505
R32319 DVSS.n8742 DVSS.n8741 2.2505
R32320 DVSS.n8740 DVSS.n8739 2.2505
R32321 DVSS.n8737 DVSS.n8718 2.2505
R32322 DVSS.n8733 DVSS.n8732 2.2505
R32323 DVSS.n8730 DVSS.n8729 2.2505
R32324 DVSS.n8728 DVSS.n8727 2.2505
R32325 DVSS.n8725 DVSS.n8722 2.2505
R32326 DVSS.n8721 DVSS.n8720 2.2505
R32327 DVSS.n9182 DVSS.n2884 2.2505
R32328 DVSS.n9181 DVSS.n9179 2.2505
R32329 DVSS.n9178 DVSS.n2980 2.2505
R32330 DVSS.n9177 DVSS.n9176 2.2505
R32331 DVSS.n9174 DVSS.n2981 2.2505
R32332 DVSS.n9172 DVSS.n9170 2.2505
R32333 DVSS.n9169 DVSS.n2983 2.2505
R32334 DVSS.n9168 DVSS.n9167 2.2505
R32335 DVSS.n9165 DVSS.n2984 2.2505
R32336 DVSS.n9163 DVSS.n9161 2.2505
R32337 DVSS.n9160 DVSS.n2986 2.2505
R32338 DVSS.n9159 DVSS.n9158 2.2505
R32339 DVSS.n9156 DVSS.n2987 2.2505
R32340 DVSS.n9154 DVSS.n9152 2.2505
R32341 DVSS.n9151 DVSS.n2989 2.2505
R32342 DVSS.n9150 DVSS.n9149 2.2505
R32343 DVSS.n9147 DVSS.n2990 2.2505
R32344 DVSS.n9145 DVSS.n9143 2.2505
R32345 DVSS.n9142 DVSS.n2992 2.2505
R32346 DVSS.n9141 DVSS.n9140 2.2505
R32347 DVSS.n9138 DVSS.n2993 2.2505
R32348 DVSS.n9136 DVSS.n9134 2.2505
R32349 DVSS.n9133 DVSS.n2995 2.2505
R32350 DVSS.n9132 DVSS.n9131 2.2505
R32351 DVSS.n9129 DVSS.n2996 2.2505
R32352 DVSS.n9127 DVSS.n9125 2.2505
R32353 DVSS.n9124 DVSS.n2998 2.2505
R32354 DVSS.n9123 DVSS.n9122 2.2505
R32355 DVSS.n9120 DVSS.n2999 2.2505
R32356 DVSS.n9118 DVSS.n9116 2.2505
R32357 DVSS.n9115 DVSS.n3001 2.2505
R32358 DVSS.n9114 DVSS.n9113 2.2505
R32359 DVSS.n9111 DVSS.n3002 2.2505
R32360 DVSS.n9109 DVSS.n9107 2.2505
R32361 DVSS.n9106 DVSS.n3004 2.2505
R32362 DVSS.n9105 DVSS.n9104 2.2505
R32363 DVSS.n9102 DVSS.n3005 2.2505
R32364 DVSS.n9100 DVSS.n9098 2.2505
R32365 DVSS.n9097 DVSS.n3007 2.2505
R32366 DVSS.n9096 DVSS.n9095 2.2505
R32367 DVSS.n9093 DVSS.n3008 2.2505
R32368 DVSS.n9091 DVSS.n9089 2.2505
R32369 DVSS.n9088 DVSS.n3010 2.2505
R32370 DVSS.n9087 DVSS.n9086 2.2505
R32371 DVSS.n9084 DVSS.n3011 2.2505
R32372 DVSS.n9082 DVSS.n9080 2.2505
R32373 DVSS.n9079 DVSS.n3013 2.2505
R32374 DVSS.n9078 DVSS.n9077 2.2505
R32375 DVSS.n9075 DVSS.n3014 2.2505
R32376 DVSS.n9073 DVSS.n9071 2.2505
R32377 DVSS.n9070 DVSS.n3016 2.2505
R32378 DVSS.n9069 DVSS.n9068 2.2505
R32379 DVSS.n9066 DVSS.n3017 2.2505
R32380 DVSS.n9064 DVSS.n9062 2.2505
R32381 DVSS.n9061 DVSS.n3019 2.2505
R32382 DVSS.n9060 DVSS.n9059 2.2505
R32383 DVSS.n9057 DVSS.n3020 2.2505
R32384 DVSS.n9055 DVSS.n9053 2.2505
R32385 DVSS.n9052 DVSS.n3022 2.2505
R32386 DVSS.n9051 DVSS.n9050 2.2505
R32387 DVSS.n9048 DVSS.n3023 2.2505
R32388 DVSS.n9046 DVSS.n9044 2.2505
R32389 DVSS.n9043 DVSS.n3025 2.2505
R32390 DVSS.n9042 DVSS.n9041 2.2505
R32391 DVSS.n9039 DVSS.n3026 2.2505
R32392 DVSS.n9037 DVSS.n9035 2.2505
R32393 DVSS.n9034 DVSS.n3028 2.2505
R32394 DVSS.n9033 DVSS.n9032 2.2505
R32395 DVSS.n9030 DVSS.n3029 2.2505
R32396 DVSS.n9028 DVSS.n9026 2.2505
R32397 DVSS.n9025 DVSS.n3031 2.2505
R32398 DVSS.n9024 DVSS.n9023 2.2505
R32399 DVSS.n9021 DVSS.n3032 2.2505
R32400 DVSS.n9019 DVSS.n9017 2.2505
R32401 DVSS.n9016 DVSS.n3034 2.2505
R32402 DVSS.n9015 DVSS.n9014 2.2505
R32403 DVSS.n9012 DVSS.n3035 2.2505
R32404 DVSS.n9010 DVSS.n9008 2.2505
R32405 DVSS.n9007 DVSS.n3037 2.2505
R32406 DVSS.n9006 DVSS.n9005 2.2505
R32407 DVSS.n9003 DVSS.n3038 2.2505
R32408 DVSS.n9001 DVSS.n8999 2.2505
R32409 DVSS.n8998 DVSS.n3039 2.2505
R32410 DVSS.n8997 DVSS.n2935 2.2505
R32411 DVSS.n9185 DVSS.n2935 2.2505
R32412 DVSS.n3039 DVSS.n2933 2.2505
R32413 DVSS.n9001 DVSS.n9000 2.2505
R32414 DVSS.n9003 DVSS.n9002 2.2505
R32415 DVSS.n9005 DVSS.n9004 2.2505
R32416 DVSS.n3037 DVSS.n3036 2.2505
R32417 DVSS.n9010 DVSS.n9009 2.2505
R32418 DVSS.n9012 DVSS.n9011 2.2505
R32419 DVSS.n9014 DVSS.n9013 2.2505
R32420 DVSS.n3034 DVSS.n3033 2.2505
R32421 DVSS.n9019 DVSS.n9018 2.2505
R32422 DVSS.n9021 DVSS.n9020 2.2505
R32423 DVSS.n9023 DVSS.n9022 2.2505
R32424 DVSS.n3031 DVSS.n3030 2.2505
R32425 DVSS.n9028 DVSS.n9027 2.2505
R32426 DVSS.n9030 DVSS.n9029 2.2505
R32427 DVSS.n9032 DVSS.n9031 2.2505
R32428 DVSS.n3028 DVSS.n3027 2.2505
R32429 DVSS.n9037 DVSS.n9036 2.2505
R32430 DVSS.n9039 DVSS.n9038 2.2505
R32431 DVSS.n9041 DVSS.n9040 2.2505
R32432 DVSS.n3025 DVSS.n3024 2.2505
R32433 DVSS.n9046 DVSS.n9045 2.2505
R32434 DVSS.n9048 DVSS.n9047 2.2505
R32435 DVSS.n9050 DVSS.n9049 2.2505
R32436 DVSS.n3022 DVSS.n3021 2.2505
R32437 DVSS.n9055 DVSS.n9054 2.2505
R32438 DVSS.n9057 DVSS.n9056 2.2505
R32439 DVSS.n9059 DVSS.n9058 2.2505
R32440 DVSS.n3019 DVSS.n3018 2.2505
R32441 DVSS.n9064 DVSS.n9063 2.2505
R32442 DVSS.n9066 DVSS.n9065 2.2505
R32443 DVSS.n9068 DVSS.n9067 2.2505
R32444 DVSS.n3016 DVSS.n3015 2.2505
R32445 DVSS.n9073 DVSS.n9072 2.2505
R32446 DVSS.n9075 DVSS.n9074 2.2505
R32447 DVSS.n9077 DVSS.n9076 2.2505
R32448 DVSS.n3013 DVSS.n3012 2.2505
R32449 DVSS.n9082 DVSS.n9081 2.2505
R32450 DVSS.n9084 DVSS.n9083 2.2505
R32451 DVSS.n9086 DVSS.n9085 2.2505
R32452 DVSS.n3010 DVSS.n3009 2.2505
R32453 DVSS.n9091 DVSS.n9090 2.2505
R32454 DVSS.n9093 DVSS.n9092 2.2505
R32455 DVSS.n9095 DVSS.n9094 2.2505
R32456 DVSS.n3007 DVSS.n3006 2.2505
R32457 DVSS.n9100 DVSS.n9099 2.2505
R32458 DVSS.n9102 DVSS.n9101 2.2505
R32459 DVSS.n9104 DVSS.n9103 2.2505
R32460 DVSS.n3004 DVSS.n3003 2.2505
R32461 DVSS.n9109 DVSS.n9108 2.2505
R32462 DVSS.n9111 DVSS.n9110 2.2505
R32463 DVSS.n9113 DVSS.n9112 2.2505
R32464 DVSS.n3001 DVSS.n3000 2.2505
R32465 DVSS.n9118 DVSS.n9117 2.2505
R32466 DVSS.n9120 DVSS.n9119 2.2505
R32467 DVSS.n9122 DVSS.n9121 2.2505
R32468 DVSS.n2998 DVSS.n2997 2.2505
R32469 DVSS.n9127 DVSS.n9126 2.2505
R32470 DVSS.n9129 DVSS.n9128 2.2505
R32471 DVSS.n9131 DVSS.n9130 2.2505
R32472 DVSS.n2995 DVSS.n2994 2.2505
R32473 DVSS.n9136 DVSS.n9135 2.2505
R32474 DVSS.n9138 DVSS.n9137 2.2505
R32475 DVSS.n9140 DVSS.n9139 2.2505
R32476 DVSS.n2992 DVSS.n2991 2.2505
R32477 DVSS.n9145 DVSS.n9144 2.2505
R32478 DVSS.n9147 DVSS.n9146 2.2505
R32479 DVSS.n9149 DVSS.n9148 2.2505
R32480 DVSS.n2989 DVSS.n2988 2.2505
R32481 DVSS.n9154 DVSS.n9153 2.2505
R32482 DVSS.n9156 DVSS.n9155 2.2505
R32483 DVSS.n9158 DVSS.n9157 2.2505
R32484 DVSS.n2986 DVSS.n2985 2.2505
R32485 DVSS.n9163 DVSS.n9162 2.2505
R32486 DVSS.n9165 DVSS.n9164 2.2505
R32487 DVSS.n9167 DVSS.n9166 2.2505
R32488 DVSS.n2983 DVSS.n2982 2.2505
R32489 DVSS.n9172 DVSS.n9171 2.2505
R32490 DVSS.n9174 DVSS.n9173 2.2505
R32491 DVSS.n9176 DVSS.n9175 2.2505
R32492 DVSS.n2980 DVSS.n2979 2.2505
R32493 DVSS.n9181 DVSS.n9180 2.2505
R32494 DVSS.n9183 DVSS.n9182 2.2505
R32495 DVSS.n9449 DVSS.n2830 2.2505
R32496 DVSS.n9451 DVSS.n9450 2.2505
R32497 DVSS.n9448 DVSS.n2832 2.2505
R32498 DVSS.n9447 DVSS.n9446 2.2505
R32499 DVSS.n9442 DVSS.n2833 2.2505
R32500 DVSS.n9438 DVSS.n9437 2.2505
R32501 DVSS.n9436 DVSS.n2834 2.2505
R32502 DVSS.n9435 DVSS.n9434 2.2505
R32503 DVSS.n9430 DVSS.n2835 2.2505
R32504 DVSS.n9426 DVSS.n9425 2.2505
R32505 DVSS.n9424 DVSS.n2836 2.2505
R32506 DVSS.n9423 DVSS.n9422 2.2505
R32507 DVSS.n9418 DVSS.n2837 2.2505
R32508 DVSS.n9414 DVSS.n9413 2.2505
R32509 DVSS.n9412 DVSS.n2838 2.2505
R32510 DVSS.n9411 DVSS.n9410 2.2505
R32511 DVSS.n9406 DVSS.n2839 2.2505
R32512 DVSS.n9402 DVSS.n9401 2.2505
R32513 DVSS.n9400 DVSS.n2840 2.2505
R32514 DVSS.n9399 DVSS.n9398 2.2505
R32515 DVSS.n9394 DVSS.n2841 2.2505
R32516 DVSS.n9390 DVSS.n9389 2.2505
R32517 DVSS.n9388 DVSS.n2842 2.2505
R32518 DVSS.n9387 DVSS.n9386 2.2505
R32519 DVSS.n9382 DVSS.n2843 2.2505
R32520 DVSS.n9378 DVSS.n9377 2.2505
R32521 DVSS.n9376 DVSS.n2844 2.2505
R32522 DVSS.n9375 DVSS.n9374 2.2505
R32523 DVSS.n9370 DVSS.n2845 2.2505
R32524 DVSS.n9366 DVSS.n9365 2.2505
R32525 DVSS.n9364 DVSS.n2846 2.2505
R32526 DVSS.n9363 DVSS.n9362 2.2505
R32527 DVSS.n9358 DVSS.n2847 2.2505
R32528 DVSS.n9354 DVSS.n9353 2.2505
R32529 DVSS.n9352 DVSS.n2848 2.2505
R32530 DVSS.n9351 DVSS.n9350 2.2505
R32531 DVSS.n9346 DVSS.n2849 2.2505
R32532 DVSS.n9342 DVSS.n9341 2.2505
R32533 DVSS.n9340 DVSS.n2850 2.2505
R32534 DVSS.n9339 DVSS.n9338 2.2505
R32535 DVSS.n9334 DVSS.n2851 2.2505
R32536 DVSS.n9330 DVSS.n9329 2.2505
R32537 DVSS.n9328 DVSS.n2852 2.2505
R32538 DVSS.n9327 DVSS.n9326 2.2505
R32539 DVSS.n9322 DVSS.n2853 2.2505
R32540 DVSS.n9318 DVSS.n9317 2.2505
R32541 DVSS.n9316 DVSS.n2854 2.2505
R32542 DVSS.n9315 DVSS.n9314 2.2505
R32543 DVSS.n9310 DVSS.n2855 2.2505
R32544 DVSS.n9306 DVSS.n9305 2.2505
R32545 DVSS.n9304 DVSS.n2856 2.2505
R32546 DVSS.n9303 DVSS.n9302 2.2505
R32547 DVSS.n9298 DVSS.n2857 2.2505
R32548 DVSS.n9294 DVSS.n9293 2.2505
R32549 DVSS.n9292 DVSS.n2858 2.2505
R32550 DVSS.n9291 DVSS.n9290 2.2505
R32551 DVSS.n9286 DVSS.n2859 2.2505
R32552 DVSS.n9282 DVSS.n9281 2.2505
R32553 DVSS.n9280 DVSS.n2860 2.2505
R32554 DVSS.n9279 DVSS.n9278 2.2505
R32555 DVSS.n9274 DVSS.n2861 2.2505
R32556 DVSS.n9270 DVSS.n9269 2.2505
R32557 DVSS.n9268 DVSS.n2862 2.2505
R32558 DVSS.n9267 DVSS.n9266 2.2505
R32559 DVSS.n9262 DVSS.n2863 2.2505
R32560 DVSS.n9258 DVSS.n9257 2.2505
R32561 DVSS.n9256 DVSS.n2864 2.2505
R32562 DVSS.n9255 DVSS.n9254 2.2505
R32563 DVSS.n9250 DVSS.n2865 2.2505
R32564 DVSS.n9246 DVSS.n9245 2.2505
R32565 DVSS.n9244 DVSS.n2866 2.2505
R32566 DVSS.n9243 DVSS.n9242 2.2505
R32567 DVSS.n9238 DVSS.n2867 2.2505
R32568 DVSS.n9234 DVSS.n9233 2.2505
R32569 DVSS.n9232 DVSS.n2868 2.2505
R32570 DVSS.n9231 DVSS.n9230 2.2505
R32571 DVSS.n9226 DVSS.n2869 2.2505
R32572 DVSS.n9222 DVSS.n9221 2.2505
R32573 DVSS.n9220 DVSS.n2870 2.2505
R32574 DVSS.n9219 DVSS.n9218 2.2505
R32575 DVSS.n9214 DVSS.n2871 2.2505
R32576 DVSS.n9210 DVSS.n9209 2.2505
R32577 DVSS.n9208 DVSS.n2874 2.2505
R32578 DVSS.n9207 DVSS.n9206 2.2505
R32579 DVSS.n9206 DVSS.n2829 2.2505
R32580 DVSS.n2874 DVSS.n2873 2.2505
R32581 DVSS.n9211 DVSS.n9210 2.2505
R32582 DVSS.n9214 DVSS.n9213 2.2505
R32583 DVSS.n9218 DVSS.n9217 2.2505
R32584 DVSS.n9215 DVSS.n2870 2.2505
R32585 DVSS.n9223 DVSS.n9222 2.2505
R32586 DVSS.n9226 DVSS.n9225 2.2505
R32587 DVSS.n9230 DVSS.n9229 2.2505
R32588 DVSS.n9227 DVSS.n2868 2.2505
R32589 DVSS.n9235 DVSS.n9234 2.2505
R32590 DVSS.n9238 DVSS.n9237 2.2505
R32591 DVSS.n9242 DVSS.n9241 2.2505
R32592 DVSS.n9239 DVSS.n2866 2.2505
R32593 DVSS.n9247 DVSS.n9246 2.2505
R32594 DVSS.n9250 DVSS.n9249 2.2505
R32595 DVSS.n9254 DVSS.n9253 2.2505
R32596 DVSS.n9251 DVSS.n2864 2.2505
R32597 DVSS.n9259 DVSS.n9258 2.2505
R32598 DVSS.n9262 DVSS.n9261 2.2505
R32599 DVSS.n9266 DVSS.n9265 2.2505
R32600 DVSS.n9263 DVSS.n2862 2.2505
R32601 DVSS.n9271 DVSS.n9270 2.2505
R32602 DVSS.n9274 DVSS.n9273 2.2505
R32603 DVSS.n9278 DVSS.n9277 2.2505
R32604 DVSS.n9275 DVSS.n2860 2.2505
R32605 DVSS.n9283 DVSS.n9282 2.2505
R32606 DVSS.n9286 DVSS.n9285 2.2505
R32607 DVSS.n9290 DVSS.n9289 2.2505
R32608 DVSS.n9287 DVSS.n2858 2.2505
R32609 DVSS.n9295 DVSS.n9294 2.2505
R32610 DVSS.n9298 DVSS.n9297 2.2505
R32611 DVSS.n9302 DVSS.n9301 2.2505
R32612 DVSS.n9299 DVSS.n2856 2.2505
R32613 DVSS.n9307 DVSS.n9306 2.2505
R32614 DVSS.n9310 DVSS.n9309 2.2505
R32615 DVSS.n9314 DVSS.n9313 2.2505
R32616 DVSS.n9311 DVSS.n2854 2.2505
R32617 DVSS.n9319 DVSS.n9318 2.2505
R32618 DVSS.n9322 DVSS.n9321 2.2505
R32619 DVSS.n9326 DVSS.n9325 2.2505
R32620 DVSS.n9323 DVSS.n2852 2.2505
R32621 DVSS.n9331 DVSS.n9330 2.2505
R32622 DVSS.n9334 DVSS.n9333 2.2505
R32623 DVSS.n9338 DVSS.n9337 2.2505
R32624 DVSS.n9335 DVSS.n2850 2.2505
R32625 DVSS.n9343 DVSS.n9342 2.2505
R32626 DVSS.n9346 DVSS.n9345 2.2505
R32627 DVSS.n9350 DVSS.n9349 2.2505
R32628 DVSS.n9347 DVSS.n2848 2.2505
R32629 DVSS.n9355 DVSS.n9354 2.2505
R32630 DVSS.n9358 DVSS.n9357 2.2505
R32631 DVSS.n9362 DVSS.n9361 2.2505
R32632 DVSS.n9359 DVSS.n2846 2.2505
R32633 DVSS.n9367 DVSS.n9366 2.2505
R32634 DVSS.n9370 DVSS.n9369 2.2505
R32635 DVSS.n9374 DVSS.n9373 2.2505
R32636 DVSS.n9371 DVSS.n2844 2.2505
R32637 DVSS.n9379 DVSS.n9378 2.2505
R32638 DVSS.n9382 DVSS.n9381 2.2505
R32639 DVSS.n9386 DVSS.n9385 2.2505
R32640 DVSS.n9383 DVSS.n2842 2.2505
R32641 DVSS.n9391 DVSS.n9390 2.2505
R32642 DVSS.n9394 DVSS.n9393 2.2505
R32643 DVSS.n9398 DVSS.n9397 2.2505
R32644 DVSS.n9395 DVSS.n2840 2.2505
R32645 DVSS.n9403 DVSS.n9402 2.2505
R32646 DVSS.n9406 DVSS.n9405 2.2505
R32647 DVSS.n9410 DVSS.n9409 2.2505
R32648 DVSS.n9407 DVSS.n2838 2.2505
R32649 DVSS.n9415 DVSS.n9414 2.2505
R32650 DVSS.n9418 DVSS.n9417 2.2505
R32651 DVSS.n9422 DVSS.n9421 2.2505
R32652 DVSS.n9419 DVSS.n2836 2.2505
R32653 DVSS.n9427 DVSS.n9426 2.2505
R32654 DVSS.n9430 DVSS.n9429 2.2505
R32655 DVSS.n9434 DVSS.n9433 2.2505
R32656 DVSS.n9431 DVSS.n2834 2.2505
R32657 DVSS.n9439 DVSS.n9438 2.2505
R32658 DVSS.n9442 DVSS.n9441 2.2505
R32659 DVSS.n9446 DVSS.n9445 2.2505
R32660 DVSS.n9443 DVSS.n2832 2.2505
R32661 DVSS.n9452 DVSS.n9451 2.2505
R32662 DVSS.n9454 DVSS.n2830 2.2505
R32663 DVSS.n9512 DVSS.n9511 2.2505
R32664 DVSS.n9513 DVSS.n9509 2.2505
R32665 DVSS.n9518 DVSS.n9514 2.2505
R32666 DVSS.n9519 DVSS.n9508 2.2505
R32667 DVSS.n9524 DVSS.n9523 2.2505
R32668 DVSS.n9525 DVSS.n9507 2.2505
R32669 DVSS.n9530 DVSS.n9526 2.2505
R32670 DVSS.n9531 DVSS.n9506 2.2505
R32671 DVSS.n9536 DVSS.n9535 2.2505
R32672 DVSS.n9537 DVSS.n9505 2.2505
R32673 DVSS.n9542 DVSS.n9538 2.2505
R32674 DVSS.n9543 DVSS.n9504 2.2505
R32675 DVSS.n9548 DVSS.n9547 2.2505
R32676 DVSS.n9549 DVSS.n9503 2.2505
R32677 DVSS.n9554 DVSS.n9550 2.2505
R32678 DVSS.n9555 DVSS.n9502 2.2505
R32679 DVSS.n9560 DVSS.n9559 2.2505
R32680 DVSS.n9561 DVSS.n9501 2.2505
R32681 DVSS.n9566 DVSS.n9562 2.2505
R32682 DVSS.n9567 DVSS.n9500 2.2505
R32683 DVSS.n9572 DVSS.n9571 2.2505
R32684 DVSS.n9573 DVSS.n9499 2.2505
R32685 DVSS.n9578 DVSS.n9574 2.2505
R32686 DVSS.n9579 DVSS.n9498 2.2505
R32687 DVSS.n9584 DVSS.n9583 2.2505
R32688 DVSS.n9585 DVSS.n9497 2.2505
R32689 DVSS.n9590 DVSS.n9586 2.2505
R32690 DVSS.n9591 DVSS.n9496 2.2505
R32691 DVSS.n9596 DVSS.n9595 2.2505
R32692 DVSS.n9597 DVSS.n9495 2.2505
R32693 DVSS.n9602 DVSS.n9598 2.2505
R32694 DVSS.n9603 DVSS.n9494 2.2505
R32695 DVSS.n9608 DVSS.n9607 2.2505
R32696 DVSS.n9609 DVSS.n9493 2.2505
R32697 DVSS.n9614 DVSS.n9610 2.2505
R32698 DVSS.n9615 DVSS.n9492 2.2505
R32699 DVSS.n9620 DVSS.n9619 2.2505
R32700 DVSS.n9621 DVSS.n9491 2.2505
R32701 DVSS.n9626 DVSS.n9622 2.2505
R32702 DVSS.n9627 DVSS.n9490 2.2505
R32703 DVSS.n9632 DVSS.n9631 2.2505
R32704 DVSS.n9633 DVSS.n9489 2.2505
R32705 DVSS.n9638 DVSS.n9634 2.2505
R32706 DVSS.n9639 DVSS.n9488 2.2505
R32707 DVSS.n9644 DVSS.n9643 2.2505
R32708 DVSS.n9645 DVSS.n9487 2.2505
R32709 DVSS.n9650 DVSS.n9646 2.2505
R32710 DVSS.n9651 DVSS.n9486 2.2505
R32711 DVSS.n9656 DVSS.n9655 2.2505
R32712 DVSS.n9657 DVSS.n9485 2.2505
R32713 DVSS.n9662 DVSS.n9658 2.2505
R32714 DVSS.n9663 DVSS.n9484 2.2505
R32715 DVSS.n9668 DVSS.n9667 2.2505
R32716 DVSS.n9669 DVSS.n9483 2.2505
R32717 DVSS.n9674 DVSS.n9670 2.2505
R32718 DVSS.n9675 DVSS.n9482 2.2505
R32719 DVSS.n9680 DVSS.n9679 2.2505
R32720 DVSS.n9681 DVSS.n9481 2.2505
R32721 DVSS.n9686 DVSS.n9682 2.2505
R32722 DVSS.n9687 DVSS.n9480 2.2505
R32723 DVSS.n9692 DVSS.n9691 2.2505
R32724 DVSS.n9693 DVSS.n9479 2.2505
R32725 DVSS.n9698 DVSS.n9694 2.2505
R32726 DVSS.n9699 DVSS.n9478 2.2505
R32727 DVSS.n9704 DVSS.n9703 2.2505
R32728 DVSS.n9705 DVSS.n9477 2.2505
R32729 DVSS.n9710 DVSS.n9706 2.2505
R32730 DVSS.n9711 DVSS.n9476 2.2505
R32731 DVSS.n9716 DVSS.n9715 2.2505
R32732 DVSS.n9717 DVSS.n9475 2.2505
R32733 DVSS.n9722 DVSS.n9718 2.2505
R32734 DVSS.n9723 DVSS.n9474 2.2505
R32735 DVSS.n9728 DVSS.n9727 2.2505
R32736 DVSS.n9729 DVSS.n9473 2.2505
R32737 DVSS.n9734 DVSS.n9730 2.2505
R32738 DVSS.n9735 DVSS.n9472 2.2505
R32739 DVSS.n9740 DVSS.n9739 2.2505
R32740 DVSS.n9741 DVSS.n9471 2.2505
R32741 DVSS.n9746 DVSS.n9742 2.2505
R32742 DVSS.n9747 DVSS.n9470 2.2505
R32743 DVSS.n9752 DVSS.n9751 2.2505
R32744 DVSS.n9753 DVSS.n9469 2.2505
R32745 DVSS.n9755 DVSS.n9754 2.2505
R32746 DVSS.n9756 DVSS.n2733 2.2505
R32747 DVSS.n9757 DVSS.n9756 2.2505
R32748 DVSS.n9755 DVSS.n9466 2.2505
R32749 DVSS.n9469 DVSS.n9468 2.2505
R32750 DVSS.n9751 DVSS.n9750 2.2505
R32751 DVSS.n9748 DVSS.n9747 2.2505
R32752 DVSS.n9746 DVSS.n9745 2.2505
R32753 DVSS.n9743 DVSS.n9471 2.2505
R32754 DVSS.n9739 DVSS.n9738 2.2505
R32755 DVSS.n9736 DVSS.n9735 2.2505
R32756 DVSS.n9734 DVSS.n9733 2.2505
R32757 DVSS.n9731 DVSS.n9473 2.2505
R32758 DVSS.n9727 DVSS.n9726 2.2505
R32759 DVSS.n9724 DVSS.n9723 2.2505
R32760 DVSS.n9722 DVSS.n9721 2.2505
R32761 DVSS.n9719 DVSS.n9475 2.2505
R32762 DVSS.n9715 DVSS.n9714 2.2505
R32763 DVSS.n9712 DVSS.n9711 2.2505
R32764 DVSS.n9710 DVSS.n9709 2.2505
R32765 DVSS.n9707 DVSS.n9477 2.2505
R32766 DVSS.n9703 DVSS.n9702 2.2505
R32767 DVSS.n9700 DVSS.n9699 2.2505
R32768 DVSS.n9698 DVSS.n9697 2.2505
R32769 DVSS.n9695 DVSS.n9479 2.2505
R32770 DVSS.n9691 DVSS.n9690 2.2505
R32771 DVSS.n9688 DVSS.n9687 2.2505
R32772 DVSS.n9686 DVSS.n9685 2.2505
R32773 DVSS.n9683 DVSS.n9481 2.2505
R32774 DVSS.n9679 DVSS.n9678 2.2505
R32775 DVSS.n9676 DVSS.n9675 2.2505
R32776 DVSS.n9674 DVSS.n9673 2.2505
R32777 DVSS.n9671 DVSS.n9483 2.2505
R32778 DVSS.n9667 DVSS.n9666 2.2505
R32779 DVSS.n9664 DVSS.n9663 2.2505
R32780 DVSS.n9662 DVSS.n9661 2.2505
R32781 DVSS.n9659 DVSS.n9485 2.2505
R32782 DVSS.n9655 DVSS.n9654 2.2505
R32783 DVSS.n9652 DVSS.n9651 2.2505
R32784 DVSS.n9650 DVSS.n9649 2.2505
R32785 DVSS.n9647 DVSS.n9487 2.2505
R32786 DVSS.n9643 DVSS.n9642 2.2505
R32787 DVSS.n9640 DVSS.n9639 2.2505
R32788 DVSS.n9638 DVSS.n9637 2.2505
R32789 DVSS.n9635 DVSS.n9489 2.2505
R32790 DVSS.n9631 DVSS.n9630 2.2505
R32791 DVSS.n9628 DVSS.n9627 2.2505
R32792 DVSS.n9626 DVSS.n9625 2.2505
R32793 DVSS.n9623 DVSS.n9491 2.2505
R32794 DVSS.n9619 DVSS.n9618 2.2505
R32795 DVSS.n9616 DVSS.n9615 2.2505
R32796 DVSS.n9614 DVSS.n9613 2.2505
R32797 DVSS.n9611 DVSS.n9493 2.2505
R32798 DVSS.n9607 DVSS.n9606 2.2505
R32799 DVSS.n9604 DVSS.n9603 2.2505
R32800 DVSS.n9602 DVSS.n9601 2.2505
R32801 DVSS.n9599 DVSS.n9495 2.2505
R32802 DVSS.n9595 DVSS.n9594 2.2505
R32803 DVSS.n9592 DVSS.n9591 2.2505
R32804 DVSS.n9590 DVSS.n9589 2.2505
R32805 DVSS.n9587 DVSS.n9497 2.2505
R32806 DVSS.n9583 DVSS.n9582 2.2505
R32807 DVSS.n9580 DVSS.n9579 2.2505
R32808 DVSS.n9578 DVSS.n9577 2.2505
R32809 DVSS.n9575 DVSS.n9499 2.2505
R32810 DVSS.n9571 DVSS.n9570 2.2505
R32811 DVSS.n9568 DVSS.n9567 2.2505
R32812 DVSS.n9566 DVSS.n9565 2.2505
R32813 DVSS.n9563 DVSS.n9501 2.2505
R32814 DVSS.n9559 DVSS.n9558 2.2505
R32815 DVSS.n9556 DVSS.n9555 2.2505
R32816 DVSS.n9554 DVSS.n9553 2.2505
R32817 DVSS.n9551 DVSS.n9503 2.2505
R32818 DVSS.n9547 DVSS.n9546 2.2505
R32819 DVSS.n9544 DVSS.n9543 2.2505
R32820 DVSS.n9542 DVSS.n9541 2.2505
R32821 DVSS.n9539 DVSS.n9505 2.2505
R32822 DVSS.n9535 DVSS.n9534 2.2505
R32823 DVSS.n9532 DVSS.n9531 2.2505
R32824 DVSS.n9530 DVSS.n9529 2.2505
R32825 DVSS.n9527 DVSS.n9507 2.2505
R32826 DVSS.n9523 DVSS.n9522 2.2505
R32827 DVSS.n9520 DVSS.n9519 2.2505
R32828 DVSS.n9518 DVSS.n9517 2.2505
R32829 DVSS.n9515 DVSS.n9509 2.2505
R32830 DVSS.n9511 DVSS.n9510 2.2505
R32831 DVSS.n10109 DVSS.n10108 2.2505
R32832 DVSS.n9777 DVSS.n9776 2.2505
R32833 DVSS.n10098 DVSS.n9778 2.2505
R32834 DVSS.n10100 DVSS.n10099 2.2505
R32835 DVSS.n10097 DVSS.n9780 2.2505
R32836 DVSS.n10096 DVSS.n10095 2.2505
R32837 DVSS.n9782 DVSS.n9781 2.2505
R32838 DVSS.n10087 DVSS.n10086 2.2505
R32839 DVSS.n10085 DVSS.n9784 2.2505
R32840 DVSS.n10084 DVSS.n10083 2.2505
R32841 DVSS.n9786 DVSS.n9785 2.2505
R32842 DVSS.n10075 DVSS.n10074 2.2505
R32843 DVSS.n10073 DVSS.n9788 2.2505
R32844 DVSS.n10072 DVSS.n10071 2.2505
R32845 DVSS.n9790 DVSS.n9789 2.2505
R32846 DVSS.n10063 DVSS.n10062 2.2505
R32847 DVSS.n10061 DVSS.n9792 2.2505
R32848 DVSS.n10060 DVSS.n10059 2.2505
R32849 DVSS.n9794 DVSS.n9793 2.2505
R32850 DVSS.n10051 DVSS.n10050 2.2505
R32851 DVSS.n10049 DVSS.n9796 2.2505
R32852 DVSS.n10048 DVSS.n10047 2.2505
R32853 DVSS.n9798 DVSS.n9797 2.2505
R32854 DVSS.n10039 DVSS.n10038 2.2505
R32855 DVSS.n10037 DVSS.n9800 2.2505
R32856 DVSS.n10036 DVSS.n10035 2.2505
R32857 DVSS.n9802 DVSS.n9801 2.2505
R32858 DVSS.n10027 DVSS.n10026 2.2505
R32859 DVSS.n10025 DVSS.n9804 2.2505
R32860 DVSS.n10024 DVSS.n10023 2.2505
R32861 DVSS.n9806 DVSS.n9805 2.2505
R32862 DVSS.n10015 DVSS.n10014 2.2505
R32863 DVSS.n10013 DVSS.n9808 2.2505
R32864 DVSS.n10012 DVSS.n10011 2.2505
R32865 DVSS.n9810 DVSS.n9809 2.2505
R32866 DVSS.n10003 DVSS.n10002 2.2505
R32867 DVSS.n10001 DVSS.n9812 2.2505
R32868 DVSS.n10000 DVSS.n9999 2.2505
R32869 DVSS.n9814 DVSS.n9813 2.2505
R32870 DVSS.n9991 DVSS.n9990 2.2505
R32871 DVSS.n9989 DVSS.n9816 2.2505
R32872 DVSS.n9988 DVSS.n9987 2.2505
R32873 DVSS.n9818 DVSS.n9817 2.2505
R32874 DVSS.n9979 DVSS.n9978 2.2505
R32875 DVSS.n9977 DVSS.n9820 2.2505
R32876 DVSS.n9976 DVSS.n9975 2.2505
R32877 DVSS.n9822 DVSS.n9821 2.2505
R32878 DVSS.n9967 DVSS.n9966 2.2505
R32879 DVSS.n9965 DVSS.n9824 2.2505
R32880 DVSS.n9964 DVSS.n9963 2.2505
R32881 DVSS.n9826 DVSS.n9825 2.2505
R32882 DVSS.n9955 DVSS.n9954 2.2505
R32883 DVSS.n9953 DVSS.n9828 2.2505
R32884 DVSS.n9952 DVSS.n9951 2.2505
R32885 DVSS.n9830 DVSS.n9829 2.2505
R32886 DVSS.n9943 DVSS.n9942 2.2505
R32887 DVSS.n9941 DVSS.n9832 2.2505
R32888 DVSS.n9940 DVSS.n9939 2.2505
R32889 DVSS.n9834 DVSS.n9833 2.2505
R32890 DVSS.n9931 DVSS.n9930 2.2505
R32891 DVSS.n9929 DVSS.n9836 2.2505
R32892 DVSS.n9928 DVSS.n9927 2.2505
R32893 DVSS.n9838 DVSS.n9837 2.2505
R32894 DVSS.n9919 DVSS.n9918 2.2505
R32895 DVSS.n9917 DVSS.n9840 2.2505
R32896 DVSS.n9916 DVSS.n9915 2.2505
R32897 DVSS.n9842 DVSS.n9841 2.2505
R32898 DVSS.n9907 DVSS.n9906 2.2505
R32899 DVSS.n9905 DVSS.n9844 2.2505
R32900 DVSS.n9904 DVSS.n9903 2.2505
R32901 DVSS.n9846 DVSS.n9845 2.2505
R32902 DVSS.n9895 DVSS.n9894 2.2505
R32903 DVSS.n9893 DVSS.n9848 2.2505
R32904 DVSS.n9892 DVSS.n9891 2.2505
R32905 DVSS.n9850 DVSS.n9849 2.2505
R32906 DVSS.n9883 DVSS.n9882 2.2505
R32907 DVSS.n9881 DVSS.n9852 2.2505
R32908 DVSS.n9880 DVSS.n9879 2.2505
R32909 DVSS.n9854 DVSS.n9853 2.2505
R32910 DVSS.n9871 DVSS.n9870 2.2505
R32911 DVSS.n9869 DVSS.n9856 2.2505
R32912 DVSS.n9868 DVSS.n9867 2.2505
R32913 DVSS.n9858 DVSS.n9857 2.2505
R32914 DVSS.n9859 DVSS.n2712 2.2505
R32915 DVSS.n9860 DVSS.n9859 2.2505
R32916 DVSS.n9862 DVSS.n9858 2.2505
R32917 DVSS.n9867 DVSS.n9866 2.2505
R32918 DVSS.n9864 DVSS.n9856 2.2505
R32919 DVSS.n9872 DVSS.n9871 2.2505
R32920 DVSS.n9874 DVSS.n9854 2.2505
R32921 DVSS.n9879 DVSS.n9878 2.2505
R32922 DVSS.n9876 DVSS.n9852 2.2505
R32923 DVSS.n9884 DVSS.n9883 2.2505
R32924 DVSS.n9886 DVSS.n9850 2.2505
R32925 DVSS.n9891 DVSS.n9890 2.2505
R32926 DVSS.n9888 DVSS.n9848 2.2505
R32927 DVSS.n9896 DVSS.n9895 2.2505
R32928 DVSS.n9898 DVSS.n9846 2.2505
R32929 DVSS.n9903 DVSS.n9902 2.2505
R32930 DVSS.n9900 DVSS.n9844 2.2505
R32931 DVSS.n9908 DVSS.n9907 2.2505
R32932 DVSS.n9910 DVSS.n9842 2.2505
R32933 DVSS.n9915 DVSS.n9914 2.2505
R32934 DVSS.n9912 DVSS.n9840 2.2505
R32935 DVSS.n9920 DVSS.n9919 2.2505
R32936 DVSS.n9922 DVSS.n9838 2.2505
R32937 DVSS.n9927 DVSS.n9926 2.2505
R32938 DVSS.n9924 DVSS.n9836 2.2505
R32939 DVSS.n9932 DVSS.n9931 2.2505
R32940 DVSS.n9934 DVSS.n9834 2.2505
R32941 DVSS.n9939 DVSS.n9938 2.2505
R32942 DVSS.n9936 DVSS.n9832 2.2505
R32943 DVSS.n9944 DVSS.n9943 2.2505
R32944 DVSS.n9946 DVSS.n9830 2.2505
R32945 DVSS.n9951 DVSS.n9950 2.2505
R32946 DVSS.n9948 DVSS.n9828 2.2505
R32947 DVSS.n9956 DVSS.n9955 2.2505
R32948 DVSS.n9958 DVSS.n9826 2.2505
R32949 DVSS.n9963 DVSS.n9962 2.2505
R32950 DVSS.n9960 DVSS.n9824 2.2505
R32951 DVSS.n9968 DVSS.n9967 2.2505
R32952 DVSS.n9970 DVSS.n9822 2.2505
R32953 DVSS.n9975 DVSS.n9974 2.2505
R32954 DVSS.n9972 DVSS.n9820 2.2505
R32955 DVSS.n9980 DVSS.n9979 2.2505
R32956 DVSS.n9982 DVSS.n9818 2.2505
R32957 DVSS.n9987 DVSS.n9986 2.2505
R32958 DVSS.n9984 DVSS.n9816 2.2505
R32959 DVSS.n9992 DVSS.n9991 2.2505
R32960 DVSS.n9994 DVSS.n9814 2.2505
R32961 DVSS.n9999 DVSS.n9998 2.2505
R32962 DVSS.n9996 DVSS.n9812 2.2505
R32963 DVSS.n10004 DVSS.n10003 2.2505
R32964 DVSS.n10006 DVSS.n9810 2.2505
R32965 DVSS.n10011 DVSS.n10010 2.2505
R32966 DVSS.n10008 DVSS.n9808 2.2505
R32967 DVSS.n10016 DVSS.n10015 2.2505
R32968 DVSS.n10018 DVSS.n9806 2.2505
R32969 DVSS.n10023 DVSS.n10022 2.2505
R32970 DVSS.n10020 DVSS.n9804 2.2505
R32971 DVSS.n10028 DVSS.n10027 2.2505
R32972 DVSS.n10030 DVSS.n9802 2.2505
R32973 DVSS.n10035 DVSS.n10034 2.2505
R32974 DVSS.n10032 DVSS.n9800 2.2505
R32975 DVSS.n10040 DVSS.n10039 2.2505
R32976 DVSS.n10042 DVSS.n9798 2.2505
R32977 DVSS.n10047 DVSS.n10046 2.2505
R32978 DVSS.n10044 DVSS.n9796 2.2505
R32979 DVSS.n10052 DVSS.n10051 2.2505
R32980 DVSS.n10054 DVSS.n9794 2.2505
R32981 DVSS.n10059 DVSS.n10058 2.2505
R32982 DVSS.n10056 DVSS.n9792 2.2505
R32983 DVSS.n10064 DVSS.n10063 2.2505
R32984 DVSS.n10066 DVSS.n9790 2.2505
R32985 DVSS.n10071 DVSS.n10070 2.2505
R32986 DVSS.n10068 DVSS.n9788 2.2505
R32987 DVSS.n10076 DVSS.n10075 2.2505
R32988 DVSS.n10078 DVSS.n9786 2.2505
R32989 DVSS.n10083 DVSS.n10082 2.2505
R32990 DVSS.n10080 DVSS.n9784 2.2505
R32991 DVSS.n10088 DVSS.n10087 2.2505
R32992 DVSS.n10090 DVSS.n9782 2.2505
R32993 DVSS.n10095 DVSS.n10094 2.2505
R32994 DVSS.n10092 DVSS.n9780 2.2505
R32995 DVSS.n10101 DVSS.n10100 2.2505
R32996 DVSS.n10103 DVSS.n9778 2.2505
R32997 DVSS.n10105 DVSS.n9777 2.2505
R32998 DVSS.n10108 DVSS.n10107 2.2505
R32999 DVSS.n10135 DVSS.n2414 2.2505
R33000 DVSS.n10137 DVSS.n10136 2.2505
R33001 DVSS.n2701 DVSS.n2416 2.2505
R33002 DVSS.n2700 DVSS.n2699 2.2505
R33003 DVSS.n2695 DVSS.n2417 2.2505
R33004 DVSS.n2691 DVSS.n2690 2.2505
R33005 DVSS.n2689 DVSS.n2418 2.2505
R33006 DVSS.n2688 DVSS.n2687 2.2505
R33007 DVSS.n2683 DVSS.n2419 2.2505
R33008 DVSS.n2679 DVSS.n2678 2.2505
R33009 DVSS.n2677 DVSS.n2420 2.2505
R33010 DVSS.n2676 DVSS.n2675 2.2505
R33011 DVSS.n2671 DVSS.n2421 2.2505
R33012 DVSS.n2667 DVSS.n2666 2.2505
R33013 DVSS.n2665 DVSS.n2422 2.2505
R33014 DVSS.n2664 DVSS.n2663 2.2505
R33015 DVSS.n2659 DVSS.n2423 2.2505
R33016 DVSS.n2655 DVSS.n2654 2.2505
R33017 DVSS.n2653 DVSS.n2424 2.2505
R33018 DVSS.n2652 DVSS.n2651 2.2505
R33019 DVSS.n2647 DVSS.n2425 2.2505
R33020 DVSS.n2643 DVSS.n2642 2.2505
R33021 DVSS.n2641 DVSS.n2426 2.2505
R33022 DVSS.n2640 DVSS.n2639 2.2505
R33023 DVSS.n2635 DVSS.n2427 2.2505
R33024 DVSS.n2631 DVSS.n2630 2.2505
R33025 DVSS.n2629 DVSS.n2428 2.2505
R33026 DVSS.n2628 DVSS.n2627 2.2505
R33027 DVSS.n2623 DVSS.n2429 2.2505
R33028 DVSS.n2619 DVSS.n2618 2.2505
R33029 DVSS.n2617 DVSS.n2430 2.2505
R33030 DVSS.n2616 DVSS.n2615 2.2505
R33031 DVSS.n2611 DVSS.n2431 2.2505
R33032 DVSS.n2607 DVSS.n2606 2.2505
R33033 DVSS.n2605 DVSS.n2432 2.2505
R33034 DVSS.n2604 DVSS.n2603 2.2505
R33035 DVSS.n2599 DVSS.n2433 2.2505
R33036 DVSS.n2595 DVSS.n2594 2.2505
R33037 DVSS.n2593 DVSS.n2434 2.2505
R33038 DVSS.n2592 DVSS.n2591 2.2505
R33039 DVSS.n2587 DVSS.n2435 2.2505
R33040 DVSS.n2583 DVSS.n2582 2.2505
R33041 DVSS.n2581 DVSS.n2436 2.2505
R33042 DVSS.n2580 DVSS.n2579 2.2505
R33043 DVSS.n2575 DVSS.n2437 2.2505
R33044 DVSS.n2571 DVSS.n2570 2.2505
R33045 DVSS.n2569 DVSS.n2438 2.2505
R33046 DVSS.n2568 DVSS.n2567 2.2505
R33047 DVSS.n2563 DVSS.n2439 2.2505
R33048 DVSS.n2559 DVSS.n2558 2.2505
R33049 DVSS.n2557 DVSS.n2440 2.2505
R33050 DVSS.n2556 DVSS.n2555 2.2505
R33051 DVSS.n2551 DVSS.n2441 2.2505
R33052 DVSS.n2547 DVSS.n2546 2.2505
R33053 DVSS.n2545 DVSS.n2442 2.2505
R33054 DVSS.n2544 DVSS.n2543 2.2505
R33055 DVSS.n2539 DVSS.n2443 2.2505
R33056 DVSS.n2535 DVSS.n2534 2.2505
R33057 DVSS.n2533 DVSS.n2444 2.2505
R33058 DVSS.n2532 DVSS.n2531 2.2505
R33059 DVSS.n2527 DVSS.n2445 2.2505
R33060 DVSS.n2523 DVSS.n2522 2.2505
R33061 DVSS.n2521 DVSS.n2446 2.2505
R33062 DVSS.n2520 DVSS.n2519 2.2505
R33063 DVSS.n2515 DVSS.n2447 2.2505
R33064 DVSS.n2511 DVSS.n2510 2.2505
R33065 DVSS.n2509 DVSS.n2448 2.2505
R33066 DVSS.n2508 DVSS.n2507 2.2505
R33067 DVSS.n2503 DVSS.n2449 2.2505
R33068 DVSS.n2499 DVSS.n2498 2.2505
R33069 DVSS.n2497 DVSS.n2450 2.2505
R33070 DVSS.n2496 DVSS.n2495 2.2505
R33071 DVSS.n2491 DVSS.n2451 2.2505
R33072 DVSS.n2487 DVSS.n2486 2.2505
R33073 DVSS.n2485 DVSS.n2452 2.2505
R33074 DVSS.n2484 DVSS.n2483 2.2505
R33075 DVSS.n2479 DVSS.n2453 2.2505
R33076 DVSS.n2475 DVSS.n2474 2.2505
R33077 DVSS.n2473 DVSS.n2454 2.2505
R33078 DVSS.n2472 DVSS.n2471 2.2505
R33079 DVSS.n2467 DVSS.n2455 2.2505
R33080 DVSS.n2463 DVSS.n2462 2.2505
R33081 DVSS.n2461 DVSS.n2458 2.2505
R33082 DVSS.n2460 DVSS.n2459 2.2505
R33083 DVSS.n2459 DVSS.n2412 2.2505
R33084 DVSS.n2458 DVSS.n2457 2.2505
R33085 DVSS.n2464 DVSS.n2463 2.2505
R33086 DVSS.n2467 DVSS.n2466 2.2505
R33087 DVSS.n2471 DVSS.n2470 2.2505
R33088 DVSS.n2468 DVSS.n2454 2.2505
R33089 DVSS.n2476 DVSS.n2475 2.2505
R33090 DVSS.n2479 DVSS.n2478 2.2505
R33091 DVSS.n2483 DVSS.n2482 2.2505
R33092 DVSS.n2480 DVSS.n2452 2.2505
R33093 DVSS.n2488 DVSS.n2487 2.2505
R33094 DVSS.n2491 DVSS.n2490 2.2505
R33095 DVSS.n2495 DVSS.n2494 2.2505
R33096 DVSS.n2492 DVSS.n2450 2.2505
R33097 DVSS.n2500 DVSS.n2499 2.2505
R33098 DVSS.n2503 DVSS.n2502 2.2505
R33099 DVSS.n2507 DVSS.n2506 2.2505
R33100 DVSS.n2504 DVSS.n2448 2.2505
R33101 DVSS.n2512 DVSS.n2511 2.2505
R33102 DVSS.n2515 DVSS.n2514 2.2505
R33103 DVSS.n2519 DVSS.n2518 2.2505
R33104 DVSS.n2516 DVSS.n2446 2.2505
R33105 DVSS.n2524 DVSS.n2523 2.2505
R33106 DVSS.n2527 DVSS.n2526 2.2505
R33107 DVSS.n2531 DVSS.n2530 2.2505
R33108 DVSS.n2528 DVSS.n2444 2.2505
R33109 DVSS.n2536 DVSS.n2535 2.2505
R33110 DVSS.n2539 DVSS.n2538 2.2505
R33111 DVSS.n2543 DVSS.n2542 2.2505
R33112 DVSS.n2540 DVSS.n2442 2.2505
R33113 DVSS.n2548 DVSS.n2547 2.2505
R33114 DVSS.n2551 DVSS.n2550 2.2505
R33115 DVSS.n2555 DVSS.n2554 2.2505
R33116 DVSS.n2552 DVSS.n2440 2.2505
R33117 DVSS.n2560 DVSS.n2559 2.2505
R33118 DVSS.n2563 DVSS.n2562 2.2505
R33119 DVSS.n2567 DVSS.n2566 2.2505
R33120 DVSS.n2564 DVSS.n2438 2.2505
R33121 DVSS.n2572 DVSS.n2571 2.2505
R33122 DVSS.n2575 DVSS.n2574 2.2505
R33123 DVSS.n2579 DVSS.n2578 2.2505
R33124 DVSS.n2576 DVSS.n2436 2.2505
R33125 DVSS.n2584 DVSS.n2583 2.2505
R33126 DVSS.n2587 DVSS.n2586 2.2505
R33127 DVSS.n2591 DVSS.n2590 2.2505
R33128 DVSS.n2588 DVSS.n2434 2.2505
R33129 DVSS.n2596 DVSS.n2595 2.2505
R33130 DVSS.n2599 DVSS.n2598 2.2505
R33131 DVSS.n2603 DVSS.n2602 2.2505
R33132 DVSS.n2600 DVSS.n2432 2.2505
R33133 DVSS.n2608 DVSS.n2607 2.2505
R33134 DVSS.n2611 DVSS.n2610 2.2505
R33135 DVSS.n2615 DVSS.n2614 2.2505
R33136 DVSS.n2612 DVSS.n2430 2.2505
R33137 DVSS.n2620 DVSS.n2619 2.2505
R33138 DVSS.n2623 DVSS.n2622 2.2505
R33139 DVSS.n2627 DVSS.n2626 2.2505
R33140 DVSS.n2624 DVSS.n2428 2.2505
R33141 DVSS.n2632 DVSS.n2631 2.2505
R33142 DVSS.n2635 DVSS.n2634 2.2505
R33143 DVSS.n2639 DVSS.n2638 2.2505
R33144 DVSS.n2636 DVSS.n2426 2.2505
R33145 DVSS.n2644 DVSS.n2643 2.2505
R33146 DVSS.n2647 DVSS.n2646 2.2505
R33147 DVSS.n2651 DVSS.n2650 2.2505
R33148 DVSS.n2648 DVSS.n2424 2.2505
R33149 DVSS.n2656 DVSS.n2655 2.2505
R33150 DVSS.n2659 DVSS.n2658 2.2505
R33151 DVSS.n2663 DVSS.n2662 2.2505
R33152 DVSS.n2660 DVSS.n2422 2.2505
R33153 DVSS.n2668 DVSS.n2667 2.2505
R33154 DVSS.n2671 DVSS.n2670 2.2505
R33155 DVSS.n2675 DVSS.n2674 2.2505
R33156 DVSS.n2672 DVSS.n2420 2.2505
R33157 DVSS.n2680 DVSS.n2679 2.2505
R33158 DVSS.n2683 DVSS.n2682 2.2505
R33159 DVSS.n2687 DVSS.n2686 2.2505
R33160 DVSS.n2684 DVSS.n2418 2.2505
R33161 DVSS.n2692 DVSS.n2691 2.2505
R33162 DVSS.n2695 DVSS.n2694 2.2505
R33163 DVSS.n2699 DVSS.n2698 2.2505
R33164 DVSS.n2696 DVSS.n2416 2.2505
R33165 DVSS.n10138 DVSS.n10137 2.2505
R33166 DVSS.n10140 DVSS.n2414 2.2505
R33167 DVSS.n10160 DVSS.n2072 2.2505
R33168 DVSS.n10162 DVSS.n10161 2.2505
R33169 DVSS.n2359 DVSS.n2074 2.2505
R33170 DVSS.n2358 DVSS.n2357 2.2505
R33171 DVSS.n2353 DVSS.n2075 2.2505
R33172 DVSS.n2349 DVSS.n2348 2.2505
R33173 DVSS.n2347 DVSS.n2076 2.2505
R33174 DVSS.n2346 DVSS.n2345 2.2505
R33175 DVSS.n2341 DVSS.n2077 2.2505
R33176 DVSS.n2337 DVSS.n2336 2.2505
R33177 DVSS.n2335 DVSS.n2078 2.2505
R33178 DVSS.n2334 DVSS.n2333 2.2505
R33179 DVSS.n2329 DVSS.n2079 2.2505
R33180 DVSS.n2325 DVSS.n2324 2.2505
R33181 DVSS.n2323 DVSS.n2080 2.2505
R33182 DVSS.n2322 DVSS.n2321 2.2505
R33183 DVSS.n2317 DVSS.n2081 2.2505
R33184 DVSS.n2313 DVSS.n2312 2.2505
R33185 DVSS.n2311 DVSS.n2082 2.2505
R33186 DVSS.n2310 DVSS.n2309 2.2505
R33187 DVSS.n2305 DVSS.n2083 2.2505
R33188 DVSS.n2301 DVSS.n2300 2.2505
R33189 DVSS.n2299 DVSS.n2084 2.2505
R33190 DVSS.n2298 DVSS.n2297 2.2505
R33191 DVSS.n2293 DVSS.n2085 2.2505
R33192 DVSS.n2289 DVSS.n2288 2.2505
R33193 DVSS.n2287 DVSS.n2086 2.2505
R33194 DVSS.n2286 DVSS.n2285 2.2505
R33195 DVSS.n2281 DVSS.n2087 2.2505
R33196 DVSS.n2277 DVSS.n2276 2.2505
R33197 DVSS.n2275 DVSS.n2088 2.2505
R33198 DVSS.n2274 DVSS.n2273 2.2505
R33199 DVSS.n2269 DVSS.n2089 2.2505
R33200 DVSS.n2265 DVSS.n2264 2.2505
R33201 DVSS.n2263 DVSS.n2090 2.2505
R33202 DVSS.n2262 DVSS.n2261 2.2505
R33203 DVSS.n2257 DVSS.n2091 2.2505
R33204 DVSS.n2253 DVSS.n2252 2.2505
R33205 DVSS.n2251 DVSS.n2092 2.2505
R33206 DVSS.n2250 DVSS.n2249 2.2505
R33207 DVSS.n2245 DVSS.n2093 2.2505
R33208 DVSS.n2241 DVSS.n2240 2.2505
R33209 DVSS.n2239 DVSS.n2094 2.2505
R33210 DVSS.n2238 DVSS.n2237 2.2505
R33211 DVSS.n2233 DVSS.n2095 2.2505
R33212 DVSS.n2229 DVSS.n2228 2.2505
R33213 DVSS.n2227 DVSS.n2096 2.2505
R33214 DVSS.n2226 DVSS.n2225 2.2505
R33215 DVSS.n2221 DVSS.n2097 2.2505
R33216 DVSS.n2217 DVSS.n2216 2.2505
R33217 DVSS.n2215 DVSS.n2098 2.2505
R33218 DVSS.n2214 DVSS.n2213 2.2505
R33219 DVSS.n2209 DVSS.n2099 2.2505
R33220 DVSS.n2205 DVSS.n2204 2.2505
R33221 DVSS.n2203 DVSS.n2100 2.2505
R33222 DVSS.n2202 DVSS.n2201 2.2505
R33223 DVSS.n2197 DVSS.n2101 2.2505
R33224 DVSS.n2193 DVSS.n2192 2.2505
R33225 DVSS.n2191 DVSS.n2102 2.2505
R33226 DVSS.n2190 DVSS.n2189 2.2505
R33227 DVSS.n2185 DVSS.n2103 2.2505
R33228 DVSS.n2181 DVSS.n2180 2.2505
R33229 DVSS.n2179 DVSS.n2104 2.2505
R33230 DVSS.n2178 DVSS.n2177 2.2505
R33231 DVSS.n2173 DVSS.n2105 2.2505
R33232 DVSS.n2169 DVSS.n2168 2.2505
R33233 DVSS.n2167 DVSS.n2106 2.2505
R33234 DVSS.n2166 DVSS.n2165 2.2505
R33235 DVSS.n2161 DVSS.n2107 2.2505
R33236 DVSS.n2157 DVSS.n2156 2.2505
R33237 DVSS.n2155 DVSS.n2108 2.2505
R33238 DVSS.n2154 DVSS.n2153 2.2505
R33239 DVSS.n2149 DVSS.n2109 2.2505
R33240 DVSS.n2145 DVSS.n2144 2.2505
R33241 DVSS.n2143 DVSS.n2110 2.2505
R33242 DVSS.n2142 DVSS.n2141 2.2505
R33243 DVSS.n2137 DVSS.n2111 2.2505
R33244 DVSS.n2133 DVSS.n2132 2.2505
R33245 DVSS.n2131 DVSS.n2112 2.2505
R33246 DVSS.n2130 DVSS.n2129 2.2505
R33247 DVSS.n2125 DVSS.n2113 2.2505
R33248 DVSS.n2121 DVSS.n2120 2.2505
R33249 DVSS.n2119 DVSS.n2116 2.2505
R33250 DVSS.n2118 DVSS.n2117 2.2505
R33251 DVSS.n2117 DVSS.n2069 2.2505
R33252 DVSS.n2116 DVSS.n2115 2.2505
R33253 DVSS.n2122 DVSS.n2121 2.2505
R33254 DVSS.n2125 DVSS.n2124 2.2505
R33255 DVSS.n2129 DVSS.n2128 2.2505
R33256 DVSS.n2126 DVSS.n2112 2.2505
R33257 DVSS.n2134 DVSS.n2133 2.2505
R33258 DVSS.n2137 DVSS.n2136 2.2505
R33259 DVSS.n2141 DVSS.n2140 2.2505
R33260 DVSS.n2138 DVSS.n2110 2.2505
R33261 DVSS.n2146 DVSS.n2145 2.2505
R33262 DVSS.n2149 DVSS.n2148 2.2505
R33263 DVSS.n2153 DVSS.n2152 2.2505
R33264 DVSS.n2150 DVSS.n2108 2.2505
R33265 DVSS.n2158 DVSS.n2157 2.2505
R33266 DVSS.n2161 DVSS.n2160 2.2505
R33267 DVSS.n2165 DVSS.n2164 2.2505
R33268 DVSS.n2162 DVSS.n2106 2.2505
R33269 DVSS.n2170 DVSS.n2169 2.2505
R33270 DVSS.n2173 DVSS.n2172 2.2505
R33271 DVSS.n2177 DVSS.n2176 2.2505
R33272 DVSS.n2174 DVSS.n2104 2.2505
R33273 DVSS.n2182 DVSS.n2181 2.2505
R33274 DVSS.n2185 DVSS.n2184 2.2505
R33275 DVSS.n2189 DVSS.n2188 2.2505
R33276 DVSS.n2186 DVSS.n2102 2.2505
R33277 DVSS.n2194 DVSS.n2193 2.2505
R33278 DVSS.n2197 DVSS.n2196 2.2505
R33279 DVSS.n2201 DVSS.n2200 2.2505
R33280 DVSS.n2198 DVSS.n2100 2.2505
R33281 DVSS.n2206 DVSS.n2205 2.2505
R33282 DVSS.n2209 DVSS.n2208 2.2505
R33283 DVSS.n2213 DVSS.n2212 2.2505
R33284 DVSS.n2210 DVSS.n2098 2.2505
R33285 DVSS.n2218 DVSS.n2217 2.2505
R33286 DVSS.n2221 DVSS.n2220 2.2505
R33287 DVSS.n2225 DVSS.n2224 2.2505
R33288 DVSS.n2222 DVSS.n2096 2.2505
R33289 DVSS.n2230 DVSS.n2229 2.2505
R33290 DVSS.n2233 DVSS.n2232 2.2505
R33291 DVSS.n2237 DVSS.n2236 2.2505
R33292 DVSS.n2234 DVSS.n2094 2.2505
R33293 DVSS.n2242 DVSS.n2241 2.2505
R33294 DVSS.n2245 DVSS.n2244 2.2505
R33295 DVSS.n2249 DVSS.n2248 2.2505
R33296 DVSS.n2246 DVSS.n2092 2.2505
R33297 DVSS.n2254 DVSS.n2253 2.2505
R33298 DVSS.n2257 DVSS.n2256 2.2505
R33299 DVSS.n2261 DVSS.n2260 2.2505
R33300 DVSS.n2258 DVSS.n2090 2.2505
R33301 DVSS.n2266 DVSS.n2265 2.2505
R33302 DVSS.n2269 DVSS.n2268 2.2505
R33303 DVSS.n2273 DVSS.n2272 2.2505
R33304 DVSS.n2270 DVSS.n2088 2.2505
R33305 DVSS.n2278 DVSS.n2277 2.2505
R33306 DVSS.n2281 DVSS.n2280 2.2505
R33307 DVSS.n2285 DVSS.n2284 2.2505
R33308 DVSS.n2282 DVSS.n2086 2.2505
R33309 DVSS.n2290 DVSS.n2289 2.2505
R33310 DVSS.n2293 DVSS.n2292 2.2505
R33311 DVSS.n2297 DVSS.n2296 2.2505
R33312 DVSS.n2294 DVSS.n2084 2.2505
R33313 DVSS.n2302 DVSS.n2301 2.2505
R33314 DVSS.n2305 DVSS.n2304 2.2505
R33315 DVSS.n2309 DVSS.n2308 2.2505
R33316 DVSS.n2306 DVSS.n2082 2.2505
R33317 DVSS.n2314 DVSS.n2313 2.2505
R33318 DVSS.n2317 DVSS.n2316 2.2505
R33319 DVSS.n2321 DVSS.n2320 2.2505
R33320 DVSS.n2318 DVSS.n2080 2.2505
R33321 DVSS.n2326 DVSS.n2325 2.2505
R33322 DVSS.n2329 DVSS.n2328 2.2505
R33323 DVSS.n2333 DVSS.n2332 2.2505
R33324 DVSS.n2330 DVSS.n2078 2.2505
R33325 DVSS.n2338 DVSS.n2337 2.2505
R33326 DVSS.n2341 DVSS.n2340 2.2505
R33327 DVSS.n2345 DVSS.n2344 2.2505
R33328 DVSS.n2342 DVSS.n2076 2.2505
R33329 DVSS.n2350 DVSS.n2349 2.2505
R33330 DVSS.n2353 DVSS.n2352 2.2505
R33331 DVSS.n2357 DVSS.n2356 2.2505
R33332 DVSS.n2354 DVSS.n2074 2.2505
R33333 DVSS.n10163 DVSS.n10162 2.2505
R33334 DVSS.n10165 DVSS.n2072 2.2505
R33335 DVSS.n10469 DVSS.n2011 2.2505
R33336 DVSS.n10471 DVSS.n10470 2.2505
R33337 DVSS.n2015 DVSS.n2014 2.2505
R33338 DVSS.n10216 DVSS.n10215 2.2505
R33339 DVSS.n10217 DVSS.n10211 2.2505
R33340 DVSS.n10222 DVSS.n10218 2.2505
R33341 DVSS.n10223 DVSS.n10210 2.2505
R33342 DVSS.n10228 DVSS.n10227 2.2505
R33343 DVSS.n10229 DVSS.n10209 2.2505
R33344 DVSS.n10234 DVSS.n10230 2.2505
R33345 DVSS.n10235 DVSS.n10208 2.2505
R33346 DVSS.n10240 DVSS.n10239 2.2505
R33347 DVSS.n10241 DVSS.n10207 2.2505
R33348 DVSS.n10246 DVSS.n10242 2.2505
R33349 DVSS.n10247 DVSS.n10206 2.2505
R33350 DVSS.n10252 DVSS.n10251 2.2505
R33351 DVSS.n10253 DVSS.n10205 2.2505
R33352 DVSS.n10258 DVSS.n10254 2.2505
R33353 DVSS.n10259 DVSS.n10204 2.2505
R33354 DVSS.n10264 DVSS.n10263 2.2505
R33355 DVSS.n10265 DVSS.n10203 2.2505
R33356 DVSS.n10270 DVSS.n10266 2.2505
R33357 DVSS.n10271 DVSS.n10202 2.2505
R33358 DVSS.n10276 DVSS.n10275 2.2505
R33359 DVSS.n10277 DVSS.n10201 2.2505
R33360 DVSS.n10282 DVSS.n10278 2.2505
R33361 DVSS.n10283 DVSS.n10200 2.2505
R33362 DVSS.n10288 DVSS.n10287 2.2505
R33363 DVSS.n10289 DVSS.n10199 2.2505
R33364 DVSS.n10294 DVSS.n10290 2.2505
R33365 DVSS.n10295 DVSS.n10198 2.2505
R33366 DVSS.n10300 DVSS.n10299 2.2505
R33367 DVSS.n10301 DVSS.n10197 2.2505
R33368 DVSS.n10306 DVSS.n10302 2.2505
R33369 DVSS.n10307 DVSS.n10196 2.2505
R33370 DVSS.n10312 DVSS.n10311 2.2505
R33371 DVSS.n10313 DVSS.n10195 2.2505
R33372 DVSS.n10318 DVSS.n10314 2.2505
R33373 DVSS.n10319 DVSS.n10194 2.2505
R33374 DVSS.n10324 DVSS.n10323 2.2505
R33375 DVSS.n10325 DVSS.n10193 2.2505
R33376 DVSS.n10330 DVSS.n10326 2.2505
R33377 DVSS.n10331 DVSS.n10192 2.2505
R33378 DVSS.n10336 DVSS.n10335 2.2505
R33379 DVSS.n10337 DVSS.n10191 2.2505
R33380 DVSS.n10342 DVSS.n10338 2.2505
R33381 DVSS.n10343 DVSS.n10190 2.2505
R33382 DVSS.n10348 DVSS.n10347 2.2505
R33383 DVSS.n10349 DVSS.n10189 2.2505
R33384 DVSS.n10354 DVSS.n10350 2.2505
R33385 DVSS.n10355 DVSS.n10188 2.2505
R33386 DVSS.n10360 DVSS.n10359 2.2505
R33387 DVSS.n10361 DVSS.n10187 2.2505
R33388 DVSS.n10366 DVSS.n10362 2.2505
R33389 DVSS.n10367 DVSS.n10186 2.2505
R33390 DVSS.n10372 DVSS.n10371 2.2505
R33391 DVSS.n10373 DVSS.n10185 2.2505
R33392 DVSS.n10378 DVSS.n10374 2.2505
R33393 DVSS.n10379 DVSS.n10184 2.2505
R33394 DVSS.n10384 DVSS.n10383 2.2505
R33395 DVSS.n10385 DVSS.n10183 2.2505
R33396 DVSS.n10390 DVSS.n10386 2.2505
R33397 DVSS.n10391 DVSS.n10182 2.2505
R33398 DVSS.n10396 DVSS.n10395 2.2505
R33399 DVSS.n10397 DVSS.n10181 2.2505
R33400 DVSS.n10402 DVSS.n10398 2.2505
R33401 DVSS.n10403 DVSS.n10180 2.2505
R33402 DVSS.n10408 DVSS.n10407 2.2505
R33403 DVSS.n10409 DVSS.n10179 2.2505
R33404 DVSS.n10414 DVSS.n10410 2.2505
R33405 DVSS.n10415 DVSS.n10178 2.2505
R33406 DVSS.n10420 DVSS.n10419 2.2505
R33407 DVSS.n10421 DVSS.n10177 2.2505
R33408 DVSS.n10426 DVSS.n10422 2.2505
R33409 DVSS.n10427 DVSS.n10176 2.2505
R33410 DVSS.n10432 DVSS.n10431 2.2505
R33411 DVSS.n10433 DVSS.n10175 2.2505
R33412 DVSS.n10438 DVSS.n10434 2.2505
R33413 DVSS.n10439 DVSS.n10174 2.2505
R33414 DVSS.n10444 DVSS.n10443 2.2505
R33415 DVSS.n10445 DVSS.n10173 2.2505
R33416 DVSS.n10450 DVSS.n10446 2.2505
R33417 DVSS.n10453 DVSS.n10172 2.2505
R33418 DVSS.n10455 DVSS.n10454 2.2505
R33419 DVSS.n10454 DVSS.n2009 2.2505
R33420 DVSS.n10453 DVSS.n10452 2.2505
R33421 DVSS.n10450 DVSS.n10449 2.2505
R33422 DVSS.n10447 DVSS.n10173 2.2505
R33423 DVSS.n10443 DVSS.n10442 2.2505
R33424 DVSS.n10440 DVSS.n10439 2.2505
R33425 DVSS.n10438 DVSS.n10437 2.2505
R33426 DVSS.n10435 DVSS.n10175 2.2505
R33427 DVSS.n10431 DVSS.n10430 2.2505
R33428 DVSS.n10428 DVSS.n10427 2.2505
R33429 DVSS.n10426 DVSS.n10425 2.2505
R33430 DVSS.n10423 DVSS.n10177 2.2505
R33431 DVSS.n10419 DVSS.n10418 2.2505
R33432 DVSS.n10416 DVSS.n10415 2.2505
R33433 DVSS.n10414 DVSS.n10413 2.2505
R33434 DVSS.n10411 DVSS.n10179 2.2505
R33435 DVSS.n10407 DVSS.n10406 2.2505
R33436 DVSS.n10404 DVSS.n10403 2.2505
R33437 DVSS.n10402 DVSS.n10401 2.2505
R33438 DVSS.n10399 DVSS.n10181 2.2505
R33439 DVSS.n10395 DVSS.n10394 2.2505
R33440 DVSS.n10392 DVSS.n10391 2.2505
R33441 DVSS.n10390 DVSS.n10389 2.2505
R33442 DVSS.n10387 DVSS.n10183 2.2505
R33443 DVSS.n10383 DVSS.n10382 2.2505
R33444 DVSS.n10380 DVSS.n10379 2.2505
R33445 DVSS.n10378 DVSS.n10377 2.2505
R33446 DVSS.n10375 DVSS.n10185 2.2505
R33447 DVSS.n10371 DVSS.n10370 2.2505
R33448 DVSS.n10368 DVSS.n10367 2.2505
R33449 DVSS.n10366 DVSS.n10365 2.2505
R33450 DVSS.n10363 DVSS.n10187 2.2505
R33451 DVSS.n10359 DVSS.n10358 2.2505
R33452 DVSS.n10356 DVSS.n10355 2.2505
R33453 DVSS.n10354 DVSS.n10353 2.2505
R33454 DVSS.n10351 DVSS.n10189 2.2505
R33455 DVSS.n10347 DVSS.n10346 2.2505
R33456 DVSS.n10344 DVSS.n10343 2.2505
R33457 DVSS.n10342 DVSS.n10341 2.2505
R33458 DVSS.n10339 DVSS.n10191 2.2505
R33459 DVSS.n10335 DVSS.n10334 2.2505
R33460 DVSS.n10332 DVSS.n10331 2.2505
R33461 DVSS.n10330 DVSS.n10329 2.2505
R33462 DVSS.n10327 DVSS.n10193 2.2505
R33463 DVSS.n10323 DVSS.n10322 2.2505
R33464 DVSS.n10320 DVSS.n10319 2.2505
R33465 DVSS.n10318 DVSS.n10317 2.2505
R33466 DVSS.n10315 DVSS.n10195 2.2505
R33467 DVSS.n10311 DVSS.n10310 2.2505
R33468 DVSS.n10308 DVSS.n10307 2.2505
R33469 DVSS.n10306 DVSS.n10305 2.2505
R33470 DVSS.n10303 DVSS.n10197 2.2505
R33471 DVSS.n10299 DVSS.n10298 2.2505
R33472 DVSS.n10296 DVSS.n10295 2.2505
R33473 DVSS.n10294 DVSS.n10293 2.2505
R33474 DVSS.n10291 DVSS.n10199 2.2505
R33475 DVSS.n10287 DVSS.n10286 2.2505
R33476 DVSS.n10284 DVSS.n10283 2.2505
R33477 DVSS.n10282 DVSS.n10281 2.2505
R33478 DVSS.n10279 DVSS.n10201 2.2505
R33479 DVSS.n10275 DVSS.n10274 2.2505
R33480 DVSS.n10272 DVSS.n10271 2.2505
R33481 DVSS.n10270 DVSS.n10269 2.2505
R33482 DVSS.n10267 DVSS.n10203 2.2505
R33483 DVSS.n10263 DVSS.n10262 2.2505
R33484 DVSS.n10260 DVSS.n10259 2.2505
R33485 DVSS.n10258 DVSS.n10257 2.2505
R33486 DVSS.n10255 DVSS.n10205 2.2505
R33487 DVSS.n10251 DVSS.n10250 2.2505
R33488 DVSS.n10248 DVSS.n10247 2.2505
R33489 DVSS.n10246 DVSS.n10245 2.2505
R33490 DVSS.n10243 DVSS.n10207 2.2505
R33491 DVSS.n10239 DVSS.n10238 2.2505
R33492 DVSS.n10236 DVSS.n10235 2.2505
R33493 DVSS.n10234 DVSS.n10233 2.2505
R33494 DVSS.n10231 DVSS.n10209 2.2505
R33495 DVSS.n10227 DVSS.n10226 2.2505
R33496 DVSS.n10224 DVSS.n10223 2.2505
R33497 DVSS.n10222 DVSS.n10221 2.2505
R33498 DVSS.n10219 DVSS.n10211 2.2505
R33499 DVSS.n10215 DVSS.n10214 2.2505
R33500 DVSS.n10212 DVSS.n2014 2.2505
R33501 DVSS.n10472 DVSS.n10471 2.2505
R33502 DVSS.n10474 DVSS.n2011 2.2505
R33503 DVSS.n1713 DVSS.n1623 2.2505
R33504 DVSS.n1715 DVSS.n1714 2.2505
R33505 DVSS.n1720 DVSS.n1716 2.2505
R33506 DVSS.n1721 DVSS.n1711 2.2505
R33507 DVSS.n1726 DVSS.n1725 2.2505
R33508 DVSS.n1727 DVSS.n1710 2.2505
R33509 DVSS.n1732 DVSS.n1728 2.2505
R33510 DVSS.n1733 DVSS.n1709 2.2505
R33511 DVSS.n1738 DVSS.n1737 2.2505
R33512 DVSS.n1739 DVSS.n1708 2.2505
R33513 DVSS.n1744 DVSS.n1740 2.2505
R33514 DVSS.n1745 DVSS.n1707 2.2505
R33515 DVSS.n1750 DVSS.n1749 2.2505
R33516 DVSS.n1751 DVSS.n1706 2.2505
R33517 DVSS.n1756 DVSS.n1752 2.2505
R33518 DVSS.n1757 DVSS.n1705 2.2505
R33519 DVSS.n1762 DVSS.n1761 2.2505
R33520 DVSS.n1763 DVSS.n1704 2.2505
R33521 DVSS.n1768 DVSS.n1764 2.2505
R33522 DVSS.n1769 DVSS.n1703 2.2505
R33523 DVSS.n1774 DVSS.n1773 2.2505
R33524 DVSS.n1775 DVSS.n1702 2.2505
R33525 DVSS.n1780 DVSS.n1776 2.2505
R33526 DVSS.n1781 DVSS.n1701 2.2505
R33527 DVSS.n1786 DVSS.n1785 2.2505
R33528 DVSS.n1787 DVSS.n1700 2.2505
R33529 DVSS.n1792 DVSS.n1788 2.2505
R33530 DVSS.n1793 DVSS.n1699 2.2505
R33531 DVSS.n1798 DVSS.n1797 2.2505
R33532 DVSS.n1799 DVSS.n1698 2.2505
R33533 DVSS.n1804 DVSS.n1800 2.2505
R33534 DVSS.n1805 DVSS.n1697 2.2505
R33535 DVSS.n1810 DVSS.n1809 2.2505
R33536 DVSS.n1811 DVSS.n1696 2.2505
R33537 DVSS.n1816 DVSS.n1812 2.2505
R33538 DVSS.n1817 DVSS.n1695 2.2505
R33539 DVSS.n1822 DVSS.n1821 2.2505
R33540 DVSS.n1823 DVSS.n1694 2.2505
R33541 DVSS.n1828 DVSS.n1824 2.2505
R33542 DVSS.n1829 DVSS.n1693 2.2505
R33543 DVSS.n1834 DVSS.n1833 2.2505
R33544 DVSS.n1835 DVSS.n1692 2.2505
R33545 DVSS.n1840 DVSS.n1836 2.2505
R33546 DVSS.n1841 DVSS.n1691 2.2505
R33547 DVSS.n1846 DVSS.n1845 2.2505
R33548 DVSS.n1847 DVSS.n1690 2.2505
R33549 DVSS.n1852 DVSS.n1848 2.2505
R33550 DVSS.n1853 DVSS.n1689 2.2505
R33551 DVSS.n1858 DVSS.n1857 2.2505
R33552 DVSS.n1859 DVSS.n1688 2.2505
R33553 DVSS.n1864 DVSS.n1860 2.2505
R33554 DVSS.n1865 DVSS.n1687 2.2505
R33555 DVSS.n1870 DVSS.n1869 2.2505
R33556 DVSS.n1871 DVSS.n1686 2.2505
R33557 DVSS.n1876 DVSS.n1872 2.2505
R33558 DVSS.n1877 DVSS.n1685 2.2505
R33559 DVSS.n1882 DVSS.n1881 2.2505
R33560 DVSS.n1883 DVSS.n1684 2.2505
R33561 DVSS.n1888 DVSS.n1884 2.2505
R33562 DVSS.n1889 DVSS.n1683 2.2505
R33563 DVSS.n1894 DVSS.n1893 2.2505
R33564 DVSS.n1895 DVSS.n1682 2.2505
R33565 DVSS.n1900 DVSS.n1896 2.2505
R33566 DVSS.n1901 DVSS.n1681 2.2505
R33567 DVSS.n1906 DVSS.n1905 2.2505
R33568 DVSS.n1907 DVSS.n1680 2.2505
R33569 DVSS.n1912 DVSS.n1908 2.2505
R33570 DVSS.n1913 DVSS.n1679 2.2505
R33571 DVSS.n1918 DVSS.n1917 2.2505
R33572 DVSS.n1919 DVSS.n1678 2.2505
R33573 DVSS.n1924 DVSS.n1920 2.2505
R33574 DVSS.n1925 DVSS.n1677 2.2505
R33575 DVSS.n1930 DVSS.n1929 2.2505
R33576 DVSS.n1931 DVSS.n1676 2.2505
R33577 DVSS.n1936 DVSS.n1932 2.2505
R33578 DVSS.n1937 DVSS.n1675 2.2505
R33579 DVSS.n1942 DVSS.n1941 2.2505
R33580 DVSS.n1943 DVSS.n1674 2.2505
R33581 DVSS.n1948 DVSS.n1944 2.2505
R33582 DVSS.n1949 DVSS.n1673 2.2505
R33583 DVSS.n1954 DVSS.n1953 2.2505
R33584 DVSS.n1955 DVSS.n1672 2.2505
R33585 DVSS.n1957 DVSS.n1956 2.2505
R33586 DVSS.n1958 DVSS.n1669 2.2505
R33587 DVSS.n1959 DVSS.n1958 2.2505
R33588 DVSS.n1957 DVSS.n1668 2.2505
R33589 DVSS.n1672 DVSS.n1671 2.2505
R33590 DVSS.n1953 DVSS.n1952 2.2505
R33591 DVSS.n1950 DVSS.n1949 2.2505
R33592 DVSS.n1948 DVSS.n1947 2.2505
R33593 DVSS.n1945 DVSS.n1674 2.2505
R33594 DVSS.n1941 DVSS.n1940 2.2505
R33595 DVSS.n1938 DVSS.n1937 2.2505
R33596 DVSS.n1936 DVSS.n1935 2.2505
R33597 DVSS.n1933 DVSS.n1676 2.2505
R33598 DVSS.n1929 DVSS.n1928 2.2505
R33599 DVSS.n1926 DVSS.n1925 2.2505
R33600 DVSS.n1924 DVSS.n1923 2.2505
R33601 DVSS.n1921 DVSS.n1678 2.2505
R33602 DVSS.n1917 DVSS.n1916 2.2505
R33603 DVSS.n1914 DVSS.n1913 2.2505
R33604 DVSS.n1912 DVSS.n1911 2.2505
R33605 DVSS.n1909 DVSS.n1680 2.2505
R33606 DVSS.n1905 DVSS.n1904 2.2505
R33607 DVSS.n1902 DVSS.n1901 2.2505
R33608 DVSS.n1900 DVSS.n1899 2.2505
R33609 DVSS.n1897 DVSS.n1682 2.2505
R33610 DVSS.n1893 DVSS.n1892 2.2505
R33611 DVSS.n1890 DVSS.n1889 2.2505
R33612 DVSS.n1888 DVSS.n1887 2.2505
R33613 DVSS.n1885 DVSS.n1684 2.2505
R33614 DVSS.n1881 DVSS.n1880 2.2505
R33615 DVSS.n1878 DVSS.n1877 2.2505
R33616 DVSS.n1876 DVSS.n1875 2.2505
R33617 DVSS.n1873 DVSS.n1686 2.2505
R33618 DVSS.n1869 DVSS.n1868 2.2505
R33619 DVSS.n1866 DVSS.n1865 2.2505
R33620 DVSS.n1864 DVSS.n1863 2.2505
R33621 DVSS.n1861 DVSS.n1688 2.2505
R33622 DVSS.n1857 DVSS.n1856 2.2505
R33623 DVSS.n1854 DVSS.n1853 2.2505
R33624 DVSS.n1852 DVSS.n1851 2.2505
R33625 DVSS.n1849 DVSS.n1690 2.2505
R33626 DVSS.n1845 DVSS.n1844 2.2505
R33627 DVSS.n1842 DVSS.n1841 2.2505
R33628 DVSS.n1840 DVSS.n1839 2.2505
R33629 DVSS.n1837 DVSS.n1692 2.2505
R33630 DVSS.n1833 DVSS.n1832 2.2505
R33631 DVSS.n1830 DVSS.n1829 2.2505
R33632 DVSS.n1828 DVSS.n1827 2.2505
R33633 DVSS.n1825 DVSS.n1694 2.2505
R33634 DVSS.n1821 DVSS.n1820 2.2505
R33635 DVSS.n1818 DVSS.n1817 2.2505
R33636 DVSS.n1816 DVSS.n1815 2.2505
R33637 DVSS.n1813 DVSS.n1696 2.2505
R33638 DVSS.n1809 DVSS.n1808 2.2505
R33639 DVSS.n1806 DVSS.n1805 2.2505
R33640 DVSS.n1804 DVSS.n1803 2.2505
R33641 DVSS.n1801 DVSS.n1698 2.2505
R33642 DVSS.n1797 DVSS.n1796 2.2505
R33643 DVSS.n1794 DVSS.n1793 2.2505
R33644 DVSS.n1792 DVSS.n1791 2.2505
R33645 DVSS.n1789 DVSS.n1700 2.2505
R33646 DVSS.n1785 DVSS.n1784 2.2505
R33647 DVSS.n1782 DVSS.n1781 2.2505
R33648 DVSS.n1780 DVSS.n1779 2.2505
R33649 DVSS.n1777 DVSS.n1702 2.2505
R33650 DVSS.n1773 DVSS.n1772 2.2505
R33651 DVSS.n1770 DVSS.n1769 2.2505
R33652 DVSS.n1768 DVSS.n1767 2.2505
R33653 DVSS.n1765 DVSS.n1704 2.2505
R33654 DVSS.n1761 DVSS.n1760 2.2505
R33655 DVSS.n1758 DVSS.n1757 2.2505
R33656 DVSS.n1756 DVSS.n1755 2.2505
R33657 DVSS.n1753 DVSS.n1706 2.2505
R33658 DVSS.n1749 DVSS.n1748 2.2505
R33659 DVSS.n1746 DVSS.n1745 2.2505
R33660 DVSS.n1744 DVSS.n1743 2.2505
R33661 DVSS.n1741 DVSS.n1708 2.2505
R33662 DVSS.n1737 DVSS.n1736 2.2505
R33663 DVSS.n1734 DVSS.n1733 2.2505
R33664 DVSS.n1732 DVSS.n1731 2.2505
R33665 DVSS.n1729 DVSS.n1710 2.2505
R33666 DVSS.n1725 DVSS.n1724 2.2505
R33667 DVSS.n1722 DVSS.n1721 2.2505
R33668 DVSS.n1720 DVSS.n1719 2.2505
R33669 DVSS.n1717 DVSS.n1714 2.2505
R33670 DVSS.n1713 DVSS.n1712 2.2505
R33671 DVSS.n1567 DVSS.n1517 2.2505
R33672 DVSS.n10750 DVSS.n10749 2.2505
R33673 DVSS.n10748 DVSS.n1569 2.2505
R33674 DVSS.n10747 DVSS.n10746 2.2505
R33675 DVSS.n10742 DVSS.n1570 2.2505
R33676 DVSS.n10738 DVSS.n10737 2.2505
R33677 DVSS.n10736 DVSS.n1571 2.2505
R33678 DVSS.n10735 DVSS.n10734 2.2505
R33679 DVSS.n10730 DVSS.n1572 2.2505
R33680 DVSS.n10726 DVSS.n10725 2.2505
R33681 DVSS.n10724 DVSS.n1573 2.2505
R33682 DVSS.n10723 DVSS.n10722 2.2505
R33683 DVSS.n10718 DVSS.n1574 2.2505
R33684 DVSS.n10714 DVSS.n10713 2.2505
R33685 DVSS.n10712 DVSS.n1575 2.2505
R33686 DVSS.n10711 DVSS.n10710 2.2505
R33687 DVSS.n10706 DVSS.n1576 2.2505
R33688 DVSS.n10702 DVSS.n10701 2.2505
R33689 DVSS.n10700 DVSS.n1577 2.2505
R33690 DVSS.n10699 DVSS.n10698 2.2505
R33691 DVSS.n10694 DVSS.n1578 2.2505
R33692 DVSS.n10690 DVSS.n10689 2.2505
R33693 DVSS.n10688 DVSS.n1579 2.2505
R33694 DVSS.n10687 DVSS.n10686 2.2505
R33695 DVSS.n10682 DVSS.n1580 2.2505
R33696 DVSS.n10678 DVSS.n10677 2.2505
R33697 DVSS.n10676 DVSS.n1581 2.2505
R33698 DVSS.n10675 DVSS.n10674 2.2505
R33699 DVSS.n10670 DVSS.n1582 2.2505
R33700 DVSS.n10666 DVSS.n10665 2.2505
R33701 DVSS.n10664 DVSS.n1583 2.2505
R33702 DVSS.n10663 DVSS.n10662 2.2505
R33703 DVSS.n10658 DVSS.n1584 2.2505
R33704 DVSS.n10654 DVSS.n10653 2.2505
R33705 DVSS.n10652 DVSS.n1585 2.2505
R33706 DVSS.n10651 DVSS.n10650 2.2505
R33707 DVSS.n10646 DVSS.n1586 2.2505
R33708 DVSS.n10642 DVSS.n10641 2.2505
R33709 DVSS.n10640 DVSS.n1587 2.2505
R33710 DVSS.n10639 DVSS.n10638 2.2505
R33711 DVSS.n10634 DVSS.n1588 2.2505
R33712 DVSS.n10630 DVSS.n10629 2.2505
R33713 DVSS.n10628 DVSS.n1589 2.2505
R33714 DVSS.n10627 DVSS.n10626 2.2505
R33715 DVSS.n10622 DVSS.n1590 2.2505
R33716 DVSS.n10618 DVSS.n10617 2.2505
R33717 DVSS.n10616 DVSS.n1591 2.2505
R33718 DVSS.n10615 DVSS.n10614 2.2505
R33719 DVSS.n10610 DVSS.n1592 2.2505
R33720 DVSS.n10606 DVSS.n10605 2.2505
R33721 DVSS.n10604 DVSS.n1593 2.2505
R33722 DVSS.n10603 DVSS.n10602 2.2505
R33723 DVSS.n10598 DVSS.n1594 2.2505
R33724 DVSS.n10594 DVSS.n10593 2.2505
R33725 DVSS.n10592 DVSS.n1595 2.2505
R33726 DVSS.n10591 DVSS.n10590 2.2505
R33727 DVSS.n10586 DVSS.n1596 2.2505
R33728 DVSS.n10582 DVSS.n10581 2.2505
R33729 DVSS.n10580 DVSS.n1597 2.2505
R33730 DVSS.n10579 DVSS.n10578 2.2505
R33731 DVSS.n10574 DVSS.n1598 2.2505
R33732 DVSS.n10570 DVSS.n10569 2.2505
R33733 DVSS.n10568 DVSS.n1599 2.2505
R33734 DVSS.n10567 DVSS.n10566 2.2505
R33735 DVSS.n10562 DVSS.n1600 2.2505
R33736 DVSS.n10558 DVSS.n10557 2.2505
R33737 DVSS.n10556 DVSS.n1601 2.2505
R33738 DVSS.n10555 DVSS.n10554 2.2505
R33739 DVSS.n10550 DVSS.n1602 2.2505
R33740 DVSS.n10546 DVSS.n10545 2.2505
R33741 DVSS.n10544 DVSS.n1603 2.2505
R33742 DVSS.n10543 DVSS.n10542 2.2505
R33743 DVSS.n10538 DVSS.n1604 2.2505
R33744 DVSS.n10534 DVSS.n10533 2.2505
R33745 DVSS.n10532 DVSS.n1605 2.2505
R33746 DVSS.n10531 DVSS.n10530 2.2505
R33747 DVSS.n10526 DVSS.n1606 2.2505
R33748 DVSS.n10522 DVSS.n10521 2.2505
R33749 DVSS.n10520 DVSS.n1607 2.2505
R33750 DVSS.n10519 DVSS.n10518 2.2505
R33751 DVSS.n10514 DVSS.n1608 2.2505
R33752 DVSS.n10510 DVSS.n10509 2.2505
R33753 DVSS.n10508 DVSS.n1611 2.2505
R33754 DVSS.n10507 DVSS.n10506 2.2505
R33755 DVSS.n10506 DVSS.n1565 2.2505
R33756 DVSS.n1611 DVSS.n1610 2.2505
R33757 DVSS.n10511 DVSS.n10510 2.2505
R33758 DVSS.n10514 DVSS.n10513 2.2505
R33759 DVSS.n10518 DVSS.n10517 2.2505
R33760 DVSS.n10515 DVSS.n1607 2.2505
R33761 DVSS.n10523 DVSS.n10522 2.2505
R33762 DVSS.n10526 DVSS.n10525 2.2505
R33763 DVSS.n10530 DVSS.n10529 2.2505
R33764 DVSS.n10527 DVSS.n1605 2.2505
R33765 DVSS.n10535 DVSS.n10534 2.2505
R33766 DVSS.n10538 DVSS.n10537 2.2505
R33767 DVSS.n10542 DVSS.n10541 2.2505
R33768 DVSS.n10539 DVSS.n1603 2.2505
R33769 DVSS.n10547 DVSS.n10546 2.2505
R33770 DVSS.n10550 DVSS.n10549 2.2505
R33771 DVSS.n10554 DVSS.n10553 2.2505
R33772 DVSS.n10551 DVSS.n1601 2.2505
R33773 DVSS.n10559 DVSS.n10558 2.2505
R33774 DVSS.n10562 DVSS.n10561 2.2505
R33775 DVSS.n10566 DVSS.n10565 2.2505
R33776 DVSS.n10563 DVSS.n1599 2.2505
R33777 DVSS.n10571 DVSS.n10570 2.2505
R33778 DVSS.n10574 DVSS.n10573 2.2505
R33779 DVSS.n10578 DVSS.n10577 2.2505
R33780 DVSS.n10575 DVSS.n1597 2.2505
R33781 DVSS.n10583 DVSS.n10582 2.2505
R33782 DVSS.n10586 DVSS.n10585 2.2505
R33783 DVSS.n10590 DVSS.n10589 2.2505
R33784 DVSS.n10587 DVSS.n1595 2.2505
R33785 DVSS.n10595 DVSS.n10594 2.2505
R33786 DVSS.n10598 DVSS.n10597 2.2505
R33787 DVSS.n10602 DVSS.n10601 2.2505
R33788 DVSS.n10599 DVSS.n1593 2.2505
R33789 DVSS.n10607 DVSS.n10606 2.2505
R33790 DVSS.n10610 DVSS.n10609 2.2505
R33791 DVSS.n10614 DVSS.n10613 2.2505
R33792 DVSS.n10611 DVSS.n1591 2.2505
R33793 DVSS.n10619 DVSS.n10618 2.2505
R33794 DVSS.n10622 DVSS.n10621 2.2505
R33795 DVSS.n10626 DVSS.n10625 2.2505
R33796 DVSS.n10623 DVSS.n1589 2.2505
R33797 DVSS.n10631 DVSS.n10630 2.2505
R33798 DVSS.n10634 DVSS.n10633 2.2505
R33799 DVSS.n10638 DVSS.n10637 2.2505
R33800 DVSS.n10635 DVSS.n1587 2.2505
R33801 DVSS.n10643 DVSS.n10642 2.2505
R33802 DVSS.n10646 DVSS.n10645 2.2505
R33803 DVSS.n10650 DVSS.n10649 2.2505
R33804 DVSS.n10647 DVSS.n1585 2.2505
R33805 DVSS.n10655 DVSS.n10654 2.2505
R33806 DVSS.n10658 DVSS.n10657 2.2505
R33807 DVSS.n10662 DVSS.n10661 2.2505
R33808 DVSS.n10659 DVSS.n1583 2.2505
R33809 DVSS.n10667 DVSS.n10666 2.2505
R33810 DVSS.n10670 DVSS.n10669 2.2505
R33811 DVSS.n10674 DVSS.n10673 2.2505
R33812 DVSS.n10671 DVSS.n1581 2.2505
R33813 DVSS.n10679 DVSS.n10678 2.2505
R33814 DVSS.n10682 DVSS.n10681 2.2505
R33815 DVSS.n10686 DVSS.n10685 2.2505
R33816 DVSS.n10683 DVSS.n1579 2.2505
R33817 DVSS.n10691 DVSS.n10690 2.2505
R33818 DVSS.n10694 DVSS.n10693 2.2505
R33819 DVSS.n10698 DVSS.n10697 2.2505
R33820 DVSS.n10695 DVSS.n1577 2.2505
R33821 DVSS.n10703 DVSS.n10702 2.2505
R33822 DVSS.n10706 DVSS.n10705 2.2505
R33823 DVSS.n10710 DVSS.n10709 2.2505
R33824 DVSS.n10707 DVSS.n1575 2.2505
R33825 DVSS.n10715 DVSS.n10714 2.2505
R33826 DVSS.n10718 DVSS.n10717 2.2505
R33827 DVSS.n10722 DVSS.n10721 2.2505
R33828 DVSS.n10719 DVSS.n1573 2.2505
R33829 DVSS.n10727 DVSS.n10726 2.2505
R33830 DVSS.n10730 DVSS.n10729 2.2505
R33831 DVSS.n10734 DVSS.n10733 2.2505
R33832 DVSS.n10731 DVSS.n1571 2.2505
R33833 DVSS.n10739 DVSS.n10738 2.2505
R33834 DVSS.n10742 DVSS.n10741 2.2505
R33835 DVSS.n10746 DVSS.n10745 2.2505
R33836 DVSS.n10743 DVSS.n1569 2.2505
R33837 DVSS.n10751 DVSS.n10750 2.2505
R33838 DVSS.n10753 DVSS.n1567 2.2505
R33839 DVSS.n10895 DVSS.n10761 2.2505
R33840 DVSS.n10897 DVSS.n10896 2.2505
R33841 DVSS.n10890 DVSS.n10889 2.2505
R33842 DVSS.n10904 DVSS.n10903 2.2505
R33843 DVSS.n10905 DVSS.n10888 2.2505
R33844 DVSS.n10907 DVSS.n10906 2.2505
R33845 DVSS.n10884 DVSS.n10883 2.2505
R33846 DVSS.n10914 DVSS.n10913 2.2505
R33847 DVSS.n10915 DVSS.n10882 2.2505
R33848 DVSS.n10917 DVSS.n10916 2.2505
R33849 DVSS.n10878 DVSS.n10877 2.2505
R33850 DVSS.n10924 DVSS.n10923 2.2505
R33851 DVSS.n10925 DVSS.n10876 2.2505
R33852 DVSS.n10927 DVSS.n10926 2.2505
R33853 DVSS.n10872 DVSS.n10871 2.2505
R33854 DVSS.n10934 DVSS.n10933 2.2505
R33855 DVSS.n10935 DVSS.n10870 2.2505
R33856 DVSS.n10937 DVSS.n10936 2.2505
R33857 DVSS.n10866 DVSS.n10865 2.2505
R33858 DVSS.n10944 DVSS.n10943 2.2505
R33859 DVSS.n10945 DVSS.n10864 2.2505
R33860 DVSS.n10947 DVSS.n10946 2.2505
R33861 DVSS.n10860 DVSS.n10859 2.2505
R33862 DVSS.n10954 DVSS.n10953 2.2505
R33863 DVSS.n10955 DVSS.n10858 2.2505
R33864 DVSS.n10957 DVSS.n10956 2.2505
R33865 DVSS.n10854 DVSS.n10853 2.2505
R33866 DVSS.n10964 DVSS.n10963 2.2505
R33867 DVSS.n10965 DVSS.n10852 2.2505
R33868 DVSS.n10967 DVSS.n10966 2.2505
R33869 DVSS.n10848 DVSS.n10847 2.2505
R33870 DVSS.n10974 DVSS.n10973 2.2505
R33871 DVSS.n10975 DVSS.n10846 2.2505
R33872 DVSS.n10977 DVSS.n10976 2.2505
R33873 DVSS.n10842 DVSS.n10841 2.2505
R33874 DVSS.n10984 DVSS.n10983 2.2505
R33875 DVSS.n10985 DVSS.n10840 2.2505
R33876 DVSS.n10987 DVSS.n10986 2.2505
R33877 DVSS.n10836 DVSS.n10835 2.2505
R33878 DVSS.n10994 DVSS.n10993 2.2505
R33879 DVSS.n10995 DVSS.n10834 2.2505
R33880 DVSS.n10997 DVSS.n10996 2.2505
R33881 DVSS.n10830 DVSS.n10829 2.2505
R33882 DVSS.n11004 DVSS.n11003 2.2505
R33883 DVSS.n11005 DVSS.n10828 2.2505
R33884 DVSS.n11007 DVSS.n11006 2.2505
R33885 DVSS.n10824 DVSS.n10823 2.2505
R33886 DVSS.n11014 DVSS.n11013 2.2505
R33887 DVSS.n11015 DVSS.n10822 2.2505
R33888 DVSS.n11017 DVSS.n11016 2.2505
R33889 DVSS.n10818 DVSS.n10817 2.2505
R33890 DVSS.n11024 DVSS.n11023 2.2505
R33891 DVSS.n11025 DVSS.n10816 2.2505
R33892 DVSS.n11027 DVSS.n11026 2.2505
R33893 DVSS.n10812 DVSS.n10811 2.2505
R33894 DVSS.n11034 DVSS.n11033 2.2505
R33895 DVSS.n11035 DVSS.n10810 2.2505
R33896 DVSS.n11037 DVSS.n11036 2.2505
R33897 DVSS.n10806 DVSS.n10805 2.2505
R33898 DVSS.n11044 DVSS.n11043 2.2505
R33899 DVSS.n11045 DVSS.n10804 2.2505
R33900 DVSS.n11047 DVSS.n11046 2.2505
R33901 DVSS.n10800 DVSS.n10799 2.2505
R33902 DVSS.n11054 DVSS.n11053 2.2505
R33903 DVSS.n11055 DVSS.n10798 2.2505
R33904 DVSS.n11057 DVSS.n11056 2.2505
R33905 DVSS.n10794 DVSS.n10793 2.2505
R33906 DVSS.n11064 DVSS.n11063 2.2505
R33907 DVSS.n11065 DVSS.n10792 2.2505
R33908 DVSS.n11067 DVSS.n11066 2.2505
R33909 DVSS.n10788 DVSS.n10787 2.2505
R33910 DVSS.n11074 DVSS.n11073 2.2505
R33911 DVSS.n11075 DVSS.n10786 2.2505
R33912 DVSS.n11077 DVSS.n11076 2.2505
R33913 DVSS.n10782 DVSS.n10781 2.2505
R33914 DVSS.n11084 DVSS.n11083 2.2505
R33915 DVSS.n11085 DVSS.n10780 2.2505
R33916 DVSS.n11087 DVSS.n11086 2.2505
R33917 DVSS.n10776 DVSS.n10775 2.2505
R33918 DVSS.n11094 DVSS.n11093 2.2505
R33919 DVSS.n11095 DVSS.n10774 2.2505
R33920 DVSS.n11097 DVSS.n11096 2.2505
R33921 DVSS.n10772 DVSS.n10771 2.2505
R33922 DVSS.n11104 DVSS.n11103 2.2505
R33923 DVSS.n11103 DVSS.n11102 2.2505
R33924 DVSS.n11100 DVSS.n10772 2.2505
R33925 DVSS.n11098 DVSS.n11097 2.2505
R33926 DVSS.n10777 DVSS.n10774 2.2505
R33927 DVSS.n11093 DVSS.n11092 2.2505
R33928 DVSS.n11090 DVSS.n10776 2.2505
R33929 DVSS.n11088 DVSS.n11087 2.2505
R33930 DVSS.n10783 DVSS.n10780 2.2505
R33931 DVSS.n11083 DVSS.n11082 2.2505
R33932 DVSS.n11080 DVSS.n10782 2.2505
R33933 DVSS.n11078 DVSS.n11077 2.2505
R33934 DVSS.n10789 DVSS.n10786 2.2505
R33935 DVSS.n11073 DVSS.n11072 2.2505
R33936 DVSS.n11070 DVSS.n10788 2.2505
R33937 DVSS.n11068 DVSS.n11067 2.2505
R33938 DVSS.n10795 DVSS.n10792 2.2505
R33939 DVSS.n11063 DVSS.n11062 2.2505
R33940 DVSS.n11060 DVSS.n10794 2.2505
R33941 DVSS.n11058 DVSS.n11057 2.2505
R33942 DVSS.n10801 DVSS.n10798 2.2505
R33943 DVSS.n11053 DVSS.n11052 2.2505
R33944 DVSS.n11050 DVSS.n10800 2.2505
R33945 DVSS.n11048 DVSS.n11047 2.2505
R33946 DVSS.n10807 DVSS.n10804 2.2505
R33947 DVSS.n11043 DVSS.n11042 2.2505
R33948 DVSS.n11040 DVSS.n10806 2.2505
R33949 DVSS.n11038 DVSS.n11037 2.2505
R33950 DVSS.n10813 DVSS.n10810 2.2505
R33951 DVSS.n11033 DVSS.n11032 2.2505
R33952 DVSS.n11030 DVSS.n10812 2.2505
R33953 DVSS.n11028 DVSS.n11027 2.2505
R33954 DVSS.n10819 DVSS.n10816 2.2505
R33955 DVSS.n11023 DVSS.n11022 2.2505
R33956 DVSS.n11020 DVSS.n10818 2.2505
R33957 DVSS.n11018 DVSS.n11017 2.2505
R33958 DVSS.n10825 DVSS.n10822 2.2505
R33959 DVSS.n11013 DVSS.n11012 2.2505
R33960 DVSS.n11010 DVSS.n10824 2.2505
R33961 DVSS.n11008 DVSS.n11007 2.2505
R33962 DVSS.n10831 DVSS.n10828 2.2505
R33963 DVSS.n11003 DVSS.n11002 2.2505
R33964 DVSS.n11000 DVSS.n10830 2.2505
R33965 DVSS.n10998 DVSS.n10997 2.2505
R33966 DVSS.n10837 DVSS.n10834 2.2505
R33967 DVSS.n10993 DVSS.n10992 2.2505
R33968 DVSS.n10990 DVSS.n10836 2.2505
R33969 DVSS.n10988 DVSS.n10987 2.2505
R33970 DVSS.n10843 DVSS.n10840 2.2505
R33971 DVSS.n10983 DVSS.n10982 2.2505
R33972 DVSS.n10980 DVSS.n10842 2.2505
R33973 DVSS.n10978 DVSS.n10977 2.2505
R33974 DVSS.n10849 DVSS.n10846 2.2505
R33975 DVSS.n10973 DVSS.n10972 2.2505
R33976 DVSS.n10970 DVSS.n10848 2.2505
R33977 DVSS.n10968 DVSS.n10967 2.2505
R33978 DVSS.n10855 DVSS.n10852 2.2505
R33979 DVSS.n10963 DVSS.n10962 2.2505
R33980 DVSS.n10960 DVSS.n10854 2.2505
R33981 DVSS.n10958 DVSS.n10957 2.2505
R33982 DVSS.n10861 DVSS.n10858 2.2505
R33983 DVSS.n10953 DVSS.n10952 2.2505
R33984 DVSS.n10950 DVSS.n10860 2.2505
R33985 DVSS.n10948 DVSS.n10947 2.2505
R33986 DVSS.n10867 DVSS.n10864 2.2505
R33987 DVSS.n10943 DVSS.n10942 2.2505
R33988 DVSS.n10940 DVSS.n10866 2.2505
R33989 DVSS.n10938 DVSS.n10937 2.2505
R33990 DVSS.n10873 DVSS.n10870 2.2505
R33991 DVSS.n10933 DVSS.n10932 2.2505
R33992 DVSS.n10930 DVSS.n10872 2.2505
R33993 DVSS.n10928 DVSS.n10927 2.2505
R33994 DVSS.n10879 DVSS.n10876 2.2505
R33995 DVSS.n10923 DVSS.n10922 2.2505
R33996 DVSS.n10920 DVSS.n10878 2.2505
R33997 DVSS.n10918 DVSS.n10917 2.2505
R33998 DVSS.n10885 DVSS.n10882 2.2505
R33999 DVSS.n10913 DVSS.n10912 2.2505
R34000 DVSS.n10910 DVSS.n10884 2.2505
R34001 DVSS.n10908 DVSS.n10907 2.2505
R34002 DVSS.n10891 DVSS.n10888 2.2505
R34003 DVSS.n10903 DVSS.n10902 2.2505
R34004 DVSS.n10900 DVSS.n10890 2.2505
R34005 DVSS.n10898 DVSS.n10897 2.2505
R34006 DVSS.n10895 DVSS.n10894 2.2505
R34007 DVSS.n13335 DVSS.n11446 2.2505
R34008 DVSS.n11445 DVSS.n11201 2.2505
R34009 DVSS.n11444 DVSS.n11443 2.2505
R34010 DVSS.n11441 DVSS.n11202 2.2505
R34011 DVSS.n11439 DVSS.n11437 2.2505
R34012 DVSS.n11436 DVSS.n11204 2.2505
R34013 DVSS.n11435 DVSS.n11434 2.2505
R34014 DVSS.n11432 DVSS.n11205 2.2505
R34015 DVSS.n11430 DVSS.n11428 2.2505
R34016 DVSS.n11427 DVSS.n11207 2.2505
R34017 DVSS.n11426 DVSS.n11425 2.2505
R34018 DVSS.n11423 DVSS.n11208 2.2505
R34019 DVSS.n11421 DVSS.n11419 2.2505
R34020 DVSS.n11418 DVSS.n11210 2.2505
R34021 DVSS.n11417 DVSS.n11416 2.2505
R34022 DVSS.n11414 DVSS.n11211 2.2505
R34023 DVSS.n11412 DVSS.n11410 2.2505
R34024 DVSS.n11409 DVSS.n11213 2.2505
R34025 DVSS.n11408 DVSS.n11407 2.2505
R34026 DVSS.n11405 DVSS.n11214 2.2505
R34027 DVSS.n11403 DVSS.n11401 2.2505
R34028 DVSS.n11400 DVSS.n11216 2.2505
R34029 DVSS.n11399 DVSS.n11398 2.2505
R34030 DVSS.n11396 DVSS.n11217 2.2505
R34031 DVSS.n11394 DVSS.n11392 2.2505
R34032 DVSS.n11391 DVSS.n11219 2.2505
R34033 DVSS.n11390 DVSS.n11389 2.2505
R34034 DVSS.n11387 DVSS.n11220 2.2505
R34035 DVSS.n11385 DVSS.n11383 2.2505
R34036 DVSS.n11382 DVSS.n11222 2.2505
R34037 DVSS.n11381 DVSS.n11380 2.2505
R34038 DVSS.n11378 DVSS.n11223 2.2505
R34039 DVSS.n11376 DVSS.n11374 2.2505
R34040 DVSS.n11373 DVSS.n11225 2.2505
R34041 DVSS.n11372 DVSS.n11371 2.2505
R34042 DVSS.n11369 DVSS.n11226 2.2505
R34043 DVSS.n11367 DVSS.n11365 2.2505
R34044 DVSS.n11364 DVSS.n11228 2.2505
R34045 DVSS.n11363 DVSS.n11362 2.2505
R34046 DVSS.n11360 DVSS.n11229 2.2505
R34047 DVSS.n11358 DVSS.n11356 2.2505
R34048 DVSS.n11355 DVSS.n11231 2.2505
R34049 DVSS.n11354 DVSS.n11353 2.2505
R34050 DVSS.n11351 DVSS.n11232 2.2505
R34051 DVSS.n11349 DVSS.n11347 2.2505
R34052 DVSS.n11346 DVSS.n11234 2.2505
R34053 DVSS.n11345 DVSS.n11344 2.2505
R34054 DVSS.n11342 DVSS.n11235 2.2505
R34055 DVSS.n11340 DVSS.n11338 2.2505
R34056 DVSS.n11337 DVSS.n11237 2.2505
R34057 DVSS.n11336 DVSS.n11335 2.2505
R34058 DVSS.n11333 DVSS.n11238 2.2505
R34059 DVSS.n11331 DVSS.n11329 2.2505
R34060 DVSS.n11328 DVSS.n11240 2.2505
R34061 DVSS.n11327 DVSS.n11326 2.2505
R34062 DVSS.n11324 DVSS.n11241 2.2505
R34063 DVSS.n11322 DVSS.n11320 2.2505
R34064 DVSS.n11319 DVSS.n11243 2.2505
R34065 DVSS.n11318 DVSS.n11317 2.2505
R34066 DVSS.n11315 DVSS.n11244 2.2505
R34067 DVSS.n11313 DVSS.n11311 2.2505
R34068 DVSS.n11310 DVSS.n11246 2.2505
R34069 DVSS.n11309 DVSS.n11308 2.2505
R34070 DVSS.n11306 DVSS.n11247 2.2505
R34071 DVSS.n11304 DVSS.n11302 2.2505
R34072 DVSS.n11301 DVSS.n11249 2.2505
R34073 DVSS.n11300 DVSS.n11299 2.2505
R34074 DVSS.n11297 DVSS.n11250 2.2505
R34075 DVSS.n11295 DVSS.n11293 2.2505
R34076 DVSS.n11292 DVSS.n11252 2.2505
R34077 DVSS.n11291 DVSS.n11290 2.2505
R34078 DVSS.n11288 DVSS.n11253 2.2505
R34079 DVSS.n11286 DVSS.n11284 2.2505
R34080 DVSS.n11283 DVSS.n11255 2.2505
R34081 DVSS.n11282 DVSS.n11281 2.2505
R34082 DVSS.n11279 DVSS.n11256 2.2505
R34083 DVSS.n11277 DVSS.n11275 2.2505
R34084 DVSS.n11274 DVSS.n11258 2.2505
R34085 DVSS.n11273 DVSS.n11272 2.2505
R34086 DVSS.n11270 DVSS.n11259 2.2505
R34087 DVSS.n11268 DVSS.n11266 2.2505
R34088 DVSS.n11265 DVSS.n11261 2.2505
R34089 DVSS.n11264 DVSS.n11263 2.2505
R34090 DVSS.n11262 DVSS.n11155 2.2505
R34091 DVSS.n13338 DVSS.n11155 2.2505
R34092 DVSS.n11263 DVSS.n11154 2.2505
R34093 DVSS.n11261 DVSS.n11260 2.2505
R34094 DVSS.n11268 DVSS.n11267 2.2505
R34095 DVSS.n11270 DVSS.n11269 2.2505
R34096 DVSS.n11272 DVSS.n11271 2.2505
R34097 DVSS.n11258 DVSS.n11257 2.2505
R34098 DVSS.n11277 DVSS.n11276 2.2505
R34099 DVSS.n11279 DVSS.n11278 2.2505
R34100 DVSS.n11281 DVSS.n11280 2.2505
R34101 DVSS.n11255 DVSS.n11254 2.2505
R34102 DVSS.n11286 DVSS.n11285 2.2505
R34103 DVSS.n11288 DVSS.n11287 2.2505
R34104 DVSS.n11290 DVSS.n11289 2.2505
R34105 DVSS.n11252 DVSS.n11251 2.2505
R34106 DVSS.n11295 DVSS.n11294 2.2505
R34107 DVSS.n11297 DVSS.n11296 2.2505
R34108 DVSS.n11299 DVSS.n11298 2.2505
R34109 DVSS.n11249 DVSS.n11248 2.2505
R34110 DVSS.n11304 DVSS.n11303 2.2505
R34111 DVSS.n11306 DVSS.n11305 2.2505
R34112 DVSS.n11308 DVSS.n11307 2.2505
R34113 DVSS.n11246 DVSS.n11245 2.2505
R34114 DVSS.n11313 DVSS.n11312 2.2505
R34115 DVSS.n11315 DVSS.n11314 2.2505
R34116 DVSS.n11317 DVSS.n11316 2.2505
R34117 DVSS.n11243 DVSS.n11242 2.2505
R34118 DVSS.n11322 DVSS.n11321 2.2505
R34119 DVSS.n11324 DVSS.n11323 2.2505
R34120 DVSS.n11326 DVSS.n11325 2.2505
R34121 DVSS.n11240 DVSS.n11239 2.2505
R34122 DVSS.n11331 DVSS.n11330 2.2505
R34123 DVSS.n11333 DVSS.n11332 2.2505
R34124 DVSS.n11335 DVSS.n11334 2.2505
R34125 DVSS.n11237 DVSS.n11236 2.2505
R34126 DVSS.n11340 DVSS.n11339 2.2505
R34127 DVSS.n11342 DVSS.n11341 2.2505
R34128 DVSS.n11344 DVSS.n11343 2.2505
R34129 DVSS.n11234 DVSS.n11233 2.2505
R34130 DVSS.n11349 DVSS.n11348 2.2505
R34131 DVSS.n11351 DVSS.n11350 2.2505
R34132 DVSS.n11353 DVSS.n11352 2.2505
R34133 DVSS.n11231 DVSS.n11230 2.2505
R34134 DVSS.n11358 DVSS.n11357 2.2505
R34135 DVSS.n11360 DVSS.n11359 2.2505
R34136 DVSS.n11362 DVSS.n11361 2.2505
R34137 DVSS.n11228 DVSS.n11227 2.2505
R34138 DVSS.n11367 DVSS.n11366 2.2505
R34139 DVSS.n11369 DVSS.n11368 2.2505
R34140 DVSS.n11371 DVSS.n11370 2.2505
R34141 DVSS.n11225 DVSS.n11224 2.2505
R34142 DVSS.n11376 DVSS.n11375 2.2505
R34143 DVSS.n11378 DVSS.n11377 2.2505
R34144 DVSS.n11380 DVSS.n11379 2.2505
R34145 DVSS.n11222 DVSS.n11221 2.2505
R34146 DVSS.n11385 DVSS.n11384 2.2505
R34147 DVSS.n11387 DVSS.n11386 2.2505
R34148 DVSS.n11389 DVSS.n11388 2.2505
R34149 DVSS.n11219 DVSS.n11218 2.2505
R34150 DVSS.n11394 DVSS.n11393 2.2505
R34151 DVSS.n11396 DVSS.n11395 2.2505
R34152 DVSS.n11398 DVSS.n11397 2.2505
R34153 DVSS.n11216 DVSS.n11215 2.2505
R34154 DVSS.n11403 DVSS.n11402 2.2505
R34155 DVSS.n11405 DVSS.n11404 2.2505
R34156 DVSS.n11407 DVSS.n11406 2.2505
R34157 DVSS.n11213 DVSS.n11212 2.2505
R34158 DVSS.n11412 DVSS.n11411 2.2505
R34159 DVSS.n11414 DVSS.n11413 2.2505
R34160 DVSS.n11416 DVSS.n11415 2.2505
R34161 DVSS.n11210 DVSS.n11209 2.2505
R34162 DVSS.n11421 DVSS.n11420 2.2505
R34163 DVSS.n11423 DVSS.n11422 2.2505
R34164 DVSS.n11425 DVSS.n11424 2.2505
R34165 DVSS.n11207 DVSS.n11206 2.2505
R34166 DVSS.n11430 DVSS.n11429 2.2505
R34167 DVSS.n11432 DVSS.n11431 2.2505
R34168 DVSS.n11434 DVSS.n11433 2.2505
R34169 DVSS.n11204 DVSS.n11203 2.2505
R34170 DVSS.n11439 DVSS.n11438 2.2505
R34171 DVSS.n11441 DVSS.n11440 2.2505
R34172 DVSS.n11443 DVSS.n11442 2.2505
R34173 DVSS.n11201 DVSS.n11200 2.2505
R34174 DVSS.n13336 DVSS.n13335 2.2505
R34175 DVSS.n13321 DVSS.n13320 2.2505
R34176 DVSS.n13319 DVSS.n11548 2.2505
R34177 DVSS.n13318 DVSS.n13317 2.2505
R34178 DVSS.n13315 DVSS.n11549 2.2505
R34179 DVSS.n13313 DVSS.n13311 2.2505
R34180 DVSS.n13310 DVSS.n11551 2.2505
R34181 DVSS.n13309 DVSS.n13308 2.2505
R34182 DVSS.n13306 DVSS.n11552 2.2505
R34183 DVSS.n13304 DVSS.n13302 2.2505
R34184 DVSS.n13301 DVSS.n11554 2.2505
R34185 DVSS.n13300 DVSS.n13299 2.2505
R34186 DVSS.n13297 DVSS.n11555 2.2505
R34187 DVSS.n13295 DVSS.n13293 2.2505
R34188 DVSS.n13292 DVSS.n11557 2.2505
R34189 DVSS.n13291 DVSS.n13290 2.2505
R34190 DVSS.n13288 DVSS.n11558 2.2505
R34191 DVSS.n13286 DVSS.n13284 2.2505
R34192 DVSS.n13283 DVSS.n11560 2.2505
R34193 DVSS.n13282 DVSS.n13281 2.2505
R34194 DVSS.n13279 DVSS.n11561 2.2505
R34195 DVSS.n13277 DVSS.n13275 2.2505
R34196 DVSS.n13274 DVSS.n11563 2.2505
R34197 DVSS.n13273 DVSS.n13272 2.2505
R34198 DVSS.n13270 DVSS.n11564 2.2505
R34199 DVSS.n13268 DVSS.n13266 2.2505
R34200 DVSS.n13265 DVSS.n11566 2.2505
R34201 DVSS.n13264 DVSS.n13263 2.2505
R34202 DVSS.n13261 DVSS.n11567 2.2505
R34203 DVSS.n13259 DVSS.n13257 2.2505
R34204 DVSS.n13256 DVSS.n11569 2.2505
R34205 DVSS.n13255 DVSS.n13254 2.2505
R34206 DVSS.n13252 DVSS.n11570 2.2505
R34207 DVSS.n13250 DVSS.n13248 2.2505
R34208 DVSS.n13247 DVSS.n11572 2.2505
R34209 DVSS.n13246 DVSS.n13245 2.2505
R34210 DVSS.n13243 DVSS.n11573 2.2505
R34211 DVSS.n13241 DVSS.n13239 2.2505
R34212 DVSS.n13238 DVSS.n11575 2.2505
R34213 DVSS.n13237 DVSS.n13236 2.2505
R34214 DVSS.n13234 DVSS.n11576 2.2505
R34215 DVSS.n13232 DVSS.n13230 2.2505
R34216 DVSS.n13229 DVSS.n11578 2.2505
R34217 DVSS.n13228 DVSS.n13227 2.2505
R34218 DVSS.n13225 DVSS.n11579 2.2505
R34219 DVSS.n13223 DVSS.n13221 2.2505
R34220 DVSS.n13220 DVSS.n11581 2.2505
R34221 DVSS.n13219 DVSS.n13218 2.2505
R34222 DVSS.n13216 DVSS.n11582 2.2505
R34223 DVSS.n13214 DVSS.n13212 2.2505
R34224 DVSS.n13211 DVSS.n11584 2.2505
R34225 DVSS.n13210 DVSS.n13209 2.2505
R34226 DVSS.n13207 DVSS.n11585 2.2505
R34227 DVSS.n13205 DVSS.n13203 2.2505
R34228 DVSS.n13202 DVSS.n11587 2.2505
R34229 DVSS.n13201 DVSS.n13200 2.2505
R34230 DVSS.n13198 DVSS.n11588 2.2505
R34231 DVSS.n13196 DVSS.n13194 2.2505
R34232 DVSS.n13193 DVSS.n11590 2.2505
R34233 DVSS.n13192 DVSS.n13191 2.2505
R34234 DVSS.n13189 DVSS.n11591 2.2505
R34235 DVSS.n13187 DVSS.n13185 2.2505
R34236 DVSS.n13184 DVSS.n11593 2.2505
R34237 DVSS.n13183 DVSS.n13182 2.2505
R34238 DVSS.n13180 DVSS.n11594 2.2505
R34239 DVSS.n13178 DVSS.n13176 2.2505
R34240 DVSS.n13175 DVSS.n11596 2.2505
R34241 DVSS.n13174 DVSS.n13173 2.2505
R34242 DVSS.n13171 DVSS.n11597 2.2505
R34243 DVSS.n13169 DVSS.n13167 2.2505
R34244 DVSS.n13166 DVSS.n11599 2.2505
R34245 DVSS.n13165 DVSS.n13164 2.2505
R34246 DVSS.n13162 DVSS.n11600 2.2505
R34247 DVSS.n13160 DVSS.n13158 2.2505
R34248 DVSS.n13157 DVSS.n11602 2.2505
R34249 DVSS.n13156 DVSS.n13155 2.2505
R34250 DVSS.n13153 DVSS.n11603 2.2505
R34251 DVSS.n13151 DVSS.n13149 2.2505
R34252 DVSS.n13148 DVSS.n11605 2.2505
R34253 DVSS.n13147 DVSS.n13146 2.2505
R34254 DVSS.n13144 DVSS.n11606 2.2505
R34255 DVSS.n13142 DVSS.n13140 2.2505
R34256 DVSS.n13139 DVSS.n11608 2.2505
R34257 DVSS.n13138 DVSS.n13137 2.2505
R34258 DVSS.n13136 DVSS.n11503 2.2505
R34259 DVSS.n13324 DVSS.n11503 2.2505
R34260 DVSS.n13137 DVSS.n11501 2.2505
R34261 DVSS.n11608 DVSS.n11607 2.2505
R34262 DVSS.n13142 DVSS.n13141 2.2505
R34263 DVSS.n13144 DVSS.n13143 2.2505
R34264 DVSS.n13146 DVSS.n13145 2.2505
R34265 DVSS.n11605 DVSS.n11604 2.2505
R34266 DVSS.n13151 DVSS.n13150 2.2505
R34267 DVSS.n13153 DVSS.n13152 2.2505
R34268 DVSS.n13155 DVSS.n13154 2.2505
R34269 DVSS.n11602 DVSS.n11601 2.2505
R34270 DVSS.n13160 DVSS.n13159 2.2505
R34271 DVSS.n13162 DVSS.n13161 2.2505
R34272 DVSS.n13164 DVSS.n13163 2.2505
R34273 DVSS.n11599 DVSS.n11598 2.2505
R34274 DVSS.n13169 DVSS.n13168 2.2505
R34275 DVSS.n13171 DVSS.n13170 2.2505
R34276 DVSS.n13173 DVSS.n13172 2.2505
R34277 DVSS.n11596 DVSS.n11595 2.2505
R34278 DVSS.n13178 DVSS.n13177 2.2505
R34279 DVSS.n13180 DVSS.n13179 2.2505
R34280 DVSS.n13182 DVSS.n13181 2.2505
R34281 DVSS.n11593 DVSS.n11592 2.2505
R34282 DVSS.n13187 DVSS.n13186 2.2505
R34283 DVSS.n13189 DVSS.n13188 2.2505
R34284 DVSS.n13191 DVSS.n13190 2.2505
R34285 DVSS.n11590 DVSS.n11589 2.2505
R34286 DVSS.n13196 DVSS.n13195 2.2505
R34287 DVSS.n13198 DVSS.n13197 2.2505
R34288 DVSS.n13200 DVSS.n13199 2.2505
R34289 DVSS.n11587 DVSS.n11586 2.2505
R34290 DVSS.n13205 DVSS.n13204 2.2505
R34291 DVSS.n13207 DVSS.n13206 2.2505
R34292 DVSS.n13209 DVSS.n13208 2.2505
R34293 DVSS.n11584 DVSS.n11583 2.2505
R34294 DVSS.n13214 DVSS.n13213 2.2505
R34295 DVSS.n13216 DVSS.n13215 2.2505
R34296 DVSS.n13218 DVSS.n13217 2.2505
R34297 DVSS.n11581 DVSS.n11580 2.2505
R34298 DVSS.n13223 DVSS.n13222 2.2505
R34299 DVSS.n13225 DVSS.n13224 2.2505
R34300 DVSS.n13227 DVSS.n13226 2.2505
R34301 DVSS.n11578 DVSS.n11577 2.2505
R34302 DVSS.n13232 DVSS.n13231 2.2505
R34303 DVSS.n13234 DVSS.n13233 2.2505
R34304 DVSS.n13236 DVSS.n13235 2.2505
R34305 DVSS.n11575 DVSS.n11574 2.2505
R34306 DVSS.n13241 DVSS.n13240 2.2505
R34307 DVSS.n13243 DVSS.n13242 2.2505
R34308 DVSS.n13245 DVSS.n13244 2.2505
R34309 DVSS.n11572 DVSS.n11571 2.2505
R34310 DVSS.n13250 DVSS.n13249 2.2505
R34311 DVSS.n13252 DVSS.n13251 2.2505
R34312 DVSS.n13254 DVSS.n13253 2.2505
R34313 DVSS.n11569 DVSS.n11568 2.2505
R34314 DVSS.n13259 DVSS.n13258 2.2505
R34315 DVSS.n13261 DVSS.n13260 2.2505
R34316 DVSS.n13263 DVSS.n13262 2.2505
R34317 DVSS.n11566 DVSS.n11565 2.2505
R34318 DVSS.n13268 DVSS.n13267 2.2505
R34319 DVSS.n13270 DVSS.n13269 2.2505
R34320 DVSS.n13272 DVSS.n13271 2.2505
R34321 DVSS.n11563 DVSS.n11562 2.2505
R34322 DVSS.n13277 DVSS.n13276 2.2505
R34323 DVSS.n13279 DVSS.n13278 2.2505
R34324 DVSS.n13281 DVSS.n13280 2.2505
R34325 DVSS.n11560 DVSS.n11559 2.2505
R34326 DVSS.n13286 DVSS.n13285 2.2505
R34327 DVSS.n13288 DVSS.n13287 2.2505
R34328 DVSS.n13290 DVSS.n13289 2.2505
R34329 DVSS.n11557 DVSS.n11556 2.2505
R34330 DVSS.n13295 DVSS.n13294 2.2505
R34331 DVSS.n13297 DVSS.n13296 2.2505
R34332 DVSS.n13299 DVSS.n13298 2.2505
R34333 DVSS.n11554 DVSS.n11553 2.2505
R34334 DVSS.n13304 DVSS.n13303 2.2505
R34335 DVSS.n13306 DVSS.n13305 2.2505
R34336 DVSS.n13308 DVSS.n13307 2.2505
R34337 DVSS.n11551 DVSS.n11550 2.2505
R34338 DVSS.n13313 DVSS.n13312 2.2505
R34339 DVSS.n13315 DVSS.n13314 2.2505
R34340 DVSS.n13317 DVSS.n13316 2.2505
R34341 DVSS.n11548 DVSS.n11547 2.2505
R34342 DVSS.n13322 DVSS.n13321 2.2505
R34343 DVSS.n7027 DVSS.n7026 2.2505
R34344 DVSS.n6695 DVSS.n6694 2.2505
R34345 DVSS.n7020 DVSS.n7019 2.2505
R34346 DVSS.n7018 DVSS.n6697 2.2505
R34347 DVSS.n7017 DVSS.n7016 2.2505
R34348 DVSS.n6699 DVSS.n6698 2.2505
R34349 DVSS.n7008 DVSS.n7007 2.2505
R34350 DVSS.n7006 DVSS.n6701 2.2505
R34351 DVSS.n7005 DVSS.n7004 2.2505
R34352 DVSS.n6703 DVSS.n6702 2.2505
R34353 DVSS.n6996 DVSS.n6995 2.2505
R34354 DVSS.n6994 DVSS.n6705 2.2505
R34355 DVSS.n6993 DVSS.n6992 2.2505
R34356 DVSS.n6707 DVSS.n6706 2.2505
R34357 DVSS.n6984 DVSS.n6983 2.2505
R34358 DVSS.n6982 DVSS.n6709 2.2505
R34359 DVSS.n6981 DVSS.n6980 2.2505
R34360 DVSS.n6711 DVSS.n6710 2.2505
R34361 DVSS.n6972 DVSS.n6971 2.2505
R34362 DVSS.n6970 DVSS.n6713 2.2505
R34363 DVSS.n6969 DVSS.n6968 2.2505
R34364 DVSS.n6715 DVSS.n6714 2.2505
R34365 DVSS.n6960 DVSS.n6959 2.2505
R34366 DVSS.n6958 DVSS.n6717 2.2505
R34367 DVSS.n6957 DVSS.n6956 2.2505
R34368 DVSS.n6719 DVSS.n6718 2.2505
R34369 DVSS.n6948 DVSS.n6947 2.2505
R34370 DVSS.n6946 DVSS.n6721 2.2505
R34371 DVSS.n6945 DVSS.n6944 2.2505
R34372 DVSS.n6723 DVSS.n6722 2.2505
R34373 DVSS.n6936 DVSS.n6935 2.2505
R34374 DVSS.n6934 DVSS.n6725 2.2505
R34375 DVSS.n6933 DVSS.n6932 2.2505
R34376 DVSS.n6727 DVSS.n6726 2.2505
R34377 DVSS.n6924 DVSS.n6923 2.2505
R34378 DVSS.n6922 DVSS.n6729 2.2505
R34379 DVSS.n6921 DVSS.n6920 2.2505
R34380 DVSS.n6731 DVSS.n6730 2.2505
R34381 DVSS.n6912 DVSS.n6911 2.2505
R34382 DVSS.n6910 DVSS.n6733 2.2505
R34383 DVSS.n6909 DVSS.n6908 2.2505
R34384 DVSS.n6735 DVSS.n6734 2.2505
R34385 DVSS.n6900 DVSS.n6899 2.2505
R34386 DVSS.n6898 DVSS.n6737 2.2505
R34387 DVSS.n6897 DVSS.n6896 2.2505
R34388 DVSS.n6739 DVSS.n6738 2.2505
R34389 DVSS.n6888 DVSS.n6887 2.2505
R34390 DVSS.n6886 DVSS.n6741 2.2505
R34391 DVSS.n6885 DVSS.n6884 2.2505
R34392 DVSS.n6743 DVSS.n6742 2.2505
R34393 DVSS.n6876 DVSS.n6875 2.2505
R34394 DVSS.n6874 DVSS.n6745 2.2505
R34395 DVSS.n6873 DVSS.n6872 2.2505
R34396 DVSS.n6747 DVSS.n6746 2.2505
R34397 DVSS.n6864 DVSS.n6863 2.2505
R34398 DVSS.n6862 DVSS.n6749 2.2505
R34399 DVSS.n6861 DVSS.n6860 2.2505
R34400 DVSS.n6751 DVSS.n6750 2.2505
R34401 DVSS.n6852 DVSS.n6851 2.2505
R34402 DVSS.n6850 DVSS.n6753 2.2505
R34403 DVSS.n6849 DVSS.n6848 2.2505
R34404 DVSS.n6755 DVSS.n6754 2.2505
R34405 DVSS.n6840 DVSS.n6839 2.2505
R34406 DVSS.n6838 DVSS.n6757 2.2505
R34407 DVSS.n6837 DVSS.n6836 2.2505
R34408 DVSS.n6759 DVSS.n6758 2.2505
R34409 DVSS.n6828 DVSS.n6827 2.2505
R34410 DVSS.n6826 DVSS.n6761 2.2505
R34411 DVSS.n6825 DVSS.n6824 2.2505
R34412 DVSS.n6763 DVSS.n6762 2.2505
R34413 DVSS.n6816 DVSS.n6815 2.2505
R34414 DVSS.n6814 DVSS.n6765 2.2505
R34415 DVSS.n6813 DVSS.n6812 2.2505
R34416 DVSS.n6767 DVSS.n6766 2.2505
R34417 DVSS.n6804 DVSS.n6803 2.2505
R34418 DVSS.n6802 DVSS.n6769 2.2505
R34419 DVSS.n6801 DVSS.n6800 2.2505
R34420 DVSS.n6771 DVSS.n6770 2.2505
R34421 DVSS.n6792 DVSS.n6791 2.2505
R34422 DVSS.n6790 DVSS.n6773 2.2505
R34423 DVSS.n6789 DVSS.n6788 2.2505
R34424 DVSS.n6775 DVSS.n6774 2.2505
R34425 DVSS.n6780 DVSS.n6779 2.2505
R34426 DVSS.n6778 DVSS.n5872 2.2505
R34427 DVSS.n6778 DVSS.n6777 2.2505
R34428 DVSS.n6781 DVSS.n6780 2.2505
R34429 DVSS.n6783 DVSS.n6775 2.2505
R34430 DVSS.n6788 DVSS.n6787 2.2505
R34431 DVSS.n6785 DVSS.n6773 2.2505
R34432 DVSS.n6793 DVSS.n6792 2.2505
R34433 DVSS.n6795 DVSS.n6771 2.2505
R34434 DVSS.n6800 DVSS.n6799 2.2505
R34435 DVSS.n6797 DVSS.n6769 2.2505
R34436 DVSS.n6805 DVSS.n6804 2.2505
R34437 DVSS.n6807 DVSS.n6767 2.2505
R34438 DVSS.n6812 DVSS.n6811 2.2505
R34439 DVSS.n6809 DVSS.n6765 2.2505
R34440 DVSS.n6817 DVSS.n6816 2.2505
R34441 DVSS.n6819 DVSS.n6763 2.2505
R34442 DVSS.n6824 DVSS.n6823 2.2505
R34443 DVSS.n6821 DVSS.n6761 2.2505
R34444 DVSS.n6829 DVSS.n6828 2.2505
R34445 DVSS.n6831 DVSS.n6759 2.2505
R34446 DVSS.n6836 DVSS.n6835 2.2505
R34447 DVSS.n6833 DVSS.n6757 2.2505
R34448 DVSS.n6841 DVSS.n6840 2.2505
R34449 DVSS.n6843 DVSS.n6755 2.2505
R34450 DVSS.n6848 DVSS.n6847 2.2505
R34451 DVSS.n6845 DVSS.n6753 2.2505
R34452 DVSS.n6853 DVSS.n6852 2.2505
R34453 DVSS.n6855 DVSS.n6751 2.2505
R34454 DVSS.n6860 DVSS.n6859 2.2505
R34455 DVSS.n6857 DVSS.n6749 2.2505
R34456 DVSS.n6865 DVSS.n6864 2.2505
R34457 DVSS.n6867 DVSS.n6747 2.2505
R34458 DVSS.n6872 DVSS.n6871 2.2505
R34459 DVSS.n6869 DVSS.n6745 2.2505
R34460 DVSS.n6877 DVSS.n6876 2.2505
R34461 DVSS.n6879 DVSS.n6743 2.2505
R34462 DVSS.n6884 DVSS.n6883 2.2505
R34463 DVSS.n6881 DVSS.n6741 2.2505
R34464 DVSS.n6889 DVSS.n6888 2.2505
R34465 DVSS.n6891 DVSS.n6739 2.2505
R34466 DVSS.n6896 DVSS.n6895 2.2505
R34467 DVSS.n6893 DVSS.n6737 2.2505
R34468 DVSS.n6901 DVSS.n6900 2.2505
R34469 DVSS.n6903 DVSS.n6735 2.2505
R34470 DVSS.n6908 DVSS.n6907 2.2505
R34471 DVSS.n6905 DVSS.n6733 2.2505
R34472 DVSS.n6913 DVSS.n6912 2.2505
R34473 DVSS.n6915 DVSS.n6731 2.2505
R34474 DVSS.n6920 DVSS.n6919 2.2505
R34475 DVSS.n6917 DVSS.n6729 2.2505
R34476 DVSS.n6925 DVSS.n6924 2.2505
R34477 DVSS.n6927 DVSS.n6727 2.2505
R34478 DVSS.n6932 DVSS.n6931 2.2505
R34479 DVSS.n6929 DVSS.n6725 2.2505
R34480 DVSS.n6937 DVSS.n6936 2.2505
R34481 DVSS.n6939 DVSS.n6723 2.2505
R34482 DVSS.n6944 DVSS.n6943 2.2505
R34483 DVSS.n6941 DVSS.n6721 2.2505
R34484 DVSS.n6949 DVSS.n6948 2.2505
R34485 DVSS.n6951 DVSS.n6719 2.2505
R34486 DVSS.n6956 DVSS.n6955 2.2505
R34487 DVSS.n6953 DVSS.n6717 2.2505
R34488 DVSS.n6961 DVSS.n6960 2.2505
R34489 DVSS.n6963 DVSS.n6715 2.2505
R34490 DVSS.n6968 DVSS.n6967 2.2505
R34491 DVSS.n6965 DVSS.n6713 2.2505
R34492 DVSS.n6973 DVSS.n6972 2.2505
R34493 DVSS.n6975 DVSS.n6711 2.2505
R34494 DVSS.n6980 DVSS.n6979 2.2505
R34495 DVSS.n6977 DVSS.n6709 2.2505
R34496 DVSS.n6985 DVSS.n6984 2.2505
R34497 DVSS.n6987 DVSS.n6707 2.2505
R34498 DVSS.n6992 DVSS.n6991 2.2505
R34499 DVSS.n6989 DVSS.n6705 2.2505
R34500 DVSS.n6997 DVSS.n6996 2.2505
R34501 DVSS.n6999 DVSS.n6703 2.2505
R34502 DVSS.n7004 DVSS.n7003 2.2505
R34503 DVSS.n7001 DVSS.n6701 2.2505
R34504 DVSS.n7009 DVSS.n7008 2.2505
R34505 DVSS.n7011 DVSS.n6699 2.2505
R34506 DVSS.n7016 DVSS.n7015 2.2505
R34507 DVSS.n7013 DVSS.n6697 2.2505
R34508 DVSS.n7021 DVSS.n7020 2.2505
R34509 DVSS.n7023 DVSS.n6695 2.2505
R34510 DVSS.n7026 DVSS.n7025 2.2505
R34511 DVSS.n6672 DVSS.n6671 2.2505
R34512 DVSS.n6239 DVSS.n6232 2.2505
R34513 DVSS.n6679 DVSS.n6678 2.2505
R34514 DVSS.n6690 DVSS.n6689 2.2505
R34515 DVSS.n5890 DVSS.n5881 2.2505
R34516 DVSS.n7033 DVSS.n7032 2.2505
R34517 DVSS.n5867 DVSS.n5866 2.2505
R34518 DVSS.n7046 DVSS.n7045 2.2505
R34519 DVSS.n7049 DVSS.n5531 2.2505
R34520 DVSS.n5574 DVSS.n5524 2.2505
R34521 DVSS.n7070 DVSS.n7069 2.2505
R34522 DVSS.n7078 DVSS.n7077 2.2505
R34523 DVSS.n5176 DVSS.n5175 2.2505
R34524 DVSS.n7089 DVSS.n7088 2.2505
R34525 DVSS.n7092 DVSS.n4840 2.2505
R34526 DVSS.n7104 DVSS.n4831 2.2505
R34527 DVSS.n7453 DVSS.n7452 2.2505
R34528 DVSS.n7460 DVSS.n7459 2.2505
R34529 DVSS.n7796 DVSS.n4817 2.2505
R34530 DVSS.n7808 DVSS.n7807 2.2505
R34531 DVSS.n7815 DVSS.n7814 2.2505
R34532 DVSS.n7817 DVSS.n4466 2.2505
R34533 DVSS.n7828 DVSS.n7827 2.2505
R34534 DVSS.n4470 DVSS.n4460 2.2505
R34535 DVSS.n7835 DVSS.n4371 2.2505
R34536 DVSS.n7839 DVSS.n7836 2.2505
R34537 DVSS.n8101 DVSS.n4361 2.2505
R34538 DVSS.n8104 DVSS.n8103 2.2505
R34539 DVSS.n8111 DVSS.n8110 2.2505
R34540 DVSS.n4014 DVSS.n3856 2.2505
R34541 DVSS.n8322 DVSS.n8321 2.2505
R34542 DVSS.n3904 DVSS.n3847 2.2505
R34543 DVSS.n8331 DVSS.n8330 2.2505
R34544 DVSS.n3849 DVSS.n3848 2.2505
R34545 DVSS.n8591 DVSS.n8590 2.2505
R34546 DVSS.n3754 DVSS.n3415 2.2505
R34547 DVSS.n3750 DVSS.n3457 2.2505
R34548 DVSS.n3406 DVSS.n3405 2.2505
R34549 DVSS.n8617 DVSS.n8616 2.2505
R34550 DVSS.n8624 DVSS.n8623 2.2505
R34551 DVSS.n8634 DVSS.n3058 2.2505
R34552 DVSS.n8971 DVSS.n8970 2.2505
R34553 DVSS.n8978 DVSS.n8977 2.2505
R34554 DVSS.n3045 DVSS.n2888 2.2505
R34555 DVSS.n9189 DVSS.n9188 2.2505
R34556 DVSS.n2936 DVSS.n2879 2.2505
R34557 DVSS.n9198 DVSS.n9197 2.2505
R34558 DVSS.n2881 DVSS.n2880 2.2505
R34559 DVSS.n9458 DVSS.n9457 2.2505
R34560 DVSS.n2782 DVSS.n2739 2.2505
R34561 DVSS.n9465 DVSS.n9464 2.2505
R34562 DVSS.n9772 DVSS.n9771 2.2505
R34563 DVSS.n2730 DVSS.n2721 2.2505
R34564 DVSS.n10115 DVSS.n10114 2.2505
R34565 DVSS.n2706 DVSS.n2705 2.2505
R34566 DVSS.n10128 DVSS.n10127 2.2505
R34567 DVSS.n10131 DVSS.n2370 2.2505
R34568 DVSS.n10142 DVSS.n2363 2.2505
R34569 DVSS.n10153 DVSS.n10152 2.2505
R34570 DVSS.n10156 DVSS.n2027 2.2505
R34571 DVSS.n2019 DVSS.n2018 2.2505
R34572 DVSS.n10462 DVSS.n10461 2.2505
R34573 DVSS.n10465 DVSS.n1967 2.2505
R34574 DVSS.n10477 DVSS.n1626 2.2505
R34575 DVSS.n10488 DVSS.n10487 2.2505
R34576 DVSS.n10495 DVSS.n10494 2.2505
R34577 DVSS.n10497 DVSS.n1521 2.2505
R34578 DVSS.n10756 DVSS.n10755 2.2505
R34579 DVSS.n1513 DVSS.n1511 2.2505
R34580 DVSS.n13358 DVSS.n13357 2.2505
R34581 DVSS.n13351 DVSS.n13350 2.2505
R34582 DVSS.n11109 DVSS.n10764 2.2505
R34583 DVSS.n11447 DVSS.n11111 2.2505
R34584 DVSS.n11450 DVSS.n11156 2.2505
R34585 DVSS.n11457 DVSS.n11455 2.2505
R34586 DVSS.n13328 DVSS.n13327 2.2505
R34587 DVSS.n11642 DVSS.n11504 2.2505
R34588 DVSS.n11644 DVSS.n11643 2.2505
R34589 DVSS.n11983 DVSS.n11982 2.2505
R34590 DVSS.n11632 DVSS.n11630 2.2505
R34591 DVSS.n13120 DVSS.n13119 2.2505
R34592 DVSS.n12337 DVSS.n11633 2.2505
R34593 DVSS.n13112 DVSS.n13111 2.2505
R34594 DVSS.n11995 DVSS.n11993 2.2505
R34595 DVSS.n12762 DVSS.n12761 2.2505
R34596 DVSS.n5985 DVSS.n5984 2.2505
R34597 DVSS.n5986 DVSS.n5982 2.2505
R34598 DVSS.n5991 DVSS.n5987 2.2505
R34599 DVSS.n5992 DVSS.n5981 2.2505
R34600 DVSS.n5997 DVSS.n5996 2.2505
R34601 DVSS.n5998 DVSS.n5980 2.2505
R34602 DVSS.n6003 DVSS.n5999 2.2505
R34603 DVSS.n6004 DVSS.n5979 2.2505
R34604 DVSS.n6009 DVSS.n6008 2.2505
R34605 DVSS.n6010 DVSS.n5978 2.2505
R34606 DVSS.n6015 DVSS.n6011 2.2505
R34607 DVSS.n6016 DVSS.n5977 2.2505
R34608 DVSS.n6021 DVSS.n6020 2.2505
R34609 DVSS.n6022 DVSS.n5976 2.2505
R34610 DVSS.n6027 DVSS.n6023 2.2505
R34611 DVSS.n6028 DVSS.n5975 2.2505
R34612 DVSS.n6033 DVSS.n6032 2.2505
R34613 DVSS.n6034 DVSS.n5974 2.2505
R34614 DVSS.n6039 DVSS.n6035 2.2505
R34615 DVSS.n6040 DVSS.n5973 2.2505
R34616 DVSS.n6045 DVSS.n6044 2.2505
R34617 DVSS.n6046 DVSS.n5972 2.2505
R34618 DVSS.n6051 DVSS.n6047 2.2505
R34619 DVSS.n6052 DVSS.n5971 2.2505
R34620 DVSS.n6057 DVSS.n6056 2.2505
R34621 DVSS.n6058 DVSS.n5970 2.2505
R34622 DVSS.n6063 DVSS.n6059 2.2505
R34623 DVSS.n6064 DVSS.n5969 2.2505
R34624 DVSS.n6069 DVSS.n6068 2.2505
R34625 DVSS.n6070 DVSS.n5968 2.2505
R34626 DVSS.n6075 DVSS.n6071 2.2505
R34627 DVSS.n6076 DVSS.n5967 2.2505
R34628 DVSS.n6081 DVSS.n6080 2.2505
R34629 DVSS.n6082 DVSS.n5966 2.2505
R34630 DVSS.n6087 DVSS.n6083 2.2505
R34631 DVSS.n6088 DVSS.n5965 2.2505
R34632 DVSS.n6093 DVSS.n6092 2.2505
R34633 DVSS.n6094 DVSS.n5964 2.2505
R34634 DVSS.n6099 DVSS.n6095 2.2505
R34635 DVSS.n6100 DVSS.n5963 2.2505
R34636 DVSS.n6105 DVSS.n6104 2.2505
R34637 DVSS.n6106 DVSS.n5962 2.2505
R34638 DVSS.n6111 DVSS.n6107 2.2505
R34639 DVSS.n6112 DVSS.n5961 2.2505
R34640 DVSS.n6117 DVSS.n6116 2.2505
R34641 DVSS.n6118 DVSS.n5960 2.2505
R34642 DVSS.n6123 DVSS.n6119 2.2505
R34643 DVSS.n6124 DVSS.n5959 2.2505
R34644 DVSS.n6129 DVSS.n6128 2.2505
R34645 DVSS.n6130 DVSS.n5958 2.2505
R34646 DVSS.n6135 DVSS.n6131 2.2505
R34647 DVSS.n6136 DVSS.n5957 2.2505
R34648 DVSS.n6141 DVSS.n6140 2.2505
R34649 DVSS.n6142 DVSS.n5956 2.2505
R34650 DVSS.n6147 DVSS.n6143 2.2505
R34651 DVSS.n6148 DVSS.n5955 2.2505
R34652 DVSS.n6153 DVSS.n6152 2.2505
R34653 DVSS.n6154 DVSS.n5954 2.2505
R34654 DVSS.n6159 DVSS.n6155 2.2505
R34655 DVSS.n6160 DVSS.n5953 2.2505
R34656 DVSS.n6165 DVSS.n6164 2.2505
R34657 DVSS.n6166 DVSS.n5952 2.2505
R34658 DVSS.n6171 DVSS.n6167 2.2505
R34659 DVSS.n6172 DVSS.n5951 2.2505
R34660 DVSS.n6177 DVSS.n6176 2.2505
R34661 DVSS.n6178 DVSS.n5950 2.2505
R34662 DVSS.n6183 DVSS.n6179 2.2505
R34663 DVSS.n6184 DVSS.n5949 2.2505
R34664 DVSS.n6189 DVSS.n6188 2.2505
R34665 DVSS.n6190 DVSS.n5948 2.2505
R34666 DVSS.n6195 DVSS.n6191 2.2505
R34667 DVSS.n6196 DVSS.n5947 2.2505
R34668 DVSS.n6201 DVSS.n6200 2.2505
R34669 DVSS.n6202 DVSS.n5946 2.2505
R34670 DVSS.n6207 DVSS.n6203 2.2505
R34671 DVSS.n6208 DVSS.n5945 2.2505
R34672 DVSS.n6213 DVSS.n6212 2.2505
R34673 DVSS.n6214 DVSS.n5944 2.2505
R34674 DVSS.n6219 DVSS.n6215 2.2505
R34675 DVSS.n6220 DVSS.n5943 2.2505
R34676 DVSS.n6225 DVSS.n6224 2.2505
R34677 DVSS.n6226 DVSS.n5942 2.2505
R34678 DVSS.n6228 DVSS.n6227 2.2505
R34679 DVSS.n5940 DVSS.n5893 2.2505
R34680 DVSS.n5940 DVSS.n5938 2.2505
R34681 DVSS.n6229 DVSS.n6228 2.2505
R34682 DVSS.n5942 DVSS.n5941 2.2505
R34683 DVSS.n6224 DVSS.n6223 2.2505
R34684 DVSS.n6221 DVSS.n6220 2.2505
R34685 DVSS.n6219 DVSS.n6218 2.2505
R34686 DVSS.n6216 DVSS.n5944 2.2505
R34687 DVSS.n6212 DVSS.n6211 2.2505
R34688 DVSS.n6209 DVSS.n6208 2.2505
R34689 DVSS.n6207 DVSS.n6206 2.2505
R34690 DVSS.n6204 DVSS.n5946 2.2505
R34691 DVSS.n6200 DVSS.n6199 2.2505
R34692 DVSS.n6197 DVSS.n6196 2.2505
R34693 DVSS.n6195 DVSS.n6194 2.2505
R34694 DVSS.n6192 DVSS.n5948 2.2505
R34695 DVSS.n6188 DVSS.n6187 2.2505
R34696 DVSS.n6185 DVSS.n6184 2.2505
R34697 DVSS.n6183 DVSS.n6182 2.2505
R34698 DVSS.n6180 DVSS.n5950 2.2505
R34699 DVSS.n6176 DVSS.n6175 2.2505
R34700 DVSS.n6173 DVSS.n6172 2.2505
R34701 DVSS.n6171 DVSS.n6170 2.2505
R34702 DVSS.n6168 DVSS.n5952 2.2505
R34703 DVSS.n6164 DVSS.n6163 2.2505
R34704 DVSS.n6161 DVSS.n6160 2.2505
R34705 DVSS.n6159 DVSS.n6158 2.2505
R34706 DVSS.n6156 DVSS.n5954 2.2505
R34707 DVSS.n6152 DVSS.n6151 2.2505
R34708 DVSS.n6149 DVSS.n6148 2.2505
R34709 DVSS.n6147 DVSS.n6146 2.2505
R34710 DVSS.n6144 DVSS.n5956 2.2505
R34711 DVSS.n6140 DVSS.n6139 2.2505
R34712 DVSS.n6137 DVSS.n6136 2.2505
R34713 DVSS.n6135 DVSS.n6134 2.2505
R34714 DVSS.n6132 DVSS.n5958 2.2505
R34715 DVSS.n6128 DVSS.n6127 2.2505
R34716 DVSS.n6125 DVSS.n6124 2.2505
R34717 DVSS.n6123 DVSS.n6122 2.2505
R34718 DVSS.n6120 DVSS.n5960 2.2505
R34719 DVSS.n6116 DVSS.n6115 2.2505
R34720 DVSS.n6113 DVSS.n6112 2.2505
R34721 DVSS.n6111 DVSS.n6110 2.2505
R34722 DVSS.n6108 DVSS.n5962 2.2505
R34723 DVSS.n6104 DVSS.n6103 2.2505
R34724 DVSS.n6101 DVSS.n6100 2.2505
R34725 DVSS.n6099 DVSS.n6098 2.2505
R34726 DVSS.n6096 DVSS.n5964 2.2505
R34727 DVSS.n6092 DVSS.n6091 2.2505
R34728 DVSS.n6089 DVSS.n6088 2.2505
R34729 DVSS.n6087 DVSS.n6086 2.2505
R34730 DVSS.n6084 DVSS.n5966 2.2505
R34731 DVSS.n6080 DVSS.n6079 2.2505
R34732 DVSS.n6077 DVSS.n6076 2.2505
R34733 DVSS.n6075 DVSS.n6074 2.2505
R34734 DVSS.n6072 DVSS.n5968 2.2505
R34735 DVSS.n6068 DVSS.n6067 2.2505
R34736 DVSS.n6065 DVSS.n6064 2.2505
R34737 DVSS.n6063 DVSS.n6062 2.2505
R34738 DVSS.n6060 DVSS.n5970 2.2505
R34739 DVSS.n6056 DVSS.n6055 2.2505
R34740 DVSS.n6053 DVSS.n6052 2.2505
R34741 DVSS.n6051 DVSS.n6050 2.2505
R34742 DVSS.n6048 DVSS.n5972 2.2505
R34743 DVSS.n6044 DVSS.n6043 2.2505
R34744 DVSS.n6041 DVSS.n6040 2.2505
R34745 DVSS.n6039 DVSS.n6038 2.2505
R34746 DVSS.n6036 DVSS.n5974 2.2505
R34747 DVSS.n6032 DVSS.n6031 2.2505
R34748 DVSS.n6029 DVSS.n6028 2.2505
R34749 DVSS.n6027 DVSS.n6026 2.2505
R34750 DVSS.n6024 DVSS.n5976 2.2505
R34751 DVSS.n6020 DVSS.n6019 2.2505
R34752 DVSS.n6017 DVSS.n6016 2.2505
R34753 DVSS.n6015 DVSS.n6014 2.2505
R34754 DVSS.n6012 DVSS.n5978 2.2505
R34755 DVSS.n6008 DVSS.n6007 2.2505
R34756 DVSS.n6005 DVSS.n6004 2.2505
R34757 DVSS.n6003 DVSS.n6002 2.2505
R34758 DVSS.n6000 DVSS.n5980 2.2505
R34759 DVSS.n5996 DVSS.n5995 2.2505
R34760 DVSS.n5993 DVSS.n5992 2.2505
R34761 DVSS.n5991 DVSS.n5990 2.2505
R34762 DVSS.n5988 DVSS.n5982 2.2505
R34763 DVSS.n5984 DVSS.n5983 2.2505
R34764 DVSS.n11978 DVSS.n11636 2.2505
R34765 DVSS.n11977 DVSS.n11975 2.2505
R34766 DVSS.n11974 DVSS.n11690 2.2505
R34767 DVSS.n11973 DVSS.n11972 2.2505
R34768 DVSS.n11968 DVSS.n11691 2.2505
R34769 DVSS.n11964 DVSS.n11963 2.2505
R34770 DVSS.n11962 DVSS.n11692 2.2505
R34771 DVSS.n11961 DVSS.n11960 2.2505
R34772 DVSS.n11956 DVSS.n11693 2.2505
R34773 DVSS.n11952 DVSS.n11951 2.2505
R34774 DVSS.n11950 DVSS.n11694 2.2505
R34775 DVSS.n11949 DVSS.n11948 2.2505
R34776 DVSS.n11944 DVSS.n11695 2.2505
R34777 DVSS.n11940 DVSS.n11939 2.2505
R34778 DVSS.n11938 DVSS.n11696 2.2505
R34779 DVSS.n11937 DVSS.n11936 2.2505
R34780 DVSS.n11932 DVSS.n11697 2.2505
R34781 DVSS.n11928 DVSS.n11927 2.2505
R34782 DVSS.n11926 DVSS.n11698 2.2505
R34783 DVSS.n11925 DVSS.n11924 2.2505
R34784 DVSS.n11920 DVSS.n11699 2.2505
R34785 DVSS.n11916 DVSS.n11915 2.2505
R34786 DVSS.n11914 DVSS.n11700 2.2505
R34787 DVSS.n11913 DVSS.n11912 2.2505
R34788 DVSS.n11908 DVSS.n11701 2.2505
R34789 DVSS.n11904 DVSS.n11903 2.2505
R34790 DVSS.n11902 DVSS.n11702 2.2505
R34791 DVSS.n11901 DVSS.n11900 2.2505
R34792 DVSS.n11896 DVSS.n11703 2.2505
R34793 DVSS.n11892 DVSS.n11891 2.2505
R34794 DVSS.n11890 DVSS.n11704 2.2505
R34795 DVSS.n11889 DVSS.n11888 2.2505
R34796 DVSS.n11884 DVSS.n11705 2.2505
R34797 DVSS.n11880 DVSS.n11879 2.2505
R34798 DVSS.n11878 DVSS.n11706 2.2505
R34799 DVSS.n11877 DVSS.n11876 2.2505
R34800 DVSS.n11872 DVSS.n11707 2.2505
R34801 DVSS.n11868 DVSS.n11867 2.2505
R34802 DVSS.n11866 DVSS.n11708 2.2505
R34803 DVSS.n11865 DVSS.n11864 2.2505
R34804 DVSS.n11860 DVSS.n11709 2.2505
R34805 DVSS.n11856 DVSS.n11855 2.2505
R34806 DVSS.n11854 DVSS.n11710 2.2505
R34807 DVSS.n11853 DVSS.n11852 2.2505
R34808 DVSS.n11848 DVSS.n11711 2.2505
R34809 DVSS.n11844 DVSS.n11843 2.2505
R34810 DVSS.n11842 DVSS.n11712 2.2505
R34811 DVSS.n11841 DVSS.n11840 2.2505
R34812 DVSS.n11836 DVSS.n11713 2.2505
R34813 DVSS.n11832 DVSS.n11831 2.2505
R34814 DVSS.n11830 DVSS.n11714 2.2505
R34815 DVSS.n11829 DVSS.n11828 2.2505
R34816 DVSS.n11824 DVSS.n11715 2.2505
R34817 DVSS.n11820 DVSS.n11819 2.2505
R34818 DVSS.n11818 DVSS.n11716 2.2505
R34819 DVSS.n11817 DVSS.n11816 2.2505
R34820 DVSS.n11812 DVSS.n11717 2.2505
R34821 DVSS.n11808 DVSS.n11807 2.2505
R34822 DVSS.n11806 DVSS.n11718 2.2505
R34823 DVSS.n11805 DVSS.n11804 2.2505
R34824 DVSS.n11800 DVSS.n11719 2.2505
R34825 DVSS.n11796 DVSS.n11795 2.2505
R34826 DVSS.n11794 DVSS.n11720 2.2505
R34827 DVSS.n11793 DVSS.n11792 2.2505
R34828 DVSS.n11788 DVSS.n11721 2.2505
R34829 DVSS.n11784 DVSS.n11783 2.2505
R34830 DVSS.n11782 DVSS.n11722 2.2505
R34831 DVSS.n11781 DVSS.n11780 2.2505
R34832 DVSS.n11776 DVSS.n11723 2.2505
R34833 DVSS.n11772 DVSS.n11771 2.2505
R34834 DVSS.n11770 DVSS.n11724 2.2505
R34835 DVSS.n11769 DVSS.n11768 2.2505
R34836 DVSS.n11764 DVSS.n11725 2.2505
R34837 DVSS.n11760 DVSS.n11759 2.2505
R34838 DVSS.n11758 DVSS.n11726 2.2505
R34839 DVSS.n11757 DVSS.n11756 2.2505
R34840 DVSS.n11752 DVSS.n11727 2.2505
R34841 DVSS.n11748 DVSS.n11747 2.2505
R34842 DVSS.n11746 DVSS.n11728 2.2505
R34843 DVSS.n11745 DVSS.n11744 2.2505
R34844 DVSS.n11740 DVSS.n11729 2.2505
R34845 DVSS.n11736 DVSS.n11735 2.2505
R34846 DVSS.n11734 DVSS.n11733 2.2505
R34847 DVSS.n11730 DVSS.n11624 2.2505
R34848 DVSS.n11730 DVSS.n11688 2.2505
R34849 DVSS.n11733 DVSS.n11732 2.2505
R34850 DVSS.n11737 DVSS.n11736 2.2505
R34851 DVSS.n11740 DVSS.n11739 2.2505
R34852 DVSS.n11744 DVSS.n11743 2.2505
R34853 DVSS.n11741 DVSS.n11728 2.2505
R34854 DVSS.n11749 DVSS.n11748 2.2505
R34855 DVSS.n11752 DVSS.n11751 2.2505
R34856 DVSS.n11756 DVSS.n11755 2.2505
R34857 DVSS.n11753 DVSS.n11726 2.2505
R34858 DVSS.n11761 DVSS.n11760 2.2505
R34859 DVSS.n11764 DVSS.n11763 2.2505
R34860 DVSS.n11768 DVSS.n11767 2.2505
R34861 DVSS.n11765 DVSS.n11724 2.2505
R34862 DVSS.n11773 DVSS.n11772 2.2505
R34863 DVSS.n11776 DVSS.n11775 2.2505
R34864 DVSS.n11780 DVSS.n11779 2.2505
R34865 DVSS.n11777 DVSS.n11722 2.2505
R34866 DVSS.n11785 DVSS.n11784 2.2505
R34867 DVSS.n11788 DVSS.n11787 2.2505
R34868 DVSS.n11792 DVSS.n11791 2.2505
R34869 DVSS.n11789 DVSS.n11720 2.2505
R34870 DVSS.n11797 DVSS.n11796 2.2505
R34871 DVSS.n11800 DVSS.n11799 2.2505
R34872 DVSS.n11804 DVSS.n11803 2.2505
R34873 DVSS.n11801 DVSS.n11718 2.2505
R34874 DVSS.n11809 DVSS.n11808 2.2505
R34875 DVSS.n11812 DVSS.n11811 2.2505
R34876 DVSS.n11816 DVSS.n11815 2.2505
R34877 DVSS.n11813 DVSS.n11716 2.2505
R34878 DVSS.n11821 DVSS.n11820 2.2505
R34879 DVSS.n11824 DVSS.n11823 2.2505
R34880 DVSS.n11828 DVSS.n11827 2.2505
R34881 DVSS.n11825 DVSS.n11714 2.2505
R34882 DVSS.n11833 DVSS.n11832 2.2505
R34883 DVSS.n11836 DVSS.n11835 2.2505
R34884 DVSS.n11840 DVSS.n11839 2.2505
R34885 DVSS.n11837 DVSS.n11712 2.2505
R34886 DVSS.n11845 DVSS.n11844 2.2505
R34887 DVSS.n11848 DVSS.n11847 2.2505
R34888 DVSS.n11852 DVSS.n11851 2.2505
R34889 DVSS.n11849 DVSS.n11710 2.2505
R34890 DVSS.n11857 DVSS.n11856 2.2505
R34891 DVSS.n11860 DVSS.n11859 2.2505
R34892 DVSS.n11864 DVSS.n11863 2.2505
R34893 DVSS.n11861 DVSS.n11708 2.2505
R34894 DVSS.n11869 DVSS.n11868 2.2505
R34895 DVSS.n11872 DVSS.n11871 2.2505
R34896 DVSS.n11876 DVSS.n11875 2.2505
R34897 DVSS.n11873 DVSS.n11706 2.2505
R34898 DVSS.n11881 DVSS.n11880 2.2505
R34899 DVSS.n11884 DVSS.n11883 2.2505
R34900 DVSS.n11888 DVSS.n11887 2.2505
R34901 DVSS.n11885 DVSS.n11704 2.2505
R34902 DVSS.n11893 DVSS.n11892 2.2505
R34903 DVSS.n11896 DVSS.n11895 2.2505
R34904 DVSS.n11900 DVSS.n11899 2.2505
R34905 DVSS.n11897 DVSS.n11702 2.2505
R34906 DVSS.n11905 DVSS.n11904 2.2505
R34907 DVSS.n11908 DVSS.n11907 2.2505
R34908 DVSS.n11912 DVSS.n11911 2.2505
R34909 DVSS.n11909 DVSS.n11700 2.2505
R34910 DVSS.n11917 DVSS.n11916 2.2505
R34911 DVSS.n11920 DVSS.n11919 2.2505
R34912 DVSS.n11924 DVSS.n11923 2.2505
R34913 DVSS.n11921 DVSS.n11698 2.2505
R34914 DVSS.n11929 DVSS.n11928 2.2505
R34915 DVSS.n11932 DVSS.n11931 2.2505
R34916 DVSS.n11936 DVSS.n11935 2.2505
R34917 DVSS.n11933 DVSS.n11696 2.2505
R34918 DVSS.n11941 DVSS.n11940 2.2505
R34919 DVSS.n11944 DVSS.n11943 2.2505
R34920 DVSS.n11948 DVSS.n11947 2.2505
R34921 DVSS.n11945 DVSS.n11694 2.2505
R34922 DVSS.n11953 DVSS.n11952 2.2505
R34923 DVSS.n11956 DVSS.n11955 2.2505
R34924 DVSS.n11960 DVSS.n11959 2.2505
R34925 DVSS.n11957 DVSS.n11692 2.2505
R34926 DVSS.n11965 DVSS.n11964 2.2505
R34927 DVSS.n11968 DVSS.n11967 2.2505
R34928 DVSS.n11972 DVSS.n11971 2.2505
R34929 DVSS.n11969 DVSS.n11690 2.2505
R34930 DVSS.n11977 DVSS.n11976 2.2505
R34931 DVSS.n11979 DVSS.n11978 2.2505
R34932 DVSS.n6673 DVSS.n6672 2.2505
R34933 DVSS.n6233 DVSS.n6232 2.2505
R34934 DVSS.n6678 DVSS.n6677 2.2505
R34935 DVSS.n6691 DVSS.n6690 2.2505
R34936 DVSS.n5883 DVSS.n5881 2.2505
R34937 DVSS.n7032 DVSS.n7031 2.2505
R34938 DVSS.n5866 DVSS.n5865 2.2505
R34939 DVSS.n7047 DVSS.n7046 2.2505
R34940 DVSS.n7050 DVSS.n7049 2.2505
R34941 DVSS.n5524 DVSS.n5523 2.2505
R34942 DVSS.n7071 DVSS.n7070 2.2505
R34943 DVSS.n7077 DVSS.n7076 2.2505
R34944 DVSS.n5175 DVSS.n5174 2.2505
R34945 DVSS.n7090 DVSS.n7089 2.2505
R34946 DVSS.n7093 DVSS.n7092 2.2505
R34947 DVSS.n4831 DVSS.n4830 2.2505
R34948 DVSS.n7454 DVSS.n7453 2.2505
R34949 DVSS.n7459 DVSS.n7458 2.2505
R34950 DVSS.n4817 DVSS.n4816 2.2505
R34951 DVSS.n7809 DVSS.n7808 2.2505
R34952 DVSS.n7814 DVSS.n7813 2.2505
R34953 DVSS.n4466 DVSS.n4464 2.2505
R34954 DVSS.n7829 DVSS.n7828 2.2505
R34955 DVSS.n4461 DVSS.n4460 2.2505
R34956 DVSS.n7835 DVSS.n7834 2.2505
R34957 DVSS.n7839 DVSS.n7838 2.2505
R34958 DVSS.n4361 DVSS.n4360 2.2505
R34959 DVSS.n8105 DVSS.n8104 2.2505
R34960 DVSS.n8110 DVSS.n8109 2.2505
R34961 DVSS.n3856 DVSS.n3854 2.2505
R34962 DVSS.n8323 DVSS.n8322 2.2505
R34963 DVSS.n3850 DVSS.n3847 2.2505
R34964 DVSS.n8330 DVSS.n8329 2.2505
R34965 DVSS.n3851 DVSS.n3849 2.2505
R34966 DVSS.n8592 DVSS.n8591 2.2505
R34967 DVSS.n3754 DVSS.n3749 2.2505
R34968 DVSS.n8597 DVSS.n3750 2.2505
R34969 DVSS.n3405 DVSS.n3404 2.2505
R34970 DVSS.n8618 DVSS.n8617 2.2505
R34971 DVSS.n8623 DVSS.n8622 2.2505
R34972 DVSS.n3058 DVSS.n3057 2.2505
R34973 DVSS.n8972 DVSS.n8971 2.2505
R34974 DVSS.n8977 DVSS.n8976 2.2505
R34975 DVSS.n2888 DVSS.n2886 2.2505
R34976 DVSS.n9190 DVSS.n9189 2.2505
R34977 DVSS.n2882 DVSS.n2879 2.2505
R34978 DVSS.n9197 DVSS.n9196 2.2505
R34979 DVSS.n2883 DVSS.n2881 2.2505
R34980 DVSS.n9459 DVSS.n9458 2.2505
R34981 DVSS.n2783 DVSS.n2782 2.2505
R34982 DVSS.n9464 DVSS.n9463 2.2505
R34983 DVSS.n9773 DVSS.n9772 2.2505
R34984 DVSS.n2723 DVSS.n2721 2.2505
R34985 DVSS.n10114 DVSS.n10113 2.2505
R34986 DVSS.n2705 DVSS.n2704 2.2505
R34987 DVSS.n10129 DVSS.n10128 2.2505
R34988 DVSS.n10132 DVSS.n10131 2.2505
R34989 DVSS.n2363 DVSS.n2362 2.2505
R34990 DVSS.n10154 DVSS.n10153 2.2505
R34991 DVSS.n10157 DVSS.n10156 2.2505
R34992 DVSS.n2018 DVSS.n2017 2.2505
R34993 DVSS.n10463 DVSS.n10462 2.2505
R34994 DVSS.n10466 DVSS.n10465 2.2505
R34995 DVSS.n1626 DVSS.n1625 2.2505
R34996 DVSS.n10489 DVSS.n10488 2.2505
R34997 DVSS.n10494 DVSS.n10493 2.2505
R34998 DVSS.n1521 DVSS.n1519 2.2505
R34999 DVSS.n10757 DVSS.n10756 2.2505
R35000 DVSS.n1515 DVSS.n1513 2.2505
R35001 DVSS.n13357 DVSS.n13356 2.2505
R35002 DVSS.n13352 DVSS.n13351 2.2505
R35003 DVSS.n10764 DVSS.n10763 2.2505
R35004 DVSS.n11448 DVSS.n11447 2.2505
R35005 DVSS.n13333 DVSS.n11450 2.2505
R35006 DVSS.n11455 DVSS.n11449 2.2505
R35007 DVSS.n13329 DVSS.n13328 2.2505
R35008 DVSS.n11642 DVSS.n11641 2.2505
R35009 DVSS.n11644 DVSS.n11638 2.2505
R35010 DVSS.n11984 DVSS.n11983 2.2505
R35011 DVSS.n11634 DVSS.n11632 2.2505
R35012 DVSS.n13119 DVSS.n13118 2.2505
R35013 DVSS.n11635 DVSS.n11633 2.2505
R35014 DVSS.n13113 DVSS.n13112 2.2505
R35015 DVSS.n11993 DVSS.n11991 2.2505
R35016 DVSS.n12763 DVSS.n12762 2.2505
R35017 DVSS.n12087 DVSS.n12044 2.2505
R35018 DVSS.n12090 DVSS.n12089 2.2505
R35019 DVSS.n12094 DVSS.n12093 2.2505
R35020 DVSS.n12097 DVSS.n12096 2.2505
R35021 DVSS.n12101 DVSS.n12100 2.2505
R35022 DVSS.n12098 DVSS.n12085 2.2505
R35023 DVSS.n12106 DVSS.n12105 2.2505
R35024 DVSS.n12109 DVSS.n12108 2.2505
R35025 DVSS.n12113 DVSS.n12112 2.2505
R35026 DVSS.n12110 DVSS.n12083 2.2505
R35027 DVSS.n12118 DVSS.n12117 2.2505
R35028 DVSS.n12121 DVSS.n12120 2.2505
R35029 DVSS.n12125 DVSS.n12124 2.2505
R35030 DVSS.n12122 DVSS.n12081 2.2505
R35031 DVSS.n12130 DVSS.n12129 2.2505
R35032 DVSS.n12133 DVSS.n12132 2.2505
R35033 DVSS.n12137 DVSS.n12136 2.2505
R35034 DVSS.n12134 DVSS.n12079 2.2505
R35035 DVSS.n12142 DVSS.n12141 2.2505
R35036 DVSS.n12145 DVSS.n12144 2.2505
R35037 DVSS.n12149 DVSS.n12148 2.2505
R35038 DVSS.n12146 DVSS.n12077 2.2505
R35039 DVSS.n12154 DVSS.n12153 2.2505
R35040 DVSS.n12157 DVSS.n12156 2.2505
R35041 DVSS.n12161 DVSS.n12160 2.2505
R35042 DVSS.n12158 DVSS.n12075 2.2505
R35043 DVSS.n12166 DVSS.n12165 2.2505
R35044 DVSS.n12169 DVSS.n12168 2.2505
R35045 DVSS.n12173 DVSS.n12172 2.2505
R35046 DVSS.n12170 DVSS.n12073 2.2505
R35047 DVSS.n12178 DVSS.n12177 2.2505
R35048 DVSS.n12181 DVSS.n12180 2.2505
R35049 DVSS.n12185 DVSS.n12184 2.2505
R35050 DVSS.n12182 DVSS.n12071 2.2505
R35051 DVSS.n12190 DVSS.n12189 2.2505
R35052 DVSS.n12193 DVSS.n12192 2.2505
R35053 DVSS.n12197 DVSS.n12196 2.2505
R35054 DVSS.n12194 DVSS.n12069 2.2505
R35055 DVSS.n12202 DVSS.n12201 2.2505
R35056 DVSS.n12205 DVSS.n12204 2.2505
R35057 DVSS.n12209 DVSS.n12208 2.2505
R35058 DVSS.n12206 DVSS.n12067 2.2505
R35059 DVSS.n12214 DVSS.n12213 2.2505
R35060 DVSS.n12217 DVSS.n12216 2.2505
R35061 DVSS.n12221 DVSS.n12220 2.2505
R35062 DVSS.n12218 DVSS.n12065 2.2505
R35063 DVSS.n12226 DVSS.n12225 2.2505
R35064 DVSS.n12229 DVSS.n12228 2.2505
R35065 DVSS.n12233 DVSS.n12232 2.2505
R35066 DVSS.n12230 DVSS.n12063 2.2505
R35067 DVSS.n12238 DVSS.n12237 2.2505
R35068 DVSS.n12241 DVSS.n12240 2.2505
R35069 DVSS.n12245 DVSS.n12244 2.2505
R35070 DVSS.n12242 DVSS.n12061 2.2505
R35071 DVSS.n12250 DVSS.n12249 2.2505
R35072 DVSS.n12253 DVSS.n12252 2.2505
R35073 DVSS.n12257 DVSS.n12256 2.2505
R35074 DVSS.n12254 DVSS.n12059 2.2505
R35075 DVSS.n12262 DVSS.n12261 2.2505
R35076 DVSS.n12265 DVSS.n12264 2.2505
R35077 DVSS.n12269 DVSS.n12268 2.2505
R35078 DVSS.n12266 DVSS.n12057 2.2505
R35079 DVSS.n12274 DVSS.n12273 2.2505
R35080 DVSS.n12277 DVSS.n12276 2.2505
R35081 DVSS.n12281 DVSS.n12280 2.2505
R35082 DVSS.n12278 DVSS.n12055 2.2505
R35083 DVSS.n12286 DVSS.n12285 2.2505
R35084 DVSS.n12289 DVSS.n12288 2.2505
R35085 DVSS.n12293 DVSS.n12292 2.2505
R35086 DVSS.n12290 DVSS.n12053 2.2505
R35087 DVSS.n12298 DVSS.n12297 2.2505
R35088 DVSS.n12301 DVSS.n12300 2.2505
R35089 DVSS.n12305 DVSS.n12304 2.2505
R35090 DVSS.n12302 DVSS.n12051 2.2505
R35091 DVSS.n12310 DVSS.n12309 2.2505
R35092 DVSS.n12313 DVSS.n12312 2.2505
R35093 DVSS.n12317 DVSS.n12316 2.2505
R35094 DVSS.n12314 DVSS.n12049 2.2505
R35095 DVSS.n12322 DVSS.n12321 2.2505
R35096 DVSS.n12325 DVSS.n12324 2.2505
R35097 DVSS.n12329 DVSS.n12328 2.2505
R35098 DVSS.n12326 DVSS.n12046 2.2505
R35099 DVSS.n12333 DVSS.n12047 2.2505
R35100 DVSS.n12335 DVSS.n12334 2.2505
R35101 DVSS.n12334 DVSS.n11988 2.2505
R35102 DVSS.n12333 DVSS.n12332 2.2505
R35103 DVSS.n12331 DVSS.n12046 2.2505
R35104 DVSS.n12330 DVSS.n12329 2.2505
R35105 DVSS.n12325 DVSS.n12048 2.2505
R35106 DVSS.n12321 DVSS.n12320 2.2505
R35107 DVSS.n12319 DVSS.n12049 2.2505
R35108 DVSS.n12318 DVSS.n12317 2.2505
R35109 DVSS.n12313 DVSS.n12050 2.2505
R35110 DVSS.n12309 DVSS.n12308 2.2505
R35111 DVSS.n12307 DVSS.n12051 2.2505
R35112 DVSS.n12306 DVSS.n12305 2.2505
R35113 DVSS.n12301 DVSS.n12052 2.2505
R35114 DVSS.n12297 DVSS.n12296 2.2505
R35115 DVSS.n12295 DVSS.n12053 2.2505
R35116 DVSS.n12294 DVSS.n12293 2.2505
R35117 DVSS.n12289 DVSS.n12054 2.2505
R35118 DVSS.n12285 DVSS.n12284 2.2505
R35119 DVSS.n12283 DVSS.n12055 2.2505
R35120 DVSS.n12282 DVSS.n12281 2.2505
R35121 DVSS.n12277 DVSS.n12056 2.2505
R35122 DVSS.n12273 DVSS.n12272 2.2505
R35123 DVSS.n12271 DVSS.n12057 2.2505
R35124 DVSS.n12270 DVSS.n12269 2.2505
R35125 DVSS.n12265 DVSS.n12058 2.2505
R35126 DVSS.n12261 DVSS.n12260 2.2505
R35127 DVSS.n12259 DVSS.n12059 2.2505
R35128 DVSS.n12258 DVSS.n12257 2.2505
R35129 DVSS.n12253 DVSS.n12060 2.2505
R35130 DVSS.n12249 DVSS.n12248 2.2505
R35131 DVSS.n12247 DVSS.n12061 2.2505
R35132 DVSS.n12246 DVSS.n12245 2.2505
R35133 DVSS.n12241 DVSS.n12062 2.2505
R35134 DVSS.n12237 DVSS.n12236 2.2505
R35135 DVSS.n12235 DVSS.n12063 2.2505
R35136 DVSS.n12234 DVSS.n12233 2.2505
R35137 DVSS.n12229 DVSS.n12064 2.2505
R35138 DVSS.n12225 DVSS.n12224 2.2505
R35139 DVSS.n12223 DVSS.n12065 2.2505
R35140 DVSS.n12222 DVSS.n12221 2.2505
R35141 DVSS.n12217 DVSS.n12066 2.2505
R35142 DVSS.n12213 DVSS.n12212 2.2505
R35143 DVSS.n12211 DVSS.n12067 2.2505
R35144 DVSS.n12210 DVSS.n12209 2.2505
R35145 DVSS.n12205 DVSS.n12068 2.2505
R35146 DVSS.n12201 DVSS.n12200 2.2505
R35147 DVSS.n12199 DVSS.n12069 2.2505
R35148 DVSS.n12198 DVSS.n12197 2.2505
R35149 DVSS.n12193 DVSS.n12070 2.2505
R35150 DVSS.n12189 DVSS.n12188 2.2505
R35151 DVSS.n12187 DVSS.n12071 2.2505
R35152 DVSS.n12186 DVSS.n12185 2.2505
R35153 DVSS.n12181 DVSS.n12072 2.2505
R35154 DVSS.n12177 DVSS.n12176 2.2505
R35155 DVSS.n12175 DVSS.n12073 2.2505
R35156 DVSS.n12174 DVSS.n12173 2.2505
R35157 DVSS.n12169 DVSS.n12074 2.2505
R35158 DVSS.n12165 DVSS.n12164 2.2505
R35159 DVSS.n12163 DVSS.n12075 2.2505
R35160 DVSS.n12162 DVSS.n12161 2.2505
R35161 DVSS.n12157 DVSS.n12076 2.2505
R35162 DVSS.n12153 DVSS.n12152 2.2505
R35163 DVSS.n12151 DVSS.n12077 2.2505
R35164 DVSS.n12150 DVSS.n12149 2.2505
R35165 DVSS.n12145 DVSS.n12078 2.2505
R35166 DVSS.n12141 DVSS.n12140 2.2505
R35167 DVSS.n12139 DVSS.n12079 2.2505
R35168 DVSS.n12138 DVSS.n12137 2.2505
R35169 DVSS.n12133 DVSS.n12080 2.2505
R35170 DVSS.n12129 DVSS.n12128 2.2505
R35171 DVSS.n12127 DVSS.n12081 2.2505
R35172 DVSS.n12126 DVSS.n12125 2.2505
R35173 DVSS.n12121 DVSS.n12082 2.2505
R35174 DVSS.n12117 DVSS.n12116 2.2505
R35175 DVSS.n12115 DVSS.n12083 2.2505
R35176 DVSS.n12114 DVSS.n12113 2.2505
R35177 DVSS.n12109 DVSS.n12084 2.2505
R35178 DVSS.n12105 DVSS.n12104 2.2505
R35179 DVSS.n12103 DVSS.n12085 2.2505
R35180 DVSS.n12102 DVSS.n12101 2.2505
R35181 DVSS.n12097 DVSS.n12086 2.2505
R35182 DVSS.n12093 DVSS.n12092 2.2505
R35183 DVSS.n12091 DVSS.n12090 2.2505
R35184 DVSS.n12087 DVSS.n12000 2.2505
R35185 DVSS.n6674 DVSS.n6673 2.2505
R35186 DVSS.n6675 DVSS.n6233 2.2505
R35187 DVSS.n6677 DVSS.n6676 2.2505
R35188 DVSS.n6692 DVSS.n6691 2.2505
R35189 DVSS.n6693 DVSS.n5883 2.2505
R35190 DVSS.n7031 DVSS.n7030 2.2505
R35191 DVSS.n7028 DVSS.n5865 2.2505
R35192 DVSS.n7047 DVSS.n5864 2.2505
R35193 DVSS.n7051 DVSS.n7050 2.2505
R35194 DVSS.n5523 DVSS.n5522 2.2505
R35195 DVSS.n7072 DVSS.n7071 2.2505
R35196 DVSS.n7076 DVSS.n7075 2.2505
R35197 DVSS.n7074 DVSS.n5174 2.2505
R35198 DVSS.n7090 DVSS.n5173 2.2505
R35199 DVSS.n7094 DVSS.n7093 2.2505
R35200 DVSS.n4830 DVSS.n4829 2.2505
R35201 DVSS.n7455 DVSS.n7454 2.2505
R35202 DVSS.n7458 DVSS.n7457 2.2505
R35203 DVSS.n4816 DVSS.n4815 2.2505
R35204 DVSS.n7810 DVSS.n7809 2.2505
R35205 DVSS.n7813 DVSS.n7812 2.2505
R35206 DVSS.n4464 DVSS.n4463 2.2505
R35207 DVSS.n7830 DVSS.n7829 2.2505
R35208 DVSS.n7832 DVSS.n4461 2.2505
R35209 DVSS.n7834 DVSS.n7833 2.2505
R35210 DVSS.n7838 DVSS.n7837 2.2505
R35211 DVSS.n4360 DVSS.n4359 2.2505
R35212 DVSS.n8106 DVSS.n8105 2.2505
R35213 DVSS.n8109 DVSS.n8108 2.2505
R35214 DVSS.n3854 DVSS.n3853 2.2505
R35215 DVSS.n8324 DVSS.n8323 2.2505
R35216 DVSS.n8326 DVSS.n3850 2.2505
R35217 DVSS.n8329 DVSS.n8328 2.2505
R35218 DVSS.n8327 DVSS.n3851 2.2505
R35219 DVSS.n8593 DVSS.n8592 2.2505
R35220 DVSS.n8594 DVSS.n3749 2.2505
R35221 DVSS.n8597 DVSS.n8596 2.2505
R35222 DVSS.n3404 DVSS.n3403 2.2505
R35223 DVSS.n8619 DVSS.n8618 2.2505
R35224 DVSS.n8622 DVSS.n8621 2.2505
R35225 DVSS.n3057 DVSS.n3056 2.2505
R35226 DVSS.n8973 DVSS.n8972 2.2505
R35227 DVSS.n8976 DVSS.n8975 2.2505
R35228 DVSS.n2886 DVSS.n2885 2.2505
R35229 DVSS.n9191 DVSS.n9190 2.2505
R35230 DVSS.n9193 DVSS.n2882 2.2505
R35231 DVSS.n9196 DVSS.n9195 2.2505
R35232 DVSS.n9194 DVSS.n2883 2.2505
R35233 DVSS.n9460 DVSS.n9459 2.2505
R35234 DVSS.n9461 DVSS.n2783 2.2505
R35235 DVSS.n9463 DVSS.n9462 2.2505
R35236 DVSS.n9774 DVSS.n9773 2.2505
R35237 DVSS.n9775 DVSS.n2723 2.2505
R35238 DVSS.n10113 DVSS.n10112 2.2505
R35239 DVSS.n10110 DVSS.n2704 2.2505
R35240 DVSS.n10129 DVSS.n2702 2.2505
R35241 DVSS.n10133 DVSS.n10132 2.2505
R35242 DVSS.n2703 DVSS.n2362 2.2505
R35243 DVSS.n10154 DVSS.n2360 2.2505
R35244 DVSS.n10158 DVSS.n10157 2.2505
R35245 DVSS.n2361 DVSS.n2017 2.2505
R35246 DVSS.n10463 DVSS.n2016 2.2505
R35247 DVSS.n10467 DVSS.n10466 2.2505
R35248 DVSS.n1625 DVSS.n1624 2.2505
R35249 DVSS.n10490 DVSS.n10489 2.2505
R35250 DVSS.n10493 DVSS.n10492 2.2505
R35251 DVSS.n1519 DVSS.n1518 2.2505
R35252 DVSS.n10758 DVSS.n10757 2.2505
R35253 DVSS.n10760 DVSS.n1515 2.2505
R35254 DVSS.n13356 DVSS.n13355 2.2505
R35255 DVSS.n13353 DVSS.n13352 2.2505
R35256 DVSS.n10763 DVSS.n10762 2.2505
R35257 DVSS.n11451 DVSS.n11448 2.2505
R35258 DVSS.n13333 DVSS.n13332 2.2505
R35259 DVSS.n13331 DVSS.n11449 2.2505
R35260 DVSS.n13330 DVSS.n13329 2.2505
R35261 DVSS.n11641 DVSS.n11640 2.2505
R35262 DVSS.n11638 DVSS.n11637 2.2505
R35263 DVSS.n11985 DVSS.n11984 2.2505
R35264 DVSS.n11987 DVSS.n11634 2.2505
R35265 DVSS.n13118 DVSS.n13117 2.2505
R35266 DVSS.n13116 DVSS.n11635 2.2505
R35267 DVSS.n13114 DVSS.n13113 2.2505
R35268 DVSS.n11991 DVSS.n11989 2.2505
R35269 DVSS.n12764 DVSS.n12763 2.2505
R35270 DVSS.n21106 DVSS.n13945 2.25007
R35271 DVSS.n21106 DVSS.n13941 2.25007
R35272 DVSS.n14076 DVSS.n14031 2.25007
R35273 DVSS.n14081 DVSS.n14031 2.25007
R35274 DVSS.n13881 DVSS.n13836 2.25007
R35275 DVSS.n13886 DVSS.n13825 2.25007
R35276 DVSS.n13737 DVSS.n13629 2.25007
R35277 DVSS.n13742 DVSS.n13629 2.25007
R35278 DVSS.n14181 DVSS.n14137 2.25007
R35279 DVSS.n14186 DVSS.n14137 2.25007
R35280 DVSS.n14276 DVSS.n14275 2.25007
R35281 DVSS.n14276 DVSS.n14274 2.25007
R35282 DVSS.n12808 DVSS.n12807 2.25007
R35283 DVSS.n12808 DVSS.n12806 2.25007
R35284 DVSS.n1000 DVSS.n999 2.25007
R35285 DVSS.n1000 DVSS.n998 2.25007
R35286 DVSS.n1082 DVSS.n1081 2.25007
R35287 DVSS.n1100 DVSS.n1078 2.25007
R35288 DVSS.n1136 DVSS.n1135 2.25007
R35289 DVSS.n1154 DVSS.n1136 2.25007
R35290 DVSS.n13006 DVSS.n13005 2.25007
R35291 DVSS.n13006 DVSS.n13004 2.25007
R35292 DVSS.n385 DVSS.n349 2.25007
R35293 DVSS.n392 DVSS.n349 2.25007
R35294 DVSS.n23218 DVSS.n16 2.25007
R35295 DVSS.n39 DVSS.n16 2.25007
R35296 DVSS.n913 DVSS.n912 2.25007
R35297 DVSS.n913 DVSS.n911 2.25007
R35298 DVSS.n22486 DVSS.n813 2.25007
R35299 DVSS.n22501 DVSS.n813 2.25007
R35300 DVSS.n248 DVSS.n217 2.25007
R35301 DVSS.n254 DVSS.n217 2.25007
R35302 DVSS.n168 DVSS.n137 2.25007
R35303 DVSS.n174 DVSS.n137 2.25007
R35304 DVSS.n102 DVSS.n72 2.25007
R35305 DVSS.n107 DVSS.n72 2.25007
R35306 DVSS.n1251 DVSS.n1250 2.25007
R35307 DVSS.n1251 DVSS.n1249 2.25007
R35308 DVSS.n1391 DVSS.n1390 2.25007
R35309 DVSS.n1391 DVSS.n1389 2.25007
R35310 DVSS.n21863 DVSS.n870 2.25007
R35311 DVSS.n21922 DVSS.n21880 2.25007
R35312 DVSS.n21631 DVSS.n21590 2.25007
R35313 DVSS.n21635 DVSS.n21590 2.25007
R35314 DVSS.n21735 DVSS.n1178 2.25007
R35315 DVSS.n21740 DVSS.n1178 2.25007
R35316 DVSS.n21951 DVSS.n1199 2.25007
R35317 DVSS.n21958 DVSS.n1199 2.25007
R35318 DVSS.n21584 DVSS.n21568 2.24982
R35319 DVSS.n20027 DVSS.n20010 2.24982
R35320 DVSS.n20166 DVSS.n14585 2.24982
R35321 DVSS.n17359 DVSS.n17358 2.24982
R35322 DVSS.n17272 DVSS.n17260 2.24982
R35323 DVSS.n17171 DVSS.n17140 2.24982
R35324 DVSS.n17169 DVSS.n17141 2.24982
R35325 DVSS.n17271 DVSS.n17261 2.24982
R35326 DVSS.n1188 DVSS.n1179 2.24982
R35327 DVSS.n20194 DVSS.n14865 2.24982
R35328 DVSS.n14650 DVSS.n14633 2.24982
R35329 DVSS.n16951 DVSS.n16941 2.24982
R35330 DVSS.n17237 DVSS.n17225 2.24982
R35331 DVSS.n17197 DVSS.n17175 2.24982
R35332 DVSS.n17459 DVSS.n17458 2.24982
R35333 DVSS.n17236 DVSS.n17226 2.24982
R35334 DVSS.n868 DVSS.n858 2.24982
R35335 DVSS.n18922 DVSS.n14517 2.24982
R35336 DVSS.n18975 DVSS.n14550 2.24982
R35337 DVSS.n17327 DVSS.n17326 2.24982
R35338 DVSS.n17387 DVSS.n17303 2.24982
R35339 DVSS.n17136 DVSS.n17121 2.24982
R35340 DVSS.n17295 DVSS.n17294 2.24982
R35341 DVSS.n17386 DVSS.n17304 2.24982
R35342 DVSS.n19503 DVSS.n19269 2.24982
R35343 DVSS.n19252 DVSS.n19251 2.24982
R35344 DVSS.n19079 DVSS.n19069 2.24982
R35345 DVSS.n19031 DVSS.n19021 2.24982
R35346 DVSS.n19170 DVSS.n19169 2.24982
R35347 DVSS.n19158 DVSS.n19156 2.24982
R35348 DVSS.n19897 DVSS.n19004 2.24982
R35349 DVSS.n19246 DVSS.n19216 2.24982
R35350 DVSS.n19620 DVSS.n19161 2.24982
R35351 DVSS.n1044 DVSS.n1042 2.24982
R35352 DVSS.n1174 DVSS.n1165 2.24982
R35353 DVSS.n12960 DVSS.n12958 2.24982
R35354 DVSS.n13092 DVSS.n13091 2.24982
R35355 DVSS.n19143 DVSS.n19141 2.24982
R35356 DVSS.n19648 DVSS.n19148 2.24982
R35357 DVSS.n1209 DVSS.n1200 2.24982
R35358 DVSS.n19100 DVSS.n19091 2.24982
R35359 DVSS.n20333 DVSS.n14854 2.24982
R35360 DVSS.n20451 DVSS.n20450 2.24982
R35361 DVSS.n17453 DVSS.n17434 2.24982
R35362 DVSS.n16937 DVSS.n16935 2.24982
R35363 DVSS.n17207 DVSS.n17199 2.24982
R35364 DVSS.n17445 DVSS.n17444 2.24982
R35365 DVSS.n17419 DVSS.n17210 2.24982
R35366 DVSS.n19314 DVSS.n19310 2.24972
R35367 DVSS.n19315 DVSS.n19309 2.24972
R35368 DVSS.n19656 DVSS.n19655 2.24972
R35369 DVSS.n19657 DVSS.n19140 2.24972
R35370 DVSS.n20049 DVSS.n20048 2.24964
R35371 DVSS.n20047 DVSS.n20040 2.24964
R35372 DVSS.n13533 DVSS.n13528 2.24964
R35373 DVSS.n13553 DVSS.n13552 2.24964
R35374 DVSS.n13533 DVSS.n13529 2.24964
R35375 DVSS.n13553 DVSS.n13551 2.24964
R35376 DVSS.n13533 DVSS.n13530 2.24964
R35377 DVSS.n13553 DVSS.n13550 2.24964
R35378 DVSS.n13533 DVSS.n13531 2.24964
R35379 DVSS.n13553 DVSS.n13549 2.24964
R35380 DVSS.n13533 DVSS.n13532 2.24964
R35381 DVSS.n13553 DVSS.n13534 2.24964
R35382 DVSS.n21096 DVSS.n13940 2.24964
R35383 DVSS.n21107 DVSS.n13938 2.24964
R35384 DVSS.n21096 DVSS.n21095 2.24964
R35385 DVSS.n21107 DVSS.n13937 2.24964
R35386 DVSS.n21096 DVSS.n21094 2.24964
R35387 DVSS.n21107 DVSS.n13936 2.24964
R35388 DVSS.n21096 DVSS.n21093 2.24964
R35389 DVSS.n21107 DVSS.n13935 2.24964
R35390 DVSS.n21096 DVSS.n21092 2.24964
R35391 DVSS.n21107 DVSS.n13934 2.24964
R35392 DVSS.n21096 DVSS.n21091 2.24964
R35393 DVSS.n21107 DVSS.n13933 2.24964
R35394 DVSS.n21096 DVSS.n21090 2.24964
R35395 DVSS.n21107 DVSS.n13932 2.24964
R35396 DVSS.n21096 DVSS.n21089 2.24964
R35397 DVSS.n21107 DVSS.n13931 2.24964
R35398 DVSS.n21096 DVSS.n21088 2.24964
R35399 DVSS.n21107 DVSS.n13930 2.24964
R35400 DVSS.n21096 DVSS.n21087 2.24964
R35401 DVSS.n21107 DVSS.n13929 2.24964
R35402 DVSS.n21096 DVSS.n13976 2.24964
R35403 DVSS.n21107 DVSS.n13928 2.24964
R35404 DVSS.n14475 DVSS.n14471 2.24964
R35405 DVSS.n20818 DVSS.n20817 2.24964
R35406 DVSS.n14475 DVSS.n14472 2.24964
R35407 DVSS.n20818 DVSS.n20816 2.24964
R35408 DVSS.n14475 DVSS.n14473 2.24964
R35409 DVSS.n20818 DVSS.n20815 2.24964
R35410 DVSS.n14475 DVSS.n14474 2.24964
R35411 DVSS.n20818 DVSS.n14482 2.24964
R35412 DVSS.n14908 DVSS.n14875 2.24964
R35413 DVSS.n14895 DVSS.n14882 2.24964
R35414 DVSS.n14908 DVSS.n14904 2.24964
R35415 DVSS.n14897 DVSS.n14882 2.24964
R35416 DVSS.n14908 DVSS.n14905 2.24964
R35417 DVSS.n14899 DVSS.n14882 2.24964
R35418 DVSS.n14908 DVSS.n14906 2.24964
R35419 DVSS.n14901 DVSS.n14882 2.24964
R35420 DVSS.n14908 DVSS.n14907 2.24964
R35421 DVSS.n14911 DVSS.n14882 2.24964
R35422 DVSS.n15296 DVSS.n15286 2.24964
R35423 DVSS.n15309 DVSS.n15307 2.24964
R35424 DVSS.n15301 DVSS.n15286 2.24964
R35425 DVSS.n15309 DVSS.n15308 2.24964
R35426 DVSS.n15303 DVSS.n15286 2.24964
R35427 DVSS.n16099 DVSS.n16074 2.24964
R35428 DVSS.n17644 DVSS.n16072 2.24964
R35429 DVSS.n16099 DVSS.n16098 2.24964
R35430 DVSS.n17644 DVSS.n16071 2.24964
R35431 DVSS.n16099 DVSS.n16097 2.24964
R35432 DVSS.n16101 DVSS.n16100 2.24964
R35433 DVSS.n17644 DVSS.n16069 2.24964
R35434 DVSS.n16255 DVSS.n16254 2.24964
R35435 DVSS.n16266 DVSS.n16265 2.24964
R35436 DVSS.n16255 DVSS.n16253 2.24964
R35437 DVSS.n16266 DVSS.n16264 2.24964
R35438 DVSS.n16255 DVSS.n16252 2.24964
R35439 DVSS.n16266 DVSS.n16263 2.24964
R35440 DVSS.n15800 DVSS.n15799 2.24964
R35441 DVSS.n15811 DVSS.n15810 2.24964
R35442 DVSS.n15800 DVSS.n15798 2.24964
R35443 DVSS.n15811 DVSS.n15809 2.24964
R35444 DVSS.n15800 DVSS.n15797 2.24964
R35445 DVSS.n15811 DVSS.n15808 2.24964
R35446 DVSS.n15800 DVSS.n15796 2.24964
R35447 DVSS.n15811 DVSS.n15807 2.24964
R35448 DVSS.n16266 DVSS.n16262 2.24964
R35449 DVSS.n17644 DVSS.n16068 2.24964
R35450 DVSS.n15299 DVSS.n15286 2.24964
R35451 DVSS.n20300 DVSS.n20213 2.24964
R35452 DVSS.n20305 DVSS.n20304 2.24964
R35453 DVSS.n13471 DVSS.n13465 2.24964
R35454 DVSS.n13501 DVSS.n13500 2.24964
R35455 DVSS.n13473 DVSS.n13465 2.24964
R35456 DVSS.n13501 DVSS.n13499 2.24964
R35457 DVSS.n13475 DVSS.n13465 2.24964
R35458 DVSS.n13501 DVSS.n13498 2.24964
R35459 DVSS.n13477 DVSS.n13465 2.24964
R35460 DVSS.n13501 DVSS.n13497 2.24964
R35461 DVSS.n13479 DVSS.n13465 2.24964
R35462 DVSS.n13501 DVSS.n13482 2.24964
R35463 DVSS.n14056 DVSS.n14055 2.24964
R35464 DVSS.n14068 DVSS.n14057 2.24964
R35465 DVSS.n14056 DVSS.n14054 2.24964
R35466 DVSS.n14068 DVSS.n14058 2.24964
R35467 DVSS.n14056 DVSS.n14053 2.24964
R35468 DVSS.n14068 DVSS.n14059 2.24964
R35469 DVSS.n14056 DVSS.n14052 2.24964
R35470 DVSS.n14068 DVSS.n14060 2.24964
R35471 DVSS.n14056 DVSS.n14051 2.24964
R35472 DVSS.n14068 DVSS.n14061 2.24964
R35473 DVSS.n14056 DVSS.n14050 2.24964
R35474 DVSS.n14068 DVSS.n14062 2.24964
R35475 DVSS.n14056 DVSS.n14049 2.24964
R35476 DVSS.n14068 DVSS.n14063 2.24964
R35477 DVSS.n14056 DVSS.n14048 2.24964
R35478 DVSS.n14068 DVSS.n14064 2.24964
R35479 DVSS.n14056 DVSS.n14047 2.24964
R35480 DVSS.n14068 DVSS.n14065 2.24964
R35481 DVSS.n14056 DVSS.n14046 2.24964
R35482 DVSS.n14068 DVSS.n14066 2.24964
R35483 DVSS.n14056 DVSS.n14045 2.24964
R35484 DVSS.n14068 DVSS.n14067 2.24964
R35485 DVSS.n14417 DVSS.n14410 2.24964
R35486 DVSS.n14444 DVSS.n14443 2.24964
R35487 DVSS.n14419 DVSS.n14410 2.24964
R35488 DVSS.n14444 DVSS.n14442 2.24964
R35489 DVSS.n14421 DVSS.n14410 2.24964
R35490 DVSS.n14444 DVSS.n14441 2.24964
R35491 DVSS.n14423 DVSS.n14410 2.24964
R35492 DVSS.n14444 DVSS.n14426 2.24964
R35493 DVSS.n14944 DVSS.n14939 2.24964
R35494 DVSS.n14992 DVSS.n14991 2.24964
R35495 DVSS.n14944 DVSS.n14940 2.24964
R35496 DVSS.n14992 DVSS.n14990 2.24964
R35497 DVSS.n14944 DVSS.n14941 2.24964
R35498 DVSS.n14992 DVSS.n14989 2.24964
R35499 DVSS.n14944 DVSS.n14942 2.24964
R35500 DVSS.n14992 DVSS.n14988 2.24964
R35501 DVSS.n14944 DVSS.n14943 2.24964
R35502 DVSS.n14992 DVSS.n14945 2.24964
R35503 DVSS.n15377 DVSS.n15374 2.24964
R35504 DVSS.n15377 DVSS.n15375 2.24964
R35505 DVSS.n15381 DVSS.n15380 2.24964
R35506 DVSS.n15377 DVSS.n15376 2.24964
R35507 DVSS.n15381 DVSS.n15379 2.24964
R35508 DVSS.n16832 DVSS.n16830 2.24964
R35509 DVSS.n16837 DVSS.n16835 2.24964
R35510 DVSS.n16832 DVSS.n16831 2.24964
R35511 DVSS.n16837 DVSS.n16834 2.24964
R35512 DVSS.n16832 DVSS.n16829 2.24964
R35513 DVSS.n16837 DVSS.n16836 2.24964
R35514 DVSS.n16832 DVSS.n16828 2.24964
R35515 DVSS.n16179 DVSS.n16152 2.24964
R35516 DVSS.n16184 DVSS.n16180 2.24964
R35517 DVSS.n16179 DVSS.n16178 2.24964
R35518 DVSS.n16184 DVSS.n16181 2.24964
R35519 DVSS.n16179 DVSS.n16177 2.24964
R35520 DVSS.n16184 DVSS.n16182 2.24964
R35521 DVSS.n15744 DVSS.n15738 2.24964
R35522 DVSS.n15756 DVSS.n15752 2.24964
R35523 DVSS.n15746 DVSS.n15738 2.24964
R35524 DVSS.n15756 DVSS.n15753 2.24964
R35525 DVSS.n15748 DVSS.n15738 2.24964
R35526 DVSS.n15756 DVSS.n15754 2.24964
R35527 DVSS.n15750 DVSS.n15738 2.24964
R35528 DVSS.n15756 DVSS.n15755 2.24964
R35529 DVSS.n16184 DVSS.n16183 2.24964
R35530 DVSS.n16837 DVSS.n16833 2.24964
R35531 DVSS.n15381 DVSS.n15378 2.24964
R35532 DVSS.n18915 DVSS.n18874 2.24964
R35533 DVSS.n18876 DVSS.n18875 2.24964
R35534 DVSS.n13591 DVSS.n13590 2.24964
R35535 DVSS.n13601 DVSS.n13600 2.24964
R35536 DVSS.n13601 DVSS.n13599 2.24964
R35537 DVSS.n13591 DVSS.n13589 2.24964
R35538 DVSS.n13601 DVSS.n13598 2.24964
R35539 DVSS.n13591 DVSS.n13588 2.24964
R35540 DVSS.n13601 DVSS.n13597 2.24964
R35541 DVSS.n13584 DVSS.n13583 2.24964
R35542 DVSS.n13582 DVSS.n13570 2.24964
R35543 DVSS.n13861 DVSS.n13860 2.24964
R35544 DVSS.n13873 DVSS.n13862 2.24964
R35545 DVSS.n13861 DVSS.n13859 2.24964
R35546 DVSS.n13873 DVSS.n13863 2.24964
R35547 DVSS.n13861 DVSS.n13858 2.24964
R35548 DVSS.n13873 DVSS.n13864 2.24964
R35549 DVSS.n13861 DVSS.n13857 2.24964
R35550 DVSS.n13873 DVSS.n13865 2.24964
R35551 DVSS.n13861 DVSS.n13856 2.24964
R35552 DVSS.n13873 DVSS.n13866 2.24964
R35553 DVSS.n13861 DVSS.n13855 2.24964
R35554 DVSS.n13873 DVSS.n13867 2.24964
R35555 DVSS.n13861 DVSS.n13854 2.24964
R35556 DVSS.n13873 DVSS.n13868 2.24964
R35557 DVSS.n13861 DVSS.n13853 2.24964
R35558 DVSS.n13873 DVSS.n13869 2.24964
R35559 DVSS.n13861 DVSS.n13852 2.24964
R35560 DVSS.n13873 DVSS.n13870 2.24964
R35561 DVSS.n13861 DVSS.n13851 2.24964
R35562 DVSS.n13873 DVSS.n13871 2.24964
R35563 DVSS.n13861 DVSS.n13850 2.24964
R35564 DVSS.n13873 DVSS.n13872 2.24964
R35565 DVSS.n20704 DVSS.n20700 2.24964
R35566 DVSS.n20722 DVSS.n20721 2.24964
R35567 DVSS.n20704 DVSS.n20701 2.24964
R35568 DVSS.n20722 DVSS.n20720 2.24964
R35569 DVSS.n20704 DVSS.n20702 2.24964
R35570 DVSS.n20722 DVSS.n20719 2.24964
R35571 DVSS.n20704 DVSS.n20703 2.24964
R35572 DVSS.n20722 DVSS.n20705 2.24964
R35573 DVSS.n18399 DVSS.n18394 2.24964
R35574 DVSS.n18432 DVSS.n18431 2.24964
R35575 DVSS.n18399 DVSS.n18395 2.24964
R35576 DVSS.n18432 DVSS.n18430 2.24964
R35577 DVSS.n18399 DVSS.n18396 2.24964
R35578 DVSS.n18432 DVSS.n18429 2.24964
R35579 DVSS.n18399 DVSS.n18397 2.24964
R35580 DVSS.n18432 DVSS.n18428 2.24964
R35581 DVSS.n18399 DVSS.n18398 2.24964
R35582 DVSS.n18432 DVSS.n18382 2.24964
R35583 DVSS.n15271 DVSS.n15239 2.24964
R35584 DVSS.n15271 DVSS.n15269 2.24964
R35585 DVSS.n15262 DVSS.n15240 2.24964
R35586 DVSS.n15271 DVSS.n15270 2.24964
R35587 DVSS.n15264 DVSS.n15240 2.24964
R35588 DVSS.n16010 DVSS.n16008 2.24964
R35589 DVSS.n16015 DVSS.n16013 2.24964
R35590 DVSS.n16010 DVSS.n16009 2.24964
R35591 DVSS.n16015 DVSS.n16012 2.24964
R35592 DVSS.n16010 DVSS.n16007 2.24964
R35593 DVSS.n16015 DVSS.n16014 2.24964
R35594 DVSS.n16010 DVSS.n16006 2.24964
R35595 DVSS.n16298 DVSS.n16292 2.24964
R35596 DVSS.n16306 DVSS.n16305 2.24964
R35597 DVSS.n15844 DVSS.n15836 2.24964
R35598 DVSS.n15850 DVSS.n15849 2.24964
R35599 DVSS.n15846 DVSS.n15836 2.24964
R35600 DVSS.n16015 DVSS.n16011 2.24964
R35601 DVSS.n15260 DVSS.n15240 2.24964
R35602 DVSS.n20337 DVSS.n14678 2.24964
R35603 DVSS.n14680 DVSS.n14679 2.24964
R35604 DVSS.n13436 DVSS.n13434 2.24964
R35605 DVSS.n21382 DVSS.n21380 2.24964
R35606 DVSS.n21382 DVSS.n21379 2.24964
R35607 DVSS.n13436 DVSS.n13433 2.24964
R35608 DVSS.n21382 DVSS.n21378 2.24964
R35609 DVSS.n13436 DVSS.n13432 2.24964
R35610 DVSS.n21382 DVSS.n21377 2.24964
R35611 DVSS.n13436 DVSS.n13435 2.24964
R35612 DVSS.n13431 DVSS.n13419 2.24964
R35613 DVSS.n14162 DVSS.n14161 2.24964
R35614 DVSS.n14174 DVSS.n14163 2.24964
R35615 DVSS.n14162 DVSS.n14160 2.24964
R35616 DVSS.n14174 DVSS.n14164 2.24964
R35617 DVSS.n14162 DVSS.n14159 2.24964
R35618 DVSS.n14174 DVSS.n14165 2.24964
R35619 DVSS.n14162 DVSS.n14158 2.24964
R35620 DVSS.n14174 DVSS.n14166 2.24964
R35621 DVSS.n14162 DVSS.n14157 2.24964
R35622 DVSS.n14174 DVSS.n14167 2.24964
R35623 DVSS.n14162 DVSS.n14156 2.24964
R35624 DVSS.n14174 DVSS.n14168 2.24964
R35625 DVSS.n14162 DVSS.n14155 2.24964
R35626 DVSS.n14174 DVSS.n14169 2.24964
R35627 DVSS.n14162 DVSS.n14154 2.24964
R35628 DVSS.n14174 DVSS.n14170 2.24964
R35629 DVSS.n14162 DVSS.n14153 2.24964
R35630 DVSS.n14174 DVSS.n14171 2.24964
R35631 DVSS.n14162 DVSS.n14152 2.24964
R35632 DVSS.n14174 DVSS.n14172 2.24964
R35633 DVSS.n14162 DVSS.n14151 2.24964
R35634 DVSS.n14174 DVSS.n14173 2.24964
R35635 DVSS.n14368 DVSS.n14361 2.24964
R35636 DVSS.n14395 DVSS.n14394 2.24964
R35637 DVSS.n14370 DVSS.n14361 2.24964
R35638 DVSS.n14395 DVSS.n14393 2.24964
R35639 DVSS.n14372 DVSS.n14361 2.24964
R35640 DVSS.n14395 DVSS.n14392 2.24964
R35641 DVSS.n14374 DVSS.n14361 2.24964
R35642 DVSS.n14395 DVSS.n14377 2.24964
R35643 DVSS.n15017 DVSS.n15012 2.24964
R35644 DVSS.n15071 DVSS.n15070 2.24964
R35645 DVSS.n15017 DVSS.n15013 2.24964
R35646 DVSS.n15071 DVSS.n15069 2.24964
R35647 DVSS.n15017 DVSS.n15014 2.24964
R35648 DVSS.n15071 DVSS.n15068 2.24964
R35649 DVSS.n15017 DVSS.n15015 2.24964
R35650 DVSS.n15071 DVSS.n15067 2.24964
R35651 DVSS.n15017 DVSS.n15016 2.24964
R35652 DVSS.n15071 DVSS.n15018 2.24964
R35653 DVSS.n15456 DVSS.n15453 2.24964
R35654 DVSS.n15456 DVSS.n15454 2.24964
R35655 DVSS.n15460 DVSS.n15459 2.24964
R35656 DVSS.n15456 DVSS.n15455 2.24964
R35657 DVSS.n15460 DVSS.n15458 2.24964
R35658 DVSS.n17535 DVSS.n17533 2.24964
R35659 DVSS.n17540 DVSS.n17538 2.24964
R35660 DVSS.n17535 DVSS.n17534 2.24964
R35661 DVSS.n17540 DVSS.n17537 2.24964
R35662 DVSS.n17535 DVSS.n17532 2.24964
R35663 DVSS.n17540 DVSS.n17539 2.24964
R35664 DVSS.n17535 DVSS.n17531 2.24964
R35665 DVSS.n15674 DVSS.n15653 2.24964
R35666 DVSS.n15671 DVSS.n15654 2.24964
R35667 DVSS.n15711 DVSS.n15690 2.24964
R35668 DVSS.n15721 DVSS.n15691 2.24964
R35669 DVSS.n15720 DVSS.n15690 2.24964
R35670 DVSS.n17540 DVSS.n17536 2.24964
R35671 DVSS.n15460 DVSS.n15457 2.24964
R35672 DVSS.n654 DVSS.n648 2.24964
R35673 DVSS.n673 DVSS.n672 2.24964
R35674 DVSS.n656 DVSS.n648 2.24964
R35675 DVSS.n658 DVSS.n648 2.24964
R35676 DVSS.n673 DVSS.n671 2.24964
R35677 DVSS.n667 DVSS.n648 2.24964
R35678 DVSS.n673 DVSS.n670 2.24964
R35679 DVSS.n612 DVSS.n609 2.24964
R35680 DVSS.n616 DVSS.n615 2.24964
R35681 DVSS.n612 DVSS.n610 2.24964
R35682 DVSS.n612 DVSS.n611 2.24964
R35683 DVSS.n616 DVSS.n614 2.24964
R35684 DVSS.n612 DVSS.n608 2.24964
R35685 DVSS.n616 DVSS.n613 2.24964
R35686 DVSS.n553 DVSS.n547 2.24964
R35687 DVSS.n566 DVSS.n565 2.24964
R35688 DVSS.n555 DVSS.n547 2.24964
R35689 DVSS.n557 DVSS.n547 2.24964
R35690 DVSS.n566 DVSS.n564 2.24964
R35691 DVSS.n560 DVSS.n547 2.24964
R35692 DVSS.n566 DVSS.n563 2.24964
R35693 DVSS.n512 DVSS.n509 2.24964
R35694 DVSS.n516 DVSS.n515 2.24964
R35695 DVSS.n512 DVSS.n510 2.24964
R35696 DVSS.n512 DVSS.n511 2.24964
R35697 DVSS.n516 DVSS.n514 2.24964
R35698 DVSS.n512 DVSS.n508 2.24964
R35699 DVSS.n516 DVSS.n513 2.24964
R35700 DVSS.n1106 DVSS.n1052 2.24964
R35701 DVSS.n1106 DVSS.n1103 2.24964
R35702 DVSS.n1084 DVSS.n1053 2.24964
R35703 DVSS.n1106 DVSS.n1104 2.24964
R35704 DVSS.n1087 DVSS.n1053 2.24964
R35705 DVSS.n1106 DVSS.n1102 2.24964
R35706 DVSS.n1089 DVSS.n1053 2.24964
R35707 DVSS.n1106 DVSS.n1105 2.24964
R35708 DVSS.n1092 DVSS.n1053 2.24964
R35709 DVSS.n1106 DVSS.n1101 2.24964
R35710 DVSS.n1094 DVSS.n1053 2.24964
R35711 DVSS.n1071 DVSS.n1053 2.24964
R35712 DVSS.n1097 DVSS.n1053 2.24964
R35713 DVSS.n1075 DVSS.n1053 2.24964
R35714 DVSS.n1099 DVSS.n1053 2.24964
R35715 DVSS.n1079 DVSS.n1053 2.24964
R35716 DVSS.n1137 DVSS.n1108 2.24964
R35717 DVSS.n1139 DVSS.n1108 2.24964
R35718 DVSS.n1164 DVSS.n1109 2.24964
R35719 DVSS.n1141 DVSS.n1108 2.24964
R35720 DVSS.n1164 DVSS.n1159 2.24964
R35721 DVSS.n1144 DVSS.n1108 2.24964
R35722 DVSS.n1164 DVSS.n1160 2.24964
R35723 DVSS.n1146 DVSS.n1108 2.24964
R35724 DVSS.n1164 DVSS.n1158 2.24964
R35725 DVSS.n1149 DVSS.n1108 2.24964
R35726 DVSS.n1164 DVSS.n1161 2.24964
R35727 DVSS.n1164 DVSS.n1157 2.24964
R35728 DVSS.n1164 DVSS.n1162 2.24964
R35729 DVSS.n1164 DVSS.n1156 2.24964
R35730 DVSS.n1164 DVSS.n1163 2.24964
R35731 DVSS.n1164 DVSS.n1155 2.24964
R35732 DVSS.n13007 DVSS.n12972 2.24964
R35733 DVSS.n13010 DVSS.n12972 2.24964
R35734 DVSS.n13009 DVSS.n12973 2.24964
R35735 DVSS.n13012 DVSS.n12972 2.24964
R35736 DVSS.n13021 DVSS.n12973 2.24964
R35737 DVSS.n13024 DVSS.n12972 2.24964
R35738 DVSS.n13023 DVSS.n12973 2.24964
R35739 DVSS.n13026 DVSS.n12972 2.24964
R35740 DVSS.n13035 DVSS.n12973 2.24964
R35741 DVSS.n13038 DVSS.n12972 2.24964
R35742 DVSS.n13037 DVSS.n12973 2.24964
R35743 DVSS.n12994 DVSS.n12973 2.24964
R35744 DVSS.n13048 DVSS.n12973 2.24964
R35745 DVSS.n12998 DVSS.n12973 2.24964
R35746 DVSS.n13057 DVSS.n12973 2.24964
R35747 DVSS.n13002 DVSS.n12973 2.24964
R35748 DVSS.n376 DVSS.n373 2.24964
R35749 DVSS.n376 DVSS.n372 2.24964
R35750 DVSS.n352 DVSS.n334 2.24964
R35751 DVSS.n376 DVSS.n374 2.24964
R35752 DVSS.n355 DVSS.n334 2.24964
R35753 DVSS.n376 DVSS.n371 2.24964
R35754 DVSS.n357 DVSS.n334 2.24964
R35755 DVSS.n376 DVSS.n375 2.24964
R35756 DVSS.n360 DVSS.n334 2.24964
R35757 DVSS.n376 DVSS.n370 2.24964
R35758 DVSS.n362 DVSS.n334 2.24964
R35759 DVSS.n339 DVSS.n334 2.24964
R35760 DVSS.n365 DVSS.n334 2.24964
R35761 DVSS.n343 DVSS.n334 2.24964
R35762 DVSS.n367 DVSS.n334 2.24964
R35763 DVSS.n347 DVSS.n334 2.24964
R35764 DVSS.n22472 DVSS.n22464 2.24964
R35765 DVSS.n22498 DVSS.n22496 2.24964
R35766 DVSS.n22472 DVSS.n22463 2.24964
R35767 DVSS.n22498 DVSS.n22497 2.24964
R35768 DVSS.n22472 DVSS.n22465 2.24964
R35769 DVSS.n22498 DVSS.n22495 2.24964
R35770 DVSS.n22472 DVSS.n22466 2.24964
R35771 DVSS.n22472 DVSS.n22467 2.24964
R35772 DVSS.n22498 DVSS.n22494 2.24964
R35773 DVSS.n22472 DVSS.n22468 2.24964
R35774 DVSS.n22472 DVSS.n22469 2.24964
R35775 DVSS.n22498 DVSS.n22493 2.24964
R35776 DVSS.n22472 DVSS.n22470 2.24964
R35777 DVSS.n22472 DVSS.n22471 2.24964
R35778 DVSS.n22498 DVSS.n22492 2.24964
R35779 DVSS.n22498 DVSS.n22491 2.24964
R35780 DVSS.n22498 DVSS.n22462 2.24964
R35781 DVSS.n239 DVSS.n231 2.24964
R35782 DVSS.n262 DVSS.n260 2.24964
R35783 DVSS.n239 DVSS.n230 2.24964
R35784 DVSS.n262 DVSS.n261 2.24964
R35785 DVSS.n239 DVSS.n232 2.24964
R35786 DVSS.n262 DVSS.n259 2.24964
R35787 DVSS.n239 DVSS.n233 2.24964
R35788 DVSS.n239 DVSS.n234 2.24964
R35789 DVSS.n262 DVSS.n258 2.24964
R35790 DVSS.n239 DVSS.n235 2.24964
R35791 DVSS.n239 DVSS.n236 2.24964
R35792 DVSS.n262 DVSS.n257 2.24964
R35793 DVSS.n239 DVSS.n237 2.24964
R35794 DVSS.n239 DVSS.n238 2.24964
R35795 DVSS.n262 DVSS.n256 2.24964
R35796 DVSS.n262 DVSS.n255 2.24964
R35797 DVSS.n262 DVSS.n229 2.24964
R35798 DVSS.n159 DVSS.n151 2.24964
R35799 DVSS.n182 DVSS.n180 2.24964
R35800 DVSS.n159 DVSS.n150 2.24964
R35801 DVSS.n182 DVSS.n181 2.24964
R35802 DVSS.n159 DVSS.n152 2.24964
R35803 DVSS.n182 DVSS.n179 2.24964
R35804 DVSS.n159 DVSS.n153 2.24964
R35805 DVSS.n159 DVSS.n154 2.24964
R35806 DVSS.n182 DVSS.n178 2.24964
R35807 DVSS.n159 DVSS.n155 2.24964
R35808 DVSS.n159 DVSS.n156 2.24964
R35809 DVSS.n182 DVSS.n177 2.24964
R35810 DVSS.n159 DVSS.n157 2.24964
R35811 DVSS.n159 DVSS.n158 2.24964
R35812 DVSS.n182 DVSS.n176 2.24964
R35813 DVSS.n182 DVSS.n175 2.24964
R35814 DVSS.n182 DVSS.n149 2.24964
R35815 DVSS.n94 DVSS.n86 2.24964
R35816 DVSS.n23172 DVSS.n23170 2.24964
R35817 DVSS.n94 DVSS.n85 2.24964
R35818 DVSS.n23172 DVSS.n23171 2.24964
R35819 DVSS.n94 DVSS.n87 2.24964
R35820 DVSS.n23172 DVSS.n23169 2.24964
R35821 DVSS.n94 DVSS.n88 2.24964
R35822 DVSS.n94 DVSS.n89 2.24964
R35823 DVSS.n23172 DVSS.n23168 2.24964
R35824 DVSS.n94 DVSS.n90 2.24964
R35825 DVSS.n94 DVSS.n91 2.24964
R35826 DVSS.n23172 DVSS.n23167 2.24964
R35827 DVSS.n94 DVSS.n92 2.24964
R35828 DVSS.n94 DVSS.n93 2.24964
R35829 DVSS.n23172 DVSS.n23166 2.24964
R35830 DVSS.n23172 DVSS.n23165 2.24964
R35831 DVSS.n23172 DVSS.n84 2.24964
R35832 DVSS.n21932 DVSS.n21923 2.24964
R35833 DVSS.n21881 DVSS.n21852 2.24964
R35834 DVSS.n21932 DVSS.n21924 2.24964
R35835 DVSS.n21890 DVSS.n21852 2.24964
R35836 DVSS.n21932 DVSS.n21925 2.24964
R35837 DVSS.n21932 DVSS.n21926 2.24964
R35838 DVSS.n21900 DVSS.n21852 2.24964
R35839 DVSS.n21932 DVSS.n21927 2.24964
R35840 DVSS.n21932 DVSS.n21928 2.24964
R35841 DVSS.n21910 DVSS.n21852 2.24964
R35842 DVSS.n21932 DVSS.n21929 2.24964
R35843 DVSS.n21932 DVSS.n21930 2.24964
R35844 DVSS.n21920 DVSS.n21852 2.24964
R35845 DVSS.n21932 DVSS.n21931 2.24964
R35846 DVSS.n21933 DVSS.n21932 2.24964
R35847 DVSS.n21942 DVSS.n21852 2.24964
R35848 DVSS.n21932 DVSS.n21851 2.24964
R35849 DVSS.n21615 DVSS.n21604 2.24964
R35850 DVSS.n21622 DVSS.n21621 2.24964
R35851 DVSS.n21615 DVSS.n21605 2.24964
R35852 DVSS.n21622 DVSS.n21620 2.24964
R35853 DVSS.n21615 DVSS.n21606 2.24964
R35854 DVSS.n21615 DVSS.n21607 2.24964
R35855 DVSS.n21622 DVSS.n21619 2.24964
R35856 DVSS.n21615 DVSS.n21608 2.24964
R35857 DVSS.n21615 DVSS.n21609 2.24964
R35858 DVSS.n21622 DVSS.n21618 2.24964
R35859 DVSS.n21615 DVSS.n21610 2.24964
R35860 DVSS.n21615 DVSS.n21611 2.24964
R35861 DVSS.n21622 DVSS.n21617 2.24964
R35862 DVSS.n21615 DVSS.n21612 2.24964
R35863 DVSS.n21615 DVSS.n21613 2.24964
R35864 DVSS.n21622 DVSS.n21616 2.24964
R35865 DVSS.n21615 DVSS.n21614 2.24964
R35866 DVSS.n21718 DVSS.n21707 2.24964
R35867 DVSS.n21725 DVSS.n21724 2.24964
R35868 DVSS.n21718 DVSS.n21708 2.24964
R35869 DVSS.n21725 DVSS.n21723 2.24964
R35870 DVSS.n21718 DVSS.n21709 2.24964
R35871 DVSS.n21718 DVSS.n21710 2.24964
R35872 DVSS.n21725 DVSS.n21722 2.24964
R35873 DVSS.n21718 DVSS.n21711 2.24964
R35874 DVSS.n21718 DVSS.n21712 2.24964
R35875 DVSS.n21725 DVSS.n21721 2.24964
R35876 DVSS.n21718 DVSS.n21713 2.24964
R35877 DVSS.n21718 DVSS.n21714 2.24964
R35878 DVSS.n21725 DVSS.n21720 2.24964
R35879 DVSS.n21718 DVSS.n21715 2.24964
R35880 DVSS.n21718 DVSS.n21716 2.24964
R35881 DVSS.n21725 DVSS.n21719 2.24964
R35882 DVSS.n21718 DVSS.n21717 2.24964
R35883 DVSS.n21811 DVSS.n21800 2.24964
R35884 DVSS.n21818 DVSS.n21817 2.24964
R35885 DVSS.n21811 DVSS.n21801 2.24964
R35886 DVSS.n21818 DVSS.n21816 2.24964
R35887 DVSS.n21811 DVSS.n21802 2.24964
R35888 DVSS.n21811 DVSS.n21803 2.24964
R35889 DVSS.n21818 DVSS.n21815 2.24964
R35890 DVSS.n21811 DVSS.n21804 2.24964
R35891 DVSS.n21811 DVSS.n21805 2.24964
R35892 DVSS.n21818 DVSS.n21814 2.24964
R35893 DVSS.n21811 DVSS.n21806 2.24964
R35894 DVSS.n21811 DVSS.n21807 2.24964
R35895 DVSS.n21818 DVSS.n21813 2.24964
R35896 DVSS.n21811 DVSS.n21808 2.24964
R35897 DVSS.n21811 DVSS.n21809 2.24964
R35898 DVSS.n21818 DVSS.n21812 2.24964
R35899 DVSS.n21811 DVSS.n21810 2.24964
R35900 DVSS.n13635 DVSS.n13630 2.24953
R35901 DVSS.n21205 DVSS.n21204 2.24953
R35902 DVSS.n13635 DVSS.n13631 2.24953
R35903 DVSS.n21205 DVSS.n21203 2.24953
R35904 DVSS.n13635 DVSS.n13632 2.24953
R35905 DVSS.n21205 DVSS.n21202 2.24953
R35906 DVSS.n13635 DVSS.n13633 2.24953
R35907 DVSS.n21205 DVSS.n21201 2.24953
R35908 DVSS.n13635 DVSS.n13634 2.24953
R35909 DVSS.n21205 DVSS.n13636 2.24953
R35910 DVSS.n21139 DVSS.n21138 2.24953
R35911 DVSS.n13758 DVSS.n13730 2.24953
R35912 DVSS.n21139 DVSS.n21137 2.24953
R35913 DVSS.n13760 DVSS.n13730 2.24953
R35914 DVSS.n21139 DVSS.n21136 2.24953
R35915 DVSS.n13762 DVSS.n13730 2.24953
R35916 DVSS.n21139 DVSS.n21135 2.24953
R35917 DVSS.n13764 DVSS.n13730 2.24953
R35918 DVSS.n21139 DVSS.n21134 2.24953
R35919 DVSS.n13766 DVSS.n13730 2.24953
R35920 DVSS.n21139 DVSS.n21133 2.24953
R35921 DVSS.n13768 DVSS.n13730 2.24953
R35922 DVSS.n21139 DVSS.n21132 2.24953
R35923 DVSS.n13770 DVSS.n13730 2.24953
R35924 DVSS.n21139 DVSS.n21131 2.24953
R35925 DVSS.n13772 DVSS.n13730 2.24953
R35926 DVSS.n21139 DVSS.n21130 2.24953
R35927 DVSS.n13774 DVSS.n13730 2.24953
R35928 DVSS.n21139 DVSS.n21129 2.24953
R35929 DVSS.n13776 DVSS.n13730 2.24953
R35930 DVSS.n21140 DVSS.n21139 2.24953
R35931 DVSS.n13778 DVSS.n13730 2.24953
R35932 DVSS.n21139 DVSS.n13729 2.24953
R35933 DVSS.n13722 DVSS.n13707 2.24953
R35934 DVSS.n13727 DVSS.n13726 2.24953
R35935 DVSS.n13707 DVSS.n13703 2.24953
R35936 DVSS.n13727 DVSS.n13725 2.24953
R35937 DVSS.n13707 DVSS.n13704 2.24953
R35938 DVSS.n13727 DVSS.n13724 2.24953
R35939 DVSS.n13707 DVSS.n13705 2.24953
R35940 DVSS.n13727 DVSS.n13723 2.24953
R35941 DVSS.n13707 DVSS.n13706 2.24953
R35942 DVSS.n13727 DVSS.n13708 2.24953
R35943 DVSS.n15170 DVSS.n15165 2.24953
R35944 DVSS.n15214 DVSS.n15213 2.24953
R35945 DVSS.n15170 DVSS.n15166 2.24953
R35946 DVSS.n15214 DVSS.n15212 2.24953
R35947 DVSS.n15170 DVSS.n15167 2.24953
R35948 DVSS.n15214 DVSS.n15211 2.24953
R35949 DVSS.n15170 DVSS.n15168 2.24953
R35950 DVSS.n15214 DVSS.n15210 2.24953
R35951 DVSS.n15170 DVSS.n15169 2.24953
R35952 DVSS.n15214 DVSS.n15171 2.24953
R35953 DVSS.n17696 DVSS.n17675 2.24953
R35954 DVSS.n17771 DVSS.n17709 2.24953
R35955 DVSS.n17699 DVSS.n17675 2.24953
R35956 DVSS.n17771 DVSS.n17708 2.24953
R35957 DVSS.n17701 DVSS.n17675 2.24953
R35958 DVSS.n17771 DVSS.n17707 2.24953
R35959 DVSS.n17703 DVSS.n17675 2.24953
R35960 DVSS.n17772 DVSS.n17771 2.24953
R35961 DVSS.n17705 DVSS.n17675 2.24953
R35962 DVSS.n17771 DVSS.n17676 2.24953
R35963 DVSS.n15957 DVSS.n15942 2.24953
R35964 DVSS.n17673 DVSS.n15962 2.24953
R35965 DVSS.n15942 DVSS.n15938 2.24953
R35966 DVSS.n17673 DVSS.n15961 2.24953
R35967 DVSS.n15942 DVSS.n15939 2.24953
R35968 DVSS.n17673 DVSS.n15960 2.24953
R35969 DVSS.n15942 DVSS.n15940 2.24953
R35970 DVSS.n17673 DVSS.n15959 2.24953
R35971 DVSS.n15942 DVSS.n15941 2.24953
R35972 DVSS.n17673 DVSS.n15943 2.24953
R35973 DVSS.n16346 DVSS.n16345 2.24953
R35974 DVSS.n16348 DVSS.n16347 2.24953
R35975 DVSS.n15891 DVSS.n15889 2.24953
R35976 DVSS.n15893 DVSS.n15892 2.24953
R35977 DVSS.n15891 DVSS.n15890 2.24953
R35978 DVSS.n18149 DVSS.n15550 2.24953
R35979 DVSS.n15571 DVSS.n15551 2.24953
R35980 DVSS.n15572 DVSS.n15550 2.24953
R35981 DVSS.n18115 DVSS.n15593 2.24953
R35982 DVSS.n18117 DVSS.n15594 2.24953
R35983 DVSS.n15512 DVSS.n15492 2.24953
R35984 DVSS.n18201 DVSS.n18198 2.24953
R35985 DVSS.n15516 DVSS.n15492 2.24953
R35986 DVSS.n18201 DVSS.n18199 2.24953
R35987 DVSS.n15518 DVSS.n15492 2.24953
R35988 DVSS.n18201 DVSS.n18200 2.24953
R35989 DVSS.n15520 DVSS.n15492 2.24953
R35990 DVSS.n18202 DVSS.n18201 2.24953
R35991 DVSS.n18203 DVSS.n15492 2.24953
R35992 DVSS.n18201 DVSS.n15491 2.24953
R35993 DVSS.n18218 DVSS.n18217 2.24953
R35994 DVSS.n18237 DVSS.n18233 2.24953
R35995 DVSS.n18218 DVSS.n18216 2.24953
R35996 DVSS.n18237 DVSS.n18234 2.24953
R35997 DVSS.n18218 DVSS.n18215 2.24953
R35998 DVSS.n18237 DVSS.n18235 2.24953
R35999 DVSS.n18218 DVSS.n18214 2.24953
R36000 DVSS.n18237 DVSS.n18236 2.24953
R36001 DVSS.n18218 DVSS.n18213 2.24953
R36002 DVSS.n18237 DVSS.n18212 2.24953
R36003 DVSS.n15092 DVSS.n15085 2.24953
R36004 DVSS.n15118 DVSS.n15114 2.24953
R36005 DVSS.n15094 DVSS.n15085 2.24953
R36006 DVSS.n15118 DVSS.n15115 2.24953
R36007 DVSS.n15096 DVSS.n15085 2.24953
R36008 DVSS.n15118 DVSS.n15116 2.24953
R36009 DVSS.n15098 DVSS.n15085 2.24953
R36010 DVSS.n15118 DVSS.n15117 2.24953
R36011 DVSS.n15100 DVSS.n15085 2.24953
R36012 DVSS.n15118 DVSS.n15102 2.24953
R36013 DVSS.n14337 DVSS.n14336 2.24953
R36014 DVSS.n20968 DVSS.n20964 2.24953
R36015 DVSS.n14337 DVSS.n14335 2.24953
R36016 DVSS.n20968 DVSS.n20965 2.24953
R36017 DVSS.n14337 DVSS.n14334 2.24953
R36018 DVSS.n20968 DVSS.n20966 2.24953
R36019 DVSS.n14337 DVSS.n14333 2.24953
R36020 DVSS.n20968 DVSS.n20967 2.24953
R36021 DVSS.n14337 DVSS.n14332 2.24953
R36022 DVSS.n20968 DVSS.n14331 2.24953
R36023 DVSS.n21054 DVSS.n14240 2.24953
R36024 DVSS.n21047 DVSS.n14295 2.24953
R36025 DVSS.n21054 DVSS.n14241 2.24953
R36026 DVSS.n21047 DVSS.n14294 2.24953
R36027 DVSS.n21054 DVSS.n14242 2.24953
R36028 DVSS.n21047 DVSS.n14293 2.24953
R36029 DVSS.n21054 DVSS.n14243 2.24953
R36030 DVSS.n21047 DVSS.n14292 2.24953
R36031 DVSS.n21054 DVSS.n14244 2.24953
R36032 DVSS.n21047 DVSS.n14291 2.24953
R36033 DVSS.n21054 DVSS.n14245 2.24953
R36034 DVSS.n21047 DVSS.n14290 2.24953
R36035 DVSS.n21054 DVSS.n14246 2.24953
R36036 DVSS.n21047 DVSS.n14289 2.24953
R36037 DVSS.n21054 DVSS.n14247 2.24953
R36038 DVSS.n21047 DVSS.n14288 2.24953
R36039 DVSS.n21054 DVSS.n14248 2.24953
R36040 DVSS.n21047 DVSS.n14287 2.24953
R36041 DVSS.n21054 DVSS.n14249 2.24953
R36042 DVSS.n21048 DVSS.n21047 2.24953
R36043 DVSS.n21054 DVSS.n14250 2.24953
R36044 DVSS.n21047 DVSS.n14252 2.24953
R36045 DVSS.n21054 DVSS.n21053 2.24953
R36046 DVSS.n13394 DVSS.n13393 2.24953
R36047 DVSS.n21422 DVSS.n21418 2.24953
R36048 DVSS.n13394 DVSS.n13392 2.24953
R36049 DVSS.n21422 DVSS.n21419 2.24953
R36050 DVSS.n13394 DVSS.n13391 2.24953
R36051 DVSS.n21422 DVSS.n21420 2.24953
R36052 DVSS.n13394 DVSS.n13390 2.24953
R36053 DVSS.n21422 DVSS.n21421 2.24953
R36054 DVSS.n13394 DVSS.n13389 2.24953
R36055 DVSS.n21422 DVSS.n13388 2.24953
R36056 DVSS.n21254 DVSS.n13572 2.24901
R36057 DVSS.n18473 DVSS.n18393 2.24901
R36058 DVSS.n13542 DVSS.n13522 2.24901
R36059 DVSS.n13548 DVSS.n13522 2.24901
R36060 DVSS.n14484 DVSS.n14465 2.24901
R36061 DVSS.n14489 DVSS.n14465 2.24901
R36062 DVSS.n20009 DVSS.n14880 2.24901
R36063 DVSS.n20009 DVSS.n14876 2.24901
R36064 DVSS.n15316 DVSS.n14903 2.24901
R36065 DVSS.n15321 DVSS.n14903 2.24901
R36066 DVSS.n17643 DVSS.n16079 2.24901
R36067 DVSS.n17643 DVSS.n16075 2.24901
R36068 DVSS.n16269 DVSS.n16096 2.24901
R36069 DVSS.n16274 DVSS.n16096 2.24901
R36070 DVSS.n13490 DVSS.n13472 2.24901
R36071 DVSS.n13496 DVSS.n13472 2.24901
R36072 DVSS.n14434 DVSS.n14416 2.24901
R36073 DVSS.n14440 DVSS.n14416 2.24901
R36074 DVSS.n14951 DVSS.n14864 2.24901
R36075 DVSS.n14987 DVSS.n14864 2.24901
R36076 DVSS.n15388 DVSS.n14938 2.24901
R36077 DVSS.n15393 DVSS.n14938 2.24901
R36078 DVSS.n16844 DVSS.n16148 2.24901
R36079 DVSS.n16849 DVSS.n16148 2.24901
R36080 DVSS.n16825 DVSS.n16157 2.24901
R36081 DVSS.n16825 DVSS.n16153 2.24901
R36082 DVSS.n13596 DVSS.n13571 2.24901
R36083 DVSS.n20714 DVSS.n14512 2.24901
R36084 DVSS.n20802 DVSS.n14512 2.24901
R36085 DVSS.n18388 DVSS.n14536 2.24901
R36086 DVSS.n18381 DVSS.n15243 2.24901
R36087 DVSS.n15268 DVSS.n15265 2.24901
R36088 DVSS.n16023 DVSS.n16000 2.24901
R36089 DVSS.n16028 DVSS.n16002 2.24901
R36090 DVSS.n16316 DVSS.n16299 2.24901
R36091 DVSS.n16636 DVSS.n16300 2.24901
R36092 DVSS.n13643 DVSS.n13624 2.24901
R36093 DVSS.n13648 DVSS.n13624 2.24901
R36094 DVSS.n21144 DVSS.n13697 2.24901
R36095 DVSS.n21144 DVSS.n13728 2.24901
R36096 DVSS.n15159 DVSS.n13702 2.24901
R36097 DVSS.n15181 DVSS.n13702 2.24901
R36098 DVSS.n17683 DVSS.n15164 2.24901
R36099 DVSS.n17688 DVSS.n15164 2.24901
R36100 DVSS.n17776 DVSS.n15932 2.24901
R36101 DVSS.n17776 DVSS.n17674 2.24901
R36102 DVSS.n16552 DVSS.n15937 2.24901
R36103 DVSS.n16557 DVSS.n15937 2.24901
R36104 DVSS.n13443 DVSS.n13420 2.24901
R36105 DVSS.n13448 DVSS.n13420 2.24901
R36106 DVSS.n14384 DVSS.n14367 2.24901
R36107 DVSS.n14389 DVSS.n14367 2.24901
R36108 DVSS.n15024 DVSS.n14853 2.24901
R36109 DVSS.n15029 DVSS.n14853 2.24901
R36110 DVSS.n15466 DVSS.n15011 2.24901
R36111 DVSS.n15461 DVSS.n15011 2.24901
R36112 DVSS.n17546 DVSS.n16895 2.24901
R36113 DVSS.n17541 DVSS.n16895 2.24901
R36114 DVSS.n15677 DVSS.n15676 2.24901
R36115 DVSS.n15677 DVSS.n15675 2.24901
R36116 DVSS.n15602 DVSS.n15589 2.24901
R36117 DVSS.n15606 DVSS.n15589 2.24901
R36118 DVSS.n15515 DVSS.n15514 2.24901
R36119 DVSS.n15515 DVSS.n15513 2.24901
R36120 DVSS.n18225 DVSS.n18207 2.24901
R36121 DVSS.n18230 DVSS.n18207 2.24901
R36122 DVSS.n15109 DVSS.n15093 2.24901
R36123 DVSS.n19951 DVSS.n15093 2.24901
R36124 DVSS.n14343 DVSS.n14326 2.24901
R36125 DVSS.n14348 DVSS.n14326 2.24901
R36126 DVSS.n13401 DVSS.n13383 2.24901
R36127 DVSS.n13406 DVSS.n13383 2.24901
R36128 DVSS.n22876 DVSS.n464 2.24901
R36129 DVSS.n479 DVSS.n464 2.24901
R36130 DVSS.n727 DVSS.n707 2.24901
R36131 DVSS.n722 DVSS.n707 2.24901
R36132 DVSS.n683 DVSS.n655 2.24901
R36133 DVSS.n22712 DVSS.n666 2.24901
R36134 DVSS.n625 DVSS.n602 2.24901
R36135 DVSS.n630 DVSS.n602 2.24901
R36136 DVSS.n575 DVSS.n554 2.24901
R36137 DVSS.n580 DVSS.n554 2.24901
R36138 DVSS.n524 DVSS.n502 2.24901
R36139 DVSS.n529 DVSS.n502 2.24901
R36140 DVSS.n15814 DVSS.n15790 2.24882
R36141 DVSS.n15819 DVSS.n15790 2.24882
R36142 DVSS.n15764 DVSS.n15743 2.24882
R36143 DVSS.n15769 DVSS.n15743 2.24882
R36144 DVSS.n15860 DVSS.n15841 2.24882
R36145 DVSS.n17862 DVSS.n15841 2.24882
R36146 DVSS.n15901 DVSS.n15883 2.24882
R36147 DVSS.n15906 DVSS.n15883 2.24882
R36148 DVSS.n18047 DVSS.n15696 2.24882
R36149 DVSS.n18047 DVSS.n15692 2.24882
R36150 DVSS.n15569 DVSS.n15568 2.24882
R36151 DVSS.n15569 DVSS.n15567 2.24882
R36152 DVSS.n12768 DVSS.n12410 2.24752
R36153 DVSS.n6404 DVSS.n6259 2.24752
R36154 DVSS.n12742 DVSS.n12553 2.24752
R36155 DVSS.n12506 DVSS.n12459 2.24752
R36156 DVSS.n12553 DVSS.n12552 2.24752
R36157 DVSS.n12506 DVSS.n12460 2.24752
R36158 DVSS.n12553 DVSS.n12551 2.24752
R36159 DVSS.n12506 DVSS.n12461 2.24752
R36160 DVSS.n12553 DVSS.n12550 2.24752
R36161 DVSS.n12506 DVSS.n12462 2.24752
R36162 DVSS.n12553 DVSS.n12549 2.24752
R36163 DVSS.n12506 DVSS.n12463 2.24752
R36164 DVSS.n12553 DVSS.n12548 2.24752
R36165 DVSS.n12506 DVSS.n12464 2.24752
R36166 DVSS.n12553 DVSS.n12547 2.24752
R36167 DVSS.n12506 DVSS.n12465 2.24752
R36168 DVSS.n12553 DVSS.n12546 2.24752
R36169 DVSS.n12506 DVSS.n12466 2.24752
R36170 DVSS.n12553 DVSS.n12545 2.24752
R36171 DVSS.n12506 DVSS.n12467 2.24752
R36172 DVSS.n12553 DVSS.n12544 2.24752
R36173 DVSS.n12506 DVSS.n12468 2.24752
R36174 DVSS.n12553 DVSS.n12543 2.24752
R36175 DVSS.n12506 DVSS.n12469 2.24752
R36176 DVSS.n12553 DVSS.n12542 2.24752
R36177 DVSS.n12506 DVSS.n12470 2.24752
R36178 DVSS.n12553 DVSS.n12541 2.24752
R36179 DVSS.n12506 DVSS.n12471 2.24752
R36180 DVSS.n12553 DVSS.n12540 2.24752
R36181 DVSS.n12506 DVSS.n12472 2.24752
R36182 DVSS.n12553 DVSS.n12539 2.24752
R36183 DVSS.n12506 DVSS.n12473 2.24752
R36184 DVSS.n12553 DVSS.n12538 2.24752
R36185 DVSS.n12506 DVSS.n12474 2.24752
R36186 DVSS.n12553 DVSS.n12537 2.24752
R36187 DVSS.n12506 DVSS.n12475 2.24752
R36188 DVSS.n12553 DVSS.n12536 2.24752
R36189 DVSS.n12506 DVSS.n12476 2.24752
R36190 DVSS.n12553 DVSS.n12535 2.24752
R36191 DVSS.n12506 DVSS.n12477 2.24752
R36192 DVSS.n12553 DVSS.n12534 2.24752
R36193 DVSS.n12506 DVSS.n12478 2.24752
R36194 DVSS.n12553 DVSS.n12533 2.24752
R36195 DVSS.n12506 DVSS.n12479 2.24752
R36196 DVSS.n12553 DVSS.n12532 2.24752
R36197 DVSS.n12506 DVSS.n12480 2.24752
R36198 DVSS.n12553 DVSS.n12531 2.24752
R36199 DVSS.n12506 DVSS.n12481 2.24752
R36200 DVSS.n12553 DVSS.n12530 2.24752
R36201 DVSS.n12506 DVSS.n12482 2.24752
R36202 DVSS.n12553 DVSS.n12529 2.24752
R36203 DVSS.n12506 DVSS.n12483 2.24752
R36204 DVSS.n12553 DVSS.n12528 2.24752
R36205 DVSS.n12506 DVSS.n12484 2.24752
R36206 DVSS.n12553 DVSS.n12527 2.24752
R36207 DVSS.n12506 DVSS.n12485 2.24752
R36208 DVSS.n12553 DVSS.n12526 2.24752
R36209 DVSS.n12506 DVSS.n12486 2.24752
R36210 DVSS.n12553 DVSS.n12525 2.24752
R36211 DVSS.n12506 DVSS.n12487 2.24752
R36212 DVSS.n12553 DVSS.n12524 2.24752
R36213 DVSS.n12506 DVSS.n12488 2.24752
R36214 DVSS.n12553 DVSS.n12523 2.24752
R36215 DVSS.n12506 DVSS.n12489 2.24752
R36216 DVSS.n12553 DVSS.n12522 2.24752
R36217 DVSS.n12506 DVSS.n12490 2.24752
R36218 DVSS.n12553 DVSS.n12521 2.24752
R36219 DVSS.n12506 DVSS.n12491 2.24752
R36220 DVSS.n12553 DVSS.n12520 2.24752
R36221 DVSS.n12506 DVSS.n12492 2.24752
R36222 DVSS.n12553 DVSS.n12519 2.24752
R36223 DVSS.n12506 DVSS.n12493 2.24752
R36224 DVSS.n12553 DVSS.n12518 2.24752
R36225 DVSS.n12506 DVSS.n12494 2.24752
R36226 DVSS.n12553 DVSS.n12517 2.24752
R36227 DVSS.n12506 DVSS.n12495 2.24752
R36228 DVSS.n12553 DVSS.n12516 2.24752
R36229 DVSS.n12506 DVSS.n12496 2.24752
R36230 DVSS.n12553 DVSS.n12515 2.24752
R36231 DVSS.n12506 DVSS.n12497 2.24752
R36232 DVSS.n12553 DVSS.n12514 2.24752
R36233 DVSS.n12506 DVSS.n12498 2.24752
R36234 DVSS.n12553 DVSS.n12513 2.24752
R36235 DVSS.n12506 DVSS.n12499 2.24752
R36236 DVSS.n12553 DVSS.n12512 2.24752
R36237 DVSS.n12506 DVSS.n12500 2.24752
R36238 DVSS.n12553 DVSS.n12511 2.24752
R36239 DVSS.n12506 DVSS.n12501 2.24752
R36240 DVSS.n12553 DVSS.n12510 2.24752
R36241 DVSS.n12506 DVSS.n12502 2.24752
R36242 DVSS.n12553 DVSS.n12509 2.24752
R36243 DVSS.n12506 DVSS.n12503 2.24752
R36244 DVSS.n12553 DVSS.n12508 2.24752
R36245 DVSS.n12506 DVSS.n12504 2.24752
R36246 DVSS.n12553 DVSS.n12507 2.24752
R36247 DVSS.n12506 DVSS.n12505 2.24752
R36248 DVSS.n12553 DVSS.n12358 2.24752
R36249 DVSS.n12506 DVSS.n12357 2.24752
R36250 DVSS.n6658 DVSS.n6657 2.24752
R36251 DVSS.n12754 DVSS.n12753 2.24752
R36252 DVSS.n6657 DVSS.n6255 2.24752
R36253 DVSS.n12755 DVSS.n12754 2.24752
R36254 DVSS.n6652 DVSS.n6650 2.24752
R36255 DVSS.n6310 DVSS.n6259 2.24752
R36256 DVSS.n6652 DVSS.n6649 2.24752
R36257 DVSS.n6312 DVSS.n6259 2.24752
R36258 DVSS.n6652 DVSS.n6648 2.24752
R36259 DVSS.n6314 DVSS.n6259 2.24752
R36260 DVSS.n6652 DVSS.n6647 2.24752
R36261 DVSS.n6316 DVSS.n6259 2.24752
R36262 DVSS.n6652 DVSS.n6646 2.24752
R36263 DVSS.n6318 DVSS.n6259 2.24752
R36264 DVSS.n6652 DVSS.n6645 2.24752
R36265 DVSS.n6320 DVSS.n6259 2.24752
R36266 DVSS.n6652 DVSS.n6644 2.24752
R36267 DVSS.n6322 DVSS.n6259 2.24752
R36268 DVSS.n6652 DVSS.n6643 2.24752
R36269 DVSS.n6324 DVSS.n6259 2.24752
R36270 DVSS.n6652 DVSS.n6642 2.24752
R36271 DVSS.n6326 DVSS.n6259 2.24752
R36272 DVSS.n6652 DVSS.n6641 2.24752
R36273 DVSS.n6328 DVSS.n6259 2.24752
R36274 DVSS.n6652 DVSS.n6640 2.24752
R36275 DVSS.n6330 DVSS.n6259 2.24752
R36276 DVSS.n6652 DVSS.n6639 2.24752
R36277 DVSS.n6332 DVSS.n6259 2.24752
R36278 DVSS.n6652 DVSS.n6638 2.24752
R36279 DVSS.n6334 DVSS.n6259 2.24752
R36280 DVSS.n6652 DVSS.n6637 2.24752
R36281 DVSS.n6336 DVSS.n6259 2.24752
R36282 DVSS.n6652 DVSS.n6636 2.24752
R36283 DVSS.n6338 DVSS.n6259 2.24752
R36284 DVSS.n6652 DVSS.n6635 2.24752
R36285 DVSS.n6340 DVSS.n6259 2.24752
R36286 DVSS.n6652 DVSS.n6634 2.24752
R36287 DVSS.n6342 DVSS.n6259 2.24752
R36288 DVSS.n6652 DVSS.n6633 2.24752
R36289 DVSS.n6344 DVSS.n6259 2.24752
R36290 DVSS.n6652 DVSS.n6632 2.24752
R36291 DVSS.n6346 DVSS.n6259 2.24752
R36292 DVSS.n6652 DVSS.n6631 2.24752
R36293 DVSS.n6348 DVSS.n6259 2.24752
R36294 DVSS.n6652 DVSS.n6630 2.24752
R36295 DVSS.n6350 DVSS.n6259 2.24752
R36296 DVSS.n6652 DVSS.n6629 2.24752
R36297 DVSS.n6352 DVSS.n6259 2.24752
R36298 DVSS.n6652 DVSS.n6628 2.24752
R36299 DVSS.n6354 DVSS.n6259 2.24752
R36300 DVSS.n6652 DVSS.n6627 2.24752
R36301 DVSS.n6356 DVSS.n6259 2.24752
R36302 DVSS.n6652 DVSS.n6626 2.24752
R36303 DVSS.n6358 DVSS.n6259 2.24752
R36304 DVSS.n6652 DVSS.n6625 2.24752
R36305 DVSS.n6360 DVSS.n6259 2.24752
R36306 DVSS.n6652 DVSS.n6624 2.24752
R36307 DVSS.n6362 DVSS.n6259 2.24752
R36308 DVSS.n6652 DVSS.n6623 2.24752
R36309 DVSS.n6364 DVSS.n6259 2.24752
R36310 DVSS.n6652 DVSS.n6622 2.24752
R36311 DVSS.n6366 DVSS.n6259 2.24752
R36312 DVSS.n6652 DVSS.n6621 2.24752
R36313 DVSS.n6368 DVSS.n6259 2.24752
R36314 DVSS.n6652 DVSS.n6620 2.24752
R36315 DVSS.n6370 DVSS.n6259 2.24752
R36316 DVSS.n6652 DVSS.n6619 2.24752
R36317 DVSS.n6372 DVSS.n6259 2.24752
R36318 DVSS.n6652 DVSS.n6618 2.24752
R36319 DVSS.n6374 DVSS.n6259 2.24752
R36320 DVSS.n6652 DVSS.n6617 2.24752
R36321 DVSS.n6376 DVSS.n6259 2.24752
R36322 DVSS.n6652 DVSS.n6616 2.24752
R36323 DVSS.n6378 DVSS.n6259 2.24752
R36324 DVSS.n6652 DVSS.n6615 2.24752
R36325 DVSS.n6380 DVSS.n6259 2.24752
R36326 DVSS.n6652 DVSS.n6614 2.24752
R36327 DVSS.n6382 DVSS.n6259 2.24752
R36328 DVSS.n6652 DVSS.n6613 2.24752
R36329 DVSS.n6384 DVSS.n6259 2.24752
R36330 DVSS.n6652 DVSS.n6612 2.24752
R36331 DVSS.n6386 DVSS.n6259 2.24752
R36332 DVSS.n6652 DVSS.n6611 2.24752
R36333 DVSS.n6388 DVSS.n6259 2.24752
R36334 DVSS.n6652 DVSS.n6610 2.24752
R36335 DVSS.n6390 DVSS.n6259 2.24752
R36336 DVSS.n6652 DVSS.n6609 2.24752
R36337 DVSS.n6392 DVSS.n6259 2.24752
R36338 DVSS.n6652 DVSS.n6608 2.24752
R36339 DVSS.n6394 DVSS.n6259 2.24752
R36340 DVSS.n6652 DVSS.n6607 2.24752
R36341 DVSS.n6396 DVSS.n6259 2.24752
R36342 DVSS.n6652 DVSS.n6606 2.24752
R36343 DVSS.n6398 DVSS.n6259 2.24752
R36344 DVSS.n6652 DVSS.n6605 2.24752
R36345 DVSS.n6400 DVSS.n6259 2.24752
R36346 DVSS.n6652 DVSS.n6604 2.24752
R36347 DVSS.n6402 DVSS.n6259 2.24752
R36348 DVSS.n6652 DVSS.n6603 2.24752
R36349 DVSS.n6652 DVSS.n6651 2.24752
R36350 DVSS.n12347 DVSS.n12346 2.24752
R36351 DVSS.n6254 DVSS.n6253 2.24752
R36352 DVSS.n12350 DVSS.n12346 2.24752
R36353 DVSS.n6253 DVSS.n6245 2.24752
R36354 DVSS.n12774 DVSS.n12345 2.24681
R36355 DVSS.n6249 DVSS.n6244 2.24681
R36356 DVSS.n6663 DVSS.n6242 2.24681
R36357 DVSS.n17366 DVSS.n17333 2.24456
R36358 DVSS.n17367 DVSS.n17366 2.24456
R36359 DVSS.n17366 DVSS.n17365 2.24456
R36360 DVSS.n17366 DVSS.n17364 2.24456
R36361 DVSS.n17366 DVSS.n17363 2.24456
R36362 DVSS.n17366 DVSS.n17362 2.24456
R36363 DVSS.n17366 DVSS.n17361 2.24456
R36364 DVSS.n17366 DVSS.n17360 2.24456
R36365 DVSS.n17357 DVSS.n17332 2.24456
R36366 DVSS.n17355 DVSS.n17332 2.24456
R36367 DVSS.n17353 DVSS.n17332 2.24456
R36368 DVSS.n17351 DVSS.n17332 2.24456
R36369 DVSS.n17349 DVSS.n17332 2.24456
R36370 DVSS.n17347 DVSS.n17332 2.24456
R36371 DVSS.n17345 DVSS.n17332 2.24456
R36372 DVSS.n17343 DVSS.n17332 2.24456
R36373 DVSS.n17408 DVSS.n17268 2.24456
R36374 DVSS.n17408 DVSS.n17267 2.24456
R36375 DVSS.n17408 DVSS.n17266 2.24456
R36376 DVSS.n17408 DVSS.n17265 2.24456
R36377 DVSS.n17408 DVSS.n17264 2.24456
R36378 DVSS.n17408 DVSS.n17263 2.24456
R36379 DVSS.n17408 DVSS.n17262 2.24456
R36380 DVSS.n17291 DVSS.n17259 2.24456
R36381 DVSS.n17289 DVSS.n17259 2.24456
R36382 DVSS.n17287 DVSS.n17259 2.24456
R36383 DVSS.n17285 DVSS.n17259 2.24456
R36384 DVSS.n17283 DVSS.n17259 2.24456
R36385 DVSS.n17281 DVSS.n17259 2.24456
R36386 DVSS.n17270 DVSS.n17259 2.24456
R36387 DVSS.n17476 DVSS.n17475 2.24456
R36388 DVSS.n17475 DVSS.n17164 2.24456
R36389 DVSS.n17475 DVSS.n17158 2.24456
R36390 DVSS.n17475 DVSS.n17154 2.24456
R36391 DVSS.n17475 DVSS.n17150 2.24456
R36392 DVSS.n17475 DVSS.n17146 2.24456
R36393 DVSS.n17475 DVSS.n17142 2.24456
R36394 DVSS.n17172 DVSS.n17138 2.24456
R36395 DVSS.n17166 DVSS.n17138 2.24456
R36396 DVSS.n17144 DVSS.n17138 2.24456
R36397 DVSS.n17148 DVSS.n17138 2.24456
R36398 DVSS.n17152 DVSS.n17138 2.24456
R36399 DVSS.n17156 DVSS.n17138 2.24456
R36400 DVSS.n17160 DVSS.n17138 2.24456
R36401 DVSS.n17162 DVSS.n17138 2.24456
R36402 DVSS.n17492 DVSS.n16949 2.24456
R36403 DVSS.n17492 DVSS.n16948 2.24456
R36404 DVSS.n17492 DVSS.n16947 2.24456
R36405 DVSS.n17492 DVSS.n16946 2.24456
R36406 DVSS.n17492 DVSS.n16945 2.24456
R36407 DVSS.n17492 DVSS.n16944 2.24456
R36408 DVSS.n17492 DVSS.n16943 2.24456
R36409 DVSS.n17492 DVSS.n16942 2.24456
R36410 DVSS.n16972 DVSS.n16940 2.24456
R36411 DVSS.n16970 DVSS.n16940 2.24456
R36412 DVSS.n16968 DVSS.n16940 2.24456
R36413 DVSS.n16966 DVSS.n16940 2.24456
R36414 DVSS.n16964 DVSS.n16940 2.24456
R36415 DVSS.n16962 DVSS.n16940 2.24456
R36416 DVSS.n16960 DVSS.n16940 2.24456
R36417 DVSS.n16950 DVSS.n16940 2.24456
R36418 DVSS.n17416 DVSS.n17233 2.24456
R36419 DVSS.n17416 DVSS.n17232 2.24456
R36420 DVSS.n17416 DVSS.n17231 2.24456
R36421 DVSS.n17416 DVSS.n17230 2.24456
R36422 DVSS.n17416 DVSS.n17229 2.24456
R36423 DVSS.n17416 DVSS.n17228 2.24456
R36424 DVSS.n17416 DVSS.n17227 2.24456
R36425 DVSS.n17256 DVSS.n17224 2.24456
R36426 DVSS.n17254 DVSS.n17224 2.24456
R36427 DVSS.n17252 DVSS.n17224 2.24456
R36428 DVSS.n17250 DVSS.n17224 2.24456
R36429 DVSS.n17248 DVSS.n17224 2.24456
R36430 DVSS.n17246 DVSS.n17224 2.24456
R36431 DVSS.n17235 DVSS.n17224 2.24456
R36432 DVSS.n17468 DVSS.n17174 2.24456
R36433 DVSS.n17468 DVSS.n17465 2.24456
R36434 DVSS.n17468 DVSS.n17464 2.24456
R36435 DVSS.n17468 DVSS.n17463 2.24456
R36436 DVSS.n17468 DVSS.n17462 2.24456
R36437 DVSS.n17468 DVSS.n17461 2.24456
R36438 DVSS.n17468 DVSS.n17460 2.24456
R36439 DVSS.n17198 DVSS.n17173 2.24456
R36440 DVSS.n17466 DVSS.n17173 2.24456
R36441 DVSS.n17193 DVSS.n17173 2.24456
R36442 DVSS.n17191 DVSS.n17173 2.24456
R36443 DVSS.n17189 DVSS.n17173 2.24456
R36444 DVSS.n17187 DVSS.n17173 2.24456
R36445 DVSS.n17185 DVSS.n17173 2.24456
R36446 DVSS.n17183 DVSS.n17173 2.24456
R36447 DVSS.n17376 DVSS.n17312 2.24456
R36448 DVSS.n17374 DVSS.n17312 2.24456
R36449 DVSS.n17324 DVSS.n17312 2.24456
R36450 DVSS.n17322 DVSS.n17312 2.24456
R36451 DVSS.n17320 DVSS.n17312 2.24456
R36452 DVSS.n17372 DVSS.n17311 2.24456
R36453 DVSS.n17373 DVSS.n17372 2.24456
R36454 DVSS.n17372 DVSS.n17331 2.24456
R36455 DVSS.n17372 DVSS.n17330 2.24456
R36456 DVSS.n17372 DVSS.n17329 2.24456
R36457 DVSS.n17372 DVSS.n17328 2.24456
R36458 DVSS.n17403 DVSS.n17308 2.24456
R36459 DVSS.n17403 DVSS.n17307 2.24456
R36460 DVSS.n17403 DVSS.n17306 2.24456
R36461 DVSS.n17403 DVSS.n17305 2.24456
R36462 DVSS.n17399 DVSS.n17302 2.24456
R36463 DVSS.n17397 DVSS.n17302 2.24456
R36464 DVSS.n17395 DVSS.n17302 2.24456
R36465 DVSS.n17385 DVSS.n17302 2.24456
R36466 DVSS.n17301 DVSS.n17120 2.24456
R36467 DVSS.n17126 DVSS.n17119 2.24456
R36468 DVSS.n17128 DVSS.n17119 2.24456
R36469 DVSS.n17130 DVSS.n17119 2.24456
R36470 DVSS.n17132 DVSS.n17119 2.24456
R36471 DVSS.n17301 DVSS.n17137 2.24456
R36472 DVSS.n17301 DVSS.n17300 2.24456
R36473 DVSS.n17301 DVSS.n17298 2.24456
R36474 DVSS.n17301 DVSS.n17297 2.24456
R36475 DVSS.n17301 DVSS.n17296 2.24456
R36476 DVSS.n17518 DVSS.n16936 2.24456
R36477 DVSS.n17515 DVSS.n16936 2.24456
R36478 DVSS.n17512 DVSS.n16936 2.24456
R36479 DVSS.n17509 DVSS.n16936 2.24456
R36480 DVSS.n17506 DVSS.n16936 2.24456
R36481 DVSS.n17517 DVSS.n16938 2.24456
R36482 DVSS.n17514 DVSS.n16938 2.24456
R36483 DVSS.n17511 DVSS.n16938 2.24456
R36484 DVSS.n17508 DVSS.n16938 2.24456
R36485 DVSS.n17505 DVSS.n16938 2.24456
R36486 DVSS.n17501 DVSS.n16938 2.24456
R36487 DVSS.n17423 DVSS.n17222 2.24456
R36488 DVSS.n17423 DVSS.n17219 2.24456
R36489 DVSS.n17423 DVSS.n17216 2.24456
R36490 DVSS.n17423 DVSS.n17213 2.24456
R36491 DVSS.n17425 DVSS.n17205 2.24456
R36492 DVSS.n17425 DVSS.n17204 2.24456
R36493 DVSS.n17425 DVSS.n17203 2.24456
R36494 DVSS.n17425 DVSS.n17202 2.24456
R36495 DVSS.n17425 DVSS.n17201 2.24456
R36496 DVSS.n17425 DVSS.n17200 2.24456
R36497 DVSS.n17452 DVSS.n17427 2.24456
R36498 DVSS.n17452 DVSS.n17449 2.24456
R36499 DVSS.n17452 DVSS.n17448 2.24456
R36500 DVSS.n17452 DVSS.n17447 2.24456
R36501 DVSS.n17452 DVSS.n17446 2.24456
R36502 DVSS.n17450 DVSS.n17426 2.24456
R36503 DVSS.n17441 DVSS.n17426 2.24456
R36504 DVSS.n17439 DVSS.n17426 2.24456
R36505 DVSS.n17437 DVSS.n17426 2.24456
R36506 DVSS.n17435 DVSS.n17426 2.24456
R36507 DVSS.n17406 DVSS.n17258 2.24456
R36508 DVSS.n17406 DVSS.n17280 2.24456
R36509 DVSS.n17369 DVSS.n17342 2.24456
R36510 DVSS.n17168 DVSS.n16081 2.24456
R36511 DVSS.n17414 DVSS.n17223 2.24456
R36512 DVSS.n17414 DVSS.n17245 2.24456
R36513 DVSS.n17490 DVSS.n16939 2.24456
R36514 DVSS.n17470 DVSS.n17195 2.24456
R36515 DVSS.n17401 DVSS.n17392 2.24456
R36516 DVSS.n17401 DVSS.n17293 2.24456
R36517 DVSS.n17401 DVSS.n17394 2.24456
R36518 DVSS.n17378 DVSS.n17318 2.24456
R36519 DVSS.n17479 DVSS.n17134 2.24456
R36520 DVSS.n17520 DVSS.n17500 2.24456
R36521 DVSS.n17503 DVSS.n16936 2.24456
R36522 DVSS.n17209 DVSS.n17208 2.24456
R36523 DVSS.n17423 DVSS.n17422 2.24456
R36524 DVSS.n17454 DVSS.n17426 2.24456
R36525 DVSS.n17456 DVSS.n17443 2.24456
R36526 DVSS.n19308 DVSS.n19307 2.24442
R36527 DVSS.n19899 DVSS.n19039 2.24442
R36528 DVSS.n19899 DVSS.n19038 2.24442
R36529 DVSS.n19899 DVSS.n19037 2.24442
R36530 DVSS.n19899 DVSS.n19036 2.24442
R36531 DVSS.n19899 DVSS.n19035 2.24442
R36532 DVSS.n19899 DVSS.n19034 2.24442
R36533 DVSS.n19899 DVSS.n19033 2.24442
R36534 DVSS.n19899 DVSS.n19032 2.24442
R36535 DVSS.n19223 DVSS.n19041 2.24442
R36536 DVSS.n19226 DVSS.n19041 2.24442
R36537 DVSS.n19229 DVSS.n19041 2.24442
R36538 DVSS.n19232 DVSS.n19041 2.24442
R36539 DVSS.n19235 DVSS.n19041 2.24442
R36540 DVSS.n19238 DVSS.n19041 2.24442
R36541 DVSS.n19241 DVSS.n19041 2.24442
R36542 DVSS.n19245 DVSS.n19041 2.24442
R36543 DVSS.n19597 DVSS.n19159 2.24442
R36544 DVSS.n19600 DVSS.n19159 2.24442
R36545 DVSS.n19603 DVSS.n19159 2.24442
R36546 DVSS.n19606 DVSS.n19159 2.24442
R36547 DVSS.n19609 DVSS.n19159 2.24442
R36548 DVSS.n19612 DVSS.n19159 2.24442
R36549 DVSS.n19615 DVSS.n19159 2.24442
R36550 DVSS.n19619 DVSS.n19159 2.24442
R36551 DVSS.n19029 DVSS.n19028 2.24442
R36552 DVSS.n19029 DVSS.n19027 2.24442
R36553 DVSS.n19029 DVSS.n19026 2.24442
R36554 DVSS.n19029 DVSS.n19025 2.24442
R36555 DVSS.n19029 DVSS.n19024 2.24442
R36556 DVSS.n19029 DVSS.n19023 2.24442
R36557 DVSS.n19029 DVSS.n19022 2.24442
R36558 DVSS.n19225 DVSS.n19171 2.24442
R36559 DVSS.n19228 DVSS.n19171 2.24442
R36560 DVSS.n19231 DVSS.n19171 2.24442
R36561 DVSS.n19234 DVSS.n19171 2.24442
R36562 DVSS.n19237 DVSS.n19171 2.24442
R36563 DVSS.n19240 DVSS.n19171 2.24442
R36564 DVSS.n19243 DVSS.n19171 2.24442
R36565 DVSS.n19599 DVSS.n19157 2.24442
R36566 DVSS.n19602 DVSS.n19157 2.24442
R36567 DVSS.n19605 DVSS.n19157 2.24442
R36568 DVSS.n19608 DVSS.n19157 2.24442
R36569 DVSS.n19611 DVSS.n19157 2.24442
R36570 DVSS.n19614 DVSS.n19157 2.24442
R36571 DVSS.n19617 DVSS.n19157 2.24442
R36572 DVSS.n19901 DVSS.n19020 2.24442
R36573 DVSS.n19249 DVSS.n19248 2.24442
R36574 DVSS.n19623 DVSS.n19622 2.24442
R36575 DVSS.n22433 DVSS.n1013 2.24442
R36576 DVSS.n1014 DVSS.n1012 2.24442
R36577 DVSS.n22383 DVSS.n1016 2.24442
R36578 DVSS.n22383 DVSS.n1051 2.24442
R36579 DVSS.n22383 DVSS.n1050 2.24442
R36580 DVSS.n22383 DVSS.n1049 2.24442
R36581 DVSS.n22383 DVSS.n1048 2.24442
R36582 DVSS.n22383 DVSS.n1047 2.24442
R36583 DVSS.n22383 DVSS.n1046 2.24442
R36584 DVSS.n22383 DVSS.n1045 2.24442
R36585 DVSS.n22369 DVSS.n22366 2.24442
R36586 DVSS.n22369 DVSS.n22364 2.24442
R36587 DVSS.n22369 DVSS.n22361 2.24442
R36588 DVSS.n22369 DVSS.n22358 2.24442
R36589 DVSS.n22369 DVSS.n22355 2.24442
R36590 DVSS.n22369 DVSS.n22352 2.24442
R36591 DVSS.n22369 DVSS.n22349 2.24442
R36592 DVSS.n22369 DVSS.n22346 2.24442
R36593 DVSS.n12970 DVSS.n12961 2.24442
R36594 DVSS.n13065 DVSS.n12961 2.24442
R36595 DVSS.n13068 DVSS.n12961 2.24442
R36596 DVSS.n13071 DVSS.n12961 2.24442
R36597 DVSS.n13074 DVSS.n12961 2.24442
R36598 DVSS.n13077 DVSS.n12961 2.24442
R36599 DVSS.n13080 DVSS.n12961 2.24442
R36600 DVSS.n13083 DVSS.n12961 2.24442
R36601 DVSS.n1027 DVSS.n1015 2.24442
R36602 DVSS.n1029 DVSS.n1015 2.24442
R36603 DVSS.n1031 DVSS.n1015 2.24442
R36604 DVSS.n1033 DVSS.n1015 2.24442
R36605 DVSS.n1035 DVSS.n1015 2.24442
R36606 DVSS.n1037 DVSS.n1015 2.24442
R36607 DVSS.n1039 DVSS.n1015 2.24442
R36608 DVSS.n22381 DVSS.n1015 2.24442
R36609 DVSS.n22371 DVSS.n1173 2.24442
R36610 DVSS.n22371 DVSS.n1172 2.24442
R36611 DVSS.n22371 DVSS.n1171 2.24442
R36612 DVSS.n22371 DVSS.n1170 2.24442
R36613 DVSS.n22371 DVSS.n1169 2.24442
R36614 DVSS.n22371 DVSS.n1168 2.24442
R36615 DVSS.n22371 DVSS.n1167 2.24442
R36616 DVSS.n22371 DVSS.n1166 2.24442
R36617 DVSS.n13064 DVSS.n12959 2.24442
R36618 DVSS.n13067 DVSS.n12959 2.24442
R36619 DVSS.n13070 DVSS.n12959 2.24442
R36620 DVSS.n13073 DVSS.n12959 2.24442
R36621 DVSS.n13076 DVSS.n12959 2.24442
R36622 DVSS.n13079 DVSS.n12959 2.24442
R36623 DVSS.n13082 DVSS.n12959 2.24442
R36624 DVSS.n13085 DVSS.n12959 2.24442
R36625 DVSS.n22385 DVSS.n1041 2.24442
R36626 DVSS.n22367 DVSS.n1153 2.24442
R36627 DVSS.n13088 DVSS.n13087 2.24442
R36628 DVSS.n13093 DVSS.n12954 2.24442
R36629 DVSS.n13093 DVSS.n12950 2.24442
R36630 DVSS.n13093 DVSS.n12946 2.24442
R36631 DVSS.n13093 DVSS.n12942 2.24442
R36632 DVSS.n13093 DVSS.n12938 2.24442
R36633 DVSS.n13093 DVSS.n12934 2.24442
R36634 DVSS.n13093 DVSS.n12930 2.24442
R36635 DVSS.n13093 DVSS.n12926 2.24442
R36636 DVSS.n12956 DVSS.n384 2.24442
R36637 DVSS.n12952 DVSS.n384 2.24442
R36638 DVSS.n12948 DVSS.n384 2.24442
R36639 DVSS.n12944 DVSS.n384 2.24442
R36640 DVSS.n12940 DVSS.n384 2.24442
R36641 DVSS.n12936 DVSS.n384 2.24442
R36642 DVSS.n12932 DVSS.n384 2.24442
R36643 DVSS.n12928 DVSS.n384 2.24442
R36644 DVSS.n12924 DVSS.n384 2.24442
R36645 DVSS.n13090 DVSS.n369 2.24442
R36646 DVSS.n19625 DVSS.n19146 2.24442
R36647 DVSS.n19628 DVSS.n19146 2.24442
R36648 DVSS.n19631 DVSS.n19146 2.24442
R36649 DVSS.n19634 DVSS.n19146 2.24442
R36650 DVSS.n19637 DVSS.n19146 2.24442
R36651 DVSS.n19640 DVSS.n19146 2.24442
R36652 DVSS.n19643 DVSS.n19146 2.24442
R36653 DVSS.n19647 DVSS.n19146 2.24442
R36654 DVSS.n19627 DVSS.n19142 2.24442
R36655 DVSS.n19630 DVSS.n19142 2.24442
R36656 DVSS.n19633 DVSS.n19142 2.24442
R36657 DVSS.n19636 DVSS.n19142 2.24442
R36658 DVSS.n19639 DVSS.n19142 2.24442
R36659 DVSS.n19642 DVSS.n19142 2.24442
R36660 DVSS.n19645 DVSS.n19142 2.24442
R36661 DVSS.n19651 DVSS.n19650 2.24442
R36662 DVSS.n19139 DVSS.n13399 2.24442
R36663 DVSS.n16461 DVSS.n16251 2.24321
R36664 DVSS.n16457 DVSS.n16251 2.24321
R36665 DVSS.n16453 DVSS.n16251 2.24321
R36666 DVSS.n16450 DVSS.n16251 2.24321
R36667 DVSS.n16446 DVSS.n16251 2.24321
R36668 DVSS.n16442 DVSS.n16251 2.24321
R36669 DVSS.n16438 DVSS.n16251 2.24321
R36670 DVSS.n16434 DVSS.n16251 2.24321
R36671 DVSS.n16430 DVSS.n16251 2.24321
R36672 DVSS.n16459 DVSS.n16426 2.24321
R36673 DVSS.n16455 DVSS.n16426 2.24321
R36674 DVSS.n16448 DVSS.n16426 2.24321
R36675 DVSS.n16444 DVSS.n16426 2.24321
R36676 DVSS.n16440 DVSS.n16426 2.24321
R36677 DVSS.n16436 DVSS.n16426 2.24321
R36678 DVSS.n16432 DVSS.n16426 2.24321
R36679 DVSS.n16428 DVSS.n16426 2.24321
R36680 DVSS.n16221 DVSS.n16176 2.24321
R36681 DVSS.n16209 DVSS.n16176 2.24321
R36682 DVSS.n16207 DVSS.n16176 2.24321
R36683 DVSS.n16205 DVSS.n16176 2.24321
R36684 DVSS.n16203 DVSS.n16176 2.24321
R36685 DVSS.n16201 DVSS.n16176 2.24321
R36686 DVSS.n16198 DVSS.n16176 2.24321
R36687 DVSS.n16196 DVSS.n16176 2.24321
R36688 DVSS.n16220 DVSS.n16219 2.24321
R36689 DVSS.n16220 DVSS.n16218 2.24321
R36690 DVSS.n16220 DVSS.n16217 2.24321
R36691 DVSS.n16220 DVSS.n16216 2.24321
R36692 DVSS.n16220 DVSS.n16215 2.24321
R36693 DVSS.n16220 DVSS.n16214 2.24321
R36694 DVSS.n16220 DVSS.n16213 2.24321
R36695 DVSS.n16220 DVSS.n16212 2.24321
R36696 DVSS.n16220 DVSS.n16211 2.24321
R36697 DVSS.n16372 DVSS.n16360 2.24321
R36698 DVSS.n16370 DVSS.n16360 2.24321
R36699 DVSS.n16368 DVSS.n16360 2.24321
R36700 DVSS.n16366 DVSS.n16360 2.24321
R36701 DVSS.n16467 DVSS.n16359 2.24321
R36702 DVSS.n16468 DVSS.n16467 2.24321
R36703 DVSS.n16467 DVSS.n16375 2.24321
R36704 DVSS.n16467 DVSS.n16374 2.24321
R36705 DVSS.n16467 DVSS.n16373 2.24321
R36706 DVSS.n16548 DVSS.n16547 2.24321
R36707 DVSS.n16548 DVSS.n16546 2.24321
R36708 DVSS.n16548 DVSS.n16545 2.24321
R36709 DVSS.n16548 DVSS.n16544 2.24321
R36710 DVSS.n16548 DVSS.n16543 2.24321
R36711 DVSS.n16542 DVSS.n16541 2.24321
R36712 DVSS.n16541 DVSS.n16483 2.24321
R36713 DVSS.n16541 DVSS.n16482 2.24321
R36714 DVSS.n16541 DVSS.n16481 2.24321
R36715 DVSS.n16541 DVSS.n16480 2.24321
R36716 DVSS.n16541 DVSS.n16479 2.24321
R36717 DVSS.n15642 DVSS.n15629 2.24321
R36718 DVSS.n15640 DVSS.n15629 2.24321
R36719 DVSS.n15638 DVSS.n15629 2.24321
R36720 DVSS.n15636 DVSS.n15629 2.24321
R36721 DVSS.n18086 DVSS.n18085 2.24321
R36722 DVSS.n18085 DVSS.n15649 2.24321
R36723 DVSS.n18085 DVSS.n15648 2.24321
R36724 DVSS.n18085 DVSS.n15647 2.24321
R36725 DVSS.n18085 DVSS.n15628 2.24321
R36726 DVSS.n18112 DVSS.n18095 2.24321
R36727 DVSS.n18112 DVSS.n18094 2.24321
R36728 DVSS.n18112 DVSS.n18093 2.24321
R36729 DVSS.n18112 DVSS.n18092 2.24321
R36730 DVSS.n18112 DVSS.n18091 2.24321
R36731 DVSS.n18107 DVSS.n18090 2.24321
R36732 DVSS.n18107 DVSS.n18106 2.24321
R36733 DVSS.n18107 DVSS.n18105 2.24321
R36734 DVSS.n18107 DVSS.n18104 2.24321
R36735 DVSS.n18107 DVSS.n18103 2.24321
R36736 DVSS.n18107 DVSS.n18102 2.24321
R36737 DVSS.n11731 DVSS.n11646 2.24164
R36738 DVSS.n11980 DVSS.n11687 2.24164
R36739 DVSS.n11738 DVSS.n11646 2.24164
R36740 DVSS.n11980 DVSS.n11686 2.24164
R36741 DVSS.n11742 DVSS.n11646 2.24164
R36742 DVSS.n11980 DVSS.n11685 2.24164
R36743 DVSS.n11750 DVSS.n11646 2.24164
R36744 DVSS.n11980 DVSS.n11684 2.24164
R36745 DVSS.n11754 DVSS.n11646 2.24164
R36746 DVSS.n11980 DVSS.n11683 2.24164
R36747 DVSS.n11762 DVSS.n11646 2.24164
R36748 DVSS.n11980 DVSS.n11682 2.24164
R36749 DVSS.n11766 DVSS.n11646 2.24164
R36750 DVSS.n11980 DVSS.n11681 2.24164
R36751 DVSS.n11774 DVSS.n11646 2.24164
R36752 DVSS.n11980 DVSS.n11680 2.24164
R36753 DVSS.n11778 DVSS.n11646 2.24164
R36754 DVSS.n11980 DVSS.n11679 2.24164
R36755 DVSS.n11786 DVSS.n11646 2.24164
R36756 DVSS.n11980 DVSS.n11678 2.24164
R36757 DVSS.n11790 DVSS.n11646 2.24164
R36758 DVSS.n11980 DVSS.n11677 2.24164
R36759 DVSS.n11798 DVSS.n11646 2.24164
R36760 DVSS.n11980 DVSS.n11676 2.24164
R36761 DVSS.n11802 DVSS.n11646 2.24164
R36762 DVSS.n11980 DVSS.n11675 2.24164
R36763 DVSS.n11810 DVSS.n11646 2.24164
R36764 DVSS.n11980 DVSS.n11674 2.24164
R36765 DVSS.n11814 DVSS.n11646 2.24164
R36766 DVSS.n11980 DVSS.n11673 2.24164
R36767 DVSS.n11822 DVSS.n11646 2.24164
R36768 DVSS.n11980 DVSS.n11672 2.24164
R36769 DVSS.n11826 DVSS.n11646 2.24164
R36770 DVSS.n11980 DVSS.n11671 2.24164
R36771 DVSS.n11834 DVSS.n11646 2.24164
R36772 DVSS.n11980 DVSS.n11670 2.24164
R36773 DVSS.n11838 DVSS.n11646 2.24164
R36774 DVSS.n11980 DVSS.n11669 2.24164
R36775 DVSS.n11846 DVSS.n11646 2.24164
R36776 DVSS.n11980 DVSS.n11668 2.24164
R36777 DVSS.n11850 DVSS.n11646 2.24164
R36778 DVSS.n11980 DVSS.n11667 2.24164
R36779 DVSS.n11858 DVSS.n11646 2.24164
R36780 DVSS.n11980 DVSS.n11666 2.24164
R36781 DVSS.n11862 DVSS.n11646 2.24164
R36782 DVSS.n11980 DVSS.n11665 2.24164
R36783 DVSS.n11870 DVSS.n11646 2.24164
R36784 DVSS.n11980 DVSS.n11664 2.24164
R36785 DVSS.n11874 DVSS.n11646 2.24164
R36786 DVSS.n11980 DVSS.n11663 2.24164
R36787 DVSS.n11882 DVSS.n11646 2.24164
R36788 DVSS.n11980 DVSS.n11662 2.24164
R36789 DVSS.n11886 DVSS.n11646 2.24164
R36790 DVSS.n11980 DVSS.n11661 2.24164
R36791 DVSS.n11894 DVSS.n11646 2.24164
R36792 DVSS.n11980 DVSS.n11660 2.24164
R36793 DVSS.n11898 DVSS.n11646 2.24164
R36794 DVSS.n11980 DVSS.n11659 2.24164
R36795 DVSS.n11906 DVSS.n11646 2.24164
R36796 DVSS.n11980 DVSS.n11658 2.24164
R36797 DVSS.n11910 DVSS.n11646 2.24164
R36798 DVSS.n11980 DVSS.n11657 2.24164
R36799 DVSS.n11918 DVSS.n11646 2.24164
R36800 DVSS.n11980 DVSS.n11656 2.24164
R36801 DVSS.n11922 DVSS.n11646 2.24164
R36802 DVSS.n11980 DVSS.n11655 2.24164
R36803 DVSS.n11930 DVSS.n11646 2.24164
R36804 DVSS.n11980 DVSS.n11654 2.24164
R36805 DVSS.n11934 DVSS.n11646 2.24164
R36806 DVSS.n11980 DVSS.n11653 2.24164
R36807 DVSS.n11942 DVSS.n11646 2.24164
R36808 DVSS.n11980 DVSS.n11652 2.24164
R36809 DVSS.n11946 DVSS.n11646 2.24164
R36810 DVSS.n11980 DVSS.n11651 2.24164
R36811 DVSS.n11954 DVSS.n11646 2.24164
R36812 DVSS.n11980 DVSS.n11650 2.24164
R36813 DVSS.n11958 DVSS.n11646 2.24164
R36814 DVSS.n11980 DVSS.n11649 2.24164
R36815 DVSS.n11966 DVSS.n11646 2.24164
R36816 DVSS.n11980 DVSS.n11648 2.24164
R36817 DVSS.n11970 DVSS.n11646 2.24164
R36818 DVSS.n11980 DVSS.n11647 2.24164
R36819 DVSS.n11689 DVSS.n11646 2.24164
R36820 DVSS.n13326 DVSS.n13325 2.24164
R36821 DVSS.n13323 DVSS.n11545 2.24164
R36822 DVSS.n13326 DVSS.n11499 2.24164
R36823 DVSS.n13323 DVSS.n11544 2.24164
R36824 DVSS.n13326 DVSS.n11498 2.24164
R36825 DVSS.n13323 DVSS.n11543 2.24164
R36826 DVSS.n13326 DVSS.n11497 2.24164
R36827 DVSS.n13323 DVSS.n11542 2.24164
R36828 DVSS.n13326 DVSS.n11496 2.24164
R36829 DVSS.n13323 DVSS.n11541 2.24164
R36830 DVSS.n13326 DVSS.n11495 2.24164
R36831 DVSS.n13323 DVSS.n11540 2.24164
R36832 DVSS.n13326 DVSS.n11494 2.24164
R36833 DVSS.n13323 DVSS.n11539 2.24164
R36834 DVSS.n13326 DVSS.n11493 2.24164
R36835 DVSS.n13323 DVSS.n11538 2.24164
R36836 DVSS.n13326 DVSS.n11492 2.24164
R36837 DVSS.n13323 DVSS.n11537 2.24164
R36838 DVSS.n13326 DVSS.n11491 2.24164
R36839 DVSS.n13323 DVSS.n11536 2.24164
R36840 DVSS.n13326 DVSS.n11490 2.24164
R36841 DVSS.n13323 DVSS.n11535 2.24164
R36842 DVSS.n13326 DVSS.n11489 2.24164
R36843 DVSS.n13323 DVSS.n11534 2.24164
R36844 DVSS.n13326 DVSS.n11488 2.24164
R36845 DVSS.n13323 DVSS.n11533 2.24164
R36846 DVSS.n13326 DVSS.n11487 2.24164
R36847 DVSS.n13323 DVSS.n11532 2.24164
R36848 DVSS.n13326 DVSS.n11486 2.24164
R36849 DVSS.n13323 DVSS.n11531 2.24164
R36850 DVSS.n13326 DVSS.n11485 2.24164
R36851 DVSS.n13323 DVSS.n11530 2.24164
R36852 DVSS.n13326 DVSS.n11484 2.24164
R36853 DVSS.n13323 DVSS.n11529 2.24164
R36854 DVSS.n13326 DVSS.n11483 2.24164
R36855 DVSS.n13323 DVSS.n11528 2.24164
R36856 DVSS.n13326 DVSS.n11482 2.24164
R36857 DVSS.n13323 DVSS.n11527 2.24164
R36858 DVSS.n13326 DVSS.n11481 2.24164
R36859 DVSS.n13323 DVSS.n11526 2.24164
R36860 DVSS.n13326 DVSS.n11480 2.24164
R36861 DVSS.n13323 DVSS.n11525 2.24164
R36862 DVSS.n13326 DVSS.n11479 2.24164
R36863 DVSS.n13323 DVSS.n11524 2.24164
R36864 DVSS.n13326 DVSS.n11478 2.24164
R36865 DVSS.n13323 DVSS.n11523 2.24164
R36866 DVSS.n13326 DVSS.n11477 2.24164
R36867 DVSS.n13323 DVSS.n11522 2.24164
R36868 DVSS.n13326 DVSS.n11476 2.24164
R36869 DVSS.n13323 DVSS.n11521 2.24164
R36870 DVSS.n13326 DVSS.n11475 2.24164
R36871 DVSS.n13323 DVSS.n11520 2.24164
R36872 DVSS.n13326 DVSS.n11474 2.24164
R36873 DVSS.n13323 DVSS.n11519 2.24164
R36874 DVSS.n13326 DVSS.n11473 2.24164
R36875 DVSS.n13323 DVSS.n11518 2.24164
R36876 DVSS.n13326 DVSS.n11472 2.24164
R36877 DVSS.n13323 DVSS.n11517 2.24164
R36878 DVSS.n13326 DVSS.n11471 2.24164
R36879 DVSS.n13323 DVSS.n11516 2.24164
R36880 DVSS.n13326 DVSS.n11470 2.24164
R36881 DVSS.n13323 DVSS.n11515 2.24164
R36882 DVSS.n13326 DVSS.n11469 2.24164
R36883 DVSS.n13323 DVSS.n11514 2.24164
R36884 DVSS.n13326 DVSS.n11468 2.24164
R36885 DVSS.n13323 DVSS.n11513 2.24164
R36886 DVSS.n13326 DVSS.n11467 2.24164
R36887 DVSS.n13323 DVSS.n11512 2.24164
R36888 DVSS.n13326 DVSS.n11466 2.24164
R36889 DVSS.n13323 DVSS.n11511 2.24164
R36890 DVSS.n13326 DVSS.n11465 2.24164
R36891 DVSS.n13323 DVSS.n11510 2.24164
R36892 DVSS.n13326 DVSS.n11464 2.24164
R36893 DVSS.n13323 DVSS.n11509 2.24164
R36894 DVSS.n13326 DVSS.n11463 2.24164
R36895 DVSS.n13323 DVSS.n11508 2.24164
R36896 DVSS.n13326 DVSS.n11462 2.24164
R36897 DVSS.n13323 DVSS.n11507 2.24164
R36898 DVSS.n13326 DVSS.n11461 2.24164
R36899 DVSS.n13323 DVSS.n11506 2.24164
R36900 DVSS.n13326 DVSS.n11460 2.24164
R36901 DVSS.n13323 DVSS.n11505 2.24164
R36902 DVSS.n13326 DVSS.n11459 2.24164
R36903 DVSS.n13340 DVSS.n13339 2.24164
R36904 DVSS.n13337 DVSS.n11197 2.24164
R36905 DVSS.n13340 DVSS.n11152 2.24164
R36906 DVSS.n13337 DVSS.n11196 2.24164
R36907 DVSS.n13340 DVSS.n11151 2.24164
R36908 DVSS.n13337 DVSS.n11195 2.24164
R36909 DVSS.n13340 DVSS.n11150 2.24164
R36910 DVSS.n13337 DVSS.n11194 2.24164
R36911 DVSS.n13340 DVSS.n11149 2.24164
R36912 DVSS.n13337 DVSS.n11193 2.24164
R36913 DVSS.n13340 DVSS.n11148 2.24164
R36914 DVSS.n13337 DVSS.n11192 2.24164
R36915 DVSS.n13340 DVSS.n11147 2.24164
R36916 DVSS.n13337 DVSS.n11191 2.24164
R36917 DVSS.n13340 DVSS.n11146 2.24164
R36918 DVSS.n13337 DVSS.n11190 2.24164
R36919 DVSS.n13340 DVSS.n11145 2.24164
R36920 DVSS.n13337 DVSS.n11189 2.24164
R36921 DVSS.n13340 DVSS.n11144 2.24164
R36922 DVSS.n13337 DVSS.n11188 2.24164
R36923 DVSS.n13340 DVSS.n11143 2.24164
R36924 DVSS.n13337 DVSS.n11187 2.24164
R36925 DVSS.n13340 DVSS.n11142 2.24164
R36926 DVSS.n13337 DVSS.n11186 2.24164
R36927 DVSS.n13340 DVSS.n11141 2.24164
R36928 DVSS.n13337 DVSS.n11185 2.24164
R36929 DVSS.n13340 DVSS.n11140 2.24164
R36930 DVSS.n13337 DVSS.n11184 2.24164
R36931 DVSS.n13340 DVSS.n11139 2.24164
R36932 DVSS.n13337 DVSS.n11183 2.24164
R36933 DVSS.n13340 DVSS.n11138 2.24164
R36934 DVSS.n13337 DVSS.n11182 2.24164
R36935 DVSS.n13340 DVSS.n11137 2.24164
R36936 DVSS.n13337 DVSS.n11181 2.24164
R36937 DVSS.n13340 DVSS.n11136 2.24164
R36938 DVSS.n13337 DVSS.n11180 2.24164
R36939 DVSS.n13340 DVSS.n11135 2.24164
R36940 DVSS.n13337 DVSS.n11179 2.24164
R36941 DVSS.n13340 DVSS.n11134 2.24164
R36942 DVSS.n13337 DVSS.n11178 2.24164
R36943 DVSS.n13340 DVSS.n11133 2.24164
R36944 DVSS.n13337 DVSS.n11177 2.24164
R36945 DVSS.n13340 DVSS.n11132 2.24164
R36946 DVSS.n13337 DVSS.n11176 2.24164
R36947 DVSS.n13340 DVSS.n11131 2.24164
R36948 DVSS.n13337 DVSS.n11175 2.24164
R36949 DVSS.n13340 DVSS.n11130 2.24164
R36950 DVSS.n13337 DVSS.n11174 2.24164
R36951 DVSS.n13340 DVSS.n11129 2.24164
R36952 DVSS.n13337 DVSS.n11173 2.24164
R36953 DVSS.n13340 DVSS.n11128 2.24164
R36954 DVSS.n13337 DVSS.n11172 2.24164
R36955 DVSS.n13340 DVSS.n11127 2.24164
R36956 DVSS.n13337 DVSS.n11171 2.24164
R36957 DVSS.n13340 DVSS.n11126 2.24164
R36958 DVSS.n13337 DVSS.n11170 2.24164
R36959 DVSS.n13340 DVSS.n11125 2.24164
R36960 DVSS.n13337 DVSS.n11169 2.24164
R36961 DVSS.n13340 DVSS.n11124 2.24164
R36962 DVSS.n13337 DVSS.n11168 2.24164
R36963 DVSS.n13340 DVSS.n11123 2.24164
R36964 DVSS.n13337 DVSS.n11167 2.24164
R36965 DVSS.n13340 DVSS.n11122 2.24164
R36966 DVSS.n13337 DVSS.n11166 2.24164
R36967 DVSS.n13340 DVSS.n11121 2.24164
R36968 DVSS.n13337 DVSS.n11165 2.24164
R36969 DVSS.n13340 DVSS.n11120 2.24164
R36970 DVSS.n13337 DVSS.n11164 2.24164
R36971 DVSS.n13340 DVSS.n11119 2.24164
R36972 DVSS.n13337 DVSS.n11163 2.24164
R36973 DVSS.n13340 DVSS.n11118 2.24164
R36974 DVSS.n13337 DVSS.n11162 2.24164
R36975 DVSS.n13340 DVSS.n11117 2.24164
R36976 DVSS.n13337 DVSS.n11161 2.24164
R36977 DVSS.n13340 DVSS.n11116 2.24164
R36978 DVSS.n13337 DVSS.n11160 2.24164
R36979 DVSS.n13340 DVSS.n11115 2.24164
R36980 DVSS.n13337 DVSS.n11159 2.24164
R36981 DVSS.n13340 DVSS.n11114 2.24164
R36982 DVSS.n13337 DVSS.n11158 2.24164
R36983 DVSS.n13340 DVSS.n11113 2.24164
R36984 DVSS.n13337 DVSS.n11157 2.24164
R36985 DVSS.n13340 DVSS.n11112 2.24164
R36986 DVSS.n11101 DVSS.n1512 2.24164
R36987 DVSS.n11099 DVSS.n10766 2.24164
R36988 DVSS.n10773 DVSS.n1512 2.24164
R36989 DVSS.n10778 DVSS.n10766 2.24164
R36990 DVSS.n11091 DVSS.n1512 2.24164
R36991 DVSS.n11089 DVSS.n10766 2.24164
R36992 DVSS.n10779 DVSS.n1512 2.24164
R36993 DVSS.n10784 DVSS.n10766 2.24164
R36994 DVSS.n11081 DVSS.n1512 2.24164
R36995 DVSS.n11079 DVSS.n10766 2.24164
R36996 DVSS.n10785 DVSS.n1512 2.24164
R36997 DVSS.n10790 DVSS.n10766 2.24164
R36998 DVSS.n11071 DVSS.n1512 2.24164
R36999 DVSS.n11069 DVSS.n10766 2.24164
R37000 DVSS.n10791 DVSS.n1512 2.24164
R37001 DVSS.n10796 DVSS.n10766 2.24164
R37002 DVSS.n11061 DVSS.n1512 2.24164
R37003 DVSS.n11059 DVSS.n10766 2.24164
R37004 DVSS.n10797 DVSS.n1512 2.24164
R37005 DVSS.n10802 DVSS.n10766 2.24164
R37006 DVSS.n11051 DVSS.n1512 2.24164
R37007 DVSS.n11049 DVSS.n10766 2.24164
R37008 DVSS.n10803 DVSS.n1512 2.24164
R37009 DVSS.n10808 DVSS.n10766 2.24164
R37010 DVSS.n11041 DVSS.n1512 2.24164
R37011 DVSS.n11039 DVSS.n10766 2.24164
R37012 DVSS.n10809 DVSS.n1512 2.24164
R37013 DVSS.n10814 DVSS.n10766 2.24164
R37014 DVSS.n11031 DVSS.n1512 2.24164
R37015 DVSS.n11029 DVSS.n10766 2.24164
R37016 DVSS.n10815 DVSS.n1512 2.24164
R37017 DVSS.n10820 DVSS.n10766 2.24164
R37018 DVSS.n11021 DVSS.n1512 2.24164
R37019 DVSS.n11019 DVSS.n10766 2.24164
R37020 DVSS.n10821 DVSS.n1512 2.24164
R37021 DVSS.n10826 DVSS.n10766 2.24164
R37022 DVSS.n11011 DVSS.n1512 2.24164
R37023 DVSS.n11009 DVSS.n10766 2.24164
R37024 DVSS.n10827 DVSS.n1512 2.24164
R37025 DVSS.n10832 DVSS.n10766 2.24164
R37026 DVSS.n11001 DVSS.n1512 2.24164
R37027 DVSS.n10999 DVSS.n10766 2.24164
R37028 DVSS.n10833 DVSS.n1512 2.24164
R37029 DVSS.n10838 DVSS.n10766 2.24164
R37030 DVSS.n10991 DVSS.n1512 2.24164
R37031 DVSS.n10989 DVSS.n10766 2.24164
R37032 DVSS.n10839 DVSS.n1512 2.24164
R37033 DVSS.n10844 DVSS.n10766 2.24164
R37034 DVSS.n10981 DVSS.n1512 2.24164
R37035 DVSS.n10979 DVSS.n10766 2.24164
R37036 DVSS.n10845 DVSS.n1512 2.24164
R37037 DVSS.n10850 DVSS.n10766 2.24164
R37038 DVSS.n10971 DVSS.n1512 2.24164
R37039 DVSS.n10969 DVSS.n10766 2.24164
R37040 DVSS.n10851 DVSS.n1512 2.24164
R37041 DVSS.n10856 DVSS.n10766 2.24164
R37042 DVSS.n10961 DVSS.n1512 2.24164
R37043 DVSS.n10959 DVSS.n10766 2.24164
R37044 DVSS.n10857 DVSS.n1512 2.24164
R37045 DVSS.n10862 DVSS.n10766 2.24164
R37046 DVSS.n10951 DVSS.n1512 2.24164
R37047 DVSS.n10949 DVSS.n10766 2.24164
R37048 DVSS.n10863 DVSS.n1512 2.24164
R37049 DVSS.n10868 DVSS.n10766 2.24164
R37050 DVSS.n10941 DVSS.n1512 2.24164
R37051 DVSS.n10939 DVSS.n10766 2.24164
R37052 DVSS.n10869 DVSS.n1512 2.24164
R37053 DVSS.n10874 DVSS.n10766 2.24164
R37054 DVSS.n10931 DVSS.n1512 2.24164
R37055 DVSS.n10929 DVSS.n10766 2.24164
R37056 DVSS.n10875 DVSS.n1512 2.24164
R37057 DVSS.n10880 DVSS.n10766 2.24164
R37058 DVSS.n10921 DVSS.n1512 2.24164
R37059 DVSS.n10919 DVSS.n10766 2.24164
R37060 DVSS.n10881 DVSS.n1512 2.24164
R37061 DVSS.n10886 DVSS.n10766 2.24164
R37062 DVSS.n10911 DVSS.n1512 2.24164
R37063 DVSS.n10909 DVSS.n10766 2.24164
R37064 DVSS.n10887 DVSS.n1512 2.24164
R37065 DVSS.n10892 DVSS.n10766 2.24164
R37066 DVSS.n10901 DVSS.n1512 2.24164
R37067 DVSS.n10899 DVSS.n10766 2.24164
R37068 DVSS.n10893 DVSS.n1512 2.24164
R37069 DVSS.n1609 DVSS.n1568 2.24164
R37070 DVSS.n10754 DVSS.n1564 2.24164
R37071 DVSS.n10512 DVSS.n1568 2.24164
R37072 DVSS.n10754 DVSS.n1563 2.24164
R37073 DVSS.n10516 DVSS.n1568 2.24164
R37074 DVSS.n10754 DVSS.n1562 2.24164
R37075 DVSS.n10524 DVSS.n1568 2.24164
R37076 DVSS.n10754 DVSS.n1561 2.24164
R37077 DVSS.n10528 DVSS.n1568 2.24164
R37078 DVSS.n10754 DVSS.n1560 2.24164
R37079 DVSS.n10536 DVSS.n1568 2.24164
R37080 DVSS.n10754 DVSS.n1559 2.24164
R37081 DVSS.n10540 DVSS.n1568 2.24164
R37082 DVSS.n10754 DVSS.n1558 2.24164
R37083 DVSS.n10548 DVSS.n1568 2.24164
R37084 DVSS.n10754 DVSS.n1557 2.24164
R37085 DVSS.n10552 DVSS.n1568 2.24164
R37086 DVSS.n10754 DVSS.n1556 2.24164
R37087 DVSS.n10560 DVSS.n1568 2.24164
R37088 DVSS.n10754 DVSS.n1555 2.24164
R37089 DVSS.n10564 DVSS.n1568 2.24164
R37090 DVSS.n10754 DVSS.n1554 2.24164
R37091 DVSS.n10572 DVSS.n1568 2.24164
R37092 DVSS.n10754 DVSS.n1553 2.24164
R37093 DVSS.n10576 DVSS.n1568 2.24164
R37094 DVSS.n10754 DVSS.n1552 2.24164
R37095 DVSS.n10584 DVSS.n1568 2.24164
R37096 DVSS.n10754 DVSS.n1551 2.24164
R37097 DVSS.n10588 DVSS.n1568 2.24164
R37098 DVSS.n10754 DVSS.n1550 2.24164
R37099 DVSS.n10596 DVSS.n1568 2.24164
R37100 DVSS.n10754 DVSS.n1549 2.24164
R37101 DVSS.n10600 DVSS.n1568 2.24164
R37102 DVSS.n10754 DVSS.n1548 2.24164
R37103 DVSS.n10608 DVSS.n1568 2.24164
R37104 DVSS.n10754 DVSS.n1547 2.24164
R37105 DVSS.n10612 DVSS.n1568 2.24164
R37106 DVSS.n10754 DVSS.n1546 2.24164
R37107 DVSS.n10620 DVSS.n1568 2.24164
R37108 DVSS.n10754 DVSS.n1545 2.24164
R37109 DVSS.n10624 DVSS.n1568 2.24164
R37110 DVSS.n10754 DVSS.n1544 2.24164
R37111 DVSS.n10632 DVSS.n1568 2.24164
R37112 DVSS.n10754 DVSS.n1543 2.24164
R37113 DVSS.n10636 DVSS.n1568 2.24164
R37114 DVSS.n10754 DVSS.n1542 2.24164
R37115 DVSS.n10644 DVSS.n1568 2.24164
R37116 DVSS.n10754 DVSS.n1541 2.24164
R37117 DVSS.n10648 DVSS.n1568 2.24164
R37118 DVSS.n10754 DVSS.n1540 2.24164
R37119 DVSS.n10656 DVSS.n1568 2.24164
R37120 DVSS.n10754 DVSS.n1539 2.24164
R37121 DVSS.n10660 DVSS.n1568 2.24164
R37122 DVSS.n10754 DVSS.n1538 2.24164
R37123 DVSS.n10668 DVSS.n1568 2.24164
R37124 DVSS.n10754 DVSS.n1537 2.24164
R37125 DVSS.n10672 DVSS.n1568 2.24164
R37126 DVSS.n10754 DVSS.n1536 2.24164
R37127 DVSS.n10680 DVSS.n1568 2.24164
R37128 DVSS.n10754 DVSS.n1535 2.24164
R37129 DVSS.n10684 DVSS.n1568 2.24164
R37130 DVSS.n10754 DVSS.n1534 2.24164
R37131 DVSS.n10692 DVSS.n1568 2.24164
R37132 DVSS.n10754 DVSS.n1533 2.24164
R37133 DVSS.n10696 DVSS.n1568 2.24164
R37134 DVSS.n10754 DVSS.n1532 2.24164
R37135 DVSS.n10704 DVSS.n1568 2.24164
R37136 DVSS.n10754 DVSS.n1531 2.24164
R37137 DVSS.n10708 DVSS.n1568 2.24164
R37138 DVSS.n10754 DVSS.n1530 2.24164
R37139 DVSS.n10716 DVSS.n1568 2.24164
R37140 DVSS.n10754 DVSS.n1529 2.24164
R37141 DVSS.n10720 DVSS.n1568 2.24164
R37142 DVSS.n10754 DVSS.n1528 2.24164
R37143 DVSS.n10728 DVSS.n1568 2.24164
R37144 DVSS.n10754 DVSS.n1527 2.24164
R37145 DVSS.n10732 DVSS.n1568 2.24164
R37146 DVSS.n10754 DVSS.n1526 2.24164
R37147 DVSS.n10740 DVSS.n1568 2.24164
R37148 DVSS.n10754 DVSS.n1525 2.24164
R37149 DVSS.n10744 DVSS.n1568 2.24164
R37150 DVSS.n10754 DVSS.n1524 2.24164
R37151 DVSS.n10752 DVSS.n1568 2.24164
R37152 DVSS.n1961 DVSS.n1960 2.24164
R37153 DVSS.n1670 DVSS.n1620 2.24164
R37154 DVSS.n1961 DVSS.n1667 2.24164
R37155 DVSS.n1951 DVSS.n1620 2.24164
R37156 DVSS.n1961 DVSS.n1666 2.24164
R37157 DVSS.n1946 DVSS.n1620 2.24164
R37158 DVSS.n1961 DVSS.n1665 2.24164
R37159 DVSS.n1939 DVSS.n1620 2.24164
R37160 DVSS.n1961 DVSS.n1664 2.24164
R37161 DVSS.n1934 DVSS.n1620 2.24164
R37162 DVSS.n1961 DVSS.n1663 2.24164
R37163 DVSS.n1927 DVSS.n1620 2.24164
R37164 DVSS.n1961 DVSS.n1662 2.24164
R37165 DVSS.n1922 DVSS.n1620 2.24164
R37166 DVSS.n1961 DVSS.n1661 2.24164
R37167 DVSS.n1915 DVSS.n1620 2.24164
R37168 DVSS.n1961 DVSS.n1660 2.24164
R37169 DVSS.n1910 DVSS.n1620 2.24164
R37170 DVSS.n1961 DVSS.n1659 2.24164
R37171 DVSS.n1903 DVSS.n1620 2.24164
R37172 DVSS.n1961 DVSS.n1658 2.24164
R37173 DVSS.n1898 DVSS.n1620 2.24164
R37174 DVSS.n1961 DVSS.n1657 2.24164
R37175 DVSS.n1891 DVSS.n1620 2.24164
R37176 DVSS.n1961 DVSS.n1656 2.24164
R37177 DVSS.n1886 DVSS.n1620 2.24164
R37178 DVSS.n1961 DVSS.n1655 2.24164
R37179 DVSS.n1879 DVSS.n1620 2.24164
R37180 DVSS.n1961 DVSS.n1654 2.24164
R37181 DVSS.n1874 DVSS.n1620 2.24164
R37182 DVSS.n1961 DVSS.n1653 2.24164
R37183 DVSS.n1867 DVSS.n1620 2.24164
R37184 DVSS.n1961 DVSS.n1652 2.24164
R37185 DVSS.n1862 DVSS.n1620 2.24164
R37186 DVSS.n1961 DVSS.n1651 2.24164
R37187 DVSS.n1855 DVSS.n1620 2.24164
R37188 DVSS.n1961 DVSS.n1650 2.24164
R37189 DVSS.n1850 DVSS.n1620 2.24164
R37190 DVSS.n1961 DVSS.n1649 2.24164
R37191 DVSS.n1843 DVSS.n1620 2.24164
R37192 DVSS.n1961 DVSS.n1648 2.24164
R37193 DVSS.n1838 DVSS.n1620 2.24164
R37194 DVSS.n1961 DVSS.n1647 2.24164
R37195 DVSS.n1831 DVSS.n1620 2.24164
R37196 DVSS.n1961 DVSS.n1646 2.24164
R37197 DVSS.n1826 DVSS.n1620 2.24164
R37198 DVSS.n1961 DVSS.n1645 2.24164
R37199 DVSS.n1819 DVSS.n1620 2.24164
R37200 DVSS.n1961 DVSS.n1644 2.24164
R37201 DVSS.n1814 DVSS.n1620 2.24164
R37202 DVSS.n1961 DVSS.n1643 2.24164
R37203 DVSS.n1807 DVSS.n1620 2.24164
R37204 DVSS.n1961 DVSS.n1642 2.24164
R37205 DVSS.n1802 DVSS.n1620 2.24164
R37206 DVSS.n1961 DVSS.n1641 2.24164
R37207 DVSS.n1795 DVSS.n1620 2.24164
R37208 DVSS.n1961 DVSS.n1640 2.24164
R37209 DVSS.n1790 DVSS.n1620 2.24164
R37210 DVSS.n1961 DVSS.n1639 2.24164
R37211 DVSS.n1783 DVSS.n1620 2.24164
R37212 DVSS.n1961 DVSS.n1638 2.24164
R37213 DVSS.n1778 DVSS.n1620 2.24164
R37214 DVSS.n1961 DVSS.n1637 2.24164
R37215 DVSS.n1771 DVSS.n1620 2.24164
R37216 DVSS.n1961 DVSS.n1636 2.24164
R37217 DVSS.n1766 DVSS.n1620 2.24164
R37218 DVSS.n1961 DVSS.n1635 2.24164
R37219 DVSS.n1759 DVSS.n1620 2.24164
R37220 DVSS.n1961 DVSS.n1634 2.24164
R37221 DVSS.n1754 DVSS.n1620 2.24164
R37222 DVSS.n1961 DVSS.n1633 2.24164
R37223 DVSS.n1747 DVSS.n1620 2.24164
R37224 DVSS.n1961 DVSS.n1632 2.24164
R37225 DVSS.n1742 DVSS.n1620 2.24164
R37226 DVSS.n1961 DVSS.n1631 2.24164
R37227 DVSS.n1735 DVSS.n1620 2.24164
R37228 DVSS.n1961 DVSS.n1630 2.24164
R37229 DVSS.n1730 DVSS.n1620 2.24164
R37230 DVSS.n1961 DVSS.n1629 2.24164
R37231 DVSS.n1723 DVSS.n1620 2.24164
R37232 DVSS.n1961 DVSS.n1628 2.24164
R37233 DVSS.n1718 DVSS.n1620 2.24164
R37234 DVSS.n1961 DVSS.n1627 2.24164
R37235 DVSS.n10451 DVSS.n2013 2.24164
R37236 DVSS.n10475 DVSS.n2008 2.24164
R37237 DVSS.n10448 DVSS.n2013 2.24164
R37238 DVSS.n10475 DVSS.n2007 2.24164
R37239 DVSS.n10441 DVSS.n2013 2.24164
R37240 DVSS.n10475 DVSS.n2006 2.24164
R37241 DVSS.n10436 DVSS.n2013 2.24164
R37242 DVSS.n10475 DVSS.n2005 2.24164
R37243 DVSS.n10429 DVSS.n2013 2.24164
R37244 DVSS.n10475 DVSS.n2004 2.24164
R37245 DVSS.n10424 DVSS.n2013 2.24164
R37246 DVSS.n10475 DVSS.n2003 2.24164
R37247 DVSS.n10417 DVSS.n2013 2.24164
R37248 DVSS.n10475 DVSS.n2002 2.24164
R37249 DVSS.n10412 DVSS.n2013 2.24164
R37250 DVSS.n10475 DVSS.n2001 2.24164
R37251 DVSS.n10405 DVSS.n2013 2.24164
R37252 DVSS.n10475 DVSS.n2000 2.24164
R37253 DVSS.n10400 DVSS.n2013 2.24164
R37254 DVSS.n10475 DVSS.n1999 2.24164
R37255 DVSS.n10393 DVSS.n2013 2.24164
R37256 DVSS.n10475 DVSS.n1998 2.24164
R37257 DVSS.n10388 DVSS.n2013 2.24164
R37258 DVSS.n10475 DVSS.n1997 2.24164
R37259 DVSS.n10381 DVSS.n2013 2.24164
R37260 DVSS.n10475 DVSS.n1996 2.24164
R37261 DVSS.n10376 DVSS.n2013 2.24164
R37262 DVSS.n10475 DVSS.n1995 2.24164
R37263 DVSS.n10369 DVSS.n2013 2.24164
R37264 DVSS.n10475 DVSS.n1994 2.24164
R37265 DVSS.n10364 DVSS.n2013 2.24164
R37266 DVSS.n10475 DVSS.n1993 2.24164
R37267 DVSS.n10357 DVSS.n2013 2.24164
R37268 DVSS.n10475 DVSS.n1992 2.24164
R37269 DVSS.n10352 DVSS.n2013 2.24164
R37270 DVSS.n10475 DVSS.n1991 2.24164
R37271 DVSS.n10345 DVSS.n2013 2.24164
R37272 DVSS.n10475 DVSS.n1990 2.24164
R37273 DVSS.n10340 DVSS.n2013 2.24164
R37274 DVSS.n10475 DVSS.n1989 2.24164
R37275 DVSS.n10333 DVSS.n2013 2.24164
R37276 DVSS.n10475 DVSS.n1988 2.24164
R37277 DVSS.n10328 DVSS.n2013 2.24164
R37278 DVSS.n10475 DVSS.n1987 2.24164
R37279 DVSS.n10321 DVSS.n2013 2.24164
R37280 DVSS.n10475 DVSS.n1986 2.24164
R37281 DVSS.n10316 DVSS.n2013 2.24164
R37282 DVSS.n10475 DVSS.n1985 2.24164
R37283 DVSS.n10309 DVSS.n2013 2.24164
R37284 DVSS.n10475 DVSS.n1984 2.24164
R37285 DVSS.n10304 DVSS.n2013 2.24164
R37286 DVSS.n10475 DVSS.n1983 2.24164
R37287 DVSS.n10297 DVSS.n2013 2.24164
R37288 DVSS.n10475 DVSS.n1982 2.24164
R37289 DVSS.n10292 DVSS.n2013 2.24164
R37290 DVSS.n10475 DVSS.n1981 2.24164
R37291 DVSS.n10285 DVSS.n2013 2.24164
R37292 DVSS.n10475 DVSS.n1980 2.24164
R37293 DVSS.n10280 DVSS.n2013 2.24164
R37294 DVSS.n10475 DVSS.n1979 2.24164
R37295 DVSS.n10273 DVSS.n2013 2.24164
R37296 DVSS.n10475 DVSS.n1978 2.24164
R37297 DVSS.n10268 DVSS.n2013 2.24164
R37298 DVSS.n10475 DVSS.n1977 2.24164
R37299 DVSS.n10261 DVSS.n2013 2.24164
R37300 DVSS.n10475 DVSS.n1976 2.24164
R37301 DVSS.n10256 DVSS.n2013 2.24164
R37302 DVSS.n10475 DVSS.n1975 2.24164
R37303 DVSS.n10249 DVSS.n2013 2.24164
R37304 DVSS.n10475 DVSS.n1974 2.24164
R37305 DVSS.n10244 DVSS.n2013 2.24164
R37306 DVSS.n10475 DVSS.n1973 2.24164
R37307 DVSS.n10237 DVSS.n2013 2.24164
R37308 DVSS.n10475 DVSS.n1972 2.24164
R37309 DVSS.n10232 DVSS.n2013 2.24164
R37310 DVSS.n10475 DVSS.n1971 2.24164
R37311 DVSS.n10225 DVSS.n2013 2.24164
R37312 DVSS.n10475 DVSS.n1970 2.24164
R37313 DVSS.n10220 DVSS.n2013 2.24164
R37314 DVSS.n10475 DVSS.n1969 2.24164
R37315 DVSS.n10213 DVSS.n2013 2.24164
R37316 DVSS.n10475 DVSS.n1968 2.24164
R37317 DVSS.n10473 DVSS.n2013 2.24164
R37318 DVSS.n2114 DVSS.n2073 2.24164
R37319 DVSS.n10166 DVSS.n2068 2.24164
R37320 DVSS.n2123 DVSS.n2073 2.24164
R37321 DVSS.n10166 DVSS.n2067 2.24164
R37322 DVSS.n2127 DVSS.n2073 2.24164
R37323 DVSS.n10166 DVSS.n2066 2.24164
R37324 DVSS.n2135 DVSS.n2073 2.24164
R37325 DVSS.n10166 DVSS.n2065 2.24164
R37326 DVSS.n2139 DVSS.n2073 2.24164
R37327 DVSS.n10166 DVSS.n2064 2.24164
R37328 DVSS.n2147 DVSS.n2073 2.24164
R37329 DVSS.n10166 DVSS.n2063 2.24164
R37330 DVSS.n2151 DVSS.n2073 2.24164
R37331 DVSS.n10166 DVSS.n2062 2.24164
R37332 DVSS.n2159 DVSS.n2073 2.24164
R37333 DVSS.n10166 DVSS.n2061 2.24164
R37334 DVSS.n2163 DVSS.n2073 2.24164
R37335 DVSS.n10166 DVSS.n2060 2.24164
R37336 DVSS.n2171 DVSS.n2073 2.24164
R37337 DVSS.n10166 DVSS.n2059 2.24164
R37338 DVSS.n2175 DVSS.n2073 2.24164
R37339 DVSS.n10166 DVSS.n2058 2.24164
R37340 DVSS.n2183 DVSS.n2073 2.24164
R37341 DVSS.n10166 DVSS.n2057 2.24164
R37342 DVSS.n2187 DVSS.n2073 2.24164
R37343 DVSS.n10166 DVSS.n2056 2.24164
R37344 DVSS.n2195 DVSS.n2073 2.24164
R37345 DVSS.n10166 DVSS.n2055 2.24164
R37346 DVSS.n2199 DVSS.n2073 2.24164
R37347 DVSS.n10166 DVSS.n2054 2.24164
R37348 DVSS.n2207 DVSS.n2073 2.24164
R37349 DVSS.n10166 DVSS.n2053 2.24164
R37350 DVSS.n2211 DVSS.n2073 2.24164
R37351 DVSS.n10166 DVSS.n2052 2.24164
R37352 DVSS.n2219 DVSS.n2073 2.24164
R37353 DVSS.n10166 DVSS.n2051 2.24164
R37354 DVSS.n2223 DVSS.n2073 2.24164
R37355 DVSS.n10166 DVSS.n2050 2.24164
R37356 DVSS.n2231 DVSS.n2073 2.24164
R37357 DVSS.n10166 DVSS.n2049 2.24164
R37358 DVSS.n2235 DVSS.n2073 2.24164
R37359 DVSS.n10166 DVSS.n2048 2.24164
R37360 DVSS.n2243 DVSS.n2073 2.24164
R37361 DVSS.n10166 DVSS.n2047 2.24164
R37362 DVSS.n2247 DVSS.n2073 2.24164
R37363 DVSS.n10166 DVSS.n2046 2.24164
R37364 DVSS.n2255 DVSS.n2073 2.24164
R37365 DVSS.n10166 DVSS.n2045 2.24164
R37366 DVSS.n2259 DVSS.n2073 2.24164
R37367 DVSS.n10166 DVSS.n2044 2.24164
R37368 DVSS.n2267 DVSS.n2073 2.24164
R37369 DVSS.n10166 DVSS.n2043 2.24164
R37370 DVSS.n2271 DVSS.n2073 2.24164
R37371 DVSS.n10166 DVSS.n2042 2.24164
R37372 DVSS.n2279 DVSS.n2073 2.24164
R37373 DVSS.n10166 DVSS.n2041 2.24164
R37374 DVSS.n2283 DVSS.n2073 2.24164
R37375 DVSS.n10166 DVSS.n2040 2.24164
R37376 DVSS.n2291 DVSS.n2073 2.24164
R37377 DVSS.n10166 DVSS.n2039 2.24164
R37378 DVSS.n2295 DVSS.n2073 2.24164
R37379 DVSS.n10166 DVSS.n2038 2.24164
R37380 DVSS.n2303 DVSS.n2073 2.24164
R37381 DVSS.n10166 DVSS.n2037 2.24164
R37382 DVSS.n2307 DVSS.n2073 2.24164
R37383 DVSS.n10166 DVSS.n2036 2.24164
R37384 DVSS.n2315 DVSS.n2073 2.24164
R37385 DVSS.n10166 DVSS.n2035 2.24164
R37386 DVSS.n2319 DVSS.n2073 2.24164
R37387 DVSS.n10166 DVSS.n2034 2.24164
R37388 DVSS.n2327 DVSS.n2073 2.24164
R37389 DVSS.n10166 DVSS.n2033 2.24164
R37390 DVSS.n2331 DVSS.n2073 2.24164
R37391 DVSS.n10166 DVSS.n2032 2.24164
R37392 DVSS.n2339 DVSS.n2073 2.24164
R37393 DVSS.n10166 DVSS.n2031 2.24164
R37394 DVSS.n2343 DVSS.n2073 2.24164
R37395 DVSS.n10166 DVSS.n2030 2.24164
R37396 DVSS.n2351 DVSS.n2073 2.24164
R37397 DVSS.n10166 DVSS.n2029 2.24164
R37398 DVSS.n2355 DVSS.n2073 2.24164
R37399 DVSS.n10166 DVSS.n2028 2.24164
R37400 DVSS.n10164 DVSS.n2073 2.24164
R37401 DVSS.n2456 DVSS.n2415 2.24164
R37402 DVSS.n10141 DVSS.n2411 2.24164
R37403 DVSS.n2465 DVSS.n2415 2.24164
R37404 DVSS.n10141 DVSS.n2410 2.24164
R37405 DVSS.n2469 DVSS.n2415 2.24164
R37406 DVSS.n10141 DVSS.n2409 2.24164
R37407 DVSS.n2477 DVSS.n2415 2.24164
R37408 DVSS.n10141 DVSS.n2408 2.24164
R37409 DVSS.n2481 DVSS.n2415 2.24164
R37410 DVSS.n10141 DVSS.n2407 2.24164
R37411 DVSS.n2489 DVSS.n2415 2.24164
R37412 DVSS.n10141 DVSS.n2406 2.24164
R37413 DVSS.n2493 DVSS.n2415 2.24164
R37414 DVSS.n10141 DVSS.n2405 2.24164
R37415 DVSS.n2501 DVSS.n2415 2.24164
R37416 DVSS.n10141 DVSS.n2404 2.24164
R37417 DVSS.n2505 DVSS.n2415 2.24164
R37418 DVSS.n10141 DVSS.n2403 2.24164
R37419 DVSS.n2513 DVSS.n2415 2.24164
R37420 DVSS.n10141 DVSS.n2402 2.24164
R37421 DVSS.n2517 DVSS.n2415 2.24164
R37422 DVSS.n10141 DVSS.n2401 2.24164
R37423 DVSS.n2525 DVSS.n2415 2.24164
R37424 DVSS.n10141 DVSS.n2400 2.24164
R37425 DVSS.n2529 DVSS.n2415 2.24164
R37426 DVSS.n10141 DVSS.n2399 2.24164
R37427 DVSS.n2537 DVSS.n2415 2.24164
R37428 DVSS.n10141 DVSS.n2398 2.24164
R37429 DVSS.n2541 DVSS.n2415 2.24164
R37430 DVSS.n10141 DVSS.n2397 2.24164
R37431 DVSS.n2549 DVSS.n2415 2.24164
R37432 DVSS.n10141 DVSS.n2396 2.24164
R37433 DVSS.n2553 DVSS.n2415 2.24164
R37434 DVSS.n10141 DVSS.n2395 2.24164
R37435 DVSS.n2561 DVSS.n2415 2.24164
R37436 DVSS.n10141 DVSS.n2394 2.24164
R37437 DVSS.n2565 DVSS.n2415 2.24164
R37438 DVSS.n10141 DVSS.n2393 2.24164
R37439 DVSS.n2573 DVSS.n2415 2.24164
R37440 DVSS.n10141 DVSS.n2392 2.24164
R37441 DVSS.n2577 DVSS.n2415 2.24164
R37442 DVSS.n10141 DVSS.n2391 2.24164
R37443 DVSS.n2585 DVSS.n2415 2.24164
R37444 DVSS.n10141 DVSS.n2390 2.24164
R37445 DVSS.n2589 DVSS.n2415 2.24164
R37446 DVSS.n10141 DVSS.n2389 2.24164
R37447 DVSS.n2597 DVSS.n2415 2.24164
R37448 DVSS.n10141 DVSS.n2388 2.24164
R37449 DVSS.n2601 DVSS.n2415 2.24164
R37450 DVSS.n10141 DVSS.n2387 2.24164
R37451 DVSS.n2609 DVSS.n2415 2.24164
R37452 DVSS.n10141 DVSS.n2386 2.24164
R37453 DVSS.n2613 DVSS.n2415 2.24164
R37454 DVSS.n10141 DVSS.n2385 2.24164
R37455 DVSS.n2621 DVSS.n2415 2.24164
R37456 DVSS.n10141 DVSS.n2384 2.24164
R37457 DVSS.n2625 DVSS.n2415 2.24164
R37458 DVSS.n10141 DVSS.n2383 2.24164
R37459 DVSS.n2633 DVSS.n2415 2.24164
R37460 DVSS.n10141 DVSS.n2382 2.24164
R37461 DVSS.n2637 DVSS.n2415 2.24164
R37462 DVSS.n10141 DVSS.n2381 2.24164
R37463 DVSS.n2645 DVSS.n2415 2.24164
R37464 DVSS.n10141 DVSS.n2380 2.24164
R37465 DVSS.n2649 DVSS.n2415 2.24164
R37466 DVSS.n10141 DVSS.n2379 2.24164
R37467 DVSS.n2657 DVSS.n2415 2.24164
R37468 DVSS.n10141 DVSS.n2378 2.24164
R37469 DVSS.n2661 DVSS.n2415 2.24164
R37470 DVSS.n10141 DVSS.n2377 2.24164
R37471 DVSS.n2669 DVSS.n2415 2.24164
R37472 DVSS.n10141 DVSS.n2376 2.24164
R37473 DVSS.n2673 DVSS.n2415 2.24164
R37474 DVSS.n10141 DVSS.n2375 2.24164
R37475 DVSS.n2681 DVSS.n2415 2.24164
R37476 DVSS.n10141 DVSS.n2374 2.24164
R37477 DVSS.n2685 DVSS.n2415 2.24164
R37478 DVSS.n10141 DVSS.n2373 2.24164
R37479 DVSS.n2693 DVSS.n2415 2.24164
R37480 DVSS.n10141 DVSS.n2372 2.24164
R37481 DVSS.n2697 DVSS.n2415 2.24164
R37482 DVSS.n10141 DVSS.n2371 2.24164
R37483 DVSS.n10139 DVSS.n2415 2.24164
R37484 DVSS.n9861 DVSS.n2718 2.24164
R37485 DVSS.n9863 DVSS.n2720 2.24164
R37486 DVSS.n9865 DVSS.n2718 2.24164
R37487 DVSS.n9855 DVSS.n2720 2.24164
R37488 DVSS.n9873 DVSS.n2718 2.24164
R37489 DVSS.n9875 DVSS.n2720 2.24164
R37490 DVSS.n9877 DVSS.n2718 2.24164
R37491 DVSS.n9851 DVSS.n2720 2.24164
R37492 DVSS.n9885 DVSS.n2718 2.24164
R37493 DVSS.n9887 DVSS.n2720 2.24164
R37494 DVSS.n9889 DVSS.n2718 2.24164
R37495 DVSS.n9847 DVSS.n2720 2.24164
R37496 DVSS.n9897 DVSS.n2718 2.24164
R37497 DVSS.n9899 DVSS.n2720 2.24164
R37498 DVSS.n9901 DVSS.n2718 2.24164
R37499 DVSS.n9843 DVSS.n2720 2.24164
R37500 DVSS.n9909 DVSS.n2718 2.24164
R37501 DVSS.n9911 DVSS.n2720 2.24164
R37502 DVSS.n9913 DVSS.n2718 2.24164
R37503 DVSS.n9839 DVSS.n2720 2.24164
R37504 DVSS.n9921 DVSS.n2718 2.24164
R37505 DVSS.n9923 DVSS.n2720 2.24164
R37506 DVSS.n9925 DVSS.n2718 2.24164
R37507 DVSS.n9835 DVSS.n2720 2.24164
R37508 DVSS.n9933 DVSS.n2718 2.24164
R37509 DVSS.n9935 DVSS.n2720 2.24164
R37510 DVSS.n9937 DVSS.n2718 2.24164
R37511 DVSS.n9831 DVSS.n2720 2.24164
R37512 DVSS.n9945 DVSS.n2718 2.24164
R37513 DVSS.n9947 DVSS.n2720 2.24164
R37514 DVSS.n9949 DVSS.n2718 2.24164
R37515 DVSS.n9827 DVSS.n2720 2.24164
R37516 DVSS.n9957 DVSS.n2718 2.24164
R37517 DVSS.n9959 DVSS.n2720 2.24164
R37518 DVSS.n9961 DVSS.n2718 2.24164
R37519 DVSS.n9823 DVSS.n2720 2.24164
R37520 DVSS.n9969 DVSS.n2718 2.24164
R37521 DVSS.n9971 DVSS.n2720 2.24164
R37522 DVSS.n9973 DVSS.n2718 2.24164
R37523 DVSS.n9819 DVSS.n2720 2.24164
R37524 DVSS.n9981 DVSS.n2718 2.24164
R37525 DVSS.n9983 DVSS.n2720 2.24164
R37526 DVSS.n9985 DVSS.n2718 2.24164
R37527 DVSS.n9815 DVSS.n2720 2.24164
R37528 DVSS.n9993 DVSS.n2718 2.24164
R37529 DVSS.n9995 DVSS.n2720 2.24164
R37530 DVSS.n9997 DVSS.n2718 2.24164
R37531 DVSS.n9811 DVSS.n2720 2.24164
R37532 DVSS.n10005 DVSS.n2718 2.24164
R37533 DVSS.n10007 DVSS.n2720 2.24164
R37534 DVSS.n10009 DVSS.n2718 2.24164
R37535 DVSS.n9807 DVSS.n2720 2.24164
R37536 DVSS.n10017 DVSS.n2718 2.24164
R37537 DVSS.n10019 DVSS.n2720 2.24164
R37538 DVSS.n10021 DVSS.n2718 2.24164
R37539 DVSS.n9803 DVSS.n2720 2.24164
R37540 DVSS.n10029 DVSS.n2718 2.24164
R37541 DVSS.n10031 DVSS.n2720 2.24164
R37542 DVSS.n10033 DVSS.n2718 2.24164
R37543 DVSS.n9799 DVSS.n2720 2.24164
R37544 DVSS.n10041 DVSS.n2718 2.24164
R37545 DVSS.n10043 DVSS.n2720 2.24164
R37546 DVSS.n10045 DVSS.n2718 2.24164
R37547 DVSS.n9795 DVSS.n2720 2.24164
R37548 DVSS.n10053 DVSS.n2718 2.24164
R37549 DVSS.n10055 DVSS.n2720 2.24164
R37550 DVSS.n10057 DVSS.n2718 2.24164
R37551 DVSS.n9791 DVSS.n2720 2.24164
R37552 DVSS.n10065 DVSS.n2718 2.24164
R37553 DVSS.n10067 DVSS.n2720 2.24164
R37554 DVSS.n10069 DVSS.n2718 2.24164
R37555 DVSS.n9787 DVSS.n2720 2.24164
R37556 DVSS.n10077 DVSS.n2718 2.24164
R37557 DVSS.n10079 DVSS.n2720 2.24164
R37558 DVSS.n10081 DVSS.n2718 2.24164
R37559 DVSS.n9783 DVSS.n2720 2.24164
R37560 DVSS.n10089 DVSS.n2718 2.24164
R37561 DVSS.n10091 DVSS.n2720 2.24164
R37562 DVSS.n10093 DVSS.n2718 2.24164
R37563 DVSS.n9779 DVSS.n2720 2.24164
R37564 DVSS.n10102 DVSS.n2718 2.24164
R37565 DVSS.n10104 DVSS.n2720 2.24164
R37566 DVSS.n10106 DVSS.n2718 2.24164
R37567 DVSS.n9759 DVSS.n9758 2.24164
R37568 DVSS.n9467 DVSS.n2728 2.24164
R37569 DVSS.n9759 DVSS.n2780 2.24164
R37570 DVSS.n9749 DVSS.n2728 2.24164
R37571 DVSS.n9759 DVSS.n2779 2.24164
R37572 DVSS.n9744 DVSS.n2728 2.24164
R37573 DVSS.n9759 DVSS.n2778 2.24164
R37574 DVSS.n9737 DVSS.n2728 2.24164
R37575 DVSS.n9759 DVSS.n2777 2.24164
R37576 DVSS.n9732 DVSS.n2728 2.24164
R37577 DVSS.n9759 DVSS.n2776 2.24164
R37578 DVSS.n9725 DVSS.n2728 2.24164
R37579 DVSS.n9759 DVSS.n2775 2.24164
R37580 DVSS.n9720 DVSS.n2728 2.24164
R37581 DVSS.n9759 DVSS.n2774 2.24164
R37582 DVSS.n9713 DVSS.n2728 2.24164
R37583 DVSS.n9759 DVSS.n2773 2.24164
R37584 DVSS.n9708 DVSS.n2728 2.24164
R37585 DVSS.n9759 DVSS.n2772 2.24164
R37586 DVSS.n9701 DVSS.n2728 2.24164
R37587 DVSS.n9759 DVSS.n2771 2.24164
R37588 DVSS.n9696 DVSS.n2728 2.24164
R37589 DVSS.n9759 DVSS.n2770 2.24164
R37590 DVSS.n9689 DVSS.n2728 2.24164
R37591 DVSS.n9759 DVSS.n2769 2.24164
R37592 DVSS.n9684 DVSS.n2728 2.24164
R37593 DVSS.n9759 DVSS.n2768 2.24164
R37594 DVSS.n9677 DVSS.n2728 2.24164
R37595 DVSS.n9759 DVSS.n2767 2.24164
R37596 DVSS.n9672 DVSS.n2728 2.24164
R37597 DVSS.n9759 DVSS.n2766 2.24164
R37598 DVSS.n9665 DVSS.n2728 2.24164
R37599 DVSS.n9759 DVSS.n2765 2.24164
R37600 DVSS.n9660 DVSS.n2728 2.24164
R37601 DVSS.n9759 DVSS.n2764 2.24164
R37602 DVSS.n9653 DVSS.n2728 2.24164
R37603 DVSS.n9759 DVSS.n2763 2.24164
R37604 DVSS.n9648 DVSS.n2728 2.24164
R37605 DVSS.n9759 DVSS.n2762 2.24164
R37606 DVSS.n9641 DVSS.n2728 2.24164
R37607 DVSS.n9759 DVSS.n2761 2.24164
R37608 DVSS.n9636 DVSS.n2728 2.24164
R37609 DVSS.n9759 DVSS.n2760 2.24164
R37610 DVSS.n9629 DVSS.n2728 2.24164
R37611 DVSS.n9759 DVSS.n2759 2.24164
R37612 DVSS.n9624 DVSS.n2728 2.24164
R37613 DVSS.n9759 DVSS.n2758 2.24164
R37614 DVSS.n9617 DVSS.n2728 2.24164
R37615 DVSS.n9759 DVSS.n2757 2.24164
R37616 DVSS.n9612 DVSS.n2728 2.24164
R37617 DVSS.n9759 DVSS.n2756 2.24164
R37618 DVSS.n9605 DVSS.n2728 2.24164
R37619 DVSS.n9759 DVSS.n2755 2.24164
R37620 DVSS.n9600 DVSS.n2728 2.24164
R37621 DVSS.n9759 DVSS.n2754 2.24164
R37622 DVSS.n9593 DVSS.n2728 2.24164
R37623 DVSS.n9759 DVSS.n2753 2.24164
R37624 DVSS.n9588 DVSS.n2728 2.24164
R37625 DVSS.n9759 DVSS.n2752 2.24164
R37626 DVSS.n9581 DVSS.n2728 2.24164
R37627 DVSS.n9759 DVSS.n2751 2.24164
R37628 DVSS.n9576 DVSS.n2728 2.24164
R37629 DVSS.n9759 DVSS.n2750 2.24164
R37630 DVSS.n9569 DVSS.n2728 2.24164
R37631 DVSS.n9759 DVSS.n2749 2.24164
R37632 DVSS.n9564 DVSS.n2728 2.24164
R37633 DVSS.n9759 DVSS.n2748 2.24164
R37634 DVSS.n9557 DVSS.n2728 2.24164
R37635 DVSS.n9759 DVSS.n2747 2.24164
R37636 DVSS.n9552 DVSS.n2728 2.24164
R37637 DVSS.n9759 DVSS.n2746 2.24164
R37638 DVSS.n9545 DVSS.n2728 2.24164
R37639 DVSS.n9759 DVSS.n2745 2.24164
R37640 DVSS.n9540 DVSS.n2728 2.24164
R37641 DVSS.n9759 DVSS.n2744 2.24164
R37642 DVSS.n9533 DVSS.n2728 2.24164
R37643 DVSS.n9759 DVSS.n2743 2.24164
R37644 DVSS.n9528 DVSS.n2728 2.24164
R37645 DVSS.n9759 DVSS.n2742 2.24164
R37646 DVSS.n9521 DVSS.n2728 2.24164
R37647 DVSS.n9759 DVSS.n2741 2.24164
R37648 DVSS.n9516 DVSS.n2728 2.24164
R37649 DVSS.n9759 DVSS.n2740 2.24164
R37650 DVSS.n2872 DVSS.n2831 2.24164
R37651 DVSS.n9455 DVSS.n2828 2.24164
R37652 DVSS.n9212 DVSS.n2831 2.24164
R37653 DVSS.n9455 DVSS.n2827 2.24164
R37654 DVSS.n9216 DVSS.n2831 2.24164
R37655 DVSS.n9455 DVSS.n2826 2.24164
R37656 DVSS.n9224 DVSS.n2831 2.24164
R37657 DVSS.n9455 DVSS.n2825 2.24164
R37658 DVSS.n9228 DVSS.n2831 2.24164
R37659 DVSS.n9455 DVSS.n2824 2.24164
R37660 DVSS.n9236 DVSS.n2831 2.24164
R37661 DVSS.n9455 DVSS.n2823 2.24164
R37662 DVSS.n9240 DVSS.n2831 2.24164
R37663 DVSS.n9455 DVSS.n2822 2.24164
R37664 DVSS.n9248 DVSS.n2831 2.24164
R37665 DVSS.n9455 DVSS.n2821 2.24164
R37666 DVSS.n9252 DVSS.n2831 2.24164
R37667 DVSS.n9455 DVSS.n2820 2.24164
R37668 DVSS.n9260 DVSS.n2831 2.24164
R37669 DVSS.n9455 DVSS.n2819 2.24164
R37670 DVSS.n9264 DVSS.n2831 2.24164
R37671 DVSS.n9455 DVSS.n2818 2.24164
R37672 DVSS.n9272 DVSS.n2831 2.24164
R37673 DVSS.n9455 DVSS.n2817 2.24164
R37674 DVSS.n9276 DVSS.n2831 2.24164
R37675 DVSS.n9455 DVSS.n2816 2.24164
R37676 DVSS.n9284 DVSS.n2831 2.24164
R37677 DVSS.n9455 DVSS.n2815 2.24164
R37678 DVSS.n9288 DVSS.n2831 2.24164
R37679 DVSS.n9455 DVSS.n2814 2.24164
R37680 DVSS.n9296 DVSS.n2831 2.24164
R37681 DVSS.n9455 DVSS.n2813 2.24164
R37682 DVSS.n9300 DVSS.n2831 2.24164
R37683 DVSS.n9455 DVSS.n2812 2.24164
R37684 DVSS.n9308 DVSS.n2831 2.24164
R37685 DVSS.n9455 DVSS.n2811 2.24164
R37686 DVSS.n9312 DVSS.n2831 2.24164
R37687 DVSS.n9455 DVSS.n2810 2.24164
R37688 DVSS.n9320 DVSS.n2831 2.24164
R37689 DVSS.n9455 DVSS.n2809 2.24164
R37690 DVSS.n9324 DVSS.n2831 2.24164
R37691 DVSS.n9455 DVSS.n2808 2.24164
R37692 DVSS.n9332 DVSS.n2831 2.24164
R37693 DVSS.n9455 DVSS.n2807 2.24164
R37694 DVSS.n9336 DVSS.n2831 2.24164
R37695 DVSS.n9455 DVSS.n2806 2.24164
R37696 DVSS.n9344 DVSS.n2831 2.24164
R37697 DVSS.n9455 DVSS.n2805 2.24164
R37698 DVSS.n9348 DVSS.n2831 2.24164
R37699 DVSS.n9455 DVSS.n2804 2.24164
R37700 DVSS.n9356 DVSS.n2831 2.24164
R37701 DVSS.n9455 DVSS.n2803 2.24164
R37702 DVSS.n9360 DVSS.n2831 2.24164
R37703 DVSS.n9455 DVSS.n2802 2.24164
R37704 DVSS.n9368 DVSS.n2831 2.24164
R37705 DVSS.n9455 DVSS.n2801 2.24164
R37706 DVSS.n9372 DVSS.n2831 2.24164
R37707 DVSS.n9455 DVSS.n2800 2.24164
R37708 DVSS.n9380 DVSS.n2831 2.24164
R37709 DVSS.n9455 DVSS.n2799 2.24164
R37710 DVSS.n9384 DVSS.n2831 2.24164
R37711 DVSS.n9455 DVSS.n2798 2.24164
R37712 DVSS.n9392 DVSS.n2831 2.24164
R37713 DVSS.n9455 DVSS.n2797 2.24164
R37714 DVSS.n9396 DVSS.n2831 2.24164
R37715 DVSS.n9455 DVSS.n2796 2.24164
R37716 DVSS.n9404 DVSS.n2831 2.24164
R37717 DVSS.n9455 DVSS.n2795 2.24164
R37718 DVSS.n9408 DVSS.n2831 2.24164
R37719 DVSS.n9455 DVSS.n2794 2.24164
R37720 DVSS.n9416 DVSS.n2831 2.24164
R37721 DVSS.n9455 DVSS.n2793 2.24164
R37722 DVSS.n9420 DVSS.n2831 2.24164
R37723 DVSS.n9455 DVSS.n2792 2.24164
R37724 DVSS.n9428 DVSS.n2831 2.24164
R37725 DVSS.n9455 DVSS.n2791 2.24164
R37726 DVSS.n9432 DVSS.n2831 2.24164
R37727 DVSS.n9455 DVSS.n2790 2.24164
R37728 DVSS.n9440 DVSS.n2831 2.24164
R37729 DVSS.n9455 DVSS.n2789 2.24164
R37730 DVSS.n9444 DVSS.n2831 2.24164
R37731 DVSS.n9455 DVSS.n2788 2.24164
R37732 DVSS.n9453 DVSS.n2831 2.24164
R37733 DVSS.n9187 DVSS.n9186 2.24164
R37734 DVSS.n9184 DVSS.n2978 2.24164
R37735 DVSS.n9187 DVSS.n2931 2.24164
R37736 DVSS.n9184 DVSS.n2977 2.24164
R37737 DVSS.n9187 DVSS.n2930 2.24164
R37738 DVSS.n9184 DVSS.n2976 2.24164
R37739 DVSS.n9187 DVSS.n2929 2.24164
R37740 DVSS.n9184 DVSS.n2975 2.24164
R37741 DVSS.n9187 DVSS.n2928 2.24164
R37742 DVSS.n9184 DVSS.n2974 2.24164
R37743 DVSS.n9187 DVSS.n2927 2.24164
R37744 DVSS.n9184 DVSS.n2973 2.24164
R37745 DVSS.n9187 DVSS.n2926 2.24164
R37746 DVSS.n9184 DVSS.n2972 2.24164
R37747 DVSS.n9187 DVSS.n2925 2.24164
R37748 DVSS.n9184 DVSS.n2971 2.24164
R37749 DVSS.n9187 DVSS.n2924 2.24164
R37750 DVSS.n9184 DVSS.n2970 2.24164
R37751 DVSS.n9187 DVSS.n2923 2.24164
R37752 DVSS.n9184 DVSS.n2969 2.24164
R37753 DVSS.n9187 DVSS.n2922 2.24164
R37754 DVSS.n9184 DVSS.n2968 2.24164
R37755 DVSS.n9187 DVSS.n2921 2.24164
R37756 DVSS.n9184 DVSS.n2967 2.24164
R37757 DVSS.n9187 DVSS.n2920 2.24164
R37758 DVSS.n9184 DVSS.n2966 2.24164
R37759 DVSS.n9187 DVSS.n2919 2.24164
R37760 DVSS.n9184 DVSS.n2965 2.24164
R37761 DVSS.n9187 DVSS.n2918 2.24164
R37762 DVSS.n9184 DVSS.n2964 2.24164
R37763 DVSS.n9187 DVSS.n2917 2.24164
R37764 DVSS.n9184 DVSS.n2963 2.24164
R37765 DVSS.n9187 DVSS.n2916 2.24164
R37766 DVSS.n9184 DVSS.n2962 2.24164
R37767 DVSS.n9187 DVSS.n2915 2.24164
R37768 DVSS.n9184 DVSS.n2961 2.24164
R37769 DVSS.n9187 DVSS.n2914 2.24164
R37770 DVSS.n9184 DVSS.n2960 2.24164
R37771 DVSS.n9187 DVSS.n2913 2.24164
R37772 DVSS.n9184 DVSS.n2959 2.24164
R37773 DVSS.n9187 DVSS.n2912 2.24164
R37774 DVSS.n9184 DVSS.n2958 2.24164
R37775 DVSS.n9187 DVSS.n2911 2.24164
R37776 DVSS.n9184 DVSS.n2957 2.24164
R37777 DVSS.n9187 DVSS.n2910 2.24164
R37778 DVSS.n9184 DVSS.n2956 2.24164
R37779 DVSS.n9187 DVSS.n2909 2.24164
R37780 DVSS.n9184 DVSS.n2955 2.24164
R37781 DVSS.n9187 DVSS.n2908 2.24164
R37782 DVSS.n9184 DVSS.n2954 2.24164
R37783 DVSS.n9187 DVSS.n2907 2.24164
R37784 DVSS.n9184 DVSS.n2953 2.24164
R37785 DVSS.n9187 DVSS.n2906 2.24164
R37786 DVSS.n9184 DVSS.n2952 2.24164
R37787 DVSS.n9187 DVSS.n2905 2.24164
R37788 DVSS.n9184 DVSS.n2951 2.24164
R37789 DVSS.n9187 DVSS.n2904 2.24164
R37790 DVSS.n9184 DVSS.n2950 2.24164
R37791 DVSS.n9187 DVSS.n2903 2.24164
R37792 DVSS.n9184 DVSS.n2949 2.24164
R37793 DVSS.n9187 DVSS.n2902 2.24164
R37794 DVSS.n9184 DVSS.n2948 2.24164
R37795 DVSS.n9187 DVSS.n2901 2.24164
R37796 DVSS.n9184 DVSS.n2947 2.24164
R37797 DVSS.n9187 DVSS.n2900 2.24164
R37798 DVSS.n9184 DVSS.n2946 2.24164
R37799 DVSS.n9187 DVSS.n2899 2.24164
R37800 DVSS.n9184 DVSS.n2945 2.24164
R37801 DVSS.n9187 DVSS.n2898 2.24164
R37802 DVSS.n9184 DVSS.n2944 2.24164
R37803 DVSS.n9187 DVSS.n2897 2.24164
R37804 DVSS.n9184 DVSS.n2943 2.24164
R37805 DVSS.n9187 DVSS.n2896 2.24164
R37806 DVSS.n9184 DVSS.n2942 2.24164
R37807 DVSS.n9187 DVSS.n2895 2.24164
R37808 DVSS.n9184 DVSS.n2941 2.24164
R37809 DVSS.n9187 DVSS.n2894 2.24164
R37810 DVSS.n9184 DVSS.n2940 2.24164
R37811 DVSS.n9187 DVSS.n2893 2.24164
R37812 DVSS.n9184 DVSS.n2939 2.24164
R37813 DVSS.n9187 DVSS.n2892 2.24164
R37814 DVSS.n9184 DVSS.n2938 2.24164
R37815 DVSS.n9187 DVSS.n2891 2.24164
R37816 DVSS.n8969 DVSS.n8968 2.24164
R37817 DVSS.n8678 DVSS.n3052 2.24164
R37818 DVSS.n8969 DVSS.n8676 2.24164
R37819 DVSS.n8959 DVSS.n3052 2.24164
R37820 DVSS.n8969 DVSS.n8675 2.24164
R37821 DVSS.n8954 DVSS.n3052 2.24164
R37822 DVSS.n8969 DVSS.n8674 2.24164
R37823 DVSS.n8947 DVSS.n3052 2.24164
R37824 DVSS.n8969 DVSS.n8673 2.24164
R37825 DVSS.n8942 DVSS.n3052 2.24164
R37826 DVSS.n8969 DVSS.n8672 2.24164
R37827 DVSS.n8935 DVSS.n3052 2.24164
R37828 DVSS.n8969 DVSS.n8671 2.24164
R37829 DVSS.n8930 DVSS.n3052 2.24164
R37830 DVSS.n8969 DVSS.n8670 2.24164
R37831 DVSS.n8923 DVSS.n3052 2.24164
R37832 DVSS.n8969 DVSS.n8669 2.24164
R37833 DVSS.n8918 DVSS.n3052 2.24164
R37834 DVSS.n8969 DVSS.n8668 2.24164
R37835 DVSS.n8911 DVSS.n3052 2.24164
R37836 DVSS.n8969 DVSS.n8667 2.24164
R37837 DVSS.n8906 DVSS.n3052 2.24164
R37838 DVSS.n8969 DVSS.n8666 2.24164
R37839 DVSS.n8899 DVSS.n3052 2.24164
R37840 DVSS.n8969 DVSS.n8665 2.24164
R37841 DVSS.n8894 DVSS.n3052 2.24164
R37842 DVSS.n8969 DVSS.n8664 2.24164
R37843 DVSS.n8887 DVSS.n3052 2.24164
R37844 DVSS.n8969 DVSS.n8663 2.24164
R37845 DVSS.n8882 DVSS.n3052 2.24164
R37846 DVSS.n8969 DVSS.n8662 2.24164
R37847 DVSS.n8875 DVSS.n3052 2.24164
R37848 DVSS.n8969 DVSS.n8661 2.24164
R37849 DVSS.n8870 DVSS.n3052 2.24164
R37850 DVSS.n8969 DVSS.n8660 2.24164
R37851 DVSS.n8863 DVSS.n3052 2.24164
R37852 DVSS.n8969 DVSS.n8659 2.24164
R37853 DVSS.n8858 DVSS.n3052 2.24164
R37854 DVSS.n8969 DVSS.n8658 2.24164
R37855 DVSS.n8851 DVSS.n3052 2.24164
R37856 DVSS.n8969 DVSS.n8657 2.24164
R37857 DVSS.n8846 DVSS.n3052 2.24164
R37858 DVSS.n8969 DVSS.n8656 2.24164
R37859 DVSS.n8839 DVSS.n3052 2.24164
R37860 DVSS.n8969 DVSS.n8655 2.24164
R37861 DVSS.n8834 DVSS.n3052 2.24164
R37862 DVSS.n8969 DVSS.n8654 2.24164
R37863 DVSS.n8827 DVSS.n3052 2.24164
R37864 DVSS.n8969 DVSS.n8653 2.24164
R37865 DVSS.n8822 DVSS.n3052 2.24164
R37866 DVSS.n8969 DVSS.n8652 2.24164
R37867 DVSS.n8815 DVSS.n3052 2.24164
R37868 DVSS.n8969 DVSS.n8651 2.24164
R37869 DVSS.n8810 DVSS.n3052 2.24164
R37870 DVSS.n8969 DVSS.n8650 2.24164
R37871 DVSS.n8803 DVSS.n3052 2.24164
R37872 DVSS.n8969 DVSS.n8649 2.24164
R37873 DVSS.n8798 DVSS.n3052 2.24164
R37874 DVSS.n8969 DVSS.n8648 2.24164
R37875 DVSS.n8791 DVSS.n3052 2.24164
R37876 DVSS.n8969 DVSS.n8647 2.24164
R37877 DVSS.n8786 DVSS.n3052 2.24164
R37878 DVSS.n8969 DVSS.n8646 2.24164
R37879 DVSS.n8779 DVSS.n3052 2.24164
R37880 DVSS.n8969 DVSS.n8645 2.24164
R37881 DVSS.n8774 DVSS.n3052 2.24164
R37882 DVSS.n8969 DVSS.n8644 2.24164
R37883 DVSS.n8767 DVSS.n3052 2.24164
R37884 DVSS.n8969 DVSS.n8643 2.24164
R37885 DVSS.n8762 DVSS.n3052 2.24164
R37886 DVSS.n8969 DVSS.n8642 2.24164
R37887 DVSS.n8755 DVSS.n3052 2.24164
R37888 DVSS.n8969 DVSS.n8641 2.24164
R37889 DVSS.n8750 DVSS.n3052 2.24164
R37890 DVSS.n8969 DVSS.n8640 2.24164
R37891 DVSS.n8743 DVSS.n3052 2.24164
R37892 DVSS.n8969 DVSS.n8639 2.24164
R37893 DVSS.n8738 DVSS.n3052 2.24164
R37894 DVSS.n8969 DVSS.n8638 2.24164
R37895 DVSS.n8731 DVSS.n3052 2.24164
R37896 DVSS.n8969 DVSS.n8637 2.24164
R37897 DVSS.n8726 DVSS.n3052 2.24164
R37898 DVSS.n8969 DVSS.n8636 2.24164
R37899 DVSS.n3154 DVSS.n3066 2.24164
R37900 DVSS.n3156 DVSS.n3059 2.24164
R37901 DVSS.n3158 DVSS.n3066 2.24164
R37902 DVSS.n3148 DVSS.n3059 2.24164
R37903 DVSS.n3166 DVSS.n3066 2.24164
R37904 DVSS.n3168 DVSS.n3059 2.24164
R37905 DVSS.n3170 DVSS.n3066 2.24164
R37906 DVSS.n3144 DVSS.n3059 2.24164
R37907 DVSS.n3178 DVSS.n3066 2.24164
R37908 DVSS.n3180 DVSS.n3059 2.24164
R37909 DVSS.n3182 DVSS.n3066 2.24164
R37910 DVSS.n3140 DVSS.n3059 2.24164
R37911 DVSS.n3190 DVSS.n3066 2.24164
R37912 DVSS.n3192 DVSS.n3059 2.24164
R37913 DVSS.n3194 DVSS.n3066 2.24164
R37914 DVSS.n3136 DVSS.n3059 2.24164
R37915 DVSS.n3202 DVSS.n3066 2.24164
R37916 DVSS.n3204 DVSS.n3059 2.24164
R37917 DVSS.n3206 DVSS.n3066 2.24164
R37918 DVSS.n3132 DVSS.n3059 2.24164
R37919 DVSS.n3214 DVSS.n3066 2.24164
R37920 DVSS.n3216 DVSS.n3059 2.24164
R37921 DVSS.n3218 DVSS.n3066 2.24164
R37922 DVSS.n3128 DVSS.n3059 2.24164
R37923 DVSS.n3226 DVSS.n3066 2.24164
R37924 DVSS.n3228 DVSS.n3059 2.24164
R37925 DVSS.n3230 DVSS.n3066 2.24164
R37926 DVSS.n3124 DVSS.n3059 2.24164
R37927 DVSS.n3238 DVSS.n3066 2.24164
R37928 DVSS.n3240 DVSS.n3059 2.24164
R37929 DVSS.n3242 DVSS.n3066 2.24164
R37930 DVSS.n3120 DVSS.n3059 2.24164
R37931 DVSS.n3250 DVSS.n3066 2.24164
R37932 DVSS.n3252 DVSS.n3059 2.24164
R37933 DVSS.n3254 DVSS.n3066 2.24164
R37934 DVSS.n3116 DVSS.n3059 2.24164
R37935 DVSS.n3262 DVSS.n3066 2.24164
R37936 DVSS.n3264 DVSS.n3059 2.24164
R37937 DVSS.n3266 DVSS.n3066 2.24164
R37938 DVSS.n3112 DVSS.n3059 2.24164
R37939 DVSS.n3274 DVSS.n3066 2.24164
R37940 DVSS.n3276 DVSS.n3059 2.24164
R37941 DVSS.n3278 DVSS.n3066 2.24164
R37942 DVSS.n3108 DVSS.n3059 2.24164
R37943 DVSS.n3286 DVSS.n3066 2.24164
R37944 DVSS.n3288 DVSS.n3059 2.24164
R37945 DVSS.n3290 DVSS.n3066 2.24164
R37946 DVSS.n3104 DVSS.n3059 2.24164
R37947 DVSS.n3298 DVSS.n3066 2.24164
R37948 DVSS.n3300 DVSS.n3059 2.24164
R37949 DVSS.n3302 DVSS.n3066 2.24164
R37950 DVSS.n3100 DVSS.n3059 2.24164
R37951 DVSS.n3310 DVSS.n3066 2.24164
R37952 DVSS.n3312 DVSS.n3059 2.24164
R37953 DVSS.n3314 DVSS.n3066 2.24164
R37954 DVSS.n3096 DVSS.n3059 2.24164
R37955 DVSS.n3322 DVSS.n3066 2.24164
R37956 DVSS.n3324 DVSS.n3059 2.24164
R37957 DVSS.n3326 DVSS.n3066 2.24164
R37958 DVSS.n3092 DVSS.n3059 2.24164
R37959 DVSS.n3334 DVSS.n3066 2.24164
R37960 DVSS.n3336 DVSS.n3059 2.24164
R37961 DVSS.n3338 DVSS.n3066 2.24164
R37962 DVSS.n3088 DVSS.n3059 2.24164
R37963 DVSS.n3346 DVSS.n3066 2.24164
R37964 DVSS.n3348 DVSS.n3059 2.24164
R37965 DVSS.n3350 DVSS.n3066 2.24164
R37966 DVSS.n3084 DVSS.n3059 2.24164
R37967 DVSS.n3358 DVSS.n3066 2.24164
R37968 DVSS.n3360 DVSS.n3059 2.24164
R37969 DVSS.n3362 DVSS.n3066 2.24164
R37970 DVSS.n3080 DVSS.n3059 2.24164
R37971 DVSS.n3370 DVSS.n3066 2.24164
R37972 DVSS.n3372 DVSS.n3059 2.24164
R37973 DVSS.n3374 DVSS.n3066 2.24164
R37974 DVSS.n3076 DVSS.n3059 2.24164
R37975 DVSS.n3382 DVSS.n3066 2.24164
R37976 DVSS.n3384 DVSS.n3059 2.24164
R37977 DVSS.n3386 DVSS.n3066 2.24164
R37978 DVSS.n3072 DVSS.n3059 2.24164
R37979 DVSS.n3395 DVSS.n3066 2.24164
R37980 DVSS.n3397 DVSS.n3059 2.24164
R37981 DVSS.n3399 DVSS.n3066 2.24164
R37982 DVSS.n8604 DVSS.n8603 2.24164
R37983 DVSS.n8601 DVSS.n3501 2.24164
R37984 DVSS.n8604 DVSS.n3456 2.24164
R37985 DVSS.n8601 DVSS.n3500 2.24164
R37986 DVSS.n8604 DVSS.n3455 2.24164
R37987 DVSS.n8601 DVSS.n3499 2.24164
R37988 DVSS.n8604 DVSS.n3454 2.24164
R37989 DVSS.n8601 DVSS.n3498 2.24164
R37990 DVSS.n8604 DVSS.n3453 2.24164
R37991 DVSS.n8601 DVSS.n3497 2.24164
R37992 DVSS.n8604 DVSS.n3452 2.24164
R37993 DVSS.n8601 DVSS.n3496 2.24164
R37994 DVSS.n8604 DVSS.n3451 2.24164
R37995 DVSS.n8601 DVSS.n3495 2.24164
R37996 DVSS.n8604 DVSS.n3450 2.24164
R37997 DVSS.n8601 DVSS.n3494 2.24164
R37998 DVSS.n8604 DVSS.n3449 2.24164
R37999 DVSS.n8601 DVSS.n3493 2.24164
R38000 DVSS.n8604 DVSS.n3448 2.24164
R38001 DVSS.n8601 DVSS.n3492 2.24164
R38002 DVSS.n8604 DVSS.n3447 2.24164
R38003 DVSS.n8601 DVSS.n3491 2.24164
R38004 DVSS.n8604 DVSS.n3446 2.24164
R38005 DVSS.n8601 DVSS.n3490 2.24164
R38006 DVSS.n8604 DVSS.n3445 2.24164
R38007 DVSS.n8601 DVSS.n3489 2.24164
R38008 DVSS.n8604 DVSS.n3444 2.24164
R38009 DVSS.n8601 DVSS.n3488 2.24164
R38010 DVSS.n8604 DVSS.n3443 2.24164
R38011 DVSS.n8601 DVSS.n3487 2.24164
R38012 DVSS.n8604 DVSS.n3442 2.24164
R38013 DVSS.n8601 DVSS.n3486 2.24164
R38014 DVSS.n8604 DVSS.n3441 2.24164
R38015 DVSS.n8601 DVSS.n3485 2.24164
R38016 DVSS.n8604 DVSS.n3440 2.24164
R38017 DVSS.n8601 DVSS.n3484 2.24164
R38018 DVSS.n8604 DVSS.n3439 2.24164
R38019 DVSS.n8601 DVSS.n3483 2.24164
R38020 DVSS.n8604 DVSS.n3438 2.24164
R38021 DVSS.n8601 DVSS.n3482 2.24164
R38022 DVSS.n8604 DVSS.n3437 2.24164
R38023 DVSS.n8601 DVSS.n3481 2.24164
R38024 DVSS.n8604 DVSS.n3436 2.24164
R38025 DVSS.n8601 DVSS.n3480 2.24164
R38026 DVSS.n8604 DVSS.n3435 2.24164
R38027 DVSS.n8601 DVSS.n3479 2.24164
R38028 DVSS.n8604 DVSS.n3434 2.24164
R38029 DVSS.n8601 DVSS.n3478 2.24164
R38030 DVSS.n8604 DVSS.n3433 2.24164
R38031 DVSS.n8601 DVSS.n3477 2.24164
R38032 DVSS.n8604 DVSS.n3432 2.24164
R38033 DVSS.n8601 DVSS.n3476 2.24164
R38034 DVSS.n8604 DVSS.n3431 2.24164
R38035 DVSS.n8601 DVSS.n3475 2.24164
R38036 DVSS.n8604 DVSS.n3430 2.24164
R38037 DVSS.n8601 DVSS.n3474 2.24164
R38038 DVSS.n8604 DVSS.n3429 2.24164
R38039 DVSS.n8601 DVSS.n3473 2.24164
R38040 DVSS.n8604 DVSS.n3428 2.24164
R38041 DVSS.n8601 DVSS.n3472 2.24164
R38042 DVSS.n8604 DVSS.n3427 2.24164
R38043 DVSS.n8601 DVSS.n3471 2.24164
R38044 DVSS.n8604 DVSS.n3426 2.24164
R38045 DVSS.n8601 DVSS.n3470 2.24164
R38046 DVSS.n8604 DVSS.n3425 2.24164
R38047 DVSS.n8601 DVSS.n3469 2.24164
R38048 DVSS.n8604 DVSS.n3424 2.24164
R38049 DVSS.n8601 DVSS.n3468 2.24164
R38050 DVSS.n8604 DVSS.n3423 2.24164
R38051 DVSS.n8601 DVSS.n3467 2.24164
R38052 DVSS.n8604 DVSS.n3422 2.24164
R38053 DVSS.n8601 DVSS.n3466 2.24164
R38054 DVSS.n8604 DVSS.n3421 2.24164
R38055 DVSS.n8601 DVSS.n3465 2.24164
R38056 DVSS.n8604 DVSS.n3420 2.24164
R38057 DVSS.n8601 DVSS.n3464 2.24164
R38058 DVSS.n8604 DVSS.n3419 2.24164
R38059 DVSS.n8601 DVSS.n3463 2.24164
R38060 DVSS.n8604 DVSS.n3418 2.24164
R38061 DVSS.n8601 DVSS.n3462 2.24164
R38062 DVSS.n8604 DVSS.n3417 2.24164
R38063 DVSS.n8601 DVSS.n3461 2.24164
R38064 DVSS.n8604 DVSS.n3416 2.24164
R38065 DVSS.n3840 DVSS.n3799 2.24164
R38066 DVSS.n8588 DVSS.n3796 2.24164
R38067 DVSS.n8345 DVSS.n3799 2.24164
R38068 DVSS.n8588 DVSS.n3795 2.24164
R38069 DVSS.n8349 DVSS.n3799 2.24164
R38070 DVSS.n8588 DVSS.n3794 2.24164
R38071 DVSS.n8357 DVSS.n3799 2.24164
R38072 DVSS.n8588 DVSS.n3793 2.24164
R38073 DVSS.n8361 DVSS.n3799 2.24164
R38074 DVSS.n8588 DVSS.n3792 2.24164
R38075 DVSS.n8369 DVSS.n3799 2.24164
R38076 DVSS.n8588 DVSS.n3791 2.24164
R38077 DVSS.n8373 DVSS.n3799 2.24164
R38078 DVSS.n8588 DVSS.n3790 2.24164
R38079 DVSS.n8381 DVSS.n3799 2.24164
R38080 DVSS.n8588 DVSS.n3789 2.24164
R38081 DVSS.n8385 DVSS.n3799 2.24164
R38082 DVSS.n8588 DVSS.n3788 2.24164
R38083 DVSS.n8393 DVSS.n3799 2.24164
R38084 DVSS.n8588 DVSS.n3787 2.24164
R38085 DVSS.n8397 DVSS.n3799 2.24164
R38086 DVSS.n8588 DVSS.n3786 2.24164
R38087 DVSS.n8405 DVSS.n3799 2.24164
R38088 DVSS.n8588 DVSS.n3785 2.24164
R38089 DVSS.n8409 DVSS.n3799 2.24164
R38090 DVSS.n8588 DVSS.n3784 2.24164
R38091 DVSS.n8417 DVSS.n3799 2.24164
R38092 DVSS.n8588 DVSS.n3783 2.24164
R38093 DVSS.n8421 DVSS.n3799 2.24164
R38094 DVSS.n8588 DVSS.n3782 2.24164
R38095 DVSS.n8429 DVSS.n3799 2.24164
R38096 DVSS.n8588 DVSS.n3781 2.24164
R38097 DVSS.n8433 DVSS.n3799 2.24164
R38098 DVSS.n8588 DVSS.n3780 2.24164
R38099 DVSS.n8441 DVSS.n3799 2.24164
R38100 DVSS.n8588 DVSS.n3779 2.24164
R38101 DVSS.n8445 DVSS.n3799 2.24164
R38102 DVSS.n8588 DVSS.n3778 2.24164
R38103 DVSS.n8453 DVSS.n3799 2.24164
R38104 DVSS.n8588 DVSS.n3777 2.24164
R38105 DVSS.n8457 DVSS.n3799 2.24164
R38106 DVSS.n8588 DVSS.n3776 2.24164
R38107 DVSS.n8465 DVSS.n3799 2.24164
R38108 DVSS.n8588 DVSS.n3775 2.24164
R38109 DVSS.n8469 DVSS.n3799 2.24164
R38110 DVSS.n8588 DVSS.n3774 2.24164
R38111 DVSS.n8477 DVSS.n3799 2.24164
R38112 DVSS.n8588 DVSS.n3773 2.24164
R38113 DVSS.n8481 DVSS.n3799 2.24164
R38114 DVSS.n8588 DVSS.n3772 2.24164
R38115 DVSS.n8489 DVSS.n3799 2.24164
R38116 DVSS.n8588 DVSS.n3771 2.24164
R38117 DVSS.n8493 DVSS.n3799 2.24164
R38118 DVSS.n8588 DVSS.n3770 2.24164
R38119 DVSS.n8501 DVSS.n3799 2.24164
R38120 DVSS.n8588 DVSS.n3769 2.24164
R38121 DVSS.n8505 DVSS.n3799 2.24164
R38122 DVSS.n8588 DVSS.n3768 2.24164
R38123 DVSS.n8513 DVSS.n3799 2.24164
R38124 DVSS.n8588 DVSS.n3767 2.24164
R38125 DVSS.n8517 DVSS.n3799 2.24164
R38126 DVSS.n8588 DVSS.n3766 2.24164
R38127 DVSS.n8525 DVSS.n3799 2.24164
R38128 DVSS.n8588 DVSS.n3765 2.24164
R38129 DVSS.n8529 DVSS.n3799 2.24164
R38130 DVSS.n8588 DVSS.n3764 2.24164
R38131 DVSS.n8537 DVSS.n3799 2.24164
R38132 DVSS.n8588 DVSS.n3763 2.24164
R38133 DVSS.n8541 DVSS.n3799 2.24164
R38134 DVSS.n8588 DVSS.n3762 2.24164
R38135 DVSS.n8549 DVSS.n3799 2.24164
R38136 DVSS.n8588 DVSS.n3761 2.24164
R38137 DVSS.n8553 DVSS.n3799 2.24164
R38138 DVSS.n8588 DVSS.n3760 2.24164
R38139 DVSS.n8561 DVSS.n3799 2.24164
R38140 DVSS.n8588 DVSS.n3759 2.24164
R38141 DVSS.n8565 DVSS.n3799 2.24164
R38142 DVSS.n8588 DVSS.n3758 2.24164
R38143 DVSS.n8573 DVSS.n3799 2.24164
R38144 DVSS.n8588 DVSS.n3757 2.24164
R38145 DVSS.n8577 DVSS.n3799 2.24164
R38146 DVSS.n8588 DVSS.n3756 2.24164
R38147 DVSS.n8586 DVSS.n3799 2.24164
R38148 DVSS.n8320 DVSS.n8319 2.24164
R38149 DVSS.n8317 DVSS.n3945 2.24164
R38150 DVSS.n8320 DVSS.n3899 2.24164
R38151 DVSS.n8317 DVSS.n3944 2.24164
R38152 DVSS.n8320 DVSS.n3898 2.24164
R38153 DVSS.n8317 DVSS.n3943 2.24164
R38154 DVSS.n8320 DVSS.n3897 2.24164
R38155 DVSS.n8317 DVSS.n3942 2.24164
R38156 DVSS.n8320 DVSS.n3896 2.24164
R38157 DVSS.n8317 DVSS.n3941 2.24164
R38158 DVSS.n8320 DVSS.n3895 2.24164
R38159 DVSS.n8317 DVSS.n3940 2.24164
R38160 DVSS.n8320 DVSS.n3894 2.24164
R38161 DVSS.n8317 DVSS.n3939 2.24164
R38162 DVSS.n8320 DVSS.n3893 2.24164
R38163 DVSS.n8317 DVSS.n3938 2.24164
R38164 DVSS.n8320 DVSS.n3892 2.24164
R38165 DVSS.n8317 DVSS.n3937 2.24164
R38166 DVSS.n8320 DVSS.n3891 2.24164
R38167 DVSS.n8317 DVSS.n3936 2.24164
R38168 DVSS.n8320 DVSS.n3890 2.24164
R38169 DVSS.n8317 DVSS.n3935 2.24164
R38170 DVSS.n8320 DVSS.n3889 2.24164
R38171 DVSS.n8317 DVSS.n3934 2.24164
R38172 DVSS.n8320 DVSS.n3888 2.24164
R38173 DVSS.n8317 DVSS.n3933 2.24164
R38174 DVSS.n8320 DVSS.n3887 2.24164
R38175 DVSS.n8317 DVSS.n3932 2.24164
R38176 DVSS.n8320 DVSS.n3886 2.24164
R38177 DVSS.n8317 DVSS.n3931 2.24164
R38178 DVSS.n8320 DVSS.n3885 2.24164
R38179 DVSS.n8317 DVSS.n3930 2.24164
R38180 DVSS.n8320 DVSS.n3884 2.24164
R38181 DVSS.n8317 DVSS.n3929 2.24164
R38182 DVSS.n8320 DVSS.n3883 2.24164
R38183 DVSS.n8317 DVSS.n3928 2.24164
R38184 DVSS.n8320 DVSS.n3882 2.24164
R38185 DVSS.n8317 DVSS.n3927 2.24164
R38186 DVSS.n8320 DVSS.n3881 2.24164
R38187 DVSS.n8317 DVSS.n3926 2.24164
R38188 DVSS.n8320 DVSS.n3880 2.24164
R38189 DVSS.n8317 DVSS.n3925 2.24164
R38190 DVSS.n8320 DVSS.n3879 2.24164
R38191 DVSS.n8317 DVSS.n3924 2.24164
R38192 DVSS.n8320 DVSS.n3878 2.24164
R38193 DVSS.n8317 DVSS.n3923 2.24164
R38194 DVSS.n8320 DVSS.n3877 2.24164
R38195 DVSS.n8317 DVSS.n3922 2.24164
R38196 DVSS.n8320 DVSS.n3876 2.24164
R38197 DVSS.n8317 DVSS.n3921 2.24164
R38198 DVSS.n8320 DVSS.n3875 2.24164
R38199 DVSS.n8317 DVSS.n3920 2.24164
R38200 DVSS.n8320 DVSS.n3874 2.24164
R38201 DVSS.n8317 DVSS.n3919 2.24164
R38202 DVSS.n8320 DVSS.n3873 2.24164
R38203 DVSS.n8317 DVSS.n3918 2.24164
R38204 DVSS.n8320 DVSS.n3872 2.24164
R38205 DVSS.n8317 DVSS.n3917 2.24164
R38206 DVSS.n8320 DVSS.n3871 2.24164
R38207 DVSS.n8317 DVSS.n3916 2.24164
R38208 DVSS.n8320 DVSS.n3870 2.24164
R38209 DVSS.n8317 DVSS.n3915 2.24164
R38210 DVSS.n8320 DVSS.n3869 2.24164
R38211 DVSS.n8317 DVSS.n3914 2.24164
R38212 DVSS.n8320 DVSS.n3868 2.24164
R38213 DVSS.n8317 DVSS.n3913 2.24164
R38214 DVSS.n8320 DVSS.n3867 2.24164
R38215 DVSS.n8317 DVSS.n3912 2.24164
R38216 DVSS.n8320 DVSS.n3866 2.24164
R38217 DVSS.n8317 DVSS.n3911 2.24164
R38218 DVSS.n8320 DVSS.n3865 2.24164
R38219 DVSS.n8317 DVSS.n3910 2.24164
R38220 DVSS.n8320 DVSS.n3864 2.24164
R38221 DVSS.n8317 DVSS.n3909 2.24164
R38222 DVSS.n8320 DVSS.n3863 2.24164
R38223 DVSS.n8317 DVSS.n3908 2.24164
R38224 DVSS.n8320 DVSS.n3862 2.24164
R38225 DVSS.n8317 DVSS.n3907 2.24164
R38226 DVSS.n8320 DVSS.n3861 2.24164
R38227 DVSS.n8317 DVSS.n3906 2.24164
R38228 DVSS.n8320 DVSS.n3860 2.24164
R38229 DVSS.n8317 DVSS.n3905 2.24164
R38230 DVSS.n8320 DVSS.n3859 2.24164
R38231 DVSS.n4110 DVSS.n4021 2.24164
R38232 DVSS.n4112 DVSS.n4022 2.24164
R38233 DVSS.n4114 DVSS.n4021 2.24164
R38234 DVSS.n4104 DVSS.n4022 2.24164
R38235 DVSS.n4122 DVSS.n4021 2.24164
R38236 DVSS.n4124 DVSS.n4022 2.24164
R38237 DVSS.n4126 DVSS.n4021 2.24164
R38238 DVSS.n4100 DVSS.n4022 2.24164
R38239 DVSS.n4134 DVSS.n4021 2.24164
R38240 DVSS.n4136 DVSS.n4022 2.24164
R38241 DVSS.n4138 DVSS.n4021 2.24164
R38242 DVSS.n4096 DVSS.n4022 2.24164
R38243 DVSS.n4146 DVSS.n4021 2.24164
R38244 DVSS.n4148 DVSS.n4022 2.24164
R38245 DVSS.n4150 DVSS.n4021 2.24164
R38246 DVSS.n4092 DVSS.n4022 2.24164
R38247 DVSS.n4158 DVSS.n4021 2.24164
R38248 DVSS.n4160 DVSS.n4022 2.24164
R38249 DVSS.n4162 DVSS.n4021 2.24164
R38250 DVSS.n4088 DVSS.n4022 2.24164
R38251 DVSS.n4170 DVSS.n4021 2.24164
R38252 DVSS.n4172 DVSS.n4022 2.24164
R38253 DVSS.n4174 DVSS.n4021 2.24164
R38254 DVSS.n4084 DVSS.n4022 2.24164
R38255 DVSS.n4182 DVSS.n4021 2.24164
R38256 DVSS.n4184 DVSS.n4022 2.24164
R38257 DVSS.n4186 DVSS.n4021 2.24164
R38258 DVSS.n4080 DVSS.n4022 2.24164
R38259 DVSS.n4194 DVSS.n4021 2.24164
R38260 DVSS.n4196 DVSS.n4022 2.24164
R38261 DVSS.n4198 DVSS.n4021 2.24164
R38262 DVSS.n4076 DVSS.n4022 2.24164
R38263 DVSS.n4206 DVSS.n4021 2.24164
R38264 DVSS.n4208 DVSS.n4022 2.24164
R38265 DVSS.n4210 DVSS.n4021 2.24164
R38266 DVSS.n4072 DVSS.n4022 2.24164
R38267 DVSS.n4218 DVSS.n4021 2.24164
R38268 DVSS.n4220 DVSS.n4022 2.24164
R38269 DVSS.n4222 DVSS.n4021 2.24164
R38270 DVSS.n4068 DVSS.n4022 2.24164
R38271 DVSS.n4230 DVSS.n4021 2.24164
R38272 DVSS.n4232 DVSS.n4022 2.24164
R38273 DVSS.n4234 DVSS.n4021 2.24164
R38274 DVSS.n4064 DVSS.n4022 2.24164
R38275 DVSS.n4242 DVSS.n4021 2.24164
R38276 DVSS.n4244 DVSS.n4022 2.24164
R38277 DVSS.n4246 DVSS.n4021 2.24164
R38278 DVSS.n4060 DVSS.n4022 2.24164
R38279 DVSS.n4254 DVSS.n4021 2.24164
R38280 DVSS.n4256 DVSS.n4022 2.24164
R38281 DVSS.n4258 DVSS.n4021 2.24164
R38282 DVSS.n4056 DVSS.n4022 2.24164
R38283 DVSS.n4266 DVSS.n4021 2.24164
R38284 DVSS.n4268 DVSS.n4022 2.24164
R38285 DVSS.n4270 DVSS.n4021 2.24164
R38286 DVSS.n4052 DVSS.n4022 2.24164
R38287 DVSS.n4278 DVSS.n4021 2.24164
R38288 DVSS.n4280 DVSS.n4022 2.24164
R38289 DVSS.n4282 DVSS.n4021 2.24164
R38290 DVSS.n4048 DVSS.n4022 2.24164
R38291 DVSS.n4290 DVSS.n4021 2.24164
R38292 DVSS.n4292 DVSS.n4022 2.24164
R38293 DVSS.n4294 DVSS.n4021 2.24164
R38294 DVSS.n4044 DVSS.n4022 2.24164
R38295 DVSS.n4302 DVSS.n4021 2.24164
R38296 DVSS.n4304 DVSS.n4022 2.24164
R38297 DVSS.n4306 DVSS.n4021 2.24164
R38298 DVSS.n4040 DVSS.n4022 2.24164
R38299 DVSS.n4314 DVSS.n4021 2.24164
R38300 DVSS.n4316 DVSS.n4022 2.24164
R38301 DVSS.n4318 DVSS.n4021 2.24164
R38302 DVSS.n4036 DVSS.n4022 2.24164
R38303 DVSS.n4326 DVSS.n4021 2.24164
R38304 DVSS.n4328 DVSS.n4022 2.24164
R38305 DVSS.n4330 DVSS.n4021 2.24164
R38306 DVSS.n4032 DVSS.n4022 2.24164
R38307 DVSS.n4338 DVSS.n4021 2.24164
R38308 DVSS.n4340 DVSS.n4022 2.24164
R38309 DVSS.n4342 DVSS.n4021 2.24164
R38310 DVSS.n4028 DVSS.n4022 2.24164
R38311 DVSS.n4351 DVSS.n4021 2.24164
R38312 DVSS.n4353 DVSS.n4022 2.24164
R38313 DVSS.n4355 DVSS.n4021 2.24164
R38314 DVSS.n8090 DVSS.n8089 2.24164
R38315 DVSS.n4415 DVSS.n4362 2.24164
R38316 DVSS.n8090 DVSS.n4412 2.24164
R38317 DVSS.n8080 DVSS.n4362 2.24164
R38318 DVSS.n8090 DVSS.n4411 2.24164
R38319 DVSS.n8075 DVSS.n4362 2.24164
R38320 DVSS.n8090 DVSS.n4410 2.24164
R38321 DVSS.n8068 DVSS.n4362 2.24164
R38322 DVSS.n8090 DVSS.n4409 2.24164
R38323 DVSS.n8063 DVSS.n4362 2.24164
R38324 DVSS.n8090 DVSS.n4408 2.24164
R38325 DVSS.n8056 DVSS.n4362 2.24164
R38326 DVSS.n8090 DVSS.n4407 2.24164
R38327 DVSS.n8051 DVSS.n4362 2.24164
R38328 DVSS.n8090 DVSS.n4406 2.24164
R38329 DVSS.n8044 DVSS.n4362 2.24164
R38330 DVSS.n8090 DVSS.n4405 2.24164
R38331 DVSS.n8039 DVSS.n4362 2.24164
R38332 DVSS.n8090 DVSS.n4404 2.24164
R38333 DVSS.n8032 DVSS.n4362 2.24164
R38334 DVSS.n8090 DVSS.n4403 2.24164
R38335 DVSS.n8027 DVSS.n4362 2.24164
R38336 DVSS.n8090 DVSS.n4402 2.24164
R38337 DVSS.n8020 DVSS.n4362 2.24164
R38338 DVSS.n8090 DVSS.n4401 2.24164
R38339 DVSS.n8015 DVSS.n4362 2.24164
R38340 DVSS.n8090 DVSS.n4400 2.24164
R38341 DVSS.n8008 DVSS.n4362 2.24164
R38342 DVSS.n8090 DVSS.n4399 2.24164
R38343 DVSS.n8003 DVSS.n4362 2.24164
R38344 DVSS.n8090 DVSS.n4398 2.24164
R38345 DVSS.n7996 DVSS.n4362 2.24164
R38346 DVSS.n8090 DVSS.n4397 2.24164
R38347 DVSS.n7991 DVSS.n4362 2.24164
R38348 DVSS.n8090 DVSS.n4396 2.24164
R38349 DVSS.n7984 DVSS.n4362 2.24164
R38350 DVSS.n8090 DVSS.n4395 2.24164
R38351 DVSS.n7979 DVSS.n4362 2.24164
R38352 DVSS.n8090 DVSS.n4394 2.24164
R38353 DVSS.n7972 DVSS.n4362 2.24164
R38354 DVSS.n8090 DVSS.n4393 2.24164
R38355 DVSS.n7967 DVSS.n4362 2.24164
R38356 DVSS.n8090 DVSS.n4392 2.24164
R38357 DVSS.n7960 DVSS.n4362 2.24164
R38358 DVSS.n8090 DVSS.n4391 2.24164
R38359 DVSS.n7955 DVSS.n4362 2.24164
R38360 DVSS.n8090 DVSS.n4390 2.24164
R38361 DVSS.n7948 DVSS.n4362 2.24164
R38362 DVSS.n8090 DVSS.n4389 2.24164
R38363 DVSS.n7943 DVSS.n4362 2.24164
R38364 DVSS.n8090 DVSS.n4388 2.24164
R38365 DVSS.n7936 DVSS.n4362 2.24164
R38366 DVSS.n8090 DVSS.n4387 2.24164
R38367 DVSS.n7931 DVSS.n4362 2.24164
R38368 DVSS.n8090 DVSS.n4386 2.24164
R38369 DVSS.n7924 DVSS.n4362 2.24164
R38370 DVSS.n8090 DVSS.n4385 2.24164
R38371 DVSS.n7919 DVSS.n4362 2.24164
R38372 DVSS.n8090 DVSS.n4384 2.24164
R38373 DVSS.n7912 DVSS.n4362 2.24164
R38374 DVSS.n8090 DVSS.n4383 2.24164
R38375 DVSS.n7907 DVSS.n4362 2.24164
R38376 DVSS.n8090 DVSS.n4382 2.24164
R38377 DVSS.n7900 DVSS.n4362 2.24164
R38378 DVSS.n8090 DVSS.n4381 2.24164
R38379 DVSS.n7895 DVSS.n4362 2.24164
R38380 DVSS.n8090 DVSS.n4380 2.24164
R38381 DVSS.n7888 DVSS.n4362 2.24164
R38382 DVSS.n8090 DVSS.n4379 2.24164
R38383 DVSS.n7883 DVSS.n4362 2.24164
R38384 DVSS.n8090 DVSS.n4378 2.24164
R38385 DVSS.n7876 DVSS.n4362 2.24164
R38386 DVSS.n8090 DVSS.n4377 2.24164
R38387 DVSS.n7871 DVSS.n4362 2.24164
R38388 DVSS.n8090 DVSS.n4376 2.24164
R38389 DVSS.n7864 DVSS.n4362 2.24164
R38390 DVSS.n8090 DVSS.n4375 2.24164
R38391 DVSS.n7859 DVSS.n4362 2.24164
R38392 DVSS.n8090 DVSS.n4374 2.24164
R38393 DVSS.n7852 DVSS.n4362 2.24164
R38394 DVSS.n8090 DVSS.n4373 2.24164
R38395 DVSS.n7847 DVSS.n4362 2.24164
R38396 DVSS.n8090 DVSS.n4372 2.24164
R38397 DVSS.n4804 DVSS.n4468 2.24164
R38398 DVSS.n4802 DVSS.n4471 2.24164
R38399 DVSS.n4476 DVSS.n4468 2.24164
R38400 DVSS.n4481 DVSS.n4471 2.24164
R38401 DVSS.n4794 DVSS.n4468 2.24164
R38402 DVSS.n4792 DVSS.n4471 2.24164
R38403 DVSS.n4482 DVSS.n4468 2.24164
R38404 DVSS.n4487 DVSS.n4471 2.24164
R38405 DVSS.n4784 DVSS.n4468 2.24164
R38406 DVSS.n4782 DVSS.n4471 2.24164
R38407 DVSS.n4488 DVSS.n4468 2.24164
R38408 DVSS.n4493 DVSS.n4471 2.24164
R38409 DVSS.n4774 DVSS.n4468 2.24164
R38410 DVSS.n4772 DVSS.n4471 2.24164
R38411 DVSS.n4494 DVSS.n4468 2.24164
R38412 DVSS.n4499 DVSS.n4471 2.24164
R38413 DVSS.n4764 DVSS.n4468 2.24164
R38414 DVSS.n4762 DVSS.n4471 2.24164
R38415 DVSS.n4500 DVSS.n4468 2.24164
R38416 DVSS.n4505 DVSS.n4471 2.24164
R38417 DVSS.n4754 DVSS.n4468 2.24164
R38418 DVSS.n4752 DVSS.n4471 2.24164
R38419 DVSS.n4506 DVSS.n4468 2.24164
R38420 DVSS.n4511 DVSS.n4471 2.24164
R38421 DVSS.n4744 DVSS.n4468 2.24164
R38422 DVSS.n4742 DVSS.n4471 2.24164
R38423 DVSS.n4512 DVSS.n4468 2.24164
R38424 DVSS.n4517 DVSS.n4471 2.24164
R38425 DVSS.n4734 DVSS.n4468 2.24164
R38426 DVSS.n4732 DVSS.n4471 2.24164
R38427 DVSS.n4518 DVSS.n4468 2.24164
R38428 DVSS.n4523 DVSS.n4471 2.24164
R38429 DVSS.n4724 DVSS.n4468 2.24164
R38430 DVSS.n4722 DVSS.n4471 2.24164
R38431 DVSS.n4524 DVSS.n4468 2.24164
R38432 DVSS.n4529 DVSS.n4471 2.24164
R38433 DVSS.n4714 DVSS.n4468 2.24164
R38434 DVSS.n4712 DVSS.n4471 2.24164
R38435 DVSS.n4530 DVSS.n4468 2.24164
R38436 DVSS.n4535 DVSS.n4471 2.24164
R38437 DVSS.n4704 DVSS.n4468 2.24164
R38438 DVSS.n4702 DVSS.n4471 2.24164
R38439 DVSS.n4536 DVSS.n4468 2.24164
R38440 DVSS.n4541 DVSS.n4471 2.24164
R38441 DVSS.n4694 DVSS.n4468 2.24164
R38442 DVSS.n4692 DVSS.n4471 2.24164
R38443 DVSS.n4542 DVSS.n4468 2.24164
R38444 DVSS.n4547 DVSS.n4471 2.24164
R38445 DVSS.n4684 DVSS.n4468 2.24164
R38446 DVSS.n4682 DVSS.n4471 2.24164
R38447 DVSS.n4548 DVSS.n4468 2.24164
R38448 DVSS.n4553 DVSS.n4471 2.24164
R38449 DVSS.n4674 DVSS.n4468 2.24164
R38450 DVSS.n4672 DVSS.n4471 2.24164
R38451 DVSS.n4554 DVSS.n4468 2.24164
R38452 DVSS.n4559 DVSS.n4471 2.24164
R38453 DVSS.n4664 DVSS.n4468 2.24164
R38454 DVSS.n4662 DVSS.n4471 2.24164
R38455 DVSS.n4560 DVSS.n4468 2.24164
R38456 DVSS.n4565 DVSS.n4471 2.24164
R38457 DVSS.n4654 DVSS.n4468 2.24164
R38458 DVSS.n4652 DVSS.n4471 2.24164
R38459 DVSS.n4566 DVSS.n4468 2.24164
R38460 DVSS.n4571 DVSS.n4471 2.24164
R38461 DVSS.n4644 DVSS.n4468 2.24164
R38462 DVSS.n4642 DVSS.n4471 2.24164
R38463 DVSS.n4572 DVSS.n4468 2.24164
R38464 DVSS.n4577 DVSS.n4471 2.24164
R38465 DVSS.n4634 DVSS.n4468 2.24164
R38466 DVSS.n4632 DVSS.n4471 2.24164
R38467 DVSS.n4578 DVSS.n4468 2.24164
R38468 DVSS.n4583 DVSS.n4471 2.24164
R38469 DVSS.n4624 DVSS.n4468 2.24164
R38470 DVSS.n4622 DVSS.n4471 2.24164
R38471 DVSS.n4584 DVSS.n4468 2.24164
R38472 DVSS.n4589 DVSS.n4471 2.24164
R38473 DVSS.n4614 DVSS.n4468 2.24164
R38474 DVSS.n4612 DVSS.n4471 2.24164
R38475 DVSS.n4590 DVSS.n4468 2.24164
R38476 DVSS.n4595 DVSS.n4471 2.24164
R38477 DVSS.n4604 DVSS.n4468 2.24164
R38478 DVSS.n4602 DVSS.n4471 2.24164
R38479 DVSS.n4596 DVSS.n4468 2.24164
R38480 DVSS.n7795 DVSS.n7794 2.24164
R38481 DVSS.n7504 DVSS.n4811 2.24164
R38482 DVSS.n7795 DVSS.n7502 2.24164
R38483 DVSS.n7785 DVSS.n4811 2.24164
R38484 DVSS.n7795 DVSS.n7501 2.24164
R38485 DVSS.n7780 DVSS.n4811 2.24164
R38486 DVSS.n7795 DVSS.n7500 2.24164
R38487 DVSS.n7773 DVSS.n4811 2.24164
R38488 DVSS.n7795 DVSS.n7499 2.24164
R38489 DVSS.n7768 DVSS.n4811 2.24164
R38490 DVSS.n7795 DVSS.n7498 2.24164
R38491 DVSS.n7761 DVSS.n4811 2.24164
R38492 DVSS.n7795 DVSS.n7497 2.24164
R38493 DVSS.n7756 DVSS.n4811 2.24164
R38494 DVSS.n7795 DVSS.n7496 2.24164
R38495 DVSS.n7749 DVSS.n4811 2.24164
R38496 DVSS.n7795 DVSS.n7495 2.24164
R38497 DVSS.n7744 DVSS.n4811 2.24164
R38498 DVSS.n7795 DVSS.n7494 2.24164
R38499 DVSS.n7737 DVSS.n4811 2.24164
R38500 DVSS.n7795 DVSS.n7493 2.24164
R38501 DVSS.n7732 DVSS.n4811 2.24164
R38502 DVSS.n7795 DVSS.n7492 2.24164
R38503 DVSS.n7725 DVSS.n4811 2.24164
R38504 DVSS.n7795 DVSS.n7491 2.24164
R38505 DVSS.n7720 DVSS.n4811 2.24164
R38506 DVSS.n7795 DVSS.n7490 2.24164
R38507 DVSS.n7713 DVSS.n4811 2.24164
R38508 DVSS.n7795 DVSS.n7489 2.24164
R38509 DVSS.n7708 DVSS.n4811 2.24164
R38510 DVSS.n7795 DVSS.n7488 2.24164
R38511 DVSS.n7701 DVSS.n4811 2.24164
R38512 DVSS.n7795 DVSS.n7487 2.24164
R38513 DVSS.n7696 DVSS.n4811 2.24164
R38514 DVSS.n7795 DVSS.n7486 2.24164
R38515 DVSS.n7689 DVSS.n4811 2.24164
R38516 DVSS.n7795 DVSS.n7485 2.24164
R38517 DVSS.n7684 DVSS.n4811 2.24164
R38518 DVSS.n7795 DVSS.n7484 2.24164
R38519 DVSS.n7677 DVSS.n4811 2.24164
R38520 DVSS.n7795 DVSS.n7483 2.24164
R38521 DVSS.n7672 DVSS.n4811 2.24164
R38522 DVSS.n7795 DVSS.n7482 2.24164
R38523 DVSS.n7665 DVSS.n4811 2.24164
R38524 DVSS.n7795 DVSS.n7481 2.24164
R38525 DVSS.n7660 DVSS.n4811 2.24164
R38526 DVSS.n7795 DVSS.n7480 2.24164
R38527 DVSS.n7653 DVSS.n4811 2.24164
R38528 DVSS.n7795 DVSS.n7479 2.24164
R38529 DVSS.n7648 DVSS.n4811 2.24164
R38530 DVSS.n7795 DVSS.n7478 2.24164
R38531 DVSS.n7641 DVSS.n4811 2.24164
R38532 DVSS.n7795 DVSS.n7477 2.24164
R38533 DVSS.n7636 DVSS.n4811 2.24164
R38534 DVSS.n7795 DVSS.n7476 2.24164
R38535 DVSS.n7629 DVSS.n4811 2.24164
R38536 DVSS.n7795 DVSS.n7475 2.24164
R38537 DVSS.n7624 DVSS.n4811 2.24164
R38538 DVSS.n7795 DVSS.n7474 2.24164
R38539 DVSS.n7617 DVSS.n4811 2.24164
R38540 DVSS.n7795 DVSS.n7473 2.24164
R38541 DVSS.n7612 DVSS.n4811 2.24164
R38542 DVSS.n7795 DVSS.n7472 2.24164
R38543 DVSS.n7605 DVSS.n4811 2.24164
R38544 DVSS.n7795 DVSS.n7471 2.24164
R38545 DVSS.n7600 DVSS.n4811 2.24164
R38546 DVSS.n7795 DVSS.n7470 2.24164
R38547 DVSS.n7593 DVSS.n4811 2.24164
R38548 DVSS.n7795 DVSS.n7469 2.24164
R38549 DVSS.n7588 DVSS.n4811 2.24164
R38550 DVSS.n7795 DVSS.n7468 2.24164
R38551 DVSS.n7581 DVSS.n4811 2.24164
R38552 DVSS.n7795 DVSS.n7467 2.24164
R38553 DVSS.n7576 DVSS.n4811 2.24164
R38554 DVSS.n7795 DVSS.n7466 2.24164
R38555 DVSS.n7569 DVSS.n4811 2.24164
R38556 DVSS.n7795 DVSS.n7465 2.24164
R38557 DVSS.n7564 DVSS.n4811 2.24164
R38558 DVSS.n7795 DVSS.n7464 2.24164
R38559 DVSS.n7557 DVSS.n4811 2.24164
R38560 DVSS.n7795 DVSS.n7463 2.24164
R38561 DVSS.n7552 DVSS.n4811 2.24164
R38562 DVSS.n7795 DVSS.n7462 2.24164
R38563 DVSS.n7441 DVSS.n4832 2.24164
R38564 DVSS.n7439 DVSS.n4825 2.24164
R38565 DVSS.n7113 DVSS.n4832 2.24164
R38566 DVSS.n7118 DVSS.n4825 2.24164
R38567 DVSS.n7431 DVSS.n4832 2.24164
R38568 DVSS.n7429 DVSS.n4825 2.24164
R38569 DVSS.n7119 DVSS.n4832 2.24164
R38570 DVSS.n7124 DVSS.n4825 2.24164
R38571 DVSS.n7421 DVSS.n4832 2.24164
R38572 DVSS.n7419 DVSS.n4825 2.24164
R38573 DVSS.n7125 DVSS.n4832 2.24164
R38574 DVSS.n7130 DVSS.n4825 2.24164
R38575 DVSS.n7411 DVSS.n4832 2.24164
R38576 DVSS.n7409 DVSS.n4825 2.24164
R38577 DVSS.n7131 DVSS.n4832 2.24164
R38578 DVSS.n7136 DVSS.n4825 2.24164
R38579 DVSS.n7401 DVSS.n4832 2.24164
R38580 DVSS.n7399 DVSS.n4825 2.24164
R38581 DVSS.n7137 DVSS.n4832 2.24164
R38582 DVSS.n7142 DVSS.n4825 2.24164
R38583 DVSS.n7391 DVSS.n4832 2.24164
R38584 DVSS.n7389 DVSS.n4825 2.24164
R38585 DVSS.n7143 DVSS.n4832 2.24164
R38586 DVSS.n7148 DVSS.n4825 2.24164
R38587 DVSS.n7381 DVSS.n4832 2.24164
R38588 DVSS.n7379 DVSS.n4825 2.24164
R38589 DVSS.n7149 DVSS.n4832 2.24164
R38590 DVSS.n7154 DVSS.n4825 2.24164
R38591 DVSS.n7371 DVSS.n4832 2.24164
R38592 DVSS.n7369 DVSS.n4825 2.24164
R38593 DVSS.n7155 DVSS.n4832 2.24164
R38594 DVSS.n7160 DVSS.n4825 2.24164
R38595 DVSS.n7361 DVSS.n4832 2.24164
R38596 DVSS.n7359 DVSS.n4825 2.24164
R38597 DVSS.n7161 DVSS.n4832 2.24164
R38598 DVSS.n7166 DVSS.n4825 2.24164
R38599 DVSS.n7351 DVSS.n4832 2.24164
R38600 DVSS.n7349 DVSS.n4825 2.24164
R38601 DVSS.n7167 DVSS.n4832 2.24164
R38602 DVSS.n7172 DVSS.n4825 2.24164
R38603 DVSS.n7341 DVSS.n4832 2.24164
R38604 DVSS.n7339 DVSS.n4825 2.24164
R38605 DVSS.n7173 DVSS.n4832 2.24164
R38606 DVSS.n7178 DVSS.n4825 2.24164
R38607 DVSS.n7331 DVSS.n4832 2.24164
R38608 DVSS.n7329 DVSS.n4825 2.24164
R38609 DVSS.n7179 DVSS.n4832 2.24164
R38610 DVSS.n7184 DVSS.n4825 2.24164
R38611 DVSS.n7321 DVSS.n4832 2.24164
R38612 DVSS.n7319 DVSS.n4825 2.24164
R38613 DVSS.n7185 DVSS.n4832 2.24164
R38614 DVSS.n7190 DVSS.n4825 2.24164
R38615 DVSS.n7311 DVSS.n4832 2.24164
R38616 DVSS.n7309 DVSS.n4825 2.24164
R38617 DVSS.n7191 DVSS.n4832 2.24164
R38618 DVSS.n7196 DVSS.n4825 2.24164
R38619 DVSS.n7301 DVSS.n4832 2.24164
R38620 DVSS.n7299 DVSS.n4825 2.24164
R38621 DVSS.n7197 DVSS.n4832 2.24164
R38622 DVSS.n7202 DVSS.n4825 2.24164
R38623 DVSS.n7291 DVSS.n4832 2.24164
R38624 DVSS.n7289 DVSS.n4825 2.24164
R38625 DVSS.n7203 DVSS.n4832 2.24164
R38626 DVSS.n7208 DVSS.n4825 2.24164
R38627 DVSS.n7281 DVSS.n4832 2.24164
R38628 DVSS.n7279 DVSS.n4825 2.24164
R38629 DVSS.n7209 DVSS.n4832 2.24164
R38630 DVSS.n7214 DVSS.n4825 2.24164
R38631 DVSS.n7271 DVSS.n4832 2.24164
R38632 DVSS.n7269 DVSS.n4825 2.24164
R38633 DVSS.n7215 DVSS.n4832 2.24164
R38634 DVSS.n7220 DVSS.n4825 2.24164
R38635 DVSS.n7261 DVSS.n4832 2.24164
R38636 DVSS.n7259 DVSS.n4825 2.24164
R38637 DVSS.n7221 DVSS.n4832 2.24164
R38638 DVSS.n7226 DVSS.n4825 2.24164
R38639 DVSS.n7251 DVSS.n4832 2.24164
R38640 DVSS.n7249 DVSS.n4825 2.24164
R38641 DVSS.n7227 DVSS.n4832 2.24164
R38642 DVSS.n7232 DVSS.n4825 2.24164
R38643 DVSS.n7241 DVSS.n4832 2.24164
R38644 DVSS.n7239 DVSS.n4825 2.24164
R38645 DVSS.n7233 DVSS.n4832 2.24164
R38646 DVSS.n4927 DVSS.n4886 2.24164
R38647 DVSS.n7102 DVSS.n4881 2.24164
R38648 DVSS.n4936 DVSS.n4886 2.24164
R38649 DVSS.n7102 DVSS.n4880 2.24164
R38650 DVSS.n4940 DVSS.n4886 2.24164
R38651 DVSS.n7102 DVSS.n4879 2.24164
R38652 DVSS.n4948 DVSS.n4886 2.24164
R38653 DVSS.n7102 DVSS.n4878 2.24164
R38654 DVSS.n4952 DVSS.n4886 2.24164
R38655 DVSS.n7102 DVSS.n4877 2.24164
R38656 DVSS.n4960 DVSS.n4886 2.24164
R38657 DVSS.n7102 DVSS.n4876 2.24164
R38658 DVSS.n4964 DVSS.n4886 2.24164
R38659 DVSS.n7102 DVSS.n4875 2.24164
R38660 DVSS.n4972 DVSS.n4886 2.24164
R38661 DVSS.n7102 DVSS.n4874 2.24164
R38662 DVSS.n4976 DVSS.n4886 2.24164
R38663 DVSS.n7102 DVSS.n4873 2.24164
R38664 DVSS.n4984 DVSS.n4886 2.24164
R38665 DVSS.n7102 DVSS.n4872 2.24164
R38666 DVSS.n4988 DVSS.n4886 2.24164
R38667 DVSS.n7102 DVSS.n4871 2.24164
R38668 DVSS.n4996 DVSS.n4886 2.24164
R38669 DVSS.n7102 DVSS.n4870 2.24164
R38670 DVSS.n5000 DVSS.n4886 2.24164
R38671 DVSS.n7102 DVSS.n4869 2.24164
R38672 DVSS.n5008 DVSS.n4886 2.24164
R38673 DVSS.n7102 DVSS.n4868 2.24164
R38674 DVSS.n5012 DVSS.n4886 2.24164
R38675 DVSS.n7102 DVSS.n4867 2.24164
R38676 DVSS.n5020 DVSS.n4886 2.24164
R38677 DVSS.n7102 DVSS.n4866 2.24164
R38678 DVSS.n5024 DVSS.n4886 2.24164
R38679 DVSS.n7102 DVSS.n4865 2.24164
R38680 DVSS.n5032 DVSS.n4886 2.24164
R38681 DVSS.n7102 DVSS.n4864 2.24164
R38682 DVSS.n5036 DVSS.n4886 2.24164
R38683 DVSS.n7102 DVSS.n4863 2.24164
R38684 DVSS.n5044 DVSS.n4886 2.24164
R38685 DVSS.n7102 DVSS.n4862 2.24164
R38686 DVSS.n5048 DVSS.n4886 2.24164
R38687 DVSS.n7102 DVSS.n4861 2.24164
R38688 DVSS.n5056 DVSS.n4886 2.24164
R38689 DVSS.n7102 DVSS.n4860 2.24164
R38690 DVSS.n5060 DVSS.n4886 2.24164
R38691 DVSS.n7102 DVSS.n4859 2.24164
R38692 DVSS.n5068 DVSS.n4886 2.24164
R38693 DVSS.n7102 DVSS.n4858 2.24164
R38694 DVSS.n5072 DVSS.n4886 2.24164
R38695 DVSS.n7102 DVSS.n4857 2.24164
R38696 DVSS.n5080 DVSS.n4886 2.24164
R38697 DVSS.n7102 DVSS.n4856 2.24164
R38698 DVSS.n5084 DVSS.n4886 2.24164
R38699 DVSS.n7102 DVSS.n4855 2.24164
R38700 DVSS.n5092 DVSS.n4886 2.24164
R38701 DVSS.n7102 DVSS.n4854 2.24164
R38702 DVSS.n5096 DVSS.n4886 2.24164
R38703 DVSS.n7102 DVSS.n4853 2.24164
R38704 DVSS.n5104 DVSS.n4886 2.24164
R38705 DVSS.n7102 DVSS.n4852 2.24164
R38706 DVSS.n5108 DVSS.n4886 2.24164
R38707 DVSS.n7102 DVSS.n4851 2.24164
R38708 DVSS.n5116 DVSS.n4886 2.24164
R38709 DVSS.n7102 DVSS.n4850 2.24164
R38710 DVSS.n5120 DVSS.n4886 2.24164
R38711 DVSS.n7102 DVSS.n4849 2.24164
R38712 DVSS.n5128 DVSS.n4886 2.24164
R38713 DVSS.n7102 DVSS.n4848 2.24164
R38714 DVSS.n5132 DVSS.n4886 2.24164
R38715 DVSS.n7102 DVSS.n4847 2.24164
R38716 DVSS.n5140 DVSS.n4886 2.24164
R38717 DVSS.n7102 DVSS.n4846 2.24164
R38718 DVSS.n5144 DVSS.n4886 2.24164
R38719 DVSS.n7102 DVSS.n4845 2.24164
R38720 DVSS.n5152 DVSS.n4886 2.24164
R38721 DVSS.n7102 DVSS.n4844 2.24164
R38722 DVSS.n5156 DVSS.n4886 2.24164
R38723 DVSS.n7102 DVSS.n4843 2.24164
R38724 DVSS.n5164 DVSS.n4886 2.24164
R38725 DVSS.n7102 DVSS.n4842 2.24164
R38726 DVSS.n5168 DVSS.n4886 2.24164
R38727 DVSS.n7102 DVSS.n4841 2.24164
R38728 DVSS.n7100 DVSS.n4886 2.24164
R38729 DVSS.n5273 DVSS.n5182 2.24164
R38730 DVSS.n5275 DVSS.n5184 2.24164
R38731 DVSS.n5277 DVSS.n5182 2.24164
R38732 DVSS.n5266 DVSS.n5184 2.24164
R38733 DVSS.n5285 DVSS.n5182 2.24164
R38734 DVSS.n5287 DVSS.n5184 2.24164
R38735 DVSS.n5289 DVSS.n5182 2.24164
R38736 DVSS.n5262 DVSS.n5184 2.24164
R38737 DVSS.n5297 DVSS.n5182 2.24164
R38738 DVSS.n5299 DVSS.n5184 2.24164
R38739 DVSS.n5301 DVSS.n5182 2.24164
R38740 DVSS.n5258 DVSS.n5184 2.24164
R38741 DVSS.n5309 DVSS.n5182 2.24164
R38742 DVSS.n5311 DVSS.n5184 2.24164
R38743 DVSS.n5313 DVSS.n5182 2.24164
R38744 DVSS.n5254 DVSS.n5184 2.24164
R38745 DVSS.n5321 DVSS.n5182 2.24164
R38746 DVSS.n5323 DVSS.n5184 2.24164
R38747 DVSS.n5325 DVSS.n5182 2.24164
R38748 DVSS.n5250 DVSS.n5184 2.24164
R38749 DVSS.n5333 DVSS.n5182 2.24164
R38750 DVSS.n5335 DVSS.n5184 2.24164
R38751 DVSS.n5337 DVSS.n5182 2.24164
R38752 DVSS.n5246 DVSS.n5184 2.24164
R38753 DVSS.n5345 DVSS.n5182 2.24164
R38754 DVSS.n5347 DVSS.n5184 2.24164
R38755 DVSS.n5349 DVSS.n5182 2.24164
R38756 DVSS.n5242 DVSS.n5184 2.24164
R38757 DVSS.n5357 DVSS.n5182 2.24164
R38758 DVSS.n5359 DVSS.n5184 2.24164
R38759 DVSS.n5361 DVSS.n5182 2.24164
R38760 DVSS.n5238 DVSS.n5184 2.24164
R38761 DVSS.n5369 DVSS.n5182 2.24164
R38762 DVSS.n5371 DVSS.n5184 2.24164
R38763 DVSS.n5373 DVSS.n5182 2.24164
R38764 DVSS.n5234 DVSS.n5184 2.24164
R38765 DVSS.n5381 DVSS.n5182 2.24164
R38766 DVSS.n5383 DVSS.n5184 2.24164
R38767 DVSS.n5385 DVSS.n5182 2.24164
R38768 DVSS.n5230 DVSS.n5184 2.24164
R38769 DVSS.n5393 DVSS.n5182 2.24164
R38770 DVSS.n5395 DVSS.n5184 2.24164
R38771 DVSS.n5397 DVSS.n5182 2.24164
R38772 DVSS.n5226 DVSS.n5184 2.24164
R38773 DVSS.n5405 DVSS.n5182 2.24164
R38774 DVSS.n5407 DVSS.n5184 2.24164
R38775 DVSS.n5409 DVSS.n5182 2.24164
R38776 DVSS.n5222 DVSS.n5184 2.24164
R38777 DVSS.n5417 DVSS.n5182 2.24164
R38778 DVSS.n5419 DVSS.n5184 2.24164
R38779 DVSS.n5421 DVSS.n5182 2.24164
R38780 DVSS.n5218 DVSS.n5184 2.24164
R38781 DVSS.n5429 DVSS.n5182 2.24164
R38782 DVSS.n5431 DVSS.n5184 2.24164
R38783 DVSS.n5433 DVSS.n5182 2.24164
R38784 DVSS.n5214 DVSS.n5184 2.24164
R38785 DVSS.n5441 DVSS.n5182 2.24164
R38786 DVSS.n5443 DVSS.n5184 2.24164
R38787 DVSS.n5445 DVSS.n5182 2.24164
R38788 DVSS.n5210 DVSS.n5184 2.24164
R38789 DVSS.n5453 DVSS.n5182 2.24164
R38790 DVSS.n5455 DVSS.n5184 2.24164
R38791 DVSS.n5457 DVSS.n5182 2.24164
R38792 DVSS.n5206 DVSS.n5184 2.24164
R38793 DVSS.n5465 DVSS.n5182 2.24164
R38794 DVSS.n5467 DVSS.n5184 2.24164
R38795 DVSS.n5469 DVSS.n5182 2.24164
R38796 DVSS.n5202 DVSS.n5184 2.24164
R38797 DVSS.n5477 DVSS.n5182 2.24164
R38798 DVSS.n5479 DVSS.n5184 2.24164
R38799 DVSS.n5481 DVSS.n5182 2.24164
R38800 DVSS.n5198 DVSS.n5184 2.24164
R38801 DVSS.n5489 DVSS.n5182 2.24164
R38802 DVSS.n5491 DVSS.n5184 2.24164
R38803 DVSS.n5493 DVSS.n5182 2.24164
R38804 DVSS.n5194 DVSS.n5184 2.24164
R38805 DVSS.n5501 DVSS.n5182 2.24164
R38806 DVSS.n5503 DVSS.n5184 2.24164
R38807 DVSS.n5505 DVSS.n5182 2.24164
R38808 DVSS.n5190 DVSS.n5184 2.24164
R38809 DVSS.n5514 DVSS.n5182 2.24164
R38810 DVSS.n5516 DVSS.n5184 2.24164
R38811 DVSS.n5518 DVSS.n5182 2.24164
R38812 DVSS.n5618 DVSS.n5577 2.24164
R38813 DVSS.n7059 DVSS.n5572 2.24164
R38814 DVSS.n5627 DVSS.n5577 2.24164
R38815 DVSS.n7059 DVSS.n5571 2.24164
R38816 DVSS.n5631 DVSS.n5577 2.24164
R38817 DVSS.n7059 DVSS.n5570 2.24164
R38818 DVSS.n5639 DVSS.n5577 2.24164
R38819 DVSS.n7059 DVSS.n5569 2.24164
R38820 DVSS.n5643 DVSS.n5577 2.24164
R38821 DVSS.n7059 DVSS.n5568 2.24164
R38822 DVSS.n5651 DVSS.n5577 2.24164
R38823 DVSS.n7059 DVSS.n5567 2.24164
R38824 DVSS.n5655 DVSS.n5577 2.24164
R38825 DVSS.n7059 DVSS.n5566 2.24164
R38826 DVSS.n5663 DVSS.n5577 2.24164
R38827 DVSS.n7059 DVSS.n5565 2.24164
R38828 DVSS.n5667 DVSS.n5577 2.24164
R38829 DVSS.n7059 DVSS.n5564 2.24164
R38830 DVSS.n5675 DVSS.n5577 2.24164
R38831 DVSS.n7059 DVSS.n5563 2.24164
R38832 DVSS.n5679 DVSS.n5577 2.24164
R38833 DVSS.n7059 DVSS.n5562 2.24164
R38834 DVSS.n5687 DVSS.n5577 2.24164
R38835 DVSS.n7059 DVSS.n5561 2.24164
R38836 DVSS.n5691 DVSS.n5577 2.24164
R38837 DVSS.n7059 DVSS.n5560 2.24164
R38838 DVSS.n5699 DVSS.n5577 2.24164
R38839 DVSS.n7059 DVSS.n5559 2.24164
R38840 DVSS.n5703 DVSS.n5577 2.24164
R38841 DVSS.n7059 DVSS.n5558 2.24164
R38842 DVSS.n5711 DVSS.n5577 2.24164
R38843 DVSS.n7059 DVSS.n5557 2.24164
R38844 DVSS.n5715 DVSS.n5577 2.24164
R38845 DVSS.n7059 DVSS.n5556 2.24164
R38846 DVSS.n5723 DVSS.n5577 2.24164
R38847 DVSS.n7059 DVSS.n5555 2.24164
R38848 DVSS.n5727 DVSS.n5577 2.24164
R38849 DVSS.n7059 DVSS.n5554 2.24164
R38850 DVSS.n5735 DVSS.n5577 2.24164
R38851 DVSS.n7059 DVSS.n5553 2.24164
R38852 DVSS.n5739 DVSS.n5577 2.24164
R38853 DVSS.n7059 DVSS.n5552 2.24164
R38854 DVSS.n5747 DVSS.n5577 2.24164
R38855 DVSS.n7059 DVSS.n5551 2.24164
R38856 DVSS.n5751 DVSS.n5577 2.24164
R38857 DVSS.n7059 DVSS.n5550 2.24164
R38858 DVSS.n5759 DVSS.n5577 2.24164
R38859 DVSS.n7059 DVSS.n5549 2.24164
R38860 DVSS.n5763 DVSS.n5577 2.24164
R38861 DVSS.n7059 DVSS.n5548 2.24164
R38862 DVSS.n5771 DVSS.n5577 2.24164
R38863 DVSS.n7059 DVSS.n5547 2.24164
R38864 DVSS.n5775 DVSS.n5577 2.24164
R38865 DVSS.n7059 DVSS.n5546 2.24164
R38866 DVSS.n5783 DVSS.n5577 2.24164
R38867 DVSS.n7059 DVSS.n5545 2.24164
R38868 DVSS.n5787 DVSS.n5577 2.24164
R38869 DVSS.n7059 DVSS.n5544 2.24164
R38870 DVSS.n5795 DVSS.n5577 2.24164
R38871 DVSS.n7059 DVSS.n5543 2.24164
R38872 DVSS.n5799 DVSS.n5577 2.24164
R38873 DVSS.n7059 DVSS.n5542 2.24164
R38874 DVSS.n5807 DVSS.n5577 2.24164
R38875 DVSS.n7059 DVSS.n5541 2.24164
R38876 DVSS.n5811 DVSS.n5577 2.24164
R38877 DVSS.n7059 DVSS.n5540 2.24164
R38878 DVSS.n5819 DVSS.n5577 2.24164
R38879 DVSS.n7059 DVSS.n5539 2.24164
R38880 DVSS.n5823 DVSS.n5577 2.24164
R38881 DVSS.n7059 DVSS.n5538 2.24164
R38882 DVSS.n5831 DVSS.n5577 2.24164
R38883 DVSS.n7059 DVSS.n5537 2.24164
R38884 DVSS.n5835 DVSS.n5577 2.24164
R38885 DVSS.n7059 DVSS.n5536 2.24164
R38886 DVSS.n5843 DVSS.n5577 2.24164
R38887 DVSS.n7059 DVSS.n5535 2.24164
R38888 DVSS.n5847 DVSS.n5577 2.24164
R38889 DVSS.n7059 DVSS.n5534 2.24164
R38890 DVSS.n5855 DVSS.n5577 2.24164
R38891 DVSS.n7059 DVSS.n5533 2.24164
R38892 DVSS.n5859 DVSS.n5577 2.24164
R38893 DVSS.n7059 DVSS.n5532 2.24164
R38894 DVSS.n7057 DVSS.n5577 2.24164
R38895 DVSS.n6776 DVSS.n5880 2.24164
R38896 DVSS.n6782 DVSS.n5878 2.24164
R38897 DVSS.n6784 DVSS.n5880 2.24164
R38898 DVSS.n6786 DVSS.n5878 2.24164
R38899 DVSS.n6772 DVSS.n5880 2.24164
R38900 DVSS.n6794 DVSS.n5878 2.24164
R38901 DVSS.n6796 DVSS.n5880 2.24164
R38902 DVSS.n6798 DVSS.n5878 2.24164
R38903 DVSS.n6768 DVSS.n5880 2.24164
R38904 DVSS.n6806 DVSS.n5878 2.24164
R38905 DVSS.n6808 DVSS.n5880 2.24164
R38906 DVSS.n6810 DVSS.n5878 2.24164
R38907 DVSS.n6764 DVSS.n5880 2.24164
R38908 DVSS.n6818 DVSS.n5878 2.24164
R38909 DVSS.n6820 DVSS.n5880 2.24164
R38910 DVSS.n6822 DVSS.n5878 2.24164
R38911 DVSS.n6760 DVSS.n5880 2.24164
R38912 DVSS.n6830 DVSS.n5878 2.24164
R38913 DVSS.n6832 DVSS.n5880 2.24164
R38914 DVSS.n6834 DVSS.n5878 2.24164
R38915 DVSS.n6756 DVSS.n5880 2.24164
R38916 DVSS.n6842 DVSS.n5878 2.24164
R38917 DVSS.n6844 DVSS.n5880 2.24164
R38918 DVSS.n6846 DVSS.n5878 2.24164
R38919 DVSS.n6752 DVSS.n5880 2.24164
R38920 DVSS.n6854 DVSS.n5878 2.24164
R38921 DVSS.n6856 DVSS.n5880 2.24164
R38922 DVSS.n6858 DVSS.n5878 2.24164
R38923 DVSS.n6748 DVSS.n5880 2.24164
R38924 DVSS.n6866 DVSS.n5878 2.24164
R38925 DVSS.n6868 DVSS.n5880 2.24164
R38926 DVSS.n6870 DVSS.n5878 2.24164
R38927 DVSS.n6744 DVSS.n5880 2.24164
R38928 DVSS.n6878 DVSS.n5878 2.24164
R38929 DVSS.n6880 DVSS.n5880 2.24164
R38930 DVSS.n6882 DVSS.n5878 2.24164
R38931 DVSS.n6740 DVSS.n5880 2.24164
R38932 DVSS.n6890 DVSS.n5878 2.24164
R38933 DVSS.n6892 DVSS.n5880 2.24164
R38934 DVSS.n6894 DVSS.n5878 2.24164
R38935 DVSS.n6736 DVSS.n5880 2.24164
R38936 DVSS.n6902 DVSS.n5878 2.24164
R38937 DVSS.n6904 DVSS.n5880 2.24164
R38938 DVSS.n6906 DVSS.n5878 2.24164
R38939 DVSS.n6732 DVSS.n5880 2.24164
R38940 DVSS.n6914 DVSS.n5878 2.24164
R38941 DVSS.n6916 DVSS.n5880 2.24164
R38942 DVSS.n6918 DVSS.n5878 2.24164
R38943 DVSS.n6728 DVSS.n5880 2.24164
R38944 DVSS.n6926 DVSS.n5878 2.24164
R38945 DVSS.n6928 DVSS.n5880 2.24164
R38946 DVSS.n6930 DVSS.n5878 2.24164
R38947 DVSS.n6724 DVSS.n5880 2.24164
R38948 DVSS.n6938 DVSS.n5878 2.24164
R38949 DVSS.n6940 DVSS.n5880 2.24164
R38950 DVSS.n6942 DVSS.n5878 2.24164
R38951 DVSS.n6720 DVSS.n5880 2.24164
R38952 DVSS.n6950 DVSS.n5878 2.24164
R38953 DVSS.n6952 DVSS.n5880 2.24164
R38954 DVSS.n6954 DVSS.n5878 2.24164
R38955 DVSS.n6716 DVSS.n5880 2.24164
R38956 DVSS.n6962 DVSS.n5878 2.24164
R38957 DVSS.n6964 DVSS.n5880 2.24164
R38958 DVSS.n6966 DVSS.n5878 2.24164
R38959 DVSS.n6712 DVSS.n5880 2.24164
R38960 DVSS.n6974 DVSS.n5878 2.24164
R38961 DVSS.n6976 DVSS.n5880 2.24164
R38962 DVSS.n6978 DVSS.n5878 2.24164
R38963 DVSS.n6708 DVSS.n5880 2.24164
R38964 DVSS.n6986 DVSS.n5878 2.24164
R38965 DVSS.n6988 DVSS.n5880 2.24164
R38966 DVSS.n6990 DVSS.n5878 2.24164
R38967 DVSS.n6704 DVSS.n5880 2.24164
R38968 DVSS.n6998 DVSS.n5878 2.24164
R38969 DVSS.n7000 DVSS.n5880 2.24164
R38970 DVSS.n7002 DVSS.n5878 2.24164
R38971 DVSS.n6700 DVSS.n5880 2.24164
R38972 DVSS.n7010 DVSS.n5878 2.24164
R38973 DVSS.n7012 DVSS.n5880 2.24164
R38974 DVSS.n7014 DVSS.n5878 2.24164
R38975 DVSS.n6696 DVSS.n5880 2.24164
R38976 DVSS.n7022 DVSS.n5878 2.24164
R38977 DVSS.n7024 DVSS.n5880 2.24164
R38978 DVSS.n12088 DVSS.n11631 2.24164
R38979 DVSS.n12336 DVSS.n12043 2.24164
R38980 DVSS.n12095 DVSS.n11631 2.24164
R38981 DVSS.n12336 DVSS.n12042 2.24164
R38982 DVSS.n12099 DVSS.n11631 2.24164
R38983 DVSS.n12336 DVSS.n12041 2.24164
R38984 DVSS.n12107 DVSS.n11631 2.24164
R38985 DVSS.n12336 DVSS.n12040 2.24164
R38986 DVSS.n12111 DVSS.n11631 2.24164
R38987 DVSS.n12336 DVSS.n12039 2.24164
R38988 DVSS.n12119 DVSS.n11631 2.24164
R38989 DVSS.n12336 DVSS.n12038 2.24164
R38990 DVSS.n12123 DVSS.n11631 2.24164
R38991 DVSS.n12336 DVSS.n12037 2.24164
R38992 DVSS.n12131 DVSS.n11631 2.24164
R38993 DVSS.n12336 DVSS.n12036 2.24164
R38994 DVSS.n12135 DVSS.n11631 2.24164
R38995 DVSS.n12336 DVSS.n12035 2.24164
R38996 DVSS.n12143 DVSS.n11631 2.24164
R38997 DVSS.n12336 DVSS.n12034 2.24164
R38998 DVSS.n12147 DVSS.n11631 2.24164
R38999 DVSS.n12336 DVSS.n12033 2.24164
R39000 DVSS.n12155 DVSS.n11631 2.24164
R39001 DVSS.n12336 DVSS.n12032 2.24164
R39002 DVSS.n12159 DVSS.n11631 2.24164
R39003 DVSS.n12336 DVSS.n12031 2.24164
R39004 DVSS.n12167 DVSS.n11631 2.24164
R39005 DVSS.n12336 DVSS.n12030 2.24164
R39006 DVSS.n12171 DVSS.n11631 2.24164
R39007 DVSS.n12336 DVSS.n12029 2.24164
R39008 DVSS.n12179 DVSS.n11631 2.24164
R39009 DVSS.n12336 DVSS.n12028 2.24164
R39010 DVSS.n12183 DVSS.n11631 2.24164
R39011 DVSS.n12336 DVSS.n12027 2.24164
R39012 DVSS.n12191 DVSS.n11631 2.24164
R39013 DVSS.n12336 DVSS.n12026 2.24164
R39014 DVSS.n12195 DVSS.n11631 2.24164
R39015 DVSS.n12336 DVSS.n12025 2.24164
R39016 DVSS.n12203 DVSS.n11631 2.24164
R39017 DVSS.n12336 DVSS.n12024 2.24164
R39018 DVSS.n12207 DVSS.n11631 2.24164
R39019 DVSS.n12336 DVSS.n12023 2.24164
R39020 DVSS.n12215 DVSS.n11631 2.24164
R39021 DVSS.n12336 DVSS.n12022 2.24164
R39022 DVSS.n12219 DVSS.n11631 2.24164
R39023 DVSS.n12336 DVSS.n12021 2.24164
R39024 DVSS.n12227 DVSS.n11631 2.24164
R39025 DVSS.n12336 DVSS.n12020 2.24164
R39026 DVSS.n12231 DVSS.n11631 2.24164
R39027 DVSS.n12336 DVSS.n12019 2.24164
R39028 DVSS.n12239 DVSS.n11631 2.24164
R39029 DVSS.n12336 DVSS.n12018 2.24164
R39030 DVSS.n12243 DVSS.n11631 2.24164
R39031 DVSS.n12336 DVSS.n12017 2.24164
R39032 DVSS.n12251 DVSS.n11631 2.24164
R39033 DVSS.n12336 DVSS.n12016 2.24164
R39034 DVSS.n12255 DVSS.n11631 2.24164
R39035 DVSS.n12336 DVSS.n12015 2.24164
R39036 DVSS.n12263 DVSS.n11631 2.24164
R39037 DVSS.n12336 DVSS.n12014 2.24164
R39038 DVSS.n12267 DVSS.n11631 2.24164
R39039 DVSS.n12336 DVSS.n12013 2.24164
R39040 DVSS.n12275 DVSS.n11631 2.24164
R39041 DVSS.n12336 DVSS.n12012 2.24164
R39042 DVSS.n12279 DVSS.n11631 2.24164
R39043 DVSS.n12336 DVSS.n12011 2.24164
R39044 DVSS.n12287 DVSS.n11631 2.24164
R39045 DVSS.n12336 DVSS.n12010 2.24164
R39046 DVSS.n12291 DVSS.n11631 2.24164
R39047 DVSS.n12336 DVSS.n12009 2.24164
R39048 DVSS.n12299 DVSS.n11631 2.24164
R39049 DVSS.n12336 DVSS.n12008 2.24164
R39050 DVSS.n12303 DVSS.n11631 2.24164
R39051 DVSS.n12336 DVSS.n12007 2.24164
R39052 DVSS.n12311 DVSS.n11631 2.24164
R39053 DVSS.n12336 DVSS.n12006 2.24164
R39054 DVSS.n12315 DVSS.n11631 2.24164
R39055 DVSS.n12336 DVSS.n12005 2.24164
R39056 DVSS.n12323 DVSS.n11631 2.24164
R39057 DVSS.n12336 DVSS.n12004 2.24164
R39058 DVSS.n12327 DVSS.n11631 2.24164
R39059 DVSS.n12336 DVSS.n12003 2.24164
R39060 DVSS.n12045 DVSS.n11631 2.24164
R39061 DVSS.n6231 DVSS.n6230 2.24164
R39062 DVSS.n5939 DVSS.n5888 2.24164
R39063 DVSS.n6231 DVSS.n5937 2.24164
R39064 DVSS.n6222 DVSS.n5888 2.24164
R39065 DVSS.n6231 DVSS.n5936 2.24164
R39066 DVSS.n6217 DVSS.n5888 2.24164
R39067 DVSS.n6231 DVSS.n5935 2.24164
R39068 DVSS.n6210 DVSS.n5888 2.24164
R39069 DVSS.n6231 DVSS.n5934 2.24164
R39070 DVSS.n6205 DVSS.n5888 2.24164
R39071 DVSS.n6231 DVSS.n5933 2.24164
R39072 DVSS.n6198 DVSS.n5888 2.24164
R39073 DVSS.n6231 DVSS.n5932 2.24164
R39074 DVSS.n6193 DVSS.n5888 2.24164
R39075 DVSS.n6231 DVSS.n5931 2.24164
R39076 DVSS.n6186 DVSS.n5888 2.24164
R39077 DVSS.n6231 DVSS.n5930 2.24164
R39078 DVSS.n6181 DVSS.n5888 2.24164
R39079 DVSS.n6231 DVSS.n5929 2.24164
R39080 DVSS.n6174 DVSS.n5888 2.24164
R39081 DVSS.n6231 DVSS.n5928 2.24164
R39082 DVSS.n6169 DVSS.n5888 2.24164
R39083 DVSS.n6231 DVSS.n5927 2.24164
R39084 DVSS.n6162 DVSS.n5888 2.24164
R39085 DVSS.n6231 DVSS.n5926 2.24164
R39086 DVSS.n6157 DVSS.n5888 2.24164
R39087 DVSS.n6231 DVSS.n5925 2.24164
R39088 DVSS.n6150 DVSS.n5888 2.24164
R39089 DVSS.n6231 DVSS.n5924 2.24164
R39090 DVSS.n6145 DVSS.n5888 2.24164
R39091 DVSS.n6231 DVSS.n5923 2.24164
R39092 DVSS.n6138 DVSS.n5888 2.24164
R39093 DVSS.n6231 DVSS.n5922 2.24164
R39094 DVSS.n6133 DVSS.n5888 2.24164
R39095 DVSS.n6231 DVSS.n5921 2.24164
R39096 DVSS.n6126 DVSS.n5888 2.24164
R39097 DVSS.n6231 DVSS.n5920 2.24164
R39098 DVSS.n6121 DVSS.n5888 2.24164
R39099 DVSS.n6231 DVSS.n5919 2.24164
R39100 DVSS.n6114 DVSS.n5888 2.24164
R39101 DVSS.n6231 DVSS.n5918 2.24164
R39102 DVSS.n6109 DVSS.n5888 2.24164
R39103 DVSS.n6231 DVSS.n5917 2.24164
R39104 DVSS.n6102 DVSS.n5888 2.24164
R39105 DVSS.n6231 DVSS.n5916 2.24164
R39106 DVSS.n6097 DVSS.n5888 2.24164
R39107 DVSS.n6231 DVSS.n5915 2.24164
R39108 DVSS.n6090 DVSS.n5888 2.24164
R39109 DVSS.n6231 DVSS.n5914 2.24164
R39110 DVSS.n6085 DVSS.n5888 2.24164
R39111 DVSS.n6231 DVSS.n5913 2.24164
R39112 DVSS.n6078 DVSS.n5888 2.24164
R39113 DVSS.n6231 DVSS.n5912 2.24164
R39114 DVSS.n6073 DVSS.n5888 2.24164
R39115 DVSS.n6231 DVSS.n5911 2.24164
R39116 DVSS.n6066 DVSS.n5888 2.24164
R39117 DVSS.n6231 DVSS.n5910 2.24164
R39118 DVSS.n6061 DVSS.n5888 2.24164
R39119 DVSS.n6231 DVSS.n5909 2.24164
R39120 DVSS.n6054 DVSS.n5888 2.24164
R39121 DVSS.n6231 DVSS.n5908 2.24164
R39122 DVSS.n6049 DVSS.n5888 2.24164
R39123 DVSS.n6231 DVSS.n5907 2.24164
R39124 DVSS.n6042 DVSS.n5888 2.24164
R39125 DVSS.n6231 DVSS.n5906 2.24164
R39126 DVSS.n6037 DVSS.n5888 2.24164
R39127 DVSS.n6231 DVSS.n5905 2.24164
R39128 DVSS.n6030 DVSS.n5888 2.24164
R39129 DVSS.n6231 DVSS.n5904 2.24164
R39130 DVSS.n6025 DVSS.n5888 2.24164
R39131 DVSS.n6231 DVSS.n5903 2.24164
R39132 DVSS.n6018 DVSS.n5888 2.24164
R39133 DVSS.n6231 DVSS.n5902 2.24164
R39134 DVSS.n6013 DVSS.n5888 2.24164
R39135 DVSS.n6231 DVSS.n5901 2.24164
R39136 DVSS.n6006 DVSS.n5888 2.24164
R39137 DVSS.n6231 DVSS.n5900 2.24164
R39138 DVSS.n6001 DVSS.n5888 2.24164
R39139 DVSS.n6231 DVSS.n5899 2.24164
R39140 DVSS.n5994 DVSS.n5888 2.24164
R39141 DVSS.n6231 DVSS.n5898 2.24164
R39142 DVSS.n5989 DVSS.n5888 2.24164
R39143 DVSS.n6231 DVSS.n5897 2.24164
R39144 DVSS.n18167 DVSS.n18166 2.24105
R39145 DVSS.n17792 DVSS.n17791 2.24048
R39146 DVSS.n17076 DVSS.n17075 2.24011
R39147 DVSS.n17075 DVSS.n17067 2.24011
R39148 DVSS.n17075 DVSS.n17068 2.24011
R39149 DVSS.n17075 DVSS.n17069 2.24011
R39150 DVSS.n17075 DVSS.n17070 2.24011
R39151 DVSS.n17075 DVSS.n17071 2.24011
R39152 DVSS.n17075 DVSS.n17072 2.24011
R39153 DVSS.n17075 DVSS.n17073 2.24011
R39154 DVSS.n17075 DVSS.n17057 2.24011
R39155 DVSS.n17034 DVSS.n15306 2.24011
R39156 DVSS.n17032 DVSS.n15306 2.24011
R39157 DVSS.n17030 DVSS.n15306 2.24011
R39158 DVSS.n17028 DVSS.n15306 2.24011
R39159 DVSS.n17026 DVSS.n15306 2.24011
R39160 DVSS.n17024 DVSS.n15306 2.24011
R39161 DVSS.n17022 DVSS.n15306 2.24011
R39162 DVSS.n17020 DVSS.n15306 2.24011
R39163 DVSS.n17018 DVSS.n15306 2.24011
R39164 DVSS.n17078 DVSS.n16843 2.24011
R39165 DVSS.n17080 DVSS.n16843 2.24011
R39166 DVSS.n17082 DVSS.n16843 2.24011
R39167 DVSS.n17084 DVSS.n16843 2.24011
R39168 DVSS.n17086 DVSS.n16843 2.24011
R39169 DVSS.n17088 DVSS.n16843 2.24011
R39170 DVSS.n17090 DVSS.n16843 2.24011
R39171 DVSS.n17092 DVSS.n16843 2.24011
R39172 DVSS.n17094 DVSS.n16843 2.24011
R39173 DVSS.n17013 DVSS.n15373 2.24011
R39174 DVSS.n17011 DVSS.n15373 2.24011
R39175 DVSS.n17009 DVSS.n15373 2.24011
R39176 DVSS.n17007 DVSS.n15373 2.24011
R39177 DVSS.n17005 DVSS.n15373 2.24011
R39178 DVSS.n17003 DVSS.n15373 2.24011
R39179 DVSS.n17001 DVSS.n15373 2.24011
R39180 DVSS.n16999 DVSS.n15373 2.24011
R39181 DVSS.n16997 DVSS.n15373 2.24011
R39182 DVSS.n17114 DVSS.n16021 2.24011
R39183 DVSS.n17102 DVSS.n16021 2.24011
R39184 DVSS.n17104 DVSS.n16021 2.24011
R39185 DVSS.n17106 DVSS.n16021 2.24011
R39186 DVSS.n17108 DVSS.n16021 2.24011
R39187 DVSS.n17110 DVSS.n16021 2.24011
R39188 DVSS.n17112 DVSS.n16021 2.24011
R39189 DVSS.n17048 DVSS.n15267 2.24011
R39190 DVSS.n17046 DVSS.n15267 2.24011
R39191 DVSS.n17044 DVSS.n15267 2.24011
R39192 DVSS.n17042 DVSS.n15267 2.24011
R39193 DVSS.n17040 DVSS.n15267 2.24011
R39194 DVSS.n17038 DVSS.n15267 2.24011
R39195 DVSS.n17530 DVSS.n16923 2.24011
R39196 DVSS.n16922 DVSS.n16900 2.24011
R39197 DVSS.n17530 DVSS.n16919 2.24011
R39198 DVSS.n17530 DVSS.n16917 2.24011
R39199 DVSS.n17530 DVSS.n16915 2.24011
R39200 DVSS.n17530 DVSS.n16913 2.24011
R39201 DVSS.n17530 DVSS.n16911 2.24011
R39202 DVSS.n16993 DVSS.n15443 2.24011
R39203 DVSS.n16991 DVSS.n15443 2.24011
R39204 DVSS.n16989 DVSS.n15443 2.24011
R39205 DVSS.n16987 DVSS.n15443 2.24011
R39206 DVSS.n16985 DVSS.n15443 2.24011
R39207 DVSS.n16983 DVSS.n15443 2.24011
R39208 DVSS.n16981 DVSS.n15443 2.24011
R39209 DVSS.n17099 DVSS.n17065 2.24011
R39210 DVSS.n17099 DVSS.n17064 2.24011
R39211 DVSS.n17099 DVSS.n17063 2.24011
R39212 DVSS.n17099 DVSS.n17062 2.24011
R39213 DVSS.n17099 DVSS.n17061 2.24011
R39214 DVSS.n17099 DVSS.n17060 2.24011
R39215 DVSS.n17099 DVSS.n17059 2.24011
R39216 DVSS.n17099 DVSS.n17058 2.24011
R39217 DVSS.n17017 DVSS.n15315 2.24011
R39218 DVSS.n17019 DVSS.n15315 2.24011
R39219 DVSS.n17021 DVSS.n15315 2.24011
R39220 DVSS.n17023 DVSS.n15315 2.24011
R39221 DVSS.n17025 DVSS.n15315 2.24011
R39222 DVSS.n17027 DVSS.n15315 2.24011
R39223 DVSS.n17029 DVSS.n15315 2.24011
R39224 DVSS.n17031 DVSS.n15315 2.24011
R39225 DVSS.n17033 DVSS.n15315 2.24011
R39226 DVSS.n17095 DVSS.n16827 2.24011
R39227 DVSS.n17093 DVSS.n16827 2.24011
R39228 DVSS.n17091 DVSS.n16827 2.24011
R39229 DVSS.n17089 DVSS.n16827 2.24011
R39230 DVSS.n17087 DVSS.n16827 2.24011
R39231 DVSS.n17085 DVSS.n16827 2.24011
R39232 DVSS.n17083 DVSS.n16827 2.24011
R39233 DVSS.n17081 DVSS.n16827 2.24011
R39234 DVSS.n17079 DVSS.n16827 2.24011
R39235 DVSS.n16996 DVSS.n15387 2.24011
R39236 DVSS.n16998 DVSS.n15387 2.24011
R39237 DVSS.n17000 DVSS.n15387 2.24011
R39238 DVSS.n17002 DVSS.n15387 2.24011
R39239 DVSS.n17004 DVSS.n15387 2.24011
R39240 DVSS.n17006 DVSS.n15387 2.24011
R39241 DVSS.n17008 DVSS.n15387 2.24011
R39242 DVSS.n17010 DVSS.n15387 2.24011
R39243 DVSS.n17012 DVSS.n15387 2.24011
R39244 DVSS.n17113 DVSS.n16005 2.24011
R39245 DVSS.n17111 DVSS.n16005 2.24011
R39246 DVSS.n17109 DVSS.n16005 2.24011
R39247 DVSS.n17107 DVSS.n16005 2.24011
R39248 DVSS.n17105 DVSS.n16005 2.24011
R39249 DVSS.n17103 DVSS.n16005 2.24011
R39250 DVSS.n17037 DVSS.n15273 2.24011
R39251 DVSS.n17039 DVSS.n15273 2.24011
R39252 DVSS.n17041 DVSS.n15273 2.24011
R39253 DVSS.n17043 DVSS.n15273 2.24011
R39254 DVSS.n17045 DVSS.n15273 2.24011
R39255 DVSS.n17047 DVSS.n15273 2.24011
R39256 DVSS.n17049 DVSS.n15273 2.24011
R39257 DVSS.n16910 DVSS.n16900 2.24011
R39258 DVSS.n16912 DVSS.n16900 2.24011
R39259 DVSS.n16914 DVSS.n16900 2.24011
R39260 DVSS.n16916 DVSS.n16900 2.24011
R39261 DVSS.n16918 DVSS.n16900 2.24011
R39262 DVSS.n16921 DVSS.n16900 2.24011
R39263 DVSS.n16982 DVSS.n15452 2.24011
R39264 DVSS.n16984 DVSS.n15452 2.24011
R39265 DVSS.n16986 DVSS.n15452 2.24011
R39266 DVSS.n16988 DVSS.n15452 2.24011
R39267 DVSS.n16990 DVSS.n15452 2.24011
R39268 DVSS.n16992 DVSS.n15452 2.24011
R39269 DVSS.n21587 DVSS.n21586 2.23787
R39270 DVSS.n21586 DVSS.n21583 2.23787
R39271 DVSS.n21586 DVSS.n21582 2.23787
R39272 DVSS.n21586 DVSS.n21581 2.23787
R39273 DVSS.n21586 DVSS.n21580 2.23787
R39274 DVSS.n21586 DVSS.n21579 2.23787
R39275 DVSS.n21586 DVSS.n21578 2.23787
R39276 DVSS.n1331 DVSS.n623 2.23787
R39277 DVSS.n1329 DVSS.n623 2.23787
R39278 DVSS.n1327 DVSS.n623 2.23787
R39279 DVSS.n1325 DVSS.n623 2.23787
R39280 DVSS.n1323 DVSS.n623 2.23787
R39281 DVSS.n1321 DVSS.n623 2.23787
R39282 DVSS.n1319 DVSS.n623 2.23787
R39283 DVSS.n1317 DVSS.n623 2.23787
R39284 DVSS.n1315 DVSS.n623 2.23787
R39285 DVSS.n1330 DVSS.n607 2.23787
R39286 DVSS.n1328 DVSS.n607 2.23787
R39287 DVSS.n1326 DVSS.n607 2.23787
R39288 DVSS.n1324 DVSS.n607 2.23787
R39289 DVSS.n1322 DVSS.n607 2.23787
R39290 DVSS.n1320 DVSS.n607 2.23787
R39291 DVSS.n1318 DVSS.n607 2.23787
R39292 DVSS.n1316 DVSS.n607 2.23787
R39293 DVSS.n1314 DVSS.n607 2.23787
R39294 DVSS.n21589 DVSS.n21576 2.23787
R39295 DVSS.n21589 DVSS.n21575 2.23787
R39296 DVSS.n21589 DVSS.n21574 2.23787
R39297 DVSS.n21589 DVSS.n21573 2.23787
R39298 DVSS.n21589 DVSS.n21572 2.23787
R39299 DVSS.n21589 DVSS.n21571 2.23787
R39300 DVSS.n21589 DVSS.n21570 2.23787
R39301 DVSS.n21589 DVSS.n21569 2.23787
R39302 DVSS.n20101 DVSS.n13947 2.23787
R39303 DVSS.n20114 DVSS.n14470 2.23787
R39304 DVSS.n20173 DVSS.n20018 2.23787
R39305 DVSS.n20673 DVSS.n14594 2.23787
R39306 DVSS.n1197 DVSS.n1177 2.23787
R39307 DVSS.n1197 DVSS.n1195 2.23787
R39308 DVSS.n1197 DVSS.n1194 2.23787
R39309 DVSS.n1197 DVSS.n1193 2.23787
R39310 DVSS.n1197 DVSS.n1192 2.23787
R39311 DVSS.n1197 DVSS.n1191 2.23787
R39312 DVSS.n1197 DVSS.n1190 2.23787
R39313 DVSS.n1197 DVSS.n1189 2.23787
R39314 DVSS.n1310 DVSS.n573 2.23787
R39315 DVSS.n1308 DVSS.n573 2.23787
R39316 DVSS.n1306 DVSS.n573 2.23787
R39317 DVSS.n1304 DVSS.n573 2.23787
R39318 DVSS.n1302 DVSS.n573 2.23787
R39319 DVSS.n1300 DVSS.n573 2.23787
R39320 DVSS.n1298 DVSS.n573 2.23787
R39321 DVSS.n1296 DVSS.n573 2.23787
R39322 DVSS.n1294 DVSS.n573 2.23787
R39323 DVSS.n1309 DVSS.n562 2.23787
R39324 DVSS.n1307 DVSS.n562 2.23787
R39325 DVSS.n1305 DVSS.n562 2.23787
R39326 DVSS.n1303 DVSS.n562 2.23787
R39327 DVSS.n1301 DVSS.n562 2.23787
R39328 DVSS.n1299 DVSS.n562 2.23787
R39329 DVSS.n1297 DVSS.n562 2.23787
R39330 DVSS.n1295 DVSS.n562 2.23787
R39331 DVSS.n1293 DVSS.n562 2.23787
R39332 DVSS.n22339 DVSS.n1187 2.23787
R39333 DVSS.n22339 DVSS.n1186 2.23787
R39334 DVSS.n22339 DVSS.n1185 2.23787
R39335 DVSS.n22339 DVSS.n1184 2.23787
R39336 DVSS.n22339 DVSS.n1183 2.23787
R39337 DVSS.n22339 DVSS.n1182 2.23787
R39338 DVSS.n22339 DVSS.n1181 2.23787
R39339 DVSS.n22339 DVSS.n1180 2.23787
R39340 DVSS.n14648 DVSS.n14631 2.23787
R39341 DVSS.n20193 DVSS.n14425 2.23787
R39342 DVSS.n22460 DVSS.n866 2.23787
R39343 DVSS.n22460 DVSS.n865 2.23787
R39344 DVSS.n22460 DVSS.n864 2.23787
R39345 DVSS.n22460 DVSS.n863 2.23787
R39346 DVSS.n22460 DVSS.n862 2.23787
R39347 DVSS.n22460 DVSS.n861 2.23787
R39348 DVSS.n22460 DVSS.n860 2.23787
R39349 DVSS.n22460 DVSS.n859 2.23787
R39350 DVSS.n1351 DVSS.n680 2.23787
R39351 DVSS.n1349 DVSS.n680 2.23787
R39352 DVSS.n1347 DVSS.n680 2.23787
R39353 DVSS.n1345 DVSS.n680 2.23787
R39354 DVSS.n1343 DVSS.n680 2.23787
R39355 DVSS.n1341 DVSS.n680 2.23787
R39356 DVSS.n1339 DVSS.n680 2.23787
R39357 DVSS.n1337 DVSS.n680 2.23787
R39358 DVSS.n1335 DVSS.n680 2.23787
R39359 DVSS.n1350 DVSS.n669 2.23787
R39360 DVSS.n1348 DVSS.n669 2.23787
R39361 DVSS.n1346 DVSS.n669 2.23787
R39362 DVSS.n1344 DVSS.n669 2.23787
R39363 DVSS.n1342 DVSS.n669 2.23787
R39364 DVSS.n1340 DVSS.n669 2.23787
R39365 DVSS.n1338 DVSS.n669 2.23787
R39366 DVSS.n1336 DVSS.n669 2.23787
R39367 DVSS.n1334 DVSS.n669 2.23787
R39368 DVSS.n22458 DVSS.n878 2.23787
R39369 DVSS.n22458 DVSS.n877 2.23787
R39370 DVSS.n22458 DVSS.n876 2.23787
R39371 DVSS.n22458 DVSS.n875 2.23787
R39372 DVSS.n22458 DVSS.n874 2.23787
R39373 DVSS.n22458 DVSS.n873 2.23787
R39374 DVSS.n22458 DVSS.n872 2.23787
R39375 DVSS.n22458 DVSS.n871 2.23787
R39376 DVSS.n20688 DVSS.n14547 2.23787
R39377 DVSS.n20699 DVSS.n14522 2.23787
R39378 DVSS.n20697 DVSS.n20696 2.23787
R39379 DVSS.n20690 DVSS.n14548 2.23787
R39380 DVSS.n19515 DVSS.n19514 2.23787
R39381 DVSS.n19515 DVSS.n19277 2.23787
R39382 DVSS.n19515 DVSS.n19276 2.23787
R39383 DVSS.n19515 DVSS.n19275 2.23787
R39384 DVSS.n19515 DVSS.n19274 2.23787
R39385 DVSS.n19515 DVSS.n19273 2.23787
R39386 DVSS.n19515 DVSS.n19272 2.23787
R39387 DVSS.n19515 DVSS.n19271 2.23787
R39388 DVSS.n19515 DVSS.n19270 2.23787
R39389 DVSS.n19592 DVSS.n19267 2.23787
R39390 DVSS.n19592 DVSS.n19265 2.23787
R39391 DVSS.n19592 DVSS.n19263 2.23787
R39392 DVSS.n19592 DVSS.n19261 2.23787
R39393 DVSS.n19592 DVSS.n19259 2.23787
R39394 DVSS.n19592 DVSS.n19257 2.23787
R39395 DVSS.n19592 DVSS.n19255 2.23787
R39396 DVSS.n19592 DVSS.n19253 2.23787
R39397 DVSS.n19089 DVSS.n19087 2.23787
R39398 DVSS.n19089 DVSS.n19086 2.23787
R39399 DVSS.n19089 DVSS.n19085 2.23787
R39400 DVSS.n19089 DVSS.n19084 2.23787
R39401 DVSS.n19089 DVSS.n19083 2.23787
R39402 DVSS.n19089 DVSS.n19082 2.23787
R39403 DVSS.n19089 DVSS.n19081 2.23787
R39404 DVSS.n19089 DVSS.n19080 2.23787
R39405 DVSS.n19512 DVSS.n19278 2.23787
R39406 DVSS.n19512 DVSS.n19511 2.23787
R39407 DVSS.n19512 DVSS.n19510 2.23787
R39408 DVSS.n19512 DVSS.n19509 2.23787
R39409 DVSS.n19512 DVSS.n19508 2.23787
R39410 DVSS.n19512 DVSS.n19507 2.23787
R39411 DVSS.n19512 DVSS.n19506 2.23787
R39412 DVSS.n19512 DVSS.n19505 2.23787
R39413 DVSS.n19266 DVSS.n19065 2.23787
R39414 DVSS.n19264 DVSS.n19065 2.23787
R39415 DVSS.n19262 DVSS.n19065 2.23787
R39416 DVSS.n19260 DVSS.n19065 2.23787
R39417 DVSS.n19258 DVSS.n19065 2.23787
R39418 DVSS.n19256 DVSS.n19065 2.23787
R39419 DVSS.n19254 DVSS.n19065 2.23787
R39420 DVSS.n19590 DVSS.n19065 2.23787
R39421 DVSS.n19850 DVSS.n19077 2.23787
R39422 DVSS.n19850 DVSS.n19076 2.23787
R39423 DVSS.n19850 DVSS.n19075 2.23787
R39424 DVSS.n19850 DVSS.n19074 2.23787
R39425 DVSS.n19850 DVSS.n19073 2.23787
R39426 DVSS.n19850 DVSS.n19072 2.23787
R39427 DVSS.n19850 DVSS.n19071 2.23787
R39428 DVSS.n19850 DVSS.n19070 2.23787
R39429 DVSS.n1218 DVSS.n1198 2.23787
R39430 DVSS.n1218 DVSS.n1216 2.23787
R39431 DVSS.n1218 DVSS.n1215 2.23787
R39432 DVSS.n1218 DVSS.n1214 2.23787
R39433 DVSS.n1218 DVSS.n1213 2.23787
R39434 DVSS.n1218 DVSS.n1212 2.23787
R39435 DVSS.n1218 DVSS.n1211 2.23787
R39436 DVSS.n1218 DVSS.n1210 2.23787
R39437 DVSS.n1290 DVSS.n523 2.23787
R39438 DVSS.n1288 DVSS.n523 2.23787
R39439 DVSS.n1286 DVSS.n523 2.23787
R39440 DVSS.n1284 DVSS.n523 2.23787
R39441 DVSS.n1282 DVSS.n523 2.23787
R39442 DVSS.n1280 DVSS.n523 2.23787
R39443 DVSS.n1278 DVSS.n523 2.23787
R39444 DVSS.n1276 DVSS.n523 2.23787
R39445 DVSS.n1274 DVSS.n523 2.23787
R39446 DVSS.n19109 DVSS.n19090 2.23787
R39447 DVSS.n19109 DVSS.n19107 2.23787
R39448 DVSS.n19109 DVSS.n19106 2.23787
R39449 DVSS.n19109 DVSS.n19105 2.23787
R39450 DVSS.n19109 DVSS.n19104 2.23787
R39451 DVSS.n19109 DVSS.n19103 2.23787
R39452 DVSS.n19109 DVSS.n19102 2.23787
R39453 DVSS.n19109 DVSS.n19101 2.23787
R39454 DVSS.n19847 DVSS.n19099 2.23787
R39455 DVSS.n19847 DVSS.n19098 2.23787
R39456 DVSS.n19847 DVSS.n19097 2.23787
R39457 DVSS.n19847 DVSS.n19096 2.23787
R39458 DVSS.n19847 DVSS.n19095 2.23787
R39459 DVSS.n19847 DVSS.n19094 2.23787
R39460 DVSS.n19847 DVSS.n19093 2.23787
R39461 DVSS.n19847 DVSS.n19092 2.23787
R39462 DVSS.n1289 DVSS.n507 2.23787
R39463 DVSS.n1287 DVSS.n507 2.23787
R39464 DVSS.n1285 DVSS.n507 2.23787
R39465 DVSS.n1283 DVSS.n507 2.23787
R39466 DVSS.n1281 DVSS.n507 2.23787
R39467 DVSS.n1279 DVSS.n507 2.23787
R39468 DVSS.n1277 DVSS.n507 2.23787
R39469 DVSS.n1275 DVSS.n507 2.23787
R39470 DVSS.n1273 DVSS.n507 2.23787
R39471 DVSS.n22336 DVSS.n1208 2.23787
R39472 DVSS.n22336 DVSS.n1207 2.23787
R39473 DVSS.n22336 DVSS.n1206 2.23787
R39474 DVSS.n22336 DVSS.n1205 2.23787
R39475 DVSS.n22336 DVSS.n1204 2.23787
R39476 DVSS.n22336 DVSS.n1203 2.23787
R39477 DVSS.n22336 DVSS.n1202 2.23787
R39478 DVSS.n22336 DVSS.n1201 2.23787
R39479 DVSS.n20358 DVSS.n14668 2.23787
R39480 DVSS.n20352 DVSS.n14376 2.23787
R39481 DVSS.n20458 DVSS.n14857 2.23787
R39482 DVSS.n20432 DVSS.n13430 2.23787
R39483 DVSS.n19193 DVSS.n19186 2.1857
R39484 DVSS.n18516 DVSS.n18515 2.1175
R39485 DVSS.n20505 DVSS.n14704 1.95638
R39486 DVSS.n20505 DVSS.n20504 1.95638
R39487 DVSS.n20469 DVSS.n14707 1.95638
R39488 DVSS.n20472 DVSS.n20469 1.95638
R39489 DVSS.n20464 DVSS.n14850 1.95638
R39490 DVSS.n20467 DVSS.n14850 1.95638
R39491 DVSS.n18999 DVSS.n13581 1.89754
R39492 DVSS.n18997 DVSS.n18583 1.89035
R39493 DVSS.n18995 DVSS.n18640 1.89035
R39494 DVSS.n18997 DVSS.n18582 1.89035
R39495 DVSS.n18995 DVSS.n18639 1.89035
R39496 DVSS.n18997 DVSS.n18581 1.89035
R39497 DVSS.n18995 DVSS.n18638 1.89035
R39498 DVSS.n18997 DVSS.n18580 1.89035
R39499 DVSS.n18995 DVSS.n18637 1.89035
R39500 DVSS.n18997 DVSS.n18579 1.89035
R39501 DVSS.n18995 DVSS.n18636 1.89035
R39502 DVSS.n18997 DVSS.n18578 1.89035
R39503 DVSS.n18995 DVSS.n18635 1.89035
R39504 DVSS.n18997 DVSS.n18577 1.89035
R39505 DVSS.n18995 DVSS.n18634 1.89035
R39506 DVSS.n18997 DVSS.n18576 1.89035
R39507 DVSS.n18995 DVSS.n18633 1.89035
R39508 DVSS.n18997 DVSS.n18575 1.89035
R39509 DVSS.n18995 DVSS.n18632 1.89035
R39510 DVSS.n18997 DVSS.n18574 1.89035
R39511 DVSS.n18995 DVSS.n18631 1.89035
R39512 DVSS.n18997 DVSS.n18573 1.89035
R39513 DVSS.n18995 DVSS.n18630 1.89035
R39514 DVSS.n18997 DVSS.n18572 1.89035
R39515 DVSS.n18995 DVSS.n18629 1.89035
R39516 DVSS.n18997 DVSS.n18571 1.89035
R39517 DVSS.n18995 DVSS.n18628 1.89035
R39518 DVSS.n18997 DVSS.n18570 1.89035
R39519 DVSS.n18995 DVSS.n18627 1.89035
R39520 DVSS.n18997 DVSS.n18569 1.89035
R39521 DVSS.n18995 DVSS.n18626 1.89035
R39522 DVSS.n18997 DVSS.n18568 1.89035
R39523 DVSS.n18995 DVSS.n18625 1.89035
R39524 DVSS.n18997 DVSS.n18567 1.89035
R39525 DVSS.n18995 DVSS.n18624 1.89035
R39526 DVSS.n18997 DVSS.n18566 1.89035
R39527 DVSS.n18995 DVSS.n18623 1.89035
R39528 DVSS.n18997 DVSS.n18565 1.89035
R39529 DVSS.n18995 DVSS.n18622 1.89035
R39530 DVSS.n18997 DVSS.n18564 1.89035
R39531 DVSS.n18995 DVSS.n18621 1.89035
R39532 DVSS.n18997 DVSS.n18563 1.89035
R39533 DVSS.n18995 DVSS.n18620 1.89035
R39534 DVSS.n18997 DVSS.n18562 1.89035
R39535 DVSS.n18995 DVSS.n18619 1.89035
R39536 DVSS.n18997 DVSS.n18561 1.89035
R39537 DVSS.n18995 DVSS.n18618 1.89035
R39538 DVSS.n18997 DVSS.n18560 1.89035
R39539 DVSS.n18995 DVSS.n18617 1.89035
R39540 DVSS.n18997 DVSS.n18559 1.89035
R39541 DVSS.n18995 DVSS.n18616 1.89035
R39542 DVSS.n18761 DVSS.n18760 1.89035
R39543 DVSS.n18995 DVSS.n18615 1.89035
R39544 DVSS.n18761 DVSS.n18759 1.89035
R39545 DVSS.n18995 DVSS.n18614 1.89035
R39546 DVSS.n18761 DVSS.n18758 1.89035
R39547 DVSS.n18995 DVSS.n18613 1.89035
R39548 DVSS.n18997 DVSS.n18555 1.89035
R39549 DVSS.n18995 DVSS.n18612 1.89035
R39550 DVSS.n18997 DVSS.n18554 1.89035
R39551 DVSS.n18995 DVSS.n18611 1.89035
R39552 DVSS.n18997 DVSS.n18553 1.89035
R39553 DVSS.n18995 DVSS.n18610 1.89035
R39554 DVSS.n18997 DVSS.n18552 1.89035
R39555 DVSS.n18995 DVSS.n18609 1.89035
R39556 DVSS.n18997 DVSS.n18551 1.89035
R39557 DVSS.n18995 DVSS.n18608 1.89035
R39558 DVSS.n18997 DVSS.n18550 1.89035
R39559 DVSS.n18995 DVSS.n18607 1.89035
R39560 DVSS.n18997 DVSS.n18549 1.89035
R39561 DVSS.n18995 DVSS.n18606 1.89035
R39562 DVSS.n18997 DVSS.n18548 1.89035
R39563 DVSS.n18995 DVSS.n18605 1.89035
R39564 DVSS.n18997 DVSS.n18547 1.89035
R39565 DVSS.n18995 DVSS.n18604 1.89035
R39566 DVSS.n18997 DVSS.n18546 1.89035
R39567 DVSS.n18995 DVSS.n18603 1.89035
R39568 DVSS.n18997 DVSS.n18545 1.89035
R39569 DVSS.n18995 DVSS.n18602 1.89035
R39570 DVSS.n18997 DVSS.n18544 1.89035
R39571 DVSS.n18995 DVSS.n18601 1.89035
R39572 DVSS.n18997 DVSS.n18543 1.89035
R39573 DVSS.n18995 DVSS.n18600 1.89035
R39574 DVSS.n18997 DVSS.n18542 1.89035
R39575 DVSS.n18995 DVSS.n18599 1.89035
R39576 DVSS.n18997 DVSS.n18541 1.89035
R39577 DVSS.n18995 DVSS.n18598 1.89035
R39578 DVSS.n18997 DVSS.n18540 1.89035
R39579 DVSS.n18995 DVSS.n18597 1.89035
R39580 DVSS.n18997 DVSS.n18539 1.89035
R39581 DVSS.n18995 DVSS.n18596 1.89035
R39582 DVSS.n18997 DVSS.n18538 1.89035
R39583 DVSS.n18995 DVSS.n18595 1.89035
R39584 DVSS.n18997 DVSS.n18537 1.89035
R39585 DVSS.n18995 DVSS.n18594 1.89035
R39586 DVSS.n18997 DVSS.n18536 1.89035
R39587 DVSS.n18995 DVSS.n18593 1.89035
R39588 DVSS.n18997 DVSS.n18535 1.89035
R39589 DVSS.n18995 DVSS.n18592 1.89035
R39590 DVSS.n18997 DVSS.n18534 1.89035
R39591 DVSS.n18995 DVSS.n18591 1.89035
R39592 DVSS.n18997 DVSS.n18533 1.89035
R39593 DVSS.n18995 DVSS.n18590 1.89035
R39594 DVSS.n18997 DVSS.n18532 1.89035
R39595 DVSS.n18995 DVSS.n18589 1.89035
R39596 DVSS.n18997 DVSS.n18531 1.89035
R39597 DVSS.n18995 DVSS.n18588 1.89035
R39598 DVSS.n18647 DVSS.n18646 1.89035
R39599 DVSS.n20474 DVSS.n14738 1.89035
R39600 DVSS.n14842 DVSS.n14705 1.89035
R39601 DVSS.n20474 DVSS.n14737 1.89035
R39602 DVSS.n14837 DVSS.n14705 1.89035
R39603 DVSS.n20474 DVSS.n14736 1.89035
R39604 DVSS.n14832 DVSS.n14705 1.89035
R39605 DVSS.n20474 DVSS.n14735 1.89035
R39606 DVSS.n14827 DVSS.n14705 1.89035
R39607 DVSS.n20474 DVSS.n14734 1.89035
R39608 DVSS.n14822 DVSS.n14705 1.89035
R39609 DVSS.n20474 DVSS.n14733 1.89035
R39610 DVSS.n14817 DVSS.n14705 1.89035
R39611 DVSS.n20474 DVSS.n14732 1.89035
R39612 DVSS.n14812 DVSS.n14705 1.89035
R39613 DVSS.n20474 DVSS.n14731 1.89035
R39614 DVSS.n14807 DVSS.n14705 1.89035
R39615 DVSS.n20474 DVSS.n14730 1.89035
R39616 DVSS.n14802 DVSS.n14705 1.89035
R39617 DVSS.n20474 DVSS.n14729 1.89035
R39618 DVSS.n14797 DVSS.n14705 1.89035
R39619 DVSS.n20474 DVSS.n14728 1.89035
R39620 DVSS.n14792 DVSS.n14705 1.89035
R39621 DVSS.n20474 DVSS.n14727 1.89035
R39622 DVSS.n14787 DVSS.n14705 1.89035
R39623 DVSS.n20474 DVSS.n14726 1.89035
R39624 DVSS.n14782 DVSS.n14705 1.89035
R39625 DVSS.n20474 DVSS.n14725 1.89035
R39626 DVSS.n14777 DVSS.n14705 1.89035
R39627 DVSS.n20474 DVSS.n14724 1.89035
R39628 DVSS.n14772 DVSS.n14705 1.89035
R39629 DVSS.n20474 DVSS.n14723 1.89035
R39630 DVSS.n14767 DVSS.n14705 1.89035
R39631 DVSS.n20474 DVSS.n14722 1.89035
R39632 DVSS.n14762 DVSS.n14705 1.89035
R39633 DVSS.n20474 DVSS.n14721 1.89035
R39634 DVSS.n14757 DVSS.n14705 1.89035
R39635 DVSS.n20474 DVSS.n14720 1.89035
R39636 DVSS.n14752 DVSS.n14705 1.89035
R39637 DVSS.n20474 DVSS.n14719 1.89035
R39638 DVSS.n14747 DVSS.n14705 1.89035
R39639 DVSS.n20474 DVSS.n14718 1.89035
R39640 DVSS.n14742 DVSS.n14705 1.89035
R39641 DVSS.n20474 DVSS.n14717 1.89035
R39642 DVSS.n20471 DVSS.n20470 1.89035
R39643 DVSS.n20474 DVSS.n14716 1.89035
R39644 DVSS.n20474 DVSS.n20473 1.89035
R39645 DVSS.n20471 DVSS.n14715 1.89035
R39646 DVSS.n20610 DVSS.n20474 1.89035
R39647 DVSS.n20608 DVSS.n14705 1.89035
R39648 DVSS.n20475 DVSS.n20474 1.89035
R39649 DVSS.n20603 DVSS.n14705 1.89035
R39650 DVSS.n20601 DVSS.n20474 1.89035
R39651 DVSS.n20477 DVSS.n14705 1.89035
R39652 DVSS.n20596 DVSS.n20474 1.89035
R39653 DVSS.n20594 DVSS.n14705 1.89035
R39654 DVSS.n20479 DVSS.n20474 1.89035
R39655 DVSS.n20589 DVSS.n14705 1.89035
R39656 DVSS.n20587 DVSS.n20474 1.89035
R39657 DVSS.n20481 DVSS.n14705 1.89035
R39658 DVSS.n20582 DVSS.n20474 1.89035
R39659 DVSS.n20580 DVSS.n14705 1.89035
R39660 DVSS.n20483 DVSS.n20474 1.89035
R39661 DVSS.n20575 DVSS.n14705 1.89035
R39662 DVSS.n20573 DVSS.n20474 1.89035
R39663 DVSS.n20485 DVSS.n14705 1.89035
R39664 DVSS.n20568 DVSS.n20474 1.89035
R39665 DVSS.n20566 DVSS.n14705 1.89035
R39666 DVSS.n20487 DVSS.n20474 1.89035
R39667 DVSS.n20561 DVSS.n14705 1.89035
R39668 DVSS.n20488 DVSS.n20474 1.89035
R39669 DVSS.n20556 DVSS.n14705 1.89035
R39670 DVSS.n20490 DVSS.n20474 1.89035
R39671 DVSS.n20551 DVSS.n14705 1.89035
R39672 DVSS.n20549 DVSS.n20474 1.89035
R39673 DVSS.n20492 DVSS.n14705 1.89035
R39674 DVSS.n20544 DVSS.n20474 1.89035
R39675 DVSS.n20542 DVSS.n14705 1.89035
R39676 DVSS.n20494 DVSS.n20474 1.89035
R39677 DVSS.n20537 DVSS.n14705 1.89035
R39678 DVSS.n20535 DVSS.n20474 1.89035
R39679 DVSS.n20496 DVSS.n14705 1.89035
R39680 DVSS.n20530 DVSS.n20474 1.89035
R39681 DVSS.n20528 DVSS.n14705 1.89035
R39682 DVSS.n20498 DVSS.n20474 1.89035
R39683 DVSS.n20523 DVSS.n14705 1.89035
R39684 DVSS.n20521 DVSS.n20474 1.89035
R39685 DVSS.n20500 DVSS.n14705 1.89035
R39686 DVSS.n20516 DVSS.n20474 1.89035
R39687 DVSS.n20514 DVSS.n14705 1.89035
R39688 DVSS.n20502 DVSS.n20474 1.89035
R39689 DVSS.n20509 DVSS.n14705 1.89035
R39690 DVSS.n13017 DVSS.n13015 1.85462
R39691 DVSS.n22377 DVSS.n22376 1.85434
R39692 DVSS.n19896 DVSS.n19895 1.85434
R39693 DVSS.n19892 DVSS.n19040 1.85434
R39694 DVSS.n19885 DVSS.n19884 1.85434
R39695 DVSS.n19883 DVSS.n19882 1.85434
R39696 DVSS.n19879 DVSS.n19047 1.85434
R39697 DVSS.n19872 DVSS.n19871 1.85434
R39698 DVSS.n19870 DVSS.n19869 1.85434
R39699 DVSS.n19866 DVSS.n19055 1.85434
R39700 DVSS.n19859 DVSS.n19858 1.85434
R39701 DVSS.n19857 DVSS.n19856 1.85434
R39702 DVSS.n19853 DVSS.n19063 1.85434
R39703 DVSS.n19588 DVSS.n19587 1.85434
R39704 DVSS.n19586 DVSS.n19585 1.85434
R39705 DVSS.n19578 DVSS.n19516 1.85434
R39706 DVSS.n19575 DVSS.n19574 1.85434
R39707 DVSS.n19573 DVSS.n19572 1.85434
R39708 DVSS.n19565 DVSS.n19525 1.85434
R39709 DVSS.n19562 DVSS.n19561 1.85434
R39710 DVSS.n19560 DVSS.n19559 1.85434
R39711 DVSS.n19552 DVSS.n19533 1.85434
R39712 DVSS.n19549 DVSS.n19548 1.85434
R39713 DVSS.n19547 DVSS.n19546 1.85434
R39714 DVSS.n664 DVSS.n663 1.85434
R39715 DVSS.n21831 DVSS.n21830 1.85434
R39716 DVSS.n21841 DVSS.n21825 1.85434
R39717 DVSS.n21845 DVSS.n21844 1.85434
R39718 DVSS.n21849 DVSS.n21848 1.85434
R39719 DVSS.n21947 DVSS.n21946 1.85434
R39720 DVSS.n21940 DVSS.n21939 1.85434
R39721 DVSS.n21918 DVSS.n21917 1.85434
R39722 DVSS.n21908 DVSS.n21907 1.85434
R39723 DVSS.n21898 DVSS.n21897 1.85434
R39724 DVSS.n21888 DVSS.n21887 1.85434
R39725 DVSS.n856 DVSS.n855 1.85434
R39726 DVSS.n848 DVSS.n847 1.85434
R39727 DVSS.n839 DVSS.n838 1.85434
R39728 DVSS.n830 DVSS.n829 1.85434
R39729 DVSS.n821 DVSS.n820 1.85434
R39730 DVSS.n22482 DVSS.n22481 1.85434
R39731 DVSS.n13043 DVSS.n13041 1.85434
R39732 DVSS.n13031 DVSS.n13029 1.85434
R39733 DVSS.n13052 DVSS.n13050 1.85434
R39734 DVSS.n19145 DVSS.n19144 1.85078
R39735 DVSS.n19890 DVSS.n19043 1.85078
R39736 DVSS.n19887 DVSS.n19046 1.85078
R39737 DVSS.n19051 DVSS.n19050 1.85078
R39738 DVSS.n19877 DVSS.n19052 1.85078
R39739 DVSS.n19874 DVSS.n19054 1.85078
R39740 DVSS.n19059 DVSS.n19058 1.85078
R39741 DVSS.n19864 DVSS.n19060 1.85078
R39742 DVSS.n19861 DVSS.n19062 1.85078
R39743 DVSS.n19067 DVSS.n19066 1.85078
R39744 DVSS.n19852 DVSS.n19068 1.85078
R39745 DVSS.n19519 DVSS.n19518 1.85078
R39746 DVSS.n19583 DVSS.n19517 1.85078
R39747 DVSS.n19580 DVSS.n19522 1.85078
R39748 DVSS.n19527 DVSS.n19526 1.85078
R39749 DVSS.n19570 DVSS.n19528 1.85078
R39750 DVSS.n19567 DVSS.n19530 1.85078
R39751 DVSS.n19535 DVSS.n19534 1.85078
R39752 DVSS.n19557 DVSS.n19536 1.85078
R39753 DVSS.n19554 DVSS.n19538 1.85078
R39754 DVSS.n19542 DVSS.n19541 1.85078
R39755 DVSS.n19545 DVSS.n19543 1.85078
R39756 DVSS.n661 DVSS.n659 1.85078
R39757 DVSS.n21833 DVSS.n21829 1.85078
R39758 DVSS.n21839 DVSS.n21828 1.85078
R39759 DVSS.n21836 DVSS.n21835 1.85078
R39760 DVSS.n21846 DVSS.n21799 1.85078
R39761 DVSS.n21950 DVSS.n21949 1.85078
R39762 DVSS.n21936 DVSS.n21934 1.85078
R39763 DVSS.n21914 DVSS.n21912 1.85078
R39764 DVSS.n21904 DVSS.n21902 1.85078
R39765 DVSS.n21894 DVSS.n21892 1.85078
R39766 DVSS.n21885 DVSS.n21883 1.85078
R39767 DVSS.n853 DVSS.n851 1.85078
R39768 DVSS.n844 DVSS.n842 1.85078
R39769 DVSS.n835 DVSS.n833 1.85078
R39770 DVSS.n826 DVSS.n824 1.85078
R39771 DVSS.n817 DVSS.n815 1.85078
R39772 DVSS.n22479 DVSS.n101 1.85078
R39773 DVSS.n13045 DVSS.n13040 1.85078
R39774 DVSS.n13033 DVSS.n13028 1.85078
R39775 DVSS.n13054 DVSS.n13049 1.85078
R39776 DVSS.n13019 DVSS.n13014 1.85078
R39777 DVSS.n13059 DVSS.n13058 1.85043
R39778 DVSS.n18157 DVSS.n18156 1.84325
R39779 DVSS.n16492 DVSS.n15542 1.84325
R39780 DVSS.n19207 DVSS.n19206 1.73383
R39781 DVSS.n19206 DVSS.n19205 1.73383
R39782 DVSS.n19176 DVSS.n19175 1.73383
R39783 DVSS.n19179 DVSS.n19176 1.73383
R39784 DVSS.n19926 DVSS.n19925 1.69374
R39785 DVSS.n18517 DVSS.n18516 1.69316
R39786 DVSS.n19904 DVSS.n19903 1.69315
R39787 DVSS.n19200 DVSS.n19199 1.69315
R39788 DVSS.n16385 DVSS.n16383 1.5284
R39789 DVSS.n15718 DVSS.n15717 1.5284
R39790 DVSS.n13096 DVSS.n12776 1.52691
R39791 DVSS.n16464 DVSS.n16463 1.5185
R39792 DVSS.n15645 DVSS.n15644 1.5185
R39793 DVSS.n19215 DVSS.n19208 1.50287
R39794 DVSS.n19215 DVSS.n19172 1.5005
R39795 DVSS.n16425 DVSS.n16424 1.5005
R39796 DVSS.n16423 DVSS.n16422 1.5005
R39797 DVSS.n16421 DVSS.n16420 1.5005
R39798 DVSS.n16419 DVSS.n16418 1.5005
R39799 DVSS.n16417 DVSS.n16313 1.5005
R39800 DVSS.n16416 DVSS.n16304 1.5005
R39801 DVSS.n16415 DVSS.n16414 1.5005
R39802 DVSS.n16413 DVSS.n16376 1.5005
R39803 DVSS.n16412 DVSS.n16411 1.5005
R39804 DVSS.n16410 DVSS.n16377 1.5005
R39805 DVSS.n16409 DVSS.n16408 1.5005
R39806 DVSS.n16407 DVSS.n16378 1.5005
R39807 DVSS.n16406 DVSS.n16405 1.5005
R39808 DVSS.n16404 DVSS.n16379 1.5005
R39809 DVSS.n16402 DVSS.n16401 1.5005
R39810 DVSS.n16400 DVSS.n16380 1.5005
R39811 DVSS.n16399 DVSS.n16398 1.5005
R39812 DVSS.n16397 DVSS.n16381 1.5005
R39813 DVSS.n16396 DVSS.n16395 1.5005
R39814 DVSS.n16394 DVSS.n16382 1.5005
R39815 DVSS.n16393 DVSS.n16392 1.5005
R39816 DVSS.n16391 DVSS.n16390 1.5005
R39817 DVSS.n16389 DVSS.n16388 1.5005
R39818 DVSS.n16387 DVSS.n16386 1.5005
R39819 DVSS.n16385 DVSS.n16384 1.5005
R39820 DVSS.n16466 DVSS.n16465 1.5005
R39821 DVSS.n22428 DVSS.n22427 1.5005
R39822 DVSS.n22426 DVSS.n22425 1.5005
R39823 DVSS.n22424 DVSS.n22423 1.5005
R39824 DVSS.n22422 DVSS.n22421 1.5005
R39825 DVSS.n22420 DVSS.n22419 1.5005
R39826 DVSS.n22418 DVSS.n22417 1.5005
R39827 DVSS.n22416 DVSS.n22415 1.5005
R39828 DVSS.n22414 DVSS.n22413 1.5005
R39829 DVSS.n22412 DVSS.n22411 1.5005
R39830 DVSS.n22410 DVSS.n22409 1.5005
R39831 DVSS.n22408 DVSS.n22407 1.5005
R39832 DVSS.n22406 DVSS.n22405 1.5005
R39833 DVSS.n22404 DVSS.n22403 1.5005
R39834 DVSS.n22402 DVSS.n22401 1.5005
R39835 DVSS.n22400 DVSS.n22399 1.5005
R39836 DVSS.n22398 DVSS.n22397 1.5005
R39837 DVSS.n22396 DVSS.n22395 1.5005
R39838 DVSS.n22394 DVSS.n22393 1.5005
R39839 DVSS.n22392 DVSS.n22391 1.5005
R39840 DVSS.n22390 DVSS.n22389 1.5005
R39841 DVSS.n22388 DVSS.n22387 1.5005
R39842 DVSS.n979 DVSS.n971 1.5005
R39843 DVSS.n22438 DVSS.n22437 1.5005
R39844 DVSS.n22440 DVSS.n22439 1.5005
R39845 DVSS.n22441 DVSS.n969 1.5005
R39846 DVSS.n22443 DVSS.n22442 1.5005
R39847 DVSS.n22445 DVSS.n22444 1.5005
R39848 DVSS.n22447 DVSS.n22446 1.5005
R39849 DVSS.n22448 DVSS.n925 1.5005
R39850 DVSS.n22450 DVSS.n22449 1.5005
R39851 DVSS.n968 DVSS.n924 1.5005
R39852 DVSS.n967 DVSS.n966 1.5005
R39853 DVSS.n965 DVSS.n964 1.5005
R39854 DVSS.n963 DVSS.n962 1.5005
R39855 DVSS.n961 DVSS.n960 1.5005
R39856 DVSS.n959 DVSS.n958 1.5005
R39857 DVSS.n957 DVSS.n956 1.5005
R39858 DVSS.n955 DVSS.n954 1.5005
R39859 DVSS.n953 DVSS.n952 1.5005
R39860 DVSS.n951 DVSS.n950 1.5005
R39861 DVSS.n949 DVSS.n948 1.5005
R39862 DVSS.n947 DVSS.n946 1.5005
R39863 DVSS.n945 DVSS.n944 1.5005
R39864 DVSS.n943 DVSS.n942 1.5005
R39865 DVSS.n941 DVSS.n940 1.5005
R39866 DVSS.n939 DVSS.n938 1.5005
R39867 DVSS.n937 DVSS.n936 1.5005
R39868 DVSS.n935 DVSS.n934 1.5005
R39869 DVSS.n933 DVSS.n932 1.5005
R39870 DVSS.n931 DVSS.n930 1.5005
R39871 DVSS.n929 DVSS.n928 1.5005
R39872 DVSS.n927 DVSS.n926 1.5005
R39873 DVSS.n889 DVSS.n880 1.5005
R39874 DVSS.n22455 DVSS.n22454 1.5005
R39875 DVSS.n881 DVSS.n879 1.5005
R39876 DVSS.n22134 DVSS.n22133 1.5005
R39877 DVSS.n22136 DVSS.n22135 1.5005
R39878 DVSS.n22138 DVSS.n22137 1.5005
R39879 DVSS.n22140 DVSS.n22139 1.5005
R39880 DVSS.n22142 DVSS.n22141 1.5005
R39881 DVSS.n22144 DVSS.n22143 1.5005
R39882 DVSS.n22146 DVSS.n22145 1.5005
R39883 DVSS.n22148 DVSS.n22147 1.5005
R39884 DVSS.n22150 DVSS.n22149 1.5005
R39885 DVSS.n22152 DVSS.n22151 1.5005
R39886 DVSS.n22154 DVSS.n22153 1.5005
R39887 DVSS.n22156 DVSS.n22155 1.5005
R39888 DVSS.n22158 DVSS.n22157 1.5005
R39889 DVSS.n22160 DVSS.n22159 1.5005
R39890 DVSS.n22162 DVSS.n22161 1.5005
R39891 DVSS.n22164 DVSS.n22163 1.5005
R39892 DVSS.n22166 DVSS.n22165 1.5005
R39893 DVSS.n22168 DVSS.n22167 1.5005
R39894 DVSS.n22170 DVSS.n22169 1.5005
R39895 DVSS.n22172 DVSS.n22171 1.5005
R39896 DVSS.n22174 DVSS.n22173 1.5005
R39897 DVSS.n22176 DVSS.n22175 1.5005
R39898 DVSS.n22178 DVSS.n22177 1.5005
R39899 DVSS.n22180 DVSS.n22179 1.5005
R39900 DVSS.n22182 DVSS.n22181 1.5005
R39901 DVSS.n22132 DVSS.n22130 1.5005
R39902 DVSS.n22131 DVSS.n1370 1.5005
R39903 DVSS.n22186 DVSS.n1362 1.5005
R39904 DVSS.n22188 DVSS.n22187 1.5005
R39905 DVSS.n22189 DVSS.n1361 1.5005
R39906 DVSS.n22191 DVSS.n22190 1.5005
R39907 DVSS.n22192 DVSS.n1360 1.5005
R39908 DVSS.n22194 DVSS.n22193 1.5005
R39909 DVSS.n22195 DVSS.n1359 1.5005
R39910 DVSS.n22197 DVSS.n22196 1.5005
R39911 DVSS.n22198 DVSS.n1358 1.5005
R39912 DVSS.n22200 DVSS.n22199 1.5005
R39913 DVSS.n22201 DVSS.n1357 1.5005
R39914 DVSS.n22203 DVSS.n22202 1.5005
R39915 DVSS.n22204 DVSS.n1356 1.5005
R39916 DVSS.n22206 DVSS.n22205 1.5005
R39917 DVSS.n22207 DVSS.n1355 1.5005
R39918 DVSS.n22209 DVSS.n22208 1.5005
R39919 DVSS.n22210 DVSS.n1354 1.5005
R39920 DVSS.n22212 DVSS.n22211 1.5005
R39921 DVSS.n22214 DVSS.n22213 1.5005
R39922 DVSS.n22216 DVSS.n22215 1.5005
R39923 DVSS.n22218 DVSS.n22217 1.5005
R39924 DVSS.n22220 DVSS.n22219 1.5005
R39925 DVSS.n22222 DVSS.n22221 1.5005
R39926 DVSS.n22224 DVSS.n22223 1.5005
R39927 DVSS.n22226 DVSS.n22225 1.5005
R39928 DVSS.n22228 DVSS.n22227 1.5005
R39929 DVSS.n22230 DVSS.n22229 1.5005
R39930 DVSS.n19420 DVSS.n1353 1.5005
R39931 DVSS.n19422 DVSS.n19421 1.5005
R39932 DVSS.n19423 DVSS.n719 1.5005
R39933 DVSS.n19424 DVSS.n712 1.5005
R39934 DVSS.n19426 DVSS.n19425 1.5005
R39935 DVSS.n19428 DVSS.n19427 1.5005
R39936 DVSS.n19429 DVSS.n19419 1.5005
R39937 DVSS.n19431 DVSS.n19430 1.5005
R39938 DVSS.n19432 DVSS.n19418 1.5005
R39939 DVSS.n19434 DVSS.n19433 1.5005
R39940 DVSS.n19435 DVSS.n19417 1.5005
R39941 DVSS.n19437 DVSS.n19436 1.5005
R39942 DVSS.n19438 DVSS.n19416 1.5005
R39943 DVSS.n19440 DVSS.n19439 1.5005
R39944 DVSS.n19441 DVSS.n19415 1.5005
R39945 DVSS.n19443 DVSS.n19442 1.5005
R39946 DVSS.n19444 DVSS.n19414 1.5005
R39947 DVSS.n19446 DVSS.n19445 1.5005
R39948 DVSS.n19447 DVSS.n19413 1.5005
R39949 DVSS.n19449 DVSS.n19448 1.5005
R39950 DVSS.n19450 DVSS.n19412 1.5005
R39951 DVSS.n19452 DVSS.n19451 1.5005
R39952 DVSS.n19453 DVSS.n19411 1.5005
R39953 DVSS.n19455 DVSS.n19454 1.5005
R39954 DVSS.n19456 DVSS.n19410 1.5005
R39955 DVSS.n19458 DVSS.n19457 1.5005
R39956 DVSS.n19459 DVSS.n19409 1.5005
R39957 DVSS.n19461 DVSS.n19460 1.5005
R39958 DVSS.n19462 DVSS.n19408 1.5005
R39959 DVSS.n19464 DVSS.n19463 1.5005
R39960 DVSS.n19465 DVSS.n19407 1.5005
R39961 DVSS.n19467 DVSS.n19466 1.5005
R39962 DVSS.n19468 DVSS.n19406 1.5005
R39963 DVSS.n19470 DVSS.n19469 1.5005
R39964 DVSS.n19471 DVSS.n19405 1.5005
R39965 DVSS.n19473 DVSS.n19472 1.5005
R39966 DVSS.n19474 DVSS.n19404 1.5005
R39967 DVSS.n19476 DVSS.n19475 1.5005
R39968 DVSS.n19477 DVSS.n19403 1.5005
R39969 DVSS.n19479 DVSS.n19478 1.5005
R39970 DVSS.n19480 DVSS.n19402 1.5005
R39971 DVSS.n19482 DVSS.n19481 1.5005
R39972 DVSS.n19483 DVSS.n19401 1.5005
R39973 DVSS.n19485 DVSS.n19484 1.5005
R39974 DVSS.n19486 DVSS.n19400 1.5005
R39975 DVSS.n19488 DVSS.n19487 1.5005
R39976 DVSS.n19489 DVSS.n19399 1.5005
R39977 DVSS.n19491 DVSS.n19490 1.5005
R39978 DVSS.n19492 DVSS.n19398 1.5005
R39979 DVSS.n19494 DVSS.n19493 1.5005
R39980 DVSS.n19495 DVSS.n19397 1.5005
R39981 DVSS.n19497 DVSS.n19496 1.5005
R39982 DVSS.n19498 DVSS.n19280 1.5005
R39983 DVSS.n19500 DVSS.n19499 1.5005
R39984 DVSS.n19396 DVSS.n19279 1.5005
R39985 DVSS.n19395 DVSS.n19394 1.5005
R39986 DVSS.n19393 DVSS.n19281 1.5005
R39987 DVSS.n19392 DVSS.n19391 1.5005
R39988 DVSS.n19390 DVSS.n19282 1.5005
R39989 DVSS.n19389 DVSS.n19388 1.5005
R39990 DVSS.n19387 DVSS.n19283 1.5005
R39991 DVSS.n19386 DVSS.n19385 1.5005
R39992 DVSS.n19384 DVSS.n19284 1.5005
R39993 DVSS.n19383 DVSS.n19382 1.5005
R39994 DVSS.n19381 DVSS.n19285 1.5005
R39995 DVSS.n19380 DVSS.n19379 1.5005
R39996 DVSS.n19378 DVSS.n19286 1.5005
R39997 DVSS.n19377 DVSS.n19376 1.5005
R39998 DVSS.n19375 DVSS.n19287 1.5005
R39999 DVSS.n19374 DVSS.n19373 1.5005
R40000 DVSS.n19372 DVSS.n19288 1.5005
R40001 DVSS.n19371 DVSS.n19370 1.5005
R40002 DVSS.n19369 DVSS.n19289 1.5005
R40003 DVSS.n19368 DVSS.n19367 1.5005
R40004 DVSS.n19366 DVSS.n19290 1.5005
R40005 DVSS.n19365 DVSS.n19364 1.5005
R40006 DVSS.n19363 DVSS.n19291 1.5005
R40007 DVSS.n19362 DVSS.n19361 1.5005
R40008 DVSS.n19360 DVSS.n19292 1.5005
R40009 DVSS.n19359 DVSS.n19358 1.5005
R40010 DVSS.n19357 DVSS.n19293 1.5005
R40011 DVSS.n19356 DVSS.n19355 1.5005
R40012 DVSS.n19354 DVSS.n19294 1.5005
R40013 DVSS.n19353 DVSS.n19352 1.5005
R40014 DVSS.n19351 DVSS.n19295 1.5005
R40015 DVSS.n19350 DVSS.n19349 1.5005
R40016 DVSS.n19348 DVSS.n19296 1.5005
R40017 DVSS.n19347 DVSS.n19346 1.5005
R40018 DVSS.n19345 DVSS.n19297 1.5005
R40019 DVSS.n19344 DVSS.n19343 1.5005
R40020 DVSS.n19342 DVSS.n19298 1.5005
R40021 DVSS.n19341 DVSS.n19340 1.5005
R40022 DVSS.n19339 DVSS.n19299 1.5005
R40023 DVSS.n19338 DVSS.n19337 1.5005
R40024 DVSS.n19336 DVSS.n19300 1.5005
R40025 DVSS.n19335 DVSS.n19334 1.5005
R40026 DVSS.n19333 DVSS.n19301 1.5005
R40027 DVSS.n19332 DVSS.n19331 1.5005
R40028 DVSS.n19330 DVSS.n19302 1.5005
R40029 DVSS.n19329 DVSS.n19328 1.5005
R40030 DVSS.n19327 DVSS.n19303 1.5005
R40031 DVSS.n19326 DVSS.n19325 1.5005
R40032 DVSS.n19324 DVSS.n19304 1.5005
R40033 DVSS.n19323 DVSS.n19322 1.5005
R40034 DVSS.n19321 DVSS.n19305 1.5005
R40035 DVSS.n19320 DVSS.n19319 1.5005
R40036 DVSS.n19318 DVSS.n19306 1.5005
R40037 DVSS.n19317 DVSS.n19316 1.5005
R40038 DVSS.n18082 DVSS.n18081 1.5005
R40039 DVSS.n15652 DVSS.n15651 1.5005
R40040 DVSS.n18075 DVSS.n18074 1.5005
R40041 DVSS.n18077 DVSS.n18076 1.5005
R40042 DVSS.n18073 DVSS.n15679 1.5005
R40043 DVSS.n18072 DVSS.n18071 1.5005
R40044 DVSS.n18070 DVSS.n15680 1.5005
R40045 DVSS.n18069 DVSS.n18068 1.5005
R40046 DVSS.n18067 DVSS.n15681 1.5005
R40047 DVSS.n18066 DVSS.n18065 1.5005
R40048 DVSS.n18064 DVSS.n15682 1.5005
R40049 DVSS.n18063 DVSS.n18062 1.5005
R40050 DVSS.n18061 DVSS.n15683 1.5005
R40051 DVSS.n18060 DVSS.n18059 1.5005
R40052 DVSS.n18058 DVSS.n18057 1.5005
R40053 DVSS.n18056 DVSS.n15685 1.5005
R40054 DVSS.n18055 DVSS.n18054 1.5005
R40055 DVSS.n18053 DVSS.n15686 1.5005
R40056 DVSS.n18052 DVSS.n18051 1.5005
R40057 DVSS.n18050 DVSS.n15687 1.5005
R40058 DVSS.n18049 DVSS.n18048 1.5005
R40059 DVSS.n15689 DVSS.n15688 1.5005
R40060 DVSS.n15713 DVSS.n15712 1.5005
R40061 DVSS.n15715 DVSS.n15714 1.5005
R40062 DVSS.n15717 DVSS.n15716 1.5005
R40063 DVSS.n18084 DVSS.n18083 1.5005
R40064 DVSS.n13097 DVSS.n13096 1.5005
R40065 DVSS.n12923 DVSS.n12819 1.5005
R40066 DVSS.n12922 DVSS.n12921 1.5005
R40067 DVSS.n12920 DVSS.n12919 1.5005
R40068 DVSS.n12918 DVSS.n12917 1.5005
R40069 DVSS.n12916 DVSS.n12915 1.5005
R40070 DVSS.n12914 DVSS.n12913 1.5005
R40071 DVSS.n12912 DVSS.n12911 1.5005
R40072 DVSS.n12910 DVSS.n12909 1.5005
R40073 DVSS.n12908 DVSS.n12907 1.5005
R40074 DVSS.n12906 DVSS.n12905 1.5005
R40075 DVSS.n12904 DVSS.n12903 1.5005
R40076 DVSS.n12902 DVSS.n12901 1.5005
R40077 DVSS.n12900 DVSS.n12899 1.5005
R40078 DVSS.n12898 DVSS.n12897 1.5005
R40079 DVSS.n12896 DVSS.n12895 1.5005
R40080 DVSS.n12894 DVSS.n12893 1.5005
R40081 DVSS.n12892 DVSS.n12891 1.5005
R40082 DVSS.n12890 DVSS.n12889 1.5005
R40083 DVSS.n12888 DVSS.n12887 1.5005
R40084 DVSS.n12886 DVSS.n12885 1.5005
R40085 DVSS.n12884 DVSS.n12883 1.5005
R40086 DVSS.n12882 DVSS.n12881 1.5005
R40087 DVSS.n12880 DVSS.n12879 1.5005
R40088 DVSS.n12878 DVSS.n12877 1.5005
R40089 DVSS.n12876 DVSS.n12875 1.5005
R40090 DVSS.n12874 DVSS.n12873 1.5005
R40091 DVSS.n12872 DVSS.n36 1.5005
R40092 DVSS.n12871 DVSS.n28 1.5005
R40093 DVSS.n12870 DVSS.n12869 1.5005
R40094 DVSS.n12868 DVSS.n12867 1.5005
R40095 DVSS.n12866 DVSS.n12865 1.5005
R40096 DVSS.n12864 DVSS.n12863 1.5005
R40097 DVSS.n12862 DVSS.n12861 1.5005
R40098 DVSS.n12860 DVSS.n12859 1.5005
R40099 DVSS.n12858 DVSS.n12857 1.5005
R40100 DVSS.n12856 DVSS.n12855 1.5005
R40101 DVSS.n12854 DVSS.n12853 1.5005
R40102 DVSS.n12852 DVSS.n12851 1.5005
R40103 DVSS.n12850 DVSS.n12849 1.5005
R40104 DVSS.n12848 DVSS.n12847 1.5005
R40105 DVSS.n12846 DVSS.n12845 1.5005
R40106 DVSS.n12844 DVSS.n12843 1.5005
R40107 DVSS.n12842 DVSS.n12841 1.5005
R40108 DVSS.n12840 DVSS.n12839 1.5005
R40109 DVSS.n12838 DVSS.n12837 1.5005
R40110 DVSS.n12836 DVSS.n12835 1.5005
R40111 DVSS.n12834 DVSS.n12833 1.5005
R40112 DVSS.n12832 DVSS.n12831 1.5005
R40113 DVSS.n12830 DVSS.n12829 1.5005
R40114 DVSS.n12828 DVSS.n12827 1.5005
R40115 DVSS.n12826 DVSS.n12825 1.5005
R40116 DVSS.n12824 DVSS.n12823 1.5005
R40117 DVSS.n12822 DVSS.n12821 1.5005
R40118 DVSS.n12820 DVSS.n1220 1.5005
R40119 DVSS.n22333 DVSS.n22332 1.5005
R40120 DVSS.n22331 DVSS.n1219 1.5005
R40121 DVSS.n22330 DVSS.n22329 1.5005
R40122 DVSS.n22328 DVSS.n22327 1.5005
R40123 DVSS.n1223 DVSS.n1222 1.5005
R40124 DVSS.n22323 DVSS.n22322 1.5005
R40125 DVSS.n22321 DVSS.n22320 1.5005
R40126 DVSS.n22319 DVSS.n22318 1.5005
R40127 DVSS.n22317 DVSS.n22316 1.5005
R40128 DVSS.n22315 DVSS.n22314 1.5005
R40129 DVSS.n22313 DVSS.n22312 1.5005
R40130 DVSS.n22311 DVSS.n22310 1.5005
R40131 DVSS.n22309 DVSS.n22308 1.5005
R40132 DVSS.n22307 DVSS.n22306 1.5005
R40133 DVSS.n22305 DVSS.n22304 1.5005
R40134 DVSS.n22303 DVSS.n22302 1.5005
R40135 DVSS.n22301 DVSS.n22300 1.5005
R40136 DVSS.n22299 DVSS.n22298 1.5005
R40137 DVSS.n22297 DVSS.n22296 1.5005
R40138 DVSS.n22295 DVSS.n22294 1.5005
R40139 DVSS.n22293 DVSS.n22292 1.5005
R40140 DVSS.n22291 DVSS.n22290 1.5005
R40141 DVSS.n22289 DVSS.n22288 1.5005
R40142 DVSS.n22287 DVSS.n22286 1.5005
R40143 DVSS.n22285 DVSS.n22284 1.5005
R40144 DVSS.n22283 DVSS.n22282 1.5005
R40145 DVSS.n22281 DVSS.n22280 1.5005
R40146 DVSS.n22279 DVSS.n22278 1.5005
R40147 DVSS.n22277 DVSS.n22276 1.5005
R40148 DVSS.n22275 DVSS.n22274 1.5005
R40149 DVSS.n22273 DVSS.n1263 1.5005
R40150 DVSS.n22272 DVSS.n22271 1.5005
R40151 DVSS.n22270 DVSS.n1264 1.5005
R40152 DVSS.n22269 DVSS.n22268 1.5005
R40153 DVSS.n22267 DVSS.n1265 1.5005
R40154 DVSS.n22266 DVSS.n22265 1.5005
R40155 DVSS.n22264 DVSS.n1266 1.5005
R40156 DVSS.n22263 DVSS.n22262 1.5005
R40157 DVSS.n22261 DVSS.n1267 1.5005
R40158 DVSS.n22260 DVSS.n22259 1.5005
R40159 DVSS.n22258 DVSS.n1268 1.5005
R40160 DVSS.n22257 DVSS.n22256 1.5005
R40161 DVSS.n22255 DVSS.n1269 1.5005
R40162 DVSS.n22254 DVSS.n22253 1.5005
R40163 DVSS.n22252 DVSS.n1270 1.5005
R40164 DVSS.n22251 DVSS.n22250 1.5005
R40165 DVSS.n22249 DVSS.n476 1.5005
R40166 DVSS.n22248 DVSS.n469 1.5005
R40167 DVSS.n22247 DVSS.n22246 1.5005
R40168 DVSS.n22245 DVSS.n22244 1.5005
R40169 DVSS.n22243 DVSS.n22242 1.5005
R40170 DVSS.n22241 DVSS.n22240 1.5005
R40171 DVSS.n22239 DVSS.n22238 1.5005
R40172 DVSS.n22237 DVSS.n22236 1.5005
R40173 DVSS.n22235 DVSS.n22234 1.5005
R40174 DVSS.n22233 DVSS.n22232 1.5005
R40175 DVSS.n19763 DVSS.n1272 1.5005
R40176 DVSS.n19765 DVSS.n19764 1.5005
R40177 DVSS.n19767 DVSS.n19766 1.5005
R40178 DVSS.n19769 DVSS.n19768 1.5005
R40179 DVSS.n19770 DVSS.n19762 1.5005
R40180 DVSS.n19772 DVSS.n19771 1.5005
R40181 DVSS.n19773 DVSS.n19761 1.5005
R40182 DVSS.n19775 DVSS.n19774 1.5005
R40183 DVSS.n19776 DVSS.n19760 1.5005
R40184 DVSS.n19778 DVSS.n19777 1.5005
R40185 DVSS.n19779 DVSS.n19759 1.5005
R40186 DVSS.n19781 DVSS.n19780 1.5005
R40187 DVSS.n19782 DVSS.n19758 1.5005
R40188 DVSS.n19784 DVSS.n19783 1.5005
R40189 DVSS.n19785 DVSS.n19757 1.5005
R40190 DVSS.n19787 DVSS.n19786 1.5005
R40191 DVSS.n19788 DVSS.n19756 1.5005
R40192 DVSS.n19790 DVSS.n19789 1.5005
R40193 DVSS.n19791 DVSS.n19755 1.5005
R40194 DVSS.n19793 DVSS.n19792 1.5005
R40195 DVSS.n19794 DVSS.n19754 1.5005
R40196 DVSS.n19796 DVSS.n19795 1.5005
R40197 DVSS.n19797 DVSS.n19753 1.5005
R40198 DVSS.n19799 DVSS.n19798 1.5005
R40199 DVSS.n19800 DVSS.n19752 1.5005
R40200 DVSS.n19802 DVSS.n19801 1.5005
R40201 DVSS.n19803 DVSS.n19751 1.5005
R40202 DVSS.n19805 DVSS.n19804 1.5005
R40203 DVSS.n19806 DVSS.n19750 1.5005
R40204 DVSS.n19808 DVSS.n19807 1.5005
R40205 DVSS.n19809 DVSS.n19749 1.5005
R40206 DVSS.n19811 DVSS.n19810 1.5005
R40207 DVSS.n19812 DVSS.n19748 1.5005
R40208 DVSS.n19814 DVSS.n19813 1.5005
R40209 DVSS.n19815 DVSS.n19747 1.5005
R40210 DVSS.n19817 DVSS.n19816 1.5005
R40211 DVSS.n19818 DVSS.n19746 1.5005
R40212 DVSS.n19820 DVSS.n19819 1.5005
R40213 DVSS.n19821 DVSS.n19745 1.5005
R40214 DVSS.n19823 DVSS.n19822 1.5005
R40215 DVSS.n19824 DVSS.n19744 1.5005
R40216 DVSS.n19826 DVSS.n19825 1.5005
R40217 DVSS.n19827 DVSS.n19743 1.5005
R40218 DVSS.n19829 DVSS.n19828 1.5005
R40219 DVSS.n19830 DVSS.n19742 1.5005
R40220 DVSS.n19832 DVSS.n19831 1.5005
R40221 DVSS.n19833 DVSS.n19741 1.5005
R40222 DVSS.n19835 DVSS.n19834 1.5005
R40223 DVSS.n19836 DVSS.n19740 1.5005
R40224 DVSS.n19838 DVSS.n19837 1.5005
R40225 DVSS.n19839 DVSS.n19739 1.5005
R40226 DVSS.n19841 DVSS.n19840 1.5005
R40227 DVSS.n19842 DVSS.n19111 1.5005
R40228 DVSS.n19844 DVSS.n19843 1.5005
R40229 DVSS.n19738 DVSS.n19110 1.5005
R40230 DVSS.n19737 DVSS.n19736 1.5005
R40231 DVSS.n19735 DVSS.n19112 1.5005
R40232 DVSS.n19734 DVSS.n19733 1.5005
R40233 DVSS.n19732 DVSS.n19113 1.5005
R40234 DVSS.n19731 DVSS.n19730 1.5005
R40235 DVSS.n19729 DVSS.n19114 1.5005
R40236 DVSS.n19728 DVSS.n19727 1.5005
R40237 DVSS.n19726 DVSS.n19115 1.5005
R40238 DVSS.n19725 DVSS.n19724 1.5005
R40239 DVSS.n19723 DVSS.n19116 1.5005
R40240 DVSS.n19722 DVSS.n19721 1.5005
R40241 DVSS.n19720 DVSS.n19117 1.5005
R40242 DVSS.n19719 DVSS.n19718 1.5005
R40243 DVSS.n19717 DVSS.n19118 1.5005
R40244 DVSS.n19716 DVSS.n19715 1.5005
R40245 DVSS.n19714 DVSS.n19119 1.5005
R40246 DVSS.n19713 DVSS.n19712 1.5005
R40247 DVSS.n19711 DVSS.n19120 1.5005
R40248 DVSS.n19710 DVSS.n19709 1.5005
R40249 DVSS.n19708 DVSS.n19121 1.5005
R40250 DVSS.n19707 DVSS.n19706 1.5005
R40251 DVSS.n19705 DVSS.n19122 1.5005
R40252 DVSS.n19704 DVSS.n19703 1.5005
R40253 DVSS.n19702 DVSS.n19123 1.5005
R40254 DVSS.n19701 DVSS.n19700 1.5005
R40255 DVSS.n19699 DVSS.n19124 1.5005
R40256 DVSS.n19698 DVSS.n19697 1.5005
R40257 DVSS.n19696 DVSS.n19125 1.5005
R40258 DVSS.n19695 DVSS.n19694 1.5005
R40259 DVSS.n19693 DVSS.n19126 1.5005
R40260 DVSS.n19692 DVSS.n19691 1.5005
R40261 DVSS.n19690 DVSS.n19127 1.5005
R40262 DVSS.n19689 DVSS.n19688 1.5005
R40263 DVSS.n19687 DVSS.n19128 1.5005
R40264 DVSS.n19686 DVSS.n19685 1.5005
R40265 DVSS.n19684 DVSS.n19129 1.5005
R40266 DVSS.n19683 DVSS.n19682 1.5005
R40267 DVSS.n19681 DVSS.n19130 1.5005
R40268 DVSS.n19680 DVSS.n19679 1.5005
R40269 DVSS.n19678 DVSS.n19131 1.5005
R40270 DVSS.n19677 DVSS.n19676 1.5005
R40271 DVSS.n19675 DVSS.n19132 1.5005
R40272 DVSS.n19674 DVSS.n19673 1.5005
R40273 DVSS.n19672 DVSS.n19133 1.5005
R40274 DVSS.n19671 DVSS.n19670 1.5005
R40275 DVSS.n19669 DVSS.n19134 1.5005
R40276 DVSS.n19668 DVSS.n19667 1.5005
R40277 DVSS.n19666 DVSS.n19135 1.5005
R40278 DVSS.n19665 DVSS.n19664 1.5005
R40279 DVSS.n19663 DVSS.n19136 1.5005
R40280 DVSS.n19662 DVSS.n19661 1.5005
R40281 DVSS.n19660 DVSS.n19137 1.5005
R40282 DVSS.n19659 DVSS.n19658 1.5005
R40283 DVSS.n19191 DVSS.n19190 1.46805
R40284 DVSS.n21162 DVSS.n21161 1.45763
R40285 DVSS.n20473 DVSS.n14710 1.42229
R40286 DVSS.n20611 DVSS.n14715 1.42229
R40287 DVSS.n20610 DVSS.n20609 1.42229
R40288 DVSS.n20609 DVSS.n20608 1.42229
R40289 DVSS.n20604 DVSS.n20475 1.42229
R40290 DVSS.n20604 DVSS.n20603 1.42229
R40291 DVSS.n20601 DVSS.n20600 1.42229
R40292 DVSS.n20600 DVSS.n20477 1.42229
R40293 DVSS.n20596 DVSS.n20595 1.42229
R40294 DVSS.n20595 DVSS.n20594 1.42229
R40295 DVSS.n20590 DVSS.n20479 1.42229
R40296 DVSS.n20590 DVSS.n20589 1.42229
R40297 DVSS.n20587 DVSS.n20586 1.42229
R40298 DVSS.n20586 DVSS.n20481 1.42229
R40299 DVSS.n20582 DVSS.n20581 1.42229
R40300 DVSS.n20581 DVSS.n20580 1.42229
R40301 DVSS.n20576 DVSS.n20483 1.42229
R40302 DVSS.n20576 DVSS.n20575 1.42229
R40303 DVSS.n20573 DVSS.n20572 1.42229
R40304 DVSS.n20572 DVSS.n20485 1.42229
R40305 DVSS.n20568 DVSS.n20567 1.42229
R40306 DVSS.n20567 DVSS.n20566 1.42229
R40307 DVSS.n20562 DVSS.n20487 1.42229
R40308 DVSS.n20562 DVSS.n20561 1.42229
R40309 DVSS.n20557 DVSS.n20488 1.42229
R40310 DVSS.n20557 DVSS.n20556 1.42229
R40311 DVSS.n20552 DVSS.n20490 1.42229
R40312 DVSS.n20552 DVSS.n20551 1.42229
R40313 DVSS.n20549 DVSS.n20548 1.42229
R40314 DVSS.n20548 DVSS.n20492 1.42229
R40315 DVSS.n20544 DVSS.n20543 1.42229
R40316 DVSS.n20543 DVSS.n20542 1.42229
R40317 DVSS.n20538 DVSS.n20494 1.42229
R40318 DVSS.n20538 DVSS.n20537 1.42229
R40319 DVSS.n20535 DVSS.n20534 1.42229
R40320 DVSS.n20534 DVSS.n20496 1.42229
R40321 DVSS.n20530 DVSS.n20529 1.42229
R40322 DVSS.n20529 DVSS.n20528 1.42229
R40323 DVSS.n20524 DVSS.n20498 1.42229
R40324 DVSS.n20524 DVSS.n20523 1.42229
R40325 DVSS.n20521 DVSS.n20520 1.42229
R40326 DVSS.n20520 DVSS.n20500 1.42229
R40327 DVSS.n20516 DVSS.n20515 1.42229
R40328 DVSS.n20515 DVSS.n20514 1.42229
R40329 DVSS.n20510 DVSS.n20502 1.42229
R40330 DVSS.n20510 DVSS.n20509 1.42229
R40331 DVSS.n14843 DVSS.n14738 1.42229
R40332 DVSS.n14843 DVSS.n14842 1.42229
R40333 DVSS.n14838 DVSS.n14737 1.42229
R40334 DVSS.n14838 DVSS.n14837 1.42229
R40335 DVSS.n14833 DVSS.n14736 1.42229
R40336 DVSS.n14833 DVSS.n14832 1.42229
R40337 DVSS.n14828 DVSS.n14735 1.42229
R40338 DVSS.n14828 DVSS.n14827 1.42229
R40339 DVSS.n14823 DVSS.n14734 1.42229
R40340 DVSS.n14823 DVSS.n14822 1.42229
R40341 DVSS.n14818 DVSS.n14733 1.42229
R40342 DVSS.n14818 DVSS.n14817 1.42229
R40343 DVSS.n14813 DVSS.n14732 1.42229
R40344 DVSS.n14813 DVSS.n14812 1.42229
R40345 DVSS.n14808 DVSS.n14731 1.42229
R40346 DVSS.n14808 DVSS.n14807 1.42229
R40347 DVSS.n14803 DVSS.n14730 1.42229
R40348 DVSS.n14803 DVSS.n14802 1.42229
R40349 DVSS.n14798 DVSS.n14729 1.42229
R40350 DVSS.n14798 DVSS.n14797 1.42229
R40351 DVSS.n14793 DVSS.n14728 1.42229
R40352 DVSS.n14793 DVSS.n14792 1.42229
R40353 DVSS.n14788 DVSS.n14727 1.42229
R40354 DVSS.n14788 DVSS.n14787 1.42229
R40355 DVSS.n14783 DVSS.n14726 1.42229
R40356 DVSS.n14783 DVSS.n14782 1.42229
R40357 DVSS.n14778 DVSS.n14725 1.42229
R40358 DVSS.n14778 DVSS.n14777 1.42229
R40359 DVSS.n14773 DVSS.n14724 1.42229
R40360 DVSS.n14773 DVSS.n14772 1.42229
R40361 DVSS.n14768 DVSS.n14723 1.42229
R40362 DVSS.n14768 DVSS.n14767 1.42229
R40363 DVSS.n14763 DVSS.n14722 1.42229
R40364 DVSS.n14763 DVSS.n14762 1.42229
R40365 DVSS.n14758 DVSS.n14721 1.42229
R40366 DVSS.n14758 DVSS.n14757 1.42229
R40367 DVSS.n14753 DVSS.n14720 1.42229
R40368 DVSS.n14753 DVSS.n14752 1.42229
R40369 DVSS.n14748 DVSS.n14719 1.42229
R40370 DVSS.n14748 DVSS.n14747 1.42229
R40371 DVSS.n14743 DVSS.n14718 1.42229
R40372 DVSS.n14743 DVSS.n14742 1.42229
R40373 DVSS.n14717 DVSS.n14712 1.42229
R40374 DVSS.n20470 DVSS.n14711 1.42229
R40375 DVSS.n20468 DVSS.n14716 1.42229
R40376 DVSS.n18763 DVSS.n18583 1.42229
R40377 DVSS.n18770 DVSS.n18640 1.42229
R40378 DVSS.n18770 DVSS.n18582 1.42229
R40379 DVSS.n18774 DVSS.n18639 1.42229
R40380 DVSS.n18774 DVSS.n18581 1.42229
R40381 DVSS.n18778 DVSS.n18638 1.42229
R40382 DVSS.n18778 DVSS.n18580 1.42229
R40383 DVSS.n18782 DVSS.n18637 1.42229
R40384 DVSS.n18782 DVSS.n18579 1.42229
R40385 DVSS.n18786 DVSS.n18636 1.42229
R40386 DVSS.n18786 DVSS.n18578 1.42229
R40387 DVSS.n18790 DVSS.n18635 1.42229
R40388 DVSS.n18790 DVSS.n18577 1.42229
R40389 DVSS.n18794 DVSS.n18634 1.42229
R40390 DVSS.n18794 DVSS.n18576 1.42229
R40391 DVSS.n18798 DVSS.n18633 1.42229
R40392 DVSS.n18798 DVSS.n18575 1.42229
R40393 DVSS.n18802 DVSS.n18632 1.42229
R40394 DVSS.n18802 DVSS.n18574 1.42229
R40395 DVSS.n18806 DVSS.n18631 1.42229
R40396 DVSS.n18806 DVSS.n18573 1.42229
R40397 DVSS.n18810 DVSS.n18630 1.42229
R40398 DVSS.n18810 DVSS.n18572 1.42229
R40399 DVSS.n18814 DVSS.n18629 1.42229
R40400 DVSS.n18814 DVSS.n18571 1.42229
R40401 DVSS.n18818 DVSS.n18628 1.42229
R40402 DVSS.n18818 DVSS.n18570 1.42229
R40403 DVSS.n18823 DVSS.n18627 1.42229
R40404 DVSS.n18823 DVSS.n18569 1.42229
R40405 DVSS.n18827 DVSS.n18626 1.42229
R40406 DVSS.n18827 DVSS.n18568 1.42229
R40407 DVSS.n18831 DVSS.n18625 1.42229
R40408 DVSS.n18831 DVSS.n18567 1.42229
R40409 DVSS.n18835 DVSS.n18624 1.42229
R40410 DVSS.n18835 DVSS.n18566 1.42229
R40411 DVSS.n18839 DVSS.n18623 1.42229
R40412 DVSS.n18839 DVSS.n18565 1.42229
R40413 DVSS.n18843 DVSS.n18622 1.42229
R40414 DVSS.n18843 DVSS.n18564 1.42229
R40415 DVSS.n18847 DVSS.n18621 1.42229
R40416 DVSS.n18847 DVSS.n18563 1.42229
R40417 DVSS.n18851 DVSS.n18620 1.42229
R40418 DVSS.n18851 DVSS.n18562 1.42229
R40419 DVSS.n18855 DVSS.n18619 1.42229
R40420 DVSS.n18855 DVSS.n18561 1.42229
R40421 DVSS.n18859 DVSS.n18618 1.42229
R40422 DVSS.n18859 DVSS.n18560 1.42229
R40423 DVSS.n18863 DVSS.n18617 1.42229
R40424 DVSS.n18863 DVSS.n18559 1.42229
R40425 DVSS.n18616 DVSS.n18558 1.42229
R40426 DVSS.n18760 DVSS.n18584 1.42229
R40427 DVSS.n18615 DVSS.n18557 1.42229
R40428 DVSS.n18759 DVSS.n18585 1.42229
R40429 DVSS.n18614 DVSS.n18556 1.42229
R40430 DVSS.n18758 DVSS.n18586 1.42229
R40431 DVSS.n18756 DVSS.n18613 1.42229
R40432 DVSS.n18756 DVSS.n18555 1.42229
R40433 DVSS.n18751 DVSS.n18612 1.42229
R40434 DVSS.n18751 DVSS.n18554 1.42229
R40435 DVSS.n18747 DVSS.n18611 1.42229
R40436 DVSS.n18747 DVSS.n18553 1.42229
R40437 DVSS.n18743 DVSS.n18610 1.42229
R40438 DVSS.n18743 DVSS.n18552 1.42229
R40439 DVSS.n18739 DVSS.n18609 1.42229
R40440 DVSS.n18739 DVSS.n18551 1.42229
R40441 DVSS.n18735 DVSS.n18608 1.42229
R40442 DVSS.n18735 DVSS.n18550 1.42229
R40443 DVSS.n18731 DVSS.n18607 1.42229
R40444 DVSS.n18731 DVSS.n18549 1.42229
R40445 DVSS.n18727 DVSS.n18606 1.42229
R40446 DVSS.n18727 DVSS.n18548 1.42229
R40447 DVSS.n18723 DVSS.n18605 1.42229
R40448 DVSS.n18723 DVSS.n18547 1.42229
R40449 DVSS.n18719 DVSS.n18604 1.42229
R40450 DVSS.n18719 DVSS.n18546 1.42229
R40451 DVSS.n18715 DVSS.n18603 1.42229
R40452 DVSS.n18715 DVSS.n18545 1.42229
R40453 DVSS.n18711 DVSS.n18602 1.42229
R40454 DVSS.n18711 DVSS.n18544 1.42229
R40455 DVSS.n18706 DVSS.n18601 1.42229
R40456 DVSS.n18706 DVSS.n18543 1.42229
R40457 DVSS.n18702 DVSS.n18600 1.42229
R40458 DVSS.n18702 DVSS.n18542 1.42229
R40459 DVSS.n18698 DVSS.n18599 1.42229
R40460 DVSS.n18698 DVSS.n18541 1.42229
R40461 DVSS.n18694 DVSS.n18598 1.42229
R40462 DVSS.n18694 DVSS.n18540 1.42229
R40463 DVSS.n18690 DVSS.n18597 1.42229
R40464 DVSS.n18690 DVSS.n18539 1.42229
R40465 DVSS.n18686 DVSS.n18596 1.42229
R40466 DVSS.n18686 DVSS.n18538 1.42229
R40467 DVSS.n18682 DVSS.n18595 1.42229
R40468 DVSS.n18682 DVSS.n18537 1.42229
R40469 DVSS.n18678 DVSS.n18594 1.42229
R40470 DVSS.n18678 DVSS.n18536 1.42229
R40471 DVSS.n18674 DVSS.n18593 1.42229
R40472 DVSS.n18674 DVSS.n18535 1.42229
R40473 DVSS.n18670 DVSS.n18592 1.42229
R40474 DVSS.n18670 DVSS.n18534 1.42229
R40475 DVSS.n18666 DVSS.n18591 1.42229
R40476 DVSS.n18666 DVSS.n18533 1.42229
R40477 DVSS.n18662 DVSS.n18590 1.42229
R40478 DVSS.n18662 DVSS.n18532 1.42229
R40479 DVSS.n18658 DVSS.n18589 1.42229
R40480 DVSS.n18658 DVSS.n18531 1.42229
R40481 DVSS.n18588 DVSS.n18530 1.42229
R40482 DVSS.n18646 DVSS.n18587 1.42229
R40483 DVSS.n18641 DVSS.n18583 1.42229
R40484 DVSS.n18763 DVSS.n18640 1.42229
R40485 DVSS.n18772 DVSS.n18639 1.42229
R40486 DVSS.n18772 DVSS.n18582 1.42229
R40487 DVSS.n18776 DVSS.n18638 1.42229
R40488 DVSS.n18776 DVSS.n18581 1.42229
R40489 DVSS.n18780 DVSS.n18637 1.42229
R40490 DVSS.n18780 DVSS.n18580 1.42229
R40491 DVSS.n18784 DVSS.n18636 1.42229
R40492 DVSS.n18784 DVSS.n18579 1.42229
R40493 DVSS.n18788 DVSS.n18635 1.42229
R40494 DVSS.n18788 DVSS.n18578 1.42229
R40495 DVSS.n18792 DVSS.n18634 1.42229
R40496 DVSS.n18792 DVSS.n18577 1.42229
R40497 DVSS.n18796 DVSS.n18633 1.42229
R40498 DVSS.n18796 DVSS.n18576 1.42229
R40499 DVSS.n18800 DVSS.n18632 1.42229
R40500 DVSS.n18800 DVSS.n18575 1.42229
R40501 DVSS.n18804 DVSS.n18631 1.42229
R40502 DVSS.n18804 DVSS.n18574 1.42229
R40503 DVSS.n18808 DVSS.n18630 1.42229
R40504 DVSS.n18808 DVSS.n18573 1.42229
R40505 DVSS.n18812 DVSS.n18629 1.42229
R40506 DVSS.n18812 DVSS.n18572 1.42229
R40507 DVSS.n18816 DVSS.n18628 1.42229
R40508 DVSS.n18816 DVSS.n18571 1.42229
R40509 DVSS.n18821 DVSS.n18627 1.42229
R40510 DVSS.n18821 DVSS.n18570 1.42229
R40511 DVSS.n18825 DVSS.n18626 1.42229
R40512 DVSS.n18825 DVSS.n18569 1.42229
R40513 DVSS.n18829 DVSS.n18625 1.42229
R40514 DVSS.n18829 DVSS.n18568 1.42229
R40515 DVSS.n18833 DVSS.n18624 1.42229
R40516 DVSS.n18833 DVSS.n18567 1.42229
R40517 DVSS.n18837 DVSS.n18623 1.42229
R40518 DVSS.n18837 DVSS.n18566 1.42229
R40519 DVSS.n18841 DVSS.n18622 1.42229
R40520 DVSS.n18841 DVSS.n18565 1.42229
R40521 DVSS.n18845 DVSS.n18621 1.42229
R40522 DVSS.n18845 DVSS.n18564 1.42229
R40523 DVSS.n18849 DVSS.n18620 1.42229
R40524 DVSS.n18849 DVSS.n18563 1.42229
R40525 DVSS.n18853 DVSS.n18619 1.42229
R40526 DVSS.n18853 DVSS.n18562 1.42229
R40527 DVSS.n18857 DVSS.n18618 1.42229
R40528 DVSS.n18857 DVSS.n18561 1.42229
R40529 DVSS.n18861 DVSS.n18617 1.42229
R40530 DVSS.n18861 DVSS.n18560 1.42229
R40531 DVSS.n18865 DVSS.n18616 1.42229
R40532 DVSS.n18865 DVSS.n18559 1.42229
R40533 DVSS.n18760 DVSS.n18558 1.42229
R40534 DVSS.n18615 DVSS.n18584 1.42229
R40535 DVSS.n18759 DVSS.n18557 1.42229
R40536 DVSS.n18614 DVSS.n18585 1.42229
R40537 DVSS.n18758 DVSS.n18556 1.42229
R40538 DVSS.n18613 DVSS.n18586 1.42229
R40539 DVSS.n18753 DVSS.n18612 1.42229
R40540 DVSS.n18753 DVSS.n18555 1.42229
R40541 DVSS.n18749 DVSS.n18611 1.42229
R40542 DVSS.n18749 DVSS.n18554 1.42229
R40543 DVSS.n18745 DVSS.n18610 1.42229
R40544 DVSS.n18745 DVSS.n18553 1.42229
R40545 DVSS.n18741 DVSS.n18609 1.42229
R40546 DVSS.n18741 DVSS.n18552 1.42229
R40547 DVSS.n18737 DVSS.n18608 1.42229
R40548 DVSS.n18737 DVSS.n18551 1.42229
R40549 DVSS.n18733 DVSS.n18607 1.42229
R40550 DVSS.n18733 DVSS.n18550 1.42229
R40551 DVSS.n18729 DVSS.n18606 1.42229
R40552 DVSS.n18729 DVSS.n18549 1.42229
R40553 DVSS.n18725 DVSS.n18605 1.42229
R40554 DVSS.n18725 DVSS.n18548 1.42229
R40555 DVSS.n18721 DVSS.n18604 1.42229
R40556 DVSS.n18721 DVSS.n18547 1.42229
R40557 DVSS.n18717 DVSS.n18603 1.42229
R40558 DVSS.n18717 DVSS.n18546 1.42229
R40559 DVSS.n18713 DVSS.n18602 1.42229
R40560 DVSS.n18713 DVSS.n18545 1.42229
R40561 DVSS.n18709 DVSS.n18601 1.42229
R40562 DVSS.n18709 DVSS.n18544 1.42229
R40563 DVSS.n18704 DVSS.n18600 1.42229
R40564 DVSS.n18704 DVSS.n18543 1.42229
R40565 DVSS.n18700 DVSS.n18599 1.42229
R40566 DVSS.n18700 DVSS.n18542 1.42229
R40567 DVSS.n18696 DVSS.n18598 1.42229
R40568 DVSS.n18696 DVSS.n18541 1.42229
R40569 DVSS.n18692 DVSS.n18597 1.42229
R40570 DVSS.n18692 DVSS.n18540 1.42229
R40571 DVSS.n18688 DVSS.n18596 1.42229
R40572 DVSS.n18688 DVSS.n18539 1.42229
R40573 DVSS.n18684 DVSS.n18595 1.42229
R40574 DVSS.n18684 DVSS.n18538 1.42229
R40575 DVSS.n18680 DVSS.n18594 1.42229
R40576 DVSS.n18680 DVSS.n18537 1.42229
R40577 DVSS.n18676 DVSS.n18593 1.42229
R40578 DVSS.n18676 DVSS.n18536 1.42229
R40579 DVSS.n18672 DVSS.n18592 1.42229
R40580 DVSS.n18672 DVSS.n18535 1.42229
R40581 DVSS.n18668 DVSS.n18591 1.42229
R40582 DVSS.n18668 DVSS.n18534 1.42229
R40583 DVSS.n18664 DVSS.n18590 1.42229
R40584 DVSS.n18664 DVSS.n18533 1.42229
R40585 DVSS.n18660 DVSS.n18589 1.42229
R40586 DVSS.n18660 DVSS.n18532 1.42229
R40587 DVSS.n18656 DVSS.n18588 1.42229
R40588 DVSS.n18656 DVSS.n18531 1.42229
R40589 DVSS.n18646 DVSS.n18530 1.42229
R40590 DVSS.n14739 DVSS.n14738 1.42229
R40591 DVSS.n14841 DVSS.n14737 1.42229
R40592 DVSS.n14842 DVSS.n14841 1.42229
R40593 DVSS.n14836 DVSS.n14736 1.42229
R40594 DVSS.n14837 DVSS.n14836 1.42229
R40595 DVSS.n14831 DVSS.n14735 1.42229
R40596 DVSS.n14832 DVSS.n14831 1.42229
R40597 DVSS.n14826 DVSS.n14734 1.42229
R40598 DVSS.n14827 DVSS.n14826 1.42229
R40599 DVSS.n14821 DVSS.n14733 1.42229
R40600 DVSS.n14822 DVSS.n14821 1.42229
R40601 DVSS.n14816 DVSS.n14732 1.42229
R40602 DVSS.n14817 DVSS.n14816 1.42229
R40603 DVSS.n14811 DVSS.n14731 1.42229
R40604 DVSS.n14812 DVSS.n14811 1.42229
R40605 DVSS.n14806 DVSS.n14730 1.42229
R40606 DVSS.n14807 DVSS.n14806 1.42229
R40607 DVSS.n14801 DVSS.n14729 1.42229
R40608 DVSS.n14802 DVSS.n14801 1.42229
R40609 DVSS.n14796 DVSS.n14728 1.42229
R40610 DVSS.n14797 DVSS.n14796 1.42229
R40611 DVSS.n14791 DVSS.n14727 1.42229
R40612 DVSS.n14792 DVSS.n14791 1.42229
R40613 DVSS.n14786 DVSS.n14726 1.42229
R40614 DVSS.n14787 DVSS.n14786 1.42229
R40615 DVSS.n14781 DVSS.n14725 1.42229
R40616 DVSS.n14782 DVSS.n14781 1.42229
R40617 DVSS.n14776 DVSS.n14724 1.42229
R40618 DVSS.n14777 DVSS.n14776 1.42229
R40619 DVSS.n14771 DVSS.n14723 1.42229
R40620 DVSS.n14772 DVSS.n14771 1.42229
R40621 DVSS.n14766 DVSS.n14722 1.42229
R40622 DVSS.n14767 DVSS.n14766 1.42229
R40623 DVSS.n14761 DVSS.n14721 1.42229
R40624 DVSS.n14762 DVSS.n14761 1.42229
R40625 DVSS.n14756 DVSS.n14720 1.42229
R40626 DVSS.n14757 DVSS.n14756 1.42229
R40627 DVSS.n14751 DVSS.n14719 1.42229
R40628 DVSS.n14752 DVSS.n14751 1.42229
R40629 DVSS.n14746 DVSS.n14718 1.42229
R40630 DVSS.n14747 DVSS.n14746 1.42229
R40631 DVSS.n14741 DVSS.n14717 1.42229
R40632 DVSS.n14742 DVSS.n14741 1.42229
R40633 DVSS.n20470 DVSS.n14712 1.42229
R40634 DVSS.n14716 DVSS.n14711 1.42229
R40635 DVSS.n20473 DVSS.n14714 1.42229
R40636 DVSS.n14715 DVSS.n14710 1.42229
R40637 DVSS.n20611 DVSS.n20610 1.42229
R40638 DVSS.n20607 DVSS.n20475 1.42229
R40639 DVSS.n20608 DVSS.n20607 1.42229
R40640 DVSS.n20602 DVSS.n20601 1.42229
R40641 DVSS.n20603 DVSS.n20602 1.42229
R40642 DVSS.n20597 DVSS.n20596 1.42229
R40643 DVSS.n20597 DVSS.n20477 1.42229
R40644 DVSS.n20593 DVSS.n20479 1.42229
R40645 DVSS.n20594 DVSS.n20593 1.42229
R40646 DVSS.n20588 DVSS.n20587 1.42229
R40647 DVSS.n20589 DVSS.n20588 1.42229
R40648 DVSS.n20583 DVSS.n20582 1.42229
R40649 DVSS.n20583 DVSS.n20481 1.42229
R40650 DVSS.n20579 DVSS.n20483 1.42229
R40651 DVSS.n20580 DVSS.n20579 1.42229
R40652 DVSS.n20574 DVSS.n20573 1.42229
R40653 DVSS.n20575 DVSS.n20574 1.42229
R40654 DVSS.n20569 DVSS.n20568 1.42229
R40655 DVSS.n20569 DVSS.n20485 1.42229
R40656 DVSS.n20565 DVSS.n20487 1.42229
R40657 DVSS.n20566 DVSS.n20565 1.42229
R40658 DVSS.n20560 DVSS.n20488 1.42229
R40659 DVSS.n20561 DVSS.n20560 1.42229
R40660 DVSS.n20555 DVSS.n20490 1.42229
R40661 DVSS.n20556 DVSS.n20555 1.42229
R40662 DVSS.n20550 DVSS.n20549 1.42229
R40663 DVSS.n20551 DVSS.n20550 1.42229
R40664 DVSS.n20545 DVSS.n20544 1.42229
R40665 DVSS.n20545 DVSS.n20492 1.42229
R40666 DVSS.n20541 DVSS.n20494 1.42229
R40667 DVSS.n20542 DVSS.n20541 1.42229
R40668 DVSS.n20536 DVSS.n20535 1.42229
R40669 DVSS.n20537 DVSS.n20536 1.42229
R40670 DVSS.n20531 DVSS.n20530 1.42229
R40671 DVSS.n20531 DVSS.n20496 1.42229
R40672 DVSS.n20527 DVSS.n20498 1.42229
R40673 DVSS.n20528 DVSS.n20527 1.42229
R40674 DVSS.n20522 DVSS.n20521 1.42229
R40675 DVSS.n20523 DVSS.n20522 1.42229
R40676 DVSS.n20517 DVSS.n20516 1.42229
R40677 DVSS.n20517 DVSS.n20500 1.42229
R40678 DVSS.n20513 DVSS.n20502 1.42229
R40679 DVSS.n20514 DVSS.n20513 1.42229
R40680 DVSS.n20509 DVSS.n20508 1.42229
R40681 DVSS.n17410 DVSS.n17053 1.35477
R40682 DVSS.n16930 DVSS.n16929 1.35477
R40683 DVSS.n19199 DVSS.n19198 1.34946
R40684 DVSS.n18169 DVSS.n18168 1.29118
R40685 DVSS.n17790 DVSS.n17789 1.29118
R40686 DVSS.n13666 DVSS.n13665 1.27407
R40687 DVSS.n19190 DVSS.n19189 1.23661
R40688 DVSS.n19192 DVSS.n19188 1.23634
R40689 DVSS.n19214 DVSS.n19003 1.17447
R40690 DVSS.n15918 DVSS.n15917 1.16121
R40691 DVSS.n18165 DVSS.n18164 1.16121
R40692 DVSS.n21447 DVSS.n21446 1.16121
R40693 DVSS.n13365 DVSS.n423 1.16121
R40694 DVSS.n16495 DVSS.n16493 1.15497
R40695 DVSS.n18158 DVSS.n18157 1.1503
R40696 DVSS.n18155 DVSS.n18154 1.14603
R40697 DVSS.n16478 DVSS.n16344 1.14075
R40698 DVSS.n18111 DVSS.n18110 1.14075
R40699 DVSS.n18158 DVSS.n15542 1.13815
R40700 DVSS.n16538 DVSS.n16537 1.1255
R40701 DVSS.n16536 DVSS.n16535 1.1255
R40702 DVSS.n16534 DVSS.n16533 1.1255
R40703 DVSS.n16532 DVSS.n16531 1.1255
R40704 DVSS.n16530 DVSS.n16529 1.1255
R40705 DVSS.n16528 DVSS.n16527 1.1255
R40706 DVSS.n16526 DVSS.n16484 1.1255
R40707 DVSS.n16525 DVSS.n16524 1.1255
R40708 DVSS.n16523 DVSS.n16485 1.1255
R40709 DVSS.n16522 DVSS.n16521 1.1255
R40710 DVSS.n16520 DVSS.n16486 1.1255
R40711 DVSS.n16519 DVSS.n16518 1.1255
R40712 DVSS.n16517 DVSS.n16487 1.1255
R40713 DVSS.n16516 DVSS.n16515 1.1255
R40714 DVSS.n16514 DVSS.n16513 1.1255
R40715 DVSS.n16512 DVSS.n16489 1.1255
R40716 DVSS.n16511 DVSS.n16510 1.1255
R40717 DVSS.n16509 DVSS.n16490 1.1255
R40718 DVSS.n16508 DVSS.n16507 1.1255
R40719 DVSS.n16506 DVSS.n16491 1.1255
R40720 DVSS.n16505 DVSS.n16504 1.1255
R40721 DVSS.n16503 DVSS.n16502 1.1255
R40722 DVSS.n16501 DVSS.n16500 1.1255
R40723 DVSS.n16499 DVSS.n16498 1.1255
R40724 DVSS.n16497 DVSS.n16496 1.1255
R40725 DVSS.n16495 DVSS.n16494 1.1255
R40726 DVSS.n16540 DVSS.n16539 1.1255
R40727 DVSS.n6670 DVSS.n6669 1.1255
R40728 DVSS.n6238 DVSS.n5896 1.1255
R40729 DVSS.n6681 DVSS.n6680 1.1255
R40730 DVSS.n6688 DVSS.n6687 1.1255
R40731 DVSS.n5889 DVSS.n5876 1.1255
R40732 DVSS.n7035 DVSS.n7034 1.1255
R40733 DVSS.n5879 DVSS.n5868 1.1255
R40734 DVSS.n7044 DVSS.n7043 1.1255
R40735 DVSS.n5869 DVSS.n5577 1.1255
R40736 DVSS.n7061 DVSS.n7060 1.1255
R40737 DVSS.n5526 DVSS.n5525 1.1255
R40738 DVSS.n7068 DVSS.n7067 1.1255
R40739 DVSS.n7080 DVSS.n7079 1.1255
R40740 DVSS.n5183 DVSS.n5177 1.1255
R40741 DVSS.n7087 DVSS.n7086 1.1255
R40742 DVSS.n4885 DVSS.n4839 1.1255
R40743 DVSS.n7106 DVSS.n7105 1.1255
R40744 DVSS.n7103 DVSS.n4833 1.1255
R40745 DVSS.n7451 DVSS.n7450 1.1255
R40746 DVSS.n7461 DVSS.n4824 1.1255
R40747 DVSS.n7798 DVSS.n7797 1.1255
R40748 DVSS.n7799 DVSS.n4818 1.1255
R40749 DVSS.n7806 DVSS.n7805 1.1255
R40750 DVSS.n7816 DVSS.n4810 1.1255
R40751 DVSS.n7819 DVSS.n7818 1.1255
R40752 DVSS.n7826 DVSS.n7825 1.1255
R40753 DVSS.n4469 DVSS.n4369 1.1255
R40754 DVSS.n8092 DVSS.n8091 1.1255
R40755 DVSS.n4413 DVSS.n4363 1.1255
R40756 DVSS.n8100 DVSS.n8099 1.1255
R40757 DVSS.n8102 DVSS.n4020 1.1255
R40758 DVSS.n8113 DVSS.n8112 1.1255
R40759 DVSS.n8120 DVSS.n4015 1.1255
R40760 DVSS.n8121 DVSS.n3858 1.1255
R40761 DVSS.n8122 DVSS.n3900 1.1255
R40762 DVSS.n8126 DVSS.n3946 1.1255
R40763 DVSS.n3846 DVSS.n3845 1.1255
R40764 DVSS.n8333 DVSS.n8332 1.1255
R40765 DVSS.n8335 DVSS.n3755 1.1255
R40766 DVSS.n8589 DVSS.n3413 1.1255
R40767 DVSS.n8606 DVSS.n8605 1.1255
R40768 DVSS.n3460 DVSS.n3407 1.1255
R40769 DVSS.n8614 DVSS.n8613 1.1255
R40770 DVSS.n8615 DVSS.n3065 1.1255
R40771 DVSS.n8626 DVSS.n8625 1.1255
R40772 DVSS.n8633 DVSS.n8632 1.1255
R40773 DVSS.n8635 DVSS.n3051 1.1255
R40774 DVSS.n8980 DVSS.n8979 1.1255
R40775 DVSS.n8987 DVSS.n3046 1.1255
R40776 DVSS.n8988 DVSS.n2890 1.1255
R40777 DVSS.n8989 DVSS.n2932 1.1255
R40778 DVSS.n8993 DVSS.n2937 1.1255
R40779 DVSS.n2878 DVSS.n2877 1.1255
R40780 DVSS.n9200 DVSS.n9199 1.1255
R40781 DVSS.n9202 DVSS.n2787 1.1255
R40782 DVSS.n9456 DVSS.n2737 1.1255
R40783 DVSS.n9761 DVSS.n9760 1.1255
R40784 DVSS.n2781 DVSS.n2731 1.1255
R40785 DVSS.n9770 DVSS.n9769 1.1255
R40786 DVSS.n2729 DVSS.n2716 1.1255
R40787 DVSS.n10117 DVSS.n10116 1.1255
R40788 DVSS.n2719 DVSS.n2707 1.1255
R40789 DVSS.n10126 DVSS.n10125 1.1255
R40790 DVSS.n2709 DVSS.n2708 1.1255
R40791 DVSS.n10144 DVSS.n10143 1.1255
R40792 DVSS.n2365 DVSS.n2364 1.1255
R40793 DVSS.n10151 DVSS.n10150 1.1255
R40794 DVSS.n10168 DVSS.n10167 1.1255
R40795 DVSS.n2070 DVSS.n2020 1.1255
R40796 DVSS.n10460 DVSS.n10459 1.1255
R40797 DVSS.n2012 DVSS.n1966 1.1255
R40798 DVSS.n10479 DVSS.n10478 1.1255
R40799 DVSS.n10476 DVSS.n1962 1.1255
R40800 DVSS.n10486 DVSS.n10485 1.1255
R40801 DVSS.n10499 DVSS.n10498 1.1255
R40802 DVSS.n10496 DVSS.n1619 1.1255
R40803 DVSS.n1615 DVSS.n1523 1.1255
R40804 DVSS.n1566 DVSS.n1509 1.1255
R40805 DVSS.n13360 DVSS.n13359 1.1255
R40806 DVSS.n10765 DVSS.n1510 1.1255
R40807 DVSS.n13349 DVSS.n13348 1.1255
R40808 DVSS.n11110 DVSS.n10768 1.1255
R40809 DVSS.n13342 DVSS.n13341 1.1255
R40810 DVSS.n11615 DVSS.n11153 1.1255
R40811 DVSS.n11616 DVSS.n11198 1.1255
R40812 DVSS.n11617 DVSS.n11458 1.1255
R40813 DVSS.n13132 DVSS.n11500 1.1255
R40814 DVSS.n13131 DVSS.n11546 1.1255
R40815 DVSS.n13130 DVSS.n11622 1.1255
R40816 DVSS.n11981 DVSS.n11621 1.1255
R40817 DVSS.n13123 DVSS.n13122 1.1255
R40818 DVSS.n13121 DVSS.n11629 1.1255
R40819 DVSS.n12339 DVSS.n12338 1.1255
R40820 DVSS.n11996 DVSS.n11994 1.1255
R40821 DVSS.n13110 DVSS.n13109 1.1255
R40822 DVSS.n12748 DVSS.n11997 1.1255
R40823 DVSS.n6669 DVSS.n6668 1.1255
R40824 DVSS.n5896 DVSS.n5895 1.1255
R40825 DVSS.n6682 DVSS.n6681 1.1255
R40826 DVSS.n6687 DVSS.n6686 1.1255
R40827 DVSS.n5876 DVSS.n5874 1.1255
R40828 DVSS.n7036 DVSS.n7035 1.1255
R40829 DVSS.n5870 DVSS.n5868 1.1255
R40830 DVSS.n7043 DVSS.n7042 1.1255
R40831 DVSS.n5871 DVSS.n5869 1.1255
R40832 DVSS.n7062 DVSS.n7061 1.1255
R40833 DVSS.n5527 DVSS.n5526 1.1255
R40834 DVSS.n7067 DVSS.n7066 1.1255
R40835 DVSS.n7081 DVSS.n7080 1.1255
R40836 DVSS.n5178 DVSS.n5177 1.1255
R40837 DVSS.n7086 DVSS.n7085 1.1255
R40838 DVSS.n4839 DVSS.n4838 1.1255
R40839 DVSS.n7107 DVSS.n7106 1.1255
R40840 DVSS.n4835 DVSS.n4833 1.1255
R40841 DVSS.n7450 DVSS.n7449 1.1255
R40842 DVSS.n7445 DVSS.n4824 1.1255
R40843 DVSS.n7798 DVSS.n4823 1.1255
R40844 DVSS.n7800 DVSS.n7799 1.1255
R40845 DVSS.n7805 DVSS.n7804 1.1255
R40846 DVSS.n4810 DVSS.n4809 1.1255
R40847 DVSS.n7820 DVSS.n7819 1.1255
R40848 DVSS.n7825 DVSS.n7824 1.1255
R40849 DVSS.n4369 DVSS.n4367 1.1255
R40850 DVSS.n8093 DVSS.n8092 1.1255
R40851 DVSS.n4364 DVSS.n4363 1.1255
R40852 DVSS.n8099 DVSS.n8098 1.1255
R40853 DVSS.n4020 DVSS.n4019 1.1255
R40854 DVSS.n8114 DVSS.n8113 1.1255
R40855 DVSS.n8120 DVSS.n8119 1.1255
R40856 DVSS.n8121 DVSS.n4012 1.1255
R40857 DVSS.n8123 DVSS.n8122 1.1255
R40858 DVSS.n8127 DVSS.n8126 1.1255
R40859 DVSS.n8125 DVSS.n3845 1.1255
R40860 DVSS.n8333 DVSS.n3844 1.1255
R40861 DVSS.n8337 DVSS.n8335 1.1255
R40862 DVSS.n3413 DVSS.n3411 1.1255
R40863 DVSS.n8607 DVSS.n8606 1.1255
R40864 DVSS.n3408 DVSS.n3407 1.1255
R40865 DVSS.n8613 DVSS.n8612 1.1255
R40866 DVSS.n3065 DVSS.n3064 1.1255
R40867 DVSS.n8627 DVSS.n8626 1.1255
R40868 DVSS.n8632 DVSS.n8631 1.1255
R40869 DVSS.n3051 DVSS.n3050 1.1255
R40870 DVSS.n8981 DVSS.n8980 1.1255
R40871 DVSS.n8987 DVSS.n8986 1.1255
R40872 DVSS.n8988 DVSS.n3043 1.1255
R40873 DVSS.n8990 DVSS.n8989 1.1255
R40874 DVSS.n8994 DVSS.n8993 1.1255
R40875 DVSS.n8992 DVSS.n2877 1.1255
R40876 DVSS.n9200 DVSS.n2876 1.1255
R40877 DVSS.n9204 DVSS.n9202 1.1255
R40878 DVSS.n2737 DVSS.n2735 1.1255
R40879 DVSS.n9762 DVSS.n9761 1.1255
R40880 DVSS.n2732 DVSS.n2731 1.1255
R40881 DVSS.n9769 DVSS.n9768 1.1255
R40882 DVSS.n2716 DVSS.n2714 1.1255
R40883 DVSS.n10118 DVSS.n10117 1.1255
R40884 DVSS.n2710 DVSS.n2707 1.1255
R40885 DVSS.n10125 DVSS.n10124 1.1255
R40886 DVSS.n2711 DVSS.n2709 1.1255
R40887 DVSS.n10145 DVSS.n10144 1.1255
R40888 DVSS.n2366 DVSS.n2365 1.1255
R40889 DVSS.n10150 DVSS.n10149 1.1255
R40890 DVSS.n10169 DVSS.n10168 1.1255
R40891 DVSS.n2022 DVSS.n2020 1.1255
R40892 DVSS.n10459 DVSS.n10458 1.1255
R40893 DVSS.n1966 DVSS.n1965 1.1255
R40894 DVSS.n10480 DVSS.n10479 1.1255
R40895 DVSS.n1963 DVSS.n1962 1.1255
R40896 DVSS.n10485 DVSS.n10484 1.1255
R40897 DVSS.n10500 DVSS.n10499 1.1255
R40898 DVSS.n1619 DVSS.n1613 1.1255
R40899 DVSS.n10504 DVSS.n1615 1.1255
R40900 DVSS.n1509 DVSS.n1507 1.1255
R40901 DVSS.n13361 DVSS.n13360 1.1255
R40902 DVSS.n1510 DVSS.n1508 1.1255
R40903 DVSS.n13348 DVSS.n13347 1.1255
R40904 DVSS.n10770 DVSS.n10768 1.1255
R40905 DVSS.n13343 DVSS.n13342 1.1255
R40906 DVSS.n11615 DVSS.n11614 1.1255
R40907 DVSS.n11616 DVSS.n11611 1.1255
R40908 DVSS.n11618 DVSS.n11617 1.1255
R40909 DVSS.n13133 DVSS.n13132 1.1255
R40910 DVSS.n13131 DVSS.n11620 1.1255
R40911 DVSS.n13130 DVSS.n13129 1.1255
R40912 DVSS.n11623 DVSS.n11621 1.1255
R40913 DVSS.n13124 DVSS.n13123 1.1255
R40914 DVSS.n11629 DVSS.n11627 1.1255
R40915 DVSS.n12340 DVSS.n12339 1.1255
R40916 DVSS.n11998 DVSS.n11996 1.1255
R40917 DVSS.n13109 DVSS.n13108 1.1255
R40918 DVSS.n11999 DVSS.n11997 1.1255
R40919 DVSS.n13106 DVSS.n11999 1.1255
R40920 DVSS.n13108 DVSS.n13107 1.1255
R40921 DVSS.n12343 DVSS.n11998 1.1255
R40922 DVSS.n12341 DVSS.n12340 1.1255
R40923 DVSS.n11627 DVSS.n11625 1.1255
R40924 DVSS.n13125 DVSS.n13124 1.1255
R40925 DVSS.n13127 DVSS.n11623 1.1255
R40926 DVSS.n13129 DVSS.n13128 1.1255
R40927 DVSS.n11620 DVSS.n11610 1.1255
R40928 DVSS.n13134 DVSS.n13133 1.1255
R40929 DVSS.n11618 DVSS.n11609 1.1255
R40930 DVSS.n11612 DVSS.n11611 1.1255
R40931 DVSS.n11614 DVSS.n11613 1.1255
R40932 DVSS.n13344 DVSS.n13343 1.1255
R40933 DVSS.n13345 DVSS.n10770 1.1255
R40934 DVSS.n13347 DVSS.n13346 1.1255
R40935 DVSS.n1508 DVSS.n1506 1.1255
R40936 DVSS.n13362 DVSS.n13361 1.1255
R40937 DVSS.n1507 DVSS.n1505 1.1255
R40938 DVSS.n10504 DVSS.n10503 1.1255
R40939 DVSS.n10502 DVSS.n1613 1.1255
R40940 DVSS.n10501 DVSS.n10500 1.1255
R40941 DVSS.n10484 DVSS.n10483 1.1255
R40942 DVSS.n10482 DVSS.n1963 1.1255
R40943 DVSS.n10481 DVSS.n10480 1.1255
R40944 DVSS.n1965 DVSS.n1964 1.1255
R40945 DVSS.n10458 DVSS.n10457 1.1255
R40946 DVSS.n10171 DVSS.n2022 1.1255
R40947 DVSS.n10170 DVSS.n10169 1.1255
R40948 DVSS.n10149 DVSS.n10148 1.1255
R40949 DVSS.n10147 DVSS.n2366 1.1255
R40950 DVSS.n10146 DVSS.n10145 1.1255
R40951 DVSS.n10122 DVSS.n2711 1.1255
R40952 DVSS.n10124 DVSS.n10123 1.1255
R40953 DVSS.n10121 DVSS.n2710 1.1255
R40954 DVSS.n10119 DVSS.n10118 1.1255
R40955 DVSS.n2714 DVSS.n2713 1.1255
R40956 DVSS.n9768 DVSS.n9767 1.1255
R40957 DVSS.n9765 DVSS.n2732 1.1255
R40958 DVSS.n9763 DVSS.n9762 1.1255
R40959 DVSS.n2735 DVSS.n2734 1.1255
R40960 DVSS.n9204 DVSS.n9203 1.1255
R40961 DVSS.n3041 DVSS.n2876 1.1255
R40962 DVSS.n8992 DVSS.n3042 1.1255
R40963 DVSS.n8995 DVSS.n8994 1.1255
R40964 DVSS.n8990 DVSS.n3040 1.1255
R40965 DVSS.n8984 DVSS.n3043 1.1255
R40966 DVSS.n8986 DVSS.n8985 1.1255
R40967 DVSS.n8982 DVSS.n8981 1.1255
R40968 DVSS.n3050 DVSS.n3049 1.1255
R40969 DVSS.n8631 DVSS.n8630 1.1255
R40970 DVSS.n8628 DVSS.n8627 1.1255
R40971 DVSS.n3064 DVSS.n3063 1.1255
R40972 DVSS.n8612 DVSS.n8611 1.1255
R40973 DVSS.n8610 DVSS.n3408 1.1255
R40974 DVSS.n8608 DVSS.n8607 1.1255
R40975 DVSS.n3411 DVSS.n3410 1.1255
R40976 DVSS.n8337 DVSS.n8336 1.1255
R40977 DVSS.n4009 DVSS.n3844 1.1255
R40978 DVSS.n8125 DVSS.n4011 1.1255
R40979 DVSS.n8128 DVSS.n8127 1.1255
R40980 DVSS.n8123 DVSS.n4008 1.1255
R40981 DVSS.n8117 DVSS.n4012 1.1255
R40982 DVSS.n8119 DVSS.n8118 1.1255
R40983 DVSS.n8115 DVSS.n8114 1.1255
R40984 DVSS.n4019 DVSS.n4018 1.1255
R40985 DVSS.n8098 DVSS.n8097 1.1255
R40986 DVSS.n8096 DVSS.n4364 1.1255
R40987 DVSS.n8094 DVSS.n8093 1.1255
R40988 DVSS.n4367 DVSS.n4366 1.1255
R40989 DVSS.n7824 DVSS.n7823 1.1255
R40990 DVSS.n7821 DVSS.n7820 1.1255
R40991 DVSS.n4809 DVSS.n4808 1.1255
R40992 DVSS.n7804 DVSS.n7803 1.1255
R40993 DVSS.n7801 DVSS.n7800 1.1255
R40994 DVSS.n4823 DVSS.n4822 1.1255
R40995 DVSS.n7446 DVSS.n7445 1.1255
R40996 DVSS.n7449 DVSS.n7448 1.1255
R40997 DVSS.n7109 DVSS.n4835 1.1255
R40998 DVSS.n7108 DVSS.n7107 1.1255
R40999 DVSS.n4838 DVSS.n4837 1.1255
R41000 DVSS.n7085 DVSS.n7084 1.1255
R41001 DVSS.n7083 DVSS.n5178 1.1255
R41002 DVSS.n7082 DVSS.n7081 1.1255
R41003 DVSS.n7066 DVSS.n7065 1.1255
R41004 DVSS.n7064 DVSS.n5527 1.1255
R41005 DVSS.n7063 DVSS.n7062 1.1255
R41006 DVSS.n7040 DVSS.n5871 1.1255
R41007 DVSS.n7042 DVSS.n7041 1.1255
R41008 DVSS.n7039 DVSS.n5870 1.1255
R41009 DVSS.n7037 DVSS.n7036 1.1255
R41010 DVSS.n5874 DVSS.n5873 1.1255
R41011 DVSS.n6686 DVSS.n6685 1.1255
R41012 DVSS.n6683 DVSS.n6682 1.1255
R41013 DVSS.n5895 DVSS.n5894 1.1255
R41014 DVSS.n6668 DVSS.n6667 1.1255
R41015 DVSS.n18154 DVSS.n18153 1.1255
R41016 DVSS.n15555 DVSS.n15546 1.1255
R41017 DVSS.n15578 DVSS.n15577 1.1255
R41018 DVSS.n15580 DVSS.n15579 1.1255
R41019 DVSS.n15581 DVSS.n15575 1.1255
R41020 DVSS.n18147 DVSS.n18146 1.1255
R41021 DVSS.n18145 DVSS.n15576 1.1255
R41022 DVSS.n18144 DVSS.n18143 1.1255
R41023 DVSS.n18142 DVSS.n15582 1.1255
R41024 DVSS.n18141 DVSS.n18140 1.1255
R41025 DVSS.n18139 DVSS.n15583 1.1255
R41026 DVSS.n18138 DVSS.n18137 1.1255
R41027 DVSS.n18136 DVSS.n18135 1.1255
R41028 DVSS.n18134 DVSS.n15585 1.1255
R41029 DVSS.n18133 DVSS.n18132 1.1255
R41030 DVSS.n18131 DVSS.n15586 1.1255
R41031 DVSS.n18130 DVSS.n18129 1.1255
R41032 DVSS.n18128 DVSS.n15587 1.1255
R41033 DVSS.n18127 DVSS.n18126 1.1255
R41034 DVSS.n18125 DVSS.n15588 1.1255
R41035 DVSS.n18124 DVSS.n18123 1.1255
R41036 DVSS.n18122 DVSS.n18121 1.1255
R41037 DVSS.n15598 DVSS.n15590 1.1255
R41038 DVSS.n18097 DVSS.n18096 1.1255
R41039 DVSS.n18099 DVSS.n18098 1.1255
R41040 DVSS.n18101 DVSS.n18100 1.1255
R41041 DVSS.n18109 DVSS.n18108 1.1255
R41042 DVSS.n14846 DVSS.n14845 1.12321
R41043 DVSS.n14845 DVSS.n14739 1.11525
R41044 DVSS.n19895 DVSS 1.09758
R41045 DVSS.n19892 DVSS 1.09758
R41046 DVSS DVSS.n19885 1.09758
R41047 DVSS.n19882 DVSS 1.09758
R41048 DVSS.n19879 DVSS 1.09758
R41049 DVSS DVSS.n19872 1.09758
R41050 DVSS.n19869 DVSS 1.09758
R41051 DVSS.n19866 DVSS 1.09758
R41052 DVSS DVSS.n19859 1.09758
R41053 DVSS.n19856 DVSS 1.09758
R41054 DVSS.n19853 DVSS 1.09758
R41055 DVSS.n19588 DVSS 1.09758
R41056 DVSS.n19585 DVSS 1.09758
R41057 DVSS DVSS.n19578 1.09758
R41058 DVSS.n19575 DVSS 1.09758
R41059 DVSS.n19572 DVSS 1.09758
R41060 DVSS DVSS.n19565 1.09758
R41061 DVSS.n19562 DVSS 1.09758
R41062 DVSS.n19559 DVSS 1.09758
R41063 DVSS DVSS.n19552 1.09758
R41064 DVSS.n19549 DVSS 1.09758
R41065 DVSS.n19546 DVSS 1.09758
R41066 DVSS.n663 DVSS 1.09758
R41067 DVSS DVSS.n21831 1.09758
R41068 DVSS.n21841 DVSS 1.09758
R41069 DVSS.n21844 DVSS 1.09758
R41070 DVSS.n21848 DVSS 1.09758
R41071 DVSS DVSS.n21947 1.09758
R41072 DVSS.n21939 DVSS 1.09758
R41073 DVSS.n21917 DVSS 1.09758
R41074 DVSS.n21907 DVSS 1.09758
R41075 DVSS.n21897 DVSS 1.09758
R41076 DVSS.n21887 DVSS 1.09758
R41077 DVSS.n855 DVSS 1.09758
R41078 DVSS.n847 DVSS 1.09758
R41079 DVSS.n838 DVSS 1.09758
R41080 DVSS.n829 DVSS 1.09758
R41081 DVSS.n820 DVSS 1.09758
R41082 DVSS.n22481 DVSS 1.09758
R41083 DVSS DVSS.n13043 1.09758
R41084 DVSS DVSS.n13031 1.09758
R41085 DVSS DVSS.n13052 1.09758
R41086 DVSS.n22376 DVSS 1.09758
R41087 DVSS DVSS.n13017 1.09723
R41088 DVSS.n18999 DVSS.n13527 1.09353
R41089 DVSS.n13059 DVSS 1.09186
R41090 DVSS.n19144 DVSS 1.09158
R41091 DVSS DVSS.n19890 1.09158
R41092 DVSS.n19887 DVSS 1.09158
R41093 DVSS.n19050 DVSS 1.09158
R41094 DVSS DVSS.n19877 1.09158
R41095 DVSS.n19874 DVSS 1.09158
R41096 DVSS.n19058 DVSS 1.09158
R41097 DVSS DVSS.n19864 1.09158
R41098 DVSS.n19861 DVSS 1.09158
R41099 DVSS.n19066 DVSS 1.09158
R41100 DVSS DVSS.n19852 1.09158
R41101 DVSS.n19519 DVSS 1.09158
R41102 DVSS DVSS.n19583 1.09158
R41103 DVSS.n19580 DVSS 1.09158
R41104 DVSS.n19526 DVSS 1.09158
R41105 DVSS DVSS.n19570 1.09158
R41106 DVSS.n19567 DVSS 1.09158
R41107 DVSS.n19534 DVSS 1.09158
R41108 DVSS DVSS.n19557 1.09158
R41109 DVSS.n19554 DVSS 1.09158
R41110 DVSS.n19541 DVSS 1.09158
R41111 DVSS DVSS.n19545 1.09158
R41112 DVSS DVSS.n661 1.09158
R41113 DVSS.n21833 DVSS 1.09158
R41114 DVSS DVSS.n21839 1.09158
R41115 DVSS.n21836 DVSS 1.09158
R41116 DVSS DVSS.n21846 1.09158
R41117 DVSS.n21949 DVSS 1.09158
R41118 DVSS DVSS.n21936 1.09158
R41119 DVSS DVSS.n21914 1.09158
R41120 DVSS DVSS.n21904 1.09158
R41121 DVSS DVSS.n21894 1.09158
R41122 DVSS DVSS.n21885 1.09158
R41123 DVSS DVSS.n853 1.09158
R41124 DVSS DVSS.n844 1.09158
R41125 DVSS DVSS.n835 1.09158
R41126 DVSS DVSS.n826 1.09158
R41127 DVSS DVSS.n817 1.09158
R41128 DVSS DVSS.n22479 1.09158
R41129 DVSS.n13045 DVSS 1.09158
R41130 DVSS.n13033 DVSS 1.09158
R41131 DVSS.n13054 DVSS 1.09158
R41132 DVSS.n13019 DVSS 1.09158
R41133 DVSS.n13662 DVSS.n13660 1.09023
R41134 DVSS.n13686 DVSS.n13685 1.06594
R41135 DVSS.n15917 DVSS.n15539 1.0621
R41136 DVSS.n18164 DVSS.n18163 1.0621
R41137 DVSS.n21446 DVSS.n21445 1.0621
R41138 DVSS.n13366 DVSS.n13365 1.0621
R41139 DVSS.n20474 DVSS.n14847 1.03912
R41140 DVSS.n17792 DVSS.n15918 1.02343
R41141 DVSS.n22636 DVSS.n734 1.02241
R41142 DVSS.n21440 DVSS.n453 1.02241
R41143 DVSS.n18166 DVSS.n18165 1.0144
R41144 DVSS.n13676 DVSS.n13673 0.994213
R41145 DVSS.n22937 DVSS.n22936 0.982731
R41146 DVSS.n21013 DVSS.n21012 0.982731
R41147 DVSS.n22585 DVSS.n22584 0.982731
R41148 DVSS.n21472 DVSS.n21447 0.959128
R41149 DVSS.n22970 DVSS.n423 0.950107
R41150 DVSS.n19209 DVSS.t167 0.913226
R41151 DVSS.n19183 DVSS.t173 0.913226
R41152 DVSS.n19182 DVSS.t188 0.913226
R41153 DVSS.n20507 DVSS.n20474 0.903572
R41154 DVSS.n12766 DVSS.n12765 0.902975
R41155 DVSS.n6653 DVSS.n6234 0.902975
R41156 DVSS.n12744 DVSS.n12555 0.9005
R41157 DVSS.n12741 DVSS.n12740 0.9005
R41158 DVSS.n12739 DVSS.n12556 0.9005
R41159 DVSS.n12738 DVSS.n12737 0.9005
R41160 DVSS.n12736 DVSS.n12557 0.9005
R41161 DVSS.n12735 DVSS.n12734 0.9005
R41162 DVSS.n12733 DVSS.n12558 0.9005
R41163 DVSS.n12732 DVSS.n12731 0.9005
R41164 DVSS.n12730 DVSS.n12559 0.9005
R41165 DVSS.n12729 DVSS.n12728 0.9005
R41166 DVSS.n12727 DVSS.n12560 0.9005
R41167 DVSS.n12726 DVSS.n12725 0.9005
R41168 DVSS.n12724 DVSS.n12561 0.9005
R41169 DVSS.n12723 DVSS.n12722 0.9005
R41170 DVSS.n12721 DVSS.n12562 0.9005
R41171 DVSS.n12720 DVSS.n12719 0.9005
R41172 DVSS.n12718 DVSS.n12563 0.9005
R41173 DVSS.n12717 DVSS.n12716 0.9005
R41174 DVSS.n12715 DVSS.n12564 0.9005
R41175 DVSS.n12714 DVSS.n12713 0.9005
R41176 DVSS.n12712 DVSS.n12565 0.9005
R41177 DVSS.n12711 DVSS.n12710 0.9005
R41178 DVSS.n12709 DVSS.n12566 0.9005
R41179 DVSS.n12708 DVSS.n12707 0.9005
R41180 DVSS.n12706 DVSS.n12567 0.9005
R41181 DVSS.n12705 DVSS.n12704 0.9005
R41182 DVSS.n12703 DVSS.n12568 0.9005
R41183 DVSS.n12702 DVSS.n12701 0.9005
R41184 DVSS.n12700 DVSS.n12569 0.9005
R41185 DVSS.n12699 DVSS.n12698 0.9005
R41186 DVSS.n12697 DVSS.n12570 0.9005
R41187 DVSS.n12696 DVSS.n12695 0.9005
R41188 DVSS.n12694 DVSS.n12571 0.9005
R41189 DVSS.n12693 DVSS.n12692 0.9005
R41190 DVSS.n12691 DVSS.n12572 0.9005
R41191 DVSS.n12690 DVSS.n12689 0.9005
R41192 DVSS.n12688 DVSS.n12573 0.9005
R41193 DVSS.n12687 DVSS.n12686 0.9005
R41194 DVSS.n12685 DVSS.n12574 0.9005
R41195 DVSS.n12684 DVSS.n12683 0.9005
R41196 DVSS.n12682 DVSS.n12575 0.9005
R41197 DVSS.n12681 DVSS.n12680 0.9005
R41198 DVSS.n12679 DVSS.n12576 0.9005
R41199 DVSS.n12678 DVSS.n12677 0.9005
R41200 DVSS.n12676 DVSS.n12577 0.9005
R41201 DVSS.n12675 DVSS.n12674 0.9005
R41202 DVSS.n12673 DVSS.n12578 0.9005
R41203 DVSS.n12672 DVSS.n12671 0.9005
R41204 DVSS.n12670 DVSS.n12579 0.9005
R41205 DVSS.n12669 DVSS.n12668 0.9005
R41206 DVSS.n12667 DVSS.n12580 0.9005
R41207 DVSS.n12666 DVSS.n12665 0.9005
R41208 DVSS.n12664 DVSS.n12581 0.9005
R41209 DVSS.n12663 DVSS.n12662 0.9005
R41210 DVSS.n12661 DVSS.n12582 0.9005
R41211 DVSS.n12660 DVSS.n12659 0.9005
R41212 DVSS.n12658 DVSS.n12583 0.9005
R41213 DVSS.n12657 DVSS.n12656 0.9005
R41214 DVSS.n12655 DVSS.n12584 0.9005
R41215 DVSS.n12654 DVSS.n12653 0.9005
R41216 DVSS.n12652 DVSS.n12585 0.9005
R41217 DVSS.n12651 DVSS.n12650 0.9005
R41218 DVSS.n12649 DVSS.n12586 0.9005
R41219 DVSS.n12648 DVSS.n12647 0.9005
R41220 DVSS.n12646 DVSS.n12587 0.9005
R41221 DVSS.n12645 DVSS.n12644 0.9005
R41222 DVSS.n12643 DVSS.n12588 0.9005
R41223 DVSS.n12642 DVSS.n12641 0.9005
R41224 DVSS.n12640 DVSS.n12589 0.9005
R41225 DVSS.n12639 DVSS.n12638 0.9005
R41226 DVSS.n12637 DVSS.n12590 0.9005
R41227 DVSS.n12636 DVSS.n12635 0.9005
R41228 DVSS.n12634 DVSS.n12591 0.9005
R41229 DVSS.n12633 DVSS.n12632 0.9005
R41230 DVSS.n12631 DVSS.n12592 0.9005
R41231 DVSS.n12630 DVSS.n12629 0.9005
R41232 DVSS.n12628 DVSS.n12593 0.9005
R41233 DVSS.n12627 DVSS.n12626 0.9005
R41234 DVSS.n12625 DVSS.n12594 0.9005
R41235 DVSS.n12624 DVSS.n12623 0.9005
R41236 DVSS.n12622 DVSS.n12595 0.9005
R41237 DVSS.n12621 DVSS.n12620 0.9005
R41238 DVSS.n12619 DVSS.n12596 0.9005
R41239 DVSS.n12618 DVSS.n12617 0.9005
R41240 DVSS.n12616 DVSS.n12597 0.9005
R41241 DVSS.n12615 DVSS.n12614 0.9005
R41242 DVSS.n12613 DVSS.n12598 0.9005
R41243 DVSS.n12612 DVSS.n12611 0.9005
R41244 DVSS.n12610 DVSS.n12599 0.9005
R41245 DVSS.n12609 DVSS.n12608 0.9005
R41246 DVSS.n12607 DVSS.n12600 0.9005
R41247 DVSS.n12606 DVSS.n12605 0.9005
R41248 DVSS.n12604 DVSS.n12601 0.9005
R41249 DVSS.n12603 DVSS.n12602 0.9005
R41250 DVSS.n12356 DVSS.n12355 0.9005
R41251 DVSS.n12771 DVSS.n12770 0.9005
R41252 DVSS.n12772 DVSS.n12353 0.9005
R41253 DVSS.n12747 DVSS.n12746 0.9005
R41254 DVSS.n12746 DVSS.n12745 0.9005
R41255 DVSS.n12744 DVSS.n12743 0.9005
R41256 DVSS.n12741 DVSS.n12411 0.9005
R41257 DVSS.n12556 DVSS.n12409 0.9005
R41258 DVSS.n12737 DVSS.n12412 0.9005
R41259 DVSS.n12736 DVSS.n12408 0.9005
R41260 DVSS.n12735 DVSS.n12413 0.9005
R41261 DVSS.n12558 DVSS.n12407 0.9005
R41262 DVSS.n12731 DVSS.n12414 0.9005
R41263 DVSS.n12730 DVSS.n12406 0.9005
R41264 DVSS.n12729 DVSS.n12415 0.9005
R41265 DVSS.n12560 DVSS.n12405 0.9005
R41266 DVSS.n12725 DVSS.n12416 0.9005
R41267 DVSS.n12724 DVSS.n12404 0.9005
R41268 DVSS.n12723 DVSS.n12417 0.9005
R41269 DVSS.n12562 DVSS.n12403 0.9005
R41270 DVSS.n12719 DVSS.n12418 0.9005
R41271 DVSS.n12718 DVSS.n12402 0.9005
R41272 DVSS.n12717 DVSS.n12419 0.9005
R41273 DVSS.n12564 DVSS.n12401 0.9005
R41274 DVSS.n12713 DVSS.n12420 0.9005
R41275 DVSS.n12712 DVSS.n12400 0.9005
R41276 DVSS.n12711 DVSS.n12421 0.9005
R41277 DVSS.n12566 DVSS.n12399 0.9005
R41278 DVSS.n12707 DVSS.n12422 0.9005
R41279 DVSS.n12706 DVSS.n12398 0.9005
R41280 DVSS.n12705 DVSS.n12423 0.9005
R41281 DVSS.n12568 DVSS.n12397 0.9005
R41282 DVSS.n12701 DVSS.n12424 0.9005
R41283 DVSS.n12700 DVSS.n12396 0.9005
R41284 DVSS.n12699 DVSS.n12425 0.9005
R41285 DVSS.n12570 DVSS.n12395 0.9005
R41286 DVSS.n12695 DVSS.n12426 0.9005
R41287 DVSS.n12694 DVSS.n12394 0.9005
R41288 DVSS.n12693 DVSS.n12427 0.9005
R41289 DVSS.n12572 DVSS.n12393 0.9005
R41290 DVSS.n12689 DVSS.n12428 0.9005
R41291 DVSS.n12688 DVSS.n12392 0.9005
R41292 DVSS.n12687 DVSS.n12429 0.9005
R41293 DVSS.n12574 DVSS.n12391 0.9005
R41294 DVSS.n12683 DVSS.n12430 0.9005
R41295 DVSS.n12682 DVSS.n12390 0.9005
R41296 DVSS.n12681 DVSS.n12431 0.9005
R41297 DVSS.n12576 DVSS.n12389 0.9005
R41298 DVSS.n12677 DVSS.n12432 0.9005
R41299 DVSS.n12676 DVSS.n12388 0.9005
R41300 DVSS.n12675 DVSS.n12433 0.9005
R41301 DVSS.n12578 DVSS.n12387 0.9005
R41302 DVSS.n12671 DVSS.n12434 0.9005
R41303 DVSS.n12670 DVSS.n12386 0.9005
R41304 DVSS.n12669 DVSS.n12435 0.9005
R41305 DVSS.n12580 DVSS.n12385 0.9005
R41306 DVSS.n12665 DVSS.n12436 0.9005
R41307 DVSS.n12664 DVSS.n12384 0.9005
R41308 DVSS.n12663 DVSS.n12437 0.9005
R41309 DVSS.n12582 DVSS.n12383 0.9005
R41310 DVSS.n12659 DVSS.n12438 0.9005
R41311 DVSS.n12658 DVSS.n12382 0.9005
R41312 DVSS.n12657 DVSS.n12439 0.9005
R41313 DVSS.n12584 DVSS.n12381 0.9005
R41314 DVSS.n12653 DVSS.n12440 0.9005
R41315 DVSS.n12652 DVSS.n12380 0.9005
R41316 DVSS.n12651 DVSS.n12441 0.9005
R41317 DVSS.n12586 DVSS.n12379 0.9005
R41318 DVSS.n12647 DVSS.n12442 0.9005
R41319 DVSS.n12646 DVSS.n12378 0.9005
R41320 DVSS.n12645 DVSS.n12443 0.9005
R41321 DVSS.n12588 DVSS.n12377 0.9005
R41322 DVSS.n12641 DVSS.n12444 0.9005
R41323 DVSS.n12640 DVSS.n12376 0.9005
R41324 DVSS.n12639 DVSS.n12445 0.9005
R41325 DVSS.n12590 DVSS.n12375 0.9005
R41326 DVSS.n12635 DVSS.n12446 0.9005
R41327 DVSS.n12634 DVSS.n12374 0.9005
R41328 DVSS.n12633 DVSS.n12447 0.9005
R41329 DVSS.n12592 DVSS.n12373 0.9005
R41330 DVSS.n12629 DVSS.n12448 0.9005
R41331 DVSS.n12628 DVSS.n12372 0.9005
R41332 DVSS.n12627 DVSS.n12449 0.9005
R41333 DVSS.n12594 DVSS.n12371 0.9005
R41334 DVSS.n12623 DVSS.n12450 0.9005
R41335 DVSS.n12622 DVSS.n12370 0.9005
R41336 DVSS.n12621 DVSS.n12451 0.9005
R41337 DVSS.n12596 DVSS.n12369 0.9005
R41338 DVSS.n12617 DVSS.n12452 0.9005
R41339 DVSS.n12616 DVSS.n12368 0.9005
R41340 DVSS.n12615 DVSS.n12453 0.9005
R41341 DVSS.n12598 DVSS.n12367 0.9005
R41342 DVSS.n12611 DVSS.n12454 0.9005
R41343 DVSS.n12610 DVSS.n12366 0.9005
R41344 DVSS.n12609 DVSS.n12455 0.9005
R41345 DVSS.n12600 DVSS.n12365 0.9005
R41346 DVSS.n12605 DVSS.n12456 0.9005
R41347 DVSS.n12604 DVSS.n12364 0.9005
R41348 DVSS.n12603 DVSS.n12457 0.9005
R41349 DVSS.n12363 DVSS.n12356 0.9005
R41350 DVSS.n12770 DVSS.n12769 0.9005
R41351 DVSS.n12362 DVSS.n12353 0.9005
R41352 DVSS.n12767 DVSS.n12766 0.9005
R41353 DVSS.n6655 DVSS.n6653 0.9005
R41354 DVSS.n6406 DVSS.n6309 0.9005
R41355 DVSS.n6308 DVSS.n6247 0.9005
R41356 DVSS.n6455 DVSS.n6311 0.9005
R41357 DVSS.n6452 DVSS.n6307 0.9005
R41358 DVSS.n6459 DVSS.n6313 0.9005
R41359 DVSS.n6460 DVSS.n6306 0.9005
R41360 DVSS.n6461 DVSS.n6315 0.9005
R41361 DVSS.n6450 DVSS.n6305 0.9005
R41362 DVSS.n6465 DVSS.n6317 0.9005
R41363 DVSS.n6466 DVSS.n6304 0.9005
R41364 DVSS.n6467 DVSS.n6319 0.9005
R41365 DVSS.n6448 DVSS.n6303 0.9005
R41366 DVSS.n6471 DVSS.n6321 0.9005
R41367 DVSS.n6472 DVSS.n6302 0.9005
R41368 DVSS.n6473 DVSS.n6323 0.9005
R41369 DVSS.n6446 DVSS.n6301 0.9005
R41370 DVSS.n6477 DVSS.n6325 0.9005
R41371 DVSS.n6478 DVSS.n6300 0.9005
R41372 DVSS.n6479 DVSS.n6327 0.9005
R41373 DVSS.n6444 DVSS.n6299 0.9005
R41374 DVSS.n6483 DVSS.n6329 0.9005
R41375 DVSS.n6484 DVSS.n6298 0.9005
R41376 DVSS.n6485 DVSS.n6331 0.9005
R41377 DVSS.n6442 DVSS.n6297 0.9005
R41378 DVSS.n6489 DVSS.n6333 0.9005
R41379 DVSS.n6490 DVSS.n6296 0.9005
R41380 DVSS.n6491 DVSS.n6335 0.9005
R41381 DVSS.n6440 DVSS.n6295 0.9005
R41382 DVSS.n6495 DVSS.n6337 0.9005
R41383 DVSS.n6496 DVSS.n6294 0.9005
R41384 DVSS.n6497 DVSS.n6339 0.9005
R41385 DVSS.n6438 DVSS.n6293 0.9005
R41386 DVSS.n6501 DVSS.n6341 0.9005
R41387 DVSS.n6502 DVSS.n6292 0.9005
R41388 DVSS.n6503 DVSS.n6343 0.9005
R41389 DVSS.n6436 DVSS.n6291 0.9005
R41390 DVSS.n6507 DVSS.n6345 0.9005
R41391 DVSS.n6508 DVSS.n6290 0.9005
R41392 DVSS.n6509 DVSS.n6347 0.9005
R41393 DVSS.n6434 DVSS.n6289 0.9005
R41394 DVSS.n6513 DVSS.n6349 0.9005
R41395 DVSS.n6514 DVSS.n6288 0.9005
R41396 DVSS.n6515 DVSS.n6351 0.9005
R41397 DVSS.n6432 DVSS.n6287 0.9005
R41398 DVSS.n6519 DVSS.n6353 0.9005
R41399 DVSS.n6520 DVSS.n6286 0.9005
R41400 DVSS.n6521 DVSS.n6355 0.9005
R41401 DVSS.n6430 DVSS.n6285 0.9005
R41402 DVSS.n6525 DVSS.n6357 0.9005
R41403 DVSS.n6526 DVSS.n6284 0.9005
R41404 DVSS.n6527 DVSS.n6359 0.9005
R41405 DVSS.n6428 DVSS.n6283 0.9005
R41406 DVSS.n6531 DVSS.n6361 0.9005
R41407 DVSS.n6532 DVSS.n6282 0.9005
R41408 DVSS.n6533 DVSS.n6363 0.9005
R41409 DVSS.n6426 DVSS.n6281 0.9005
R41410 DVSS.n6537 DVSS.n6365 0.9005
R41411 DVSS.n6538 DVSS.n6280 0.9005
R41412 DVSS.n6539 DVSS.n6367 0.9005
R41413 DVSS.n6424 DVSS.n6279 0.9005
R41414 DVSS.n6543 DVSS.n6369 0.9005
R41415 DVSS.n6544 DVSS.n6278 0.9005
R41416 DVSS.n6545 DVSS.n6371 0.9005
R41417 DVSS.n6422 DVSS.n6277 0.9005
R41418 DVSS.n6549 DVSS.n6373 0.9005
R41419 DVSS.n6550 DVSS.n6276 0.9005
R41420 DVSS.n6551 DVSS.n6375 0.9005
R41421 DVSS.n6420 DVSS.n6275 0.9005
R41422 DVSS.n6555 DVSS.n6377 0.9005
R41423 DVSS.n6556 DVSS.n6274 0.9005
R41424 DVSS.n6557 DVSS.n6379 0.9005
R41425 DVSS.n6418 DVSS.n6273 0.9005
R41426 DVSS.n6561 DVSS.n6381 0.9005
R41427 DVSS.n6562 DVSS.n6272 0.9005
R41428 DVSS.n6563 DVSS.n6383 0.9005
R41429 DVSS.n6416 DVSS.n6271 0.9005
R41430 DVSS.n6567 DVSS.n6385 0.9005
R41431 DVSS.n6568 DVSS.n6270 0.9005
R41432 DVSS.n6569 DVSS.n6387 0.9005
R41433 DVSS.n6414 DVSS.n6269 0.9005
R41434 DVSS.n6573 DVSS.n6389 0.9005
R41435 DVSS.n6574 DVSS.n6268 0.9005
R41436 DVSS.n6575 DVSS.n6391 0.9005
R41437 DVSS.n6412 DVSS.n6267 0.9005
R41438 DVSS.n6579 DVSS.n6393 0.9005
R41439 DVSS.n6580 DVSS.n6266 0.9005
R41440 DVSS.n6581 DVSS.n6395 0.9005
R41441 DVSS.n6410 DVSS.n6265 0.9005
R41442 DVSS.n6585 DVSS.n6397 0.9005
R41443 DVSS.n6586 DVSS.n6264 0.9005
R41444 DVSS.n6587 DVSS.n6399 0.9005
R41445 DVSS.n6408 DVSS.n6263 0.9005
R41446 DVSS.n6591 DVSS.n6401 0.9005
R41447 DVSS.n6592 DVSS.n6262 0.9005
R41448 DVSS.n6593 DVSS.n6403 0.9005
R41449 DVSS.n6405 DVSS.n6261 0.9005
R41450 DVSS.n6601 DVSS.n6600 0.9005
R41451 DVSS.n6596 DVSS.n6260 0.9005
R41452 DVSS.n6454 DVSS.n6247 0.9005
R41453 DVSS.n6456 DVSS.n6455 0.9005
R41454 DVSS.n6457 DVSS.n6452 0.9005
R41455 DVSS.n6459 DVSS.n6458 0.9005
R41456 DVSS.n6460 DVSS.n6451 0.9005
R41457 DVSS.n6462 DVSS.n6461 0.9005
R41458 DVSS.n6463 DVSS.n6450 0.9005
R41459 DVSS.n6465 DVSS.n6464 0.9005
R41460 DVSS.n6466 DVSS.n6449 0.9005
R41461 DVSS.n6468 DVSS.n6467 0.9005
R41462 DVSS.n6469 DVSS.n6448 0.9005
R41463 DVSS.n6471 DVSS.n6470 0.9005
R41464 DVSS.n6472 DVSS.n6447 0.9005
R41465 DVSS.n6474 DVSS.n6473 0.9005
R41466 DVSS.n6475 DVSS.n6446 0.9005
R41467 DVSS.n6477 DVSS.n6476 0.9005
R41468 DVSS.n6478 DVSS.n6445 0.9005
R41469 DVSS.n6480 DVSS.n6479 0.9005
R41470 DVSS.n6481 DVSS.n6444 0.9005
R41471 DVSS.n6483 DVSS.n6482 0.9005
R41472 DVSS.n6484 DVSS.n6443 0.9005
R41473 DVSS.n6486 DVSS.n6485 0.9005
R41474 DVSS.n6487 DVSS.n6442 0.9005
R41475 DVSS.n6489 DVSS.n6488 0.9005
R41476 DVSS.n6490 DVSS.n6441 0.9005
R41477 DVSS.n6492 DVSS.n6491 0.9005
R41478 DVSS.n6493 DVSS.n6440 0.9005
R41479 DVSS.n6495 DVSS.n6494 0.9005
R41480 DVSS.n6496 DVSS.n6439 0.9005
R41481 DVSS.n6498 DVSS.n6497 0.9005
R41482 DVSS.n6499 DVSS.n6438 0.9005
R41483 DVSS.n6501 DVSS.n6500 0.9005
R41484 DVSS.n6502 DVSS.n6437 0.9005
R41485 DVSS.n6504 DVSS.n6503 0.9005
R41486 DVSS.n6505 DVSS.n6436 0.9005
R41487 DVSS.n6507 DVSS.n6506 0.9005
R41488 DVSS.n6508 DVSS.n6435 0.9005
R41489 DVSS.n6510 DVSS.n6509 0.9005
R41490 DVSS.n6511 DVSS.n6434 0.9005
R41491 DVSS.n6513 DVSS.n6512 0.9005
R41492 DVSS.n6514 DVSS.n6433 0.9005
R41493 DVSS.n6516 DVSS.n6515 0.9005
R41494 DVSS.n6517 DVSS.n6432 0.9005
R41495 DVSS.n6519 DVSS.n6518 0.9005
R41496 DVSS.n6520 DVSS.n6431 0.9005
R41497 DVSS.n6522 DVSS.n6521 0.9005
R41498 DVSS.n6523 DVSS.n6430 0.9005
R41499 DVSS.n6525 DVSS.n6524 0.9005
R41500 DVSS.n6526 DVSS.n6429 0.9005
R41501 DVSS.n6528 DVSS.n6527 0.9005
R41502 DVSS.n6529 DVSS.n6428 0.9005
R41503 DVSS.n6531 DVSS.n6530 0.9005
R41504 DVSS.n6532 DVSS.n6427 0.9005
R41505 DVSS.n6534 DVSS.n6533 0.9005
R41506 DVSS.n6535 DVSS.n6426 0.9005
R41507 DVSS.n6537 DVSS.n6536 0.9005
R41508 DVSS.n6538 DVSS.n6425 0.9005
R41509 DVSS.n6540 DVSS.n6539 0.9005
R41510 DVSS.n6541 DVSS.n6424 0.9005
R41511 DVSS.n6543 DVSS.n6542 0.9005
R41512 DVSS.n6544 DVSS.n6423 0.9005
R41513 DVSS.n6546 DVSS.n6545 0.9005
R41514 DVSS.n6547 DVSS.n6422 0.9005
R41515 DVSS.n6549 DVSS.n6548 0.9005
R41516 DVSS.n6550 DVSS.n6421 0.9005
R41517 DVSS.n6552 DVSS.n6551 0.9005
R41518 DVSS.n6553 DVSS.n6420 0.9005
R41519 DVSS.n6555 DVSS.n6554 0.9005
R41520 DVSS.n6556 DVSS.n6419 0.9005
R41521 DVSS.n6558 DVSS.n6557 0.9005
R41522 DVSS.n6559 DVSS.n6418 0.9005
R41523 DVSS.n6561 DVSS.n6560 0.9005
R41524 DVSS.n6562 DVSS.n6417 0.9005
R41525 DVSS.n6564 DVSS.n6563 0.9005
R41526 DVSS.n6565 DVSS.n6416 0.9005
R41527 DVSS.n6567 DVSS.n6566 0.9005
R41528 DVSS.n6568 DVSS.n6415 0.9005
R41529 DVSS.n6570 DVSS.n6569 0.9005
R41530 DVSS.n6571 DVSS.n6414 0.9005
R41531 DVSS.n6573 DVSS.n6572 0.9005
R41532 DVSS.n6574 DVSS.n6413 0.9005
R41533 DVSS.n6576 DVSS.n6575 0.9005
R41534 DVSS.n6577 DVSS.n6412 0.9005
R41535 DVSS.n6579 DVSS.n6578 0.9005
R41536 DVSS.n6580 DVSS.n6411 0.9005
R41537 DVSS.n6582 DVSS.n6581 0.9005
R41538 DVSS.n6583 DVSS.n6410 0.9005
R41539 DVSS.n6585 DVSS.n6584 0.9005
R41540 DVSS.n6586 DVSS.n6409 0.9005
R41541 DVSS.n6588 DVSS.n6587 0.9005
R41542 DVSS.n6589 DVSS.n6408 0.9005
R41543 DVSS.n6591 DVSS.n6590 0.9005
R41544 DVSS.n6592 DVSS.n6407 0.9005
R41545 DVSS.n6594 DVSS.n6593 0.9005
R41546 DVSS.n6595 DVSS.n6405 0.9005
R41547 DVSS.n6600 DVSS.n6599 0.9005
R41548 DVSS.n6598 DVSS.n6406 0.9005
R41549 DVSS.n6597 DVSS.n6596 0.9005
R41550 DVSS.n21156 DVSS.n13683 0.826598
R41551 DVSS.n21154 DVSS.n13685 0.825923
R41552 DVSS.n22961 DVSS.n425 0.805246
R41553 DVSS.n22960 DVSS.n427 0.805246
R41554 DVSS.n20986 DVSS.n14312 0.805246
R41555 DVSS.n21462 DVSS.n21461 0.805246
R41556 DVSS.n21463 DVSS.n21449 0.805246
R41557 DVSS.n22637 DVSS.n22636 0.800929
R41558 DVSS.n22885 DVSS.n453 0.800929
R41559 DVSS.n20985 DVSS.n20984 0.800919
R41560 DVSS.n21439 DVSS.n21438 0.800919
R41561 DVSS.n18526 DVSS.n15146 0.769676
R41562 DVSS.n19916 DVSS.n15140 0.769676
R41563 DVSS.n19192 DVSS.n19191 0.766266
R41564 DVSS.n14845 DVSS.n14844 0.764199
R41565 DVSS.n17786 DVSS.n17785 0.763161
R41566 DVSS.n18173 DVSS.n18172 0.763161
R41567 DVSS.n19903 DVSS.n19003 0.753658
R41568 DVSS.n13104 DVSS.n12354 0.7505
R41569 DVSS.n12752 DVSS.n12344 0.7505
R41570 DVSS.n12749 DVSS.n12349 0.7505
R41571 DVSS.n12759 DVSS.n12345 0.7505
R41572 DVSS.n6665 DVSS.n6248 0.7505
R41573 DVSS.n6659 DVSS.n6243 0.7505
R41574 DVSS.n6663 DVSS.n6662 0.7505
R41575 DVSS.n6660 DVSS.n6244 0.7505
R41576 DVSS.n16934 DVSS.n16928 0.743357
R41577 DVSS.n17525 DVSS.n16928 0.743357
R41578 DVSS.n17381 DVSS.n16975 0.743357
R41579 DVSS.n17484 DVSS.n16975 0.743357
R41580 DVSS.n17485 DVSS.n17052 0.743357
R41581 DVSS.n17485 DVSS.n17484 0.743357
R41582 DVSS.n17524 DVSS.n17523 0.743357
R41583 DVSS.n17525 DVSS.n17524 0.743357
R41584 DVSS.n17117 DVSS.n17054 0.743357
R41585 DVSS.n17484 DVSS.n17054 0.743357
R41586 DVSS.n17527 DVSS.n17526 0.743357
R41587 DVSS.n17526 DVSS.n17525 0.743357
R41588 DVSS.n16932 DVSS.n16927 0.743357
R41589 DVSS.n17525 DVSS.n16927 0.743357
R41590 DVSS.n17483 DVSS.n17482 0.743357
R41591 DVSS.n17484 DVSS.n17483 0.743357
R41592 DVSS.n18166 DVSS.n15535 0.739761
R41593 DVSS.n17793 DVSS.n17792 0.739479
R41594 DVSS.n19197 DVSS.n19196 0.735895
R41595 DVSS.n21440 DVSS.n21439 0.721313
R41596 DVSS.n20469 DVSS.n20468 0.686775
R41597 DVSS.n18996 DVSS.n18587 0.685361
R41598 DVSS.n18167 DVSS.n15534 0.680043
R41599 DVSS.n19927 DVSS.n19926 0.680043
R41600 DVSS.n17791 DVSS.n15919 0.679786
R41601 DVSS.n18516 DVSS.n18497 0.679786
R41602 DVSS.n22971 DVSS.n22970 0.667713
R41603 DVSS.n21473 DVSS.n21472 0.667713
R41604 DVSS.n21162 DVSS.n13681 0.661953
R41605 DVSS.n19212 DVSS.n19211 0.650781
R41606 DVSS.n19208 DVSS.n19174 0.650781
R41607 DVSS.n19194 DVSS.n19185 0.650781
R41608 DVSS.n19213 DVSS.n19209 0.650642
R41609 DVSS.n19195 DVSS.n19183 0.650642
R41610 DVSS.n13663 DVSS.n734 0.645111
R41611 DVSS.n18163 DVSS.n18162 0.64349
R41612 DVSS.n21444 DVSS.n13366 0.64349
R41613 DVSS.n19198 DVSS.n19182 0.641169
R41614 DVSS.n17791 DVSS.n17790 0.640826
R41615 DVSS.n18168 DVSS.n18167 0.640249
R41616 DVSS.n19213 DVSS.n19212 0.610577
R41617 DVSS.n18162 DVSS.n15539 0.599112
R41618 DVSS.n21445 DVSS.n21444 0.599112
R41619 DVSS.n21013 DVSS.n21010 0.596931
R41620 DVSS.n19207 DVSS.n19175 0.585639
R41621 DVSS.n19211 DVSS.n19210 0.585514
R41622 DVSS.n19174 DVSS.n19173 0.585514
R41623 DVSS.n19188 DVSS.n19187 0.585514
R41624 DVSS.n19185 DVSS.n19184 0.585514
R41625 DVSS.n19195 DVSS.n19194 0.578395
R41626 DVSS.n14579 DVSS 0.557375
R41627 DVSS.n14579 DVSS 0.557375
R41628 DVSS.n14623 DVSS 0.557375
R41629 DVSS.n14623 DVSS 0.557375
R41630 DVSS.n20640 DVSS 0.557375
R41631 DVSS.n20640 DVSS 0.557375
R41632 DVSS.n19194 DVSS.n19193 0.547605
R41633 DVSS.n19198 DVSS.n19197 0.515144
R41634 DVSS.n17793 DVSS.n15916 0.505984
R41635 DVSS.n18001 DVSS.n15535 0.505984
R41636 DVSS.n17798 DVSS.n17797 0.5005
R41637 DVSS.n17799 DVSS.n15915 0.5005
R41638 DVSS.n17802 DVSS.n17800 0.5005
R41639 DVSS.n17804 DVSS.n15913 0.5005
R41640 DVSS.n17807 DVSS.n17806 0.5005
R41641 DVSS.n17808 DVSS.n15912 0.5005
R41642 DVSS.n17811 DVSS.n17809 0.5005
R41643 DVSS.n17813 DVSS.n15910 0.5005
R41644 DVSS.n17816 DVSS.n17815 0.5005
R41645 DVSS.n17817 DVSS.n15909 0.5005
R41646 DVSS.n17819 DVSS.n17818 0.5005
R41647 DVSS.n15877 DVSS.n15876 0.5005
R41648 DVSS.n17826 DVSS.n17825 0.5005
R41649 DVSS.n17827 DVSS.n15875 0.5005
R41650 DVSS.n17830 DVSS.n17829 0.5005
R41651 DVSS.n17828 DVSS.n15873 0.5005
R41652 DVSS.n17834 DVSS.n15872 0.5005
R41653 DVSS.n17837 DVSS.n17836 0.5005
R41654 DVSS.n17838 DVSS.n15871 0.5005
R41655 DVSS.n17841 DVSS.n17839 0.5005
R41656 DVSS.n17843 DVSS.n15869 0.5005
R41657 DVSS.n17846 DVSS.n17845 0.5005
R41658 DVSS.n17847 DVSS.n15868 0.5005
R41659 DVSS.n17850 DVSS.n17848 0.5005
R41660 DVSS.n17852 DVSS.n15866 0.5005
R41661 DVSS.n17855 DVSS.n17854 0.5005
R41662 DVSS.n17856 DVSS.n15865 0.5005
R41663 DVSS.n17858 DVSS.n17857 0.5005
R41664 DVSS.n15835 DVSS.n15834 0.5005
R41665 DVSS.n17868 DVSS.n17867 0.5005
R41666 DVSS.n17869 DVSS.n15833 0.5005
R41667 DVSS.n17872 DVSS.n17871 0.5005
R41668 DVSS.n17870 DVSS.n15830 0.5005
R41669 DVSS.n17876 DVSS.n15831 0.5005
R41670 DVSS.n17878 DVSS.n15829 0.5005
R41671 DVSS.n17881 DVSS.n17880 0.5005
R41672 DVSS.n17882 DVSS.n15828 0.5005
R41673 DVSS.n17885 DVSS.n17883 0.5005
R41674 DVSS.n17887 DVSS.n15826 0.5005
R41675 DVSS.n17890 DVSS.n17889 0.5005
R41676 DVSS.n17891 DVSS.n15825 0.5005
R41677 DVSS.n17894 DVSS.n17892 0.5005
R41678 DVSS.n17896 DVSS.n15823 0.5005
R41679 DVSS.n17899 DVSS.n17898 0.5005
R41680 DVSS.n17900 DVSS.n15822 0.5005
R41681 DVSS.n17904 DVSS.n17901 0.5005
R41682 DVSS.n17903 DVSS.n17902 0.5005
R41683 DVSS.n15784 DVSS.n15783 0.5005
R41684 DVSS.n17912 DVSS.n17911 0.5005
R41685 DVSS.n17913 DVSS.n15782 0.5005
R41686 DVSS.n17916 DVSS.n17915 0.5005
R41687 DVSS.n17914 DVSS.n15780 0.5005
R41688 DVSS.n17920 DVSS.n15779 0.5005
R41689 DVSS.n17923 DVSS.n17922 0.5005
R41690 DVSS.n17924 DVSS.n15778 0.5005
R41691 DVSS.n17927 DVSS.n17925 0.5005
R41692 DVSS.n17929 DVSS.n15776 0.5005
R41693 DVSS.n17932 DVSS.n17931 0.5005
R41694 DVSS.n17933 DVSS.n15775 0.5005
R41695 DVSS.n17936 DVSS.n17934 0.5005
R41696 DVSS.n17938 DVSS.n15773 0.5005
R41697 DVSS.n17941 DVSS.n17940 0.5005
R41698 DVSS.n17942 DVSS.n15772 0.5005
R41699 DVSS.n17944 DVSS.n17943 0.5005
R41700 DVSS.n15737 DVSS.n15736 0.5005
R41701 DVSS.n17952 DVSS.n17951 0.5005
R41702 DVSS.n17953 DVSS.n15735 0.5005
R41703 DVSS.n17956 DVSS.n17955 0.5005
R41704 DVSS.n17954 DVSS.n15732 0.5005
R41705 DVSS.n17960 DVSS.n15733 0.5005
R41706 DVSS.n17962 DVSS.n15731 0.5005
R41707 DVSS.n17965 DVSS.n17964 0.5005
R41708 DVSS.n17966 DVSS.n15730 0.5005
R41709 DVSS.n17969 DVSS.n17967 0.5005
R41710 DVSS.n17971 DVSS.n15728 0.5005
R41711 DVSS.n17974 DVSS.n17973 0.5005
R41712 DVSS.n17975 DVSS.n15727 0.5005
R41713 DVSS.n18042 DVSS.n17976 0.5005
R41714 DVSS.n18041 DVSS.n17977 0.5005
R41715 DVSS.n18039 DVSS.n17978 0.5005
R41716 DVSS.n18037 DVSS.n17979 0.5005
R41717 DVSS.n18035 DVSS.n17980 0.5005
R41718 DVSS.n18033 DVSS.n17981 0.5005
R41719 DVSS.n18032 DVSS.n17982 0.5005
R41720 DVSS.n18031 DVSS.n17983 0.5005
R41721 DVSS.n17986 DVSS.n17984 0.5005
R41722 DVSS.n18027 DVSS.n17987 0.5005
R41723 DVSS.n18026 DVSS.n17988 0.5005
R41724 DVSS.n18025 DVSS.n17989 0.5005
R41725 DVSS.n18023 DVSS.n17990 0.5005
R41726 DVSS.n18021 DVSS.n17991 0.5005
R41727 DVSS.n18019 DVSS.n17992 0.5005
R41728 DVSS.n18017 DVSS.n17993 0.5005
R41729 DVSS.n18015 DVSS.n17994 0.5005
R41730 DVSS.n18013 DVSS.n17995 0.5005
R41731 DVSS.n18011 DVSS.n17996 0.5005
R41732 DVSS.n18009 DVSS.n17997 0.5005
R41733 DVSS.n18007 DVSS.n17998 0.5005
R41734 DVSS.n18005 DVSS.n17999 0.5005
R41735 DVSS.n18003 DVSS.n18000 0.5005
R41736 DVSS.n18002 DVSS.n15570 0.5005
R41737 DVSS.n17795 DVSS.n17794 0.5005
R41738 DVSS.n17797 DVSS.n17796 0.5005
R41739 DVSS.n15915 DVSS.n15914 0.5005
R41740 DVSS.n17802 DVSS.n17801 0.5005
R41741 DVSS.n17804 DVSS.n17803 0.5005
R41742 DVSS.n17806 DVSS.n17805 0.5005
R41743 DVSS.n15912 DVSS.n15911 0.5005
R41744 DVSS.n17811 DVSS.n17810 0.5005
R41745 DVSS.n17813 DVSS.n17812 0.5005
R41746 DVSS.n17815 DVSS.n17814 0.5005
R41747 DVSS.n15909 DVSS.n15908 0.5005
R41748 DVSS.n17820 DVSS.n17819 0.5005
R41749 DVSS.n15878 DVSS.n15877 0.5005
R41750 DVSS.n17825 DVSS.n17824 0.5005
R41751 DVSS.n15875 DVSS.n15874 0.5005
R41752 DVSS.n17831 DVSS.n17830 0.5005
R41753 DVSS.n17832 DVSS.n15873 0.5005
R41754 DVSS.n17834 DVSS.n17833 0.5005
R41755 DVSS.n17836 DVSS.n17835 0.5005
R41756 DVSS.n15871 DVSS.n15870 0.5005
R41757 DVSS.n17841 DVSS.n17840 0.5005
R41758 DVSS.n17843 DVSS.n17842 0.5005
R41759 DVSS.n17845 DVSS.n17844 0.5005
R41760 DVSS.n15868 DVSS.n15867 0.5005
R41761 DVSS.n17850 DVSS.n17849 0.5005
R41762 DVSS.n17852 DVSS.n17851 0.5005
R41763 DVSS.n17854 DVSS.n17853 0.5005
R41764 DVSS.n15865 DVSS.n15864 0.5005
R41765 DVSS.n17859 DVSS.n17858 0.5005
R41766 DVSS.n17861 DVSS.n15835 0.5005
R41767 DVSS.n17867 DVSS.n17866 0.5005
R41768 DVSS.n15833 DVSS.n15832 0.5005
R41769 DVSS.n17873 DVSS.n17872 0.5005
R41770 DVSS.n17874 DVSS.n15830 0.5005
R41771 DVSS.n17876 DVSS.n17875 0.5005
R41772 DVSS.n17878 DVSS.n17877 0.5005
R41773 DVSS.n17880 DVSS.n17879 0.5005
R41774 DVSS.n15828 DVSS.n15827 0.5005
R41775 DVSS.n17885 DVSS.n17884 0.5005
R41776 DVSS.n17887 DVSS.n17886 0.5005
R41777 DVSS.n17889 DVSS.n17888 0.5005
R41778 DVSS.n15825 DVSS.n15824 0.5005
R41779 DVSS.n17894 DVSS.n17893 0.5005
R41780 DVSS.n17896 DVSS.n17895 0.5005
R41781 DVSS.n17898 DVSS.n17897 0.5005
R41782 DVSS.n15822 DVSS.n15821 0.5005
R41783 DVSS.n17905 DVSS.n17904 0.5005
R41784 DVSS.n17903 DVSS.n15785 0.5005
R41785 DVSS.n17909 DVSS.n15784 0.5005
R41786 DVSS.n17911 DVSS.n17910 0.5005
R41787 DVSS.n15782 DVSS.n15781 0.5005
R41788 DVSS.n17917 DVSS.n17916 0.5005
R41789 DVSS.n17918 DVSS.n15780 0.5005
R41790 DVSS.n17920 DVSS.n17919 0.5005
R41791 DVSS.n17922 DVSS.n17921 0.5005
R41792 DVSS.n15778 DVSS.n15777 0.5005
R41793 DVSS.n17927 DVSS.n17926 0.5005
R41794 DVSS.n17929 DVSS.n17928 0.5005
R41795 DVSS.n17931 DVSS.n17930 0.5005
R41796 DVSS.n15775 DVSS.n15774 0.5005
R41797 DVSS.n17936 DVSS.n17935 0.5005
R41798 DVSS.n17938 DVSS.n17937 0.5005
R41799 DVSS.n17940 DVSS.n17939 0.5005
R41800 DVSS.n15772 DVSS.n15771 0.5005
R41801 DVSS.n17945 DVSS.n17944 0.5005
R41802 DVSS.n17946 DVSS.n15737 0.5005
R41803 DVSS.n17951 DVSS.n17950 0.5005
R41804 DVSS.n15735 DVSS.n15734 0.5005
R41805 DVSS.n17957 DVSS.n17956 0.5005
R41806 DVSS.n17958 DVSS.n15732 0.5005
R41807 DVSS.n17960 DVSS.n17959 0.5005
R41808 DVSS.n17962 DVSS.n17961 0.5005
R41809 DVSS.n17964 DVSS.n17963 0.5005
R41810 DVSS.n15730 DVSS.n15729 0.5005
R41811 DVSS.n17969 DVSS.n17968 0.5005
R41812 DVSS.n17971 DVSS.n17970 0.5005
R41813 DVSS.n17973 DVSS.n17972 0.5005
R41814 DVSS.n15727 DVSS.n15726 0.5005
R41815 DVSS.n18043 DVSS.n18042 0.5005
R41816 DVSS.n18041 DVSS.n18040 0.5005
R41817 DVSS.n18039 DVSS.n18038 0.5005
R41818 DVSS.n18037 DVSS.n18036 0.5005
R41819 DVSS.n18035 DVSS.n18034 0.5005
R41820 DVSS.n18033 DVSS.n15703 0.5005
R41821 DVSS.n18032 DVSS.n15708 0.5005
R41822 DVSS.n18031 DVSS.n18030 0.5005
R41823 DVSS.n18029 DVSS.n17984 0.5005
R41824 DVSS.n18028 DVSS.n18027 0.5005
R41825 DVSS.n18026 DVSS.n17985 0.5005
R41826 DVSS.n18025 DVSS.n18024 0.5005
R41827 DVSS.n18023 DVSS.n18022 0.5005
R41828 DVSS.n18021 DVSS.n18020 0.5005
R41829 DVSS.n18019 DVSS.n18018 0.5005
R41830 DVSS.n18017 DVSS.n18016 0.5005
R41831 DVSS.n18015 DVSS.n18014 0.5005
R41832 DVSS.n18013 DVSS.n18012 0.5005
R41833 DVSS.n18011 DVSS.n18010 0.5005
R41834 DVSS.n18009 DVSS.n18008 0.5005
R41835 DVSS.n18007 DVSS.n18006 0.5005
R41836 DVSS.n18005 DVSS.n18004 0.5005
R41837 DVSS.n18003 DVSS.n15563 0.5005
R41838 DVSS.n19215 DVSS.n19214 0.5005
R41839 DVSS.n22639 DVSS.n22638 0.455549
R41840 DVSS.n22884 DVSS.n22883 0.455549
R41841 DVSS.n16567 DVSS.n15919 0.455549
R41842 DVSS.n16739 DVSS.n15534 0.455549
R41843 DVSS.n17784 DVSS.n17783 0.455549
R41844 DVSS.n18177 DVSS.n18174 0.455549
R41845 DVSS.n17722 DVSS.n17719 0.455549
R41846 DVSS.n18251 DVSS.n18248 0.455549
R41847 DVSS.n18497 DVSS.n18496 0.455549
R41848 DVSS.n19930 DVSS.n19927 0.455549
R41849 DVSS.n21152 DVSS.n21151 0.455549
R41850 DVSS.n20983 DVSS.n20982 0.455549
R41851 DVSS.n21180 DVSS.n13658 0.455549
R41852 DVSS.n21437 DVSS.n21436 0.455549
R41853 DVSS.n22882 DVSS.n22881 0.4505
R41854 DVSS.n457 DVSS.n456 0.4505
R41855 DVSS.n22872 DVSS.n22871 0.4505
R41856 DVSS.n22870 DVSS.n22869 0.4505
R41857 DVSS.n22868 DVSS.n484 0.4505
R41858 DVSS.n22866 DVSS.n22864 0.4505
R41859 DVSS.n22863 DVSS.n486 0.4505
R41860 DVSS.n22862 DVSS.n22861 0.4505
R41861 DVSS.n22859 DVSS.n487 0.4505
R41862 DVSS.n22857 DVSS.n22855 0.4505
R41863 DVSS.n22854 DVSS.n489 0.4505
R41864 DVSS.n22853 DVSS.n22852 0.4505
R41865 DVSS.n22850 DVSS.n490 0.4505
R41866 DVSS.n22844 DVSS.n491 0.4505
R41867 DVSS.n22846 DVSS.n22845 0.4505
R41868 DVSS.n22843 DVSS.n493 0.4505
R41869 DVSS.n22842 DVSS.n22841 0.4505
R41870 DVSS.n495 DVSS.n494 0.4505
R41871 DVSS.n22835 DVSS.n22834 0.4505
R41872 DVSS.n22669 DVSS.n22668 0.4505
R41873 DVSS.n22667 DVSS.n732 0.4505
R41874 DVSS.n22666 DVSS.n22665 0.4505
R41875 DVSS.n22663 DVSS.n22640 0.4505
R41876 DVSS.n22661 DVSS.n22659 0.4505
R41877 DVSS.n22658 DVSS.n22642 0.4505
R41878 DVSS.n22657 DVSS.n22656 0.4505
R41879 DVSS.n22654 DVSS.n22643 0.4505
R41880 DVSS.n22652 DVSS.n22650 0.4505
R41881 DVSS.n22649 DVSS.n22645 0.4505
R41882 DVSS.n22648 DVSS.n22647 0.4505
R41883 DVSS.n700 DVSS.n699 0.4505
R41884 DVSS.n22676 DVSS.n22675 0.4505
R41885 DVSS.n22677 DVSS.n698 0.4505
R41886 DVSS.n22680 DVSS.n22679 0.4505
R41887 DVSS.n22678 DVSS.n696 0.4505
R41888 DVSS.n22684 DVSS.n695 0.4505
R41889 DVSS.n22687 DVSS.n22686 0.4505
R41890 DVSS.n22688 DVSS.n694 0.4505
R41891 DVSS.n22691 DVSS.n22689 0.4505
R41892 DVSS.n22693 DVSS.n692 0.4505
R41893 DVSS.n22696 DVSS.n22695 0.4505
R41894 DVSS.n22697 DVSS.n691 0.4505
R41895 DVSS.n22700 DVSS.n22698 0.4505
R41896 DVSS.n22702 DVSS.n689 0.4505
R41897 DVSS.n22705 DVSS.n22704 0.4505
R41898 DVSS.n22706 DVSS.n688 0.4505
R41899 DVSS.n22708 DVSS.n22707 0.4505
R41900 DVSS.n647 DVSS.n646 0.4505
R41901 DVSS.n22718 DVSS.n22717 0.4505
R41902 DVSS.n22719 DVSS.n645 0.4505
R41903 DVSS.n22722 DVSS.n22721 0.4505
R41904 DVSS.n22720 DVSS.n642 0.4505
R41905 DVSS.n22726 DVSS.n643 0.4505
R41906 DVSS.n22728 DVSS.n641 0.4505
R41907 DVSS.n22731 DVSS.n22730 0.4505
R41908 DVSS.n22732 DVSS.n640 0.4505
R41909 DVSS.n22735 DVSS.n22733 0.4505
R41910 DVSS.n22737 DVSS.n638 0.4505
R41911 DVSS.n22740 DVSS.n22739 0.4505
R41912 DVSS.n22741 DVSS.n637 0.4505
R41913 DVSS.n22744 DVSS.n22742 0.4505
R41914 DVSS.n22746 DVSS.n635 0.4505
R41915 DVSS.n22749 DVSS.n22748 0.4505
R41916 DVSS.n22750 DVSS.n633 0.4505
R41917 DVSS.n22753 DVSS.n22752 0.4505
R41918 DVSS.n22751 DVSS.n634 0.4505
R41919 DVSS.n595 DVSS.n594 0.4505
R41920 DVSS.n22761 DVSS.n22760 0.4505
R41921 DVSS.n22762 DVSS.n593 0.4505
R41922 DVSS.n22765 DVSS.n22764 0.4505
R41923 DVSS.n22763 DVSS.n591 0.4505
R41924 DVSS.n22769 DVSS.n590 0.4505
R41925 DVSS.n22772 DVSS.n22771 0.4505
R41926 DVSS.n22773 DVSS.n589 0.4505
R41927 DVSS.n22776 DVSS.n22774 0.4505
R41928 DVSS.n22778 DVSS.n587 0.4505
R41929 DVSS.n22781 DVSS.n22780 0.4505
R41930 DVSS.n22782 DVSS.n586 0.4505
R41931 DVSS.n22785 DVSS.n22783 0.4505
R41932 DVSS.n22787 DVSS.n584 0.4505
R41933 DVSS.n22790 DVSS.n22789 0.4505
R41934 DVSS.n22791 DVSS.n583 0.4505
R41935 DVSS.n22793 DVSS.n22792 0.4505
R41936 DVSS.n546 DVSS.n545 0.4505
R41937 DVSS.n22801 DVSS.n22800 0.4505
R41938 DVSS.n22802 DVSS.n544 0.4505
R41939 DVSS.n22805 DVSS.n22804 0.4505
R41940 DVSS.n22803 DVSS.n541 0.4505
R41941 DVSS.n22809 DVSS.n542 0.4505
R41942 DVSS.n22811 DVSS.n540 0.4505
R41943 DVSS.n22814 DVSS.n22813 0.4505
R41944 DVSS.n22815 DVSS.n539 0.4505
R41945 DVSS.n22818 DVSS.n22816 0.4505
R41946 DVSS.n22820 DVSS.n537 0.4505
R41947 DVSS.n22823 DVSS.n22822 0.4505
R41948 DVSS.n22824 DVSS.n536 0.4505
R41949 DVSS.n22827 DVSS.n22825 0.4505
R41950 DVSS.n22829 DVSS.n534 0.4505
R41951 DVSS.n22832 DVSS.n22831 0.4505
R41952 DVSS.n22833 DVSS.n533 0.4505
R41953 DVSS.n16740 DVSS.n16737 0.4505
R41954 DVSS.n16743 DVSS.n16741 0.4505
R41955 DVSS.n16745 DVSS.n16736 0.4505
R41956 DVSS.n16748 DVSS.n16747 0.4505
R41957 DVSS.n16749 DVSS.n16735 0.4505
R41958 DVSS.n16752 DVSS.n16750 0.4505
R41959 DVSS.n16754 DVSS.n16733 0.4505
R41960 DVSS.n16757 DVSS.n16756 0.4505
R41961 DVSS.n16758 DVSS.n16732 0.4505
R41962 DVSS.n16761 DVSS.n16759 0.4505
R41963 DVSS.n16763 DVSS.n16730 0.4505
R41964 DVSS.n16766 DVSS.n16765 0.4505
R41965 DVSS.n16767 DVSS.n16729 0.4505
R41966 DVSS.n16769 DVSS.n16768 0.4505
R41967 DVSS.n16727 DVSS.n16726 0.4505
R41968 DVSS.n16774 DVSS.n16773 0.4505
R41969 DVSS.n16775 DVSS.n16725 0.4505
R41970 DVSS.n16777 DVSS.n16776 0.4505
R41971 DVSS.n16779 DVSS.n16724 0.4505
R41972 DVSS.n16572 DVSS.n16571 0.4505
R41973 DVSS.n16573 DVSS.n16566 0.4505
R41974 DVSS.n16576 DVSS.n16574 0.4505
R41975 DVSS.n16578 DVSS.n16564 0.4505
R41976 DVSS.n16581 DVSS.n16580 0.4505
R41977 DVSS.n16582 DVSS.n16563 0.4505
R41978 DVSS.n16585 DVSS.n16583 0.4505
R41979 DVSS.n16587 DVSS.n16561 0.4505
R41980 DVSS.n16590 DVSS.n16589 0.4505
R41981 DVSS.n16591 DVSS.n16560 0.4505
R41982 DVSS.n16593 DVSS.n16592 0.4505
R41983 DVSS.n16333 DVSS.n16332 0.4505
R41984 DVSS.n16600 DVSS.n16599 0.4505
R41985 DVSS.n16601 DVSS.n16331 0.4505
R41986 DVSS.n16604 DVSS.n16603 0.4505
R41987 DVSS.n16602 DVSS.n16329 0.4505
R41988 DVSS.n16608 DVSS.n16328 0.4505
R41989 DVSS.n16611 DVSS.n16610 0.4505
R41990 DVSS.n16612 DVSS.n16327 0.4505
R41991 DVSS.n16615 DVSS.n16613 0.4505
R41992 DVSS.n16617 DVSS.n16325 0.4505
R41993 DVSS.n16620 DVSS.n16619 0.4505
R41994 DVSS.n16621 DVSS.n16324 0.4505
R41995 DVSS.n16624 DVSS.n16622 0.4505
R41996 DVSS.n16626 DVSS.n16322 0.4505
R41997 DVSS.n16629 DVSS.n16628 0.4505
R41998 DVSS.n16630 DVSS.n16321 0.4505
R41999 DVSS.n16632 DVSS.n16631 0.4505
R42000 DVSS.n16291 DVSS.n16290 0.4505
R42001 DVSS.n16642 DVSS.n16641 0.4505
R42002 DVSS.n16643 DVSS.n16289 0.4505
R42003 DVSS.n16646 DVSS.n16645 0.4505
R42004 DVSS.n16644 DVSS.n16286 0.4505
R42005 DVSS.n16650 DVSS.n16287 0.4505
R42006 DVSS.n16652 DVSS.n16285 0.4505
R42007 DVSS.n16655 DVSS.n16654 0.4505
R42008 DVSS.n16656 DVSS.n16284 0.4505
R42009 DVSS.n16659 DVSS.n16657 0.4505
R42010 DVSS.n16661 DVSS.n16282 0.4505
R42011 DVSS.n16664 DVSS.n16663 0.4505
R42012 DVSS.n16665 DVSS.n16281 0.4505
R42013 DVSS.n16668 DVSS.n16666 0.4505
R42014 DVSS.n16670 DVSS.n16279 0.4505
R42015 DVSS.n16673 DVSS.n16672 0.4505
R42016 DVSS.n16674 DVSS.n16277 0.4505
R42017 DVSS.n16677 DVSS.n16676 0.4505
R42018 DVSS.n16675 DVSS.n16278 0.4505
R42019 DVSS.n16240 DVSS.n16239 0.4505
R42020 DVSS.n16685 DVSS.n16684 0.4505
R42021 DVSS.n16686 DVSS.n16238 0.4505
R42022 DVSS.n16688 DVSS.n16687 0.4505
R42023 DVSS.n16236 DVSS.n16235 0.4505
R42024 DVSS.n16693 DVSS.n16692 0.4505
R42025 DVSS.n16694 DVSS.n16234 0.4505
R42026 DVSS.n16697 DVSS.n16695 0.4505
R42027 DVSS.n16699 DVSS.n16232 0.4505
R42028 DVSS.n16702 DVSS.n16701 0.4505
R42029 DVSS.n16703 DVSS.n16231 0.4505
R42030 DVSS.n16706 DVSS.n16704 0.4505
R42031 DVSS.n16708 DVSS.n16229 0.4505
R42032 DVSS.n16711 DVSS.n16710 0.4505
R42033 DVSS.n16712 DVSS.n16226 0.4505
R42034 DVSS.n16820 DVSS.n16819 0.4505
R42035 DVSS.n16818 DVSS.n16228 0.4505
R42036 DVSS.n16817 DVSS.n16816 0.4505
R42037 DVSS.n16814 DVSS.n16713 0.4505
R42038 DVSS.n16813 DVSS.n16812 0.4505
R42039 DVSS.n16811 DVSS.n16714 0.4505
R42040 DVSS.n16810 DVSS.n16809 0.4505
R42041 DVSS.n16805 DVSS.n16715 0.4505
R42042 DVSS.n16804 DVSS.n16802 0.4505
R42043 DVSS.n16801 DVSS.n16717 0.4505
R42044 DVSS.n16800 DVSS.n16799 0.4505
R42045 DVSS.n16797 DVSS.n16718 0.4505
R42046 DVSS.n16795 DVSS.n16793 0.4505
R42047 DVSS.n16792 DVSS.n16720 0.4505
R42048 DVSS.n16791 DVSS.n16790 0.4505
R42049 DVSS.n16788 DVSS.n16721 0.4505
R42050 DVSS.n16786 DVSS.n16784 0.4505
R42051 DVSS.n16783 DVSS.n16723 0.4505
R42052 DVSS.n16782 DVSS.n16781 0.4505
R42053 DVSS.n16738 DVSS.n15613 0.4505
R42054 DVSS.n16737 DVSS.n15608 0.4505
R42055 DVSS.n16743 DVSS.n16742 0.4505
R42056 DVSS.n16745 DVSS.n16744 0.4505
R42057 DVSS.n16747 DVSS.n16746 0.4505
R42058 DVSS.n16735 DVSS.n16734 0.4505
R42059 DVSS.n16752 DVSS.n16751 0.4505
R42060 DVSS.n16754 DVSS.n16753 0.4505
R42061 DVSS.n16756 DVSS.n16755 0.4505
R42062 DVSS.n16732 DVSS.n16731 0.4505
R42063 DVSS.n16761 DVSS.n16760 0.4505
R42064 DVSS.n16763 DVSS.n16762 0.4505
R42065 DVSS.n16765 DVSS.n16764 0.4505
R42066 DVSS.n16729 DVSS.n16728 0.4505
R42067 DVSS.n16770 DVSS.n16769 0.4505
R42068 DVSS.n16771 DVSS.n16727 0.4505
R42069 DVSS.n16773 DVSS.n16772 0.4505
R42070 DVSS.n16725 DVSS.n15673 0.4505
R42071 DVSS.n16777 DVSS.n15668 0.4505
R42072 DVSS.n16779 DVSS.n16778 0.4505
R42073 DVSS.n16569 DVSS.n16568 0.4505
R42074 DVSS.n16571 DVSS.n16570 0.4505
R42075 DVSS.n16566 DVSS.n16565 0.4505
R42076 DVSS.n16576 DVSS.n16575 0.4505
R42077 DVSS.n16578 DVSS.n16577 0.4505
R42078 DVSS.n16580 DVSS.n16579 0.4505
R42079 DVSS.n16563 DVSS.n16562 0.4505
R42080 DVSS.n16585 DVSS.n16584 0.4505
R42081 DVSS.n16587 DVSS.n16586 0.4505
R42082 DVSS.n16589 DVSS.n16588 0.4505
R42083 DVSS.n16560 DVSS.n16559 0.4505
R42084 DVSS.n16594 DVSS.n16593 0.4505
R42085 DVSS.n16334 DVSS.n16333 0.4505
R42086 DVSS.n16599 DVSS.n16598 0.4505
R42087 DVSS.n16331 DVSS.n16330 0.4505
R42088 DVSS.n16605 DVSS.n16604 0.4505
R42089 DVSS.n16606 DVSS.n16329 0.4505
R42090 DVSS.n16608 DVSS.n16607 0.4505
R42091 DVSS.n16610 DVSS.n16609 0.4505
R42092 DVSS.n16327 DVSS.n16326 0.4505
R42093 DVSS.n16615 DVSS.n16614 0.4505
R42094 DVSS.n16617 DVSS.n16616 0.4505
R42095 DVSS.n16619 DVSS.n16618 0.4505
R42096 DVSS.n16324 DVSS.n16323 0.4505
R42097 DVSS.n16624 DVSS.n16623 0.4505
R42098 DVSS.n16626 DVSS.n16625 0.4505
R42099 DVSS.n16628 DVSS.n16627 0.4505
R42100 DVSS.n16321 DVSS.n16320 0.4505
R42101 DVSS.n16633 DVSS.n16632 0.4505
R42102 DVSS.n16635 DVSS.n16291 0.4505
R42103 DVSS.n16641 DVSS.n16640 0.4505
R42104 DVSS.n16289 DVSS.n16288 0.4505
R42105 DVSS.n16647 DVSS.n16646 0.4505
R42106 DVSS.n16648 DVSS.n16286 0.4505
R42107 DVSS.n16650 DVSS.n16649 0.4505
R42108 DVSS.n16652 DVSS.n16651 0.4505
R42109 DVSS.n16654 DVSS.n16653 0.4505
R42110 DVSS.n16284 DVSS.n16283 0.4505
R42111 DVSS.n16659 DVSS.n16658 0.4505
R42112 DVSS.n16661 DVSS.n16660 0.4505
R42113 DVSS.n16663 DVSS.n16662 0.4505
R42114 DVSS.n16281 DVSS.n16280 0.4505
R42115 DVSS.n16668 DVSS.n16667 0.4505
R42116 DVSS.n16670 DVSS.n16669 0.4505
R42117 DVSS.n16672 DVSS.n16671 0.4505
R42118 DVSS.n16277 DVSS.n16276 0.4505
R42119 DVSS.n16678 DVSS.n16677 0.4505
R42120 DVSS.n16278 DVSS.n16241 0.4505
R42121 DVSS.n16682 DVSS.n16240 0.4505
R42122 DVSS.n16684 DVSS.n16683 0.4505
R42123 DVSS.n16238 DVSS.n16237 0.4505
R42124 DVSS.n16689 DVSS.n16688 0.4505
R42125 DVSS.n16690 DVSS.n16236 0.4505
R42126 DVSS.n16692 DVSS.n16691 0.4505
R42127 DVSS.n16234 DVSS.n16233 0.4505
R42128 DVSS.n16697 DVSS.n16696 0.4505
R42129 DVSS.n16699 DVSS.n16698 0.4505
R42130 DVSS.n16701 DVSS.n16700 0.4505
R42131 DVSS.n16231 DVSS.n16230 0.4505
R42132 DVSS.n16706 DVSS.n16705 0.4505
R42133 DVSS.n16708 DVSS.n16707 0.4505
R42134 DVSS.n16710 DVSS.n16709 0.4505
R42135 DVSS.n16226 DVSS.n16225 0.4505
R42136 DVSS.n16821 DVSS.n16820 0.4505
R42137 DVSS.n16228 DVSS.n16227 0.4505
R42138 DVSS.n16816 DVSS.n16815 0.4505
R42139 DVSS.n16814 DVSS.n16165 0.4505
R42140 DVSS.n16813 DVSS.n16171 0.4505
R42141 DVSS.n16806 DVSS.n16714 0.4505
R42142 DVSS.n16809 DVSS.n16808 0.4505
R42143 DVSS.n16807 DVSS.n16805 0.4505
R42144 DVSS.n16804 DVSS.n16803 0.4505
R42145 DVSS.n16717 DVSS.n16716 0.4505
R42146 DVSS.n16799 DVSS.n16798 0.4505
R42147 DVSS.n16797 DVSS.n16796 0.4505
R42148 DVSS.n16795 DVSS.n16794 0.4505
R42149 DVSS.n16720 DVSS.n16719 0.4505
R42150 DVSS.n16790 DVSS.n16789 0.4505
R42151 DVSS.n16788 DVSS.n16787 0.4505
R42152 DVSS.n16786 DVSS.n16785 0.4505
R42153 DVSS.n16723 DVSS.n16722 0.4505
R42154 DVSS.n16781 DVSS.n16780 0.4505
R42155 DVSS.n18178 DVSS.n15531 0.4505
R42156 DVSS.n18181 DVSS.n18179 0.4505
R42157 DVSS.n18184 DVSS.n18183 0.4505
R42158 DVSS.n18185 DVSS.n15529 0.4505
R42159 DVSS.n18188 DVSS.n18186 0.4505
R42160 DVSS.n18190 DVSS.n15527 0.4505
R42161 DVSS.n18193 DVSS.n18192 0.4505
R42162 DVSS.n18194 DVSS.n15525 0.4505
R42163 DVSS.n18196 DVSS.n18195 0.4505
R42164 DVSS.n15526 DVSS.n15523 0.4505
R42165 DVSS.n17566 DVSS.n17564 0.4505
R42166 DVSS.n17567 DVSS.n17563 0.4505
R42167 DVSS.n17569 DVSS.n17568 0.4505
R42168 DVSS.n17570 DVSS.n17561 0.4505
R42169 DVSS.n17572 DVSS.n17571 0.4505
R42170 DVSS.n17562 DVSS.n17558 0.4505
R42171 DVSS.n17576 DVSS.n17559 0.4505
R42172 DVSS.n17578 DVSS.n17557 0.4505
R42173 DVSS.n17581 DVSS.n17580 0.4505
R42174 DVSS.n17782 DVSS.n17781 0.4505
R42175 DVSS.n15925 DVSS.n15924 0.4505
R42176 DVSS.n15971 DVSS.n15969 0.4505
R42177 DVSS.n15974 DVSS.n15973 0.4505
R42178 DVSS.n15975 DVSS.n15968 0.4505
R42179 DVSS.n15978 DVSS.n15976 0.4505
R42180 DVSS.n15980 DVSS.n15966 0.4505
R42181 DVSS.n15983 DVSS.n15982 0.4505
R42182 DVSS.n15984 DVSS.n15963 0.4505
R42183 DVSS.n17671 DVSS.n17670 0.4505
R42184 DVSS.n17669 DVSS.n15965 0.4505
R42185 DVSS.n17668 DVSS.n17667 0.4505
R42186 DVSS.n17666 DVSS.n15985 0.4505
R42187 DVSS.n17665 DVSS.n15987 0.4505
R42188 DVSS.n15990 DVSS.n15986 0.4505
R42189 DVSS.n17661 DVSS.n17660 0.4505
R42190 DVSS.n17659 DVSS.n15989 0.4505
R42191 DVSS.n17658 DVSS.n17657 0.4505
R42192 DVSS.n15992 DVSS.n15991 0.4505
R42193 DVSS.n16042 DVSS.n16040 0.4505
R42194 DVSS.n16045 DVSS.n16044 0.4505
R42195 DVSS.n16046 DVSS.n16039 0.4505
R42196 DVSS.n16049 DVSS.n16047 0.4505
R42197 DVSS.n16051 DVSS.n16037 0.4505
R42198 DVSS.n16054 DVSS.n16053 0.4505
R42199 DVSS.n16055 DVSS.n16036 0.4505
R42200 DVSS.n16058 DVSS.n16056 0.4505
R42201 DVSS.n16060 DVSS.n16034 0.4505
R42202 DVSS.n16063 DVSS.n16062 0.4505
R42203 DVSS.n16064 DVSS.n16032 0.4505
R42204 DVSS.n17651 DVSS.n17650 0.4505
R42205 DVSS.n17649 DVSS.n16033 0.4505
R42206 DVSS.n17648 DVSS.n17647 0.4505
R42207 DVSS.n16066 DVSS.n16065 0.4505
R42208 DVSS.n16113 DVSS.n16112 0.4505
R42209 DVSS.n16116 DVSS.n16114 0.4505
R42210 DVSS.n16118 DVSS.n16111 0.4505
R42211 DVSS.n16121 DVSS.n16120 0.4505
R42212 DVSS.n16122 DVSS.n16110 0.4505
R42213 DVSS.n16125 DVSS.n16123 0.4505
R42214 DVSS.n16127 DVSS.n16108 0.4505
R42215 DVSS.n16130 DVSS.n16129 0.4505
R42216 DVSS.n16131 DVSS.n16105 0.4505
R42217 DVSS.n17638 DVSS.n17637 0.4505
R42218 DVSS.n17636 DVSS.n16107 0.4505
R42219 DVSS.n17635 DVSS.n17634 0.4505
R42220 DVSS.n17632 DVSS.n16132 0.4505
R42221 DVSS.n17631 DVSS.n17630 0.4505
R42222 DVSS.n17629 DVSS.n16133 0.4505
R42223 DVSS.n17628 DVSS.n17627 0.4505
R42224 DVSS.n16135 DVSS.n16134 0.4505
R42225 DVSS.n17623 DVSS.n17622 0.4505
R42226 DVSS.n17621 DVSS.n16138 0.4505
R42227 DVSS.n17620 DVSS.n17619 0.4505
R42228 DVSS.n16140 DVSS.n16139 0.4505
R42229 DVSS.n16864 DVSS.n16862 0.4505
R42230 DVSS.n16867 DVSS.n16866 0.4505
R42231 DVSS.n16868 DVSS.n16861 0.4505
R42232 DVSS.n16871 DVSS.n16869 0.4505
R42233 DVSS.n16873 DVSS.n16859 0.4505
R42234 DVSS.n16876 DVSS.n16875 0.4505
R42235 DVSS.n16877 DVSS.n16858 0.4505
R42236 DVSS.n16880 DVSS.n16878 0.4505
R42237 DVSS.n16882 DVSS.n16856 0.4505
R42238 DVSS.n16885 DVSS.n16884 0.4505
R42239 DVSS.n16886 DVSS.n16854 0.4505
R42240 DVSS.n17613 DVSS.n17612 0.4505
R42241 DVSS.n17611 DVSS.n16855 0.4505
R42242 DVSS.n17610 DVSS.n17609 0.4505
R42243 DVSS.n16888 DVSS.n16887 0.4505
R42244 DVSS.n17550 DVSS.n17547 0.4505
R42245 DVSS.n17602 DVSS.n17601 0.4505
R42246 DVSS.n17600 DVSS.n17549 0.4505
R42247 DVSS.n17599 DVSS.n17598 0.4505
R42248 DVSS.n17596 DVSS.n17551 0.4505
R42249 DVSS.n17594 DVSS.n17592 0.4505
R42250 DVSS.n17591 DVSS.n17553 0.4505
R42251 DVSS.n17590 DVSS.n17589 0.4505
R42252 DVSS.n17587 DVSS.n17554 0.4505
R42253 DVSS.n17585 DVSS.n17583 0.4505
R42254 DVSS.n17582 DVSS.n17556 0.4505
R42255 DVSS.n18176 DVSS.n18175 0.4505
R42256 DVSS.n15531 DVSS.n15530 0.4505
R42257 DVSS.n18181 DVSS.n18180 0.4505
R42258 DVSS.n18183 DVSS.n18182 0.4505
R42259 DVSS.n15529 DVSS.n15528 0.4505
R42260 DVSS.n18188 DVSS.n18187 0.4505
R42261 DVSS.n18190 DVSS.n18189 0.4505
R42262 DVSS.n18192 DVSS.n18191 0.4505
R42263 DVSS.n15525 DVSS.n15524 0.4505
R42264 DVSS.n18197 DVSS.n18196 0.4505
R42265 DVSS.n15523 DVSS.n15522 0.4505
R42266 DVSS.n17566 DVSS.n17565 0.4505
R42267 DVSS.n17567 DVSS.n15511 0.4505
R42268 DVSS.n17568 DVSS.n15505 0.4505
R42269 DVSS.n17561 DVSS.n17560 0.4505
R42270 DVSS.n17573 DVSS.n17572 0.4505
R42271 DVSS.n17574 DVSS.n17558 0.4505
R42272 DVSS.n17576 DVSS.n17575 0.4505
R42273 DVSS.n17578 DVSS.n17577 0.4505
R42274 DVSS.n17580 DVSS.n17579 0.4505
R42275 DVSS.n15923 DVSS.n15922 0.4505
R42276 DVSS.n17781 DVSS.n17780 0.4505
R42277 DVSS.n15948 DVSS.n15925 0.4505
R42278 DVSS.n15971 DVSS.n15970 0.4505
R42279 DVSS.n15973 DVSS.n15972 0.4505
R42280 DVSS.n15968 DVSS.n15967 0.4505
R42281 DVSS.n15978 DVSS.n15977 0.4505
R42282 DVSS.n15980 DVSS.n15979 0.4505
R42283 DVSS.n15982 DVSS.n15981 0.4505
R42284 DVSS.n15963 DVSS.n15958 0.4505
R42285 DVSS.n17672 DVSS.n17671 0.4505
R42286 DVSS.n15965 DVSS.n15964 0.4505
R42287 DVSS.n17667 DVSS.n15955 0.4505
R42288 DVSS.n17666 DVSS.n15956 0.4505
R42289 DVSS.n17665 DVSS.n17664 0.4505
R42290 DVSS.n17663 DVSS.n15986 0.4505
R42291 DVSS.n17662 DVSS.n17661 0.4505
R42292 DVSS.n15989 DVSS.n15988 0.4505
R42293 DVSS.n17657 DVSS.n17656 0.4505
R42294 DVSS.n15999 DVSS.n15992 0.4505
R42295 DVSS.n16042 DVSS.n16041 0.4505
R42296 DVSS.n16044 DVSS.n16043 0.4505
R42297 DVSS.n16039 DVSS.n16038 0.4505
R42298 DVSS.n16049 DVSS.n16048 0.4505
R42299 DVSS.n16051 DVSS.n16050 0.4505
R42300 DVSS.n16053 DVSS.n16052 0.4505
R42301 DVSS.n16036 DVSS.n16035 0.4505
R42302 DVSS.n16058 DVSS.n16057 0.4505
R42303 DVSS.n16060 DVSS.n16059 0.4505
R42304 DVSS.n16062 DVSS.n16061 0.4505
R42305 DVSS.n16032 DVSS.n16030 0.4505
R42306 DVSS.n17652 DVSS.n17651 0.4505
R42307 DVSS.n16033 DVSS.n16031 0.4505
R42308 DVSS.n17647 DVSS.n17646 0.4505
R42309 DVSS.n17645 DVSS.n16066 0.4505
R42310 DVSS.n16112 DVSS.n16073 0.4505
R42311 DVSS.n16116 DVSS.n16115 0.4505
R42312 DVSS.n16118 DVSS.n16117 0.4505
R42313 DVSS.n16120 DVSS.n16119 0.4505
R42314 DVSS.n16110 DVSS.n16109 0.4505
R42315 DVSS.n16125 DVSS.n16124 0.4505
R42316 DVSS.n16127 DVSS.n16126 0.4505
R42317 DVSS.n16129 DVSS.n16128 0.4505
R42318 DVSS.n16105 DVSS.n16104 0.4505
R42319 DVSS.n17639 DVSS.n17638 0.4505
R42320 DVSS.n16107 DVSS.n16106 0.4505
R42321 DVSS.n17634 DVSS.n17633 0.4505
R42322 DVSS.n17632 DVSS.n16087 0.4505
R42323 DVSS.n17631 DVSS.n16093 0.4505
R42324 DVSS.n16136 DVSS.n16133 0.4505
R42325 DVSS.n17627 DVSS.n17626 0.4505
R42326 DVSS.n17625 DVSS.n16135 0.4505
R42327 DVSS.n17624 DVSS.n17623 0.4505
R42328 DVSS.n16138 DVSS.n16137 0.4505
R42329 DVSS.n17619 DVSS.n17618 0.4505
R42330 DVSS.n16147 DVSS.n16140 0.4505
R42331 DVSS.n16864 DVSS.n16863 0.4505
R42332 DVSS.n16866 DVSS.n16865 0.4505
R42333 DVSS.n16861 DVSS.n16860 0.4505
R42334 DVSS.n16871 DVSS.n16870 0.4505
R42335 DVSS.n16873 DVSS.n16872 0.4505
R42336 DVSS.n16875 DVSS.n16874 0.4505
R42337 DVSS.n16858 DVSS.n16857 0.4505
R42338 DVSS.n16880 DVSS.n16879 0.4505
R42339 DVSS.n16882 DVSS.n16881 0.4505
R42340 DVSS.n16884 DVSS.n16883 0.4505
R42341 DVSS.n16854 DVSS.n16852 0.4505
R42342 DVSS.n17614 DVSS.n17613 0.4505
R42343 DVSS.n16855 DVSS.n16853 0.4505
R42344 DVSS.n17609 DVSS.n17608 0.4505
R42345 DVSS.n17607 DVSS.n16888 0.4505
R42346 DVSS.n17547 DVSS.n16894 0.4505
R42347 DVSS.n17603 DVSS.n17602 0.4505
R42348 DVSS.n17549 DVSS.n17548 0.4505
R42349 DVSS.n17598 DVSS.n17597 0.4505
R42350 DVSS.n17596 DVSS.n17595 0.4505
R42351 DVSS.n17594 DVSS.n17593 0.4505
R42352 DVSS.n17553 DVSS.n17552 0.4505
R42353 DVSS.n17589 DVSS.n17588 0.4505
R42354 DVSS.n17587 DVSS.n17586 0.4505
R42355 DVSS.n17585 DVSS.n17584 0.4505
R42356 DVSS.n17556 DVSS.n17555 0.4505
R42357 DVSS.n18252 DVSS.n18247 0.4505
R42358 DVSS.n18255 DVSS.n18253 0.4505
R42359 DVSS.n18257 DVSS.n18245 0.4505
R42360 DVSS.n18260 DVSS.n18259 0.4505
R42361 DVSS.n18261 DVSS.n18244 0.4505
R42362 DVSS.n18264 DVSS.n18262 0.4505
R42363 DVSS.n18266 DVSS.n18242 0.4505
R42364 DVSS.n18269 DVSS.n18268 0.4505
R42365 DVSS.n18270 DVSS.n18240 0.4505
R42366 DVSS.n18272 DVSS.n18271 0.4505
R42367 DVSS.n18241 DVSS.n18238 0.4505
R42368 DVSS.n15484 DVSS.n15483 0.4505
R42369 DVSS.n18279 DVSS.n18278 0.4505
R42370 DVSS.n18280 DVSS.n15481 0.4505
R42371 DVSS.n18282 DVSS.n18281 0.4505
R42372 DVSS.n15482 DVSS.n15478 0.4505
R42373 DVSS.n18286 DVSS.n15479 0.4505
R42374 DVSS.n18288 DVSS.n15477 0.4505
R42375 DVSS.n18291 DVSS.n18290 0.4505
R42376 DVSS.n17723 DVSS.n17718 0.4505
R42377 DVSS.n17726 DVSS.n17724 0.4505
R42378 DVSS.n17728 DVSS.n17716 0.4505
R42379 DVSS.n17731 DVSS.n17730 0.4505
R42380 DVSS.n17732 DVSS.n17715 0.4505
R42381 DVSS.n17735 DVSS.n17733 0.4505
R42382 DVSS.n17737 DVSS.n17713 0.4505
R42383 DVSS.n17740 DVSS.n17739 0.4505
R42384 DVSS.n17741 DVSS.n17710 0.4505
R42385 DVSS.n17769 DVSS.n17768 0.4505
R42386 DVSS.n17767 DVSS.n17712 0.4505
R42387 DVSS.n17766 DVSS.n17765 0.4505
R42388 DVSS.n17764 DVSS.n17742 0.4505
R42389 DVSS.n17763 DVSS.n17744 0.4505
R42390 DVSS.n17747 DVSS.n17743 0.4505
R42391 DVSS.n17759 DVSS.n17758 0.4505
R42392 DVSS.n17757 DVSS.n17746 0.4505
R42393 DVSS.n17756 DVSS.n17755 0.4505
R42394 DVSS.n17753 DVSS.n17748 0.4505
R42395 DVSS.n17751 DVSS.n17749 0.4505
R42396 DVSS.n15278 DVSS.n15275 0.4505
R42397 DVSS.n18376 DVSS.n18375 0.4505
R42398 DVSS.n18374 DVSS.n15277 0.4505
R42399 DVSS.n18373 DVSS.n18372 0.4505
R42400 DVSS.n18370 DVSS.n15279 0.4505
R42401 DVSS.n18368 DVSS.n18366 0.4505
R42402 DVSS.n18365 DVSS.n15281 0.4505
R42403 DVSS.n18364 DVSS.n18363 0.4505
R42404 DVSS.n18361 DVSS.n15282 0.4505
R42405 DVSS.n18359 DVSS.n18358 0.4505
R42406 DVSS.n18357 DVSS.n15283 0.4505
R42407 DVSS.n18356 DVSS.n18355 0.4505
R42408 DVSS.n15285 DVSS.n15284 0.4505
R42409 DVSS.n18351 DVSS.n18350 0.4505
R42410 DVSS.n18349 DVSS.n15287 0.4505
R42411 DVSS.n18348 DVSS.n18347 0.4505
R42412 DVSS.n15289 DVSS.n15288 0.4505
R42413 DVSS.n15336 DVSS.n15335 0.4505
R42414 DVSS.n15337 DVSS.n15333 0.4505
R42415 DVSS.n15340 DVSS.n15338 0.4505
R42416 DVSS.n15342 DVSS.n15331 0.4505
R42417 DVSS.n15345 DVSS.n15344 0.4505
R42418 DVSS.n15346 DVSS.n15330 0.4505
R42419 DVSS.n15349 DVSS.n15347 0.4505
R42420 DVSS.n15351 DVSS.n15328 0.4505
R42421 DVSS.n15354 DVSS.n15353 0.4505
R42422 DVSS.n15355 DVSS.n15326 0.4505
R42423 DVSS.n18341 DVSS.n18340 0.4505
R42424 DVSS.n18339 DVSS.n15327 0.4505
R42425 DVSS.n18338 DVSS.n18337 0.4505
R42426 DVSS.n15357 DVSS.n15356 0.4505
R42427 DVSS.n18333 DVSS.n18332 0.4505
R42428 DVSS.n18331 DVSS.n15359 0.4505
R42429 DVSS.n18330 DVSS.n18329 0.4505
R42430 DVSS.n15361 DVSS.n15360 0.4505
R42431 DVSS.n15408 DVSS.n15406 0.4505
R42432 DVSS.n15411 DVSS.n15410 0.4505
R42433 DVSS.n15412 DVSS.n15405 0.4505
R42434 DVSS.n15415 DVSS.n15413 0.4505
R42435 DVSS.n15417 DVSS.n15403 0.4505
R42436 DVSS.n15420 DVSS.n15419 0.4505
R42437 DVSS.n15421 DVSS.n15402 0.4505
R42438 DVSS.n15424 DVSS.n15422 0.4505
R42439 DVSS.n15426 DVSS.n15400 0.4505
R42440 DVSS.n15429 DVSS.n15428 0.4505
R42441 DVSS.n15430 DVSS.n15398 0.4505
R42442 DVSS.n18323 DVSS.n18322 0.4505
R42443 DVSS.n18321 DVSS.n15399 0.4505
R42444 DVSS.n18320 DVSS.n18319 0.4505
R42445 DVSS.n15432 DVSS.n15431 0.4505
R42446 DVSS.n15470 DVSS.n15467 0.4505
R42447 DVSS.n18312 DVSS.n18311 0.4505
R42448 DVSS.n18310 DVSS.n15469 0.4505
R42449 DVSS.n18309 DVSS.n18308 0.4505
R42450 DVSS.n18306 DVSS.n15471 0.4505
R42451 DVSS.n18304 DVSS.n18302 0.4505
R42452 DVSS.n18301 DVSS.n15473 0.4505
R42453 DVSS.n18300 DVSS.n18299 0.4505
R42454 DVSS.n18297 DVSS.n15474 0.4505
R42455 DVSS.n18295 DVSS.n18293 0.4505
R42456 DVSS.n18292 DVSS.n15476 0.4505
R42457 DVSS.n18250 DVSS.n18249 0.4505
R42458 DVSS.n18247 DVSS.n18246 0.4505
R42459 DVSS.n18255 DVSS.n18254 0.4505
R42460 DVSS.n18257 DVSS.n18256 0.4505
R42461 DVSS.n18259 DVSS.n18258 0.4505
R42462 DVSS.n18244 DVSS.n18243 0.4505
R42463 DVSS.n18264 DVSS.n18263 0.4505
R42464 DVSS.n18266 DVSS.n18265 0.4505
R42465 DVSS.n18268 DVSS.n18267 0.4505
R42466 DVSS.n18240 DVSS.n18239 0.4505
R42467 DVSS.n18273 DVSS.n18272 0.4505
R42468 DVSS.n18238 DVSS.n18232 0.4505
R42469 DVSS.n15490 DVSS.n15484 0.4505
R42470 DVSS.n18278 DVSS.n18277 0.4505
R42471 DVSS.n15481 DVSS.n15480 0.4505
R42472 DVSS.n18283 DVSS.n18282 0.4505
R42473 DVSS.n18284 DVSS.n15478 0.4505
R42474 DVSS.n18286 DVSS.n18285 0.4505
R42475 DVSS.n18288 DVSS.n18287 0.4505
R42476 DVSS.n18290 DVSS.n18289 0.4505
R42477 DVSS.n17721 DVSS.n17720 0.4505
R42478 DVSS.n17718 DVSS.n17717 0.4505
R42479 DVSS.n17726 DVSS.n17725 0.4505
R42480 DVSS.n17728 DVSS.n17727 0.4505
R42481 DVSS.n17730 DVSS.n17729 0.4505
R42482 DVSS.n17715 DVSS.n17714 0.4505
R42483 DVSS.n17735 DVSS.n17734 0.4505
R42484 DVSS.n17737 DVSS.n17736 0.4505
R42485 DVSS.n17739 DVSS.n17738 0.4505
R42486 DVSS.n17710 DVSS.n17706 0.4505
R42487 DVSS.n17770 DVSS.n17769 0.4505
R42488 DVSS.n17712 DVSS.n17711 0.4505
R42489 DVSS.n17765 DVSS.n17691 0.4505
R42490 DVSS.n17764 DVSS.n17698 0.4505
R42491 DVSS.n17763 DVSS.n17762 0.4505
R42492 DVSS.n17761 DVSS.n17743 0.4505
R42493 DVSS.n17760 DVSS.n17759 0.4505
R42494 DVSS.n17746 DVSS.n17745 0.4505
R42495 DVSS.n17755 DVSS.n17754 0.4505
R42496 DVSS.n17753 DVSS.n17752 0.4505
R42497 DVSS.n17751 DVSS.n17750 0.4505
R42498 DVSS.n15275 DVSS.n15274 0.4505
R42499 DVSS.n18377 DVSS.n18376 0.4505
R42500 DVSS.n15277 DVSS.n15276 0.4505
R42501 DVSS.n18372 DVSS.n18371 0.4505
R42502 DVSS.n18370 DVSS.n18369 0.4505
R42503 DVSS.n18368 DVSS.n18367 0.4505
R42504 DVSS.n15281 DVSS.n15280 0.4505
R42505 DVSS.n18363 DVSS.n18362 0.4505
R42506 DVSS.n18361 DVSS.n18360 0.4505
R42507 DVSS.n18359 DVSS.n15253 0.4505
R42508 DVSS.n15283 DVSS.n15259 0.4505
R42509 DVSS.n18355 DVSS.n18354 0.4505
R42510 DVSS.n18353 DVSS.n15285 0.4505
R42511 DVSS.n18352 DVSS.n18351 0.4505
R42512 DVSS.n15290 DVSS.n15287 0.4505
R42513 DVSS.n18347 DVSS.n18346 0.4505
R42514 DVSS.n15298 DVSS.n15289 0.4505
R42515 DVSS.n15335 DVSS.n15334 0.4505
R42516 DVSS.n15333 DVSS.n15332 0.4505
R42517 DVSS.n15340 DVSS.n15339 0.4505
R42518 DVSS.n15342 DVSS.n15341 0.4505
R42519 DVSS.n15344 DVSS.n15343 0.4505
R42520 DVSS.n15330 DVSS.n15329 0.4505
R42521 DVSS.n15349 DVSS.n15348 0.4505
R42522 DVSS.n15351 DVSS.n15350 0.4505
R42523 DVSS.n15353 DVSS.n15352 0.4505
R42524 DVSS.n15326 DVSS.n15324 0.4505
R42525 DVSS.n18342 DVSS.n18341 0.4505
R42526 DVSS.n15327 DVSS.n15325 0.4505
R42527 DVSS.n18337 DVSS.n18336 0.4505
R42528 DVSS.n18335 DVSS.n15357 0.4505
R42529 DVSS.n18334 DVSS.n18333 0.4505
R42530 DVSS.n15359 DVSS.n15358 0.4505
R42531 DVSS.n18329 DVSS.n18328 0.4505
R42532 DVSS.n15368 DVSS.n15361 0.4505
R42533 DVSS.n15408 DVSS.n15407 0.4505
R42534 DVSS.n15410 DVSS.n15409 0.4505
R42535 DVSS.n15405 DVSS.n15404 0.4505
R42536 DVSS.n15415 DVSS.n15414 0.4505
R42537 DVSS.n15417 DVSS.n15416 0.4505
R42538 DVSS.n15419 DVSS.n15418 0.4505
R42539 DVSS.n15402 DVSS.n15401 0.4505
R42540 DVSS.n15424 DVSS.n15423 0.4505
R42541 DVSS.n15426 DVSS.n15425 0.4505
R42542 DVSS.n15428 DVSS.n15427 0.4505
R42543 DVSS.n15398 DVSS.n15396 0.4505
R42544 DVSS.n18324 DVSS.n18323 0.4505
R42545 DVSS.n15399 DVSS.n15397 0.4505
R42546 DVSS.n18319 DVSS.n18318 0.4505
R42547 DVSS.n18317 DVSS.n15432 0.4505
R42548 DVSS.n15467 DVSS.n15438 0.4505
R42549 DVSS.n18313 DVSS.n18312 0.4505
R42550 DVSS.n15469 DVSS.n15468 0.4505
R42551 DVSS.n18308 DVSS.n18307 0.4505
R42552 DVSS.n18306 DVSS.n18305 0.4505
R42553 DVSS.n18304 DVSS.n18303 0.4505
R42554 DVSS.n15473 DVSS.n15472 0.4505
R42555 DVSS.n18299 DVSS.n18298 0.4505
R42556 DVSS.n18297 DVSS.n18296 0.4505
R42557 DVSS.n18295 DVSS.n18294 0.4505
R42558 DVSS.n15476 DVSS.n15475 0.4505
R42559 DVSS.n19931 DVSS.n15125 0.4505
R42560 DVSS.n19934 DVSS.n19932 0.4505
R42561 DVSS.n19937 DVSS.n19936 0.4505
R42562 DVSS.n19938 DVSS.n15123 0.4505
R42563 DVSS.n19941 DVSS.n19939 0.4505
R42564 DVSS.n19943 DVSS.n15121 0.4505
R42565 DVSS.n19946 DVSS.n19945 0.4505
R42566 DVSS.n19947 DVSS.n15120 0.4505
R42567 DVSS.n19949 DVSS.n19948 0.4505
R42568 DVSS.n15083 DVSS.n15082 0.4505
R42569 DVSS.n19957 DVSS.n19956 0.4505
R42570 DVSS.n19958 DVSS.n15081 0.4505
R42571 DVSS.n19960 DVSS.n19959 0.4505
R42572 DVSS.n15079 DVSS.n15078 0.4505
R42573 DVSS.n19965 DVSS.n19964 0.4505
R42574 DVSS.n19966 DVSS.n15036 0.4505
R42575 DVSS.n19968 DVSS.n19967 0.4505
R42576 DVSS.n15077 DVSS.n15035 0.4505
R42577 DVSS.n15076 DVSS.n15075 0.4505
R42578 DVSS.n18495 DVSS.n18494 0.4505
R42579 DVSS.n15152 DVSS.n15151 0.4505
R42580 DVSS.n15196 DVSS.n15195 0.4505
R42581 DVSS.n15197 DVSS.n15193 0.4505
R42582 DVSS.n15200 DVSS.n15198 0.4505
R42583 DVSS.n15202 DVSS.n15191 0.4505
R42584 DVSS.n15205 DVSS.n15204 0.4505
R42585 DVSS.n15206 DVSS.n15190 0.4505
R42586 DVSS.n15208 DVSS.n15207 0.4505
R42587 DVSS.n15216 DVSS.n15188 0.4505
R42588 DVSS.n15219 DVSS.n15218 0.4505
R42589 DVSS.n15220 DVSS.n15186 0.4505
R42590 DVSS.n18488 DVSS.n18487 0.4505
R42591 DVSS.n18486 DVSS.n15187 0.4505
R42592 DVSS.n18485 DVSS.n18484 0.4505
R42593 DVSS.n15222 DVSS.n15221 0.4505
R42594 DVSS.n18480 DVSS.n18479 0.4505
R42595 DVSS.n18478 DVSS.n15224 0.4505
R42596 DVSS.n18477 DVSS.n18476 0.4505
R42597 DVSS.n15226 DVSS.n15225 0.4505
R42598 DVSS.n18412 DVSS.n18411 0.4505
R42599 DVSS.n18413 DVSS.n18409 0.4505
R42600 DVSS.n18416 DVSS.n18414 0.4505
R42601 DVSS.n18418 DVSS.n18407 0.4505
R42602 DVSS.n18421 DVSS.n18420 0.4505
R42603 DVSS.n18422 DVSS.n18406 0.4505
R42604 DVSS.n18425 DVSS.n18423 0.4505
R42605 DVSS.n18426 DVSS.n18404 0.4505
R42606 DVSS.n18436 DVSS.n18435 0.4505
R42607 DVSS.n18437 DVSS.n18402 0.4505
R42608 DVSS.n18470 DVSS.n18469 0.4505
R42609 DVSS.n18468 DVSS.n18403 0.4505
R42610 DVSS.n18467 DVSS.n18466 0.4505
R42611 DVSS.n18463 DVSS.n18438 0.4505
R42612 DVSS.n18462 DVSS.n18460 0.4505
R42613 DVSS.n18459 DVSS.n18440 0.4505
R42614 DVSS.n18458 DVSS.n18457 0.4505
R42615 DVSS.n18455 DVSS.n18441 0.4505
R42616 DVSS.n18453 DVSS.n18451 0.4505
R42617 DVSS.n18450 DVSS.n18443 0.4505
R42618 DVSS.n18449 DVSS.n18448 0.4505
R42619 DVSS.n18446 DVSS.n18444 0.4505
R42620 DVSS.n14917 DVSS.n14914 0.4505
R42621 DVSS.n20004 DVSS.n20003 0.4505
R42622 DVSS.n20002 DVSS.n14916 0.4505
R42623 DVSS.n20001 DVSS.n20000 0.4505
R42624 DVSS.n19998 DVSS.n14918 0.4505
R42625 DVSS.n19997 DVSS.n19996 0.4505
R42626 DVSS.n19995 DVSS.n14919 0.4505
R42627 DVSS.n19994 DVSS.n19993 0.4505
R42628 DVSS.n14921 DVSS.n14920 0.4505
R42629 DVSS.n19989 DVSS.n19988 0.4505
R42630 DVSS.n19987 DVSS.n14924 0.4505
R42631 DVSS.n19986 DVSS.n19985 0.4505
R42632 DVSS.n14926 DVSS.n14925 0.4505
R42633 DVSS.n14970 DVSS.n14968 0.4505
R42634 DVSS.n14973 DVSS.n14972 0.4505
R42635 DVSS.n14974 DVSS.n14967 0.4505
R42636 DVSS.n14977 DVSS.n14975 0.4505
R42637 DVSS.n14979 DVSS.n14965 0.4505
R42638 DVSS.n14982 DVSS.n14981 0.4505
R42639 DVSS.n14983 DVSS.n14964 0.4505
R42640 DVSS.n14986 DVSS.n14984 0.4505
R42641 DVSS.n14994 DVSS.n14962 0.4505
R42642 DVSS.n14997 DVSS.n14996 0.4505
R42643 DVSS.n14998 DVSS.n14960 0.4505
R42644 DVSS.n19979 DVSS.n19978 0.4505
R42645 DVSS.n19977 DVSS.n14961 0.4505
R42646 DVSS.n19976 DVSS.n19975 0.4505
R42647 DVSS.n15000 DVSS.n14999 0.4505
R42648 DVSS.n15045 DVSS.n15044 0.4505
R42649 DVSS.n15048 DVSS.n15046 0.4505
R42650 DVSS.n15050 DVSS.n15043 0.4505
R42651 DVSS.n15053 DVSS.n15052 0.4505
R42652 DVSS.n15054 DVSS.n15042 0.4505
R42653 DVSS.n15057 DVSS.n15055 0.4505
R42654 DVSS.n15059 DVSS.n15040 0.4505
R42655 DVSS.n15062 DVSS.n15061 0.4505
R42656 DVSS.n15063 DVSS.n15039 0.4505
R42657 DVSS.n15065 DVSS.n15064 0.4505
R42658 DVSS.n15073 DVSS.n15037 0.4505
R42659 DVSS.n19929 DVSS.n19928 0.4505
R42660 DVSS.n15125 DVSS.n15124 0.4505
R42661 DVSS.n19934 DVSS.n19933 0.4505
R42662 DVSS.n19936 DVSS.n19935 0.4505
R42663 DVSS.n15123 DVSS.n15122 0.4505
R42664 DVSS.n19941 DVSS.n19940 0.4505
R42665 DVSS.n19943 DVSS.n19942 0.4505
R42666 DVSS.n19945 DVSS.n19944 0.4505
R42667 DVSS.n15120 DVSS.n15119 0.4505
R42668 DVSS.n19950 DVSS.n19949 0.4505
R42669 DVSS.n15091 DVSS.n15083 0.4505
R42670 DVSS.n19956 DVSS.n19955 0.4505
R42671 DVSS.n15084 DVSS.n15081 0.4505
R42672 DVSS.n19961 DVSS.n19960 0.4505
R42673 DVSS.n19962 DVSS.n15079 0.4505
R42674 DVSS.n19964 DVSS.n19963 0.4505
R42675 DVSS.n15036 DVSS.n15034 0.4505
R42676 DVSS.n19969 DVSS.n19968 0.4505
R42677 DVSS.n15035 DVSS.n15033 0.4505
R42678 DVSS.n15075 DVSS.n15074 0.4505
R42679 DVSS.n15150 DVSS.n15149 0.4505
R42680 DVSS.n18494 DVSS.n18493 0.4505
R42681 DVSS.n15176 DVSS.n15152 0.4505
R42682 DVSS.n15195 DVSS.n15194 0.4505
R42683 DVSS.n15193 DVSS.n15192 0.4505
R42684 DVSS.n15200 DVSS.n15199 0.4505
R42685 DVSS.n15202 DVSS.n15201 0.4505
R42686 DVSS.n15204 DVSS.n15203 0.4505
R42687 DVSS.n15190 DVSS.n15189 0.4505
R42688 DVSS.n15209 DVSS.n15208 0.4505
R42689 DVSS.n15216 DVSS.n15215 0.4505
R42690 DVSS.n15218 DVSS.n15217 0.4505
R42691 DVSS.n15186 DVSS.n15184 0.4505
R42692 DVSS.n18489 DVSS.n18488 0.4505
R42693 DVSS.n15187 DVSS.n15185 0.4505
R42694 DVSS.n18484 DVSS.n18483 0.4505
R42695 DVSS.n18482 DVSS.n15222 0.4505
R42696 DVSS.n18481 DVSS.n18480 0.4505
R42697 DVSS.n15227 DVSS.n15224 0.4505
R42698 DVSS.n18476 DVSS.n18475 0.4505
R42699 DVSS.n15234 DVSS.n15226 0.4505
R42700 DVSS.n18411 DVSS.n18410 0.4505
R42701 DVSS.n18409 DVSS.n18408 0.4505
R42702 DVSS.n18416 DVSS.n18415 0.4505
R42703 DVSS.n18418 DVSS.n18417 0.4505
R42704 DVSS.n18420 DVSS.n18419 0.4505
R42705 DVSS.n18406 DVSS.n18405 0.4505
R42706 DVSS.n18425 DVSS.n18424 0.4505
R42707 DVSS.n18427 DVSS.n18426 0.4505
R42708 DVSS.n18435 DVSS.n18434 0.4505
R42709 DVSS.n18402 DVSS.n18400 0.4505
R42710 DVSS.n18471 DVSS.n18470 0.4505
R42711 DVSS.n18403 DVSS.n18401 0.4505
R42712 DVSS.n18466 DVSS.n18465 0.4505
R42713 DVSS.n18464 DVSS.n18463 0.4505
R42714 DVSS.n18462 DVSS.n18461 0.4505
R42715 DVSS.n18440 DVSS.n18439 0.4505
R42716 DVSS.n18457 DVSS.n18456 0.4505
R42717 DVSS.n18455 DVSS.n18454 0.4505
R42718 DVSS.n18453 DVSS.n18452 0.4505
R42719 DVSS.n18443 DVSS.n18442 0.4505
R42720 DVSS.n18448 DVSS.n18447 0.4505
R42721 DVSS.n18446 DVSS.n18445 0.4505
R42722 DVSS.n14914 DVSS.n14913 0.4505
R42723 DVSS.n20005 DVSS.n20004 0.4505
R42724 DVSS.n14916 DVSS.n14915 0.4505
R42725 DVSS.n20000 DVSS.n19999 0.4505
R42726 DVSS.n19998 DVSS.n14888 0.4505
R42727 DVSS.n19997 DVSS.n14894 0.4505
R42728 DVSS.n14922 DVSS.n14919 0.4505
R42729 DVSS.n19993 DVSS.n19992 0.4505
R42730 DVSS.n19991 DVSS.n14921 0.4505
R42731 DVSS.n19990 DVSS.n19989 0.4505
R42732 DVSS.n14924 DVSS.n14923 0.4505
R42733 DVSS.n19985 DVSS.n19984 0.4505
R42734 DVSS.n14933 DVSS.n14926 0.4505
R42735 DVSS.n14970 DVSS.n14969 0.4505
R42736 DVSS.n14972 DVSS.n14971 0.4505
R42737 DVSS.n14967 DVSS.n14966 0.4505
R42738 DVSS.n14977 DVSS.n14976 0.4505
R42739 DVSS.n14979 DVSS.n14978 0.4505
R42740 DVSS.n14981 DVSS.n14980 0.4505
R42741 DVSS.n14964 DVSS.n14963 0.4505
R42742 DVSS.n14986 DVSS.n14985 0.4505
R42743 DVSS.n14994 DVSS.n14993 0.4505
R42744 DVSS.n14996 DVSS.n14995 0.4505
R42745 DVSS.n14960 DVSS.n14958 0.4505
R42746 DVSS.n19980 DVSS.n19979 0.4505
R42747 DVSS.n14961 DVSS.n14959 0.4505
R42748 DVSS.n19975 DVSS.n19974 0.4505
R42749 DVSS.n19973 DVSS.n15000 0.4505
R42750 DVSS.n15044 DVSS.n15006 0.4505
R42751 DVSS.n15048 DVSS.n15047 0.4505
R42752 DVSS.n15050 DVSS.n15049 0.4505
R42753 DVSS.n15052 DVSS.n15051 0.4505
R42754 DVSS.n15042 DVSS.n15041 0.4505
R42755 DVSS.n15057 DVSS.n15056 0.4505
R42756 DVSS.n15059 DVSS.n15058 0.4505
R42757 DVSS.n15061 DVSS.n15060 0.4505
R42758 DVSS.n15039 DVSS.n15038 0.4505
R42759 DVSS.n15066 DVSS.n15065 0.4505
R42760 DVSS.n15073 DVSS.n15072 0.4505
R42761 DVSS.n20981 DVSS.n20980 0.4505
R42762 DVSS.n14319 DVSS.n14318 0.4505
R42763 DVSS.n20949 DVSS.n20948 0.4505
R42764 DVSS.n20952 DVSS.n20950 0.4505
R42765 DVSS.n20954 DVSS.n20946 0.4505
R42766 DVSS.n20957 DVSS.n20956 0.4505
R42767 DVSS.n20958 DVSS.n20945 0.4505
R42768 DVSS.n20961 DVSS.n20959 0.4505
R42769 DVSS.n20962 DVSS.n20943 0.4505
R42770 DVSS.n20971 DVSS.n20970 0.4505
R42771 DVSS.n20972 DVSS.n14354 0.4505
R42772 DVSS.n20974 DVSS.n20973 0.4505
R42773 DVSS.n20942 DVSS.n14352 0.4505
R42774 DVSS.n20941 DVSS.n20940 0.4505
R42775 DVSS.n14356 DVSS.n14355 0.4505
R42776 DVSS.n20936 DVSS.n20935 0.4505
R42777 DVSS.n20934 DVSS.n14358 0.4505
R42778 DVSS.n20933 DVSS.n20932 0.4505
R42779 DVSS.n14360 DVSS.n14359 0.4505
R42780 DVSS.n21150 DVSS.n21149 0.4505
R42781 DVSS.n13690 DVSS.n13689 0.4505
R42782 DVSS.n20745 DVSS.n20743 0.4505
R42783 DVSS.n20747 DVSS.n20742 0.4505
R42784 DVSS.n20750 DVSS.n20749 0.4505
R42785 DVSS.n20751 DVSS.n20741 0.4505
R42786 DVSS.n20754 DVSS.n20752 0.4505
R42787 DVSS.n20756 DVSS.n20739 0.4505
R42788 DVSS.n20759 DVSS.n20758 0.4505
R42789 DVSS.n20760 DVSS.n20738 0.4505
R42790 DVSS.n20763 DVSS.n20761 0.4505
R42791 DVSS.n20764 DVSS.n20736 0.4505
R42792 DVSS.n20766 DVSS.n20765 0.4505
R42793 DVSS.n20767 DVSS.n20735 0.4505
R42794 DVSS.n20770 DVSS.n20769 0.4505
R42795 DVSS.n20768 DVSS.n20732 0.4505
R42796 DVSS.n20774 DVSS.n20733 0.4505
R42797 DVSS.n20776 DVSS.n20731 0.4505
R42798 DVSS.n20779 DVSS.n20778 0.4505
R42799 DVSS.n20780 DVSS.n20730 0.4505
R42800 DVSS.n20783 DVSS.n20781 0.4505
R42801 DVSS.n20785 DVSS.n20728 0.4505
R42802 DVSS.n20788 DVSS.n20787 0.4505
R42803 DVSS.n20789 DVSS.n20727 0.4505
R42804 DVSS.n20792 DVSS.n20790 0.4505
R42805 DVSS.n20794 DVSS.n20725 0.4505
R42806 DVSS.n20797 DVSS.n20796 0.4505
R42807 DVSS.n20798 DVSS.n20724 0.4505
R42808 DVSS.n20800 DVSS.n20799 0.4505
R42809 DVSS.n14505 DVSS.n14504 0.4505
R42810 DVSS.n20808 DVSS.n20807 0.4505
R42811 DVSS.n20809 DVSS.n14503 0.4505
R42812 DVSS.n20812 DVSS.n20811 0.4505
R42813 DVSS.n20810 DVSS.n14501 0.4505
R42814 DVSS.n20820 DVSS.n14500 0.4505
R42815 DVSS.n20823 DVSS.n20822 0.4505
R42816 DVSS.n20824 DVSS.n14499 0.4505
R42817 DVSS.n20827 DVSS.n20825 0.4505
R42818 DVSS.n20829 DVSS.n14497 0.4505
R42819 DVSS.n20832 DVSS.n20831 0.4505
R42820 DVSS.n20833 DVSS.n14496 0.4505
R42821 DVSS.n20836 DVSS.n20834 0.4505
R42822 DVSS.n20838 DVSS.n14494 0.4505
R42823 DVSS.n20841 DVSS.n20840 0.4505
R42824 DVSS.n20842 DVSS.n14492 0.4505
R42825 DVSS.n20845 DVSS.n20844 0.4505
R42826 DVSS.n20843 DVSS.n14493 0.4505
R42827 DVSS.n14458 DVSS.n14457 0.4505
R42828 DVSS.n20853 DVSS.n20852 0.4505
R42829 DVSS.n20854 DVSS.n14456 0.4505
R42830 DVSS.n20857 DVSS.n20856 0.4505
R42831 DVSS.n20855 DVSS.n14454 0.4505
R42832 DVSS.n20861 DVSS.n14453 0.4505
R42833 DVSS.n20864 DVSS.n20863 0.4505
R42834 DVSS.n20865 DVSS.n14452 0.4505
R42835 DVSS.n20868 DVSS.n20866 0.4505
R42836 DVSS.n20870 DVSS.n14450 0.4505
R42837 DVSS.n20873 DVSS.n20872 0.4505
R42838 DVSS.n20874 DVSS.n14449 0.4505
R42839 DVSS.n20877 DVSS.n20875 0.4505
R42840 DVSS.n20879 DVSS.n14447 0.4505
R42841 DVSS.n20882 DVSS.n20881 0.4505
R42842 DVSS.n20883 DVSS.n14446 0.4505
R42843 DVSS.n20885 DVSS.n20884 0.4505
R42844 DVSS.n14409 DVSS.n14408 0.4505
R42845 DVSS.n20893 DVSS.n20892 0.4505
R42846 DVSS.n20894 DVSS.n14407 0.4505
R42847 DVSS.n20897 DVSS.n20896 0.4505
R42848 DVSS.n20895 DVSS.n14405 0.4505
R42849 DVSS.n20901 DVSS.n14404 0.4505
R42850 DVSS.n20904 DVSS.n20903 0.4505
R42851 DVSS.n20905 DVSS.n14403 0.4505
R42852 DVSS.n20908 DVSS.n20906 0.4505
R42853 DVSS.n20910 DVSS.n14401 0.4505
R42854 DVSS.n20913 DVSS.n20912 0.4505
R42855 DVSS.n20914 DVSS.n14400 0.4505
R42856 DVSS.n20917 DVSS.n20915 0.4505
R42857 DVSS.n20919 DVSS.n14398 0.4505
R42858 DVSS.n20922 DVSS.n20921 0.4505
R42859 DVSS.n20923 DVSS.n14397 0.4505
R42860 DVSS.n20925 DVSS.n20924 0.4505
R42861 DVSS.n14317 DVSS.n14316 0.4505
R42862 DVSS.n20980 DVSS.n20979 0.4505
R42863 DVSS.n14342 DVSS.n14319 0.4505
R42864 DVSS.n20948 DVSS.n20947 0.4505
R42865 DVSS.n20952 DVSS.n20951 0.4505
R42866 DVSS.n20954 DVSS.n20953 0.4505
R42867 DVSS.n20956 DVSS.n20955 0.4505
R42868 DVSS.n20945 DVSS.n20944 0.4505
R42869 DVSS.n20961 DVSS.n20960 0.4505
R42870 DVSS.n20963 DVSS.n20962 0.4505
R42871 DVSS.n20970 DVSS.n20969 0.4505
R42872 DVSS.n14354 DVSS.n14353 0.4505
R42873 DVSS.n20975 DVSS.n20974 0.4505
R42874 DVSS.n14352 DVSS.n14351 0.4505
R42875 DVSS.n20940 DVSS.n20939 0.4505
R42876 DVSS.n20938 DVSS.n14356 0.4505
R42877 DVSS.n20937 DVSS.n20936 0.4505
R42878 DVSS.n14358 DVSS.n14357 0.4505
R42879 DVSS.n20932 DVSS.n20931 0.4505
R42880 DVSS.n20927 DVSS.n14360 0.4505
R42881 DVSS.n13688 DVSS.n13687 0.4505
R42882 DVSS.n21149 DVSS.n21148 0.4505
R42883 DVSS.n13713 DVSS.n13690 0.4505
R42884 DVSS.n20745 DVSS.n20744 0.4505
R42885 DVSS.n20747 DVSS.n20746 0.4505
R42886 DVSS.n20749 DVSS.n20748 0.4505
R42887 DVSS.n20741 DVSS.n20740 0.4505
R42888 DVSS.n20754 DVSS.n20753 0.4505
R42889 DVSS.n20756 DVSS.n20755 0.4505
R42890 DVSS.n20758 DVSS.n20757 0.4505
R42891 DVSS.n20738 DVSS.n20737 0.4505
R42892 DVSS.n20763 DVSS.n20762 0.4505
R42893 DVSS.n20764 DVSS.n13720 0.4505
R42894 DVSS.n20765 DVSS.n13721 0.4505
R42895 DVSS.n20735 DVSS.n20734 0.4505
R42896 DVSS.n20771 DVSS.n20770 0.4505
R42897 DVSS.n20772 DVSS.n20732 0.4505
R42898 DVSS.n20774 DVSS.n20773 0.4505
R42899 DVSS.n20776 DVSS.n20775 0.4505
R42900 DVSS.n20778 DVSS.n20777 0.4505
R42901 DVSS.n20730 DVSS.n20729 0.4505
R42902 DVSS.n20783 DVSS.n20782 0.4505
R42903 DVSS.n20785 DVSS.n20784 0.4505
R42904 DVSS.n20787 DVSS.n20786 0.4505
R42905 DVSS.n20727 DVSS.n20726 0.4505
R42906 DVSS.n20792 DVSS.n20791 0.4505
R42907 DVSS.n20794 DVSS.n20793 0.4505
R42908 DVSS.n20796 DVSS.n20795 0.4505
R42909 DVSS.n20724 DVSS.n20723 0.4505
R42910 DVSS.n20801 DVSS.n20800 0.4505
R42911 DVSS.n14506 DVSS.n14505 0.4505
R42912 DVSS.n20807 DVSS.n20806 0.4505
R42913 DVSS.n14503 DVSS.n14502 0.4505
R42914 DVSS.n20813 DVSS.n20812 0.4505
R42915 DVSS.n20814 DVSS.n14501 0.4505
R42916 DVSS.n20820 DVSS.n20819 0.4505
R42917 DVSS.n20822 DVSS.n20821 0.4505
R42918 DVSS.n14499 DVSS.n14498 0.4505
R42919 DVSS.n20827 DVSS.n20826 0.4505
R42920 DVSS.n20829 DVSS.n20828 0.4505
R42921 DVSS.n20831 DVSS.n20830 0.4505
R42922 DVSS.n14496 DVSS.n14495 0.4505
R42923 DVSS.n20836 DVSS.n20835 0.4505
R42924 DVSS.n20838 DVSS.n20837 0.4505
R42925 DVSS.n20840 DVSS.n20839 0.4505
R42926 DVSS.n14492 DVSS.n14491 0.4505
R42927 DVSS.n20846 DVSS.n20845 0.4505
R42928 DVSS.n14493 DVSS.n14459 0.4505
R42929 DVSS.n20850 DVSS.n14458 0.4505
R42930 DVSS.n20852 DVSS.n20851 0.4505
R42931 DVSS.n14456 DVSS.n14455 0.4505
R42932 DVSS.n20858 DVSS.n20857 0.4505
R42933 DVSS.n20859 DVSS.n14454 0.4505
R42934 DVSS.n20861 DVSS.n20860 0.4505
R42935 DVSS.n20863 DVSS.n20862 0.4505
R42936 DVSS.n14452 DVSS.n14451 0.4505
R42937 DVSS.n20868 DVSS.n20867 0.4505
R42938 DVSS.n20870 DVSS.n20869 0.4505
R42939 DVSS.n20872 DVSS.n20871 0.4505
R42940 DVSS.n14449 DVSS.n14448 0.4505
R42941 DVSS.n20877 DVSS.n20876 0.4505
R42942 DVSS.n20879 DVSS.n20878 0.4505
R42943 DVSS.n20881 DVSS.n20880 0.4505
R42944 DVSS.n14446 DVSS.n14445 0.4505
R42945 DVSS.n20886 DVSS.n20885 0.4505
R42946 DVSS.n20887 DVSS.n14409 0.4505
R42947 DVSS.n20892 DVSS.n20891 0.4505
R42948 DVSS.n14407 DVSS.n14406 0.4505
R42949 DVSS.n20898 DVSS.n20897 0.4505
R42950 DVSS.n20899 DVSS.n14405 0.4505
R42951 DVSS.n20901 DVSS.n20900 0.4505
R42952 DVSS.n20903 DVSS.n20902 0.4505
R42953 DVSS.n14403 DVSS.n14402 0.4505
R42954 DVSS.n20908 DVSS.n20907 0.4505
R42955 DVSS.n20910 DVSS.n20909 0.4505
R42956 DVSS.n20912 DVSS.n20911 0.4505
R42957 DVSS.n14400 DVSS.n14399 0.4505
R42958 DVSS.n20917 DVSS.n20916 0.4505
R42959 DVSS.n20919 DVSS.n20918 0.4505
R42960 DVSS.n20921 DVSS.n20920 0.4505
R42961 DVSS.n14397 DVSS.n14396 0.4505
R42962 DVSS.n20926 DVSS.n20925 0.4505
R42963 DVSS.n21358 DVSS.n21356 0.4505
R42964 DVSS.n21360 DVSS.n13456 0.4505
R42965 DVSS.n21363 DVSS.n21362 0.4505
R42966 DVSS.n21364 DVSS.n13455 0.4505
R42967 DVSS.n21367 DVSS.n21365 0.4505
R42968 DVSS.n21369 DVSS.n13453 0.4505
R42969 DVSS.n21372 DVSS.n21371 0.4505
R42970 DVSS.n21373 DVSS.n13452 0.4505
R42971 DVSS.n21375 DVSS.n21374 0.4505
R42972 DVSS.n13418 DVSS.n13417 0.4505
R42973 DVSS.n21387 DVSS.n21386 0.4505
R42974 DVSS.n21388 DVSS.n13416 0.4505
R42975 DVSS.n21390 DVSS.n21389 0.4505
R42976 DVSS.n13414 DVSS.n13413 0.4505
R42977 DVSS.n21395 DVSS.n21394 0.4505
R42978 DVSS.n21396 DVSS.n13410 0.4505
R42979 DVSS.n21428 DVSS.n21427 0.4505
R42980 DVSS.n21426 DVSS.n13412 0.4505
R42981 DVSS.n21425 DVSS.n21424 0.4505
R42982 DVSS.n21416 DVSS.n21397 0.4505
R42983 DVSS.n21415 DVSS.n21413 0.4505
R42984 DVSS.n21412 DVSS.n21399 0.4505
R42985 DVSS.n21411 DVSS.n21410 0.4505
R42986 DVSS.n21408 DVSS.n21400 0.4505
R42987 DVSS.n21406 DVSS.n21404 0.4505
R42988 DVSS.n21403 DVSS.n21402 0.4505
R42989 DVSS.n13376 DVSS.n13375 0.4505
R42990 DVSS.n21435 DVSS.n21434 0.4505
R42991 DVSS.n21185 DVSS.n21184 0.4505
R42992 DVSS.n21186 DVSS.n13657 0.4505
R42993 DVSS.n21189 DVSS.n21187 0.4505
R42994 DVSS.n21191 DVSS.n13655 0.4505
R42995 DVSS.n21194 DVSS.n21193 0.4505
R42996 DVSS.n21195 DVSS.n13654 0.4505
R42997 DVSS.n21198 DVSS.n21196 0.4505
R42998 DVSS.n21200 DVSS.n13652 0.4505
R42999 DVSS.n21208 DVSS.n21207 0.4505
R43000 DVSS.n21209 DVSS.n13651 0.4505
R43001 DVSS.n21211 DVSS.n21210 0.4505
R43002 DVSS.n13617 DVSS.n13616 0.4505
R43003 DVSS.n21218 DVSS.n21217 0.4505
R43004 DVSS.n21219 DVSS.n13615 0.4505
R43005 DVSS.n21222 DVSS.n21221 0.4505
R43006 DVSS.n21220 DVSS.n13613 0.4505
R43007 DVSS.n21226 DVSS.n13612 0.4505
R43008 DVSS.n21229 DVSS.n21228 0.4505
R43009 DVSS.n21230 DVSS.n13611 0.4505
R43010 DVSS.n21233 DVSS.n21231 0.4505
R43011 DVSS.n21235 DVSS.n13609 0.4505
R43012 DVSS.n21238 DVSS.n21237 0.4505
R43013 DVSS.n21239 DVSS.n13608 0.4505
R43014 DVSS.n21242 DVSS.n21240 0.4505
R43015 DVSS.n21244 DVSS.n13606 0.4505
R43016 DVSS.n21247 DVSS.n21246 0.4505
R43017 DVSS.n21248 DVSS.n13605 0.4505
R43018 DVSS.n21250 DVSS.n21249 0.4505
R43019 DVSS.n13569 DVSS.n13568 0.4505
R43020 DVSS.n21260 DVSS.n21259 0.4505
R43021 DVSS.n21261 DVSS.n13567 0.4505
R43022 DVSS.n21264 DVSS.n21263 0.4505
R43023 DVSS.n21262 DVSS.n13564 0.4505
R43024 DVSS.n21268 DVSS.n13565 0.4505
R43025 DVSS.n21270 DVSS.n13563 0.4505
R43026 DVSS.n21273 DVSS.n21272 0.4505
R43027 DVSS.n21274 DVSS.n13562 0.4505
R43028 DVSS.n21277 DVSS.n21275 0.4505
R43029 DVSS.n21279 DVSS.n13560 0.4505
R43030 DVSS.n21282 DVSS.n21281 0.4505
R43031 DVSS.n21283 DVSS.n13559 0.4505
R43032 DVSS.n21286 DVSS.n21284 0.4505
R43033 DVSS.n21288 DVSS.n13557 0.4505
R43034 DVSS.n21291 DVSS.n21290 0.4505
R43035 DVSS.n21292 DVSS.n13555 0.4505
R43036 DVSS.n21295 DVSS.n21294 0.4505
R43037 DVSS.n21293 DVSS.n13556 0.4505
R43038 DVSS.n13515 DVSS.n13514 0.4505
R43039 DVSS.n21303 DVSS.n21302 0.4505
R43040 DVSS.n21304 DVSS.n13513 0.4505
R43041 DVSS.n21307 DVSS.n21306 0.4505
R43042 DVSS.n21305 DVSS.n13511 0.4505
R43043 DVSS.n21311 DVSS.n13510 0.4505
R43044 DVSS.n21314 DVSS.n21313 0.4505
R43045 DVSS.n21315 DVSS.n13509 0.4505
R43046 DVSS.n21318 DVSS.n21316 0.4505
R43047 DVSS.n21320 DVSS.n13507 0.4505
R43048 DVSS.n21323 DVSS.n21322 0.4505
R43049 DVSS.n21324 DVSS.n13506 0.4505
R43050 DVSS.n21327 DVSS.n21325 0.4505
R43051 DVSS.n21329 DVSS.n13504 0.4505
R43052 DVSS.n21332 DVSS.n21331 0.4505
R43053 DVSS.n21333 DVSS.n13503 0.4505
R43054 DVSS.n21335 DVSS.n21334 0.4505
R43055 DVSS.n13464 DVSS.n13463 0.4505
R43056 DVSS.n21343 DVSS.n21342 0.4505
R43057 DVSS.n21344 DVSS.n13462 0.4505
R43058 DVSS.n21347 DVSS.n21346 0.4505
R43059 DVSS.n21345 DVSS.n13460 0.4505
R43060 DVSS.n21351 DVSS.n13459 0.4505
R43061 DVSS.n21354 DVSS.n21353 0.4505
R43062 DVSS.n21355 DVSS.n13458 0.4505
R43063 DVSS.n13374 DVSS.n13373 0.4505
R43064 DVSS.n21434 DVSS.n21433 0.4505
R43065 DVSS.n13400 DVSS.n13376 0.4505
R43066 DVSS.n21402 DVSS.n21401 0.4505
R43067 DVSS.n21406 DVSS.n21405 0.4505
R43068 DVSS.n21408 DVSS.n21407 0.4505
R43069 DVSS.n21410 DVSS.n21409 0.4505
R43070 DVSS.n21399 DVSS.n21398 0.4505
R43071 DVSS.n21415 DVSS.n21414 0.4505
R43072 DVSS.n21417 DVSS.n21416 0.4505
R43073 DVSS.n21424 DVSS.n21423 0.4505
R43074 DVSS.n13412 DVSS.n13411 0.4505
R43075 DVSS.n21429 DVSS.n21428 0.4505
R43076 DVSS.n13410 DVSS.n13409 0.4505
R43077 DVSS.n21394 DVSS.n21393 0.4505
R43078 DVSS.n21392 DVSS.n13414 0.4505
R43079 DVSS.n21391 DVSS.n21390 0.4505
R43080 DVSS.n13416 DVSS.n13415 0.4505
R43081 DVSS.n21386 DVSS.n21385 0.4505
R43082 DVSS.n21381 DVSS.n13418 0.4505
R43083 DVSS.n21376 DVSS.n21375 0.4505
R43084 DVSS.n13452 DVSS.n13451 0.4505
R43085 DVSS.n21371 DVSS.n21370 0.4505
R43086 DVSS.n21369 DVSS.n21368 0.4505
R43087 DVSS.n21367 DVSS.n21366 0.4505
R43088 DVSS.n13455 DVSS.n13454 0.4505
R43089 DVSS.n21362 DVSS.n21361 0.4505
R43090 DVSS.n21360 DVSS.n21359 0.4505
R43091 DVSS.n21358 DVSS.n21357 0.4505
R43092 DVSS.n21182 DVSS.n21181 0.4505
R43093 DVSS.n21184 DVSS.n21183 0.4505
R43094 DVSS.n13657 DVSS.n13656 0.4505
R43095 DVSS.n21189 DVSS.n21188 0.4505
R43096 DVSS.n21191 DVSS.n21190 0.4505
R43097 DVSS.n21193 DVSS.n21192 0.4505
R43098 DVSS.n13654 DVSS.n13653 0.4505
R43099 DVSS.n21198 DVSS.n21197 0.4505
R43100 DVSS.n21200 DVSS.n21199 0.4505
R43101 DVSS.n21207 DVSS.n21206 0.4505
R43102 DVSS.n13651 DVSS.n13650 0.4505
R43103 DVSS.n21212 DVSS.n21211 0.4505
R43104 DVSS.n13618 DVSS.n13617 0.4505
R43105 DVSS.n21217 DVSS.n21216 0.4505
R43106 DVSS.n13615 DVSS.n13614 0.4505
R43107 DVSS.n21223 DVSS.n21222 0.4505
R43108 DVSS.n21224 DVSS.n13613 0.4505
R43109 DVSS.n21226 DVSS.n21225 0.4505
R43110 DVSS.n21228 DVSS.n21227 0.4505
R43111 DVSS.n13611 DVSS.n13610 0.4505
R43112 DVSS.n21233 DVSS.n21232 0.4505
R43113 DVSS.n21235 DVSS.n21234 0.4505
R43114 DVSS.n21237 DVSS.n21236 0.4505
R43115 DVSS.n13608 DVSS.n13607 0.4505
R43116 DVSS.n21242 DVSS.n21241 0.4505
R43117 DVSS.n21244 DVSS.n21243 0.4505
R43118 DVSS.n21246 DVSS.n21245 0.4505
R43119 DVSS.n13605 DVSS.n13604 0.4505
R43120 DVSS.n21251 DVSS.n21250 0.4505
R43121 DVSS.n21253 DVSS.n13569 0.4505
R43122 DVSS.n21259 DVSS.n21258 0.4505
R43123 DVSS.n13567 DVSS.n13566 0.4505
R43124 DVSS.n21265 DVSS.n21264 0.4505
R43125 DVSS.n21266 DVSS.n13564 0.4505
R43126 DVSS.n21268 DVSS.n21267 0.4505
R43127 DVSS.n21270 DVSS.n21269 0.4505
R43128 DVSS.n21272 DVSS.n21271 0.4505
R43129 DVSS.n13562 DVSS.n13561 0.4505
R43130 DVSS.n21277 DVSS.n21276 0.4505
R43131 DVSS.n21279 DVSS.n21278 0.4505
R43132 DVSS.n21281 DVSS.n21280 0.4505
R43133 DVSS.n13559 DVSS.n13558 0.4505
R43134 DVSS.n21286 DVSS.n21285 0.4505
R43135 DVSS.n21288 DVSS.n21287 0.4505
R43136 DVSS.n21290 DVSS.n21289 0.4505
R43137 DVSS.n13555 DVSS.n13554 0.4505
R43138 DVSS.n21296 DVSS.n21295 0.4505
R43139 DVSS.n13556 DVSS.n13516 0.4505
R43140 DVSS.n21300 DVSS.n13515 0.4505
R43141 DVSS.n21302 DVSS.n21301 0.4505
R43142 DVSS.n13513 DVSS.n13512 0.4505
R43143 DVSS.n21308 DVSS.n21307 0.4505
R43144 DVSS.n21309 DVSS.n13511 0.4505
R43145 DVSS.n21311 DVSS.n21310 0.4505
R43146 DVSS.n21313 DVSS.n21312 0.4505
R43147 DVSS.n13509 DVSS.n13508 0.4505
R43148 DVSS.n21318 DVSS.n21317 0.4505
R43149 DVSS.n21320 DVSS.n21319 0.4505
R43150 DVSS.n21322 DVSS.n21321 0.4505
R43151 DVSS.n13506 DVSS.n13505 0.4505
R43152 DVSS.n21327 DVSS.n21326 0.4505
R43153 DVSS.n21329 DVSS.n21328 0.4505
R43154 DVSS.n21331 DVSS.n21330 0.4505
R43155 DVSS.n13503 DVSS.n13502 0.4505
R43156 DVSS.n21336 DVSS.n21335 0.4505
R43157 DVSS.n21337 DVSS.n13464 0.4505
R43158 DVSS.n21342 DVSS.n21341 0.4505
R43159 DVSS.n13462 DVSS.n13461 0.4505
R43160 DVSS.n21348 DVSS.n21347 0.4505
R43161 DVSS.n21349 DVSS.n13460 0.4505
R43162 DVSS.n21351 DVSS.n21350 0.4505
R43163 DVSS.n21353 DVSS.n21352 0.4505
R43164 DVSS.n13458 DVSS.n13457 0.4505
R43165 DVSS.n455 DVSS.n454 0.4505
R43166 DVSS.n22881 DVSS.n22880 0.4505
R43167 DVSS.n22875 DVSS.n457 0.4505
R43168 DVSS.n22873 DVSS.n22872 0.4505
R43169 DVSS.n22869 DVSS.n483 0.4505
R43170 DVSS.n22868 DVSS.n22867 0.4505
R43171 DVSS.n22866 DVSS.n22865 0.4505
R43172 DVSS.n486 DVSS.n485 0.4505
R43173 DVSS.n22861 DVSS.n22860 0.4505
R43174 DVSS.n22859 DVSS.n22858 0.4505
R43175 DVSS.n22857 DVSS.n22856 0.4505
R43176 DVSS.n489 DVSS.n488 0.4505
R43177 DVSS.n22852 DVSS.n22851 0.4505
R43178 DVSS.n22850 DVSS.n22849 0.4505
R43179 DVSS.n22848 DVSS.n491 0.4505
R43180 DVSS.n22847 DVSS.n22846 0.4505
R43181 DVSS.n493 DVSS.n492 0.4505
R43182 DVSS.n22841 DVSS.n22840 0.4505
R43183 DVSS.n496 DVSS.n495 0.4505
R43184 DVSS.n22836 DVSS.n22835 0.4505
R43185 DVSS.n730 DVSS.n729 0.4505
R43186 DVSS.n22670 DVSS.n22669 0.4505
R43187 DVSS.n732 DVSS.n731 0.4505
R43188 DVSS.n22665 DVSS.n22664 0.4505
R43189 DVSS.n22663 DVSS.n22662 0.4505
R43190 DVSS.n22661 DVSS.n22660 0.4505
R43191 DVSS.n22642 DVSS.n22641 0.4505
R43192 DVSS.n22656 DVSS.n22655 0.4505
R43193 DVSS.n22654 DVSS.n22653 0.4505
R43194 DVSS.n22652 DVSS.n22651 0.4505
R43195 DVSS.n22645 DVSS.n22644 0.4505
R43196 DVSS.n22647 DVSS.n22646 0.4505
R43197 DVSS.n701 DVSS.n700 0.4505
R43198 DVSS.n22675 DVSS.n22674 0.4505
R43199 DVSS.n698 DVSS.n697 0.4505
R43200 DVSS.n22681 DVSS.n22680 0.4505
R43201 DVSS.n22682 DVSS.n696 0.4505
R43202 DVSS.n22684 DVSS.n22683 0.4505
R43203 DVSS.n22686 DVSS.n22685 0.4505
R43204 DVSS.n694 DVSS.n693 0.4505
R43205 DVSS.n22691 DVSS.n22690 0.4505
R43206 DVSS.n22693 DVSS.n22692 0.4505
R43207 DVSS.n22695 DVSS.n22694 0.4505
R43208 DVSS.n691 DVSS.n690 0.4505
R43209 DVSS.n22700 DVSS.n22699 0.4505
R43210 DVSS.n22702 DVSS.n22701 0.4505
R43211 DVSS.n22704 DVSS.n22703 0.4505
R43212 DVSS.n688 DVSS.n687 0.4505
R43213 DVSS.n22709 DVSS.n22708 0.4505
R43214 DVSS.n22711 DVSS.n647 0.4505
R43215 DVSS.n22717 DVSS.n22716 0.4505
R43216 DVSS.n645 DVSS.n644 0.4505
R43217 DVSS.n22723 DVSS.n22722 0.4505
R43218 DVSS.n22724 DVSS.n642 0.4505
R43219 DVSS.n22726 DVSS.n22725 0.4505
R43220 DVSS.n22728 DVSS.n22727 0.4505
R43221 DVSS.n22730 DVSS.n22729 0.4505
R43222 DVSS.n640 DVSS.n639 0.4505
R43223 DVSS.n22735 DVSS.n22734 0.4505
R43224 DVSS.n22737 DVSS.n22736 0.4505
R43225 DVSS.n22739 DVSS.n22738 0.4505
R43226 DVSS.n637 DVSS.n636 0.4505
R43227 DVSS.n22744 DVSS.n22743 0.4505
R43228 DVSS.n22746 DVSS.n22745 0.4505
R43229 DVSS.n22748 DVSS.n22747 0.4505
R43230 DVSS.n633 DVSS.n632 0.4505
R43231 DVSS.n22754 DVSS.n22753 0.4505
R43232 DVSS.n634 DVSS.n596 0.4505
R43233 DVSS.n22758 DVSS.n595 0.4505
R43234 DVSS.n22760 DVSS.n22759 0.4505
R43235 DVSS.n593 DVSS.n592 0.4505
R43236 DVSS.n22766 DVSS.n22765 0.4505
R43237 DVSS.n22767 DVSS.n591 0.4505
R43238 DVSS.n22769 DVSS.n22768 0.4505
R43239 DVSS.n22771 DVSS.n22770 0.4505
R43240 DVSS.n589 DVSS.n588 0.4505
R43241 DVSS.n22776 DVSS.n22775 0.4505
R43242 DVSS.n22778 DVSS.n22777 0.4505
R43243 DVSS.n22780 DVSS.n22779 0.4505
R43244 DVSS.n586 DVSS.n585 0.4505
R43245 DVSS.n22785 DVSS.n22784 0.4505
R43246 DVSS.n22787 DVSS.n22786 0.4505
R43247 DVSS.n22789 DVSS.n22788 0.4505
R43248 DVSS.n583 DVSS.n582 0.4505
R43249 DVSS.n22794 DVSS.n22793 0.4505
R43250 DVSS.n22795 DVSS.n546 0.4505
R43251 DVSS.n22800 DVSS.n22799 0.4505
R43252 DVSS.n544 DVSS.n543 0.4505
R43253 DVSS.n22806 DVSS.n22805 0.4505
R43254 DVSS.n22807 DVSS.n541 0.4505
R43255 DVSS.n22809 DVSS.n22808 0.4505
R43256 DVSS.n22811 DVSS.n22810 0.4505
R43257 DVSS.n22813 DVSS.n22812 0.4505
R43258 DVSS.n539 DVSS.n538 0.4505
R43259 DVSS.n22818 DVSS.n22817 0.4505
R43260 DVSS.n22820 DVSS.n22819 0.4505
R43261 DVSS.n22822 DVSS.n22821 0.4505
R43262 DVSS.n536 DVSS.n535 0.4505
R43263 DVSS.n22827 DVSS.n22826 0.4505
R43264 DVSS.n22829 DVSS.n22828 0.4505
R43265 DVSS.n22831 DVSS.n22830 0.4505
R43266 DVSS.n533 DVSS.n532 0.4505
R43267 DVSS.n19203 DVSS.n13481 0.417781
R43268 DVSS.n19904 DVSS.n19002 0.416947
R43269 DVSS.n19200 DVSS.n19181 0.416947
R43270 DVSS.n22230 DVSS.n1352 0.404033
R43271 DVSS.n22233 DVSS.n1271 0.404033
R43272 DVSS.n22457 DVSS.n22456 0.404033
R43273 DVSS.n22335 DVSS.n22334 0.404033
R43274 DVSS.n19513 DVSS.n19501 0.404033
R43275 DVSS.n19846 DVSS.n19845 0.404033
R43276 DVSS.n19214 DVSS.n19213 0.400763
R43277 DVSS.n19202 DVSS.n19200 0.371929
R43278 DVSS.n19202 DVSS.n19201 0.371929
R43279 DVSS.n19905 DVSS.n19904 0.371929
R43280 DVSS.n19906 DVSS.n19905 0.371929
R43281 DVSS.n15541 DVSS 0.367475
R43282 DVSS.n18174 DVSS.n18173 0.355011
R43283 DVSS.n18248 DVSS.n15140 0.355011
R43284 DVSS.n20984 DVSS.n20983 0.355011
R43285 DVSS.n21438 DVSS.n21437 0.355011
R43286 DVSS.n22885 DVSS.n22884 0.355011
R43287 DVSS.n17785 DVSS.n17784 0.354754
R43288 DVSS.n17719 DVSS.n15146 0.354754
R43289 DVSS.n21153 DVSS.n21152 0.354754
R43290 DVSS.n21180 DVSS.n21179 0.354754
R43291 DVSS.n22638 DVSS.n22637 0.354754
R43292 DVSS.n19191 DVSS.n19186 0.343668
R43293 DVSS.n13681 DVSS.n13680 0.335693
R43294 DVSS.n19210 DVSS.t196 0.3281
R43295 DVSS.n19210 DVSS.t186 0.3281
R43296 DVSS.n19173 DVSS.t179 0.3281
R43297 DVSS.n19173 DVSS.t198 0.3281
R43298 DVSS.n19187 DVSS.t163 0.3281
R43299 DVSS.n19187 DVSS.t181 0.3281
R43300 DVSS.n19190 DVSS.t183 0.3281
R43301 DVSS.n19190 DVSS.t177 0.3281
R43302 DVSS.n19184 DVSS.t165 0.3281
R43303 DVSS.n19184 DVSS.t171 0.3281
R43304 DVSS.n19903 DVSS.n19902 0.321929
R43305 DVSS.n19199 DVSS.n19147 0.321929
R43306 DVSS.n21146 DVSS.n13702 0.320711
R43307 DVSS.n19953 DVSS.n14326 0.320711
R43308 DVSS.n15540 DVSS.t191 0.312926
R43309 DVSS.n15540 DVSS.t193 0.312926
R43310 DVSS.n15584 DVSS.t192 0.312926
R43311 DVSS.n16488 DVSS.t194 0.312926
R43312 DVSS.n16403 DVSS.t193 0.312926
R43313 DVSS.n16403 DVSS.t194 0.312926
R43314 DVSS.n15684 DVSS.t192 0.312926
R43315 DVSS.n15684 DVSS.t191 0.312926
R43316 DVSS.n21154 DVSS.n21153 0.292137
R43317 DVSS.n13682 DVSS.n13681 0.285184
R43318 DVSS.n16195 DVSS.n15645 0.264133
R43319 DVSS.n16464 DVSS.n16462 0.264133
R43320 DVSS.n21171 DVSS.n21170 0.258595
R43321 DVSS.n17798 DVSS.n15916 0.256847
R43322 DVSS.n18001 DVSS.n18000 0.256847
R43323 DVSS.n17786 DVSS.n15144 0.252283
R43324 DVSS.n18172 DVSS.n15141 0.252283
R43325 DVSS.n18507 DVSS.n13686 0.247099
R43326 DVSS.n21214 DVSS.n13629 0.244637
R43327 DVSS.n14251 DVSS.n13383 0.244637
R43328 DVSS.n22628 DVSS.n22627 0.243721
R43329 DVSS.n22894 DVSS.n22893 0.243721
R43330 DVSS.n19196 DVSS.n19160 0.237342
R43331 DVSS.n22668 DVSS.n22639 0.231338
R43332 DVSS.n22883 DVSS.n22882 0.231338
R43333 DVSS.n16572 DVSS.n16567 0.231338
R43334 DVSS.n16740 DVSS.n16739 0.231338
R43335 DVSS.n17783 DVSS.n17782 0.231338
R43336 DVSS.n18178 DVSS.n18177 0.231338
R43337 DVSS.n17723 DVSS.n17722 0.231338
R43338 DVSS.n18252 DVSS.n18251 0.231338
R43339 DVSS.n18496 DVSS.n18495 0.231338
R43340 DVSS.n19931 DVSS.n19930 0.231338
R43341 DVSS.n21151 DVSS.n21150 0.231338
R43342 DVSS.n20982 DVSS.n20981 0.231338
R43343 DVSS.n21185 DVSS.n13658 0.231338
R43344 DVSS.n21436 DVSS.n21435 0.231338
R43345 DVSS.n22973 DVSS.n22972 0.229958
R43346 DVSS.n13663 DVSS.n13662 0.221772
R43347 DVSS.n19314 DVSS.n19012 0.220853
R43348 DVSS.n19653 DVSS.n19652 0.220853
R43349 DVSS.n22432 DVSS.n22386 0.220853
R43350 DVSS.n1409 DVSS.n1408 0.218146
R43351 DVSS.n22570 DVSS.n22569 0.218146
R43352 DVSS.n21475 DVSS.n21474 0.218146
R43353 DVSS.n13788 DVSS.n13787 0.217409
R43354 DVSS.n21026 DVSS.n14308 0.217409
R43355 DVSS.n21991 DVSS.n21988 0.217409
R43356 DVSS.n23224 DVSS.n3 0.217409
R43357 DVSS.n14228 DVSS.n14227 0.214786
R43358 DVSS.n21030 DVSS.n14307 0.214786
R43359 DVSS.n21032 DVSS.n14306 0.214786
R43360 DVSS.n21034 DVSS.n14305 0.214786
R43361 DVSS.n21036 DVSS.n14304 0.214786
R43362 DVSS.n21038 DVSS.n14303 0.214786
R43363 DVSS.n21040 DVSS.n14302 0.214786
R43364 DVSS.n21042 DVSS.n14301 0.214786
R43365 DVSS.n21044 DVSS.n14300 0.214786
R43366 DVSS.n21045 DVSS.n14299 0.214786
R43367 DVSS.n14298 DVSS.n14296 0.214786
R43368 DVSS.n14297 DVSS.n14238 0.214786
R43369 DVSS.n21056 DVSS.n14237 0.214786
R43370 DVSS.n21057 DVSS.n14236 0.214786
R43371 DVSS.n14235 DVSS.n14233 0.214786
R43372 DVSS.n21061 DVSS.n14232 0.214786
R43373 DVSS.n21062 DVSS.n14231 0.214786
R43374 DVSS.n21063 DVSS.n14230 0.214786
R43375 DVSS.n14229 DVSS.n14192 0.214786
R43376 DVSS.n13793 DVSS.n13792 0.214786
R43377 DVSS.n13794 DVSS.n13786 0.214786
R43378 DVSS.n13797 DVSS.n13795 0.214786
R43379 DVSS.n13799 DVSS.n13784 0.214786
R43380 DVSS.n13802 DVSS.n13801 0.214786
R43381 DVSS.n13803 DVSS.n13783 0.214786
R43382 DVSS.n13806 DVSS.n13804 0.214786
R43383 DVSS.n13808 DVSS.n13781 0.214786
R43384 DVSS.n13811 DVSS.n13810 0.214786
R43385 DVSS.n13812 DVSS.n13780 0.214786
R43386 DVSS.n21127 DVSS.n13813 0.214786
R43387 DVSS.n21126 DVSS.n13814 0.214786
R43388 DVSS.n21125 DVSS.n13815 0.214786
R43389 DVSS.n21124 DVSS.n13816 0.214786
R43390 DVSS.n13819 DVSS.n13817 0.214786
R43391 DVSS.n21120 DVSS.n13820 0.214786
R43392 DVSS.n21119 DVSS.n13821 0.214786
R43393 DVSS.n21118 DVSS.n13822 0.214786
R43394 DVSS.n13897 DVSS.n13823 0.214786
R43395 DVSS.n13900 DVSS.n13898 0.214786
R43396 DVSS.n13903 DVSS.n13902 0.214786
R43397 DVSS.n13904 DVSS.n13896 0.214786
R43398 DVSS.n13907 DVSS.n13905 0.214786
R43399 DVSS.n13909 DVSS.n13894 0.214786
R43400 DVSS.n13912 DVSS.n13911 0.214786
R43401 DVSS.n13913 DVSS.n13893 0.214786
R43402 DVSS.n13916 DVSS.n13914 0.214786
R43403 DVSS.n13918 DVSS.n13891 0.214786
R43404 DVSS.n13921 DVSS.n13920 0.214786
R43405 DVSS.n13922 DVSS.n13890 0.214786
R43406 DVSS.n21112 DVSS.n13923 0.214786
R43407 DVSS.n21111 DVSS.n13924 0.214786
R43408 DVSS.n21110 DVSS.n13925 0.214786
R43409 DVSS.n13987 DVSS.n13926 0.214786
R43410 DVSS.n13988 DVSS.n13986 0.214786
R43411 DVSS.n13991 DVSS.n13989 0.214786
R43412 DVSS.n13993 DVSS.n13985 0.214786
R43413 DVSS.n13996 DVSS.n13995 0.214786
R43414 DVSS.n13997 DVSS.n13984 0.214786
R43415 DVSS.n14000 DVSS.n13998 0.214786
R43416 DVSS.n14002 DVSS.n13982 0.214786
R43417 DVSS.n14005 DVSS.n14004 0.214786
R43418 DVSS.n14006 DVSS.n13981 0.214786
R43419 DVSS.n21101 DVSS.n14007 0.214786
R43420 DVSS.n21100 DVSS.n14008 0.214786
R43421 DVSS.n21098 DVSS.n14009 0.214786
R43422 DVSS.n21086 DVSS.n14010 0.214786
R43423 DVSS.n21085 DVSS.n14011 0.214786
R43424 DVSS.n21084 DVSS.n14012 0.214786
R43425 DVSS.n14015 DVSS.n14013 0.214786
R43426 DVSS.n21080 DVSS.n14016 0.214786
R43427 DVSS.n21079 DVSS.n14017 0.214786
R43428 DVSS.n21078 DVSS.n14018 0.214786
R43429 DVSS.n14094 DVSS.n14019 0.214786
R43430 DVSS.n14097 DVSS.n14095 0.214786
R43431 DVSS.n14099 DVSS.n14093 0.214786
R43432 DVSS.n14102 DVSS.n14101 0.214786
R43433 DVSS.n14103 DVSS.n14092 0.214786
R43434 DVSS.n14106 DVSS.n14104 0.214786
R43435 DVSS.n14108 DVSS.n14090 0.214786
R43436 DVSS.n14111 DVSS.n14110 0.214786
R43437 DVSS.n14112 DVSS.n14089 0.214786
R43438 DVSS.n14115 DVSS.n14113 0.214786
R43439 DVSS.n14117 DVSS.n14087 0.214786
R43440 DVSS.n14120 DVSS.n14119 0.214786
R43441 DVSS.n14121 DVSS.n14086 0.214786
R43442 DVSS.n21072 DVSS.n14122 0.214786
R43443 DVSS.n21071 DVSS.n14123 0.214786
R43444 DVSS.n21070 DVSS.n14124 0.214786
R43445 DVSS.n14201 DVSS.n14125 0.214786
R43446 DVSS.n14202 DVSS.n14200 0.214786
R43447 DVSS.n14205 DVSS.n14203 0.214786
R43448 DVSS.n14207 DVSS.n14199 0.214786
R43449 DVSS.n14210 DVSS.n14209 0.214786
R43450 DVSS.n14211 DVSS.n14198 0.214786
R43451 DVSS.n14214 DVSS.n14212 0.214786
R43452 DVSS.n14216 DVSS.n14196 0.214786
R43453 DVSS.n14219 DVSS.n14218 0.214786
R43454 DVSS.n14220 DVSS.n14195 0.214786
R43455 DVSS.n14223 DVSS.n14221 0.214786
R43456 DVSS.n14225 DVSS.n14193 0.214786
R43457 DVSS.n21028 DVSS.n21027 0.214786
R43458 DVSS.n21030 DVSS.n21029 0.214786
R43459 DVSS.n21032 DVSS.n21031 0.214786
R43460 DVSS.n21034 DVSS.n21033 0.214786
R43461 DVSS.n21036 DVSS.n21035 0.214786
R43462 DVSS.n21038 DVSS.n21037 0.214786
R43463 DVSS.n21040 DVSS.n21039 0.214786
R43464 DVSS.n21042 DVSS.n21041 0.214786
R43465 DVSS.n21044 DVSS.n21043 0.214786
R43466 DVSS.n21046 DVSS.n21045 0.214786
R43467 DVSS.n14296 DVSS.n14277 0.214786
R43468 DVSS.n14239 DVSS.n14238 0.214786
R43469 DVSS.n21056 DVSS.n21055 0.214786
R43470 DVSS.n21058 DVSS.n21057 0.214786
R43471 DVSS.n21059 DVSS.n14233 0.214786
R43472 DVSS.n21061 DVSS.n21060 0.214786
R43473 DVSS.n21062 DVSS.n14191 0.214786
R43474 DVSS.n21064 DVSS.n21063 0.214786
R43475 DVSS.n14192 DVSS.n14190 0.214786
R43476 DVSS.n14227 DVSS.n14226 0.214786
R43477 DVSS.n13790 DVSS.n13789 0.214786
R43478 DVSS.n13792 DVSS.n13791 0.214786
R43479 DVSS.n13786 DVSS.n13785 0.214786
R43480 DVSS.n13797 DVSS.n13796 0.214786
R43481 DVSS.n13799 DVSS.n13798 0.214786
R43482 DVSS.n13801 DVSS.n13800 0.214786
R43483 DVSS.n13783 DVSS.n13782 0.214786
R43484 DVSS.n13806 DVSS.n13805 0.214786
R43485 DVSS.n13808 DVSS.n13807 0.214786
R43486 DVSS.n13810 DVSS.n13809 0.214786
R43487 DVSS.n13780 DVSS.n13779 0.214786
R43488 DVSS.n21128 DVSS.n21127 0.214786
R43489 DVSS.n21126 DVSS.n13745 0.214786
R43490 DVSS.n21125 DVSS.n13757 0.214786
R43491 DVSS.n21124 DVSS.n21123 0.214786
R43492 DVSS.n21122 DVSS.n13817 0.214786
R43493 DVSS.n21121 DVSS.n21120 0.214786
R43494 DVSS.n21119 DVSS.n13818 0.214786
R43495 DVSS.n21118 DVSS.n21117 0.214786
R43496 DVSS.n13837 DVSS.n13823 0.214786
R43497 DVSS.n13900 DVSS.n13899 0.214786
R43498 DVSS.n13902 DVSS.n13901 0.214786
R43499 DVSS.n13896 DVSS.n13895 0.214786
R43500 DVSS.n13907 DVSS.n13906 0.214786
R43501 DVSS.n13909 DVSS.n13908 0.214786
R43502 DVSS.n13911 DVSS.n13910 0.214786
R43503 DVSS.n13893 DVSS.n13892 0.214786
R43504 DVSS.n13916 DVSS.n13915 0.214786
R43505 DVSS.n13918 DVSS.n13917 0.214786
R43506 DVSS.n13920 DVSS.n13919 0.214786
R43507 DVSS.n13890 DVSS.n13888 0.214786
R43508 DVSS.n21113 DVSS.n21112 0.214786
R43509 DVSS.n21111 DVSS.n13889 0.214786
R43510 DVSS.n21110 DVSS.n21109 0.214786
R43511 DVSS.n21108 DVSS.n13926 0.214786
R43512 DVSS.n13986 DVSS.n13939 0.214786
R43513 DVSS.n13991 DVSS.n13990 0.214786
R43514 DVSS.n13993 DVSS.n13992 0.214786
R43515 DVSS.n13995 DVSS.n13994 0.214786
R43516 DVSS.n13984 DVSS.n13983 0.214786
R43517 DVSS.n14000 DVSS.n13999 0.214786
R43518 DVSS.n14002 DVSS.n14001 0.214786
R43519 DVSS.n14004 DVSS.n14003 0.214786
R43520 DVSS.n13981 DVSS.n13980 0.214786
R43521 DVSS.n21102 DVSS.n21101 0.214786
R43522 DVSS.n21100 DVSS.n21099 0.214786
R43523 DVSS.n21098 DVSS.n21097 0.214786
R43524 DVSS.n21086 DVSS.n13953 0.214786
R43525 DVSS.n21085 DVSS.n13965 0.214786
R43526 DVSS.n21084 DVSS.n21083 0.214786
R43527 DVSS.n21082 DVSS.n14013 0.214786
R43528 DVSS.n21081 DVSS.n21080 0.214786
R43529 DVSS.n21079 DVSS.n14014 0.214786
R43530 DVSS.n21078 DVSS.n21077 0.214786
R43531 DVSS.n14032 DVSS.n14019 0.214786
R43532 DVSS.n14097 DVSS.n14096 0.214786
R43533 DVSS.n14099 DVSS.n14098 0.214786
R43534 DVSS.n14101 DVSS.n14100 0.214786
R43535 DVSS.n14092 DVSS.n14091 0.214786
R43536 DVSS.n14106 DVSS.n14105 0.214786
R43537 DVSS.n14108 DVSS.n14107 0.214786
R43538 DVSS.n14110 DVSS.n14109 0.214786
R43539 DVSS.n14089 DVSS.n14088 0.214786
R43540 DVSS.n14115 DVSS.n14114 0.214786
R43541 DVSS.n14117 DVSS.n14116 0.214786
R43542 DVSS.n14119 DVSS.n14118 0.214786
R43543 DVSS.n14086 DVSS.n14084 0.214786
R43544 DVSS.n21073 DVSS.n21072 0.214786
R43545 DVSS.n21071 DVSS.n14085 0.214786
R43546 DVSS.n21070 DVSS.n21069 0.214786
R43547 DVSS.n21068 DVSS.n14125 0.214786
R43548 DVSS.n14200 DVSS.n14138 0.214786
R43549 DVSS.n14205 DVSS.n14204 0.214786
R43550 DVSS.n14207 DVSS.n14206 0.214786
R43551 DVSS.n14209 DVSS.n14208 0.214786
R43552 DVSS.n14198 DVSS.n14197 0.214786
R43553 DVSS.n14214 DVSS.n14213 0.214786
R43554 DVSS.n14216 DVSS.n14215 0.214786
R43555 DVSS.n14218 DVSS.n14217 0.214786
R43556 DVSS.n14195 DVSS.n14194 0.214786
R43557 DVSS.n14223 DVSS.n14222 0.214786
R43558 DVSS.n14225 DVSS.n14224 0.214786
R43559 DVSS.n1407 DVSS.n1405 0.214786
R43560 DVSS.n21990 DVSS.n21989 0.214786
R43561 DVSS.n21987 DVSS.n21986 0.214786
R43562 DVSS.n21994 DVSS.n21985 0.214786
R43563 DVSS.n21995 DVSS.n21984 0.214786
R43564 DVSS.n21996 DVSS.n21983 0.214786
R43565 DVSS.n21981 DVSS.n21980 0.214786
R43566 DVSS.n22000 DVSS.n21979 0.214786
R43567 DVSS.n22001 DVSS.n21978 0.214786
R43568 DVSS.n22002 DVSS.n21977 0.214786
R43569 DVSS.n21975 DVSS.n21974 0.214786
R43570 DVSS.n22006 DVSS.n21973 0.214786
R43571 DVSS.n22007 DVSS.n21972 0.214786
R43572 DVSS.n22008 DVSS.n1252 0.214786
R43573 DVSS.n21969 DVSS.n1238 0.214786
R43574 DVSS.n22012 DVSS.n21968 0.214786
R43575 DVSS.n22014 DVSS.n21967 0.214786
R43576 DVSS.n22015 DVSS.n21966 0.214786
R43577 DVSS.n21965 DVSS.n21775 0.214786
R43578 DVSS.n22019 DVSS.n21774 0.214786
R43579 DVSS.n22020 DVSS.n21773 0.214786
R43580 DVSS.n22021 DVSS.n21772 0.214786
R43581 DVSS.n21960 DVSS.n21770 0.214786
R43582 DVSS.n22025 DVSS.n21769 0.214786
R43583 DVSS.n22026 DVSS.n21768 0.214786
R43584 DVSS.n22027 DVSS.n21767 0.214786
R43585 DVSS.n21956 DVSS.n21765 0.214786
R43586 DVSS.n22031 DVSS.n21764 0.214786
R43587 DVSS.n22032 DVSS.n21763 0.214786
R43588 DVSS.n22033 DVSS.n21762 0.214786
R43589 DVSS.n21953 DVSS.n21760 0.214786
R43590 DVSS.n22037 DVSS.n21759 0.214786
R43591 DVSS.n22038 DVSS.n21758 0.214786
R43592 DVSS.n22039 DVSS.n21757 0.214786
R43593 DVSS.n21746 DVSS.n21744 0.214786
R43594 DVSS.n22044 DVSS.n22043 0.214786
R43595 DVSS.n21745 DVSS.n21743 0.214786
R43596 DVSS.n21753 DVSS.n21752 0.214786
R43597 DVSS.n21751 DVSS.n21750 0.214786
R43598 DVSS.n21749 DVSS.n21694 0.214786
R43599 DVSS.n22049 DVSS.n22048 0.214786
R43600 DVSS.n21726 DVSS.n21680 0.214786
R43601 DVSS.n22053 DVSS.n21679 0.214786
R43602 DVSS.n22054 DVSS.n21678 0.214786
R43603 DVSS.n22055 DVSS.n21677 0.214786
R43604 DVSS.n21737 DVSS.n21675 0.214786
R43605 DVSS.n22059 DVSS.n21674 0.214786
R43606 DVSS.n22060 DVSS.n21673 0.214786
R43607 DVSS.n22061 DVSS.n21672 0.214786
R43608 DVSS.n21731 DVSS.n21670 0.214786
R43609 DVSS.n22065 DVSS.n21669 0.214786
R43610 DVSS.n22066 DVSS.n21668 0.214786
R43611 DVSS.n22067 DVSS.n21667 0.214786
R43612 DVSS.n21641 DVSS.n21639 0.214786
R43613 DVSS.n22072 DVSS.n22071 0.214786
R43614 DVSS.n21640 DVSS.n21638 0.214786
R43615 DVSS.n21663 DVSS.n21662 0.214786
R43616 DVSS.n21661 DVSS.n21660 0.214786
R43617 DVSS.n21659 DVSS.n21645 0.214786
R43618 DVSS.n21644 DVSS.n21643 0.214786
R43619 DVSS.n21655 DVSS.n21654 0.214786
R43620 DVSS.n21653 DVSS.n21652 0.214786
R43621 DVSS.n21651 DVSS.n21648 0.214786
R43622 DVSS.n21647 DVSS.n21591 0.214786
R43623 DVSS.n22078 DVSS.n22077 0.214786
R43624 DVSS.n22081 DVSS.n1462 0.214786
R43625 DVSS.n22082 DVSS.n1461 0.214786
R43626 DVSS.n22083 DVSS.n1460 0.214786
R43627 DVSS.n21627 DVSS.n1458 0.214786
R43628 DVSS.n22087 DVSS.n1457 0.214786
R43629 DVSS.n22088 DVSS.n1456 0.214786
R43630 DVSS.n22089 DVSS.n1455 0.214786
R43631 DVSS.n21870 DVSS.n1453 0.214786
R43632 DVSS.n22093 DVSS.n1452 0.214786
R43633 DVSS.n22094 DVSS.n1451 0.214786
R43634 DVSS.n22095 DVSS.n1450 0.214786
R43635 DVSS.n21866 DVSS.n1448 0.214786
R43636 DVSS.n22099 DVSS.n1447 0.214786
R43637 DVSS.n22100 DVSS.n1446 0.214786
R43638 DVSS.n22101 DVSS.n1445 0.214786
R43639 DVSS.n21862 DVSS.n1443 0.214786
R43640 DVSS.n22105 DVSS.n1442 0.214786
R43641 DVSS.n22106 DVSS.n1441 0.214786
R43642 DVSS.n22107 DVSS.n1440 0.214786
R43643 DVSS.n21859 DVSS.n1438 0.214786
R43644 DVSS.n22111 DVSS.n1437 0.214786
R43645 DVSS.n22112 DVSS.n1436 0.214786
R43646 DVSS.n22113 DVSS.n1435 0.214786
R43647 DVSS.n1395 DVSS.n1393 0.214786
R43648 DVSS.n22119 DVSS.n22118 0.214786
R43649 DVSS.n1394 DVSS.n1378 0.214786
R43650 DVSS.n1431 DVSS.n1430 0.214786
R43651 DVSS.n1429 DVSS.n1428 0.214786
R43652 DVSS.n1427 DVSS.n1399 0.214786
R43653 DVSS.n1398 DVSS.n1397 0.214786
R43654 DVSS.n1423 DVSS.n1422 0.214786
R43655 DVSS.n1421 DVSS.n1420 0.214786
R43656 DVSS.n1419 DVSS.n1403 0.214786
R43657 DVSS.n1402 DVSS.n1401 0.214786
R43658 DVSS.n1415 DVSS.n1414 0.214786
R43659 DVSS.n1413 DVSS.n1412 0.214786
R43660 DVSS.n1411 DVSS.n1406 0.214786
R43661 DVSS.n1411 DVSS.n1410 0.214786
R43662 DVSS.n1413 DVSS.n1404 0.214786
R43663 DVSS.n1416 DVSS.n1415 0.214786
R43664 DVSS.n1417 DVSS.n1402 0.214786
R43665 DVSS.n1419 DVSS.n1418 0.214786
R43666 DVSS.n1421 DVSS.n1400 0.214786
R43667 DVSS.n1424 DVSS.n1423 0.214786
R43668 DVSS.n1425 DVSS.n1398 0.214786
R43669 DVSS.n1427 DVSS.n1426 0.214786
R43670 DVSS.n1429 DVSS.n1396 0.214786
R43671 DVSS.n1432 DVSS.n1431 0.214786
R43672 DVSS.n1433 DVSS.n1394 0.214786
R43673 DVSS.n22118 DVSS.n22117 0.214786
R43674 DVSS.n22116 DVSS.n1395 0.214786
R43675 DVSS.n22114 DVSS.n22113 0.214786
R43676 DVSS.n22112 DVSS.n1434 0.214786
R43677 DVSS.n22111 DVSS.n22110 0.214786
R43678 DVSS.n22109 DVSS.n1438 0.214786
R43679 DVSS.n22108 DVSS.n22107 0.214786
R43680 DVSS.n22106 DVSS.n1439 0.214786
R43681 DVSS.n22105 DVSS.n22104 0.214786
R43682 DVSS.n22103 DVSS.n1443 0.214786
R43683 DVSS.n22102 DVSS.n22101 0.214786
R43684 DVSS.n22100 DVSS.n1444 0.214786
R43685 DVSS.n22099 DVSS.n22098 0.214786
R43686 DVSS.n22097 DVSS.n1448 0.214786
R43687 DVSS.n22096 DVSS.n22095 0.214786
R43688 DVSS.n22094 DVSS.n1449 0.214786
R43689 DVSS.n22093 DVSS.n22092 0.214786
R43690 DVSS.n22091 DVSS.n1453 0.214786
R43691 DVSS.n22090 DVSS.n22089 0.214786
R43692 DVSS.n22088 DVSS.n1454 0.214786
R43693 DVSS.n22087 DVSS.n22086 0.214786
R43694 DVSS.n22085 DVSS.n1458 0.214786
R43695 DVSS.n22084 DVSS.n22083 0.214786
R43696 DVSS.n22082 DVSS.n1459 0.214786
R43697 DVSS.n22081 DVSS.n22080 0.214786
R43698 DVSS.n22079 DVSS.n22078 0.214786
R43699 DVSS.n21649 DVSS.n21647 0.214786
R43700 DVSS.n21651 DVSS.n21650 0.214786
R43701 DVSS.n21653 DVSS.n21646 0.214786
R43702 DVSS.n21656 DVSS.n21655 0.214786
R43703 DVSS.n21657 DVSS.n21644 0.214786
R43704 DVSS.n21659 DVSS.n21658 0.214786
R43705 DVSS.n21661 DVSS.n21642 0.214786
R43706 DVSS.n21664 DVSS.n21663 0.214786
R43707 DVSS.n21665 DVSS.n21640 0.214786
R43708 DVSS.n22071 DVSS.n22070 0.214786
R43709 DVSS.n22069 DVSS.n21641 0.214786
R43710 DVSS.n22068 DVSS.n22067 0.214786
R43711 DVSS.n22066 DVSS.n21666 0.214786
R43712 DVSS.n22065 DVSS.n22064 0.214786
R43713 DVSS.n22063 DVSS.n21670 0.214786
R43714 DVSS.n22062 DVSS.n22061 0.214786
R43715 DVSS.n22060 DVSS.n21671 0.214786
R43716 DVSS.n22059 DVSS.n22058 0.214786
R43717 DVSS.n22057 DVSS.n21675 0.214786
R43718 DVSS.n22056 DVSS.n22055 0.214786
R43719 DVSS.n22054 DVSS.n21676 0.214786
R43720 DVSS.n22053 DVSS.n22052 0.214786
R43721 DVSS.n22051 DVSS.n21680 0.214786
R43722 DVSS.n22050 DVSS.n22049 0.214786
R43723 DVSS.n21749 DVSS.n21748 0.214786
R43724 DVSS.n21751 DVSS.n21747 0.214786
R43725 DVSS.n21754 DVSS.n21753 0.214786
R43726 DVSS.n21755 DVSS.n21745 0.214786
R43727 DVSS.n22043 DVSS.n22042 0.214786
R43728 DVSS.n22041 DVSS.n21746 0.214786
R43729 DVSS.n22040 DVSS.n22039 0.214786
R43730 DVSS.n22038 DVSS.n21756 0.214786
R43731 DVSS.n22037 DVSS.n22036 0.214786
R43732 DVSS.n22035 DVSS.n21760 0.214786
R43733 DVSS.n22034 DVSS.n22033 0.214786
R43734 DVSS.n22032 DVSS.n21761 0.214786
R43735 DVSS.n22031 DVSS.n22030 0.214786
R43736 DVSS.n22029 DVSS.n21765 0.214786
R43737 DVSS.n22028 DVSS.n22027 0.214786
R43738 DVSS.n22026 DVSS.n21766 0.214786
R43739 DVSS.n22025 DVSS.n22024 0.214786
R43740 DVSS.n22023 DVSS.n21770 0.214786
R43741 DVSS.n22022 DVSS.n22021 0.214786
R43742 DVSS.n22020 DVSS.n21771 0.214786
R43743 DVSS.n22019 DVSS.n22018 0.214786
R43744 DVSS.n22017 DVSS.n21775 0.214786
R43745 DVSS.n22016 DVSS.n22015 0.214786
R43746 DVSS.n22014 DVSS.n21776 0.214786
R43747 DVSS.n22012 DVSS.n22011 0.214786
R43748 DVSS.n22010 DVSS.n21969 0.214786
R43749 DVSS.n22009 DVSS.n22008 0.214786
R43750 DVSS.n22007 DVSS.n21971 0.214786
R43751 DVSS.n22006 DVSS.n22005 0.214786
R43752 DVSS.n22004 DVSS.n21975 0.214786
R43753 DVSS.n22003 DVSS.n22002 0.214786
R43754 DVSS.n22001 DVSS.n21976 0.214786
R43755 DVSS.n22000 DVSS.n21999 0.214786
R43756 DVSS.n21998 DVSS.n21981 0.214786
R43757 DVSS.n21997 DVSS.n21996 0.214786
R43758 DVSS.n21995 DVSS.n21982 0.214786
R43759 DVSS.n21994 DVSS.n21993 0.214786
R43760 DVSS.n21992 DVSS.n21987 0.214786
R43761 DVSS.n23223 DVSS.n23222 0.214786
R43762 DVSS.n4 DVSS.n2 0.214786
R43763 DVSS.n23227 DVSS.n1 0.214786
R43764 DVSS.n23216 DVSS.n0 0.214786
R43765 DVSS.n23215 DVSS.n23214 0.214786
R43766 DVSS.n44 DVSS.n43 0.214786
R43767 DVSS.n23209 DVSS.n23208 0.214786
R43768 DVSS.n23207 DVSS.n23206 0.214786
R43769 DVSS.n23205 DVSS.n48 0.214786
R43770 DVSS.n47 DVSS.n46 0.214786
R43771 DVSS.n23201 DVSS.n23200 0.214786
R43772 DVSS.n23199 DVSS.n23198 0.214786
R43773 DVSS.n23197 DVSS.n51 0.214786
R43774 DVSS.n23191 DVSS.n50 0.214786
R43775 DVSS.n23193 DVSS.n23192 0.214786
R43776 DVSS.n23189 DVSS.n23188 0.214786
R43777 DVSS.n57 DVSS.n56 0.214786
R43778 DVSS.n23184 DVSS.n23183 0.214786
R43779 DVSS.n60 DVSS.n59 0.214786
R43780 DVSS.n23179 DVSS.n23178 0.214786
R43781 DVSS.n111 DVSS.n110 0.214786
R43782 DVSS.n23174 DVSS.n23173 0.214786
R43783 DVSS.n23164 DVSS.n23163 0.214786
R43784 DVSS.n23162 DVSS.n115 0.214786
R43785 DVSS.n114 DVSS.n113 0.214786
R43786 DVSS.n23158 DVSS.n23157 0.214786
R43787 DVSS.n23156 DVSS.n23155 0.214786
R43788 DVSS.n23154 DVSS.n119 0.214786
R43789 DVSS.n118 DVSS.n117 0.214786
R43790 DVSS.n23150 DVSS.n23149 0.214786
R43791 DVSS.n23148 DVSS.n23147 0.214786
R43792 DVSS.n23146 DVSS.n122 0.214786
R43793 DVSS.n23140 DVSS.n121 0.214786
R43794 DVSS.n23142 DVSS.n23141 0.214786
R43795 DVSS.n23139 DVSS.n124 0.214786
R43796 DVSS.n185 DVSS.n125 0.214786
R43797 DVSS.n23135 DVSS.n23134 0.214786
R43798 DVSS.n184 DVSS.n183 0.214786
R43799 DVSS.n23129 DVSS.n23128 0.214786
R43800 DVSS.n23126 DVSS.n191 0.214786
R43801 DVSS.n190 DVSS.n189 0.214786
R43802 DVSS.n23122 DVSS.n23121 0.214786
R43803 DVSS.n23120 DVSS.n23119 0.214786
R43804 DVSS.n23118 DVSS.n195 0.214786
R43805 DVSS.n194 DVSS.n193 0.214786
R43806 DVSS.n23114 DVSS.n23113 0.214786
R43807 DVSS.n23112 DVSS.n23111 0.214786
R43808 DVSS.n23110 DVSS.n198 0.214786
R43809 DVSS.n23104 DVSS.n197 0.214786
R43810 DVSS.n23106 DVSS.n23105 0.214786
R43811 DVSS.n23103 DVSS.n200 0.214786
R43812 DVSS.n23102 DVSS.n23101 0.214786
R43813 DVSS.n202 DVSS.n201 0.214786
R43814 DVSS.n23097 DVSS.n23096 0.214786
R43815 DVSS.n205 DVSS.n204 0.214786
R43816 DVSS.n23092 DVSS.n23091 0.214786
R43817 DVSS.n264 DVSS.n263 0.214786
R43818 DVSS.n23087 DVSS.n23086 0.214786
R43819 DVSS.n23085 DVSS.n23084 0.214786
R43820 DVSS.n23083 DVSS.n268 0.214786
R43821 DVSS.n267 DVSS.n266 0.214786
R43822 DVSS.n23079 DVSS.n23078 0.214786
R43823 DVSS.n23077 DVSS.n23076 0.214786
R43824 DVSS.n23074 DVSS.n274 0.214786
R43825 DVSS.n273 DVSS.n272 0.214786
R43826 DVSS.n22513 DVSS.n22512 0.214786
R43827 DVSS.n22516 DVSS.n22511 0.214786
R43828 DVSS.n22517 DVSS.n22510 0.214786
R43829 DVSS.n22518 DVSS.n22509 0.214786
R43830 DVSS.n22508 DVSS.n22506 0.214786
R43831 DVSS.n22522 DVSS.n22505 0.214786
R43832 DVSS.n22523 DVSS.n801 0.214786
R43833 DVSS.n22524 DVSS.n800 0.214786
R43834 DVSS.n22499 DVSS.n798 0.214786
R43835 DVSS.n22528 DVSS.n797 0.214786
R43836 DVSS.n22529 DVSS.n796 0.214786
R43837 DVSS.n22530 DVSS.n795 0.214786
R43838 DVSS.n22488 DVSS.n793 0.214786
R43839 DVSS.n22534 DVSS.n792 0.214786
R43840 DVSS.n22535 DVSS.n791 0.214786
R43841 DVSS.n22536 DVSS.n790 0.214786
R43842 DVSS.n22484 DVSS.n788 0.214786
R43843 DVSS.n22540 DVSS.n787 0.214786
R43844 DVSS.n22541 DVSS.n786 0.214786
R43845 DVSS.n22542 DVSS.n785 0.214786
R43846 DVSS.n784 DVSS.n781 0.214786
R43847 DVSS.n22546 DVSS.n780 0.214786
R43848 DVSS.n22548 DVSS.n777 0.214786
R43849 DVSS.n22549 DVSS.n776 0.214786
R43850 DVSS.n890 DVSS.n774 0.214786
R43851 DVSS.n22553 DVSS.n773 0.214786
R43852 DVSS.n22554 DVSS.n772 0.214786
R43853 DVSS.n22555 DVSS.n771 0.214786
R43854 DVSS.n894 DVSS.n769 0.214786
R43855 DVSS.n22559 DVSS.n768 0.214786
R43856 DVSS.n22560 DVSS.n767 0.214786
R43857 DVSS.n22561 DVSS.n766 0.214786
R43858 DVSS.n897 DVSS.n764 0.214786
R43859 DVSS.n22565 DVSS.n763 0.214786
R43860 DVSS.n22566 DVSS.n762 0.214786
R43861 DVSS.n22567 DVSS.n761 0.214786
R43862 DVSS.n759 DVSS.n758 0.214786
R43863 DVSS.n22568 DVSS.n22567 0.214786
R43864 DVSS.n22566 DVSS.n760 0.214786
R43865 DVSS.n22565 DVSS.n22564 0.214786
R43866 DVSS.n22563 DVSS.n764 0.214786
R43867 DVSS.n22562 DVSS.n22561 0.214786
R43868 DVSS.n22560 DVSS.n765 0.214786
R43869 DVSS.n22559 DVSS.n22558 0.214786
R43870 DVSS.n22557 DVSS.n769 0.214786
R43871 DVSS.n22556 DVSS.n22555 0.214786
R43872 DVSS.n22554 DVSS.n770 0.214786
R43873 DVSS.n22553 DVSS.n22552 0.214786
R43874 DVSS.n22551 DVSS.n774 0.214786
R43875 DVSS.n22550 DVSS.n22549 0.214786
R43876 DVSS.n22548 DVSS.n775 0.214786
R43877 DVSS.n22546 DVSS.n22545 0.214786
R43878 DVSS.n22544 DVSS.n781 0.214786
R43879 DVSS.n22543 DVSS.n22542 0.214786
R43880 DVSS.n22541 DVSS.n783 0.214786
R43881 DVSS.n22540 DVSS.n22539 0.214786
R43882 DVSS.n22538 DVSS.n788 0.214786
R43883 DVSS.n22537 DVSS.n22536 0.214786
R43884 DVSS.n22535 DVSS.n789 0.214786
R43885 DVSS.n22534 DVSS.n22533 0.214786
R43886 DVSS.n22532 DVSS.n793 0.214786
R43887 DVSS.n22531 DVSS.n22530 0.214786
R43888 DVSS.n22529 DVSS.n794 0.214786
R43889 DVSS.n22528 DVSS.n22527 0.214786
R43890 DVSS.n22526 DVSS.n798 0.214786
R43891 DVSS.n22525 DVSS.n22524 0.214786
R43892 DVSS.n22523 DVSS.n799 0.214786
R43893 DVSS.n22522 DVSS.n22521 0.214786
R43894 DVSS.n22520 DVSS.n22506 0.214786
R43895 DVSS.n22519 DVSS.n22518 0.214786
R43896 DVSS.n22517 DVSS.n22507 0.214786
R43897 DVSS.n22516 DVSS.n22515 0.214786
R43898 DVSS.n22514 DVSS.n22513 0.214786
R43899 DVSS.n275 DVSS.n273 0.214786
R43900 DVSS.n23074 DVSS.n23073 0.214786
R43901 DVSS.n23077 DVSS.n269 0.214786
R43902 DVSS.n23080 DVSS.n23079 0.214786
R43903 DVSS.n23081 DVSS.n267 0.214786
R43904 DVSS.n23083 DVSS.n23082 0.214786
R43905 DVSS.n23085 DVSS.n265 0.214786
R43906 DVSS.n23088 DVSS.n23087 0.214786
R43907 DVSS.n23089 DVSS.n264 0.214786
R43908 DVSS.n23091 DVSS.n23090 0.214786
R43909 DVSS.n204 DVSS.n203 0.214786
R43910 DVSS.n23098 DVSS.n23097 0.214786
R43911 DVSS.n23099 DVSS.n202 0.214786
R43912 DVSS.n23101 DVSS.n23100 0.214786
R43913 DVSS.n200 DVSS.n199 0.214786
R43914 DVSS.n23107 DVSS.n23106 0.214786
R43915 DVSS.n23108 DVSS.n197 0.214786
R43916 DVSS.n23110 DVSS.n23109 0.214786
R43917 DVSS.n23112 DVSS.n196 0.214786
R43918 DVSS.n23115 DVSS.n23114 0.214786
R43919 DVSS.n23116 DVSS.n194 0.214786
R43920 DVSS.n23118 DVSS.n23117 0.214786
R43921 DVSS.n23120 DVSS.n192 0.214786
R43922 DVSS.n23123 DVSS.n23122 0.214786
R43923 DVSS.n23124 DVSS.n190 0.214786
R43924 DVSS.n23126 DVSS.n23125 0.214786
R43925 DVSS.n23130 DVSS.n23129 0.214786
R43926 DVSS.n23131 DVSS.n184 0.214786
R43927 DVSS.n23134 DVSS.n23133 0.214786
R43928 DVSS.n23132 DVSS.n185 0.214786
R43929 DVSS.n124 DVSS.n123 0.214786
R43930 DVSS.n23143 DVSS.n23142 0.214786
R43931 DVSS.n23144 DVSS.n121 0.214786
R43932 DVSS.n23146 DVSS.n23145 0.214786
R43933 DVSS.n23148 DVSS.n120 0.214786
R43934 DVSS.n23151 DVSS.n23150 0.214786
R43935 DVSS.n23152 DVSS.n118 0.214786
R43936 DVSS.n23154 DVSS.n23153 0.214786
R43937 DVSS.n23156 DVSS.n116 0.214786
R43938 DVSS.n23159 DVSS.n23158 0.214786
R43939 DVSS.n23160 DVSS.n114 0.214786
R43940 DVSS.n23162 DVSS.n23161 0.214786
R43941 DVSS.n23164 DVSS.n112 0.214786
R43942 DVSS.n23175 DVSS.n23174 0.214786
R43943 DVSS.n23176 DVSS.n111 0.214786
R43944 DVSS.n23178 DVSS.n23177 0.214786
R43945 DVSS.n59 DVSS.n58 0.214786
R43946 DVSS.n23185 DVSS.n23184 0.214786
R43947 DVSS.n23186 DVSS.n57 0.214786
R43948 DVSS.n23188 DVSS.n23187 0.214786
R43949 DVSS.n23194 DVSS.n23193 0.214786
R43950 DVSS.n23195 DVSS.n50 0.214786
R43951 DVSS.n23197 DVSS.n23196 0.214786
R43952 DVSS.n23199 DVSS.n49 0.214786
R43953 DVSS.n23202 DVSS.n23201 0.214786
R43954 DVSS.n23203 DVSS.n47 0.214786
R43955 DVSS.n23205 DVSS.n23204 0.214786
R43956 DVSS.n23207 DVSS.n45 0.214786
R43957 DVSS.n23210 DVSS.n23209 0.214786
R43958 DVSS.n23211 DVSS.n44 0.214786
R43959 DVSS.n23214 DVSS.n23213 0.214786
R43960 DVSS.n23212 DVSS.n0 0.214786
R43961 DVSS.n23227 DVSS.n23226 0.214786
R43962 DVSS.n23225 DVSS.n2 0.214786
R43963 DVSS.n421 DVSS.n420 0.214786
R43964 DVSS.n12784 DVSS.n419 0.214786
R43965 DVSS.n22976 DVSS.n418 0.214786
R43966 DVSS.n22977 DVSS.n417 0.214786
R43967 DVSS.n22978 DVSS.n416 0.214786
R43968 DVSS.n12788 DVSS.n414 0.214786
R43969 DVSS.n22982 DVSS.n413 0.214786
R43970 DVSS.n22983 DVSS.n412 0.214786
R43971 DVSS.n22984 DVSS.n411 0.214786
R43972 DVSS.n12791 DVSS.n409 0.214786
R43973 DVSS.n22988 DVSS.n408 0.214786
R43974 DVSS.n22989 DVSS.n407 0.214786
R43975 DVSS.n22990 DVSS.n406 0.214786
R43976 DVSS.n12794 DVSS.n404 0.214786
R43977 DVSS.n22994 DVSS.n403 0.214786
R43978 DVSS.n22996 DVSS.n402 0.214786
R43979 DVSS.n398 DVSS.n396 0.214786
R43980 DVSS.n23001 DVSS.n23000 0.214786
R43981 DVSS.n397 DVSS.n395 0.214786
R43982 DVSS.n350 DVSS.n333 0.214786
R43983 DVSS.n21476 DVSS.n987 0.214786
R43984 DVSS.n21477 DVSS.n1001 0.214786
R43985 DVSS.n21479 DVSS.n21478 0.214786
R43986 DVSS.n1497 DVSS.n1496 0.214786
R43987 DVSS.n21483 DVSS.n1498 0.214786
R43988 DVSS.n21485 DVSS.n21484 0.214786
R43989 DVSS.n21487 DVSS.n21486 0.214786
R43990 DVSS.n1493 DVSS.n1492 0.214786
R43991 DVSS.n21491 DVSS.n1494 0.214786
R43992 DVSS.n21493 DVSS.n21492 0.214786
R43993 DVSS.n21495 DVSS.n21494 0.214786
R43994 DVSS.n1489 DVSS.n1488 0.214786
R43995 DVSS.n21499 DVSS.n1490 0.214786
R43996 DVSS.n21501 DVSS.n21500 0.214786
R43997 DVSS.n21503 DVSS.n21502 0.214786
R43998 DVSS.n21509 DVSS.n21508 0.214786
R43999 DVSS.n21510 DVSS.n1483 0.214786
R44000 DVSS.n21512 DVSS.n21511 0.214786
R44001 DVSS.n21514 DVSS.n21513 0.214786
R44002 DVSS.n1480 DVSS.n1479 0.214786
R44003 DVSS.n21518 DVSS.n1481 0.214786
R44004 DVSS.n21520 DVSS.n21519 0.214786
R44005 DVSS.n21522 DVSS.n21521 0.214786
R44006 DVSS.n1476 DVSS.n1475 0.214786
R44007 DVSS.n21526 DVSS.n1477 0.214786
R44008 DVSS.n21528 DVSS.n21527 0.214786
R44009 DVSS.n21530 DVSS.n21529 0.214786
R44010 DVSS.n1472 DVSS.n1471 0.214786
R44011 DVSS.n21534 DVSS.n1473 0.214786
R44012 DVSS.n21536 DVSS.n21535 0.214786
R44013 DVSS.n21537 DVSS.n1067 0.214786
R44014 DVSS.n1469 DVSS.n1083 0.214786
R44015 DVSS.n21543 DVSS.n21542 0.214786
R44016 DVSS.n21544 DVSS.n1468 0.214786
R44017 DVSS.n21546 DVSS.n21545 0.214786
R44018 DVSS.n21548 DVSS.n21547 0.214786
R44019 DVSS.n1465 DVSS.n1464 0.214786
R44020 DVSS.n21552 DVSS.n1466 0.214786
R44021 DVSS.n21554 DVSS.n21553 0.214786
R44022 DVSS.n23069 DVSS.n279 0.214786
R44023 DVSS.n23068 DVSS.n280 0.214786
R44024 DVSS.n23067 DVSS.n281 0.214786
R44025 DVSS.n1120 DVSS.n282 0.214786
R44026 DVSS.n23063 DVSS.n284 0.214786
R44027 DVSS.n23062 DVSS.n285 0.214786
R44028 DVSS.n23061 DVSS.n286 0.214786
R44029 DVSS.n1123 DVSS.n287 0.214786
R44030 DVSS.n23057 DVSS.n289 0.214786
R44031 DVSS.n23056 DVSS.n290 0.214786
R44032 DVSS.n23055 DVSS.n291 0.214786
R44033 DVSS.n294 DVSS.n292 0.214786
R44034 DVSS.n23051 DVSS.n295 0.214786
R44035 DVSS.n23050 DVSS.n296 0.214786
R44036 DVSS.n23049 DVSS.n297 0.214786
R44037 DVSS.n12980 DVSS.n298 0.214786
R44038 DVSS.n23045 DVSS.n300 0.214786
R44039 DVSS.n23044 DVSS.n301 0.214786
R44040 DVSS.n23043 DVSS.n302 0.214786
R44041 DVSS.n12983 DVSS.n303 0.214786
R44042 DVSS.n23039 DVSS.n305 0.214786
R44043 DVSS.n23038 DVSS.n306 0.214786
R44044 DVSS.n23037 DVSS.n307 0.214786
R44045 DVSS.n12986 DVSS.n308 0.214786
R44046 DVSS.n23032 DVSS.n310 0.214786
R44047 DVSS.n23031 DVSS.n311 0.214786
R44048 DVSS.n23030 DVSS.n312 0.214786
R44049 DVSS.n12990 DVSS.n313 0.214786
R44050 DVSS.n23026 DVSS.n315 0.214786
R44051 DVSS.n23025 DVSS.n316 0.214786
R44052 DVSS.n23024 DVSS.n317 0.214786
R44053 DVSS.n382 DVSS.n318 0.214786
R44054 DVSS.n23020 DVSS.n320 0.214786
R44055 DVSS.n23019 DVSS.n321 0.214786
R44056 DVSS.n23018 DVSS.n322 0.214786
R44057 DVSS.n388 DVSS.n323 0.214786
R44058 DVSS.n23014 DVSS.n325 0.214786
R44059 DVSS.n23013 DVSS.n326 0.214786
R44060 DVSS.n23012 DVSS.n327 0.214786
R44061 DVSS.n391 DVSS.n328 0.214786
R44062 DVSS.n23008 DVSS.n330 0.214786
R44063 DVSS.n23007 DVSS.n331 0.214786
R44064 DVSS.n22974 DVSS.n419 0.214786
R44065 DVSS.n22976 DVSS.n22975 0.214786
R44066 DVSS.n22977 DVSS.n415 0.214786
R44067 DVSS.n22979 DVSS.n22978 0.214786
R44068 DVSS.n22980 DVSS.n414 0.214786
R44069 DVSS.n22982 DVSS.n22981 0.214786
R44070 DVSS.n22983 DVSS.n410 0.214786
R44071 DVSS.n22985 DVSS.n22984 0.214786
R44072 DVSS.n22986 DVSS.n409 0.214786
R44073 DVSS.n22988 DVSS.n22987 0.214786
R44074 DVSS.n22989 DVSS.n405 0.214786
R44075 DVSS.n22991 DVSS.n22990 0.214786
R44076 DVSS.n22992 DVSS.n404 0.214786
R44077 DVSS.n22994 DVSS.n22993 0.214786
R44078 DVSS.n22997 DVSS.n22996 0.214786
R44079 DVSS.n22998 DVSS.n398 0.214786
R44080 DVSS.n23000 DVSS.n22999 0.214786
R44081 DVSS.n400 DVSS.n397 0.214786
R44082 DVSS.n399 DVSS.n333 0.214786
R44083 DVSS.n21477 DVSS.n1499 0.214786
R44084 DVSS.n21480 DVSS.n21479 0.214786
R44085 DVSS.n21481 DVSS.n1497 0.214786
R44086 DVSS.n21483 DVSS.n21482 0.214786
R44087 DVSS.n21485 DVSS.n1495 0.214786
R44088 DVSS.n21488 DVSS.n21487 0.214786
R44089 DVSS.n21489 DVSS.n1493 0.214786
R44090 DVSS.n21491 DVSS.n21490 0.214786
R44091 DVSS.n21493 DVSS.n1491 0.214786
R44092 DVSS.n21496 DVSS.n21495 0.214786
R44093 DVSS.n21497 DVSS.n1489 0.214786
R44094 DVSS.n21499 DVSS.n21498 0.214786
R44095 DVSS.n21500 DVSS.n1487 0.214786
R44096 DVSS.n21504 DVSS.n21503 0.214786
R44097 DVSS.n21508 DVSS.n21507 0.214786
R44098 DVSS.n21506 DVSS.n1483 0.214786
R44099 DVSS.n21512 DVSS.n1482 0.214786
R44100 DVSS.n21515 DVSS.n21514 0.214786
R44101 DVSS.n21516 DVSS.n1480 0.214786
R44102 DVSS.n21518 DVSS.n21517 0.214786
R44103 DVSS.n21520 DVSS.n1478 0.214786
R44104 DVSS.n21523 DVSS.n21522 0.214786
R44105 DVSS.n21524 DVSS.n1476 0.214786
R44106 DVSS.n21526 DVSS.n21525 0.214786
R44107 DVSS.n21528 DVSS.n1474 0.214786
R44108 DVSS.n21531 DVSS.n21530 0.214786
R44109 DVSS.n21532 DVSS.n1472 0.214786
R44110 DVSS.n21534 DVSS.n21533 0.214786
R44111 DVSS.n21536 DVSS.n1470 0.214786
R44112 DVSS.n21538 DVSS.n21537 0.214786
R44113 DVSS.n21539 DVSS.n1469 0.214786
R44114 DVSS.n21542 DVSS.n21541 0.214786
R44115 DVSS.n21540 DVSS.n1468 0.214786
R44116 DVSS.n21546 DVSS.n1467 0.214786
R44117 DVSS.n21549 DVSS.n21548 0.214786
R44118 DVSS.n21550 DVSS.n1465 0.214786
R44119 DVSS.n21552 DVSS.n21551 0.214786
R44120 DVSS.n21553 DVSS.n277 0.214786
R44121 DVSS.n23070 DVSS.n23069 0.214786
R44122 DVSS.n23068 DVSS.n278 0.214786
R44123 DVSS.n23067 DVSS.n23066 0.214786
R44124 DVSS.n23065 DVSS.n282 0.214786
R44125 DVSS.n23064 DVSS.n23063 0.214786
R44126 DVSS.n23062 DVSS.n283 0.214786
R44127 DVSS.n23061 DVSS.n23060 0.214786
R44128 DVSS.n23059 DVSS.n287 0.214786
R44129 DVSS.n23058 DVSS.n23057 0.214786
R44130 DVSS.n23056 DVSS.n288 0.214786
R44131 DVSS.n23055 DVSS.n23054 0.214786
R44132 DVSS.n23053 DVSS.n292 0.214786
R44133 DVSS.n23052 DVSS.n23051 0.214786
R44134 DVSS.n23050 DVSS.n293 0.214786
R44135 DVSS.n23049 DVSS.n23048 0.214786
R44136 DVSS.n23047 DVSS.n298 0.214786
R44137 DVSS.n23046 DVSS.n23045 0.214786
R44138 DVSS.n23044 DVSS.n299 0.214786
R44139 DVSS.n23043 DVSS.n23042 0.214786
R44140 DVSS.n23041 DVSS.n303 0.214786
R44141 DVSS.n23040 DVSS.n23039 0.214786
R44142 DVSS.n23038 DVSS.n304 0.214786
R44143 DVSS.n23037 DVSS.n23036 0.214786
R44144 DVSS.n23035 DVSS.n308 0.214786
R44145 DVSS.n23033 DVSS.n23032 0.214786
R44146 DVSS.n23031 DVSS.n309 0.214786
R44147 DVSS.n23030 DVSS.n23029 0.214786
R44148 DVSS.n23028 DVSS.n313 0.214786
R44149 DVSS.n23027 DVSS.n23026 0.214786
R44150 DVSS.n23025 DVSS.n314 0.214786
R44151 DVSS.n23024 DVSS.n23023 0.214786
R44152 DVSS.n23022 DVSS.n318 0.214786
R44153 DVSS.n23021 DVSS.n23020 0.214786
R44154 DVSS.n23019 DVSS.n319 0.214786
R44155 DVSS.n23018 DVSS.n23017 0.214786
R44156 DVSS.n23016 DVSS.n323 0.214786
R44157 DVSS.n23015 DVSS.n23014 0.214786
R44158 DVSS.n23013 DVSS.n324 0.214786
R44159 DVSS.n23012 DVSS.n23011 0.214786
R44160 DVSS.n23010 DVSS.n328 0.214786
R44161 DVSS.n23009 DVSS.n23008 0.214786
R44162 DVSS.n23007 DVSS.n329 0.214786
R44163 DVSS.n23006 DVSS.n332 0.214786
R44164 DVSS.n23006 DVSS.n23005 0.214786
R44165 DVSS.n21172 DVSS.n13665 0.209612
R44166 DVSS.n1333 DVSS.n1332 0.20887
R44167 DVSS.n1292 DVSS.n1291 0.20887
R44168 DVSS.n22459 DVSS.n869 0.20887
R44169 DVSS.n22338 DVSS.n22337 0.20887
R44170 DVSS.n19503 DVSS.n19502 0.20887
R44171 DVSS.n19849 DVSS.n19848 0.20887
R44172 DVSS.n13095 DVSS.n13094 0.202266
R44173 DVSS.n20848 DVSS.n14470 0.201178
R44174 DVSS.n20889 DVSS.n14425 0.201178
R44175 DVSS.n20804 DVSS.n20699 0.201178
R44176 DVSS.n20929 DVSS.n14376 0.201178
R44177 DVSS.n21161 DVSS.n21160 0.199543
R44178 DVSS.n17036 DVSS.n17035 0.189014
R44179 DVSS.n16995 DVSS.n16994 0.189014
R44180 DVSS.n17101 DVSS.n17100 0.189014
R44181 DVSS.n17077 DVSS.n16909 0.189014
R44182 DVSS.n18820 DVSS.t189 0.187174
R44183 DVSS.n18708 DVSS.t168 0.187174
R44184 DVSS.n14578 DVSS.t169 0.187174
R44185 DVSS.n14578 DVSS.t168 0.187174
R44186 DVSS.n14577 DVSS.t0 0.187174
R44187 DVSS.n14577 DVSS.t189 0.187174
R44188 DVSS.n14622 DVSS.t174 0.187174
R44189 DVSS.n14622 DVSS.t169 0.187174
R44190 DVSS.n14621 DVSS.t1 0.187174
R44191 DVSS.n14621 DVSS.t0 0.187174
R44192 DVSS.n14662 DVSS.t175 0.187174
R44193 DVSS.n14662 DVSS.t174 0.187174
R44194 DVSS.n14661 DVSS.t184 0.187174
R44195 DVSS.n14661 DVSS.t1 0.187174
R44196 DVSS.n20489 DVSS.t175 0.187174
R44197 DVSS.n14740 DVSS.t184 0.187174
R44198 DVSS.n1313 DVSS.n1312 0.186859
R44199 DVSS.n1312 DVSS.n1311 0.186859
R44200 DVSS.n22341 DVSS.n1176 0.186859
R44201 DVSS.n22341 DVSS.n22340 0.186859
R44202 DVSS.n19594 DVSS.n19593 0.186859
R44203 DVSS.n19594 DVSS.n19078 0.186859
R44204 DVSS.n18526 DVSS.n18525 0.183303
R44205 DVSS.n19917 DVSS.n19916 0.183303
R44206 DVSS.n19003 DVSS.n19001 0.17981
R44207 DVSS.n19001 DVSS.n18998 0.17981
R44208 DVSS.n19204 DVSS.n19203 0.173833
R44209 DVSS.n19189 DVSS.n19186 0.172918
R44210 DVSS.n21463 DVSS.n21462 0.17013
R44211 DVSS.n22961 DVSS.n22960 0.16989
R44212 DVSS.n21026 DVSS.n21025 0.159572
R44213 DVSS.n22972 DVSS.n22971 0.159572
R44214 DVSS.n22950 DVSS.n3 0.159572
R44215 DVSS.n21988 DVSS.n442 0.159572
R44216 DVSS.n13788 DVSS.n13682 0.159452
R44217 DVSS.n21474 DVSS.n21473 0.159452
R44218 DVSS.n22571 DVSS.n22570 0.159452
R44219 DVSS.n1408 DVSS.n744 0.159452
R44220 DVSS.n18511 DVSS.n18510 0.159115
R44221 DVSS.n13677 DVSS.n13669 0.159115
R44222 DVSS.n18515 DVSS.n18498 0.158395
R44223 DVSS.n18511 DVSS.n18498 0.158395
R44224 DVSS.n21169 DVSS.n13669 0.158395
R44225 DVSS.n21170 DVSS.n21169 0.158395
R44226 DVSS.n17016 DVSS.n17015 0.154959
R44227 DVSS.n17015 DVSS.n17014 0.154959
R44228 DVSS.n17098 DVSS.n17097 0.154959
R44229 DVSS.n17097 DVSS.n17096 0.154959
R44230 DVSS.n15918 DVSS.n15888 0.154827
R44231 DVSS.n15917 DVSS.n15848 0.154827
R44232 DVSS.n15795 DVSS.n15539 0.154827
R44233 DVSS.n18163 DVSS.n15538 0.154827
R44234 DVSS.n18164 DVSS.n15537 0.154827
R44235 DVSS.n18165 DVSS.n15536 0.154827
R44236 DVSS.n21447 DVSS.n1501 0.154827
R44237 DVSS.n21446 DVSS.n1502 0.154827
R44238 DVSS.n21445 DVSS.n1503 0.154827
R44239 DVSS.n13366 DVSS.n1504 0.154827
R44240 DVSS.n13365 DVSS.n13364 0.154827
R44241 DVSS.n13101 DVSS.n423 0.154827
R44242 DVSS.n20986 DVSS.n20985 0.150957
R44243 DVSS.n21157 DVSS.n21155 0.15089
R44244 DVSS.n21161 DVSS.n13682 0.149792
R44245 DVSS.n19209 DVSS 0.149572
R44246 DVSS.n19183 DVSS 0.149572
R44247 DVSS.n19182 DVSS 0.149572
R44248 DVSS.n19211 DVSS 0.149479
R44249 DVSS.n19174 DVSS 0.149479
R44250 DVSS.n19188 DVSS 0.149479
R44251 DVSS.n19185 DVSS 0.149479
R44252 DVSS.n17383 DVSS.n17053 0.148831
R44253 DVSS.n17424 DVSS.n16929 0.148831
R44254 DVSS.n17787 DVSS.n17786 0.146974
R44255 DVSS.n18172 DVSS.n18171 0.146974
R44256 DVSS.n21153 DVSS.n13686 0.146893
R44257 DVSS.n19000 DVSS.n18999 0.144944
R44258 DVSS.n19178 DVSS.n19000 0.144944
R44259 DVSS.n20469 DVSS.n14714 0.137755
R44260 DVSS DVSS.n16471 0.131883
R44261 DVSS DVSS.n18089 0.131883
R44262 DVSS.n21106 DVSS.n13947 0.130407
R44263 DVSS.n14631 DVSS.n14031 0.130407
R44264 DVSS.n20688 DVSS.n13836 0.130407
R44265 DVSS.n14668 DVSS.n14137 0.130407
R44266 DVSS.n18527 DVSS.n18526 0.122586
R44267 DVSS.n19916 DVSS.n19915 0.122586
R44268 DVSS.n22974 DVSS.n22973 0.114699
R44269 DVSS.n21175 DVSS.n13664 0.114607
R44270 DVSS.n17481 DVSS.n17117 0.113608
R44271 DVSS.n17382 DVSS.n17117 0.113608
R44272 DVSS.n17380 DVSS.n17052 0.113608
R44273 DVSS.n17052 DVSS.n17051 0.113608
R44274 DVSS.n17523 DVSS.n16933 0.113608
R44275 DVSS.n17523 DVSS.n17522 0.113608
R44276 DVSS.n17522 DVSS.n16934 0.113608
R44277 DVSS.n16979 DVSS.n16934 0.113608
R44278 DVSS.n17382 DVSS.n17381 0.113608
R44279 DVSS.n17381 DVSS.n17380 0.113608
R44280 DVSS.n17528 DVSS.n17527 0.113608
R44281 DVSS.n17527 DVSS.n16924 0.113608
R44282 DVSS.n16932 DVSS.n16924 0.113608
R44283 DVSS.n16933 DVSS.n16932 0.113608
R44284 DVSS.n17482 DVSS.n17116 0.113608
R44285 DVSS.n17482 DVSS.n17481 0.113608
R44286 DVSS.n17405 DVSS.n17404 0.111803
R44287 DVSS.n17418 DVSS.n17417 0.111803
R44288 DVSS.n17371 DVSS.n17370 0.111803
R44289 DVSS.n17494 DVSS.n17493 0.111803
R44290 DVSS.n17478 DVSS.n17477 0.111803
R44291 DVSS.n17469 DVSS.n17457 0.111803
R44292 DVSS.n21475 DVSS.n1499 0.110647
R44293 DVSS.n22569 DVSS.n22568 0.110647
R44294 DVSS.n1410 DVSS.n1409 0.110647
R44295 DVSS.n23225 DVSS.n23224 0.110634
R44296 DVSS.n21992 DVSS.n21991 0.110634
R44297 DVSS.n13793 DVSS.n13787 0.110634
R44298 DVSS.n14308 DVSS.n14307 0.110634
R44299 DVSS.n19197 DVSS.n19177 0.108833
R44300 DVSS.n19180 DVSS.n19177 0.108833
R44301 DVSS.n16493 DVSS.n15899 0.106064
R44302 DVSS.n18155 DVSS.n15545 0.105653
R44303 DVSS.n19900 DVSS.n19030 0.104685
R44304 DVSS.n19626 DVSS.n19624 0.104685
R44305 DVSS.n22384 DVSS.n1043 0.104685
R44306 DVSS.n13091 DVSS.n13089 0.104685
R44307 DVSS.n22965 DVSS.n425 0.100706
R44308 DVSS.n22966 DVSS.n22965 0.100706
R44309 DVSS.n22967 DVSS.n22966 0.100706
R44310 DVSS.n22967 DVSS.n422 0.100706
R44311 DVSS.n22937 DVSS.n433 0.100706
R44312 DVSS.n22942 DVSS.n433 0.100706
R44313 DVSS.n22943 DVSS.n22942 0.100706
R44314 DVSS.n22944 DVSS.n22943 0.100706
R44315 DVSS.n22944 DVSS.n431 0.100706
R44316 DVSS.n22948 DVSS.n431 0.100706
R44317 DVSS.n22949 DVSS.n22948 0.100706
R44318 DVSS.n22951 DVSS.n429 0.100706
R44319 DVSS.n22955 DVSS.n429 0.100706
R44320 DVSS.n22956 DVSS.n22955 0.100706
R44321 DVSS.n22956 DVSS.n427 0.100706
R44322 DVSS.n22895 DVSS.n448 0.100706
R44323 DVSS.n22900 DVSS.n448 0.100706
R44324 DVSS.n22901 DVSS.n22900 0.100706
R44325 DVSS.n22902 DVSS.n22901 0.100706
R44326 DVSS.n22902 DVSS.n446 0.100706
R44327 DVSS.n22906 DVSS.n446 0.100706
R44328 DVSS.n22907 DVSS.n22906 0.100706
R44329 DVSS.n22908 DVSS.n22907 0.100706
R44330 DVSS.n22908 DVSS.n444 0.100706
R44331 DVSS.n22912 DVSS.n444 0.100706
R44332 DVSS.n22913 DVSS.n22912 0.100706
R44333 DVSS.n22917 DVSS.n22916 0.100706
R44334 DVSS.n22917 DVSS.n440 0.100706
R44335 DVSS.n22921 DVSS.n440 0.100706
R44336 DVSS.n22922 DVSS.n22921 0.100706
R44337 DVSS.n22923 DVSS.n22922 0.100706
R44338 DVSS.n22923 DVSS.n438 0.100706
R44339 DVSS.n22927 DVSS.n438 0.100706
R44340 DVSS.n22928 DVSS.n22927 0.100706
R44341 DVSS.n22929 DVSS.n22928 0.100706
R44342 DVSS.n22929 DVSS.n436 0.100706
R44343 DVSS.n22934 DVSS.n436 0.100706
R44344 DVSS.n18169 DVSS.n15532 0.100706
R44345 DVSS.n18173 DVSS.n15532 0.100706
R44346 DVSS.n17789 DVSS.n15921 0.100706
R44347 DVSS.n17785 DVSS.n15921 0.100706
R44348 DVSS.n19918 DVSS.n15140 0.100706
R44349 DVSS.n19919 DVSS.n19918 0.100706
R44350 DVSS.n19920 DVSS.n19919 0.100706
R44351 DVSS.n19920 DVSS.n15138 0.100706
R44352 DVSS.n19924 DVSS.n15138 0.100706
R44353 DVSS.n18524 DVSS.n15146 0.100706
R44354 DVSS.n18524 DVSS.n18523 0.100706
R44355 DVSS.n18523 DVSS.n18522 0.100706
R44356 DVSS.n18522 DVSS.n15148 0.100706
R44357 DVSS.n18518 DVSS.n15148 0.100706
R44358 DVSS.n15135 DVSS.n15127 0.100706
R44359 DVSS.n15130 DVSS.n15127 0.100706
R44360 DVSS.n15130 DVSS.n15129 0.100706
R44361 DVSS.n15129 DVSS.n14315 0.100706
R44362 DVSS.n20984 DVSS.n14315 0.100706
R44363 DVSS.n18508 DVSS.n18507 0.100706
R44364 DVSS.n20990 DVSS.n14312 0.100706
R44365 DVSS.n20991 DVSS.n20990 0.100706
R44366 DVSS.n20992 DVSS.n20991 0.100706
R44367 DVSS.n20992 DVSS.n14309 0.100706
R44368 DVSS.n21024 DVSS.n14310 0.100706
R44369 DVSS.n21020 DVSS.n14310 0.100706
R44370 DVSS.n21020 DVSS.n21019 0.100706
R44371 DVSS.n21019 DVSS.n21018 0.100706
R44372 DVSS.n21018 DVSS.n20996 0.100706
R44373 DVSS.n21011 DVSS.n20996 0.100706
R44374 DVSS.n21012 DVSS.n21011 0.100706
R44375 DVSS.n21160 DVSS.n13683 0.100706
R44376 DVSS.n13680 DVSS.n13676 0.100706
R44377 DVSS.n21008 DVSS.n21000 0.100706
R44378 DVSS.n21003 DVSS.n21000 0.100706
R44379 DVSS.n21003 DVSS.n21002 0.100706
R44380 DVSS.n21002 DVSS.n13372 0.100706
R44381 DVSS.n21438 DVSS.n13372 0.100706
R44382 DVSS.n13666 DVSS.n13659 0.100706
R44383 DVSS.n21179 DVSS.n13659 0.100706
R44384 DVSS.n21179 DVSS.n13660 0.100706
R44385 DVSS.n22886 DVSS.n22885 0.100706
R44386 DVSS.n22887 DVSS.n22886 0.100706
R44387 DVSS.n22887 DVSS.n451 0.100706
R44388 DVSS.n22892 DVSS.n451 0.100706
R44389 DVSS.n22637 DVSS.n733 0.100706
R44390 DVSS.n22633 DVSS.n733 0.100706
R44391 DVSS.n22633 DVSS.n22632 0.100706
R44392 DVSS.n22632 DVSS.n736 0.100706
R44393 DVSS.n22626 DVSS.n738 0.100706
R44394 DVSS.n22621 DVSS.n738 0.100706
R44395 DVSS.n22621 DVSS.n22620 0.100706
R44396 DVSS.n22620 DVSS.n22619 0.100706
R44397 DVSS.n22619 DVSS.n740 0.100706
R44398 DVSS.n22615 DVSS.n740 0.100706
R44399 DVSS.n22615 DVSS.n22614 0.100706
R44400 DVSS.n22614 DVSS.n22613 0.100706
R44401 DVSS.n22613 DVSS.n742 0.100706
R44402 DVSS.n22609 DVSS.n742 0.100706
R44403 DVSS.n22609 DVSS.n22608 0.100706
R44404 DVSS.n22605 DVSS.n22604 0.100706
R44405 DVSS.n22604 DVSS.n746 0.100706
R44406 DVSS.n22600 DVSS.n746 0.100706
R44407 DVSS.n22600 DVSS.n22599 0.100706
R44408 DVSS.n22599 DVSS.n22598 0.100706
R44409 DVSS.n22598 DVSS.n748 0.100706
R44410 DVSS.n22594 DVSS.n748 0.100706
R44411 DVSS.n22594 DVSS.n22593 0.100706
R44412 DVSS.n22593 DVSS.n22592 0.100706
R44413 DVSS.n22592 DVSS.n750 0.100706
R44414 DVSS.n22587 DVSS.n750 0.100706
R44415 DVSS.n22584 DVSS.n753 0.100706
R44416 DVSS.n22579 DVSS.n753 0.100706
R44417 DVSS.n22579 DVSS.n22578 0.100706
R44418 DVSS.n22578 DVSS.n22577 0.100706
R44419 DVSS.n22577 DVSS.n755 0.100706
R44420 DVSS.n22573 DVSS.n755 0.100706
R44421 DVSS.n22573 DVSS.n22572 0.100706
R44422 DVSS.n21455 DVSS.n757 0.100706
R44423 DVSS.n21456 DVSS.n21455 0.100706
R44424 DVSS.n21456 DVSS.n21452 0.100706
R44425 DVSS.n21461 DVSS.n21452 0.100706
R44426 DVSS.n21467 DVSS.n21449 0.100706
R44427 DVSS.n21468 DVSS.n21467 0.100706
R44428 DVSS.n21469 DVSS.n21468 0.100706
R44429 DVSS.n21469 DVSS.n1500 0.100706
R44430 DVSS.n18159 DVSS.n15541 0.0975237
R44431 DVSS.n19596 DVSS.n19250 0.0936793
R44432 DVSS.n19598 DVSS.n19596 0.0936793
R44433 DVSS.n22370 DVSS.n22343 0.0936793
R44434 DVSS.n22343 DVSS.n1175 0.0936793
R44435 DVSS.n17776 DVSS.n17775 0.0933421
R44436 DVSS.n18491 DVSS.n15164 0.0933421
R44437 DVSS.n18207 DVSS.n18206 0.0933421
R44438 DVSS.n18275 DVSS.n15093 0.0933421
R44439 DVSS DVSS.t53 0.092694
R44440 DVSS DVSS.t121 0.092694
R44441 DVSS DVSS.t157 0.092694
R44442 DVSS DVSS.t61 0.092694
R44443 DVSS DVSS.t67 0.092694
R44444 DVSS DVSS.t155 0.092694
R44445 DVSS DVSS.t21 0.092694
R44446 DVSS DVSS.t65 0.092694
R44447 DVSS.n21383 DVSS.n13430 0.0921244
R44448 DVSS.n20173 DVSS.n20009 0.091861
R44449 DVSS.n20316 DVSS.n14864 0.091861
R44450 DVSS.n20697 DVSS.n14536 0.091861
R44451 DVSS.n20458 DVSS.n14853 0.091861
R44452 DVSS.n17412 DVSS.n17409 0.0916968
R44453 DVSS.n17413 DVSS.n17412 0.0916968
R44454 DVSS.n17488 DVSS.n16974 0.0916968
R44455 DVSS.n17489 DVSS.n17488 0.0916968
R44456 DVSS.n17474 DVSS.n17473 0.0916968
R44457 DVSS.n17473 DVSS.n17471 0.0916968
R44458 DVSS.n20673 DVSS.n13527 0.0908951
R44459 DVSS.n20647 DVSS.n13481 0.0908951
R44460 DVSS.n14548 DVSS.n13581 0.0908951
R44461 DVSS.n21174 DVSS.n13665 0.0901892
R44462 DVSS.n21173 DVSS.n13664 0.08969
R44463 DVSS.n13671 DVSS.n13668 0.08969
R44464 DVSS.n21168 DVSS.n21167 0.08969
R44465 DVSS.n21166 DVSS.n13670 0.08969
R44466 DVSS.n21165 DVSS.n21164 0.08969
R44467 DVSS.n21163 DVSS.n13672 0.08969
R44468 DVSS.n18501 DVSS.n13674 0.08969
R44469 DVSS.n18503 DVSS.n18502 0.08969
R44470 DVSS.n18504 DVSS.n18500 0.08969
R44471 DVSS.n18513 DVSS.n18512 0.08969
R44472 DVSS.n16243 DVSS.n15790 0.0865927
R44473 DVSS.n16167 DVSS.n15743 0.0865927
R44474 DVSS.n20007 DVSS.n14903 0.0865488
R44475 DVSS.n19982 DVSS.n14938 0.0865488
R44476 DVSS.n18473 DVSS.n18381 0.0865488
R44477 DVSS.n19971 DVSS.n15011 0.0865488
R44478 DVSS.n17790 DVSS.n15920 0.0785115
R44479 DVSS.n18168 DVSS.n15533 0.0785115
R44480 DVSS.n22586 DVSS.n22585 0.0776868
R44481 DVSS.n22936 DVSS.n22935 0.0776868
R44482 DVSS.n13679 DVSS.n13678 0.0758488
R44483 DVSS.n21466 DVSS.n21450 0.0758488
R44484 DVSS.n21460 DVSS.n21459 0.0758488
R44485 DVSS.n22583 DVSS.n22582 0.0758488
R44486 DVSS.n22589 DVSS.n22588 0.0758488
R44487 DVSS.n22607 DVSS.n22606 0.0758488
R44488 DVSS.n22625 DVSS.n22624 0.0758488
R44489 DVSS.n22631 DVSS.n22630 0.0758488
R44490 DVSS.n21159 DVSS.n21158 0.0758488
R44491 DVSS.n18506 DVSS.n18505 0.0758488
R44492 DVSS.n15134 DVSS.n15133 0.0758488
R44493 DVSS.n20989 DVSS.n14313 0.0758488
R44494 DVSS.n20998 DVSS.n20997 0.0758488
R44495 DVSS.n21007 DVSS.n21006 0.0758488
R44496 DVSS.n22891 DVSS.n22890 0.0758488
R44497 DVSS.n22897 DVSS.n22896 0.0758488
R44498 DVSS.n22915 DVSS.n22914 0.0758488
R44499 DVSS.n22933 DVSS.n22932 0.0758488
R44500 DVSS.n22939 DVSS.n22938 0.0758488
R44501 DVSS.n22958 DVSS.n22957 0.0758488
R44502 DVSS.n22964 DVSS.n426 0.0758488
R44503 DVSS.n18992 DVSS.n18647 0.0758261
R44504 DVSS.n20618 DVSS.n14703 0.0758261
R44505 DVSS.n18768 DVSS.n18767 0.0758261
R44506 DVSS.n20465 DVSS.n20463 0.0758261
R44507 DVSS.n21472 DVSS.n21471 0.0758118
R44508 DVSS.n22970 DVSS.n22969 0.0758118
R44509 DVSS.n21176 DVSS.n13662 0.0745984
R44510 DVSS.n16472 DVSS 0.0734261
R44511 DVSS.n18113 DVSS 0.0734261
R44512 DVSS.n19313 DVSS.n13624 0.0727368
R44513 DVSS.n21431 DVSS.n13399 0.0727368
R44514 DVSS.n18159 DVSS.n18158 0.0702987
R44515 DVSS.n21010 DVSS.n21009 0.068
R44516 DVSS.n15812 DVSS.n15542 0.0651698
R44517 DVSS.n18157 DVSS.n15543 0.0651698
R44518 DVSS.n16492 DVSS.n15857 0.0651698
R44519 DVSS.n18156 DVSS.n15544 0.0651698
R44520 DVSS.n13052 DVSS.n13051 0.0640746
R44521 DVSS.n13031 DVSS.n13030 0.0640746
R44522 DVSS.n13043 DVSS.n13042 0.0640746
R44523 DVSS.n22481 DVSS.n246 0.0640746
R44524 DVSS.n820 DVSS.n819 0.0640746
R44525 DVSS.n829 DVSS.n828 0.0640746
R44526 DVSS.n838 DVSS.n837 0.0640746
R44527 DVSS.n847 DVSS.n846 0.0640746
R44528 DVSS.n855 DVSS.n854 0.0640746
R44529 DVSS.n21887 DVSS.n21886 0.0640746
R44530 DVSS.n21897 DVSS.n21896 0.0640746
R44531 DVSS.n21907 DVSS.n21906 0.0640746
R44532 DVSS.n21917 DVSS.n21916 0.0640746
R44533 DVSS.n21939 DVSS.n21938 0.0640746
R44534 DVSS.n21947 DVSS.n21629 0.0640746
R44535 DVSS.n21848 DVSS.n21603 0.0640746
R44536 DVSS.n21844 DVSS.n21843 0.0640746
R44537 DVSS.n21842 DVSS.n21841 0.0640746
R44538 DVSS.n21831 DVSS.n21827 0.0640746
R44539 DVSS.n663 DVSS.n662 0.0640746
R44540 DVSS.n19546 DVSS.n19539 0.0640746
R44541 DVSS.n19550 DVSS.n19549 0.0640746
R44542 DVSS.n19552 DVSS.n19551 0.0640746
R44543 DVSS.n19559 DVSS.n19531 0.0640746
R44544 DVSS.n19563 DVSS.n19562 0.0640746
R44545 DVSS.n19565 DVSS.n19564 0.0640746
R44546 DVSS.n19572 DVSS.n19523 0.0640746
R44547 DVSS.n19576 DVSS.n19575 0.0640746
R44548 DVSS.n19578 DVSS.n19577 0.0640746
R44549 DVSS.n19585 DVSS.n19268 0.0640746
R44550 DVSS.n19589 DVSS.n19588 0.0640746
R44551 DVSS.n19854 DVSS.n19853 0.0640746
R44552 DVSS.n19856 DVSS.n19855 0.0640746
R44553 DVSS.n19859 DVSS.n19057 0.0640746
R44554 DVSS.n19867 DVSS.n19866 0.0640746
R44555 DVSS.n19869 DVSS.n19868 0.0640746
R44556 DVSS.n19872 DVSS.n19049 0.0640746
R44557 DVSS.n19880 DVSS.n19879 0.0640746
R44558 DVSS.n19882 DVSS.n19881 0.0640746
R44559 DVSS.n19885 DVSS.n19042 0.0640746
R44560 DVSS.n19893 DVSS.n19892 0.0640746
R44561 DVSS.n19895 DVSS.n19894 0.0640746
R44562 DVSS.n13020 DVSS.n13019 0.0640746
R44563 DVSS.n13055 DVSS.n13054 0.0640746
R44564 DVSS.n13034 DVSS.n13033 0.0640746
R44565 DVSS.n13046 DVSS.n13045 0.0640746
R44566 DVSS.n22479 DVSS.n166 0.0640746
R44567 DVSS.n817 DVSS.n816 0.0640746
R44568 DVSS.n826 DVSS.n825 0.0640746
R44569 DVSS.n835 DVSS.n834 0.0640746
R44570 DVSS.n844 DVSS.n843 0.0640746
R44571 DVSS.n853 DVSS.n852 0.0640746
R44572 DVSS.n21885 DVSS.n21884 0.0640746
R44573 DVSS.n21894 DVSS.n21893 0.0640746
R44574 DVSS.n21904 DVSS.n21903 0.0640746
R44575 DVSS.n21914 DVSS.n21913 0.0640746
R44576 DVSS.n21936 DVSS.n21935 0.0640746
R44577 DVSS.n21949 DVSS.n21733 0.0640746
R44578 DVSS.n21846 DVSS.n21706 0.0640746
R44579 DVSS.n21837 DVSS.n21836 0.0640746
R44580 DVSS.n21839 DVSS.n21838 0.0640746
R44581 DVSS.n21834 DVSS.n21833 0.0640746
R44582 DVSS.n661 DVSS.n660 0.0640746
R44583 DVSS.n19545 DVSS.n19544 0.0640746
R44584 DVSS.n19541 DVSS.n19537 0.0640746
R44585 DVSS.n19555 DVSS.n19554 0.0640746
R44586 DVSS.n19557 DVSS.n19556 0.0640746
R44587 DVSS.n19534 DVSS.n19529 0.0640746
R44588 DVSS.n19568 DVSS.n19567 0.0640746
R44589 DVSS.n19570 DVSS.n19569 0.0640746
R44590 DVSS.n19526 DVSS.n19521 0.0640746
R44591 DVSS.n19581 DVSS.n19580 0.0640746
R44592 DVSS.n19583 DVSS.n19582 0.0640746
R44593 DVSS.n19520 DVSS.n19519 0.0640746
R44594 DVSS.n19852 DVSS.n19851 0.0640746
R44595 DVSS.n19066 DVSS.n19061 0.0640746
R44596 DVSS.n19862 DVSS.n19861 0.0640746
R44597 DVSS.n19864 DVSS.n19863 0.0640746
R44598 DVSS.n19058 DVSS.n19053 0.0640746
R44599 DVSS.n19875 DVSS.n19874 0.0640746
R44600 DVSS.n19877 DVSS.n19876 0.0640746
R44601 DVSS.n19050 DVSS.n19045 0.0640746
R44602 DVSS.n19888 DVSS.n19887 0.0640746
R44603 DVSS.n19890 DVSS.n19889 0.0640746
R44604 DVSS.n19144 DVSS.n19044 0.0640746
R44605 DVSS.n22376 DVSS.n22375 0.0640746
R44606 DVSS.n13017 DVSS.n13016 0.0638464
R44607 DVSS.n13060 DVSS.n13059 0.0638464
R44608 DVSS.n21466 DVSS.n21465 0.0618953
R44609 DVSS.n22964 DVSS.n22963 0.0618953
R44610 DVSS.n18515 DVSS.n18514 0.061538
R44611 DVSS.n18514 DVSS.n18513 0.060427
R44612 DVSS DVSS.n19891 0.059934
R44613 DVSS DVSS.n19886 0.059934
R44614 DVSS DVSS.n19048 0.059934
R44615 DVSS DVSS.n19878 0.059934
R44616 DVSS DVSS.n19873 0.059934
R44617 DVSS DVSS.n19056 0.059934
R44618 DVSS DVSS.n19865 0.059934
R44619 DVSS DVSS.n19860 0.059934
R44620 DVSS DVSS.n19064 0.059934
R44621 DVSS DVSS.n19584 0.059934
R44622 DVSS DVSS.n19579 0.059934
R44623 DVSS DVSS.n19524 0.059934
R44624 DVSS DVSS.n19571 0.059934
R44625 DVSS DVSS.n19566 0.059934
R44626 DVSS DVSS.n19532 0.059934
R44627 DVSS DVSS.n19558 0.059934
R44628 DVSS DVSS.n19553 0.059934
R44629 DVSS DVSS.n19540 0.059934
R44630 DVSS DVSS.n21832 0.059934
R44631 DVSS DVSS.n21840 0.059934
R44632 DVSS DVSS.n21826 0.059934
R44633 DVSS DVSS.n21847 0.059934
R44634 DVSS DVSS.n21948 0.059934
R44635 DVSS DVSS.n21937 0.059934
R44636 DVSS DVSS.n21915 0.059934
R44637 DVSS DVSS.n21905 0.059934
R44638 DVSS DVSS.n21895 0.059934
R44639 DVSS DVSS.n845 0.059934
R44640 DVSS DVSS.n836 0.059934
R44641 DVSS DVSS.n827 0.059934
R44642 DVSS DVSS.n818 0.059934
R44643 DVSS DVSS.n22480 0.059934
R44644 DVSS DVSS.n13044 0.059934
R44645 DVSS DVSS.n13032 0.059934
R44646 DVSS DVSS.n13053 0.059934
R44647 DVSS DVSS.n13018 0.059934
R44648 DVSS.n21464 DVSS.n21463 0.0574993
R44649 DVSS.n22962 DVSS.n22961 0.0574993
R44650 DVSS.n18663 DVSS.n18661 0.0568736
R44651 DVSS.n18661 DVSS.n18659 0.0568736
R44652 DVSS.n18659 DVSS.n18657 0.0568736
R44653 DVSS.n18773 DVSS.n18771 0.0568736
R44654 DVSS.n18775 DVSS.n18773 0.0568736
R44655 DVSS.n22583 DVSS.n752 0.056314
R44656 DVSS.n22938 DVSS.n434 0.056314
R44657 DVSS.n18992 DVSS.n18991 0.0562609
R44658 DVSS.n18991 DVSS.n18990 0.0562609
R44659 DVSS.n20686 DVSS.n14568 0.0562609
R44660 DVSS.n20676 DVSS.n14568 0.0562609
R44661 DVSS.n20676 DVSS.n20675 0.0562609
R44662 DVSS.n20671 DVSS.n14603 0.0562609
R44663 DVSS.n20661 DVSS.n14603 0.0562609
R44664 DVSS.n20661 DVSS.n20660 0.0562609
R44665 DVSS.n20660 DVSS.n20659 0.0562609
R44666 DVSS.n20659 DVSS.n14616 0.0562609
R44667 DVSS.n20645 DVSS.n14652 0.0562609
R44668 DVSS.n20634 DVSS.n14652 0.0562609
R44669 DVSS.n20634 DVSS.n20633 0.0562609
R44670 DVSS.n20620 DVSS.n20619 0.0562609
R44671 DVSS.n20619 DVSS.n20618 0.0562609
R44672 DVSS.n18767 DVSS.n18766 0.0562609
R44673 DVSS.n18766 DVSS.n18764 0.0562609
R44674 DVSS.n20105 DVSS.n14535 0.0562609
R44675 DVSS.n20106 DVSS.n20105 0.0562609
R44676 DVSS.n20107 DVSS.n20106 0.0562609
R44677 DVSS.n20177 DVSS.n20175 0.0562609
R44678 DVSS.n20178 DVSS.n20177 0.0562609
R44679 DVSS.n20180 DVSS.n20178 0.0562609
R44680 DVSS.n20181 DVSS.n20180 0.0562609
R44681 DVSS.n20183 DVSS.n20181 0.0562609
R44682 DVSS.n20320 DVSS.n20318 0.0562609
R44683 DVSS.n20321 DVSS.n20320 0.0562609
R44684 DVSS.n20323 DVSS.n20321 0.0562609
R44685 DVSS.n20462 DVSS.n20460 0.0562609
R44686 DVSS.n20463 DVSS.n20462 0.0562609
R44687 DVSS.n15533 DVSS.n15141 0.055378
R44688 DVSS.n19915 DVSS.n15137 0.055378
R44689 DVSS.n15920 DVSS.n15144 0.055378
R44690 DVSS.n18527 DVSS.n15145 0.055378
R44691 DVSS.n21462 DVSS.n21451 0.0551556
R44692 DVSS.n22960 DVSS.n22959 0.0551556
R44693 DVSS.n22630 DVSS.n22629 0.0549186
R44694 DVSS.n22891 DVSS.n450 0.0549186
R44695 DVSS.n1351 DVSS.n1350 0.0540178
R44696 DVSS.n1349 DVSS.n1348 0.0540178
R44697 DVSS.n1347 DVSS.n1346 0.0540178
R44698 DVSS.n1345 DVSS.n1344 0.0540178
R44699 DVSS.n1343 DVSS.n1342 0.0540178
R44700 DVSS.n1341 DVSS.n1340 0.0540178
R44701 DVSS.n1339 DVSS.n1338 0.0540178
R44702 DVSS.n1337 DVSS.n1336 0.0540178
R44703 DVSS.n1335 DVSS.n1334 0.0540178
R44704 DVSS.n1331 DVSS.n1330 0.0540178
R44705 DVSS.n1329 DVSS.n1328 0.0540178
R44706 DVSS.n1327 DVSS.n1326 0.0540178
R44707 DVSS.n1325 DVSS.n1324 0.0540178
R44708 DVSS.n1323 DVSS.n1322 0.0540178
R44709 DVSS.n1321 DVSS.n1320 0.0540178
R44710 DVSS.n1319 DVSS.n1318 0.0540178
R44711 DVSS.n1317 DVSS.n1316 0.0540178
R44712 DVSS.n1315 DVSS.n1314 0.0540178
R44713 DVSS.n1310 DVSS.n1309 0.0540178
R44714 DVSS.n1308 DVSS.n1307 0.0540178
R44715 DVSS.n1306 DVSS.n1305 0.0540178
R44716 DVSS.n1304 DVSS.n1303 0.0540178
R44717 DVSS.n1302 DVSS.n1301 0.0540178
R44718 DVSS.n1300 DVSS.n1299 0.0540178
R44719 DVSS.n1298 DVSS.n1297 0.0540178
R44720 DVSS.n1296 DVSS.n1295 0.0540178
R44721 DVSS.n1294 DVSS.n1293 0.0540178
R44722 DVSS.n1290 DVSS.n1289 0.0540178
R44723 DVSS.n1288 DVSS.n1287 0.0540178
R44724 DVSS.n1286 DVSS.n1285 0.0540178
R44725 DVSS.n1284 DVSS.n1283 0.0540178
R44726 DVSS.n1282 DVSS.n1281 0.0540178
R44727 DVSS.n1280 DVSS.n1279 0.0540178
R44728 DVSS.n1278 DVSS.n1277 0.0540178
R44729 DVSS.n1276 DVSS.n1275 0.0540178
R44730 DVSS.n1274 DVSS.n1273 0.0540178
R44731 DVSS.n878 DVSS.n866 0.0540178
R44732 DVSS.n877 DVSS.n865 0.0540178
R44733 DVSS.n876 DVSS.n864 0.0540178
R44734 DVSS.n875 DVSS.n863 0.0540178
R44735 DVSS.n874 DVSS.n862 0.0540178
R44736 DVSS.n873 DVSS.n861 0.0540178
R44737 DVSS.n872 DVSS.n860 0.0540178
R44738 DVSS.n871 DVSS.n859 0.0540178
R44739 DVSS.n21587 DVSS.n21575 0.0540178
R44740 DVSS.n21583 DVSS.n21574 0.0540178
R44741 DVSS.n21582 DVSS.n21573 0.0540178
R44742 DVSS.n21581 DVSS.n21572 0.0540178
R44743 DVSS.n21580 DVSS.n21571 0.0540178
R44744 DVSS.n21579 DVSS.n21570 0.0540178
R44745 DVSS.n21578 DVSS.n21569 0.0540178
R44746 DVSS.n1187 DVSS.n1177 0.0540178
R44747 DVSS.n1195 DVSS.n1186 0.0540178
R44748 DVSS.n1194 DVSS.n1185 0.0540178
R44749 DVSS.n1193 DVSS.n1184 0.0540178
R44750 DVSS.n1192 DVSS.n1183 0.0540178
R44751 DVSS.n1191 DVSS.n1182 0.0540178
R44752 DVSS.n1190 DVSS.n1181 0.0540178
R44753 DVSS.n1189 DVSS.n1180 0.0540178
R44754 DVSS.n1208 DVSS.n1198 0.0540178
R44755 DVSS.n1216 DVSS.n1207 0.0540178
R44756 DVSS.n1215 DVSS.n1206 0.0540178
R44757 DVSS.n1214 DVSS.n1205 0.0540178
R44758 DVSS.n1213 DVSS.n1204 0.0540178
R44759 DVSS.n1212 DVSS.n1203 0.0540178
R44760 DVSS.n1211 DVSS.n1202 0.0540178
R44761 DVSS.n1210 DVSS.n1201 0.0540178
R44762 DVSS.n21583 DVSS.n21575 0.0540178
R44763 DVSS.n21582 DVSS.n21574 0.0540178
R44764 DVSS.n21581 DVSS.n21573 0.0540178
R44765 DVSS.n21580 DVSS.n21572 0.0540178
R44766 DVSS.n21579 DVSS.n21571 0.0540178
R44767 DVSS.n21578 DVSS.n21570 0.0540178
R44768 DVSS.n1330 DVSS.n1329 0.0540178
R44769 DVSS.n1328 DVSS.n1327 0.0540178
R44770 DVSS.n1326 DVSS.n1325 0.0540178
R44771 DVSS.n1324 DVSS.n1323 0.0540178
R44772 DVSS.n1322 DVSS.n1321 0.0540178
R44773 DVSS.n1320 DVSS.n1319 0.0540178
R44774 DVSS.n1318 DVSS.n1317 0.0540178
R44775 DVSS.n1316 DVSS.n1315 0.0540178
R44776 DVSS.n1195 DVSS.n1187 0.0540178
R44777 DVSS.n1194 DVSS.n1186 0.0540178
R44778 DVSS.n1193 DVSS.n1185 0.0540178
R44779 DVSS.n1192 DVSS.n1184 0.0540178
R44780 DVSS.n1191 DVSS.n1183 0.0540178
R44781 DVSS.n1190 DVSS.n1182 0.0540178
R44782 DVSS.n1189 DVSS.n1181 0.0540178
R44783 DVSS.n1309 DVSS.n1308 0.0540178
R44784 DVSS.n1307 DVSS.n1306 0.0540178
R44785 DVSS.n1305 DVSS.n1304 0.0540178
R44786 DVSS.n1303 DVSS.n1302 0.0540178
R44787 DVSS.n1301 DVSS.n1300 0.0540178
R44788 DVSS.n1299 DVSS.n1298 0.0540178
R44789 DVSS.n1297 DVSS.n1296 0.0540178
R44790 DVSS.n1295 DVSS.n1294 0.0540178
R44791 DVSS.n878 DVSS.n865 0.0540178
R44792 DVSS.n877 DVSS.n864 0.0540178
R44793 DVSS.n876 DVSS.n863 0.0540178
R44794 DVSS.n875 DVSS.n862 0.0540178
R44795 DVSS.n874 DVSS.n861 0.0540178
R44796 DVSS.n873 DVSS.n860 0.0540178
R44797 DVSS.n872 DVSS.n859 0.0540178
R44798 DVSS.n1350 DVSS.n1349 0.0540178
R44799 DVSS.n1348 DVSS.n1347 0.0540178
R44800 DVSS.n1346 DVSS.n1345 0.0540178
R44801 DVSS.n1344 DVSS.n1343 0.0540178
R44802 DVSS.n1342 DVSS.n1341 0.0540178
R44803 DVSS.n1340 DVSS.n1339 0.0540178
R44804 DVSS.n1338 DVSS.n1337 0.0540178
R44805 DVSS.n1336 DVSS.n1335 0.0540178
R44806 DVSS.n19514 DVSS.n19278 0.0540178
R44807 DVSS.n19511 DVSS.n19277 0.0540178
R44808 DVSS.n19510 DVSS.n19276 0.0540178
R44809 DVSS.n19509 DVSS.n19275 0.0540178
R44810 DVSS.n19508 DVSS.n19274 0.0540178
R44811 DVSS.n19507 DVSS.n19273 0.0540178
R44812 DVSS.n19506 DVSS.n19272 0.0540178
R44813 DVSS.n19505 DVSS.n19271 0.0540178
R44814 DVSS.n19267 DVSS.n19266 0.0540178
R44815 DVSS.n19265 DVSS.n19264 0.0540178
R44816 DVSS.n19263 DVSS.n19262 0.0540178
R44817 DVSS.n19261 DVSS.n19260 0.0540178
R44818 DVSS.n19259 DVSS.n19258 0.0540178
R44819 DVSS.n19257 DVSS.n19256 0.0540178
R44820 DVSS.n19255 DVSS.n19254 0.0540178
R44821 DVSS.n19590 DVSS.n19253 0.0540178
R44822 DVSS.n19087 DVSS.n19077 0.0540178
R44823 DVSS.n19086 DVSS.n19076 0.0540178
R44824 DVSS.n19085 DVSS.n19075 0.0540178
R44825 DVSS.n19084 DVSS.n19074 0.0540178
R44826 DVSS.n19083 DVSS.n19073 0.0540178
R44827 DVSS.n19082 DVSS.n19072 0.0540178
R44828 DVSS.n19081 DVSS.n19071 0.0540178
R44829 DVSS.n19080 DVSS.n19070 0.0540178
R44830 DVSS.n19099 DVSS.n19090 0.0540178
R44831 DVSS.n19107 DVSS.n19098 0.0540178
R44832 DVSS.n19106 DVSS.n19097 0.0540178
R44833 DVSS.n19105 DVSS.n19096 0.0540178
R44834 DVSS.n19104 DVSS.n19095 0.0540178
R44835 DVSS.n19103 DVSS.n19094 0.0540178
R44836 DVSS.n19102 DVSS.n19093 0.0540178
R44837 DVSS.n19101 DVSS.n19092 0.0540178
R44838 DVSS.n19278 DVSS.n19277 0.0540178
R44839 DVSS.n19511 DVSS.n19276 0.0540178
R44840 DVSS.n19510 DVSS.n19275 0.0540178
R44841 DVSS.n19509 DVSS.n19274 0.0540178
R44842 DVSS.n19508 DVSS.n19273 0.0540178
R44843 DVSS.n19507 DVSS.n19272 0.0540178
R44844 DVSS.n19506 DVSS.n19271 0.0540178
R44845 DVSS.n19505 DVSS.n19270 0.0540178
R44846 DVSS.n19266 DVSS.n19265 0.0540178
R44847 DVSS.n19264 DVSS.n19263 0.0540178
R44848 DVSS.n19262 DVSS.n19261 0.0540178
R44849 DVSS.n19260 DVSS.n19259 0.0540178
R44850 DVSS.n19258 DVSS.n19257 0.0540178
R44851 DVSS.n19256 DVSS.n19255 0.0540178
R44852 DVSS.n19254 DVSS.n19253 0.0540178
R44853 DVSS.n19086 DVSS.n19077 0.0540178
R44854 DVSS.n19085 DVSS.n19076 0.0540178
R44855 DVSS.n19084 DVSS.n19075 0.0540178
R44856 DVSS.n19083 DVSS.n19074 0.0540178
R44857 DVSS.n19082 DVSS.n19073 0.0540178
R44858 DVSS.n19081 DVSS.n19072 0.0540178
R44859 DVSS.n19080 DVSS.n19071 0.0540178
R44860 DVSS.n1216 DVSS.n1208 0.0540178
R44861 DVSS.n1215 DVSS.n1207 0.0540178
R44862 DVSS.n1214 DVSS.n1206 0.0540178
R44863 DVSS.n1213 DVSS.n1205 0.0540178
R44864 DVSS.n1212 DVSS.n1204 0.0540178
R44865 DVSS.n1211 DVSS.n1203 0.0540178
R44866 DVSS.n1210 DVSS.n1202 0.0540178
R44867 DVSS.n1289 DVSS.n1288 0.0540178
R44868 DVSS.n1287 DVSS.n1286 0.0540178
R44869 DVSS.n1285 DVSS.n1284 0.0540178
R44870 DVSS.n1283 DVSS.n1282 0.0540178
R44871 DVSS.n1281 DVSS.n1280 0.0540178
R44872 DVSS.n1279 DVSS.n1278 0.0540178
R44873 DVSS.n1277 DVSS.n1276 0.0540178
R44874 DVSS.n1275 DVSS.n1274 0.0540178
R44875 DVSS.n19107 DVSS.n19099 0.0540178
R44876 DVSS.n19106 DVSS.n19098 0.0540178
R44877 DVSS.n19105 DVSS.n19097 0.0540178
R44878 DVSS.n19104 DVSS.n19096 0.0540178
R44879 DVSS.n19103 DVSS.n19095 0.0540178
R44880 DVSS.n19102 DVSS.n19094 0.0540178
R44881 DVSS.n19101 DVSS.n19093 0.0540178
R44882 DVSS.n14650 DVSS.n14649 0.0533261
R44883 DVSS.n20315 DVSS.n20194 0.0533261
R44884 DVSS.n868 DVSS.n867 0.0533261
R44885 DVSS.n22459 DVSS.n868 0.0533261
R44886 DVSS.n21588 DVSS.n21577 0.0533261
R44887 DVSS.n21585 DVSS.n21584 0.0533261
R44888 DVSS.n21584 DVSS.n1176 0.0533261
R44889 DVSS.n1196 DVSS.n1188 0.0533261
R44890 DVSS.n22338 DVSS.n1188 0.0533261
R44891 DVSS.n1217 DVSS.n1209 0.0533261
R44892 DVSS.n22335 DVSS.n1209 0.0533261
R44893 DVSS.n19504 DVSS.n19503 0.0533261
R44894 DVSS.n19591 DVSS.n19251 0.0533261
R44895 DVSS.n19593 DVSS.n19251 0.0533261
R44896 DVSS.n19088 DVSS.n19079 0.0533261
R44897 DVSS.n19849 DVSS.n19079 0.0533261
R44898 DVSS.n19108 DVSS.n19100 0.0533261
R44899 DVSS.n19846 DVSS.n19100 0.0533261
R44900 DVSS.n16222 DVSS.n15541 0.0528794
R44901 DVSS.n16427 DVSS.n15541 0.0528794
R44902 DVSS.n18506 DVSS.n13684 0.0521279
R44903 DVSS.n15133 DVSS.n15132 0.0521279
R44904 DVSS.n21006 DVSS.n21005 0.0521279
R44905 DVSS.n21158 DVSS.n21157 0.0507326
R44906 DVSS.n20987 DVSS.n14313 0.0507326
R44907 DVSS.n22971 DVSS.n422 0.0506031
R44908 DVSS.n22950 DVSS.n22949 0.0506031
R44909 DVSS.n22951 DVSS.n22950 0.0506031
R44910 DVSS.n22913 DVSS.n442 0.0506031
R44911 DVSS.n22916 DVSS.n442 0.0506031
R44912 DVSS.n21025 DVSS.n14309 0.0506031
R44913 DVSS.n21025 DVSS.n21024 0.0506031
R44914 DVSS.n22608 DVSS.n744 0.0506031
R44915 DVSS.n22605 DVSS.n744 0.0506031
R44916 DVSS.n22572 DVSS.n22571 0.0506031
R44917 DVSS.n22571 DVSS.n757 0.0506031
R44918 DVSS.n21473 DVSS.n1500 0.0506031
R44919 DVSS.n14559 DVSS.n14549 0.0503913
R44920 DVSS.n14562 DVSS.n14561 0.0503913
R44921 DVSS.n20674 DVSS.n14584 0.0503913
R44922 DVSS.n20123 DVSS.n14595 0.0503913
R44923 DVSS.n20310 DVSS.n14647 0.0503913
R44924 DVSS.n20646 DVSS.n14651 0.0503913
R44925 DVSS.n20430 DVSS.n20429 0.0503913
R44926 DVSS.n20356 DVSS.n20341 0.0503913
R44927 DVSS.n14538 DVSS.n14528 0.0503913
R44928 DVSS.n14540 DVSS.n14529 0.0503913
R44929 DVSS.n20110 DVSS.n20019 0.0503913
R44930 DVSS.n20112 DVSS.n20020 0.0503913
R44931 DVSS.n20195 DVSS.n20192 0.0503913
R44932 DVSS.n20317 DVSS.n14863 0.0503913
R44933 DVSS.n20363 DVSS.n20330 0.0503913
R44934 DVSS.n20350 DVSS.n20331 0.0503913
R44935 DVSS.n21172 DVSS.n21171 0.0503
R44936 DVSS.n19249 DVSS.n19215 0.0495829
R44937 DVSS.n19623 DVSS.n19160 0.0495829
R44938 DVSS.n19902 DVSS.n19901 0.0495829
R44939 DVSS.n19651 DVSS.n19147 0.0495829
R44940 DVSS.n20987 DVSS.n20986 0.0495306
R44941 DVSS.n20985 DVSS.n14314 0.0490001
R44942 DVSS.n21439 DVSS.n13371 0.0490001
R44943 DVSS.n22636 DVSS.n22635 0.0489295
R44944 DVSS.n453 DVSS.n452 0.0489295
R44945 DVSS.n18777 DVSS.n18775 0.0479692
R44946 DVSS.n21459 DVSS.n21458 0.0479419
R44947 DVSS.n22588 DVSS.n751 0.0479419
R44948 DVSS.n22933 DVSS.n435 0.0479419
R44949 DVSS.n22957 DVSS.n428 0.0479419
R44950 DVSS.n18903 DVSS.n14555 0.0474565
R44951 DVSS.n18943 DVSS.n14554 0.0474565
R44952 DVSS.n20125 DVSS.n14591 0.0474565
R44953 DVSS.n20672 DVSS.n20671 0.0474565
R44954 DVSS.n14630 DVSS.n14616 0.0474565
R44955 DVSS.n20202 DVSS.n14635 0.0474565
R44956 DVSS.n20428 DVSS.n20359 0.0474565
R44957 DVSS.n20446 DVSS.n20445 0.0474565
R44958 DVSS.n18888 DVSS.n14524 0.0474565
R44959 DVSS.n18947 DVSS.n14521 0.0474565
R44960 DVSS.n20098 DVSS.n20016 0.0474565
R44961 DVSS.n20175 DVSS.n20174 0.0474565
R44962 DVSS.n20185 DVSS.n20183 0.0474565
R44963 DVSS.n20204 DVSS.n14867 0.0474565
R44964 DVSS.n20365 DVSS.n14858 0.0474565
R44965 DVSS.n20344 DVSS.n14855 0.0474565
R44966 DVSS.n22231 DVSS.n1312 0.0457174
R44967 DVSS.n22342 DVSS.n22341 0.0457174
R44968 DVSS.n19595 DVSS.n19594 0.0457174
R44969 DVSS.n21174 DVSS.n21173 0.0455
R44970 DVSS.n17048 DVSS.n17047 0.0450718
R44971 DVSS.n17046 DVSS.n17045 0.0450718
R44972 DVSS.n17044 DVSS.n17043 0.0450718
R44973 DVSS.n17042 DVSS.n17041 0.0450718
R44974 DVSS.n17040 DVSS.n17039 0.0450718
R44975 DVSS.n17038 DVSS.n17037 0.0450718
R44976 DVSS.n17034 DVSS.n17033 0.0450718
R44977 DVSS.n17032 DVSS.n17031 0.0450718
R44978 DVSS.n17030 DVSS.n17029 0.0450718
R44979 DVSS.n17028 DVSS.n17027 0.0450718
R44980 DVSS.n17026 DVSS.n17025 0.0450718
R44981 DVSS.n17024 DVSS.n17023 0.0450718
R44982 DVSS.n17022 DVSS.n17021 0.0450718
R44983 DVSS.n17020 DVSS.n17019 0.0450718
R44984 DVSS.n17018 DVSS.n17017 0.0450718
R44985 DVSS.n17013 DVSS.n17012 0.0450718
R44986 DVSS.n17011 DVSS.n17010 0.0450718
R44987 DVSS.n17009 DVSS.n17008 0.0450718
R44988 DVSS.n17007 DVSS.n17006 0.0450718
R44989 DVSS.n17005 DVSS.n17004 0.0450718
R44990 DVSS.n17003 DVSS.n17002 0.0450718
R44991 DVSS.n17001 DVSS.n17000 0.0450718
R44992 DVSS.n16999 DVSS.n16998 0.0450718
R44993 DVSS.n16997 DVSS.n16996 0.0450718
R44994 DVSS.n16993 DVSS.n16992 0.0450718
R44995 DVSS.n16991 DVSS.n16990 0.0450718
R44996 DVSS.n16989 DVSS.n16988 0.0450718
R44997 DVSS.n16987 DVSS.n16986 0.0450718
R44998 DVSS.n16985 DVSS.n16984 0.0450718
R44999 DVSS.n16983 DVSS.n16982 0.0450718
R45000 DVSS.n17113 DVSS.n17112 0.0450718
R45001 DVSS.n17112 DVSS.n17111 0.0450718
R45002 DVSS.n17111 DVSS.n17110 0.0450718
R45003 DVSS.n17110 DVSS.n17109 0.0450718
R45004 DVSS.n17109 DVSS.n17108 0.0450718
R45005 DVSS.n17108 DVSS.n17107 0.0450718
R45006 DVSS.n17107 DVSS.n17106 0.0450718
R45007 DVSS.n17106 DVSS.n17105 0.0450718
R45008 DVSS.n17105 DVSS.n17104 0.0450718
R45009 DVSS.n17104 DVSS.n17103 0.0450718
R45010 DVSS.n17103 DVSS.n17102 0.0450718
R45011 DVSS.n17073 DVSS.n17065 0.0450718
R45012 DVSS.n17073 DVSS.n17064 0.0450718
R45013 DVSS.n17072 DVSS.n17064 0.0450718
R45014 DVSS.n17072 DVSS.n17063 0.0450718
R45015 DVSS.n17071 DVSS.n17063 0.0450718
R45016 DVSS.n17071 DVSS.n17062 0.0450718
R45017 DVSS.n17070 DVSS.n17062 0.0450718
R45018 DVSS.n17070 DVSS.n17061 0.0450718
R45019 DVSS.n17069 DVSS.n17061 0.0450718
R45020 DVSS.n17069 DVSS.n17060 0.0450718
R45021 DVSS.n17068 DVSS.n17060 0.0450718
R45022 DVSS.n17068 DVSS.n17059 0.0450718
R45023 DVSS.n17067 DVSS.n17059 0.0450718
R45024 DVSS.n17067 DVSS.n17058 0.0450718
R45025 DVSS.n17076 DVSS.n17058 0.0450718
R45026 DVSS.n17095 DVSS.n17094 0.0450718
R45027 DVSS.n17094 DVSS.n17093 0.0450718
R45028 DVSS.n17093 DVSS.n17092 0.0450718
R45029 DVSS.n17092 DVSS.n17091 0.0450718
R45030 DVSS.n17091 DVSS.n17090 0.0450718
R45031 DVSS.n17090 DVSS.n17089 0.0450718
R45032 DVSS.n17089 DVSS.n17088 0.0450718
R45033 DVSS.n17088 DVSS.n17087 0.0450718
R45034 DVSS.n17087 DVSS.n17086 0.0450718
R45035 DVSS.n17086 DVSS.n17085 0.0450718
R45036 DVSS.n17085 DVSS.n17084 0.0450718
R45037 DVSS.n17084 DVSS.n17083 0.0450718
R45038 DVSS.n17083 DVSS.n17082 0.0450718
R45039 DVSS.n17082 DVSS.n17081 0.0450718
R45040 DVSS.n17081 DVSS.n17080 0.0450718
R45041 DVSS.n17080 DVSS.n17079 0.0450718
R45042 DVSS.n17079 DVSS.n17078 0.0450718
R45043 DVSS.n16911 DVSS.n16910 0.0450718
R45044 DVSS.n16912 DVSS.n16911 0.0450718
R45045 DVSS.n16913 DVSS.n16912 0.0450718
R45046 DVSS.n16914 DVSS.n16913 0.0450718
R45047 DVSS.n16915 DVSS.n16914 0.0450718
R45048 DVSS.n16916 DVSS.n16915 0.0450718
R45049 DVSS.n16917 DVSS.n16916 0.0450718
R45050 DVSS.n16918 DVSS.n16917 0.0450718
R45051 DVSS.n16919 DVSS.n16918 0.0450718
R45052 DVSS.n16921 DVSS.n16919 0.0450718
R45053 DVSS.n16923 DVSS.n16921 0.0450718
R45054 DVSS.n16923 DVSS.n16922 0.0450718
R45055 DVSS.n17019 DVSS.n17018 0.0450718
R45056 DVSS.n17021 DVSS.n17020 0.0450718
R45057 DVSS.n17023 DVSS.n17022 0.0450718
R45058 DVSS.n17025 DVSS.n17024 0.0450718
R45059 DVSS.n17027 DVSS.n17026 0.0450718
R45060 DVSS.n17029 DVSS.n17028 0.0450718
R45061 DVSS.n17031 DVSS.n17030 0.0450718
R45062 DVSS.n17033 DVSS.n17032 0.0450718
R45063 DVSS.n16998 DVSS.n16997 0.0450718
R45064 DVSS.n17000 DVSS.n16999 0.0450718
R45065 DVSS.n17002 DVSS.n17001 0.0450718
R45066 DVSS.n17004 DVSS.n17003 0.0450718
R45067 DVSS.n17006 DVSS.n17005 0.0450718
R45068 DVSS.n17008 DVSS.n17007 0.0450718
R45069 DVSS.n17010 DVSS.n17009 0.0450718
R45070 DVSS.n17012 DVSS.n17011 0.0450718
R45071 DVSS.n17114 DVSS.n17113 0.0450718
R45072 DVSS.n17039 DVSS.n17038 0.0450718
R45073 DVSS.n17041 DVSS.n17040 0.0450718
R45074 DVSS.n17043 DVSS.n17042 0.0450718
R45075 DVSS.n17045 DVSS.n17044 0.0450718
R45076 DVSS.n17047 DVSS.n17046 0.0450718
R45077 DVSS.n17049 DVSS.n17048 0.0450718
R45078 DVSS.n16982 DVSS.n16981 0.0450718
R45079 DVSS.n16984 DVSS.n16983 0.0450718
R45080 DVSS.n16986 DVSS.n16985 0.0450718
R45081 DVSS.n16988 DVSS.n16987 0.0450718
R45082 DVSS.n16990 DVSS.n16989 0.0450718
R45083 DVSS.n16992 DVSS.n16991 0.0450718
R45084 DVSS.n18901 DVSS.n14558 0.0445217
R45085 DVSS.n18945 DVSS.n14563 0.0445217
R45086 DVSS.n20084 DVSS.n14596 0.0445217
R45087 DVSS.n20166 DVSS.n14602 0.0445217
R45088 DVSS.n20649 DVSS.n20648 0.0445217
R45089 DVSS.n20200 DVSS.n14646 0.0445217
R45090 DVSS.n20417 DVSS.n20416 0.0445217
R45091 DVSS.n20448 DVSS.n20447 0.0445217
R45092 DVSS.n18893 DVSS.n14527 0.0445217
R45093 DVSS.n18951 DVSS.n14530 0.0445217
R45094 DVSS.n20096 DVSS.n20021 0.0445217
R45095 DVSS.n20027 DVSS.n14874 0.0445217
R45096 DVSS.n20184 DVSS.n14873 0.0445217
R45097 DVSS.n20231 DVSS.n20191 0.0445217
R45098 DVSS.n20371 DVSS.n20329 0.0445217
R45099 DVSS.n20457 DVSS.n20332 0.0445217
R45100 DVSS.n17074 DVSS.n17066 0.0442838
R45101 DVSS.n21170 DVSS.n13668 0.04343
R45102 DVSS.n21169 DVSS.n21168 0.04343
R45103 DVSS.n13670 DVSS.n13669 0.04343
R45104 DVSS.n18512 DVSS.n18511 0.04343
R45105 DVSS.n18499 DVSS.n18498 0.04343
R45106 DVSS.n18665 DVSS.n18663 0.0424895
R45107 DVSS.n13679 DVSS.n13675 0.0423605
R45108 DVSS.n21015 DVSS.n20997 0.0423605
R45109 DVSS.n1501 DVSS.n1000 0.0422789
R45110 DVSS.n13101 DVSS.n13100 0.0422789
R45111 DVSS.n18890 DVSS.n14556 0.041587
R45112 DVSS.n18961 DVSS.n14553 0.041587
R45113 DVSS.n20086 DVSS.n14590 0.041587
R45114 DVSS.n20167 DVSS.n14601 0.041587
R45115 DVSS.n14641 DVSS.n14632 0.041587
R45116 DVSS.n20292 DVSS.n14636 0.041587
R45117 DVSS.n20418 DVSS.n20415 0.041587
R45118 DVSS.n20452 DVSS.n20451 0.041587
R45119 DVSS.n18895 DVSS.n14525 0.041587
R45120 DVSS.n18949 DVSS.n14520 0.041587
R45121 DVSS.n20090 DVSS.n20015 0.041587
R45122 DVSS.n20172 DVSS.n20171 0.041587
R45123 DVSS.n20262 DVSS.n20186 0.041587
R45124 DVSS.n20233 DVSS.n14868 0.041587
R45125 DVSS.n20373 DVSS.n14859 0.041587
R45126 DVSS.n20456 DVSS.n20333 0.041587
R45127 DVSS.n21164 DVSS.n13673 0.04037
R45128 DVSS.n21163 DVSS.n21162 0.04037
R45129 DVSS.n21156 DVSS.n13674 0.04037
R45130 DVSS.n18503 DVSS.n13685 0.04037
R45131 DVSS.n18509 DVSS.n18504 0.04037
R45132 DVSS.n21014 DVSS.n21013 0.040062
R45133 DVSS DVSS.n14577 0.039875
R45134 DVSS DVSS.n14578 0.039875
R45135 DVSS DVSS.n14621 0.039875
R45136 DVSS DVSS.n14622 0.039875
R45137 DVSS DVSS.n14661 0.039875
R45138 DVSS DVSS.n14662 0.039875
R45139 DVSS DVSS.n15540 0.039875
R45140 DVSS.n22606 DVSS.n745 0.0395698
R45141 DVSS.n22915 DVSS.n441 0.0395698
R45142 DVSS.n18657 DVSS.n18655 0.0395659
R45143 DVSS.n18771 DVSS.n18769 0.0395659
R45144 DVSS.n1503 DVSS.n1136 0.0392219
R45145 DVSS.n13006 DVSS.n1504 0.0392219
R45146 DVSS.n1502 DVSS.n1082 0.0392219
R45147 DVSS.n13364 DVSS.n349 0.0392219
R45148 DVSS.n18504 DVSS.n18503 0.0389615
R45149 DVSS.n18503 DVSS.n13674 0.0389615
R45150 DVSS.n21164 DVSS.n13670 0.0389615
R45151 DVSS.n21465 DVSS.n21464 0.0389615
R45152 DVSS.n21458 DVSS.n21451 0.0389615
R45153 DVSS.n22581 DVSS.n752 0.0389615
R45154 DVSS.n22590 DVSS.n751 0.0389615
R45155 DVSS.n745 DVSS.n743 0.0389615
R45156 DVSS.n22623 DVSS.n737 0.0389615
R45157 DVSS.n22629 DVSS.n735 0.0389615
R45158 DVSS.n21173 DVSS.n13668 0.0389615
R45159 DVSS.n21168 DVSS.n13670 0.0389615
R45160 DVSS.n21168 DVSS.n13668 0.0389615
R45161 DVSS.n21163 DVSS.n13674 0.0389615
R45162 DVSS.n21164 DVSS.n21163 0.0389615
R45163 DVSS.n18512 DVSS.n18499 0.0389615
R45164 DVSS.n18512 DVSS.n18504 0.0389615
R45165 DVSS.n15132 DVSS.n15126 0.0389615
R45166 DVSS.n20988 DVSS.n20987 0.0389615
R45167 DVSS.n21015 DVSS.n21014 0.0389615
R45168 DVSS.n21005 DVSS.n20999 0.0389615
R45169 DVSS.n22889 DVSS.n450 0.0389615
R45170 DVSS.n22898 DVSS.n449 0.0389615
R45171 DVSS.n443 DVSS.n441 0.0389615
R45172 DVSS.n22931 DVSS.n435 0.0389615
R45173 DVSS.n22940 DVSS.n434 0.0389615
R45174 DVSS.n22959 DVSS.n428 0.0389615
R45175 DVSS.n22963 DVSS.n22962 0.0389615
R45176 DVSS.n18648 DVSS.n14557 0.0386522
R45177 DVSS.n18963 DVSS.n14564 0.0386522
R45178 DVSS.n20135 DVSS.n14597 0.0386522
R45179 DVSS.n20164 DVSS.n14586 0.0386522
R45180 DVSS.n20268 DVSS.n14640 0.0386522
R45181 DVSS.n20294 DVSS.n14645 0.0386522
R45182 DVSS.n20414 DVSS.n20413 0.0386522
R45183 DVSS.n20449 DVSS.n14702 0.0386522
R45184 DVSS.n18891 DVSS.n14526 0.0386522
R45185 DVSS.n18941 DVSS.n14531 0.0386522
R45186 DVSS.n20088 DVSS.n20022 0.0386522
R45187 DVSS.n20026 DVSS.n20011 0.0386522
R45188 DVSS.n20266 DVSS.n14872 0.0386522
R45189 DVSS.n20235 DVSS.n20190 0.0386522
R45190 DVSS.n20379 DVSS.n20328 0.0386522
R45191 DVSS.n20459 DVSS.n14852 0.0386522
R45192 DVSS.n11734 DVSS.n11624 0.0380882
R45193 DVSS.n11735 DVSS.n11734 0.0380882
R45194 DVSS.n11735 DVSS.n11729 0.0380882
R45195 DVSS.n11745 DVSS.n11729 0.0380882
R45196 DVSS.n11746 DVSS.n11745 0.0380882
R45197 DVSS.n11747 DVSS.n11746 0.0380882
R45198 DVSS.n11747 DVSS.n11727 0.0380882
R45199 DVSS.n11757 DVSS.n11727 0.0380882
R45200 DVSS.n11758 DVSS.n11757 0.0380882
R45201 DVSS.n11759 DVSS.n11758 0.0380882
R45202 DVSS.n11759 DVSS.n11725 0.0380882
R45203 DVSS.n11769 DVSS.n11725 0.0380882
R45204 DVSS.n11770 DVSS.n11769 0.0380882
R45205 DVSS.n11771 DVSS.n11770 0.0380882
R45206 DVSS.n11771 DVSS.n11723 0.0380882
R45207 DVSS.n11781 DVSS.n11723 0.0380882
R45208 DVSS.n11782 DVSS.n11781 0.0380882
R45209 DVSS.n11783 DVSS.n11782 0.0380882
R45210 DVSS.n11783 DVSS.n11721 0.0380882
R45211 DVSS.n11793 DVSS.n11721 0.0380882
R45212 DVSS.n11794 DVSS.n11793 0.0380882
R45213 DVSS.n11795 DVSS.n11794 0.0380882
R45214 DVSS.n11795 DVSS.n11719 0.0380882
R45215 DVSS.n11805 DVSS.n11719 0.0380882
R45216 DVSS.n11806 DVSS.n11805 0.0380882
R45217 DVSS.n11807 DVSS.n11806 0.0380882
R45218 DVSS.n11807 DVSS.n11717 0.0380882
R45219 DVSS.n11817 DVSS.n11717 0.0380882
R45220 DVSS.n11818 DVSS.n11817 0.0380882
R45221 DVSS.n11819 DVSS.n11818 0.0380882
R45222 DVSS.n11819 DVSS.n11715 0.0380882
R45223 DVSS.n11829 DVSS.n11715 0.0380882
R45224 DVSS.n11830 DVSS.n11829 0.0380882
R45225 DVSS.n11831 DVSS.n11830 0.0380882
R45226 DVSS.n11831 DVSS.n11713 0.0380882
R45227 DVSS.n11841 DVSS.n11713 0.0380882
R45228 DVSS.n11842 DVSS.n11841 0.0380882
R45229 DVSS.n11843 DVSS.n11842 0.0380882
R45230 DVSS.n11843 DVSS.n11711 0.0380882
R45231 DVSS.n11853 DVSS.n11711 0.0380882
R45232 DVSS.n11854 DVSS.n11853 0.0380882
R45233 DVSS.n11855 DVSS.n11854 0.0380882
R45234 DVSS.n11855 DVSS.n11709 0.0380882
R45235 DVSS.n11865 DVSS.n11709 0.0380882
R45236 DVSS.n11866 DVSS.n11865 0.0380882
R45237 DVSS.n11867 DVSS.n11866 0.0380882
R45238 DVSS.n11867 DVSS.n11707 0.0380882
R45239 DVSS.n11877 DVSS.n11707 0.0380882
R45240 DVSS.n11878 DVSS.n11877 0.0380882
R45241 DVSS.n11879 DVSS.n11878 0.0380882
R45242 DVSS.n11879 DVSS.n11705 0.0380882
R45243 DVSS.n11889 DVSS.n11705 0.0380882
R45244 DVSS.n11890 DVSS.n11889 0.0380882
R45245 DVSS.n11891 DVSS.n11890 0.0380882
R45246 DVSS.n11891 DVSS.n11703 0.0380882
R45247 DVSS.n11901 DVSS.n11703 0.0380882
R45248 DVSS.n11902 DVSS.n11901 0.0380882
R45249 DVSS.n11903 DVSS.n11902 0.0380882
R45250 DVSS.n11903 DVSS.n11701 0.0380882
R45251 DVSS.n11913 DVSS.n11701 0.0380882
R45252 DVSS.n11914 DVSS.n11913 0.0380882
R45253 DVSS.n11915 DVSS.n11914 0.0380882
R45254 DVSS.n11915 DVSS.n11699 0.0380882
R45255 DVSS.n11925 DVSS.n11699 0.0380882
R45256 DVSS.n11926 DVSS.n11925 0.0380882
R45257 DVSS.n11927 DVSS.n11926 0.0380882
R45258 DVSS.n11927 DVSS.n11697 0.0380882
R45259 DVSS.n11937 DVSS.n11697 0.0380882
R45260 DVSS.n11938 DVSS.n11937 0.0380882
R45261 DVSS.n11939 DVSS.n11938 0.0380882
R45262 DVSS.n11939 DVSS.n11695 0.0380882
R45263 DVSS.n11949 DVSS.n11695 0.0380882
R45264 DVSS.n11950 DVSS.n11949 0.0380882
R45265 DVSS.n11951 DVSS.n11950 0.0380882
R45266 DVSS.n11951 DVSS.n11693 0.0380882
R45267 DVSS.n11961 DVSS.n11693 0.0380882
R45268 DVSS.n11962 DVSS.n11961 0.0380882
R45269 DVSS.n11963 DVSS.n11962 0.0380882
R45270 DVSS.n11963 DVSS.n11691 0.0380882
R45271 DVSS.n11973 DVSS.n11691 0.0380882
R45272 DVSS.n11974 DVSS.n11973 0.0380882
R45273 DVSS.n11975 DVSS.n11974 0.0380882
R45274 DVSS.n11975 DVSS.n11636 0.0380882
R45275 DVSS.n5623 DVSS.n5622 0.0380882
R45276 DVSS.n5624 DVSS.n5623 0.0380882
R45277 DVSS.n5624 DVSS.n5617 0.0380882
R45278 DVSS.n5634 DVSS.n5617 0.0380882
R45279 DVSS.n5635 DVSS.n5634 0.0380882
R45280 DVSS.n5636 DVSS.n5635 0.0380882
R45281 DVSS.n5636 DVSS.n5615 0.0380882
R45282 DVSS.n5646 DVSS.n5615 0.0380882
R45283 DVSS.n5647 DVSS.n5646 0.0380882
R45284 DVSS.n5648 DVSS.n5647 0.0380882
R45285 DVSS.n5648 DVSS.n5613 0.0380882
R45286 DVSS.n5658 DVSS.n5613 0.0380882
R45287 DVSS.n5659 DVSS.n5658 0.0380882
R45288 DVSS.n5660 DVSS.n5659 0.0380882
R45289 DVSS.n5660 DVSS.n5611 0.0380882
R45290 DVSS.n5670 DVSS.n5611 0.0380882
R45291 DVSS.n5671 DVSS.n5670 0.0380882
R45292 DVSS.n5672 DVSS.n5671 0.0380882
R45293 DVSS.n5672 DVSS.n5609 0.0380882
R45294 DVSS.n5682 DVSS.n5609 0.0380882
R45295 DVSS.n5683 DVSS.n5682 0.0380882
R45296 DVSS.n5684 DVSS.n5683 0.0380882
R45297 DVSS.n5684 DVSS.n5607 0.0380882
R45298 DVSS.n5694 DVSS.n5607 0.0380882
R45299 DVSS.n5695 DVSS.n5694 0.0380882
R45300 DVSS.n5696 DVSS.n5695 0.0380882
R45301 DVSS.n5696 DVSS.n5605 0.0380882
R45302 DVSS.n5706 DVSS.n5605 0.0380882
R45303 DVSS.n5707 DVSS.n5706 0.0380882
R45304 DVSS.n5708 DVSS.n5707 0.0380882
R45305 DVSS.n5708 DVSS.n5603 0.0380882
R45306 DVSS.n5718 DVSS.n5603 0.0380882
R45307 DVSS.n5719 DVSS.n5718 0.0380882
R45308 DVSS.n5720 DVSS.n5719 0.0380882
R45309 DVSS.n5720 DVSS.n5601 0.0380882
R45310 DVSS.n5730 DVSS.n5601 0.0380882
R45311 DVSS.n5731 DVSS.n5730 0.0380882
R45312 DVSS.n5732 DVSS.n5731 0.0380882
R45313 DVSS.n5732 DVSS.n5599 0.0380882
R45314 DVSS.n5742 DVSS.n5599 0.0380882
R45315 DVSS.n5743 DVSS.n5742 0.0380882
R45316 DVSS.n5744 DVSS.n5743 0.0380882
R45317 DVSS.n5744 DVSS.n5597 0.0380882
R45318 DVSS.n5754 DVSS.n5597 0.0380882
R45319 DVSS.n5755 DVSS.n5754 0.0380882
R45320 DVSS.n5756 DVSS.n5755 0.0380882
R45321 DVSS.n5756 DVSS.n5595 0.0380882
R45322 DVSS.n5766 DVSS.n5595 0.0380882
R45323 DVSS.n5767 DVSS.n5766 0.0380882
R45324 DVSS.n5768 DVSS.n5767 0.0380882
R45325 DVSS.n5768 DVSS.n5593 0.0380882
R45326 DVSS.n5778 DVSS.n5593 0.0380882
R45327 DVSS.n5779 DVSS.n5778 0.0380882
R45328 DVSS.n5780 DVSS.n5779 0.0380882
R45329 DVSS.n5780 DVSS.n5591 0.0380882
R45330 DVSS.n5790 DVSS.n5591 0.0380882
R45331 DVSS.n5791 DVSS.n5790 0.0380882
R45332 DVSS.n5792 DVSS.n5791 0.0380882
R45333 DVSS.n5792 DVSS.n5589 0.0380882
R45334 DVSS.n5802 DVSS.n5589 0.0380882
R45335 DVSS.n5803 DVSS.n5802 0.0380882
R45336 DVSS.n5804 DVSS.n5803 0.0380882
R45337 DVSS.n5804 DVSS.n5587 0.0380882
R45338 DVSS.n5814 DVSS.n5587 0.0380882
R45339 DVSS.n5815 DVSS.n5814 0.0380882
R45340 DVSS.n5816 DVSS.n5815 0.0380882
R45341 DVSS.n5816 DVSS.n5585 0.0380882
R45342 DVSS.n5826 DVSS.n5585 0.0380882
R45343 DVSS.n5827 DVSS.n5826 0.0380882
R45344 DVSS.n5828 DVSS.n5827 0.0380882
R45345 DVSS.n5828 DVSS.n5583 0.0380882
R45346 DVSS.n5838 DVSS.n5583 0.0380882
R45347 DVSS.n5839 DVSS.n5838 0.0380882
R45348 DVSS.n5840 DVSS.n5839 0.0380882
R45349 DVSS.n5840 DVSS.n5581 0.0380882
R45350 DVSS.n5850 DVSS.n5581 0.0380882
R45351 DVSS.n5851 DVSS.n5850 0.0380882
R45352 DVSS.n5852 DVSS.n5851 0.0380882
R45353 DVSS.n5852 DVSS.n5579 0.0380882
R45354 DVSS.n5862 DVSS.n5579 0.0380882
R45355 DVSS.n5863 DVSS.n5862 0.0380882
R45356 DVSS.n7054 DVSS.n5863 0.0380882
R45357 DVSS.n7054 DVSS.n7053 0.0380882
R45358 DVSS.n5621 DVSS.n5620 0.0380882
R45359 DVSS.n5625 DVSS.n5620 0.0380882
R45360 DVSS.n5629 DVSS.n5625 0.0380882
R45361 DVSS.n5633 DVSS.n5629 0.0380882
R45362 DVSS.n5633 DVSS.n5616 0.0380882
R45363 DVSS.n5637 DVSS.n5616 0.0380882
R45364 DVSS.n5641 DVSS.n5637 0.0380882
R45365 DVSS.n5645 DVSS.n5641 0.0380882
R45366 DVSS.n5645 DVSS.n5614 0.0380882
R45367 DVSS.n5649 DVSS.n5614 0.0380882
R45368 DVSS.n5653 DVSS.n5649 0.0380882
R45369 DVSS.n5657 DVSS.n5653 0.0380882
R45370 DVSS.n5657 DVSS.n5612 0.0380882
R45371 DVSS.n5661 DVSS.n5612 0.0380882
R45372 DVSS.n5665 DVSS.n5661 0.0380882
R45373 DVSS.n5669 DVSS.n5665 0.0380882
R45374 DVSS.n5669 DVSS.n5610 0.0380882
R45375 DVSS.n5673 DVSS.n5610 0.0380882
R45376 DVSS.n5677 DVSS.n5673 0.0380882
R45377 DVSS.n5681 DVSS.n5677 0.0380882
R45378 DVSS.n5681 DVSS.n5608 0.0380882
R45379 DVSS.n5685 DVSS.n5608 0.0380882
R45380 DVSS.n5689 DVSS.n5685 0.0380882
R45381 DVSS.n5693 DVSS.n5689 0.0380882
R45382 DVSS.n5693 DVSS.n5606 0.0380882
R45383 DVSS.n5697 DVSS.n5606 0.0380882
R45384 DVSS.n5701 DVSS.n5697 0.0380882
R45385 DVSS.n5705 DVSS.n5701 0.0380882
R45386 DVSS.n5705 DVSS.n5604 0.0380882
R45387 DVSS.n5709 DVSS.n5604 0.0380882
R45388 DVSS.n5713 DVSS.n5709 0.0380882
R45389 DVSS.n5717 DVSS.n5713 0.0380882
R45390 DVSS.n5717 DVSS.n5602 0.0380882
R45391 DVSS.n5721 DVSS.n5602 0.0380882
R45392 DVSS.n5725 DVSS.n5721 0.0380882
R45393 DVSS.n5729 DVSS.n5725 0.0380882
R45394 DVSS.n5729 DVSS.n5600 0.0380882
R45395 DVSS.n5733 DVSS.n5600 0.0380882
R45396 DVSS.n5737 DVSS.n5733 0.0380882
R45397 DVSS.n5741 DVSS.n5737 0.0380882
R45398 DVSS.n5741 DVSS.n5598 0.0380882
R45399 DVSS.n5745 DVSS.n5598 0.0380882
R45400 DVSS.n5749 DVSS.n5745 0.0380882
R45401 DVSS.n5753 DVSS.n5749 0.0380882
R45402 DVSS.n5753 DVSS.n5596 0.0380882
R45403 DVSS.n5757 DVSS.n5596 0.0380882
R45404 DVSS.n5761 DVSS.n5757 0.0380882
R45405 DVSS.n5765 DVSS.n5761 0.0380882
R45406 DVSS.n5765 DVSS.n5594 0.0380882
R45407 DVSS.n5769 DVSS.n5594 0.0380882
R45408 DVSS.n5773 DVSS.n5769 0.0380882
R45409 DVSS.n5777 DVSS.n5773 0.0380882
R45410 DVSS.n5777 DVSS.n5592 0.0380882
R45411 DVSS.n5781 DVSS.n5592 0.0380882
R45412 DVSS.n5785 DVSS.n5781 0.0380882
R45413 DVSS.n5789 DVSS.n5785 0.0380882
R45414 DVSS.n5789 DVSS.n5590 0.0380882
R45415 DVSS.n5793 DVSS.n5590 0.0380882
R45416 DVSS.n5797 DVSS.n5793 0.0380882
R45417 DVSS.n5801 DVSS.n5797 0.0380882
R45418 DVSS.n5801 DVSS.n5588 0.0380882
R45419 DVSS.n5805 DVSS.n5588 0.0380882
R45420 DVSS.n5809 DVSS.n5805 0.0380882
R45421 DVSS.n5813 DVSS.n5809 0.0380882
R45422 DVSS.n5813 DVSS.n5586 0.0380882
R45423 DVSS.n5817 DVSS.n5586 0.0380882
R45424 DVSS.n5821 DVSS.n5817 0.0380882
R45425 DVSS.n5825 DVSS.n5821 0.0380882
R45426 DVSS.n5825 DVSS.n5584 0.0380882
R45427 DVSS.n5829 DVSS.n5584 0.0380882
R45428 DVSS.n5833 DVSS.n5829 0.0380882
R45429 DVSS.n5837 DVSS.n5833 0.0380882
R45430 DVSS.n5837 DVSS.n5582 0.0380882
R45431 DVSS.n5841 DVSS.n5582 0.0380882
R45432 DVSS.n5845 DVSS.n5841 0.0380882
R45433 DVSS.n5849 DVSS.n5845 0.0380882
R45434 DVSS.n5849 DVSS.n5580 0.0380882
R45435 DVSS.n5853 DVSS.n5580 0.0380882
R45436 DVSS.n5857 DVSS.n5853 0.0380882
R45437 DVSS.n5861 DVSS.n5857 0.0380882
R45438 DVSS.n5861 DVSS.n5578 0.0380882
R45439 DVSS.n7055 DVSS.n5578 0.0380882
R45440 DVSS.n7055 DVSS.n5576 0.0380882
R45441 DVSS.n5270 DVSS.n5268 0.0380882
R45442 DVSS.n5280 DVSS.n5268 0.0380882
R45443 DVSS.n5281 DVSS.n5280 0.0380882
R45444 DVSS.n5282 DVSS.n5281 0.0380882
R45445 DVSS.n5282 DVSS.n5264 0.0380882
R45446 DVSS.n5292 DVSS.n5264 0.0380882
R45447 DVSS.n5293 DVSS.n5292 0.0380882
R45448 DVSS.n5294 DVSS.n5293 0.0380882
R45449 DVSS.n5294 DVSS.n5260 0.0380882
R45450 DVSS.n5304 DVSS.n5260 0.0380882
R45451 DVSS.n5305 DVSS.n5304 0.0380882
R45452 DVSS.n5306 DVSS.n5305 0.0380882
R45453 DVSS.n5306 DVSS.n5256 0.0380882
R45454 DVSS.n5316 DVSS.n5256 0.0380882
R45455 DVSS.n5317 DVSS.n5316 0.0380882
R45456 DVSS.n5318 DVSS.n5317 0.0380882
R45457 DVSS.n5318 DVSS.n5252 0.0380882
R45458 DVSS.n5328 DVSS.n5252 0.0380882
R45459 DVSS.n5329 DVSS.n5328 0.0380882
R45460 DVSS.n5330 DVSS.n5329 0.0380882
R45461 DVSS.n5330 DVSS.n5248 0.0380882
R45462 DVSS.n5340 DVSS.n5248 0.0380882
R45463 DVSS.n5341 DVSS.n5340 0.0380882
R45464 DVSS.n5342 DVSS.n5341 0.0380882
R45465 DVSS.n5342 DVSS.n5244 0.0380882
R45466 DVSS.n5352 DVSS.n5244 0.0380882
R45467 DVSS.n5353 DVSS.n5352 0.0380882
R45468 DVSS.n5354 DVSS.n5353 0.0380882
R45469 DVSS.n5354 DVSS.n5240 0.0380882
R45470 DVSS.n5364 DVSS.n5240 0.0380882
R45471 DVSS.n5365 DVSS.n5364 0.0380882
R45472 DVSS.n5366 DVSS.n5365 0.0380882
R45473 DVSS.n5366 DVSS.n5236 0.0380882
R45474 DVSS.n5376 DVSS.n5236 0.0380882
R45475 DVSS.n5377 DVSS.n5376 0.0380882
R45476 DVSS.n5378 DVSS.n5377 0.0380882
R45477 DVSS.n5378 DVSS.n5232 0.0380882
R45478 DVSS.n5388 DVSS.n5232 0.0380882
R45479 DVSS.n5389 DVSS.n5388 0.0380882
R45480 DVSS.n5390 DVSS.n5389 0.0380882
R45481 DVSS.n5390 DVSS.n5228 0.0380882
R45482 DVSS.n5400 DVSS.n5228 0.0380882
R45483 DVSS.n5401 DVSS.n5400 0.0380882
R45484 DVSS.n5402 DVSS.n5401 0.0380882
R45485 DVSS.n5402 DVSS.n5224 0.0380882
R45486 DVSS.n5412 DVSS.n5224 0.0380882
R45487 DVSS.n5413 DVSS.n5412 0.0380882
R45488 DVSS.n5414 DVSS.n5413 0.0380882
R45489 DVSS.n5414 DVSS.n5220 0.0380882
R45490 DVSS.n5424 DVSS.n5220 0.0380882
R45491 DVSS.n5425 DVSS.n5424 0.0380882
R45492 DVSS.n5426 DVSS.n5425 0.0380882
R45493 DVSS.n5426 DVSS.n5216 0.0380882
R45494 DVSS.n5436 DVSS.n5216 0.0380882
R45495 DVSS.n5437 DVSS.n5436 0.0380882
R45496 DVSS.n5438 DVSS.n5437 0.0380882
R45497 DVSS.n5438 DVSS.n5212 0.0380882
R45498 DVSS.n5448 DVSS.n5212 0.0380882
R45499 DVSS.n5449 DVSS.n5448 0.0380882
R45500 DVSS.n5450 DVSS.n5449 0.0380882
R45501 DVSS.n5450 DVSS.n5208 0.0380882
R45502 DVSS.n5460 DVSS.n5208 0.0380882
R45503 DVSS.n5461 DVSS.n5460 0.0380882
R45504 DVSS.n5462 DVSS.n5461 0.0380882
R45505 DVSS.n5462 DVSS.n5204 0.0380882
R45506 DVSS.n5472 DVSS.n5204 0.0380882
R45507 DVSS.n5473 DVSS.n5472 0.0380882
R45508 DVSS.n5474 DVSS.n5473 0.0380882
R45509 DVSS.n5474 DVSS.n5200 0.0380882
R45510 DVSS.n5484 DVSS.n5200 0.0380882
R45511 DVSS.n5485 DVSS.n5484 0.0380882
R45512 DVSS.n5486 DVSS.n5485 0.0380882
R45513 DVSS.n5486 DVSS.n5196 0.0380882
R45514 DVSS.n5496 DVSS.n5196 0.0380882
R45515 DVSS.n5497 DVSS.n5496 0.0380882
R45516 DVSS.n5498 DVSS.n5497 0.0380882
R45517 DVSS.n5498 DVSS.n5192 0.0380882
R45518 DVSS.n5508 DVSS.n5192 0.0380882
R45519 DVSS.n5509 DVSS.n5508 0.0380882
R45520 DVSS.n5511 DVSS.n5509 0.0380882
R45521 DVSS.n5511 DVSS.n5510 0.0380882
R45522 DVSS.n5510 DVSS.n5187 0.0380882
R45523 DVSS.n5521 DVSS.n5187 0.0380882
R45524 DVSS.n5271 DVSS.n5269 0.0380882
R45525 DVSS.n5279 DVSS.n5269 0.0380882
R45526 DVSS.n5279 DVSS.n5267 0.0380882
R45527 DVSS.n5283 DVSS.n5267 0.0380882
R45528 DVSS.n5283 DVSS.n5265 0.0380882
R45529 DVSS.n5291 DVSS.n5265 0.0380882
R45530 DVSS.n5291 DVSS.n5263 0.0380882
R45531 DVSS.n5295 DVSS.n5263 0.0380882
R45532 DVSS.n5295 DVSS.n5261 0.0380882
R45533 DVSS.n5303 DVSS.n5261 0.0380882
R45534 DVSS.n5303 DVSS.n5259 0.0380882
R45535 DVSS.n5307 DVSS.n5259 0.0380882
R45536 DVSS.n5307 DVSS.n5257 0.0380882
R45537 DVSS.n5315 DVSS.n5257 0.0380882
R45538 DVSS.n5315 DVSS.n5255 0.0380882
R45539 DVSS.n5319 DVSS.n5255 0.0380882
R45540 DVSS.n5319 DVSS.n5253 0.0380882
R45541 DVSS.n5327 DVSS.n5253 0.0380882
R45542 DVSS.n5327 DVSS.n5251 0.0380882
R45543 DVSS.n5331 DVSS.n5251 0.0380882
R45544 DVSS.n5331 DVSS.n5249 0.0380882
R45545 DVSS.n5339 DVSS.n5249 0.0380882
R45546 DVSS.n5339 DVSS.n5247 0.0380882
R45547 DVSS.n5343 DVSS.n5247 0.0380882
R45548 DVSS.n5343 DVSS.n5245 0.0380882
R45549 DVSS.n5351 DVSS.n5245 0.0380882
R45550 DVSS.n5351 DVSS.n5243 0.0380882
R45551 DVSS.n5355 DVSS.n5243 0.0380882
R45552 DVSS.n5355 DVSS.n5241 0.0380882
R45553 DVSS.n5363 DVSS.n5241 0.0380882
R45554 DVSS.n5363 DVSS.n5239 0.0380882
R45555 DVSS.n5367 DVSS.n5239 0.0380882
R45556 DVSS.n5367 DVSS.n5237 0.0380882
R45557 DVSS.n5375 DVSS.n5237 0.0380882
R45558 DVSS.n5375 DVSS.n5235 0.0380882
R45559 DVSS.n5379 DVSS.n5235 0.0380882
R45560 DVSS.n5379 DVSS.n5233 0.0380882
R45561 DVSS.n5387 DVSS.n5233 0.0380882
R45562 DVSS.n5387 DVSS.n5231 0.0380882
R45563 DVSS.n5391 DVSS.n5231 0.0380882
R45564 DVSS.n5391 DVSS.n5229 0.0380882
R45565 DVSS.n5399 DVSS.n5229 0.0380882
R45566 DVSS.n5399 DVSS.n5227 0.0380882
R45567 DVSS.n5403 DVSS.n5227 0.0380882
R45568 DVSS.n5403 DVSS.n5225 0.0380882
R45569 DVSS.n5411 DVSS.n5225 0.0380882
R45570 DVSS.n5411 DVSS.n5223 0.0380882
R45571 DVSS.n5415 DVSS.n5223 0.0380882
R45572 DVSS.n5415 DVSS.n5221 0.0380882
R45573 DVSS.n5423 DVSS.n5221 0.0380882
R45574 DVSS.n5423 DVSS.n5219 0.0380882
R45575 DVSS.n5427 DVSS.n5219 0.0380882
R45576 DVSS.n5427 DVSS.n5217 0.0380882
R45577 DVSS.n5435 DVSS.n5217 0.0380882
R45578 DVSS.n5435 DVSS.n5215 0.0380882
R45579 DVSS.n5439 DVSS.n5215 0.0380882
R45580 DVSS.n5439 DVSS.n5213 0.0380882
R45581 DVSS.n5447 DVSS.n5213 0.0380882
R45582 DVSS.n5447 DVSS.n5211 0.0380882
R45583 DVSS.n5451 DVSS.n5211 0.0380882
R45584 DVSS.n5451 DVSS.n5209 0.0380882
R45585 DVSS.n5459 DVSS.n5209 0.0380882
R45586 DVSS.n5459 DVSS.n5207 0.0380882
R45587 DVSS.n5463 DVSS.n5207 0.0380882
R45588 DVSS.n5463 DVSS.n5205 0.0380882
R45589 DVSS.n5471 DVSS.n5205 0.0380882
R45590 DVSS.n5471 DVSS.n5203 0.0380882
R45591 DVSS.n5475 DVSS.n5203 0.0380882
R45592 DVSS.n5475 DVSS.n5201 0.0380882
R45593 DVSS.n5483 DVSS.n5201 0.0380882
R45594 DVSS.n5483 DVSS.n5199 0.0380882
R45595 DVSS.n5487 DVSS.n5199 0.0380882
R45596 DVSS.n5487 DVSS.n5197 0.0380882
R45597 DVSS.n5495 DVSS.n5197 0.0380882
R45598 DVSS.n5495 DVSS.n5195 0.0380882
R45599 DVSS.n5499 DVSS.n5195 0.0380882
R45600 DVSS.n5499 DVSS.n5193 0.0380882
R45601 DVSS.n5507 DVSS.n5193 0.0380882
R45602 DVSS.n5507 DVSS.n5191 0.0380882
R45603 DVSS.n5512 DVSS.n5191 0.0380882
R45604 DVSS.n5512 DVSS.n5189 0.0380882
R45605 DVSS.n5189 DVSS.n5188 0.0380882
R45606 DVSS.n5520 DVSS.n5188 0.0380882
R45607 DVSS.n4932 DVSS.n4931 0.0380882
R45608 DVSS.n4933 DVSS.n4932 0.0380882
R45609 DVSS.n4933 DVSS.n4926 0.0380882
R45610 DVSS.n4943 DVSS.n4926 0.0380882
R45611 DVSS.n4944 DVSS.n4943 0.0380882
R45612 DVSS.n4945 DVSS.n4944 0.0380882
R45613 DVSS.n4945 DVSS.n4924 0.0380882
R45614 DVSS.n4955 DVSS.n4924 0.0380882
R45615 DVSS.n4956 DVSS.n4955 0.0380882
R45616 DVSS.n4957 DVSS.n4956 0.0380882
R45617 DVSS.n4957 DVSS.n4922 0.0380882
R45618 DVSS.n4967 DVSS.n4922 0.0380882
R45619 DVSS.n4968 DVSS.n4967 0.0380882
R45620 DVSS.n4969 DVSS.n4968 0.0380882
R45621 DVSS.n4969 DVSS.n4920 0.0380882
R45622 DVSS.n4979 DVSS.n4920 0.0380882
R45623 DVSS.n4980 DVSS.n4979 0.0380882
R45624 DVSS.n4981 DVSS.n4980 0.0380882
R45625 DVSS.n4981 DVSS.n4918 0.0380882
R45626 DVSS.n4991 DVSS.n4918 0.0380882
R45627 DVSS.n4992 DVSS.n4991 0.0380882
R45628 DVSS.n4993 DVSS.n4992 0.0380882
R45629 DVSS.n4993 DVSS.n4916 0.0380882
R45630 DVSS.n5003 DVSS.n4916 0.0380882
R45631 DVSS.n5004 DVSS.n5003 0.0380882
R45632 DVSS.n5005 DVSS.n5004 0.0380882
R45633 DVSS.n5005 DVSS.n4914 0.0380882
R45634 DVSS.n5015 DVSS.n4914 0.0380882
R45635 DVSS.n5016 DVSS.n5015 0.0380882
R45636 DVSS.n5017 DVSS.n5016 0.0380882
R45637 DVSS.n5017 DVSS.n4912 0.0380882
R45638 DVSS.n5027 DVSS.n4912 0.0380882
R45639 DVSS.n5028 DVSS.n5027 0.0380882
R45640 DVSS.n5029 DVSS.n5028 0.0380882
R45641 DVSS.n5029 DVSS.n4910 0.0380882
R45642 DVSS.n5039 DVSS.n4910 0.0380882
R45643 DVSS.n5040 DVSS.n5039 0.0380882
R45644 DVSS.n5041 DVSS.n5040 0.0380882
R45645 DVSS.n5041 DVSS.n4908 0.0380882
R45646 DVSS.n5051 DVSS.n4908 0.0380882
R45647 DVSS.n5052 DVSS.n5051 0.0380882
R45648 DVSS.n5053 DVSS.n5052 0.0380882
R45649 DVSS.n5053 DVSS.n4906 0.0380882
R45650 DVSS.n5063 DVSS.n4906 0.0380882
R45651 DVSS.n5064 DVSS.n5063 0.0380882
R45652 DVSS.n5065 DVSS.n5064 0.0380882
R45653 DVSS.n5065 DVSS.n4904 0.0380882
R45654 DVSS.n5075 DVSS.n4904 0.0380882
R45655 DVSS.n5076 DVSS.n5075 0.0380882
R45656 DVSS.n5077 DVSS.n5076 0.0380882
R45657 DVSS.n5077 DVSS.n4902 0.0380882
R45658 DVSS.n5087 DVSS.n4902 0.0380882
R45659 DVSS.n5088 DVSS.n5087 0.0380882
R45660 DVSS.n5089 DVSS.n5088 0.0380882
R45661 DVSS.n5089 DVSS.n4900 0.0380882
R45662 DVSS.n5099 DVSS.n4900 0.0380882
R45663 DVSS.n5100 DVSS.n5099 0.0380882
R45664 DVSS.n5101 DVSS.n5100 0.0380882
R45665 DVSS.n5101 DVSS.n4898 0.0380882
R45666 DVSS.n5111 DVSS.n4898 0.0380882
R45667 DVSS.n5112 DVSS.n5111 0.0380882
R45668 DVSS.n5113 DVSS.n5112 0.0380882
R45669 DVSS.n5113 DVSS.n4896 0.0380882
R45670 DVSS.n5123 DVSS.n4896 0.0380882
R45671 DVSS.n5124 DVSS.n5123 0.0380882
R45672 DVSS.n5125 DVSS.n5124 0.0380882
R45673 DVSS.n5125 DVSS.n4894 0.0380882
R45674 DVSS.n5135 DVSS.n4894 0.0380882
R45675 DVSS.n5136 DVSS.n5135 0.0380882
R45676 DVSS.n5137 DVSS.n5136 0.0380882
R45677 DVSS.n5137 DVSS.n4892 0.0380882
R45678 DVSS.n5147 DVSS.n4892 0.0380882
R45679 DVSS.n5148 DVSS.n5147 0.0380882
R45680 DVSS.n5149 DVSS.n5148 0.0380882
R45681 DVSS.n5149 DVSS.n4890 0.0380882
R45682 DVSS.n5159 DVSS.n4890 0.0380882
R45683 DVSS.n5160 DVSS.n5159 0.0380882
R45684 DVSS.n5161 DVSS.n5160 0.0380882
R45685 DVSS.n5161 DVSS.n4888 0.0380882
R45686 DVSS.n5171 DVSS.n4888 0.0380882
R45687 DVSS.n5172 DVSS.n5171 0.0380882
R45688 DVSS.n7097 DVSS.n5172 0.0380882
R45689 DVSS.n7097 DVSS.n7096 0.0380882
R45690 DVSS.n4930 DVSS.n4929 0.0380882
R45691 DVSS.n4934 DVSS.n4929 0.0380882
R45692 DVSS.n4938 DVSS.n4934 0.0380882
R45693 DVSS.n4942 DVSS.n4938 0.0380882
R45694 DVSS.n4942 DVSS.n4925 0.0380882
R45695 DVSS.n4946 DVSS.n4925 0.0380882
R45696 DVSS.n4950 DVSS.n4946 0.0380882
R45697 DVSS.n4954 DVSS.n4950 0.0380882
R45698 DVSS.n4954 DVSS.n4923 0.0380882
R45699 DVSS.n4958 DVSS.n4923 0.0380882
R45700 DVSS.n4962 DVSS.n4958 0.0380882
R45701 DVSS.n4966 DVSS.n4962 0.0380882
R45702 DVSS.n4966 DVSS.n4921 0.0380882
R45703 DVSS.n4970 DVSS.n4921 0.0380882
R45704 DVSS.n4974 DVSS.n4970 0.0380882
R45705 DVSS.n4978 DVSS.n4974 0.0380882
R45706 DVSS.n4978 DVSS.n4919 0.0380882
R45707 DVSS.n4982 DVSS.n4919 0.0380882
R45708 DVSS.n4986 DVSS.n4982 0.0380882
R45709 DVSS.n4990 DVSS.n4986 0.0380882
R45710 DVSS.n4990 DVSS.n4917 0.0380882
R45711 DVSS.n4994 DVSS.n4917 0.0380882
R45712 DVSS.n4998 DVSS.n4994 0.0380882
R45713 DVSS.n5002 DVSS.n4998 0.0380882
R45714 DVSS.n5002 DVSS.n4915 0.0380882
R45715 DVSS.n5006 DVSS.n4915 0.0380882
R45716 DVSS.n5010 DVSS.n5006 0.0380882
R45717 DVSS.n5014 DVSS.n5010 0.0380882
R45718 DVSS.n5014 DVSS.n4913 0.0380882
R45719 DVSS.n5018 DVSS.n4913 0.0380882
R45720 DVSS.n5022 DVSS.n5018 0.0380882
R45721 DVSS.n5026 DVSS.n5022 0.0380882
R45722 DVSS.n5026 DVSS.n4911 0.0380882
R45723 DVSS.n5030 DVSS.n4911 0.0380882
R45724 DVSS.n5034 DVSS.n5030 0.0380882
R45725 DVSS.n5038 DVSS.n5034 0.0380882
R45726 DVSS.n5038 DVSS.n4909 0.0380882
R45727 DVSS.n5042 DVSS.n4909 0.0380882
R45728 DVSS.n5046 DVSS.n5042 0.0380882
R45729 DVSS.n5050 DVSS.n5046 0.0380882
R45730 DVSS.n5050 DVSS.n4907 0.0380882
R45731 DVSS.n5054 DVSS.n4907 0.0380882
R45732 DVSS.n5058 DVSS.n5054 0.0380882
R45733 DVSS.n5062 DVSS.n5058 0.0380882
R45734 DVSS.n5062 DVSS.n4905 0.0380882
R45735 DVSS.n5066 DVSS.n4905 0.0380882
R45736 DVSS.n5070 DVSS.n5066 0.0380882
R45737 DVSS.n5074 DVSS.n5070 0.0380882
R45738 DVSS.n5074 DVSS.n4903 0.0380882
R45739 DVSS.n5078 DVSS.n4903 0.0380882
R45740 DVSS.n5082 DVSS.n5078 0.0380882
R45741 DVSS.n5086 DVSS.n5082 0.0380882
R45742 DVSS.n5086 DVSS.n4901 0.0380882
R45743 DVSS.n5090 DVSS.n4901 0.0380882
R45744 DVSS.n5094 DVSS.n5090 0.0380882
R45745 DVSS.n5098 DVSS.n5094 0.0380882
R45746 DVSS.n5098 DVSS.n4899 0.0380882
R45747 DVSS.n5102 DVSS.n4899 0.0380882
R45748 DVSS.n5106 DVSS.n5102 0.0380882
R45749 DVSS.n5110 DVSS.n5106 0.0380882
R45750 DVSS.n5110 DVSS.n4897 0.0380882
R45751 DVSS.n5114 DVSS.n4897 0.0380882
R45752 DVSS.n5118 DVSS.n5114 0.0380882
R45753 DVSS.n5122 DVSS.n5118 0.0380882
R45754 DVSS.n5122 DVSS.n4895 0.0380882
R45755 DVSS.n5126 DVSS.n4895 0.0380882
R45756 DVSS.n5130 DVSS.n5126 0.0380882
R45757 DVSS.n5134 DVSS.n5130 0.0380882
R45758 DVSS.n5134 DVSS.n4893 0.0380882
R45759 DVSS.n5138 DVSS.n4893 0.0380882
R45760 DVSS.n5142 DVSS.n5138 0.0380882
R45761 DVSS.n5146 DVSS.n5142 0.0380882
R45762 DVSS.n5146 DVSS.n4891 0.0380882
R45763 DVSS.n5150 DVSS.n4891 0.0380882
R45764 DVSS.n5154 DVSS.n5150 0.0380882
R45765 DVSS.n5158 DVSS.n5154 0.0380882
R45766 DVSS.n5158 DVSS.n4889 0.0380882
R45767 DVSS.n5162 DVSS.n4889 0.0380882
R45768 DVSS.n5166 DVSS.n5162 0.0380882
R45769 DVSS.n5170 DVSS.n5166 0.0380882
R45770 DVSS.n5170 DVSS.n4887 0.0380882
R45771 DVSS.n7098 DVSS.n4887 0.0380882
R45772 DVSS.n7098 DVSS.n4884 0.0380882
R45773 DVSS.n7444 DVSS.n7111 0.0380882
R45774 DVSS.n7436 DVSS.n7111 0.0380882
R45775 DVSS.n7436 DVSS.n7435 0.0380882
R45776 DVSS.n7435 DVSS.n7434 0.0380882
R45777 DVSS.n7434 DVSS.n7115 0.0380882
R45778 DVSS.n7426 DVSS.n7115 0.0380882
R45779 DVSS.n7426 DVSS.n7425 0.0380882
R45780 DVSS.n7425 DVSS.n7424 0.0380882
R45781 DVSS.n7424 DVSS.n7121 0.0380882
R45782 DVSS.n7416 DVSS.n7121 0.0380882
R45783 DVSS.n7416 DVSS.n7415 0.0380882
R45784 DVSS.n7415 DVSS.n7414 0.0380882
R45785 DVSS.n7414 DVSS.n7127 0.0380882
R45786 DVSS.n7406 DVSS.n7127 0.0380882
R45787 DVSS.n7406 DVSS.n7405 0.0380882
R45788 DVSS.n7405 DVSS.n7404 0.0380882
R45789 DVSS.n7404 DVSS.n7133 0.0380882
R45790 DVSS.n7396 DVSS.n7133 0.0380882
R45791 DVSS.n7396 DVSS.n7395 0.0380882
R45792 DVSS.n7395 DVSS.n7394 0.0380882
R45793 DVSS.n7394 DVSS.n7139 0.0380882
R45794 DVSS.n7386 DVSS.n7139 0.0380882
R45795 DVSS.n7386 DVSS.n7385 0.0380882
R45796 DVSS.n7385 DVSS.n7384 0.0380882
R45797 DVSS.n7384 DVSS.n7145 0.0380882
R45798 DVSS.n7376 DVSS.n7145 0.0380882
R45799 DVSS.n7376 DVSS.n7375 0.0380882
R45800 DVSS.n7375 DVSS.n7374 0.0380882
R45801 DVSS.n7374 DVSS.n7151 0.0380882
R45802 DVSS.n7366 DVSS.n7151 0.0380882
R45803 DVSS.n7366 DVSS.n7365 0.0380882
R45804 DVSS.n7365 DVSS.n7364 0.0380882
R45805 DVSS.n7364 DVSS.n7157 0.0380882
R45806 DVSS.n7356 DVSS.n7157 0.0380882
R45807 DVSS.n7356 DVSS.n7355 0.0380882
R45808 DVSS.n7355 DVSS.n7354 0.0380882
R45809 DVSS.n7354 DVSS.n7163 0.0380882
R45810 DVSS.n7346 DVSS.n7163 0.0380882
R45811 DVSS.n7346 DVSS.n7345 0.0380882
R45812 DVSS.n7345 DVSS.n7344 0.0380882
R45813 DVSS.n7344 DVSS.n7169 0.0380882
R45814 DVSS.n7336 DVSS.n7169 0.0380882
R45815 DVSS.n7336 DVSS.n7335 0.0380882
R45816 DVSS.n7335 DVSS.n7334 0.0380882
R45817 DVSS.n7334 DVSS.n7175 0.0380882
R45818 DVSS.n7326 DVSS.n7175 0.0380882
R45819 DVSS.n7326 DVSS.n7325 0.0380882
R45820 DVSS.n7325 DVSS.n7324 0.0380882
R45821 DVSS.n7324 DVSS.n7181 0.0380882
R45822 DVSS.n7316 DVSS.n7181 0.0380882
R45823 DVSS.n7316 DVSS.n7315 0.0380882
R45824 DVSS.n7315 DVSS.n7314 0.0380882
R45825 DVSS.n7314 DVSS.n7187 0.0380882
R45826 DVSS.n7306 DVSS.n7187 0.0380882
R45827 DVSS.n7306 DVSS.n7305 0.0380882
R45828 DVSS.n7305 DVSS.n7304 0.0380882
R45829 DVSS.n7304 DVSS.n7193 0.0380882
R45830 DVSS.n7296 DVSS.n7193 0.0380882
R45831 DVSS.n7296 DVSS.n7295 0.0380882
R45832 DVSS.n7295 DVSS.n7294 0.0380882
R45833 DVSS.n7294 DVSS.n7199 0.0380882
R45834 DVSS.n7286 DVSS.n7199 0.0380882
R45835 DVSS.n7286 DVSS.n7285 0.0380882
R45836 DVSS.n7285 DVSS.n7284 0.0380882
R45837 DVSS.n7284 DVSS.n7205 0.0380882
R45838 DVSS.n7276 DVSS.n7205 0.0380882
R45839 DVSS.n7276 DVSS.n7275 0.0380882
R45840 DVSS.n7275 DVSS.n7274 0.0380882
R45841 DVSS.n7274 DVSS.n7211 0.0380882
R45842 DVSS.n7266 DVSS.n7211 0.0380882
R45843 DVSS.n7266 DVSS.n7265 0.0380882
R45844 DVSS.n7265 DVSS.n7264 0.0380882
R45845 DVSS.n7264 DVSS.n7217 0.0380882
R45846 DVSS.n7256 DVSS.n7217 0.0380882
R45847 DVSS.n7256 DVSS.n7255 0.0380882
R45848 DVSS.n7255 DVSS.n7254 0.0380882
R45849 DVSS.n7254 DVSS.n7223 0.0380882
R45850 DVSS.n7246 DVSS.n7223 0.0380882
R45851 DVSS.n7246 DVSS.n7245 0.0380882
R45852 DVSS.n7245 DVSS.n7244 0.0380882
R45853 DVSS.n7244 DVSS.n7229 0.0380882
R45854 DVSS.n7236 DVSS.n7229 0.0380882
R45855 DVSS.n7236 DVSS.n4828 0.0380882
R45856 DVSS.n7443 DVSS.n7112 0.0380882
R45857 DVSS.n7437 DVSS.n7112 0.0380882
R45858 DVSS.n7437 DVSS.n7114 0.0380882
R45859 DVSS.n7433 DVSS.n7114 0.0380882
R45860 DVSS.n7433 DVSS.n7116 0.0380882
R45861 DVSS.n7427 DVSS.n7116 0.0380882
R45862 DVSS.n7427 DVSS.n7120 0.0380882
R45863 DVSS.n7423 DVSS.n7120 0.0380882
R45864 DVSS.n7423 DVSS.n7122 0.0380882
R45865 DVSS.n7417 DVSS.n7122 0.0380882
R45866 DVSS.n7417 DVSS.n7126 0.0380882
R45867 DVSS.n7413 DVSS.n7126 0.0380882
R45868 DVSS.n7413 DVSS.n7128 0.0380882
R45869 DVSS.n7407 DVSS.n7128 0.0380882
R45870 DVSS.n7407 DVSS.n7132 0.0380882
R45871 DVSS.n7403 DVSS.n7132 0.0380882
R45872 DVSS.n7403 DVSS.n7134 0.0380882
R45873 DVSS.n7397 DVSS.n7134 0.0380882
R45874 DVSS.n7397 DVSS.n7138 0.0380882
R45875 DVSS.n7393 DVSS.n7138 0.0380882
R45876 DVSS.n7393 DVSS.n7140 0.0380882
R45877 DVSS.n7387 DVSS.n7140 0.0380882
R45878 DVSS.n7387 DVSS.n7144 0.0380882
R45879 DVSS.n7383 DVSS.n7144 0.0380882
R45880 DVSS.n7383 DVSS.n7146 0.0380882
R45881 DVSS.n7377 DVSS.n7146 0.0380882
R45882 DVSS.n7377 DVSS.n7150 0.0380882
R45883 DVSS.n7373 DVSS.n7150 0.0380882
R45884 DVSS.n7373 DVSS.n7152 0.0380882
R45885 DVSS.n7367 DVSS.n7152 0.0380882
R45886 DVSS.n7367 DVSS.n7156 0.0380882
R45887 DVSS.n7363 DVSS.n7156 0.0380882
R45888 DVSS.n7363 DVSS.n7158 0.0380882
R45889 DVSS.n7357 DVSS.n7158 0.0380882
R45890 DVSS.n7357 DVSS.n7162 0.0380882
R45891 DVSS.n7353 DVSS.n7162 0.0380882
R45892 DVSS.n7353 DVSS.n7164 0.0380882
R45893 DVSS.n7347 DVSS.n7164 0.0380882
R45894 DVSS.n7347 DVSS.n7168 0.0380882
R45895 DVSS.n7343 DVSS.n7168 0.0380882
R45896 DVSS.n7343 DVSS.n7170 0.0380882
R45897 DVSS.n7337 DVSS.n7170 0.0380882
R45898 DVSS.n7337 DVSS.n7174 0.0380882
R45899 DVSS.n7333 DVSS.n7174 0.0380882
R45900 DVSS.n7333 DVSS.n7176 0.0380882
R45901 DVSS.n7327 DVSS.n7176 0.0380882
R45902 DVSS.n7327 DVSS.n7180 0.0380882
R45903 DVSS.n7323 DVSS.n7180 0.0380882
R45904 DVSS.n7323 DVSS.n7182 0.0380882
R45905 DVSS.n7317 DVSS.n7182 0.0380882
R45906 DVSS.n7317 DVSS.n7186 0.0380882
R45907 DVSS.n7313 DVSS.n7186 0.0380882
R45908 DVSS.n7313 DVSS.n7188 0.0380882
R45909 DVSS.n7307 DVSS.n7188 0.0380882
R45910 DVSS.n7307 DVSS.n7192 0.0380882
R45911 DVSS.n7303 DVSS.n7192 0.0380882
R45912 DVSS.n7303 DVSS.n7194 0.0380882
R45913 DVSS.n7297 DVSS.n7194 0.0380882
R45914 DVSS.n7297 DVSS.n7198 0.0380882
R45915 DVSS.n7293 DVSS.n7198 0.0380882
R45916 DVSS.n7293 DVSS.n7200 0.0380882
R45917 DVSS.n7287 DVSS.n7200 0.0380882
R45918 DVSS.n7287 DVSS.n7204 0.0380882
R45919 DVSS.n7283 DVSS.n7204 0.0380882
R45920 DVSS.n7283 DVSS.n7206 0.0380882
R45921 DVSS.n7277 DVSS.n7206 0.0380882
R45922 DVSS.n7277 DVSS.n7210 0.0380882
R45923 DVSS.n7273 DVSS.n7210 0.0380882
R45924 DVSS.n7273 DVSS.n7212 0.0380882
R45925 DVSS.n7267 DVSS.n7212 0.0380882
R45926 DVSS.n7267 DVSS.n7216 0.0380882
R45927 DVSS.n7263 DVSS.n7216 0.0380882
R45928 DVSS.n7263 DVSS.n7218 0.0380882
R45929 DVSS.n7257 DVSS.n7218 0.0380882
R45930 DVSS.n7257 DVSS.n7222 0.0380882
R45931 DVSS.n7253 DVSS.n7222 0.0380882
R45932 DVSS.n7253 DVSS.n7224 0.0380882
R45933 DVSS.n7247 DVSS.n7224 0.0380882
R45934 DVSS.n7247 DVSS.n7228 0.0380882
R45935 DVSS.n7243 DVSS.n7228 0.0380882
R45936 DVSS.n7243 DVSS.n7230 0.0380882
R45937 DVSS.n7237 DVSS.n7230 0.0380882
R45938 DVSS.n7237 DVSS.n7235 0.0380882
R45939 DVSS.n7790 DVSS.n4821 0.0380882
R45940 DVSS.n7790 DVSS.n7789 0.0380882
R45941 DVSS.n7789 DVSS.n7788 0.0380882
R45942 DVSS.n7788 DVSS.n7507 0.0380882
R45943 DVSS.n7778 DVSS.n7507 0.0380882
R45944 DVSS.n7778 DVSS.n7777 0.0380882
R45945 DVSS.n7777 DVSS.n7776 0.0380882
R45946 DVSS.n7776 DVSS.n7509 0.0380882
R45947 DVSS.n7766 DVSS.n7509 0.0380882
R45948 DVSS.n7766 DVSS.n7765 0.0380882
R45949 DVSS.n7765 DVSS.n7764 0.0380882
R45950 DVSS.n7764 DVSS.n7511 0.0380882
R45951 DVSS.n7754 DVSS.n7511 0.0380882
R45952 DVSS.n7754 DVSS.n7753 0.0380882
R45953 DVSS.n7753 DVSS.n7752 0.0380882
R45954 DVSS.n7752 DVSS.n7513 0.0380882
R45955 DVSS.n7742 DVSS.n7513 0.0380882
R45956 DVSS.n7742 DVSS.n7741 0.0380882
R45957 DVSS.n7741 DVSS.n7740 0.0380882
R45958 DVSS.n7740 DVSS.n7515 0.0380882
R45959 DVSS.n7730 DVSS.n7515 0.0380882
R45960 DVSS.n7730 DVSS.n7729 0.0380882
R45961 DVSS.n7729 DVSS.n7728 0.0380882
R45962 DVSS.n7728 DVSS.n7517 0.0380882
R45963 DVSS.n7718 DVSS.n7517 0.0380882
R45964 DVSS.n7718 DVSS.n7717 0.0380882
R45965 DVSS.n7717 DVSS.n7716 0.0380882
R45966 DVSS.n7716 DVSS.n7519 0.0380882
R45967 DVSS.n7706 DVSS.n7519 0.0380882
R45968 DVSS.n7706 DVSS.n7705 0.0380882
R45969 DVSS.n7705 DVSS.n7704 0.0380882
R45970 DVSS.n7704 DVSS.n7521 0.0380882
R45971 DVSS.n7694 DVSS.n7521 0.0380882
R45972 DVSS.n7694 DVSS.n7693 0.0380882
R45973 DVSS.n7693 DVSS.n7692 0.0380882
R45974 DVSS.n7692 DVSS.n7523 0.0380882
R45975 DVSS.n7682 DVSS.n7523 0.0380882
R45976 DVSS.n7682 DVSS.n7681 0.0380882
R45977 DVSS.n7681 DVSS.n7680 0.0380882
R45978 DVSS.n7680 DVSS.n7525 0.0380882
R45979 DVSS.n7670 DVSS.n7525 0.0380882
R45980 DVSS.n7670 DVSS.n7669 0.0380882
R45981 DVSS.n7669 DVSS.n7668 0.0380882
R45982 DVSS.n7668 DVSS.n7527 0.0380882
R45983 DVSS.n7658 DVSS.n7527 0.0380882
R45984 DVSS.n7658 DVSS.n7657 0.0380882
R45985 DVSS.n7657 DVSS.n7656 0.0380882
R45986 DVSS.n7656 DVSS.n7529 0.0380882
R45987 DVSS.n7646 DVSS.n7529 0.0380882
R45988 DVSS.n7646 DVSS.n7645 0.0380882
R45989 DVSS.n7645 DVSS.n7644 0.0380882
R45990 DVSS.n7644 DVSS.n7531 0.0380882
R45991 DVSS.n7634 DVSS.n7531 0.0380882
R45992 DVSS.n7634 DVSS.n7633 0.0380882
R45993 DVSS.n7633 DVSS.n7632 0.0380882
R45994 DVSS.n7632 DVSS.n7533 0.0380882
R45995 DVSS.n7622 DVSS.n7533 0.0380882
R45996 DVSS.n7622 DVSS.n7621 0.0380882
R45997 DVSS.n7621 DVSS.n7620 0.0380882
R45998 DVSS.n7620 DVSS.n7535 0.0380882
R45999 DVSS.n7610 DVSS.n7535 0.0380882
R46000 DVSS.n7610 DVSS.n7609 0.0380882
R46001 DVSS.n7609 DVSS.n7608 0.0380882
R46002 DVSS.n7608 DVSS.n7537 0.0380882
R46003 DVSS.n7598 DVSS.n7537 0.0380882
R46004 DVSS.n7598 DVSS.n7597 0.0380882
R46005 DVSS.n7597 DVSS.n7596 0.0380882
R46006 DVSS.n7596 DVSS.n7539 0.0380882
R46007 DVSS.n7586 DVSS.n7539 0.0380882
R46008 DVSS.n7586 DVSS.n7585 0.0380882
R46009 DVSS.n7585 DVSS.n7584 0.0380882
R46010 DVSS.n7584 DVSS.n7541 0.0380882
R46011 DVSS.n7574 DVSS.n7541 0.0380882
R46012 DVSS.n7574 DVSS.n7573 0.0380882
R46013 DVSS.n7573 DVSS.n7572 0.0380882
R46014 DVSS.n7572 DVSS.n7543 0.0380882
R46015 DVSS.n7562 DVSS.n7543 0.0380882
R46016 DVSS.n7562 DVSS.n7561 0.0380882
R46017 DVSS.n7561 DVSS.n7560 0.0380882
R46018 DVSS.n7560 DVSS.n7545 0.0380882
R46019 DVSS.n7550 DVSS.n7545 0.0380882
R46020 DVSS.n7550 DVSS.n7549 0.0380882
R46021 DVSS.n7549 DVSS.n4814 0.0380882
R46022 DVSS.n7792 DVSS.n7791 0.0380882
R46023 DVSS.n7791 DVSS.n7506 0.0380882
R46024 DVSS.n7787 DVSS.n7506 0.0380882
R46025 DVSS.n7787 DVSS.n7783 0.0380882
R46026 DVSS.n7783 DVSS.n7782 0.0380882
R46027 DVSS.n7782 DVSS.n7508 0.0380882
R46028 DVSS.n7775 DVSS.n7508 0.0380882
R46029 DVSS.n7775 DVSS.n7771 0.0380882
R46030 DVSS.n7771 DVSS.n7770 0.0380882
R46031 DVSS.n7770 DVSS.n7510 0.0380882
R46032 DVSS.n7763 DVSS.n7510 0.0380882
R46033 DVSS.n7763 DVSS.n7759 0.0380882
R46034 DVSS.n7759 DVSS.n7758 0.0380882
R46035 DVSS.n7758 DVSS.n7512 0.0380882
R46036 DVSS.n7751 DVSS.n7512 0.0380882
R46037 DVSS.n7751 DVSS.n7747 0.0380882
R46038 DVSS.n7747 DVSS.n7746 0.0380882
R46039 DVSS.n7746 DVSS.n7514 0.0380882
R46040 DVSS.n7739 DVSS.n7514 0.0380882
R46041 DVSS.n7739 DVSS.n7735 0.0380882
R46042 DVSS.n7735 DVSS.n7734 0.0380882
R46043 DVSS.n7734 DVSS.n7516 0.0380882
R46044 DVSS.n7727 DVSS.n7516 0.0380882
R46045 DVSS.n7727 DVSS.n7723 0.0380882
R46046 DVSS.n7723 DVSS.n7722 0.0380882
R46047 DVSS.n7722 DVSS.n7518 0.0380882
R46048 DVSS.n7715 DVSS.n7518 0.0380882
R46049 DVSS.n7715 DVSS.n7711 0.0380882
R46050 DVSS.n7711 DVSS.n7710 0.0380882
R46051 DVSS.n7710 DVSS.n7520 0.0380882
R46052 DVSS.n7703 DVSS.n7520 0.0380882
R46053 DVSS.n7703 DVSS.n7699 0.0380882
R46054 DVSS.n7699 DVSS.n7698 0.0380882
R46055 DVSS.n7698 DVSS.n7522 0.0380882
R46056 DVSS.n7691 DVSS.n7522 0.0380882
R46057 DVSS.n7691 DVSS.n7687 0.0380882
R46058 DVSS.n7687 DVSS.n7686 0.0380882
R46059 DVSS.n7686 DVSS.n7524 0.0380882
R46060 DVSS.n7679 DVSS.n7524 0.0380882
R46061 DVSS.n7679 DVSS.n7675 0.0380882
R46062 DVSS.n7675 DVSS.n7674 0.0380882
R46063 DVSS.n7674 DVSS.n7526 0.0380882
R46064 DVSS.n7667 DVSS.n7526 0.0380882
R46065 DVSS.n7667 DVSS.n7663 0.0380882
R46066 DVSS.n7663 DVSS.n7662 0.0380882
R46067 DVSS.n7662 DVSS.n7528 0.0380882
R46068 DVSS.n7655 DVSS.n7528 0.0380882
R46069 DVSS.n7655 DVSS.n7651 0.0380882
R46070 DVSS.n7651 DVSS.n7650 0.0380882
R46071 DVSS.n7650 DVSS.n7530 0.0380882
R46072 DVSS.n7643 DVSS.n7530 0.0380882
R46073 DVSS.n7643 DVSS.n7639 0.0380882
R46074 DVSS.n7639 DVSS.n7638 0.0380882
R46075 DVSS.n7638 DVSS.n7532 0.0380882
R46076 DVSS.n7631 DVSS.n7532 0.0380882
R46077 DVSS.n7631 DVSS.n7627 0.0380882
R46078 DVSS.n7627 DVSS.n7626 0.0380882
R46079 DVSS.n7626 DVSS.n7534 0.0380882
R46080 DVSS.n7619 DVSS.n7534 0.0380882
R46081 DVSS.n7619 DVSS.n7615 0.0380882
R46082 DVSS.n7615 DVSS.n7614 0.0380882
R46083 DVSS.n7614 DVSS.n7536 0.0380882
R46084 DVSS.n7607 DVSS.n7536 0.0380882
R46085 DVSS.n7607 DVSS.n7603 0.0380882
R46086 DVSS.n7603 DVSS.n7602 0.0380882
R46087 DVSS.n7602 DVSS.n7538 0.0380882
R46088 DVSS.n7595 DVSS.n7538 0.0380882
R46089 DVSS.n7595 DVSS.n7591 0.0380882
R46090 DVSS.n7591 DVSS.n7590 0.0380882
R46091 DVSS.n7590 DVSS.n7540 0.0380882
R46092 DVSS.n7583 DVSS.n7540 0.0380882
R46093 DVSS.n7583 DVSS.n7579 0.0380882
R46094 DVSS.n7579 DVSS.n7578 0.0380882
R46095 DVSS.n7578 DVSS.n7542 0.0380882
R46096 DVSS.n7571 DVSS.n7542 0.0380882
R46097 DVSS.n7571 DVSS.n7567 0.0380882
R46098 DVSS.n7567 DVSS.n7566 0.0380882
R46099 DVSS.n7566 DVSS.n7544 0.0380882
R46100 DVSS.n7559 DVSS.n7544 0.0380882
R46101 DVSS.n7559 DVSS.n7555 0.0380882
R46102 DVSS.n7555 DVSS.n7554 0.0380882
R46103 DVSS.n7554 DVSS.n7548 0.0380882
R46104 DVSS.n7548 DVSS.n7547 0.0380882
R46105 DVSS.n4807 DVSS.n4474 0.0380882
R46106 DVSS.n4799 DVSS.n4474 0.0380882
R46107 DVSS.n4799 DVSS.n4798 0.0380882
R46108 DVSS.n4798 DVSS.n4797 0.0380882
R46109 DVSS.n4797 DVSS.n4478 0.0380882
R46110 DVSS.n4789 DVSS.n4478 0.0380882
R46111 DVSS.n4789 DVSS.n4788 0.0380882
R46112 DVSS.n4788 DVSS.n4787 0.0380882
R46113 DVSS.n4787 DVSS.n4484 0.0380882
R46114 DVSS.n4779 DVSS.n4484 0.0380882
R46115 DVSS.n4779 DVSS.n4778 0.0380882
R46116 DVSS.n4778 DVSS.n4777 0.0380882
R46117 DVSS.n4777 DVSS.n4490 0.0380882
R46118 DVSS.n4769 DVSS.n4490 0.0380882
R46119 DVSS.n4769 DVSS.n4768 0.0380882
R46120 DVSS.n4768 DVSS.n4767 0.0380882
R46121 DVSS.n4767 DVSS.n4496 0.0380882
R46122 DVSS.n4759 DVSS.n4496 0.0380882
R46123 DVSS.n4759 DVSS.n4758 0.0380882
R46124 DVSS.n4758 DVSS.n4757 0.0380882
R46125 DVSS.n4757 DVSS.n4502 0.0380882
R46126 DVSS.n4749 DVSS.n4502 0.0380882
R46127 DVSS.n4749 DVSS.n4748 0.0380882
R46128 DVSS.n4748 DVSS.n4747 0.0380882
R46129 DVSS.n4747 DVSS.n4508 0.0380882
R46130 DVSS.n4739 DVSS.n4508 0.0380882
R46131 DVSS.n4739 DVSS.n4738 0.0380882
R46132 DVSS.n4738 DVSS.n4737 0.0380882
R46133 DVSS.n4737 DVSS.n4514 0.0380882
R46134 DVSS.n4729 DVSS.n4514 0.0380882
R46135 DVSS.n4729 DVSS.n4728 0.0380882
R46136 DVSS.n4728 DVSS.n4727 0.0380882
R46137 DVSS.n4727 DVSS.n4520 0.0380882
R46138 DVSS.n4719 DVSS.n4520 0.0380882
R46139 DVSS.n4719 DVSS.n4718 0.0380882
R46140 DVSS.n4718 DVSS.n4717 0.0380882
R46141 DVSS.n4717 DVSS.n4526 0.0380882
R46142 DVSS.n4709 DVSS.n4526 0.0380882
R46143 DVSS.n4709 DVSS.n4708 0.0380882
R46144 DVSS.n4708 DVSS.n4707 0.0380882
R46145 DVSS.n4707 DVSS.n4532 0.0380882
R46146 DVSS.n4699 DVSS.n4532 0.0380882
R46147 DVSS.n4699 DVSS.n4698 0.0380882
R46148 DVSS.n4698 DVSS.n4697 0.0380882
R46149 DVSS.n4697 DVSS.n4538 0.0380882
R46150 DVSS.n4689 DVSS.n4538 0.0380882
R46151 DVSS.n4689 DVSS.n4688 0.0380882
R46152 DVSS.n4688 DVSS.n4687 0.0380882
R46153 DVSS.n4687 DVSS.n4544 0.0380882
R46154 DVSS.n4679 DVSS.n4544 0.0380882
R46155 DVSS.n4679 DVSS.n4678 0.0380882
R46156 DVSS.n4678 DVSS.n4677 0.0380882
R46157 DVSS.n4677 DVSS.n4550 0.0380882
R46158 DVSS.n4669 DVSS.n4550 0.0380882
R46159 DVSS.n4669 DVSS.n4668 0.0380882
R46160 DVSS.n4668 DVSS.n4667 0.0380882
R46161 DVSS.n4667 DVSS.n4556 0.0380882
R46162 DVSS.n4659 DVSS.n4556 0.0380882
R46163 DVSS.n4659 DVSS.n4658 0.0380882
R46164 DVSS.n4658 DVSS.n4657 0.0380882
R46165 DVSS.n4657 DVSS.n4562 0.0380882
R46166 DVSS.n4649 DVSS.n4562 0.0380882
R46167 DVSS.n4649 DVSS.n4648 0.0380882
R46168 DVSS.n4648 DVSS.n4647 0.0380882
R46169 DVSS.n4647 DVSS.n4568 0.0380882
R46170 DVSS.n4639 DVSS.n4568 0.0380882
R46171 DVSS.n4639 DVSS.n4638 0.0380882
R46172 DVSS.n4638 DVSS.n4637 0.0380882
R46173 DVSS.n4637 DVSS.n4574 0.0380882
R46174 DVSS.n4629 DVSS.n4574 0.0380882
R46175 DVSS.n4629 DVSS.n4628 0.0380882
R46176 DVSS.n4628 DVSS.n4627 0.0380882
R46177 DVSS.n4627 DVSS.n4580 0.0380882
R46178 DVSS.n4619 DVSS.n4580 0.0380882
R46179 DVSS.n4619 DVSS.n4618 0.0380882
R46180 DVSS.n4618 DVSS.n4617 0.0380882
R46181 DVSS.n4617 DVSS.n4586 0.0380882
R46182 DVSS.n4609 DVSS.n4586 0.0380882
R46183 DVSS.n4609 DVSS.n4608 0.0380882
R46184 DVSS.n4608 DVSS.n4607 0.0380882
R46185 DVSS.n4607 DVSS.n4592 0.0380882
R46186 DVSS.n4599 DVSS.n4592 0.0380882
R46187 DVSS.n4599 DVSS.n4462 0.0380882
R46188 DVSS.n4806 DVSS.n4475 0.0380882
R46189 DVSS.n4800 DVSS.n4475 0.0380882
R46190 DVSS.n4800 DVSS.n4477 0.0380882
R46191 DVSS.n4796 DVSS.n4477 0.0380882
R46192 DVSS.n4796 DVSS.n4479 0.0380882
R46193 DVSS.n4790 DVSS.n4479 0.0380882
R46194 DVSS.n4790 DVSS.n4483 0.0380882
R46195 DVSS.n4786 DVSS.n4483 0.0380882
R46196 DVSS.n4786 DVSS.n4485 0.0380882
R46197 DVSS.n4780 DVSS.n4485 0.0380882
R46198 DVSS.n4780 DVSS.n4489 0.0380882
R46199 DVSS.n4776 DVSS.n4489 0.0380882
R46200 DVSS.n4776 DVSS.n4491 0.0380882
R46201 DVSS.n4770 DVSS.n4491 0.0380882
R46202 DVSS.n4770 DVSS.n4495 0.0380882
R46203 DVSS.n4766 DVSS.n4495 0.0380882
R46204 DVSS.n4766 DVSS.n4497 0.0380882
R46205 DVSS.n4760 DVSS.n4497 0.0380882
R46206 DVSS.n4760 DVSS.n4501 0.0380882
R46207 DVSS.n4756 DVSS.n4501 0.0380882
R46208 DVSS.n4756 DVSS.n4503 0.0380882
R46209 DVSS.n4750 DVSS.n4503 0.0380882
R46210 DVSS.n4750 DVSS.n4507 0.0380882
R46211 DVSS.n4746 DVSS.n4507 0.0380882
R46212 DVSS.n4746 DVSS.n4509 0.0380882
R46213 DVSS.n4740 DVSS.n4509 0.0380882
R46214 DVSS.n4740 DVSS.n4513 0.0380882
R46215 DVSS.n4736 DVSS.n4513 0.0380882
R46216 DVSS.n4736 DVSS.n4515 0.0380882
R46217 DVSS.n4730 DVSS.n4515 0.0380882
R46218 DVSS.n4730 DVSS.n4519 0.0380882
R46219 DVSS.n4726 DVSS.n4519 0.0380882
R46220 DVSS.n4726 DVSS.n4521 0.0380882
R46221 DVSS.n4720 DVSS.n4521 0.0380882
R46222 DVSS.n4720 DVSS.n4525 0.0380882
R46223 DVSS.n4716 DVSS.n4525 0.0380882
R46224 DVSS.n4716 DVSS.n4527 0.0380882
R46225 DVSS.n4710 DVSS.n4527 0.0380882
R46226 DVSS.n4710 DVSS.n4531 0.0380882
R46227 DVSS.n4706 DVSS.n4531 0.0380882
R46228 DVSS.n4706 DVSS.n4533 0.0380882
R46229 DVSS.n4700 DVSS.n4533 0.0380882
R46230 DVSS.n4700 DVSS.n4537 0.0380882
R46231 DVSS.n4696 DVSS.n4537 0.0380882
R46232 DVSS.n4696 DVSS.n4539 0.0380882
R46233 DVSS.n4690 DVSS.n4539 0.0380882
R46234 DVSS.n4690 DVSS.n4543 0.0380882
R46235 DVSS.n4686 DVSS.n4543 0.0380882
R46236 DVSS.n4686 DVSS.n4545 0.0380882
R46237 DVSS.n4680 DVSS.n4545 0.0380882
R46238 DVSS.n4680 DVSS.n4549 0.0380882
R46239 DVSS.n4676 DVSS.n4549 0.0380882
R46240 DVSS.n4676 DVSS.n4551 0.0380882
R46241 DVSS.n4670 DVSS.n4551 0.0380882
R46242 DVSS.n4670 DVSS.n4555 0.0380882
R46243 DVSS.n4666 DVSS.n4555 0.0380882
R46244 DVSS.n4666 DVSS.n4557 0.0380882
R46245 DVSS.n4660 DVSS.n4557 0.0380882
R46246 DVSS.n4660 DVSS.n4561 0.0380882
R46247 DVSS.n4656 DVSS.n4561 0.0380882
R46248 DVSS.n4656 DVSS.n4563 0.0380882
R46249 DVSS.n4650 DVSS.n4563 0.0380882
R46250 DVSS.n4650 DVSS.n4567 0.0380882
R46251 DVSS.n4646 DVSS.n4567 0.0380882
R46252 DVSS.n4646 DVSS.n4569 0.0380882
R46253 DVSS.n4640 DVSS.n4569 0.0380882
R46254 DVSS.n4640 DVSS.n4573 0.0380882
R46255 DVSS.n4636 DVSS.n4573 0.0380882
R46256 DVSS.n4636 DVSS.n4575 0.0380882
R46257 DVSS.n4630 DVSS.n4575 0.0380882
R46258 DVSS.n4630 DVSS.n4579 0.0380882
R46259 DVSS.n4626 DVSS.n4579 0.0380882
R46260 DVSS.n4626 DVSS.n4581 0.0380882
R46261 DVSS.n4620 DVSS.n4581 0.0380882
R46262 DVSS.n4620 DVSS.n4585 0.0380882
R46263 DVSS.n4616 DVSS.n4585 0.0380882
R46264 DVSS.n4616 DVSS.n4587 0.0380882
R46265 DVSS.n4610 DVSS.n4587 0.0380882
R46266 DVSS.n4610 DVSS.n4591 0.0380882
R46267 DVSS.n4606 DVSS.n4591 0.0380882
R46268 DVSS.n4606 DVSS.n4593 0.0380882
R46269 DVSS.n4600 DVSS.n4593 0.0380882
R46270 DVSS.n4600 DVSS.n4598 0.0380882
R46271 DVSS.n8085 DVSS.n4365 0.0380882
R46272 DVSS.n8085 DVSS.n8084 0.0380882
R46273 DVSS.n8084 DVSS.n8083 0.0380882
R46274 DVSS.n8083 DVSS.n4418 0.0380882
R46275 DVSS.n8073 DVSS.n4418 0.0380882
R46276 DVSS.n8073 DVSS.n8072 0.0380882
R46277 DVSS.n8072 DVSS.n8071 0.0380882
R46278 DVSS.n8071 DVSS.n4420 0.0380882
R46279 DVSS.n8061 DVSS.n4420 0.0380882
R46280 DVSS.n8061 DVSS.n8060 0.0380882
R46281 DVSS.n8060 DVSS.n8059 0.0380882
R46282 DVSS.n8059 DVSS.n4422 0.0380882
R46283 DVSS.n8049 DVSS.n4422 0.0380882
R46284 DVSS.n8049 DVSS.n8048 0.0380882
R46285 DVSS.n8048 DVSS.n8047 0.0380882
R46286 DVSS.n8047 DVSS.n4424 0.0380882
R46287 DVSS.n8037 DVSS.n4424 0.0380882
R46288 DVSS.n8037 DVSS.n8036 0.0380882
R46289 DVSS.n8036 DVSS.n8035 0.0380882
R46290 DVSS.n8035 DVSS.n4426 0.0380882
R46291 DVSS.n8025 DVSS.n4426 0.0380882
R46292 DVSS.n8025 DVSS.n8024 0.0380882
R46293 DVSS.n8024 DVSS.n8023 0.0380882
R46294 DVSS.n8023 DVSS.n4428 0.0380882
R46295 DVSS.n8013 DVSS.n4428 0.0380882
R46296 DVSS.n8013 DVSS.n8012 0.0380882
R46297 DVSS.n8012 DVSS.n8011 0.0380882
R46298 DVSS.n8011 DVSS.n4430 0.0380882
R46299 DVSS.n8001 DVSS.n4430 0.0380882
R46300 DVSS.n8001 DVSS.n8000 0.0380882
R46301 DVSS.n8000 DVSS.n7999 0.0380882
R46302 DVSS.n7999 DVSS.n4432 0.0380882
R46303 DVSS.n7989 DVSS.n4432 0.0380882
R46304 DVSS.n7989 DVSS.n7988 0.0380882
R46305 DVSS.n7988 DVSS.n7987 0.0380882
R46306 DVSS.n7987 DVSS.n4434 0.0380882
R46307 DVSS.n7977 DVSS.n4434 0.0380882
R46308 DVSS.n7977 DVSS.n7976 0.0380882
R46309 DVSS.n7976 DVSS.n7975 0.0380882
R46310 DVSS.n7975 DVSS.n4436 0.0380882
R46311 DVSS.n7965 DVSS.n4436 0.0380882
R46312 DVSS.n7965 DVSS.n7964 0.0380882
R46313 DVSS.n7964 DVSS.n7963 0.0380882
R46314 DVSS.n7963 DVSS.n4438 0.0380882
R46315 DVSS.n7953 DVSS.n4438 0.0380882
R46316 DVSS.n7953 DVSS.n7952 0.0380882
R46317 DVSS.n7952 DVSS.n7951 0.0380882
R46318 DVSS.n7951 DVSS.n4440 0.0380882
R46319 DVSS.n7941 DVSS.n4440 0.0380882
R46320 DVSS.n7941 DVSS.n7940 0.0380882
R46321 DVSS.n7940 DVSS.n7939 0.0380882
R46322 DVSS.n7939 DVSS.n4442 0.0380882
R46323 DVSS.n7929 DVSS.n4442 0.0380882
R46324 DVSS.n7929 DVSS.n7928 0.0380882
R46325 DVSS.n7928 DVSS.n7927 0.0380882
R46326 DVSS.n7927 DVSS.n4444 0.0380882
R46327 DVSS.n7917 DVSS.n4444 0.0380882
R46328 DVSS.n7917 DVSS.n7916 0.0380882
R46329 DVSS.n7916 DVSS.n7915 0.0380882
R46330 DVSS.n7915 DVSS.n4446 0.0380882
R46331 DVSS.n7905 DVSS.n4446 0.0380882
R46332 DVSS.n7905 DVSS.n7904 0.0380882
R46333 DVSS.n7904 DVSS.n7903 0.0380882
R46334 DVSS.n7903 DVSS.n4448 0.0380882
R46335 DVSS.n7893 DVSS.n4448 0.0380882
R46336 DVSS.n7893 DVSS.n7892 0.0380882
R46337 DVSS.n7892 DVSS.n7891 0.0380882
R46338 DVSS.n7891 DVSS.n4450 0.0380882
R46339 DVSS.n7881 DVSS.n4450 0.0380882
R46340 DVSS.n7881 DVSS.n7880 0.0380882
R46341 DVSS.n7880 DVSS.n7879 0.0380882
R46342 DVSS.n7879 DVSS.n4452 0.0380882
R46343 DVSS.n7869 DVSS.n4452 0.0380882
R46344 DVSS.n7869 DVSS.n7868 0.0380882
R46345 DVSS.n7868 DVSS.n7867 0.0380882
R46346 DVSS.n7867 DVSS.n4454 0.0380882
R46347 DVSS.n7857 DVSS.n4454 0.0380882
R46348 DVSS.n7857 DVSS.n7856 0.0380882
R46349 DVSS.n7856 DVSS.n7855 0.0380882
R46350 DVSS.n7855 DVSS.n4456 0.0380882
R46351 DVSS.n7845 DVSS.n4456 0.0380882
R46352 DVSS.n7845 DVSS.n7844 0.0380882
R46353 DVSS.n7844 DVSS.n7843 0.0380882
R46354 DVSS.n8087 DVSS.n8086 0.0380882
R46355 DVSS.n8086 DVSS.n4417 0.0380882
R46356 DVSS.n8082 DVSS.n4417 0.0380882
R46357 DVSS.n8082 DVSS.n8078 0.0380882
R46358 DVSS.n8078 DVSS.n8077 0.0380882
R46359 DVSS.n8077 DVSS.n4419 0.0380882
R46360 DVSS.n8070 DVSS.n4419 0.0380882
R46361 DVSS.n8070 DVSS.n8066 0.0380882
R46362 DVSS.n8066 DVSS.n8065 0.0380882
R46363 DVSS.n8065 DVSS.n4421 0.0380882
R46364 DVSS.n8058 DVSS.n4421 0.0380882
R46365 DVSS.n8058 DVSS.n8054 0.0380882
R46366 DVSS.n8054 DVSS.n8053 0.0380882
R46367 DVSS.n8053 DVSS.n4423 0.0380882
R46368 DVSS.n8046 DVSS.n4423 0.0380882
R46369 DVSS.n8046 DVSS.n8042 0.0380882
R46370 DVSS.n8042 DVSS.n8041 0.0380882
R46371 DVSS.n8041 DVSS.n4425 0.0380882
R46372 DVSS.n8034 DVSS.n4425 0.0380882
R46373 DVSS.n8034 DVSS.n8030 0.0380882
R46374 DVSS.n8030 DVSS.n8029 0.0380882
R46375 DVSS.n8029 DVSS.n4427 0.0380882
R46376 DVSS.n8022 DVSS.n4427 0.0380882
R46377 DVSS.n8022 DVSS.n8018 0.0380882
R46378 DVSS.n8018 DVSS.n8017 0.0380882
R46379 DVSS.n8017 DVSS.n4429 0.0380882
R46380 DVSS.n8010 DVSS.n4429 0.0380882
R46381 DVSS.n8010 DVSS.n8006 0.0380882
R46382 DVSS.n8006 DVSS.n8005 0.0380882
R46383 DVSS.n8005 DVSS.n4431 0.0380882
R46384 DVSS.n7998 DVSS.n4431 0.0380882
R46385 DVSS.n7998 DVSS.n7994 0.0380882
R46386 DVSS.n7994 DVSS.n7993 0.0380882
R46387 DVSS.n7993 DVSS.n4433 0.0380882
R46388 DVSS.n7986 DVSS.n4433 0.0380882
R46389 DVSS.n7986 DVSS.n7982 0.0380882
R46390 DVSS.n7982 DVSS.n7981 0.0380882
R46391 DVSS.n7981 DVSS.n4435 0.0380882
R46392 DVSS.n7974 DVSS.n4435 0.0380882
R46393 DVSS.n7974 DVSS.n7970 0.0380882
R46394 DVSS.n7970 DVSS.n7969 0.0380882
R46395 DVSS.n7969 DVSS.n4437 0.0380882
R46396 DVSS.n7962 DVSS.n4437 0.0380882
R46397 DVSS.n7962 DVSS.n7958 0.0380882
R46398 DVSS.n7958 DVSS.n7957 0.0380882
R46399 DVSS.n7957 DVSS.n4439 0.0380882
R46400 DVSS.n7950 DVSS.n4439 0.0380882
R46401 DVSS.n7950 DVSS.n7946 0.0380882
R46402 DVSS.n7946 DVSS.n7945 0.0380882
R46403 DVSS.n7945 DVSS.n4441 0.0380882
R46404 DVSS.n7938 DVSS.n4441 0.0380882
R46405 DVSS.n7938 DVSS.n7934 0.0380882
R46406 DVSS.n7934 DVSS.n7933 0.0380882
R46407 DVSS.n7933 DVSS.n4443 0.0380882
R46408 DVSS.n7926 DVSS.n4443 0.0380882
R46409 DVSS.n7926 DVSS.n7922 0.0380882
R46410 DVSS.n7922 DVSS.n7921 0.0380882
R46411 DVSS.n7921 DVSS.n4445 0.0380882
R46412 DVSS.n7914 DVSS.n4445 0.0380882
R46413 DVSS.n7914 DVSS.n7910 0.0380882
R46414 DVSS.n7910 DVSS.n7909 0.0380882
R46415 DVSS.n7909 DVSS.n4447 0.0380882
R46416 DVSS.n7902 DVSS.n4447 0.0380882
R46417 DVSS.n7902 DVSS.n7898 0.0380882
R46418 DVSS.n7898 DVSS.n7897 0.0380882
R46419 DVSS.n7897 DVSS.n4449 0.0380882
R46420 DVSS.n7890 DVSS.n4449 0.0380882
R46421 DVSS.n7890 DVSS.n7886 0.0380882
R46422 DVSS.n7886 DVSS.n7885 0.0380882
R46423 DVSS.n7885 DVSS.n4451 0.0380882
R46424 DVSS.n7878 DVSS.n4451 0.0380882
R46425 DVSS.n7878 DVSS.n7874 0.0380882
R46426 DVSS.n7874 DVSS.n7873 0.0380882
R46427 DVSS.n7873 DVSS.n4453 0.0380882
R46428 DVSS.n7866 DVSS.n4453 0.0380882
R46429 DVSS.n7866 DVSS.n7862 0.0380882
R46430 DVSS.n7862 DVSS.n7861 0.0380882
R46431 DVSS.n7861 DVSS.n4455 0.0380882
R46432 DVSS.n7854 DVSS.n4455 0.0380882
R46433 DVSS.n7854 DVSS.n7850 0.0380882
R46434 DVSS.n7850 DVSS.n7849 0.0380882
R46435 DVSS.n7849 DVSS.n4457 0.0380882
R46436 DVSS.n7842 DVSS.n4457 0.0380882
R46437 DVSS.n4106 DVSS.n4017 0.0380882
R46438 DVSS.n4117 DVSS.n4106 0.0380882
R46439 DVSS.n4118 DVSS.n4117 0.0380882
R46440 DVSS.n4119 DVSS.n4118 0.0380882
R46441 DVSS.n4119 DVSS.n4102 0.0380882
R46442 DVSS.n4129 DVSS.n4102 0.0380882
R46443 DVSS.n4130 DVSS.n4129 0.0380882
R46444 DVSS.n4131 DVSS.n4130 0.0380882
R46445 DVSS.n4131 DVSS.n4098 0.0380882
R46446 DVSS.n4141 DVSS.n4098 0.0380882
R46447 DVSS.n4142 DVSS.n4141 0.0380882
R46448 DVSS.n4143 DVSS.n4142 0.0380882
R46449 DVSS.n4143 DVSS.n4094 0.0380882
R46450 DVSS.n4153 DVSS.n4094 0.0380882
R46451 DVSS.n4154 DVSS.n4153 0.0380882
R46452 DVSS.n4155 DVSS.n4154 0.0380882
R46453 DVSS.n4155 DVSS.n4090 0.0380882
R46454 DVSS.n4165 DVSS.n4090 0.0380882
R46455 DVSS.n4166 DVSS.n4165 0.0380882
R46456 DVSS.n4167 DVSS.n4166 0.0380882
R46457 DVSS.n4167 DVSS.n4086 0.0380882
R46458 DVSS.n4177 DVSS.n4086 0.0380882
R46459 DVSS.n4178 DVSS.n4177 0.0380882
R46460 DVSS.n4179 DVSS.n4178 0.0380882
R46461 DVSS.n4179 DVSS.n4082 0.0380882
R46462 DVSS.n4189 DVSS.n4082 0.0380882
R46463 DVSS.n4190 DVSS.n4189 0.0380882
R46464 DVSS.n4191 DVSS.n4190 0.0380882
R46465 DVSS.n4191 DVSS.n4078 0.0380882
R46466 DVSS.n4201 DVSS.n4078 0.0380882
R46467 DVSS.n4202 DVSS.n4201 0.0380882
R46468 DVSS.n4203 DVSS.n4202 0.0380882
R46469 DVSS.n4203 DVSS.n4074 0.0380882
R46470 DVSS.n4213 DVSS.n4074 0.0380882
R46471 DVSS.n4214 DVSS.n4213 0.0380882
R46472 DVSS.n4215 DVSS.n4214 0.0380882
R46473 DVSS.n4215 DVSS.n4070 0.0380882
R46474 DVSS.n4225 DVSS.n4070 0.0380882
R46475 DVSS.n4226 DVSS.n4225 0.0380882
R46476 DVSS.n4227 DVSS.n4226 0.0380882
R46477 DVSS.n4227 DVSS.n4066 0.0380882
R46478 DVSS.n4237 DVSS.n4066 0.0380882
R46479 DVSS.n4238 DVSS.n4237 0.0380882
R46480 DVSS.n4239 DVSS.n4238 0.0380882
R46481 DVSS.n4239 DVSS.n4062 0.0380882
R46482 DVSS.n4249 DVSS.n4062 0.0380882
R46483 DVSS.n4250 DVSS.n4249 0.0380882
R46484 DVSS.n4251 DVSS.n4250 0.0380882
R46485 DVSS.n4251 DVSS.n4058 0.0380882
R46486 DVSS.n4261 DVSS.n4058 0.0380882
R46487 DVSS.n4262 DVSS.n4261 0.0380882
R46488 DVSS.n4263 DVSS.n4262 0.0380882
R46489 DVSS.n4263 DVSS.n4054 0.0380882
R46490 DVSS.n4273 DVSS.n4054 0.0380882
R46491 DVSS.n4274 DVSS.n4273 0.0380882
R46492 DVSS.n4275 DVSS.n4274 0.0380882
R46493 DVSS.n4275 DVSS.n4050 0.0380882
R46494 DVSS.n4285 DVSS.n4050 0.0380882
R46495 DVSS.n4286 DVSS.n4285 0.0380882
R46496 DVSS.n4287 DVSS.n4286 0.0380882
R46497 DVSS.n4287 DVSS.n4046 0.0380882
R46498 DVSS.n4297 DVSS.n4046 0.0380882
R46499 DVSS.n4298 DVSS.n4297 0.0380882
R46500 DVSS.n4299 DVSS.n4298 0.0380882
R46501 DVSS.n4299 DVSS.n4042 0.0380882
R46502 DVSS.n4309 DVSS.n4042 0.0380882
R46503 DVSS.n4310 DVSS.n4309 0.0380882
R46504 DVSS.n4311 DVSS.n4310 0.0380882
R46505 DVSS.n4311 DVSS.n4038 0.0380882
R46506 DVSS.n4321 DVSS.n4038 0.0380882
R46507 DVSS.n4322 DVSS.n4321 0.0380882
R46508 DVSS.n4323 DVSS.n4322 0.0380882
R46509 DVSS.n4323 DVSS.n4034 0.0380882
R46510 DVSS.n4333 DVSS.n4034 0.0380882
R46511 DVSS.n4334 DVSS.n4333 0.0380882
R46512 DVSS.n4335 DVSS.n4334 0.0380882
R46513 DVSS.n4335 DVSS.n4030 0.0380882
R46514 DVSS.n4345 DVSS.n4030 0.0380882
R46515 DVSS.n4346 DVSS.n4345 0.0380882
R46516 DVSS.n4348 DVSS.n4346 0.0380882
R46517 DVSS.n4348 DVSS.n4347 0.0380882
R46518 DVSS.n4347 DVSS.n4025 0.0380882
R46519 DVSS.n4358 DVSS.n4025 0.0380882
R46520 DVSS.n4108 DVSS.n4107 0.0380882
R46521 DVSS.n4116 DVSS.n4107 0.0380882
R46522 DVSS.n4116 DVSS.n4105 0.0380882
R46523 DVSS.n4120 DVSS.n4105 0.0380882
R46524 DVSS.n4120 DVSS.n4103 0.0380882
R46525 DVSS.n4128 DVSS.n4103 0.0380882
R46526 DVSS.n4128 DVSS.n4101 0.0380882
R46527 DVSS.n4132 DVSS.n4101 0.0380882
R46528 DVSS.n4132 DVSS.n4099 0.0380882
R46529 DVSS.n4140 DVSS.n4099 0.0380882
R46530 DVSS.n4140 DVSS.n4097 0.0380882
R46531 DVSS.n4144 DVSS.n4097 0.0380882
R46532 DVSS.n4144 DVSS.n4095 0.0380882
R46533 DVSS.n4152 DVSS.n4095 0.0380882
R46534 DVSS.n4152 DVSS.n4093 0.0380882
R46535 DVSS.n4156 DVSS.n4093 0.0380882
R46536 DVSS.n4156 DVSS.n4091 0.0380882
R46537 DVSS.n4164 DVSS.n4091 0.0380882
R46538 DVSS.n4164 DVSS.n4089 0.0380882
R46539 DVSS.n4168 DVSS.n4089 0.0380882
R46540 DVSS.n4168 DVSS.n4087 0.0380882
R46541 DVSS.n4176 DVSS.n4087 0.0380882
R46542 DVSS.n4176 DVSS.n4085 0.0380882
R46543 DVSS.n4180 DVSS.n4085 0.0380882
R46544 DVSS.n4180 DVSS.n4083 0.0380882
R46545 DVSS.n4188 DVSS.n4083 0.0380882
R46546 DVSS.n4188 DVSS.n4081 0.0380882
R46547 DVSS.n4192 DVSS.n4081 0.0380882
R46548 DVSS.n4192 DVSS.n4079 0.0380882
R46549 DVSS.n4200 DVSS.n4079 0.0380882
R46550 DVSS.n4200 DVSS.n4077 0.0380882
R46551 DVSS.n4204 DVSS.n4077 0.0380882
R46552 DVSS.n4204 DVSS.n4075 0.0380882
R46553 DVSS.n4212 DVSS.n4075 0.0380882
R46554 DVSS.n4212 DVSS.n4073 0.0380882
R46555 DVSS.n4216 DVSS.n4073 0.0380882
R46556 DVSS.n4216 DVSS.n4071 0.0380882
R46557 DVSS.n4224 DVSS.n4071 0.0380882
R46558 DVSS.n4224 DVSS.n4069 0.0380882
R46559 DVSS.n4228 DVSS.n4069 0.0380882
R46560 DVSS.n4228 DVSS.n4067 0.0380882
R46561 DVSS.n4236 DVSS.n4067 0.0380882
R46562 DVSS.n4236 DVSS.n4065 0.0380882
R46563 DVSS.n4240 DVSS.n4065 0.0380882
R46564 DVSS.n4240 DVSS.n4063 0.0380882
R46565 DVSS.n4248 DVSS.n4063 0.0380882
R46566 DVSS.n4248 DVSS.n4061 0.0380882
R46567 DVSS.n4252 DVSS.n4061 0.0380882
R46568 DVSS.n4252 DVSS.n4059 0.0380882
R46569 DVSS.n4260 DVSS.n4059 0.0380882
R46570 DVSS.n4260 DVSS.n4057 0.0380882
R46571 DVSS.n4264 DVSS.n4057 0.0380882
R46572 DVSS.n4264 DVSS.n4055 0.0380882
R46573 DVSS.n4272 DVSS.n4055 0.0380882
R46574 DVSS.n4272 DVSS.n4053 0.0380882
R46575 DVSS.n4276 DVSS.n4053 0.0380882
R46576 DVSS.n4276 DVSS.n4051 0.0380882
R46577 DVSS.n4284 DVSS.n4051 0.0380882
R46578 DVSS.n4284 DVSS.n4049 0.0380882
R46579 DVSS.n4288 DVSS.n4049 0.0380882
R46580 DVSS.n4288 DVSS.n4047 0.0380882
R46581 DVSS.n4296 DVSS.n4047 0.0380882
R46582 DVSS.n4296 DVSS.n4045 0.0380882
R46583 DVSS.n4300 DVSS.n4045 0.0380882
R46584 DVSS.n4300 DVSS.n4043 0.0380882
R46585 DVSS.n4308 DVSS.n4043 0.0380882
R46586 DVSS.n4308 DVSS.n4041 0.0380882
R46587 DVSS.n4312 DVSS.n4041 0.0380882
R46588 DVSS.n4312 DVSS.n4039 0.0380882
R46589 DVSS.n4320 DVSS.n4039 0.0380882
R46590 DVSS.n4320 DVSS.n4037 0.0380882
R46591 DVSS.n4324 DVSS.n4037 0.0380882
R46592 DVSS.n4324 DVSS.n4035 0.0380882
R46593 DVSS.n4332 DVSS.n4035 0.0380882
R46594 DVSS.n4332 DVSS.n4033 0.0380882
R46595 DVSS.n4336 DVSS.n4033 0.0380882
R46596 DVSS.n4336 DVSS.n4031 0.0380882
R46597 DVSS.n4344 DVSS.n4031 0.0380882
R46598 DVSS.n4344 DVSS.n4029 0.0380882
R46599 DVSS.n4349 DVSS.n4029 0.0380882
R46600 DVSS.n4349 DVSS.n4027 0.0380882
R46601 DVSS.n4027 DVSS.n4026 0.0380882
R46602 DVSS.n4357 DVSS.n4026 0.0380882
R46603 DVSS.n8131 DVSS.n8130 0.0380882
R46604 DVSS.n8132 DVSS.n8131 0.0380882
R46605 DVSS.n8132 DVSS.n4006 0.0380882
R46606 DVSS.n8139 DVSS.n4006 0.0380882
R46607 DVSS.n8140 DVSS.n8139 0.0380882
R46608 DVSS.n8141 DVSS.n8140 0.0380882
R46609 DVSS.n8141 DVSS.n4003 0.0380882
R46610 DVSS.n8148 DVSS.n4003 0.0380882
R46611 DVSS.n8149 DVSS.n8148 0.0380882
R46612 DVSS.n8150 DVSS.n8149 0.0380882
R46613 DVSS.n8150 DVSS.n4000 0.0380882
R46614 DVSS.n8157 DVSS.n4000 0.0380882
R46615 DVSS.n8158 DVSS.n8157 0.0380882
R46616 DVSS.n8159 DVSS.n8158 0.0380882
R46617 DVSS.n8159 DVSS.n3997 0.0380882
R46618 DVSS.n8166 DVSS.n3997 0.0380882
R46619 DVSS.n8167 DVSS.n8166 0.0380882
R46620 DVSS.n8168 DVSS.n8167 0.0380882
R46621 DVSS.n8168 DVSS.n3994 0.0380882
R46622 DVSS.n8175 DVSS.n3994 0.0380882
R46623 DVSS.n8176 DVSS.n8175 0.0380882
R46624 DVSS.n8177 DVSS.n8176 0.0380882
R46625 DVSS.n8177 DVSS.n3991 0.0380882
R46626 DVSS.n8184 DVSS.n3991 0.0380882
R46627 DVSS.n8185 DVSS.n8184 0.0380882
R46628 DVSS.n8186 DVSS.n8185 0.0380882
R46629 DVSS.n8186 DVSS.n3988 0.0380882
R46630 DVSS.n8193 DVSS.n3988 0.0380882
R46631 DVSS.n8194 DVSS.n8193 0.0380882
R46632 DVSS.n8195 DVSS.n8194 0.0380882
R46633 DVSS.n8195 DVSS.n3985 0.0380882
R46634 DVSS.n8202 DVSS.n3985 0.0380882
R46635 DVSS.n8203 DVSS.n8202 0.0380882
R46636 DVSS.n8204 DVSS.n8203 0.0380882
R46637 DVSS.n8204 DVSS.n3982 0.0380882
R46638 DVSS.n8211 DVSS.n3982 0.0380882
R46639 DVSS.n8212 DVSS.n8211 0.0380882
R46640 DVSS.n8213 DVSS.n8212 0.0380882
R46641 DVSS.n8213 DVSS.n3979 0.0380882
R46642 DVSS.n8220 DVSS.n3979 0.0380882
R46643 DVSS.n8221 DVSS.n8220 0.0380882
R46644 DVSS.n8222 DVSS.n8221 0.0380882
R46645 DVSS.n8222 DVSS.n3976 0.0380882
R46646 DVSS.n8229 DVSS.n3976 0.0380882
R46647 DVSS.n8230 DVSS.n8229 0.0380882
R46648 DVSS.n8231 DVSS.n8230 0.0380882
R46649 DVSS.n8231 DVSS.n3973 0.0380882
R46650 DVSS.n8238 DVSS.n3973 0.0380882
R46651 DVSS.n8239 DVSS.n8238 0.0380882
R46652 DVSS.n8240 DVSS.n8239 0.0380882
R46653 DVSS.n8240 DVSS.n3970 0.0380882
R46654 DVSS.n8247 DVSS.n3970 0.0380882
R46655 DVSS.n8248 DVSS.n8247 0.0380882
R46656 DVSS.n8249 DVSS.n8248 0.0380882
R46657 DVSS.n8249 DVSS.n3967 0.0380882
R46658 DVSS.n8256 DVSS.n3967 0.0380882
R46659 DVSS.n8257 DVSS.n8256 0.0380882
R46660 DVSS.n8258 DVSS.n8257 0.0380882
R46661 DVSS.n8258 DVSS.n3964 0.0380882
R46662 DVSS.n8265 DVSS.n3964 0.0380882
R46663 DVSS.n8266 DVSS.n8265 0.0380882
R46664 DVSS.n8267 DVSS.n8266 0.0380882
R46665 DVSS.n8267 DVSS.n3961 0.0380882
R46666 DVSS.n8274 DVSS.n3961 0.0380882
R46667 DVSS.n8275 DVSS.n8274 0.0380882
R46668 DVSS.n8276 DVSS.n8275 0.0380882
R46669 DVSS.n8276 DVSS.n3958 0.0380882
R46670 DVSS.n8283 DVSS.n3958 0.0380882
R46671 DVSS.n8284 DVSS.n8283 0.0380882
R46672 DVSS.n8285 DVSS.n8284 0.0380882
R46673 DVSS.n8285 DVSS.n3955 0.0380882
R46674 DVSS.n8292 DVSS.n3955 0.0380882
R46675 DVSS.n8293 DVSS.n8292 0.0380882
R46676 DVSS.n8294 DVSS.n8293 0.0380882
R46677 DVSS.n8294 DVSS.n3952 0.0380882
R46678 DVSS.n8301 DVSS.n3952 0.0380882
R46679 DVSS.n8302 DVSS.n8301 0.0380882
R46680 DVSS.n8303 DVSS.n8302 0.0380882
R46681 DVSS.n8303 DVSS.n3949 0.0380882
R46682 DVSS.n8310 DVSS.n3949 0.0380882
R46683 DVSS.n8311 DVSS.n8310 0.0380882
R46684 DVSS.n8312 DVSS.n8311 0.0380882
R46685 DVSS.n8312 DVSS.n3852 0.0380882
R46686 DVSS.n4007 DVSS.n3903 0.0380882
R46687 DVSS.n8134 DVSS.n4007 0.0380882
R46688 DVSS.n8136 DVSS.n8134 0.0380882
R46689 DVSS.n8138 DVSS.n8136 0.0380882
R46690 DVSS.n8138 DVSS.n4005 0.0380882
R46691 DVSS.n8143 DVSS.n4005 0.0380882
R46692 DVSS.n8145 DVSS.n8143 0.0380882
R46693 DVSS.n8147 DVSS.n8145 0.0380882
R46694 DVSS.n8147 DVSS.n4002 0.0380882
R46695 DVSS.n8152 DVSS.n4002 0.0380882
R46696 DVSS.n8154 DVSS.n8152 0.0380882
R46697 DVSS.n8156 DVSS.n8154 0.0380882
R46698 DVSS.n8156 DVSS.n3999 0.0380882
R46699 DVSS.n8161 DVSS.n3999 0.0380882
R46700 DVSS.n8163 DVSS.n8161 0.0380882
R46701 DVSS.n8165 DVSS.n8163 0.0380882
R46702 DVSS.n8165 DVSS.n3996 0.0380882
R46703 DVSS.n8170 DVSS.n3996 0.0380882
R46704 DVSS.n8172 DVSS.n8170 0.0380882
R46705 DVSS.n8174 DVSS.n8172 0.0380882
R46706 DVSS.n8174 DVSS.n3993 0.0380882
R46707 DVSS.n8179 DVSS.n3993 0.0380882
R46708 DVSS.n8181 DVSS.n8179 0.0380882
R46709 DVSS.n8183 DVSS.n8181 0.0380882
R46710 DVSS.n8183 DVSS.n3990 0.0380882
R46711 DVSS.n8188 DVSS.n3990 0.0380882
R46712 DVSS.n8190 DVSS.n8188 0.0380882
R46713 DVSS.n8192 DVSS.n8190 0.0380882
R46714 DVSS.n8192 DVSS.n3987 0.0380882
R46715 DVSS.n8197 DVSS.n3987 0.0380882
R46716 DVSS.n8199 DVSS.n8197 0.0380882
R46717 DVSS.n8201 DVSS.n8199 0.0380882
R46718 DVSS.n8201 DVSS.n3984 0.0380882
R46719 DVSS.n8206 DVSS.n3984 0.0380882
R46720 DVSS.n8208 DVSS.n8206 0.0380882
R46721 DVSS.n8210 DVSS.n8208 0.0380882
R46722 DVSS.n8210 DVSS.n3981 0.0380882
R46723 DVSS.n8215 DVSS.n3981 0.0380882
R46724 DVSS.n8217 DVSS.n8215 0.0380882
R46725 DVSS.n8219 DVSS.n8217 0.0380882
R46726 DVSS.n8219 DVSS.n3978 0.0380882
R46727 DVSS.n8224 DVSS.n3978 0.0380882
R46728 DVSS.n8226 DVSS.n8224 0.0380882
R46729 DVSS.n8228 DVSS.n8226 0.0380882
R46730 DVSS.n8228 DVSS.n3975 0.0380882
R46731 DVSS.n8233 DVSS.n3975 0.0380882
R46732 DVSS.n8235 DVSS.n8233 0.0380882
R46733 DVSS.n8237 DVSS.n8235 0.0380882
R46734 DVSS.n8237 DVSS.n3972 0.0380882
R46735 DVSS.n8242 DVSS.n3972 0.0380882
R46736 DVSS.n8244 DVSS.n8242 0.0380882
R46737 DVSS.n8246 DVSS.n8244 0.0380882
R46738 DVSS.n8246 DVSS.n3969 0.0380882
R46739 DVSS.n8251 DVSS.n3969 0.0380882
R46740 DVSS.n8253 DVSS.n8251 0.0380882
R46741 DVSS.n8255 DVSS.n8253 0.0380882
R46742 DVSS.n8255 DVSS.n3966 0.0380882
R46743 DVSS.n8260 DVSS.n3966 0.0380882
R46744 DVSS.n8262 DVSS.n8260 0.0380882
R46745 DVSS.n8264 DVSS.n8262 0.0380882
R46746 DVSS.n8264 DVSS.n3963 0.0380882
R46747 DVSS.n8269 DVSS.n3963 0.0380882
R46748 DVSS.n8271 DVSS.n8269 0.0380882
R46749 DVSS.n8273 DVSS.n8271 0.0380882
R46750 DVSS.n8273 DVSS.n3960 0.0380882
R46751 DVSS.n8278 DVSS.n3960 0.0380882
R46752 DVSS.n8280 DVSS.n8278 0.0380882
R46753 DVSS.n8282 DVSS.n8280 0.0380882
R46754 DVSS.n8282 DVSS.n3957 0.0380882
R46755 DVSS.n8287 DVSS.n3957 0.0380882
R46756 DVSS.n8289 DVSS.n8287 0.0380882
R46757 DVSS.n8291 DVSS.n8289 0.0380882
R46758 DVSS.n8291 DVSS.n3954 0.0380882
R46759 DVSS.n8296 DVSS.n3954 0.0380882
R46760 DVSS.n8298 DVSS.n8296 0.0380882
R46761 DVSS.n8300 DVSS.n8298 0.0380882
R46762 DVSS.n8300 DVSS.n3951 0.0380882
R46763 DVSS.n8305 DVSS.n3951 0.0380882
R46764 DVSS.n8307 DVSS.n8305 0.0380882
R46765 DVSS.n8309 DVSS.n8307 0.0380882
R46766 DVSS.n8309 DVSS.n3948 0.0380882
R46767 DVSS.n8314 DVSS.n3948 0.0380882
R46768 DVSS.n8315 DVSS.n8314 0.0380882
R46769 DVSS.n8341 DVSS.n8340 0.0380882
R46770 DVSS.n8342 DVSS.n8341 0.0380882
R46771 DVSS.n8342 DVSS.n3839 0.0380882
R46772 DVSS.n8352 DVSS.n3839 0.0380882
R46773 DVSS.n8353 DVSS.n8352 0.0380882
R46774 DVSS.n8354 DVSS.n8353 0.0380882
R46775 DVSS.n8354 DVSS.n3837 0.0380882
R46776 DVSS.n8364 DVSS.n3837 0.0380882
R46777 DVSS.n8365 DVSS.n8364 0.0380882
R46778 DVSS.n8366 DVSS.n8365 0.0380882
R46779 DVSS.n8366 DVSS.n3835 0.0380882
R46780 DVSS.n8376 DVSS.n3835 0.0380882
R46781 DVSS.n8377 DVSS.n8376 0.0380882
R46782 DVSS.n8378 DVSS.n8377 0.0380882
R46783 DVSS.n8378 DVSS.n3833 0.0380882
R46784 DVSS.n8388 DVSS.n3833 0.0380882
R46785 DVSS.n8389 DVSS.n8388 0.0380882
R46786 DVSS.n8390 DVSS.n8389 0.0380882
R46787 DVSS.n8390 DVSS.n3831 0.0380882
R46788 DVSS.n8400 DVSS.n3831 0.0380882
R46789 DVSS.n8401 DVSS.n8400 0.0380882
R46790 DVSS.n8402 DVSS.n8401 0.0380882
R46791 DVSS.n8402 DVSS.n3829 0.0380882
R46792 DVSS.n8412 DVSS.n3829 0.0380882
R46793 DVSS.n8413 DVSS.n8412 0.0380882
R46794 DVSS.n8414 DVSS.n8413 0.0380882
R46795 DVSS.n8414 DVSS.n3827 0.0380882
R46796 DVSS.n8424 DVSS.n3827 0.0380882
R46797 DVSS.n8425 DVSS.n8424 0.0380882
R46798 DVSS.n8426 DVSS.n8425 0.0380882
R46799 DVSS.n8426 DVSS.n3825 0.0380882
R46800 DVSS.n8436 DVSS.n3825 0.0380882
R46801 DVSS.n8437 DVSS.n8436 0.0380882
R46802 DVSS.n8438 DVSS.n8437 0.0380882
R46803 DVSS.n8438 DVSS.n3823 0.0380882
R46804 DVSS.n8448 DVSS.n3823 0.0380882
R46805 DVSS.n8449 DVSS.n8448 0.0380882
R46806 DVSS.n8450 DVSS.n8449 0.0380882
R46807 DVSS.n8450 DVSS.n3821 0.0380882
R46808 DVSS.n8460 DVSS.n3821 0.0380882
R46809 DVSS.n8461 DVSS.n8460 0.0380882
R46810 DVSS.n8462 DVSS.n8461 0.0380882
R46811 DVSS.n8462 DVSS.n3819 0.0380882
R46812 DVSS.n8472 DVSS.n3819 0.0380882
R46813 DVSS.n8473 DVSS.n8472 0.0380882
R46814 DVSS.n8474 DVSS.n8473 0.0380882
R46815 DVSS.n8474 DVSS.n3817 0.0380882
R46816 DVSS.n8484 DVSS.n3817 0.0380882
R46817 DVSS.n8485 DVSS.n8484 0.0380882
R46818 DVSS.n8486 DVSS.n8485 0.0380882
R46819 DVSS.n8486 DVSS.n3815 0.0380882
R46820 DVSS.n8496 DVSS.n3815 0.0380882
R46821 DVSS.n8497 DVSS.n8496 0.0380882
R46822 DVSS.n8498 DVSS.n8497 0.0380882
R46823 DVSS.n8498 DVSS.n3813 0.0380882
R46824 DVSS.n8508 DVSS.n3813 0.0380882
R46825 DVSS.n8509 DVSS.n8508 0.0380882
R46826 DVSS.n8510 DVSS.n8509 0.0380882
R46827 DVSS.n8510 DVSS.n3811 0.0380882
R46828 DVSS.n8520 DVSS.n3811 0.0380882
R46829 DVSS.n8521 DVSS.n8520 0.0380882
R46830 DVSS.n8522 DVSS.n8521 0.0380882
R46831 DVSS.n8522 DVSS.n3809 0.0380882
R46832 DVSS.n8532 DVSS.n3809 0.0380882
R46833 DVSS.n8533 DVSS.n8532 0.0380882
R46834 DVSS.n8534 DVSS.n8533 0.0380882
R46835 DVSS.n8534 DVSS.n3807 0.0380882
R46836 DVSS.n8544 DVSS.n3807 0.0380882
R46837 DVSS.n8545 DVSS.n8544 0.0380882
R46838 DVSS.n8546 DVSS.n8545 0.0380882
R46839 DVSS.n8546 DVSS.n3805 0.0380882
R46840 DVSS.n8556 DVSS.n3805 0.0380882
R46841 DVSS.n8557 DVSS.n8556 0.0380882
R46842 DVSS.n8558 DVSS.n8557 0.0380882
R46843 DVSS.n8558 DVSS.n3803 0.0380882
R46844 DVSS.n8568 DVSS.n3803 0.0380882
R46845 DVSS.n8569 DVSS.n8568 0.0380882
R46846 DVSS.n8570 DVSS.n8569 0.0380882
R46847 DVSS.n8570 DVSS.n3801 0.0380882
R46848 DVSS.n8580 DVSS.n3801 0.0380882
R46849 DVSS.n8581 DVSS.n8580 0.0380882
R46850 DVSS.n8583 DVSS.n8581 0.0380882
R46851 DVSS.n8583 DVSS.n8582 0.0380882
R46852 DVSS.n8339 DVSS.n3842 0.0380882
R46853 DVSS.n8343 DVSS.n3842 0.0380882
R46854 DVSS.n8347 DVSS.n8343 0.0380882
R46855 DVSS.n8351 DVSS.n8347 0.0380882
R46856 DVSS.n8351 DVSS.n3838 0.0380882
R46857 DVSS.n8355 DVSS.n3838 0.0380882
R46858 DVSS.n8359 DVSS.n8355 0.0380882
R46859 DVSS.n8363 DVSS.n8359 0.0380882
R46860 DVSS.n8363 DVSS.n3836 0.0380882
R46861 DVSS.n8367 DVSS.n3836 0.0380882
R46862 DVSS.n8371 DVSS.n8367 0.0380882
R46863 DVSS.n8375 DVSS.n8371 0.0380882
R46864 DVSS.n8375 DVSS.n3834 0.0380882
R46865 DVSS.n8379 DVSS.n3834 0.0380882
R46866 DVSS.n8383 DVSS.n8379 0.0380882
R46867 DVSS.n8387 DVSS.n8383 0.0380882
R46868 DVSS.n8387 DVSS.n3832 0.0380882
R46869 DVSS.n8391 DVSS.n3832 0.0380882
R46870 DVSS.n8395 DVSS.n8391 0.0380882
R46871 DVSS.n8399 DVSS.n8395 0.0380882
R46872 DVSS.n8399 DVSS.n3830 0.0380882
R46873 DVSS.n8403 DVSS.n3830 0.0380882
R46874 DVSS.n8407 DVSS.n8403 0.0380882
R46875 DVSS.n8411 DVSS.n8407 0.0380882
R46876 DVSS.n8411 DVSS.n3828 0.0380882
R46877 DVSS.n8415 DVSS.n3828 0.0380882
R46878 DVSS.n8419 DVSS.n8415 0.0380882
R46879 DVSS.n8423 DVSS.n8419 0.0380882
R46880 DVSS.n8423 DVSS.n3826 0.0380882
R46881 DVSS.n8427 DVSS.n3826 0.0380882
R46882 DVSS.n8431 DVSS.n8427 0.0380882
R46883 DVSS.n8435 DVSS.n8431 0.0380882
R46884 DVSS.n8435 DVSS.n3824 0.0380882
R46885 DVSS.n8439 DVSS.n3824 0.0380882
R46886 DVSS.n8443 DVSS.n8439 0.0380882
R46887 DVSS.n8447 DVSS.n8443 0.0380882
R46888 DVSS.n8447 DVSS.n3822 0.0380882
R46889 DVSS.n8451 DVSS.n3822 0.0380882
R46890 DVSS.n8455 DVSS.n8451 0.0380882
R46891 DVSS.n8459 DVSS.n8455 0.0380882
R46892 DVSS.n8459 DVSS.n3820 0.0380882
R46893 DVSS.n8463 DVSS.n3820 0.0380882
R46894 DVSS.n8467 DVSS.n8463 0.0380882
R46895 DVSS.n8471 DVSS.n8467 0.0380882
R46896 DVSS.n8471 DVSS.n3818 0.0380882
R46897 DVSS.n8475 DVSS.n3818 0.0380882
R46898 DVSS.n8479 DVSS.n8475 0.0380882
R46899 DVSS.n8483 DVSS.n8479 0.0380882
R46900 DVSS.n8483 DVSS.n3816 0.0380882
R46901 DVSS.n8487 DVSS.n3816 0.0380882
R46902 DVSS.n8491 DVSS.n8487 0.0380882
R46903 DVSS.n8495 DVSS.n8491 0.0380882
R46904 DVSS.n8495 DVSS.n3814 0.0380882
R46905 DVSS.n8499 DVSS.n3814 0.0380882
R46906 DVSS.n8503 DVSS.n8499 0.0380882
R46907 DVSS.n8507 DVSS.n8503 0.0380882
R46908 DVSS.n8507 DVSS.n3812 0.0380882
R46909 DVSS.n8511 DVSS.n3812 0.0380882
R46910 DVSS.n8515 DVSS.n8511 0.0380882
R46911 DVSS.n8519 DVSS.n8515 0.0380882
R46912 DVSS.n8519 DVSS.n3810 0.0380882
R46913 DVSS.n8523 DVSS.n3810 0.0380882
R46914 DVSS.n8527 DVSS.n8523 0.0380882
R46915 DVSS.n8531 DVSS.n8527 0.0380882
R46916 DVSS.n8531 DVSS.n3808 0.0380882
R46917 DVSS.n8535 DVSS.n3808 0.0380882
R46918 DVSS.n8539 DVSS.n8535 0.0380882
R46919 DVSS.n8543 DVSS.n8539 0.0380882
R46920 DVSS.n8543 DVSS.n3806 0.0380882
R46921 DVSS.n8547 DVSS.n3806 0.0380882
R46922 DVSS.n8551 DVSS.n8547 0.0380882
R46923 DVSS.n8555 DVSS.n8551 0.0380882
R46924 DVSS.n8555 DVSS.n3804 0.0380882
R46925 DVSS.n8559 DVSS.n3804 0.0380882
R46926 DVSS.n8563 DVSS.n8559 0.0380882
R46927 DVSS.n8567 DVSS.n8563 0.0380882
R46928 DVSS.n8567 DVSS.n3802 0.0380882
R46929 DVSS.n8571 DVSS.n3802 0.0380882
R46930 DVSS.n8575 DVSS.n8571 0.0380882
R46931 DVSS.n8579 DVSS.n8575 0.0380882
R46932 DVSS.n8579 DVSS.n3800 0.0380882
R46933 DVSS.n8584 DVSS.n3800 0.0380882
R46934 DVSS.n8584 DVSS.n3798 0.0380882
R46935 DVSS.n3566 DVSS.n3409 0.0380882
R46936 DVSS.n3567 DVSS.n3566 0.0380882
R46937 DVSS.n3568 DVSS.n3567 0.0380882
R46938 DVSS.n3568 DVSS.n3562 0.0380882
R46939 DVSS.n3575 DVSS.n3562 0.0380882
R46940 DVSS.n3576 DVSS.n3575 0.0380882
R46941 DVSS.n3577 DVSS.n3576 0.0380882
R46942 DVSS.n3577 DVSS.n3559 0.0380882
R46943 DVSS.n3584 DVSS.n3559 0.0380882
R46944 DVSS.n3585 DVSS.n3584 0.0380882
R46945 DVSS.n3586 DVSS.n3585 0.0380882
R46946 DVSS.n3586 DVSS.n3556 0.0380882
R46947 DVSS.n3593 DVSS.n3556 0.0380882
R46948 DVSS.n3594 DVSS.n3593 0.0380882
R46949 DVSS.n3595 DVSS.n3594 0.0380882
R46950 DVSS.n3595 DVSS.n3553 0.0380882
R46951 DVSS.n3602 DVSS.n3553 0.0380882
R46952 DVSS.n3603 DVSS.n3602 0.0380882
R46953 DVSS.n3604 DVSS.n3603 0.0380882
R46954 DVSS.n3604 DVSS.n3550 0.0380882
R46955 DVSS.n3611 DVSS.n3550 0.0380882
R46956 DVSS.n3612 DVSS.n3611 0.0380882
R46957 DVSS.n3613 DVSS.n3612 0.0380882
R46958 DVSS.n3613 DVSS.n3547 0.0380882
R46959 DVSS.n3620 DVSS.n3547 0.0380882
R46960 DVSS.n3621 DVSS.n3620 0.0380882
R46961 DVSS.n3622 DVSS.n3621 0.0380882
R46962 DVSS.n3622 DVSS.n3544 0.0380882
R46963 DVSS.n3629 DVSS.n3544 0.0380882
R46964 DVSS.n3630 DVSS.n3629 0.0380882
R46965 DVSS.n3631 DVSS.n3630 0.0380882
R46966 DVSS.n3631 DVSS.n3541 0.0380882
R46967 DVSS.n3638 DVSS.n3541 0.0380882
R46968 DVSS.n3639 DVSS.n3638 0.0380882
R46969 DVSS.n3640 DVSS.n3639 0.0380882
R46970 DVSS.n3640 DVSS.n3538 0.0380882
R46971 DVSS.n3647 DVSS.n3538 0.0380882
R46972 DVSS.n3648 DVSS.n3647 0.0380882
R46973 DVSS.n3649 DVSS.n3648 0.0380882
R46974 DVSS.n3649 DVSS.n3535 0.0380882
R46975 DVSS.n3656 DVSS.n3535 0.0380882
R46976 DVSS.n3657 DVSS.n3656 0.0380882
R46977 DVSS.n3658 DVSS.n3657 0.0380882
R46978 DVSS.n3658 DVSS.n3532 0.0380882
R46979 DVSS.n3665 DVSS.n3532 0.0380882
R46980 DVSS.n3666 DVSS.n3665 0.0380882
R46981 DVSS.n3667 DVSS.n3666 0.0380882
R46982 DVSS.n3667 DVSS.n3529 0.0380882
R46983 DVSS.n3674 DVSS.n3529 0.0380882
R46984 DVSS.n3675 DVSS.n3674 0.0380882
R46985 DVSS.n3676 DVSS.n3675 0.0380882
R46986 DVSS.n3676 DVSS.n3526 0.0380882
R46987 DVSS.n3683 DVSS.n3526 0.0380882
R46988 DVSS.n3684 DVSS.n3683 0.0380882
R46989 DVSS.n3685 DVSS.n3684 0.0380882
R46990 DVSS.n3685 DVSS.n3523 0.0380882
R46991 DVSS.n3692 DVSS.n3523 0.0380882
R46992 DVSS.n3693 DVSS.n3692 0.0380882
R46993 DVSS.n3694 DVSS.n3693 0.0380882
R46994 DVSS.n3694 DVSS.n3520 0.0380882
R46995 DVSS.n3701 DVSS.n3520 0.0380882
R46996 DVSS.n3702 DVSS.n3701 0.0380882
R46997 DVSS.n3703 DVSS.n3702 0.0380882
R46998 DVSS.n3703 DVSS.n3517 0.0380882
R46999 DVSS.n3710 DVSS.n3517 0.0380882
R47000 DVSS.n3711 DVSS.n3710 0.0380882
R47001 DVSS.n3712 DVSS.n3711 0.0380882
R47002 DVSS.n3712 DVSS.n3514 0.0380882
R47003 DVSS.n3719 DVSS.n3514 0.0380882
R47004 DVSS.n3720 DVSS.n3719 0.0380882
R47005 DVSS.n3721 DVSS.n3720 0.0380882
R47006 DVSS.n3721 DVSS.n3511 0.0380882
R47007 DVSS.n3728 DVSS.n3511 0.0380882
R47008 DVSS.n3729 DVSS.n3728 0.0380882
R47009 DVSS.n3730 DVSS.n3729 0.0380882
R47010 DVSS.n3730 DVSS.n3508 0.0380882
R47011 DVSS.n3737 DVSS.n3508 0.0380882
R47012 DVSS.n3738 DVSS.n3737 0.0380882
R47013 DVSS.n3739 DVSS.n3738 0.0380882
R47014 DVSS.n3739 DVSS.n3505 0.0380882
R47015 DVSS.n3746 DVSS.n3505 0.0380882
R47016 DVSS.n3747 DVSS.n3746 0.0380882
R47017 DVSS.n3748 DVSS.n3747 0.0380882
R47018 DVSS.n3565 DVSS.n3459 0.0380882
R47019 DVSS.n3565 DVSS.n3564 0.0380882
R47020 DVSS.n3570 DVSS.n3564 0.0380882
R47021 DVSS.n3572 DVSS.n3570 0.0380882
R47022 DVSS.n3574 DVSS.n3572 0.0380882
R47023 DVSS.n3574 DVSS.n3561 0.0380882
R47024 DVSS.n3579 DVSS.n3561 0.0380882
R47025 DVSS.n3581 DVSS.n3579 0.0380882
R47026 DVSS.n3583 DVSS.n3581 0.0380882
R47027 DVSS.n3583 DVSS.n3558 0.0380882
R47028 DVSS.n3588 DVSS.n3558 0.0380882
R47029 DVSS.n3590 DVSS.n3588 0.0380882
R47030 DVSS.n3592 DVSS.n3590 0.0380882
R47031 DVSS.n3592 DVSS.n3555 0.0380882
R47032 DVSS.n3597 DVSS.n3555 0.0380882
R47033 DVSS.n3599 DVSS.n3597 0.0380882
R47034 DVSS.n3601 DVSS.n3599 0.0380882
R47035 DVSS.n3601 DVSS.n3552 0.0380882
R47036 DVSS.n3606 DVSS.n3552 0.0380882
R47037 DVSS.n3608 DVSS.n3606 0.0380882
R47038 DVSS.n3610 DVSS.n3608 0.0380882
R47039 DVSS.n3610 DVSS.n3549 0.0380882
R47040 DVSS.n3615 DVSS.n3549 0.0380882
R47041 DVSS.n3617 DVSS.n3615 0.0380882
R47042 DVSS.n3619 DVSS.n3617 0.0380882
R47043 DVSS.n3619 DVSS.n3546 0.0380882
R47044 DVSS.n3624 DVSS.n3546 0.0380882
R47045 DVSS.n3626 DVSS.n3624 0.0380882
R47046 DVSS.n3628 DVSS.n3626 0.0380882
R47047 DVSS.n3628 DVSS.n3543 0.0380882
R47048 DVSS.n3633 DVSS.n3543 0.0380882
R47049 DVSS.n3635 DVSS.n3633 0.0380882
R47050 DVSS.n3637 DVSS.n3635 0.0380882
R47051 DVSS.n3637 DVSS.n3540 0.0380882
R47052 DVSS.n3642 DVSS.n3540 0.0380882
R47053 DVSS.n3644 DVSS.n3642 0.0380882
R47054 DVSS.n3646 DVSS.n3644 0.0380882
R47055 DVSS.n3646 DVSS.n3537 0.0380882
R47056 DVSS.n3651 DVSS.n3537 0.0380882
R47057 DVSS.n3653 DVSS.n3651 0.0380882
R47058 DVSS.n3655 DVSS.n3653 0.0380882
R47059 DVSS.n3655 DVSS.n3534 0.0380882
R47060 DVSS.n3660 DVSS.n3534 0.0380882
R47061 DVSS.n3662 DVSS.n3660 0.0380882
R47062 DVSS.n3664 DVSS.n3662 0.0380882
R47063 DVSS.n3664 DVSS.n3531 0.0380882
R47064 DVSS.n3669 DVSS.n3531 0.0380882
R47065 DVSS.n3671 DVSS.n3669 0.0380882
R47066 DVSS.n3673 DVSS.n3671 0.0380882
R47067 DVSS.n3673 DVSS.n3528 0.0380882
R47068 DVSS.n3678 DVSS.n3528 0.0380882
R47069 DVSS.n3680 DVSS.n3678 0.0380882
R47070 DVSS.n3682 DVSS.n3680 0.0380882
R47071 DVSS.n3682 DVSS.n3525 0.0380882
R47072 DVSS.n3687 DVSS.n3525 0.0380882
R47073 DVSS.n3689 DVSS.n3687 0.0380882
R47074 DVSS.n3691 DVSS.n3689 0.0380882
R47075 DVSS.n3691 DVSS.n3522 0.0380882
R47076 DVSS.n3696 DVSS.n3522 0.0380882
R47077 DVSS.n3698 DVSS.n3696 0.0380882
R47078 DVSS.n3700 DVSS.n3698 0.0380882
R47079 DVSS.n3700 DVSS.n3519 0.0380882
R47080 DVSS.n3705 DVSS.n3519 0.0380882
R47081 DVSS.n3707 DVSS.n3705 0.0380882
R47082 DVSS.n3709 DVSS.n3707 0.0380882
R47083 DVSS.n3709 DVSS.n3516 0.0380882
R47084 DVSS.n3714 DVSS.n3516 0.0380882
R47085 DVSS.n3716 DVSS.n3714 0.0380882
R47086 DVSS.n3718 DVSS.n3716 0.0380882
R47087 DVSS.n3718 DVSS.n3513 0.0380882
R47088 DVSS.n3723 DVSS.n3513 0.0380882
R47089 DVSS.n3725 DVSS.n3723 0.0380882
R47090 DVSS.n3727 DVSS.n3725 0.0380882
R47091 DVSS.n3727 DVSS.n3510 0.0380882
R47092 DVSS.n3732 DVSS.n3510 0.0380882
R47093 DVSS.n3734 DVSS.n3732 0.0380882
R47094 DVSS.n3736 DVSS.n3734 0.0380882
R47095 DVSS.n3736 DVSS.n3507 0.0380882
R47096 DVSS.n3741 DVSS.n3507 0.0380882
R47097 DVSS.n3743 DVSS.n3741 0.0380882
R47098 DVSS.n3745 DVSS.n3743 0.0380882
R47099 DVSS.n3745 DVSS.n3504 0.0380882
R47100 DVSS.n8599 DVSS.n3504 0.0380882
R47101 DVSS.n3150 DVSS.n3062 0.0380882
R47102 DVSS.n3161 DVSS.n3150 0.0380882
R47103 DVSS.n3162 DVSS.n3161 0.0380882
R47104 DVSS.n3163 DVSS.n3162 0.0380882
R47105 DVSS.n3163 DVSS.n3146 0.0380882
R47106 DVSS.n3173 DVSS.n3146 0.0380882
R47107 DVSS.n3174 DVSS.n3173 0.0380882
R47108 DVSS.n3175 DVSS.n3174 0.0380882
R47109 DVSS.n3175 DVSS.n3142 0.0380882
R47110 DVSS.n3185 DVSS.n3142 0.0380882
R47111 DVSS.n3186 DVSS.n3185 0.0380882
R47112 DVSS.n3187 DVSS.n3186 0.0380882
R47113 DVSS.n3187 DVSS.n3138 0.0380882
R47114 DVSS.n3197 DVSS.n3138 0.0380882
R47115 DVSS.n3198 DVSS.n3197 0.0380882
R47116 DVSS.n3199 DVSS.n3198 0.0380882
R47117 DVSS.n3199 DVSS.n3134 0.0380882
R47118 DVSS.n3209 DVSS.n3134 0.0380882
R47119 DVSS.n3210 DVSS.n3209 0.0380882
R47120 DVSS.n3211 DVSS.n3210 0.0380882
R47121 DVSS.n3211 DVSS.n3130 0.0380882
R47122 DVSS.n3221 DVSS.n3130 0.0380882
R47123 DVSS.n3222 DVSS.n3221 0.0380882
R47124 DVSS.n3223 DVSS.n3222 0.0380882
R47125 DVSS.n3223 DVSS.n3126 0.0380882
R47126 DVSS.n3233 DVSS.n3126 0.0380882
R47127 DVSS.n3234 DVSS.n3233 0.0380882
R47128 DVSS.n3235 DVSS.n3234 0.0380882
R47129 DVSS.n3235 DVSS.n3122 0.0380882
R47130 DVSS.n3245 DVSS.n3122 0.0380882
R47131 DVSS.n3246 DVSS.n3245 0.0380882
R47132 DVSS.n3247 DVSS.n3246 0.0380882
R47133 DVSS.n3247 DVSS.n3118 0.0380882
R47134 DVSS.n3257 DVSS.n3118 0.0380882
R47135 DVSS.n3258 DVSS.n3257 0.0380882
R47136 DVSS.n3259 DVSS.n3258 0.0380882
R47137 DVSS.n3259 DVSS.n3114 0.0380882
R47138 DVSS.n3269 DVSS.n3114 0.0380882
R47139 DVSS.n3270 DVSS.n3269 0.0380882
R47140 DVSS.n3271 DVSS.n3270 0.0380882
R47141 DVSS.n3271 DVSS.n3110 0.0380882
R47142 DVSS.n3281 DVSS.n3110 0.0380882
R47143 DVSS.n3282 DVSS.n3281 0.0380882
R47144 DVSS.n3283 DVSS.n3282 0.0380882
R47145 DVSS.n3283 DVSS.n3106 0.0380882
R47146 DVSS.n3293 DVSS.n3106 0.0380882
R47147 DVSS.n3294 DVSS.n3293 0.0380882
R47148 DVSS.n3295 DVSS.n3294 0.0380882
R47149 DVSS.n3295 DVSS.n3102 0.0380882
R47150 DVSS.n3305 DVSS.n3102 0.0380882
R47151 DVSS.n3306 DVSS.n3305 0.0380882
R47152 DVSS.n3307 DVSS.n3306 0.0380882
R47153 DVSS.n3307 DVSS.n3098 0.0380882
R47154 DVSS.n3317 DVSS.n3098 0.0380882
R47155 DVSS.n3318 DVSS.n3317 0.0380882
R47156 DVSS.n3319 DVSS.n3318 0.0380882
R47157 DVSS.n3319 DVSS.n3094 0.0380882
R47158 DVSS.n3329 DVSS.n3094 0.0380882
R47159 DVSS.n3330 DVSS.n3329 0.0380882
R47160 DVSS.n3331 DVSS.n3330 0.0380882
R47161 DVSS.n3331 DVSS.n3090 0.0380882
R47162 DVSS.n3341 DVSS.n3090 0.0380882
R47163 DVSS.n3342 DVSS.n3341 0.0380882
R47164 DVSS.n3343 DVSS.n3342 0.0380882
R47165 DVSS.n3343 DVSS.n3086 0.0380882
R47166 DVSS.n3353 DVSS.n3086 0.0380882
R47167 DVSS.n3354 DVSS.n3353 0.0380882
R47168 DVSS.n3355 DVSS.n3354 0.0380882
R47169 DVSS.n3355 DVSS.n3082 0.0380882
R47170 DVSS.n3365 DVSS.n3082 0.0380882
R47171 DVSS.n3366 DVSS.n3365 0.0380882
R47172 DVSS.n3367 DVSS.n3366 0.0380882
R47173 DVSS.n3367 DVSS.n3078 0.0380882
R47174 DVSS.n3377 DVSS.n3078 0.0380882
R47175 DVSS.n3378 DVSS.n3377 0.0380882
R47176 DVSS.n3379 DVSS.n3378 0.0380882
R47177 DVSS.n3379 DVSS.n3074 0.0380882
R47178 DVSS.n3389 DVSS.n3074 0.0380882
R47179 DVSS.n3390 DVSS.n3389 0.0380882
R47180 DVSS.n3392 DVSS.n3390 0.0380882
R47181 DVSS.n3392 DVSS.n3391 0.0380882
R47182 DVSS.n3391 DVSS.n3069 0.0380882
R47183 DVSS.n3402 DVSS.n3069 0.0380882
R47184 DVSS.n3152 DVSS.n3151 0.0380882
R47185 DVSS.n3160 DVSS.n3151 0.0380882
R47186 DVSS.n3160 DVSS.n3149 0.0380882
R47187 DVSS.n3164 DVSS.n3149 0.0380882
R47188 DVSS.n3164 DVSS.n3147 0.0380882
R47189 DVSS.n3172 DVSS.n3147 0.0380882
R47190 DVSS.n3172 DVSS.n3145 0.0380882
R47191 DVSS.n3176 DVSS.n3145 0.0380882
R47192 DVSS.n3176 DVSS.n3143 0.0380882
R47193 DVSS.n3184 DVSS.n3143 0.0380882
R47194 DVSS.n3184 DVSS.n3141 0.0380882
R47195 DVSS.n3188 DVSS.n3141 0.0380882
R47196 DVSS.n3188 DVSS.n3139 0.0380882
R47197 DVSS.n3196 DVSS.n3139 0.0380882
R47198 DVSS.n3196 DVSS.n3137 0.0380882
R47199 DVSS.n3200 DVSS.n3137 0.0380882
R47200 DVSS.n3200 DVSS.n3135 0.0380882
R47201 DVSS.n3208 DVSS.n3135 0.0380882
R47202 DVSS.n3208 DVSS.n3133 0.0380882
R47203 DVSS.n3212 DVSS.n3133 0.0380882
R47204 DVSS.n3212 DVSS.n3131 0.0380882
R47205 DVSS.n3220 DVSS.n3131 0.0380882
R47206 DVSS.n3220 DVSS.n3129 0.0380882
R47207 DVSS.n3224 DVSS.n3129 0.0380882
R47208 DVSS.n3224 DVSS.n3127 0.0380882
R47209 DVSS.n3232 DVSS.n3127 0.0380882
R47210 DVSS.n3232 DVSS.n3125 0.0380882
R47211 DVSS.n3236 DVSS.n3125 0.0380882
R47212 DVSS.n3236 DVSS.n3123 0.0380882
R47213 DVSS.n3244 DVSS.n3123 0.0380882
R47214 DVSS.n3244 DVSS.n3121 0.0380882
R47215 DVSS.n3248 DVSS.n3121 0.0380882
R47216 DVSS.n3248 DVSS.n3119 0.0380882
R47217 DVSS.n3256 DVSS.n3119 0.0380882
R47218 DVSS.n3256 DVSS.n3117 0.0380882
R47219 DVSS.n3260 DVSS.n3117 0.0380882
R47220 DVSS.n3260 DVSS.n3115 0.0380882
R47221 DVSS.n3268 DVSS.n3115 0.0380882
R47222 DVSS.n3268 DVSS.n3113 0.0380882
R47223 DVSS.n3272 DVSS.n3113 0.0380882
R47224 DVSS.n3272 DVSS.n3111 0.0380882
R47225 DVSS.n3280 DVSS.n3111 0.0380882
R47226 DVSS.n3280 DVSS.n3109 0.0380882
R47227 DVSS.n3284 DVSS.n3109 0.0380882
R47228 DVSS.n3284 DVSS.n3107 0.0380882
R47229 DVSS.n3292 DVSS.n3107 0.0380882
R47230 DVSS.n3292 DVSS.n3105 0.0380882
R47231 DVSS.n3296 DVSS.n3105 0.0380882
R47232 DVSS.n3296 DVSS.n3103 0.0380882
R47233 DVSS.n3304 DVSS.n3103 0.0380882
R47234 DVSS.n3304 DVSS.n3101 0.0380882
R47235 DVSS.n3308 DVSS.n3101 0.0380882
R47236 DVSS.n3308 DVSS.n3099 0.0380882
R47237 DVSS.n3316 DVSS.n3099 0.0380882
R47238 DVSS.n3316 DVSS.n3097 0.0380882
R47239 DVSS.n3320 DVSS.n3097 0.0380882
R47240 DVSS.n3320 DVSS.n3095 0.0380882
R47241 DVSS.n3328 DVSS.n3095 0.0380882
R47242 DVSS.n3328 DVSS.n3093 0.0380882
R47243 DVSS.n3332 DVSS.n3093 0.0380882
R47244 DVSS.n3332 DVSS.n3091 0.0380882
R47245 DVSS.n3340 DVSS.n3091 0.0380882
R47246 DVSS.n3340 DVSS.n3089 0.0380882
R47247 DVSS.n3344 DVSS.n3089 0.0380882
R47248 DVSS.n3344 DVSS.n3087 0.0380882
R47249 DVSS.n3352 DVSS.n3087 0.0380882
R47250 DVSS.n3352 DVSS.n3085 0.0380882
R47251 DVSS.n3356 DVSS.n3085 0.0380882
R47252 DVSS.n3356 DVSS.n3083 0.0380882
R47253 DVSS.n3364 DVSS.n3083 0.0380882
R47254 DVSS.n3364 DVSS.n3081 0.0380882
R47255 DVSS.n3368 DVSS.n3081 0.0380882
R47256 DVSS.n3368 DVSS.n3079 0.0380882
R47257 DVSS.n3376 DVSS.n3079 0.0380882
R47258 DVSS.n3376 DVSS.n3077 0.0380882
R47259 DVSS.n3380 DVSS.n3077 0.0380882
R47260 DVSS.n3380 DVSS.n3075 0.0380882
R47261 DVSS.n3388 DVSS.n3075 0.0380882
R47262 DVSS.n3388 DVSS.n3073 0.0380882
R47263 DVSS.n3393 DVSS.n3073 0.0380882
R47264 DVSS.n3393 DVSS.n3071 0.0380882
R47265 DVSS.n3071 DVSS.n3070 0.0380882
R47266 DVSS.n3401 DVSS.n3070 0.0380882
R47267 DVSS.n8964 DVSS.n3048 0.0380882
R47268 DVSS.n8964 DVSS.n8963 0.0380882
R47269 DVSS.n8963 DVSS.n8962 0.0380882
R47270 DVSS.n8962 DVSS.n8681 0.0380882
R47271 DVSS.n8952 DVSS.n8681 0.0380882
R47272 DVSS.n8952 DVSS.n8951 0.0380882
R47273 DVSS.n8951 DVSS.n8950 0.0380882
R47274 DVSS.n8950 DVSS.n8683 0.0380882
R47275 DVSS.n8940 DVSS.n8683 0.0380882
R47276 DVSS.n8940 DVSS.n8939 0.0380882
R47277 DVSS.n8939 DVSS.n8938 0.0380882
R47278 DVSS.n8938 DVSS.n8685 0.0380882
R47279 DVSS.n8928 DVSS.n8685 0.0380882
R47280 DVSS.n8928 DVSS.n8927 0.0380882
R47281 DVSS.n8927 DVSS.n8926 0.0380882
R47282 DVSS.n8926 DVSS.n8687 0.0380882
R47283 DVSS.n8916 DVSS.n8687 0.0380882
R47284 DVSS.n8916 DVSS.n8915 0.0380882
R47285 DVSS.n8915 DVSS.n8914 0.0380882
R47286 DVSS.n8914 DVSS.n8689 0.0380882
R47287 DVSS.n8904 DVSS.n8689 0.0380882
R47288 DVSS.n8904 DVSS.n8903 0.0380882
R47289 DVSS.n8903 DVSS.n8902 0.0380882
R47290 DVSS.n8902 DVSS.n8691 0.0380882
R47291 DVSS.n8892 DVSS.n8691 0.0380882
R47292 DVSS.n8892 DVSS.n8891 0.0380882
R47293 DVSS.n8891 DVSS.n8890 0.0380882
R47294 DVSS.n8890 DVSS.n8693 0.0380882
R47295 DVSS.n8880 DVSS.n8693 0.0380882
R47296 DVSS.n8880 DVSS.n8879 0.0380882
R47297 DVSS.n8879 DVSS.n8878 0.0380882
R47298 DVSS.n8878 DVSS.n8695 0.0380882
R47299 DVSS.n8868 DVSS.n8695 0.0380882
R47300 DVSS.n8868 DVSS.n8867 0.0380882
R47301 DVSS.n8867 DVSS.n8866 0.0380882
R47302 DVSS.n8866 DVSS.n8697 0.0380882
R47303 DVSS.n8856 DVSS.n8697 0.0380882
R47304 DVSS.n8856 DVSS.n8855 0.0380882
R47305 DVSS.n8855 DVSS.n8854 0.0380882
R47306 DVSS.n8854 DVSS.n8699 0.0380882
R47307 DVSS.n8844 DVSS.n8699 0.0380882
R47308 DVSS.n8844 DVSS.n8843 0.0380882
R47309 DVSS.n8843 DVSS.n8842 0.0380882
R47310 DVSS.n8842 DVSS.n8701 0.0380882
R47311 DVSS.n8832 DVSS.n8701 0.0380882
R47312 DVSS.n8832 DVSS.n8831 0.0380882
R47313 DVSS.n8831 DVSS.n8830 0.0380882
R47314 DVSS.n8830 DVSS.n8703 0.0380882
R47315 DVSS.n8820 DVSS.n8703 0.0380882
R47316 DVSS.n8820 DVSS.n8819 0.0380882
R47317 DVSS.n8819 DVSS.n8818 0.0380882
R47318 DVSS.n8818 DVSS.n8705 0.0380882
R47319 DVSS.n8808 DVSS.n8705 0.0380882
R47320 DVSS.n8808 DVSS.n8807 0.0380882
R47321 DVSS.n8807 DVSS.n8806 0.0380882
R47322 DVSS.n8806 DVSS.n8707 0.0380882
R47323 DVSS.n8796 DVSS.n8707 0.0380882
R47324 DVSS.n8796 DVSS.n8795 0.0380882
R47325 DVSS.n8795 DVSS.n8794 0.0380882
R47326 DVSS.n8794 DVSS.n8709 0.0380882
R47327 DVSS.n8784 DVSS.n8709 0.0380882
R47328 DVSS.n8784 DVSS.n8783 0.0380882
R47329 DVSS.n8783 DVSS.n8782 0.0380882
R47330 DVSS.n8782 DVSS.n8711 0.0380882
R47331 DVSS.n8772 DVSS.n8711 0.0380882
R47332 DVSS.n8772 DVSS.n8771 0.0380882
R47333 DVSS.n8771 DVSS.n8770 0.0380882
R47334 DVSS.n8770 DVSS.n8713 0.0380882
R47335 DVSS.n8760 DVSS.n8713 0.0380882
R47336 DVSS.n8760 DVSS.n8759 0.0380882
R47337 DVSS.n8759 DVSS.n8758 0.0380882
R47338 DVSS.n8758 DVSS.n8715 0.0380882
R47339 DVSS.n8748 DVSS.n8715 0.0380882
R47340 DVSS.n8748 DVSS.n8747 0.0380882
R47341 DVSS.n8747 DVSS.n8746 0.0380882
R47342 DVSS.n8746 DVSS.n8717 0.0380882
R47343 DVSS.n8736 DVSS.n8717 0.0380882
R47344 DVSS.n8736 DVSS.n8735 0.0380882
R47345 DVSS.n8735 DVSS.n8734 0.0380882
R47346 DVSS.n8734 DVSS.n8719 0.0380882
R47347 DVSS.n8724 DVSS.n8719 0.0380882
R47348 DVSS.n8724 DVSS.n8723 0.0380882
R47349 DVSS.n8723 DVSS.n3055 0.0380882
R47350 DVSS.n8966 DVSS.n8965 0.0380882
R47351 DVSS.n8965 DVSS.n8680 0.0380882
R47352 DVSS.n8961 DVSS.n8680 0.0380882
R47353 DVSS.n8961 DVSS.n8957 0.0380882
R47354 DVSS.n8957 DVSS.n8956 0.0380882
R47355 DVSS.n8956 DVSS.n8682 0.0380882
R47356 DVSS.n8949 DVSS.n8682 0.0380882
R47357 DVSS.n8949 DVSS.n8945 0.0380882
R47358 DVSS.n8945 DVSS.n8944 0.0380882
R47359 DVSS.n8944 DVSS.n8684 0.0380882
R47360 DVSS.n8937 DVSS.n8684 0.0380882
R47361 DVSS.n8937 DVSS.n8933 0.0380882
R47362 DVSS.n8933 DVSS.n8932 0.0380882
R47363 DVSS.n8932 DVSS.n8686 0.0380882
R47364 DVSS.n8925 DVSS.n8686 0.0380882
R47365 DVSS.n8925 DVSS.n8921 0.0380882
R47366 DVSS.n8921 DVSS.n8920 0.0380882
R47367 DVSS.n8920 DVSS.n8688 0.0380882
R47368 DVSS.n8913 DVSS.n8688 0.0380882
R47369 DVSS.n8913 DVSS.n8909 0.0380882
R47370 DVSS.n8909 DVSS.n8908 0.0380882
R47371 DVSS.n8908 DVSS.n8690 0.0380882
R47372 DVSS.n8901 DVSS.n8690 0.0380882
R47373 DVSS.n8901 DVSS.n8897 0.0380882
R47374 DVSS.n8897 DVSS.n8896 0.0380882
R47375 DVSS.n8896 DVSS.n8692 0.0380882
R47376 DVSS.n8889 DVSS.n8692 0.0380882
R47377 DVSS.n8889 DVSS.n8885 0.0380882
R47378 DVSS.n8885 DVSS.n8884 0.0380882
R47379 DVSS.n8884 DVSS.n8694 0.0380882
R47380 DVSS.n8877 DVSS.n8694 0.0380882
R47381 DVSS.n8877 DVSS.n8873 0.0380882
R47382 DVSS.n8873 DVSS.n8872 0.0380882
R47383 DVSS.n8872 DVSS.n8696 0.0380882
R47384 DVSS.n8865 DVSS.n8696 0.0380882
R47385 DVSS.n8865 DVSS.n8861 0.0380882
R47386 DVSS.n8861 DVSS.n8860 0.0380882
R47387 DVSS.n8860 DVSS.n8698 0.0380882
R47388 DVSS.n8853 DVSS.n8698 0.0380882
R47389 DVSS.n8853 DVSS.n8849 0.0380882
R47390 DVSS.n8849 DVSS.n8848 0.0380882
R47391 DVSS.n8848 DVSS.n8700 0.0380882
R47392 DVSS.n8841 DVSS.n8700 0.0380882
R47393 DVSS.n8841 DVSS.n8837 0.0380882
R47394 DVSS.n8837 DVSS.n8836 0.0380882
R47395 DVSS.n8836 DVSS.n8702 0.0380882
R47396 DVSS.n8829 DVSS.n8702 0.0380882
R47397 DVSS.n8829 DVSS.n8825 0.0380882
R47398 DVSS.n8825 DVSS.n8824 0.0380882
R47399 DVSS.n8824 DVSS.n8704 0.0380882
R47400 DVSS.n8817 DVSS.n8704 0.0380882
R47401 DVSS.n8817 DVSS.n8813 0.0380882
R47402 DVSS.n8813 DVSS.n8812 0.0380882
R47403 DVSS.n8812 DVSS.n8706 0.0380882
R47404 DVSS.n8805 DVSS.n8706 0.0380882
R47405 DVSS.n8805 DVSS.n8801 0.0380882
R47406 DVSS.n8801 DVSS.n8800 0.0380882
R47407 DVSS.n8800 DVSS.n8708 0.0380882
R47408 DVSS.n8793 DVSS.n8708 0.0380882
R47409 DVSS.n8793 DVSS.n8789 0.0380882
R47410 DVSS.n8789 DVSS.n8788 0.0380882
R47411 DVSS.n8788 DVSS.n8710 0.0380882
R47412 DVSS.n8781 DVSS.n8710 0.0380882
R47413 DVSS.n8781 DVSS.n8777 0.0380882
R47414 DVSS.n8777 DVSS.n8776 0.0380882
R47415 DVSS.n8776 DVSS.n8712 0.0380882
R47416 DVSS.n8769 DVSS.n8712 0.0380882
R47417 DVSS.n8769 DVSS.n8765 0.0380882
R47418 DVSS.n8765 DVSS.n8764 0.0380882
R47419 DVSS.n8764 DVSS.n8714 0.0380882
R47420 DVSS.n8757 DVSS.n8714 0.0380882
R47421 DVSS.n8757 DVSS.n8753 0.0380882
R47422 DVSS.n8753 DVSS.n8752 0.0380882
R47423 DVSS.n8752 DVSS.n8716 0.0380882
R47424 DVSS.n8745 DVSS.n8716 0.0380882
R47425 DVSS.n8745 DVSS.n8741 0.0380882
R47426 DVSS.n8741 DVSS.n8740 0.0380882
R47427 DVSS.n8740 DVSS.n8718 0.0380882
R47428 DVSS.n8733 DVSS.n8718 0.0380882
R47429 DVSS.n8733 DVSS.n8729 0.0380882
R47430 DVSS.n8729 DVSS.n8728 0.0380882
R47431 DVSS.n8728 DVSS.n8722 0.0380882
R47432 DVSS.n8722 DVSS.n8721 0.0380882
R47433 DVSS.n8998 DVSS.n8997 0.0380882
R47434 DVSS.n8999 DVSS.n8998 0.0380882
R47435 DVSS.n8999 DVSS.n3038 0.0380882
R47436 DVSS.n9006 DVSS.n3038 0.0380882
R47437 DVSS.n9007 DVSS.n9006 0.0380882
R47438 DVSS.n9008 DVSS.n9007 0.0380882
R47439 DVSS.n9008 DVSS.n3035 0.0380882
R47440 DVSS.n9015 DVSS.n3035 0.0380882
R47441 DVSS.n9016 DVSS.n9015 0.0380882
R47442 DVSS.n9017 DVSS.n9016 0.0380882
R47443 DVSS.n9017 DVSS.n3032 0.0380882
R47444 DVSS.n9024 DVSS.n3032 0.0380882
R47445 DVSS.n9025 DVSS.n9024 0.0380882
R47446 DVSS.n9026 DVSS.n9025 0.0380882
R47447 DVSS.n9026 DVSS.n3029 0.0380882
R47448 DVSS.n9033 DVSS.n3029 0.0380882
R47449 DVSS.n9034 DVSS.n9033 0.0380882
R47450 DVSS.n9035 DVSS.n9034 0.0380882
R47451 DVSS.n9035 DVSS.n3026 0.0380882
R47452 DVSS.n9042 DVSS.n3026 0.0380882
R47453 DVSS.n9043 DVSS.n9042 0.0380882
R47454 DVSS.n9044 DVSS.n9043 0.0380882
R47455 DVSS.n9044 DVSS.n3023 0.0380882
R47456 DVSS.n9051 DVSS.n3023 0.0380882
R47457 DVSS.n9052 DVSS.n9051 0.0380882
R47458 DVSS.n9053 DVSS.n9052 0.0380882
R47459 DVSS.n9053 DVSS.n3020 0.0380882
R47460 DVSS.n9060 DVSS.n3020 0.0380882
R47461 DVSS.n9061 DVSS.n9060 0.0380882
R47462 DVSS.n9062 DVSS.n9061 0.0380882
R47463 DVSS.n9062 DVSS.n3017 0.0380882
R47464 DVSS.n9069 DVSS.n3017 0.0380882
R47465 DVSS.n9070 DVSS.n9069 0.0380882
R47466 DVSS.n9071 DVSS.n9070 0.0380882
R47467 DVSS.n9071 DVSS.n3014 0.0380882
R47468 DVSS.n9078 DVSS.n3014 0.0380882
R47469 DVSS.n9079 DVSS.n9078 0.0380882
R47470 DVSS.n9080 DVSS.n9079 0.0380882
R47471 DVSS.n9080 DVSS.n3011 0.0380882
R47472 DVSS.n9087 DVSS.n3011 0.0380882
R47473 DVSS.n9088 DVSS.n9087 0.0380882
R47474 DVSS.n9089 DVSS.n9088 0.0380882
R47475 DVSS.n9089 DVSS.n3008 0.0380882
R47476 DVSS.n9096 DVSS.n3008 0.0380882
R47477 DVSS.n9097 DVSS.n9096 0.0380882
R47478 DVSS.n9098 DVSS.n9097 0.0380882
R47479 DVSS.n9098 DVSS.n3005 0.0380882
R47480 DVSS.n9105 DVSS.n3005 0.0380882
R47481 DVSS.n9106 DVSS.n9105 0.0380882
R47482 DVSS.n9107 DVSS.n9106 0.0380882
R47483 DVSS.n9107 DVSS.n3002 0.0380882
R47484 DVSS.n9114 DVSS.n3002 0.0380882
R47485 DVSS.n9115 DVSS.n9114 0.0380882
R47486 DVSS.n9116 DVSS.n9115 0.0380882
R47487 DVSS.n9116 DVSS.n2999 0.0380882
R47488 DVSS.n9123 DVSS.n2999 0.0380882
R47489 DVSS.n9124 DVSS.n9123 0.0380882
R47490 DVSS.n9125 DVSS.n9124 0.0380882
R47491 DVSS.n9125 DVSS.n2996 0.0380882
R47492 DVSS.n9132 DVSS.n2996 0.0380882
R47493 DVSS.n9133 DVSS.n9132 0.0380882
R47494 DVSS.n9134 DVSS.n9133 0.0380882
R47495 DVSS.n9134 DVSS.n2993 0.0380882
R47496 DVSS.n9141 DVSS.n2993 0.0380882
R47497 DVSS.n9142 DVSS.n9141 0.0380882
R47498 DVSS.n9143 DVSS.n9142 0.0380882
R47499 DVSS.n9143 DVSS.n2990 0.0380882
R47500 DVSS.n9150 DVSS.n2990 0.0380882
R47501 DVSS.n9151 DVSS.n9150 0.0380882
R47502 DVSS.n9152 DVSS.n9151 0.0380882
R47503 DVSS.n9152 DVSS.n2987 0.0380882
R47504 DVSS.n9159 DVSS.n2987 0.0380882
R47505 DVSS.n9160 DVSS.n9159 0.0380882
R47506 DVSS.n9161 DVSS.n9160 0.0380882
R47507 DVSS.n9161 DVSS.n2984 0.0380882
R47508 DVSS.n9168 DVSS.n2984 0.0380882
R47509 DVSS.n9169 DVSS.n9168 0.0380882
R47510 DVSS.n9170 DVSS.n9169 0.0380882
R47511 DVSS.n9170 DVSS.n2981 0.0380882
R47512 DVSS.n9177 DVSS.n2981 0.0380882
R47513 DVSS.n9178 DVSS.n9177 0.0380882
R47514 DVSS.n9179 DVSS.n9178 0.0380882
R47515 DVSS.n9179 DVSS.n2884 0.0380882
R47516 DVSS.n3039 DVSS.n2935 0.0380882
R47517 DVSS.n9001 DVSS.n3039 0.0380882
R47518 DVSS.n9003 DVSS.n9001 0.0380882
R47519 DVSS.n9005 DVSS.n9003 0.0380882
R47520 DVSS.n9005 DVSS.n3037 0.0380882
R47521 DVSS.n9010 DVSS.n3037 0.0380882
R47522 DVSS.n9012 DVSS.n9010 0.0380882
R47523 DVSS.n9014 DVSS.n9012 0.0380882
R47524 DVSS.n9014 DVSS.n3034 0.0380882
R47525 DVSS.n9019 DVSS.n3034 0.0380882
R47526 DVSS.n9021 DVSS.n9019 0.0380882
R47527 DVSS.n9023 DVSS.n9021 0.0380882
R47528 DVSS.n9023 DVSS.n3031 0.0380882
R47529 DVSS.n9028 DVSS.n3031 0.0380882
R47530 DVSS.n9030 DVSS.n9028 0.0380882
R47531 DVSS.n9032 DVSS.n9030 0.0380882
R47532 DVSS.n9032 DVSS.n3028 0.0380882
R47533 DVSS.n9037 DVSS.n3028 0.0380882
R47534 DVSS.n9039 DVSS.n9037 0.0380882
R47535 DVSS.n9041 DVSS.n9039 0.0380882
R47536 DVSS.n9041 DVSS.n3025 0.0380882
R47537 DVSS.n9046 DVSS.n3025 0.0380882
R47538 DVSS.n9048 DVSS.n9046 0.0380882
R47539 DVSS.n9050 DVSS.n9048 0.0380882
R47540 DVSS.n9050 DVSS.n3022 0.0380882
R47541 DVSS.n9055 DVSS.n3022 0.0380882
R47542 DVSS.n9057 DVSS.n9055 0.0380882
R47543 DVSS.n9059 DVSS.n9057 0.0380882
R47544 DVSS.n9059 DVSS.n3019 0.0380882
R47545 DVSS.n9064 DVSS.n3019 0.0380882
R47546 DVSS.n9066 DVSS.n9064 0.0380882
R47547 DVSS.n9068 DVSS.n9066 0.0380882
R47548 DVSS.n9068 DVSS.n3016 0.0380882
R47549 DVSS.n9073 DVSS.n3016 0.0380882
R47550 DVSS.n9075 DVSS.n9073 0.0380882
R47551 DVSS.n9077 DVSS.n9075 0.0380882
R47552 DVSS.n9077 DVSS.n3013 0.0380882
R47553 DVSS.n9082 DVSS.n3013 0.0380882
R47554 DVSS.n9084 DVSS.n9082 0.0380882
R47555 DVSS.n9086 DVSS.n9084 0.0380882
R47556 DVSS.n9086 DVSS.n3010 0.0380882
R47557 DVSS.n9091 DVSS.n3010 0.0380882
R47558 DVSS.n9093 DVSS.n9091 0.0380882
R47559 DVSS.n9095 DVSS.n9093 0.0380882
R47560 DVSS.n9095 DVSS.n3007 0.0380882
R47561 DVSS.n9100 DVSS.n3007 0.0380882
R47562 DVSS.n9102 DVSS.n9100 0.0380882
R47563 DVSS.n9104 DVSS.n9102 0.0380882
R47564 DVSS.n9104 DVSS.n3004 0.0380882
R47565 DVSS.n9109 DVSS.n3004 0.0380882
R47566 DVSS.n9111 DVSS.n9109 0.0380882
R47567 DVSS.n9113 DVSS.n9111 0.0380882
R47568 DVSS.n9113 DVSS.n3001 0.0380882
R47569 DVSS.n9118 DVSS.n3001 0.0380882
R47570 DVSS.n9120 DVSS.n9118 0.0380882
R47571 DVSS.n9122 DVSS.n9120 0.0380882
R47572 DVSS.n9122 DVSS.n2998 0.0380882
R47573 DVSS.n9127 DVSS.n2998 0.0380882
R47574 DVSS.n9129 DVSS.n9127 0.0380882
R47575 DVSS.n9131 DVSS.n9129 0.0380882
R47576 DVSS.n9131 DVSS.n2995 0.0380882
R47577 DVSS.n9136 DVSS.n2995 0.0380882
R47578 DVSS.n9138 DVSS.n9136 0.0380882
R47579 DVSS.n9140 DVSS.n9138 0.0380882
R47580 DVSS.n9140 DVSS.n2992 0.0380882
R47581 DVSS.n9145 DVSS.n2992 0.0380882
R47582 DVSS.n9147 DVSS.n9145 0.0380882
R47583 DVSS.n9149 DVSS.n9147 0.0380882
R47584 DVSS.n9149 DVSS.n2989 0.0380882
R47585 DVSS.n9154 DVSS.n2989 0.0380882
R47586 DVSS.n9156 DVSS.n9154 0.0380882
R47587 DVSS.n9158 DVSS.n9156 0.0380882
R47588 DVSS.n9158 DVSS.n2986 0.0380882
R47589 DVSS.n9163 DVSS.n2986 0.0380882
R47590 DVSS.n9165 DVSS.n9163 0.0380882
R47591 DVSS.n9167 DVSS.n9165 0.0380882
R47592 DVSS.n9167 DVSS.n2983 0.0380882
R47593 DVSS.n9172 DVSS.n2983 0.0380882
R47594 DVSS.n9174 DVSS.n9172 0.0380882
R47595 DVSS.n9176 DVSS.n9174 0.0380882
R47596 DVSS.n9176 DVSS.n2980 0.0380882
R47597 DVSS.n9181 DVSS.n2980 0.0380882
R47598 DVSS.n9182 DVSS.n9181 0.0380882
R47599 DVSS.n9208 DVSS.n9207 0.0380882
R47600 DVSS.n9209 DVSS.n9208 0.0380882
R47601 DVSS.n9209 DVSS.n2871 0.0380882
R47602 DVSS.n9219 DVSS.n2871 0.0380882
R47603 DVSS.n9220 DVSS.n9219 0.0380882
R47604 DVSS.n9221 DVSS.n9220 0.0380882
R47605 DVSS.n9221 DVSS.n2869 0.0380882
R47606 DVSS.n9231 DVSS.n2869 0.0380882
R47607 DVSS.n9232 DVSS.n9231 0.0380882
R47608 DVSS.n9233 DVSS.n9232 0.0380882
R47609 DVSS.n9233 DVSS.n2867 0.0380882
R47610 DVSS.n9243 DVSS.n2867 0.0380882
R47611 DVSS.n9244 DVSS.n9243 0.0380882
R47612 DVSS.n9245 DVSS.n9244 0.0380882
R47613 DVSS.n9245 DVSS.n2865 0.0380882
R47614 DVSS.n9255 DVSS.n2865 0.0380882
R47615 DVSS.n9256 DVSS.n9255 0.0380882
R47616 DVSS.n9257 DVSS.n9256 0.0380882
R47617 DVSS.n9257 DVSS.n2863 0.0380882
R47618 DVSS.n9267 DVSS.n2863 0.0380882
R47619 DVSS.n9268 DVSS.n9267 0.0380882
R47620 DVSS.n9269 DVSS.n9268 0.0380882
R47621 DVSS.n9269 DVSS.n2861 0.0380882
R47622 DVSS.n9279 DVSS.n2861 0.0380882
R47623 DVSS.n9280 DVSS.n9279 0.0380882
R47624 DVSS.n9281 DVSS.n9280 0.0380882
R47625 DVSS.n9281 DVSS.n2859 0.0380882
R47626 DVSS.n9291 DVSS.n2859 0.0380882
R47627 DVSS.n9292 DVSS.n9291 0.0380882
R47628 DVSS.n9293 DVSS.n9292 0.0380882
R47629 DVSS.n9293 DVSS.n2857 0.0380882
R47630 DVSS.n9303 DVSS.n2857 0.0380882
R47631 DVSS.n9304 DVSS.n9303 0.0380882
R47632 DVSS.n9305 DVSS.n9304 0.0380882
R47633 DVSS.n9305 DVSS.n2855 0.0380882
R47634 DVSS.n9315 DVSS.n2855 0.0380882
R47635 DVSS.n9316 DVSS.n9315 0.0380882
R47636 DVSS.n9317 DVSS.n9316 0.0380882
R47637 DVSS.n9317 DVSS.n2853 0.0380882
R47638 DVSS.n9327 DVSS.n2853 0.0380882
R47639 DVSS.n9328 DVSS.n9327 0.0380882
R47640 DVSS.n9329 DVSS.n9328 0.0380882
R47641 DVSS.n9329 DVSS.n2851 0.0380882
R47642 DVSS.n9339 DVSS.n2851 0.0380882
R47643 DVSS.n9340 DVSS.n9339 0.0380882
R47644 DVSS.n9341 DVSS.n9340 0.0380882
R47645 DVSS.n9341 DVSS.n2849 0.0380882
R47646 DVSS.n9351 DVSS.n2849 0.0380882
R47647 DVSS.n9352 DVSS.n9351 0.0380882
R47648 DVSS.n9353 DVSS.n9352 0.0380882
R47649 DVSS.n9353 DVSS.n2847 0.0380882
R47650 DVSS.n9363 DVSS.n2847 0.0380882
R47651 DVSS.n9364 DVSS.n9363 0.0380882
R47652 DVSS.n9365 DVSS.n9364 0.0380882
R47653 DVSS.n9365 DVSS.n2845 0.0380882
R47654 DVSS.n9375 DVSS.n2845 0.0380882
R47655 DVSS.n9376 DVSS.n9375 0.0380882
R47656 DVSS.n9377 DVSS.n9376 0.0380882
R47657 DVSS.n9377 DVSS.n2843 0.0380882
R47658 DVSS.n9387 DVSS.n2843 0.0380882
R47659 DVSS.n9388 DVSS.n9387 0.0380882
R47660 DVSS.n9389 DVSS.n9388 0.0380882
R47661 DVSS.n9389 DVSS.n2841 0.0380882
R47662 DVSS.n9399 DVSS.n2841 0.0380882
R47663 DVSS.n9400 DVSS.n9399 0.0380882
R47664 DVSS.n9401 DVSS.n9400 0.0380882
R47665 DVSS.n9401 DVSS.n2839 0.0380882
R47666 DVSS.n9411 DVSS.n2839 0.0380882
R47667 DVSS.n9412 DVSS.n9411 0.0380882
R47668 DVSS.n9413 DVSS.n9412 0.0380882
R47669 DVSS.n9413 DVSS.n2837 0.0380882
R47670 DVSS.n9423 DVSS.n2837 0.0380882
R47671 DVSS.n9424 DVSS.n9423 0.0380882
R47672 DVSS.n9425 DVSS.n9424 0.0380882
R47673 DVSS.n9425 DVSS.n2835 0.0380882
R47674 DVSS.n9435 DVSS.n2835 0.0380882
R47675 DVSS.n9436 DVSS.n9435 0.0380882
R47676 DVSS.n9437 DVSS.n9436 0.0380882
R47677 DVSS.n9437 DVSS.n2833 0.0380882
R47678 DVSS.n9447 DVSS.n2833 0.0380882
R47679 DVSS.n9448 DVSS.n9447 0.0380882
R47680 DVSS.n9450 DVSS.n9448 0.0380882
R47681 DVSS.n9450 DVSS.n9449 0.0380882
R47682 DVSS.n9206 DVSS.n2874 0.0380882
R47683 DVSS.n9210 DVSS.n2874 0.0380882
R47684 DVSS.n9214 DVSS.n9210 0.0380882
R47685 DVSS.n9218 DVSS.n9214 0.0380882
R47686 DVSS.n9218 DVSS.n2870 0.0380882
R47687 DVSS.n9222 DVSS.n2870 0.0380882
R47688 DVSS.n9226 DVSS.n9222 0.0380882
R47689 DVSS.n9230 DVSS.n9226 0.0380882
R47690 DVSS.n9230 DVSS.n2868 0.0380882
R47691 DVSS.n9234 DVSS.n2868 0.0380882
R47692 DVSS.n9238 DVSS.n9234 0.0380882
R47693 DVSS.n9242 DVSS.n9238 0.0380882
R47694 DVSS.n9242 DVSS.n2866 0.0380882
R47695 DVSS.n9246 DVSS.n2866 0.0380882
R47696 DVSS.n9250 DVSS.n9246 0.0380882
R47697 DVSS.n9254 DVSS.n9250 0.0380882
R47698 DVSS.n9254 DVSS.n2864 0.0380882
R47699 DVSS.n9258 DVSS.n2864 0.0380882
R47700 DVSS.n9262 DVSS.n9258 0.0380882
R47701 DVSS.n9266 DVSS.n9262 0.0380882
R47702 DVSS.n9266 DVSS.n2862 0.0380882
R47703 DVSS.n9270 DVSS.n2862 0.0380882
R47704 DVSS.n9274 DVSS.n9270 0.0380882
R47705 DVSS.n9278 DVSS.n9274 0.0380882
R47706 DVSS.n9278 DVSS.n2860 0.0380882
R47707 DVSS.n9282 DVSS.n2860 0.0380882
R47708 DVSS.n9286 DVSS.n9282 0.0380882
R47709 DVSS.n9290 DVSS.n9286 0.0380882
R47710 DVSS.n9290 DVSS.n2858 0.0380882
R47711 DVSS.n9294 DVSS.n2858 0.0380882
R47712 DVSS.n9298 DVSS.n9294 0.0380882
R47713 DVSS.n9302 DVSS.n9298 0.0380882
R47714 DVSS.n9302 DVSS.n2856 0.0380882
R47715 DVSS.n9306 DVSS.n2856 0.0380882
R47716 DVSS.n9310 DVSS.n9306 0.0380882
R47717 DVSS.n9314 DVSS.n9310 0.0380882
R47718 DVSS.n9314 DVSS.n2854 0.0380882
R47719 DVSS.n9318 DVSS.n2854 0.0380882
R47720 DVSS.n9322 DVSS.n9318 0.0380882
R47721 DVSS.n9326 DVSS.n9322 0.0380882
R47722 DVSS.n9326 DVSS.n2852 0.0380882
R47723 DVSS.n9330 DVSS.n2852 0.0380882
R47724 DVSS.n9334 DVSS.n9330 0.0380882
R47725 DVSS.n9338 DVSS.n9334 0.0380882
R47726 DVSS.n9338 DVSS.n2850 0.0380882
R47727 DVSS.n9342 DVSS.n2850 0.0380882
R47728 DVSS.n9346 DVSS.n9342 0.0380882
R47729 DVSS.n9350 DVSS.n9346 0.0380882
R47730 DVSS.n9350 DVSS.n2848 0.0380882
R47731 DVSS.n9354 DVSS.n2848 0.0380882
R47732 DVSS.n9358 DVSS.n9354 0.0380882
R47733 DVSS.n9362 DVSS.n9358 0.0380882
R47734 DVSS.n9362 DVSS.n2846 0.0380882
R47735 DVSS.n9366 DVSS.n2846 0.0380882
R47736 DVSS.n9370 DVSS.n9366 0.0380882
R47737 DVSS.n9374 DVSS.n9370 0.0380882
R47738 DVSS.n9374 DVSS.n2844 0.0380882
R47739 DVSS.n9378 DVSS.n2844 0.0380882
R47740 DVSS.n9382 DVSS.n9378 0.0380882
R47741 DVSS.n9386 DVSS.n9382 0.0380882
R47742 DVSS.n9386 DVSS.n2842 0.0380882
R47743 DVSS.n9390 DVSS.n2842 0.0380882
R47744 DVSS.n9394 DVSS.n9390 0.0380882
R47745 DVSS.n9398 DVSS.n9394 0.0380882
R47746 DVSS.n9398 DVSS.n2840 0.0380882
R47747 DVSS.n9402 DVSS.n2840 0.0380882
R47748 DVSS.n9406 DVSS.n9402 0.0380882
R47749 DVSS.n9410 DVSS.n9406 0.0380882
R47750 DVSS.n9410 DVSS.n2838 0.0380882
R47751 DVSS.n9414 DVSS.n2838 0.0380882
R47752 DVSS.n9418 DVSS.n9414 0.0380882
R47753 DVSS.n9422 DVSS.n9418 0.0380882
R47754 DVSS.n9422 DVSS.n2836 0.0380882
R47755 DVSS.n9426 DVSS.n2836 0.0380882
R47756 DVSS.n9430 DVSS.n9426 0.0380882
R47757 DVSS.n9434 DVSS.n9430 0.0380882
R47758 DVSS.n9434 DVSS.n2834 0.0380882
R47759 DVSS.n9438 DVSS.n2834 0.0380882
R47760 DVSS.n9442 DVSS.n9438 0.0380882
R47761 DVSS.n9446 DVSS.n9442 0.0380882
R47762 DVSS.n9446 DVSS.n2832 0.0380882
R47763 DVSS.n9451 DVSS.n2832 0.0380882
R47764 DVSS.n9451 DVSS.n2830 0.0380882
R47765 DVSS.n9754 DVSS.n2733 0.0380882
R47766 DVSS.n9754 DVSS.n9753 0.0380882
R47767 DVSS.n9753 DVSS.n9752 0.0380882
R47768 DVSS.n9752 DVSS.n9470 0.0380882
R47769 DVSS.n9742 DVSS.n9470 0.0380882
R47770 DVSS.n9742 DVSS.n9741 0.0380882
R47771 DVSS.n9741 DVSS.n9740 0.0380882
R47772 DVSS.n9740 DVSS.n9472 0.0380882
R47773 DVSS.n9730 DVSS.n9472 0.0380882
R47774 DVSS.n9730 DVSS.n9729 0.0380882
R47775 DVSS.n9729 DVSS.n9728 0.0380882
R47776 DVSS.n9728 DVSS.n9474 0.0380882
R47777 DVSS.n9718 DVSS.n9474 0.0380882
R47778 DVSS.n9718 DVSS.n9717 0.0380882
R47779 DVSS.n9717 DVSS.n9716 0.0380882
R47780 DVSS.n9716 DVSS.n9476 0.0380882
R47781 DVSS.n9706 DVSS.n9476 0.0380882
R47782 DVSS.n9706 DVSS.n9705 0.0380882
R47783 DVSS.n9705 DVSS.n9704 0.0380882
R47784 DVSS.n9704 DVSS.n9478 0.0380882
R47785 DVSS.n9694 DVSS.n9478 0.0380882
R47786 DVSS.n9694 DVSS.n9693 0.0380882
R47787 DVSS.n9693 DVSS.n9692 0.0380882
R47788 DVSS.n9692 DVSS.n9480 0.0380882
R47789 DVSS.n9682 DVSS.n9480 0.0380882
R47790 DVSS.n9682 DVSS.n9681 0.0380882
R47791 DVSS.n9681 DVSS.n9680 0.0380882
R47792 DVSS.n9680 DVSS.n9482 0.0380882
R47793 DVSS.n9670 DVSS.n9482 0.0380882
R47794 DVSS.n9670 DVSS.n9669 0.0380882
R47795 DVSS.n9669 DVSS.n9668 0.0380882
R47796 DVSS.n9668 DVSS.n9484 0.0380882
R47797 DVSS.n9658 DVSS.n9484 0.0380882
R47798 DVSS.n9658 DVSS.n9657 0.0380882
R47799 DVSS.n9657 DVSS.n9656 0.0380882
R47800 DVSS.n9656 DVSS.n9486 0.0380882
R47801 DVSS.n9646 DVSS.n9486 0.0380882
R47802 DVSS.n9646 DVSS.n9645 0.0380882
R47803 DVSS.n9645 DVSS.n9644 0.0380882
R47804 DVSS.n9644 DVSS.n9488 0.0380882
R47805 DVSS.n9634 DVSS.n9488 0.0380882
R47806 DVSS.n9634 DVSS.n9633 0.0380882
R47807 DVSS.n9633 DVSS.n9632 0.0380882
R47808 DVSS.n9632 DVSS.n9490 0.0380882
R47809 DVSS.n9622 DVSS.n9490 0.0380882
R47810 DVSS.n9622 DVSS.n9621 0.0380882
R47811 DVSS.n9621 DVSS.n9620 0.0380882
R47812 DVSS.n9620 DVSS.n9492 0.0380882
R47813 DVSS.n9610 DVSS.n9492 0.0380882
R47814 DVSS.n9610 DVSS.n9609 0.0380882
R47815 DVSS.n9609 DVSS.n9608 0.0380882
R47816 DVSS.n9608 DVSS.n9494 0.0380882
R47817 DVSS.n9598 DVSS.n9494 0.0380882
R47818 DVSS.n9598 DVSS.n9597 0.0380882
R47819 DVSS.n9597 DVSS.n9596 0.0380882
R47820 DVSS.n9596 DVSS.n9496 0.0380882
R47821 DVSS.n9586 DVSS.n9496 0.0380882
R47822 DVSS.n9586 DVSS.n9585 0.0380882
R47823 DVSS.n9585 DVSS.n9584 0.0380882
R47824 DVSS.n9584 DVSS.n9498 0.0380882
R47825 DVSS.n9574 DVSS.n9498 0.0380882
R47826 DVSS.n9574 DVSS.n9573 0.0380882
R47827 DVSS.n9573 DVSS.n9572 0.0380882
R47828 DVSS.n9572 DVSS.n9500 0.0380882
R47829 DVSS.n9562 DVSS.n9500 0.0380882
R47830 DVSS.n9562 DVSS.n9561 0.0380882
R47831 DVSS.n9561 DVSS.n9560 0.0380882
R47832 DVSS.n9560 DVSS.n9502 0.0380882
R47833 DVSS.n9550 DVSS.n9502 0.0380882
R47834 DVSS.n9550 DVSS.n9549 0.0380882
R47835 DVSS.n9549 DVSS.n9548 0.0380882
R47836 DVSS.n9548 DVSS.n9504 0.0380882
R47837 DVSS.n9538 DVSS.n9504 0.0380882
R47838 DVSS.n9538 DVSS.n9537 0.0380882
R47839 DVSS.n9537 DVSS.n9536 0.0380882
R47840 DVSS.n9536 DVSS.n9506 0.0380882
R47841 DVSS.n9526 DVSS.n9506 0.0380882
R47842 DVSS.n9526 DVSS.n9525 0.0380882
R47843 DVSS.n9525 DVSS.n9524 0.0380882
R47844 DVSS.n9524 DVSS.n9508 0.0380882
R47845 DVSS.n9514 DVSS.n9508 0.0380882
R47846 DVSS.n9514 DVSS.n9513 0.0380882
R47847 DVSS.n9513 DVSS.n9512 0.0380882
R47848 DVSS.n9756 DVSS.n9755 0.0380882
R47849 DVSS.n9755 DVSS.n9469 0.0380882
R47850 DVSS.n9751 DVSS.n9469 0.0380882
R47851 DVSS.n9751 DVSS.n9747 0.0380882
R47852 DVSS.n9747 DVSS.n9746 0.0380882
R47853 DVSS.n9746 DVSS.n9471 0.0380882
R47854 DVSS.n9739 DVSS.n9471 0.0380882
R47855 DVSS.n9739 DVSS.n9735 0.0380882
R47856 DVSS.n9735 DVSS.n9734 0.0380882
R47857 DVSS.n9734 DVSS.n9473 0.0380882
R47858 DVSS.n9727 DVSS.n9473 0.0380882
R47859 DVSS.n9727 DVSS.n9723 0.0380882
R47860 DVSS.n9723 DVSS.n9722 0.0380882
R47861 DVSS.n9722 DVSS.n9475 0.0380882
R47862 DVSS.n9715 DVSS.n9475 0.0380882
R47863 DVSS.n9715 DVSS.n9711 0.0380882
R47864 DVSS.n9711 DVSS.n9710 0.0380882
R47865 DVSS.n9710 DVSS.n9477 0.0380882
R47866 DVSS.n9703 DVSS.n9477 0.0380882
R47867 DVSS.n9703 DVSS.n9699 0.0380882
R47868 DVSS.n9699 DVSS.n9698 0.0380882
R47869 DVSS.n9698 DVSS.n9479 0.0380882
R47870 DVSS.n9691 DVSS.n9479 0.0380882
R47871 DVSS.n9691 DVSS.n9687 0.0380882
R47872 DVSS.n9687 DVSS.n9686 0.0380882
R47873 DVSS.n9686 DVSS.n9481 0.0380882
R47874 DVSS.n9679 DVSS.n9481 0.0380882
R47875 DVSS.n9679 DVSS.n9675 0.0380882
R47876 DVSS.n9675 DVSS.n9674 0.0380882
R47877 DVSS.n9674 DVSS.n9483 0.0380882
R47878 DVSS.n9667 DVSS.n9483 0.0380882
R47879 DVSS.n9667 DVSS.n9663 0.0380882
R47880 DVSS.n9663 DVSS.n9662 0.0380882
R47881 DVSS.n9662 DVSS.n9485 0.0380882
R47882 DVSS.n9655 DVSS.n9485 0.0380882
R47883 DVSS.n9655 DVSS.n9651 0.0380882
R47884 DVSS.n9651 DVSS.n9650 0.0380882
R47885 DVSS.n9650 DVSS.n9487 0.0380882
R47886 DVSS.n9643 DVSS.n9487 0.0380882
R47887 DVSS.n9643 DVSS.n9639 0.0380882
R47888 DVSS.n9639 DVSS.n9638 0.0380882
R47889 DVSS.n9638 DVSS.n9489 0.0380882
R47890 DVSS.n9631 DVSS.n9489 0.0380882
R47891 DVSS.n9631 DVSS.n9627 0.0380882
R47892 DVSS.n9627 DVSS.n9626 0.0380882
R47893 DVSS.n9626 DVSS.n9491 0.0380882
R47894 DVSS.n9619 DVSS.n9491 0.0380882
R47895 DVSS.n9619 DVSS.n9615 0.0380882
R47896 DVSS.n9615 DVSS.n9614 0.0380882
R47897 DVSS.n9614 DVSS.n9493 0.0380882
R47898 DVSS.n9607 DVSS.n9493 0.0380882
R47899 DVSS.n9607 DVSS.n9603 0.0380882
R47900 DVSS.n9603 DVSS.n9602 0.0380882
R47901 DVSS.n9602 DVSS.n9495 0.0380882
R47902 DVSS.n9595 DVSS.n9495 0.0380882
R47903 DVSS.n9595 DVSS.n9591 0.0380882
R47904 DVSS.n9591 DVSS.n9590 0.0380882
R47905 DVSS.n9590 DVSS.n9497 0.0380882
R47906 DVSS.n9583 DVSS.n9497 0.0380882
R47907 DVSS.n9583 DVSS.n9579 0.0380882
R47908 DVSS.n9579 DVSS.n9578 0.0380882
R47909 DVSS.n9578 DVSS.n9499 0.0380882
R47910 DVSS.n9571 DVSS.n9499 0.0380882
R47911 DVSS.n9571 DVSS.n9567 0.0380882
R47912 DVSS.n9567 DVSS.n9566 0.0380882
R47913 DVSS.n9566 DVSS.n9501 0.0380882
R47914 DVSS.n9559 DVSS.n9501 0.0380882
R47915 DVSS.n9559 DVSS.n9555 0.0380882
R47916 DVSS.n9555 DVSS.n9554 0.0380882
R47917 DVSS.n9554 DVSS.n9503 0.0380882
R47918 DVSS.n9547 DVSS.n9503 0.0380882
R47919 DVSS.n9547 DVSS.n9543 0.0380882
R47920 DVSS.n9543 DVSS.n9542 0.0380882
R47921 DVSS.n9542 DVSS.n9505 0.0380882
R47922 DVSS.n9535 DVSS.n9505 0.0380882
R47923 DVSS.n9535 DVSS.n9531 0.0380882
R47924 DVSS.n9531 DVSS.n9530 0.0380882
R47925 DVSS.n9530 DVSS.n9507 0.0380882
R47926 DVSS.n9523 DVSS.n9507 0.0380882
R47927 DVSS.n9523 DVSS.n9519 0.0380882
R47928 DVSS.n9519 DVSS.n9518 0.0380882
R47929 DVSS.n9518 DVSS.n9509 0.0380882
R47930 DVSS.n9511 DVSS.n9509 0.0380882
R47931 DVSS.n9857 DVSS.n2712 0.0380882
R47932 DVSS.n9868 DVSS.n9857 0.0380882
R47933 DVSS.n9869 DVSS.n9868 0.0380882
R47934 DVSS.n9870 DVSS.n9869 0.0380882
R47935 DVSS.n9870 DVSS.n9853 0.0380882
R47936 DVSS.n9880 DVSS.n9853 0.0380882
R47937 DVSS.n9881 DVSS.n9880 0.0380882
R47938 DVSS.n9882 DVSS.n9881 0.0380882
R47939 DVSS.n9882 DVSS.n9849 0.0380882
R47940 DVSS.n9892 DVSS.n9849 0.0380882
R47941 DVSS.n9893 DVSS.n9892 0.0380882
R47942 DVSS.n9894 DVSS.n9893 0.0380882
R47943 DVSS.n9894 DVSS.n9845 0.0380882
R47944 DVSS.n9904 DVSS.n9845 0.0380882
R47945 DVSS.n9905 DVSS.n9904 0.0380882
R47946 DVSS.n9906 DVSS.n9905 0.0380882
R47947 DVSS.n9906 DVSS.n9841 0.0380882
R47948 DVSS.n9916 DVSS.n9841 0.0380882
R47949 DVSS.n9917 DVSS.n9916 0.0380882
R47950 DVSS.n9918 DVSS.n9917 0.0380882
R47951 DVSS.n9918 DVSS.n9837 0.0380882
R47952 DVSS.n9928 DVSS.n9837 0.0380882
R47953 DVSS.n9929 DVSS.n9928 0.0380882
R47954 DVSS.n9930 DVSS.n9929 0.0380882
R47955 DVSS.n9930 DVSS.n9833 0.0380882
R47956 DVSS.n9940 DVSS.n9833 0.0380882
R47957 DVSS.n9941 DVSS.n9940 0.0380882
R47958 DVSS.n9942 DVSS.n9941 0.0380882
R47959 DVSS.n9942 DVSS.n9829 0.0380882
R47960 DVSS.n9952 DVSS.n9829 0.0380882
R47961 DVSS.n9953 DVSS.n9952 0.0380882
R47962 DVSS.n9954 DVSS.n9953 0.0380882
R47963 DVSS.n9954 DVSS.n9825 0.0380882
R47964 DVSS.n9964 DVSS.n9825 0.0380882
R47965 DVSS.n9965 DVSS.n9964 0.0380882
R47966 DVSS.n9966 DVSS.n9965 0.0380882
R47967 DVSS.n9966 DVSS.n9821 0.0380882
R47968 DVSS.n9976 DVSS.n9821 0.0380882
R47969 DVSS.n9977 DVSS.n9976 0.0380882
R47970 DVSS.n9978 DVSS.n9977 0.0380882
R47971 DVSS.n9978 DVSS.n9817 0.0380882
R47972 DVSS.n9988 DVSS.n9817 0.0380882
R47973 DVSS.n9989 DVSS.n9988 0.0380882
R47974 DVSS.n9990 DVSS.n9989 0.0380882
R47975 DVSS.n9990 DVSS.n9813 0.0380882
R47976 DVSS.n10000 DVSS.n9813 0.0380882
R47977 DVSS.n10001 DVSS.n10000 0.0380882
R47978 DVSS.n10002 DVSS.n10001 0.0380882
R47979 DVSS.n10002 DVSS.n9809 0.0380882
R47980 DVSS.n10012 DVSS.n9809 0.0380882
R47981 DVSS.n10013 DVSS.n10012 0.0380882
R47982 DVSS.n10014 DVSS.n10013 0.0380882
R47983 DVSS.n10014 DVSS.n9805 0.0380882
R47984 DVSS.n10024 DVSS.n9805 0.0380882
R47985 DVSS.n10025 DVSS.n10024 0.0380882
R47986 DVSS.n10026 DVSS.n10025 0.0380882
R47987 DVSS.n10026 DVSS.n9801 0.0380882
R47988 DVSS.n10036 DVSS.n9801 0.0380882
R47989 DVSS.n10037 DVSS.n10036 0.0380882
R47990 DVSS.n10038 DVSS.n10037 0.0380882
R47991 DVSS.n10038 DVSS.n9797 0.0380882
R47992 DVSS.n10048 DVSS.n9797 0.0380882
R47993 DVSS.n10049 DVSS.n10048 0.0380882
R47994 DVSS.n10050 DVSS.n10049 0.0380882
R47995 DVSS.n10050 DVSS.n9793 0.0380882
R47996 DVSS.n10060 DVSS.n9793 0.0380882
R47997 DVSS.n10061 DVSS.n10060 0.0380882
R47998 DVSS.n10062 DVSS.n10061 0.0380882
R47999 DVSS.n10062 DVSS.n9789 0.0380882
R48000 DVSS.n10072 DVSS.n9789 0.0380882
R48001 DVSS.n10073 DVSS.n10072 0.0380882
R48002 DVSS.n10074 DVSS.n10073 0.0380882
R48003 DVSS.n10074 DVSS.n9785 0.0380882
R48004 DVSS.n10084 DVSS.n9785 0.0380882
R48005 DVSS.n10085 DVSS.n10084 0.0380882
R48006 DVSS.n10086 DVSS.n10085 0.0380882
R48007 DVSS.n10086 DVSS.n9781 0.0380882
R48008 DVSS.n10096 DVSS.n9781 0.0380882
R48009 DVSS.n10097 DVSS.n10096 0.0380882
R48010 DVSS.n10099 DVSS.n10097 0.0380882
R48011 DVSS.n10099 DVSS.n10098 0.0380882
R48012 DVSS.n10098 DVSS.n9776 0.0380882
R48013 DVSS.n10109 DVSS.n9776 0.0380882
R48014 DVSS.n9859 DVSS.n9858 0.0380882
R48015 DVSS.n9867 DVSS.n9858 0.0380882
R48016 DVSS.n9867 DVSS.n9856 0.0380882
R48017 DVSS.n9871 DVSS.n9856 0.0380882
R48018 DVSS.n9871 DVSS.n9854 0.0380882
R48019 DVSS.n9879 DVSS.n9854 0.0380882
R48020 DVSS.n9879 DVSS.n9852 0.0380882
R48021 DVSS.n9883 DVSS.n9852 0.0380882
R48022 DVSS.n9883 DVSS.n9850 0.0380882
R48023 DVSS.n9891 DVSS.n9850 0.0380882
R48024 DVSS.n9891 DVSS.n9848 0.0380882
R48025 DVSS.n9895 DVSS.n9848 0.0380882
R48026 DVSS.n9895 DVSS.n9846 0.0380882
R48027 DVSS.n9903 DVSS.n9846 0.0380882
R48028 DVSS.n9903 DVSS.n9844 0.0380882
R48029 DVSS.n9907 DVSS.n9844 0.0380882
R48030 DVSS.n9907 DVSS.n9842 0.0380882
R48031 DVSS.n9915 DVSS.n9842 0.0380882
R48032 DVSS.n9915 DVSS.n9840 0.0380882
R48033 DVSS.n9919 DVSS.n9840 0.0380882
R48034 DVSS.n9919 DVSS.n9838 0.0380882
R48035 DVSS.n9927 DVSS.n9838 0.0380882
R48036 DVSS.n9927 DVSS.n9836 0.0380882
R48037 DVSS.n9931 DVSS.n9836 0.0380882
R48038 DVSS.n9931 DVSS.n9834 0.0380882
R48039 DVSS.n9939 DVSS.n9834 0.0380882
R48040 DVSS.n9939 DVSS.n9832 0.0380882
R48041 DVSS.n9943 DVSS.n9832 0.0380882
R48042 DVSS.n9943 DVSS.n9830 0.0380882
R48043 DVSS.n9951 DVSS.n9830 0.0380882
R48044 DVSS.n9951 DVSS.n9828 0.0380882
R48045 DVSS.n9955 DVSS.n9828 0.0380882
R48046 DVSS.n9955 DVSS.n9826 0.0380882
R48047 DVSS.n9963 DVSS.n9826 0.0380882
R48048 DVSS.n9963 DVSS.n9824 0.0380882
R48049 DVSS.n9967 DVSS.n9824 0.0380882
R48050 DVSS.n9967 DVSS.n9822 0.0380882
R48051 DVSS.n9975 DVSS.n9822 0.0380882
R48052 DVSS.n9975 DVSS.n9820 0.0380882
R48053 DVSS.n9979 DVSS.n9820 0.0380882
R48054 DVSS.n9979 DVSS.n9818 0.0380882
R48055 DVSS.n9987 DVSS.n9818 0.0380882
R48056 DVSS.n9987 DVSS.n9816 0.0380882
R48057 DVSS.n9991 DVSS.n9816 0.0380882
R48058 DVSS.n9991 DVSS.n9814 0.0380882
R48059 DVSS.n9999 DVSS.n9814 0.0380882
R48060 DVSS.n9999 DVSS.n9812 0.0380882
R48061 DVSS.n10003 DVSS.n9812 0.0380882
R48062 DVSS.n10003 DVSS.n9810 0.0380882
R48063 DVSS.n10011 DVSS.n9810 0.0380882
R48064 DVSS.n10011 DVSS.n9808 0.0380882
R48065 DVSS.n10015 DVSS.n9808 0.0380882
R48066 DVSS.n10015 DVSS.n9806 0.0380882
R48067 DVSS.n10023 DVSS.n9806 0.0380882
R48068 DVSS.n10023 DVSS.n9804 0.0380882
R48069 DVSS.n10027 DVSS.n9804 0.0380882
R48070 DVSS.n10027 DVSS.n9802 0.0380882
R48071 DVSS.n10035 DVSS.n9802 0.0380882
R48072 DVSS.n10035 DVSS.n9800 0.0380882
R48073 DVSS.n10039 DVSS.n9800 0.0380882
R48074 DVSS.n10039 DVSS.n9798 0.0380882
R48075 DVSS.n10047 DVSS.n9798 0.0380882
R48076 DVSS.n10047 DVSS.n9796 0.0380882
R48077 DVSS.n10051 DVSS.n9796 0.0380882
R48078 DVSS.n10051 DVSS.n9794 0.0380882
R48079 DVSS.n10059 DVSS.n9794 0.0380882
R48080 DVSS.n10059 DVSS.n9792 0.0380882
R48081 DVSS.n10063 DVSS.n9792 0.0380882
R48082 DVSS.n10063 DVSS.n9790 0.0380882
R48083 DVSS.n10071 DVSS.n9790 0.0380882
R48084 DVSS.n10071 DVSS.n9788 0.0380882
R48085 DVSS.n10075 DVSS.n9788 0.0380882
R48086 DVSS.n10075 DVSS.n9786 0.0380882
R48087 DVSS.n10083 DVSS.n9786 0.0380882
R48088 DVSS.n10083 DVSS.n9784 0.0380882
R48089 DVSS.n10087 DVSS.n9784 0.0380882
R48090 DVSS.n10087 DVSS.n9782 0.0380882
R48091 DVSS.n10095 DVSS.n9782 0.0380882
R48092 DVSS.n10095 DVSS.n9780 0.0380882
R48093 DVSS.n10100 DVSS.n9780 0.0380882
R48094 DVSS.n10100 DVSS.n9778 0.0380882
R48095 DVSS.n9778 DVSS.n9777 0.0380882
R48096 DVSS.n10108 DVSS.n9777 0.0380882
R48097 DVSS.n2461 DVSS.n2460 0.0380882
R48098 DVSS.n2462 DVSS.n2461 0.0380882
R48099 DVSS.n2462 DVSS.n2455 0.0380882
R48100 DVSS.n2472 DVSS.n2455 0.0380882
R48101 DVSS.n2473 DVSS.n2472 0.0380882
R48102 DVSS.n2474 DVSS.n2473 0.0380882
R48103 DVSS.n2474 DVSS.n2453 0.0380882
R48104 DVSS.n2484 DVSS.n2453 0.0380882
R48105 DVSS.n2485 DVSS.n2484 0.0380882
R48106 DVSS.n2486 DVSS.n2485 0.0380882
R48107 DVSS.n2486 DVSS.n2451 0.0380882
R48108 DVSS.n2496 DVSS.n2451 0.0380882
R48109 DVSS.n2497 DVSS.n2496 0.0380882
R48110 DVSS.n2498 DVSS.n2497 0.0380882
R48111 DVSS.n2498 DVSS.n2449 0.0380882
R48112 DVSS.n2508 DVSS.n2449 0.0380882
R48113 DVSS.n2509 DVSS.n2508 0.0380882
R48114 DVSS.n2510 DVSS.n2509 0.0380882
R48115 DVSS.n2510 DVSS.n2447 0.0380882
R48116 DVSS.n2520 DVSS.n2447 0.0380882
R48117 DVSS.n2521 DVSS.n2520 0.0380882
R48118 DVSS.n2522 DVSS.n2521 0.0380882
R48119 DVSS.n2522 DVSS.n2445 0.0380882
R48120 DVSS.n2532 DVSS.n2445 0.0380882
R48121 DVSS.n2533 DVSS.n2532 0.0380882
R48122 DVSS.n2534 DVSS.n2533 0.0380882
R48123 DVSS.n2534 DVSS.n2443 0.0380882
R48124 DVSS.n2544 DVSS.n2443 0.0380882
R48125 DVSS.n2545 DVSS.n2544 0.0380882
R48126 DVSS.n2546 DVSS.n2545 0.0380882
R48127 DVSS.n2546 DVSS.n2441 0.0380882
R48128 DVSS.n2556 DVSS.n2441 0.0380882
R48129 DVSS.n2557 DVSS.n2556 0.0380882
R48130 DVSS.n2558 DVSS.n2557 0.0380882
R48131 DVSS.n2558 DVSS.n2439 0.0380882
R48132 DVSS.n2568 DVSS.n2439 0.0380882
R48133 DVSS.n2569 DVSS.n2568 0.0380882
R48134 DVSS.n2570 DVSS.n2569 0.0380882
R48135 DVSS.n2570 DVSS.n2437 0.0380882
R48136 DVSS.n2580 DVSS.n2437 0.0380882
R48137 DVSS.n2581 DVSS.n2580 0.0380882
R48138 DVSS.n2582 DVSS.n2581 0.0380882
R48139 DVSS.n2582 DVSS.n2435 0.0380882
R48140 DVSS.n2592 DVSS.n2435 0.0380882
R48141 DVSS.n2593 DVSS.n2592 0.0380882
R48142 DVSS.n2594 DVSS.n2593 0.0380882
R48143 DVSS.n2594 DVSS.n2433 0.0380882
R48144 DVSS.n2604 DVSS.n2433 0.0380882
R48145 DVSS.n2605 DVSS.n2604 0.0380882
R48146 DVSS.n2606 DVSS.n2605 0.0380882
R48147 DVSS.n2606 DVSS.n2431 0.0380882
R48148 DVSS.n2616 DVSS.n2431 0.0380882
R48149 DVSS.n2617 DVSS.n2616 0.0380882
R48150 DVSS.n2618 DVSS.n2617 0.0380882
R48151 DVSS.n2618 DVSS.n2429 0.0380882
R48152 DVSS.n2628 DVSS.n2429 0.0380882
R48153 DVSS.n2629 DVSS.n2628 0.0380882
R48154 DVSS.n2630 DVSS.n2629 0.0380882
R48155 DVSS.n2630 DVSS.n2427 0.0380882
R48156 DVSS.n2640 DVSS.n2427 0.0380882
R48157 DVSS.n2641 DVSS.n2640 0.0380882
R48158 DVSS.n2642 DVSS.n2641 0.0380882
R48159 DVSS.n2642 DVSS.n2425 0.0380882
R48160 DVSS.n2652 DVSS.n2425 0.0380882
R48161 DVSS.n2653 DVSS.n2652 0.0380882
R48162 DVSS.n2654 DVSS.n2653 0.0380882
R48163 DVSS.n2654 DVSS.n2423 0.0380882
R48164 DVSS.n2664 DVSS.n2423 0.0380882
R48165 DVSS.n2665 DVSS.n2664 0.0380882
R48166 DVSS.n2666 DVSS.n2665 0.0380882
R48167 DVSS.n2666 DVSS.n2421 0.0380882
R48168 DVSS.n2676 DVSS.n2421 0.0380882
R48169 DVSS.n2677 DVSS.n2676 0.0380882
R48170 DVSS.n2678 DVSS.n2677 0.0380882
R48171 DVSS.n2678 DVSS.n2419 0.0380882
R48172 DVSS.n2688 DVSS.n2419 0.0380882
R48173 DVSS.n2689 DVSS.n2688 0.0380882
R48174 DVSS.n2690 DVSS.n2689 0.0380882
R48175 DVSS.n2690 DVSS.n2417 0.0380882
R48176 DVSS.n2700 DVSS.n2417 0.0380882
R48177 DVSS.n2701 DVSS.n2700 0.0380882
R48178 DVSS.n10136 DVSS.n2701 0.0380882
R48179 DVSS.n10136 DVSS.n10135 0.0380882
R48180 DVSS.n2459 DVSS.n2458 0.0380882
R48181 DVSS.n2463 DVSS.n2458 0.0380882
R48182 DVSS.n2467 DVSS.n2463 0.0380882
R48183 DVSS.n2471 DVSS.n2467 0.0380882
R48184 DVSS.n2471 DVSS.n2454 0.0380882
R48185 DVSS.n2475 DVSS.n2454 0.0380882
R48186 DVSS.n2479 DVSS.n2475 0.0380882
R48187 DVSS.n2483 DVSS.n2479 0.0380882
R48188 DVSS.n2483 DVSS.n2452 0.0380882
R48189 DVSS.n2487 DVSS.n2452 0.0380882
R48190 DVSS.n2491 DVSS.n2487 0.0380882
R48191 DVSS.n2495 DVSS.n2491 0.0380882
R48192 DVSS.n2495 DVSS.n2450 0.0380882
R48193 DVSS.n2499 DVSS.n2450 0.0380882
R48194 DVSS.n2503 DVSS.n2499 0.0380882
R48195 DVSS.n2507 DVSS.n2503 0.0380882
R48196 DVSS.n2507 DVSS.n2448 0.0380882
R48197 DVSS.n2511 DVSS.n2448 0.0380882
R48198 DVSS.n2515 DVSS.n2511 0.0380882
R48199 DVSS.n2519 DVSS.n2515 0.0380882
R48200 DVSS.n2519 DVSS.n2446 0.0380882
R48201 DVSS.n2523 DVSS.n2446 0.0380882
R48202 DVSS.n2527 DVSS.n2523 0.0380882
R48203 DVSS.n2531 DVSS.n2527 0.0380882
R48204 DVSS.n2531 DVSS.n2444 0.0380882
R48205 DVSS.n2535 DVSS.n2444 0.0380882
R48206 DVSS.n2539 DVSS.n2535 0.0380882
R48207 DVSS.n2543 DVSS.n2539 0.0380882
R48208 DVSS.n2543 DVSS.n2442 0.0380882
R48209 DVSS.n2547 DVSS.n2442 0.0380882
R48210 DVSS.n2551 DVSS.n2547 0.0380882
R48211 DVSS.n2555 DVSS.n2551 0.0380882
R48212 DVSS.n2555 DVSS.n2440 0.0380882
R48213 DVSS.n2559 DVSS.n2440 0.0380882
R48214 DVSS.n2563 DVSS.n2559 0.0380882
R48215 DVSS.n2567 DVSS.n2563 0.0380882
R48216 DVSS.n2567 DVSS.n2438 0.0380882
R48217 DVSS.n2571 DVSS.n2438 0.0380882
R48218 DVSS.n2575 DVSS.n2571 0.0380882
R48219 DVSS.n2579 DVSS.n2575 0.0380882
R48220 DVSS.n2579 DVSS.n2436 0.0380882
R48221 DVSS.n2583 DVSS.n2436 0.0380882
R48222 DVSS.n2587 DVSS.n2583 0.0380882
R48223 DVSS.n2591 DVSS.n2587 0.0380882
R48224 DVSS.n2591 DVSS.n2434 0.0380882
R48225 DVSS.n2595 DVSS.n2434 0.0380882
R48226 DVSS.n2599 DVSS.n2595 0.0380882
R48227 DVSS.n2603 DVSS.n2599 0.0380882
R48228 DVSS.n2603 DVSS.n2432 0.0380882
R48229 DVSS.n2607 DVSS.n2432 0.0380882
R48230 DVSS.n2611 DVSS.n2607 0.0380882
R48231 DVSS.n2615 DVSS.n2611 0.0380882
R48232 DVSS.n2615 DVSS.n2430 0.0380882
R48233 DVSS.n2619 DVSS.n2430 0.0380882
R48234 DVSS.n2623 DVSS.n2619 0.0380882
R48235 DVSS.n2627 DVSS.n2623 0.0380882
R48236 DVSS.n2627 DVSS.n2428 0.0380882
R48237 DVSS.n2631 DVSS.n2428 0.0380882
R48238 DVSS.n2635 DVSS.n2631 0.0380882
R48239 DVSS.n2639 DVSS.n2635 0.0380882
R48240 DVSS.n2639 DVSS.n2426 0.0380882
R48241 DVSS.n2643 DVSS.n2426 0.0380882
R48242 DVSS.n2647 DVSS.n2643 0.0380882
R48243 DVSS.n2651 DVSS.n2647 0.0380882
R48244 DVSS.n2651 DVSS.n2424 0.0380882
R48245 DVSS.n2655 DVSS.n2424 0.0380882
R48246 DVSS.n2659 DVSS.n2655 0.0380882
R48247 DVSS.n2663 DVSS.n2659 0.0380882
R48248 DVSS.n2663 DVSS.n2422 0.0380882
R48249 DVSS.n2667 DVSS.n2422 0.0380882
R48250 DVSS.n2671 DVSS.n2667 0.0380882
R48251 DVSS.n2675 DVSS.n2671 0.0380882
R48252 DVSS.n2675 DVSS.n2420 0.0380882
R48253 DVSS.n2679 DVSS.n2420 0.0380882
R48254 DVSS.n2683 DVSS.n2679 0.0380882
R48255 DVSS.n2687 DVSS.n2683 0.0380882
R48256 DVSS.n2687 DVSS.n2418 0.0380882
R48257 DVSS.n2691 DVSS.n2418 0.0380882
R48258 DVSS.n2695 DVSS.n2691 0.0380882
R48259 DVSS.n2699 DVSS.n2695 0.0380882
R48260 DVSS.n2699 DVSS.n2416 0.0380882
R48261 DVSS.n10137 DVSS.n2416 0.0380882
R48262 DVSS.n10137 DVSS.n2414 0.0380882
R48263 DVSS.n2119 DVSS.n2118 0.0380882
R48264 DVSS.n2120 DVSS.n2119 0.0380882
R48265 DVSS.n2120 DVSS.n2113 0.0380882
R48266 DVSS.n2130 DVSS.n2113 0.0380882
R48267 DVSS.n2131 DVSS.n2130 0.0380882
R48268 DVSS.n2132 DVSS.n2131 0.0380882
R48269 DVSS.n2132 DVSS.n2111 0.0380882
R48270 DVSS.n2142 DVSS.n2111 0.0380882
R48271 DVSS.n2143 DVSS.n2142 0.0380882
R48272 DVSS.n2144 DVSS.n2143 0.0380882
R48273 DVSS.n2144 DVSS.n2109 0.0380882
R48274 DVSS.n2154 DVSS.n2109 0.0380882
R48275 DVSS.n2155 DVSS.n2154 0.0380882
R48276 DVSS.n2156 DVSS.n2155 0.0380882
R48277 DVSS.n2156 DVSS.n2107 0.0380882
R48278 DVSS.n2166 DVSS.n2107 0.0380882
R48279 DVSS.n2167 DVSS.n2166 0.0380882
R48280 DVSS.n2168 DVSS.n2167 0.0380882
R48281 DVSS.n2168 DVSS.n2105 0.0380882
R48282 DVSS.n2178 DVSS.n2105 0.0380882
R48283 DVSS.n2179 DVSS.n2178 0.0380882
R48284 DVSS.n2180 DVSS.n2179 0.0380882
R48285 DVSS.n2180 DVSS.n2103 0.0380882
R48286 DVSS.n2190 DVSS.n2103 0.0380882
R48287 DVSS.n2191 DVSS.n2190 0.0380882
R48288 DVSS.n2192 DVSS.n2191 0.0380882
R48289 DVSS.n2192 DVSS.n2101 0.0380882
R48290 DVSS.n2202 DVSS.n2101 0.0380882
R48291 DVSS.n2203 DVSS.n2202 0.0380882
R48292 DVSS.n2204 DVSS.n2203 0.0380882
R48293 DVSS.n2204 DVSS.n2099 0.0380882
R48294 DVSS.n2214 DVSS.n2099 0.0380882
R48295 DVSS.n2215 DVSS.n2214 0.0380882
R48296 DVSS.n2216 DVSS.n2215 0.0380882
R48297 DVSS.n2216 DVSS.n2097 0.0380882
R48298 DVSS.n2226 DVSS.n2097 0.0380882
R48299 DVSS.n2227 DVSS.n2226 0.0380882
R48300 DVSS.n2228 DVSS.n2227 0.0380882
R48301 DVSS.n2228 DVSS.n2095 0.0380882
R48302 DVSS.n2238 DVSS.n2095 0.0380882
R48303 DVSS.n2239 DVSS.n2238 0.0380882
R48304 DVSS.n2240 DVSS.n2239 0.0380882
R48305 DVSS.n2240 DVSS.n2093 0.0380882
R48306 DVSS.n2250 DVSS.n2093 0.0380882
R48307 DVSS.n2251 DVSS.n2250 0.0380882
R48308 DVSS.n2252 DVSS.n2251 0.0380882
R48309 DVSS.n2252 DVSS.n2091 0.0380882
R48310 DVSS.n2262 DVSS.n2091 0.0380882
R48311 DVSS.n2263 DVSS.n2262 0.0380882
R48312 DVSS.n2264 DVSS.n2263 0.0380882
R48313 DVSS.n2264 DVSS.n2089 0.0380882
R48314 DVSS.n2274 DVSS.n2089 0.0380882
R48315 DVSS.n2275 DVSS.n2274 0.0380882
R48316 DVSS.n2276 DVSS.n2275 0.0380882
R48317 DVSS.n2276 DVSS.n2087 0.0380882
R48318 DVSS.n2286 DVSS.n2087 0.0380882
R48319 DVSS.n2287 DVSS.n2286 0.0380882
R48320 DVSS.n2288 DVSS.n2287 0.0380882
R48321 DVSS.n2288 DVSS.n2085 0.0380882
R48322 DVSS.n2298 DVSS.n2085 0.0380882
R48323 DVSS.n2299 DVSS.n2298 0.0380882
R48324 DVSS.n2300 DVSS.n2299 0.0380882
R48325 DVSS.n2300 DVSS.n2083 0.0380882
R48326 DVSS.n2310 DVSS.n2083 0.0380882
R48327 DVSS.n2311 DVSS.n2310 0.0380882
R48328 DVSS.n2312 DVSS.n2311 0.0380882
R48329 DVSS.n2312 DVSS.n2081 0.0380882
R48330 DVSS.n2322 DVSS.n2081 0.0380882
R48331 DVSS.n2323 DVSS.n2322 0.0380882
R48332 DVSS.n2324 DVSS.n2323 0.0380882
R48333 DVSS.n2324 DVSS.n2079 0.0380882
R48334 DVSS.n2334 DVSS.n2079 0.0380882
R48335 DVSS.n2335 DVSS.n2334 0.0380882
R48336 DVSS.n2336 DVSS.n2335 0.0380882
R48337 DVSS.n2336 DVSS.n2077 0.0380882
R48338 DVSS.n2346 DVSS.n2077 0.0380882
R48339 DVSS.n2347 DVSS.n2346 0.0380882
R48340 DVSS.n2348 DVSS.n2347 0.0380882
R48341 DVSS.n2348 DVSS.n2075 0.0380882
R48342 DVSS.n2358 DVSS.n2075 0.0380882
R48343 DVSS.n2359 DVSS.n2358 0.0380882
R48344 DVSS.n10161 DVSS.n2359 0.0380882
R48345 DVSS.n10161 DVSS.n10160 0.0380882
R48346 DVSS.n2117 DVSS.n2116 0.0380882
R48347 DVSS.n2121 DVSS.n2116 0.0380882
R48348 DVSS.n2125 DVSS.n2121 0.0380882
R48349 DVSS.n2129 DVSS.n2125 0.0380882
R48350 DVSS.n2129 DVSS.n2112 0.0380882
R48351 DVSS.n2133 DVSS.n2112 0.0380882
R48352 DVSS.n2137 DVSS.n2133 0.0380882
R48353 DVSS.n2141 DVSS.n2137 0.0380882
R48354 DVSS.n2141 DVSS.n2110 0.0380882
R48355 DVSS.n2145 DVSS.n2110 0.0380882
R48356 DVSS.n2149 DVSS.n2145 0.0380882
R48357 DVSS.n2153 DVSS.n2149 0.0380882
R48358 DVSS.n2153 DVSS.n2108 0.0380882
R48359 DVSS.n2157 DVSS.n2108 0.0380882
R48360 DVSS.n2161 DVSS.n2157 0.0380882
R48361 DVSS.n2165 DVSS.n2161 0.0380882
R48362 DVSS.n2165 DVSS.n2106 0.0380882
R48363 DVSS.n2169 DVSS.n2106 0.0380882
R48364 DVSS.n2173 DVSS.n2169 0.0380882
R48365 DVSS.n2177 DVSS.n2173 0.0380882
R48366 DVSS.n2177 DVSS.n2104 0.0380882
R48367 DVSS.n2181 DVSS.n2104 0.0380882
R48368 DVSS.n2185 DVSS.n2181 0.0380882
R48369 DVSS.n2189 DVSS.n2185 0.0380882
R48370 DVSS.n2189 DVSS.n2102 0.0380882
R48371 DVSS.n2193 DVSS.n2102 0.0380882
R48372 DVSS.n2197 DVSS.n2193 0.0380882
R48373 DVSS.n2201 DVSS.n2197 0.0380882
R48374 DVSS.n2201 DVSS.n2100 0.0380882
R48375 DVSS.n2205 DVSS.n2100 0.0380882
R48376 DVSS.n2209 DVSS.n2205 0.0380882
R48377 DVSS.n2213 DVSS.n2209 0.0380882
R48378 DVSS.n2213 DVSS.n2098 0.0380882
R48379 DVSS.n2217 DVSS.n2098 0.0380882
R48380 DVSS.n2221 DVSS.n2217 0.0380882
R48381 DVSS.n2225 DVSS.n2221 0.0380882
R48382 DVSS.n2225 DVSS.n2096 0.0380882
R48383 DVSS.n2229 DVSS.n2096 0.0380882
R48384 DVSS.n2233 DVSS.n2229 0.0380882
R48385 DVSS.n2237 DVSS.n2233 0.0380882
R48386 DVSS.n2237 DVSS.n2094 0.0380882
R48387 DVSS.n2241 DVSS.n2094 0.0380882
R48388 DVSS.n2245 DVSS.n2241 0.0380882
R48389 DVSS.n2249 DVSS.n2245 0.0380882
R48390 DVSS.n2249 DVSS.n2092 0.0380882
R48391 DVSS.n2253 DVSS.n2092 0.0380882
R48392 DVSS.n2257 DVSS.n2253 0.0380882
R48393 DVSS.n2261 DVSS.n2257 0.0380882
R48394 DVSS.n2261 DVSS.n2090 0.0380882
R48395 DVSS.n2265 DVSS.n2090 0.0380882
R48396 DVSS.n2269 DVSS.n2265 0.0380882
R48397 DVSS.n2273 DVSS.n2269 0.0380882
R48398 DVSS.n2273 DVSS.n2088 0.0380882
R48399 DVSS.n2277 DVSS.n2088 0.0380882
R48400 DVSS.n2281 DVSS.n2277 0.0380882
R48401 DVSS.n2285 DVSS.n2281 0.0380882
R48402 DVSS.n2285 DVSS.n2086 0.0380882
R48403 DVSS.n2289 DVSS.n2086 0.0380882
R48404 DVSS.n2293 DVSS.n2289 0.0380882
R48405 DVSS.n2297 DVSS.n2293 0.0380882
R48406 DVSS.n2297 DVSS.n2084 0.0380882
R48407 DVSS.n2301 DVSS.n2084 0.0380882
R48408 DVSS.n2305 DVSS.n2301 0.0380882
R48409 DVSS.n2309 DVSS.n2305 0.0380882
R48410 DVSS.n2309 DVSS.n2082 0.0380882
R48411 DVSS.n2313 DVSS.n2082 0.0380882
R48412 DVSS.n2317 DVSS.n2313 0.0380882
R48413 DVSS.n2321 DVSS.n2317 0.0380882
R48414 DVSS.n2321 DVSS.n2080 0.0380882
R48415 DVSS.n2325 DVSS.n2080 0.0380882
R48416 DVSS.n2329 DVSS.n2325 0.0380882
R48417 DVSS.n2333 DVSS.n2329 0.0380882
R48418 DVSS.n2333 DVSS.n2078 0.0380882
R48419 DVSS.n2337 DVSS.n2078 0.0380882
R48420 DVSS.n2341 DVSS.n2337 0.0380882
R48421 DVSS.n2345 DVSS.n2341 0.0380882
R48422 DVSS.n2345 DVSS.n2076 0.0380882
R48423 DVSS.n2349 DVSS.n2076 0.0380882
R48424 DVSS.n2353 DVSS.n2349 0.0380882
R48425 DVSS.n2357 DVSS.n2353 0.0380882
R48426 DVSS.n2357 DVSS.n2074 0.0380882
R48427 DVSS.n10162 DVSS.n2074 0.0380882
R48428 DVSS.n10162 DVSS.n2072 0.0380882
R48429 DVSS.n10455 DVSS.n10172 0.0380882
R48430 DVSS.n10446 DVSS.n10172 0.0380882
R48431 DVSS.n10446 DVSS.n10445 0.0380882
R48432 DVSS.n10445 DVSS.n10444 0.0380882
R48433 DVSS.n10444 DVSS.n10174 0.0380882
R48434 DVSS.n10434 DVSS.n10174 0.0380882
R48435 DVSS.n10434 DVSS.n10433 0.0380882
R48436 DVSS.n10433 DVSS.n10432 0.0380882
R48437 DVSS.n10432 DVSS.n10176 0.0380882
R48438 DVSS.n10422 DVSS.n10176 0.0380882
R48439 DVSS.n10422 DVSS.n10421 0.0380882
R48440 DVSS.n10421 DVSS.n10420 0.0380882
R48441 DVSS.n10420 DVSS.n10178 0.0380882
R48442 DVSS.n10410 DVSS.n10178 0.0380882
R48443 DVSS.n10410 DVSS.n10409 0.0380882
R48444 DVSS.n10409 DVSS.n10408 0.0380882
R48445 DVSS.n10408 DVSS.n10180 0.0380882
R48446 DVSS.n10398 DVSS.n10180 0.0380882
R48447 DVSS.n10398 DVSS.n10397 0.0380882
R48448 DVSS.n10397 DVSS.n10396 0.0380882
R48449 DVSS.n10396 DVSS.n10182 0.0380882
R48450 DVSS.n10386 DVSS.n10182 0.0380882
R48451 DVSS.n10386 DVSS.n10385 0.0380882
R48452 DVSS.n10385 DVSS.n10384 0.0380882
R48453 DVSS.n10384 DVSS.n10184 0.0380882
R48454 DVSS.n10374 DVSS.n10184 0.0380882
R48455 DVSS.n10374 DVSS.n10373 0.0380882
R48456 DVSS.n10373 DVSS.n10372 0.0380882
R48457 DVSS.n10372 DVSS.n10186 0.0380882
R48458 DVSS.n10362 DVSS.n10186 0.0380882
R48459 DVSS.n10362 DVSS.n10361 0.0380882
R48460 DVSS.n10361 DVSS.n10360 0.0380882
R48461 DVSS.n10360 DVSS.n10188 0.0380882
R48462 DVSS.n10350 DVSS.n10188 0.0380882
R48463 DVSS.n10350 DVSS.n10349 0.0380882
R48464 DVSS.n10349 DVSS.n10348 0.0380882
R48465 DVSS.n10348 DVSS.n10190 0.0380882
R48466 DVSS.n10338 DVSS.n10190 0.0380882
R48467 DVSS.n10338 DVSS.n10337 0.0380882
R48468 DVSS.n10337 DVSS.n10336 0.0380882
R48469 DVSS.n10336 DVSS.n10192 0.0380882
R48470 DVSS.n10326 DVSS.n10192 0.0380882
R48471 DVSS.n10326 DVSS.n10325 0.0380882
R48472 DVSS.n10325 DVSS.n10324 0.0380882
R48473 DVSS.n10324 DVSS.n10194 0.0380882
R48474 DVSS.n10314 DVSS.n10194 0.0380882
R48475 DVSS.n10314 DVSS.n10313 0.0380882
R48476 DVSS.n10313 DVSS.n10312 0.0380882
R48477 DVSS.n10312 DVSS.n10196 0.0380882
R48478 DVSS.n10302 DVSS.n10196 0.0380882
R48479 DVSS.n10302 DVSS.n10301 0.0380882
R48480 DVSS.n10301 DVSS.n10300 0.0380882
R48481 DVSS.n10300 DVSS.n10198 0.0380882
R48482 DVSS.n10290 DVSS.n10198 0.0380882
R48483 DVSS.n10290 DVSS.n10289 0.0380882
R48484 DVSS.n10289 DVSS.n10288 0.0380882
R48485 DVSS.n10288 DVSS.n10200 0.0380882
R48486 DVSS.n10278 DVSS.n10200 0.0380882
R48487 DVSS.n10278 DVSS.n10277 0.0380882
R48488 DVSS.n10277 DVSS.n10276 0.0380882
R48489 DVSS.n10276 DVSS.n10202 0.0380882
R48490 DVSS.n10266 DVSS.n10202 0.0380882
R48491 DVSS.n10266 DVSS.n10265 0.0380882
R48492 DVSS.n10265 DVSS.n10264 0.0380882
R48493 DVSS.n10264 DVSS.n10204 0.0380882
R48494 DVSS.n10254 DVSS.n10204 0.0380882
R48495 DVSS.n10254 DVSS.n10253 0.0380882
R48496 DVSS.n10253 DVSS.n10252 0.0380882
R48497 DVSS.n10252 DVSS.n10206 0.0380882
R48498 DVSS.n10242 DVSS.n10206 0.0380882
R48499 DVSS.n10242 DVSS.n10241 0.0380882
R48500 DVSS.n10241 DVSS.n10240 0.0380882
R48501 DVSS.n10240 DVSS.n10208 0.0380882
R48502 DVSS.n10230 DVSS.n10208 0.0380882
R48503 DVSS.n10230 DVSS.n10229 0.0380882
R48504 DVSS.n10229 DVSS.n10228 0.0380882
R48505 DVSS.n10228 DVSS.n10210 0.0380882
R48506 DVSS.n10218 DVSS.n10210 0.0380882
R48507 DVSS.n10218 DVSS.n10217 0.0380882
R48508 DVSS.n10217 DVSS.n10216 0.0380882
R48509 DVSS.n10216 DVSS.n2015 0.0380882
R48510 DVSS.n10470 DVSS.n2015 0.0380882
R48511 DVSS.n10470 DVSS.n10469 0.0380882
R48512 DVSS.n10454 DVSS.n10453 0.0380882
R48513 DVSS.n10453 DVSS.n10450 0.0380882
R48514 DVSS.n10450 DVSS.n10173 0.0380882
R48515 DVSS.n10443 DVSS.n10173 0.0380882
R48516 DVSS.n10443 DVSS.n10439 0.0380882
R48517 DVSS.n10439 DVSS.n10438 0.0380882
R48518 DVSS.n10438 DVSS.n10175 0.0380882
R48519 DVSS.n10431 DVSS.n10175 0.0380882
R48520 DVSS.n10431 DVSS.n10427 0.0380882
R48521 DVSS.n10427 DVSS.n10426 0.0380882
R48522 DVSS.n10426 DVSS.n10177 0.0380882
R48523 DVSS.n10419 DVSS.n10177 0.0380882
R48524 DVSS.n10419 DVSS.n10415 0.0380882
R48525 DVSS.n10415 DVSS.n10414 0.0380882
R48526 DVSS.n10414 DVSS.n10179 0.0380882
R48527 DVSS.n10407 DVSS.n10179 0.0380882
R48528 DVSS.n10407 DVSS.n10403 0.0380882
R48529 DVSS.n10403 DVSS.n10402 0.0380882
R48530 DVSS.n10402 DVSS.n10181 0.0380882
R48531 DVSS.n10395 DVSS.n10181 0.0380882
R48532 DVSS.n10395 DVSS.n10391 0.0380882
R48533 DVSS.n10391 DVSS.n10390 0.0380882
R48534 DVSS.n10390 DVSS.n10183 0.0380882
R48535 DVSS.n10383 DVSS.n10183 0.0380882
R48536 DVSS.n10383 DVSS.n10379 0.0380882
R48537 DVSS.n10379 DVSS.n10378 0.0380882
R48538 DVSS.n10378 DVSS.n10185 0.0380882
R48539 DVSS.n10371 DVSS.n10185 0.0380882
R48540 DVSS.n10371 DVSS.n10367 0.0380882
R48541 DVSS.n10367 DVSS.n10366 0.0380882
R48542 DVSS.n10366 DVSS.n10187 0.0380882
R48543 DVSS.n10359 DVSS.n10187 0.0380882
R48544 DVSS.n10359 DVSS.n10355 0.0380882
R48545 DVSS.n10355 DVSS.n10354 0.0380882
R48546 DVSS.n10354 DVSS.n10189 0.0380882
R48547 DVSS.n10347 DVSS.n10189 0.0380882
R48548 DVSS.n10347 DVSS.n10343 0.0380882
R48549 DVSS.n10343 DVSS.n10342 0.0380882
R48550 DVSS.n10342 DVSS.n10191 0.0380882
R48551 DVSS.n10335 DVSS.n10191 0.0380882
R48552 DVSS.n10335 DVSS.n10331 0.0380882
R48553 DVSS.n10331 DVSS.n10330 0.0380882
R48554 DVSS.n10330 DVSS.n10193 0.0380882
R48555 DVSS.n10323 DVSS.n10193 0.0380882
R48556 DVSS.n10323 DVSS.n10319 0.0380882
R48557 DVSS.n10319 DVSS.n10318 0.0380882
R48558 DVSS.n10318 DVSS.n10195 0.0380882
R48559 DVSS.n10311 DVSS.n10195 0.0380882
R48560 DVSS.n10311 DVSS.n10307 0.0380882
R48561 DVSS.n10307 DVSS.n10306 0.0380882
R48562 DVSS.n10306 DVSS.n10197 0.0380882
R48563 DVSS.n10299 DVSS.n10197 0.0380882
R48564 DVSS.n10299 DVSS.n10295 0.0380882
R48565 DVSS.n10295 DVSS.n10294 0.0380882
R48566 DVSS.n10294 DVSS.n10199 0.0380882
R48567 DVSS.n10287 DVSS.n10199 0.0380882
R48568 DVSS.n10287 DVSS.n10283 0.0380882
R48569 DVSS.n10283 DVSS.n10282 0.0380882
R48570 DVSS.n10282 DVSS.n10201 0.0380882
R48571 DVSS.n10275 DVSS.n10201 0.0380882
R48572 DVSS.n10275 DVSS.n10271 0.0380882
R48573 DVSS.n10271 DVSS.n10270 0.0380882
R48574 DVSS.n10270 DVSS.n10203 0.0380882
R48575 DVSS.n10263 DVSS.n10203 0.0380882
R48576 DVSS.n10263 DVSS.n10259 0.0380882
R48577 DVSS.n10259 DVSS.n10258 0.0380882
R48578 DVSS.n10258 DVSS.n10205 0.0380882
R48579 DVSS.n10251 DVSS.n10205 0.0380882
R48580 DVSS.n10251 DVSS.n10247 0.0380882
R48581 DVSS.n10247 DVSS.n10246 0.0380882
R48582 DVSS.n10246 DVSS.n10207 0.0380882
R48583 DVSS.n10239 DVSS.n10207 0.0380882
R48584 DVSS.n10239 DVSS.n10235 0.0380882
R48585 DVSS.n10235 DVSS.n10234 0.0380882
R48586 DVSS.n10234 DVSS.n10209 0.0380882
R48587 DVSS.n10227 DVSS.n10209 0.0380882
R48588 DVSS.n10227 DVSS.n10223 0.0380882
R48589 DVSS.n10223 DVSS.n10222 0.0380882
R48590 DVSS.n10222 DVSS.n10211 0.0380882
R48591 DVSS.n10215 DVSS.n10211 0.0380882
R48592 DVSS.n10215 DVSS.n2014 0.0380882
R48593 DVSS.n10471 DVSS.n2014 0.0380882
R48594 DVSS.n10471 DVSS.n2011 0.0380882
R48595 DVSS.n1956 DVSS.n1669 0.0380882
R48596 DVSS.n1956 DVSS.n1955 0.0380882
R48597 DVSS.n1955 DVSS.n1954 0.0380882
R48598 DVSS.n1954 DVSS.n1673 0.0380882
R48599 DVSS.n1944 DVSS.n1673 0.0380882
R48600 DVSS.n1944 DVSS.n1943 0.0380882
R48601 DVSS.n1943 DVSS.n1942 0.0380882
R48602 DVSS.n1942 DVSS.n1675 0.0380882
R48603 DVSS.n1932 DVSS.n1675 0.0380882
R48604 DVSS.n1932 DVSS.n1931 0.0380882
R48605 DVSS.n1931 DVSS.n1930 0.0380882
R48606 DVSS.n1930 DVSS.n1677 0.0380882
R48607 DVSS.n1920 DVSS.n1677 0.0380882
R48608 DVSS.n1920 DVSS.n1919 0.0380882
R48609 DVSS.n1919 DVSS.n1918 0.0380882
R48610 DVSS.n1918 DVSS.n1679 0.0380882
R48611 DVSS.n1908 DVSS.n1679 0.0380882
R48612 DVSS.n1908 DVSS.n1907 0.0380882
R48613 DVSS.n1907 DVSS.n1906 0.0380882
R48614 DVSS.n1906 DVSS.n1681 0.0380882
R48615 DVSS.n1896 DVSS.n1681 0.0380882
R48616 DVSS.n1896 DVSS.n1895 0.0380882
R48617 DVSS.n1895 DVSS.n1894 0.0380882
R48618 DVSS.n1894 DVSS.n1683 0.0380882
R48619 DVSS.n1884 DVSS.n1683 0.0380882
R48620 DVSS.n1884 DVSS.n1883 0.0380882
R48621 DVSS.n1883 DVSS.n1882 0.0380882
R48622 DVSS.n1882 DVSS.n1685 0.0380882
R48623 DVSS.n1872 DVSS.n1685 0.0380882
R48624 DVSS.n1872 DVSS.n1871 0.0380882
R48625 DVSS.n1871 DVSS.n1870 0.0380882
R48626 DVSS.n1870 DVSS.n1687 0.0380882
R48627 DVSS.n1860 DVSS.n1687 0.0380882
R48628 DVSS.n1860 DVSS.n1859 0.0380882
R48629 DVSS.n1859 DVSS.n1858 0.0380882
R48630 DVSS.n1858 DVSS.n1689 0.0380882
R48631 DVSS.n1848 DVSS.n1689 0.0380882
R48632 DVSS.n1848 DVSS.n1847 0.0380882
R48633 DVSS.n1847 DVSS.n1846 0.0380882
R48634 DVSS.n1846 DVSS.n1691 0.0380882
R48635 DVSS.n1836 DVSS.n1691 0.0380882
R48636 DVSS.n1836 DVSS.n1835 0.0380882
R48637 DVSS.n1835 DVSS.n1834 0.0380882
R48638 DVSS.n1834 DVSS.n1693 0.0380882
R48639 DVSS.n1824 DVSS.n1693 0.0380882
R48640 DVSS.n1824 DVSS.n1823 0.0380882
R48641 DVSS.n1823 DVSS.n1822 0.0380882
R48642 DVSS.n1822 DVSS.n1695 0.0380882
R48643 DVSS.n1812 DVSS.n1695 0.0380882
R48644 DVSS.n1812 DVSS.n1811 0.0380882
R48645 DVSS.n1811 DVSS.n1810 0.0380882
R48646 DVSS.n1810 DVSS.n1697 0.0380882
R48647 DVSS.n1800 DVSS.n1697 0.0380882
R48648 DVSS.n1800 DVSS.n1799 0.0380882
R48649 DVSS.n1799 DVSS.n1798 0.0380882
R48650 DVSS.n1798 DVSS.n1699 0.0380882
R48651 DVSS.n1788 DVSS.n1699 0.0380882
R48652 DVSS.n1788 DVSS.n1787 0.0380882
R48653 DVSS.n1787 DVSS.n1786 0.0380882
R48654 DVSS.n1786 DVSS.n1701 0.0380882
R48655 DVSS.n1776 DVSS.n1701 0.0380882
R48656 DVSS.n1776 DVSS.n1775 0.0380882
R48657 DVSS.n1775 DVSS.n1774 0.0380882
R48658 DVSS.n1774 DVSS.n1703 0.0380882
R48659 DVSS.n1764 DVSS.n1703 0.0380882
R48660 DVSS.n1764 DVSS.n1763 0.0380882
R48661 DVSS.n1763 DVSS.n1762 0.0380882
R48662 DVSS.n1762 DVSS.n1705 0.0380882
R48663 DVSS.n1752 DVSS.n1705 0.0380882
R48664 DVSS.n1752 DVSS.n1751 0.0380882
R48665 DVSS.n1751 DVSS.n1750 0.0380882
R48666 DVSS.n1750 DVSS.n1707 0.0380882
R48667 DVSS.n1740 DVSS.n1707 0.0380882
R48668 DVSS.n1740 DVSS.n1739 0.0380882
R48669 DVSS.n1739 DVSS.n1738 0.0380882
R48670 DVSS.n1738 DVSS.n1709 0.0380882
R48671 DVSS.n1728 DVSS.n1709 0.0380882
R48672 DVSS.n1728 DVSS.n1727 0.0380882
R48673 DVSS.n1727 DVSS.n1726 0.0380882
R48674 DVSS.n1726 DVSS.n1711 0.0380882
R48675 DVSS.n1716 DVSS.n1711 0.0380882
R48676 DVSS.n1716 DVSS.n1715 0.0380882
R48677 DVSS.n1715 DVSS.n1623 0.0380882
R48678 DVSS.n1958 DVSS.n1957 0.0380882
R48679 DVSS.n1957 DVSS.n1672 0.0380882
R48680 DVSS.n1953 DVSS.n1672 0.0380882
R48681 DVSS.n1953 DVSS.n1949 0.0380882
R48682 DVSS.n1949 DVSS.n1948 0.0380882
R48683 DVSS.n1948 DVSS.n1674 0.0380882
R48684 DVSS.n1941 DVSS.n1674 0.0380882
R48685 DVSS.n1941 DVSS.n1937 0.0380882
R48686 DVSS.n1937 DVSS.n1936 0.0380882
R48687 DVSS.n1936 DVSS.n1676 0.0380882
R48688 DVSS.n1929 DVSS.n1676 0.0380882
R48689 DVSS.n1929 DVSS.n1925 0.0380882
R48690 DVSS.n1925 DVSS.n1924 0.0380882
R48691 DVSS.n1924 DVSS.n1678 0.0380882
R48692 DVSS.n1917 DVSS.n1678 0.0380882
R48693 DVSS.n1917 DVSS.n1913 0.0380882
R48694 DVSS.n1913 DVSS.n1912 0.0380882
R48695 DVSS.n1912 DVSS.n1680 0.0380882
R48696 DVSS.n1905 DVSS.n1680 0.0380882
R48697 DVSS.n1905 DVSS.n1901 0.0380882
R48698 DVSS.n1901 DVSS.n1900 0.0380882
R48699 DVSS.n1900 DVSS.n1682 0.0380882
R48700 DVSS.n1893 DVSS.n1682 0.0380882
R48701 DVSS.n1893 DVSS.n1889 0.0380882
R48702 DVSS.n1889 DVSS.n1888 0.0380882
R48703 DVSS.n1888 DVSS.n1684 0.0380882
R48704 DVSS.n1881 DVSS.n1684 0.0380882
R48705 DVSS.n1881 DVSS.n1877 0.0380882
R48706 DVSS.n1877 DVSS.n1876 0.0380882
R48707 DVSS.n1876 DVSS.n1686 0.0380882
R48708 DVSS.n1869 DVSS.n1686 0.0380882
R48709 DVSS.n1869 DVSS.n1865 0.0380882
R48710 DVSS.n1865 DVSS.n1864 0.0380882
R48711 DVSS.n1864 DVSS.n1688 0.0380882
R48712 DVSS.n1857 DVSS.n1688 0.0380882
R48713 DVSS.n1857 DVSS.n1853 0.0380882
R48714 DVSS.n1853 DVSS.n1852 0.0380882
R48715 DVSS.n1852 DVSS.n1690 0.0380882
R48716 DVSS.n1845 DVSS.n1690 0.0380882
R48717 DVSS.n1845 DVSS.n1841 0.0380882
R48718 DVSS.n1841 DVSS.n1840 0.0380882
R48719 DVSS.n1840 DVSS.n1692 0.0380882
R48720 DVSS.n1833 DVSS.n1692 0.0380882
R48721 DVSS.n1833 DVSS.n1829 0.0380882
R48722 DVSS.n1829 DVSS.n1828 0.0380882
R48723 DVSS.n1828 DVSS.n1694 0.0380882
R48724 DVSS.n1821 DVSS.n1694 0.0380882
R48725 DVSS.n1821 DVSS.n1817 0.0380882
R48726 DVSS.n1817 DVSS.n1816 0.0380882
R48727 DVSS.n1816 DVSS.n1696 0.0380882
R48728 DVSS.n1809 DVSS.n1696 0.0380882
R48729 DVSS.n1809 DVSS.n1805 0.0380882
R48730 DVSS.n1805 DVSS.n1804 0.0380882
R48731 DVSS.n1804 DVSS.n1698 0.0380882
R48732 DVSS.n1797 DVSS.n1698 0.0380882
R48733 DVSS.n1797 DVSS.n1793 0.0380882
R48734 DVSS.n1793 DVSS.n1792 0.0380882
R48735 DVSS.n1792 DVSS.n1700 0.0380882
R48736 DVSS.n1785 DVSS.n1700 0.0380882
R48737 DVSS.n1785 DVSS.n1781 0.0380882
R48738 DVSS.n1781 DVSS.n1780 0.0380882
R48739 DVSS.n1780 DVSS.n1702 0.0380882
R48740 DVSS.n1773 DVSS.n1702 0.0380882
R48741 DVSS.n1773 DVSS.n1769 0.0380882
R48742 DVSS.n1769 DVSS.n1768 0.0380882
R48743 DVSS.n1768 DVSS.n1704 0.0380882
R48744 DVSS.n1761 DVSS.n1704 0.0380882
R48745 DVSS.n1761 DVSS.n1757 0.0380882
R48746 DVSS.n1757 DVSS.n1756 0.0380882
R48747 DVSS.n1756 DVSS.n1706 0.0380882
R48748 DVSS.n1749 DVSS.n1706 0.0380882
R48749 DVSS.n1749 DVSS.n1745 0.0380882
R48750 DVSS.n1745 DVSS.n1744 0.0380882
R48751 DVSS.n1744 DVSS.n1708 0.0380882
R48752 DVSS.n1737 DVSS.n1708 0.0380882
R48753 DVSS.n1737 DVSS.n1733 0.0380882
R48754 DVSS.n1733 DVSS.n1732 0.0380882
R48755 DVSS.n1732 DVSS.n1710 0.0380882
R48756 DVSS.n1725 DVSS.n1710 0.0380882
R48757 DVSS.n1725 DVSS.n1721 0.0380882
R48758 DVSS.n1721 DVSS.n1720 0.0380882
R48759 DVSS.n1720 DVSS.n1714 0.0380882
R48760 DVSS.n1714 DVSS.n1713 0.0380882
R48761 DVSS.n10508 DVSS.n10507 0.0380882
R48762 DVSS.n10509 DVSS.n10508 0.0380882
R48763 DVSS.n10509 DVSS.n1608 0.0380882
R48764 DVSS.n10519 DVSS.n1608 0.0380882
R48765 DVSS.n10520 DVSS.n10519 0.0380882
R48766 DVSS.n10521 DVSS.n10520 0.0380882
R48767 DVSS.n10521 DVSS.n1606 0.0380882
R48768 DVSS.n10531 DVSS.n1606 0.0380882
R48769 DVSS.n10532 DVSS.n10531 0.0380882
R48770 DVSS.n10533 DVSS.n10532 0.0380882
R48771 DVSS.n10533 DVSS.n1604 0.0380882
R48772 DVSS.n10543 DVSS.n1604 0.0380882
R48773 DVSS.n10544 DVSS.n10543 0.0380882
R48774 DVSS.n10545 DVSS.n10544 0.0380882
R48775 DVSS.n10545 DVSS.n1602 0.0380882
R48776 DVSS.n10555 DVSS.n1602 0.0380882
R48777 DVSS.n10556 DVSS.n10555 0.0380882
R48778 DVSS.n10557 DVSS.n10556 0.0380882
R48779 DVSS.n10557 DVSS.n1600 0.0380882
R48780 DVSS.n10567 DVSS.n1600 0.0380882
R48781 DVSS.n10568 DVSS.n10567 0.0380882
R48782 DVSS.n10569 DVSS.n10568 0.0380882
R48783 DVSS.n10569 DVSS.n1598 0.0380882
R48784 DVSS.n10579 DVSS.n1598 0.0380882
R48785 DVSS.n10580 DVSS.n10579 0.0380882
R48786 DVSS.n10581 DVSS.n10580 0.0380882
R48787 DVSS.n10581 DVSS.n1596 0.0380882
R48788 DVSS.n10591 DVSS.n1596 0.0380882
R48789 DVSS.n10592 DVSS.n10591 0.0380882
R48790 DVSS.n10593 DVSS.n10592 0.0380882
R48791 DVSS.n10593 DVSS.n1594 0.0380882
R48792 DVSS.n10603 DVSS.n1594 0.0380882
R48793 DVSS.n10604 DVSS.n10603 0.0380882
R48794 DVSS.n10605 DVSS.n10604 0.0380882
R48795 DVSS.n10605 DVSS.n1592 0.0380882
R48796 DVSS.n10615 DVSS.n1592 0.0380882
R48797 DVSS.n10616 DVSS.n10615 0.0380882
R48798 DVSS.n10617 DVSS.n10616 0.0380882
R48799 DVSS.n10617 DVSS.n1590 0.0380882
R48800 DVSS.n10627 DVSS.n1590 0.0380882
R48801 DVSS.n10628 DVSS.n10627 0.0380882
R48802 DVSS.n10629 DVSS.n10628 0.0380882
R48803 DVSS.n10629 DVSS.n1588 0.0380882
R48804 DVSS.n10639 DVSS.n1588 0.0380882
R48805 DVSS.n10640 DVSS.n10639 0.0380882
R48806 DVSS.n10641 DVSS.n10640 0.0380882
R48807 DVSS.n10641 DVSS.n1586 0.0380882
R48808 DVSS.n10651 DVSS.n1586 0.0380882
R48809 DVSS.n10652 DVSS.n10651 0.0380882
R48810 DVSS.n10653 DVSS.n10652 0.0380882
R48811 DVSS.n10653 DVSS.n1584 0.0380882
R48812 DVSS.n10663 DVSS.n1584 0.0380882
R48813 DVSS.n10664 DVSS.n10663 0.0380882
R48814 DVSS.n10665 DVSS.n10664 0.0380882
R48815 DVSS.n10665 DVSS.n1582 0.0380882
R48816 DVSS.n10675 DVSS.n1582 0.0380882
R48817 DVSS.n10676 DVSS.n10675 0.0380882
R48818 DVSS.n10677 DVSS.n10676 0.0380882
R48819 DVSS.n10677 DVSS.n1580 0.0380882
R48820 DVSS.n10687 DVSS.n1580 0.0380882
R48821 DVSS.n10688 DVSS.n10687 0.0380882
R48822 DVSS.n10689 DVSS.n10688 0.0380882
R48823 DVSS.n10689 DVSS.n1578 0.0380882
R48824 DVSS.n10699 DVSS.n1578 0.0380882
R48825 DVSS.n10700 DVSS.n10699 0.0380882
R48826 DVSS.n10701 DVSS.n10700 0.0380882
R48827 DVSS.n10701 DVSS.n1576 0.0380882
R48828 DVSS.n10711 DVSS.n1576 0.0380882
R48829 DVSS.n10712 DVSS.n10711 0.0380882
R48830 DVSS.n10713 DVSS.n10712 0.0380882
R48831 DVSS.n10713 DVSS.n1574 0.0380882
R48832 DVSS.n10723 DVSS.n1574 0.0380882
R48833 DVSS.n10724 DVSS.n10723 0.0380882
R48834 DVSS.n10725 DVSS.n10724 0.0380882
R48835 DVSS.n10725 DVSS.n1572 0.0380882
R48836 DVSS.n10735 DVSS.n1572 0.0380882
R48837 DVSS.n10736 DVSS.n10735 0.0380882
R48838 DVSS.n10737 DVSS.n10736 0.0380882
R48839 DVSS.n10737 DVSS.n1570 0.0380882
R48840 DVSS.n10747 DVSS.n1570 0.0380882
R48841 DVSS.n10748 DVSS.n10747 0.0380882
R48842 DVSS.n10749 DVSS.n10748 0.0380882
R48843 DVSS.n10749 DVSS.n1517 0.0380882
R48844 DVSS.n10506 DVSS.n1611 0.0380882
R48845 DVSS.n10510 DVSS.n1611 0.0380882
R48846 DVSS.n10514 DVSS.n10510 0.0380882
R48847 DVSS.n10518 DVSS.n10514 0.0380882
R48848 DVSS.n10518 DVSS.n1607 0.0380882
R48849 DVSS.n10522 DVSS.n1607 0.0380882
R48850 DVSS.n10526 DVSS.n10522 0.0380882
R48851 DVSS.n10530 DVSS.n10526 0.0380882
R48852 DVSS.n10530 DVSS.n1605 0.0380882
R48853 DVSS.n10534 DVSS.n1605 0.0380882
R48854 DVSS.n10538 DVSS.n10534 0.0380882
R48855 DVSS.n10542 DVSS.n10538 0.0380882
R48856 DVSS.n10542 DVSS.n1603 0.0380882
R48857 DVSS.n10546 DVSS.n1603 0.0380882
R48858 DVSS.n10550 DVSS.n10546 0.0380882
R48859 DVSS.n10554 DVSS.n10550 0.0380882
R48860 DVSS.n10554 DVSS.n1601 0.0380882
R48861 DVSS.n10558 DVSS.n1601 0.0380882
R48862 DVSS.n10562 DVSS.n10558 0.0380882
R48863 DVSS.n10566 DVSS.n10562 0.0380882
R48864 DVSS.n10566 DVSS.n1599 0.0380882
R48865 DVSS.n10570 DVSS.n1599 0.0380882
R48866 DVSS.n10574 DVSS.n10570 0.0380882
R48867 DVSS.n10578 DVSS.n10574 0.0380882
R48868 DVSS.n10578 DVSS.n1597 0.0380882
R48869 DVSS.n10582 DVSS.n1597 0.0380882
R48870 DVSS.n10586 DVSS.n10582 0.0380882
R48871 DVSS.n10590 DVSS.n10586 0.0380882
R48872 DVSS.n10590 DVSS.n1595 0.0380882
R48873 DVSS.n10594 DVSS.n1595 0.0380882
R48874 DVSS.n10598 DVSS.n10594 0.0380882
R48875 DVSS.n10602 DVSS.n10598 0.0380882
R48876 DVSS.n10602 DVSS.n1593 0.0380882
R48877 DVSS.n10606 DVSS.n1593 0.0380882
R48878 DVSS.n10610 DVSS.n10606 0.0380882
R48879 DVSS.n10614 DVSS.n10610 0.0380882
R48880 DVSS.n10614 DVSS.n1591 0.0380882
R48881 DVSS.n10618 DVSS.n1591 0.0380882
R48882 DVSS.n10622 DVSS.n10618 0.0380882
R48883 DVSS.n10626 DVSS.n10622 0.0380882
R48884 DVSS.n10626 DVSS.n1589 0.0380882
R48885 DVSS.n10630 DVSS.n1589 0.0380882
R48886 DVSS.n10634 DVSS.n10630 0.0380882
R48887 DVSS.n10638 DVSS.n10634 0.0380882
R48888 DVSS.n10638 DVSS.n1587 0.0380882
R48889 DVSS.n10642 DVSS.n1587 0.0380882
R48890 DVSS.n10646 DVSS.n10642 0.0380882
R48891 DVSS.n10650 DVSS.n10646 0.0380882
R48892 DVSS.n10650 DVSS.n1585 0.0380882
R48893 DVSS.n10654 DVSS.n1585 0.0380882
R48894 DVSS.n10658 DVSS.n10654 0.0380882
R48895 DVSS.n10662 DVSS.n10658 0.0380882
R48896 DVSS.n10662 DVSS.n1583 0.0380882
R48897 DVSS.n10666 DVSS.n1583 0.0380882
R48898 DVSS.n10670 DVSS.n10666 0.0380882
R48899 DVSS.n10674 DVSS.n10670 0.0380882
R48900 DVSS.n10674 DVSS.n1581 0.0380882
R48901 DVSS.n10678 DVSS.n1581 0.0380882
R48902 DVSS.n10682 DVSS.n10678 0.0380882
R48903 DVSS.n10686 DVSS.n10682 0.0380882
R48904 DVSS.n10686 DVSS.n1579 0.0380882
R48905 DVSS.n10690 DVSS.n1579 0.0380882
R48906 DVSS.n10694 DVSS.n10690 0.0380882
R48907 DVSS.n10698 DVSS.n10694 0.0380882
R48908 DVSS.n10698 DVSS.n1577 0.0380882
R48909 DVSS.n10702 DVSS.n1577 0.0380882
R48910 DVSS.n10706 DVSS.n10702 0.0380882
R48911 DVSS.n10710 DVSS.n10706 0.0380882
R48912 DVSS.n10710 DVSS.n1575 0.0380882
R48913 DVSS.n10714 DVSS.n1575 0.0380882
R48914 DVSS.n10718 DVSS.n10714 0.0380882
R48915 DVSS.n10722 DVSS.n10718 0.0380882
R48916 DVSS.n10722 DVSS.n1573 0.0380882
R48917 DVSS.n10726 DVSS.n1573 0.0380882
R48918 DVSS.n10730 DVSS.n10726 0.0380882
R48919 DVSS.n10734 DVSS.n10730 0.0380882
R48920 DVSS.n10734 DVSS.n1571 0.0380882
R48921 DVSS.n10738 DVSS.n1571 0.0380882
R48922 DVSS.n10742 DVSS.n10738 0.0380882
R48923 DVSS.n10746 DVSS.n10742 0.0380882
R48924 DVSS.n10746 DVSS.n1569 0.0380882
R48925 DVSS.n10750 DVSS.n1569 0.0380882
R48926 DVSS.n10750 DVSS.n1567 0.0380882
R48927 DVSS.n11104 DVSS.n10771 0.0380882
R48928 DVSS.n11096 DVSS.n10771 0.0380882
R48929 DVSS.n11096 DVSS.n11095 0.0380882
R48930 DVSS.n11095 DVSS.n11094 0.0380882
R48931 DVSS.n11094 DVSS.n10775 0.0380882
R48932 DVSS.n11086 DVSS.n10775 0.0380882
R48933 DVSS.n11086 DVSS.n11085 0.0380882
R48934 DVSS.n11085 DVSS.n11084 0.0380882
R48935 DVSS.n11084 DVSS.n10781 0.0380882
R48936 DVSS.n11076 DVSS.n10781 0.0380882
R48937 DVSS.n11076 DVSS.n11075 0.0380882
R48938 DVSS.n11075 DVSS.n11074 0.0380882
R48939 DVSS.n11074 DVSS.n10787 0.0380882
R48940 DVSS.n11066 DVSS.n10787 0.0380882
R48941 DVSS.n11066 DVSS.n11065 0.0380882
R48942 DVSS.n11065 DVSS.n11064 0.0380882
R48943 DVSS.n11064 DVSS.n10793 0.0380882
R48944 DVSS.n11056 DVSS.n10793 0.0380882
R48945 DVSS.n11056 DVSS.n11055 0.0380882
R48946 DVSS.n11055 DVSS.n11054 0.0380882
R48947 DVSS.n11054 DVSS.n10799 0.0380882
R48948 DVSS.n11046 DVSS.n10799 0.0380882
R48949 DVSS.n11046 DVSS.n11045 0.0380882
R48950 DVSS.n11045 DVSS.n11044 0.0380882
R48951 DVSS.n11044 DVSS.n10805 0.0380882
R48952 DVSS.n11036 DVSS.n10805 0.0380882
R48953 DVSS.n11036 DVSS.n11035 0.0380882
R48954 DVSS.n11035 DVSS.n11034 0.0380882
R48955 DVSS.n11034 DVSS.n10811 0.0380882
R48956 DVSS.n11026 DVSS.n10811 0.0380882
R48957 DVSS.n11026 DVSS.n11025 0.0380882
R48958 DVSS.n11025 DVSS.n11024 0.0380882
R48959 DVSS.n11024 DVSS.n10817 0.0380882
R48960 DVSS.n11016 DVSS.n10817 0.0380882
R48961 DVSS.n11016 DVSS.n11015 0.0380882
R48962 DVSS.n11015 DVSS.n11014 0.0380882
R48963 DVSS.n11014 DVSS.n10823 0.0380882
R48964 DVSS.n11006 DVSS.n10823 0.0380882
R48965 DVSS.n11006 DVSS.n11005 0.0380882
R48966 DVSS.n11005 DVSS.n11004 0.0380882
R48967 DVSS.n11004 DVSS.n10829 0.0380882
R48968 DVSS.n10996 DVSS.n10829 0.0380882
R48969 DVSS.n10996 DVSS.n10995 0.0380882
R48970 DVSS.n10995 DVSS.n10994 0.0380882
R48971 DVSS.n10994 DVSS.n10835 0.0380882
R48972 DVSS.n10986 DVSS.n10835 0.0380882
R48973 DVSS.n10986 DVSS.n10985 0.0380882
R48974 DVSS.n10985 DVSS.n10984 0.0380882
R48975 DVSS.n10984 DVSS.n10841 0.0380882
R48976 DVSS.n10976 DVSS.n10841 0.0380882
R48977 DVSS.n10976 DVSS.n10975 0.0380882
R48978 DVSS.n10975 DVSS.n10974 0.0380882
R48979 DVSS.n10974 DVSS.n10847 0.0380882
R48980 DVSS.n10966 DVSS.n10847 0.0380882
R48981 DVSS.n10966 DVSS.n10965 0.0380882
R48982 DVSS.n10965 DVSS.n10964 0.0380882
R48983 DVSS.n10964 DVSS.n10853 0.0380882
R48984 DVSS.n10956 DVSS.n10853 0.0380882
R48985 DVSS.n10956 DVSS.n10955 0.0380882
R48986 DVSS.n10955 DVSS.n10954 0.0380882
R48987 DVSS.n10954 DVSS.n10859 0.0380882
R48988 DVSS.n10946 DVSS.n10859 0.0380882
R48989 DVSS.n10946 DVSS.n10945 0.0380882
R48990 DVSS.n10945 DVSS.n10944 0.0380882
R48991 DVSS.n10944 DVSS.n10865 0.0380882
R48992 DVSS.n10936 DVSS.n10865 0.0380882
R48993 DVSS.n10936 DVSS.n10935 0.0380882
R48994 DVSS.n10935 DVSS.n10934 0.0380882
R48995 DVSS.n10934 DVSS.n10871 0.0380882
R48996 DVSS.n10926 DVSS.n10871 0.0380882
R48997 DVSS.n10926 DVSS.n10925 0.0380882
R48998 DVSS.n10925 DVSS.n10924 0.0380882
R48999 DVSS.n10924 DVSS.n10877 0.0380882
R49000 DVSS.n10916 DVSS.n10877 0.0380882
R49001 DVSS.n10916 DVSS.n10915 0.0380882
R49002 DVSS.n10915 DVSS.n10914 0.0380882
R49003 DVSS.n10914 DVSS.n10883 0.0380882
R49004 DVSS.n10906 DVSS.n10883 0.0380882
R49005 DVSS.n10906 DVSS.n10905 0.0380882
R49006 DVSS.n10905 DVSS.n10904 0.0380882
R49007 DVSS.n10904 DVSS.n10889 0.0380882
R49008 DVSS.n10896 DVSS.n10889 0.0380882
R49009 DVSS.n10896 DVSS.n10761 0.0380882
R49010 DVSS.n11103 DVSS.n10772 0.0380882
R49011 DVSS.n11097 DVSS.n10772 0.0380882
R49012 DVSS.n11097 DVSS.n10774 0.0380882
R49013 DVSS.n11093 DVSS.n10774 0.0380882
R49014 DVSS.n11093 DVSS.n10776 0.0380882
R49015 DVSS.n11087 DVSS.n10776 0.0380882
R49016 DVSS.n11087 DVSS.n10780 0.0380882
R49017 DVSS.n11083 DVSS.n10780 0.0380882
R49018 DVSS.n11083 DVSS.n10782 0.0380882
R49019 DVSS.n11077 DVSS.n10782 0.0380882
R49020 DVSS.n11077 DVSS.n10786 0.0380882
R49021 DVSS.n11073 DVSS.n10786 0.0380882
R49022 DVSS.n11073 DVSS.n10788 0.0380882
R49023 DVSS.n11067 DVSS.n10788 0.0380882
R49024 DVSS.n11067 DVSS.n10792 0.0380882
R49025 DVSS.n11063 DVSS.n10792 0.0380882
R49026 DVSS.n11063 DVSS.n10794 0.0380882
R49027 DVSS.n11057 DVSS.n10794 0.0380882
R49028 DVSS.n11057 DVSS.n10798 0.0380882
R49029 DVSS.n11053 DVSS.n10798 0.0380882
R49030 DVSS.n11053 DVSS.n10800 0.0380882
R49031 DVSS.n11047 DVSS.n10800 0.0380882
R49032 DVSS.n11047 DVSS.n10804 0.0380882
R49033 DVSS.n11043 DVSS.n10804 0.0380882
R49034 DVSS.n11043 DVSS.n10806 0.0380882
R49035 DVSS.n11037 DVSS.n10806 0.0380882
R49036 DVSS.n11037 DVSS.n10810 0.0380882
R49037 DVSS.n11033 DVSS.n10810 0.0380882
R49038 DVSS.n11033 DVSS.n10812 0.0380882
R49039 DVSS.n11027 DVSS.n10812 0.0380882
R49040 DVSS.n11027 DVSS.n10816 0.0380882
R49041 DVSS.n11023 DVSS.n10816 0.0380882
R49042 DVSS.n11023 DVSS.n10818 0.0380882
R49043 DVSS.n11017 DVSS.n10818 0.0380882
R49044 DVSS.n11017 DVSS.n10822 0.0380882
R49045 DVSS.n11013 DVSS.n10822 0.0380882
R49046 DVSS.n11013 DVSS.n10824 0.0380882
R49047 DVSS.n11007 DVSS.n10824 0.0380882
R49048 DVSS.n11007 DVSS.n10828 0.0380882
R49049 DVSS.n11003 DVSS.n10828 0.0380882
R49050 DVSS.n11003 DVSS.n10830 0.0380882
R49051 DVSS.n10997 DVSS.n10830 0.0380882
R49052 DVSS.n10997 DVSS.n10834 0.0380882
R49053 DVSS.n10993 DVSS.n10834 0.0380882
R49054 DVSS.n10993 DVSS.n10836 0.0380882
R49055 DVSS.n10987 DVSS.n10836 0.0380882
R49056 DVSS.n10987 DVSS.n10840 0.0380882
R49057 DVSS.n10983 DVSS.n10840 0.0380882
R49058 DVSS.n10983 DVSS.n10842 0.0380882
R49059 DVSS.n10977 DVSS.n10842 0.0380882
R49060 DVSS.n10977 DVSS.n10846 0.0380882
R49061 DVSS.n10973 DVSS.n10846 0.0380882
R49062 DVSS.n10973 DVSS.n10848 0.0380882
R49063 DVSS.n10967 DVSS.n10848 0.0380882
R49064 DVSS.n10967 DVSS.n10852 0.0380882
R49065 DVSS.n10963 DVSS.n10852 0.0380882
R49066 DVSS.n10963 DVSS.n10854 0.0380882
R49067 DVSS.n10957 DVSS.n10854 0.0380882
R49068 DVSS.n10957 DVSS.n10858 0.0380882
R49069 DVSS.n10953 DVSS.n10858 0.0380882
R49070 DVSS.n10953 DVSS.n10860 0.0380882
R49071 DVSS.n10947 DVSS.n10860 0.0380882
R49072 DVSS.n10947 DVSS.n10864 0.0380882
R49073 DVSS.n10943 DVSS.n10864 0.0380882
R49074 DVSS.n10943 DVSS.n10866 0.0380882
R49075 DVSS.n10937 DVSS.n10866 0.0380882
R49076 DVSS.n10937 DVSS.n10870 0.0380882
R49077 DVSS.n10933 DVSS.n10870 0.0380882
R49078 DVSS.n10933 DVSS.n10872 0.0380882
R49079 DVSS.n10927 DVSS.n10872 0.0380882
R49080 DVSS.n10927 DVSS.n10876 0.0380882
R49081 DVSS.n10923 DVSS.n10876 0.0380882
R49082 DVSS.n10923 DVSS.n10878 0.0380882
R49083 DVSS.n10917 DVSS.n10878 0.0380882
R49084 DVSS.n10917 DVSS.n10882 0.0380882
R49085 DVSS.n10913 DVSS.n10882 0.0380882
R49086 DVSS.n10913 DVSS.n10884 0.0380882
R49087 DVSS.n10907 DVSS.n10884 0.0380882
R49088 DVSS.n10907 DVSS.n10888 0.0380882
R49089 DVSS.n10903 DVSS.n10888 0.0380882
R49090 DVSS.n10903 DVSS.n10890 0.0380882
R49091 DVSS.n10897 DVSS.n10890 0.0380882
R49092 DVSS.n10897 DVSS.n10895 0.0380882
R49093 DVSS.n11264 DVSS.n11262 0.0380882
R49094 DVSS.n11265 DVSS.n11264 0.0380882
R49095 DVSS.n11266 DVSS.n11265 0.0380882
R49096 DVSS.n11266 DVSS.n11259 0.0380882
R49097 DVSS.n11273 DVSS.n11259 0.0380882
R49098 DVSS.n11274 DVSS.n11273 0.0380882
R49099 DVSS.n11275 DVSS.n11274 0.0380882
R49100 DVSS.n11275 DVSS.n11256 0.0380882
R49101 DVSS.n11282 DVSS.n11256 0.0380882
R49102 DVSS.n11283 DVSS.n11282 0.0380882
R49103 DVSS.n11284 DVSS.n11283 0.0380882
R49104 DVSS.n11284 DVSS.n11253 0.0380882
R49105 DVSS.n11291 DVSS.n11253 0.0380882
R49106 DVSS.n11292 DVSS.n11291 0.0380882
R49107 DVSS.n11293 DVSS.n11292 0.0380882
R49108 DVSS.n11293 DVSS.n11250 0.0380882
R49109 DVSS.n11300 DVSS.n11250 0.0380882
R49110 DVSS.n11301 DVSS.n11300 0.0380882
R49111 DVSS.n11302 DVSS.n11301 0.0380882
R49112 DVSS.n11302 DVSS.n11247 0.0380882
R49113 DVSS.n11309 DVSS.n11247 0.0380882
R49114 DVSS.n11310 DVSS.n11309 0.0380882
R49115 DVSS.n11311 DVSS.n11310 0.0380882
R49116 DVSS.n11311 DVSS.n11244 0.0380882
R49117 DVSS.n11318 DVSS.n11244 0.0380882
R49118 DVSS.n11319 DVSS.n11318 0.0380882
R49119 DVSS.n11320 DVSS.n11319 0.0380882
R49120 DVSS.n11320 DVSS.n11241 0.0380882
R49121 DVSS.n11327 DVSS.n11241 0.0380882
R49122 DVSS.n11328 DVSS.n11327 0.0380882
R49123 DVSS.n11329 DVSS.n11328 0.0380882
R49124 DVSS.n11329 DVSS.n11238 0.0380882
R49125 DVSS.n11336 DVSS.n11238 0.0380882
R49126 DVSS.n11337 DVSS.n11336 0.0380882
R49127 DVSS.n11338 DVSS.n11337 0.0380882
R49128 DVSS.n11338 DVSS.n11235 0.0380882
R49129 DVSS.n11345 DVSS.n11235 0.0380882
R49130 DVSS.n11346 DVSS.n11345 0.0380882
R49131 DVSS.n11347 DVSS.n11346 0.0380882
R49132 DVSS.n11347 DVSS.n11232 0.0380882
R49133 DVSS.n11354 DVSS.n11232 0.0380882
R49134 DVSS.n11355 DVSS.n11354 0.0380882
R49135 DVSS.n11356 DVSS.n11355 0.0380882
R49136 DVSS.n11356 DVSS.n11229 0.0380882
R49137 DVSS.n11363 DVSS.n11229 0.0380882
R49138 DVSS.n11364 DVSS.n11363 0.0380882
R49139 DVSS.n11365 DVSS.n11364 0.0380882
R49140 DVSS.n11365 DVSS.n11226 0.0380882
R49141 DVSS.n11372 DVSS.n11226 0.0380882
R49142 DVSS.n11373 DVSS.n11372 0.0380882
R49143 DVSS.n11374 DVSS.n11373 0.0380882
R49144 DVSS.n11374 DVSS.n11223 0.0380882
R49145 DVSS.n11381 DVSS.n11223 0.0380882
R49146 DVSS.n11382 DVSS.n11381 0.0380882
R49147 DVSS.n11383 DVSS.n11382 0.0380882
R49148 DVSS.n11383 DVSS.n11220 0.0380882
R49149 DVSS.n11390 DVSS.n11220 0.0380882
R49150 DVSS.n11391 DVSS.n11390 0.0380882
R49151 DVSS.n11392 DVSS.n11391 0.0380882
R49152 DVSS.n11392 DVSS.n11217 0.0380882
R49153 DVSS.n11399 DVSS.n11217 0.0380882
R49154 DVSS.n11400 DVSS.n11399 0.0380882
R49155 DVSS.n11401 DVSS.n11400 0.0380882
R49156 DVSS.n11401 DVSS.n11214 0.0380882
R49157 DVSS.n11408 DVSS.n11214 0.0380882
R49158 DVSS.n11409 DVSS.n11408 0.0380882
R49159 DVSS.n11410 DVSS.n11409 0.0380882
R49160 DVSS.n11410 DVSS.n11211 0.0380882
R49161 DVSS.n11417 DVSS.n11211 0.0380882
R49162 DVSS.n11418 DVSS.n11417 0.0380882
R49163 DVSS.n11419 DVSS.n11418 0.0380882
R49164 DVSS.n11419 DVSS.n11208 0.0380882
R49165 DVSS.n11426 DVSS.n11208 0.0380882
R49166 DVSS.n11427 DVSS.n11426 0.0380882
R49167 DVSS.n11428 DVSS.n11427 0.0380882
R49168 DVSS.n11428 DVSS.n11205 0.0380882
R49169 DVSS.n11435 DVSS.n11205 0.0380882
R49170 DVSS.n11436 DVSS.n11435 0.0380882
R49171 DVSS.n11437 DVSS.n11436 0.0380882
R49172 DVSS.n11437 DVSS.n11202 0.0380882
R49173 DVSS.n11444 DVSS.n11202 0.0380882
R49174 DVSS.n11445 DVSS.n11444 0.0380882
R49175 DVSS.n11446 DVSS.n11445 0.0380882
R49176 DVSS.n11263 DVSS.n11155 0.0380882
R49177 DVSS.n11263 DVSS.n11261 0.0380882
R49178 DVSS.n11268 DVSS.n11261 0.0380882
R49179 DVSS.n11270 DVSS.n11268 0.0380882
R49180 DVSS.n11272 DVSS.n11270 0.0380882
R49181 DVSS.n11272 DVSS.n11258 0.0380882
R49182 DVSS.n11277 DVSS.n11258 0.0380882
R49183 DVSS.n11279 DVSS.n11277 0.0380882
R49184 DVSS.n11281 DVSS.n11279 0.0380882
R49185 DVSS.n11281 DVSS.n11255 0.0380882
R49186 DVSS.n11286 DVSS.n11255 0.0380882
R49187 DVSS.n11288 DVSS.n11286 0.0380882
R49188 DVSS.n11290 DVSS.n11288 0.0380882
R49189 DVSS.n11290 DVSS.n11252 0.0380882
R49190 DVSS.n11295 DVSS.n11252 0.0380882
R49191 DVSS.n11297 DVSS.n11295 0.0380882
R49192 DVSS.n11299 DVSS.n11297 0.0380882
R49193 DVSS.n11299 DVSS.n11249 0.0380882
R49194 DVSS.n11304 DVSS.n11249 0.0380882
R49195 DVSS.n11306 DVSS.n11304 0.0380882
R49196 DVSS.n11308 DVSS.n11306 0.0380882
R49197 DVSS.n11308 DVSS.n11246 0.0380882
R49198 DVSS.n11313 DVSS.n11246 0.0380882
R49199 DVSS.n11315 DVSS.n11313 0.0380882
R49200 DVSS.n11317 DVSS.n11315 0.0380882
R49201 DVSS.n11317 DVSS.n11243 0.0380882
R49202 DVSS.n11322 DVSS.n11243 0.0380882
R49203 DVSS.n11324 DVSS.n11322 0.0380882
R49204 DVSS.n11326 DVSS.n11324 0.0380882
R49205 DVSS.n11326 DVSS.n11240 0.0380882
R49206 DVSS.n11331 DVSS.n11240 0.0380882
R49207 DVSS.n11333 DVSS.n11331 0.0380882
R49208 DVSS.n11335 DVSS.n11333 0.0380882
R49209 DVSS.n11335 DVSS.n11237 0.0380882
R49210 DVSS.n11340 DVSS.n11237 0.0380882
R49211 DVSS.n11342 DVSS.n11340 0.0380882
R49212 DVSS.n11344 DVSS.n11342 0.0380882
R49213 DVSS.n11344 DVSS.n11234 0.0380882
R49214 DVSS.n11349 DVSS.n11234 0.0380882
R49215 DVSS.n11351 DVSS.n11349 0.0380882
R49216 DVSS.n11353 DVSS.n11351 0.0380882
R49217 DVSS.n11353 DVSS.n11231 0.0380882
R49218 DVSS.n11358 DVSS.n11231 0.0380882
R49219 DVSS.n11360 DVSS.n11358 0.0380882
R49220 DVSS.n11362 DVSS.n11360 0.0380882
R49221 DVSS.n11362 DVSS.n11228 0.0380882
R49222 DVSS.n11367 DVSS.n11228 0.0380882
R49223 DVSS.n11369 DVSS.n11367 0.0380882
R49224 DVSS.n11371 DVSS.n11369 0.0380882
R49225 DVSS.n11371 DVSS.n11225 0.0380882
R49226 DVSS.n11376 DVSS.n11225 0.0380882
R49227 DVSS.n11378 DVSS.n11376 0.0380882
R49228 DVSS.n11380 DVSS.n11378 0.0380882
R49229 DVSS.n11380 DVSS.n11222 0.0380882
R49230 DVSS.n11385 DVSS.n11222 0.0380882
R49231 DVSS.n11387 DVSS.n11385 0.0380882
R49232 DVSS.n11389 DVSS.n11387 0.0380882
R49233 DVSS.n11389 DVSS.n11219 0.0380882
R49234 DVSS.n11394 DVSS.n11219 0.0380882
R49235 DVSS.n11396 DVSS.n11394 0.0380882
R49236 DVSS.n11398 DVSS.n11396 0.0380882
R49237 DVSS.n11398 DVSS.n11216 0.0380882
R49238 DVSS.n11403 DVSS.n11216 0.0380882
R49239 DVSS.n11405 DVSS.n11403 0.0380882
R49240 DVSS.n11407 DVSS.n11405 0.0380882
R49241 DVSS.n11407 DVSS.n11213 0.0380882
R49242 DVSS.n11412 DVSS.n11213 0.0380882
R49243 DVSS.n11414 DVSS.n11412 0.0380882
R49244 DVSS.n11416 DVSS.n11414 0.0380882
R49245 DVSS.n11416 DVSS.n11210 0.0380882
R49246 DVSS.n11421 DVSS.n11210 0.0380882
R49247 DVSS.n11423 DVSS.n11421 0.0380882
R49248 DVSS.n11425 DVSS.n11423 0.0380882
R49249 DVSS.n11425 DVSS.n11207 0.0380882
R49250 DVSS.n11430 DVSS.n11207 0.0380882
R49251 DVSS.n11432 DVSS.n11430 0.0380882
R49252 DVSS.n11434 DVSS.n11432 0.0380882
R49253 DVSS.n11434 DVSS.n11204 0.0380882
R49254 DVSS.n11439 DVSS.n11204 0.0380882
R49255 DVSS.n11441 DVSS.n11439 0.0380882
R49256 DVSS.n11443 DVSS.n11441 0.0380882
R49257 DVSS.n11443 DVSS.n11201 0.0380882
R49258 DVSS.n13335 DVSS.n11201 0.0380882
R49259 DVSS.n13138 DVSS.n13136 0.0380882
R49260 DVSS.n13139 DVSS.n13138 0.0380882
R49261 DVSS.n13140 DVSS.n13139 0.0380882
R49262 DVSS.n13140 DVSS.n11606 0.0380882
R49263 DVSS.n13147 DVSS.n11606 0.0380882
R49264 DVSS.n13148 DVSS.n13147 0.0380882
R49265 DVSS.n13149 DVSS.n13148 0.0380882
R49266 DVSS.n13149 DVSS.n11603 0.0380882
R49267 DVSS.n13156 DVSS.n11603 0.0380882
R49268 DVSS.n13157 DVSS.n13156 0.0380882
R49269 DVSS.n13158 DVSS.n13157 0.0380882
R49270 DVSS.n13158 DVSS.n11600 0.0380882
R49271 DVSS.n13165 DVSS.n11600 0.0380882
R49272 DVSS.n13166 DVSS.n13165 0.0380882
R49273 DVSS.n13167 DVSS.n13166 0.0380882
R49274 DVSS.n13167 DVSS.n11597 0.0380882
R49275 DVSS.n13174 DVSS.n11597 0.0380882
R49276 DVSS.n13175 DVSS.n13174 0.0380882
R49277 DVSS.n13176 DVSS.n13175 0.0380882
R49278 DVSS.n13176 DVSS.n11594 0.0380882
R49279 DVSS.n13183 DVSS.n11594 0.0380882
R49280 DVSS.n13184 DVSS.n13183 0.0380882
R49281 DVSS.n13185 DVSS.n13184 0.0380882
R49282 DVSS.n13185 DVSS.n11591 0.0380882
R49283 DVSS.n13192 DVSS.n11591 0.0380882
R49284 DVSS.n13193 DVSS.n13192 0.0380882
R49285 DVSS.n13194 DVSS.n13193 0.0380882
R49286 DVSS.n13194 DVSS.n11588 0.0380882
R49287 DVSS.n13201 DVSS.n11588 0.0380882
R49288 DVSS.n13202 DVSS.n13201 0.0380882
R49289 DVSS.n13203 DVSS.n13202 0.0380882
R49290 DVSS.n13203 DVSS.n11585 0.0380882
R49291 DVSS.n13210 DVSS.n11585 0.0380882
R49292 DVSS.n13211 DVSS.n13210 0.0380882
R49293 DVSS.n13212 DVSS.n13211 0.0380882
R49294 DVSS.n13212 DVSS.n11582 0.0380882
R49295 DVSS.n13219 DVSS.n11582 0.0380882
R49296 DVSS.n13220 DVSS.n13219 0.0380882
R49297 DVSS.n13221 DVSS.n13220 0.0380882
R49298 DVSS.n13221 DVSS.n11579 0.0380882
R49299 DVSS.n13228 DVSS.n11579 0.0380882
R49300 DVSS.n13229 DVSS.n13228 0.0380882
R49301 DVSS.n13230 DVSS.n13229 0.0380882
R49302 DVSS.n13230 DVSS.n11576 0.0380882
R49303 DVSS.n13237 DVSS.n11576 0.0380882
R49304 DVSS.n13238 DVSS.n13237 0.0380882
R49305 DVSS.n13239 DVSS.n13238 0.0380882
R49306 DVSS.n13239 DVSS.n11573 0.0380882
R49307 DVSS.n13246 DVSS.n11573 0.0380882
R49308 DVSS.n13247 DVSS.n13246 0.0380882
R49309 DVSS.n13248 DVSS.n13247 0.0380882
R49310 DVSS.n13248 DVSS.n11570 0.0380882
R49311 DVSS.n13255 DVSS.n11570 0.0380882
R49312 DVSS.n13256 DVSS.n13255 0.0380882
R49313 DVSS.n13257 DVSS.n13256 0.0380882
R49314 DVSS.n13257 DVSS.n11567 0.0380882
R49315 DVSS.n13264 DVSS.n11567 0.0380882
R49316 DVSS.n13265 DVSS.n13264 0.0380882
R49317 DVSS.n13266 DVSS.n13265 0.0380882
R49318 DVSS.n13266 DVSS.n11564 0.0380882
R49319 DVSS.n13273 DVSS.n11564 0.0380882
R49320 DVSS.n13274 DVSS.n13273 0.0380882
R49321 DVSS.n13275 DVSS.n13274 0.0380882
R49322 DVSS.n13275 DVSS.n11561 0.0380882
R49323 DVSS.n13282 DVSS.n11561 0.0380882
R49324 DVSS.n13283 DVSS.n13282 0.0380882
R49325 DVSS.n13284 DVSS.n13283 0.0380882
R49326 DVSS.n13284 DVSS.n11558 0.0380882
R49327 DVSS.n13291 DVSS.n11558 0.0380882
R49328 DVSS.n13292 DVSS.n13291 0.0380882
R49329 DVSS.n13293 DVSS.n13292 0.0380882
R49330 DVSS.n13293 DVSS.n11555 0.0380882
R49331 DVSS.n13300 DVSS.n11555 0.0380882
R49332 DVSS.n13301 DVSS.n13300 0.0380882
R49333 DVSS.n13302 DVSS.n13301 0.0380882
R49334 DVSS.n13302 DVSS.n11552 0.0380882
R49335 DVSS.n13309 DVSS.n11552 0.0380882
R49336 DVSS.n13310 DVSS.n13309 0.0380882
R49337 DVSS.n13311 DVSS.n13310 0.0380882
R49338 DVSS.n13311 DVSS.n11549 0.0380882
R49339 DVSS.n13318 DVSS.n11549 0.0380882
R49340 DVSS.n13319 DVSS.n13318 0.0380882
R49341 DVSS.n13320 DVSS.n13319 0.0380882
R49342 DVSS.n13137 DVSS.n11503 0.0380882
R49343 DVSS.n13137 DVSS.n11608 0.0380882
R49344 DVSS.n13142 DVSS.n11608 0.0380882
R49345 DVSS.n13144 DVSS.n13142 0.0380882
R49346 DVSS.n13146 DVSS.n13144 0.0380882
R49347 DVSS.n13146 DVSS.n11605 0.0380882
R49348 DVSS.n13151 DVSS.n11605 0.0380882
R49349 DVSS.n13153 DVSS.n13151 0.0380882
R49350 DVSS.n13155 DVSS.n13153 0.0380882
R49351 DVSS.n13155 DVSS.n11602 0.0380882
R49352 DVSS.n13160 DVSS.n11602 0.0380882
R49353 DVSS.n13162 DVSS.n13160 0.0380882
R49354 DVSS.n13164 DVSS.n13162 0.0380882
R49355 DVSS.n13164 DVSS.n11599 0.0380882
R49356 DVSS.n13169 DVSS.n11599 0.0380882
R49357 DVSS.n13171 DVSS.n13169 0.0380882
R49358 DVSS.n13173 DVSS.n13171 0.0380882
R49359 DVSS.n13173 DVSS.n11596 0.0380882
R49360 DVSS.n13178 DVSS.n11596 0.0380882
R49361 DVSS.n13180 DVSS.n13178 0.0380882
R49362 DVSS.n13182 DVSS.n13180 0.0380882
R49363 DVSS.n13182 DVSS.n11593 0.0380882
R49364 DVSS.n13187 DVSS.n11593 0.0380882
R49365 DVSS.n13189 DVSS.n13187 0.0380882
R49366 DVSS.n13191 DVSS.n13189 0.0380882
R49367 DVSS.n13191 DVSS.n11590 0.0380882
R49368 DVSS.n13196 DVSS.n11590 0.0380882
R49369 DVSS.n13198 DVSS.n13196 0.0380882
R49370 DVSS.n13200 DVSS.n13198 0.0380882
R49371 DVSS.n13200 DVSS.n11587 0.0380882
R49372 DVSS.n13205 DVSS.n11587 0.0380882
R49373 DVSS.n13207 DVSS.n13205 0.0380882
R49374 DVSS.n13209 DVSS.n13207 0.0380882
R49375 DVSS.n13209 DVSS.n11584 0.0380882
R49376 DVSS.n13214 DVSS.n11584 0.0380882
R49377 DVSS.n13216 DVSS.n13214 0.0380882
R49378 DVSS.n13218 DVSS.n13216 0.0380882
R49379 DVSS.n13218 DVSS.n11581 0.0380882
R49380 DVSS.n13223 DVSS.n11581 0.0380882
R49381 DVSS.n13225 DVSS.n13223 0.0380882
R49382 DVSS.n13227 DVSS.n13225 0.0380882
R49383 DVSS.n13227 DVSS.n11578 0.0380882
R49384 DVSS.n13232 DVSS.n11578 0.0380882
R49385 DVSS.n13234 DVSS.n13232 0.0380882
R49386 DVSS.n13236 DVSS.n13234 0.0380882
R49387 DVSS.n13236 DVSS.n11575 0.0380882
R49388 DVSS.n13241 DVSS.n11575 0.0380882
R49389 DVSS.n13243 DVSS.n13241 0.0380882
R49390 DVSS.n13245 DVSS.n13243 0.0380882
R49391 DVSS.n13245 DVSS.n11572 0.0380882
R49392 DVSS.n13250 DVSS.n11572 0.0380882
R49393 DVSS.n13252 DVSS.n13250 0.0380882
R49394 DVSS.n13254 DVSS.n13252 0.0380882
R49395 DVSS.n13254 DVSS.n11569 0.0380882
R49396 DVSS.n13259 DVSS.n11569 0.0380882
R49397 DVSS.n13261 DVSS.n13259 0.0380882
R49398 DVSS.n13263 DVSS.n13261 0.0380882
R49399 DVSS.n13263 DVSS.n11566 0.0380882
R49400 DVSS.n13268 DVSS.n11566 0.0380882
R49401 DVSS.n13270 DVSS.n13268 0.0380882
R49402 DVSS.n13272 DVSS.n13270 0.0380882
R49403 DVSS.n13272 DVSS.n11563 0.0380882
R49404 DVSS.n13277 DVSS.n11563 0.0380882
R49405 DVSS.n13279 DVSS.n13277 0.0380882
R49406 DVSS.n13281 DVSS.n13279 0.0380882
R49407 DVSS.n13281 DVSS.n11560 0.0380882
R49408 DVSS.n13286 DVSS.n11560 0.0380882
R49409 DVSS.n13288 DVSS.n13286 0.0380882
R49410 DVSS.n13290 DVSS.n13288 0.0380882
R49411 DVSS.n13290 DVSS.n11557 0.0380882
R49412 DVSS.n13295 DVSS.n11557 0.0380882
R49413 DVSS.n13297 DVSS.n13295 0.0380882
R49414 DVSS.n13299 DVSS.n13297 0.0380882
R49415 DVSS.n13299 DVSS.n11554 0.0380882
R49416 DVSS.n13304 DVSS.n11554 0.0380882
R49417 DVSS.n13306 DVSS.n13304 0.0380882
R49418 DVSS.n13308 DVSS.n13306 0.0380882
R49419 DVSS.n13308 DVSS.n11551 0.0380882
R49420 DVSS.n13313 DVSS.n11551 0.0380882
R49421 DVSS.n13315 DVSS.n13313 0.0380882
R49422 DVSS.n13317 DVSS.n13315 0.0380882
R49423 DVSS.n13317 DVSS.n11548 0.0380882
R49424 DVSS.n13321 DVSS.n11548 0.0380882
R49425 DVSS.n6779 DVSS.n5872 0.0380882
R49426 DVSS.n6779 DVSS.n6774 0.0380882
R49427 DVSS.n6789 DVSS.n6774 0.0380882
R49428 DVSS.n6790 DVSS.n6789 0.0380882
R49429 DVSS.n6791 DVSS.n6790 0.0380882
R49430 DVSS.n6791 DVSS.n6770 0.0380882
R49431 DVSS.n6801 DVSS.n6770 0.0380882
R49432 DVSS.n6802 DVSS.n6801 0.0380882
R49433 DVSS.n6803 DVSS.n6802 0.0380882
R49434 DVSS.n6803 DVSS.n6766 0.0380882
R49435 DVSS.n6813 DVSS.n6766 0.0380882
R49436 DVSS.n6814 DVSS.n6813 0.0380882
R49437 DVSS.n6815 DVSS.n6814 0.0380882
R49438 DVSS.n6815 DVSS.n6762 0.0380882
R49439 DVSS.n6825 DVSS.n6762 0.0380882
R49440 DVSS.n6826 DVSS.n6825 0.0380882
R49441 DVSS.n6827 DVSS.n6826 0.0380882
R49442 DVSS.n6827 DVSS.n6758 0.0380882
R49443 DVSS.n6837 DVSS.n6758 0.0380882
R49444 DVSS.n6838 DVSS.n6837 0.0380882
R49445 DVSS.n6839 DVSS.n6838 0.0380882
R49446 DVSS.n6839 DVSS.n6754 0.0380882
R49447 DVSS.n6849 DVSS.n6754 0.0380882
R49448 DVSS.n6850 DVSS.n6849 0.0380882
R49449 DVSS.n6851 DVSS.n6850 0.0380882
R49450 DVSS.n6851 DVSS.n6750 0.0380882
R49451 DVSS.n6861 DVSS.n6750 0.0380882
R49452 DVSS.n6862 DVSS.n6861 0.0380882
R49453 DVSS.n6863 DVSS.n6862 0.0380882
R49454 DVSS.n6863 DVSS.n6746 0.0380882
R49455 DVSS.n6873 DVSS.n6746 0.0380882
R49456 DVSS.n6874 DVSS.n6873 0.0380882
R49457 DVSS.n6875 DVSS.n6874 0.0380882
R49458 DVSS.n6875 DVSS.n6742 0.0380882
R49459 DVSS.n6885 DVSS.n6742 0.0380882
R49460 DVSS.n6886 DVSS.n6885 0.0380882
R49461 DVSS.n6887 DVSS.n6886 0.0380882
R49462 DVSS.n6887 DVSS.n6738 0.0380882
R49463 DVSS.n6897 DVSS.n6738 0.0380882
R49464 DVSS.n6898 DVSS.n6897 0.0380882
R49465 DVSS.n6899 DVSS.n6898 0.0380882
R49466 DVSS.n6899 DVSS.n6734 0.0380882
R49467 DVSS.n6909 DVSS.n6734 0.0380882
R49468 DVSS.n6910 DVSS.n6909 0.0380882
R49469 DVSS.n6911 DVSS.n6910 0.0380882
R49470 DVSS.n6911 DVSS.n6730 0.0380882
R49471 DVSS.n6921 DVSS.n6730 0.0380882
R49472 DVSS.n6922 DVSS.n6921 0.0380882
R49473 DVSS.n6923 DVSS.n6922 0.0380882
R49474 DVSS.n6923 DVSS.n6726 0.0380882
R49475 DVSS.n6933 DVSS.n6726 0.0380882
R49476 DVSS.n6934 DVSS.n6933 0.0380882
R49477 DVSS.n6935 DVSS.n6934 0.0380882
R49478 DVSS.n6935 DVSS.n6722 0.0380882
R49479 DVSS.n6945 DVSS.n6722 0.0380882
R49480 DVSS.n6946 DVSS.n6945 0.0380882
R49481 DVSS.n6947 DVSS.n6946 0.0380882
R49482 DVSS.n6947 DVSS.n6718 0.0380882
R49483 DVSS.n6957 DVSS.n6718 0.0380882
R49484 DVSS.n6958 DVSS.n6957 0.0380882
R49485 DVSS.n6959 DVSS.n6958 0.0380882
R49486 DVSS.n6959 DVSS.n6714 0.0380882
R49487 DVSS.n6969 DVSS.n6714 0.0380882
R49488 DVSS.n6970 DVSS.n6969 0.0380882
R49489 DVSS.n6971 DVSS.n6970 0.0380882
R49490 DVSS.n6971 DVSS.n6710 0.0380882
R49491 DVSS.n6981 DVSS.n6710 0.0380882
R49492 DVSS.n6982 DVSS.n6981 0.0380882
R49493 DVSS.n6983 DVSS.n6982 0.0380882
R49494 DVSS.n6983 DVSS.n6706 0.0380882
R49495 DVSS.n6993 DVSS.n6706 0.0380882
R49496 DVSS.n6994 DVSS.n6993 0.0380882
R49497 DVSS.n6995 DVSS.n6994 0.0380882
R49498 DVSS.n6995 DVSS.n6702 0.0380882
R49499 DVSS.n7005 DVSS.n6702 0.0380882
R49500 DVSS.n7006 DVSS.n7005 0.0380882
R49501 DVSS.n7007 DVSS.n7006 0.0380882
R49502 DVSS.n7007 DVSS.n6698 0.0380882
R49503 DVSS.n7017 DVSS.n6698 0.0380882
R49504 DVSS.n7018 DVSS.n7017 0.0380882
R49505 DVSS.n7019 DVSS.n7018 0.0380882
R49506 DVSS.n7019 DVSS.n6694 0.0380882
R49507 DVSS.n7027 DVSS.n6694 0.0380882
R49508 DVSS.n6780 DVSS.n6778 0.0380882
R49509 DVSS.n6780 DVSS.n6775 0.0380882
R49510 DVSS.n6788 DVSS.n6775 0.0380882
R49511 DVSS.n6788 DVSS.n6773 0.0380882
R49512 DVSS.n6792 DVSS.n6773 0.0380882
R49513 DVSS.n6792 DVSS.n6771 0.0380882
R49514 DVSS.n6800 DVSS.n6771 0.0380882
R49515 DVSS.n6800 DVSS.n6769 0.0380882
R49516 DVSS.n6804 DVSS.n6769 0.0380882
R49517 DVSS.n6804 DVSS.n6767 0.0380882
R49518 DVSS.n6812 DVSS.n6767 0.0380882
R49519 DVSS.n6812 DVSS.n6765 0.0380882
R49520 DVSS.n6816 DVSS.n6765 0.0380882
R49521 DVSS.n6816 DVSS.n6763 0.0380882
R49522 DVSS.n6824 DVSS.n6763 0.0380882
R49523 DVSS.n6824 DVSS.n6761 0.0380882
R49524 DVSS.n6828 DVSS.n6761 0.0380882
R49525 DVSS.n6828 DVSS.n6759 0.0380882
R49526 DVSS.n6836 DVSS.n6759 0.0380882
R49527 DVSS.n6836 DVSS.n6757 0.0380882
R49528 DVSS.n6840 DVSS.n6757 0.0380882
R49529 DVSS.n6840 DVSS.n6755 0.0380882
R49530 DVSS.n6848 DVSS.n6755 0.0380882
R49531 DVSS.n6848 DVSS.n6753 0.0380882
R49532 DVSS.n6852 DVSS.n6753 0.0380882
R49533 DVSS.n6852 DVSS.n6751 0.0380882
R49534 DVSS.n6860 DVSS.n6751 0.0380882
R49535 DVSS.n6860 DVSS.n6749 0.0380882
R49536 DVSS.n6864 DVSS.n6749 0.0380882
R49537 DVSS.n6864 DVSS.n6747 0.0380882
R49538 DVSS.n6872 DVSS.n6747 0.0380882
R49539 DVSS.n6872 DVSS.n6745 0.0380882
R49540 DVSS.n6876 DVSS.n6745 0.0380882
R49541 DVSS.n6876 DVSS.n6743 0.0380882
R49542 DVSS.n6884 DVSS.n6743 0.0380882
R49543 DVSS.n6884 DVSS.n6741 0.0380882
R49544 DVSS.n6888 DVSS.n6741 0.0380882
R49545 DVSS.n6888 DVSS.n6739 0.0380882
R49546 DVSS.n6896 DVSS.n6739 0.0380882
R49547 DVSS.n6896 DVSS.n6737 0.0380882
R49548 DVSS.n6900 DVSS.n6737 0.0380882
R49549 DVSS.n6900 DVSS.n6735 0.0380882
R49550 DVSS.n6908 DVSS.n6735 0.0380882
R49551 DVSS.n6908 DVSS.n6733 0.0380882
R49552 DVSS.n6912 DVSS.n6733 0.0380882
R49553 DVSS.n6912 DVSS.n6731 0.0380882
R49554 DVSS.n6920 DVSS.n6731 0.0380882
R49555 DVSS.n6920 DVSS.n6729 0.0380882
R49556 DVSS.n6924 DVSS.n6729 0.0380882
R49557 DVSS.n6924 DVSS.n6727 0.0380882
R49558 DVSS.n6932 DVSS.n6727 0.0380882
R49559 DVSS.n6932 DVSS.n6725 0.0380882
R49560 DVSS.n6936 DVSS.n6725 0.0380882
R49561 DVSS.n6936 DVSS.n6723 0.0380882
R49562 DVSS.n6944 DVSS.n6723 0.0380882
R49563 DVSS.n6944 DVSS.n6721 0.0380882
R49564 DVSS.n6948 DVSS.n6721 0.0380882
R49565 DVSS.n6948 DVSS.n6719 0.0380882
R49566 DVSS.n6956 DVSS.n6719 0.0380882
R49567 DVSS.n6956 DVSS.n6717 0.0380882
R49568 DVSS.n6960 DVSS.n6717 0.0380882
R49569 DVSS.n6960 DVSS.n6715 0.0380882
R49570 DVSS.n6968 DVSS.n6715 0.0380882
R49571 DVSS.n6968 DVSS.n6713 0.0380882
R49572 DVSS.n6972 DVSS.n6713 0.0380882
R49573 DVSS.n6972 DVSS.n6711 0.0380882
R49574 DVSS.n6980 DVSS.n6711 0.0380882
R49575 DVSS.n6980 DVSS.n6709 0.0380882
R49576 DVSS.n6984 DVSS.n6709 0.0380882
R49577 DVSS.n6984 DVSS.n6707 0.0380882
R49578 DVSS.n6992 DVSS.n6707 0.0380882
R49579 DVSS.n6992 DVSS.n6705 0.0380882
R49580 DVSS.n6996 DVSS.n6705 0.0380882
R49581 DVSS.n6996 DVSS.n6703 0.0380882
R49582 DVSS.n7004 DVSS.n6703 0.0380882
R49583 DVSS.n7004 DVSS.n6701 0.0380882
R49584 DVSS.n7008 DVSS.n6701 0.0380882
R49585 DVSS.n7008 DVSS.n6699 0.0380882
R49586 DVSS.n7016 DVSS.n6699 0.0380882
R49587 DVSS.n7016 DVSS.n6697 0.0380882
R49588 DVSS.n7020 DVSS.n6697 0.0380882
R49589 DVSS.n7020 DVSS.n6695 0.0380882
R49590 DVSS.n7026 DVSS.n6695 0.0380882
R49591 DVSS.n6227 DVSS.n5893 0.0380882
R49592 DVSS.n6227 DVSS.n6226 0.0380882
R49593 DVSS.n6226 DVSS.n6225 0.0380882
R49594 DVSS.n6225 DVSS.n5943 0.0380882
R49595 DVSS.n6215 DVSS.n5943 0.0380882
R49596 DVSS.n6215 DVSS.n6214 0.0380882
R49597 DVSS.n6214 DVSS.n6213 0.0380882
R49598 DVSS.n6213 DVSS.n5945 0.0380882
R49599 DVSS.n6203 DVSS.n5945 0.0380882
R49600 DVSS.n6203 DVSS.n6202 0.0380882
R49601 DVSS.n6202 DVSS.n6201 0.0380882
R49602 DVSS.n6201 DVSS.n5947 0.0380882
R49603 DVSS.n6191 DVSS.n5947 0.0380882
R49604 DVSS.n6191 DVSS.n6190 0.0380882
R49605 DVSS.n6190 DVSS.n6189 0.0380882
R49606 DVSS.n6189 DVSS.n5949 0.0380882
R49607 DVSS.n6179 DVSS.n5949 0.0380882
R49608 DVSS.n6179 DVSS.n6178 0.0380882
R49609 DVSS.n6178 DVSS.n6177 0.0380882
R49610 DVSS.n6177 DVSS.n5951 0.0380882
R49611 DVSS.n6167 DVSS.n5951 0.0380882
R49612 DVSS.n6167 DVSS.n6166 0.0380882
R49613 DVSS.n6166 DVSS.n6165 0.0380882
R49614 DVSS.n6165 DVSS.n5953 0.0380882
R49615 DVSS.n6155 DVSS.n5953 0.0380882
R49616 DVSS.n6155 DVSS.n6154 0.0380882
R49617 DVSS.n6154 DVSS.n6153 0.0380882
R49618 DVSS.n6153 DVSS.n5955 0.0380882
R49619 DVSS.n6143 DVSS.n5955 0.0380882
R49620 DVSS.n6143 DVSS.n6142 0.0380882
R49621 DVSS.n6142 DVSS.n6141 0.0380882
R49622 DVSS.n6141 DVSS.n5957 0.0380882
R49623 DVSS.n6131 DVSS.n5957 0.0380882
R49624 DVSS.n6131 DVSS.n6130 0.0380882
R49625 DVSS.n6130 DVSS.n6129 0.0380882
R49626 DVSS.n6129 DVSS.n5959 0.0380882
R49627 DVSS.n6119 DVSS.n5959 0.0380882
R49628 DVSS.n6119 DVSS.n6118 0.0380882
R49629 DVSS.n6118 DVSS.n6117 0.0380882
R49630 DVSS.n6117 DVSS.n5961 0.0380882
R49631 DVSS.n6107 DVSS.n5961 0.0380882
R49632 DVSS.n6107 DVSS.n6106 0.0380882
R49633 DVSS.n6106 DVSS.n6105 0.0380882
R49634 DVSS.n6105 DVSS.n5963 0.0380882
R49635 DVSS.n6095 DVSS.n5963 0.0380882
R49636 DVSS.n6095 DVSS.n6094 0.0380882
R49637 DVSS.n6094 DVSS.n6093 0.0380882
R49638 DVSS.n6093 DVSS.n5965 0.0380882
R49639 DVSS.n6083 DVSS.n5965 0.0380882
R49640 DVSS.n6083 DVSS.n6082 0.0380882
R49641 DVSS.n6082 DVSS.n6081 0.0380882
R49642 DVSS.n6081 DVSS.n5967 0.0380882
R49643 DVSS.n6071 DVSS.n5967 0.0380882
R49644 DVSS.n6071 DVSS.n6070 0.0380882
R49645 DVSS.n6070 DVSS.n6069 0.0380882
R49646 DVSS.n6069 DVSS.n5969 0.0380882
R49647 DVSS.n6059 DVSS.n5969 0.0380882
R49648 DVSS.n6059 DVSS.n6058 0.0380882
R49649 DVSS.n6058 DVSS.n6057 0.0380882
R49650 DVSS.n6057 DVSS.n5971 0.0380882
R49651 DVSS.n6047 DVSS.n5971 0.0380882
R49652 DVSS.n6047 DVSS.n6046 0.0380882
R49653 DVSS.n6046 DVSS.n6045 0.0380882
R49654 DVSS.n6045 DVSS.n5973 0.0380882
R49655 DVSS.n6035 DVSS.n5973 0.0380882
R49656 DVSS.n6035 DVSS.n6034 0.0380882
R49657 DVSS.n6034 DVSS.n6033 0.0380882
R49658 DVSS.n6033 DVSS.n5975 0.0380882
R49659 DVSS.n6023 DVSS.n5975 0.0380882
R49660 DVSS.n6023 DVSS.n6022 0.0380882
R49661 DVSS.n6022 DVSS.n6021 0.0380882
R49662 DVSS.n6021 DVSS.n5977 0.0380882
R49663 DVSS.n6011 DVSS.n5977 0.0380882
R49664 DVSS.n6011 DVSS.n6010 0.0380882
R49665 DVSS.n6010 DVSS.n6009 0.0380882
R49666 DVSS.n6009 DVSS.n5979 0.0380882
R49667 DVSS.n5999 DVSS.n5979 0.0380882
R49668 DVSS.n5999 DVSS.n5998 0.0380882
R49669 DVSS.n5998 DVSS.n5997 0.0380882
R49670 DVSS.n5997 DVSS.n5981 0.0380882
R49671 DVSS.n5987 DVSS.n5981 0.0380882
R49672 DVSS.n5987 DVSS.n5986 0.0380882
R49673 DVSS.n5986 DVSS.n5985 0.0380882
R49674 DVSS.n6228 DVSS.n5940 0.0380882
R49675 DVSS.n6228 DVSS.n5942 0.0380882
R49676 DVSS.n6224 DVSS.n5942 0.0380882
R49677 DVSS.n6224 DVSS.n6220 0.0380882
R49678 DVSS.n6220 DVSS.n6219 0.0380882
R49679 DVSS.n6219 DVSS.n5944 0.0380882
R49680 DVSS.n6212 DVSS.n5944 0.0380882
R49681 DVSS.n6212 DVSS.n6208 0.0380882
R49682 DVSS.n6208 DVSS.n6207 0.0380882
R49683 DVSS.n6207 DVSS.n5946 0.0380882
R49684 DVSS.n6200 DVSS.n5946 0.0380882
R49685 DVSS.n6200 DVSS.n6196 0.0380882
R49686 DVSS.n6196 DVSS.n6195 0.0380882
R49687 DVSS.n6195 DVSS.n5948 0.0380882
R49688 DVSS.n6188 DVSS.n5948 0.0380882
R49689 DVSS.n6188 DVSS.n6184 0.0380882
R49690 DVSS.n6184 DVSS.n6183 0.0380882
R49691 DVSS.n6183 DVSS.n5950 0.0380882
R49692 DVSS.n6176 DVSS.n5950 0.0380882
R49693 DVSS.n6176 DVSS.n6172 0.0380882
R49694 DVSS.n6172 DVSS.n6171 0.0380882
R49695 DVSS.n6171 DVSS.n5952 0.0380882
R49696 DVSS.n6164 DVSS.n5952 0.0380882
R49697 DVSS.n6164 DVSS.n6160 0.0380882
R49698 DVSS.n6160 DVSS.n6159 0.0380882
R49699 DVSS.n6159 DVSS.n5954 0.0380882
R49700 DVSS.n6152 DVSS.n5954 0.0380882
R49701 DVSS.n6152 DVSS.n6148 0.0380882
R49702 DVSS.n6148 DVSS.n6147 0.0380882
R49703 DVSS.n6147 DVSS.n5956 0.0380882
R49704 DVSS.n6140 DVSS.n5956 0.0380882
R49705 DVSS.n6140 DVSS.n6136 0.0380882
R49706 DVSS.n6136 DVSS.n6135 0.0380882
R49707 DVSS.n6135 DVSS.n5958 0.0380882
R49708 DVSS.n6128 DVSS.n5958 0.0380882
R49709 DVSS.n6128 DVSS.n6124 0.0380882
R49710 DVSS.n6124 DVSS.n6123 0.0380882
R49711 DVSS.n6123 DVSS.n5960 0.0380882
R49712 DVSS.n6116 DVSS.n5960 0.0380882
R49713 DVSS.n6116 DVSS.n6112 0.0380882
R49714 DVSS.n6112 DVSS.n6111 0.0380882
R49715 DVSS.n6111 DVSS.n5962 0.0380882
R49716 DVSS.n6104 DVSS.n5962 0.0380882
R49717 DVSS.n6104 DVSS.n6100 0.0380882
R49718 DVSS.n6100 DVSS.n6099 0.0380882
R49719 DVSS.n6099 DVSS.n5964 0.0380882
R49720 DVSS.n6092 DVSS.n5964 0.0380882
R49721 DVSS.n6092 DVSS.n6088 0.0380882
R49722 DVSS.n6088 DVSS.n6087 0.0380882
R49723 DVSS.n6087 DVSS.n5966 0.0380882
R49724 DVSS.n6080 DVSS.n5966 0.0380882
R49725 DVSS.n6080 DVSS.n6076 0.0380882
R49726 DVSS.n6076 DVSS.n6075 0.0380882
R49727 DVSS.n6075 DVSS.n5968 0.0380882
R49728 DVSS.n6068 DVSS.n5968 0.0380882
R49729 DVSS.n6068 DVSS.n6064 0.0380882
R49730 DVSS.n6064 DVSS.n6063 0.0380882
R49731 DVSS.n6063 DVSS.n5970 0.0380882
R49732 DVSS.n6056 DVSS.n5970 0.0380882
R49733 DVSS.n6056 DVSS.n6052 0.0380882
R49734 DVSS.n6052 DVSS.n6051 0.0380882
R49735 DVSS.n6051 DVSS.n5972 0.0380882
R49736 DVSS.n6044 DVSS.n5972 0.0380882
R49737 DVSS.n6044 DVSS.n6040 0.0380882
R49738 DVSS.n6040 DVSS.n6039 0.0380882
R49739 DVSS.n6039 DVSS.n5974 0.0380882
R49740 DVSS.n6032 DVSS.n5974 0.0380882
R49741 DVSS.n6032 DVSS.n6028 0.0380882
R49742 DVSS.n6028 DVSS.n6027 0.0380882
R49743 DVSS.n6027 DVSS.n5976 0.0380882
R49744 DVSS.n6020 DVSS.n5976 0.0380882
R49745 DVSS.n6020 DVSS.n6016 0.0380882
R49746 DVSS.n6016 DVSS.n6015 0.0380882
R49747 DVSS.n6015 DVSS.n5978 0.0380882
R49748 DVSS.n6008 DVSS.n5978 0.0380882
R49749 DVSS.n6008 DVSS.n6004 0.0380882
R49750 DVSS.n6004 DVSS.n6003 0.0380882
R49751 DVSS.n6003 DVSS.n5980 0.0380882
R49752 DVSS.n5996 DVSS.n5980 0.0380882
R49753 DVSS.n5996 DVSS.n5992 0.0380882
R49754 DVSS.n5992 DVSS.n5991 0.0380882
R49755 DVSS.n5991 DVSS.n5982 0.0380882
R49756 DVSS.n5984 DVSS.n5982 0.0380882
R49757 DVSS.n11733 DVSS.n11730 0.0380882
R49758 DVSS.n11736 DVSS.n11733 0.0380882
R49759 DVSS.n11740 DVSS.n11736 0.0380882
R49760 DVSS.n11744 DVSS.n11740 0.0380882
R49761 DVSS.n11744 DVSS.n11728 0.0380882
R49762 DVSS.n11748 DVSS.n11728 0.0380882
R49763 DVSS.n11752 DVSS.n11748 0.0380882
R49764 DVSS.n11756 DVSS.n11752 0.0380882
R49765 DVSS.n11756 DVSS.n11726 0.0380882
R49766 DVSS.n11760 DVSS.n11726 0.0380882
R49767 DVSS.n11764 DVSS.n11760 0.0380882
R49768 DVSS.n11768 DVSS.n11764 0.0380882
R49769 DVSS.n11768 DVSS.n11724 0.0380882
R49770 DVSS.n11772 DVSS.n11724 0.0380882
R49771 DVSS.n11776 DVSS.n11772 0.0380882
R49772 DVSS.n11780 DVSS.n11776 0.0380882
R49773 DVSS.n11780 DVSS.n11722 0.0380882
R49774 DVSS.n11784 DVSS.n11722 0.0380882
R49775 DVSS.n11788 DVSS.n11784 0.0380882
R49776 DVSS.n11792 DVSS.n11788 0.0380882
R49777 DVSS.n11792 DVSS.n11720 0.0380882
R49778 DVSS.n11796 DVSS.n11720 0.0380882
R49779 DVSS.n11800 DVSS.n11796 0.0380882
R49780 DVSS.n11804 DVSS.n11800 0.0380882
R49781 DVSS.n11804 DVSS.n11718 0.0380882
R49782 DVSS.n11808 DVSS.n11718 0.0380882
R49783 DVSS.n11812 DVSS.n11808 0.0380882
R49784 DVSS.n11816 DVSS.n11812 0.0380882
R49785 DVSS.n11816 DVSS.n11716 0.0380882
R49786 DVSS.n11820 DVSS.n11716 0.0380882
R49787 DVSS.n11824 DVSS.n11820 0.0380882
R49788 DVSS.n11828 DVSS.n11824 0.0380882
R49789 DVSS.n11828 DVSS.n11714 0.0380882
R49790 DVSS.n11832 DVSS.n11714 0.0380882
R49791 DVSS.n11836 DVSS.n11832 0.0380882
R49792 DVSS.n11840 DVSS.n11836 0.0380882
R49793 DVSS.n11840 DVSS.n11712 0.0380882
R49794 DVSS.n11844 DVSS.n11712 0.0380882
R49795 DVSS.n11848 DVSS.n11844 0.0380882
R49796 DVSS.n11852 DVSS.n11848 0.0380882
R49797 DVSS.n11852 DVSS.n11710 0.0380882
R49798 DVSS.n11856 DVSS.n11710 0.0380882
R49799 DVSS.n11860 DVSS.n11856 0.0380882
R49800 DVSS.n11864 DVSS.n11860 0.0380882
R49801 DVSS.n11864 DVSS.n11708 0.0380882
R49802 DVSS.n11868 DVSS.n11708 0.0380882
R49803 DVSS.n11872 DVSS.n11868 0.0380882
R49804 DVSS.n11876 DVSS.n11872 0.0380882
R49805 DVSS.n11876 DVSS.n11706 0.0380882
R49806 DVSS.n11880 DVSS.n11706 0.0380882
R49807 DVSS.n11884 DVSS.n11880 0.0380882
R49808 DVSS.n11888 DVSS.n11884 0.0380882
R49809 DVSS.n11888 DVSS.n11704 0.0380882
R49810 DVSS.n11892 DVSS.n11704 0.0380882
R49811 DVSS.n11896 DVSS.n11892 0.0380882
R49812 DVSS.n11900 DVSS.n11896 0.0380882
R49813 DVSS.n11900 DVSS.n11702 0.0380882
R49814 DVSS.n11904 DVSS.n11702 0.0380882
R49815 DVSS.n11908 DVSS.n11904 0.0380882
R49816 DVSS.n11912 DVSS.n11908 0.0380882
R49817 DVSS.n11912 DVSS.n11700 0.0380882
R49818 DVSS.n11916 DVSS.n11700 0.0380882
R49819 DVSS.n11920 DVSS.n11916 0.0380882
R49820 DVSS.n11924 DVSS.n11920 0.0380882
R49821 DVSS.n11924 DVSS.n11698 0.0380882
R49822 DVSS.n11928 DVSS.n11698 0.0380882
R49823 DVSS.n11932 DVSS.n11928 0.0380882
R49824 DVSS.n11936 DVSS.n11932 0.0380882
R49825 DVSS.n11936 DVSS.n11696 0.0380882
R49826 DVSS.n11940 DVSS.n11696 0.0380882
R49827 DVSS.n11944 DVSS.n11940 0.0380882
R49828 DVSS.n11948 DVSS.n11944 0.0380882
R49829 DVSS.n11948 DVSS.n11694 0.0380882
R49830 DVSS.n11952 DVSS.n11694 0.0380882
R49831 DVSS.n11956 DVSS.n11952 0.0380882
R49832 DVSS.n11960 DVSS.n11956 0.0380882
R49833 DVSS.n11960 DVSS.n11692 0.0380882
R49834 DVSS.n11964 DVSS.n11692 0.0380882
R49835 DVSS.n11968 DVSS.n11964 0.0380882
R49836 DVSS.n11972 DVSS.n11968 0.0380882
R49837 DVSS.n11972 DVSS.n11690 0.0380882
R49838 DVSS.n11977 DVSS.n11690 0.0380882
R49839 DVSS.n11978 DVSS.n11977 0.0380882
R49840 DVSS.n12090 DVSS.n12087 0.0380882
R49841 DVSS.n12093 DVSS.n12090 0.0380882
R49842 DVSS.n12097 DVSS.n12093 0.0380882
R49843 DVSS.n12101 DVSS.n12097 0.0380882
R49844 DVSS.n12101 DVSS.n12085 0.0380882
R49845 DVSS.n12105 DVSS.n12085 0.0380882
R49846 DVSS.n12109 DVSS.n12105 0.0380882
R49847 DVSS.n12113 DVSS.n12109 0.0380882
R49848 DVSS.n12113 DVSS.n12083 0.0380882
R49849 DVSS.n12117 DVSS.n12083 0.0380882
R49850 DVSS.n12121 DVSS.n12117 0.0380882
R49851 DVSS.n12125 DVSS.n12121 0.0380882
R49852 DVSS.n12125 DVSS.n12081 0.0380882
R49853 DVSS.n12129 DVSS.n12081 0.0380882
R49854 DVSS.n12133 DVSS.n12129 0.0380882
R49855 DVSS.n12137 DVSS.n12133 0.0380882
R49856 DVSS.n12137 DVSS.n12079 0.0380882
R49857 DVSS.n12141 DVSS.n12079 0.0380882
R49858 DVSS.n12145 DVSS.n12141 0.0380882
R49859 DVSS.n12149 DVSS.n12145 0.0380882
R49860 DVSS.n12149 DVSS.n12077 0.0380882
R49861 DVSS.n12153 DVSS.n12077 0.0380882
R49862 DVSS.n12157 DVSS.n12153 0.0380882
R49863 DVSS.n12161 DVSS.n12157 0.0380882
R49864 DVSS.n12161 DVSS.n12075 0.0380882
R49865 DVSS.n12165 DVSS.n12075 0.0380882
R49866 DVSS.n12169 DVSS.n12165 0.0380882
R49867 DVSS.n12173 DVSS.n12169 0.0380882
R49868 DVSS.n12173 DVSS.n12073 0.0380882
R49869 DVSS.n12177 DVSS.n12073 0.0380882
R49870 DVSS.n12181 DVSS.n12177 0.0380882
R49871 DVSS.n12185 DVSS.n12181 0.0380882
R49872 DVSS.n12185 DVSS.n12071 0.0380882
R49873 DVSS.n12189 DVSS.n12071 0.0380882
R49874 DVSS.n12193 DVSS.n12189 0.0380882
R49875 DVSS.n12197 DVSS.n12193 0.0380882
R49876 DVSS.n12197 DVSS.n12069 0.0380882
R49877 DVSS.n12201 DVSS.n12069 0.0380882
R49878 DVSS.n12205 DVSS.n12201 0.0380882
R49879 DVSS.n12209 DVSS.n12205 0.0380882
R49880 DVSS.n12209 DVSS.n12067 0.0380882
R49881 DVSS.n12213 DVSS.n12067 0.0380882
R49882 DVSS.n12217 DVSS.n12213 0.0380882
R49883 DVSS.n12221 DVSS.n12217 0.0380882
R49884 DVSS.n12221 DVSS.n12065 0.0380882
R49885 DVSS.n12225 DVSS.n12065 0.0380882
R49886 DVSS.n12229 DVSS.n12225 0.0380882
R49887 DVSS.n12233 DVSS.n12229 0.0380882
R49888 DVSS.n12233 DVSS.n12063 0.0380882
R49889 DVSS.n12237 DVSS.n12063 0.0380882
R49890 DVSS.n12241 DVSS.n12237 0.0380882
R49891 DVSS.n12245 DVSS.n12241 0.0380882
R49892 DVSS.n12245 DVSS.n12061 0.0380882
R49893 DVSS.n12249 DVSS.n12061 0.0380882
R49894 DVSS.n12253 DVSS.n12249 0.0380882
R49895 DVSS.n12257 DVSS.n12253 0.0380882
R49896 DVSS.n12257 DVSS.n12059 0.0380882
R49897 DVSS.n12261 DVSS.n12059 0.0380882
R49898 DVSS.n12265 DVSS.n12261 0.0380882
R49899 DVSS.n12269 DVSS.n12265 0.0380882
R49900 DVSS.n12269 DVSS.n12057 0.0380882
R49901 DVSS.n12273 DVSS.n12057 0.0380882
R49902 DVSS.n12277 DVSS.n12273 0.0380882
R49903 DVSS.n12281 DVSS.n12277 0.0380882
R49904 DVSS.n12281 DVSS.n12055 0.0380882
R49905 DVSS.n12285 DVSS.n12055 0.0380882
R49906 DVSS.n12289 DVSS.n12285 0.0380882
R49907 DVSS.n12293 DVSS.n12289 0.0380882
R49908 DVSS.n12293 DVSS.n12053 0.0380882
R49909 DVSS.n12297 DVSS.n12053 0.0380882
R49910 DVSS.n12301 DVSS.n12297 0.0380882
R49911 DVSS.n12305 DVSS.n12301 0.0380882
R49912 DVSS.n12305 DVSS.n12051 0.0380882
R49913 DVSS.n12309 DVSS.n12051 0.0380882
R49914 DVSS.n12313 DVSS.n12309 0.0380882
R49915 DVSS.n12317 DVSS.n12313 0.0380882
R49916 DVSS.n12317 DVSS.n12049 0.0380882
R49917 DVSS.n12321 DVSS.n12049 0.0380882
R49918 DVSS.n12325 DVSS.n12321 0.0380882
R49919 DVSS.n12329 DVSS.n12325 0.0380882
R49920 DVSS.n12329 DVSS.n12046 0.0380882
R49921 DVSS.n12333 DVSS.n12046 0.0380882
R49922 DVSS.n12334 DVSS.n12333 0.0380882
R49923 DVSS.n12091 DVSS.n12000 0.0380882
R49924 DVSS.n12092 DVSS.n12091 0.0380882
R49925 DVSS.n12092 DVSS.n12086 0.0380882
R49926 DVSS.n12102 DVSS.n12086 0.0380882
R49927 DVSS.n12103 DVSS.n12102 0.0380882
R49928 DVSS.n12104 DVSS.n12103 0.0380882
R49929 DVSS.n12104 DVSS.n12084 0.0380882
R49930 DVSS.n12114 DVSS.n12084 0.0380882
R49931 DVSS.n12115 DVSS.n12114 0.0380882
R49932 DVSS.n12116 DVSS.n12115 0.0380882
R49933 DVSS.n12116 DVSS.n12082 0.0380882
R49934 DVSS.n12126 DVSS.n12082 0.0380882
R49935 DVSS.n12127 DVSS.n12126 0.0380882
R49936 DVSS.n12128 DVSS.n12127 0.0380882
R49937 DVSS.n12128 DVSS.n12080 0.0380882
R49938 DVSS.n12138 DVSS.n12080 0.0380882
R49939 DVSS.n12139 DVSS.n12138 0.0380882
R49940 DVSS.n12140 DVSS.n12139 0.0380882
R49941 DVSS.n12140 DVSS.n12078 0.0380882
R49942 DVSS.n12150 DVSS.n12078 0.0380882
R49943 DVSS.n12151 DVSS.n12150 0.0380882
R49944 DVSS.n12152 DVSS.n12151 0.0380882
R49945 DVSS.n12152 DVSS.n12076 0.0380882
R49946 DVSS.n12162 DVSS.n12076 0.0380882
R49947 DVSS.n12163 DVSS.n12162 0.0380882
R49948 DVSS.n12164 DVSS.n12163 0.0380882
R49949 DVSS.n12164 DVSS.n12074 0.0380882
R49950 DVSS.n12174 DVSS.n12074 0.0380882
R49951 DVSS.n12175 DVSS.n12174 0.0380882
R49952 DVSS.n12176 DVSS.n12175 0.0380882
R49953 DVSS.n12176 DVSS.n12072 0.0380882
R49954 DVSS.n12186 DVSS.n12072 0.0380882
R49955 DVSS.n12187 DVSS.n12186 0.0380882
R49956 DVSS.n12188 DVSS.n12187 0.0380882
R49957 DVSS.n12188 DVSS.n12070 0.0380882
R49958 DVSS.n12198 DVSS.n12070 0.0380882
R49959 DVSS.n12199 DVSS.n12198 0.0380882
R49960 DVSS.n12200 DVSS.n12199 0.0380882
R49961 DVSS.n12200 DVSS.n12068 0.0380882
R49962 DVSS.n12210 DVSS.n12068 0.0380882
R49963 DVSS.n12211 DVSS.n12210 0.0380882
R49964 DVSS.n12212 DVSS.n12211 0.0380882
R49965 DVSS.n12212 DVSS.n12066 0.0380882
R49966 DVSS.n12222 DVSS.n12066 0.0380882
R49967 DVSS.n12223 DVSS.n12222 0.0380882
R49968 DVSS.n12224 DVSS.n12223 0.0380882
R49969 DVSS.n12224 DVSS.n12064 0.0380882
R49970 DVSS.n12234 DVSS.n12064 0.0380882
R49971 DVSS.n12235 DVSS.n12234 0.0380882
R49972 DVSS.n12236 DVSS.n12235 0.0380882
R49973 DVSS.n12236 DVSS.n12062 0.0380882
R49974 DVSS.n12246 DVSS.n12062 0.0380882
R49975 DVSS.n12247 DVSS.n12246 0.0380882
R49976 DVSS.n12248 DVSS.n12247 0.0380882
R49977 DVSS.n12248 DVSS.n12060 0.0380882
R49978 DVSS.n12258 DVSS.n12060 0.0380882
R49979 DVSS.n12259 DVSS.n12258 0.0380882
R49980 DVSS.n12260 DVSS.n12259 0.0380882
R49981 DVSS.n12260 DVSS.n12058 0.0380882
R49982 DVSS.n12270 DVSS.n12058 0.0380882
R49983 DVSS.n12271 DVSS.n12270 0.0380882
R49984 DVSS.n12272 DVSS.n12271 0.0380882
R49985 DVSS.n12272 DVSS.n12056 0.0380882
R49986 DVSS.n12282 DVSS.n12056 0.0380882
R49987 DVSS.n12283 DVSS.n12282 0.0380882
R49988 DVSS.n12284 DVSS.n12283 0.0380882
R49989 DVSS.n12284 DVSS.n12054 0.0380882
R49990 DVSS.n12294 DVSS.n12054 0.0380882
R49991 DVSS.n12295 DVSS.n12294 0.0380882
R49992 DVSS.n12296 DVSS.n12295 0.0380882
R49993 DVSS.n12296 DVSS.n12052 0.0380882
R49994 DVSS.n12306 DVSS.n12052 0.0380882
R49995 DVSS.n12307 DVSS.n12306 0.0380882
R49996 DVSS.n12308 DVSS.n12307 0.0380882
R49997 DVSS.n12308 DVSS.n12050 0.0380882
R49998 DVSS.n12318 DVSS.n12050 0.0380882
R49999 DVSS.n12319 DVSS.n12318 0.0380882
R50000 DVSS.n12320 DVSS.n12319 0.0380882
R50001 DVSS.n12320 DVSS.n12048 0.0380882
R50002 DVSS.n12330 DVSS.n12048 0.0380882
R50003 DVSS.n12331 DVSS.n12330 0.0380882
R50004 DVSS.n12332 DVSS.n12331 0.0380882
R50005 DVSS.n12332 DVSS.n11988 0.0380882
R50006 DVSS.n18927 DVSS.n14552 0.0357174
R50007 DVSS.n20687 DVSS.n20686 0.0357174
R50008 DVSS.n20137 DVSS.n14589 0.0357174
R50009 DVSS.n20034 DVSS.n14600 0.0357174
R50010 DVSS.n20253 DVSS.n14642 0.0357174
R50011 DVSS.n20290 DVSS.n14637 0.0357174
R50012 DVSS.n20633 DVSS.n20632 0.0357174
R50013 DVSS.n20412 DVSS.n20376 0.0357174
R50014 DVSS.n18939 DVSS.n14519 0.0357174
R50015 DVSS.n20698 DVSS.n14535 0.0357174
R50016 DVSS.n20082 DVSS.n20014 0.0357174
R50017 DVSS.n20036 DVSS.n20025 0.0357174
R50018 DVSS.n20264 DVSS.n20187 0.0357174
R50019 DVSS.n20241 DVSS.n14869 0.0357174
R50020 DVSS.n20325 DVSS.n20323 0.0357174
R50021 DVSS.n20381 DVSS.n14860 0.0357174
R50022 DVSS.n22585 DVSS.n752 0.034437
R50023 DVSS.n22936 DVSS.n434 0.034437
R50024 DVSS.n22625 DVSS.n737 0.0339884
R50025 DVSS.n22896 DVSS.n449 0.0339884
R50026 DVSS.n19915 DVSS.n19914 0.0337188
R50027 DVSS.n18528 DVSS.n18527 0.0337188
R50028 DVSS.n18528 DVSS.n15144 0.0337188
R50029 DVSS.n19914 DVSS.n15141 0.0337188
R50030 DVSS.n13018 DVSS.t85 0.03326
R50031 DVSS.n13018 DVSS.t5 0.03326
R50032 DVSS.n19891 DVSS.t51 0.03326
R50033 DVSS.n19891 DVSS.t141 0.03326
R50034 DVSS.n19886 DVSS.t25 0.03326
R50035 DVSS.n19886 DVSS.t153 0.03326
R50036 DVSS.n19048 DVSS.t73 0.03326
R50037 DVSS.n19048 DVSS.t15 0.03326
R50038 DVSS.n19878 DVSS.t101 0.03326
R50039 DVSS.n19878 DVSS.t143 0.03326
R50040 DVSS.n19873 DVSS.t113 0.03326
R50041 DVSS.n19873 DVSS.t3 0.03326
R50042 DVSS.n19056 DVSS.t133 0.03326
R50043 DVSS.n19056 DVSS.t17 0.03326
R50044 DVSS.n19865 DVSS.t103 0.03326
R50045 DVSS.n19865 DVSS.t77 0.03326
R50046 DVSS.n19860 DVSS.t123 0.03326
R50047 DVSS.n19860 DVSS.t89 0.03326
R50048 DVSS.n19064 DVSS.t135 0.03326
R50049 DVSS.n19064 DVSS.t57 0.03326
R50050 DVSS.n19584 DVSS.t35 0.03326
R50051 DVSS.n19584 DVSS.t91 0.03326
R50052 DVSS.n19579 DVSS.t55 0.03326
R50053 DVSS.n19579 DVSS.t109 0.03326
R50054 DVSS.n19524 DVSS.t27 0.03326
R50055 DVSS.n19524 DVSS.t43 0.03326
R50056 DVSS.n19571 DVSS.t137 0.03326
R50057 DVSS.n19571 DVSS.t59 0.03326
R50058 DVSS.n19566 DVSS.t145 0.03326
R50059 DVSS.n19566 DVSS.t79 0.03326
R50060 DVSS.n19532 DVSS.t7 0.03326
R50061 DVSS.n19532 DVSS.t93 0.03326
R50062 DVSS.n19558 DVSS.t23 0.03326
R50063 DVSS.n19558 DVSS.t117 0.03326
R50064 DVSS.n19553 DVSS.t159 0.03326
R50065 DVSS.n19553 DVSS.t127 0.03326
R50066 DVSS.n19540 DVSS.t39 0.03326
R50067 DVSS.n19540 DVSS.t147 0.03326
R50068 DVSS.n21832 DVSS.t75 0.03326
R50069 DVSS.n21832 DVSS.t131 0.03326
R50070 DVSS.n21840 DVSS.t105 0.03326
R50071 DVSS.n21840 DVSS.t19 0.03326
R50072 DVSS.n21826 DVSS.t115 0.03326
R50073 DVSS.n21826 DVSS.t29 0.03326
R50074 DVSS.n21847 DVSS.t87 0.03326
R50075 DVSS.n21847 DVSS.t45 0.03326
R50076 DVSS.n21948 DVSS.t107 0.03326
R50077 DVSS.n21948 DVSS.t63 0.03326
R50078 DVSS.n21937 DVSS.t125 0.03326
R50079 DVSS.n21937 DVSS.t37 0.03326
R50080 DVSS.n21915 DVSS.t11 0.03326
R50081 DVSS.n21915 DVSS.t47 0.03326
R50082 DVSS.n21905 DVSS.t31 0.03326
R50083 DVSS.n21905 DVSS.t81 0.03326
R50084 DVSS.n21895 DVSS.t161 0.03326
R50085 DVSS.n21895 DVSS.t95 0.03326
R50086 DVSS.n845 DVSS.t119 0.03326
R50087 DVSS.n845 DVSS.t83 0.03326
R50088 DVSS.n836 DVSS.t139 0.03326
R50089 DVSS.n836 DVSS.t49 0.03326
R50090 DVSS.n827 DVSS.t149 0.03326
R50091 DVSS.n827 DVSS.t69 0.03326
R50092 DVSS.n818 DVSS.t9 0.03326
R50093 DVSS.n818 DVSS.t97 0.03326
R50094 DVSS.n22480 DVSS.t13 0.03326
R50095 DVSS.n22480 DVSS.t111 0.03326
R50096 DVSS.n13044 DVSS.t33 0.03326
R50097 DVSS.n13044 DVSS.t129 0.03326
R50098 DVSS.n13032 DVSS.t41 0.03326
R50099 DVSS.n13032 DVSS.t99 0.03326
R50100 DVSS.n13053 DVSS.t71 0.03326
R50101 DVSS.n13053 DVSS.t151 0.03326
R50102 DVSS.n21174 DVSS.n13667 0.0329
R50103 DVSS.n13667 DVSS.n13661 0.0329
R50104 DVSS.n21178 DVSS.n13661 0.0329
R50105 DVSS.n21178 DVSS.n21177 0.0329
R50106 DVSS.n18525 DVSS.n15147 0.0329
R50107 DVSS.n18521 DVSS.n15147 0.0329
R50108 DVSS.n18521 DVSS.n18520 0.0329
R50109 DVSS.n18520 DVSS.n18519 0.0329
R50110 DVSS.n17788 DVSS.n17787 0.0329
R50111 DVSS.n18171 DVSS.n18170 0.0329
R50112 DVSS.n19917 DVSS.n15139 0.0329
R50113 DVSS.n19921 DVSS.n15139 0.0329
R50114 DVSS.n19922 DVSS.n19921 0.0329
R50115 DVSS.n19923 DVSS.n19922 0.0329
R50116 DVSS.n18929 DVSS.n14565 0.0327826
R50117 DVSS.n18975 DVSS.n14567 0.0327826
R50118 DVSS.n20069 DVSS.n14598 0.0327826
R50119 DVSS.n20032 DVSS.n14587 0.0327826
R50120 DVSS.n20255 DVSS.n14639 0.0327826
R50121 DVSS.n20239 DVSS.n14644 0.0327826
R50122 DVSS.n20631 DVSS.n14669 0.0327826
R50123 DVSS.n20401 DVSS.n20400 0.0327826
R50124 DVSS.n18933 DVSS.n14532 0.0327826
R50125 DVSS.n18922 DVSS.n14534 0.0327826
R50126 DVSS.n20080 DVSS.n20023 0.0327826
R50127 DVSS.n20065 DVSS.n20012 0.0327826
R50128 DVSS.n20259 DVSS.n14871 0.0327826
R50129 DVSS.n20243 DVSS.n20189 0.0327826
R50130 DVSS.n20324 DVSS.n14862 0.0327826
R50131 DVSS.n20391 DVSS.n20327 0.0327826
R50132 DVSS.n17051 DVSS.n17050 0.032527
R50133 DVSS.n16980 DVSS.n16979 0.032527
R50134 DVSS.n17116 DVSS.n17115 0.032527
R50135 DVSS.n17528 DVSS.n16920 0.032527
R50136 DVSS.n6675 DVSS.n6674 0.03245
R50137 DVSS.n6676 DVSS.n6675 0.03245
R50138 DVSS.n6693 DVSS.n6692 0.03245
R50139 DVSS.n7030 DVSS.n6693 0.03245
R50140 DVSS.n7028 DVSS.n5864 0.03245
R50141 DVSS.n7051 DVSS.n5522 0.03245
R50142 DVSS.n7072 DVSS.n5522 0.03245
R50143 DVSS.n7075 DVSS.n7074 0.03245
R50144 DVSS.n7074 DVSS.n5173 0.03245
R50145 DVSS.n7094 DVSS.n4829 0.03245
R50146 DVSS.n7455 DVSS.n4829 0.03245
R50147 DVSS.n7457 DVSS.n4815 0.03245
R50148 DVSS.n7810 DVSS.n4815 0.03245
R50149 DVSS.n7812 DVSS.n4463 0.03245
R50150 DVSS.n7830 DVSS.n4463 0.03245
R50151 DVSS.n7833 DVSS.n7832 0.03245
R50152 DVSS.n7837 DVSS.n4359 0.03245
R50153 DVSS.n8106 DVSS.n4359 0.03245
R50154 DVSS.n8108 DVSS.n3853 0.03245
R50155 DVSS.n8324 DVSS.n3853 0.03245
R50156 DVSS.n8328 DVSS.n8326 0.03245
R50157 DVSS.n8328 DVSS.n8327 0.03245
R50158 DVSS.n8594 DVSS.n8593 0.03245
R50159 DVSS.n8596 DVSS.n8594 0.03245
R50160 DVSS.n8619 DVSS.n3403 0.03245
R50161 DVSS.n8621 DVSS.n3056 0.03245
R50162 DVSS.n8973 DVSS.n3056 0.03245
R50163 DVSS.n8975 DVSS.n2885 0.03245
R50164 DVSS.n9191 DVSS.n2885 0.03245
R50165 DVSS.n9195 DVSS.n9193 0.03245
R50166 DVSS.n9195 DVSS.n9194 0.03245
R50167 DVSS.n9461 DVSS.n9460 0.03245
R50168 DVSS.n9462 DVSS.n9461 0.03245
R50169 DVSS.n9775 DVSS.n9774 0.03245
R50170 DVSS.n10112 DVSS.n9775 0.03245
R50171 DVSS.n10110 DVSS.n2702 0.03245
R50172 DVSS.n10133 DVSS.n2703 0.03245
R50173 DVSS.n2703 DVSS.n2360 0.03245
R50174 DVSS.n10158 DVSS.n2361 0.03245
R50175 DVSS.n2361 DVSS.n2016 0.03245
R50176 DVSS.n10467 DVSS.n1624 0.03245
R50177 DVSS.n10490 DVSS.n1624 0.03245
R50178 DVSS.n10492 DVSS.n1518 0.03245
R50179 DVSS.n10758 DVSS.n1518 0.03245
R50180 DVSS.n13355 DVSS.n10760 0.03245
R50181 DVSS.n13353 DVSS.n10762 0.03245
R50182 DVSS.n11451 DVSS.n10762 0.03245
R50183 DVSS.n13332 DVSS.n13331 0.03245
R50184 DVSS.n13331 DVSS.n13330 0.03245
R50185 DVSS.n11640 DVSS.n11637 0.03245
R50186 DVSS.n11985 DVSS.n11637 0.03245
R50187 DVSS.n13117 DVSS.n11987 0.03245
R50188 DVSS.n13117 DVSS.n13116 0.03245
R50189 DVSS.n13114 DVSS.n11989 0.03245
R50190 DVSS.n12764 DVSS.n11989 0.03245
R50191 DVSS.n17259 DVSS.n17138 0.0320219
R50192 DVSS.n17224 DVSS.n17173 0.0320219
R50193 DVSS.n17302 DVSS.n17301 0.0320219
R50194 DVSS.n17426 DVSS.n17425 0.0320219
R50195 DVSS.n7052 DVSS.n5864 0.031775
R50196 DVSS.n13126 DVSS.n11624 0.0317353
R50197 DVSS.n5622 DVSS.n5528 0.0317353
R50198 DVSS.n5270 DVSS.n5179 0.0317353
R50199 DVSS.n4931 DVSS.n4837 0.0317353
R50200 DVSS.n7447 DVSS.n7444 0.0317353
R50201 DVSS.n7802 DVSS.n4821 0.0317353
R50202 DVSS.n7822 DVSS.n4807 0.0317353
R50203 DVSS.n8095 DVSS.n4365 0.0317353
R50204 DVSS.n8116 DVSS.n4017 0.0317353
R50205 DVSS.n8130 DVSS.n8129 0.0317353
R50206 DVSS.n8340 DVSS.n3843 0.0317353
R50207 DVSS.n8609 DVSS.n3409 0.0317353
R50208 DVSS.n8629 DVSS.n3062 0.0317353
R50209 DVSS.n8983 DVSS.n3048 0.0317353
R50210 DVSS.n8997 DVSS.n8996 0.0317353
R50211 DVSS.n9207 DVSS.n2875 0.0317353
R50212 DVSS.n9764 DVSS.n2733 0.0317353
R50213 DVSS.n10120 DVSS.n2712 0.0317353
R50214 DVSS.n2460 DVSS.n2367 0.0317353
R50215 DVSS.n2118 DVSS.n2024 0.0317353
R50216 DVSS.n10456 DVSS.n10455 0.0317353
R50217 DVSS.n1669 DVSS.n1616 0.0317353
R50218 DVSS.n10507 DVSS.n1612 0.0317353
R50219 DVSS.n11105 DVSS.n11104 0.0317353
R50220 DVSS.n11262 DVSS.n11106 0.0317353
R50221 DVSS.n13136 DVSS.n13135 0.0317353
R50222 DVSS.n7038 DVSS.n5872 0.0317353
R50223 DVSS.n6684 DVSS.n5893 0.0317353
R50224 DVSS.n12342 DVSS.n12000 0.0317353
R50225 DVSS.n17406 DVSS.n15305 0.0316707
R50226 DVSS.n17414 DVSS.n15372 0.0316707
R50227 DVSS.n17401 DVSS.n15266 0.0316707
R50228 DVSS.n17209 DVSS.n15442 0.0316707
R50229 DVSS.n8620 DVSS.n8619 0.031325
R50230 DVSS.n22624 DVSS.n22623 0.0311977
R50231 DVSS.n22898 DVSS.n22897 0.0311977
R50232 DVSS.n18517 DVSS.n15145 0.0311
R50233 DVSS.n19925 DVSS.n15137 0.0311
R50234 DVSS.n10111 DVSS.n10110 0.030875
R50235 DVSS.n13355 DVSS.n13354 0.030875
R50236 DVSS.n7832 DVSS.n7831 0.030425
R50237 DVSS.n18973 DVSS.n14551 0.0298478
R50238 DVSS.n18976 DVSS.n14566 0.0298478
R50239 DVSS.n20071 DVSS.n14588 0.0298478
R50240 DVSS.n20149 DVSS.n14599 0.0298478
R50241 DVSS.n20278 DVSS.n14643 0.0298478
R50242 DVSS.n20237 DVSS.n14638 0.0298478
R50243 DVSS.n20397 DVSS.n20396 0.0298478
R50244 DVSS.n20402 DVSS.n20399 0.0298478
R50245 DVSS.n18931 DVSS.n14518 0.0298478
R50246 DVSS.n18923 DVSS.n14533 0.0298478
R50247 DVSS.n20075 DVSS.n20013 0.0298478
R50248 DVSS.n20067 DVSS.n20024 0.0298478
R50249 DVSS.n20257 DVSS.n20188 0.0298478
R50250 DVSS.n20249 DVSS.n14870 0.0298478
R50251 DVSS.n20387 DVSS.n20326 0.0298478
R50252 DVSS.n20393 DVSS.n14861 0.0298478
R50253 DVSS.n17015 DVSS.n16976 0.0293889
R50254 DVSS.n16976 DVSS.t190 0.0293889
R50255 DVSS.n17097 DVSS.n16925 0.0293889
R50256 DVSS.t190 DVSS.n16925 0.0293889
R50257 DVSS.n7833 DVSS.n4458 0.028625
R50258 DVSS.n6672 DVSS.n6232 0.0284039
R50259 DVSS.n6678 DVSS.n6232 0.0284039
R50260 DVSS.n6690 DVSS.n5881 0.0284039
R50261 DVSS.n7032 DVSS.n5881 0.0284039
R50262 DVSS.n7046 DVSS.n5866 0.0284039
R50263 DVSS.n7049 DVSS.n5524 0.0284039
R50264 DVSS.n7070 DVSS.n5524 0.0284039
R50265 DVSS.n7077 DVSS.n5175 0.0284039
R50266 DVSS.n7089 DVSS.n5175 0.0284039
R50267 DVSS.n7092 DVSS.n4831 0.0284039
R50268 DVSS.n7453 DVSS.n4831 0.0284039
R50269 DVSS.n7459 DVSS.n4817 0.0284039
R50270 DVSS.n7808 DVSS.n4817 0.0284039
R50271 DVSS.n7814 DVSS.n4466 0.0284039
R50272 DVSS.n7828 DVSS.n4466 0.0284039
R50273 DVSS.n7835 DVSS.n4460 0.0284039
R50274 DVSS.n7839 DVSS.n4361 0.0284039
R50275 DVSS.n8104 DVSS.n4361 0.0284039
R50276 DVSS.n8110 DVSS.n3856 0.0284039
R50277 DVSS.n8322 DVSS.n3856 0.0284039
R50278 DVSS.n8330 DVSS.n3847 0.0284039
R50279 DVSS.n8330 DVSS.n3849 0.0284039
R50280 DVSS.n8591 DVSS.n3754 0.0284039
R50281 DVSS.n3754 DVSS.n3750 0.0284039
R50282 DVSS.n8617 DVSS.n3405 0.0284039
R50283 DVSS.n8623 DVSS.n3058 0.0284039
R50284 DVSS.n8971 DVSS.n3058 0.0284039
R50285 DVSS.n8977 DVSS.n2888 0.0284039
R50286 DVSS.n9189 DVSS.n2888 0.0284039
R50287 DVSS.n9197 DVSS.n2879 0.0284039
R50288 DVSS.n9197 DVSS.n2881 0.0284039
R50289 DVSS.n9458 DVSS.n2782 0.0284039
R50290 DVSS.n9464 DVSS.n2782 0.0284039
R50291 DVSS.n9772 DVSS.n2721 0.0284039
R50292 DVSS.n10114 DVSS.n2721 0.0284039
R50293 DVSS.n10128 DVSS.n2705 0.0284039
R50294 DVSS.n10131 DVSS.n2363 0.0284039
R50295 DVSS.n10153 DVSS.n2363 0.0284039
R50296 DVSS.n10156 DVSS.n2018 0.0284039
R50297 DVSS.n10462 DVSS.n2018 0.0284039
R50298 DVSS.n10465 DVSS.n1626 0.0284039
R50299 DVSS.n10488 DVSS.n1626 0.0284039
R50300 DVSS.n10494 DVSS.n1521 0.0284039
R50301 DVSS.n10756 DVSS.n1521 0.0284039
R50302 DVSS.n13357 DVSS.n1513 0.0284039
R50303 DVSS.n13351 DVSS.n10764 0.0284039
R50304 DVSS.n11447 DVSS.n10764 0.0284039
R50305 DVSS.n11455 DVSS.n11450 0.0284039
R50306 DVSS.n13328 DVSS.n11455 0.0284039
R50307 DVSS.n11644 DVSS.n11642 0.0284039
R50308 DVSS.n11983 DVSS.n11644 0.0284039
R50309 DVSS.n13119 DVSS.n11632 0.0284039
R50310 DVSS.n13119 DVSS.n11633 0.0284039
R50311 DVSS.n13112 DVSS.n11993 0.0284039
R50312 DVSS.n12762 DVSS.n11993 0.0284039
R50313 DVSS.n6673 DVSS.n6233 0.0284039
R50314 DVSS.n6677 DVSS.n6233 0.0284039
R50315 DVSS.n6691 DVSS.n5883 0.0284039
R50316 DVSS.n7031 DVSS.n5883 0.0284039
R50317 DVSS.n7047 DVSS.n5865 0.0284039
R50318 DVSS.n7050 DVSS.n5523 0.0284039
R50319 DVSS.n7071 DVSS.n5523 0.0284039
R50320 DVSS.n7076 DVSS.n5174 0.0284039
R50321 DVSS.n7090 DVSS.n5174 0.0284039
R50322 DVSS.n7093 DVSS.n4830 0.0284039
R50323 DVSS.n7454 DVSS.n4830 0.0284039
R50324 DVSS.n7458 DVSS.n4816 0.0284039
R50325 DVSS.n7809 DVSS.n4816 0.0284039
R50326 DVSS.n7813 DVSS.n4464 0.0284039
R50327 DVSS.n7829 DVSS.n4464 0.0284039
R50328 DVSS.n7834 DVSS.n4461 0.0284039
R50329 DVSS.n7838 DVSS.n4360 0.0284039
R50330 DVSS.n8105 DVSS.n4360 0.0284039
R50331 DVSS.n8109 DVSS.n3854 0.0284039
R50332 DVSS.n8323 DVSS.n3854 0.0284039
R50333 DVSS.n8329 DVSS.n3850 0.0284039
R50334 DVSS.n8329 DVSS.n3851 0.0284039
R50335 DVSS.n8592 DVSS.n3749 0.0284039
R50336 DVSS.n8597 DVSS.n3749 0.0284039
R50337 DVSS.n8618 DVSS.n3404 0.0284039
R50338 DVSS.n8622 DVSS.n3057 0.0284039
R50339 DVSS.n8972 DVSS.n3057 0.0284039
R50340 DVSS.n8976 DVSS.n2886 0.0284039
R50341 DVSS.n9190 DVSS.n2886 0.0284039
R50342 DVSS.n9196 DVSS.n2882 0.0284039
R50343 DVSS.n9196 DVSS.n2883 0.0284039
R50344 DVSS.n9459 DVSS.n2783 0.0284039
R50345 DVSS.n9463 DVSS.n2783 0.0284039
R50346 DVSS.n9773 DVSS.n2723 0.0284039
R50347 DVSS.n10113 DVSS.n2723 0.0284039
R50348 DVSS.n10129 DVSS.n2704 0.0284039
R50349 DVSS.n10132 DVSS.n2362 0.0284039
R50350 DVSS.n10154 DVSS.n2362 0.0284039
R50351 DVSS.n10157 DVSS.n2017 0.0284039
R50352 DVSS.n10463 DVSS.n2017 0.0284039
R50353 DVSS.n10466 DVSS.n1625 0.0284039
R50354 DVSS.n10489 DVSS.n1625 0.0284039
R50355 DVSS.n10493 DVSS.n1519 0.0284039
R50356 DVSS.n10757 DVSS.n1519 0.0284039
R50357 DVSS.n13356 DVSS.n1515 0.0284039
R50358 DVSS.n13352 DVSS.n10763 0.0284039
R50359 DVSS.n11448 DVSS.n10763 0.0284039
R50360 DVSS.n13333 DVSS.n11449 0.0284039
R50361 DVSS.n13329 DVSS.n11449 0.0284039
R50362 DVSS.n11641 DVSS.n11638 0.0284039
R50363 DVSS.n11984 DVSS.n11638 0.0284039
R50364 DVSS.n13118 DVSS.n11634 0.0284039
R50365 DVSS.n13118 DVSS.n11635 0.0284039
R50366 DVSS.n13113 DVSS.n11991 0.0284039
R50367 DVSS.n12763 DVSS.n11991 0.0284039
R50368 DVSS.n16387 DVSS.n16385 0.0284
R50369 DVSS.n16389 DVSS.n16387 0.0284
R50370 DVSS.n16391 DVSS.n16389 0.0284
R50371 DVSS.n16392 DVSS.n16391 0.0284
R50372 DVSS.n16392 DVSS.n16382 0.0284
R50373 DVSS.n16396 DVSS.n16382 0.0284
R50374 DVSS.n16397 DVSS.n16396 0.0284
R50375 DVSS.n16398 DVSS.n16397 0.0284
R50376 DVSS.n16398 DVSS.n16380 0.0284
R50377 DVSS.n16402 DVSS.n16380 0.0284
R50378 DVSS.n16405 DVSS.n16404 0.0284
R50379 DVSS.n16409 DVSS.n16378 0.0284
R50380 DVSS.n16410 DVSS.n16409 0.0284
R50381 DVSS.n16411 DVSS.n16410 0.0284
R50382 DVSS.n16411 DVSS.n16376 0.0284
R50383 DVSS.n16415 DVSS.n16376 0.0284
R50384 DVSS.n16416 DVSS.n16415 0.0284
R50385 DVSS.n16417 DVSS.n16416 0.0284
R50386 DVSS.n16419 DVSS.n16417 0.0284
R50387 DVSS.n16421 DVSS.n16419 0.0284
R50388 DVSS.n16423 DVSS.n16421 0.0284
R50389 DVSS.n16425 DVSS.n16423 0.0284
R50390 DVSS.n16465 DVSS.n16425 0.0284
R50391 DVSS.n15717 DVSS.n15715 0.0284
R50392 DVSS.n15715 DVSS.n15713 0.0284
R50393 DVSS.n15713 DVSS.n15688 0.0284
R50394 DVSS.n18049 DVSS.n15688 0.0284
R50395 DVSS.n18050 DVSS.n18049 0.0284
R50396 DVSS.n18051 DVSS.n18050 0.0284
R50397 DVSS.n18051 DVSS.n15686 0.0284
R50398 DVSS.n18055 DVSS.n15686 0.0284
R50399 DVSS.n18056 DVSS.n18055 0.0284
R50400 DVSS.n18057 DVSS.n18056 0.0284
R50401 DVSS.n18061 DVSS.n18060 0.0284
R50402 DVSS.n18062 DVSS.n15682 0.0284
R50403 DVSS.n18066 DVSS.n15682 0.0284
R50404 DVSS.n18067 DVSS.n18066 0.0284
R50405 DVSS.n18068 DVSS.n18067 0.0284
R50406 DVSS.n18068 DVSS.n15680 0.0284
R50407 DVSS.n18072 DVSS.n15680 0.0284
R50408 DVSS.n18073 DVSS.n18072 0.0284
R50409 DVSS.n18076 DVSS.n18073 0.0284
R50410 DVSS.n18076 DVSS.n18075 0.0284
R50411 DVSS.n18075 DVSS.n15651 0.0284
R50412 DVSS.n18082 DVSS.n15651 0.0284
R50413 DVSS.n18083 DVSS.n18082 0.0284
R50414 DVSS.n18655 DVSS.n18654 0.0283804
R50415 DVSS.n18655 DVSS.n18647 0.0283804
R50416 DVSS.n20503 DVSS.n14703 0.0283804
R50417 DVSS.n18769 DVSS.n18762 0.0283804
R50418 DVSS.n18769 DVSS.n18768 0.0283804
R50419 DVSS.n20466 DVSS.n20465 0.0283804
R50420 DVSS.n10134 DVSS.n2702 0.028175
R50421 DVSS.n10760 DVSS.n10759 0.028175
R50422 DVSS.n7046 DVSS.n5575 0.0278144
R50423 DVSS.n7048 DVSS.n7047 0.0278144
R50424 DVSS.n8595 DVSS.n3403 0.027725
R50425 DVSS.n8617 DVSS.n3067 0.0274214
R50426 DVSS.n8618 DVSS.n3068 0.0274214
R50427 DVSS.n7029 DVSS.n7028 0.027275
R50428 DVSS.n20690 DVSS.n20689 0.0272589
R50429 DVSS.n14560 DVSS.n14547 0.0272589
R50430 DVSS.n14594 DVSS.n14593 0.0272589
R50431 DVSS.n20101 DVSS.n14592 0.0272589
R50432 DVSS.n14648 DVSS.n14634 0.0272589
R50433 DVSS.n20432 DVSS.n20431 0.0272589
R50434 DVSS.n20358 DVSS.n20357 0.0272589
R50435 DVSS.n20696 DVSS.n14523 0.0272589
R50436 DVSS.n14537 DVSS.n14522 0.0272589
R50437 DVSS.n20109 DVSS.n20018 0.0272589
R50438 DVSS.n20114 DVSS.n20017 0.0272589
R50439 DVSS.n20193 DVSS.n14866 0.0272589
R50440 DVSS.n20362 DVSS.n14857 0.0272589
R50441 DVSS.n20352 DVSS.n14856 0.0272589
R50442 DVSS.n21577 DVSS.n21576 0.0272589
R50443 DVSS.n21588 DVSS.n21587 0.0272589
R50444 DVSS.n1332 DVSS.n1331 0.0272589
R50445 DVSS.n1314 DVSS.n1313 0.0272589
R50446 DVSS.n21576 DVSS.n869 0.0272589
R50447 DVSS.n21585 DVSS.n21569 0.0272589
R50448 DVSS.n20102 DVSS.n20101 0.0272589
R50449 DVSS.n20115 DVSS.n20114 0.0272589
R50450 DVSS.n20115 DVSS.n20018 0.0272589
R50451 DVSS.n20102 DVSS.n14594 0.0272589
R50452 DVSS.n22340 DVSS.n1177 0.0272589
R50453 DVSS.n1311 DVSS.n1310 0.0272589
R50454 DVSS.n1293 DVSS.n1292 0.0272589
R50455 DVSS.n1196 DVSS.n1180 0.0272589
R50456 DVSS.n14649 DVSS.n14648 0.0272589
R50457 DVSS.n20315 DVSS.n20193 0.0272589
R50458 DVSS.n22457 DVSS.n866 0.0272589
R50459 DVSS.n1352 DVSS.n1351 0.0272589
R50460 DVSS.n1334 DVSS.n1333 0.0272589
R50461 DVSS.n871 DVSS.n867 0.0272589
R50462 DVSS.n20691 DVSS.n14547 0.0272589
R50463 DVSS.n20695 DVSS.n14522 0.0272589
R50464 DVSS.n20696 DVSS.n20695 0.0272589
R50465 DVSS.n20691 DVSS.n20690 0.0272589
R50466 DVSS.n19504 DVSS.n19270 0.0272589
R50467 DVSS.n19514 DVSS.n19513 0.0272589
R50468 DVSS.n19502 DVSS.n19267 0.0272589
R50469 DVSS.n19087 DVSS.n19078 0.0272589
R50470 DVSS.n19591 DVSS.n19590 0.0272589
R50471 DVSS.n19088 DVSS.n19070 0.0272589
R50472 DVSS.n22337 DVSS.n1198 0.0272589
R50473 DVSS.n1291 DVSS.n1290 0.0272589
R50474 DVSS.n19848 DVSS.n19090 0.0272589
R50475 DVSS.n19108 DVSS.n19092 0.0272589
R50476 DVSS.n1273 DVSS.n1271 0.0272589
R50477 DVSS.n1217 DVSS.n1201 0.0272589
R50478 DVSS.n20433 DVSS.n20358 0.0272589
R50479 DVSS.n20353 DVSS.n20352 0.0272589
R50480 DVSS.n20353 DVSS.n14857 0.0272589
R50481 DVSS.n20433 DVSS.n20432 0.0272589
R50482 DVSS.n16464 DVSS.n16365 0.0271238
R50483 DVSS.n18087 DVSS.n15645 0.0271238
R50484 DVSS.n2722 DVSS.n2705 0.0270284
R50485 DVSS.n13357 DVSS.n1514 0.0270284
R50486 DVSS.n2724 DVSS.n2704 0.0270284
R50487 DVSS.n13356 DVSS.n1516 0.0270284
R50488 DVSS.n18978 DVSS.n14551 0.026913
R50489 DVSS.n18978 DVSS.n14566 0.026913
R50490 DVSS.n20147 DVSS.n14588 0.026913
R50491 DVSS.n20147 DVSS.n14599 0.026913
R50492 DVSS.n20280 DVSS.n14643 0.026913
R50493 DVSS.n20280 DVSS.n14638 0.026913
R50494 DVSS.n20398 DVSS.n20397 0.026913
R50495 DVSS.n20399 DVSS.n20398 0.026913
R50496 DVSS.n18925 DVSS.n14518 0.026913
R50497 DVSS.n18925 DVSS.n14533 0.026913
R50498 DVSS.n20073 DVSS.n20013 0.026913
R50499 DVSS.n20073 DVSS.n20024 0.026913
R50500 DVSS.n20251 DVSS.n20188 0.026913
R50501 DVSS.n20251 DVSS.n14870 0.026913
R50502 DVSS.n20389 DVSS.n20326 0.026913
R50503 DVSS.n20389 DVSS.n14861 0.026913
R50504 DVSS.n19316 DVSS.n19306 0.026913
R50505 DVSS.n19320 DVSS.n19306 0.026913
R50506 DVSS.n19321 DVSS.n19320 0.026913
R50507 DVSS.n19322 DVSS.n19321 0.026913
R50508 DVSS.n19322 DVSS.n19304 0.026913
R50509 DVSS.n19326 DVSS.n19304 0.026913
R50510 DVSS.n19327 DVSS.n19326 0.026913
R50511 DVSS.n19328 DVSS.n19327 0.026913
R50512 DVSS.n19328 DVSS.n19302 0.026913
R50513 DVSS.n19332 DVSS.n19302 0.026913
R50514 DVSS.n19333 DVSS.n19332 0.026913
R50515 DVSS.n19334 DVSS.n19333 0.026913
R50516 DVSS.n19334 DVSS.n19300 0.026913
R50517 DVSS.n19338 DVSS.n19300 0.026913
R50518 DVSS.n19339 DVSS.n19338 0.026913
R50519 DVSS.n19340 DVSS.n19339 0.026913
R50520 DVSS.n19340 DVSS.n19298 0.026913
R50521 DVSS.n19344 DVSS.n19298 0.026913
R50522 DVSS.n19345 DVSS.n19344 0.026913
R50523 DVSS.n19346 DVSS.n19345 0.026913
R50524 DVSS.n19346 DVSS.n19296 0.026913
R50525 DVSS.n19350 DVSS.n19296 0.026913
R50526 DVSS.n19351 DVSS.n19350 0.026913
R50527 DVSS.n19352 DVSS.n19351 0.026913
R50528 DVSS.n19352 DVSS.n19294 0.026913
R50529 DVSS.n19356 DVSS.n19294 0.026913
R50530 DVSS.n19357 DVSS.n19356 0.026913
R50531 DVSS.n19358 DVSS.n19357 0.026913
R50532 DVSS.n19358 DVSS.n19292 0.026913
R50533 DVSS.n19362 DVSS.n19292 0.026913
R50534 DVSS.n19363 DVSS.n19362 0.026913
R50535 DVSS.n19364 DVSS.n19363 0.026913
R50536 DVSS.n19364 DVSS.n19290 0.026913
R50537 DVSS.n19368 DVSS.n19290 0.026913
R50538 DVSS.n19369 DVSS.n19368 0.026913
R50539 DVSS.n19370 DVSS.n19369 0.026913
R50540 DVSS.n19370 DVSS.n19288 0.026913
R50541 DVSS.n19374 DVSS.n19288 0.026913
R50542 DVSS.n19375 DVSS.n19374 0.026913
R50543 DVSS.n19376 DVSS.n19375 0.026913
R50544 DVSS.n19376 DVSS.n19286 0.026913
R50545 DVSS.n19380 DVSS.n19286 0.026913
R50546 DVSS.n19381 DVSS.n19380 0.026913
R50547 DVSS.n19382 DVSS.n19381 0.026913
R50548 DVSS.n19382 DVSS.n19284 0.026913
R50549 DVSS.n19386 DVSS.n19284 0.026913
R50550 DVSS.n19387 DVSS.n19386 0.026913
R50551 DVSS.n19388 DVSS.n19387 0.026913
R50552 DVSS.n19388 DVSS.n19282 0.026913
R50553 DVSS.n19392 DVSS.n19282 0.026913
R50554 DVSS.n19393 DVSS.n19392 0.026913
R50555 DVSS.n19394 DVSS.n19393 0.026913
R50556 DVSS.n19394 DVSS.n19279 0.026913
R50557 DVSS.n19500 DVSS.n19280 0.026913
R50558 DVSS.n19496 DVSS.n19280 0.026913
R50559 DVSS.n19496 DVSS.n19495 0.026913
R50560 DVSS.n19495 DVSS.n19494 0.026913
R50561 DVSS.n19494 DVSS.n19398 0.026913
R50562 DVSS.n19490 DVSS.n19398 0.026913
R50563 DVSS.n19490 DVSS.n19489 0.026913
R50564 DVSS.n19489 DVSS.n19488 0.026913
R50565 DVSS.n19488 DVSS.n19400 0.026913
R50566 DVSS.n19484 DVSS.n19400 0.026913
R50567 DVSS.n19484 DVSS.n19483 0.026913
R50568 DVSS.n19483 DVSS.n19482 0.026913
R50569 DVSS.n19482 DVSS.n19402 0.026913
R50570 DVSS.n19478 DVSS.n19402 0.026913
R50571 DVSS.n19478 DVSS.n19477 0.026913
R50572 DVSS.n19477 DVSS.n19476 0.026913
R50573 DVSS.n19476 DVSS.n19404 0.026913
R50574 DVSS.n19472 DVSS.n19404 0.026913
R50575 DVSS.n19472 DVSS.n19471 0.026913
R50576 DVSS.n19471 DVSS.n19470 0.026913
R50577 DVSS.n19470 DVSS.n19406 0.026913
R50578 DVSS.n19466 DVSS.n19406 0.026913
R50579 DVSS.n19466 DVSS.n19465 0.026913
R50580 DVSS.n19465 DVSS.n19464 0.026913
R50581 DVSS.n19464 DVSS.n19408 0.026913
R50582 DVSS.n19460 DVSS.n19408 0.026913
R50583 DVSS.n19460 DVSS.n19459 0.026913
R50584 DVSS.n19459 DVSS.n19458 0.026913
R50585 DVSS.n19458 DVSS.n19410 0.026913
R50586 DVSS.n19454 DVSS.n19410 0.026913
R50587 DVSS.n19454 DVSS.n19453 0.026913
R50588 DVSS.n19453 DVSS.n19452 0.026913
R50589 DVSS.n19452 DVSS.n19412 0.026913
R50590 DVSS.n19448 DVSS.n19412 0.026913
R50591 DVSS.n19448 DVSS.n19447 0.026913
R50592 DVSS.n19447 DVSS.n19446 0.026913
R50593 DVSS.n19446 DVSS.n19414 0.026913
R50594 DVSS.n19442 DVSS.n19414 0.026913
R50595 DVSS.n19442 DVSS.n19441 0.026913
R50596 DVSS.n19441 DVSS.n19440 0.026913
R50597 DVSS.n19440 DVSS.n19416 0.026913
R50598 DVSS.n19436 DVSS.n19416 0.026913
R50599 DVSS.n19436 DVSS.n19435 0.026913
R50600 DVSS.n19435 DVSS.n19434 0.026913
R50601 DVSS.n19434 DVSS.n19418 0.026913
R50602 DVSS.n19430 DVSS.n19418 0.026913
R50603 DVSS.n19430 DVSS.n19429 0.026913
R50604 DVSS.n19429 DVSS.n19428 0.026913
R50605 DVSS.n19428 DVSS.n19425 0.026913
R50606 DVSS.n19425 DVSS.n19424 0.026913
R50607 DVSS.n19424 DVSS.n19423 0.026913
R50608 DVSS.n19423 DVSS.n19422 0.026913
R50609 DVSS.n19422 DVSS.n1353 0.026913
R50610 DVSS.n22230 DVSS.n1353 0.026913
R50611 DVSS.n22230 DVSS.n22228 0.026913
R50612 DVSS.n22228 DVSS.n22226 0.026913
R50613 DVSS.n22226 DVSS.n22224 0.026913
R50614 DVSS.n22224 DVSS.n22222 0.026913
R50615 DVSS.n22222 DVSS.n22220 0.026913
R50616 DVSS.n22220 DVSS.n22218 0.026913
R50617 DVSS.n22218 DVSS.n22215 0.026913
R50618 DVSS.n22215 DVSS.n22214 0.026913
R50619 DVSS.n22214 DVSS.n22212 0.026913
R50620 DVSS.n22212 DVSS.n1354 0.026913
R50621 DVSS.n22208 DVSS.n1354 0.026913
R50622 DVSS.n22208 DVSS.n22207 0.026913
R50623 DVSS.n22207 DVSS.n22206 0.026913
R50624 DVSS.n22206 DVSS.n1356 0.026913
R50625 DVSS.n22202 DVSS.n1356 0.026913
R50626 DVSS.n22202 DVSS.n22201 0.026913
R50627 DVSS.n22201 DVSS.n22200 0.026913
R50628 DVSS.n22200 DVSS.n1358 0.026913
R50629 DVSS.n22196 DVSS.n1358 0.026913
R50630 DVSS.n22196 DVSS.n22195 0.026913
R50631 DVSS.n22195 DVSS.n22194 0.026913
R50632 DVSS.n22194 DVSS.n1360 0.026913
R50633 DVSS.n22190 DVSS.n1360 0.026913
R50634 DVSS.n22190 DVSS.n22189 0.026913
R50635 DVSS.n22189 DVSS.n22188 0.026913
R50636 DVSS.n22188 DVSS.n1362 0.026913
R50637 DVSS.n22131 DVSS.n1362 0.026913
R50638 DVSS.n22132 DVSS.n22131 0.026913
R50639 DVSS.n22181 DVSS.n22132 0.026913
R50640 DVSS.n22181 DVSS.n22180 0.026913
R50641 DVSS.n22180 DVSS.n22178 0.026913
R50642 DVSS.n22178 DVSS.n22175 0.026913
R50643 DVSS.n22175 DVSS.n22174 0.026913
R50644 DVSS.n22174 DVSS.n22172 0.026913
R50645 DVSS.n22172 DVSS.n22170 0.026913
R50646 DVSS.n22170 DVSS.n22168 0.026913
R50647 DVSS.n22168 DVSS.n22166 0.026913
R50648 DVSS.n22166 DVSS.n22164 0.026913
R50649 DVSS.n22164 DVSS.n22162 0.026913
R50650 DVSS.n22162 DVSS.n22159 0.026913
R50651 DVSS.n22159 DVSS.n22158 0.026913
R50652 DVSS.n22158 DVSS.n22156 0.026913
R50653 DVSS.n22156 DVSS.n22154 0.026913
R50654 DVSS.n22154 DVSS.n22152 0.026913
R50655 DVSS.n22152 DVSS.n22150 0.026913
R50656 DVSS.n22150 DVSS.n22148 0.026913
R50657 DVSS.n22148 DVSS.n22146 0.026913
R50658 DVSS.n22146 DVSS.n22143 0.026913
R50659 DVSS.n22143 DVSS.n22142 0.026913
R50660 DVSS.n22142 DVSS.n22140 0.026913
R50661 DVSS.n22140 DVSS.n22138 0.026913
R50662 DVSS.n22138 DVSS.n22136 0.026913
R50663 DVSS.n22136 DVSS.n22134 0.026913
R50664 DVSS.n22134 DVSS.n879 0.026913
R50665 DVSS.n22455 DVSS.n880 0.026913
R50666 DVSS.n927 DVSS.n880 0.026913
R50667 DVSS.n929 DVSS.n927 0.026913
R50668 DVSS.n931 DVSS.n929 0.026913
R50669 DVSS.n933 DVSS.n931 0.026913
R50670 DVSS.n935 DVSS.n933 0.026913
R50671 DVSS.n937 DVSS.n935 0.026913
R50672 DVSS.n939 DVSS.n937 0.026913
R50673 DVSS.n940 DVSS.n939 0.026913
R50674 DVSS.n943 DVSS.n940 0.026913
R50675 DVSS.n945 DVSS.n943 0.026913
R50676 DVSS.n947 DVSS.n945 0.026913
R50677 DVSS.n949 DVSS.n947 0.026913
R50678 DVSS.n951 DVSS.n949 0.026913
R50679 DVSS.n953 DVSS.n951 0.026913
R50680 DVSS.n954 DVSS.n953 0.026913
R50681 DVSS.n957 DVSS.n954 0.026913
R50682 DVSS.n959 DVSS.n957 0.026913
R50683 DVSS.n961 DVSS.n959 0.026913
R50684 DVSS.n963 DVSS.n961 0.026913
R50685 DVSS.n965 DVSS.n963 0.026913
R50686 DVSS.n967 DVSS.n965 0.026913
R50687 DVSS.n968 DVSS.n967 0.026913
R50688 DVSS.n22449 DVSS.n968 0.026913
R50689 DVSS.n22449 DVSS.n22448 0.026913
R50690 DVSS.n22448 DVSS.n22447 0.026913
R50691 DVSS.n22447 DVSS.n22445 0.026913
R50692 DVSS.n22445 DVSS.n22443 0.026913
R50693 DVSS.n22443 DVSS.n969 0.026913
R50694 DVSS.n22439 DVSS.n969 0.026913
R50695 DVSS.n22439 DVSS.n22438 0.026913
R50696 DVSS.n22438 DVSS.n971 0.026913
R50697 DVSS.n22387 DVSS.n971 0.026913
R50698 DVSS.n22390 DVSS.n22387 0.026913
R50699 DVSS.n22392 DVSS.n22390 0.026913
R50700 DVSS.n22394 DVSS.n22392 0.026913
R50701 DVSS.n22396 DVSS.n22394 0.026913
R50702 DVSS.n22398 DVSS.n22396 0.026913
R50703 DVSS.n22400 DVSS.n22398 0.026913
R50704 DVSS.n22402 DVSS.n22400 0.026913
R50705 DVSS.n22403 DVSS.n22402 0.026913
R50706 DVSS.n22406 DVSS.n22403 0.026913
R50707 DVSS.n22408 DVSS.n22406 0.026913
R50708 DVSS.n22410 DVSS.n22408 0.026913
R50709 DVSS.n22412 DVSS.n22410 0.026913
R50710 DVSS.n22414 DVSS.n22412 0.026913
R50711 DVSS.n22416 DVSS.n22414 0.026913
R50712 DVSS.n22418 DVSS.n22416 0.026913
R50713 DVSS.n22419 DVSS.n22418 0.026913
R50714 DVSS.n22422 DVSS.n22419 0.026913
R50715 DVSS.n22424 DVSS.n22422 0.026913
R50716 DVSS.n22426 DVSS.n22424 0.026913
R50717 DVSS.n22428 DVSS.n22426 0.026913
R50718 DVSS.n19315 DVSS.n19314 0.026913
R50719 DVSS.n19898 DVSS.n19897 0.026913
R50720 DVSS.n19900 DVSS.n19021 0.026913
R50721 DVSS.n19247 DVSS.n19246 0.026913
R50722 DVSS.n19250 DVSS.n19169 0.026913
R50723 DVSS.n19621 DVSS.n19620 0.026913
R50724 DVSS.n19624 DVSS.n19156 0.026913
R50725 DVSS.n19649 DVSS.n19648 0.026913
R50726 DVSS.n19652 DVSS.n19141 0.026913
R50727 DVSS.n19657 DVSS.n19656 0.026913
R50728 DVSS.n19658 DVSS.n19137 0.026913
R50729 DVSS.n19662 DVSS.n19137 0.026913
R50730 DVSS.n19663 DVSS.n19662 0.026913
R50731 DVSS.n19664 DVSS.n19663 0.026913
R50732 DVSS.n19664 DVSS.n19135 0.026913
R50733 DVSS.n19668 DVSS.n19135 0.026913
R50734 DVSS.n19669 DVSS.n19668 0.026913
R50735 DVSS.n19670 DVSS.n19669 0.026913
R50736 DVSS.n19670 DVSS.n19133 0.026913
R50737 DVSS.n19674 DVSS.n19133 0.026913
R50738 DVSS.n19675 DVSS.n19674 0.026913
R50739 DVSS.n19676 DVSS.n19675 0.026913
R50740 DVSS.n19676 DVSS.n19131 0.026913
R50741 DVSS.n19680 DVSS.n19131 0.026913
R50742 DVSS.n19681 DVSS.n19680 0.026913
R50743 DVSS.n19682 DVSS.n19681 0.026913
R50744 DVSS.n19682 DVSS.n19129 0.026913
R50745 DVSS.n19686 DVSS.n19129 0.026913
R50746 DVSS.n19687 DVSS.n19686 0.026913
R50747 DVSS.n19688 DVSS.n19687 0.026913
R50748 DVSS.n19688 DVSS.n19127 0.026913
R50749 DVSS.n19692 DVSS.n19127 0.026913
R50750 DVSS.n19693 DVSS.n19692 0.026913
R50751 DVSS.n19694 DVSS.n19693 0.026913
R50752 DVSS.n19694 DVSS.n19125 0.026913
R50753 DVSS.n19698 DVSS.n19125 0.026913
R50754 DVSS.n19699 DVSS.n19698 0.026913
R50755 DVSS.n19700 DVSS.n19699 0.026913
R50756 DVSS.n19700 DVSS.n19123 0.026913
R50757 DVSS.n19704 DVSS.n19123 0.026913
R50758 DVSS.n19705 DVSS.n19704 0.026913
R50759 DVSS.n19706 DVSS.n19705 0.026913
R50760 DVSS.n19706 DVSS.n19121 0.026913
R50761 DVSS.n19710 DVSS.n19121 0.026913
R50762 DVSS.n19711 DVSS.n19710 0.026913
R50763 DVSS.n19712 DVSS.n19711 0.026913
R50764 DVSS.n19712 DVSS.n19119 0.026913
R50765 DVSS.n19716 DVSS.n19119 0.026913
R50766 DVSS.n19717 DVSS.n19716 0.026913
R50767 DVSS.n19718 DVSS.n19717 0.026913
R50768 DVSS.n19718 DVSS.n19117 0.026913
R50769 DVSS.n19722 DVSS.n19117 0.026913
R50770 DVSS.n19723 DVSS.n19722 0.026913
R50771 DVSS.n19724 DVSS.n19723 0.026913
R50772 DVSS.n19724 DVSS.n19115 0.026913
R50773 DVSS.n19728 DVSS.n19115 0.026913
R50774 DVSS.n19729 DVSS.n19728 0.026913
R50775 DVSS.n19730 DVSS.n19729 0.026913
R50776 DVSS.n19730 DVSS.n19113 0.026913
R50777 DVSS.n19734 DVSS.n19113 0.026913
R50778 DVSS.n19735 DVSS.n19734 0.026913
R50779 DVSS.n19736 DVSS.n19735 0.026913
R50780 DVSS.n19736 DVSS.n19110 0.026913
R50781 DVSS.n19844 DVSS.n19111 0.026913
R50782 DVSS.n19840 DVSS.n19111 0.026913
R50783 DVSS.n19840 DVSS.n19839 0.026913
R50784 DVSS.n19839 DVSS.n19838 0.026913
R50785 DVSS.n19838 DVSS.n19740 0.026913
R50786 DVSS.n19834 DVSS.n19740 0.026913
R50787 DVSS.n19834 DVSS.n19833 0.026913
R50788 DVSS.n19833 DVSS.n19832 0.026913
R50789 DVSS.n19832 DVSS.n19742 0.026913
R50790 DVSS.n19828 DVSS.n19742 0.026913
R50791 DVSS.n19828 DVSS.n19827 0.026913
R50792 DVSS.n19827 DVSS.n19826 0.026913
R50793 DVSS.n19826 DVSS.n19744 0.026913
R50794 DVSS.n19822 DVSS.n19744 0.026913
R50795 DVSS.n19822 DVSS.n19821 0.026913
R50796 DVSS.n19821 DVSS.n19820 0.026913
R50797 DVSS.n19820 DVSS.n19746 0.026913
R50798 DVSS.n19816 DVSS.n19746 0.026913
R50799 DVSS.n19816 DVSS.n19815 0.026913
R50800 DVSS.n19815 DVSS.n19814 0.026913
R50801 DVSS.n19814 DVSS.n19748 0.026913
R50802 DVSS.n19810 DVSS.n19748 0.026913
R50803 DVSS.n19810 DVSS.n19809 0.026913
R50804 DVSS.n19809 DVSS.n19808 0.026913
R50805 DVSS.n19808 DVSS.n19750 0.026913
R50806 DVSS.n19804 DVSS.n19750 0.026913
R50807 DVSS.n19804 DVSS.n19803 0.026913
R50808 DVSS.n19803 DVSS.n19802 0.026913
R50809 DVSS.n19802 DVSS.n19752 0.026913
R50810 DVSS.n19798 DVSS.n19752 0.026913
R50811 DVSS.n19798 DVSS.n19797 0.026913
R50812 DVSS.n19797 DVSS.n19796 0.026913
R50813 DVSS.n19796 DVSS.n19754 0.026913
R50814 DVSS.n19792 DVSS.n19754 0.026913
R50815 DVSS.n19792 DVSS.n19791 0.026913
R50816 DVSS.n19791 DVSS.n19790 0.026913
R50817 DVSS.n19790 DVSS.n19756 0.026913
R50818 DVSS.n19786 DVSS.n19756 0.026913
R50819 DVSS.n19786 DVSS.n19785 0.026913
R50820 DVSS.n19785 DVSS.n19784 0.026913
R50821 DVSS.n19784 DVSS.n19758 0.026913
R50822 DVSS.n19780 DVSS.n19758 0.026913
R50823 DVSS.n19780 DVSS.n19779 0.026913
R50824 DVSS.n19779 DVSS.n19778 0.026913
R50825 DVSS.n19778 DVSS.n19760 0.026913
R50826 DVSS.n19774 DVSS.n19760 0.026913
R50827 DVSS.n19774 DVSS.n19773 0.026913
R50828 DVSS.n19773 DVSS.n19772 0.026913
R50829 DVSS.n19772 DVSS.n19762 0.026913
R50830 DVSS.n19768 DVSS.n19762 0.026913
R50831 DVSS.n19768 DVSS.n19767 0.026913
R50832 DVSS.n19767 DVSS.n19765 0.026913
R50833 DVSS.n19765 DVSS.n1272 0.026913
R50834 DVSS.n22233 DVSS.n1272 0.026913
R50835 DVSS.n22235 DVSS.n22233 0.026913
R50836 DVSS.n22237 DVSS.n22235 0.026913
R50837 DVSS.n22239 DVSS.n22237 0.026913
R50838 DVSS.n22241 DVSS.n22239 0.026913
R50839 DVSS.n22243 DVSS.n22241 0.026913
R50840 DVSS.n22244 DVSS.n22243 0.026913
R50841 DVSS.n22247 DVSS.n22244 0.026913
R50842 DVSS.n22248 DVSS.n22247 0.026913
R50843 DVSS.n22249 DVSS.n22248 0.026913
R50844 DVSS.n22251 DVSS.n22249 0.026913
R50845 DVSS.n22252 DVSS.n22251 0.026913
R50846 DVSS.n22253 DVSS.n22252 0.026913
R50847 DVSS.n22253 DVSS.n1269 0.026913
R50848 DVSS.n22257 DVSS.n1269 0.026913
R50849 DVSS.n22258 DVSS.n22257 0.026913
R50850 DVSS.n22259 DVSS.n22258 0.026913
R50851 DVSS.n22259 DVSS.n1267 0.026913
R50852 DVSS.n22263 DVSS.n1267 0.026913
R50853 DVSS.n22264 DVSS.n22263 0.026913
R50854 DVSS.n22265 DVSS.n22264 0.026913
R50855 DVSS.n22265 DVSS.n1265 0.026913
R50856 DVSS.n22269 DVSS.n1265 0.026913
R50857 DVSS.n22270 DVSS.n22269 0.026913
R50858 DVSS.n22271 DVSS.n22270 0.026913
R50859 DVSS.n22271 DVSS.n1263 0.026913
R50860 DVSS.n22275 DVSS.n1263 0.026913
R50861 DVSS.n22277 DVSS.n22275 0.026913
R50862 DVSS.n22279 DVSS.n22277 0.026913
R50863 DVSS.n22281 DVSS.n22279 0.026913
R50864 DVSS.n22283 DVSS.n22281 0.026913
R50865 DVSS.n22284 DVSS.n22283 0.026913
R50866 DVSS.n22287 DVSS.n22284 0.026913
R50867 DVSS.n22289 DVSS.n22287 0.026913
R50868 DVSS.n22291 DVSS.n22289 0.026913
R50869 DVSS.n22293 DVSS.n22291 0.026913
R50870 DVSS.n22295 DVSS.n22293 0.026913
R50871 DVSS.n22297 DVSS.n22295 0.026913
R50872 DVSS.n22299 DVSS.n22297 0.026913
R50873 DVSS.n22300 DVSS.n22299 0.026913
R50874 DVSS.n22303 DVSS.n22300 0.026913
R50875 DVSS.n22305 DVSS.n22303 0.026913
R50876 DVSS.n22307 DVSS.n22305 0.026913
R50877 DVSS.n22309 DVSS.n22307 0.026913
R50878 DVSS.n22311 DVSS.n22309 0.026913
R50879 DVSS.n22313 DVSS.n22311 0.026913
R50880 DVSS.n22315 DVSS.n22313 0.026913
R50881 DVSS.n22316 DVSS.n22315 0.026913
R50882 DVSS.n22319 DVSS.n22316 0.026913
R50883 DVSS.n22321 DVSS.n22319 0.026913
R50884 DVSS.n22322 DVSS.n22321 0.026913
R50885 DVSS.n22322 DVSS.n1222 0.026913
R50886 DVSS.n22328 DVSS.n1222 0.026913
R50887 DVSS.n22329 DVSS.n22328 0.026913
R50888 DVSS.n22329 DVSS.n1219 0.026913
R50889 DVSS.n22333 DVSS.n1220 0.026913
R50890 DVSS.n12822 DVSS.n1220 0.026913
R50891 DVSS.n12824 DVSS.n12822 0.026913
R50892 DVSS.n12826 DVSS.n12824 0.026913
R50893 DVSS.n12828 DVSS.n12826 0.026913
R50894 DVSS.n12830 DVSS.n12828 0.026913
R50895 DVSS.n12832 DVSS.n12830 0.026913
R50896 DVSS.n12834 DVSS.n12832 0.026913
R50897 DVSS.n12835 DVSS.n12834 0.026913
R50898 DVSS.n12838 DVSS.n12835 0.026913
R50899 DVSS.n12840 DVSS.n12838 0.026913
R50900 DVSS.n12842 DVSS.n12840 0.026913
R50901 DVSS.n12844 DVSS.n12842 0.026913
R50902 DVSS.n12846 DVSS.n12844 0.026913
R50903 DVSS.n12848 DVSS.n12846 0.026913
R50904 DVSS.n12849 DVSS.n12848 0.026913
R50905 DVSS.n12852 DVSS.n12849 0.026913
R50906 DVSS.n12854 DVSS.n12852 0.026913
R50907 DVSS.n12856 DVSS.n12854 0.026913
R50908 DVSS.n12858 DVSS.n12856 0.026913
R50909 DVSS.n12860 DVSS.n12858 0.026913
R50910 DVSS.n12862 DVSS.n12860 0.026913
R50911 DVSS.n12864 DVSS.n12862 0.026913
R50912 DVSS.n12865 DVSS.n12864 0.026913
R50913 DVSS.n12868 DVSS.n12865 0.026913
R50914 DVSS.n12870 DVSS.n12868 0.026913
R50915 DVSS.n12871 DVSS.n12870 0.026913
R50916 DVSS.n12872 DVSS.n12871 0.026913
R50917 DVSS.n12873 DVSS.n12872 0.026913
R50918 DVSS.n12876 DVSS.n12873 0.026913
R50919 DVSS.n12878 DVSS.n12876 0.026913
R50920 DVSS.n12880 DVSS.n12878 0.026913
R50921 DVSS.n12881 DVSS.n12880 0.026913
R50922 DVSS.n12884 DVSS.n12881 0.026913
R50923 DVSS.n12886 DVSS.n12884 0.026913
R50924 DVSS.n12888 DVSS.n12886 0.026913
R50925 DVSS.n12890 DVSS.n12888 0.026913
R50926 DVSS.n12892 DVSS.n12890 0.026913
R50927 DVSS.n12894 DVSS.n12892 0.026913
R50928 DVSS.n12896 DVSS.n12894 0.026913
R50929 DVSS.n12897 DVSS.n12896 0.026913
R50930 DVSS.n12900 DVSS.n12897 0.026913
R50931 DVSS.n12902 DVSS.n12900 0.026913
R50932 DVSS.n12904 DVSS.n12902 0.026913
R50933 DVSS.n12906 DVSS.n12904 0.026913
R50934 DVSS.n12908 DVSS.n12906 0.026913
R50935 DVSS.n12910 DVSS.n12908 0.026913
R50936 DVSS.n12912 DVSS.n12910 0.026913
R50937 DVSS.n12913 DVSS.n12912 0.026913
R50938 DVSS.n12916 DVSS.n12913 0.026913
R50939 DVSS.n12918 DVSS.n12916 0.026913
R50940 DVSS.n12920 DVSS.n12918 0.026913
R50941 DVSS.n12922 DVSS.n12920 0.026913
R50942 DVSS.n12923 DVSS.n12922 0.026913
R50943 DVSS.n22384 DVSS.n1042 0.026913
R50944 DVSS.n22370 DVSS.n1174 0.026913
R50945 DVSS.n13089 DVSS.n12958 0.026913
R50946 DVSS.n4467 DVSS.n4460 0.0266354
R50947 DVSS.n4465 DVSS.n4461 0.0266354
R50948 DVSS.n17402 DVSS.n17386 0.0263511
R50949 DVSS.n17402 DVSS.n17387 0.0263511
R50950 DVSS.n17407 DVSS.n17271 0.0263511
R50951 DVSS.n17407 DVSS.n17272 0.0263511
R50952 DVSS.n17415 DVSS.n17236 0.0263511
R50953 DVSS.n17415 DVSS.n17237 0.0263511
R50954 DVSS.n17420 DVSS.n17419 0.0263511
R50955 DVSS.n17326 DVSS.n17319 0.0263511
R50956 DVSS.n17358 DVSS.n17344 0.0263511
R50957 DVSS.n17491 DVSS.n16951 0.0263511
R50958 DVSS.n17294 DVSS.n17135 0.0263511
R50959 DVSS.n17136 DVSS.n17135 0.0263511
R50960 DVSS.n17170 DVSS.n17169 0.0263511
R50961 DVSS.n17171 DVSS.n17170 0.0263511
R50962 DVSS.n17458 DVSS.n17196 0.0263511
R50963 DVSS.n17197 DVSS.n17196 0.0263511
R50964 DVSS.n17455 DVSS.n17444 0.0263511
R50965 DVSS.n7073 DVSS.n7072 0.025925
R50966 DVSS.n11986 DVSS.n11636 0.0259118
R50967 DVSS.n7053 DVSS.n7052 0.0259118
R50968 DVSS.n7073 DVSS.n5521 0.0259118
R50969 DVSS.n7096 DVSS.n7095 0.0259118
R50970 DVSS.n7456 DVSS.n4828 0.0259118
R50971 DVSS.n7811 DVSS.n4814 0.0259118
R50972 DVSS.n7831 DVSS.n4462 0.0259118
R50973 DVSS.n7843 DVSS.n4458 0.0259118
R50974 DVSS.n8107 DVSS.n4358 0.0259118
R50975 DVSS.n8325 DVSS.n3852 0.0259118
R50976 DVSS.n8582 DVSS.n3751 0.0259118
R50977 DVSS.n8595 DVSS.n3748 0.0259118
R50978 DVSS.n8620 DVSS.n3402 0.0259118
R50979 DVSS.n8974 DVSS.n3055 0.0259118
R50980 DVSS.n9192 DVSS.n2884 0.0259118
R50981 DVSS.n9449 DVSS.n2784 0.0259118
R50982 DVSS.n9512 DVSS.n2725 0.0259118
R50983 DVSS.n10111 DVSS.n10109 0.0259118
R50984 DVSS.n10135 DVSS.n10134 0.0259118
R50985 DVSS.n10160 DVSS.n10159 0.0259118
R50986 DVSS.n10469 DVSS.n10468 0.0259118
R50987 DVSS.n10491 DVSS.n1623 0.0259118
R50988 DVSS.n10759 DVSS.n1517 0.0259118
R50989 DVSS.n13354 DVSS.n10761 0.0259118
R50990 DVSS.n11452 DVSS.n11446 0.0259118
R50991 DVSS.n13320 DVSS.n11453 0.0259118
R50992 DVSS.n7029 DVSS.n7027 0.0259118
R50993 DVSS.n5985 DVSS.n5885 0.0259118
R50994 DVSS.n13115 DVSS.n11988 0.0259118
R50995 DVSS.n21175 DVSS.n13663 0.0258846
R50996 DVSS.n22607 DVSS.n743 0.0256163
R50997 DVSS.n22914 DVSS.n443 0.0256163
R50998 DVSS.n8974 DVSS.n8973 0.025475
R50999 DVSS.n13115 DVSS.n13114 0.025475
R51000 DVSS.n13104 DVSS.n12353 0.0251375
R51001 DVSS.n12362 DVSS.n12354 0.0251375
R51002 DVSS.n6665 DVSS.n6247 0.0251375
R51003 DVSS.n6308 DVSS.n6248 0.0251375
R51004 DVSS.n7840 DVSS.n7835 0.0250633
R51005 DVSS.n7834 DVSS.n4459 0.0250633
R51006 DVSS.n9774 DVSS.n2725 0.025025
R51007 DVSS.n11452 DVSS.n11451 0.025025
R51008 DVSS.n10128 DVSS.n2413 0.0246703
R51009 DVSS.n1522 DVSS.n1513 0.0246703
R51010 DVSS.n10130 DVSS.n10129 0.0246703
R51011 DVSS.n1520 DVSS.n1515 0.0246703
R51012 DVSS.n7812 DVSS.n7811 0.024575
R51013 DVSS.n3502 DVSS.n3405 0.0242773
R51014 DVSS.n8598 DVSS.n3404 0.0242773
R51015 DVSS.n16497 DVSS.n16495 0.0241441
R51016 DVSS.n16499 DVSS.n16497 0.0241441
R51017 DVSS.n16501 DVSS.n16499 0.0241441
R51018 DVSS.n16503 DVSS.n16501 0.0241441
R51019 DVSS.n16505 DVSS.n16503 0.0241441
R51020 DVSS.n16506 DVSS.n16505 0.0241441
R51021 DVSS.n16507 DVSS.n16506 0.0241441
R51022 DVSS.n16507 DVSS.n16490 0.0241441
R51023 DVSS.n16511 DVSS.n16490 0.0241441
R51024 DVSS.n16512 DVSS.n16511 0.0241441
R51025 DVSS.n16513 DVSS.n16512 0.0241441
R51026 DVSS.n16517 DVSS.n16516 0.0241441
R51027 DVSS.n16518 DVSS.n16486 0.0241441
R51028 DVSS.n16522 DVSS.n16486 0.0241441
R51029 DVSS.n16523 DVSS.n16522 0.0241441
R51030 DVSS.n16524 DVSS.n16523 0.0241441
R51031 DVSS.n16524 DVSS.n16484 0.0241441
R51032 DVSS.n16528 DVSS.n16484 0.0241441
R51033 DVSS.n16530 DVSS.n16528 0.0241441
R51034 DVSS.n16532 DVSS.n16530 0.0241441
R51035 DVSS.n16534 DVSS.n16532 0.0241441
R51036 DVSS.n16536 DVSS.n16534 0.0241441
R51037 DVSS.n16538 DVSS.n16536 0.0241441
R51038 DVSS.n16539 DVSS.n16538 0.0241441
R51039 DVSS.n18154 DVSS.n15546 0.0241441
R51040 DVSS.n15578 DVSS.n15546 0.0241441
R51041 DVSS.n15580 DVSS.n15578 0.0241441
R51042 DVSS.n15581 DVSS.n15580 0.0241441
R51043 DVSS.n18146 DVSS.n15581 0.0241441
R51044 DVSS.n18146 DVSS.n18145 0.0241441
R51045 DVSS.n18145 DVSS.n18144 0.0241441
R51046 DVSS.n18144 DVSS.n15582 0.0241441
R51047 DVSS.n18140 DVSS.n15582 0.0241441
R51048 DVSS.n18140 DVSS.n18139 0.0241441
R51049 DVSS.n18139 DVSS.n18138 0.0241441
R51050 DVSS.n18135 DVSS.n18134 0.0241441
R51051 DVSS.n18133 DVSS.n15586 0.0241441
R51052 DVSS.n18129 DVSS.n15586 0.0241441
R51053 DVSS.n18129 DVSS.n18128 0.0241441
R51054 DVSS.n18128 DVSS.n18127 0.0241441
R51055 DVSS.n18127 DVSS.n15588 0.0241441
R51056 DVSS.n18123 DVSS.n15588 0.0241441
R51057 DVSS.n18123 DVSS.n18122 0.0241441
R51058 DVSS.n18122 DVSS.n15590 0.0241441
R51059 DVSS.n18097 DVSS.n15590 0.0241441
R51060 DVSS.n18099 DVSS.n18097 0.0241441
R51061 DVSS.n18101 DVSS.n18099 0.0241441
R51062 DVSS.n18109 DVSS.n18101 0.0241441
R51063 DVSS.n18973 DVSS.n14565 0.0239783
R51064 DVSS.n18976 DVSS.n18975 0.0239783
R51065 DVSS.n20071 DVSS.n14598 0.0239783
R51066 DVSS.n20149 DVSS.n14587 0.0239783
R51067 DVSS.n20278 DVSS.n14639 0.0239783
R51068 DVSS.n20237 DVSS.n14644 0.0239783
R51069 DVSS.n20396 DVSS.n14669 0.0239783
R51070 DVSS.n20402 DVSS.n20401 0.0239783
R51071 DVSS.n18931 DVSS.n14532 0.0239783
R51072 DVSS.n18923 DVSS.n18922 0.0239783
R51073 DVSS.n20075 DVSS.n20023 0.0239783
R51074 DVSS.n20067 DVSS.n20012 0.0239783
R51075 DVSS.n20257 DVSS.n14871 0.0239783
R51076 DVSS.n20249 DVSS.n20189 0.0239783
R51077 DVSS.n20387 DVSS.n14862 0.0239783
R51078 DVSS.n20393 DVSS.n20327 0.0239783
R51079 DVSS.n5882 DVSS.n5866 0.0238843
R51080 DVSS.n5884 DVSS.n5865 0.0238843
R51081 DVSS.n16549 DVSS.n16478 0.0230723
R51082 DVSS.n18110 DVSS.n15622 0.0230723
R51083 DVSS.n13678 DVSS.n13677 0.0228256
R51084 DVSS.n21014 DVSS.n20998 0.0228256
R51085 DVSS.n17050 DVSS.n17049 0.0227859
R51086 DVSS.n17035 DVSS.n17034 0.0227859
R51087 DVSS.n17014 DVSS.n17013 0.0227859
R51088 DVSS.n16994 DVSS.n16993 0.0227859
R51089 DVSS.n17115 DVSS.n17114 0.0227859
R51090 DVSS.n17102 DVSS.n17101 0.0227859
R51091 DVSS.n17066 DVSS.n17057 0.0227859
R51092 DVSS.n17098 DVSS.n17076 0.0227859
R51093 DVSS.n17078 DVSS.n17077 0.0227859
R51094 DVSS.n17074 DVSS.n17065 0.0227859
R51095 DVSS.n17017 DVSS.n17016 0.0227859
R51096 DVSS.n17100 DVSS.n17057 0.0227859
R51097 DVSS.n17096 DVSS.n17095 0.0227859
R51098 DVSS.n16996 DVSS.n16995 0.0227859
R51099 DVSS.n17037 DVSS.n17036 0.0227859
R51100 DVSS.n16910 DVSS.n16909 0.0227859
R51101 DVSS.n16922 DVSS.n16920 0.0227859
R51102 DVSS.n16981 DVSS.n16980 0.0227859
R51103 DVSS DVSS.n16378 0.022775
R51104 DVSS.n18062 DVSS 0.022775
R51105 DVSS.n8107 DVSS.n8106 0.022775
R51106 DVSS.n7070 DVSS.n5185 0.0227052
R51107 DVSS.n7071 DVSS.n5186 0.0227052
R51108 DVSS.n16403 DVSS.n16402 0.02255
R51109 DVSS.n18057 DVSS.n15684 0.02255
R51110 DVSS.n10159 DVSS.n2360 0.022325
R51111 DVSS.n10492 DVSS.n10491 0.022325
R51112 DVSS.n8971 DVSS.n3053 0.0223122
R51113 DVSS.n13112 DVSS.n11992 0.0223122
R51114 DVSS.n8972 DVSS.n3054 0.0223122
R51115 DVSS.n13113 DVSS.n11990 0.0223122
R51116 DVSS.n19894 DVSS.n19041 0.0221878
R51117 DVSS.n19159 DVSS.n19044 0.0221878
R51118 DVSS.n19899 DVSS.n19896 0.0221878
R51119 DVSS.n19146 DVSS.n19145 0.0221878
R51120 DVSS.n19894 DVSS.n19893 0.0219244
R51121 DVSS.n19893 DVSS.n19042 0.0219244
R51122 DVSS.n19881 DVSS.n19042 0.0219244
R51123 DVSS.n19881 DVSS.n19880 0.0219244
R51124 DVSS.n19880 DVSS.n19049 0.0219244
R51125 DVSS.n19868 DVSS.n19049 0.0219244
R51126 DVSS.n19868 DVSS.n19867 0.0219244
R51127 DVSS.n19867 DVSS.n19057 0.0219244
R51128 DVSS.n19855 DVSS.n19057 0.0219244
R51129 DVSS.n19855 DVSS.n19854 0.0219244
R51130 DVSS.n19589 DVSS.n19268 0.0219244
R51131 DVSS.n19577 DVSS.n19268 0.0219244
R51132 DVSS.n19577 DVSS.n19576 0.0219244
R51133 DVSS.n19576 DVSS.n19523 0.0219244
R51134 DVSS.n19564 DVSS.n19523 0.0219244
R51135 DVSS.n19564 DVSS.n19563 0.0219244
R51136 DVSS.n19563 DVSS.n19531 0.0219244
R51137 DVSS.n19551 DVSS.n19531 0.0219244
R51138 DVSS.n19551 DVSS.n19550 0.0219244
R51139 DVSS.n19550 DVSS.n19539 0.0219244
R51140 DVSS.n21842 DVSS.n21827 0.0219244
R51141 DVSS.n21843 DVSS.n21842 0.0219244
R51142 DVSS.n21843 DVSS.n21603 0.0219244
R51143 DVSS.n19889 DVSS.n19044 0.0219244
R51144 DVSS.n19889 DVSS.n19888 0.0219244
R51145 DVSS.n19888 DVSS.n19045 0.0219244
R51146 DVSS.n19876 DVSS.n19045 0.0219244
R51147 DVSS.n19876 DVSS.n19875 0.0219244
R51148 DVSS.n19875 DVSS.n19053 0.0219244
R51149 DVSS.n19863 DVSS.n19053 0.0219244
R51150 DVSS.n19863 DVSS.n19862 0.0219244
R51151 DVSS.n19862 DVSS.n19061 0.0219244
R51152 DVSS.n19851 DVSS.n19061 0.0219244
R51153 DVSS.n19582 DVSS.n19520 0.0219244
R51154 DVSS.n19582 DVSS.n19581 0.0219244
R51155 DVSS.n19581 DVSS.n19521 0.0219244
R51156 DVSS.n19569 DVSS.n19521 0.0219244
R51157 DVSS.n19569 DVSS.n19568 0.0219244
R51158 DVSS.n19568 DVSS.n19529 0.0219244
R51159 DVSS.n19556 DVSS.n19529 0.0219244
R51160 DVSS.n19556 DVSS.n19555 0.0219244
R51161 DVSS.n19555 DVSS.n19537 0.0219244
R51162 DVSS.n19544 DVSS.n19537 0.0219244
R51163 DVSS.n21838 DVSS.n21834 0.0219244
R51164 DVSS.n21838 DVSS.n21837 0.0219244
R51165 DVSS.n21837 DVSS.n21706 0.0219244
R51166 DVSS.n19896 DVSS.n19040 0.0219244
R51167 DVSS.n19884 DVSS.n19040 0.0219244
R51168 DVSS.n19884 DVSS.n19883 0.0219244
R51169 DVSS.n19883 DVSS.n19047 0.0219244
R51170 DVSS.n19871 DVSS.n19047 0.0219244
R51171 DVSS.n19871 DVSS.n19870 0.0219244
R51172 DVSS.n19870 DVSS.n19055 0.0219244
R51173 DVSS.n19858 DVSS.n19055 0.0219244
R51174 DVSS.n19858 DVSS.n19857 0.0219244
R51175 DVSS.n19857 DVSS.n19063 0.0219244
R51176 DVSS.n19587 DVSS.n19586 0.0219244
R51177 DVSS.n19586 DVSS.n19516 0.0219244
R51178 DVSS.n19574 DVSS.n19516 0.0219244
R51179 DVSS.n19574 DVSS.n19573 0.0219244
R51180 DVSS.n19573 DVSS.n19525 0.0219244
R51181 DVSS.n19561 DVSS.n19525 0.0219244
R51182 DVSS.n19561 DVSS.n19560 0.0219244
R51183 DVSS.n19560 DVSS.n19533 0.0219244
R51184 DVSS.n19548 DVSS.n19533 0.0219244
R51185 DVSS.n19548 DVSS.n19547 0.0219244
R51186 DVSS.n21830 DVSS.n21825 0.0219244
R51187 DVSS.n21845 DVSS.n21825 0.0219244
R51188 DVSS.n21849 DVSS.n21845 0.0219244
R51189 DVSS.n19145 DVSS.n19043 0.0219244
R51190 DVSS.n19046 DVSS.n19043 0.0219244
R51191 DVSS.n19051 DVSS.n19046 0.0219244
R51192 DVSS.n19052 DVSS.n19051 0.0219244
R51193 DVSS.n19054 DVSS.n19052 0.0219244
R51194 DVSS.n19059 DVSS.n19054 0.0219244
R51195 DVSS.n19060 DVSS.n19059 0.0219244
R51196 DVSS.n19062 DVSS.n19060 0.0219244
R51197 DVSS.n19067 DVSS.n19062 0.0219244
R51198 DVSS.n19068 DVSS.n19067 0.0219244
R51199 DVSS.n19518 DVSS.n19517 0.0219244
R51200 DVSS.n19522 DVSS.n19517 0.0219244
R51201 DVSS.n19527 DVSS.n19522 0.0219244
R51202 DVSS.n19528 DVSS.n19527 0.0219244
R51203 DVSS.n19530 DVSS.n19528 0.0219244
R51204 DVSS.n19535 DVSS.n19530 0.0219244
R51205 DVSS.n19536 DVSS.n19535 0.0219244
R51206 DVSS.n19538 DVSS.n19536 0.0219244
R51207 DVSS.n19542 DVSS.n19538 0.0219244
R51208 DVSS.n19543 DVSS.n19542 0.0219244
R51209 DVSS.n21829 DVSS.n21828 0.0219244
R51210 DVSS.n21835 DVSS.n21828 0.0219244
R51211 DVSS.n21835 DVSS.n21799 0.0219244
R51212 DVSS.n9772 DVSS.n2727 0.0219192
R51213 DVSS.n11447 DVSS.n11199 0.0219192
R51214 DVSS.n9773 DVSS.n2726 0.0219192
R51215 DVSS.n13334 DVSS.n11448 0.0219192
R51216 DVSS.n8593 DVSS.n3751 0.021875
R51217 DVSS.n21176 DVSS.n21175 0.02156
R51218 DVSS.n21173 DVSS.n21172 0.02156
R51219 DVSS.n7814 DVSS.n4812 0.0215262
R51220 DVSS.n7813 DVSS.n4813 0.0215262
R51221 DVSS.n6692 DVSS.n5885 0.021425
R51222 DVSS.n18929 DVSS.n14552 0.0210435
R51223 DVSS.n20687 DVSS.n14567 0.0210435
R51224 DVSS.n20069 DVSS.n14589 0.0210435
R51225 DVSS.n20032 DVSS.n14600 0.0210435
R51226 DVSS.n20255 DVSS.n14642 0.0210435
R51227 DVSS.n20239 DVSS.n14637 0.0210435
R51228 DVSS.n20632 DVSS.n20631 0.0210435
R51229 DVSS.n20400 DVSS.n20376 0.0210435
R51230 DVSS.n18933 DVSS.n14519 0.0210435
R51231 DVSS.n20698 DVSS.n14534 0.0210435
R51232 DVSS.n20080 DVSS.n20014 0.0210435
R51233 DVSS.n20065 DVSS.n20025 0.0210435
R51234 DVSS.n20259 DVSS.n20187 0.0210435
R51235 DVSS.n20243 DVSS.n14869 0.0210435
R51236 DVSS.n20325 DVSS.n20324 0.0210435
R51237 DVSS.n20391 DVSS.n14860 0.0210435
R51238 DVSS.n21177 DVSS.n21176 0.0209
R51239 DVSS.n17488 DVSS.n17487 0.0202719
R51240 DVSS.n17487 DVSS.t190 0.0202719
R51241 DVSS.n17412 DVSS.n17411 0.0202719
R51242 DVSS.n17411 DVSS.t190 0.0202719
R51243 DVSS.n17473 DVSS.n17472 0.0202719
R51244 DVSS.n17472 DVSS.t190 0.0202719
R51245 DVSS.n7095 DVSS.n5173 0.020075
R51246 DVSS.n8104 DVSS.n4023 0.0199541
R51247 DVSS.n8105 DVSS.n4024 0.0199541
R51248 DVSS.n19854 DVSS.n19065 0.0199049
R51249 DVSS.n19592 DVSS.n19589 0.0199049
R51250 DVSS.n19851 DVSS.n19850 0.0199049
R51251 DVSS.n19520 DVSS.n19089 0.0199049
R51252 DVSS.n19512 DVSS.n19063 0.0199049
R51253 DVSS.n19587 DVSS.n19515 0.0199049
R51254 DVSS.n19847 DVSS.n19068 0.0199049
R51255 DVSS.n19518 DVSS.n19109 0.0199049
R51256 DVSS DVSS.n16192 0.0198891
R51257 DVSS.n16452 DVSS 0.0198891
R51258 DVSS.n5619 DVSS.n5618 0.019716
R51259 DVSS.n5626 DVSS.n5572 0.019716
R51260 DVSS.n5627 DVSS.n5626 0.019716
R51261 DVSS.n5632 DVSS.n5571 0.019716
R51262 DVSS.n5632 DVSS.n5631 0.019716
R51263 DVSS.n5638 DVSS.n5570 0.019716
R51264 DVSS.n5639 DVSS.n5638 0.019716
R51265 DVSS.n5644 DVSS.n5569 0.019716
R51266 DVSS.n5644 DVSS.n5643 0.019716
R51267 DVSS.n5650 DVSS.n5568 0.019716
R51268 DVSS.n5651 DVSS.n5650 0.019716
R51269 DVSS.n5656 DVSS.n5567 0.019716
R51270 DVSS.n5656 DVSS.n5655 0.019716
R51271 DVSS.n5662 DVSS.n5566 0.019716
R51272 DVSS.n5663 DVSS.n5662 0.019716
R51273 DVSS.n5668 DVSS.n5565 0.019716
R51274 DVSS.n5668 DVSS.n5667 0.019716
R51275 DVSS.n5674 DVSS.n5564 0.019716
R51276 DVSS.n5675 DVSS.n5674 0.019716
R51277 DVSS.n5680 DVSS.n5563 0.019716
R51278 DVSS.n5680 DVSS.n5679 0.019716
R51279 DVSS.n5686 DVSS.n5562 0.019716
R51280 DVSS.n5687 DVSS.n5686 0.019716
R51281 DVSS.n5692 DVSS.n5561 0.019716
R51282 DVSS.n5692 DVSS.n5691 0.019716
R51283 DVSS.n5698 DVSS.n5560 0.019716
R51284 DVSS.n5699 DVSS.n5698 0.019716
R51285 DVSS.n5704 DVSS.n5559 0.019716
R51286 DVSS.n5704 DVSS.n5703 0.019716
R51287 DVSS.n5710 DVSS.n5558 0.019716
R51288 DVSS.n5711 DVSS.n5710 0.019716
R51289 DVSS.n5716 DVSS.n5557 0.019716
R51290 DVSS.n5716 DVSS.n5715 0.019716
R51291 DVSS.n5722 DVSS.n5556 0.019716
R51292 DVSS.n5723 DVSS.n5722 0.019716
R51293 DVSS.n5728 DVSS.n5555 0.019716
R51294 DVSS.n5728 DVSS.n5727 0.019716
R51295 DVSS.n5734 DVSS.n5554 0.019716
R51296 DVSS.n5735 DVSS.n5734 0.019716
R51297 DVSS.n5740 DVSS.n5553 0.019716
R51298 DVSS.n5740 DVSS.n5739 0.019716
R51299 DVSS.n5746 DVSS.n5552 0.019716
R51300 DVSS.n5747 DVSS.n5746 0.019716
R51301 DVSS.n5752 DVSS.n5551 0.019716
R51302 DVSS.n5752 DVSS.n5751 0.019716
R51303 DVSS.n5758 DVSS.n5550 0.019716
R51304 DVSS.n5759 DVSS.n5758 0.019716
R51305 DVSS.n5764 DVSS.n5549 0.019716
R51306 DVSS.n5764 DVSS.n5763 0.019716
R51307 DVSS.n5770 DVSS.n5548 0.019716
R51308 DVSS.n5771 DVSS.n5770 0.019716
R51309 DVSS.n5776 DVSS.n5547 0.019716
R51310 DVSS.n5776 DVSS.n5775 0.019716
R51311 DVSS.n5782 DVSS.n5546 0.019716
R51312 DVSS.n5783 DVSS.n5782 0.019716
R51313 DVSS.n5788 DVSS.n5545 0.019716
R51314 DVSS.n5788 DVSS.n5787 0.019716
R51315 DVSS.n5794 DVSS.n5544 0.019716
R51316 DVSS.n5795 DVSS.n5794 0.019716
R51317 DVSS.n5800 DVSS.n5543 0.019716
R51318 DVSS.n5800 DVSS.n5799 0.019716
R51319 DVSS.n5806 DVSS.n5542 0.019716
R51320 DVSS.n5807 DVSS.n5806 0.019716
R51321 DVSS.n5812 DVSS.n5541 0.019716
R51322 DVSS.n5812 DVSS.n5811 0.019716
R51323 DVSS.n5818 DVSS.n5540 0.019716
R51324 DVSS.n5819 DVSS.n5818 0.019716
R51325 DVSS.n5824 DVSS.n5539 0.019716
R51326 DVSS.n5824 DVSS.n5823 0.019716
R51327 DVSS.n5830 DVSS.n5538 0.019716
R51328 DVSS.n5831 DVSS.n5830 0.019716
R51329 DVSS.n5836 DVSS.n5537 0.019716
R51330 DVSS.n5836 DVSS.n5835 0.019716
R51331 DVSS.n5842 DVSS.n5536 0.019716
R51332 DVSS.n5843 DVSS.n5842 0.019716
R51333 DVSS.n5848 DVSS.n5535 0.019716
R51334 DVSS.n5848 DVSS.n5847 0.019716
R51335 DVSS.n5854 DVSS.n5534 0.019716
R51336 DVSS.n5855 DVSS.n5854 0.019716
R51337 DVSS.n5860 DVSS.n5533 0.019716
R51338 DVSS.n5860 DVSS.n5859 0.019716
R51339 DVSS.n7056 DVSS.n5532 0.019716
R51340 DVSS.n7057 DVSS.n7056 0.019716
R51341 DVSS.n5274 DVSS.n5273 0.019716
R51342 DVSS.n5278 DVSS.n5275 0.019716
R51343 DVSS.n5278 DVSS.n5277 0.019716
R51344 DVSS.n5284 DVSS.n5266 0.019716
R51345 DVSS.n5285 DVSS.n5284 0.019716
R51346 DVSS.n5290 DVSS.n5287 0.019716
R51347 DVSS.n5290 DVSS.n5289 0.019716
R51348 DVSS.n5296 DVSS.n5262 0.019716
R51349 DVSS.n5297 DVSS.n5296 0.019716
R51350 DVSS.n5302 DVSS.n5299 0.019716
R51351 DVSS.n5302 DVSS.n5301 0.019716
R51352 DVSS.n5308 DVSS.n5258 0.019716
R51353 DVSS.n5309 DVSS.n5308 0.019716
R51354 DVSS.n5314 DVSS.n5311 0.019716
R51355 DVSS.n5314 DVSS.n5313 0.019716
R51356 DVSS.n5320 DVSS.n5254 0.019716
R51357 DVSS.n5321 DVSS.n5320 0.019716
R51358 DVSS.n5326 DVSS.n5323 0.019716
R51359 DVSS.n5326 DVSS.n5325 0.019716
R51360 DVSS.n5332 DVSS.n5250 0.019716
R51361 DVSS.n5333 DVSS.n5332 0.019716
R51362 DVSS.n5338 DVSS.n5335 0.019716
R51363 DVSS.n5338 DVSS.n5337 0.019716
R51364 DVSS.n5344 DVSS.n5246 0.019716
R51365 DVSS.n5345 DVSS.n5344 0.019716
R51366 DVSS.n5350 DVSS.n5347 0.019716
R51367 DVSS.n5350 DVSS.n5349 0.019716
R51368 DVSS.n5356 DVSS.n5242 0.019716
R51369 DVSS.n5357 DVSS.n5356 0.019716
R51370 DVSS.n5362 DVSS.n5359 0.019716
R51371 DVSS.n5362 DVSS.n5361 0.019716
R51372 DVSS.n5368 DVSS.n5238 0.019716
R51373 DVSS.n5369 DVSS.n5368 0.019716
R51374 DVSS.n5374 DVSS.n5371 0.019716
R51375 DVSS.n5374 DVSS.n5373 0.019716
R51376 DVSS.n5380 DVSS.n5234 0.019716
R51377 DVSS.n5381 DVSS.n5380 0.019716
R51378 DVSS.n5386 DVSS.n5383 0.019716
R51379 DVSS.n5386 DVSS.n5385 0.019716
R51380 DVSS.n5392 DVSS.n5230 0.019716
R51381 DVSS.n5393 DVSS.n5392 0.019716
R51382 DVSS.n5398 DVSS.n5395 0.019716
R51383 DVSS.n5398 DVSS.n5397 0.019716
R51384 DVSS.n5404 DVSS.n5226 0.019716
R51385 DVSS.n5405 DVSS.n5404 0.019716
R51386 DVSS.n5410 DVSS.n5407 0.019716
R51387 DVSS.n5410 DVSS.n5409 0.019716
R51388 DVSS.n5416 DVSS.n5222 0.019716
R51389 DVSS.n5417 DVSS.n5416 0.019716
R51390 DVSS.n5422 DVSS.n5419 0.019716
R51391 DVSS.n5422 DVSS.n5421 0.019716
R51392 DVSS.n5428 DVSS.n5218 0.019716
R51393 DVSS.n5429 DVSS.n5428 0.019716
R51394 DVSS.n5434 DVSS.n5431 0.019716
R51395 DVSS.n5434 DVSS.n5433 0.019716
R51396 DVSS.n5440 DVSS.n5214 0.019716
R51397 DVSS.n5441 DVSS.n5440 0.019716
R51398 DVSS.n5446 DVSS.n5443 0.019716
R51399 DVSS.n5446 DVSS.n5445 0.019716
R51400 DVSS.n5452 DVSS.n5210 0.019716
R51401 DVSS.n5453 DVSS.n5452 0.019716
R51402 DVSS.n5458 DVSS.n5455 0.019716
R51403 DVSS.n5458 DVSS.n5457 0.019716
R51404 DVSS.n5464 DVSS.n5206 0.019716
R51405 DVSS.n5465 DVSS.n5464 0.019716
R51406 DVSS.n5470 DVSS.n5467 0.019716
R51407 DVSS.n5470 DVSS.n5469 0.019716
R51408 DVSS.n5476 DVSS.n5202 0.019716
R51409 DVSS.n5477 DVSS.n5476 0.019716
R51410 DVSS.n5482 DVSS.n5479 0.019716
R51411 DVSS.n5482 DVSS.n5481 0.019716
R51412 DVSS.n5488 DVSS.n5198 0.019716
R51413 DVSS.n5489 DVSS.n5488 0.019716
R51414 DVSS.n5494 DVSS.n5491 0.019716
R51415 DVSS.n5494 DVSS.n5493 0.019716
R51416 DVSS.n5500 DVSS.n5194 0.019716
R51417 DVSS.n5501 DVSS.n5500 0.019716
R51418 DVSS.n5506 DVSS.n5503 0.019716
R51419 DVSS.n5506 DVSS.n5505 0.019716
R51420 DVSS.n5513 DVSS.n5190 0.019716
R51421 DVSS.n5514 DVSS.n5513 0.019716
R51422 DVSS.n5517 DVSS.n5516 0.019716
R51423 DVSS.n5518 DVSS.n5517 0.019716
R51424 DVSS.n4928 DVSS.n4927 0.019716
R51425 DVSS.n4935 DVSS.n4881 0.019716
R51426 DVSS.n4936 DVSS.n4935 0.019716
R51427 DVSS.n4941 DVSS.n4880 0.019716
R51428 DVSS.n4941 DVSS.n4940 0.019716
R51429 DVSS.n4947 DVSS.n4879 0.019716
R51430 DVSS.n4948 DVSS.n4947 0.019716
R51431 DVSS.n4953 DVSS.n4878 0.019716
R51432 DVSS.n4953 DVSS.n4952 0.019716
R51433 DVSS.n4959 DVSS.n4877 0.019716
R51434 DVSS.n4960 DVSS.n4959 0.019716
R51435 DVSS.n4965 DVSS.n4876 0.019716
R51436 DVSS.n4965 DVSS.n4964 0.019716
R51437 DVSS.n4971 DVSS.n4875 0.019716
R51438 DVSS.n4972 DVSS.n4971 0.019716
R51439 DVSS.n4977 DVSS.n4874 0.019716
R51440 DVSS.n4977 DVSS.n4976 0.019716
R51441 DVSS.n4983 DVSS.n4873 0.019716
R51442 DVSS.n4984 DVSS.n4983 0.019716
R51443 DVSS.n4989 DVSS.n4872 0.019716
R51444 DVSS.n4989 DVSS.n4988 0.019716
R51445 DVSS.n4995 DVSS.n4871 0.019716
R51446 DVSS.n4996 DVSS.n4995 0.019716
R51447 DVSS.n5001 DVSS.n4870 0.019716
R51448 DVSS.n5001 DVSS.n5000 0.019716
R51449 DVSS.n5007 DVSS.n4869 0.019716
R51450 DVSS.n5008 DVSS.n5007 0.019716
R51451 DVSS.n5013 DVSS.n4868 0.019716
R51452 DVSS.n5013 DVSS.n5012 0.019716
R51453 DVSS.n5019 DVSS.n4867 0.019716
R51454 DVSS.n5020 DVSS.n5019 0.019716
R51455 DVSS.n5025 DVSS.n4866 0.019716
R51456 DVSS.n5025 DVSS.n5024 0.019716
R51457 DVSS.n5031 DVSS.n4865 0.019716
R51458 DVSS.n5032 DVSS.n5031 0.019716
R51459 DVSS.n5037 DVSS.n4864 0.019716
R51460 DVSS.n5037 DVSS.n5036 0.019716
R51461 DVSS.n5043 DVSS.n4863 0.019716
R51462 DVSS.n5044 DVSS.n5043 0.019716
R51463 DVSS.n5049 DVSS.n4862 0.019716
R51464 DVSS.n5049 DVSS.n5048 0.019716
R51465 DVSS.n5055 DVSS.n4861 0.019716
R51466 DVSS.n5056 DVSS.n5055 0.019716
R51467 DVSS.n5061 DVSS.n4860 0.019716
R51468 DVSS.n5061 DVSS.n5060 0.019716
R51469 DVSS.n5067 DVSS.n4859 0.019716
R51470 DVSS.n5068 DVSS.n5067 0.019716
R51471 DVSS.n5073 DVSS.n4858 0.019716
R51472 DVSS.n5073 DVSS.n5072 0.019716
R51473 DVSS.n5079 DVSS.n4857 0.019716
R51474 DVSS.n5080 DVSS.n5079 0.019716
R51475 DVSS.n5085 DVSS.n4856 0.019716
R51476 DVSS.n5085 DVSS.n5084 0.019716
R51477 DVSS.n5091 DVSS.n4855 0.019716
R51478 DVSS.n5092 DVSS.n5091 0.019716
R51479 DVSS.n5097 DVSS.n4854 0.019716
R51480 DVSS.n5097 DVSS.n5096 0.019716
R51481 DVSS.n5103 DVSS.n4853 0.019716
R51482 DVSS.n5104 DVSS.n5103 0.019716
R51483 DVSS.n5109 DVSS.n4852 0.019716
R51484 DVSS.n5109 DVSS.n5108 0.019716
R51485 DVSS.n5115 DVSS.n4851 0.019716
R51486 DVSS.n5116 DVSS.n5115 0.019716
R51487 DVSS.n5121 DVSS.n4850 0.019716
R51488 DVSS.n5121 DVSS.n5120 0.019716
R51489 DVSS.n5127 DVSS.n4849 0.019716
R51490 DVSS.n5128 DVSS.n5127 0.019716
R51491 DVSS.n5133 DVSS.n4848 0.019716
R51492 DVSS.n5133 DVSS.n5132 0.019716
R51493 DVSS.n5139 DVSS.n4847 0.019716
R51494 DVSS.n5140 DVSS.n5139 0.019716
R51495 DVSS.n5145 DVSS.n4846 0.019716
R51496 DVSS.n5145 DVSS.n5144 0.019716
R51497 DVSS.n5151 DVSS.n4845 0.019716
R51498 DVSS.n5152 DVSS.n5151 0.019716
R51499 DVSS.n5157 DVSS.n4844 0.019716
R51500 DVSS.n5157 DVSS.n5156 0.019716
R51501 DVSS.n5163 DVSS.n4843 0.019716
R51502 DVSS.n5164 DVSS.n5163 0.019716
R51503 DVSS.n5169 DVSS.n4842 0.019716
R51504 DVSS.n5169 DVSS.n5168 0.019716
R51505 DVSS.n7099 DVSS.n4841 0.019716
R51506 DVSS.n7100 DVSS.n7099 0.019716
R51507 DVSS.n7441 DVSS.n7440 0.019716
R51508 DVSS.n7439 DVSS.n7438 0.019716
R51509 DVSS.n7438 DVSS.n7113 0.019716
R51510 DVSS.n7432 DVSS.n7118 0.019716
R51511 DVSS.n7432 DVSS.n7431 0.019716
R51512 DVSS.n7429 DVSS.n7428 0.019716
R51513 DVSS.n7428 DVSS.n7119 0.019716
R51514 DVSS.n7422 DVSS.n7124 0.019716
R51515 DVSS.n7422 DVSS.n7421 0.019716
R51516 DVSS.n7419 DVSS.n7418 0.019716
R51517 DVSS.n7418 DVSS.n7125 0.019716
R51518 DVSS.n7412 DVSS.n7130 0.019716
R51519 DVSS.n7412 DVSS.n7411 0.019716
R51520 DVSS.n7409 DVSS.n7408 0.019716
R51521 DVSS.n7408 DVSS.n7131 0.019716
R51522 DVSS.n7402 DVSS.n7136 0.019716
R51523 DVSS.n7402 DVSS.n7401 0.019716
R51524 DVSS.n7399 DVSS.n7398 0.019716
R51525 DVSS.n7398 DVSS.n7137 0.019716
R51526 DVSS.n7392 DVSS.n7142 0.019716
R51527 DVSS.n7392 DVSS.n7391 0.019716
R51528 DVSS.n7389 DVSS.n7388 0.019716
R51529 DVSS.n7388 DVSS.n7143 0.019716
R51530 DVSS.n7382 DVSS.n7148 0.019716
R51531 DVSS.n7382 DVSS.n7381 0.019716
R51532 DVSS.n7379 DVSS.n7378 0.019716
R51533 DVSS.n7378 DVSS.n7149 0.019716
R51534 DVSS.n7372 DVSS.n7154 0.019716
R51535 DVSS.n7372 DVSS.n7371 0.019716
R51536 DVSS.n7369 DVSS.n7368 0.019716
R51537 DVSS.n7368 DVSS.n7155 0.019716
R51538 DVSS.n7362 DVSS.n7160 0.019716
R51539 DVSS.n7362 DVSS.n7361 0.019716
R51540 DVSS.n7359 DVSS.n7358 0.019716
R51541 DVSS.n7358 DVSS.n7161 0.019716
R51542 DVSS.n7352 DVSS.n7166 0.019716
R51543 DVSS.n7352 DVSS.n7351 0.019716
R51544 DVSS.n7349 DVSS.n7348 0.019716
R51545 DVSS.n7348 DVSS.n7167 0.019716
R51546 DVSS.n7342 DVSS.n7172 0.019716
R51547 DVSS.n7342 DVSS.n7341 0.019716
R51548 DVSS.n7339 DVSS.n7338 0.019716
R51549 DVSS.n7338 DVSS.n7173 0.019716
R51550 DVSS.n7332 DVSS.n7178 0.019716
R51551 DVSS.n7332 DVSS.n7331 0.019716
R51552 DVSS.n7329 DVSS.n7328 0.019716
R51553 DVSS.n7328 DVSS.n7179 0.019716
R51554 DVSS.n7322 DVSS.n7184 0.019716
R51555 DVSS.n7322 DVSS.n7321 0.019716
R51556 DVSS.n7319 DVSS.n7318 0.019716
R51557 DVSS.n7318 DVSS.n7185 0.019716
R51558 DVSS.n7312 DVSS.n7190 0.019716
R51559 DVSS.n7312 DVSS.n7311 0.019716
R51560 DVSS.n7309 DVSS.n7308 0.019716
R51561 DVSS.n7308 DVSS.n7191 0.019716
R51562 DVSS.n7302 DVSS.n7196 0.019716
R51563 DVSS.n7302 DVSS.n7301 0.019716
R51564 DVSS.n7299 DVSS.n7298 0.019716
R51565 DVSS.n7298 DVSS.n7197 0.019716
R51566 DVSS.n7292 DVSS.n7202 0.019716
R51567 DVSS.n7292 DVSS.n7291 0.019716
R51568 DVSS.n7289 DVSS.n7288 0.019716
R51569 DVSS.n7288 DVSS.n7203 0.019716
R51570 DVSS.n7282 DVSS.n7208 0.019716
R51571 DVSS.n7282 DVSS.n7281 0.019716
R51572 DVSS.n7279 DVSS.n7278 0.019716
R51573 DVSS.n7278 DVSS.n7209 0.019716
R51574 DVSS.n7272 DVSS.n7214 0.019716
R51575 DVSS.n7272 DVSS.n7271 0.019716
R51576 DVSS.n7269 DVSS.n7268 0.019716
R51577 DVSS.n7268 DVSS.n7215 0.019716
R51578 DVSS.n7262 DVSS.n7220 0.019716
R51579 DVSS.n7262 DVSS.n7261 0.019716
R51580 DVSS.n7259 DVSS.n7258 0.019716
R51581 DVSS.n7258 DVSS.n7221 0.019716
R51582 DVSS.n7252 DVSS.n7226 0.019716
R51583 DVSS.n7252 DVSS.n7251 0.019716
R51584 DVSS.n7249 DVSS.n7248 0.019716
R51585 DVSS.n7248 DVSS.n7227 0.019716
R51586 DVSS.n7242 DVSS.n7232 0.019716
R51587 DVSS.n7242 DVSS.n7241 0.019716
R51588 DVSS.n7239 DVSS.n7238 0.019716
R51589 DVSS.n7238 DVSS.n7233 0.019716
R51590 DVSS.n7794 DVSS.n7503 0.019716
R51591 DVSS.n7505 DVSS.n7504 0.019716
R51592 DVSS.n7505 DVSS.n7502 0.019716
R51593 DVSS.n7785 DVSS.n7784 0.019716
R51594 DVSS.n7784 DVSS.n7501 0.019716
R51595 DVSS.n7780 DVSS.n7779 0.019716
R51596 DVSS.n7779 DVSS.n7500 0.019716
R51597 DVSS.n7773 DVSS.n7772 0.019716
R51598 DVSS.n7772 DVSS.n7499 0.019716
R51599 DVSS.n7768 DVSS.n7767 0.019716
R51600 DVSS.n7767 DVSS.n7498 0.019716
R51601 DVSS.n7761 DVSS.n7760 0.019716
R51602 DVSS.n7760 DVSS.n7497 0.019716
R51603 DVSS.n7756 DVSS.n7755 0.019716
R51604 DVSS.n7755 DVSS.n7496 0.019716
R51605 DVSS.n7749 DVSS.n7748 0.019716
R51606 DVSS.n7748 DVSS.n7495 0.019716
R51607 DVSS.n7744 DVSS.n7743 0.019716
R51608 DVSS.n7743 DVSS.n7494 0.019716
R51609 DVSS.n7737 DVSS.n7736 0.019716
R51610 DVSS.n7736 DVSS.n7493 0.019716
R51611 DVSS.n7732 DVSS.n7731 0.019716
R51612 DVSS.n7731 DVSS.n7492 0.019716
R51613 DVSS.n7725 DVSS.n7724 0.019716
R51614 DVSS.n7724 DVSS.n7491 0.019716
R51615 DVSS.n7720 DVSS.n7719 0.019716
R51616 DVSS.n7719 DVSS.n7490 0.019716
R51617 DVSS.n7713 DVSS.n7712 0.019716
R51618 DVSS.n7712 DVSS.n7489 0.019716
R51619 DVSS.n7708 DVSS.n7707 0.019716
R51620 DVSS.n7707 DVSS.n7488 0.019716
R51621 DVSS.n7701 DVSS.n7700 0.019716
R51622 DVSS.n7700 DVSS.n7487 0.019716
R51623 DVSS.n7696 DVSS.n7695 0.019716
R51624 DVSS.n7695 DVSS.n7486 0.019716
R51625 DVSS.n7689 DVSS.n7688 0.019716
R51626 DVSS.n7688 DVSS.n7485 0.019716
R51627 DVSS.n7684 DVSS.n7683 0.019716
R51628 DVSS.n7683 DVSS.n7484 0.019716
R51629 DVSS.n7677 DVSS.n7676 0.019716
R51630 DVSS.n7676 DVSS.n7483 0.019716
R51631 DVSS.n7672 DVSS.n7671 0.019716
R51632 DVSS.n7671 DVSS.n7482 0.019716
R51633 DVSS.n7665 DVSS.n7664 0.019716
R51634 DVSS.n7664 DVSS.n7481 0.019716
R51635 DVSS.n7660 DVSS.n7659 0.019716
R51636 DVSS.n7659 DVSS.n7480 0.019716
R51637 DVSS.n7653 DVSS.n7652 0.019716
R51638 DVSS.n7652 DVSS.n7479 0.019716
R51639 DVSS.n7648 DVSS.n7647 0.019716
R51640 DVSS.n7647 DVSS.n7478 0.019716
R51641 DVSS.n7641 DVSS.n7640 0.019716
R51642 DVSS.n7640 DVSS.n7477 0.019716
R51643 DVSS.n7636 DVSS.n7635 0.019716
R51644 DVSS.n7635 DVSS.n7476 0.019716
R51645 DVSS.n7629 DVSS.n7628 0.019716
R51646 DVSS.n7628 DVSS.n7475 0.019716
R51647 DVSS.n7624 DVSS.n7623 0.019716
R51648 DVSS.n7623 DVSS.n7474 0.019716
R51649 DVSS.n7617 DVSS.n7616 0.019716
R51650 DVSS.n7616 DVSS.n7473 0.019716
R51651 DVSS.n7612 DVSS.n7611 0.019716
R51652 DVSS.n7611 DVSS.n7472 0.019716
R51653 DVSS.n7605 DVSS.n7604 0.019716
R51654 DVSS.n7604 DVSS.n7471 0.019716
R51655 DVSS.n7600 DVSS.n7599 0.019716
R51656 DVSS.n7599 DVSS.n7470 0.019716
R51657 DVSS.n7593 DVSS.n7592 0.019716
R51658 DVSS.n7592 DVSS.n7469 0.019716
R51659 DVSS.n7588 DVSS.n7587 0.019716
R51660 DVSS.n7587 DVSS.n7468 0.019716
R51661 DVSS.n7581 DVSS.n7580 0.019716
R51662 DVSS.n7580 DVSS.n7467 0.019716
R51663 DVSS.n7576 DVSS.n7575 0.019716
R51664 DVSS.n7575 DVSS.n7466 0.019716
R51665 DVSS.n7569 DVSS.n7568 0.019716
R51666 DVSS.n7568 DVSS.n7465 0.019716
R51667 DVSS.n7564 DVSS.n7563 0.019716
R51668 DVSS.n7563 DVSS.n7464 0.019716
R51669 DVSS.n7557 DVSS.n7556 0.019716
R51670 DVSS.n7556 DVSS.n7463 0.019716
R51671 DVSS.n7552 DVSS.n7551 0.019716
R51672 DVSS.n7551 DVSS.n7462 0.019716
R51673 DVSS.n4804 DVSS.n4803 0.019716
R51674 DVSS.n4802 DVSS.n4801 0.019716
R51675 DVSS.n4801 DVSS.n4476 0.019716
R51676 DVSS.n4795 DVSS.n4481 0.019716
R51677 DVSS.n4795 DVSS.n4794 0.019716
R51678 DVSS.n4792 DVSS.n4791 0.019716
R51679 DVSS.n4791 DVSS.n4482 0.019716
R51680 DVSS.n4785 DVSS.n4487 0.019716
R51681 DVSS.n4785 DVSS.n4784 0.019716
R51682 DVSS.n4782 DVSS.n4781 0.019716
R51683 DVSS.n4781 DVSS.n4488 0.019716
R51684 DVSS.n4775 DVSS.n4493 0.019716
R51685 DVSS.n4775 DVSS.n4774 0.019716
R51686 DVSS.n4772 DVSS.n4771 0.019716
R51687 DVSS.n4771 DVSS.n4494 0.019716
R51688 DVSS.n4765 DVSS.n4499 0.019716
R51689 DVSS.n4765 DVSS.n4764 0.019716
R51690 DVSS.n4762 DVSS.n4761 0.019716
R51691 DVSS.n4761 DVSS.n4500 0.019716
R51692 DVSS.n4755 DVSS.n4505 0.019716
R51693 DVSS.n4755 DVSS.n4754 0.019716
R51694 DVSS.n4752 DVSS.n4751 0.019716
R51695 DVSS.n4751 DVSS.n4506 0.019716
R51696 DVSS.n4745 DVSS.n4511 0.019716
R51697 DVSS.n4745 DVSS.n4744 0.019716
R51698 DVSS.n4742 DVSS.n4741 0.019716
R51699 DVSS.n4741 DVSS.n4512 0.019716
R51700 DVSS.n4735 DVSS.n4517 0.019716
R51701 DVSS.n4735 DVSS.n4734 0.019716
R51702 DVSS.n4732 DVSS.n4731 0.019716
R51703 DVSS.n4731 DVSS.n4518 0.019716
R51704 DVSS.n4725 DVSS.n4523 0.019716
R51705 DVSS.n4725 DVSS.n4724 0.019716
R51706 DVSS.n4722 DVSS.n4721 0.019716
R51707 DVSS.n4721 DVSS.n4524 0.019716
R51708 DVSS.n4715 DVSS.n4529 0.019716
R51709 DVSS.n4715 DVSS.n4714 0.019716
R51710 DVSS.n4712 DVSS.n4711 0.019716
R51711 DVSS.n4711 DVSS.n4530 0.019716
R51712 DVSS.n4705 DVSS.n4535 0.019716
R51713 DVSS.n4705 DVSS.n4704 0.019716
R51714 DVSS.n4702 DVSS.n4701 0.019716
R51715 DVSS.n4701 DVSS.n4536 0.019716
R51716 DVSS.n4695 DVSS.n4541 0.019716
R51717 DVSS.n4695 DVSS.n4694 0.019716
R51718 DVSS.n4692 DVSS.n4691 0.019716
R51719 DVSS.n4691 DVSS.n4542 0.019716
R51720 DVSS.n4685 DVSS.n4547 0.019716
R51721 DVSS.n4685 DVSS.n4684 0.019716
R51722 DVSS.n4682 DVSS.n4681 0.019716
R51723 DVSS.n4681 DVSS.n4548 0.019716
R51724 DVSS.n4675 DVSS.n4553 0.019716
R51725 DVSS.n4675 DVSS.n4674 0.019716
R51726 DVSS.n4672 DVSS.n4671 0.019716
R51727 DVSS.n4671 DVSS.n4554 0.019716
R51728 DVSS.n4665 DVSS.n4559 0.019716
R51729 DVSS.n4665 DVSS.n4664 0.019716
R51730 DVSS.n4662 DVSS.n4661 0.019716
R51731 DVSS.n4661 DVSS.n4560 0.019716
R51732 DVSS.n4655 DVSS.n4565 0.019716
R51733 DVSS.n4655 DVSS.n4654 0.019716
R51734 DVSS.n4652 DVSS.n4651 0.019716
R51735 DVSS.n4651 DVSS.n4566 0.019716
R51736 DVSS.n4645 DVSS.n4571 0.019716
R51737 DVSS.n4645 DVSS.n4644 0.019716
R51738 DVSS.n4642 DVSS.n4641 0.019716
R51739 DVSS.n4641 DVSS.n4572 0.019716
R51740 DVSS.n4635 DVSS.n4577 0.019716
R51741 DVSS.n4635 DVSS.n4634 0.019716
R51742 DVSS.n4632 DVSS.n4631 0.019716
R51743 DVSS.n4631 DVSS.n4578 0.019716
R51744 DVSS.n4625 DVSS.n4583 0.019716
R51745 DVSS.n4625 DVSS.n4624 0.019716
R51746 DVSS.n4622 DVSS.n4621 0.019716
R51747 DVSS.n4621 DVSS.n4584 0.019716
R51748 DVSS.n4615 DVSS.n4589 0.019716
R51749 DVSS.n4615 DVSS.n4614 0.019716
R51750 DVSS.n4612 DVSS.n4611 0.019716
R51751 DVSS.n4611 DVSS.n4590 0.019716
R51752 DVSS.n4605 DVSS.n4595 0.019716
R51753 DVSS.n4605 DVSS.n4604 0.019716
R51754 DVSS.n4602 DVSS.n4601 0.019716
R51755 DVSS.n4601 DVSS.n4596 0.019716
R51756 DVSS.n8089 DVSS.n4414 0.019716
R51757 DVSS.n4416 DVSS.n4415 0.019716
R51758 DVSS.n4416 DVSS.n4412 0.019716
R51759 DVSS.n8080 DVSS.n8079 0.019716
R51760 DVSS.n8079 DVSS.n4411 0.019716
R51761 DVSS.n8075 DVSS.n8074 0.019716
R51762 DVSS.n8074 DVSS.n4410 0.019716
R51763 DVSS.n8068 DVSS.n8067 0.019716
R51764 DVSS.n8067 DVSS.n4409 0.019716
R51765 DVSS.n8063 DVSS.n8062 0.019716
R51766 DVSS.n8062 DVSS.n4408 0.019716
R51767 DVSS.n8056 DVSS.n8055 0.019716
R51768 DVSS.n8055 DVSS.n4407 0.019716
R51769 DVSS.n8051 DVSS.n8050 0.019716
R51770 DVSS.n8050 DVSS.n4406 0.019716
R51771 DVSS.n8044 DVSS.n8043 0.019716
R51772 DVSS.n8043 DVSS.n4405 0.019716
R51773 DVSS.n8039 DVSS.n8038 0.019716
R51774 DVSS.n8038 DVSS.n4404 0.019716
R51775 DVSS.n8032 DVSS.n8031 0.019716
R51776 DVSS.n8031 DVSS.n4403 0.019716
R51777 DVSS.n8027 DVSS.n8026 0.019716
R51778 DVSS.n8026 DVSS.n4402 0.019716
R51779 DVSS.n8020 DVSS.n8019 0.019716
R51780 DVSS.n8019 DVSS.n4401 0.019716
R51781 DVSS.n8015 DVSS.n8014 0.019716
R51782 DVSS.n8014 DVSS.n4400 0.019716
R51783 DVSS.n8008 DVSS.n8007 0.019716
R51784 DVSS.n8007 DVSS.n4399 0.019716
R51785 DVSS.n8003 DVSS.n8002 0.019716
R51786 DVSS.n8002 DVSS.n4398 0.019716
R51787 DVSS.n7996 DVSS.n7995 0.019716
R51788 DVSS.n7995 DVSS.n4397 0.019716
R51789 DVSS.n7991 DVSS.n7990 0.019716
R51790 DVSS.n7990 DVSS.n4396 0.019716
R51791 DVSS.n7984 DVSS.n7983 0.019716
R51792 DVSS.n7983 DVSS.n4395 0.019716
R51793 DVSS.n7979 DVSS.n7978 0.019716
R51794 DVSS.n7978 DVSS.n4394 0.019716
R51795 DVSS.n7972 DVSS.n7971 0.019716
R51796 DVSS.n7971 DVSS.n4393 0.019716
R51797 DVSS.n7967 DVSS.n7966 0.019716
R51798 DVSS.n7966 DVSS.n4392 0.019716
R51799 DVSS.n7960 DVSS.n7959 0.019716
R51800 DVSS.n7959 DVSS.n4391 0.019716
R51801 DVSS.n7955 DVSS.n7954 0.019716
R51802 DVSS.n7954 DVSS.n4390 0.019716
R51803 DVSS.n7948 DVSS.n7947 0.019716
R51804 DVSS.n7947 DVSS.n4389 0.019716
R51805 DVSS.n7943 DVSS.n7942 0.019716
R51806 DVSS.n7942 DVSS.n4388 0.019716
R51807 DVSS.n7936 DVSS.n7935 0.019716
R51808 DVSS.n7935 DVSS.n4387 0.019716
R51809 DVSS.n7931 DVSS.n7930 0.019716
R51810 DVSS.n7930 DVSS.n4386 0.019716
R51811 DVSS.n7924 DVSS.n7923 0.019716
R51812 DVSS.n7923 DVSS.n4385 0.019716
R51813 DVSS.n7919 DVSS.n7918 0.019716
R51814 DVSS.n7918 DVSS.n4384 0.019716
R51815 DVSS.n7912 DVSS.n7911 0.019716
R51816 DVSS.n7911 DVSS.n4383 0.019716
R51817 DVSS.n7907 DVSS.n7906 0.019716
R51818 DVSS.n7906 DVSS.n4382 0.019716
R51819 DVSS.n7900 DVSS.n7899 0.019716
R51820 DVSS.n7899 DVSS.n4381 0.019716
R51821 DVSS.n7895 DVSS.n7894 0.019716
R51822 DVSS.n7894 DVSS.n4380 0.019716
R51823 DVSS.n7888 DVSS.n7887 0.019716
R51824 DVSS.n7887 DVSS.n4379 0.019716
R51825 DVSS.n7883 DVSS.n7882 0.019716
R51826 DVSS.n7882 DVSS.n4378 0.019716
R51827 DVSS.n7876 DVSS.n7875 0.019716
R51828 DVSS.n7875 DVSS.n4377 0.019716
R51829 DVSS.n7871 DVSS.n7870 0.019716
R51830 DVSS.n7870 DVSS.n4376 0.019716
R51831 DVSS.n7864 DVSS.n7863 0.019716
R51832 DVSS.n7863 DVSS.n4375 0.019716
R51833 DVSS.n7859 DVSS.n7858 0.019716
R51834 DVSS.n7858 DVSS.n4374 0.019716
R51835 DVSS.n7852 DVSS.n7851 0.019716
R51836 DVSS.n7851 DVSS.n4373 0.019716
R51837 DVSS.n7847 DVSS.n7846 0.019716
R51838 DVSS.n7846 DVSS.n4372 0.019716
R51839 DVSS.n4111 DVSS.n4110 0.019716
R51840 DVSS.n4115 DVSS.n4112 0.019716
R51841 DVSS.n4115 DVSS.n4114 0.019716
R51842 DVSS.n4121 DVSS.n4104 0.019716
R51843 DVSS.n4122 DVSS.n4121 0.019716
R51844 DVSS.n4127 DVSS.n4124 0.019716
R51845 DVSS.n4127 DVSS.n4126 0.019716
R51846 DVSS.n4133 DVSS.n4100 0.019716
R51847 DVSS.n4134 DVSS.n4133 0.019716
R51848 DVSS.n4139 DVSS.n4136 0.019716
R51849 DVSS.n4139 DVSS.n4138 0.019716
R51850 DVSS.n4145 DVSS.n4096 0.019716
R51851 DVSS.n4146 DVSS.n4145 0.019716
R51852 DVSS.n4151 DVSS.n4148 0.019716
R51853 DVSS.n4151 DVSS.n4150 0.019716
R51854 DVSS.n4157 DVSS.n4092 0.019716
R51855 DVSS.n4158 DVSS.n4157 0.019716
R51856 DVSS.n4163 DVSS.n4160 0.019716
R51857 DVSS.n4163 DVSS.n4162 0.019716
R51858 DVSS.n4169 DVSS.n4088 0.019716
R51859 DVSS.n4170 DVSS.n4169 0.019716
R51860 DVSS.n4175 DVSS.n4172 0.019716
R51861 DVSS.n4175 DVSS.n4174 0.019716
R51862 DVSS.n4181 DVSS.n4084 0.019716
R51863 DVSS.n4182 DVSS.n4181 0.019716
R51864 DVSS.n4187 DVSS.n4184 0.019716
R51865 DVSS.n4187 DVSS.n4186 0.019716
R51866 DVSS.n4193 DVSS.n4080 0.019716
R51867 DVSS.n4194 DVSS.n4193 0.019716
R51868 DVSS.n4199 DVSS.n4196 0.019716
R51869 DVSS.n4199 DVSS.n4198 0.019716
R51870 DVSS.n4205 DVSS.n4076 0.019716
R51871 DVSS.n4206 DVSS.n4205 0.019716
R51872 DVSS.n4211 DVSS.n4208 0.019716
R51873 DVSS.n4211 DVSS.n4210 0.019716
R51874 DVSS.n4217 DVSS.n4072 0.019716
R51875 DVSS.n4218 DVSS.n4217 0.019716
R51876 DVSS.n4223 DVSS.n4220 0.019716
R51877 DVSS.n4223 DVSS.n4222 0.019716
R51878 DVSS.n4229 DVSS.n4068 0.019716
R51879 DVSS.n4230 DVSS.n4229 0.019716
R51880 DVSS.n4235 DVSS.n4232 0.019716
R51881 DVSS.n4235 DVSS.n4234 0.019716
R51882 DVSS.n4241 DVSS.n4064 0.019716
R51883 DVSS.n4242 DVSS.n4241 0.019716
R51884 DVSS.n4247 DVSS.n4244 0.019716
R51885 DVSS.n4247 DVSS.n4246 0.019716
R51886 DVSS.n4253 DVSS.n4060 0.019716
R51887 DVSS.n4254 DVSS.n4253 0.019716
R51888 DVSS.n4259 DVSS.n4256 0.019716
R51889 DVSS.n4259 DVSS.n4258 0.019716
R51890 DVSS.n4265 DVSS.n4056 0.019716
R51891 DVSS.n4266 DVSS.n4265 0.019716
R51892 DVSS.n4271 DVSS.n4268 0.019716
R51893 DVSS.n4271 DVSS.n4270 0.019716
R51894 DVSS.n4277 DVSS.n4052 0.019716
R51895 DVSS.n4278 DVSS.n4277 0.019716
R51896 DVSS.n4283 DVSS.n4280 0.019716
R51897 DVSS.n4283 DVSS.n4282 0.019716
R51898 DVSS.n4289 DVSS.n4048 0.019716
R51899 DVSS.n4290 DVSS.n4289 0.019716
R51900 DVSS.n4295 DVSS.n4292 0.019716
R51901 DVSS.n4295 DVSS.n4294 0.019716
R51902 DVSS.n4301 DVSS.n4044 0.019716
R51903 DVSS.n4302 DVSS.n4301 0.019716
R51904 DVSS.n4307 DVSS.n4304 0.019716
R51905 DVSS.n4307 DVSS.n4306 0.019716
R51906 DVSS.n4313 DVSS.n4040 0.019716
R51907 DVSS.n4314 DVSS.n4313 0.019716
R51908 DVSS.n4319 DVSS.n4316 0.019716
R51909 DVSS.n4319 DVSS.n4318 0.019716
R51910 DVSS.n4325 DVSS.n4036 0.019716
R51911 DVSS.n4326 DVSS.n4325 0.019716
R51912 DVSS.n4331 DVSS.n4328 0.019716
R51913 DVSS.n4331 DVSS.n4330 0.019716
R51914 DVSS.n4337 DVSS.n4032 0.019716
R51915 DVSS.n4338 DVSS.n4337 0.019716
R51916 DVSS.n4343 DVSS.n4340 0.019716
R51917 DVSS.n4343 DVSS.n4342 0.019716
R51918 DVSS.n4350 DVSS.n4028 0.019716
R51919 DVSS.n4351 DVSS.n4350 0.019716
R51920 DVSS.n4354 DVSS.n4353 0.019716
R51921 DVSS.n4355 DVSS.n4354 0.019716
R51922 DVSS.n8319 DVSS.n3901 0.019716
R51923 DVSS.n8133 DVSS.n3945 0.019716
R51924 DVSS.n8133 DVSS.n3899 0.019716
R51925 DVSS.n8137 DVSS.n3944 0.019716
R51926 DVSS.n8137 DVSS.n3898 0.019716
R51927 DVSS.n8142 DVSS.n3943 0.019716
R51928 DVSS.n8142 DVSS.n3897 0.019716
R51929 DVSS.n8146 DVSS.n3942 0.019716
R51930 DVSS.n8146 DVSS.n3896 0.019716
R51931 DVSS.n8151 DVSS.n3941 0.019716
R51932 DVSS.n8151 DVSS.n3895 0.019716
R51933 DVSS.n8155 DVSS.n3940 0.019716
R51934 DVSS.n8155 DVSS.n3894 0.019716
R51935 DVSS.n8160 DVSS.n3939 0.019716
R51936 DVSS.n8160 DVSS.n3893 0.019716
R51937 DVSS.n8164 DVSS.n3938 0.019716
R51938 DVSS.n8164 DVSS.n3892 0.019716
R51939 DVSS.n8169 DVSS.n3937 0.019716
R51940 DVSS.n8169 DVSS.n3891 0.019716
R51941 DVSS.n8173 DVSS.n3936 0.019716
R51942 DVSS.n8173 DVSS.n3890 0.019716
R51943 DVSS.n8178 DVSS.n3935 0.019716
R51944 DVSS.n8178 DVSS.n3889 0.019716
R51945 DVSS.n8182 DVSS.n3934 0.019716
R51946 DVSS.n8182 DVSS.n3888 0.019716
R51947 DVSS.n8187 DVSS.n3933 0.019716
R51948 DVSS.n8187 DVSS.n3887 0.019716
R51949 DVSS.n8191 DVSS.n3932 0.019716
R51950 DVSS.n8191 DVSS.n3886 0.019716
R51951 DVSS.n8196 DVSS.n3931 0.019716
R51952 DVSS.n8196 DVSS.n3885 0.019716
R51953 DVSS.n8200 DVSS.n3930 0.019716
R51954 DVSS.n8200 DVSS.n3884 0.019716
R51955 DVSS.n8205 DVSS.n3929 0.019716
R51956 DVSS.n8205 DVSS.n3883 0.019716
R51957 DVSS.n8209 DVSS.n3928 0.019716
R51958 DVSS.n8209 DVSS.n3882 0.019716
R51959 DVSS.n8214 DVSS.n3927 0.019716
R51960 DVSS.n8214 DVSS.n3881 0.019716
R51961 DVSS.n8218 DVSS.n3926 0.019716
R51962 DVSS.n8218 DVSS.n3880 0.019716
R51963 DVSS.n8223 DVSS.n3925 0.019716
R51964 DVSS.n8223 DVSS.n3879 0.019716
R51965 DVSS.n8227 DVSS.n3924 0.019716
R51966 DVSS.n8227 DVSS.n3878 0.019716
R51967 DVSS.n8232 DVSS.n3923 0.019716
R51968 DVSS.n8232 DVSS.n3877 0.019716
R51969 DVSS.n8236 DVSS.n3922 0.019716
R51970 DVSS.n8236 DVSS.n3876 0.019716
R51971 DVSS.n8241 DVSS.n3921 0.019716
R51972 DVSS.n8241 DVSS.n3875 0.019716
R51973 DVSS.n8245 DVSS.n3920 0.019716
R51974 DVSS.n8245 DVSS.n3874 0.019716
R51975 DVSS.n8250 DVSS.n3919 0.019716
R51976 DVSS.n8250 DVSS.n3873 0.019716
R51977 DVSS.n8254 DVSS.n3918 0.019716
R51978 DVSS.n8254 DVSS.n3872 0.019716
R51979 DVSS.n8259 DVSS.n3917 0.019716
R51980 DVSS.n8259 DVSS.n3871 0.019716
R51981 DVSS.n8263 DVSS.n3916 0.019716
R51982 DVSS.n8263 DVSS.n3870 0.019716
R51983 DVSS.n8268 DVSS.n3915 0.019716
R51984 DVSS.n8268 DVSS.n3869 0.019716
R51985 DVSS.n8272 DVSS.n3914 0.019716
R51986 DVSS.n8272 DVSS.n3868 0.019716
R51987 DVSS.n8277 DVSS.n3913 0.019716
R51988 DVSS.n8277 DVSS.n3867 0.019716
R51989 DVSS.n8281 DVSS.n3912 0.019716
R51990 DVSS.n8281 DVSS.n3866 0.019716
R51991 DVSS.n8286 DVSS.n3911 0.019716
R51992 DVSS.n8286 DVSS.n3865 0.019716
R51993 DVSS.n8290 DVSS.n3910 0.019716
R51994 DVSS.n8290 DVSS.n3864 0.019716
R51995 DVSS.n8295 DVSS.n3909 0.019716
R51996 DVSS.n8295 DVSS.n3863 0.019716
R51997 DVSS.n8299 DVSS.n3908 0.019716
R51998 DVSS.n8299 DVSS.n3862 0.019716
R51999 DVSS.n8304 DVSS.n3907 0.019716
R52000 DVSS.n8304 DVSS.n3861 0.019716
R52001 DVSS.n8308 DVSS.n3906 0.019716
R52002 DVSS.n8308 DVSS.n3860 0.019716
R52003 DVSS.n8313 DVSS.n3905 0.019716
R52004 DVSS.n8313 DVSS.n3859 0.019716
R52005 DVSS.n3841 DVSS.n3840 0.019716
R52006 DVSS.n8344 DVSS.n3796 0.019716
R52007 DVSS.n8345 DVSS.n8344 0.019716
R52008 DVSS.n8350 DVSS.n3795 0.019716
R52009 DVSS.n8350 DVSS.n8349 0.019716
R52010 DVSS.n8356 DVSS.n3794 0.019716
R52011 DVSS.n8357 DVSS.n8356 0.019716
R52012 DVSS.n8362 DVSS.n3793 0.019716
R52013 DVSS.n8362 DVSS.n8361 0.019716
R52014 DVSS.n8368 DVSS.n3792 0.019716
R52015 DVSS.n8369 DVSS.n8368 0.019716
R52016 DVSS.n8374 DVSS.n3791 0.019716
R52017 DVSS.n8374 DVSS.n8373 0.019716
R52018 DVSS.n8380 DVSS.n3790 0.019716
R52019 DVSS.n8381 DVSS.n8380 0.019716
R52020 DVSS.n8386 DVSS.n3789 0.019716
R52021 DVSS.n8386 DVSS.n8385 0.019716
R52022 DVSS.n8392 DVSS.n3788 0.019716
R52023 DVSS.n8393 DVSS.n8392 0.019716
R52024 DVSS.n8398 DVSS.n3787 0.019716
R52025 DVSS.n8398 DVSS.n8397 0.019716
R52026 DVSS.n8404 DVSS.n3786 0.019716
R52027 DVSS.n8405 DVSS.n8404 0.019716
R52028 DVSS.n8410 DVSS.n3785 0.019716
R52029 DVSS.n8410 DVSS.n8409 0.019716
R52030 DVSS.n8416 DVSS.n3784 0.019716
R52031 DVSS.n8417 DVSS.n8416 0.019716
R52032 DVSS.n8422 DVSS.n3783 0.019716
R52033 DVSS.n8422 DVSS.n8421 0.019716
R52034 DVSS.n8428 DVSS.n3782 0.019716
R52035 DVSS.n8429 DVSS.n8428 0.019716
R52036 DVSS.n8434 DVSS.n3781 0.019716
R52037 DVSS.n8434 DVSS.n8433 0.019716
R52038 DVSS.n8440 DVSS.n3780 0.019716
R52039 DVSS.n8441 DVSS.n8440 0.019716
R52040 DVSS.n8446 DVSS.n3779 0.019716
R52041 DVSS.n8446 DVSS.n8445 0.019716
R52042 DVSS.n8452 DVSS.n3778 0.019716
R52043 DVSS.n8453 DVSS.n8452 0.019716
R52044 DVSS.n8458 DVSS.n3777 0.019716
R52045 DVSS.n8458 DVSS.n8457 0.019716
R52046 DVSS.n8464 DVSS.n3776 0.019716
R52047 DVSS.n8465 DVSS.n8464 0.019716
R52048 DVSS.n8470 DVSS.n3775 0.019716
R52049 DVSS.n8470 DVSS.n8469 0.019716
R52050 DVSS.n8476 DVSS.n3774 0.019716
R52051 DVSS.n8477 DVSS.n8476 0.019716
R52052 DVSS.n8482 DVSS.n3773 0.019716
R52053 DVSS.n8482 DVSS.n8481 0.019716
R52054 DVSS.n8488 DVSS.n3772 0.019716
R52055 DVSS.n8489 DVSS.n8488 0.019716
R52056 DVSS.n8494 DVSS.n3771 0.019716
R52057 DVSS.n8494 DVSS.n8493 0.019716
R52058 DVSS.n8500 DVSS.n3770 0.019716
R52059 DVSS.n8501 DVSS.n8500 0.019716
R52060 DVSS.n8506 DVSS.n3769 0.019716
R52061 DVSS.n8506 DVSS.n8505 0.019716
R52062 DVSS.n8512 DVSS.n3768 0.019716
R52063 DVSS.n8513 DVSS.n8512 0.019716
R52064 DVSS.n8518 DVSS.n3767 0.019716
R52065 DVSS.n8518 DVSS.n8517 0.019716
R52066 DVSS.n8524 DVSS.n3766 0.019716
R52067 DVSS.n8525 DVSS.n8524 0.019716
R52068 DVSS.n8530 DVSS.n3765 0.019716
R52069 DVSS.n8530 DVSS.n8529 0.019716
R52070 DVSS.n8536 DVSS.n3764 0.019716
R52071 DVSS.n8537 DVSS.n8536 0.019716
R52072 DVSS.n8542 DVSS.n3763 0.019716
R52073 DVSS.n8542 DVSS.n8541 0.019716
R52074 DVSS.n8548 DVSS.n3762 0.019716
R52075 DVSS.n8549 DVSS.n8548 0.019716
R52076 DVSS.n8554 DVSS.n3761 0.019716
R52077 DVSS.n8554 DVSS.n8553 0.019716
R52078 DVSS.n8560 DVSS.n3760 0.019716
R52079 DVSS.n8561 DVSS.n8560 0.019716
R52080 DVSS.n8566 DVSS.n3759 0.019716
R52081 DVSS.n8566 DVSS.n8565 0.019716
R52082 DVSS.n8572 DVSS.n3758 0.019716
R52083 DVSS.n8573 DVSS.n8572 0.019716
R52084 DVSS.n8578 DVSS.n3757 0.019716
R52085 DVSS.n8578 DVSS.n8577 0.019716
R52086 DVSS.n8585 DVSS.n3756 0.019716
R52087 DVSS.n8586 DVSS.n8585 0.019716
R52088 DVSS.n8603 DVSS.n3458 0.019716
R52089 DVSS.n3563 DVSS.n3501 0.019716
R52090 DVSS.n3563 DVSS.n3456 0.019716
R52091 DVSS.n3571 DVSS.n3500 0.019716
R52092 DVSS.n3571 DVSS.n3455 0.019716
R52093 DVSS.n3560 DVSS.n3499 0.019716
R52094 DVSS.n3560 DVSS.n3454 0.019716
R52095 DVSS.n3580 DVSS.n3498 0.019716
R52096 DVSS.n3580 DVSS.n3453 0.019716
R52097 DVSS.n3557 DVSS.n3497 0.019716
R52098 DVSS.n3557 DVSS.n3452 0.019716
R52099 DVSS.n3589 DVSS.n3496 0.019716
R52100 DVSS.n3589 DVSS.n3451 0.019716
R52101 DVSS.n3554 DVSS.n3495 0.019716
R52102 DVSS.n3554 DVSS.n3450 0.019716
R52103 DVSS.n3598 DVSS.n3494 0.019716
R52104 DVSS.n3598 DVSS.n3449 0.019716
R52105 DVSS.n3551 DVSS.n3493 0.019716
R52106 DVSS.n3551 DVSS.n3448 0.019716
R52107 DVSS.n3607 DVSS.n3492 0.019716
R52108 DVSS.n3607 DVSS.n3447 0.019716
R52109 DVSS.n3548 DVSS.n3491 0.019716
R52110 DVSS.n3548 DVSS.n3446 0.019716
R52111 DVSS.n3616 DVSS.n3490 0.019716
R52112 DVSS.n3616 DVSS.n3445 0.019716
R52113 DVSS.n3545 DVSS.n3489 0.019716
R52114 DVSS.n3545 DVSS.n3444 0.019716
R52115 DVSS.n3625 DVSS.n3488 0.019716
R52116 DVSS.n3625 DVSS.n3443 0.019716
R52117 DVSS.n3542 DVSS.n3487 0.019716
R52118 DVSS.n3542 DVSS.n3442 0.019716
R52119 DVSS.n3634 DVSS.n3486 0.019716
R52120 DVSS.n3634 DVSS.n3441 0.019716
R52121 DVSS.n3539 DVSS.n3485 0.019716
R52122 DVSS.n3539 DVSS.n3440 0.019716
R52123 DVSS.n3643 DVSS.n3484 0.019716
R52124 DVSS.n3643 DVSS.n3439 0.019716
R52125 DVSS.n3536 DVSS.n3483 0.019716
R52126 DVSS.n3536 DVSS.n3438 0.019716
R52127 DVSS.n3652 DVSS.n3482 0.019716
R52128 DVSS.n3652 DVSS.n3437 0.019716
R52129 DVSS.n3533 DVSS.n3481 0.019716
R52130 DVSS.n3533 DVSS.n3436 0.019716
R52131 DVSS.n3661 DVSS.n3480 0.019716
R52132 DVSS.n3661 DVSS.n3435 0.019716
R52133 DVSS.n3530 DVSS.n3479 0.019716
R52134 DVSS.n3530 DVSS.n3434 0.019716
R52135 DVSS.n3670 DVSS.n3478 0.019716
R52136 DVSS.n3670 DVSS.n3433 0.019716
R52137 DVSS.n3527 DVSS.n3477 0.019716
R52138 DVSS.n3527 DVSS.n3432 0.019716
R52139 DVSS.n3679 DVSS.n3476 0.019716
R52140 DVSS.n3679 DVSS.n3431 0.019716
R52141 DVSS.n3524 DVSS.n3475 0.019716
R52142 DVSS.n3524 DVSS.n3430 0.019716
R52143 DVSS.n3688 DVSS.n3474 0.019716
R52144 DVSS.n3688 DVSS.n3429 0.019716
R52145 DVSS.n3521 DVSS.n3473 0.019716
R52146 DVSS.n3521 DVSS.n3428 0.019716
R52147 DVSS.n3697 DVSS.n3472 0.019716
R52148 DVSS.n3697 DVSS.n3427 0.019716
R52149 DVSS.n3518 DVSS.n3471 0.019716
R52150 DVSS.n3518 DVSS.n3426 0.019716
R52151 DVSS.n3706 DVSS.n3470 0.019716
R52152 DVSS.n3706 DVSS.n3425 0.019716
R52153 DVSS.n3515 DVSS.n3469 0.019716
R52154 DVSS.n3515 DVSS.n3424 0.019716
R52155 DVSS.n3715 DVSS.n3468 0.019716
R52156 DVSS.n3715 DVSS.n3423 0.019716
R52157 DVSS.n3512 DVSS.n3467 0.019716
R52158 DVSS.n3512 DVSS.n3422 0.019716
R52159 DVSS.n3724 DVSS.n3466 0.019716
R52160 DVSS.n3724 DVSS.n3421 0.019716
R52161 DVSS.n3509 DVSS.n3465 0.019716
R52162 DVSS.n3509 DVSS.n3420 0.019716
R52163 DVSS.n3733 DVSS.n3464 0.019716
R52164 DVSS.n3733 DVSS.n3419 0.019716
R52165 DVSS.n3506 DVSS.n3463 0.019716
R52166 DVSS.n3506 DVSS.n3418 0.019716
R52167 DVSS.n3742 DVSS.n3462 0.019716
R52168 DVSS.n3742 DVSS.n3417 0.019716
R52169 DVSS.n3503 DVSS.n3461 0.019716
R52170 DVSS.n3503 DVSS.n3416 0.019716
R52171 DVSS.n3155 DVSS.n3154 0.019716
R52172 DVSS.n3159 DVSS.n3156 0.019716
R52173 DVSS.n3159 DVSS.n3158 0.019716
R52174 DVSS.n3165 DVSS.n3148 0.019716
R52175 DVSS.n3166 DVSS.n3165 0.019716
R52176 DVSS.n3171 DVSS.n3168 0.019716
R52177 DVSS.n3171 DVSS.n3170 0.019716
R52178 DVSS.n3177 DVSS.n3144 0.019716
R52179 DVSS.n3178 DVSS.n3177 0.019716
R52180 DVSS.n3183 DVSS.n3180 0.019716
R52181 DVSS.n3183 DVSS.n3182 0.019716
R52182 DVSS.n3189 DVSS.n3140 0.019716
R52183 DVSS.n3190 DVSS.n3189 0.019716
R52184 DVSS.n3195 DVSS.n3192 0.019716
R52185 DVSS.n3195 DVSS.n3194 0.019716
R52186 DVSS.n3201 DVSS.n3136 0.019716
R52187 DVSS.n3202 DVSS.n3201 0.019716
R52188 DVSS.n3207 DVSS.n3204 0.019716
R52189 DVSS.n3207 DVSS.n3206 0.019716
R52190 DVSS.n3213 DVSS.n3132 0.019716
R52191 DVSS.n3214 DVSS.n3213 0.019716
R52192 DVSS.n3219 DVSS.n3216 0.019716
R52193 DVSS.n3219 DVSS.n3218 0.019716
R52194 DVSS.n3225 DVSS.n3128 0.019716
R52195 DVSS.n3226 DVSS.n3225 0.019716
R52196 DVSS.n3231 DVSS.n3228 0.019716
R52197 DVSS.n3231 DVSS.n3230 0.019716
R52198 DVSS.n3237 DVSS.n3124 0.019716
R52199 DVSS.n3238 DVSS.n3237 0.019716
R52200 DVSS.n3243 DVSS.n3240 0.019716
R52201 DVSS.n3243 DVSS.n3242 0.019716
R52202 DVSS.n3249 DVSS.n3120 0.019716
R52203 DVSS.n3250 DVSS.n3249 0.019716
R52204 DVSS.n3255 DVSS.n3252 0.019716
R52205 DVSS.n3255 DVSS.n3254 0.019716
R52206 DVSS.n3261 DVSS.n3116 0.019716
R52207 DVSS.n3262 DVSS.n3261 0.019716
R52208 DVSS.n3267 DVSS.n3264 0.019716
R52209 DVSS.n3267 DVSS.n3266 0.019716
R52210 DVSS.n3273 DVSS.n3112 0.019716
R52211 DVSS.n3274 DVSS.n3273 0.019716
R52212 DVSS.n3279 DVSS.n3276 0.019716
R52213 DVSS.n3279 DVSS.n3278 0.019716
R52214 DVSS.n3285 DVSS.n3108 0.019716
R52215 DVSS.n3286 DVSS.n3285 0.019716
R52216 DVSS.n3291 DVSS.n3288 0.019716
R52217 DVSS.n3291 DVSS.n3290 0.019716
R52218 DVSS.n3297 DVSS.n3104 0.019716
R52219 DVSS.n3298 DVSS.n3297 0.019716
R52220 DVSS.n3303 DVSS.n3300 0.019716
R52221 DVSS.n3303 DVSS.n3302 0.019716
R52222 DVSS.n3309 DVSS.n3100 0.019716
R52223 DVSS.n3310 DVSS.n3309 0.019716
R52224 DVSS.n3315 DVSS.n3312 0.019716
R52225 DVSS.n3315 DVSS.n3314 0.019716
R52226 DVSS.n3321 DVSS.n3096 0.019716
R52227 DVSS.n3322 DVSS.n3321 0.019716
R52228 DVSS.n3327 DVSS.n3324 0.019716
R52229 DVSS.n3327 DVSS.n3326 0.019716
R52230 DVSS.n3333 DVSS.n3092 0.019716
R52231 DVSS.n3334 DVSS.n3333 0.019716
R52232 DVSS.n3339 DVSS.n3336 0.019716
R52233 DVSS.n3339 DVSS.n3338 0.019716
R52234 DVSS.n3345 DVSS.n3088 0.019716
R52235 DVSS.n3346 DVSS.n3345 0.019716
R52236 DVSS.n3351 DVSS.n3348 0.019716
R52237 DVSS.n3351 DVSS.n3350 0.019716
R52238 DVSS.n3357 DVSS.n3084 0.019716
R52239 DVSS.n3358 DVSS.n3357 0.019716
R52240 DVSS.n3363 DVSS.n3360 0.019716
R52241 DVSS.n3363 DVSS.n3362 0.019716
R52242 DVSS.n3369 DVSS.n3080 0.019716
R52243 DVSS.n3370 DVSS.n3369 0.019716
R52244 DVSS.n3375 DVSS.n3372 0.019716
R52245 DVSS.n3375 DVSS.n3374 0.019716
R52246 DVSS.n3381 DVSS.n3076 0.019716
R52247 DVSS.n3382 DVSS.n3381 0.019716
R52248 DVSS.n3387 DVSS.n3384 0.019716
R52249 DVSS.n3387 DVSS.n3386 0.019716
R52250 DVSS.n3394 DVSS.n3072 0.019716
R52251 DVSS.n3395 DVSS.n3394 0.019716
R52252 DVSS.n3398 DVSS.n3397 0.019716
R52253 DVSS.n3399 DVSS.n3398 0.019716
R52254 DVSS.n8968 DVSS.n8677 0.019716
R52255 DVSS.n8679 DVSS.n8678 0.019716
R52256 DVSS.n8679 DVSS.n8676 0.019716
R52257 DVSS.n8959 DVSS.n8958 0.019716
R52258 DVSS.n8958 DVSS.n8675 0.019716
R52259 DVSS.n8954 DVSS.n8953 0.019716
R52260 DVSS.n8953 DVSS.n8674 0.019716
R52261 DVSS.n8947 DVSS.n8946 0.019716
R52262 DVSS.n8946 DVSS.n8673 0.019716
R52263 DVSS.n8942 DVSS.n8941 0.019716
R52264 DVSS.n8941 DVSS.n8672 0.019716
R52265 DVSS.n8935 DVSS.n8934 0.019716
R52266 DVSS.n8934 DVSS.n8671 0.019716
R52267 DVSS.n8930 DVSS.n8929 0.019716
R52268 DVSS.n8929 DVSS.n8670 0.019716
R52269 DVSS.n8923 DVSS.n8922 0.019716
R52270 DVSS.n8922 DVSS.n8669 0.019716
R52271 DVSS.n8918 DVSS.n8917 0.019716
R52272 DVSS.n8917 DVSS.n8668 0.019716
R52273 DVSS.n8911 DVSS.n8910 0.019716
R52274 DVSS.n8910 DVSS.n8667 0.019716
R52275 DVSS.n8906 DVSS.n8905 0.019716
R52276 DVSS.n8905 DVSS.n8666 0.019716
R52277 DVSS.n8899 DVSS.n8898 0.019716
R52278 DVSS.n8898 DVSS.n8665 0.019716
R52279 DVSS.n8894 DVSS.n8893 0.019716
R52280 DVSS.n8893 DVSS.n8664 0.019716
R52281 DVSS.n8887 DVSS.n8886 0.019716
R52282 DVSS.n8886 DVSS.n8663 0.019716
R52283 DVSS.n8882 DVSS.n8881 0.019716
R52284 DVSS.n8881 DVSS.n8662 0.019716
R52285 DVSS.n8875 DVSS.n8874 0.019716
R52286 DVSS.n8874 DVSS.n8661 0.019716
R52287 DVSS.n8870 DVSS.n8869 0.019716
R52288 DVSS.n8869 DVSS.n8660 0.019716
R52289 DVSS.n8863 DVSS.n8862 0.019716
R52290 DVSS.n8862 DVSS.n8659 0.019716
R52291 DVSS.n8858 DVSS.n8857 0.019716
R52292 DVSS.n8857 DVSS.n8658 0.019716
R52293 DVSS.n8851 DVSS.n8850 0.019716
R52294 DVSS.n8850 DVSS.n8657 0.019716
R52295 DVSS.n8846 DVSS.n8845 0.019716
R52296 DVSS.n8845 DVSS.n8656 0.019716
R52297 DVSS.n8839 DVSS.n8838 0.019716
R52298 DVSS.n8838 DVSS.n8655 0.019716
R52299 DVSS.n8834 DVSS.n8833 0.019716
R52300 DVSS.n8833 DVSS.n8654 0.019716
R52301 DVSS.n8827 DVSS.n8826 0.019716
R52302 DVSS.n8826 DVSS.n8653 0.019716
R52303 DVSS.n8822 DVSS.n8821 0.019716
R52304 DVSS.n8821 DVSS.n8652 0.019716
R52305 DVSS.n8815 DVSS.n8814 0.019716
R52306 DVSS.n8814 DVSS.n8651 0.019716
R52307 DVSS.n8810 DVSS.n8809 0.019716
R52308 DVSS.n8809 DVSS.n8650 0.019716
R52309 DVSS.n8803 DVSS.n8802 0.019716
R52310 DVSS.n8802 DVSS.n8649 0.019716
R52311 DVSS.n8798 DVSS.n8797 0.019716
R52312 DVSS.n8797 DVSS.n8648 0.019716
R52313 DVSS.n8791 DVSS.n8790 0.019716
R52314 DVSS.n8790 DVSS.n8647 0.019716
R52315 DVSS.n8786 DVSS.n8785 0.019716
R52316 DVSS.n8785 DVSS.n8646 0.019716
R52317 DVSS.n8779 DVSS.n8778 0.019716
R52318 DVSS.n8778 DVSS.n8645 0.019716
R52319 DVSS.n8774 DVSS.n8773 0.019716
R52320 DVSS.n8773 DVSS.n8644 0.019716
R52321 DVSS.n8767 DVSS.n8766 0.019716
R52322 DVSS.n8766 DVSS.n8643 0.019716
R52323 DVSS.n8762 DVSS.n8761 0.019716
R52324 DVSS.n8761 DVSS.n8642 0.019716
R52325 DVSS.n8755 DVSS.n8754 0.019716
R52326 DVSS.n8754 DVSS.n8641 0.019716
R52327 DVSS.n8750 DVSS.n8749 0.019716
R52328 DVSS.n8749 DVSS.n8640 0.019716
R52329 DVSS.n8743 DVSS.n8742 0.019716
R52330 DVSS.n8742 DVSS.n8639 0.019716
R52331 DVSS.n8738 DVSS.n8737 0.019716
R52332 DVSS.n8737 DVSS.n8638 0.019716
R52333 DVSS.n8731 DVSS.n8730 0.019716
R52334 DVSS.n8730 DVSS.n8637 0.019716
R52335 DVSS.n8726 DVSS.n8725 0.019716
R52336 DVSS.n8725 DVSS.n8636 0.019716
R52337 DVSS.n9186 DVSS.n2933 0.019716
R52338 DVSS.n9000 DVSS.n2978 0.019716
R52339 DVSS.n9000 DVSS.n2931 0.019716
R52340 DVSS.n9004 DVSS.n2977 0.019716
R52341 DVSS.n9004 DVSS.n2930 0.019716
R52342 DVSS.n9009 DVSS.n2976 0.019716
R52343 DVSS.n9009 DVSS.n2929 0.019716
R52344 DVSS.n9013 DVSS.n2975 0.019716
R52345 DVSS.n9013 DVSS.n2928 0.019716
R52346 DVSS.n9018 DVSS.n2974 0.019716
R52347 DVSS.n9018 DVSS.n2927 0.019716
R52348 DVSS.n9022 DVSS.n2973 0.019716
R52349 DVSS.n9022 DVSS.n2926 0.019716
R52350 DVSS.n9027 DVSS.n2972 0.019716
R52351 DVSS.n9027 DVSS.n2925 0.019716
R52352 DVSS.n9031 DVSS.n2971 0.019716
R52353 DVSS.n9031 DVSS.n2924 0.019716
R52354 DVSS.n9036 DVSS.n2970 0.019716
R52355 DVSS.n9036 DVSS.n2923 0.019716
R52356 DVSS.n9040 DVSS.n2969 0.019716
R52357 DVSS.n9040 DVSS.n2922 0.019716
R52358 DVSS.n9045 DVSS.n2968 0.019716
R52359 DVSS.n9045 DVSS.n2921 0.019716
R52360 DVSS.n9049 DVSS.n2967 0.019716
R52361 DVSS.n9049 DVSS.n2920 0.019716
R52362 DVSS.n9054 DVSS.n2966 0.019716
R52363 DVSS.n9054 DVSS.n2919 0.019716
R52364 DVSS.n9058 DVSS.n2965 0.019716
R52365 DVSS.n9058 DVSS.n2918 0.019716
R52366 DVSS.n9063 DVSS.n2964 0.019716
R52367 DVSS.n9063 DVSS.n2917 0.019716
R52368 DVSS.n9067 DVSS.n2963 0.019716
R52369 DVSS.n9067 DVSS.n2916 0.019716
R52370 DVSS.n9072 DVSS.n2962 0.019716
R52371 DVSS.n9072 DVSS.n2915 0.019716
R52372 DVSS.n9076 DVSS.n2961 0.019716
R52373 DVSS.n9076 DVSS.n2914 0.019716
R52374 DVSS.n9081 DVSS.n2960 0.019716
R52375 DVSS.n9081 DVSS.n2913 0.019716
R52376 DVSS.n9085 DVSS.n2959 0.019716
R52377 DVSS.n9085 DVSS.n2912 0.019716
R52378 DVSS.n9090 DVSS.n2958 0.019716
R52379 DVSS.n9090 DVSS.n2911 0.019716
R52380 DVSS.n9094 DVSS.n2957 0.019716
R52381 DVSS.n9094 DVSS.n2910 0.019716
R52382 DVSS.n9099 DVSS.n2956 0.019716
R52383 DVSS.n9099 DVSS.n2909 0.019716
R52384 DVSS.n9103 DVSS.n2955 0.019716
R52385 DVSS.n9103 DVSS.n2908 0.019716
R52386 DVSS.n9108 DVSS.n2954 0.019716
R52387 DVSS.n9108 DVSS.n2907 0.019716
R52388 DVSS.n9112 DVSS.n2953 0.019716
R52389 DVSS.n9112 DVSS.n2906 0.019716
R52390 DVSS.n9117 DVSS.n2952 0.019716
R52391 DVSS.n9117 DVSS.n2905 0.019716
R52392 DVSS.n9121 DVSS.n2951 0.019716
R52393 DVSS.n9121 DVSS.n2904 0.019716
R52394 DVSS.n9126 DVSS.n2950 0.019716
R52395 DVSS.n9126 DVSS.n2903 0.019716
R52396 DVSS.n9130 DVSS.n2949 0.019716
R52397 DVSS.n9130 DVSS.n2902 0.019716
R52398 DVSS.n9135 DVSS.n2948 0.019716
R52399 DVSS.n9135 DVSS.n2901 0.019716
R52400 DVSS.n9139 DVSS.n2947 0.019716
R52401 DVSS.n9139 DVSS.n2900 0.019716
R52402 DVSS.n9144 DVSS.n2946 0.019716
R52403 DVSS.n9144 DVSS.n2899 0.019716
R52404 DVSS.n9148 DVSS.n2945 0.019716
R52405 DVSS.n9148 DVSS.n2898 0.019716
R52406 DVSS.n9153 DVSS.n2944 0.019716
R52407 DVSS.n9153 DVSS.n2897 0.019716
R52408 DVSS.n9157 DVSS.n2943 0.019716
R52409 DVSS.n9157 DVSS.n2896 0.019716
R52410 DVSS.n9162 DVSS.n2942 0.019716
R52411 DVSS.n9162 DVSS.n2895 0.019716
R52412 DVSS.n9166 DVSS.n2941 0.019716
R52413 DVSS.n9166 DVSS.n2894 0.019716
R52414 DVSS.n9171 DVSS.n2940 0.019716
R52415 DVSS.n9171 DVSS.n2893 0.019716
R52416 DVSS.n9175 DVSS.n2939 0.019716
R52417 DVSS.n9175 DVSS.n2892 0.019716
R52418 DVSS.n9180 DVSS.n2938 0.019716
R52419 DVSS.n9180 DVSS.n2891 0.019716
R52420 DVSS.n2873 DVSS.n2872 0.019716
R52421 DVSS.n9211 DVSS.n2828 0.019716
R52422 DVSS.n9212 DVSS.n9211 0.019716
R52423 DVSS.n9217 DVSS.n2827 0.019716
R52424 DVSS.n9217 DVSS.n9216 0.019716
R52425 DVSS.n9223 DVSS.n2826 0.019716
R52426 DVSS.n9224 DVSS.n9223 0.019716
R52427 DVSS.n9229 DVSS.n2825 0.019716
R52428 DVSS.n9229 DVSS.n9228 0.019716
R52429 DVSS.n9235 DVSS.n2824 0.019716
R52430 DVSS.n9236 DVSS.n9235 0.019716
R52431 DVSS.n9241 DVSS.n2823 0.019716
R52432 DVSS.n9241 DVSS.n9240 0.019716
R52433 DVSS.n9247 DVSS.n2822 0.019716
R52434 DVSS.n9248 DVSS.n9247 0.019716
R52435 DVSS.n9253 DVSS.n2821 0.019716
R52436 DVSS.n9253 DVSS.n9252 0.019716
R52437 DVSS.n9259 DVSS.n2820 0.019716
R52438 DVSS.n9260 DVSS.n9259 0.019716
R52439 DVSS.n9265 DVSS.n2819 0.019716
R52440 DVSS.n9265 DVSS.n9264 0.019716
R52441 DVSS.n9271 DVSS.n2818 0.019716
R52442 DVSS.n9272 DVSS.n9271 0.019716
R52443 DVSS.n9277 DVSS.n2817 0.019716
R52444 DVSS.n9277 DVSS.n9276 0.019716
R52445 DVSS.n9283 DVSS.n2816 0.019716
R52446 DVSS.n9284 DVSS.n9283 0.019716
R52447 DVSS.n9289 DVSS.n2815 0.019716
R52448 DVSS.n9289 DVSS.n9288 0.019716
R52449 DVSS.n9295 DVSS.n2814 0.019716
R52450 DVSS.n9296 DVSS.n9295 0.019716
R52451 DVSS.n9301 DVSS.n2813 0.019716
R52452 DVSS.n9301 DVSS.n9300 0.019716
R52453 DVSS.n9307 DVSS.n2812 0.019716
R52454 DVSS.n9308 DVSS.n9307 0.019716
R52455 DVSS.n9313 DVSS.n2811 0.019716
R52456 DVSS.n9313 DVSS.n9312 0.019716
R52457 DVSS.n9319 DVSS.n2810 0.019716
R52458 DVSS.n9320 DVSS.n9319 0.019716
R52459 DVSS.n9325 DVSS.n2809 0.019716
R52460 DVSS.n9325 DVSS.n9324 0.019716
R52461 DVSS.n9331 DVSS.n2808 0.019716
R52462 DVSS.n9332 DVSS.n9331 0.019716
R52463 DVSS.n9337 DVSS.n2807 0.019716
R52464 DVSS.n9337 DVSS.n9336 0.019716
R52465 DVSS.n9343 DVSS.n2806 0.019716
R52466 DVSS.n9344 DVSS.n9343 0.019716
R52467 DVSS.n9349 DVSS.n2805 0.019716
R52468 DVSS.n9349 DVSS.n9348 0.019716
R52469 DVSS.n9355 DVSS.n2804 0.019716
R52470 DVSS.n9356 DVSS.n9355 0.019716
R52471 DVSS.n9361 DVSS.n2803 0.019716
R52472 DVSS.n9361 DVSS.n9360 0.019716
R52473 DVSS.n9367 DVSS.n2802 0.019716
R52474 DVSS.n9368 DVSS.n9367 0.019716
R52475 DVSS.n9373 DVSS.n2801 0.019716
R52476 DVSS.n9373 DVSS.n9372 0.019716
R52477 DVSS.n9379 DVSS.n2800 0.019716
R52478 DVSS.n9380 DVSS.n9379 0.019716
R52479 DVSS.n9385 DVSS.n2799 0.019716
R52480 DVSS.n9385 DVSS.n9384 0.019716
R52481 DVSS.n9391 DVSS.n2798 0.019716
R52482 DVSS.n9392 DVSS.n9391 0.019716
R52483 DVSS.n9397 DVSS.n2797 0.019716
R52484 DVSS.n9397 DVSS.n9396 0.019716
R52485 DVSS.n9403 DVSS.n2796 0.019716
R52486 DVSS.n9404 DVSS.n9403 0.019716
R52487 DVSS.n9409 DVSS.n2795 0.019716
R52488 DVSS.n9409 DVSS.n9408 0.019716
R52489 DVSS.n9415 DVSS.n2794 0.019716
R52490 DVSS.n9416 DVSS.n9415 0.019716
R52491 DVSS.n9421 DVSS.n2793 0.019716
R52492 DVSS.n9421 DVSS.n9420 0.019716
R52493 DVSS.n9427 DVSS.n2792 0.019716
R52494 DVSS.n9428 DVSS.n9427 0.019716
R52495 DVSS.n9433 DVSS.n2791 0.019716
R52496 DVSS.n9433 DVSS.n9432 0.019716
R52497 DVSS.n9439 DVSS.n2790 0.019716
R52498 DVSS.n9440 DVSS.n9439 0.019716
R52499 DVSS.n9445 DVSS.n2789 0.019716
R52500 DVSS.n9445 DVSS.n9444 0.019716
R52501 DVSS.n9452 DVSS.n2788 0.019716
R52502 DVSS.n9453 DVSS.n9452 0.019716
R52503 DVSS.n9758 DVSS.n9466 0.019716
R52504 DVSS.n9468 DVSS.n9467 0.019716
R52505 DVSS.n9468 DVSS.n2780 0.019716
R52506 DVSS.n9749 DVSS.n9748 0.019716
R52507 DVSS.n9748 DVSS.n2779 0.019716
R52508 DVSS.n9744 DVSS.n9743 0.019716
R52509 DVSS.n9743 DVSS.n2778 0.019716
R52510 DVSS.n9737 DVSS.n9736 0.019716
R52511 DVSS.n9736 DVSS.n2777 0.019716
R52512 DVSS.n9732 DVSS.n9731 0.019716
R52513 DVSS.n9731 DVSS.n2776 0.019716
R52514 DVSS.n9725 DVSS.n9724 0.019716
R52515 DVSS.n9724 DVSS.n2775 0.019716
R52516 DVSS.n9720 DVSS.n9719 0.019716
R52517 DVSS.n9719 DVSS.n2774 0.019716
R52518 DVSS.n9713 DVSS.n9712 0.019716
R52519 DVSS.n9712 DVSS.n2773 0.019716
R52520 DVSS.n9708 DVSS.n9707 0.019716
R52521 DVSS.n9707 DVSS.n2772 0.019716
R52522 DVSS.n9701 DVSS.n9700 0.019716
R52523 DVSS.n9700 DVSS.n2771 0.019716
R52524 DVSS.n9696 DVSS.n9695 0.019716
R52525 DVSS.n9695 DVSS.n2770 0.019716
R52526 DVSS.n9689 DVSS.n9688 0.019716
R52527 DVSS.n9688 DVSS.n2769 0.019716
R52528 DVSS.n9684 DVSS.n9683 0.019716
R52529 DVSS.n9683 DVSS.n2768 0.019716
R52530 DVSS.n9677 DVSS.n9676 0.019716
R52531 DVSS.n9676 DVSS.n2767 0.019716
R52532 DVSS.n9672 DVSS.n9671 0.019716
R52533 DVSS.n9671 DVSS.n2766 0.019716
R52534 DVSS.n9665 DVSS.n9664 0.019716
R52535 DVSS.n9664 DVSS.n2765 0.019716
R52536 DVSS.n9660 DVSS.n9659 0.019716
R52537 DVSS.n9659 DVSS.n2764 0.019716
R52538 DVSS.n9653 DVSS.n9652 0.019716
R52539 DVSS.n9652 DVSS.n2763 0.019716
R52540 DVSS.n9648 DVSS.n9647 0.019716
R52541 DVSS.n9647 DVSS.n2762 0.019716
R52542 DVSS.n9641 DVSS.n9640 0.019716
R52543 DVSS.n9640 DVSS.n2761 0.019716
R52544 DVSS.n9636 DVSS.n9635 0.019716
R52545 DVSS.n9635 DVSS.n2760 0.019716
R52546 DVSS.n9629 DVSS.n9628 0.019716
R52547 DVSS.n9628 DVSS.n2759 0.019716
R52548 DVSS.n9624 DVSS.n9623 0.019716
R52549 DVSS.n9623 DVSS.n2758 0.019716
R52550 DVSS.n9617 DVSS.n9616 0.019716
R52551 DVSS.n9616 DVSS.n2757 0.019716
R52552 DVSS.n9612 DVSS.n9611 0.019716
R52553 DVSS.n9611 DVSS.n2756 0.019716
R52554 DVSS.n9605 DVSS.n9604 0.019716
R52555 DVSS.n9604 DVSS.n2755 0.019716
R52556 DVSS.n9600 DVSS.n9599 0.019716
R52557 DVSS.n9599 DVSS.n2754 0.019716
R52558 DVSS.n9593 DVSS.n9592 0.019716
R52559 DVSS.n9592 DVSS.n2753 0.019716
R52560 DVSS.n9588 DVSS.n9587 0.019716
R52561 DVSS.n9587 DVSS.n2752 0.019716
R52562 DVSS.n9581 DVSS.n9580 0.019716
R52563 DVSS.n9580 DVSS.n2751 0.019716
R52564 DVSS.n9576 DVSS.n9575 0.019716
R52565 DVSS.n9575 DVSS.n2750 0.019716
R52566 DVSS.n9569 DVSS.n9568 0.019716
R52567 DVSS.n9568 DVSS.n2749 0.019716
R52568 DVSS.n9564 DVSS.n9563 0.019716
R52569 DVSS.n9563 DVSS.n2748 0.019716
R52570 DVSS.n9557 DVSS.n9556 0.019716
R52571 DVSS.n9556 DVSS.n2747 0.019716
R52572 DVSS.n9552 DVSS.n9551 0.019716
R52573 DVSS.n9551 DVSS.n2746 0.019716
R52574 DVSS.n9545 DVSS.n9544 0.019716
R52575 DVSS.n9544 DVSS.n2745 0.019716
R52576 DVSS.n9540 DVSS.n9539 0.019716
R52577 DVSS.n9539 DVSS.n2744 0.019716
R52578 DVSS.n9533 DVSS.n9532 0.019716
R52579 DVSS.n9532 DVSS.n2743 0.019716
R52580 DVSS.n9528 DVSS.n9527 0.019716
R52581 DVSS.n9527 DVSS.n2742 0.019716
R52582 DVSS.n9521 DVSS.n9520 0.019716
R52583 DVSS.n9520 DVSS.n2741 0.019716
R52584 DVSS.n9516 DVSS.n9515 0.019716
R52585 DVSS.n9515 DVSS.n2740 0.019716
R52586 DVSS.n9862 DVSS.n9861 0.019716
R52587 DVSS.n9866 DVSS.n9863 0.019716
R52588 DVSS.n9866 DVSS.n9865 0.019716
R52589 DVSS.n9872 DVSS.n9855 0.019716
R52590 DVSS.n9873 DVSS.n9872 0.019716
R52591 DVSS.n9878 DVSS.n9875 0.019716
R52592 DVSS.n9878 DVSS.n9877 0.019716
R52593 DVSS.n9884 DVSS.n9851 0.019716
R52594 DVSS.n9885 DVSS.n9884 0.019716
R52595 DVSS.n9890 DVSS.n9887 0.019716
R52596 DVSS.n9890 DVSS.n9889 0.019716
R52597 DVSS.n9896 DVSS.n9847 0.019716
R52598 DVSS.n9897 DVSS.n9896 0.019716
R52599 DVSS.n9902 DVSS.n9899 0.019716
R52600 DVSS.n9902 DVSS.n9901 0.019716
R52601 DVSS.n9908 DVSS.n9843 0.019716
R52602 DVSS.n9909 DVSS.n9908 0.019716
R52603 DVSS.n9914 DVSS.n9911 0.019716
R52604 DVSS.n9914 DVSS.n9913 0.019716
R52605 DVSS.n9920 DVSS.n9839 0.019716
R52606 DVSS.n9921 DVSS.n9920 0.019716
R52607 DVSS.n9926 DVSS.n9923 0.019716
R52608 DVSS.n9926 DVSS.n9925 0.019716
R52609 DVSS.n9932 DVSS.n9835 0.019716
R52610 DVSS.n9933 DVSS.n9932 0.019716
R52611 DVSS.n9938 DVSS.n9935 0.019716
R52612 DVSS.n9938 DVSS.n9937 0.019716
R52613 DVSS.n9944 DVSS.n9831 0.019716
R52614 DVSS.n9945 DVSS.n9944 0.019716
R52615 DVSS.n9950 DVSS.n9947 0.019716
R52616 DVSS.n9950 DVSS.n9949 0.019716
R52617 DVSS.n9956 DVSS.n9827 0.019716
R52618 DVSS.n9957 DVSS.n9956 0.019716
R52619 DVSS.n9962 DVSS.n9959 0.019716
R52620 DVSS.n9962 DVSS.n9961 0.019716
R52621 DVSS.n9968 DVSS.n9823 0.019716
R52622 DVSS.n9969 DVSS.n9968 0.019716
R52623 DVSS.n9974 DVSS.n9971 0.019716
R52624 DVSS.n9974 DVSS.n9973 0.019716
R52625 DVSS.n9980 DVSS.n9819 0.019716
R52626 DVSS.n9981 DVSS.n9980 0.019716
R52627 DVSS.n9986 DVSS.n9983 0.019716
R52628 DVSS.n9986 DVSS.n9985 0.019716
R52629 DVSS.n9992 DVSS.n9815 0.019716
R52630 DVSS.n9993 DVSS.n9992 0.019716
R52631 DVSS.n9998 DVSS.n9995 0.019716
R52632 DVSS.n9998 DVSS.n9997 0.019716
R52633 DVSS.n10004 DVSS.n9811 0.019716
R52634 DVSS.n10005 DVSS.n10004 0.019716
R52635 DVSS.n10010 DVSS.n10007 0.019716
R52636 DVSS.n10010 DVSS.n10009 0.019716
R52637 DVSS.n10016 DVSS.n9807 0.019716
R52638 DVSS.n10017 DVSS.n10016 0.019716
R52639 DVSS.n10022 DVSS.n10019 0.019716
R52640 DVSS.n10022 DVSS.n10021 0.019716
R52641 DVSS.n10028 DVSS.n9803 0.019716
R52642 DVSS.n10029 DVSS.n10028 0.019716
R52643 DVSS.n10034 DVSS.n10031 0.019716
R52644 DVSS.n10034 DVSS.n10033 0.019716
R52645 DVSS.n10040 DVSS.n9799 0.019716
R52646 DVSS.n10041 DVSS.n10040 0.019716
R52647 DVSS.n10046 DVSS.n10043 0.019716
R52648 DVSS.n10046 DVSS.n10045 0.019716
R52649 DVSS.n10052 DVSS.n9795 0.019716
R52650 DVSS.n10053 DVSS.n10052 0.019716
R52651 DVSS.n10058 DVSS.n10055 0.019716
R52652 DVSS.n10058 DVSS.n10057 0.019716
R52653 DVSS.n10064 DVSS.n9791 0.019716
R52654 DVSS.n10065 DVSS.n10064 0.019716
R52655 DVSS.n10070 DVSS.n10067 0.019716
R52656 DVSS.n10070 DVSS.n10069 0.019716
R52657 DVSS.n10076 DVSS.n9787 0.019716
R52658 DVSS.n10077 DVSS.n10076 0.019716
R52659 DVSS.n10082 DVSS.n10079 0.019716
R52660 DVSS.n10082 DVSS.n10081 0.019716
R52661 DVSS.n10088 DVSS.n9783 0.019716
R52662 DVSS.n10089 DVSS.n10088 0.019716
R52663 DVSS.n10094 DVSS.n10091 0.019716
R52664 DVSS.n10094 DVSS.n10093 0.019716
R52665 DVSS.n10101 DVSS.n9779 0.019716
R52666 DVSS.n10102 DVSS.n10101 0.019716
R52667 DVSS.n10105 DVSS.n10104 0.019716
R52668 DVSS.n10106 DVSS.n10105 0.019716
R52669 DVSS.n2457 DVSS.n2456 0.019716
R52670 DVSS.n2464 DVSS.n2411 0.019716
R52671 DVSS.n2465 DVSS.n2464 0.019716
R52672 DVSS.n2470 DVSS.n2410 0.019716
R52673 DVSS.n2470 DVSS.n2469 0.019716
R52674 DVSS.n2476 DVSS.n2409 0.019716
R52675 DVSS.n2477 DVSS.n2476 0.019716
R52676 DVSS.n2482 DVSS.n2408 0.019716
R52677 DVSS.n2482 DVSS.n2481 0.019716
R52678 DVSS.n2488 DVSS.n2407 0.019716
R52679 DVSS.n2489 DVSS.n2488 0.019716
R52680 DVSS.n2494 DVSS.n2406 0.019716
R52681 DVSS.n2494 DVSS.n2493 0.019716
R52682 DVSS.n2500 DVSS.n2405 0.019716
R52683 DVSS.n2501 DVSS.n2500 0.019716
R52684 DVSS.n2506 DVSS.n2404 0.019716
R52685 DVSS.n2506 DVSS.n2505 0.019716
R52686 DVSS.n2512 DVSS.n2403 0.019716
R52687 DVSS.n2513 DVSS.n2512 0.019716
R52688 DVSS.n2518 DVSS.n2402 0.019716
R52689 DVSS.n2518 DVSS.n2517 0.019716
R52690 DVSS.n2524 DVSS.n2401 0.019716
R52691 DVSS.n2525 DVSS.n2524 0.019716
R52692 DVSS.n2530 DVSS.n2400 0.019716
R52693 DVSS.n2530 DVSS.n2529 0.019716
R52694 DVSS.n2536 DVSS.n2399 0.019716
R52695 DVSS.n2537 DVSS.n2536 0.019716
R52696 DVSS.n2542 DVSS.n2398 0.019716
R52697 DVSS.n2542 DVSS.n2541 0.019716
R52698 DVSS.n2548 DVSS.n2397 0.019716
R52699 DVSS.n2549 DVSS.n2548 0.019716
R52700 DVSS.n2554 DVSS.n2396 0.019716
R52701 DVSS.n2554 DVSS.n2553 0.019716
R52702 DVSS.n2560 DVSS.n2395 0.019716
R52703 DVSS.n2561 DVSS.n2560 0.019716
R52704 DVSS.n2566 DVSS.n2394 0.019716
R52705 DVSS.n2566 DVSS.n2565 0.019716
R52706 DVSS.n2572 DVSS.n2393 0.019716
R52707 DVSS.n2573 DVSS.n2572 0.019716
R52708 DVSS.n2578 DVSS.n2392 0.019716
R52709 DVSS.n2578 DVSS.n2577 0.019716
R52710 DVSS.n2584 DVSS.n2391 0.019716
R52711 DVSS.n2585 DVSS.n2584 0.019716
R52712 DVSS.n2590 DVSS.n2390 0.019716
R52713 DVSS.n2590 DVSS.n2589 0.019716
R52714 DVSS.n2596 DVSS.n2389 0.019716
R52715 DVSS.n2597 DVSS.n2596 0.019716
R52716 DVSS.n2602 DVSS.n2388 0.019716
R52717 DVSS.n2602 DVSS.n2601 0.019716
R52718 DVSS.n2608 DVSS.n2387 0.019716
R52719 DVSS.n2609 DVSS.n2608 0.019716
R52720 DVSS.n2614 DVSS.n2386 0.019716
R52721 DVSS.n2614 DVSS.n2613 0.019716
R52722 DVSS.n2620 DVSS.n2385 0.019716
R52723 DVSS.n2621 DVSS.n2620 0.019716
R52724 DVSS.n2626 DVSS.n2384 0.019716
R52725 DVSS.n2626 DVSS.n2625 0.019716
R52726 DVSS.n2632 DVSS.n2383 0.019716
R52727 DVSS.n2633 DVSS.n2632 0.019716
R52728 DVSS.n2638 DVSS.n2382 0.019716
R52729 DVSS.n2638 DVSS.n2637 0.019716
R52730 DVSS.n2644 DVSS.n2381 0.019716
R52731 DVSS.n2645 DVSS.n2644 0.019716
R52732 DVSS.n2650 DVSS.n2380 0.019716
R52733 DVSS.n2650 DVSS.n2649 0.019716
R52734 DVSS.n2656 DVSS.n2379 0.019716
R52735 DVSS.n2657 DVSS.n2656 0.019716
R52736 DVSS.n2662 DVSS.n2378 0.019716
R52737 DVSS.n2662 DVSS.n2661 0.019716
R52738 DVSS.n2668 DVSS.n2377 0.019716
R52739 DVSS.n2669 DVSS.n2668 0.019716
R52740 DVSS.n2674 DVSS.n2376 0.019716
R52741 DVSS.n2674 DVSS.n2673 0.019716
R52742 DVSS.n2680 DVSS.n2375 0.019716
R52743 DVSS.n2681 DVSS.n2680 0.019716
R52744 DVSS.n2686 DVSS.n2374 0.019716
R52745 DVSS.n2686 DVSS.n2685 0.019716
R52746 DVSS.n2692 DVSS.n2373 0.019716
R52747 DVSS.n2693 DVSS.n2692 0.019716
R52748 DVSS.n2698 DVSS.n2372 0.019716
R52749 DVSS.n2698 DVSS.n2697 0.019716
R52750 DVSS.n10138 DVSS.n2371 0.019716
R52751 DVSS.n10139 DVSS.n10138 0.019716
R52752 DVSS.n2115 DVSS.n2114 0.019716
R52753 DVSS.n2122 DVSS.n2068 0.019716
R52754 DVSS.n2123 DVSS.n2122 0.019716
R52755 DVSS.n2128 DVSS.n2067 0.019716
R52756 DVSS.n2128 DVSS.n2127 0.019716
R52757 DVSS.n2134 DVSS.n2066 0.019716
R52758 DVSS.n2135 DVSS.n2134 0.019716
R52759 DVSS.n2140 DVSS.n2065 0.019716
R52760 DVSS.n2140 DVSS.n2139 0.019716
R52761 DVSS.n2146 DVSS.n2064 0.019716
R52762 DVSS.n2147 DVSS.n2146 0.019716
R52763 DVSS.n2152 DVSS.n2063 0.019716
R52764 DVSS.n2152 DVSS.n2151 0.019716
R52765 DVSS.n2158 DVSS.n2062 0.019716
R52766 DVSS.n2159 DVSS.n2158 0.019716
R52767 DVSS.n2164 DVSS.n2061 0.019716
R52768 DVSS.n2164 DVSS.n2163 0.019716
R52769 DVSS.n2170 DVSS.n2060 0.019716
R52770 DVSS.n2171 DVSS.n2170 0.019716
R52771 DVSS.n2176 DVSS.n2059 0.019716
R52772 DVSS.n2176 DVSS.n2175 0.019716
R52773 DVSS.n2182 DVSS.n2058 0.019716
R52774 DVSS.n2183 DVSS.n2182 0.019716
R52775 DVSS.n2188 DVSS.n2057 0.019716
R52776 DVSS.n2188 DVSS.n2187 0.019716
R52777 DVSS.n2194 DVSS.n2056 0.019716
R52778 DVSS.n2195 DVSS.n2194 0.019716
R52779 DVSS.n2200 DVSS.n2055 0.019716
R52780 DVSS.n2200 DVSS.n2199 0.019716
R52781 DVSS.n2206 DVSS.n2054 0.019716
R52782 DVSS.n2207 DVSS.n2206 0.019716
R52783 DVSS.n2212 DVSS.n2053 0.019716
R52784 DVSS.n2212 DVSS.n2211 0.019716
R52785 DVSS.n2218 DVSS.n2052 0.019716
R52786 DVSS.n2219 DVSS.n2218 0.019716
R52787 DVSS.n2224 DVSS.n2051 0.019716
R52788 DVSS.n2224 DVSS.n2223 0.019716
R52789 DVSS.n2230 DVSS.n2050 0.019716
R52790 DVSS.n2231 DVSS.n2230 0.019716
R52791 DVSS.n2236 DVSS.n2049 0.019716
R52792 DVSS.n2236 DVSS.n2235 0.019716
R52793 DVSS.n2242 DVSS.n2048 0.019716
R52794 DVSS.n2243 DVSS.n2242 0.019716
R52795 DVSS.n2248 DVSS.n2047 0.019716
R52796 DVSS.n2248 DVSS.n2247 0.019716
R52797 DVSS.n2254 DVSS.n2046 0.019716
R52798 DVSS.n2255 DVSS.n2254 0.019716
R52799 DVSS.n2260 DVSS.n2045 0.019716
R52800 DVSS.n2260 DVSS.n2259 0.019716
R52801 DVSS.n2266 DVSS.n2044 0.019716
R52802 DVSS.n2267 DVSS.n2266 0.019716
R52803 DVSS.n2272 DVSS.n2043 0.019716
R52804 DVSS.n2272 DVSS.n2271 0.019716
R52805 DVSS.n2278 DVSS.n2042 0.019716
R52806 DVSS.n2279 DVSS.n2278 0.019716
R52807 DVSS.n2284 DVSS.n2041 0.019716
R52808 DVSS.n2284 DVSS.n2283 0.019716
R52809 DVSS.n2290 DVSS.n2040 0.019716
R52810 DVSS.n2291 DVSS.n2290 0.019716
R52811 DVSS.n2296 DVSS.n2039 0.019716
R52812 DVSS.n2296 DVSS.n2295 0.019716
R52813 DVSS.n2302 DVSS.n2038 0.019716
R52814 DVSS.n2303 DVSS.n2302 0.019716
R52815 DVSS.n2308 DVSS.n2037 0.019716
R52816 DVSS.n2308 DVSS.n2307 0.019716
R52817 DVSS.n2314 DVSS.n2036 0.019716
R52818 DVSS.n2315 DVSS.n2314 0.019716
R52819 DVSS.n2320 DVSS.n2035 0.019716
R52820 DVSS.n2320 DVSS.n2319 0.019716
R52821 DVSS.n2326 DVSS.n2034 0.019716
R52822 DVSS.n2327 DVSS.n2326 0.019716
R52823 DVSS.n2332 DVSS.n2033 0.019716
R52824 DVSS.n2332 DVSS.n2331 0.019716
R52825 DVSS.n2338 DVSS.n2032 0.019716
R52826 DVSS.n2339 DVSS.n2338 0.019716
R52827 DVSS.n2344 DVSS.n2031 0.019716
R52828 DVSS.n2344 DVSS.n2343 0.019716
R52829 DVSS.n2350 DVSS.n2030 0.019716
R52830 DVSS.n2351 DVSS.n2350 0.019716
R52831 DVSS.n2356 DVSS.n2029 0.019716
R52832 DVSS.n2356 DVSS.n2355 0.019716
R52833 DVSS.n10163 DVSS.n2028 0.019716
R52834 DVSS.n10164 DVSS.n10163 0.019716
R52835 DVSS.n10452 DVSS.n10451 0.019716
R52836 DVSS.n10449 DVSS.n2008 0.019716
R52837 DVSS.n10449 DVSS.n10448 0.019716
R52838 DVSS.n10442 DVSS.n2007 0.019716
R52839 DVSS.n10442 DVSS.n10441 0.019716
R52840 DVSS.n10437 DVSS.n2006 0.019716
R52841 DVSS.n10437 DVSS.n10436 0.019716
R52842 DVSS.n10430 DVSS.n2005 0.019716
R52843 DVSS.n10430 DVSS.n10429 0.019716
R52844 DVSS.n10425 DVSS.n2004 0.019716
R52845 DVSS.n10425 DVSS.n10424 0.019716
R52846 DVSS.n10418 DVSS.n2003 0.019716
R52847 DVSS.n10418 DVSS.n10417 0.019716
R52848 DVSS.n10413 DVSS.n2002 0.019716
R52849 DVSS.n10413 DVSS.n10412 0.019716
R52850 DVSS.n10406 DVSS.n2001 0.019716
R52851 DVSS.n10406 DVSS.n10405 0.019716
R52852 DVSS.n10401 DVSS.n2000 0.019716
R52853 DVSS.n10401 DVSS.n10400 0.019716
R52854 DVSS.n10394 DVSS.n1999 0.019716
R52855 DVSS.n10394 DVSS.n10393 0.019716
R52856 DVSS.n10389 DVSS.n1998 0.019716
R52857 DVSS.n10389 DVSS.n10388 0.019716
R52858 DVSS.n10382 DVSS.n1997 0.019716
R52859 DVSS.n10382 DVSS.n10381 0.019716
R52860 DVSS.n10377 DVSS.n1996 0.019716
R52861 DVSS.n10377 DVSS.n10376 0.019716
R52862 DVSS.n10370 DVSS.n1995 0.019716
R52863 DVSS.n10370 DVSS.n10369 0.019716
R52864 DVSS.n10365 DVSS.n1994 0.019716
R52865 DVSS.n10365 DVSS.n10364 0.019716
R52866 DVSS.n10358 DVSS.n1993 0.019716
R52867 DVSS.n10358 DVSS.n10357 0.019716
R52868 DVSS.n10353 DVSS.n1992 0.019716
R52869 DVSS.n10353 DVSS.n10352 0.019716
R52870 DVSS.n10346 DVSS.n1991 0.019716
R52871 DVSS.n10346 DVSS.n10345 0.019716
R52872 DVSS.n10341 DVSS.n1990 0.019716
R52873 DVSS.n10341 DVSS.n10340 0.019716
R52874 DVSS.n10334 DVSS.n1989 0.019716
R52875 DVSS.n10334 DVSS.n10333 0.019716
R52876 DVSS.n10329 DVSS.n1988 0.019716
R52877 DVSS.n10329 DVSS.n10328 0.019716
R52878 DVSS.n10322 DVSS.n1987 0.019716
R52879 DVSS.n10322 DVSS.n10321 0.019716
R52880 DVSS.n10317 DVSS.n1986 0.019716
R52881 DVSS.n10317 DVSS.n10316 0.019716
R52882 DVSS.n10310 DVSS.n1985 0.019716
R52883 DVSS.n10310 DVSS.n10309 0.019716
R52884 DVSS.n10305 DVSS.n1984 0.019716
R52885 DVSS.n10305 DVSS.n10304 0.019716
R52886 DVSS.n10298 DVSS.n1983 0.019716
R52887 DVSS.n10298 DVSS.n10297 0.019716
R52888 DVSS.n10293 DVSS.n1982 0.019716
R52889 DVSS.n10293 DVSS.n10292 0.019716
R52890 DVSS.n10286 DVSS.n1981 0.019716
R52891 DVSS.n10286 DVSS.n10285 0.019716
R52892 DVSS.n10281 DVSS.n1980 0.019716
R52893 DVSS.n10281 DVSS.n10280 0.019716
R52894 DVSS.n10274 DVSS.n1979 0.019716
R52895 DVSS.n10274 DVSS.n10273 0.019716
R52896 DVSS.n10269 DVSS.n1978 0.019716
R52897 DVSS.n10269 DVSS.n10268 0.019716
R52898 DVSS.n10262 DVSS.n1977 0.019716
R52899 DVSS.n10262 DVSS.n10261 0.019716
R52900 DVSS.n10257 DVSS.n1976 0.019716
R52901 DVSS.n10257 DVSS.n10256 0.019716
R52902 DVSS.n10250 DVSS.n1975 0.019716
R52903 DVSS.n10250 DVSS.n10249 0.019716
R52904 DVSS.n10245 DVSS.n1974 0.019716
R52905 DVSS.n10245 DVSS.n10244 0.019716
R52906 DVSS.n10238 DVSS.n1973 0.019716
R52907 DVSS.n10238 DVSS.n10237 0.019716
R52908 DVSS.n10233 DVSS.n1972 0.019716
R52909 DVSS.n10233 DVSS.n10232 0.019716
R52910 DVSS.n10226 DVSS.n1971 0.019716
R52911 DVSS.n10226 DVSS.n10225 0.019716
R52912 DVSS.n10221 DVSS.n1970 0.019716
R52913 DVSS.n10221 DVSS.n10220 0.019716
R52914 DVSS.n10214 DVSS.n1969 0.019716
R52915 DVSS.n10214 DVSS.n10213 0.019716
R52916 DVSS.n10472 DVSS.n1968 0.019716
R52917 DVSS.n10473 DVSS.n10472 0.019716
R52918 DVSS.n1960 DVSS.n1668 0.019716
R52919 DVSS.n1671 DVSS.n1670 0.019716
R52920 DVSS.n1671 DVSS.n1667 0.019716
R52921 DVSS.n1951 DVSS.n1950 0.019716
R52922 DVSS.n1950 DVSS.n1666 0.019716
R52923 DVSS.n1946 DVSS.n1945 0.019716
R52924 DVSS.n1945 DVSS.n1665 0.019716
R52925 DVSS.n1939 DVSS.n1938 0.019716
R52926 DVSS.n1938 DVSS.n1664 0.019716
R52927 DVSS.n1934 DVSS.n1933 0.019716
R52928 DVSS.n1933 DVSS.n1663 0.019716
R52929 DVSS.n1927 DVSS.n1926 0.019716
R52930 DVSS.n1926 DVSS.n1662 0.019716
R52931 DVSS.n1922 DVSS.n1921 0.019716
R52932 DVSS.n1921 DVSS.n1661 0.019716
R52933 DVSS.n1915 DVSS.n1914 0.019716
R52934 DVSS.n1914 DVSS.n1660 0.019716
R52935 DVSS.n1910 DVSS.n1909 0.019716
R52936 DVSS.n1909 DVSS.n1659 0.019716
R52937 DVSS.n1903 DVSS.n1902 0.019716
R52938 DVSS.n1902 DVSS.n1658 0.019716
R52939 DVSS.n1898 DVSS.n1897 0.019716
R52940 DVSS.n1897 DVSS.n1657 0.019716
R52941 DVSS.n1891 DVSS.n1890 0.019716
R52942 DVSS.n1890 DVSS.n1656 0.019716
R52943 DVSS.n1886 DVSS.n1885 0.019716
R52944 DVSS.n1885 DVSS.n1655 0.019716
R52945 DVSS.n1879 DVSS.n1878 0.019716
R52946 DVSS.n1878 DVSS.n1654 0.019716
R52947 DVSS.n1874 DVSS.n1873 0.019716
R52948 DVSS.n1873 DVSS.n1653 0.019716
R52949 DVSS.n1867 DVSS.n1866 0.019716
R52950 DVSS.n1866 DVSS.n1652 0.019716
R52951 DVSS.n1862 DVSS.n1861 0.019716
R52952 DVSS.n1861 DVSS.n1651 0.019716
R52953 DVSS.n1855 DVSS.n1854 0.019716
R52954 DVSS.n1854 DVSS.n1650 0.019716
R52955 DVSS.n1850 DVSS.n1849 0.019716
R52956 DVSS.n1849 DVSS.n1649 0.019716
R52957 DVSS.n1843 DVSS.n1842 0.019716
R52958 DVSS.n1842 DVSS.n1648 0.019716
R52959 DVSS.n1838 DVSS.n1837 0.019716
R52960 DVSS.n1837 DVSS.n1647 0.019716
R52961 DVSS.n1831 DVSS.n1830 0.019716
R52962 DVSS.n1830 DVSS.n1646 0.019716
R52963 DVSS.n1826 DVSS.n1825 0.019716
R52964 DVSS.n1825 DVSS.n1645 0.019716
R52965 DVSS.n1819 DVSS.n1818 0.019716
R52966 DVSS.n1818 DVSS.n1644 0.019716
R52967 DVSS.n1814 DVSS.n1813 0.019716
R52968 DVSS.n1813 DVSS.n1643 0.019716
R52969 DVSS.n1807 DVSS.n1806 0.019716
R52970 DVSS.n1806 DVSS.n1642 0.019716
R52971 DVSS.n1802 DVSS.n1801 0.019716
R52972 DVSS.n1801 DVSS.n1641 0.019716
R52973 DVSS.n1795 DVSS.n1794 0.019716
R52974 DVSS.n1794 DVSS.n1640 0.019716
R52975 DVSS.n1790 DVSS.n1789 0.019716
R52976 DVSS.n1789 DVSS.n1639 0.019716
R52977 DVSS.n1783 DVSS.n1782 0.019716
R52978 DVSS.n1782 DVSS.n1638 0.019716
R52979 DVSS.n1778 DVSS.n1777 0.019716
R52980 DVSS.n1777 DVSS.n1637 0.019716
R52981 DVSS.n1771 DVSS.n1770 0.019716
R52982 DVSS.n1770 DVSS.n1636 0.019716
R52983 DVSS.n1766 DVSS.n1765 0.019716
R52984 DVSS.n1765 DVSS.n1635 0.019716
R52985 DVSS.n1759 DVSS.n1758 0.019716
R52986 DVSS.n1758 DVSS.n1634 0.019716
R52987 DVSS.n1754 DVSS.n1753 0.019716
R52988 DVSS.n1753 DVSS.n1633 0.019716
R52989 DVSS.n1747 DVSS.n1746 0.019716
R52990 DVSS.n1746 DVSS.n1632 0.019716
R52991 DVSS.n1742 DVSS.n1741 0.019716
R52992 DVSS.n1741 DVSS.n1631 0.019716
R52993 DVSS.n1735 DVSS.n1734 0.019716
R52994 DVSS.n1734 DVSS.n1630 0.019716
R52995 DVSS.n1730 DVSS.n1729 0.019716
R52996 DVSS.n1729 DVSS.n1629 0.019716
R52997 DVSS.n1723 DVSS.n1722 0.019716
R52998 DVSS.n1722 DVSS.n1628 0.019716
R52999 DVSS.n1718 DVSS.n1717 0.019716
R53000 DVSS.n1717 DVSS.n1627 0.019716
R53001 DVSS.n1610 DVSS.n1609 0.019716
R53002 DVSS.n10511 DVSS.n1564 0.019716
R53003 DVSS.n10512 DVSS.n10511 0.019716
R53004 DVSS.n10517 DVSS.n1563 0.019716
R53005 DVSS.n10517 DVSS.n10516 0.019716
R53006 DVSS.n10523 DVSS.n1562 0.019716
R53007 DVSS.n10524 DVSS.n10523 0.019716
R53008 DVSS.n10529 DVSS.n1561 0.019716
R53009 DVSS.n10529 DVSS.n10528 0.019716
R53010 DVSS.n10535 DVSS.n1560 0.019716
R53011 DVSS.n10536 DVSS.n10535 0.019716
R53012 DVSS.n10541 DVSS.n1559 0.019716
R53013 DVSS.n10541 DVSS.n10540 0.019716
R53014 DVSS.n10547 DVSS.n1558 0.019716
R53015 DVSS.n10548 DVSS.n10547 0.019716
R53016 DVSS.n10553 DVSS.n1557 0.019716
R53017 DVSS.n10553 DVSS.n10552 0.019716
R53018 DVSS.n10559 DVSS.n1556 0.019716
R53019 DVSS.n10560 DVSS.n10559 0.019716
R53020 DVSS.n10565 DVSS.n1555 0.019716
R53021 DVSS.n10565 DVSS.n10564 0.019716
R53022 DVSS.n10571 DVSS.n1554 0.019716
R53023 DVSS.n10572 DVSS.n10571 0.019716
R53024 DVSS.n10577 DVSS.n1553 0.019716
R53025 DVSS.n10577 DVSS.n10576 0.019716
R53026 DVSS.n10583 DVSS.n1552 0.019716
R53027 DVSS.n10584 DVSS.n10583 0.019716
R53028 DVSS.n10589 DVSS.n1551 0.019716
R53029 DVSS.n10589 DVSS.n10588 0.019716
R53030 DVSS.n10595 DVSS.n1550 0.019716
R53031 DVSS.n10596 DVSS.n10595 0.019716
R53032 DVSS.n10601 DVSS.n1549 0.019716
R53033 DVSS.n10601 DVSS.n10600 0.019716
R53034 DVSS.n10607 DVSS.n1548 0.019716
R53035 DVSS.n10608 DVSS.n10607 0.019716
R53036 DVSS.n10613 DVSS.n1547 0.019716
R53037 DVSS.n10613 DVSS.n10612 0.019716
R53038 DVSS.n10619 DVSS.n1546 0.019716
R53039 DVSS.n10620 DVSS.n10619 0.019716
R53040 DVSS.n10625 DVSS.n1545 0.019716
R53041 DVSS.n10625 DVSS.n10624 0.019716
R53042 DVSS.n10631 DVSS.n1544 0.019716
R53043 DVSS.n10632 DVSS.n10631 0.019716
R53044 DVSS.n10637 DVSS.n1543 0.019716
R53045 DVSS.n10637 DVSS.n10636 0.019716
R53046 DVSS.n10643 DVSS.n1542 0.019716
R53047 DVSS.n10644 DVSS.n10643 0.019716
R53048 DVSS.n10649 DVSS.n1541 0.019716
R53049 DVSS.n10649 DVSS.n10648 0.019716
R53050 DVSS.n10655 DVSS.n1540 0.019716
R53051 DVSS.n10656 DVSS.n10655 0.019716
R53052 DVSS.n10661 DVSS.n1539 0.019716
R53053 DVSS.n10661 DVSS.n10660 0.019716
R53054 DVSS.n10667 DVSS.n1538 0.019716
R53055 DVSS.n10668 DVSS.n10667 0.019716
R53056 DVSS.n10673 DVSS.n1537 0.019716
R53057 DVSS.n10673 DVSS.n10672 0.019716
R53058 DVSS.n10679 DVSS.n1536 0.019716
R53059 DVSS.n10680 DVSS.n10679 0.019716
R53060 DVSS.n10685 DVSS.n1535 0.019716
R53061 DVSS.n10685 DVSS.n10684 0.019716
R53062 DVSS.n10691 DVSS.n1534 0.019716
R53063 DVSS.n10692 DVSS.n10691 0.019716
R53064 DVSS.n10697 DVSS.n1533 0.019716
R53065 DVSS.n10697 DVSS.n10696 0.019716
R53066 DVSS.n10703 DVSS.n1532 0.019716
R53067 DVSS.n10704 DVSS.n10703 0.019716
R53068 DVSS.n10709 DVSS.n1531 0.019716
R53069 DVSS.n10709 DVSS.n10708 0.019716
R53070 DVSS.n10715 DVSS.n1530 0.019716
R53071 DVSS.n10716 DVSS.n10715 0.019716
R53072 DVSS.n10721 DVSS.n1529 0.019716
R53073 DVSS.n10721 DVSS.n10720 0.019716
R53074 DVSS.n10727 DVSS.n1528 0.019716
R53075 DVSS.n10728 DVSS.n10727 0.019716
R53076 DVSS.n10733 DVSS.n1527 0.019716
R53077 DVSS.n10733 DVSS.n10732 0.019716
R53078 DVSS.n10739 DVSS.n1526 0.019716
R53079 DVSS.n10740 DVSS.n10739 0.019716
R53080 DVSS.n10745 DVSS.n1525 0.019716
R53081 DVSS.n10745 DVSS.n10744 0.019716
R53082 DVSS.n10751 DVSS.n1524 0.019716
R53083 DVSS.n10752 DVSS.n10751 0.019716
R53084 DVSS.n11101 DVSS.n11100 0.019716
R53085 DVSS.n11099 DVSS.n11098 0.019716
R53086 DVSS.n11098 DVSS.n10773 0.019716
R53087 DVSS.n11092 DVSS.n10778 0.019716
R53088 DVSS.n11092 DVSS.n11091 0.019716
R53089 DVSS.n11089 DVSS.n11088 0.019716
R53090 DVSS.n11088 DVSS.n10779 0.019716
R53091 DVSS.n11082 DVSS.n10784 0.019716
R53092 DVSS.n11082 DVSS.n11081 0.019716
R53093 DVSS.n11079 DVSS.n11078 0.019716
R53094 DVSS.n11078 DVSS.n10785 0.019716
R53095 DVSS.n11072 DVSS.n10790 0.019716
R53096 DVSS.n11072 DVSS.n11071 0.019716
R53097 DVSS.n11069 DVSS.n11068 0.019716
R53098 DVSS.n11068 DVSS.n10791 0.019716
R53099 DVSS.n11062 DVSS.n10796 0.019716
R53100 DVSS.n11062 DVSS.n11061 0.019716
R53101 DVSS.n11059 DVSS.n11058 0.019716
R53102 DVSS.n11058 DVSS.n10797 0.019716
R53103 DVSS.n11052 DVSS.n10802 0.019716
R53104 DVSS.n11052 DVSS.n11051 0.019716
R53105 DVSS.n11049 DVSS.n11048 0.019716
R53106 DVSS.n11048 DVSS.n10803 0.019716
R53107 DVSS.n11042 DVSS.n10808 0.019716
R53108 DVSS.n11042 DVSS.n11041 0.019716
R53109 DVSS.n11039 DVSS.n11038 0.019716
R53110 DVSS.n11038 DVSS.n10809 0.019716
R53111 DVSS.n11032 DVSS.n10814 0.019716
R53112 DVSS.n11032 DVSS.n11031 0.019716
R53113 DVSS.n11029 DVSS.n11028 0.019716
R53114 DVSS.n11028 DVSS.n10815 0.019716
R53115 DVSS.n11022 DVSS.n10820 0.019716
R53116 DVSS.n11022 DVSS.n11021 0.019716
R53117 DVSS.n11019 DVSS.n11018 0.019716
R53118 DVSS.n11018 DVSS.n10821 0.019716
R53119 DVSS.n11012 DVSS.n10826 0.019716
R53120 DVSS.n11012 DVSS.n11011 0.019716
R53121 DVSS.n11009 DVSS.n11008 0.019716
R53122 DVSS.n11008 DVSS.n10827 0.019716
R53123 DVSS.n11002 DVSS.n10832 0.019716
R53124 DVSS.n11002 DVSS.n11001 0.019716
R53125 DVSS.n10999 DVSS.n10998 0.019716
R53126 DVSS.n10998 DVSS.n10833 0.019716
R53127 DVSS.n10992 DVSS.n10838 0.019716
R53128 DVSS.n10992 DVSS.n10991 0.019716
R53129 DVSS.n10989 DVSS.n10988 0.019716
R53130 DVSS.n10988 DVSS.n10839 0.019716
R53131 DVSS.n10982 DVSS.n10844 0.019716
R53132 DVSS.n10982 DVSS.n10981 0.019716
R53133 DVSS.n10979 DVSS.n10978 0.019716
R53134 DVSS.n10978 DVSS.n10845 0.019716
R53135 DVSS.n10972 DVSS.n10850 0.019716
R53136 DVSS.n10972 DVSS.n10971 0.019716
R53137 DVSS.n10969 DVSS.n10968 0.019716
R53138 DVSS.n10968 DVSS.n10851 0.019716
R53139 DVSS.n10962 DVSS.n10856 0.019716
R53140 DVSS.n10962 DVSS.n10961 0.019716
R53141 DVSS.n10959 DVSS.n10958 0.019716
R53142 DVSS.n10958 DVSS.n10857 0.019716
R53143 DVSS.n10952 DVSS.n10862 0.019716
R53144 DVSS.n10952 DVSS.n10951 0.019716
R53145 DVSS.n10949 DVSS.n10948 0.019716
R53146 DVSS.n10948 DVSS.n10863 0.019716
R53147 DVSS.n10942 DVSS.n10868 0.019716
R53148 DVSS.n10942 DVSS.n10941 0.019716
R53149 DVSS.n10939 DVSS.n10938 0.019716
R53150 DVSS.n10938 DVSS.n10869 0.019716
R53151 DVSS.n10932 DVSS.n10874 0.019716
R53152 DVSS.n10932 DVSS.n10931 0.019716
R53153 DVSS.n10929 DVSS.n10928 0.019716
R53154 DVSS.n10928 DVSS.n10875 0.019716
R53155 DVSS.n10922 DVSS.n10880 0.019716
R53156 DVSS.n10922 DVSS.n10921 0.019716
R53157 DVSS.n10919 DVSS.n10918 0.019716
R53158 DVSS.n10918 DVSS.n10881 0.019716
R53159 DVSS.n10912 DVSS.n10886 0.019716
R53160 DVSS.n10912 DVSS.n10911 0.019716
R53161 DVSS.n10909 DVSS.n10908 0.019716
R53162 DVSS.n10908 DVSS.n10887 0.019716
R53163 DVSS.n10902 DVSS.n10892 0.019716
R53164 DVSS.n10902 DVSS.n10901 0.019716
R53165 DVSS.n10899 DVSS.n10898 0.019716
R53166 DVSS.n10898 DVSS.n10893 0.019716
R53167 DVSS.n13339 DVSS.n11154 0.019716
R53168 DVSS.n11260 DVSS.n11197 0.019716
R53169 DVSS.n11260 DVSS.n11152 0.019716
R53170 DVSS.n11269 DVSS.n11196 0.019716
R53171 DVSS.n11269 DVSS.n11151 0.019716
R53172 DVSS.n11257 DVSS.n11195 0.019716
R53173 DVSS.n11257 DVSS.n11150 0.019716
R53174 DVSS.n11278 DVSS.n11194 0.019716
R53175 DVSS.n11278 DVSS.n11149 0.019716
R53176 DVSS.n11254 DVSS.n11193 0.019716
R53177 DVSS.n11254 DVSS.n11148 0.019716
R53178 DVSS.n11287 DVSS.n11192 0.019716
R53179 DVSS.n11287 DVSS.n11147 0.019716
R53180 DVSS.n11251 DVSS.n11191 0.019716
R53181 DVSS.n11251 DVSS.n11146 0.019716
R53182 DVSS.n11296 DVSS.n11190 0.019716
R53183 DVSS.n11296 DVSS.n11145 0.019716
R53184 DVSS.n11248 DVSS.n11189 0.019716
R53185 DVSS.n11248 DVSS.n11144 0.019716
R53186 DVSS.n11305 DVSS.n11188 0.019716
R53187 DVSS.n11305 DVSS.n11143 0.019716
R53188 DVSS.n11245 DVSS.n11187 0.019716
R53189 DVSS.n11245 DVSS.n11142 0.019716
R53190 DVSS.n11314 DVSS.n11186 0.019716
R53191 DVSS.n11314 DVSS.n11141 0.019716
R53192 DVSS.n11242 DVSS.n11185 0.019716
R53193 DVSS.n11242 DVSS.n11140 0.019716
R53194 DVSS.n11323 DVSS.n11184 0.019716
R53195 DVSS.n11323 DVSS.n11139 0.019716
R53196 DVSS.n11239 DVSS.n11183 0.019716
R53197 DVSS.n11239 DVSS.n11138 0.019716
R53198 DVSS.n11332 DVSS.n11182 0.019716
R53199 DVSS.n11332 DVSS.n11137 0.019716
R53200 DVSS.n11236 DVSS.n11181 0.019716
R53201 DVSS.n11236 DVSS.n11136 0.019716
R53202 DVSS.n11341 DVSS.n11180 0.019716
R53203 DVSS.n11341 DVSS.n11135 0.019716
R53204 DVSS.n11233 DVSS.n11179 0.019716
R53205 DVSS.n11233 DVSS.n11134 0.019716
R53206 DVSS.n11350 DVSS.n11178 0.019716
R53207 DVSS.n11350 DVSS.n11133 0.019716
R53208 DVSS.n11230 DVSS.n11177 0.019716
R53209 DVSS.n11230 DVSS.n11132 0.019716
R53210 DVSS.n11359 DVSS.n11176 0.019716
R53211 DVSS.n11359 DVSS.n11131 0.019716
R53212 DVSS.n11227 DVSS.n11175 0.019716
R53213 DVSS.n11227 DVSS.n11130 0.019716
R53214 DVSS.n11368 DVSS.n11174 0.019716
R53215 DVSS.n11368 DVSS.n11129 0.019716
R53216 DVSS.n11224 DVSS.n11173 0.019716
R53217 DVSS.n11224 DVSS.n11128 0.019716
R53218 DVSS.n11377 DVSS.n11172 0.019716
R53219 DVSS.n11377 DVSS.n11127 0.019716
R53220 DVSS.n11221 DVSS.n11171 0.019716
R53221 DVSS.n11221 DVSS.n11126 0.019716
R53222 DVSS.n11386 DVSS.n11170 0.019716
R53223 DVSS.n11386 DVSS.n11125 0.019716
R53224 DVSS.n11218 DVSS.n11169 0.019716
R53225 DVSS.n11218 DVSS.n11124 0.019716
R53226 DVSS.n11395 DVSS.n11168 0.019716
R53227 DVSS.n11395 DVSS.n11123 0.019716
R53228 DVSS.n11215 DVSS.n11167 0.019716
R53229 DVSS.n11215 DVSS.n11122 0.019716
R53230 DVSS.n11404 DVSS.n11166 0.019716
R53231 DVSS.n11404 DVSS.n11121 0.019716
R53232 DVSS.n11212 DVSS.n11165 0.019716
R53233 DVSS.n11212 DVSS.n11120 0.019716
R53234 DVSS.n11413 DVSS.n11164 0.019716
R53235 DVSS.n11413 DVSS.n11119 0.019716
R53236 DVSS.n11209 DVSS.n11163 0.019716
R53237 DVSS.n11209 DVSS.n11118 0.019716
R53238 DVSS.n11422 DVSS.n11162 0.019716
R53239 DVSS.n11422 DVSS.n11117 0.019716
R53240 DVSS.n11206 DVSS.n11161 0.019716
R53241 DVSS.n11206 DVSS.n11116 0.019716
R53242 DVSS.n11431 DVSS.n11160 0.019716
R53243 DVSS.n11431 DVSS.n11115 0.019716
R53244 DVSS.n11203 DVSS.n11159 0.019716
R53245 DVSS.n11203 DVSS.n11114 0.019716
R53246 DVSS.n11440 DVSS.n11158 0.019716
R53247 DVSS.n11440 DVSS.n11113 0.019716
R53248 DVSS.n11200 DVSS.n11157 0.019716
R53249 DVSS.n11200 DVSS.n11112 0.019716
R53250 DVSS.n13325 DVSS.n11501 0.019716
R53251 DVSS.n11607 DVSS.n11545 0.019716
R53252 DVSS.n11607 DVSS.n11499 0.019716
R53253 DVSS.n13143 DVSS.n11544 0.019716
R53254 DVSS.n13143 DVSS.n11498 0.019716
R53255 DVSS.n11604 DVSS.n11543 0.019716
R53256 DVSS.n11604 DVSS.n11497 0.019716
R53257 DVSS.n13152 DVSS.n11542 0.019716
R53258 DVSS.n13152 DVSS.n11496 0.019716
R53259 DVSS.n11601 DVSS.n11541 0.019716
R53260 DVSS.n11601 DVSS.n11495 0.019716
R53261 DVSS.n13161 DVSS.n11540 0.019716
R53262 DVSS.n13161 DVSS.n11494 0.019716
R53263 DVSS.n11598 DVSS.n11539 0.019716
R53264 DVSS.n11598 DVSS.n11493 0.019716
R53265 DVSS.n13170 DVSS.n11538 0.019716
R53266 DVSS.n13170 DVSS.n11492 0.019716
R53267 DVSS.n11595 DVSS.n11537 0.019716
R53268 DVSS.n11595 DVSS.n11491 0.019716
R53269 DVSS.n13179 DVSS.n11536 0.019716
R53270 DVSS.n13179 DVSS.n11490 0.019716
R53271 DVSS.n11592 DVSS.n11535 0.019716
R53272 DVSS.n11592 DVSS.n11489 0.019716
R53273 DVSS.n13188 DVSS.n11534 0.019716
R53274 DVSS.n13188 DVSS.n11488 0.019716
R53275 DVSS.n11589 DVSS.n11533 0.019716
R53276 DVSS.n11589 DVSS.n11487 0.019716
R53277 DVSS.n13197 DVSS.n11532 0.019716
R53278 DVSS.n13197 DVSS.n11486 0.019716
R53279 DVSS.n11586 DVSS.n11531 0.019716
R53280 DVSS.n11586 DVSS.n11485 0.019716
R53281 DVSS.n13206 DVSS.n11530 0.019716
R53282 DVSS.n13206 DVSS.n11484 0.019716
R53283 DVSS.n11583 DVSS.n11529 0.019716
R53284 DVSS.n11583 DVSS.n11483 0.019716
R53285 DVSS.n13215 DVSS.n11528 0.019716
R53286 DVSS.n13215 DVSS.n11482 0.019716
R53287 DVSS.n11580 DVSS.n11527 0.019716
R53288 DVSS.n11580 DVSS.n11481 0.019716
R53289 DVSS.n13224 DVSS.n11526 0.019716
R53290 DVSS.n13224 DVSS.n11480 0.019716
R53291 DVSS.n11577 DVSS.n11525 0.019716
R53292 DVSS.n11577 DVSS.n11479 0.019716
R53293 DVSS.n13233 DVSS.n11524 0.019716
R53294 DVSS.n13233 DVSS.n11478 0.019716
R53295 DVSS.n11574 DVSS.n11523 0.019716
R53296 DVSS.n11574 DVSS.n11477 0.019716
R53297 DVSS.n13242 DVSS.n11522 0.019716
R53298 DVSS.n13242 DVSS.n11476 0.019716
R53299 DVSS.n11571 DVSS.n11521 0.019716
R53300 DVSS.n11571 DVSS.n11475 0.019716
R53301 DVSS.n13251 DVSS.n11520 0.019716
R53302 DVSS.n13251 DVSS.n11474 0.019716
R53303 DVSS.n11568 DVSS.n11519 0.019716
R53304 DVSS.n11568 DVSS.n11473 0.019716
R53305 DVSS.n13260 DVSS.n11518 0.019716
R53306 DVSS.n13260 DVSS.n11472 0.019716
R53307 DVSS.n11565 DVSS.n11517 0.019716
R53308 DVSS.n11565 DVSS.n11471 0.019716
R53309 DVSS.n13269 DVSS.n11516 0.019716
R53310 DVSS.n13269 DVSS.n11470 0.019716
R53311 DVSS.n11562 DVSS.n11515 0.019716
R53312 DVSS.n11562 DVSS.n11469 0.019716
R53313 DVSS.n13278 DVSS.n11514 0.019716
R53314 DVSS.n13278 DVSS.n11468 0.019716
R53315 DVSS.n11559 DVSS.n11513 0.019716
R53316 DVSS.n11559 DVSS.n11467 0.019716
R53317 DVSS.n13287 DVSS.n11512 0.019716
R53318 DVSS.n13287 DVSS.n11466 0.019716
R53319 DVSS.n11556 DVSS.n11511 0.019716
R53320 DVSS.n11556 DVSS.n11465 0.019716
R53321 DVSS.n13296 DVSS.n11510 0.019716
R53322 DVSS.n13296 DVSS.n11464 0.019716
R53323 DVSS.n11553 DVSS.n11509 0.019716
R53324 DVSS.n11553 DVSS.n11463 0.019716
R53325 DVSS.n13305 DVSS.n11508 0.019716
R53326 DVSS.n13305 DVSS.n11462 0.019716
R53327 DVSS.n11550 DVSS.n11507 0.019716
R53328 DVSS.n11550 DVSS.n11461 0.019716
R53329 DVSS.n13314 DVSS.n11506 0.019716
R53330 DVSS.n13314 DVSS.n11460 0.019716
R53331 DVSS.n11547 DVSS.n11505 0.019716
R53332 DVSS.n11547 DVSS.n11459 0.019716
R53333 DVSS.n11732 DVSS.n11731 0.019716
R53334 DVSS.n11737 DVSS.n11687 0.019716
R53335 DVSS.n11738 DVSS.n11737 0.019716
R53336 DVSS.n11743 DVSS.n11686 0.019716
R53337 DVSS.n11743 DVSS.n11742 0.019716
R53338 DVSS.n11749 DVSS.n11685 0.019716
R53339 DVSS.n11750 DVSS.n11749 0.019716
R53340 DVSS.n11755 DVSS.n11684 0.019716
R53341 DVSS.n11755 DVSS.n11754 0.019716
R53342 DVSS.n11761 DVSS.n11683 0.019716
R53343 DVSS.n11762 DVSS.n11761 0.019716
R53344 DVSS.n11767 DVSS.n11682 0.019716
R53345 DVSS.n11767 DVSS.n11766 0.019716
R53346 DVSS.n11773 DVSS.n11681 0.019716
R53347 DVSS.n11774 DVSS.n11773 0.019716
R53348 DVSS.n11779 DVSS.n11680 0.019716
R53349 DVSS.n11779 DVSS.n11778 0.019716
R53350 DVSS.n11785 DVSS.n11679 0.019716
R53351 DVSS.n11786 DVSS.n11785 0.019716
R53352 DVSS.n11791 DVSS.n11678 0.019716
R53353 DVSS.n11791 DVSS.n11790 0.019716
R53354 DVSS.n11797 DVSS.n11677 0.019716
R53355 DVSS.n11798 DVSS.n11797 0.019716
R53356 DVSS.n11803 DVSS.n11676 0.019716
R53357 DVSS.n11803 DVSS.n11802 0.019716
R53358 DVSS.n11809 DVSS.n11675 0.019716
R53359 DVSS.n11810 DVSS.n11809 0.019716
R53360 DVSS.n11815 DVSS.n11674 0.019716
R53361 DVSS.n11815 DVSS.n11814 0.019716
R53362 DVSS.n11821 DVSS.n11673 0.019716
R53363 DVSS.n11822 DVSS.n11821 0.019716
R53364 DVSS.n11827 DVSS.n11672 0.019716
R53365 DVSS.n11827 DVSS.n11826 0.019716
R53366 DVSS.n11833 DVSS.n11671 0.019716
R53367 DVSS.n11834 DVSS.n11833 0.019716
R53368 DVSS.n11839 DVSS.n11670 0.019716
R53369 DVSS.n11839 DVSS.n11838 0.019716
R53370 DVSS.n11845 DVSS.n11669 0.019716
R53371 DVSS.n11846 DVSS.n11845 0.019716
R53372 DVSS.n11851 DVSS.n11668 0.019716
R53373 DVSS.n11851 DVSS.n11850 0.019716
R53374 DVSS.n11857 DVSS.n11667 0.019716
R53375 DVSS.n11858 DVSS.n11857 0.019716
R53376 DVSS.n11863 DVSS.n11666 0.019716
R53377 DVSS.n11863 DVSS.n11862 0.019716
R53378 DVSS.n11869 DVSS.n11665 0.019716
R53379 DVSS.n11870 DVSS.n11869 0.019716
R53380 DVSS.n11875 DVSS.n11664 0.019716
R53381 DVSS.n11875 DVSS.n11874 0.019716
R53382 DVSS.n11881 DVSS.n11663 0.019716
R53383 DVSS.n11882 DVSS.n11881 0.019716
R53384 DVSS.n11887 DVSS.n11662 0.019716
R53385 DVSS.n11887 DVSS.n11886 0.019716
R53386 DVSS.n11893 DVSS.n11661 0.019716
R53387 DVSS.n11894 DVSS.n11893 0.019716
R53388 DVSS.n11899 DVSS.n11660 0.019716
R53389 DVSS.n11899 DVSS.n11898 0.019716
R53390 DVSS.n11905 DVSS.n11659 0.019716
R53391 DVSS.n11906 DVSS.n11905 0.019716
R53392 DVSS.n11911 DVSS.n11658 0.019716
R53393 DVSS.n11911 DVSS.n11910 0.019716
R53394 DVSS.n11917 DVSS.n11657 0.019716
R53395 DVSS.n11918 DVSS.n11917 0.019716
R53396 DVSS.n11923 DVSS.n11656 0.019716
R53397 DVSS.n11923 DVSS.n11922 0.019716
R53398 DVSS.n11929 DVSS.n11655 0.019716
R53399 DVSS.n11930 DVSS.n11929 0.019716
R53400 DVSS.n11935 DVSS.n11654 0.019716
R53401 DVSS.n11935 DVSS.n11934 0.019716
R53402 DVSS.n11941 DVSS.n11653 0.019716
R53403 DVSS.n11942 DVSS.n11941 0.019716
R53404 DVSS.n11947 DVSS.n11652 0.019716
R53405 DVSS.n11947 DVSS.n11946 0.019716
R53406 DVSS.n11953 DVSS.n11651 0.019716
R53407 DVSS.n11954 DVSS.n11953 0.019716
R53408 DVSS.n11959 DVSS.n11650 0.019716
R53409 DVSS.n11959 DVSS.n11958 0.019716
R53410 DVSS.n11965 DVSS.n11649 0.019716
R53411 DVSS.n11966 DVSS.n11965 0.019716
R53412 DVSS.n11971 DVSS.n11648 0.019716
R53413 DVSS.n11971 DVSS.n11970 0.019716
R53414 DVSS.n11976 DVSS.n11647 0.019716
R53415 DVSS.n11976 DVSS.n11689 0.019716
R53416 DVSS.n11731 DVSS.n11688 0.019716
R53417 DVSS.n11732 DVSS.n11687 0.019716
R53418 DVSS.n11739 DVSS.n11686 0.019716
R53419 DVSS.n11739 DVSS.n11738 0.019716
R53420 DVSS.n11741 DVSS.n11685 0.019716
R53421 DVSS.n11742 DVSS.n11741 0.019716
R53422 DVSS.n11751 DVSS.n11684 0.019716
R53423 DVSS.n11751 DVSS.n11750 0.019716
R53424 DVSS.n11753 DVSS.n11683 0.019716
R53425 DVSS.n11754 DVSS.n11753 0.019716
R53426 DVSS.n11763 DVSS.n11682 0.019716
R53427 DVSS.n11763 DVSS.n11762 0.019716
R53428 DVSS.n11765 DVSS.n11681 0.019716
R53429 DVSS.n11766 DVSS.n11765 0.019716
R53430 DVSS.n11775 DVSS.n11680 0.019716
R53431 DVSS.n11775 DVSS.n11774 0.019716
R53432 DVSS.n11777 DVSS.n11679 0.019716
R53433 DVSS.n11778 DVSS.n11777 0.019716
R53434 DVSS.n11787 DVSS.n11678 0.019716
R53435 DVSS.n11787 DVSS.n11786 0.019716
R53436 DVSS.n11789 DVSS.n11677 0.019716
R53437 DVSS.n11790 DVSS.n11789 0.019716
R53438 DVSS.n11799 DVSS.n11676 0.019716
R53439 DVSS.n11799 DVSS.n11798 0.019716
R53440 DVSS.n11801 DVSS.n11675 0.019716
R53441 DVSS.n11802 DVSS.n11801 0.019716
R53442 DVSS.n11811 DVSS.n11674 0.019716
R53443 DVSS.n11811 DVSS.n11810 0.019716
R53444 DVSS.n11813 DVSS.n11673 0.019716
R53445 DVSS.n11814 DVSS.n11813 0.019716
R53446 DVSS.n11823 DVSS.n11672 0.019716
R53447 DVSS.n11823 DVSS.n11822 0.019716
R53448 DVSS.n11825 DVSS.n11671 0.019716
R53449 DVSS.n11826 DVSS.n11825 0.019716
R53450 DVSS.n11835 DVSS.n11670 0.019716
R53451 DVSS.n11835 DVSS.n11834 0.019716
R53452 DVSS.n11837 DVSS.n11669 0.019716
R53453 DVSS.n11838 DVSS.n11837 0.019716
R53454 DVSS.n11847 DVSS.n11668 0.019716
R53455 DVSS.n11847 DVSS.n11846 0.019716
R53456 DVSS.n11849 DVSS.n11667 0.019716
R53457 DVSS.n11850 DVSS.n11849 0.019716
R53458 DVSS.n11859 DVSS.n11666 0.019716
R53459 DVSS.n11859 DVSS.n11858 0.019716
R53460 DVSS.n11861 DVSS.n11665 0.019716
R53461 DVSS.n11862 DVSS.n11861 0.019716
R53462 DVSS.n11871 DVSS.n11664 0.019716
R53463 DVSS.n11871 DVSS.n11870 0.019716
R53464 DVSS.n11873 DVSS.n11663 0.019716
R53465 DVSS.n11874 DVSS.n11873 0.019716
R53466 DVSS.n11883 DVSS.n11662 0.019716
R53467 DVSS.n11883 DVSS.n11882 0.019716
R53468 DVSS.n11885 DVSS.n11661 0.019716
R53469 DVSS.n11886 DVSS.n11885 0.019716
R53470 DVSS.n11895 DVSS.n11660 0.019716
R53471 DVSS.n11895 DVSS.n11894 0.019716
R53472 DVSS.n11897 DVSS.n11659 0.019716
R53473 DVSS.n11898 DVSS.n11897 0.019716
R53474 DVSS.n11907 DVSS.n11658 0.019716
R53475 DVSS.n11907 DVSS.n11906 0.019716
R53476 DVSS.n11909 DVSS.n11657 0.019716
R53477 DVSS.n11910 DVSS.n11909 0.019716
R53478 DVSS.n11919 DVSS.n11656 0.019716
R53479 DVSS.n11919 DVSS.n11918 0.019716
R53480 DVSS.n11921 DVSS.n11655 0.019716
R53481 DVSS.n11922 DVSS.n11921 0.019716
R53482 DVSS.n11931 DVSS.n11654 0.019716
R53483 DVSS.n11931 DVSS.n11930 0.019716
R53484 DVSS.n11933 DVSS.n11653 0.019716
R53485 DVSS.n11934 DVSS.n11933 0.019716
R53486 DVSS.n11943 DVSS.n11652 0.019716
R53487 DVSS.n11943 DVSS.n11942 0.019716
R53488 DVSS.n11945 DVSS.n11651 0.019716
R53489 DVSS.n11946 DVSS.n11945 0.019716
R53490 DVSS.n11955 DVSS.n11650 0.019716
R53491 DVSS.n11955 DVSS.n11954 0.019716
R53492 DVSS.n11957 DVSS.n11649 0.019716
R53493 DVSS.n11958 DVSS.n11957 0.019716
R53494 DVSS.n11967 DVSS.n11648 0.019716
R53495 DVSS.n11967 DVSS.n11966 0.019716
R53496 DVSS.n11969 DVSS.n11647 0.019716
R53497 DVSS.n11970 DVSS.n11969 0.019716
R53498 DVSS.n11979 DVSS.n11689 0.019716
R53499 DVSS.n13325 DVSS.n13324 0.019716
R53500 DVSS.n11545 DVSS.n11501 0.019716
R53501 DVSS.n13141 DVSS.n11544 0.019716
R53502 DVSS.n13141 DVSS.n11499 0.019716
R53503 DVSS.n13145 DVSS.n11543 0.019716
R53504 DVSS.n13145 DVSS.n11498 0.019716
R53505 DVSS.n13150 DVSS.n11542 0.019716
R53506 DVSS.n13150 DVSS.n11497 0.019716
R53507 DVSS.n13154 DVSS.n11541 0.019716
R53508 DVSS.n13154 DVSS.n11496 0.019716
R53509 DVSS.n13159 DVSS.n11540 0.019716
R53510 DVSS.n13159 DVSS.n11495 0.019716
R53511 DVSS.n13163 DVSS.n11539 0.019716
R53512 DVSS.n13163 DVSS.n11494 0.019716
R53513 DVSS.n13168 DVSS.n11538 0.019716
R53514 DVSS.n13168 DVSS.n11493 0.019716
R53515 DVSS.n13172 DVSS.n11537 0.019716
R53516 DVSS.n13172 DVSS.n11492 0.019716
R53517 DVSS.n13177 DVSS.n11536 0.019716
R53518 DVSS.n13177 DVSS.n11491 0.019716
R53519 DVSS.n13181 DVSS.n11535 0.019716
R53520 DVSS.n13181 DVSS.n11490 0.019716
R53521 DVSS.n13186 DVSS.n11534 0.019716
R53522 DVSS.n13186 DVSS.n11489 0.019716
R53523 DVSS.n13190 DVSS.n11533 0.019716
R53524 DVSS.n13190 DVSS.n11488 0.019716
R53525 DVSS.n13195 DVSS.n11532 0.019716
R53526 DVSS.n13195 DVSS.n11487 0.019716
R53527 DVSS.n13199 DVSS.n11531 0.019716
R53528 DVSS.n13199 DVSS.n11486 0.019716
R53529 DVSS.n13204 DVSS.n11530 0.019716
R53530 DVSS.n13204 DVSS.n11485 0.019716
R53531 DVSS.n13208 DVSS.n11529 0.019716
R53532 DVSS.n13208 DVSS.n11484 0.019716
R53533 DVSS.n13213 DVSS.n11528 0.019716
R53534 DVSS.n13213 DVSS.n11483 0.019716
R53535 DVSS.n13217 DVSS.n11527 0.019716
R53536 DVSS.n13217 DVSS.n11482 0.019716
R53537 DVSS.n13222 DVSS.n11526 0.019716
R53538 DVSS.n13222 DVSS.n11481 0.019716
R53539 DVSS.n13226 DVSS.n11525 0.019716
R53540 DVSS.n13226 DVSS.n11480 0.019716
R53541 DVSS.n13231 DVSS.n11524 0.019716
R53542 DVSS.n13231 DVSS.n11479 0.019716
R53543 DVSS.n13235 DVSS.n11523 0.019716
R53544 DVSS.n13235 DVSS.n11478 0.019716
R53545 DVSS.n13240 DVSS.n11522 0.019716
R53546 DVSS.n13240 DVSS.n11477 0.019716
R53547 DVSS.n13244 DVSS.n11521 0.019716
R53548 DVSS.n13244 DVSS.n11476 0.019716
R53549 DVSS.n13249 DVSS.n11520 0.019716
R53550 DVSS.n13249 DVSS.n11475 0.019716
R53551 DVSS.n13253 DVSS.n11519 0.019716
R53552 DVSS.n13253 DVSS.n11474 0.019716
R53553 DVSS.n13258 DVSS.n11518 0.019716
R53554 DVSS.n13258 DVSS.n11473 0.019716
R53555 DVSS.n13262 DVSS.n11517 0.019716
R53556 DVSS.n13262 DVSS.n11472 0.019716
R53557 DVSS.n13267 DVSS.n11516 0.019716
R53558 DVSS.n13267 DVSS.n11471 0.019716
R53559 DVSS.n13271 DVSS.n11515 0.019716
R53560 DVSS.n13271 DVSS.n11470 0.019716
R53561 DVSS.n13276 DVSS.n11514 0.019716
R53562 DVSS.n13276 DVSS.n11469 0.019716
R53563 DVSS.n13280 DVSS.n11513 0.019716
R53564 DVSS.n13280 DVSS.n11468 0.019716
R53565 DVSS.n13285 DVSS.n11512 0.019716
R53566 DVSS.n13285 DVSS.n11467 0.019716
R53567 DVSS.n13289 DVSS.n11511 0.019716
R53568 DVSS.n13289 DVSS.n11466 0.019716
R53569 DVSS.n13294 DVSS.n11510 0.019716
R53570 DVSS.n13294 DVSS.n11465 0.019716
R53571 DVSS.n13298 DVSS.n11509 0.019716
R53572 DVSS.n13298 DVSS.n11464 0.019716
R53573 DVSS.n13303 DVSS.n11508 0.019716
R53574 DVSS.n13303 DVSS.n11463 0.019716
R53575 DVSS.n13307 DVSS.n11507 0.019716
R53576 DVSS.n13307 DVSS.n11462 0.019716
R53577 DVSS.n13312 DVSS.n11506 0.019716
R53578 DVSS.n13312 DVSS.n11461 0.019716
R53579 DVSS.n13316 DVSS.n11505 0.019716
R53580 DVSS.n13316 DVSS.n11460 0.019716
R53581 DVSS.n13322 DVSS.n11459 0.019716
R53582 DVSS.n13339 DVSS.n13338 0.019716
R53583 DVSS.n11197 DVSS.n11154 0.019716
R53584 DVSS.n11267 DVSS.n11196 0.019716
R53585 DVSS.n11267 DVSS.n11152 0.019716
R53586 DVSS.n11271 DVSS.n11195 0.019716
R53587 DVSS.n11271 DVSS.n11151 0.019716
R53588 DVSS.n11276 DVSS.n11194 0.019716
R53589 DVSS.n11276 DVSS.n11150 0.019716
R53590 DVSS.n11280 DVSS.n11193 0.019716
R53591 DVSS.n11280 DVSS.n11149 0.019716
R53592 DVSS.n11285 DVSS.n11192 0.019716
R53593 DVSS.n11285 DVSS.n11148 0.019716
R53594 DVSS.n11289 DVSS.n11191 0.019716
R53595 DVSS.n11289 DVSS.n11147 0.019716
R53596 DVSS.n11294 DVSS.n11190 0.019716
R53597 DVSS.n11294 DVSS.n11146 0.019716
R53598 DVSS.n11298 DVSS.n11189 0.019716
R53599 DVSS.n11298 DVSS.n11145 0.019716
R53600 DVSS.n11303 DVSS.n11188 0.019716
R53601 DVSS.n11303 DVSS.n11144 0.019716
R53602 DVSS.n11307 DVSS.n11187 0.019716
R53603 DVSS.n11307 DVSS.n11143 0.019716
R53604 DVSS.n11312 DVSS.n11186 0.019716
R53605 DVSS.n11312 DVSS.n11142 0.019716
R53606 DVSS.n11316 DVSS.n11185 0.019716
R53607 DVSS.n11316 DVSS.n11141 0.019716
R53608 DVSS.n11321 DVSS.n11184 0.019716
R53609 DVSS.n11321 DVSS.n11140 0.019716
R53610 DVSS.n11325 DVSS.n11183 0.019716
R53611 DVSS.n11325 DVSS.n11139 0.019716
R53612 DVSS.n11330 DVSS.n11182 0.019716
R53613 DVSS.n11330 DVSS.n11138 0.019716
R53614 DVSS.n11334 DVSS.n11181 0.019716
R53615 DVSS.n11334 DVSS.n11137 0.019716
R53616 DVSS.n11339 DVSS.n11180 0.019716
R53617 DVSS.n11339 DVSS.n11136 0.019716
R53618 DVSS.n11343 DVSS.n11179 0.019716
R53619 DVSS.n11343 DVSS.n11135 0.019716
R53620 DVSS.n11348 DVSS.n11178 0.019716
R53621 DVSS.n11348 DVSS.n11134 0.019716
R53622 DVSS.n11352 DVSS.n11177 0.019716
R53623 DVSS.n11352 DVSS.n11133 0.019716
R53624 DVSS.n11357 DVSS.n11176 0.019716
R53625 DVSS.n11357 DVSS.n11132 0.019716
R53626 DVSS.n11361 DVSS.n11175 0.019716
R53627 DVSS.n11361 DVSS.n11131 0.019716
R53628 DVSS.n11366 DVSS.n11174 0.019716
R53629 DVSS.n11366 DVSS.n11130 0.019716
R53630 DVSS.n11370 DVSS.n11173 0.019716
R53631 DVSS.n11370 DVSS.n11129 0.019716
R53632 DVSS.n11375 DVSS.n11172 0.019716
R53633 DVSS.n11375 DVSS.n11128 0.019716
R53634 DVSS.n11379 DVSS.n11171 0.019716
R53635 DVSS.n11379 DVSS.n11127 0.019716
R53636 DVSS.n11384 DVSS.n11170 0.019716
R53637 DVSS.n11384 DVSS.n11126 0.019716
R53638 DVSS.n11388 DVSS.n11169 0.019716
R53639 DVSS.n11388 DVSS.n11125 0.019716
R53640 DVSS.n11393 DVSS.n11168 0.019716
R53641 DVSS.n11393 DVSS.n11124 0.019716
R53642 DVSS.n11397 DVSS.n11167 0.019716
R53643 DVSS.n11397 DVSS.n11123 0.019716
R53644 DVSS.n11402 DVSS.n11166 0.019716
R53645 DVSS.n11402 DVSS.n11122 0.019716
R53646 DVSS.n11406 DVSS.n11165 0.019716
R53647 DVSS.n11406 DVSS.n11121 0.019716
R53648 DVSS.n11411 DVSS.n11164 0.019716
R53649 DVSS.n11411 DVSS.n11120 0.019716
R53650 DVSS.n11415 DVSS.n11163 0.019716
R53651 DVSS.n11415 DVSS.n11119 0.019716
R53652 DVSS.n11420 DVSS.n11162 0.019716
R53653 DVSS.n11420 DVSS.n11118 0.019716
R53654 DVSS.n11424 DVSS.n11161 0.019716
R53655 DVSS.n11424 DVSS.n11117 0.019716
R53656 DVSS.n11429 DVSS.n11160 0.019716
R53657 DVSS.n11429 DVSS.n11116 0.019716
R53658 DVSS.n11433 DVSS.n11159 0.019716
R53659 DVSS.n11433 DVSS.n11115 0.019716
R53660 DVSS.n11438 DVSS.n11158 0.019716
R53661 DVSS.n11438 DVSS.n11114 0.019716
R53662 DVSS.n11442 DVSS.n11157 0.019716
R53663 DVSS.n11442 DVSS.n11113 0.019716
R53664 DVSS.n13336 DVSS.n11112 0.019716
R53665 DVSS.n11102 DVSS.n11101 0.019716
R53666 DVSS.n11100 DVSS.n11099 0.019716
R53667 DVSS.n10778 DVSS.n10777 0.019716
R53668 DVSS.n10777 DVSS.n10773 0.019716
R53669 DVSS.n11090 DVSS.n11089 0.019716
R53670 DVSS.n11091 DVSS.n11090 0.019716
R53671 DVSS.n10784 DVSS.n10783 0.019716
R53672 DVSS.n10783 DVSS.n10779 0.019716
R53673 DVSS.n11080 DVSS.n11079 0.019716
R53674 DVSS.n11081 DVSS.n11080 0.019716
R53675 DVSS.n10790 DVSS.n10789 0.019716
R53676 DVSS.n10789 DVSS.n10785 0.019716
R53677 DVSS.n11070 DVSS.n11069 0.019716
R53678 DVSS.n11071 DVSS.n11070 0.019716
R53679 DVSS.n10796 DVSS.n10795 0.019716
R53680 DVSS.n10795 DVSS.n10791 0.019716
R53681 DVSS.n11060 DVSS.n11059 0.019716
R53682 DVSS.n11061 DVSS.n11060 0.019716
R53683 DVSS.n10802 DVSS.n10801 0.019716
R53684 DVSS.n10801 DVSS.n10797 0.019716
R53685 DVSS.n11050 DVSS.n11049 0.019716
R53686 DVSS.n11051 DVSS.n11050 0.019716
R53687 DVSS.n10808 DVSS.n10807 0.019716
R53688 DVSS.n10807 DVSS.n10803 0.019716
R53689 DVSS.n11040 DVSS.n11039 0.019716
R53690 DVSS.n11041 DVSS.n11040 0.019716
R53691 DVSS.n10814 DVSS.n10813 0.019716
R53692 DVSS.n10813 DVSS.n10809 0.019716
R53693 DVSS.n11030 DVSS.n11029 0.019716
R53694 DVSS.n11031 DVSS.n11030 0.019716
R53695 DVSS.n10820 DVSS.n10819 0.019716
R53696 DVSS.n10819 DVSS.n10815 0.019716
R53697 DVSS.n11020 DVSS.n11019 0.019716
R53698 DVSS.n11021 DVSS.n11020 0.019716
R53699 DVSS.n10826 DVSS.n10825 0.019716
R53700 DVSS.n10825 DVSS.n10821 0.019716
R53701 DVSS.n11010 DVSS.n11009 0.019716
R53702 DVSS.n11011 DVSS.n11010 0.019716
R53703 DVSS.n10832 DVSS.n10831 0.019716
R53704 DVSS.n10831 DVSS.n10827 0.019716
R53705 DVSS.n11000 DVSS.n10999 0.019716
R53706 DVSS.n11001 DVSS.n11000 0.019716
R53707 DVSS.n10838 DVSS.n10837 0.019716
R53708 DVSS.n10837 DVSS.n10833 0.019716
R53709 DVSS.n10990 DVSS.n10989 0.019716
R53710 DVSS.n10991 DVSS.n10990 0.019716
R53711 DVSS.n10844 DVSS.n10843 0.019716
R53712 DVSS.n10843 DVSS.n10839 0.019716
R53713 DVSS.n10980 DVSS.n10979 0.019716
R53714 DVSS.n10981 DVSS.n10980 0.019716
R53715 DVSS.n10850 DVSS.n10849 0.019716
R53716 DVSS.n10849 DVSS.n10845 0.019716
R53717 DVSS.n10970 DVSS.n10969 0.019716
R53718 DVSS.n10971 DVSS.n10970 0.019716
R53719 DVSS.n10856 DVSS.n10855 0.019716
R53720 DVSS.n10855 DVSS.n10851 0.019716
R53721 DVSS.n10960 DVSS.n10959 0.019716
R53722 DVSS.n10961 DVSS.n10960 0.019716
R53723 DVSS.n10862 DVSS.n10861 0.019716
R53724 DVSS.n10861 DVSS.n10857 0.019716
R53725 DVSS.n10950 DVSS.n10949 0.019716
R53726 DVSS.n10951 DVSS.n10950 0.019716
R53727 DVSS.n10868 DVSS.n10867 0.019716
R53728 DVSS.n10867 DVSS.n10863 0.019716
R53729 DVSS.n10940 DVSS.n10939 0.019716
R53730 DVSS.n10941 DVSS.n10940 0.019716
R53731 DVSS.n10874 DVSS.n10873 0.019716
R53732 DVSS.n10873 DVSS.n10869 0.019716
R53733 DVSS.n10930 DVSS.n10929 0.019716
R53734 DVSS.n10931 DVSS.n10930 0.019716
R53735 DVSS.n10880 DVSS.n10879 0.019716
R53736 DVSS.n10879 DVSS.n10875 0.019716
R53737 DVSS.n10920 DVSS.n10919 0.019716
R53738 DVSS.n10921 DVSS.n10920 0.019716
R53739 DVSS.n10886 DVSS.n10885 0.019716
R53740 DVSS.n10885 DVSS.n10881 0.019716
R53741 DVSS.n10910 DVSS.n10909 0.019716
R53742 DVSS.n10911 DVSS.n10910 0.019716
R53743 DVSS.n10892 DVSS.n10891 0.019716
R53744 DVSS.n10891 DVSS.n10887 0.019716
R53745 DVSS.n10900 DVSS.n10899 0.019716
R53746 DVSS.n10901 DVSS.n10900 0.019716
R53747 DVSS.n10894 DVSS.n10893 0.019716
R53748 DVSS.n1609 DVSS.n1565 0.019716
R53749 DVSS.n1610 DVSS.n1564 0.019716
R53750 DVSS.n10513 DVSS.n1563 0.019716
R53751 DVSS.n10513 DVSS.n10512 0.019716
R53752 DVSS.n10515 DVSS.n1562 0.019716
R53753 DVSS.n10516 DVSS.n10515 0.019716
R53754 DVSS.n10525 DVSS.n1561 0.019716
R53755 DVSS.n10525 DVSS.n10524 0.019716
R53756 DVSS.n10527 DVSS.n1560 0.019716
R53757 DVSS.n10528 DVSS.n10527 0.019716
R53758 DVSS.n10537 DVSS.n1559 0.019716
R53759 DVSS.n10537 DVSS.n10536 0.019716
R53760 DVSS.n10539 DVSS.n1558 0.019716
R53761 DVSS.n10540 DVSS.n10539 0.019716
R53762 DVSS.n10549 DVSS.n1557 0.019716
R53763 DVSS.n10549 DVSS.n10548 0.019716
R53764 DVSS.n10551 DVSS.n1556 0.019716
R53765 DVSS.n10552 DVSS.n10551 0.019716
R53766 DVSS.n10561 DVSS.n1555 0.019716
R53767 DVSS.n10561 DVSS.n10560 0.019716
R53768 DVSS.n10563 DVSS.n1554 0.019716
R53769 DVSS.n10564 DVSS.n10563 0.019716
R53770 DVSS.n10573 DVSS.n1553 0.019716
R53771 DVSS.n10573 DVSS.n10572 0.019716
R53772 DVSS.n10575 DVSS.n1552 0.019716
R53773 DVSS.n10576 DVSS.n10575 0.019716
R53774 DVSS.n10585 DVSS.n1551 0.019716
R53775 DVSS.n10585 DVSS.n10584 0.019716
R53776 DVSS.n10587 DVSS.n1550 0.019716
R53777 DVSS.n10588 DVSS.n10587 0.019716
R53778 DVSS.n10597 DVSS.n1549 0.019716
R53779 DVSS.n10597 DVSS.n10596 0.019716
R53780 DVSS.n10599 DVSS.n1548 0.019716
R53781 DVSS.n10600 DVSS.n10599 0.019716
R53782 DVSS.n10609 DVSS.n1547 0.019716
R53783 DVSS.n10609 DVSS.n10608 0.019716
R53784 DVSS.n10611 DVSS.n1546 0.019716
R53785 DVSS.n10612 DVSS.n10611 0.019716
R53786 DVSS.n10621 DVSS.n1545 0.019716
R53787 DVSS.n10621 DVSS.n10620 0.019716
R53788 DVSS.n10623 DVSS.n1544 0.019716
R53789 DVSS.n10624 DVSS.n10623 0.019716
R53790 DVSS.n10633 DVSS.n1543 0.019716
R53791 DVSS.n10633 DVSS.n10632 0.019716
R53792 DVSS.n10635 DVSS.n1542 0.019716
R53793 DVSS.n10636 DVSS.n10635 0.019716
R53794 DVSS.n10645 DVSS.n1541 0.019716
R53795 DVSS.n10645 DVSS.n10644 0.019716
R53796 DVSS.n10647 DVSS.n1540 0.019716
R53797 DVSS.n10648 DVSS.n10647 0.019716
R53798 DVSS.n10657 DVSS.n1539 0.019716
R53799 DVSS.n10657 DVSS.n10656 0.019716
R53800 DVSS.n10659 DVSS.n1538 0.019716
R53801 DVSS.n10660 DVSS.n10659 0.019716
R53802 DVSS.n10669 DVSS.n1537 0.019716
R53803 DVSS.n10669 DVSS.n10668 0.019716
R53804 DVSS.n10671 DVSS.n1536 0.019716
R53805 DVSS.n10672 DVSS.n10671 0.019716
R53806 DVSS.n10681 DVSS.n1535 0.019716
R53807 DVSS.n10681 DVSS.n10680 0.019716
R53808 DVSS.n10683 DVSS.n1534 0.019716
R53809 DVSS.n10684 DVSS.n10683 0.019716
R53810 DVSS.n10693 DVSS.n1533 0.019716
R53811 DVSS.n10693 DVSS.n10692 0.019716
R53812 DVSS.n10695 DVSS.n1532 0.019716
R53813 DVSS.n10696 DVSS.n10695 0.019716
R53814 DVSS.n10705 DVSS.n1531 0.019716
R53815 DVSS.n10705 DVSS.n10704 0.019716
R53816 DVSS.n10707 DVSS.n1530 0.019716
R53817 DVSS.n10708 DVSS.n10707 0.019716
R53818 DVSS.n10717 DVSS.n1529 0.019716
R53819 DVSS.n10717 DVSS.n10716 0.019716
R53820 DVSS.n10719 DVSS.n1528 0.019716
R53821 DVSS.n10720 DVSS.n10719 0.019716
R53822 DVSS.n10729 DVSS.n1527 0.019716
R53823 DVSS.n10729 DVSS.n10728 0.019716
R53824 DVSS.n10731 DVSS.n1526 0.019716
R53825 DVSS.n10732 DVSS.n10731 0.019716
R53826 DVSS.n10741 DVSS.n1525 0.019716
R53827 DVSS.n10741 DVSS.n10740 0.019716
R53828 DVSS.n10743 DVSS.n1524 0.019716
R53829 DVSS.n10744 DVSS.n10743 0.019716
R53830 DVSS.n10753 DVSS.n10752 0.019716
R53831 DVSS.n1960 DVSS.n1959 0.019716
R53832 DVSS.n1670 DVSS.n1668 0.019716
R53833 DVSS.n1952 DVSS.n1951 0.019716
R53834 DVSS.n1952 DVSS.n1667 0.019716
R53835 DVSS.n1947 DVSS.n1946 0.019716
R53836 DVSS.n1947 DVSS.n1666 0.019716
R53837 DVSS.n1940 DVSS.n1939 0.019716
R53838 DVSS.n1940 DVSS.n1665 0.019716
R53839 DVSS.n1935 DVSS.n1934 0.019716
R53840 DVSS.n1935 DVSS.n1664 0.019716
R53841 DVSS.n1928 DVSS.n1927 0.019716
R53842 DVSS.n1928 DVSS.n1663 0.019716
R53843 DVSS.n1923 DVSS.n1922 0.019716
R53844 DVSS.n1923 DVSS.n1662 0.019716
R53845 DVSS.n1916 DVSS.n1915 0.019716
R53846 DVSS.n1916 DVSS.n1661 0.019716
R53847 DVSS.n1911 DVSS.n1910 0.019716
R53848 DVSS.n1911 DVSS.n1660 0.019716
R53849 DVSS.n1904 DVSS.n1903 0.019716
R53850 DVSS.n1904 DVSS.n1659 0.019716
R53851 DVSS.n1899 DVSS.n1898 0.019716
R53852 DVSS.n1899 DVSS.n1658 0.019716
R53853 DVSS.n1892 DVSS.n1891 0.019716
R53854 DVSS.n1892 DVSS.n1657 0.019716
R53855 DVSS.n1887 DVSS.n1886 0.019716
R53856 DVSS.n1887 DVSS.n1656 0.019716
R53857 DVSS.n1880 DVSS.n1879 0.019716
R53858 DVSS.n1880 DVSS.n1655 0.019716
R53859 DVSS.n1875 DVSS.n1874 0.019716
R53860 DVSS.n1875 DVSS.n1654 0.019716
R53861 DVSS.n1868 DVSS.n1867 0.019716
R53862 DVSS.n1868 DVSS.n1653 0.019716
R53863 DVSS.n1863 DVSS.n1862 0.019716
R53864 DVSS.n1863 DVSS.n1652 0.019716
R53865 DVSS.n1856 DVSS.n1855 0.019716
R53866 DVSS.n1856 DVSS.n1651 0.019716
R53867 DVSS.n1851 DVSS.n1850 0.019716
R53868 DVSS.n1851 DVSS.n1650 0.019716
R53869 DVSS.n1844 DVSS.n1843 0.019716
R53870 DVSS.n1844 DVSS.n1649 0.019716
R53871 DVSS.n1839 DVSS.n1838 0.019716
R53872 DVSS.n1839 DVSS.n1648 0.019716
R53873 DVSS.n1832 DVSS.n1831 0.019716
R53874 DVSS.n1832 DVSS.n1647 0.019716
R53875 DVSS.n1827 DVSS.n1826 0.019716
R53876 DVSS.n1827 DVSS.n1646 0.019716
R53877 DVSS.n1820 DVSS.n1819 0.019716
R53878 DVSS.n1820 DVSS.n1645 0.019716
R53879 DVSS.n1815 DVSS.n1814 0.019716
R53880 DVSS.n1815 DVSS.n1644 0.019716
R53881 DVSS.n1808 DVSS.n1807 0.019716
R53882 DVSS.n1808 DVSS.n1643 0.019716
R53883 DVSS.n1803 DVSS.n1802 0.019716
R53884 DVSS.n1803 DVSS.n1642 0.019716
R53885 DVSS.n1796 DVSS.n1795 0.019716
R53886 DVSS.n1796 DVSS.n1641 0.019716
R53887 DVSS.n1791 DVSS.n1790 0.019716
R53888 DVSS.n1791 DVSS.n1640 0.019716
R53889 DVSS.n1784 DVSS.n1783 0.019716
R53890 DVSS.n1784 DVSS.n1639 0.019716
R53891 DVSS.n1779 DVSS.n1778 0.019716
R53892 DVSS.n1779 DVSS.n1638 0.019716
R53893 DVSS.n1772 DVSS.n1771 0.019716
R53894 DVSS.n1772 DVSS.n1637 0.019716
R53895 DVSS.n1767 DVSS.n1766 0.019716
R53896 DVSS.n1767 DVSS.n1636 0.019716
R53897 DVSS.n1760 DVSS.n1759 0.019716
R53898 DVSS.n1760 DVSS.n1635 0.019716
R53899 DVSS.n1755 DVSS.n1754 0.019716
R53900 DVSS.n1755 DVSS.n1634 0.019716
R53901 DVSS.n1748 DVSS.n1747 0.019716
R53902 DVSS.n1748 DVSS.n1633 0.019716
R53903 DVSS.n1743 DVSS.n1742 0.019716
R53904 DVSS.n1743 DVSS.n1632 0.019716
R53905 DVSS.n1736 DVSS.n1735 0.019716
R53906 DVSS.n1736 DVSS.n1631 0.019716
R53907 DVSS.n1731 DVSS.n1730 0.019716
R53908 DVSS.n1731 DVSS.n1630 0.019716
R53909 DVSS.n1724 DVSS.n1723 0.019716
R53910 DVSS.n1724 DVSS.n1629 0.019716
R53911 DVSS.n1719 DVSS.n1718 0.019716
R53912 DVSS.n1719 DVSS.n1628 0.019716
R53913 DVSS.n1712 DVSS.n1627 0.019716
R53914 DVSS.n10451 DVSS.n2009 0.019716
R53915 DVSS.n10452 DVSS.n2008 0.019716
R53916 DVSS.n10447 DVSS.n2007 0.019716
R53917 DVSS.n10448 DVSS.n10447 0.019716
R53918 DVSS.n10440 DVSS.n2006 0.019716
R53919 DVSS.n10441 DVSS.n10440 0.019716
R53920 DVSS.n10435 DVSS.n2005 0.019716
R53921 DVSS.n10436 DVSS.n10435 0.019716
R53922 DVSS.n10428 DVSS.n2004 0.019716
R53923 DVSS.n10429 DVSS.n10428 0.019716
R53924 DVSS.n10423 DVSS.n2003 0.019716
R53925 DVSS.n10424 DVSS.n10423 0.019716
R53926 DVSS.n10416 DVSS.n2002 0.019716
R53927 DVSS.n10417 DVSS.n10416 0.019716
R53928 DVSS.n10411 DVSS.n2001 0.019716
R53929 DVSS.n10412 DVSS.n10411 0.019716
R53930 DVSS.n10404 DVSS.n2000 0.019716
R53931 DVSS.n10405 DVSS.n10404 0.019716
R53932 DVSS.n10399 DVSS.n1999 0.019716
R53933 DVSS.n10400 DVSS.n10399 0.019716
R53934 DVSS.n10392 DVSS.n1998 0.019716
R53935 DVSS.n10393 DVSS.n10392 0.019716
R53936 DVSS.n10387 DVSS.n1997 0.019716
R53937 DVSS.n10388 DVSS.n10387 0.019716
R53938 DVSS.n10380 DVSS.n1996 0.019716
R53939 DVSS.n10381 DVSS.n10380 0.019716
R53940 DVSS.n10375 DVSS.n1995 0.019716
R53941 DVSS.n10376 DVSS.n10375 0.019716
R53942 DVSS.n10368 DVSS.n1994 0.019716
R53943 DVSS.n10369 DVSS.n10368 0.019716
R53944 DVSS.n10363 DVSS.n1993 0.019716
R53945 DVSS.n10364 DVSS.n10363 0.019716
R53946 DVSS.n10356 DVSS.n1992 0.019716
R53947 DVSS.n10357 DVSS.n10356 0.019716
R53948 DVSS.n10351 DVSS.n1991 0.019716
R53949 DVSS.n10352 DVSS.n10351 0.019716
R53950 DVSS.n10344 DVSS.n1990 0.019716
R53951 DVSS.n10345 DVSS.n10344 0.019716
R53952 DVSS.n10339 DVSS.n1989 0.019716
R53953 DVSS.n10340 DVSS.n10339 0.019716
R53954 DVSS.n10332 DVSS.n1988 0.019716
R53955 DVSS.n10333 DVSS.n10332 0.019716
R53956 DVSS.n10327 DVSS.n1987 0.019716
R53957 DVSS.n10328 DVSS.n10327 0.019716
R53958 DVSS.n10320 DVSS.n1986 0.019716
R53959 DVSS.n10321 DVSS.n10320 0.019716
R53960 DVSS.n10315 DVSS.n1985 0.019716
R53961 DVSS.n10316 DVSS.n10315 0.019716
R53962 DVSS.n10308 DVSS.n1984 0.019716
R53963 DVSS.n10309 DVSS.n10308 0.019716
R53964 DVSS.n10303 DVSS.n1983 0.019716
R53965 DVSS.n10304 DVSS.n10303 0.019716
R53966 DVSS.n10296 DVSS.n1982 0.019716
R53967 DVSS.n10297 DVSS.n10296 0.019716
R53968 DVSS.n10291 DVSS.n1981 0.019716
R53969 DVSS.n10292 DVSS.n10291 0.019716
R53970 DVSS.n10284 DVSS.n1980 0.019716
R53971 DVSS.n10285 DVSS.n10284 0.019716
R53972 DVSS.n10279 DVSS.n1979 0.019716
R53973 DVSS.n10280 DVSS.n10279 0.019716
R53974 DVSS.n10272 DVSS.n1978 0.019716
R53975 DVSS.n10273 DVSS.n10272 0.019716
R53976 DVSS.n10267 DVSS.n1977 0.019716
R53977 DVSS.n10268 DVSS.n10267 0.019716
R53978 DVSS.n10260 DVSS.n1976 0.019716
R53979 DVSS.n10261 DVSS.n10260 0.019716
R53980 DVSS.n10255 DVSS.n1975 0.019716
R53981 DVSS.n10256 DVSS.n10255 0.019716
R53982 DVSS.n10248 DVSS.n1974 0.019716
R53983 DVSS.n10249 DVSS.n10248 0.019716
R53984 DVSS.n10243 DVSS.n1973 0.019716
R53985 DVSS.n10244 DVSS.n10243 0.019716
R53986 DVSS.n10236 DVSS.n1972 0.019716
R53987 DVSS.n10237 DVSS.n10236 0.019716
R53988 DVSS.n10231 DVSS.n1971 0.019716
R53989 DVSS.n10232 DVSS.n10231 0.019716
R53990 DVSS.n10224 DVSS.n1970 0.019716
R53991 DVSS.n10225 DVSS.n10224 0.019716
R53992 DVSS.n10219 DVSS.n1969 0.019716
R53993 DVSS.n10220 DVSS.n10219 0.019716
R53994 DVSS.n10212 DVSS.n1968 0.019716
R53995 DVSS.n10213 DVSS.n10212 0.019716
R53996 DVSS.n10474 DVSS.n10473 0.019716
R53997 DVSS.n2114 DVSS.n2069 0.019716
R53998 DVSS.n2115 DVSS.n2068 0.019716
R53999 DVSS.n2124 DVSS.n2067 0.019716
R54000 DVSS.n2124 DVSS.n2123 0.019716
R54001 DVSS.n2126 DVSS.n2066 0.019716
R54002 DVSS.n2127 DVSS.n2126 0.019716
R54003 DVSS.n2136 DVSS.n2065 0.019716
R54004 DVSS.n2136 DVSS.n2135 0.019716
R54005 DVSS.n2138 DVSS.n2064 0.019716
R54006 DVSS.n2139 DVSS.n2138 0.019716
R54007 DVSS.n2148 DVSS.n2063 0.019716
R54008 DVSS.n2148 DVSS.n2147 0.019716
R54009 DVSS.n2150 DVSS.n2062 0.019716
R54010 DVSS.n2151 DVSS.n2150 0.019716
R54011 DVSS.n2160 DVSS.n2061 0.019716
R54012 DVSS.n2160 DVSS.n2159 0.019716
R54013 DVSS.n2162 DVSS.n2060 0.019716
R54014 DVSS.n2163 DVSS.n2162 0.019716
R54015 DVSS.n2172 DVSS.n2059 0.019716
R54016 DVSS.n2172 DVSS.n2171 0.019716
R54017 DVSS.n2174 DVSS.n2058 0.019716
R54018 DVSS.n2175 DVSS.n2174 0.019716
R54019 DVSS.n2184 DVSS.n2057 0.019716
R54020 DVSS.n2184 DVSS.n2183 0.019716
R54021 DVSS.n2186 DVSS.n2056 0.019716
R54022 DVSS.n2187 DVSS.n2186 0.019716
R54023 DVSS.n2196 DVSS.n2055 0.019716
R54024 DVSS.n2196 DVSS.n2195 0.019716
R54025 DVSS.n2198 DVSS.n2054 0.019716
R54026 DVSS.n2199 DVSS.n2198 0.019716
R54027 DVSS.n2208 DVSS.n2053 0.019716
R54028 DVSS.n2208 DVSS.n2207 0.019716
R54029 DVSS.n2210 DVSS.n2052 0.019716
R54030 DVSS.n2211 DVSS.n2210 0.019716
R54031 DVSS.n2220 DVSS.n2051 0.019716
R54032 DVSS.n2220 DVSS.n2219 0.019716
R54033 DVSS.n2222 DVSS.n2050 0.019716
R54034 DVSS.n2223 DVSS.n2222 0.019716
R54035 DVSS.n2232 DVSS.n2049 0.019716
R54036 DVSS.n2232 DVSS.n2231 0.019716
R54037 DVSS.n2234 DVSS.n2048 0.019716
R54038 DVSS.n2235 DVSS.n2234 0.019716
R54039 DVSS.n2244 DVSS.n2047 0.019716
R54040 DVSS.n2244 DVSS.n2243 0.019716
R54041 DVSS.n2246 DVSS.n2046 0.019716
R54042 DVSS.n2247 DVSS.n2246 0.019716
R54043 DVSS.n2256 DVSS.n2045 0.019716
R54044 DVSS.n2256 DVSS.n2255 0.019716
R54045 DVSS.n2258 DVSS.n2044 0.019716
R54046 DVSS.n2259 DVSS.n2258 0.019716
R54047 DVSS.n2268 DVSS.n2043 0.019716
R54048 DVSS.n2268 DVSS.n2267 0.019716
R54049 DVSS.n2270 DVSS.n2042 0.019716
R54050 DVSS.n2271 DVSS.n2270 0.019716
R54051 DVSS.n2280 DVSS.n2041 0.019716
R54052 DVSS.n2280 DVSS.n2279 0.019716
R54053 DVSS.n2282 DVSS.n2040 0.019716
R54054 DVSS.n2283 DVSS.n2282 0.019716
R54055 DVSS.n2292 DVSS.n2039 0.019716
R54056 DVSS.n2292 DVSS.n2291 0.019716
R54057 DVSS.n2294 DVSS.n2038 0.019716
R54058 DVSS.n2295 DVSS.n2294 0.019716
R54059 DVSS.n2304 DVSS.n2037 0.019716
R54060 DVSS.n2304 DVSS.n2303 0.019716
R54061 DVSS.n2306 DVSS.n2036 0.019716
R54062 DVSS.n2307 DVSS.n2306 0.019716
R54063 DVSS.n2316 DVSS.n2035 0.019716
R54064 DVSS.n2316 DVSS.n2315 0.019716
R54065 DVSS.n2318 DVSS.n2034 0.019716
R54066 DVSS.n2319 DVSS.n2318 0.019716
R54067 DVSS.n2328 DVSS.n2033 0.019716
R54068 DVSS.n2328 DVSS.n2327 0.019716
R54069 DVSS.n2330 DVSS.n2032 0.019716
R54070 DVSS.n2331 DVSS.n2330 0.019716
R54071 DVSS.n2340 DVSS.n2031 0.019716
R54072 DVSS.n2340 DVSS.n2339 0.019716
R54073 DVSS.n2342 DVSS.n2030 0.019716
R54074 DVSS.n2343 DVSS.n2342 0.019716
R54075 DVSS.n2352 DVSS.n2029 0.019716
R54076 DVSS.n2352 DVSS.n2351 0.019716
R54077 DVSS.n2354 DVSS.n2028 0.019716
R54078 DVSS.n2355 DVSS.n2354 0.019716
R54079 DVSS.n10165 DVSS.n10164 0.019716
R54080 DVSS.n2456 DVSS.n2412 0.019716
R54081 DVSS.n2457 DVSS.n2411 0.019716
R54082 DVSS.n2466 DVSS.n2410 0.019716
R54083 DVSS.n2466 DVSS.n2465 0.019716
R54084 DVSS.n2468 DVSS.n2409 0.019716
R54085 DVSS.n2469 DVSS.n2468 0.019716
R54086 DVSS.n2478 DVSS.n2408 0.019716
R54087 DVSS.n2478 DVSS.n2477 0.019716
R54088 DVSS.n2480 DVSS.n2407 0.019716
R54089 DVSS.n2481 DVSS.n2480 0.019716
R54090 DVSS.n2490 DVSS.n2406 0.019716
R54091 DVSS.n2490 DVSS.n2489 0.019716
R54092 DVSS.n2492 DVSS.n2405 0.019716
R54093 DVSS.n2493 DVSS.n2492 0.019716
R54094 DVSS.n2502 DVSS.n2404 0.019716
R54095 DVSS.n2502 DVSS.n2501 0.019716
R54096 DVSS.n2504 DVSS.n2403 0.019716
R54097 DVSS.n2505 DVSS.n2504 0.019716
R54098 DVSS.n2514 DVSS.n2402 0.019716
R54099 DVSS.n2514 DVSS.n2513 0.019716
R54100 DVSS.n2516 DVSS.n2401 0.019716
R54101 DVSS.n2517 DVSS.n2516 0.019716
R54102 DVSS.n2526 DVSS.n2400 0.019716
R54103 DVSS.n2526 DVSS.n2525 0.019716
R54104 DVSS.n2528 DVSS.n2399 0.019716
R54105 DVSS.n2529 DVSS.n2528 0.019716
R54106 DVSS.n2538 DVSS.n2398 0.019716
R54107 DVSS.n2538 DVSS.n2537 0.019716
R54108 DVSS.n2540 DVSS.n2397 0.019716
R54109 DVSS.n2541 DVSS.n2540 0.019716
R54110 DVSS.n2550 DVSS.n2396 0.019716
R54111 DVSS.n2550 DVSS.n2549 0.019716
R54112 DVSS.n2552 DVSS.n2395 0.019716
R54113 DVSS.n2553 DVSS.n2552 0.019716
R54114 DVSS.n2562 DVSS.n2394 0.019716
R54115 DVSS.n2562 DVSS.n2561 0.019716
R54116 DVSS.n2564 DVSS.n2393 0.019716
R54117 DVSS.n2565 DVSS.n2564 0.019716
R54118 DVSS.n2574 DVSS.n2392 0.019716
R54119 DVSS.n2574 DVSS.n2573 0.019716
R54120 DVSS.n2576 DVSS.n2391 0.019716
R54121 DVSS.n2577 DVSS.n2576 0.019716
R54122 DVSS.n2586 DVSS.n2390 0.019716
R54123 DVSS.n2586 DVSS.n2585 0.019716
R54124 DVSS.n2588 DVSS.n2389 0.019716
R54125 DVSS.n2589 DVSS.n2588 0.019716
R54126 DVSS.n2598 DVSS.n2388 0.019716
R54127 DVSS.n2598 DVSS.n2597 0.019716
R54128 DVSS.n2600 DVSS.n2387 0.019716
R54129 DVSS.n2601 DVSS.n2600 0.019716
R54130 DVSS.n2610 DVSS.n2386 0.019716
R54131 DVSS.n2610 DVSS.n2609 0.019716
R54132 DVSS.n2612 DVSS.n2385 0.019716
R54133 DVSS.n2613 DVSS.n2612 0.019716
R54134 DVSS.n2622 DVSS.n2384 0.019716
R54135 DVSS.n2622 DVSS.n2621 0.019716
R54136 DVSS.n2624 DVSS.n2383 0.019716
R54137 DVSS.n2625 DVSS.n2624 0.019716
R54138 DVSS.n2634 DVSS.n2382 0.019716
R54139 DVSS.n2634 DVSS.n2633 0.019716
R54140 DVSS.n2636 DVSS.n2381 0.019716
R54141 DVSS.n2637 DVSS.n2636 0.019716
R54142 DVSS.n2646 DVSS.n2380 0.019716
R54143 DVSS.n2646 DVSS.n2645 0.019716
R54144 DVSS.n2648 DVSS.n2379 0.019716
R54145 DVSS.n2649 DVSS.n2648 0.019716
R54146 DVSS.n2658 DVSS.n2378 0.019716
R54147 DVSS.n2658 DVSS.n2657 0.019716
R54148 DVSS.n2660 DVSS.n2377 0.019716
R54149 DVSS.n2661 DVSS.n2660 0.019716
R54150 DVSS.n2670 DVSS.n2376 0.019716
R54151 DVSS.n2670 DVSS.n2669 0.019716
R54152 DVSS.n2672 DVSS.n2375 0.019716
R54153 DVSS.n2673 DVSS.n2672 0.019716
R54154 DVSS.n2682 DVSS.n2374 0.019716
R54155 DVSS.n2682 DVSS.n2681 0.019716
R54156 DVSS.n2684 DVSS.n2373 0.019716
R54157 DVSS.n2685 DVSS.n2684 0.019716
R54158 DVSS.n2694 DVSS.n2372 0.019716
R54159 DVSS.n2694 DVSS.n2693 0.019716
R54160 DVSS.n2696 DVSS.n2371 0.019716
R54161 DVSS.n2697 DVSS.n2696 0.019716
R54162 DVSS.n10140 DVSS.n10139 0.019716
R54163 DVSS.n9861 DVSS.n9860 0.019716
R54164 DVSS.n9863 DVSS.n9862 0.019716
R54165 DVSS.n9864 DVSS.n9855 0.019716
R54166 DVSS.n9865 DVSS.n9864 0.019716
R54167 DVSS.n9875 DVSS.n9874 0.019716
R54168 DVSS.n9874 DVSS.n9873 0.019716
R54169 DVSS.n9876 DVSS.n9851 0.019716
R54170 DVSS.n9877 DVSS.n9876 0.019716
R54171 DVSS.n9887 DVSS.n9886 0.019716
R54172 DVSS.n9886 DVSS.n9885 0.019716
R54173 DVSS.n9888 DVSS.n9847 0.019716
R54174 DVSS.n9889 DVSS.n9888 0.019716
R54175 DVSS.n9899 DVSS.n9898 0.019716
R54176 DVSS.n9898 DVSS.n9897 0.019716
R54177 DVSS.n9900 DVSS.n9843 0.019716
R54178 DVSS.n9901 DVSS.n9900 0.019716
R54179 DVSS.n9911 DVSS.n9910 0.019716
R54180 DVSS.n9910 DVSS.n9909 0.019716
R54181 DVSS.n9912 DVSS.n9839 0.019716
R54182 DVSS.n9913 DVSS.n9912 0.019716
R54183 DVSS.n9923 DVSS.n9922 0.019716
R54184 DVSS.n9922 DVSS.n9921 0.019716
R54185 DVSS.n9924 DVSS.n9835 0.019716
R54186 DVSS.n9925 DVSS.n9924 0.019716
R54187 DVSS.n9935 DVSS.n9934 0.019716
R54188 DVSS.n9934 DVSS.n9933 0.019716
R54189 DVSS.n9936 DVSS.n9831 0.019716
R54190 DVSS.n9937 DVSS.n9936 0.019716
R54191 DVSS.n9947 DVSS.n9946 0.019716
R54192 DVSS.n9946 DVSS.n9945 0.019716
R54193 DVSS.n9948 DVSS.n9827 0.019716
R54194 DVSS.n9949 DVSS.n9948 0.019716
R54195 DVSS.n9959 DVSS.n9958 0.019716
R54196 DVSS.n9958 DVSS.n9957 0.019716
R54197 DVSS.n9960 DVSS.n9823 0.019716
R54198 DVSS.n9961 DVSS.n9960 0.019716
R54199 DVSS.n9971 DVSS.n9970 0.019716
R54200 DVSS.n9970 DVSS.n9969 0.019716
R54201 DVSS.n9972 DVSS.n9819 0.019716
R54202 DVSS.n9973 DVSS.n9972 0.019716
R54203 DVSS.n9983 DVSS.n9982 0.019716
R54204 DVSS.n9982 DVSS.n9981 0.019716
R54205 DVSS.n9984 DVSS.n9815 0.019716
R54206 DVSS.n9985 DVSS.n9984 0.019716
R54207 DVSS.n9995 DVSS.n9994 0.019716
R54208 DVSS.n9994 DVSS.n9993 0.019716
R54209 DVSS.n9996 DVSS.n9811 0.019716
R54210 DVSS.n9997 DVSS.n9996 0.019716
R54211 DVSS.n10007 DVSS.n10006 0.019716
R54212 DVSS.n10006 DVSS.n10005 0.019716
R54213 DVSS.n10008 DVSS.n9807 0.019716
R54214 DVSS.n10009 DVSS.n10008 0.019716
R54215 DVSS.n10019 DVSS.n10018 0.019716
R54216 DVSS.n10018 DVSS.n10017 0.019716
R54217 DVSS.n10020 DVSS.n9803 0.019716
R54218 DVSS.n10021 DVSS.n10020 0.019716
R54219 DVSS.n10031 DVSS.n10030 0.019716
R54220 DVSS.n10030 DVSS.n10029 0.019716
R54221 DVSS.n10032 DVSS.n9799 0.019716
R54222 DVSS.n10033 DVSS.n10032 0.019716
R54223 DVSS.n10043 DVSS.n10042 0.019716
R54224 DVSS.n10042 DVSS.n10041 0.019716
R54225 DVSS.n10044 DVSS.n9795 0.019716
R54226 DVSS.n10045 DVSS.n10044 0.019716
R54227 DVSS.n10055 DVSS.n10054 0.019716
R54228 DVSS.n10054 DVSS.n10053 0.019716
R54229 DVSS.n10056 DVSS.n9791 0.019716
R54230 DVSS.n10057 DVSS.n10056 0.019716
R54231 DVSS.n10067 DVSS.n10066 0.019716
R54232 DVSS.n10066 DVSS.n10065 0.019716
R54233 DVSS.n10068 DVSS.n9787 0.019716
R54234 DVSS.n10069 DVSS.n10068 0.019716
R54235 DVSS.n10079 DVSS.n10078 0.019716
R54236 DVSS.n10078 DVSS.n10077 0.019716
R54237 DVSS.n10080 DVSS.n9783 0.019716
R54238 DVSS.n10081 DVSS.n10080 0.019716
R54239 DVSS.n10091 DVSS.n10090 0.019716
R54240 DVSS.n10090 DVSS.n10089 0.019716
R54241 DVSS.n10092 DVSS.n9779 0.019716
R54242 DVSS.n10093 DVSS.n10092 0.019716
R54243 DVSS.n10104 DVSS.n10103 0.019716
R54244 DVSS.n10103 DVSS.n10102 0.019716
R54245 DVSS.n10107 DVSS.n10106 0.019716
R54246 DVSS.n9758 DVSS.n9757 0.019716
R54247 DVSS.n9467 DVSS.n9466 0.019716
R54248 DVSS.n9750 DVSS.n9749 0.019716
R54249 DVSS.n9750 DVSS.n2780 0.019716
R54250 DVSS.n9745 DVSS.n9744 0.019716
R54251 DVSS.n9745 DVSS.n2779 0.019716
R54252 DVSS.n9738 DVSS.n9737 0.019716
R54253 DVSS.n9738 DVSS.n2778 0.019716
R54254 DVSS.n9733 DVSS.n9732 0.019716
R54255 DVSS.n9733 DVSS.n2777 0.019716
R54256 DVSS.n9726 DVSS.n9725 0.019716
R54257 DVSS.n9726 DVSS.n2776 0.019716
R54258 DVSS.n9721 DVSS.n9720 0.019716
R54259 DVSS.n9721 DVSS.n2775 0.019716
R54260 DVSS.n9714 DVSS.n9713 0.019716
R54261 DVSS.n9714 DVSS.n2774 0.019716
R54262 DVSS.n9709 DVSS.n9708 0.019716
R54263 DVSS.n9709 DVSS.n2773 0.019716
R54264 DVSS.n9702 DVSS.n9701 0.019716
R54265 DVSS.n9702 DVSS.n2772 0.019716
R54266 DVSS.n9697 DVSS.n9696 0.019716
R54267 DVSS.n9697 DVSS.n2771 0.019716
R54268 DVSS.n9690 DVSS.n9689 0.019716
R54269 DVSS.n9690 DVSS.n2770 0.019716
R54270 DVSS.n9685 DVSS.n9684 0.019716
R54271 DVSS.n9685 DVSS.n2769 0.019716
R54272 DVSS.n9678 DVSS.n9677 0.019716
R54273 DVSS.n9678 DVSS.n2768 0.019716
R54274 DVSS.n9673 DVSS.n9672 0.019716
R54275 DVSS.n9673 DVSS.n2767 0.019716
R54276 DVSS.n9666 DVSS.n9665 0.019716
R54277 DVSS.n9666 DVSS.n2766 0.019716
R54278 DVSS.n9661 DVSS.n9660 0.019716
R54279 DVSS.n9661 DVSS.n2765 0.019716
R54280 DVSS.n9654 DVSS.n9653 0.019716
R54281 DVSS.n9654 DVSS.n2764 0.019716
R54282 DVSS.n9649 DVSS.n9648 0.019716
R54283 DVSS.n9649 DVSS.n2763 0.019716
R54284 DVSS.n9642 DVSS.n9641 0.019716
R54285 DVSS.n9642 DVSS.n2762 0.019716
R54286 DVSS.n9637 DVSS.n9636 0.019716
R54287 DVSS.n9637 DVSS.n2761 0.019716
R54288 DVSS.n9630 DVSS.n9629 0.019716
R54289 DVSS.n9630 DVSS.n2760 0.019716
R54290 DVSS.n9625 DVSS.n9624 0.019716
R54291 DVSS.n9625 DVSS.n2759 0.019716
R54292 DVSS.n9618 DVSS.n9617 0.019716
R54293 DVSS.n9618 DVSS.n2758 0.019716
R54294 DVSS.n9613 DVSS.n9612 0.019716
R54295 DVSS.n9613 DVSS.n2757 0.019716
R54296 DVSS.n9606 DVSS.n9605 0.019716
R54297 DVSS.n9606 DVSS.n2756 0.019716
R54298 DVSS.n9601 DVSS.n9600 0.019716
R54299 DVSS.n9601 DVSS.n2755 0.019716
R54300 DVSS.n9594 DVSS.n9593 0.019716
R54301 DVSS.n9594 DVSS.n2754 0.019716
R54302 DVSS.n9589 DVSS.n9588 0.019716
R54303 DVSS.n9589 DVSS.n2753 0.019716
R54304 DVSS.n9582 DVSS.n9581 0.019716
R54305 DVSS.n9582 DVSS.n2752 0.019716
R54306 DVSS.n9577 DVSS.n9576 0.019716
R54307 DVSS.n9577 DVSS.n2751 0.019716
R54308 DVSS.n9570 DVSS.n9569 0.019716
R54309 DVSS.n9570 DVSS.n2750 0.019716
R54310 DVSS.n9565 DVSS.n9564 0.019716
R54311 DVSS.n9565 DVSS.n2749 0.019716
R54312 DVSS.n9558 DVSS.n9557 0.019716
R54313 DVSS.n9558 DVSS.n2748 0.019716
R54314 DVSS.n9553 DVSS.n9552 0.019716
R54315 DVSS.n9553 DVSS.n2747 0.019716
R54316 DVSS.n9546 DVSS.n9545 0.019716
R54317 DVSS.n9546 DVSS.n2746 0.019716
R54318 DVSS.n9541 DVSS.n9540 0.019716
R54319 DVSS.n9541 DVSS.n2745 0.019716
R54320 DVSS.n9534 DVSS.n9533 0.019716
R54321 DVSS.n9534 DVSS.n2744 0.019716
R54322 DVSS.n9529 DVSS.n9528 0.019716
R54323 DVSS.n9529 DVSS.n2743 0.019716
R54324 DVSS.n9522 DVSS.n9521 0.019716
R54325 DVSS.n9522 DVSS.n2742 0.019716
R54326 DVSS.n9517 DVSS.n9516 0.019716
R54327 DVSS.n9517 DVSS.n2741 0.019716
R54328 DVSS.n9510 DVSS.n2740 0.019716
R54329 DVSS.n2872 DVSS.n2829 0.019716
R54330 DVSS.n2873 DVSS.n2828 0.019716
R54331 DVSS.n9213 DVSS.n2827 0.019716
R54332 DVSS.n9213 DVSS.n9212 0.019716
R54333 DVSS.n9215 DVSS.n2826 0.019716
R54334 DVSS.n9216 DVSS.n9215 0.019716
R54335 DVSS.n9225 DVSS.n2825 0.019716
R54336 DVSS.n9225 DVSS.n9224 0.019716
R54337 DVSS.n9227 DVSS.n2824 0.019716
R54338 DVSS.n9228 DVSS.n9227 0.019716
R54339 DVSS.n9237 DVSS.n2823 0.019716
R54340 DVSS.n9237 DVSS.n9236 0.019716
R54341 DVSS.n9239 DVSS.n2822 0.019716
R54342 DVSS.n9240 DVSS.n9239 0.019716
R54343 DVSS.n9249 DVSS.n2821 0.019716
R54344 DVSS.n9249 DVSS.n9248 0.019716
R54345 DVSS.n9251 DVSS.n2820 0.019716
R54346 DVSS.n9252 DVSS.n9251 0.019716
R54347 DVSS.n9261 DVSS.n2819 0.019716
R54348 DVSS.n9261 DVSS.n9260 0.019716
R54349 DVSS.n9263 DVSS.n2818 0.019716
R54350 DVSS.n9264 DVSS.n9263 0.019716
R54351 DVSS.n9273 DVSS.n2817 0.019716
R54352 DVSS.n9273 DVSS.n9272 0.019716
R54353 DVSS.n9275 DVSS.n2816 0.019716
R54354 DVSS.n9276 DVSS.n9275 0.019716
R54355 DVSS.n9285 DVSS.n2815 0.019716
R54356 DVSS.n9285 DVSS.n9284 0.019716
R54357 DVSS.n9287 DVSS.n2814 0.019716
R54358 DVSS.n9288 DVSS.n9287 0.019716
R54359 DVSS.n9297 DVSS.n2813 0.019716
R54360 DVSS.n9297 DVSS.n9296 0.019716
R54361 DVSS.n9299 DVSS.n2812 0.019716
R54362 DVSS.n9300 DVSS.n9299 0.019716
R54363 DVSS.n9309 DVSS.n2811 0.019716
R54364 DVSS.n9309 DVSS.n9308 0.019716
R54365 DVSS.n9311 DVSS.n2810 0.019716
R54366 DVSS.n9312 DVSS.n9311 0.019716
R54367 DVSS.n9321 DVSS.n2809 0.019716
R54368 DVSS.n9321 DVSS.n9320 0.019716
R54369 DVSS.n9323 DVSS.n2808 0.019716
R54370 DVSS.n9324 DVSS.n9323 0.019716
R54371 DVSS.n9333 DVSS.n2807 0.019716
R54372 DVSS.n9333 DVSS.n9332 0.019716
R54373 DVSS.n9335 DVSS.n2806 0.019716
R54374 DVSS.n9336 DVSS.n9335 0.019716
R54375 DVSS.n9345 DVSS.n2805 0.019716
R54376 DVSS.n9345 DVSS.n9344 0.019716
R54377 DVSS.n9347 DVSS.n2804 0.019716
R54378 DVSS.n9348 DVSS.n9347 0.019716
R54379 DVSS.n9357 DVSS.n2803 0.019716
R54380 DVSS.n9357 DVSS.n9356 0.019716
R54381 DVSS.n9359 DVSS.n2802 0.019716
R54382 DVSS.n9360 DVSS.n9359 0.019716
R54383 DVSS.n9369 DVSS.n2801 0.019716
R54384 DVSS.n9369 DVSS.n9368 0.019716
R54385 DVSS.n9371 DVSS.n2800 0.019716
R54386 DVSS.n9372 DVSS.n9371 0.019716
R54387 DVSS.n9381 DVSS.n2799 0.019716
R54388 DVSS.n9381 DVSS.n9380 0.019716
R54389 DVSS.n9383 DVSS.n2798 0.019716
R54390 DVSS.n9384 DVSS.n9383 0.019716
R54391 DVSS.n9393 DVSS.n2797 0.019716
R54392 DVSS.n9393 DVSS.n9392 0.019716
R54393 DVSS.n9395 DVSS.n2796 0.019716
R54394 DVSS.n9396 DVSS.n9395 0.019716
R54395 DVSS.n9405 DVSS.n2795 0.019716
R54396 DVSS.n9405 DVSS.n9404 0.019716
R54397 DVSS.n9407 DVSS.n2794 0.019716
R54398 DVSS.n9408 DVSS.n9407 0.019716
R54399 DVSS.n9417 DVSS.n2793 0.019716
R54400 DVSS.n9417 DVSS.n9416 0.019716
R54401 DVSS.n9419 DVSS.n2792 0.019716
R54402 DVSS.n9420 DVSS.n9419 0.019716
R54403 DVSS.n9429 DVSS.n2791 0.019716
R54404 DVSS.n9429 DVSS.n9428 0.019716
R54405 DVSS.n9431 DVSS.n2790 0.019716
R54406 DVSS.n9432 DVSS.n9431 0.019716
R54407 DVSS.n9441 DVSS.n2789 0.019716
R54408 DVSS.n9441 DVSS.n9440 0.019716
R54409 DVSS.n9443 DVSS.n2788 0.019716
R54410 DVSS.n9444 DVSS.n9443 0.019716
R54411 DVSS.n9454 DVSS.n9453 0.019716
R54412 DVSS.n9186 DVSS.n9185 0.019716
R54413 DVSS.n2978 DVSS.n2933 0.019716
R54414 DVSS.n9002 DVSS.n2977 0.019716
R54415 DVSS.n9002 DVSS.n2931 0.019716
R54416 DVSS.n3036 DVSS.n2976 0.019716
R54417 DVSS.n3036 DVSS.n2930 0.019716
R54418 DVSS.n9011 DVSS.n2975 0.019716
R54419 DVSS.n9011 DVSS.n2929 0.019716
R54420 DVSS.n3033 DVSS.n2974 0.019716
R54421 DVSS.n3033 DVSS.n2928 0.019716
R54422 DVSS.n9020 DVSS.n2973 0.019716
R54423 DVSS.n9020 DVSS.n2927 0.019716
R54424 DVSS.n3030 DVSS.n2972 0.019716
R54425 DVSS.n3030 DVSS.n2926 0.019716
R54426 DVSS.n9029 DVSS.n2971 0.019716
R54427 DVSS.n9029 DVSS.n2925 0.019716
R54428 DVSS.n3027 DVSS.n2970 0.019716
R54429 DVSS.n3027 DVSS.n2924 0.019716
R54430 DVSS.n9038 DVSS.n2969 0.019716
R54431 DVSS.n9038 DVSS.n2923 0.019716
R54432 DVSS.n3024 DVSS.n2968 0.019716
R54433 DVSS.n3024 DVSS.n2922 0.019716
R54434 DVSS.n9047 DVSS.n2967 0.019716
R54435 DVSS.n9047 DVSS.n2921 0.019716
R54436 DVSS.n3021 DVSS.n2966 0.019716
R54437 DVSS.n3021 DVSS.n2920 0.019716
R54438 DVSS.n9056 DVSS.n2965 0.019716
R54439 DVSS.n9056 DVSS.n2919 0.019716
R54440 DVSS.n3018 DVSS.n2964 0.019716
R54441 DVSS.n3018 DVSS.n2918 0.019716
R54442 DVSS.n9065 DVSS.n2963 0.019716
R54443 DVSS.n9065 DVSS.n2917 0.019716
R54444 DVSS.n3015 DVSS.n2962 0.019716
R54445 DVSS.n3015 DVSS.n2916 0.019716
R54446 DVSS.n9074 DVSS.n2961 0.019716
R54447 DVSS.n9074 DVSS.n2915 0.019716
R54448 DVSS.n3012 DVSS.n2960 0.019716
R54449 DVSS.n3012 DVSS.n2914 0.019716
R54450 DVSS.n9083 DVSS.n2959 0.019716
R54451 DVSS.n9083 DVSS.n2913 0.019716
R54452 DVSS.n3009 DVSS.n2958 0.019716
R54453 DVSS.n3009 DVSS.n2912 0.019716
R54454 DVSS.n9092 DVSS.n2957 0.019716
R54455 DVSS.n9092 DVSS.n2911 0.019716
R54456 DVSS.n3006 DVSS.n2956 0.019716
R54457 DVSS.n3006 DVSS.n2910 0.019716
R54458 DVSS.n9101 DVSS.n2955 0.019716
R54459 DVSS.n9101 DVSS.n2909 0.019716
R54460 DVSS.n3003 DVSS.n2954 0.019716
R54461 DVSS.n3003 DVSS.n2908 0.019716
R54462 DVSS.n9110 DVSS.n2953 0.019716
R54463 DVSS.n9110 DVSS.n2907 0.019716
R54464 DVSS.n3000 DVSS.n2952 0.019716
R54465 DVSS.n3000 DVSS.n2906 0.019716
R54466 DVSS.n9119 DVSS.n2951 0.019716
R54467 DVSS.n9119 DVSS.n2905 0.019716
R54468 DVSS.n2997 DVSS.n2950 0.019716
R54469 DVSS.n2997 DVSS.n2904 0.019716
R54470 DVSS.n9128 DVSS.n2949 0.019716
R54471 DVSS.n9128 DVSS.n2903 0.019716
R54472 DVSS.n2994 DVSS.n2948 0.019716
R54473 DVSS.n2994 DVSS.n2902 0.019716
R54474 DVSS.n9137 DVSS.n2947 0.019716
R54475 DVSS.n9137 DVSS.n2901 0.019716
R54476 DVSS.n2991 DVSS.n2946 0.019716
R54477 DVSS.n2991 DVSS.n2900 0.019716
R54478 DVSS.n9146 DVSS.n2945 0.019716
R54479 DVSS.n9146 DVSS.n2899 0.019716
R54480 DVSS.n2988 DVSS.n2944 0.019716
R54481 DVSS.n2988 DVSS.n2898 0.019716
R54482 DVSS.n9155 DVSS.n2943 0.019716
R54483 DVSS.n9155 DVSS.n2897 0.019716
R54484 DVSS.n2985 DVSS.n2942 0.019716
R54485 DVSS.n2985 DVSS.n2896 0.019716
R54486 DVSS.n9164 DVSS.n2941 0.019716
R54487 DVSS.n9164 DVSS.n2895 0.019716
R54488 DVSS.n2982 DVSS.n2940 0.019716
R54489 DVSS.n2982 DVSS.n2894 0.019716
R54490 DVSS.n9173 DVSS.n2939 0.019716
R54491 DVSS.n9173 DVSS.n2893 0.019716
R54492 DVSS.n2979 DVSS.n2938 0.019716
R54493 DVSS.n2979 DVSS.n2892 0.019716
R54494 DVSS.n9183 DVSS.n2891 0.019716
R54495 DVSS.n8968 DVSS.n8967 0.019716
R54496 DVSS.n8678 DVSS.n8677 0.019716
R54497 DVSS.n8960 DVSS.n8959 0.019716
R54498 DVSS.n8960 DVSS.n8676 0.019716
R54499 DVSS.n8955 DVSS.n8954 0.019716
R54500 DVSS.n8955 DVSS.n8675 0.019716
R54501 DVSS.n8948 DVSS.n8947 0.019716
R54502 DVSS.n8948 DVSS.n8674 0.019716
R54503 DVSS.n8943 DVSS.n8942 0.019716
R54504 DVSS.n8943 DVSS.n8673 0.019716
R54505 DVSS.n8936 DVSS.n8935 0.019716
R54506 DVSS.n8936 DVSS.n8672 0.019716
R54507 DVSS.n8931 DVSS.n8930 0.019716
R54508 DVSS.n8931 DVSS.n8671 0.019716
R54509 DVSS.n8924 DVSS.n8923 0.019716
R54510 DVSS.n8924 DVSS.n8670 0.019716
R54511 DVSS.n8919 DVSS.n8918 0.019716
R54512 DVSS.n8919 DVSS.n8669 0.019716
R54513 DVSS.n8912 DVSS.n8911 0.019716
R54514 DVSS.n8912 DVSS.n8668 0.019716
R54515 DVSS.n8907 DVSS.n8906 0.019716
R54516 DVSS.n8907 DVSS.n8667 0.019716
R54517 DVSS.n8900 DVSS.n8899 0.019716
R54518 DVSS.n8900 DVSS.n8666 0.019716
R54519 DVSS.n8895 DVSS.n8894 0.019716
R54520 DVSS.n8895 DVSS.n8665 0.019716
R54521 DVSS.n8888 DVSS.n8887 0.019716
R54522 DVSS.n8888 DVSS.n8664 0.019716
R54523 DVSS.n8883 DVSS.n8882 0.019716
R54524 DVSS.n8883 DVSS.n8663 0.019716
R54525 DVSS.n8876 DVSS.n8875 0.019716
R54526 DVSS.n8876 DVSS.n8662 0.019716
R54527 DVSS.n8871 DVSS.n8870 0.019716
R54528 DVSS.n8871 DVSS.n8661 0.019716
R54529 DVSS.n8864 DVSS.n8863 0.019716
R54530 DVSS.n8864 DVSS.n8660 0.019716
R54531 DVSS.n8859 DVSS.n8858 0.019716
R54532 DVSS.n8859 DVSS.n8659 0.019716
R54533 DVSS.n8852 DVSS.n8851 0.019716
R54534 DVSS.n8852 DVSS.n8658 0.019716
R54535 DVSS.n8847 DVSS.n8846 0.019716
R54536 DVSS.n8847 DVSS.n8657 0.019716
R54537 DVSS.n8840 DVSS.n8839 0.019716
R54538 DVSS.n8840 DVSS.n8656 0.019716
R54539 DVSS.n8835 DVSS.n8834 0.019716
R54540 DVSS.n8835 DVSS.n8655 0.019716
R54541 DVSS.n8828 DVSS.n8827 0.019716
R54542 DVSS.n8828 DVSS.n8654 0.019716
R54543 DVSS.n8823 DVSS.n8822 0.019716
R54544 DVSS.n8823 DVSS.n8653 0.019716
R54545 DVSS.n8816 DVSS.n8815 0.019716
R54546 DVSS.n8816 DVSS.n8652 0.019716
R54547 DVSS.n8811 DVSS.n8810 0.019716
R54548 DVSS.n8811 DVSS.n8651 0.019716
R54549 DVSS.n8804 DVSS.n8803 0.019716
R54550 DVSS.n8804 DVSS.n8650 0.019716
R54551 DVSS.n8799 DVSS.n8798 0.019716
R54552 DVSS.n8799 DVSS.n8649 0.019716
R54553 DVSS.n8792 DVSS.n8791 0.019716
R54554 DVSS.n8792 DVSS.n8648 0.019716
R54555 DVSS.n8787 DVSS.n8786 0.019716
R54556 DVSS.n8787 DVSS.n8647 0.019716
R54557 DVSS.n8780 DVSS.n8779 0.019716
R54558 DVSS.n8780 DVSS.n8646 0.019716
R54559 DVSS.n8775 DVSS.n8774 0.019716
R54560 DVSS.n8775 DVSS.n8645 0.019716
R54561 DVSS.n8768 DVSS.n8767 0.019716
R54562 DVSS.n8768 DVSS.n8644 0.019716
R54563 DVSS.n8763 DVSS.n8762 0.019716
R54564 DVSS.n8763 DVSS.n8643 0.019716
R54565 DVSS.n8756 DVSS.n8755 0.019716
R54566 DVSS.n8756 DVSS.n8642 0.019716
R54567 DVSS.n8751 DVSS.n8750 0.019716
R54568 DVSS.n8751 DVSS.n8641 0.019716
R54569 DVSS.n8744 DVSS.n8743 0.019716
R54570 DVSS.n8744 DVSS.n8640 0.019716
R54571 DVSS.n8739 DVSS.n8738 0.019716
R54572 DVSS.n8739 DVSS.n8639 0.019716
R54573 DVSS.n8732 DVSS.n8731 0.019716
R54574 DVSS.n8732 DVSS.n8638 0.019716
R54575 DVSS.n8727 DVSS.n8726 0.019716
R54576 DVSS.n8727 DVSS.n8637 0.019716
R54577 DVSS.n8720 DVSS.n8636 0.019716
R54578 DVSS.n3154 DVSS.n3153 0.019716
R54579 DVSS.n3156 DVSS.n3155 0.019716
R54580 DVSS.n3157 DVSS.n3148 0.019716
R54581 DVSS.n3158 DVSS.n3157 0.019716
R54582 DVSS.n3168 DVSS.n3167 0.019716
R54583 DVSS.n3167 DVSS.n3166 0.019716
R54584 DVSS.n3169 DVSS.n3144 0.019716
R54585 DVSS.n3170 DVSS.n3169 0.019716
R54586 DVSS.n3180 DVSS.n3179 0.019716
R54587 DVSS.n3179 DVSS.n3178 0.019716
R54588 DVSS.n3181 DVSS.n3140 0.019716
R54589 DVSS.n3182 DVSS.n3181 0.019716
R54590 DVSS.n3192 DVSS.n3191 0.019716
R54591 DVSS.n3191 DVSS.n3190 0.019716
R54592 DVSS.n3193 DVSS.n3136 0.019716
R54593 DVSS.n3194 DVSS.n3193 0.019716
R54594 DVSS.n3204 DVSS.n3203 0.019716
R54595 DVSS.n3203 DVSS.n3202 0.019716
R54596 DVSS.n3205 DVSS.n3132 0.019716
R54597 DVSS.n3206 DVSS.n3205 0.019716
R54598 DVSS.n3216 DVSS.n3215 0.019716
R54599 DVSS.n3215 DVSS.n3214 0.019716
R54600 DVSS.n3217 DVSS.n3128 0.019716
R54601 DVSS.n3218 DVSS.n3217 0.019716
R54602 DVSS.n3228 DVSS.n3227 0.019716
R54603 DVSS.n3227 DVSS.n3226 0.019716
R54604 DVSS.n3229 DVSS.n3124 0.019716
R54605 DVSS.n3230 DVSS.n3229 0.019716
R54606 DVSS.n3240 DVSS.n3239 0.019716
R54607 DVSS.n3239 DVSS.n3238 0.019716
R54608 DVSS.n3241 DVSS.n3120 0.019716
R54609 DVSS.n3242 DVSS.n3241 0.019716
R54610 DVSS.n3252 DVSS.n3251 0.019716
R54611 DVSS.n3251 DVSS.n3250 0.019716
R54612 DVSS.n3253 DVSS.n3116 0.019716
R54613 DVSS.n3254 DVSS.n3253 0.019716
R54614 DVSS.n3264 DVSS.n3263 0.019716
R54615 DVSS.n3263 DVSS.n3262 0.019716
R54616 DVSS.n3265 DVSS.n3112 0.019716
R54617 DVSS.n3266 DVSS.n3265 0.019716
R54618 DVSS.n3276 DVSS.n3275 0.019716
R54619 DVSS.n3275 DVSS.n3274 0.019716
R54620 DVSS.n3277 DVSS.n3108 0.019716
R54621 DVSS.n3278 DVSS.n3277 0.019716
R54622 DVSS.n3288 DVSS.n3287 0.019716
R54623 DVSS.n3287 DVSS.n3286 0.019716
R54624 DVSS.n3289 DVSS.n3104 0.019716
R54625 DVSS.n3290 DVSS.n3289 0.019716
R54626 DVSS.n3300 DVSS.n3299 0.019716
R54627 DVSS.n3299 DVSS.n3298 0.019716
R54628 DVSS.n3301 DVSS.n3100 0.019716
R54629 DVSS.n3302 DVSS.n3301 0.019716
R54630 DVSS.n3312 DVSS.n3311 0.019716
R54631 DVSS.n3311 DVSS.n3310 0.019716
R54632 DVSS.n3313 DVSS.n3096 0.019716
R54633 DVSS.n3314 DVSS.n3313 0.019716
R54634 DVSS.n3324 DVSS.n3323 0.019716
R54635 DVSS.n3323 DVSS.n3322 0.019716
R54636 DVSS.n3325 DVSS.n3092 0.019716
R54637 DVSS.n3326 DVSS.n3325 0.019716
R54638 DVSS.n3336 DVSS.n3335 0.019716
R54639 DVSS.n3335 DVSS.n3334 0.019716
R54640 DVSS.n3337 DVSS.n3088 0.019716
R54641 DVSS.n3338 DVSS.n3337 0.019716
R54642 DVSS.n3348 DVSS.n3347 0.019716
R54643 DVSS.n3347 DVSS.n3346 0.019716
R54644 DVSS.n3349 DVSS.n3084 0.019716
R54645 DVSS.n3350 DVSS.n3349 0.019716
R54646 DVSS.n3360 DVSS.n3359 0.019716
R54647 DVSS.n3359 DVSS.n3358 0.019716
R54648 DVSS.n3361 DVSS.n3080 0.019716
R54649 DVSS.n3362 DVSS.n3361 0.019716
R54650 DVSS.n3372 DVSS.n3371 0.019716
R54651 DVSS.n3371 DVSS.n3370 0.019716
R54652 DVSS.n3373 DVSS.n3076 0.019716
R54653 DVSS.n3374 DVSS.n3373 0.019716
R54654 DVSS.n3384 DVSS.n3383 0.019716
R54655 DVSS.n3383 DVSS.n3382 0.019716
R54656 DVSS.n3385 DVSS.n3072 0.019716
R54657 DVSS.n3386 DVSS.n3385 0.019716
R54658 DVSS.n3397 DVSS.n3396 0.019716
R54659 DVSS.n3396 DVSS.n3395 0.019716
R54660 DVSS.n3400 DVSS.n3399 0.019716
R54661 DVSS.n8603 DVSS.n8602 0.019716
R54662 DVSS.n3501 DVSS.n3458 0.019716
R54663 DVSS.n3569 DVSS.n3500 0.019716
R54664 DVSS.n3569 DVSS.n3456 0.019716
R54665 DVSS.n3573 DVSS.n3499 0.019716
R54666 DVSS.n3573 DVSS.n3455 0.019716
R54667 DVSS.n3578 DVSS.n3498 0.019716
R54668 DVSS.n3578 DVSS.n3454 0.019716
R54669 DVSS.n3582 DVSS.n3497 0.019716
R54670 DVSS.n3582 DVSS.n3453 0.019716
R54671 DVSS.n3587 DVSS.n3496 0.019716
R54672 DVSS.n3587 DVSS.n3452 0.019716
R54673 DVSS.n3591 DVSS.n3495 0.019716
R54674 DVSS.n3591 DVSS.n3451 0.019716
R54675 DVSS.n3596 DVSS.n3494 0.019716
R54676 DVSS.n3596 DVSS.n3450 0.019716
R54677 DVSS.n3600 DVSS.n3493 0.019716
R54678 DVSS.n3600 DVSS.n3449 0.019716
R54679 DVSS.n3605 DVSS.n3492 0.019716
R54680 DVSS.n3605 DVSS.n3448 0.019716
R54681 DVSS.n3609 DVSS.n3491 0.019716
R54682 DVSS.n3609 DVSS.n3447 0.019716
R54683 DVSS.n3614 DVSS.n3490 0.019716
R54684 DVSS.n3614 DVSS.n3446 0.019716
R54685 DVSS.n3618 DVSS.n3489 0.019716
R54686 DVSS.n3618 DVSS.n3445 0.019716
R54687 DVSS.n3623 DVSS.n3488 0.019716
R54688 DVSS.n3623 DVSS.n3444 0.019716
R54689 DVSS.n3627 DVSS.n3487 0.019716
R54690 DVSS.n3627 DVSS.n3443 0.019716
R54691 DVSS.n3632 DVSS.n3486 0.019716
R54692 DVSS.n3632 DVSS.n3442 0.019716
R54693 DVSS.n3636 DVSS.n3485 0.019716
R54694 DVSS.n3636 DVSS.n3441 0.019716
R54695 DVSS.n3641 DVSS.n3484 0.019716
R54696 DVSS.n3641 DVSS.n3440 0.019716
R54697 DVSS.n3645 DVSS.n3483 0.019716
R54698 DVSS.n3645 DVSS.n3439 0.019716
R54699 DVSS.n3650 DVSS.n3482 0.019716
R54700 DVSS.n3650 DVSS.n3438 0.019716
R54701 DVSS.n3654 DVSS.n3481 0.019716
R54702 DVSS.n3654 DVSS.n3437 0.019716
R54703 DVSS.n3659 DVSS.n3480 0.019716
R54704 DVSS.n3659 DVSS.n3436 0.019716
R54705 DVSS.n3663 DVSS.n3479 0.019716
R54706 DVSS.n3663 DVSS.n3435 0.019716
R54707 DVSS.n3668 DVSS.n3478 0.019716
R54708 DVSS.n3668 DVSS.n3434 0.019716
R54709 DVSS.n3672 DVSS.n3477 0.019716
R54710 DVSS.n3672 DVSS.n3433 0.019716
R54711 DVSS.n3677 DVSS.n3476 0.019716
R54712 DVSS.n3677 DVSS.n3432 0.019716
R54713 DVSS.n3681 DVSS.n3475 0.019716
R54714 DVSS.n3681 DVSS.n3431 0.019716
R54715 DVSS.n3686 DVSS.n3474 0.019716
R54716 DVSS.n3686 DVSS.n3430 0.019716
R54717 DVSS.n3690 DVSS.n3473 0.019716
R54718 DVSS.n3690 DVSS.n3429 0.019716
R54719 DVSS.n3695 DVSS.n3472 0.019716
R54720 DVSS.n3695 DVSS.n3428 0.019716
R54721 DVSS.n3699 DVSS.n3471 0.019716
R54722 DVSS.n3699 DVSS.n3427 0.019716
R54723 DVSS.n3704 DVSS.n3470 0.019716
R54724 DVSS.n3704 DVSS.n3426 0.019716
R54725 DVSS.n3708 DVSS.n3469 0.019716
R54726 DVSS.n3708 DVSS.n3425 0.019716
R54727 DVSS.n3713 DVSS.n3468 0.019716
R54728 DVSS.n3713 DVSS.n3424 0.019716
R54729 DVSS.n3717 DVSS.n3467 0.019716
R54730 DVSS.n3717 DVSS.n3423 0.019716
R54731 DVSS.n3722 DVSS.n3466 0.019716
R54732 DVSS.n3722 DVSS.n3422 0.019716
R54733 DVSS.n3726 DVSS.n3465 0.019716
R54734 DVSS.n3726 DVSS.n3421 0.019716
R54735 DVSS.n3731 DVSS.n3464 0.019716
R54736 DVSS.n3731 DVSS.n3420 0.019716
R54737 DVSS.n3735 DVSS.n3463 0.019716
R54738 DVSS.n3735 DVSS.n3419 0.019716
R54739 DVSS.n3740 DVSS.n3462 0.019716
R54740 DVSS.n3740 DVSS.n3418 0.019716
R54741 DVSS.n3744 DVSS.n3461 0.019716
R54742 DVSS.n3744 DVSS.n3417 0.019716
R54743 DVSS.n8600 DVSS.n3416 0.019716
R54744 DVSS.n3840 DVSS.n3797 0.019716
R54745 DVSS.n3841 DVSS.n3796 0.019716
R54746 DVSS.n8346 DVSS.n3795 0.019716
R54747 DVSS.n8346 DVSS.n8345 0.019716
R54748 DVSS.n8348 DVSS.n3794 0.019716
R54749 DVSS.n8349 DVSS.n8348 0.019716
R54750 DVSS.n8358 DVSS.n3793 0.019716
R54751 DVSS.n8358 DVSS.n8357 0.019716
R54752 DVSS.n8360 DVSS.n3792 0.019716
R54753 DVSS.n8361 DVSS.n8360 0.019716
R54754 DVSS.n8370 DVSS.n3791 0.019716
R54755 DVSS.n8370 DVSS.n8369 0.019716
R54756 DVSS.n8372 DVSS.n3790 0.019716
R54757 DVSS.n8373 DVSS.n8372 0.019716
R54758 DVSS.n8382 DVSS.n3789 0.019716
R54759 DVSS.n8382 DVSS.n8381 0.019716
R54760 DVSS.n8384 DVSS.n3788 0.019716
R54761 DVSS.n8385 DVSS.n8384 0.019716
R54762 DVSS.n8394 DVSS.n3787 0.019716
R54763 DVSS.n8394 DVSS.n8393 0.019716
R54764 DVSS.n8396 DVSS.n3786 0.019716
R54765 DVSS.n8397 DVSS.n8396 0.019716
R54766 DVSS.n8406 DVSS.n3785 0.019716
R54767 DVSS.n8406 DVSS.n8405 0.019716
R54768 DVSS.n8408 DVSS.n3784 0.019716
R54769 DVSS.n8409 DVSS.n8408 0.019716
R54770 DVSS.n8418 DVSS.n3783 0.019716
R54771 DVSS.n8418 DVSS.n8417 0.019716
R54772 DVSS.n8420 DVSS.n3782 0.019716
R54773 DVSS.n8421 DVSS.n8420 0.019716
R54774 DVSS.n8430 DVSS.n3781 0.019716
R54775 DVSS.n8430 DVSS.n8429 0.019716
R54776 DVSS.n8432 DVSS.n3780 0.019716
R54777 DVSS.n8433 DVSS.n8432 0.019716
R54778 DVSS.n8442 DVSS.n3779 0.019716
R54779 DVSS.n8442 DVSS.n8441 0.019716
R54780 DVSS.n8444 DVSS.n3778 0.019716
R54781 DVSS.n8445 DVSS.n8444 0.019716
R54782 DVSS.n8454 DVSS.n3777 0.019716
R54783 DVSS.n8454 DVSS.n8453 0.019716
R54784 DVSS.n8456 DVSS.n3776 0.019716
R54785 DVSS.n8457 DVSS.n8456 0.019716
R54786 DVSS.n8466 DVSS.n3775 0.019716
R54787 DVSS.n8466 DVSS.n8465 0.019716
R54788 DVSS.n8468 DVSS.n3774 0.019716
R54789 DVSS.n8469 DVSS.n8468 0.019716
R54790 DVSS.n8478 DVSS.n3773 0.019716
R54791 DVSS.n8478 DVSS.n8477 0.019716
R54792 DVSS.n8480 DVSS.n3772 0.019716
R54793 DVSS.n8481 DVSS.n8480 0.019716
R54794 DVSS.n8490 DVSS.n3771 0.019716
R54795 DVSS.n8490 DVSS.n8489 0.019716
R54796 DVSS.n8492 DVSS.n3770 0.019716
R54797 DVSS.n8493 DVSS.n8492 0.019716
R54798 DVSS.n8502 DVSS.n3769 0.019716
R54799 DVSS.n8502 DVSS.n8501 0.019716
R54800 DVSS.n8504 DVSS.n3768 0.019716
R54801 DVSS.n8505 DVSS.n8504 0.019716
R54802 DVSS.n8514 DVSS.n3767 0.019716
R54803 DVSS.n8514 DVSS.n8513 0.019716
R54804 DVSS.n8516 DVSS.n3766 0.019716
R54805 DVSS.n8517 DVSS.n8516 0.019716
R54806 DVSS.n8526 DVSS.n3765 0.019716
R54807 DVSS.n8526 DVSS.n8525 0.019716
R54808 DVSS.n8528 DVSS.n3764 0.019716
R54809 DVSS.n8529 DVSS.n8528 0.019716
R54810 DVSS.n8538 DVSS.n3763 0.019716
R54811 DVSS.n8538 DVSS.n8537 0.019716
R54812 DVSS.n8540 DVSS.n3762 0.019716
R54813 DVSS.n8541 DVSS.n8540 0.019716
R54814 DVSS.n8550 DVSS.n3761 0.019716
R54815 DVSS.n8550 DVSS.n8549 0.019716
R54816 DVSS.n8552 DVSS.n3760 0.019716
R54817 DVSS.n8553 DVSS.n8552 0.019716
R54818 DVSS.n8562 DVSS.n3759 0.019716
R54819 DVSS.n8562 DVSS.n8561 0.019716
R54820 DVSS.n8564 DVSS.n3758 0.019716
R54821 DVSS.n8565 DVSS.n8564 0.019716
R54822 DVSS.n8574 DVSS.n3757 0.019716
R54823 DVSS.n8574 DVSS.n8573 0.019716
R54824 DVSS.n8576 DVSS.n3756 0.019716
R54825 DVSS.n8577 DVSS.n8576 0.019716
R54826 DVSS.n8587 DVSS.n8586 0.019716
R54827 DVSS.n8319 DVSS.n8318 0.019716
R54828 DVSS.n3945 DVSS.n3901 0.019716
R54829 DVSS.n8135 DVSS.n3944 0.019716
R54830 DVSS.n8135 DVSS.n3899 0.019716
R54831 DVSS.n4004 DVSS.n3943 0.019716
R54832 DVSS.n4004 DVSS.n3898 0.019716
R54833 DVSS.n8144 DVSS.n3942 0.019716
R54834 DVSS.n8144 DVSS.n3897 0.019716
R54835 DVSS.n4001 DVSS.n3941 0.019716
R54836 DVSS.n4001 DVSS.n3896 0.019716
R54837 DVSS.n8153 DVSS.n3940 0.019716
R54838 DVSS.n8153 DVSS.n3895 0.019716
R54839 DVSS.n3998 DVSS.n3939 0.019716
R54840 DVSS.n3998 DVSS.n3894 0.019716
R54841 DVSS.n8162 DVSS.n3938 0.019716
R54842 DVSS.n8162 DVSS.n3893 0.019716
R54843 DVSS.n3995 DVSS.n3937 0.019716
R54844 DVSS.n3995 DVSS.n3892 0.019716
R54845 DVSS.n8171 DVSS.n3936 0.019716
R54846 DVSS.n8171 DVSS.n3891 0.019716
R54847 DVSS.n3992 DVSS.n3935 0.019716
R54848 DVSS.n3992 DVSS.n3890 0.019716
R54849 DVSS.n8180 DVSS.n3934 0.019716
R54850 DVSS.n8180 DVSS.n3889 0.019716
R54851 DVSS.n3989 DVSS.n3933 0.019716
R54852 DVSS.n3989 DVSS.n3888 0.019716
R54853 DVSS.n8189 DVSS.n3932 0.019716
R54854 DVSS.n8189 DVSS.n3887 0.019716
R54855 DVSS.n3986 DVSS.n3931 0.019716
R54856 DVSS.n3986 DVSS.n3886 0.019716
R54857 DVSS.n8198 DVSS.n3930 0.019716
R54858 DVSS.n8198 DVSS.n3885 0.019716
R54859 DVSS.n3983 DVSS.n3929 0.019716
R54860 DVSS.n3983 DVSS.n3884 0.019716
R54861 DVSS.n8207 DVSS.n3928 0.019716
R54862 DVSS.n8207 DVSS.n3883 0.019716
R54863 DVSS.n3980 DVSS.n3927 0.019716
R54864 DVSS.n3980 DVSS.n3882 0.019716
R54865 DVSS.n8216 DVSS.n3926 0.019716
R54866 DVSS.n8216 DVSS.n3881 0.019716
R54867 DVSS.n3977 DVSS.n3925 0.019716
R54868 DVSS.n3977 DVSS.n3880 0.019716
R54869 DVSS.n8225 DVSS.n3924 0.019716
R54870 DVSS.n8225 DVSS.n3879 0.019716
R54871 DVSS.n3974 DVSS.n3923 0.019716
R54872 DVSS.n3974 DVSS.n3878 0.019716
R54873 DVSS.n8234 DVSS.n3922 0.019716
R54874 DVSS.n8234 DVSS.n3877 0.019716
R54875 DVSS.n3971 DVSS.n3921 0.019716
R54876 DVSS.n3971 DVSS.n3876 0.019716
R54877 DVSS.n8243 DVSS.n3920 0.019716
R54878 DVSS.n8243 DVSS.n3875 0.019716
R54879 DVSS.n3968 DVSS.n3919 0.019716
R54880 DVSS.n3968 DVSS.n3874 0.019716
R54881 DVSS.n8252 DVSS.n3918 0.019716
R54882 DVSS.n8252 DVSS.n3873 0.019716
R54883 DVSS.n3965 DVSS.n3917 0.019716
R54884 DVSS.n3965 DVSS.n3872 0.019716
R54885 DVSS.n8261 DVSS.n3916 0.019716
R54886 DVSS.n8261 DVSS.n3871 0.019716
R54887 DVSS.n3962 DVSS.n3915 0.019716
R54888 DVSS.n3962 DVSS.n3870 0.019716
R54889 DVSS.n8270 DVSS.n3914 0.019716
R54890 DVSS.n8270 DVSS.n3869 0.019716
R54891 DVSS.n3959 DVSS.n3913 0.019716
R54892 DVSS.n3959 DVSS.n3868 0.019716
R54893 DVSS.n8279 DVSS.n3912 0.019716
R54894 DVSS.n8279 DVSS.n3867 0.019716
R54895 DVSS.n3956 DVSS.n3911 0.019716
R54896 DVSS.n3956 DVSS.n3866 0.019716
R54897 DVSS.n8288 DVSS.n3910 0.019716
R54898 DVSS.n8288 DVSS.n3865 0.019716
R54899 DVSS.n3953 DVSS.n3909 0.019716
R54900 DVSS.n3953 DVSS.n3864 0.019716
R54901 DVSS.n8297 DVSS.n3908 0.019716
R54902 DVSS.n8297 DVSS.n3863 0.019716
R54903 DVSS.n3950 DVSS.n3907 0.019716
R54904 DVSS.n3950 DVSS.n3862 0.019716
R54905 DVSS.n8306 DVSS.n3906 0.019716
R54906 DVSS.n8306 DVSS.n3861 0.019716
R54907 DVSS.n3947 DVSS.n3905 0.019716
R54908 DVSS.n3947 DVSS.n3860 0.019716
R54909 DVSS.n8316 DVSS.n3859 0.019716
R54910 DVSS.n4110 DVSS.n4109 0.019716
R54911 DVSS.n4112 DVSS.n4111 0.019716
R54912 DVSS.n4113 DVSS.n4104 0.019716
R54913 DVSS.n4114 DVSS.n4113 0.019716
R54914 DVSS.n4124 DVSS.n4123 0.019716
R54915 DVSS.n4123 DVSS.n4122 0.019716
R54916 DVSS.n4125 DVSS.n4100 0.019716
R54917 DVSS.n4126 DVSS.n4125 0.019716
R54918 DVSS.n4136 DVSS.n4135 0.019716
R54919 DVSS.n4135 DVSS.n4134 0.019716
R54920 DVSS.n4137 DVSS.n4096 0.019716
R54921 DVSS.n4138 DVSS.n4137 0.019716
R54922 DVSS.n4148 DVSS.n4147 0.019716
R54923 DVSS.n4147 DVSS.n4146 0.019716
R54924 DVSS.n4149 DVSS.n4092 0.019716
R54925 DVSS.n4150 DVSS.n4149 0.019716
R54926 DVSS.n4160 DVSS.n4159 0.019716
R54927 DVSS.n4159 DVSS.n4158 0.019716
R54928 DVSS.n4161 DVSS.n4088 0.019716
R54929 DVSS.n4162 DVSS.n4161 0.019716
R54930 DVSS.n4172 DVSS.n4171 0.019716
R54931 DVSS.n4171 DVSS.n4170 0.019716
R54932 DVSS.n4173 DVSS.n4084 0.019716
R54933 DVSS.n4174 DVSS.n4173 0.019716
R54934 DVSS.n4184 DVSS.n4183 0.019716
R54935 DVSS.n4183 DVSS.n4182 0.019716
R54936 DVSS.n4185 DVSS.n4080 0.019716
R54937 DVSS.n4186 DVSS.n4185 0.019716
R54938 DVSS.n4196 DVSS.n4195 0.019716
R54939 DVSS.n4195 DVSS.n4194 0.019716
R54940 DVSS.n4197 DVSS.n4076 0.019716
R54941 DVSS.n4198 DVSS.n4197 0.019716
R54942 DVSS.n4208 DVSS.n4207 0.019716
R54943 DVSS.n4207 DVSS.n4206 0.019716
R54944 DVSS.n4209 DVSS.n4072 0.019716
R54945 DVSS.n4210 DVSS.n4209 0.019716
R54946 DVSS.n4220 DVSS.n4219 0.019716
R54947 DVSS.n4219 DVSS.n4218 0.019716
R54948 DVSS.n4221 DVSS.n4068 0.019716
R54949 DVSS.n4222 DVSS.n4221 0.019716
R54950 DVSS.n4232 DVSS.n4231 0.019716
R54951 DVSS.n4231 DVSS.n4230 0.019716
R54952 DVSS.n4233 DVSS.n4064 0.019716
R54953 DVSS.n4234 DVSS.n4233 0.019716
R54954 DVSS.n4244 DVSS.n4243 0.019716
R54955 DVSS.n4243 DVSS.n4242 0.019716
R54956 DVSS.n4245 DVSS.n4060 0.019716
R54957 DVSS.n4246 DVSS.n4245 0.019716
R54958 DVSS.n4256 DVSS.n4255 0.019716
R54959 DVSS.n4255 DVSS.n4254 0.019716
R54960 DVSS.n4257 DVSS.n4056 0.019716
R54961 DVSS.n4258 DVSS.n4257 0.019716
R54962 DVSS.n4268 DVSS.n4267 0.019716
R54963 DVSS.n4267 DVSS.n4266 0.019716
R54964 DVSS.n4269 DVSS.n4052 0.019716
R54965 DVSS.n4270 DVSS.n4269 0.019716
R54966 DVSS.n4280 DVSS.n4279 0.019716
R54967 DVSS.n4279 DVSS.n4278 0.019716
R54968 DVSS.n4281 DVSS.n4048 0.019716
R54969 DVSS.n4282 DVSS.n4281 0.019716
R54970 DVSS.n4292 DVSS.n4291 0.019716
R54971 DVSS.n4291 DVSS.n4290 0.019716
R54972 DVSS.n4293 DVSS.n4044 0.019716
R54973 DVSS.n4294 DVSS.n4293 0.019716
R54974 DVSS.n4304 DVSS.n4303 0.019716
R54975 DVSS.n4303 DVSS.n4302 0.019716
R54976 DVSS.n4305 DVSS.n4040 0.019716
R54977 DVSS.n4306 DVSS.n4305 0.019716
R54978 DVSS.n4316 DVSS.n4315 0.019716
R54979 DVSS.n4315 DVSS.n4314 0.019716
R54980 DVSS.n4317 DVSS.n4036 0.019716
R54981 DVSS.n4318 DVSS.n4317 0.019716
R54982 DVSS.n4328 DVSS.n4327 0.019716
R54983 DVSS.n4327 DVSS.n4326 0.019716
R54984 DVSS.n4329 DVSS.n4032 0.019716
R54985 DVSS.n4330 DVSS.n4329 0.019716
R54986 DVSS.n4340 DVSS.n4339 0.019716
R54987 DVSS.n4339 DVSS.n4338 0.019716
R54988 DVSS.n4341 DVSS.n4028 0.019716
R54989 DVSS.n4342 DVSS.n4341 0.019716
R54990 DVSS.n4353 DVSS.n4352 0.019716
R54991 DVSS.n4352 DVSS.n4351 0.019716
R54992 DVSS.n4356 DVSS.n4355 0.019716
R54993 DVSS.n8089 DVSS.n8088 0.019716
R54994 DVSS.n4415 DVSS.n4414 0.019716
R54995 DVSS.n8081 DVSS.n8080 0.019716
R54996 DVSS.n8081 DVSS.n4412 0.019716
R54997 DVSS.n8076 DVSS.n8075 0.019716
R54998 DVSS.n8076 DVSS.n4411 0.019716
R54999 DVSS.n8069 DVSS.n8068 0.019716
R55000 DVSS.n8069 DVSS.n4410 0.019716
R55001 DVSS.n8064 DVSS.n8063 0.019716
R55002 DVSS.n8064 DVSS.n4409 0.019716
R55003 DVSS.n8057 DVSS.n8056 0.019716
R55004 DVSS.n8057 DVSS.n4408 0.019716
R55005 DVSS.n8052 DVSS.n8051 0.019716
R55006 DVSS.n8052 DVSS.n4407 0.019716
R55007 DVSS.n8045 DVSS.n8044 0.019716
R55008 DVSS.n8045 DVSS.n4406 0.019716
R55009 DVSS.n8040 DVSS.n8039 0.019716
R55010 DVSS.n8040 DVSS.n4405 0.019716
R55011 DVSS.n8033 DVSS.n8032 0.019716
R55012 DVSS.n8033 DVSS.n4404 0.019716
R55013 DVSS.n8028 DVSS.n8027 0.019716
R55014 DVSS.n8028 DVSS.n4403 0.019716
R55015 DVSS.n8021 DVSS.n8020 0.019716
R55016 DVSS.n8021 DVSS.n4402 0.019716
R55017 DVSS.n8016 DVSS.n8015 0.019716
R55018 DVSS.n8016 DVSS.n4401 0.019716
R55019 DVSS.n8009 DVSS.n8008 0.019716
R55020 DVSS.n8009 DVSS.n4400 0.019716
R55021 DVSS.n8004 DVSS.n8003 0.019716
R55022 DVSS.n8004 DVSS.n4399 0.019716
R55023 DVSS.n7997 DVSS.n7996 0.019716
R55024 DVSS.n7997 DVSS.n4398 0.019716
R55025 DVSS.n7992 DVSS.n7991 0.019716
R55026 DVSS.n7992 DVSS.n4397 0.019716
R55027 DVSS.n7985 DVSS.n7984 0.019716
R55028 DVSS.n7985 DVSS.n4396 0.019716
R55029 DVSS.n7980 DVSS.n7979 0.019716
R55030 DVSS.n7980 DVSS.n4395 0.019716
R55031 DVSS.n7973 DVSS.n7972 0.019716
R55032 DVSS.n7973 DVSS.n4394 0.019716
R55033 DVSS.n7968 DVSS.n7967 0.019716
R55034 DVSS.n7968 DVSS.n4393 0.019716
R55035 DVSS.n7961 DVSS.n7960 0.019716
R55036 DVSS.n7961 DVSS.n4392 0.019716
R55037 DVSS.n7956 DVSS.n7955 0.019716
R55038 DVSS.n7956 DVSS.n4391 0.019716
R55039 DVSS.n7949 DVSS.n7948 0.019716
R55040 DVSS.n7949 DVSS.n4390 0.019716
R55041 DVSS.n7944 DVSS.n7943 0.019716
R55042 DVSS.n7944 DVSS.n4389 0.019716
R55043 DVSS.n7937 DVSS.n7936 0.019716
R55044 DVSS.n7937 DVSS.n4388 0.019716
R55045 DVSS.n7932 DVSS.n7931 0.019716
R55046 DVSS.n7932 DVSS.n4387 0.019716
R55047 DVSS.n7925 DVSS.n7924 0.019716
R55048 DVSS.n7925 DVSS.n4386 0.019716
R55049 DVSS.n7920 DVSS.n7919 0.019716
R55050 DVSS.n7920 DVSS.n4385 0.019716
R55051 DVSS.n7913 DVSS.n7912 0.019716
R55052 DVSS.n7913 DVSS.n4384 0.019716
R55053 DVSS.n7908 DVSS.n7907 0.019716
R55054 DVSS.n7908 DVSS.n4383 0.019716
R55055 DVSS.n7901 DVSS.n7900 0.019716
R55056 DVSS.n7901 DVSS.n4382 0.019716
R55057 DVSS.n7896 DVSS.n7895 0.019716
R55058 DVSS.n7896 DVSS.n4381 0.019716
R55059 DVSS.n7889 DVSS.n7888 0.019716
R55060 DVSS.n7889 DVSS.n4380 0.019716
R55061 DVSS.n7884 DVSS.n7883 0.019716
R55062 DVSS.n7884 DVSS.n4379 0.019716
R55063 DVSS.n7877 DVSS.n7876 0.019716
R55064 DVSS.n7877 DVSS.n4378 0.019716
R55065 DVSS.n7872 DVSS.n7871 0.019716
R55066 DVSS.n7872 DVSS.n4377 0.019716
R55067 DVSS.n7865 DVSS.n7864 0.019716
R55068 DVSS.n7865 DVSS.n4376 0.019716
R55069 DVSS.n7860 DVSS.n7859 0.019716
R55070 DVSS.n7860 DVSS.n4375 0.019716
R55071 DVSS.n7853 DVSS.n7852 0.019716
R55072 DVSS.n7853 DVSS.n4374 0.019716
R55073 DVSS.n7848 DVSS.n7847 0.019716
R55074 DVSS.n7848 DVSS.n4373 0.019716
R55075 DVSS.n7841 DVSS.n4372 0.019716
R55076 DVSS.n4805 DVSS.n4804 0.019716
R55077 DVSS.n4803 DVSS.n4802 0.019716
R55078 DVSS.n4481 DVSS.n4480 0.019716
R55079 DVSS.n4480 DVSS.n4476 0.019716
R55080 DVSS.n4793 DVSS.n4792 0.019716
R55081 DVSS.n4794 DVSS.n4793 0.019716
R55082 DVSS.n4487 DVSS.n4486 0.019716
R55083 DVSS.n4486 DVSS.n4482 0.019716
R55084 DVSS.n4783 DVSS.n4782 0.019716
R55085 DVSS.n4784 DVSS.n4783 0.019716
R55086 DVSS.n4493 DVSS.n4492 0.019716
R55087 DVSS.n4492 DVSS.n4488 0.019716
R55088 DVSS.n4773 DVSS.n4772 0.019716
R55089 DVSS.n4774 DVSS.n4773 0.019716
R55090 DVSS.n4499 DVSS.n4498 0.019716
R55091 DVSS.n4498 DVSS.n4494 0.019716
R55092 DVSS.n4763 DVSS.n4762 0.019716
R55093 DVSS.n4764 DVSS.n4763 0.019716
R55094 DVSS.n4505 DVSS.n4504 0.019716
R55095 DVSS.n4504 DVSS.n4500 0.019716
R55096 DVSS.n4753 DVSS.n4752 0.019716
R55097 DVSS.n4754 DVSS.n4753 0.019716
R55098 DVSS.n4511 DVSS.n4510 0.019716
R55099 DVSS.n4510 DVSS.n4506 0.019716
R55100 DVSS.n4743 DVSS.n4742 0.019716
R55101 DVSS.n4744 DVSS.n4743 0.019716
R55102 DVSS.n4517 DVSS.n4516 0.019716
R55103 DVSS.n4516 DVSS.n4512 0.019716
R55104 DVSS.n4733 DVSS.n4732 0.019716
R55105 DVSS.n4734 DVSS.n4733 0.019716
R55106 DVSS.n4523 DVSS.n4522 0.019716
R55107 DVSS.n4522 DVSS.n4518 0.019716
R55108 DVSS.n4723 DVSS.n4722 0.019716
R55109 DVSS.n4724 DVSS.n4723 0.019716
R55110 DVSS.n4529 DVSS.n4528 0.019716
R55111 DVSS.n4528 DVSS.n4524 0.019716
R55112 DVSS.n4713 DVSS.n4712 0.019716
R55113 DVSS.n4714 DVSS.n4713 0.019716
R55114 DVSS.n4535 DVSS.n4534 0.019716
R55115 DVSS.n4534 DVSS.n4530 0.019716
R55116 DVSS.n4703 DVSS.n4702 0.019716
R55117 DVSS.n4704 DVSS.n4703 0.019716
R55118 DVSS.n4541 DVSS.n4540 0.019716
R55119 DVSS.n4540 DVSS.n4536 0.019716
R55120 DVSS.n4693 DVSS.n4692 0.019716
R55121 DVSS.n4694 DVSS.n4693 0.019716
R55122 DVSS.n4547 DVSS.n4546 0.019716
R55123 DVSS.n4546 DVSS.n4542 0.019716
R55124 DVSS.n4683 DVSS.n4682 0.019716
R55125 DVSS.n4684 DVSS.n4683 0.019716
R55126 DVSS.n4553 DVSS.n4552 0.019716
R55127 DVSS.n4552 DVSS.n4548 0.019716
R55128 DVSS.n4673 DVSS.n4672 0.019716
R55129 DVSS.n4674 DVSS.n4673 0.019716
R55130 DVSS.n4559 DVSS.n4558 0.019716
R55131 DVSS.n4558 DVSS.n4554 0.019716
R55132 DVSS.n4663 DVSS.n4662 0.019716
R55133 DVSS.n4664 DVSS.n4663 0.019716
R55134 DVSS.n4565 DVSS.n4564 0.019716
R55135 DVSS.n4564 DVSS.n4560 0.019716
R55136 DVSS.n4653 DVSS.n4652 0.019716
R55137 DVSS.n4654 DVSS.n4653 0.019716
R55138 DVSS.n4571 DVSS.n4570 0.019716
R55139 DVSS.n4570 DVSS.n4566 0.019716
R55140 DVSS.n4643 DVSS.n4642 0.019716
R55141 DVSS.n4644 DVSS.n4643 0.019716
R55142 DVSS.n4577 DVSS.n4576 0.019716
R55143 DVSS.n4576 DVSS.n4572 0.019716
R55144 DVSS.n4633 DVSS.n4632 0.019716
R55145 DVSS.n4634 DVSS.n4633 0.019716
R55146 DVSS.n4583 DVSS.n4582 0.019716
R55147 DVSS.n4582 DVSS.n4578 0.019716
R55148 DVSS.n4623 DVSS.n4622 0.019716
R55149 DVSS.n4624 DVSS.n4623 0.019716
R55150 DVSS.n4589 DVSS.n4588 0.019716
R55151 DVSS.n4588 DVSS.n4584 0.019716
R55152 DVSS.n4613 DVSS.n4612 0.019716
R55153 DVSS.n4614 DVSS.n4613 0.019716
R55154 DVSS.n4595 DVSS.n4594 0.019716
R55155 DVSS.n4594 DVSS.n4590 0.019716
R55156 DVSS.n4603 DVSS.n4602 0.019716
R55157 DVSS.n4604 DVSS.n4603 0.019716
R55158 DVSS.n4597 DVSS.n4596 0.019716
R55159 DVSS.n7794 DVSS.n7793 0.019716
R55160 DVSS.n7504 DVSS.n7503 0.019716
R55161 DVSS.n7786 DVSS.n7785 0.019716
R55162 DVSS.n7786 DVSS.n7502 0.019716
R55163 DVSS.n7781 DVSS.n7780 0.019716
R55164 DVSS.n7781 DVSS.n7501 0.019716
R55165 DVSS.n7774 DVSS.n7773 0.019716
R55166 DVSS.n7774 DVSS.n7500 0.019716
R55167 DVSS.n7769 DVSS.n7768 0.019716
R55168 DVSS.n7769 DVSS.n7499 0.019716
R55169 DVSS.n7762 DVSS.n7761 0.019716
R55170 DVSS.n7762 DVSS.n7498 0.019716
R55171 DVSS.n7757 DVSS.n7756 0.019716
R55172 DVSS.n7757 DVSS.n7497 0.019716
R55173 DVSS.n7750 DVSS.n7749 0.019716
R55174 DVSS.n7750 DVSS.n7496 0.019716
R55175 DVSS.n7745 DVSS.n7744 0.019716
R55176 DVSS.n7745 DVSS.n7495 0.019716
R55177 DVSS.n7738 DVSS.n7737 0.019716
R55178 DVSS.n7738 DVSS.n7494 0.019716
R55179 DVSS.n7733 DVSS.n7732 0.019716
R55180 DVSS.n7733 DVSS.n7493 0.019716
R55181 DVSS.n7726 DVSS.n7725 0.019716
R55182 DVSS.n7726 DVSS.n7492 0.019716
R55183 DVSS.n7721 DVSS.n7720 0.019716
R55184 DVSS.n7721 DVSS.n7491 0.019716
R55185 DVSS.n7714 DVSS.n7713 0.019716
R55186 DVSS.n7714 DVSS.n7490 0.019716
R55187 DVSS.n7709 DVSS.n7708 0.019716
R55188 DVSS.n7709 DVSS.n7489 0.019716
R55189 DVSS.n7702 DVSS.n7701 0.019716
R55190 DVSS.n7702 DVSS.n7488 0.019716
R55191 DVSS.n7697 DVSS.n7696 0.019716
R55192 DVSS.n7697 DVSS.n7487 0.019716
R55193 DVSS.n7690 DVSS.n7689 0.019716
R55194 DVSS.n7690 DVSS.n7486 0.019716
R55195 DVSS.n7685 DVSS.n7684 0.019716
R55196 DVSS.n7685 DVSS.n7485 0.019716
R55197 DVSS.n7678 DVSS.n7677 0.019716
R55198 DVSS.n7678 DVSS.n7484 0.019716
R55199 DVSS.n7673 DVSS.n7672 0.019716
R55200 DVSS.n7673 DVSS.n7483 0.019716
R55201 DVSS.n7666 DVSS.n7665 0.019716
R55202 DVSS.n7666 DVSS.n7482 0.019716
R55203 DVSS.n7661 DVSS.n7660 0.019716
R55204 DVSS.n7661 DVSS.n7481 0.019716
R55205 DVSS.n7654 DVSS.n7653 0.019716
R55206 DVSS.n7654 DVSS.n7480 0.019716
R55207 DVSS.n7649 DVSS.n7648 0.019716
R55208 DVSS.n7649 DVSS.n7479 0.019716
R55209 DVSS.n7642 DVSS.n7641 0.019716
R55210 DVSS.n7642 DVSS.n7478 0.019716
R55211 DVSS.n7637 DVSS.n7636 0.019716
R55212 DVSS.n7637 DVSS.n7477 0.019716
R55213 DVSS.n7630 DVSS.n7629 0.019716
R55214 DVSS.n7630 DVSS.n7476 0.019716
R55215 DVSS.n7625 DVSS.n7624 0.019716
R55216 DVSS.n7625 DVSS.n7475 0.019716
R55217 DVSS.n7618 DVSS.n7617 0.019716
R55218 DVSS.n7618 DVSS.n7474 0.019716
R55219 DVSS.n7613 DVSS.n7612 0.019716
R55220 DVSS.n7613 DVSS.n7473 0.019716
R55221 DVSS.n7606 DVSS.n7605 0.019716
R55222 DVSS.n7606 DVSS.n7472 0.019716
R55223 DVSS.n7601 DVSS.n7600 0.019716
R55224 DVSS.n7601 DVSS.n7471 0.019716
R55225 DVSS.n7594 DVSS.n7593 0.019716
R55226 DVSS.n7594 DVSS.n7470 0.019716
R55227 DVSS.n7589 DVSS.n7588 0.019716
R55228 DVSS.n7589 DVSS.n7469 0.019716
R55229 DVSS.n7582 DVSS.n7581 0.019716
R55230 DVSS.n7582 DVSS.n7468 0.019716
R55231 DVSS.n7577 DVSS.n7576 0.019716
R55232 DVSS.n7577 DVSS.n7467 0.019716
R55233 DVSS.n7570 DVSS.n7569 0.019716
R55234 DVSS.n7570 DVSS.n7466 0.019716
R55235 DVSS.n7565 DVSS.n7564 0.019716
R55236 DVSS.n7565 DVSS.n7465 0.019716
R55237 DVSS.n7558 DVSS.n7557 0.019716
R55238 DVSS.n7558 DVSS.n7464 0.019716
R55239 DVSS.n7553 DVSS.n7552 0.019716
R55240 DVSS.n7553 DVSS.n7463 0.019716
R55241 DVSS.n7546 DVSS.n7462 0.019716
R55242 DVSS.n7442 DVSS.n7441 0.019716
R55243 DVSS.n7440 DVSS.n7439 0.019716
R55244 DVSS.n7118 DVSS.n7117 0.019716
R55245 DVSS.n7117 DVSS.n7113 0.019716
R55246 DVSS.n7430 DVSS.n7429 0.019716
R55247 DVSS.n7431 DVSS.n7430 0.019716
R55248 DVSS.n7124 DVSS.n7123 0.019716
R55249 DVSS.n7123 DVSS.n7119 0.019716
R55250 DVSS.n7420 DVSS.n7419 0.019716
R55251 DVSS.n7421 DVSS.n7420 0.019716
R55252 DVSS.n7130 DVSS.n7129 0.019716
R55253 DVSS.n7129 DVSS.n7125 0.019716
R55254 DVSS.n7410 DVSS.n7409 0.019716
R55255 DVSS.n7411 DVSS.n7410 0.019716
R55256 DVSS.n7136 DVSS.n7135 0.019716
R55257 DVSS.n7135 DVSS.n7131 0.019716
R55258 DVSS.n7400 DVSS.n7399 0.019716
R55259 DVSS.n7401 DVSS.n7400 0.019716
R55260 DVSS.n7142 DVSS.n7141 0.019716
R55261 DVSS.n7141 DVSS.n7137 0.019716
R55262 DVSS.n7390 DVSS.n7389 0.019716
R55263 DVSS.n7391 DVSS.n7390 0.019716
R55264 DVSS.n7148 DVSS.n7147 0.019716
R55265 DVSS.n7147 DVSS.n7143 0.019716
R55266 DVSS.n7380 DVSS.n7379 0.019716
R55267 DVSS.n7381 DVSS.n7380 0.019716
R55268 DVSS.n7154 DVSS.n7153 0.019716
R55269 DVSS.n7153 DVSS.n7149 0.019716
R55270 DVSS.n7370 DVSS.n7369 0.019716
R55271 DVSS.n7371 DVSS.n7370 0.019716
R55272 DVSS.n7160 DVSS.n7159 0.019716
R55273 DVSS.n7159 DVSS.n7155 0.019716
R55274 DVSS.n7360 DVSS.n7359 0.019716
R55275 DVSS.n7361 DVSS.n7360 0.019716
R55276 DVSS.n7166 DVSS.n7165 0.019716
R55277 DVSS.n7165 DVSS.n7161 0.019716
R55278 DVSS.n7350 DVSS.n7349 0.019716
R55279 DVSS.n7351 DVSS.n7350 0.019716
R55280 DVSS.n7172 DVSS.n7171 0.019716
R55281 DVSS.n7171 DVSS.n7167 0.019716
R55282 DVSS.n7340 DVSS.n7339 0.019716
R55283 DVSS.n7341 DVSS.n7340 0.019716
R55284 DVSS.n7178 DVSS.n7177 0.019716
R55285 DVSS.n7177 DVSS.n7173 0.019716
R55286 DVSS.n7330 DVSS.n7329 0.019716
R55287 DVSS.n7331 DVSS.n7330 0.019716
R55288 DVSS.n7184 DVSS.n7183 0.019716
R55289 DVSS.n7183 DVSS.n7179 0.019716
R55290 DVSS.n7320 DVSS.n7319 0.019716
R55291 DVSS.n7321 DVSS.n7320 0.019716
R55292 DVSS.n7190 DVSS.n7189 0.019716
R55293 DVSS.n7189 DVSS.n7185 0.019716
R55294 DVSS.n7310 DVSS.n7309 0.019716
R55295 DVSS.n7311 DVSS.n7310 0.019716
R55296 DVSS.n7196 DVSS.n7195 0.019716
R55297 DVSS.n7195 DVSS.n7191 0.019716
R55298 DVSS.n7300 DVSS.n7299 0.019716
R55299 DVSS.n7301 DVSS.n7300 0.019716
R55300 DVSS.n7202 DVSS.n7201 0.019716
R55301 DVSS.n7201 DVSS.n7197 0.019716
R55302 DVSS.n7290 DVSS.n7289 0.019716
R55303 DVSS.n7291 DVSS.n7290 0.019716
R55304 DVSS.n7208 DVSS.n7207 0.019716
R55305 DVSS.n7207 DVSS.n7203 0.019716
R55306 DVSS.n7280 DVSS.n7279 0.019716
R55307 DVSS.n7281 DVSS.n7280 0.019716
R55308 DVSS.n7214 DVSS.n7213 0.019716
R55309 DVSS.n7213 DVSS.n7209 0.019716
R55310 DVSS.n7270 DVSS.n7269 0.019716
R55311 DVSS.n7271 DVSS.n7270 0.019716
R55312 DVSS.n7220 DVSS.n7219 0.019716
R55313 DVSS.n7219 DVSS.n7215 0.019716
R55314 DVSS.n7260 DVSS.n7259 0.019716
R55315 DVSS.n7261 DVSS.n7260 0.019716
R55316 DVSS.n7226 DVSS.n7225 0.019716
R55317 DVSS.n7225 DVSS.n7221 0.019716
R55318 DVSS.n7250 DVSS.n7249 0.019716
R55319 DVSS.n7251 DVSS.n7250 0.019716
R55320 DVSS.n7232 DVSS.n7231 0.019716
R55321 DVSS.n7231 DVSS.n7227 0.019716
R55322 DVSS.n7240 DVSS.n7239 0.019716
R55323 DVSS.n7241 DVSS.n7240 0.019716
R55324 DVSS.n7234 DVSS.n7233 0.019716
R55325 DVSS.n4927 DVSS.n4882 0.019716
R55326 DVSS.n4928 DVSS.n4881 0.019716
R55327 DVSS.n4937 DVSS.n4880 0.019716
R55328 DVSS.n4937 DVSS.n4936 0.019716
R55329 DVSS.n4939 DVSS.n4879 0.019716
R55330 DVSS.n4940 DVSS.n4939 0.019716
R55331 DVSS.n4949 DVSS.n4878 0.019716
R55332 DVSS.n4949 DVSS.n4948 0.019716
R55333 DVSS.n4951 DVSS.n4877 0.019716
R55334 DVSS.n4952 DVSS.n4951 0.019716
R55335 DVSS.n4961 DVSS.n4876 0.019716
R55336 DVSS.n4961 DVSS.n4960 0.019716
R55337 DVSS.n4963 DVSS.n4875 0.019716
R55338 DVSS.n4964 DVSS.n4963 0.019716
R55339 DVSS.n4973 DVSS.n4874 0.019716
R55340 DVSS.n4973 DVSS.n4972 0.019716
R55341 DVSS.n4975 DVSS.n4873 0.019716
R55342 DVSS.n4976 DVSS.n4975 0.019716
R55343 DVSS.n4985 DVSS.n4872 0.019716
R55344 DVSS.n4985 DVSS.n4984 0.019716
R55345 DVSS.n4987 DVSS.n4871 0.019716
R55346 DVSS.n4988 DVSS.n4987 0.019716
R55347 DVSS.n4997 DVSS.n4870 0.019716
R55348 DVSS.n4997 DVSS.n4996 0.019716
R55349 DVSS.n4999 DVSS.n4869 0.019716
R55350 DVSS.n5000 DVSS.n4999 0.019716
R55351 DVSS.n5009 DVSS.n4868 0.019716
R55352 DVSS.n5009 DVSS.n5008 0.019716
R55353 DVSS.n5011 DVSS.n4867 0.019716
R55354 DVSS.n5012 DVSS.n5011 0.019716
R55355 DVSS.n5021 DVSS.n4866 0.019716
R55356 DVSS.n5021 DVSS.n5020 0.019716
R55357 DVSS.n5023 DVSS.n4865 0.019716
R55358 DVSS.n5024 DVSS.n5023 0.019716
R55359 DVSS.n5033 DVSS.n4864 0.019716
R55360 DVSS.n5033 DVSS.n5032 0.019716
R55361 DVSS.n5035 DVSS.n4863 0.019716
R55362 DVSS.n5036 DVSS.n5035 0.019716
R55363 DVSS.n5045 DVSS.n4862 0.019716
R55364 DVSS.n5045 DVSS.n5044 0.019716
R55365 DVSS.n5047 DVSS.n4861 0.019716
R55366 DVSS.n5048 DVSS.n5047 0.019716
R55367 DVSS.n5057 DVSS.n4860 0.019716
R55368 DVSS.n5057 DVSS.n5056 0.019716
R55369 DVSS.n5059 DVSS.n4859 0.019716
R55370 DVSS.n5060 DVSS.n5059 0.019716
R55371 DVSS.n5069 DVSS.n4858 0.019716
R55372 DVSS.n5069 DVSS.n5068 0.019716
R55373 DVSS.n5071 DVSS.n4857 0.019716
R55374 DVSS.n5072 DVSS.n5071 0.019716
R55375 DVSS.n5081 DVSS.n4856 0.019716
R55376 DVSS.n5081 DVSS.n5080 0.019716
R55377 DVSS.n5083 DVSS.n4855 0.019716
R55378 DVSS.n5084 DVSS.n5083 0.019716
R55379 DVSS.n5093 DVSS.n4854 0.019716
R55380 DVSS.n5093 DVSS.n5092 0.019716
R55381 DVSS.n5095 DVSS.n4853 0.019716
R55382 DVSS.n5096 DVSS.n5095 0.019716
R55383 DVSS.n5105 DVSS.n4852 0.019716
R55384 DVSS.n5105 DVSS.n5104 0.019716
R55385 DVSS.n5107 DVSS.n4851 0.019716
R55386 DVSS.n5108 DVSS.n5107 0.019716
R55387 DVSS.n5117 DVSS.n4850 0.019716
R55388 DVSS.n5117 DVSS.n5116 0.019716
R55389 DVSS.n5119 DVSS.n4849 0.019716
R55390 DVSS.n5120 DVSS.n5119 0.019716
R55391 DVSS.n5129 DVSS.n4848 0.019716
R55392 DVSS.n5129 DVSS.n5128 0.019716
R55393 DVSS.n5131 DVSS.n4847 0.019716
R55394 DVSS.n5132 DVSS.n5131 0.019716
R55395 DVSS.n5141 DVSS.n4846 0.019716
R55396 DVSS.n5141 DVSS.n5140 0.019716
R55397 DVSS.n5143 DVSS.n4845 0.019716
R55398 DVSS.n5144 DVSS.n5143 0.019716
R55399 DVSS.n5153 DVSS.n4844 0.019716
R55400 DVSS.n5153 DVSS.n5152 0.019716
R55401 DVSS.n5155 DVSS.n4843 0.019716
R55402 DVSS.n5156 DVSS.n5155 0.019716
R55403 DVSS.n5165 DVSS.n4842 0.019716
R55404 DVSS.n5165 DVSS.n5164 0.019716
R55405 DVSS.n5167 DVSS.n4841 0.019716
R55406 DVSS.n5168 DVSS.n5167 0.019716
R55407 DVSS.n7101 DVSS.n7100 0.019716
R55408 DVSS.n5273 DVSS.n5272 0.019716
R55409 DVSS.n5275 DVSS.n5274 0.019716
R55410 DVSS.n5276 DVSS.n5266 0.019716
R55411 DVSS.n5277 DVSS.n5276 0.019716
R55412 DVSS.n5287 DVSS.n5286 0.019716
R55413 DVSS.n5286 DVSS.n5285 0.019716
R55414 DVSS.n5288 DVSS.n5262 0.019716
R55415 DVSS.n5289 DVSS.n5288 0.019716
R55416 DVSS.n5299 DVSS.n5298 0.019716
R55417 DVSS.n5298 DVSS.n5297 0.019716
R55418 DVSS.n5300 DVSS.n5258 0.019716
R55419 DVSS.n5301 DVSS.n5300 0.019716
R55420 DVSS.n5311 DVSS.n5310 0.019716
R55421 DVSS.n5310 DVSS.n5309 0.019716
R55422 DVSS.n5312 DVSS.n5254 0.019716
R55423 DVSS.n5313 DVSS.n5312 0.019716
R55424 DVSS.n5323 DVSS.n5322 0.019716
R55425 DVSS.n5322 DVSS.n5321 0.019716
R55426 DVSS.n5324 DVSS.n5250 0.019716
R55427 DVSS.n5325 DVSS.n5324 0.019716
R55428 DVSS.n5335 DVSS.n5334 0.019716
R55429 DVSS.n5334 DVSS.n5333 0.019716
R55430 DVSS.n5336 DVSS.n5246 0.019716
R55431 DVSS.n5337 DVSS.n5336 0.019716
R55432 DVSS.n5347 DVSS.n5346 0.019716
R55433 DVSS.n5346 DVSS.n5345 0.019716
R55434 DVSS.n5348 DVSS.n5242 0.019716
R55435 DVSS.n5349 DVSS.n5348 0.019716
R55436 DVSS.n5359 DVSS.n5358 0.019716
R55437 DVSS.n5358 DVSS.n5357 0.019716
R55438 DVSS.n5360 DVSS.n5238 0.019716
R55439 DVSS.n5361 DVSS.n5360 0.019716
R55440 DVSS.n5371 DVSS.n5370 0.019716
R55441 DVSS.n5370 DVSS.n5369 0.019716
R55442 DVSS.n5372 DVSS.n5234 0.019716
R55443 DVSS.n5373 DVSS.n5372 0.019716
R55444 DVSS.n5383 DVSS.n5382 0.019716
R55445 DVSS.n5382 DVSS.n5381 0.019716
R55446 DVSS.n5384 DVSS.n5230 0.019716
R55447 DVSS.n5385 DVSS.n5384 0.019716
R55448 DVSS.n5395 DVSS.n5394 0.019716
R55449 DVSS.n5394 DVSS.n5393 0.019716
R55450 DVSS.n5396 DVSS.n5226 0.019716
R55451 DVSS.n5397 DVSS.n5396 0.019716
R55452 DVSS.n5407 DVSS.n5406 0.019716
R55453 DVSS.n5406 DVSS.n5405 0.019716
R55454 DVSS.n5408 DVSS.n5222 0.019716
R55455 DVSS.n5409 DVSS.n5408 0.019716
R55456 DVSS.n5419 DVSS.n5418 0.019716
R55457 DVSS.n5418 DVSS.n5417 0.019716
R55458 DVSS.n5420 DVSS.n5218 0.019716
R55459 DVSS.n5421 DVSS.n5420 0.019716
R55460 DVSS.n5431 DVSS.n5430 0.019716
R55461 DVSS.n5430 DVSS.n5429 0.019716
R55462 DVSS.n5432 DVSS.n5214 0.019716
R55463 DVSS.n5433 DVSS.n5432 0.019716
R55464 DVSS.n5443 DVSS.n5442 0.019716
R55465 DVSS.n5442 DVSS.n5441 0.019716
R55466 DVSS.n5444 DVSS.n5210 0.019716
R55467 DVSS.n5445 DVSS.n5444 0.019716
R55468 DVSS.n5455 DVSS.n5454 0.019716
R55469 DVSS.n5454 DVSS.n5453 0.019716
R55470 DVSS.n5456 DVSS.n5206 0.019716
R55471 DVSS.n5457 DVSS.n5456 0.019716
R55472 DVSS.n5467 DVSS.n5466 0.019716
R55473 DVSS.n5466 DVSS.n5465 0.019716
R55474 DVSS.n5468 DVSS.n5202 0.019716
R55475 DVSS.n5469 DVSS.n5468 0.019716
R55476 DVSS.n5479 DVSS.n5478 0.019716
R55477 DVSS.n5478 DVSS.n5477 0.019716
R55478 DVSS.n5480 DVSS.n5198 0.019716
R55479 DVSS.n5481 DVSS.n5480 0.019716
R55480 DVSS.n5491 DVSS.n5490 0.019716
R55481 DVSS.n5490 DVSS.n5489 0.019716
R55482 DVSS.n5492 DVSS.n5194 0.019716
R55483 DVSS.n5493 DVSS.n5492 0.019716
R55484 DVSS.n5503 DVSS.n5502 0.019716
R55485 DVSS.n5502 DVSS.n5501 0.019716
R55486 DVSS.n5504 DVSS.n5190 0.019716
R55487 DVSS.n5505 DVSS.n5504 0.019716
R55488 DVSS.n5516 DVSS.n5515 0.019716
R55489 DVSS.n5515 DVSS.n5514 0.019716
R55490 DVSS.n5519 DVSS.n5518 0.019716
R55491 DVSS.n5618 DVSS.n5573 0.019716
R55492 DVSS.n5619 DVSS.n5572 0.019716
R55493 DVSS.n5628 DVSS.n5571 0.019716
R55494 DVSS.n5628 DVSS.n5627 0.019716
R55495 DVSS.n5630 DVSS.n5570 0.019716
R55496 DVSS.n5631 DVSS.n5630 0.019716
R55497 DVSS.n5640 DVSS.n5569 0.019716
R55498 DVSS.n5640 DVSS.n5639 0.019716
R55499 DVSS.n5642 DVSS.n5568 0.019716
R55500 DVSS.n5643 DVSS.n5642 0.019716
R55501 DVSS.n5652 DVSS.n5567 0.019716
R55502 DVSS.n5652 DVSS.n5651 0.019716
R55503 DVSS.n5654 DVSS.n5566 0.019716
R55504 DVSS.n5655 DVSS.n5654 0.019716
R55505 DVSS.n5664 DVSS.n5565 0.019716
R55506 DVSS.n5664 DVSS.n5663 0.019716
R55507 DVSS.n5666 DVSS.n5564 0.019716
R55508 DVSS.n5667 DVSS.n5666 0.019716
R55509 DVSS.n5676 DVSS.n5563 0.019716
R55510 DVSS.n5676 DVSS.n5675 0.019716
R55511 DVSS.n5678 DVSS.n5562 0.019716
R55512 DVSS.n5679 DVSS.n5678 0.019716
R55513 DVSS.n5688 DVSS.n5561 0.019716
R55514 DVSS.n5688 DVSS.n5687 0.019716
R55515 DVSS.n5690 DVSS.n5560 0.019716
R55516 DVSS.n5691 DVSS.n5690 0.019716
R55517 DVSS.n5700 DVSS.n5559 0.019716
R55518 DVSS.n5700 DVSS.n5699 0.019716
R55519 DVSS.n5702 DVSS.n5558 0.019716
R55520 DVSS.n5703 DVSS.n5702 0.019716
R55521 DVSS.n5712 DVSS.n5557 0.019716
R55522 DVSS.n5712 DVSS.n5711 0.019716
R55523 DVSS.n5714 DVSS.n5556 0.019716
R55524 DVSS.n5715 DVSS.n5714 0.019716
R55525 DVSS.n5724 DVSS.n5555 0.019716
R55526 DVSS.n5724 DVSS.n5723 0.019716
R55527 DVSS.n5726 DVSS.n5554 0.019716
R55528 DVSS.n5727 DVSS.n5726 0.019716
R55529 DVSS.n5736 DVSS.n5553 0.019716
R55530 DVSS.n5736 DVSS.n5735 0.019716
R55531 DVSS.n5738 DVSS.n5552 0.019716
R55532 DVSS.n5739 DVSS.n5738 0.019716
R55533 DVSS.n5748 DVSS.n5551 0.019716
R55534 DVSS.n5748 DVSS.n5747 0.019716
R55535 DVSS.n5750 DVSS.n5550 0.019716
R55536 DVSS.n5751 DVSS.n5750 0.019716
R55537 DVSS.n5760 DVSS.n5549 0.019716
R55538 DVSS.n5760 DVSS.n5759 0.019716
R55539 DVSS.n5762 DVSS.n5548 0.019716
R55540 DVSS.n5763 DVSS.n5762 0.019716
R55541 DVSS.n5772 DVSS.n5547 0.019716
R55542 DVSS.n5772 DVSS.n5771 0.019716
R55543 DVSS.n5774 DVSS.n5546 0.019716
R55544 DVSS.n5775 DVSS.n5774 0.019716
R55545 DVSS.n5784 DVSS.n5545 0.019716
R55546 DVSS.n5784 DVSS.n5783 0.019716
R55547 DVSS.n5786 DVSS.n5544 0.019716
R55548 DVSS.n5787 DVSS.n5786 0.019716
R55549 DVSS.n5796 DVSS.n5543 0.019716
R55550 DVSS.n5796 DVSS.n5795 0.019716
R55551 DVSS.n5798 DVSS.n5542 0.019716
R55552 DVSS.n5799 DVSS.n5798 0.019716
R55553 DVSS.n5808 DVSS.n5541 0.019716
R55554 DVSS.n5808 DVSS.n5807 0.019716
R55555 DVSS.n5810 DVSS.n5540 0.019716
R55556 DVSS.n5811 DVSS.n5810 0.019716
R55557 DVSS.n5820 DVSS.n5539 0.019716
R55558 DVSS.n5820 DVSS.n5819 0.019716
R55559 DVSS.n5822 DVSS.n5538 0.019716
R55560 DVSS.n5823 DVSS.n5822 0.019716
R55561 DVSS.n5832 DVSS.n5537 0.019716
R55562 DVSS.n5832 DVSS.n5831 0.019716
R55563 DVSS.n5834 DVSS.n5536 0.019716
R55564 DVSS.n5835 DVSS.n5834 0.019716
R55565 DVSS.n5844 DVSS.n5535 0.019716
R55566 DVSS.n5844 DVSS.n5843 0.019716
R55567 DVSS.n5846 DVSS.n5534 0.019716
R55568 DVSS.n5847 DVSS.n5846 0.019716
R55569 DVSS.n5856 DVSS.n5533 0.019716
R55570 DVSS.n5856 DVSS.n5855 0.019716
R55571 DVSS.n5858 DVSS.n5532 0.019716
R55572 DVSS.n5859 DVSS.n5858 0.019716
R55573 DVSS.n7058 DVSS.n7057 0.019716
R55574 DVSS.n6781 DVSS.n6776 0.019716
R55575 DVSS.n6782 DVSS.n6781 0.019716
R55576 DVSS.n6787 DVSS.n6784 0.019716
R55577 DVSS.n6787 DVSS.n6786 0.019716
R55578 DVSS.n6793 DVSS.n6772 0.019716
R55579 DVSS.n6794 DVSS.n6793 0.019716
R55580 DVSS.n6799 DVSS.n6796 0.019716
R55581 DVSS.n6799 DVSS.n6798 0.019716
R55582 DVSS.n6805 DVSS.n6768 0.019716
R55583 DVSS.n6806 DVSS.n6805 0.019716
R55584 DVSS.n6811 DVSS.n6808 0.019716
R55585 DVSS.n6811 DVSS.n6810 0.019716
R55586 DVSS.n6817 DVSS.n6764 0.019716
R55587 DVSS.n6818 DVSS.n6817 0.019716
R55588 DVSS.n6823 DVSS.n6820 0.019716
R55589 DVSS.n6823 DVSS.n6822 0.019716
R55590 DVSS.n6829 DVSS.n6760 0.019716
R55591 DVSS.n6830 DVSS.n6829 0.019716
R55592 DVSS.n6835 DVSS.n6832 0.019716
R55593 DVSS.n6835 DVSS.n6834 0.019716
R55594 DVSS.n6841 DVSS.n6756 0.019716
R55595 DVSS.n6842 DVSS.n6841 0.019716
R55596 DVSS.n6847 DVSS.n6844 0.019716
R55597 DVSS.n6847 DVSS.n6846 0.019716
R55598 DVSS.n6853 DVSS.n6752 0.019716
R55599 DVSS.n6854 DVSS.n6853 0.019716
R55600 DVSS.n6859 DVSS.n6856 0.019716
R55601 DVSS.n6859 DVSS.n6858 0.019716
R55602 DVSS.n6865 DVSS.n6748 0.019716
R55603 DVSS.n6866 DVSS.n6865 0.019716
R55604 DVSS.n6871 DVSS.n6868 0.019716
R55605 DVSS.n6871 DVSS.n6870 0.019716
R55606 DVSS.n6877 DVSS.n6744 0.019716
R55607 DVSS.n6878 DVSS.n6877 0.019716
R55608 DVSS.n6883 DVSS.n6880 0.019716
R55609 DVSS.n6883 DVSS.n6882 0.019716
R55610 DVSS.n6889 DVSS.n6740 0.019716
R55611 DVSS.n6890 DVSS.n6889 0.019716
R55612 DVSS.n6895 DVSS.n6892 0.019716
R55613 DVSS.n6895 DVSS.n6894 0.019716
R55614 DVSS.n6901 DVSS.n6736 0.019716
R55615 DVSS.n6902 DVSS.n6901 0.019716
R55616 DVSS.n6907 DVSS.n6904 0.019716
R55617 DVSS.n6907 DVSS.n6906 0.019716
R55618 DVSS.n6913 DVSS.n6732 0.019716
R55619 DVSS.n6914 DVSS.n6913 0.019716
R55620 DVSS.n6919 DVSS.n6916 0.019716
R55621 DVSS.n6919 DVSS.n6918 0.019716
R55622 DVSS.n6925 DVSS.n6728 0.019716
R55623 DVSS.n6926 DVSS.n6925 0.019716
R55624 DVSS.n6931 DVSS.n6928 0.019716
R55625 DVSS.n6931 DVSS.n6930 0.019716
R55626 DVSS.n6937 DVSS.n6724 0.019716
R55627 DVSS.n6938 DVSS.n6937 0.019716
R55628 DVSS.n6943 DVSS.n6940 0.019716
R55629 DVSS.n6943 DVSS.n6942 0.019716
R55630 DVSS.n6949 DVSS.n6720 0.019716
R55631 DVSS.n6950 DVSS.n6949 0.019716
R55632 DVSS.n6955 DVSS.n6952 0.019716
R55633 DVSS.n6955 DVSS.n6954 0.019716
R55634 DVSS.n6961 DVSS.n6716 0.019716
R55635 DVSS.n6962 DVSS.n6961 0.019716
R55636 DVSS.n6967 DVSS.n6964 0.019716
R55637 DVSS.n6967 DVSS.n6966 0.019716
R55638 DVSS.n6973 DVSS.n6712 0.019716
R55639 DVSS.n6974 DVSS.n6973 0.019716
R55640 DVSS.n6979 DVSS.n6976 0.019716
R55641 DVSS.n6979 DVSS.n6978 0.019716
R55642 DVSS.n6985 DVSS.n6708 0.019716
R55643 DVSS.n6986 DVSS.n6985 0.019716
R55644 DVSS.n6991 DVSS.n6988 0.019716
R55645 DVSS.n6991 DVSS.n6990 0.019716
R55646 DVSS.n6997 DVSS.n6704 0.019716
R55647 DVSS.n6998 DVSS.n6997 0.019716
R55648 DVSS.n7003 DVSS.n7000 0.019716
R55649 DVSS.n7003 DVSS.n7002 0.019716
R55650 DVSS.n7009 DVSS.n6700 0.019716
R55651 DVSS.n7010 DVSS.n7009 0.019716
R55652 DVSS.n7015 DVSS.n7012 0.019716
R55653 DVSS.n7015 DVSS.n7014 0.019716
R55654 DVSS.n7021 DVSS.n6696 0.019716
R55655 DVSS.n7022 DVSS.n7021 0.019716
R55656 DVSS.n7025 DVSS.n7024 0.019716
R55657 DVSS.n6777 DVSS.n6776 0.019716
R55658 DVSS.n6784 DVSS.n6783 0.019716
R55659 DVSS.n6783 DVSS.n6782 0.019716
R55660 DVSS.n6785 DVSS.n6772 0.019716
R55661 DVSS.n6786 DVSS.n6785 0.019716
R55662 DVSS.n6796 DVSS.n6795 0.019716
R55663 DVSS.n6795 DVSS.n6794 0.019716
R55664 DVSS.n6797 DVSS.n6768 0.019716
R55665 DVSS.n6798 DVSS.n6797 0.019716
R55666 DVSS.n6808 DVSS.n6807 0.019716
R55667 DVSS.n6807 DVSS.n6806 0.019716
R55668 DVSS.n6809 DVSS.n6764 0.019716
R55669 DVSS.n6810 DVSS.n6809 0.019716
R55670 DVSS.n6820 DVSS.n6819 0.019716
R55671 DVSS.n6819 DVSS.n6818 0.019716
R55672 DVSS.n6821 DVSS.n6760 0.019716
R55673 DVSS.n6822 DVSS.n6821 0.019716
R55674 DVSS.n6832 DVSS.n6831 0.019716
R55675 DVSS.n6831 DVSS.n6830 0.019716
R55676 DVSS.n6833 DVSS.n6756 0.019716
R55677 DVSS.n6834 DVSS.n6833 0.019716
R55678 DVSS.n6844 DVSS.n6843 0.019716
R55679 DVSS.n6843 DVSS.n6842 0.019716
R55680 DVSS.n6845 DVSS.n6752 0.019716
R55681 DVSS.n6846 DVSS.n6845 0.019716
R55682 DVSS.n6856 DVSS.n6855 0.019716
R55683 DVSS.n6855 DVSS.n6854 0.019716
R55684 DVSS.n6857 DVSS.n6748 0.019716
R55685 DVSS.n6858 DVSS.n6857 0.019716
R55686 DVSS.n6868 DVSS.n6867 0.019716
R55687 DVSS.n6867 DVSS.n6866 0.019716
R55688 DVSS.n6869 DVSS.n6744 0.019716
R55689 DVSS.n6870 DVSS.n6869 0.019716
R55690 DVSS.n6880 DVSS.n6879 0.019716
R55691 DVSS.n6879 DVSS.n6878 0.019716
R55692 DVSS.n6881 DVSS.n6740 0.019716
R55693 DVSS.n6882 DVSS.n6881 0.019716
R55694 DVSS.n6892 DVSS.n6891 0.019716
R55695 DVSS.n6891 DVSS.n6890 0.019716
R55696 DVSS.n6893 DVSS.n6736 0.019716
R55697 DVSS.n6894 DVSS.n6893 0.019716
R55698 DVSS.n6904 DVSS.n6903 0.019716
R55699 DVSS.n6903 DVSS.n6902 0.019716
R55700 DVSS.n6905 DVSS.n6732 0.019716
R55701 DVSS.n6906 DVSS.n6905 0.019716
R55702 DVSS.n6916 DVSS.n6915 0.019716
R55703 DVSS.n6915 DVSS.n6914 0.019716
R55704 DVSS.n6917 DVSS.n6728 0.019716
R55705 DVSS.n6918 DVSS.n6917 0.019716
R55706 DVSS.n6928 DVSS.n6927 0.019716
R55707 DVSS.n6927 DVSS.n6926 0.019716
R55708 DVSS.n6929 DVSS.n6724 0.019716
R55709 DVSS.n6930 DVSS.n6929 0.019716
R55710 DVSS.n6940 DVSS.n6939 0.019716
R55711 DVSS.n6939 DVSS.n6938 0.019716
R55712 DVSS.n6941 DVSS.n6720 0.019716
R55713 DVSS.n6942 DVSS.n6941 0.019716
R55714 DVSS.n6952 DVSS.n6951 0.019716
R55715 DVSS.n6951 DVSS.n6950 0.019716
R55716 DVSS.n6953 DVSS.n6716 0.019716
R55717 DVSS.n6954 DVSS.n6953 0.019716
R55718 DVSS.n6964 DVSS.n6963 0.019716
R55719 DVSS.n6963 DVSS.n6962 0.019716
R55720 DVSS.n6965 DVSS.n6712 0.019716
R55721 DVSS.n6966 DVSS.n6965 0.019716
R55722 DVSS.n6976 DVSS.n6975 0.019716
R55723 DVSS.n6975 DVSS.n6974 0.019716
R55724 DVSS.n6977 DVSS.n6708 0.019716
R55725 DVSS.n6978 DVSS.n6977 0.019716
R55726 DVSS.n6988 DVSS.n6987 0.019716
R55727 DVSS.n6987 DVSS.n6986 0.019716
R55728 DVSS.n6989 DVSS.n6704 0.019716
R55729 DVSS.n6990 DVSS.n6989 0.019716
R55730 DVSS.n7000 DVSS.n6999 0.019716
R55731 DVSS.n6999 DVSS.n6998 0.019716
R55732 DVSS.n7001 DVSS.n6700 0.019716
R55733 DVSS.n7002 DVSS.n7001 0.019716
R55734 DVSS.n7012 DVSS.n7011 0.019716
R55735 DVSS.n7011 DVSS.n7010 0.019716
R55736 DVSS.n7013 DVSS.n6696 0.019716
R55737 DVSS.n7014 DVSS.n7013 0.019716
R55738 DVSS.n7024 DVSS.n7023 0.019716
R55739 DVSS.n7023 DVSS.n7022 0.019716
R55740 DVSS.n12088 DVSS.n12044 0.019716
R55741 DVSS.n12094 DVSS.n12043 0.019716
R55742 DVSS.n12095 DVSS.n12094 0.019716
R55743 DVSS.n12100 DVSS.n12042 0.019716
R55744 DVSS.n12100 DVSS.n12099 0.019716
R55745 DVSS.n12106 DVSS.n12041 0.019716
R55746 DVSS.n12107 DVSS.n12106 0.019716
R55747 DVSS.n12112 DVSS.n12040 0.019716
R55748 DVSS.n12112 DVSS.n12111 0.019716
R55749 DVSS.n12118 DVSS.n12039 0.019716
R55750 DVSS.n12119 DVSS.n12118 0.019716
R55751 DVSS.n12124 DVSS.n12038 0.019716
R55752 DVSS.n12124 DVSS.n12123 0.019716
R55753 DVSS.n12130 DVSS.n12037 0.019716
R55754 DVSS.n12131 DVSS.n12130 0.019716
R55755 DVSS.n12136 DVSS.n12036 0.019716
R55756 DVSS.n12136 DVSS.n12135 0.019716
R55757 DVSS.n12142 DVSS.n12035 0.019716
R55758 DVSS.n12143 DVSS.n12142 0.019716
R55759 DVSS.n12148 DVSS.n12034 0.019716
R55760 DVSS.n12148 DVSS.n12147 0.019716
R55761 DVSS.n12154 DVSS.n12033 0.019716
R55762 DVSS.n12155 DVSS.n12154 0.019716
R55763 DVSS.n12160 DVSS.n12032 0.019716
R55764 DVSS.n12160 DVSS.n12159 0.019716
R55765 DVSS.n12166 DVSS.n12031 0.019716
R55766 DVSS.n12167 DVSS.n12166 0.019716
R55767 DVSS.n12172 DVSS.n12030 0.019716
R55768 DVSS.n12172 DVSS.n12171 0.019716
R55769 DVSS.n12178 DVSS.n12029 0.019716
R55770 DVSS.n12179 DVSS.n12178 0.019716
R55771 DVSS.n12184 DVSS.n12028 0.019716
R55772 DVSS.n12184 DVSS.n12183 0.019716
R55773 DVSS.n12190 DVSS.n12027 0.019716
R55774 DVSS.n12191 DVSS.n12190 0.019716
R55775 DVSS.n12196 DVSS.n12026 0.019716
R55776 DVSS.n12196 DVSS.n12195 0.019716
R55777 DVSS.n12202 DVSS.n12025 0.019716
R55778 DVSS.n12203 DVSS.n12202 0.019716
R55779 DVSS.n12208 DVSS.n12024 0.019716
R55780 DVSS.n12208 DVSS.n12207 0.019716
R55781 DVSS.n12214 DVSS.n12023 0.019716
R55782 DVSS.n12215 DVSS.n12214 0.019716
R55783 DVSS.n12220 DVSS.n12022 0.019716
R55784 DVSS.n12220 DVSS.n12219 0.019716
R55785 DVSS.n12226 DVSS.n12021 0.019716
R55786 DVSS.n12227 DVSS.n12226 0.019716
R55787 DVSS.n12232 DVSS.n12020 0.019716
R55788 DVSS.n12232 DVSS.n12231 0.019716
R55789 DVSS.n12238 DVSS.n12019 0.019716
R55790 DVSS.n12239 DVSS.n12238 0.019716
R55791 DVSS.n12244 DVSS.n12018 0.019716
R55792 DVSS.n12244 DVSS.n12243 0.019716
R55793 DVSS.n12250 DVSS.n12017 0.019716
R55794 DVSS.n12251 DVSS.n12250 0.019716
R55795 DVSS.n12256 DVSS.n12016 0.019716
R55796 DVSS.n12256 DVSS.n12255 0.019716
R55797 DVSS.n12262 DVSS.n12015 0.019716
R55798 DVSS.n12263 DVSS.n12262 0.019716
R55799 DVSS.n12268 DVSS.n12014 0.019716
R55800 DVSS.n12268 DVSS.n12267 0.019716
R55801 DVSS.n12274 DVSS.n12013 0.019716
R55802 DVSS.n12275 DVSS.n12274 0.019716
R55803 DVSS.n12280 DVSS.n12012 0.019716
R55804 DVSS.n12280 DVSS.n12279 0.019716
R55805 DVSS.n12286 DVSS.n12011 0.019716
R55806 DVSS.n12287 DVSS.n12286 0.019716
R55807 DVSS.n12292 DVSS.n12010 0.019716
R55808 DVSS.n12292 DVSS.n12291 0.019716
R55809 DVSS.n12298 DVSS.n12009 0.019716
R55810 DVSS.n12299 DVSS.n12298 0.019716
R55811 DVSS.n12304 DVSS.n12008 0.019716
R55812 DVSS.n12304 DVSS.n12303 0.019716
R55813 DVSS.n12310 DVSS.n12007 0.019716
R55814 DVSS.n12311 DVSS.n12310 0.019716
R55815 DVSS.n12316 DVSS.n12006 0.019716
R55816 DVSS.n12316 DVSS.n12315 0.019716
R55817 DVSS.n12322 DVSS.n12005 0.019716
R55818 DVSS.n12323 DVSS.n12322 0.019716
R55819 DVSS.n12328 DVSS.n12004 0.019716
R55820 DVSS.n12328 DVSS.n12327 0.019716
R55821 DVSS.n12047 DVSS.n12003 0.019716
R55822 DVSS.n12047 DVSS.n12045 0.019716
R55823 DVSS.n12089 DVSS.n12043 0.019716
R55824 DVSS.n12089 DVSS.n12088 0.019716
R55825 DVSS.n12096 DVSS.n12042 0.019716
R55826 DVSS.n12096 DVSS.n12095 0.019716
R55827 DVSS.n12098 DVSS.n12041 0.019716
R55828 DVSS.n12099 DVSS.n12098 0.019716
R55829 DVSS.n12108 DVSS.n12040 0.019716
R55830 DVSS.n12108 DVSS.n12107 0.019716
R55831 DVSS.n12110 DVSS.n12039 0.019716
R55832 DVSS.n12111 DVSS.n12110 0.019716
R55833 DVSS.n12120 DVSS.n12038 0.019716
R55834 DVSS.n12120 DVSS.n12119 0.019716
R55835 DVSS.n12122 DVSS.n12037 0.019716
R55836 DVSS.n12123 DVSS.n12122 0.019716
R55837 DVSS.n12132 DVSS.n12036 0.019716
R55838 DVSS.n12132 DVSS.n12131 0.019716
R55839 DVSS.n12134 DVSS.n12035 0.019716
R55840 DVSS.n12135 DVSS.n12134 0.019716
R55841 DVSS.n12144 DVSS.n12034 0.019716
R55842 DVSS.n12144 DVSS.n12143 0.019716
R55843 DVSS.n12146 DVSS.n12033 0.019716
R55844 DVSS.n12147 DVSS.n12146 0.019716
R55845 DVSS.n12156 DVSS.n12032 0.019716
R55846 DVSS.n12156 DVSS.n12155 0.019716
R55847 DVSS.n12158 DVSS.n12031 0.019716
R55848 DVSS.n12159 DVSS.n12158 0.019716
R55849 DVSS.n12168 DVSS.n12030 0.019716
R55850 DVSS.n12168 DVSS.n12167 0.019716
R55851 DVSS.n12170 DVSS.n12029 0.019716
R55852 DVSS.n12171 DVSS.n12170 0.019716
R55853 DVSS.n12180 DVSS.n12028 0.019716
R55854 DVSS.n12180 DVSS.n12179 0.019716
R55855 DVSS.n12182 DVSS.n12027 0.019716
R55856 DVSS.n12183 DVSS.n12182 0.019716
R55857 DVSS.n12192 DVSS.n12026 0.019716
R55858 DVSS.n12192 DVSS.n12191 0.019716
R55859 DVSS.n12194 DVSS.n12025 0.019716
R55860 DVSS.n12195 DVSS.n12194 0.019716
R55861 DVSS.n12204 DVSS.n12024 0.019716
R55862 DVSS.n12204 DVSS.n12203 0.019716
R55863 DVSS.n12206 DVSS.n12023 0.019716
R55864 DVSS.n12207 DVSS.n12206 0.019716
R55865 DVSS.n12216 DVSS.n12022 0.019716
R55866 DVSS.n12216 DVSS.n12215 0.019716
R55867 DVSS.n12218 DVSS.n12021 0.019716
R55868 DVSS.n12219 DVSS.n12218 0.019716
R55869 DVSS.n12228 DVSS.n12020 0.019716
R55870 DVSS.n12228 DVSS.n12227 0.019716
R55871 DVSS.n12230 DVSS.n12019 0.019716
R55872 DVSS.n12231 DVSS.n12230 0.019716
R55873 DVSS.n12240 DVSS.n12018 0.019716
R55874 DVSS.n12240 DVSS.n12239 0.019716
R55875 DVSS.n12242 DVSS.n12017 0.019716
R55876 DVSS.n12243 DVSS.n12242 0.019716
R55877 DVSS.n12252 DVSS.n12016 0.019716
R55878 DVSS.n12252 DVSS.n12251 0.019716
R55879 DVSS.n12254 DVSS.n12015 0.019716
R55880 DVSS.n12255 DVSS.n12254 0.019716
R55881 DVSS.n12264 DVSS.n12014 0.019716
R55882 DVSS.n12264 DVSS.n12263 0.019716
R55883 DVSS.n12266 DVSS.n12013 0.019716
R55884 DVSS.n12267 DVSS.n12266 0.019716
R55885 DVSS.n12276 DVSS.n12012 0.019716
R55886 DVSS.n12276 DVSS.n12275 0.019716
R55887 DVSS.n12278 DVSS.n12011 0.019716
R55888 DVSS.n12279 DVSS.n12278 0.019716
R55889 DVSS.n12288 DVSS.n12010 0.019716
R55890 DVSS.n12288 DVSS.n12287 0.019716
R55891 DVSS.n12290 DVSS.n12009 0.019716
R55892 DVSS.n12291 DVSS.n12290 0.019716
R55893 DVSS.n12300 DVSS.n12008 0.019716
R55894 DVSS.n12300 DVSS.n12299 0.019716
R55895 DVSS.n12302 DVSS.n12007 0.019716
R55896 DVSS.n12303 DVSS.n12302 0.019716
R55897 DVSS.n12312 DVSS.n12006 0.019716
R55898 DVSS.n12312 DVSS.n12311 0.019716
R55899 DVSS.n12314 DVSS.n12005 0.019716
R55900 DVSS.n12315 DVSS.n12314 0.019716
R55901 DVSS.n12324 DVSS.n12004 0.019716
R55902 DVSS.n12324 DVSS.n12323 0.019716
R55903 DVSS.n12326 DVSS.n12003 0.019716
R55904 DVSS.n12327 DVSS.n12326 0.019716
R55905 DVSS.n12335 DVSS.n12045 0.019716
R55906 DVSS.n6230 DVSS.n5938 0.019716
R55907 DVSS.n5941 DVSS.n5939 0.019716
R55908 DVSS.n5941 DVSS.n5937 0.019716
R55909 DVSS.n6222 DVSS.n6221 0.019716
R55910 DVSS.n6221 DVSS.n5936 0.019716
R55911 DVSS.n6217 DVSS.n6216 0.019716
R55912 DVSS.n6216 DVSS.n5935 0.019716
R55913 DVSS.n6210 DVSS.n6209 0.019716
R55914 DVSS.n6209 DVSS.n5934 0.019716
R55915 DVSS.n6205 DVSS.n6204 0.019716
R55916 DVSS.n6204 DVSS.n5933 0.019716
R55917 DVSS.n6198 DVSS.n6197 0.019716
R55918 DVSS.n6197 DVSS.n5932 0.019716
R55919 DVSS.n6193 DVSS.n6192 0.019716
R55920 DVSS.n6192 DVSS.n5931 0.019716
R55921 DVSS.n6186 DVSS.n6185 0.019716
R55922 DVSS.n6185 DVSS.n5930 0.019716
R55923 DVSS.n6181 DVSS.n6180 0.019716
R55924 DVSS.n6180 DVSS.n5929 0.019716
R55925 DVSS.n6174 DVSS.n6173 0.019716
R55926 DVSS.n6173 DVSS.n5928 0.019716
R55927 DVSS.n6169 DVSS.n6168 0.019716
R55928 DVSS.n6168 DVSS.n5927 0.019716
R55929 DVSS.n6162 DVSS.n6161 0.019716
R55930 DVSS.n6161 DVSS.n5926 0.019716
R55931 DVSS.n6157 DVSS.n6156 0.019716
R55932 DVSS.n6156 DVSS.n5925 0.019716
R55933 DVSS.n6150 DVSS.n6149 0.019716
R55934 DVSS.n6149 DVSS.n5924 0.019716
R55935 DVSS.n6145 DVSS.n6144 0.019716
R55936 DVSS.n6144 DVSS.n5923 0.019716
R55937 DVSS.n6138 DVSS.n6137 0.019716
R55938 DVSS.n6137 DVSS.n5922 0.019716
R55939 DVSS.n6133 DVSS.n6132 0.019716
R55940 DVSS.n6132 DVSS.n5921 0.019716
R55941 DVSS.n6126 DVSS.n6125 0.019716
R55942 DVSS.n6125 DVSS.n5920 0.019716
R55943 DVSS.n6121 DVSS.n6120 0.019716
R55944 DVSS.n6120 DVSS.n5919 0.019716
R55945 DVSS.n6114 DVSS.n6113 0.019716
R55946 DVSS.n6113 DVSS.n5918 0.019716
R55947 DVSS.n6109 DVSS.n6108 0.019716
R55948 DVSS.n6108 DVSS.n5917 0.019716
R55949 DVSS.n6102 DVSS.n6101 0.019716
R55950 DVSS.n6101 DVSS.n5916 0.019716
R55951 DVSS.n6097 DVSS.n6096 0.019716
R55952 DVSS.n6096 DVSS.n5915 0.019716
R55953 DVSS.n6090 DVSS.n6089 0.019716
R55954 DVSS.n6089 DVSS.n5914 0.019716
R55955 DVSS.n6085 DVSS.n6084 0.019716
R55956 DVSS.n6084 DVSS.n5913 0.019716
R55957 DVSS.n6078 DVSS.n6077 0.019716
R55958 DVSS.n6077 DVSS.n5912 0.019716
R55959 DVSS.n6073 DVSS.n6072 0.019716
R55960 DVSS.n6072 DVSS.n5911 0.019716
R55961 DVSS.n6066 DVSS.n6065 0.019716
R55962 DVSS.n6065 DVSS.n5910 0.019716
R55963 DVSS.n6061 DVSS.n6060 0.019716
R55964 DVSS.n6060 DVSS.n5909 0.019716
R55965 DVSS.n6054 DVSS.n6053 0.019716
R55966 DVSS.n6053 DVSS.n5908 0.019716
R55967 DVSS.n6049 DVSS.n6048 0.019716
R55968 DVSS.n6048 DVSS.n5907 0.019716
R55969 DVSS.n6042 DVSS.n6041 0.019716
R55970 DVSS.n6041 DVSS.n5906 0.019716
R55971 DVSS.n6037 DVSS.n6036 0.019716
R55972 DVSS.n6036 DVSS.n5905 0.019716
R55973 DVSS.n6030 DVSS.n6029 0.019716
R55974 DVSS.n6029 DVSS.n5904 0.019716
R55975 DVSS.n6025 DVSS.n6024 0.019716
R55976 DVSS.n6024 DVSS.n5903 0.019716
R55977 DVSS.n6018 DVSS.n6017 0.019716
R55978 DVSS.n6017 DVSS.n5902 0.019716
R55979 DVSS.n6013 DVSS.n6012 0.019716
R55980 DVSS.n6012 DVSS.n5901 0.019716
R55981 DVSS.n6006 DVSS.n6005 0.019716
R55982 DVSS.n6005 DVSS.n5900 0.019716
R55983 DVSS.n6001 DVSS.n6000 0.019716
R55984 DVSS.n6000 DVSS.n5899 0.019716
R55985 DVSS.n5994 DVSS.n5993 0.019716
R55986 DVSS.n5993 DVSS.n5898 0.019716
R55987 DVSS.n5989 DVSS.n5988 0.019716
R55988 DVSS.n5988 DVSS.n5897 0.019716
R55989 DVSS.n6229 DVSS.n5939 0.019716
R55990 DVSS.n6230 DVSS.n6229 0.019716
R55991 DVSS.n6223 DVSS.n6222 0.019716
R55992 DVSS.n6223 DVSS.n5937 0.019716
R55993 DVSS.n6218 DVSS.n6217 0.019716
R55994 DVSS.n6218 DVSS.n5936 0.019716
R55995 DVSS.n6211 DVSS.n6210 0.019716
R55996 DVSS.n6211 DVSS.n5935 0.019716
R55997 DVSS.n6206 DVSS.n6205 0.019716
R55998 DVSS.n6206 DVSS.n5934 0.019716
R55999 DVSS.n6199 DVSS.n6198 0.019716
R56000 DVSS.n6199 DVSS.n5933 0.019716
R56001 DVSS.n6194 DVSS.n6193 0.019716
R56002 DVSS.n6194 DVSS.n5932 0.019716
R56003 DVSS.n6187 DVSS.n6186 0.019716
R56004 DVSS.n6187 DVSS.n5931 0.019716
R56005 DVSS.n6182 DVSS.n6181 0.019716
R56006 DVSS.n6182 DVSS.n5930 0.019716
R56007 DVSS.n6175 DVSS.n6174 0.019716
R56008 DVSS.n6175 DVSS.n5929 0.019716
R56009 DVSS.n6170 DVSS.n6169 0.019716
R56010 DVSS.n6170 DVSS.n5928 0.019716
R56011 DVSS.n6163 DVSS.n6162 0.019716
R56012 DVSS.n6163 DVSS.n5927 0.019716
R56013 DVSS.n6158 DVSS.n6157 0.019716
R56014 DVSS.n6158 DVSS.n5926 0.019716
R56015 DVSS.n6151 DVSS.n6150 0.019716
R56016 DVSS.n6151 DVSS.n5925 0.019716
R56017 DVSS.n6146 DVSS.n6145 0.019716
R56018 DVSS.n6146 DVSS.n5924 0.019716
R56019 DVSS.n6139 DVSS.n6138 0.019716
R56020 DVSS.n6139 DVSS.n5923 0.019716
R56021 DVSS.n6134 DVSS.n6133 0.019716
R56022 DVSS.n6134 DVSS.n5922 0.019716
R56023 DVSS.n6127 DVSS.n6126 0.019716
R56024 DVSS.n6127 DVSS.n5921 0.019716
R56025 DVSS.n6122 DVSS.n6121 0.019716
R56026 DVSS.n6122 DVSS.n5920 0.019716
R56027 DVSS.n6115 DVSS.n6114 0.019716
R56028 DVSS.n6115 DVSS.n5919 0.019716
R56029 DVSS.n6110 DVSS.n6109 0.019716
R56030 DVSS.n6110 DVSS.n5918 0.019716
R56031 DVSS.n6103 DVSS.n6102 0.019716
R56032 DVSS.n6103 DVSS.n5917 0.019716
R56033 DVSS.n6098 DVSS.n6097 0.019716
R56034 DVSS.n6098 DVSS.n5916 0.019716
R56035 DVSS.n6091 DVSS.n6090 0.019716
R56036 DVSS.n6091 DVSS.n5915 0.019716
R56037 DVSS.n6086 DVSS.n6085 0.019716
R56038 DVSS.n6086 DVSS.n5914 0.019716
R56039 DVSS.n6079 DVSS.n6078 0.019716
R56040 DVSS.n6079 DVSS.n5913 0.019716
R56041 DVSS.n6074 DVSS.n6073 0.019716
R56042 DVSS.n6074 DVSS.n5912 0.019716
R56043 DVSS.n6067 DVSS.n6066 0.019716
R56044 DVSS.n6067 DVSS.n5911 0.019716
R56045 DVSS.n6062 DVSS.n6061 0.019716
R56046 DVSS.n6062 DVSS.n5910 0.019716
R56047 DVSS.n6055 DVSS.n6054 0.019716
R56048 DVSS.n6055 DVSS.n5909 0.019716
R56049 DVSS.n6050 DVSS.n6049 0.019716
R56050 DVSS.n6050 DVSS.n5908 0.019716
R56051 DVSS.n6043 DVSS.n6042 0.019716
R56052 DVSS.n6043 DVSS.n5907 0.019716
R56053 DVSS.n6038 DVSS.n6037 0.019716
R56054 DVSS.n6038 DVSS.n5906 0.019716
R56055 DVSS.n6031 DVSS.n6030 0.019716
R56056 DVSS.n6031 DVSS.n5905 0.019716
R56057 DVSS.n6026 DVSS.n6025 0.019716
R56058 DVSS.n6026 DVSS.n5904 0.019716
R56059 DVSS.n6019 DVSS.n6018 0.019716
R56060 DVSS.n6019 DVSS.n5903 0.019716
R56061 DVSS.n6014 DVSS.n6013 0.019716
R56062 DVSS.n6014 DVSS.n5902 0.019716
R56063 DVSS.n6007 DVSS.n6006 0.019716
R56064 DVSS.n6007 DVSS.n5901 0.019716
R56065 DVSS.n6002 DVSS.n6001 0.019716
R56066 DVSS.n6002 DVSS.n5900 0.019716
R56067 DVSS.n5995 DVSS.n5994 0.019716
R56068 DVSS.n5995 DVSS.n5899 0.019716
R56069 DVSS.n5990 DVSS.n5989 0.019716
R56070 DVSS.n5990 DVSS.n5898 0.019716
R56071 DVSS.n5983 DVSS.n5897 0.019716
R56072 DVSS.n19215 DVSS.n13522 0.0196854
R56073 DVSS.n19160 DVSS.n13472 0.0196854
R56074 DVSS.n19902 DVSS.n13576 0.0196854
R56075 DVSS.n19147 DVSS.n13425 0.0196854
R56076 DVSS.n9192 DVSS.n9191 0.019625
R56077 DVSS.n11987 DVSS.n11986 0.019625
R56078 DVSS.n13095 DVSS.n12923 0.0195761
R56079 DVSS.n10153 DVSS.n2071 0.0195611
R56080 DVSS.n10494 DVSS.n1621 0.0195611
R56081 DVSS.n10155 DVSS.n10154 0.0195611
R56082 DVSS.n10493 DVSS.n1622 0.0195611
R56083 DVSS.n19175 DVSS.n19172 0.0194474
R56084 DVSS.n17382 DVSS.n17309 0.0194096
R56085 DVSS.n17207 DVSS.n16933 0.0194096
R56086 DVSS.n17380 DVSS.n17379 0.0194096
R56087 DVSS.n17522 DVSS.n16935 0.0194096
R56088 DVSS.n17481 DVSS.n17480 0.0194096
R56089 DVSS.n17453 DVSS.n16924 0.0194096
R56090 DVSS.n16518 DVSS 0.0193771
R56091 DVSS DVSS.n18133 0.0193771
R56092 DVSS.n18867 DVSS.n18761 0.0192079
R56093 DVSS.n16513 DVSS.n16488 0.0191864
R56094 DVSS.n18138 DVSS.n15584 0.0191864
R56095 DVSS.n9460 DVSS.n2784 0.019175
R56096 DVSS.n13330 DVSS.n11453 0.019175
R56097 DVSS.n8591 DVSS.n3753 0.0191681
R56098 DVSS.n8592 DVSS.n3752 0.0191681
R56099 DVSS.n18513 DVSS.n18500 0.019095
R56100 DVSS.n18501 DVSS.n13672 0.019095
R56101 DVSS.n21165 DVSS.n13672 0.019095
R56102 DVSS.n21167 DVSS.n13671 0.019095
R56103 DVSS.n13671 DVSS.n13664 0.019095
R56104 DVSS.n21166 DVSS.n21165 0.019095
R56105 DVSS.n21167 DVSS.n21166 0.019095
R56106 DVSS.n18502 DVSS.n18500 0.019095
R56107 DVSS.n18502 DVSS.n18501 0.019095
R56108 DVSS.n20613 DVSS.n20612 0.0188287
R56109 DVSS.n6690 DVSS.n5887 0.0187751
R56110 DVSS.n6691 DVSS.n5886 0.0187751
R56111 DVSS.n7457 DVSS.n7456 0.018725
R56112 DVSS.n19189 DVSS 0.0186516
R56113 DVSS.n18990 DVSS.n14557 0.0181087
R56114 DVSS.n18927 DVSS.n14564 0.0181087
R56115 DVSS.n20137 DVSS.n14597 0.0181087
R56116 DVSS.n20034 DVSS.n14586 0.0181087
R56117 DVSS.n20253 DVSS.n14640 0.0181087
R56118 DVSS.n20290 DVSS.n14645 0.0181087
R56119 DVSS.n20413 DVSS.n20412 0.0181087
R56120 DVSS.n20620 DVSS.n14702 0.0181087
R56121 DVSS.n18764 DVSS.n14526 0.0181087
R56122 DVSS.n18939 DVSS.n14531 0.0181087
R56123 DVSS.n20082 DVSS.n20022 0.0181087
R56124 DVSS.n20036 DVSS.n20011 0.0181087
R56125 DVSS.n20264 DVSS.n14872 0.0181087
R56126 DVSS.n20241 DVSS.n20190 0.0181087
R56127 DVSS.n20381 DVSS.n20328 0.0181087
R56128 DVSS.n20460 DVSS.n20459 0.0181087
R56129 DVSS.n14844 DVSS.n14840 0.0180085
R56130 DVSS.n14840 DVSS.n14839 0.0180085
R56131 DVSS.n14839 DVSS.n14835 0.0180085
R56132 DVSS.n14835 DVSS.n14834 0.0180085
R56133 DVSS.n14834 DVSS.n14830 0.0180085
R56134 DVSS.n14830 DVSS.n14829 0.0180085
R56135 DVSS.n14829 DVSS.n14825 0.0180085
R56136 DVSS.n14825 DVSS.n14824 0.0180085
R56137 DVSS.n14824 DVSS.n14820 0.0180085
R56138 DVSS.n14820 DVSS.n14819 0.0180085
R56139 DVSS.n14819 DVSS.n14815 0.0180085
R56140 DVSS.n14815 DVSS.n14814 0.0180085
R56141 DVSS.n14814 DVSS.n14810 0.0180085
R56142 DVSS.n14810 DVSS.n14809 0.0180085
R56143 DVSS.n14809 DVSS.n14805 0.0180085
R56144 DVSS.n14805 DVSS.n14804 0.0180085
R56145 DVSS.n14804 DVSS.n14800 0.0180085
R56146 DVSS.n14800 DVSS.n14799 0.0180085
R56147 DVSS.n14795 DVSS.n14794 0.0180085
R56148 DVSS.n14790 DVSS.n14789 0.0180085
R56149 DVSS.n14789 DVSS.n14785 0.0180085
R56150 DVSS.n14785 DVSS.n14784 0.0180085
R56151 DVSS.n14784 DVSS.n14780 0.0180085
R56152 DVSS.n14780 DVSS.n14779 0.0180085
R56153 DVSS.n14779 DVSS.n14775 0.0180085
R56154 DVSS.n14775 DVSS.n14774 0.0180085
R56155 DVSS.n14774 DVSS.n14770 0.0180085
R56156 DVSS.n14770 DVSS.n14769 0.0180085
R56157 DVSS.n14769 DVSS.n14765 0.0180085
R56158 DVSS.n14765 DVSS.n14764 0.0180085
R56159 DVSS.n14764 DVSS.n14760 0.0180085
R56160 DVSS.n14760 DVSS.n14759 0.0180085
R56161 DVSS.n14759 DVSS.n14755 0.0180085
R56162 DVSS.n14755 DVSS.n14754 0.0180085
R56163 DVSS.n14754 DVSS.n14750 0.0180085
R56164 DVSS.n14750 DVSS.n14749 0.0180085
R56165 DVSS.n14749 DVSS.n14745 0.0180085
R56166 DVSS.n14745 DVSS.n14744 0.0180085
R56167 DVSS.n14744 DVSS.n14708 0.0180085
R56168 DVSS.n20606 DVSS.n14709 0.0180085
R56169 DVSS.n20606 DVSS.n20605 0.0180085
R56170 DVSS.n20605 DVSS.n20476 0.0180085
R56171 DVSS.n20599 DVSS.n20476 0.0180085
R56172 DVSS.n20599 DVSS.n20598 0.0180085
R56173 DVSS.n20598 DVSS.n20478 0.0180085
R56174 DVSS.n20592 DVSS.n20478 0.0180085
R56175 DVSS.n20592 DVSS.n20591 0.0180085
R56176 DVSS.n20591 DVSS.n20480 0.0180085
R56177 DVSS.n20585 DVSS.n20480 0.0180085
R56178 DVSS.n20585 DVSS.n20584 0.0180085
R56179 DVSS.n20584 DVSS.n20482 0.0180085
R56180 DVSS.n20578 DVSS.n20482 0.0180085
R56181 DVSS.n20578 DVSS.n20577 0.0180085
R56182 DVSS.n20577 DVSS.n20484 0.0180085
R56183 DVSS.n20571 DVSS.n20484 0.0180085
R56184 DVSS.n20571 DVSS.n20570 0.0180085
R56185 DVSS.n20570 DVSS.n20486 0.0180085
R56186 DVSS.n20564 DVSS.n20486 0.0180085
R56187 DVSS.n20564 DVSS.n20563 0.0180085
R56188 DVSS.n20559 DVSS.n20558 0.0180085
R56189 DVSS.n20554 DVSS.n20553 0.0180085
R56190 DVSS.n20553 DVSS.n20491 0.0180085
R56191 DVSS.n20547 DVSS.n20491 0.0180085
R56192 DVSS.n20547 DVSS.n20546 0.0180085
R56193 DVSS.n20546 DVSS.n20493 0.0180085
R56194 DVSS.n20540 DVSS.n20493 0.0180085
R56195 DVSS.n20540 DVSS.n20539 0.0180085
R56196 DVSS.n20539 DVSS.n20495 0.0180085
R56197 DVSS.n20533 DVSS.n20495 0.0180085
R56198 DVSS.n20533 DVSS.n20532 0.0180085
R56199 DVSS.n20532 DVSS.n20497 0.0180085
R56200 DVSS.n20526 DVSS.n20497 0.0180085
R56201 DVSS.n20526 DVSS.n20525 0.0180085
R56202 DVSS.n20525 DVSS.n20499 0.0180085
R56203 DVSS.n20519 DVSS.n20499 0.0180085
R56204 DVSS.n20519 DVSS.n20518 0.0180085
R56205 DVSS.n20518 DVSS.n20501 0.0180085
R56206 DVSS.n20512 DVSS.n20501 0.0180085
R56207 DVSS.n20512 DVSS.n20511 0.0180085
R56208 DVSS.n18754 DVSS.n18752 0.0178311
R56209 DVSS.n18752 DVSS.n18750 0.0178311
R56210 DVSS.n18750 DVSS.n18748 0.0178311
R56211 DVSS.n18748 DVSS.n18746 0.0178311
R56212 DVSS.n18746 DVSS.n18744 0.0178311
R56213 DVSS.n18744 DVSS.n18742 0.0178311
R56214 DVSS.n18742 DVSS.n18740 0.0178311
R56215 DVSS.n18740 DVSS.n18738 0.0178311
R56216 DVSS.n18738 DVSS.n18736 0.0178311
R56217 DVSS.n18736 DVSS.n18734 0.0178311
R56218 DVSS.n18734 DVSS.n18732 0.0178311
R56219 DVSS.n18732 DVSS.n18730 0.0178311
R56220 DVSS.n18730 DVSS.n18728 0.0178311
R56221 DVSS.n18728 DVSS.n18726 0.0178311
R56222 DVSS.n18726 DVSS.n18724 0.0178311
R56223 DVSS.n18724 DVSS.n18722 0.0178311
R56224 DVSS.n18722 DVSS.n18720 0.0178311
R56225 DVSS.n18720 DVSS.n18718 0.0178311
R56226 DVSS.n18718 DVSS.n18716 0.0178311
R56227 DVSS.n18716 DVSS.n18714 0.0178311
R56228 DVSS.n18712 DVSS.n18710 0.0178311
R56229 DVSS.n18707 DVSS.n18705 0.0178311
R56230 DVSS.n18705 DVSS.n18703 0.0178311
R56231 DVSS.n18703 DVSS.n18701 0.0178311
R56232 DVSS.n18701 DVSS.n18699 0.0178311
R56233 DVSS.n18699 DVSS.n18697 0.0178311
R56234 DVSS.n18697 DVSS.n18695 0.0178311
R56235 DVSS.n18695 DVSS.n18693 0.0178311
R56236 DVSS.n18693 DVSS.n18691 0.0178311
R56237 DVSS.n18691 DVSS.n18689 0.0178311
R56238 DVSS.n18689 DVSS.n18687 0.0178311
R56239 DVSS.n18687 DVSS.n18685 0.0178311
R56240 DVSS.n18685 DVSS.n18683 0.0178311
R56241 DVSS.n18683 DVSS.n18681 0.0178311
R56242 DVSS.n18681 DVSS.n18679 0.0178311
R56243 DVSS.n18679 DVSS.n18677 0.0178311
R56244 DVSS.n18677 DVSS.n18675 0.0178311
R56245 DVSS.n18675 DVSS.n18673 0.0178311
R56246 DVSS.n18673 DVSS.n18671 0.0178311
R56247 DVSS.n18671 DVSS.n18669 0.0178311
R56248 DVSS.n18669 DVSS.n18667 0.0178311
R56249 DVSS.n18667 DVSS.n18665 0.0178311
R56250 DVSS.n18779 DVSS.n18777 0.0178311
R56251 DVSS.n18781 DVSS.n18779 0.0178311
R56252 DVSS.n18783 DVSS.n18781 0.0178311
R56253 DVSS.n18785 DVSS.n18783 0.0178311
R56254 DVSS.n18787 DVSS.n18785 0.0178311
R56255 DVSS.n18789 DVSS.n18787 0.0178311
R56256 DVSS.n18791 DVSS.n18789 0.0178311
R56257 DVSS.n18793 DVSS.n18791 0.0178311
R56258 DVSS.n18795 DVSS.n18793 0.0178311
R56259 DVSS.n18797 DVSS.n18795 0.0178311
R56260 DVSS.n18799 DVSS.n18797 0.0178311
R56261 DVSS.n18801 DVSS.n18799 0.0178311
R56262 DVSS.n18803 DVSS.n18801 0.0178311
R56263 DVSS.n18805 DVSS.n18803 0.0178311
R56264 DVSS.n18807 DVSS.n18805 0.0178311
R56265 DVSS.n18809 DVSS.n18807 0.0178311
R56266 DVSS.n18811 DVSS.n18809 0.0178311
R56267 DVSS.n18813 DVSS.n18811 0.0178311
R56268 DVSS.n18815 DVSS.n18813 0.0178311
R56269 DVSS.n18817 DVSS.n18815 0.0178311
R56270 DVSS.n18819 DVSS.n18817 0.0178311
R56271 DVSS.n18824 DVSS.n18822 0.0178311
R56272 DVSS.n18828 DVSS.n18826 0.0178311
R56273 DVSS.n18830 DVSS.n18828 0.0178311
R56274 DVSS.n18832 DVSS.n18830 0.0178311
R56275 DVSS.n18834 DVSS.n18832 0.0178311
R56276 DVSS.n18836 DVSS.n18834 0.0178311
R56277 DVSS.n18838 DVSS.n18836 0.0178311
R56278 DVSS.n18840 DVSS.n18838 0.0178311
R56279 DVSS.n18842 DVSS.n18840 0.0178311
R56280 DVSS.n18844 DVSS.n18842 0.0178311
R56281 DVSS.n18846 DVSS.n18844 0.0178311
R56282 DVSS.n18848 DVSS.n18846 0.0178311
R56283 DVSS.n18850 DVSS.n18848 0.0178311
R56284 DVSS.n18852 DVSS.n18850 0.0178311
R56285 DVSS.n18854 DVSS.n18852 0.0178311
R56286 DVSS.n18856 DVSS.n18854 0.0178311
R56287 DVSS.n18858 DVSS.n18856 0.0178311
R56288 DVSS.n18860 DVSS.n18858 0.0178311
R56289 DVSS.n18862 DVSS.n18860 0.0178311
R56290 DVSS.n18864 DVSS.n18862 0.0178311
R56291 DVSS.n18866 DVSS.n18864 0.0178311
R56292 DVSS.n22074 DVSS.n21603 0.0177537
R56293 DVSS.n22046 DVSS.n21706 0.0177537
R56294 DVSS.n21850 DVSS.n21849 0.0177537
R56295 DVSS.n21963 DVSS.n21799 0.0177537
R56296 DVSS.n7089 DVSS.n4883 0.0175961
R56297 DVSS.n7091 DVSS.n7090 0.0175961
R56298 DVSS.n17778 DVSS.n15937 0.0175526
R56299 DVSS.n18118 DVSS.n15515 0.0175526
R56300 DVSS.n6664 DVSS.n6253 0.017282
R56301 DVSS.n6667 DVSS.n6666 0.017282
R56302 DVSS.n6667 DVSS.n5894 0.017282
R56303 DVSS.n6683 DVSS.n5894 0.017282
R56304 DVSS.n6685 DVSS.n5873 0.017282
R56305 DVSS.n7037 DVSS.n5873 0.017282
R56306 DVSS.n7041 DVSS.n7039 0.017282
R56307 DVSS.n7041 DVSS.n7040 0.017282
R56308 DVSS.n7064 DVSS.n7063 0.017282
R56309 DVSS.n7065 DVSS.n7064 0.017282
R56310 DVSS.n7083 DVSS.n7082 0.017282
R56311 DVSS.n7084 DVSS.n7083 0.017282
R56312 DVSS.n7084 DVSS.n4837 0.017282
R56313 DVSS.n7108 DVSS.n4837 0.017282
R56314 DVSS.n7109 DVSS.n7108 0.017282
R56315 DVSS.n7446 DVSS.n4822 0.017282
R56316 DVSS.n7801 DVSS.n4822 0.017282
R56317 DVSS.n7803 DVSS.n4808 0.017282
R56318 DVSS.n7821 DVSS.n4808 0.017282
R56319 DVSS.n7823 DVSS.n4366 0.017282
R56320 DVSS.n8094 DVSS.n4366 0.017282
R56321 DVSS.n8097 DVSS.n8096 0.017282
R56322 DVSS.n8097 DVSS.n4018 0.017282
R56323 DVSS.n8115 DVSS.n4018 0.017282
R56324 DVSS.n8118 DVSS.n8117 0.017282
R56325 DVSS.n8117 DVSS.n4008 0.017282
R56326 DVSS.n8128 DVSS.n4011 0.017282
R56327 DVSS.n8336 DVSS.n3410 0.017282
R56328 DVSS.n8608 DVSS.n3410 0.017282
R56329 DVSS.n8611 DVSS.n8610 0.017282
R56330 DVSS.n8611 DVSS.n3063 0.017282
R56331 DVSS.n8628 DVSS.n3063 0.017282
R56332 DVSS.n8630 DVSS.n3049 0.017282
R56333 DVSS.n8982 DVSS.n3049 0.017282
R56334 DVSS.n8985 DVSS.n8984 0.017282
R56335 DVSS.n8984 DVSS.n3040 0.017282
R56336 DVSS.n8995 DVSS.n3042 0.017282
R56337 DVSS.n3042 DVSS.n3041 0.017282
R56338 DVSS.n9203 DVSS.n2734 0.017282
R56339 DVSS.n9763 DVSS.n2734 0.017282
R56340 DVSS.n9767 DVSS.n9765 0.017282
R56341 DVSS.n10119 DVSS.n2713 0.017282
R56342 DVSS.n10123 DVSS.n10121 0.017282
R56343 DVSS.n10123 DVSS.n10122 0.017282
R56344 DVSS.n10147 DVSS.n10146 0.017282
R56345 DVSS.n10148 DVSS.n10147 0.017282
R56346 DVSS.n10171 DVSS.n10170 0.017282
R56347 DVSS.n10457 DVSS.n10171 0.017282
R56348 DVSS.n10481 DVSS.n1964 0.017282
R56349 DVSS.n10482 DVSS.n10481 0.017282
R56350 DVSS.n10483 DVSS.n10482 0.017282
R56351 DVSS.n10502 DVSS.n10501 0.017282
R56352 DVSS.n10503 DVSS.n10502 0.017282
R56353 DVSS.n13362 DVSS.n1506 0.017282
R56354 DVSS.n13346 DVSS.n13345 0.017282
R56355 DVSS.n13345 DVSS.n13344 0.017282
R56356 DVSS.n11613 DVSS.n11612 0.017282
R56357 DVSS.n11612 DVSS.n11609 0.017282
R56358 DVSS.n13134 DVSS.n11610 0.017282
R56359 DVSS.n13128 DVSS.n11610 0.017282
R56360 DVSS.n13128 DVSS.n13127 0.017282
R56361 DVSS.n13125 DVSS.n11625 0.017282
R56362 DVSS.n12341 DVSS.n11625 0.017282
R56363 DVSS.n13107 DVSS.n12343 0.017282
R56364 DVSS.n13107 DVSS.n13106 0.017282
R56365 DVSS.n13106 DVSS.n13105 0.017282
R56366 DVSS.n13105 DVSS.n12346 0.017282
R56367 DVSS.n13103 DVSS.n12346 0.017282
R56368 DVSS.n21144 DVSS.n21143 0.0172684
R56369 DVSS.n20977 DVSS.n14276 0.0172684
R56370 DVSS.n21460 DVSS.n21451 0.0172442
R56371 DVSS.n22590 DVSS.n22589 0.0172442
R56372 DVSS.n22932 DVSS.n22931 0.0172442
R56373 DVSS.n22959 DVSS.n22958 0.0172442
R56374 DVSS.n9189 DVSS.n2889 0.0172031
R56375 DVSS.n11645 DVSS.n11632 0.0172031
R56376 DVSS.n9190 DVSS.n2887 0.0172031
R56377 DVSS.n11639 DVSS.n11634 0.0172031
R56378 DVSS.n18162 DVSS.n18161 0.0171667
R56379 DVSS.n18161 DVSS.n18160 0.0171667
R56380 DVSS.n21444 DVSS.n21443 0.0171667
R56381 DVSS.n21443 DVSS.n21442 0.0171667
R56382 DVSS.n19501 DVSS.n19279 0.0171304
R56383 DVSS.n22456 DVSS.n22455 0.0171304
R56384 DVSS.n19845 DVSS.n19110 0.0171304
R56385 DVSS.n22334 DVSS.n22333 0.0171304
R56386 DVSS.n20613 DVSS.n14708 0.017087
R56387 DVSS.n8325 DVSS.n8324 0.016925
R56388 DVSS.n18867 DVSS.n18866 0.0169189
R56389 DVSS.n9458 DVSS.n2786 0.01681
R56390 DVSS.n13328 DVSS.n11456 0.01681
R56391 DVSS.n9459 DVSS.n2785 0.01681
R56392 DVSS.n13329 DVSS.n11454 0.01681
R56393 DVSS.n8630 DVSS.n8629 0.0167406
R56394 DVSS.n13135 DVSS.n11609 0.0167406
R56395 DVSS.n16549 DVSS.n16542 0.0165729
R56396 DVSS.n16547 DVSS.n16477 0.0165729
R56397 DVSS.n16483 DVSS.n16477 0.0165729
R56398 DVSS.n16546 DVSS.n16476 0.0165729
R56399 DVSS.n16482 DVSS.n16476 0.0165729
R56400 DVSS.n16545 DVSS.n16475 0.0165729
R56401 DVSS.n16481 DVSS.n16475 0.0165729
R56402 DVSS.n16544 DVSS.n16474 0.0165729
R56403 DVSS.n16480 DVSS.n16474 0.0165729
R56404 DVSS.n16543 DVSS.n16473 0.0165729
R56405 DVSS.n16479 DVSS.n16473 0.0165729
R56406 DVSS.n16471 DVSS.n16359 0.0165729
R56407 DVSS.n16469 DVSS.n16372 0.0165729
R56408 DVSS.n16469 DVSS.n16468 0.0165729
R56409 DVSS.n16371 DVSS.n16370 0.0165729
R56410 DVSS.n16375 DVSS.n16371 0.0165729
R56411 DVSS.n16369 DVSS.n16368 0.0165729
R56412 DVSS.n16374 DVSS.n16369 0.0165729
R56413 DVSS.n16367 DVSS.n16366 0.0165729
R56414 DVSS.n16373 DVSS.n16367 0.0165729
R56415 DVSS.n18087 DVSS.n18086 0.0165729
R56416 DVSS.n15643 DVSS.n15642 0.0165729
R56417 DVSS.n15649 DVSS.n15643 0.0165729
R56418 DVSS.n15641 DVSS.n15640 0.0165729
R56419 DVSS.n15648 DVSS.n15641 0.0165729
R56420 DVSS.n15639 DVSS.n15638 0.0165729
R56421 DVSS.n15647 DVSS.n15639 0.0165729
R56422 DVSS.n15637 DVSS.n15636 0.0165729
R56423 DVSS.n15637 DVSS.n15628 0.0165729
R56424 DVSS.n18113 DVSS.n18090 0.0165729
R56425 DVSS.n18095 DVSS.n15627 0.0165729
R56426 DVSS.n18106 DVSS.n15627 0.0165729
R56427 DVSS.n18094 DVSS.n15626 0.0165729
R56428 DVSS.n18105 DVSS.n15626 0.0165729
R56429 DVSS.n18093 DVSS.n15625 0.0165729
R56430 DVSS.n18104 DVSS.n15625 0.0165729
R56431 DVSS.n18092 DVSS.n15624 0.0165729
R56432 DVSS.n18103 DVSS.n15624 0.0165729
R56433 DVSS.n18091 DVSS.n15623 0.0165729
R56434 DVSS.n18102 DVSS.n15623 0.0165729
R56435 DVSS.n16221 DVSS.n16186 0.0165729
R56436 DVSS.n16219 DVSS.n16186 0.0165729
R56437 DVSS.n16209 DVSS.n16187 0.0165729
R56438 DVSS.n16218 DVSS.n16187 0.0165729
R56439 DVSS.n16207 DVSS.n16188 0.0165729
R56440 DVSS.n16217 DVSS.n16188 0.0165729
R56441 DVSS.n16205 DVSS.n16189 0.0165729
R56442 DVSS.n16216 DVSS.n16189 0.0165729
R56443 DVSS.n16203 DVSS.n16190 0.0165729
R56444 DVSS.n16215 DVSS.n16190 0.0165729
R56445 DVSS.n16201 DVSS.n16191 0.0165729
R56446 DVSS.n16214 DVSS.n16191 0.0165729
R56447 DVSS.n16213 DVSS.n16192 0.0165729
R56448 DVSS.n16198 DVSS.n16193 0.0165729
R56449 DVSS.n16212 DVSS.n16193 0.0165729
R56450 DVSS.n16196 DVSS.n16194 0.0165729
R56451 DVSS.n16211 DVSS.n16194 0.0165729
R56452 DVSS.n16461 DVSS.n16460 0.0165729
R56453 DVSS.n16460 DVSS.n16459 0.0165729
R56454 DVSS.n16457 DVSS.n16456 0.0165729
R56455 DVSS.n16456 DVSS.n16455 0.0165729
R56456 DVSS.n16453 DVSS.n16452 0.0165729
R56457 DVSS.n16450 DVSS.n16449 0.0165729
R56458 DVSS.n16449 DVSS.n16448 0.0165729
R56459 DVSS.n16446 DVSS.n16445 0.0165729
R56460 DVSS.n16445 DVSS.n16444 0.0165729
R56461 DVSS.n16442 DVSS.n16441 0.0165729
R56462 DVSS.n16441 DVSS.n16440 0.0165729
R56463 DVSS.n16438 DVSS.n16437 0.0165729
R56464 DVSS.n16437 DVSS.n16436 0.0165729
R56465 DVSS.n16434 DVSS.n16433 0.0165729
R56466 DVSS.n16433 DVSS.n16432 0.0165729
R56467 DVSS.n16430 DVSS.n16429 0.0165729
R56468 DVSS.n16429 DVSS.n16428 0.0165729
R56469 DVSS.n16462 DVSS.n16461 0.0165729
R56470 DVSS.n16458 DVSS.n16457 0.0165729
R56471 DVSS.n16454 DVSS.n16453 0.0165729
R56472 DVSS.n16451 DVSS.n16450 0.0165729
R56473 DVSS.n16447 DVSS.n16446 0.0165729
R56474 DVSS.n16443 DVSS.n16442 0.0165729
R56475 DVSS.n16439 DVSS.n16438 0.0165729
R56476 DVSS.n16435 DVSS.n16434 0.0165729
R56477 DVSS.n16431 DVSS.n16430 0.0165729
R56478 DVSS.n16459 DVSS.n16458 0.0165729
R56479 DVSS.n16455 DVSS.n16454 0.0165729
R56480 DVSS.n16448 DVSS.n16447 0.0165729
R56481 DVSS.n16444 DVSS.n16443 0.0165729
R56482 DVSS.n16440 DVSS.n16439 0.0165729
R56483 DVSS.n16436 DVSS.n16435 0.0165729
R56484 DVSS.n16432 DVSS.n16431 0.0165729
R56485 DVSS.n16428 DVSS.n16427 0.0165729
R56486 DVSS.n16222 DVSS.n16221 0.0165729
R56487 DVSS.n16210 DVSS.n16209 0.0165729
R56488 DVSS.n16208 DVSS.n16207 0.0165729
R56489 DVSS.n16206 DVSS.n16205 0.0165729
R56490 DVSS.n16204 DVSS.n16203 0.0165729
R56491 DVSS.n16202 DVSS.n16201 0.0165729
R56492 DVSS.n16199 DVSS.n16198 0.0165729
R56493 DVSS.n16197 DVSS.n16196 0.0165729
R56494 DVSS.n16219 DVSS.n16210 0.0165729
R56495 DVSS.n16218 DVSS.n16208 0.0165729
R56496 DVSS.n16217 DVSS.n16206 0.0165729
R56497 DVSS.n16216 DVSS.n16204 0.0165729
R56498 DVSS.n16215 DVSS.n16202 0.0165729
R56499 DVSS.n16214 DVSS.n16200 0.0165729
R56500 DVSS.n16213 DVSS.n16199 0.0165729
R56501 DVSS.n16212 DVSS.n16197 0.0165729
R56502 DVSS.n16211 DVSS.n16195 0.0165729
R56503 DVSS.n16372 DVSS.n16361 0.0165729
R56504 DVSS.n16370 DVSS.n16362 0.0165729
R56505 DVSS.n16368 DVSS.n16363 0.0165729
R56506 DVSS.n16366 DVSS.n16364 0.0165729
R56507 DVSS.n16361 DVSS.n16359 0.0165729
R56508 DVSS.n16468 DVSS.n16362 0.0165729
R56509 DVSS.n16375 DVSS.n16363 0.0165729
R56510 DVSS.n16374 DVSS.n16364 0.0165729
R56511 DVSS.n16373 DVSS.n16365 0.0165729
R56512 DVSS.n16547 DVSS.n16354 0.0165729
R56513 DVSS.n16546 DVSS.n16355 0.0165729
R56514 DVSS.n16545 DVSS.n16356 0.0165729
R56515 DVSS.n16544 DVSS.n16357 0.0165729
R56516 DVSS.n16543 DVSS.n16358 0.0165729
R56517 DVSS.n16542 DVSS.n16354 0.0165729
R56518 DVSS.n16483 DVSS.n16355 0.0165729
R56519 DVSS.n16482 DVSS.n16356 0.0165729
R56520 DVSS.n16481 DVSS.n16357 0.0165729
R56521 DVSS.n16480 DVSS.n16358 0.0165729
R56522 DVSS.n16479 DVSS.n16472 0.0165729
R56523 DVSS.n15642 DVSS.n15631 0.0165729
R56524 DVSS.n15640 DVSS.n15632 0.0165729
R56525 DVSS.n15638 DVSS.n15633 0.0165729
R56526 DVSS.n15636 DVSS.n15634 0.0165729
R56527 DVSS.n18086 DVSS.n15631 0.0165729
R56528 DVSS.n15649 DVSS.n15632 0.0165729
R56529 DVSS.n15648 DVSS.n15633 0.0165729
R56530 DVSS.n15647 DVSS.n15634 0.0165729
R56531 DVSS.n18089 DVSS.n15628 0.0165729
R56532 DVSS.n18095 DVSS.n15617 0.0165729
R56533 DVSS.n18094 DVSS.n15618 0.0165729
R56534 DVSS.n18093 DVSS.n15619 0.0165729
R56535 DVSS.n18092 DVSS.n15620 0.0165729
R56536 DVSS.n18091 DVSS.n15621 0.0165729
R56537 DVSS.n18090 DVSS.n15617 0.0165729
R56538 DVSS.n18106 DVSS.n15618 0.0165729
R56539 DVSS.n18105 DVSS.n15619 0.0165729
R56540 DVSS.n18104 DVSS.n15620 0.0165729
R56541 DVSS.n18103 DVSS.n15621 0.0165729
R56542 DVSS.n18102 DVSS.n15622 0.0165729
R56543 DVSS.n10468 DVSS.n2016 0.016475
R56544 DVSS.n10468 DVSS.n10467 0.016475
R56545 DVSS.n6453 DVSS.n6253 0.0164699
R56546 DVSS.n7459 DVSS.n4826 0.016417
R56547 DVSS.n7458 DVSS.n4827 0.016417
R56548 DVSS.n20563 DVSS 0.0163191
R56549 DVSS.n17641 DVSS.n16096 0.0163049
R56550 DVSS.n16826 DVSS.n16825 0.0163049
R56551 DVSS.n16299 DVSS.n16004 0.0163049
R56552 DVSS.n16899 DVSS.n15677 0.0163049
R56553 DVSS.n6252 DVSS.n6251 0.0161992
R56554 DVSS.n9764 DVSS.n9763 0.0161992
R56555 DVSS.n10501 DVSS.n1616 0.0161992
R56556 DVSS.n18714 DVSS 0.0161588
R56557 DVSS.n8326 DVSS.n8325 0.016025
R56558 DVSS.n19193 DVSS.n19192 0.0158947
R56559 DVSS.n1151 DVSS.n217 0.015778
R56560 DVSS.n13047 DVSS.n137 0.015778
R56561 DVSS.n1096 DVSS.n813 0.015778
R56562 DVSS.n364 DVSS.n72 0.015778
R56563 DVSS.n13369 DVSS.n734 0.015774
R56564 DVSS.n21441 DVSS.n21440 0.015774
R56565 DVSS.n6685 DVSS.n6684 0.0156579
R56566 DVSS.n8095 DVSS.n8094 0.0156579
R56567 DVSS.n18514 DVSS.n18499 0.0155703
R56568 DVSS.n6669 DVSS.n5896 0.0154799
R56569 DVSS.n6681 DVSS.n5896 0.0154799
R56570 DVSS.n6687 DVSS.n5876 0.0154799
R56571 DVSS.n7035 DVSS.n5876 0.0154799
R56572 DVSS.n7043 DVSS.n5868 0.0154799
R56573 DVSS.n7043 DVSS.n5869 0.0154799
R56574 DVSS.n7061 DVSS.n5526 0.0154799
R56575 DVSS.n7067 DVSS.n5526 0.0154799
R56576 DVSS.n7080 DVSS.n5177 0.0154799
R56577 DVSS.n7086 DVSS.n5177 0.0154799
R56578 DVSS.n7086 DVSS.n4839 0.0154799
R56579 DVSS.n7106 DVSS.n4839 0.0154799
R56580 DVSS.n7106 DVSS.n4833 0.0154799
R56581 DVSS.n7450 DVSS.n4833 0.0154799
R56582 DVSS.n7798 DVSS.n4824 0.0154799
R56583 DVSS.n7799 DVSS.n7798 0.0154799
R56584 DVSS.n7805 DVSS.n4810 0.0154799
R56585 DVSS.n7819 DVSS.n4810 0.0154799
R56586 DVSS.n7825 DVSS.n4369 0.0154799
R56587 DVSS.n8092 DVSS.n4369 0.0154799
R56588 DVSS.n8099 DVSS.n4363 0.0154799
R56589 DVSS.n8099 DVSS.n4020 0.0154799
R56590 DVSS.n8113 DVSS.n4020 0.0154799
R56591 DVSS.n8121 DVSS.n8120 0.0154799
R56592 DVSS.n8122 DVSS.n8121 0.0154799
R56593 DVSS.n8126 DVSS.n3845 0.0154799
R56594 DVSS.n8333 DVSS.n3845 0.0154799
R56595 DVSS.n8335 DVSS.n3413 0.0154799
R56596 DVSS.n8606 DVSS.n3413 0.0154799
R56597 DVSS.n8613 DVSS.n3407 0.0154799
R56598 DVSS.n8613 DVSS.n3065 0.0154799
R56599 DVSS.n8626 DVSS.n3065 0.0154799
R56600 DVSS.n8632 DVSS.n3051 0.0154799
R56601 DVSS.n8980 DVSS.n3051 0.0154799
R56602 DVSS.n8988 DVSS.n8987 0.0154799
R56603 DVSS.n8989 DVSS.n8988 0.0154799
R56604 DVSS.n8993 DVSS.n2877 0.0154799
R56605 DVSS.n9200 DVSS.n2877 0.0154799
R56606 DVSS.n9202 DVSS.n2737 0.0154799
R56607 DVSS.n9761 DVSS.n2737 0.0154799
R56608 DVSS.n9769 DVSS.n2731 0.0154799
R56609 DVSS.n9769 DVSS.n2716 0.0154799
R56610 DVSS.n10117 DVSS.n2716 0.0154799
R56611 DVSS.n10125 DVSS.n2707 0.0154799
R56612 DVSS.n10125 DVSS.n2709 0.0154799
R56613 DVSS.n10144 DVSS.n2365 0.0154799
R56614 DVSS.n10150 DVSS.n2365 0.0154799
R56615 DVSS.n10168 DVSS.n2020 0.0154799
R56616 DVSS.n10459 DVSS.n2020 0.0154799
R56617 DVSS.n10479 DVSS.n1966 0.0154799
R56618 DVSS.n10479 DVSS.n1962 0.0154799
R56619 DVSS.n10485 DVSS.n1962 0.0154799
R56620 DVSS.n10499 DVSS.n1619 0.0154799
R56621 DVSS.n1619 DVSS.n1615 0.0154799
R56622 DVSS.n13360 DVSS.n1509 0.0154799
R56623 DVSS.n13360 DVSS.n1510 0.0154799
R56624 DVSS.n13348 DVSS.n10768 0.0154799
R56625 DVSS.n13342 DVSS.n10768 0.0154799
R56626 DVSS.n11616 DVSS.n11615 0.0154799
R56627 DVSS.n11617 DVSS.n11616 0.0154799
R56628 DVSS.n13132 DVSS.n13131 0.0154799
R56629 DVSS.n13131 DVSS.n13130 0.0154799
R56630 DVSS.n13130 DVSS.n11621 0.0154799
R56631 DVSS.n13123 DVSS.n11629 0.0154799
R56632 DVSS.n12339 DVSS.n11629 0.0154799
R56633 DVSS.n13109 DVSS.n11996 0.0154799
R56634 DVSS.n13109 DVSS.n11997 0.0154799
R56635 DVSS.n6668 DVSS.n5895 0.0154799
R56636 DVSS.n6682 DVSS.n5895 0.0154799
R56637 DVSS.n6686 DVSS.n5874 0.0154799
R56638 DVSS.n7036 DVSS.n5874 0.0154799
R56639 DVSS.n7042 DVSS.n5870 0.0154799
R56640 DVSS.n7042 DVSS.n5871 0.0154799
R56641 DVSS.n7062 DVSS.n5527 0.0154799
R56642 DVSS.n7066 DVSS.n5527 0.0154799
R56643 DVSS.n7081 DVSS.n5178 0.0154799
R56644 DVSS.n7085 DVSS.n5178 0.0154799
R56645 DVSS.n7085 DVSS.n4838 0.0154799
R56646 DVSS.n7107 DVSS.n4838 0.0154799
R56647 DVSS.n7107 DVSS.n4835 0.0154799
R56648 DVSS.n7449 DVSS.n4835 0.0154799
R56649 DVSS.n7445 DVSS.n4823 0.0154799
R56650 DVSS.n7800 DVSS.n4823 0.0154799
R56651 DVSS.n7804 DVSS.n4809 0.0154799
R56652 DVSS.n7820 DVSS.n4809 0.0154799
R56653 DVSS.n7824 DVSS.n4367 0.0154799
R56654 DVSS.n8093 DVSS.n4367 0.0154799
R56655 DVSS.n8098 DVSS.n4364 0.0154799
R56656 DVSS.n8098 DVSS.n4019 0.0154799
R56657 DVSS.n8114 DVSS.n4019 0.0154799
R56658 DVSS.n8119 DVSS.n4012 0.0154799
R56659 DVSS.n8123 DVSS.n4012 0.0154799
R56660 DVSS.n8127 DVSS.n8125 0.0154799
R56661 DVSS.n8125 DVSS.n3844 0.0154799
R56662 DVSS.n8337 DVSS.n3411 0.0154799
R56663 DVSS.n8607 DVSS.n3411 0.0154799
R56664 DVSS.n8612 DVSS.n3408 0.0154799
R56665 DVSS.n8612 DVSS.n3064 0.0154799
R56666 DVSS.n8627 DVSS.n3064 0.0154799
R56667 DVSS.n8631 DVSS.n3050 0.0154799
R56668 DVSS.n8981 DVSS.n3050 0.0154799
R56669 DVSS.n8986 DVSS.n3043 0.0154799
R56670 DVSS.n8990 DVSS.n3043 0.0154799
R56671 DVSS.n8994 DVSS.n8992 0.0154799
R56672 DVSS.n8992 DVSS.n2876 0.0154799
R56673 DVSS.n9204 DVSS.n2735 0.0154799
R56674 DVSS.n9762 DVSS.n2735 0.0154799
R56675 DVSS.n9768 DVSS.n2732 0.0154799
R56676 DVSS.n9768 DVSS.n2714 0.0154799
R56677 DVSS.n10118 DVSS.n2714 0.0154799
R56678 DVSS.n10124 DVSS.n2710 0.0154799
R56679 DVSS.n10124 DVSS.n2711 0.0154799
R56680 DVSS.n10145 DVSS.n2366 0.0154799
R56681 DVSS.n10149 DVSS.n2366 0.0154799
R56682 DVSS.n10169 DVSS.n2022 0.0154799
R56683 DVSS.n10458 DVSS.n2022 0.0154799
R56684 DVSS.n10480 DVSS.n1965 0.0154799
R56685 DVSS.n10480 DVSS.n1963 0.0154799
R56686 DVSS.n10484 DVSS.n1963 0.0154799
R56687 DVSS.n10500 DVSS.n1613 0.0154799
R56688 DVSS.n10504 DVSS.n1613 0.0154799
R56689 DVSS.n13361 DVSS.n1507 0.0154799
R56690 DVSS.n13361 DVSS.n1508 0.0154799
R56691 DVSS.n13347 DVSS.n10770 0.0154799
R56692 DVSS.n13343 DVSS.n10770 0.0154799
R56693 DVSS.n11614 DVSS.n11611 0.0154799
R56694 DVSS.n11618 DVSS.n11611 0.0154799
R56695 DVSS.n13133 DVSS.n11620 0.0154799
R56696 DVSS.n13129 DVSS.n11620 0.0154799
R56697 DVSS.n13129 DVSS.n11623 0.0154799
R56698 DVSS.n13124 DVSS.n11627 0.0154799
R56699 DVSS.n12340 DVSS.n11627 0.0154799
R56700 DVSS.n13108 DVSS.n11998 0.0154799
R56701 DVSS.n13108 DVSS.n11999 0.0154799
R56702 DVSS.n18648 DVSS.n14556 0.0151739
R56703 DVSS.n18963 DVSS.n14553 0.0151739
R56704 DVSS.n20135 DVSS.n14590 0.0151739
R56705 DVSS.n20164 DVSS.n14601 0.0151739
R56706 DVSS.n20268 DVSS.n14641 0.0151739
R56707 DVSS.n20294 DVSS.n14636 0.0151739
R56708 DVSS.n20415 DVSS.n20414 0.0151739
R56709 DVSS.n20451 DVSS.n20449 0.0151739
R56710 DVSS.n18891 DVSS.n14525 0.0151739
R56711 DVSS.n18941 DVSS.n14520 0.0151739
R56712 DVSS.n20088 DVSS.n20015 0.0151739
R56713 DVSS.n20172 DVSS.n20026 0.0151739
R56714 DVSS.n20266 DVSS.n20186 0.0151739
R56715 DVSS.n20235 DVSS.n14868 0.0151739
R56716 DVSS.n20379 DVSS.n14859 0.0151739
R56717 DVSS.n20333 DVSS.n14852 0.0151739
R56718 DVSS.n8118 DVSS.n8116 0.0151165
R56719 DVSS.n8632 DVSS.n3060 0.0149966
R56720 DVSS.n11617 DVSS.n11502 0.0149966
R56721 DVSS.n8631 DVSS.n3061 0.0149966
R56722 DVSS.n11619 DVSS.n11618 0.0149966
R56723 DVSS.n18869 DVSS.n18868 0.0149101
R56724 DVSS.n18986 DVSS.n18869 0.0149101
R56725 DVSS.n18907 DVSS.n18884 0.0149101
R56726 DVSS.n18917 DVSS.n14576 0.0149101
R56727 DVSS.n20682 DVSS.n14576 0.0149101
R56728 DVSS.n20682 DVSS.n20681 0.0149101
R56729 DVSS.n20681 DVSS.n20680 0.0149101
R56730 DVSS.n20131 DVSS.n20052 0.0149101
R56731 DVSS.n20078 DVSS.n20052 0.0149101
R56732 DVSS.n20667 DVSS.n14611 0.0149101
R56733 DVSS.n20667 DVSS.n20666 0.0149101
R56734 DVSS.n20666 DVSS.n20665 0.0149101
R56735 DVSS.n20655 DVSS.n14624 0.0149101
R56736 DVSS.n20655 DVSS.n20654 0.0149101
R56737 DVSS.n20654 DVSS.n20653 0.0149101
R56738 DVSS.n20298 DVSS.n20225 0.0149101
R56739 DVSS.n20298 DVSS.n20226 0.0149101
R56740 DVSS.n20639 DVSS.n20638 0.0149101
R56741 DVSS.n20638 DVSS.n14663 0.0149101
R56742 DVSS.n20627 DVSS.n14663 0.0149101
R56743 DVSS.n20627 DVSS.n14676 0.0149101
R56744 DVSS.n20441 DVSS.n20440 0.0149101
R56745 DVSS.n20624 DVSS.n14694 0.0149101
R56746 DVSS.n20614 DVSS.n14694 0.0149101
R56747 DVSS.n8322 DVSS.n3857 0.014845
R56748 DVSS.n8323 DVSS.n3855 0.014845
R56749 DVSS.n12751 DVSS.n11997 0.014755
R56750 DVSS.n12348 DVSS.n11999 0.014755
R56751 DVSS.n20613 DVSS.n14709 0.0146297
R56752 DVSS.n10121 DVSS.n10120 0.0145752
R56753 DVSS.n10457 DVSS.n10456 0.0145752
R56754 DVSS.n9761 DVSS.n2738 0.0145134
R56755 DVSS.n10499 DVSS.n1618 0.0145134
R56756 DVSS.n9762 DVSS.n2736 0.0145134
R56757 DVSS.n10500 DVSS.n1617 0.0145134
R56758 DVSS.n18867 DVSS.n18754 0.0144865
R56759 DVSS.n21159 DVSS.n13675 0.0144535
R56760 DVSS.n20989 DVSS.n20988 0.0144535
R56761 DVSS.n10462 DVSS.n2010 0.014452
R56762 DVSS.n10465 DVSS.n2010 0.014452
R56763 DVSS.n10464 DVSS.n10463 0.014452
R56764 DVSS.n10466 DVSS.n10464 0.014452
R56765 DVSS.n12772 DVSS.n12771 0.01445
R56766 DVSS.n12771 DVSS.n12355 0.01445
R56767 DVSS.n12602 DVSS.n12355 0.01445
R56768 DVSS.n12602 DVSS.n12601 0.01445
R56769 DVSS.n12606 DVSS.n12601 0.01445
R56770 DVSS.n12607 DVSS.n12606 0.01445
R56771 DVSS.n12608 DVSS.n12607 0.01445
R56772 DVSS.n12608 DVSS.n12599 0.01445
R56773 DVSS.n12612 DVSS.n12599 0.01445
R56774 DVSS.n12613 DVSS.n12612 0.01445
R56775 DVSS.n12614 DVSS.n12613 0.01445
R56776 DVSS.n12614 DVSS.n12597 0.01445
R56777 DVSS.n12618 DVSS.n12597 0.01445
R56778 DVSS.n12619 DVSS.n12618 0.01445
R56779 DVSS.n12620 DVSS.n12619 0.01445
R56780 DVSS.n12620 DVSS.n12595 0.01445
R56781 DVSS.n12624 DVSS.n12595 0.01445
R56782 DVSS.n12625 DVSS.n12624 0.01445
R56783 DVSS.n12626 DVSS.n12625 0.01445
R56784 DVSS.n12626 DVSS.n12593 0.01445
R56785 DVSS.n12630 DVSS.n12593 0.01445
R56786 DVSS.n12631 DVSS.n12630 0.01445
R56787 DVSS.n12632 DVSS.n12631 0.01445
R56788 DVSS.n12632 DVSS.n12591 0.01445
R56789 DVSS.n12636 DVSS.n12591 0.01445
R56790 DVSS.n12637 DVSS.n12636 0.01445
R56791 DVSS.n12638 DVSS.n12637 0.01445
R56792 DVSS.n12638 DVSS.n12589 0.01445
R56793 DVSS.n12642 DVSS.n12589 0.01445
R56794 DVSS.n12643 DVSS.n12642 0.01445
R56795 DVSS.n12644 DVSS.n12643 0.01445
R56796 DVSS.n12644 DVSS.n12587 0.01445
R56797 DVSS.n12648 DVSS.n12587 0.01445
R56798 DVSS.n12649 DVSS.n12648 0.01445
R56799 DVSS.n12650 DVSS.n12649 0.01445
R56800 DVSS.n12650 DVSS.n12585 0.01445
R56801 DVSS.n12654 DVSS.n12585 0.01445
R56802 DVSS.n12655 DVSS.n12654 0.01445
R56803 DVSS.n12656 DVSS.n12655 0.01445
R56804 DVSS.n12656 DVSS.n12583 0.01445
R56805 DVSS.n12660 DVSS.n12583 0.01445
R56806 DVSS.n12661 DVSS.n12660 0.01445
R56807 DVSS.n12662 DVSS.n12661 0.01445
R56808 DVSS.n12662 DVSS.n12581 0.01445
R56809 DVSS.n12666 DVSS.n12581 0.01445
R56810 DVSS.n12667 DVSS.n12666 0.01445
R56811 DVSS.n12668 DVSS.n12667 0.01445
R56812 DVSS.n12668 DVSS.n12579 0.01445
R56813 DVSS.n12672 DVSS.n12579 0.01445
R56814 DVSS.n12673 DVSS.n12672 0.01445
R56815 DVSS.n12674 DVSS.n12673 0.01445
R56816 DVSS.n12674 DVSS.n12577 0.01445
R56817 DVSS.n12678 DVSS.n12577 0.01445
R56818 DVSS.n12679 DVSS.n12678 0.01445
R56819 DVSS.n12680 DVSS.n12679 0.01445
R56820 DVSS.n12680 DVSS.n12575 0.01445
R56821 DVSS.n12684 DVSS.n12575 0.01445
R56822 DVSS.n12685 DVSS.n12684 0.01445
R56823 DVSS.n12686 DVSS.n12685 0.01445
R56824 DVSS.n12686 DVSS.n12573 0.01445
R56825 DVSS.n12690 DVSS.n12573 0.01445
R56826 DVSS.n12691 DVSS.n12690 0.01445
R56827 DVSS.n12692 DVSS.n12691 0.01445
R56828 DVSS.n12692 DVSS.n12571 0.01445
R56829 DVSS.n12696 DVSS.n12571 0.01445
R56830 DVSS.n12697 DVSS.n12696 0.01445
R56831 DVSS.n12698 DVSS.n12697 0.01445
R56832 DVSS.n12698 DVSS.n12569 0.01445
R56833 DVSS.n12702 DVSS.n12569 0.01445
R56834 DVSS.n12703 DVSS.n12702 0.01445
R56835 DVSS.n12704 DVSS.n12703 0.01445
R56836 DVSS.n12704 DVSS.n12567 0.01445
R56837 DVSS.n12708 DVSS.n12567 0.01445
R56838 DVSS.n12709 DVSS.n12708 0.01445
R56839 DVSS.n12710 DVSS.n12709 0.01445
R56840 DVSS.n12710 DVSS.n12565 0.01445
R56841 DVSS.n12714 DVSS.n12565 0.01445
R56842 DVSS.n12715 DVSS.n12714 0.01445
R56843 DVSS.n12716 DVSS.n12715 0.01445
R56844 DVSS.n12716 DVSS.n12563 0.01445
R56845 DVSS.n12720 DVSS.n12563 0.01445
R56846 DVSS.n12721 DVSS.n12720 0.01445
R56847 DVSS.n12722 DVSS.n12721 0.01445
R56848 DVSS.n12722 DVSS.n12561 0.01445
R56849 DVSS.n12726 DVSS.n12561 0.01445
R56850 DVSS.n12727 DVSS.n12726 0.01445
R56851 DVSS.n12728 DVSS.n12727 0.01445
R56852 DVSS.n12728 DVSS.n12559 0.01445
R56853 DVSS.n12732 DVSS.n12559 0.01445
R56854 DVSS.n12733 DVSS.n12732 0.01445
R56855 DVSS.n12734 DVSS.n12733 0.01445
R56856 DVSS.n12734 DVSS.n12557 0.01445
R56857 DVSS.n12738 DVSS.n12557 0.01445
R56858 DVSS.n12739 DVSS.n12738 0.01445
R56859 DVSS.n12740 DVSS.n12739 0.01445
R56860 DVSS.n12740 DVSS.n12555 0.01445
R56861 DVSS.n12747 DVSS.n12555 0.01445
R56862 DVSS.n12770 DVSS.n12353 0.01445
R56863 DVSS.n12770 DVSS.n12356 0.01445
R56864 DVSS.n12603 DVSS.n12356 0.01445
R56865 DVSS.n12604 DVSS.n12603 0.01445
R56866 DVSS.n12605 DVSS.n12604 0.01445
R56867 DVSS.n12605 DVSS.n12600 0.01445
R56868 DVSS.n12609 DVSS.n12600 0.01445
R56869 DVSS.n12610 DVSS.n12609 0.01445
R56870 DVSS.n12611 DVSS.n12610 0.01445
R56871 DVSS.n12611 DVSS.n12598 0.01445
R56872 DVSS.n12615 DVSS.n12598 0.01445
R56873 DVSS.n12616 DVSS.n12615 0.01445
R56874 DVSS.n12617 DVSS.n12616 0.01445
R56875 DVSS.n12617 DVSS.n12596 0.01445
R56876 DVSS.n12621 DVSS.n12596 0.01445
R56877 DVSS.n12622 DVSS.n12621 0.01445
R56878 DVSS.n12623 DVSS.n12622 0.01445
R56879 DVSS.n12623 DVSS.n12594 0.01445
R56880 DVSS.n12627 DVSS.n12594 0.01445
R56881 DVSS.n12628 DVSS.n12627 0.01445
R56882 DVSS.n12629 DVSS.n12628 0.01445
R56883 DVSS.n12629 DVSS.n12592 0.01445
R56884 DVSS.n12633 DVSS.n12592 0.01445
R56885 DVSS.n12634 DVSS.n12633 0.01445
R56886 DVSS.n12635 DVSS.n12634 0.01445
R56887 DVSS.n12635 DVSS.n12590 0.01445
R56888 DVSS.n12639 DVSS.n12590 0.01445
R56889 DVSS.n12640 DVSS.n12639 0.01445
R56890 DVSS.n12641 DVSS.n12640 0.01445
R56891 DVSS.n12641 DVSS.n12588 0.01445
R56892 DVSS.n12645 DVSS.n12588 0.01445
R56893 DVSS.n12646 DVSS.n12645 0.01445
R56894 DVSS.n12647 DVSS.n12646 0.01445
R56895 DVSS.n12647 DVSS.n12586 0.01445
R56896 DVSS.n12651 DVSS.n12586 0.01445
R56897 DVSS.n12652 DVSS.n12651 0.01445
R56898 DVSS.n12653 DVSS.n12652 0.01445
R56899 DVSS.n12653 DVSS.n12584 0.01445
R56900 DVSS.n12657 DVSS.n12584 0.01445
R56901 DVSS.n12658 DVSS.n12657 0.01445
R56902 DVSS.n12659 DVSS.n12658 0.01445
R56903 DVSS.n12659 DVSS.n12582 0.01445
R56904 DVSS.n12663 DVSS.n12582 0.01445
R56905 DVSS.n12664 DVSS.n12663 0.01445
R56906 DVSS.n12665 DVSS.n12664 0.01445
R56907 DVSS.n12665 DVSS.n12580 0.01445
R56908 DVSS.n12669 DVSS.n12580 0.01445
R56909 DVSS.n12670 DVSS.n12669 0.01445
R56910 DVSS.n12671 DVSS.n12670 0.01445
R56911 DVSS.n12671 DVSS.n12578 0.01445
R56912 DVSS.n12675 DVSS.n12578 0.01445
R56913 DVSS.n12676 DVSS.n12675 0.01445
R56914 DVSS.n12677 DVSS.n12676 0.01445
R56915 DVSS.n12677 DVSS.n12576 0.01445
R56916 DVSS.n12681 DVSS.n12576 0.01445
R56917 DVSS.n12682 DVSS.n12681 0.01445
R56918 DVSS.n12683 DVSS.n12682 0.01445
R56919 DVSS.n12683 DVSS.n12574 0.01445
R56920 DVSS.n12687 DVSS.n12574 0.01445
R56921 DVSS.n12688 DVSS.n12687 0.01445
R56922 DVSS.n12689 DVSS.n12688 0.01445
R56923 DVSS.n12689 DVSS.n12572 0.01445
R56924 DVSS.n12693 DVSS.n12572 0.01445
R56925 DVSS.n12694 DVSS.n12693 0.01445
R56926 DVSS.n12695 DVSS.n12694 0.01445
R56927 DVSS.n12695 DVSS.n12570 0.01445
R56928 DVSS.n12699 DVSS.n12570 0.01445
R56929 DVSS.n12700 DVSS.n12699 0.01445
R56930 DVSS.n12701 DVSS.n12700 0.01445
R56931 DVSS.n12701 DVSS.n12568 0.01445
R56932 DVSS.n12705 DVSS.n12568 0.01445
R56933 DVSS.n12706 DVSS.n12705 0.01445
R56934 DVSS.n12707 DVSS.n12706 0.01445
R56935 DVSS.n12707 DVSS.n12566 0.01445
R56936 DVSS.n12711 DVSS.n12566 0.01445
R56937 DVSS.n12712 DVSS.n12711 0.01445
R56938 DVSS.n12713 DVSS.n12712 0.01445
R56939 DVSS.n12713 DVSS.n12564 0.01445
R56940 DVSS.n12717 DVSS.n12564 0.01445
R56941 DVSS.n12718 DVSS.n12717 0.01445
R56942 DVSS.n12719 DVSS.n12718 0.01445
R56943 DVSS.n12719 DVSS.n12562 0.01445
R56944 DVSS.n12723 DVSS.n12562 0.01445
R56945 DVSS.n12724 DVSS.n12723 0.01445
R56946 DVSS.n12725 DVSS.n12724 0.01445
R56947 DVSS.n12725 DVSS.n12560 0.01445
R56948 DVSS.n12729 DVSS.n12560 0.01445
R56949 DVSS.n12730 DVSS.n12729 0.01445
R56950 DVSS.n12731 DVSS.n12730 0.01445
R56951 DVSS.n12731 DVSS.n12558 0.01445
R56952 DVSS.n12735 DVSS.n12558 0.01445
R56953 DVSS.n12736 DVSS.n12735 0.01445
R56954 DVSS.n12737 DVSS.n12736 0.01445
R56955 DVSS.n12737 DVSS.n12556 0.01445
R56956 DVSS.n12741 DVSS.n12556 0.01445
R56957 DVSS.n12744 DVSS.n12741 0.01445
R56958 DVSS.n12746 DVSS.n12744 0.01445
R56959 DVSS.n6455 DVSS.n6247 0.01445
R56960 DVSS.n6455 DVSS.n6452 0.01445
R56961 DVSS.n6459 DVSS.n6452 0.01445
R56962 DVSS.n6460 DVSS.n6459 0.01445
R56963 DVSS.n6461 DVSS.n6460 0.01445
R56964 DVSS.n6461 DVSS.n6450 0.01445
R56965 DVSS.n6465 DVSS.n6450 0.01445
R56966 DVSS.n6466 DVSS.n6465 0.01445
R56967 DVSS.n6467 DVSS.n6466 0.01445
R56968 DVSS.n6467 DVSS.n6448 0.01445
R56969 DVSS.n6471 DVSS.n6448 0.01445
R56970 DVSS.n6472 DVSS.n6471 0.01445
R56971 DVSS.n6473 DVSS.n6472 0.01445
R56972 DVSS.n6473 DVSS.n6446 0.01445
R56973 DVSS.n6477 DVSS.n6446 0.01445
R56974 DVSS.n6478 DVSS.n6477 0.01445
R56975 DVSS.n6479 DVSS.n6478 0.01445
R56976 DVSS.n6479 DVSS.n6444 0.01445
R56977 DVSS.n6483 DVSS.n6444 0.01445
R56978 DVSS.n6484 DVSS.n6483 0.01445
R56979 DVSS.n6485 DVSS.n6484 0.01445
R56980 DVSS.n6485 DVSS.n6442 0.01445
R56981 DVSS.n6489 DVSS.n6442 0.01445
R56982 DVSS.n6490 DVSS.n6489 0.01445
R56983 DVSS.n6491 DVSS.n6490 0.01445
R56984 DVSS.n6491 DVSS.n6440 0.01445
R56985 DVSS.n6495 DVSS.n6440 0.01445
R56986 DVSS.n6496 DVSS.n6495 0.01445
R56987 DVSS.n6497 DVSS.n6496 0.01445
R56988 DVSS.n6497 DVSS.n6438 0.01445
R56989 DVSS.n6501 DVSS.n6438 0.01445
R56990 DVSS.n6502 DVSS.n6501 0.01445
R56991 DVSS.n6503 DVSS.n6502 0.01445
R56992 DVSS.n6503 DVSS.n6436 0.01445
R56993 DVSS.n6507 DVSS.n6436 0.01445
R56994 DVSS.n6508 DVSS.n6507 0.01445
R56995 DVSS.n6509 DVSS.n6508 0.01445
R56996 DVSS.n6509 DVSS.n6434 0.01445
R56997 DVSS.n6513 DVSS.n6434 0.01445
R56998 DVSS.n6514 DVSS.n6513 0.01445
R56999 DVSS.n6515 DVSS.n6514 0.01445
R57000 DVSS.n6515 DVSS.n6432 0.01445
R57001 DVSS.n6519 DVSS.n6432 0.01445
R57002 DVSS.n6520 DVSS.n6519 0.01445
R57003 DVSS.n6521 DVSS.n6520 0.01445
R57004 DVSS.n6521 DVSS.n6430 0.01445
R57005 DVSS.n6525 DVSS.n6430 0.01445
R57006 DVSS.n6526 DVSS.n6525 0.01445
R57007 DVSS.n6527 DVSS.n6526 0.01445
R57008 DVSS.n6527 DVSS.n6428 0.01445
R57009 DVSS.n6531 DVSS.n6428 0.01445
R57010 DVSS.n6532 DVSS.n6531 0.01445
R57011 DVSS.n6533 DVSS.n6532 0.01445
R57012 DVSS.n6533 DVSS.n6426 0.01445
R57013 DVSS.n6537 DVSS.n6426 0.01445
R57014 DVSS.n6538 DVSS.n6537 0.01445
R57015 DVSS.n6539 DVSS.n6538 0.01445
R57016 DVSS.n6539 DVSS.n6424 0.01445
R57017 DVSS.n6543 DVSS.n6424 0.01445
R57018 DVSS.n6544 DVSS.n6543 0.01445
R57019 DVSS.n6545 DVSS.n6544 0.01445
R57020 DVSS.n6545 DVSS.n6422 0.01445
R57021 DVSS.n6549 DVSS.n6422 0.01445
R57022 DVSS.n6550 DVSS.n6549 0.01445
R57023 DVSS.n6551 DVSS.n6550 0.01445
R57024 DVSS.n6551 DVSS.n6420 0.01445
R57025 DVSS.n6555 DVSS.n6420 0.01445
R57026 DVSS.n6556 DVSS.n6555 0.01445
R57027 DVSS.n6557 DVSS.n6556 0.01445
R57028 DVSS.n6557 DVSS.n6418 0.01445
R57029 DVSS.n6561 DVSS.n6418 0.01445
R57030 DVSS.n6562 DVSS.n6561 0.01445
R57031 DVSS.n6563 DVSS.n6562 0.01445
R57032 DVSS.n6563 DVSS.n6416 0.01445
R57033 DVSS.n6567 DVSS.n6416 0.01445
R57034 DVSS.n6568 DVSS.n6567 0.01445
R57035 DVSS.n6569 DVSS.n6568 0.01445
R57036 DVSS.n6569 DVSS.n6414 0.01445
R57037 DVSS.n6573 DVSS.n6414 0.01445
R57038 DVSS.n6574 DVSS.n6573 0.01445
R57039 DVSS.n6575 DVSS.n6574 0.01445
R57040 DVSS.n6575 DVSS.n6412 0.01445
R57041 DVSS.n6579 DVSS.n6412 0.01445
R57042 DVSS.n6580 DVSS.n6579 0.01445
R57043 DVSS.n6581 DVSS.n6580 0.01445
R57044 DVSS.n6581 DVSS.n6410 0.01445
R57045 DVSS.n6585 DVSS.n6410 0.01445
R57046 DVSS.n6586 DVSS.n6585 0.01445
R57047 DVSS.n6587 DVSS.n6586 0.01445
R57048 DVSS.n6587 DVSS.n6408 0.01445
R57049 DVSS.n6591 DVSS.n6408 0.01445
R57050 DVSS.n6592 DVSS.n6591 0.01445
R57051 DVSS.n6593 DVSS.n6592 0.01445
R57052 DVSS.n6593 DVSS.n6405 0.01445
R57053 DVSS.n6600 DVSS.n6405 0.01445
R57054 DVSS.n6600 DVSS.n6406 0.01445
R57055 DVSS.n6596 DVSS.n6406 0.01445
R57056 DVSS.n6456 DVSS.n6454 0.01445
R57057 DVSS.n6457 DVSS.n6456 0.01445
R57058 DVSS.n6458 DVSS.n6457 0.01445
R57059 DVSS.n6458 DVSS.n6451 0.01445
R57060 DVSS.n6462 DVSS.n6451 0.01445
R57061 DVSS.n6463 DVSS.n6462 0.01445
R57062 DVSS.n6464 DVSS.n6463 0.01445
R57063 DVSS.n6464 DVSS.n6449 0.01445
R57064 DVSS.n6468 DVSS.n6449 0.01445
R57065 DVSS.n6469 DVSS.n6468 0.01445
R57066 DVSS.n6470 DVSS.n6469 0.01445
R57067 DVSS.n6470 DVSS.n6447 0.01445
R57068 DVSS.n6474 DVSS.n6447 0.01445
R57069 DVSS.n6475 DVSS.n6474 0.01445
R57070 DVSS.n6476 DVSS.n6475 0.01445
R57071 DVSS.n6476 DVSS.n6445 0.01445
R57072 DVSS.n6480 DVSS.n6445 0.01445
R57073 DVSS.n6481 DVSS.n6480 0.01445
R57074 DVSS.n6482 DVSS.n6481 0.01445
R57075 DVSS.n6482 DVSS.n6443 0.01445
R57076 DVSS.n6486 DVSS.n6443 0.01445
R57077 DVSS.n6487 DVSS.n6486 0.01445
R57078 DVSS.n6488 DVSS.n6487 0.01445
R57079 DVSS.n6488 DVSS.n6441 0.01445
R57080 DVSS.n6492 DVSS.n6441 0.01445
R57081 DVSS.n6493 DVSS.n6492 0.01445
R57082 DVSS.n6494 DVSS.n6493 0.01445
R57083 DVSS.n6494 DVSS.n6439 0.01445
R57084 DVSS.n6498 DVSS.n6439 0.01445
R57085 DVSS.n6499 DVSS.n6498 0.01445
R57086 DVSS.n6500 DVSS.n6499 0.01445
R57087 DVSS.n6500 DVSS.n6437 0.01445
R57088 DVSS.n6504 DVSS.n6437 0.01445
R57089 DVSS.n6505 DVSS.n6504 0.01445
R57090 DVSS.n6506 DVSS.n6505 0.01445
R57091 DVSS.n6506 DVSS.n6435 0.01445
R57092 DVSS.n6510 DVSS.n6435 0.01445
R57093 DVSS.n6511 DVSS.n6510 0.01445
R57094 DVSS.n6512 DVSS.n6511 0.01445
R57095 DVSS.n6512 DVSS.n6433 0.01445
R57096 DVSS.n6516 DVSS.n6433 0.01445
R57097 DVSS.n6517 DVSS.n6516 0.01445
R57098 DVSS.n6518 DVSS.n6517 0.01445
R57099 DVSS.n6518 DVSS.n6431 0.01445
R57100 DVSS.n6522 DVSS.n6431 0.01445
R57101 DVSS.n6523 DVSS.n6522 0.01445
R57102 DVSS.n6524 DVSS.n6523 0.01445
R57103 DVSS.n6524 DVSS.n6429 0.01445
R57104 DVSS.n6528 DVSS.n6429 0.01445
R57105 DVSS.n6529 DVSS.n6528 0.01445
R57106 DVSS.n6530 DVSS.n6529 0.01445
R57107 DVSS.n6530 DVSS.n6427 0.01445
R57108 DVSS.n6534 DVSS.n6427 0.01445
R57109 DVSS.n6535 DVSS.n6534 0.01445
R57110 DVSS.n6536 DVSS.n6535 0.01445
R57111 DVSS.n6536 DVSS.n6425 0.01445
R57112 DVSS.n6540 DVSS.n6425 0.01445
R57113 DVSS.n6541 DVSS.n6540 0.01445
R57114 DVSS.n6542 DVSS.n6541 0.01445
R57115 DVSS.n6542 DVSS.n6423 0.01445
R57116 DVSS.n6546 DVSS.n6423 0.01445
R57117 DVSS.n6547 DVSS.n6546 0.01445
R57118 DVSS.n6548 DVSS.n6547 0.01445
R57119 DVSS.n6548 DVSS.n6421 0.01445
R57120 DVSS.n6552 DVSS.n6421 0.01445
R57121 DVSS.n6553 DVSS.n6552 0.01445
R57122 DVSS.n6554 DVSS.n6553 0.01445
R57123 DVSS.n6554 DVSS.n6419 0.01445
R57124 DVSS.n6558 DVSS.n6419 0.01445
R57125 DVSS.n6559 DVSS.n6558 0.01445
R57126 DVSS.n6560 DVSS.n6559 0.01445
R57127 DVSS.n6560 DVSS.n6417 0.01445
R57128 DVSS.n6564 DVSS.n6417 0.01445
R57129 DVSS.n6565 DVSS.n6564 0.01445
R57130 DVSS.n6566 DVSS.n6565 0.01445
R57131 DVSS.n6566 DVSS.n6415 0.01445
R57132 DVSS.n6570 DVSS.n6415 0.01445
R57133 DVSS.n6571 DVSS.n6570 0.01445
R57134 DVSS.n6572 DVSS.n6571 0.01445
R57135 DVSS.n6572 DVSS.n6413 0.01445
R57136 DVSS.n6576 DVSS.n6413 0.01445
R57137 DVSS.n6577 DVSS.n6576 0.01445
R57138 DVSS.n6578 DVSS.n6577 0.01445
R57139 DVSS.n6578 DVSS.n6411 0.01445
R57140 DVSS.n6582 DVSS.n6411 0.01445
R57141 DVSS.n6583 DVSS.n6582 0.01445
R57142 DVSS.n6584 DVSS.n6583 0.01445
R57143 DVSS.n6584 DVSS.n6409 0.01445
R57144 DVSS.n6588 DVSS.n6409 0.01445
R57145 DVSS.n6589 DVSS.n6588 0.01445
R57146 DVSS.n6590 DVSS.n6589 0.01445
R57147 DVSS.n6590 DVSS.n6407 0.01445
R57148 DVSS.n6594 DVSS.n6407 0.01445
R57149 DVSS.n6595 DVSS.n6594 0.01445
R57150 DVSS.n6599 DVSS.n6595 0.01445
R57151 DVSS.n6599 DVSS.n6598 0.01445
R57152 DVSS.n6598 DVSS.n6597 0.01445
R57153 DVSS.n18909 DVSS.n18880 0.0144045
R57154 DVSS.n20348 DVSS.n14691 0.0144045
R57155 DVSS.n12775 DVSS.n12773 0.0143045
R57156 DVSS.n22627 DVSS.n737 0.014281
R57157 DVSS.n22894 DVSS.n449 0.014281
R57158 DVSS.n7456 DVSS.n7455 0.014225
R57159 DVSS.n19315 DVSS.n19308 0.0141679
R57160 DVSS.n19039 DVSS.n19011 0.0141679
R57161 DVSS.n19028 DVSS.n19011 0.0141679
R57162 DVSS.n19038 DVSS.n19010 0.0141679
R57163 DVSS.n19027 DVSS.n19010 0.0141679
R57164 DVSS.n19037 DVSS.n19009 0.0141679
R57165 DVSS.n19026 DVSS.n19009 0.0141679
R57166 DVSS.n19036 DVSS.n19008 0.0141679
R57167 DVSS.n19025 DVSS.n19008 0.0141679
R57168 DVSS.n19035 DVSS.n19007 0.0141679
R57169 DVSS.n19024 DVSS.n19007 0.0141679
R57170 DVSS.n19034 DVSS.n19006 0.0141679
R57171 DVSS.n19023 DVSS.n19006 0.0141679
R57172 DVSS.n19033 DVSS.n19005 0.0141679
R57173 DVSS.n19022 DVSS.n19005 0.0141679
R57174 DVSS.n19897 DVSS.n19032 0.0141679
R57175 DVSS.n19898 DVSS.n19020 0.0141679
R57176 DVSS.n19224 DVSS.n19223 0.0141679
R57177 DVSS.n19225 DVSS.n19224 0.0141679
R57178 DVSS.n19226 DVSS.n19222 0.0141679
R57179 DVSS.n19228 DVSS.n19222 0.0141679
R57180 DVSS.n19229 DVSS.n19221 0.0141679
R57181 DVSS.n19231 DVSS.n19221 0.0141679
R57182 DVSS.n19232 DVSS.n19220 0.0141679
R57183 DVSS.n19234 DVSS.n19220 0.0141679
R57184 DVSS.n19235 DVSS.n19219 0.0141679
R57185 DVSS.n19237 DVSS.n19219 0.0141679
R57186 DVSS.n19238 DVSS.n19218 0.0141679
R57187 DVSS.n19240 DVSS.n19218 0.0141679
R57188 DVSS.n19241 DVSS.n19217 0.0141679
R57189 DVSS.n19243 DVSS.n19217 0.0141679
R57190 DVSS.n19246 DVSS.n19245 0.0141679
R57191 DVSS.n19248 DVSS.n19247 0.0141679
R57192 DVSS.n19597 DVSS.n19168 0.0141679
R57193 DVSS.n19599 DVSS.n19168 0.0141679
R57194 DVSS.n19600 DVSS.n19167 0.0141679
R57195 DVSS.n19602 DVSS.n19167 0.0141679
R57196 DVSS.n19603 DVSS.n19166 0.0141679
R57197 DVSS.n19605 DVSS.n19166 0.0141679
R57198 DVSS.n19606 DVSS.n19165 0.0141679
R57199 DVSS.n19608 DVSS.n19165 0.0141679
R57200 DVSS.n19609 DVSS.n19164 0.0141679
R57201 DVSS.n19611 DVSS.n19164 0.0141679
R57202 DVSS.n19612 DVSS.n19163 0.0141679
R57203 DVSS.n19614 DVSS.n19163 0.0141679
R57204 DVSS.n19615 DVSS.n19162 0.0141679
R57205 DVSS.n19617 DVSS.n19162 0.0141679
R57206 DVSS.n19620 DVSS.n19619 0.0141679
R57207 DVSS.n19622 DVSS.n19621 0.0141679
R57208 DVSS.n19625 DVSS.n19155 0.0141679
R57209 DVSS.n19627 DVSS.n19155 0.0141679
R57210 DVSS.n19628 DVSS.n19154 0.0141679
R57211 DVSS.n19630 DVSS.n19154 0.0141679
R57212 DVSS.n19631 DVSS.n19153 0.0141679
R57213 DVSS.n19633 DVSS.n19153 0.0141679
R57214 DVSS.n19634 DVSS.n19152 0.0141679
R57215 DVSS.n19636 DVSS.n19152 0.0141679
R57216 DVSS.n19637 DVSS.n19151 0.0141679
R57217 DVSS.n19639 DVSS.n19151 0.0141679
R57218 DVSS.n19640 DVSS.n19150 0.0141679
R57219 DVSS.n19642 DVSS.n19150 0.0141679
R57220 DVSS.n19643 DVSS.n19149 0.0141679
R57221 DVSS.n19645 DVSS.n19149 0.0141679
R57222 DVSS.n19648 DVSS.n19647 0.0141679
R57223 DVSS.n19650 DVSS.n19649 0.0141679
R57224 DVSS.n19657 DVSS.n19139 0.0141679
R57225 DVSS.n19312 DVSS.n19308 0.0141679
R57226 DVSS.n19039 DVSS.n19012 0.0141679
R57227 DVSS.n19038 DVSS.n19013 0.0141679
R57228 DVSS.n19037 DVSS.n19014 0.0141679
R57229 DVSS.n19036 DVSS.n19015 0.0141679
R57230 DVSS.n19035 DVSS.n19016 0.0141679
R57231 DVSS.n19034 DVSS.n19017 0.0141679
R57232 DVSS.n19033 DVSS.n19018 0.0141679
R57233 DVSS.n19032 DVSS.n19019 0.0141679
R57234 DVSS.n19223 DVSS.n19030 0.0141679
R57235 DVSS.n19227 DVSS.n19226 0.0141679
R57236 DVSS.n19230 DVSS.n19229 0.0141679
R57237 DVSS.n19233 DVSS.n19232 0.0141679
R57238 DVSS.n19236 DVSS.n19235 0.0141679
R57239 DVSS.n19239 DVSS.n19238 0.0141679
R57240 DVSS.n19242 DVSS.n19241 0.0141679
R57241 DVSS.n19245 DVSS.n19244 0.0141679
R57242 DVSS.n19598 DVSS.n19597 0.0141679
R57243 DVSS.n19601 DVSS.n19600 0.0141679
R57244 DVSS.n19604 DVSS.n19603 0.0141679
R57245 DVSS.n19607 DVSS.n19606 0.0141679
R57246 DVSS.n19610 DVSS.n19609 0.0141679
R57247 DVSS.n19613 DVSS.n19612 0.0141679
R57248 DVSS.n19616 DVSS.n19615 0.0141679
R57249 DVSS.n19619 DVSS.n19618 0.0141679
R57250 DVSS.n19028 DVSS.n19013 0.0141679
R57251 DVSS.n19027 DVSS.n19014 0.0141679
R57252 DVSS.n19026 DVSS.n19015 0.0141679
R57253 DVSS.n19025 DVSS.n19016 0.0141679
R57254 DVSS.n19024 DVSS.n19017 0.0141679
R57255 DVSS.n19023 DVSS.n19018 0.0141679
R57256 DVSS.n19022 DVSS.n19019 0.0141679
R57257 DVSS.n19227 DVSS.n19225 0.0141679
R57258 DVSS.n19230 DVSS.n19228 0.0141679
R57259 DVSS.n19233 DVSS.n19231 0.0141679
R57260 DVSS.n19236 DVSS.n19234 0.0141679
R57261 DVSS.n19239 DVSS.n19237 0.0141679
R57262 DVSS.n19242 DVSS.n19240 0.0141679
R57263 DVSS.n19244 DVSS.n19243 0.0141679
R57264 DVSS.n19601 DVSS.n19599 0.0141679
R57265 DVSS.n19604 DVSS.n19602 0.0141679
R57266 DVSS.n19607 DVSS.n19605 0.0141679
R57267 DVSS.n19610 DVSS.n19608 0.0141679
R57268 DVSS.n19613 DVSS.n19611 0.0141679
R57269 DVSS.n19616 DVSS.n19614 0.0141679
R57270 DVSS.n19618 DVSS.n19617 0.0141679
R57271 DVSS.n19021 DVSS.n19020 0.0141679
R57272 DVSS.n19248 DVSS.n19169 0.0141679
R57273 DVSS.n19622 DVSS.n19156 0.0141679
R57274 DVSS.n22429 DVSS.n1013 0.0141679
R57275 DVSS.n22429 DVSS.n1014 0.0141679
R57276 DVSS.n1025 DVSS.n1016 0.0141679
R57277 DVSS.n1027 DVSS.n1025 0.0141679
R57278 DVSS.n1051 DVSS.n1024 0.0141679
R57279 DVSS.n1029 DVSS.n1024 0.0141679
R57280 DVSS.n1050 DVSS.n1023 0.0141679
R57281 DVSS.n1031 DVSS.n1023 0.0141679
R57282 DVSS.n1049 DVSS.n1022 0.0141679
R57283 DVSS.n1033 DVSS.n1022 0.0141679
R57284 DVSS.n1048 DVSS.n1021 0.0141679
R57285 DVSS.n1035 DVSS.n1021 0.0141679
R57286 DVSS.n1047 DVSS.n1020 0.0141679
R57287 DVSS.n1037 DVSS.n1020 0.0141679
R57288 DVSS.n1046 DVSS.n1019 0.0141679
R57289 DVSS.n1039 DVSS.n1019 0.0141679
R57290 DVSS.n1045 DVSS.n1018 0.0141679
R57291 DVSS.n22381 DVSS.n1018 0.0141679
R57292 DVSS.n22382 DVSS.n1041 0.0141679
R57293 DVSS.n22366 DVSS.n22365 0.0141679
R57294 DVSS.n22365 DVSS.n1173 0.0141679
R57295 DVSS.n22364 DVSS.n22362 0.0141679
R57296 DVSS.n22362 DVSS.n1172 0.0141679
R57297 DVSS.n22361 DVSS.n22359 0.0141679
R57298 DVSS.n22359 DVSS.n1171 0.0141679
R57299 DVSS.n22358 DVSS.n22356 0.0141679
R57300 DVSS.n22356 DVSS.n1170 0.0141679
R57301 DVSS.n22355 DVSS.n22353 0.0141679
R57302 DVSS.n22353 DVSS.n1169 0.0141679
R57303 DVSS.n22352 DVSS.n22350 0.0141679
R57304 DVSS.n22350 DVSS.n1168 0.0141679
R57305 DVSS.n22349 DVSS.n22347 0.0141679
R57306 DVSS.n22347 DVSS.n1167 0.0141679
R57307 DVSS.n22346 DVSS.n22344 0.0141679
R57308 DVSS.n22344 DVSS.n1166 0.0141679
R57309 DVSS.n22368 DVSS.n22367 0.0141679
R57310 DVSS.n12971 DVSS.n12970 0.0141679
R57311 DVSS.n13064 DVSS.n12971 0.0141679
R57312 DVSS.n13065 DVSS.n12969 0.0141679
R57313 DVSS.n13067 DVSS.n12969 0.0141679
R57314 DVSS.n13068 DVSS.n12968 0.0141679
R57315 DVSS.n13070 DVSS.n12968 0.0141679
R57316 DVSS.n13071 DVSS.n12967 0.0141679
R57317 DVSS.n13073 DVSS.n12967 0.0141679
R57318 DVSS.n13074 DVSS.n12966 0.0141679
R57319 DVSS.n13076 DVSS.n12966 0.0141679
R57320 DVSS.n13077 DVSS.n12965 0.0141679
R57321 DVSS.n13079 DVSS.n12965 0.0141679
R57322 DVSS.n13080 DVSS.n12964 0.0141679
R57323 DVSS.n13082 DVSS.n12964 0.0141679
R57324 DVSS.n13083 DVSS.n12963 0.0141679
R57325 DVSS.n13085 DVSS.n12963 0.0141679
R57326 DVSS.n13087 DVSS.n13086 0.0141679
R57327 DVSS.n13090 DVSS.n12957 0.0141679
R57328 DVSS.n12957 DVSS.n12956 0.0141679
R57329 DVSS.n12954 DVSS.n12953 0.0141679
R57330 DVSS.n12953 DVSS.n12952 0.0141679
R57331 DVSS.n12950 DVSS.n12949 0.0141679
R57332 DVSS.n12949 DVSS.n12948 0.0141679
R57333 DVSS.n12946 DVSS.n12945 0.0141679
R57334 DVSS.n12945 DVSS.n12944 0.0141679
R57335 DVSS.n12942 DVSS.n12941 0.0141679
R57336 DVSS.n12941 DVSS.n12940 0.0141679
R57337 DVSS.n12938 DVSS.n12937 0.0141679
R57338 DVSS.n12937 DVSS.n12936 0.0141679
R57339 DVSS.n12934 DVSS.n12933 0.0141679
R57340 DVSS.n12933 DVSS.n12932 0.0141679
R57341 DVSS.n12930 DVSS.n12929 0.0141679
R57342 DVSS.n12929 DVSS.n12928 0.0141679
R57343 DVSS.n12926 DVSS.n12925 0.0141679
R57344 DVSS.n12925 DVSS.n12924 0.0141679
R57345 DVSS.n22430 DVSS.n1013 0.0141679
R57346 DVSS.n22432 DVSS.n1014 0.0141679
R57347 DVSS.n22386 DVSS.n1016 0.0141679
R57348 DVSS.n1051 DVSS.n1028 0.0141679
R57349 DVSS.n1050 DVSS.n1030 0.0141679
R57350 DVSS.n1049 DVSS.n1032 0.0141679
R57351 DVSS.n1048 DVSS.n1034 0.0141679
R57352 DVSS.n1047 DVSS.n1036 0.0141679
R57353 DVSS.n1046 DVSS.n1038 0.0141679
R57354 DVSS.n1045 DVSS.n1040 0.0141679
R57355 DVSS.n22366 DVSS.n1043 0.0141679
R57356 DVSS.n22364 DVSS.n22363 0.0141679
R57357 DVSS.n22361 DVSS.n22360 0.0141679
R57358 DVSS.n22358 DVSS.n22357 0.0141679
R57359 DVSS.n22355 DVSS.n22354 0.0141679
R57360 DVSS.n22352 DVSS.n22351 0.0141679
R57361 DVSS.n22349 DVSS.n22348 0.0141679
R57362 DVSS.n22346 DVSS.n22345 0.0141679
R57363 DVSS.n12970 DVSS.n1175 0.0141679
R57364 DVSS.n13066 DVSS.n13065 0.0141679
R57365 DVSS.n13069 DVSS.n13068 0.0141679
R57366 DVSS.n13072 DVSS.n13071 0.0141679
R57367 DVSS.n13075 DVSS.n13074 0.0141679
R57368 DVSS.n13078 DVSS.n13077 0.0141679
R57369 DVSS.n13081 DVSS.n13080 0.0141679
R57370 DVSS.n13084 DVSS.n13083 0.0141679
R57371 DVSS.n1028 DVSS.n1027 0.0141679
R57372 DVSS.n1030 DVSS.n1029 0.0141679
R57373 DVSS.n1032 DVSS.n1031 0.0141679
R57374 DVSS.n1034 DVSS.n1033 0.0141679
R57375 DVSS.n1036 DVSS.n1035 0.0141679
R57376 DVSS.n1038 DVSS.n1037 0.0141679
R57377 DVSS.n1040 DVSS.n1039 0.0141679
R57378 DVSS.n22382 DVSS.n22381 0.0141679
R57379 DVSS.n22363 DVSS.n1173 0.0141679
R57380 DVSS.n22360 DVSS.n1172 0.0141679
R57381 DVSS.n22357 DVSS.n1171 0.0141679
R57382 DVSS.n22354 DVSS.n1170 0.0141679
R57383 DVSS.n22351 DVSS.n1169 0.0141679
R57384 DVSS.n22348 DVSS.n1168 0.0141679
R57385 DVSS.n22345 DVSS.n1167 0.0141679
R57386 DVSS.n22368 DVSS.n1166 0.0141679
R57387 DVSS.n13066 DVSS.n13064 0.0141679
R57388 DVSS.n13069 DVSS.n13067 0.0141679
R57389 DVSS.n13072 DVSS.n13070 0.0141679
R57390 DVSS.n13075 DVSS.n13073 0.0141679
R57391 DVSS.n13078 DVSS.n13076 0.0141679
R57392 DVSS.n13081 DVSS.n13079 0.0141679
R57393 DVSS.n13084 DVSS.n13082 0.0141679
R57394 DVSS.n13086 DVSS.n13085 0.0141679
R57395 DVSS.n1042 DVSS.n1041 0.0141679
R57396 DVSS.n22367 DVSS.n1174 0.0141679
R57397 DVSS.n13087 DVSS.n12958 0.0141679
R57398 DVSS.n12955 DVSS.n12954 0.0141679
R57399 DVSS.n12951 DVSS.n12950 0.0141679
R57400 DVSS.n12947 DVSS.n12946 0.0141679
R57401 DVSS.n12943 DVSS.n12942 0.0141679
R57402 DVSS.n12939 DVSS.n12938 0.0141679
R57403 DVSS.n12935 DVSS.n12934 0.0141679
R57404 DVSS.n12931 DVSS.n12930 0.0141679
R57405 DVSS.n12927 DVSS.n12926 0.0141679
R57406 DVSS.n12956 DVSS.n12955 0.0141679
R57407 DVSS.n12952 DVSS.n12951 0.0141679
R57408 DVSS.n12948 DVSS.n12947 0.0141679
R57409 DVSS.n12944 DVSS.n12943 0.0141679
R57410 DVSS.n12940 DVSS.n12939 0.0141679
R57411 DVSS.n12936 DVSS.n12935 0.0141679
R57412 DVSS.n12932 DVSS.n12931 0.0141679
R57413 DVSS.n12928 DVSS.n12927 0.0141679
R57414 DVSS.n13094 DVSS.n12924 0.0141679
R57415 DVSS.n13091 DVSS.n13090 0.0141679
R57416 DVSS.n19626 DVSS.n19625 0.0141679
R57417 DVSS.n19629 DVSS.n19628 0.0141679
R57418 DVSS.n19632 DVSS.n19631 0.0141679
R57419 DVSS.n19635 DVSS.n19634 0.0141679
R57420 DVSS.n19638 DVSS.n19637 0.0141679
R57421 DVSS.n19641 DVSS.n19640 0.0141679
R57422 DVSS.n19644 DVSS.n19643 0.0141679
R57423 DVSS.n19647 DVSS.n19646 0.0141679
R57424 DVSS.n19629 DVSS.n19627 0.0141679
R57425 DVSS.n19632 DVSS.n19630 0.0141679
R57426 DVSS.n19635 DVSS.n19633 0.0141679
R57427 DVSS.n19638 DVSS.n19636 0.0141679
R57428 DVSS.n19641 DVSS.n19639 0.0141679
R57429 DVSS.n19644 DVSS.n19642 0.0141679
R57430 DVSS.n19646 DVSS.n19645 0.0141679
R57431 DVSS.n19650 DVSS.n19141 0.0141679
R57432 DVSS.n19653 DVSS.n19139 0.0141679
R57433 DVSS.n18908 DVSS.n18883 0.0141517
R57434 DVSS.n20438 DVSS.n14680 0.0141517
R57435 DVSS.n3857 DVSS.n3847 0.014059
R57436 DVSS.n3855 DVSS.n3850 0.014059
R57437 DVSS.n8609 DVSS.n8608 0.0140338
R57438 DVSS.n13126 DVSS.n13125 0.0140338
R57439 DVSS.n13102 DVSS.n12351 0.0140338
R57440 DVSS.n6687 DVSS.n5891 0.0140302
R57441 DVSS.n8092 DVSS.n4370 0.0140302
R57442 DVSS.n6686 DVSS.n5892 0.0140302
R57443 DVSS.n8093 DVSS.n4368 0.0140302
R57444 DVSS.n17388 DVSS.n17308 0.0138885
R57445 DVSS.n17399 DVSS.n17388 0.0138885
R57446 DVSS.n17389 DVSS.n17307 0.0138885
R57447 DVSS.n17397 DVSS.n17389 0.0138885
R57448 DVSS.n17390 DVSS.n17306 0.0138885
R57449 DVSS.n17395 DVSS.n17390 0.0138885
R57450 DVSS.n17393 DVSS.n17305 0.0138885
R57451 DVSS.n17386 DVSS.n17385 0.0138885
R57452 DVSS.n17273 DVSS.n17268 0.0138885
R57453 DVSS.n17291 DVSS.n17273 0.0138885
R57454 DVSS.n17274 DVSS.n17267 0.0138885
R57455 DVSS.n17289 DVSS.n17274 0.0138885
R57456 DVSS.n17275 DVSS.n17266 0.0138885
R57457 DVSS.n17287 DVSS.n17275 0.0138885
R57458 DVSS.n17276 DVSS.n17265 0.0138885
R57459 DVSS.n17285 DVSS.n17276 0.0138885
R57460 DVSS.n17277 DVSS.n17264 0.0138885
R57461 DVSS.n17283 DVSS.n17277 0.0138885
R57462 DVSS.n17278 DVSS.n17263 0.0138885
R57463 DVSS.n17281 DVSS.n17278 0.0138885
R57464 DVSS.n17279 DVSS.n17262 0.0138885
R57465 DVSS.n17271 DVSS.n17270 0.0138885
R57466 DVSS.n17238 DVSS.n17233 0.0138885
R57467 DVSS.n17256 DVSS.n17238 0.0138885
R57468 DVSS.n17239 DVSS.n17232 0.0138885
R57469 DVSS.n17254 DVSS.n17239 0.0138885
R57470 DVSS.n17240 DVSS.n17231 0.0138885
R57471 DVSS.n17252 DVSS.n17240 0.0138885
R57472 DVSS.n17241 DVSS.n17230 0.0138885
R57473 DVSS.n17250 DVSS.n17241 0.0138885
R57474 DVSS.n17242 DVSS.n17229 0.0138885
R57475 DVSS.n17248 DVSS.n17242 0.0138885
R57476 DVSS.n17243 DVSS.n17228 0.0138885
R57477 DVSS.n17246 DVSS.n17243 0.0138885
R57478 DVSS.n17244 DVSS.n17227 0.0138885
R57479 DVSS.n17236 DVSS.n17235 0.0138885
R57480 DVSS.n17220 DVSS.n17205 0.0138885
R57481 DVSS.n17222 DVSS.n17220 0.0138885
R57482 DVSS.n17217 DVSS.n17204 0.0138885
R57483 DVSS.n17219 DVSS.n17217 0.0138885
R57484 DVSS.n17214 DVSS.n17203 0.0138885
R57485 DVSS.n17216 DVSS.n17214 0.0138885
R57486 DVSS.n17211 DVSS.n17202 0.0138885
R57487 DVSS.n17213 DVSS.n17211 0.0138885
R57488 DVSS.n17419 DVSS.n17201 0.0138885
R57489 DVSS.n17421 DVSS.n17200 0.0138885
R57490 DVSS.n17379 DVSS.n17311 0.0138885
R57491 DVSS.n17376 DVSS.n17313 0.0138885
R57492 DVSS.n17373 DVSS.n17313 0.0138885
R57493 DVSS.n17374 DVSS.n17314 0.0138885
R57494 DVSS.n17331 DVSS.n17314 0.0138885
R57495 DVSS.n17324 DVSS.n17315 0.0138885
R57496 DVSS.n17330 DVSS.n17315 0.0138885
R57497 DVSS.n17322 DVSS.n17316 0.0138885
R57498 DVSS.n17329 DVSS.n17316 0.0138885
R57499 DVSS.n17320 DVSS.n17317 0.0138885
R57500 DVSS.n17328 DVSS.n17317 0.0138885
R57501 DVSS.n17334 DVSS.n17333 0.0138885
R57502 DVSS.n17357 DVSS.n17334 0.0138885
R57503 DVSS.n17367 DVSS.n17335 0.0138885
R57504 DVSS.n17355 DVSS.n17335 0.0138885
R57505 DVSS.n17365 DVSS.n17336 0.0138885
R57506 DVSS.n17353 DVSS.n17336 0.0138885
R57507 DVSS.n17364 DVSS.n17337 0.0138885
R57508 DVSS.n17351 DVSS.n17337 0.0138885
R57509 DVSS.n17363 DVSS.n17338 0.0138885
R57510 DVSS.n17349 DVSS.n17338 0.0138885
R57511 DVSS.n17362 DVSS.n17339 0.0138885
R57512 DVSS.n17347 DVSS.n17339 0.0138885
R57513 DVSS.n17361 DVSS.n17340 0.0138885
R57514 DVSS.n17345 DVSS.n17340 0.0138885
R57515 DVSS.n17360 DVSS.n17341 0.0138885
R57516 DVSS.n17343 DVSS.n17341 0.0138885
R57517 DVSS.n16952 DVSS.n16949 0.0138885
R57518 DVSS.n16972 DVSS.n16952 0.0138885
R57519 DVSS.n16953 DVSS.n16948 0.0138885
R57520 DVSS.n16970 DVSS.n16953 0.0138885
R57521 DVSS.n16954 DVSS.n16947 0.0138885
R57522 DVSS.n16968 DVSS.n16954 0.0138885
R57523 DVSS.n16955 DVSS.n16946 0.0138885
R57524 DVSS.n16966 DVSS.n16955 0.0138885
R57525 DVSS.n16956 DVSS.n16945 0.0138885
R57526 DVSS.n16964 DVSS.n16956 0.0138885
R57527 DVSS.n16957 DVSS.n16944 0.0138885
R57528 DVSS.n16962 DVSS.n16957 0.0138885
R57529 DVSS.n16958 DVSS.n16943 0.0138885
R57530 DVSS.n16960 DVSS.n16958 0.0138885
R57531 DVSS.n16959 DVSS.n16942 0.0138885
R57532 DVSS.n16959 DVSS.n16950 0.0138885
R57533 DVSS.n17519 DVSS.n17517 0.0138885
R57534 DVSS.n17519 DVSS.n17518 0.0138885
R57535 DVSS.n17516 DVSS.n17514 0.0138885
R57536 DVSS.n17516 DVSS.n17515 0.0138885
R57537 DVSS.n17513 DVSS.n17511 0.0138885
R57538 DVSS.n17513 DVSS.n17512 0.0138885
R57539 DVSS.n17510 DVSS.n17508 0.0138885
R57540 DVSS.n17510 DVSS.n17509 0.0138885
R57541 DVSS.n17507 DVSS.n17505 0.0138885
R57542 DVSS.n17507 DVSS.n17506 0.0138885
R57543 DVSS.n17504 DVSS.n17501 0.0138885
R57544 DVSS.n17480 DVSS.n17120 0.0138885
R57545 DVSS.n17126 DVSS.n17125 0.0138885
R57546 DVSS.n17296 DVSS.n17125 0.0138885
R57547 DVSS.n17128 DVSS.n17124 0.0138885
R57548 DVSS.n17297 DVSS.n17124 0.0138885
R57549 DVSS.n17130 DVSS.n17123 0.0138885
R57550 DVSS.n17298 DVSS.n17123 0.0138885
R57551 DVSS.n17132 DVSS.n17122 0.0138885
R57552 DVSS.n17300 DVSS.n17122 0.0138885
R57553 DVSS.n17137 DVSS.n17136 0.0138885
R57554 DVSS.n17476 DVSS.n17139 0.0138885
R57555 DVSS.n17162 DVSS.n17139 0.0138885
R57556 DVSS.n17164 DVSS.n17161 0.0138885
R57557 DVSS.n17161 DVSS.n17160 0.0138885
R57558 DVSS.n17158 DVSS.n17157 0.0138885
R57559 DVSS.n17157 DVSS.n17156 0.0138885
R57560 DVSS.n17154 DVSS.n17153 0.0138885
R57561 DVSS.n17153 DVSS.n17152 0.0138885
R57562 DVSS.n17150 DVSS.n17149 0.0138885
R57563 DVSS.n17149 DVSS.n17148 0.0138885
R57564 DVSS.n17146 DVSS.n17145 0.0138885
R57565 DVSS.n17145 DVSS.n17144 0.0138885
R57566 DVSS.n17165 DVSS.n17142 0.0138885
R57567 DVSS.n17166 DVSS.n17165 0.0138885
R57568 DVSS.n17172 DVSS.n17171 0.0138885
R57569 DVSS.n17182 DVSS.n17174 0.0138885
R57570 DVSS.n17183 DVSS.n17182 0.0138885
R57571 DVSS.n17465 DVSS.n17181 0.0138885
R57572 DVSS.n17185 DVSS.n17181 0.0138885
R57573 DVSS.n17464 DVSS.n17180 0.0138885
R57574 DVSS.n17187 DVSS.n17180 0.0138885
R57575 DVSS.n17463 DVSS.n17179 0.0138885
R57576 DVSS.n17189 DVSS.n17179 0.0138885
R57577 DVSS.n17462 DVSS.n17178 0.0138885
R57578 DVSS.n17191 DVSS.n17178 0.0138885
R57579 DVSS.n17461 DVSS.n17177 0.0138885
R57580 DVSS.n17193 DVSS.n17177 0.0138885
R57581 DVSS.n17460 DVSS.n17176 0.0138885
R57582 DVSS.n17466 DVSS.n17176 0.0138885
R57583 DVSS.n17198 DVSS.n17197 0.0138885
R57584 DVSS.n17432 DVSS.n17427 0.0138885
R57585 DVSS.n17435 DVSS.n17432 0.0138885
R57586 DVSS.n17449 DVSS.n17431 0.0138885
R57587 DVSS.n17437 DVSS.n17431 0.0138885
R57588 DVSS.n17448 DVSS.n17430 0.0138885
R57589 DVSS.n17439 DVSS.n17430 0.0138885
R57590 DVSS.n17447 DVSS.n17429 0.0138885
R57591 DVSS.n17441 DVSS.n17429 0.0138885
R57592 DVSS.n17446 DVSS.n17428 0.0138885
R57593 DVSS.n17450 DVSS.n17428 0.0138885
R57594 DVSS.n17370 DVSS.n17333 0.0138885
R57595 DVSS.n17368 DVSS.n17367 0.0138885
R57596 DVSS.n17365 DVSS.n17356 0.0138885
R57597 DVSS.n17364 DVSS.n17354 0.0138885
R57598 DVSS.n17363 DVSS.n17352 0.0138885
R57599 DVSS.n17362 DVSS.n17350 0.0138885
R57600 DVSS.n17361 DVSS.n17348 0.0138885
R57601 DVSS.n17360 DVSS.n17346 0.0138885
R57602 DVSS.n17368 DVSS.n17357 0.0138885
R57603 DVSS.n17356 DVSS.n17355 0.0138885
R57604 DVSS.n17354 DVSS.n17353 0.0138885
R57605 DVSS.n17352 DVSS.n17351 0.0138885
R57606 DVSS.n17350 DVSS.n17349 0.0138885
R57607 DVSS.n17348 DVSS.n17347 0.0138885
R57608 DVSS.n17346 DVSS.n17345 0.0138885
R57609 DVSS.n17344 DVSS.n17343 0.0138885
R57610 DVSS.n17405 DVSS.n17268 0.0138885
R57611 DVSS.n17292 DVSS.n17267 0.0138885
R57612 DVSS.n17290 DVSS.n17266 0.0138885
R57613 DVSS.n17288 DVSS.n17265 0.0138885
R57614 DVSS.n17286 DVSS.n17264 0.0138885
R57615 DVSS.n17284 DVSS.n17263 0.0138885
R57616 DVSS.n17282 DVSS.n17262 0.0138885
R57617 DVSS.n17292 DVSS.n17291 0.0138885
R57618 DVSS.n17290 DVSS.n17289 0.0138885
R57619 DVSS.n17288 DVSS.n17287 0.0138885
R57620 DVSS.n17286 DVSS.n17285 0.0138885
R57621 DVSS.n17284 DVSS.n17283 0.0138885
R57622 DVSS.n17282 DVSS.n17281 0.0138885
R57623 DVSS.n17270 DVSS.n17269 0.0138885
R57624 DVSS.n17477 DVSS.n17476 0.0138885
R57625 DVSS.n17164 DVSS.n17163 0.0138885
R57626 DVSS.n17159 DVSS.n17158 0.0138885
R57627 DVSS.n17155 DVSS.n17154 0.0138885
R57628 DVSS.n17151 DVSS.n17150 0.0138885
R57629 DVSS.n17147 DVSS.n17146 0.0138885
R57630 DVSS.n17143 DVSS.n17142 0.0138885
R57631 DVSS.n17474 DVSS.n17172 0.0138885
R57632 DVSS.n17167 DVSS.n17166 0.0138885
R57633 DVSS.n17144 DVSS.n17143 0.0138885
R57634 DVSS.n17148 DVSS.n17147 0.0138885
R57635 DVSS.n17152 DVSS.n17151 0.0138885
R57636 DVSS.n17156 DVSS.n17155 0.0138885
R57637 DVSS.n17160 DVSS.n17159 0.0138885
R57638 DVSS.n17163 DVSS.n17162 0.0138885
R57639 DVSS.n17489 DVSS.n16949 0.0138885
R57640 DVSS.n16973 DVSS.n16948 0.0138885
R57641 DVSS.n16971 DVSS.n16947 0.0138885
R57642 DVSS.n16969 DVSS.n16946 0.0138885
R57643 DVSS.n16967 DVSS.n16945 0.0138885
R57644 DVSS.n16965 DVSS.n16944 0.0138885
R57645 DVSS.n16963 DVSS.n16943 0.0138885
R57646 DVSS.n16961 DVSS.n16942 0.0138885
R57647 DVSS.n16973 DVSS.n16972 0.0138885
R57648 DVSS.n16971 DVSS.n16970 0.0138885
R57649 DVSS.n16969 DVSS.n16968 0.0138885
R57650 DVSS.n16967 DVSS.n16966 0.0138885
R57651 DVSS.n16965 DVSS.n16964 0.0138885
R57652 DVSS.n16963 DVSS.n16962 0.0138885
R57653 DVSS.n16961 DVSS.n16960 0.0138885
R57654 DVSS.n17491 DVSS.n16950 0.0138885
R57655 DVSS.n17413 DVSS.n17233 0.0138885
R57656 DVSS.n17257 DVSS.n17232 0.0138885
R57657 DVSS.n17255 DVSS.n17231 0.0138885
R57658 DVSS.n17253 DVSS.n17230 0.0138885
R57659 DVSS.n17251 DVSS.n17229 0.0138885
R57660 DVSS.n17249 DVSS.n17228 0.0138885
R57661 DVSS.n17247 DVSS.n17227 0.0138885
R57662 DVSS.n17257 DVSS.n17256 0.0138885
R57663 DVSS.n17255 DVSS.n17254 0.0138885
R57664 DVSS.n17253 DVSS.n17252 0.0138885
R57665 DVSS.n17251 DVSS.n17250 0.0138885
R57666 DVSS.n17249 DVSS.n17248 0.0138885
R57667 DVSS.n17247 DVSS.n17246 0.0138885
R57668 DVSS.n17235 DVSS.n17234 0.0138885
R57669 DVSS.n17471 DVSS.n17174 0.0138885
R57670 DVSS.n17465 DVSS.n17184 0.0138885
R57671 DVSS.n17464 DVSS.n17186 0.0138885
R57672 DVSS.n17463 DVSS.n17188 0.0138885
R57673 DVSS.n17462 DVSS.n17190 0.0138885
R57674 DVSS.n17461 DVSS.n17192 0.0138885
R57675 DVSS.n17460 DVSS.n17194 0.0138885
R57676 DVSS.n17469 DVSS.n17198 0.0138885
R57677 DVSS.n17467 DVSS.n17466 0.0138885
R57678 DVSS.n17194 DVSS.n17193 0.0138885
R57679 DVSS.n17192 DVSS.n17191 0.0138885
R57680 DVSS.n17190 DVSS.n17189 0.0138885
R57681 DVSS.n17188 DVSS.n17187 0.0138885
R57682 DVSS.n17186 DVSS.n17185 0.0138885
R57683 DVSS.n17184 DVSS.n17183 0.0138885
R57684 DVSS.n17377 DVSS.n17376 0.0138885
R57685 DVSS.n17375 DVSS.n17374 0.0138885
R57686 DVSS.n17325 DVSS.n17324 0.0138885
R57687 DVSS.n17323 DVSS.n17322 0.0138885
R57688 DVSS.n17321 DVSS.n17320 0.0138885
R57689 DVSS.n17377 DVSS.n17311 0.0138885
R57690 DVSS.n17375 DVSS.n17373 0.0138885
R57691 DVSS.n17331 DVSS.n17325 0.0138885
R57692 DVSS.n17330 DVSS.n17323 0.0138885
R57693 DVSS.n17329 DVSS.n17321 0.0138885
R57694 DVSS.n17328 DVSS.n17319 0.0138885
R57695 DVSS.n17391 DVSS.n17308 0.0138885
R57696 DVSS.n17400 DVSS.n17307 0.0138885
R57697 DVSS.n17398 DVSS.n17306 0.0138885
R57698 DVSS.n17396 DVSS.n17305 0.0138885
R57699 DVSS.n17400 DVSS.n17399 0.0138885
R57700 DVSS.n17398 DVSS.n17397 0.0138885
R57701 DVSS.n17396 DVSS.n17395 0.0138885
R57702 DVSS.n17385 DVSS.n17384 0.0138885
R57703 DVSS.n17127 DVSS.n17126 0.0138885
R57704 DVSS.n17129 DVSS.n17128 0.0138885
R57705 DVSS.n17131 DVSS.n17130 0.0138885
R57706 DVSS.n17133 DVSS.n17132 0.0138885
R57707 DVSS.n17478 DVSS.n17137 0.0138885
R57708 DVSS.n17300 DVSS.n17299 0.0138885
R57709 DVSS.n17298 DVSS.n17133 0.0138885
R57710 DVSS.n17297 DVSS.n17131 0.0138885
R57711 DVSS.n17296 DVSS.n17129 0.0138885
R57712 DVSS.n17127 DVSS.n17120 0.0138885
R57713 DVSS.n17518 DVSS.n17495 0.0138885
R57714 DVSS.n17515 DVSS.n17496 0.0138885
R57715 DVSS.n17512 DVSS.n17497 0.0138885
R57716 DVSS.n17509 DVSS.n17498 0.0138885
R57717 DVSS.n17506 DVSS.n17499 0.0138885
R57718 DVSS.n17517 DVSS.n17494 0.0138885
R57719 DVSS.n17514 DVSS.n17495 0.0138885
R57720 DVSS.n17511 DVSS.n17496 0.0138885
R57721 DVSS.n17508 DVSS.n17497 0.0138885
R57722 DVSS.n17505 DVSS.n17498 0.0138885
R57723 DVSS.n17501 DVSS.n17499 0.0138885
R57724 DVSS.n17222 DVSS.n17221 0.0138885
R57725 DVSS.n17219 DVSS.n17218 0.0138885
R57726 DVSS.n17216 DVSS.n17215 0.0138885
R57727 DVSS.n17213 DVSS.n17212 0.0138885
R57728 DVSS.n17418 DVSS.n17205 0.0138885
R57729 DVSS.n17221 DVSS.n17204 0.0138885
R57730 DVSS.n17218 DVSS.n17203 0.0138885
R57731 DVSS.n17215 DVSS.n17202 0.0138885
R57732 DVSS.n17212 DVSS.n17201 0.0138885
R57733 DVSS.n17420 DVSS.n17200 0.0138885
R57734 DVSS.n17457 DVSS.n17427 0.0138885
R57735 DVSS.n17449 DVSS.n17436 0.0138885
R57736 DVSS.n17448 DVSS.n17438 0.0138885
R57737 DVSS.n17447 DVSS.n17440 0.0138885
R57738 DVSS.n17446 DVSS.n17442 0.0138885
R57739 DVSS.n17451 DVSS.n17450 0.0138885
R57740 DVSS.n17442 DVSS.n17441 0.0138885
R57741 DVSS.n17440 DVSS.n17439 0.0138885
R57742 DVSS.n17438 DVSS.n17437 0.0138885
R57743 DVSS.n17436 DVSS.n17435 0.0138885
R57744 DVSS.n17392 DVSS.n17309 0.0138885
R57745 DVSS.n17394 DVSS.n17384 0.0138885
R57746 DVSS.n17404 DVSS.n17293 0.0138885
R57747 DVSS.n17280 DVSS.n17269 0.0138885
R57748 DVSS.n17409 DVSS.n17258 0.0138885
R57749 DVSS.n17245 DVSS.n17234 0.0138885
R57750 DVSS.n17417 DVSS.n17223 0.0138885
R57751 DVSS.n17422 DVSS.n17206 0.0138885
R57752 DVSS.n17208 DVSS.n17206 0.0138885
R57753 DVSS.n17371 DVSS.n17318 0.0138885
R57754 DVSS.n17342 DVSS.n16974 0.0138885
R57755 DVSS.n17493 DVSS.n16939 0.0138885
R57756 DVSS.n17503 DVSS.n17502 0.0138885
R57757 DVSS.n17502 DVSS.n17500 0.0138885
R57758 DVSS.n17299 DVSS.n17134 0.0138885
R57759 DVSS.n17168 DVSS.n17167 0.0138885
R57760 DVSS.n17467 DVSS.n17195 0.0138885
R57761 DVSS.n17451 DVSS.n17443 0.0138885
R57762 DVSS.n17454 DVSS.n17453 0.0138885
R57763 DVSS.n17272 DVSS.n17258 0.0138885
R57764 DVSS.n17280 DVSS.n17279 0.0138885
R57765 DVSS.n17358 DVSS.n17342 0.0138885
R57766 DVSS.n17169 DVSS.n17168 0.0138885
R57767 DVSS.n17237 DVSS.n17223 0.0138885
R57768 DVSS.n17245 DVSS.n17244 0.0138885
R57769 DVSS.n16951 DVSS.n16939 0.0138885
R57770 DVSS.n17458 DVSS.n17195 0.0138885
R57771 DVSS.n17387 DVSS.n17293 0.0138885
R57772 DVSS.n17394 DVSS.n17393 0.0138885
R57773 DVSS.n17392 DVSS.n17391 0.0138885
R57774 DVSS.n17326 DVSS.n17318 0.0138885
R57775 DVSS.n17294 DVSS.n17134 0.0138885
R57776 DVSS.n17500 DVSS.n16935 0.0138885
R57777 DVSS.n17504 DVSS.n17503 0.0138885
R57778 DVSS.n17208 DVSS.n17207 0.0138885
R57779 DVSS.n17422 DVSS.n17421 0.0138885
R57780 DVSS.n17455 DVSS.n17454 0.0138885
R57781 DVSS.n17444 DVSS.n17443 0.0138885
R57782 DVSS.n14790 DVSS 0.0138618
R57783 DVSS.n9194 DVSS.n2784 0.013775
R57784 DVSS.n11640 DVSS.n11453 0.013775
R57785 DVSS.n18826 DVSS 0.0137264
R57786 DVSS.n18982 DVSS.n18915 0.0136461
R57787 DVSS.n20129 DVSS.n20059 0.0136461
R57788 DVSS.n20141 DVSS.n20060 0.0136461
R57789 DVSS.n20286 DVSS.n20216 0.0136461
R57790 DVSS.n20215 DVSS.n20214 0.0136461
R57791 DVSS.n20383 DVSS.n14686 0.0136461
R57792 DVSS.n17822 DVSS.n15888 0.0135737
R57793 DVSS.n15564 DVSS.n15536 0.0135737
R57794 DVSS.n8120 DVSS.n4013 0.013547
R57795 DVSS.n8119 DVSS.n4016 0.013547
R57796 DVSS.n19196 DVSS.n19195 0.0135263
R57797 DVSS.n7065 DVSS.n5179 0.0134925
R57798 DVSS.n7447 DVSS.n7446 0.0134925
R57799 DVSS.n20641 DVSS.n20640 0.0133933
R57800 DVSS.n9193 DVSS.n9192 0.013325
R57801 DVSS.n11986 DVSS.n11985 0.013325
R57802 DVSS.n21470 DVSS.n21448 0.0131563
R57803 DVSS.n21471 DVSS.n21470 0.0131563
R57804 DVSS.n22580 DVSS.n754 0.0131563
R57805 DVSS.n22576 DVSS.n754 0.0131563
R57806 DVSS.n22576 DVSS.n22575 0.0131563
R57807 DVSS.n22575 DVSS.n22574 0.0131563
R57808 DVSS.n22574 DVSS.n756 0.0131563
R57809 DVSS.n21453 DVSS.n756 0.0131563
R57810 DVSS.n21454 DVSS.n21453 0.0131563
R57811 DVSS.n21457 DVSS.n21454 0.0131563
R57812 DVSS.n22603 DVSS.n22602 0.0131563
R57813 DVSS.n22602 DVSS.n22601 0.0131563
R57814 DVSS.n22601 DVSS.n747 0.0131563
R57815 DVSS.n22597 DVSS.n747 0.0131563
R57816 DVSS.n22597 DVSS.n22596 0.0131563
R57817 DVSS.n22596 DVSS.n22595 0.0131563
R57818 DVSS.n22595 DVSS.n749 0.0131563
R57819 DVSS.n22591 DVSS.n749 0.0131563
R57820 DVSS.n22622 DVSS.n739 0.0131563
R57821 DVSS.n22618 DVSS.n739 0.0131563
R57822 DVSS.n22618 DVSS.n22617 0.0131563
R57823 DVSS.n22617 DVSS.n22616 0.0131563
R57824 DVSS.n22616 DVSS.n741 0.0131563
R57825 DVSS.n22612 DVSS.n741 0.0131563
R57826 DVSS.n22612 DVSS.n22611 0.0131563
R57827 DVSS.n22611 DVSS.n22610 0.0131563
R57828 DVSS.n22635 DVSS.n22634 0.0131563
R57829 DVSS.n15131 DVSS.n15128 0.0131563
R57830 DVSS.n15128 DVSS.n14314 0.0131563
R57831 DVSS.n20993 DVSS.n14311 0.0131563
R57832 DVSS.n20994 DVSS.n20993 0.0131563
R57833 DVSS.n21023 DVSS.n20994 0.0131563
R57834 DVSS.n21023 DVSS.n21022 0.0131563
R57835 DVSS.n21022 DVSS.n21021 0.0131563
R57836 DVSS.n21021 DVSS.n20995 0.0131563
R57837 DVSS.n21017 DVSS.n20995 0.0131563
R57838 DVSS.n21017 DVSS.n21016 0.0131563
R57839 DVSS.n21004 DVSS.n21001 0.0131563
R57840 DVSS.n21001 DVSS.n13371 0.0131563
R57841 DVSS.n22888 DVSS.n452 0.0131563
R57842 DVSS.n22899 DVSS.n447 0.0131563
R57843 DVSS.n22903 DVSS.n447 0.0131563
R57844 DVSS.n22904 DVSS.n22903 0.0131563
R57845 DVSS.n22905 DVSS.n22904 0.0131563
R57846 DVSS.n22905 DVSS.n445 0.0131563
R57847 DVSS.n22909 DVSS.n445 0.0131563
R57848 DVSS.n22910 DVSS.n22909 0.0131563
R57849 DVSS.n22911 DVSS.n22910 0.0131563
R57850 DVSS.n22919 DVSS.n22918 0.0131563
R57851 DVSS.n22920 DVSS.n22919 0.0131563
R57852 DVSS.n22920 DVSS.n439 0.0131563
R57853 DVSS.n22924 DVSS.n439 0.0131563
R57854 DVSS.n22925 DVSS.n22924 0.0131563
R57855 DVSS.n22926 DVSS.n22925 0.0131563
R57856 DVSS.n22926 DVSS.n437 0.0131563
R57857 DVSS.n22930 DVSS.n437 0.0131563
R57858 DVSS.n22941 DVSS.n432 0.0131563
R57859 DVSS.n22945 DVSS.n432 0.0131563
R57860 DVSS.n22946 DVSS.n22945 0.0131563
R57861 DVSS.n22947 DVSS.n22946 0.0131563
R57862 DVSS.n22947 DVSS.n430 0.0131563
R57863 DVSS.n22952 DVSS.n430 0.0131563
R57864 DVSS.n22953 DVSS.n22952 0.0131563
R57865 DVSS.n22954 DVSS.n22953 0.0131563
R57866 DVSS.n22968 DVSS.n424 0.0131563
R57867 DVSS.n22969 DVSS.n22968 0.0131563
R57868 DVSS.n18953 DVSS.n18910 0.0131404
R57869 DVSS.n20346 DVSS.n14681 0.0131404
R57870 DVSS.n2717 DVSS.n2707 0.0130638
R57871 DVSS.n10459 DVSS.n2021 0.0130638
R57872 DVSS.n2715 DVSS.n2710 0.0130638
R57873 DVSS.n10458 DVSS.n2023 0.0130638
R57874 DVSS.n18510 DVSS.n18505 0.0130581
R57875 DVSS.n15134 DVSS.n15126 0.0130581
R57876 DVSS.n21007 DVSS.n20999 0.0130581
R57877 DVSS.n8985 DVSS.n8983 0.0129511
R57878 DVSS.n13344 DVSS.n11106 0.0129511
R57879 DVSS.n18897 DVSS.n18881 0.0128876
R57880 DVSS.n20338 DVSS.n14692 0.0128876
R57881 DVSS.n7095 DVSS.n7094 0.012875
R57882 DVSS.n6669 DVSS.n6240 0.0128221
R57883 DVSS.n6668 DVSS.n6241 0.0128221
R57884 DVSS.n14799 DVSS.n14740 0.0127867
R57885 DVSS.n18820 DVSS.n18819 0.0126622
R57886 DVSS.n20055 DVSS.n14579 0.0126348
R57887 DVSS.n17907 DVSS.n15795 0.0126171
R57888 DVSS.n17948 DVSS.n15538 0.0126171
R57889 DVSS.n17864 DVSS.n15848 0.0126171
R57890 DVSS.n18045 DVSS.n15537 0.0126171
R57891 DVSS.n8606 DVSS.n3414 0.0125805
R57892 DVSS.n13123 DVSS.n11628 0.0125805
R57893 DVSS.n8607 DVSS.n3412 0.0125805
R57894 DVSS.n13124 DVSS.n11626 0.0125805
R57895 DVSS.n7453 DVSS.n4826 0.0124869
R57896 DVSS.n7454 DVSS.n4827 0.0124869
R57897 DVSS.n3041 DVSS.n2875 0.0124098
R57898 DVSS.n1612 DVSS.n1505 0.0124098
R57899 DVSS.n18983 DVSS.n18914 0.012382
R57900 DVSS.n20094 DVSS.n20053 0.012382
R57901 DVSS.n20306 DVSS.n20208 0.012382
R57902 DVSS.n20385 DVSS.n14685 0.012382
R57903 DVSS.n16200 DVSS 0.012365
R57904 DVSS DVSS.n16451 0.012365
R57905 DVSS.n12349 DVSS.n12348 0.0123125
R57906 DVSS.n12751 DVSS.n12749 0.0123125
R57907 DVSS.n6663 DVSS.n6241 0.0123125
R57908 DVSS.n6662 DVSS.n6240 0.0123125
R57909 DVSS.n17051 DVSS.n16977 0.0122568
R57910 DVSS.n16979 DVSS.n16978 0.0122568
R57911 DVSS.n17116 DVSS.n17056 0.0122568
R57912 DVSS.n17529 DVSS.n17528 0.0122568
R57913 DVSS.n18890 DVSS.n14558 0.0122391
R57914 DVSS.n18961 DVSS.n14563 0.0122391
R57915 DVSS.n20086 DVSS.n14596 0.0122391
R57916 DVSS.n20167 DVSS.n20166 0.0122391
R57917 DVSS.n20648 DVSS.n14632 0.0122391
R57918 DVSS.n20292 DVSS.n14646 0.0122391
R57919 DVSS.n20418 DVSS.n20417 0.0122391
R57920 DVSS.n20452 DVSS.n20448 0.0122391
R57921 DVSS.n18895 DVSS.n14527 0.0122391
R57922 DVSS.n18949 DVSS.n14530 0.0122391
R57923 DVSS.n20090 DVSS.n20021 0.0122391
R57924 DVSS.n20171 DVSS.n20027 0.0122391
R57925 DVSS.n20262 DVSS.n14873 0.0122391
R57926 DVSS.n20233 DVSS.n20191 0.0122391
R57927 DVSS.n20373 DVSS.n20329 0.0122391
R57928 DVSS.n20457 DVSS.n20456 0.0122391
R57929 DVSS.n7067 DVSS.n5181 0.0120973
R57930 DVSS.n4834 DVSS.n4824 0.0120973
R57931 DVSS.n7066 DVSS.n5180 0.0120973
R57932 DVSS.n7445 DVSS.n4836 0.0120973
R57933 DVSS.n2881 DVSS.n2786 0.0120939
R57934 DVSS.n11642 DVSS.n11456 0.0120939
R57935 DVSS.n2883 DVSS.n2785 0.0120939
R57936 DVSS.n11641 DVSS.n11454 0.0120939
R57937 DVSS.n12765 DVSS.n12747 0.011975
R57938 DVSS.n6597 DVSS.n6234 0.011975
R57939 DVSS.n22586 DVSS.n751 0.0119373
R57940 DVSS.n22935 DVSS.n435 0.0119373
R57941 DVSS.n19914 DVSS.n19913 0.0119115
R57942 DVSS.n18529 DVSS.n18528 0.0119115
R57943 DVSS.n18955 DVSS.n18879 0.0118764
R57944 DVSS.n20157 DVSS.n20156 0.0118764
R57945 DVSS.n20220 DVSS.n14625 0.0118764
R57946 DVSS.n20424 DVSS.n14690 0.0118764
R57947 DVSS.n7039 DVSS.n7038 0.0118684
R57948 DVSS.n7822 DVSS.n7821 0.0118684
R57949 DVSS.n22581 DVSS.n22580 0.01175
R57950 DVSS.n22941 DVSS.n22940 0.01175
R57951 DVSS.n2889 DVSS.n2879 0.0117009
R57952 DVSS.n11983 DVSS.n11645 0.0117009
R57953 DVSS.n2887 DVSS.n2882 0.0117009
R57954 DVSS.n11984 DVSS.n11639 0.0117009
R57955 DVSS.n18882 DVSS.n18872 0.0116236
R57956 DVSS.n20337 DVSS.n14693 0.0116236
R57957 DVSS.n8987 DVSS.n3044 0.0116141
R57958 DVSS.n13342 DVSS.n11108 0.0116141
R57959 DVSS.n8986 DVSS.n3047 0.0116141
R57960 DVSS.n13343 DVSS.n11107 0.0116141
R57961 DVSS.n6676 DVSS.n5885 0.011525
R57962 DVSS.n22634 DVSS.n735 0.0115156
R57963 DVSS.n22889 DVSS.n22888 0.0115156
R57964 DVSS.n4011 DVSS.n4010 0.0114624
R57965 DVSS.n8129 DVSS.n8128 0.0113271
R57966 DVSS.n7092 DVSS.n4883 0.0113079
R57967 DVSS.n7093 DVSS.n7091 0.0113079
R57968 DVSS.n9201 DVSS.n9200 0.0111309
R57969 DVSS.n1614 DVSS.n1509 0.0111309
R57970 DVSS.n9205 DVSS.n2876 0.0111309
R57971 DVSS.n10505 DVSS.n1507 0.0111309
R57972 DVSS.n18969 DVSS.n18876 0.011118
R57973 DVSS.n20092 DVSS.n20058 0.011118
R57974 DVSS.n20062 DVSS.n20061 0.011118
R57975 DVSS.n20247 DVSS.n20217 0.011118
R57976 DVSS.n20305 DVSS.n20210 0.011118
R57977 DVSS.n20406 DVSS.n14687 0.011118
R57978 DVSS.n8327 DVSS.n3751 0.011075
R57979 DVSS.n15136 DVSS.n15126 0.0110469
R57980 DVSS.n21009 DVSS.n20999 0.0110469
R57981 DVSS.n20988 DVSS.n14311 0.0108125
R57982 DVSS.n10146 DVSS.n2367 0.0107857
R57983 DVSS.n10148 DVSS.n2024 0.0107857
R57984 DVSS.n22629 DVSS.n22628 0.0107654
R57985 DVSS.n22893 DVSS.n450 0.0107654
R57986 DVSS.n22231 DVSS.n22230 0.0106562
R57987 DVSS.n22233 DVSS.n22231 0.0106562
R57988 DVSS.n5877 DVSS.n5868 0.0106477
R57989 DVSS.n7819 DVSS.n4472 0.0106477
R57990 DVSS.n5875 DVSS.n5870 0.0106477
R57991 DVSS.n7820 DVSS.n4473 0.0106477
R57992 DVSS.n10159 DVSS.n10158 0.010625
R57993 DVSS.n10491 DVSS.n10490 0.010625
R57994 DVSS.n18957 DVSS.n18911 0.0106124
R57995 DVSS.n20049 DVSS.n20044 0.0106124
R57996 DVSS.n20261 DVSS.n20221 0.0106124
R57997 DVSS.n20422 DVSS.n14682 0.0106124
R57998 DVSS.n5621 DVSS.n5529 0.0105588
R57999 DVSS.n7048 DVSS.n5576 0.0105588
R58000 DVSS.n5573 DVSS.n5530 0.0105588
R58001 DVSS.n7058 DVSS.n5575 0.0105588
R58002 DVSS.n5271 DVSS.n5180 0.0105588
R58003 DVSS.n5520 DVSS.n5186 0.0105588
R58004 DVSS.n5272 DVSS.n5181 0.0105588
R58005 DVSS.n5519 DVSS.n5185 0.0105588
R58006 DVSS.n4930 DVSS.n4838 0.0105588
R58007 DVSS.n7091 DVSS.n4884 0.0105588
R58008 DVSS.n4882 DVSS.n4839 0.0105588
R58009 DVSS.n7101 DVSS.n4883 0.0105588
R58010 DVSS.n7443 DVSS.n4836 0.0105588
R58011 DVSS.n7235 DVSS.n4827 0.0105588
R58012 DVSS.n7442 DVSS.n4834 0.0105588
R58013 DVSS.n7234 DVSS.n4826 0.0105588
R58014 DVSS.n7792 DVSS.n4820 0.0105588
R58015 DVSS.n7547 DVSS.n4813 0.0105588
R58016 DVSS.n7793 DVSS.n4819 0.0105588
R58017 DVSS.n7546 DVSS.n4812 0.0105588
R58018 DVSS.n4806 DVSS.n4473 0.0105588
R58019 DVSS.n4598 DVSS.n4465 0.0105588
R58020 DVSS.n4805 DVSS.n4472 0.0105588
R58021 DVSS.n4597 DVSS.n4467 0.0105588
R58022 DVSS.n8087 DVSS.n4368 0.0105588
R58023 DVSS.n7842 DVSS.n4459 0.0105588
R58024 DVSS.n8088 DVSS.n4370 0.0105588
R58025 DVSS.n7841 DVSS.n7840 0.0105588
R58026 DVSS.n4108 DVSS.n4016 0.0105588
R58027 DVSS.n4357 DVSS.n4024 0.0105588
R58028 DVSS.n4109 DVSS.n4013 0.0105588
R58029 DVSS.n4356 DVSS.n4023 0.0105588
R58030 DVSS.n8124 DVSS.n3903 0.0105588
R58031 DVSS.n8315 DVSS.n3855 0.0105588
R58032 DVSS.n8318 DVSS.n3902 0.0105588
R58033 DVSS.n8316 DVSS.n3857 0.0105588
R58034 DVSS.n8339 DVSS.n8338 0.0105588
R58035 DVSS.n3798 DVSS.n3752 0.0105588
R58036 DVSS.n8334 DVSS.n3797 0.0105588
R58037 DVSS.n8587 DVSS.n3753 0.0105588
R58038 DVSS.n3459 DVSS.n3412 0.0105588
R58039 DVSS.n8599 DVSS.n8598 0.0105588
R58040 DVSS.n8602 DVSS.n3414 0.0105588
R58041 DVSS.n8600 DVSS.n3502 0.0105588
R58042 DVSS.n3152 DVSS.n3061 0.0105588
R58043 DVSS.n3401 DVSS.n3068 0.0105588
R58044 DVSS.n3153 DVSS.n3060 0.0105588
R58045 DVSS.n3400 DVSS.n3067 0.0105588
R58046 DVSS.n8966 DVSS.n3047 0.0105588
R58047 DVSS.n8721 DVSS.n3054 0.0105588
R58048 DVSS.n8967 DVSS.n3044 0.0105588
R58049 DVSS.n8720 DVSS.n3053 0.0105588
R58050 DVSS.n8991 DVSS.n2935 0.0105588
R58051 DVSS.n9182 DVSS.n2887 0.0105588
R58052 DVSS.n9185 DVSS.n2934 0.0105588
R58053 DVSS.n9183 DVSS.n2889 0.0105588
R58054 DVSS.n9206 DVSS.n9205 0.0105588
R58055 DVSS.n2830 DVSS.n2785 0.0105588
R58056 DVSS.n9201 DVSS.n2829 0.0105588
R58057 DVSS.n9454 DVSS.n2786 0.0105588
R58058 DVSS.n9756 DVSS.n2736 0.0105588
R58059 DVSS.n9511 DVSS.n2726 0.0105588
R58060 DVSS.n9757 DVSS.n2738 0.0105588
R58061 DVSS.n9510 DVSS.n2727 0.0105588
R58062 DVSS.n9859 DVSS.n2715 0.0105588
R58063 DVSS.n10108 DVSS.n2724 0.0105588
R58064 DVSS.n9860 DVSS.n2717 0.0105588
R58065 DVSS.n10107 DVSS.n2722 0.0105588
R58066 DVSS.n2459 DVSS.n2368 0.0105588
R58067 DVSS.n10130 DVSS.n2414 0.0105588
R58068 DVSS.n2412 DVSS.n2369 0.0105588
R58069 DVSS.n10140 DVSS.n2413 0.0105588
R58070 DVSS.n2117 DVSS.n2025 0.0105588
R58071 DVSS.n10155 DVSS.n2072 0.0105588
R58072 DVSS.n2069 DVSS.n2026 0.0105588
R58073 DVSS.n10165 DVSS.n2071 0.0105588
R58074 DVSS.n10454 DVSS.n2023 0.0105588
R58075 DVSS.n10464 DVSS.n2011 0.0105588
R58076 DVSS.n2021 DVSS.n2009 0.0105588
R58077 DVSS.n10474 DVSS.n2010 0.0105588
R58078 DVSS.n1958 DVSS.n1617 0.0105588
R58079 DVSS.n1713 DVSS.n1622 0.0105588
R58080 DVSS.n1959 DVSS.n1618 0.0105588
R58081 DVSS.n1712 DVSS.n1621 0.0105588
R58082 DVSS.n10506 DVSS.n10505 0.0105588
R58083 DVSS.n1567 DVSS.n1520 0.0105588
R58084 DVSS.n1614 DVSS.n1565 0.0105588
R58085 DVSS.n10753 DVSS.n1522 0.0105588
R58086 DVSS.n11103 DVSS.n10769 0.0105588
R58087 DVSS.n10895 DVSS.n1516 0.0105588
R58088 DVSS.n11102 DVSS.n10767 0.0105588
R58089 DVSS.n10894 DVSS.n1514 0.0105588
R58090 DVSS.n11155 DVSS.n11107 0.0105588
R58091 DVSS.n13335 DVSS.n13334 0.0105588
R58092 DVSS.n13338 DVSS.n11108 0.0105588
R58093 DVSS.n13336 DVSS.n11199 0.0105588
R58094 DVSS.n11619 DVSS.n11503 0.0105588
R58095 DVSS.n13321 DVSS.n11454 0.0105588
R58096 DVSS.n13324 DVSS.n11502 0.0105588
R58097 DVSS.n13322 DVSS.n11456 0.0105588
R58098 DVSS.n11688 DVSS.n11628 0.0105588
R58099 DVSS.n11979 DVSS.n11645 0.0105588
R58100 DVSS.n6778 DVSS.n5875 0.0105588
R58101 DVSS.n7026 DVSS.n5884 0.0105588
R58102 DVSS.n6777 DVSS.n5877 0.0105588
R58103 DVSS.n7025 DVSS.n5882 0.0105588
R58104 DVSS.n12044 DVSS.n12002 0.0105588
R58105 DVSS.n12335 DVSS.n11992 0.0105588
R58106 DVSS.n5938 DVSS.n5891 0.0105588
R58107 DVSS.n5983 DVSS.n5887 0.0105588
R58108 DVSS.n5940 DVSS.n5892 0.0105588
R58109 DVSS.n5984 DVSS.n5886 0.0105588
R58110 DVSS.n11730 DVSS.n11626 0.0105588
R58111 DVSS.n11978 DVSS.n11639 0.0105588
R58112 DVSS.n12087 DVSS.n12001 0.0105588
R58113 DVSS.n12334 DVSS.n11990 0.0105588
R58114 DVSS.n17797 DVSS.n17795 0.0105
R58115 DVSS.n17797 DVSS.n15915 0.0105
R58116 DVSS.n17802 DVSS.n15915 0.0105
R58117 DVSS.n17804 DVSS.n17802 0.0105
R58118 DVSS.n17806 DVSS.n17804 0.0105
R58119 DVSS.n17806 DVSS.n15912 0.0105
R58120 DVSS.n17811 DVSS.n15912 0.0105
R58121 DVSS.n17813 DVSS.n17811 0.0105
R58122 DVSS.n17815 DVSS.n17813 0.0105
R58123 DVSS.n17815 DVSS.n15909 0.0105
R58124 DVSS.n17819 DVSS.n15909 0.0105
R58125 DVSS.n17819 DVSS.n15877 0.0105
R58126 DVSS.n17825 DVSS.n15877 0.0105
R58127 DVSS.n17825 DVSS.n15875 0.0105
R58128 DVSS.n17830 DVSS.n15875 0.0105
R58129 DVSS.n17830 DVSS.n15873 0.0105
R58130 DVSS.n17834 DVSS.n15873 0.0105
R58131 DVSS.n17836 DVSS.n17834 0.0105
R58132 DVSS.n17836 DVSS.n15871 0.0105
R58133 DVSS.n17841 DVSS.n15871 0.0105
R58134 DVSS.n17843 DVSS.n17841 0.0105
R58135 DVSS.n17845 DVSS.n17843 0.0105
R58136 DVSS.n17845 DVSS.n15868 0.0105
R58137 DVSS.n17850 DVSS.n15868 0.0105
R58138 DVSS.n17852 DVSS.n17850 0.0105
R58139 DVSS.n17854 DVSS.n17852 0.0105
R58140 DVSS.n17854 DVSS.n15865 0.0105
R58141 DVSS.n17858 DVSS.n15865 0.0105
R58142 DVSS.n17858 DVSS.n15835 0.0105
R58143 DVSS.n17867 DVSS.n15835 0.0105
R58144 DVSS.n17867 DVSS.n15833 0.0105
R58145 DVSS.n17872 DVSS.n15833 0.0105
R58146 DVSS.n17872 DVSS.n15830 0.0105
R58147 DVSS.n17876 DVSS.n15830 0.0105
R58148 DVSS.n17878 DVSS.n17876 0.0105
R58149 DVSS.n17880 DVSS.n17878 0.0105
R58150 DVSS.n17880 DVSS.n15828 0.0105
R58151 DVSS.n17885 DVSS.n15828 0.0105
R58152 DVSS.n17887 DVSS.n17885 0.0105
R58153 DVSS.n17889 DVSS.n17887 0.0105
R58154 DVSS.n17889 DVSS.n15825 0.0105
R58155 DVSS.n17894 DVSS.n15825 0.0105
R58156 DVSS.n17896 DVSS.n17894 0.0105
R58157 DVSS.n17898 DVSS.n17896 0.0105
R58158 DVSS.n17898 DVSS.n15822 0.0105
R58159 DVSS.n17904 DVSS.n15822 0.0105
R58160 DVSS.n17904 DVSS.n17903 0.0105
R58161 DVSS.n17903 DVSS.n15784 0.0105
R58162 DVSS.n17911 DVSS.n15784 0.0105
R58163 DVSS.n17911 DVSS.n15782 0.0105
R58164 DVSS.n17916 DVSS.n15782 0.0105
R58165 DVSS.n17916 DVSS.n15780 0.0105
R58166 DVSS.n17920 DVSS.n15780 0.0105
R58167 DVSS.n17922 DVSS.n17920 0.0105
R58168 DVSS.n17922 DVSS.n15778 0.0105
R58169 DVSS.n17927 DVSS.n15778 0.0105
R58170 DVSS.n17929 DVSS.n17927 0.0105
R58171 DVSS.n17931 DVSS.n17929 0.0105
R58172 DVSS.n17931 DVSS.n15775 0.0105
R58173 DVSS.n17936 DVSS.n15775 0.0105
R58174 DVSS.n17938 DVSS.n17936 0.0105
R58175 DVSS.n17940 DVSS.n17938 0.0105
R58176 DVSS.n17940 DVSS.n15772 0.0105
R58177 DVSS.n17944 DVSS.n15772 0.0105
R58178 DVSS.n17944 DVSS.n15737 0.0105
R58179 DVSS.n17951 DVSS.n15737 0.0105
R58180 DVSS.n17951 DVSS.n15735 0.0105
R58181 DVSS.n17956 DVSS.n15735 0.0105
R58182 DVSS.n17956 DVSS.n15732 0.0105
R58183 DVSS.n17960 DVSS.n15732 0.0105
R58184 DVSS.n17962 DVSS.n17960 0.0105
R58185 DVSS.n17964 DVSS.n17962 0.0105
R58186 DVSS.n17964 DVSS.n15730 0.0105
R58187 DVSS.n17969 DVSS.n15730 0.0105
R58188 DVSS.n17971 DVSS.n17969 0.0105
R58189 DVSS.n17973 DVSS.n17971 0.0105
R58190 DVSS.n17973 DVSS.n15727 0.0105
R58191 DVSS.n18042 DVSS.n15727 0.0105
R58192 DVSS.n18042 DVSS.n18041 0.0105
R58193 DVSS.n18041 DVSS.n18039 0.0105
R58194 DVSS.n18039 DVSS.n18037 0.0105
R58195 DVSS.n18037 DVSS.n18035 0.0105
R58196 DVSS.n18035 DVSS.n18033 0.0105
R58197 DVSS.n18033 DVSS.n18032 0.0105
R58198 DVSS.n18032 DVSS.n18031 0.0105
R58199 DVSS.n18031 DVSS.n17984 0.0105
R58200 DVSS.n18027 DVSS.n17984 0.0105
R58201 DVSS.n18027 DVSS.n18026 0.0105
R58202 DVSS.n18026 DVSS.n18025 0.0105
R58203 DVSS.n18025 DVSS.n18023 0.0105
R58204 DVSS.n18023 DVSS.n18021 0.0105
R58205 DVSS.n18021 DVSS.n18019 0.0105
R58206 DVSS.n18019 DVSS.n18017 0.0105
R58207 DVSS.n18017 DVSS.n18015 0.0105
R58208 DVSS.n18015 DVSS.n18013 0.0105
R58209 DVSS.n18013 DVSS.n18011 0.0105
R58210 DVSS.n18011 DVSS.n18009 0.0105
R58211 DVSS.n18007 DVSS.n18005 0.0105
R58212 DVSS.n18005 DVSS.n18003 0.0105
R58213 DVSS.n18003 DVSS.n18002 0.0105
R58214 DVSS.n17794 DVSS.n17793 0.0105
R58215 DVSS.n17824 DVSS.n15874 0.0105
R58216 DVSS.n17831 DVSS.n15874 0.0105
R58217 DVSS.n17832 DVSS.n17831 0.0105
R58218 DVSS.n17833 DVSS.n17832 0.0105
R58219 DVSS.n17873 DVSS.n15832 0.0105
R58220 DVSS.n17874 DVSS.n17873 0.0105
R58221 DVSS.n17875 DVSS.n17874 0.0105
R58222 DVSS.n17910 DVSS.n17909 0.0105
R58223 DVSS.n17910 DVSS.n15781 0.0105
R58224 DVSS.n17917 DVSS.n15781 0.0105
R58225 DVSS.n17918 DVSS.n17917 0.0105
R58226 DVSS.n17919 DVSS.n17918 0.0105
R58227 DVSS.n17957 DVSS.n15734 0.0105
R58228 DVSS.n17958 DVSS.n17957 0.0105
R58229 DVSS.n17959 DVSS.n17958 0.0105
R58230 DVSS.n18030 DVSS.n15708 0.0105
R58231 DVSS.n18030 DVSS.n18029 0.0105
R58232 DVSS.n18029 DVSS.n18028 0.0105
R58233 DVSS.n18028 DVSS.n17985 0.0105
R58234 DVSS.n15570 DVSS.n15535 0.0105
R58235 DVSS.n16465 DVSS.n16464 0.0104
R58236 DVSS.n18083 DVSS.n15645 0.0104
R58237 DVSS.n13363 DVSS.n1505 0.0103797
R58238 DVSS.n18986 DVSS.n18985 0.0103596
R58239 DVSS.n20625 DVSS.n20624 0.0103596
R58240 DVSS.n22973 DVSS.n420 0.0103531
R58241 DVSS.n22591 DVSS.n22590 0.0103438
R58242 DVSS.n22931 DVSS.n22930 0.0103438
R58243 DVSS.n20554 DVSS.n20489 0.0103294
R58244 DVSS.n19501 DVSS.n19500 0.0102826
R58245 DVSS.n22456 DVSS.n879 0.0102826
R58246 DVSS.n19845 DVSS.n19844 0.0102826
R58247 DVSS.n22334 DVSS.n1219 0.0102826
R58248 DVSS.n22631 DVSS.n735 0.0102674
R58249 DVSS.n22890 DVSS.n22889 0.0102674
R58250 DVSS.n4009 DVSS.n3843 0.0102444
R58251 DVSS.n12343 DVSS.n12342 0.0102444
R58252 DVSS.n18708 DVSS.n18707 0.0102297
R58253 DVSS.n8108 DVSS.n8107 0.010175
R58254 DVSS.n12765 DVSS.n12764 0.010175
R58255 DVSS.n8126 DVSS.n3902 0.0101644
R58256 DVSS.n8127 DVSS.n8124 0.0101644
R58257 DVSS.n6678 DVSS.n5887 0.0101288
R58258 DVSS.n6677 DVSS.n5886 0.0101288
R58259 DVSS DVSS.n20051 0.0101067
R58260 DVSS.n18967 DVSS.n18913 0.00985393
R58261 DVSS.n20119 DVSS.n20054 0.00985393
R58262 DVSS.n20153 DVSS.n20050 0.00985393
R58263 DVSS.n20245 DVSS.n20223 0.00985393
R58264 DVSS.n20302 DVSS.n20301 0.00985393
R58265 DVSS.n20408 DVSS.n14684 0.00985393
R58266 DVSS.n3849 DVSS.n3753 0.00973581
R58267 DVSS.n3851 DVSS.n3752 0.00973581
R58268 DVSS.n7040 DVSS.n5528 0.00970301
R58269 DVSS.n7803 DVSS.n7802 0.00970301
R58270 DVSS.n10144 DVSS.n2369 0.00968121
R58271 DVSS.n10150 DVSS.n2026 0.00968121
R58272 DVSS.n10145 DVSS.n2368 0.00968121
R58273 DVSS.n10149 DVSS.n2025 0.00968121
R58274 DVSS.n22669 DVSS.n730 0.00962857
R58275 DVSS.n22669 DVSS.n732 0.00962857
R58276 DVSS.n22665 DVSS.n732 0.00962857
R58277 DVSS.n22665 DVSS.n22663 0.00962857
R58278 DVSS.n22663 DVSS.n22661 0.00962857
R58279 DVSS.n22661 DVSS.n22642 0.00962857
R58280 DVSS.n22656 DVSS.n22642 0.00962857
R58281 DVSS.n22656 DVSS.n22654 0.00962857
R58282 DVSS.n22654 DVSS.n22652 0.00962857
R58283 DVSS.n22652 DVSS.n22645 0.00962857
R58284 DVSS.n22647 DVSS.n22645 0.00962857
R58285 DVSS.n22647 DVSS.n700 0.00962857
R58286 DVSS.n22675 DVSS.n700 0.00962857
R58287 DVSS.n22675 DVSS.n698 0.00962857
R58288 DVSS.n22680 DVSS.n698 0.00962857
R58289 DVSS.n22680 DVSS.n696 0.00962857
R58290 DVSS.n22684 DVSS.n696 0.00962857
R58291 DVSS.n22686 DVSS.n22684 0.00962857
R58292 DVSS.n22686 DVSS.n694 0.00962857
R58293 DVSS.n22691 DVSS.n694 0.00962857
R58294 DVSS.n22693 DVSS.n22691 0.00962857
R58295 DVSS.n22695 DVSS.n22693 0.00962857
R58296 DVSS.n22695 DVSS.n691 0.00962857
R58297 DVSS.n22700 DVSS.n691 0.00962857
R58298 DVSS.n22702 DVSS.n22700 0.00962857
R58299 DVSS.n22704 DVSS.n22702 0.00962857
R58300 DVSS.n22704 DVSS.n688 0.00962857
R58301 DVSS.n22708 DVSS.n688 0.00962857
R58302 DVSS.n22708 DVSS.n647 0.00962857
R58303 DVSS.n22717 DVSS.n647 0.00962857
R58304 DVSS.n22717 DVSS.n645 0.00962857
R58305 DVSS.n22722 DVSS.n645 0.00962857
R58306 DVSS.n22722 DVSS.n642 0.00962857
R58307 DVSS.n22726 DVSS.n642 0.00962857
R58308 DVSS.n22728 DVSS.n22726 0.00962857
R58309 DVSS.n22730 DVSS.n22728 0.00962857
R58310 DVSS.n22730 DVSS.n640 0.00962857
R58311 DVSS.n22735 DVSS.n640 0.00962857
R58312 DVSS.n22737 DVSS.n22735 0.00962857
R58313 DVSS.n22739 DVSS.n22737 0.00962857
R58314 DVSS.n22739 DVSS.n637 0.00962857
R58315 DVSS.n22744 DVSS.n637 0.00962857
R58316 DVSS.n22746 DVSS.n22744 0.00962857
R58317 DVSS.n22748 DVSS.n22746 0.00962857
R58318 DVSS.n22748 DVSS.n633 0.00962857
R58319 DVSS.n22753 DVSS.n633 0.00962857
R58320 DVSS.n22753 DVSS.n634 0.00962857
R58321 DVSS.n634 DVSS.n595 0.00962857
R58322 DVSS.n22760 DVSS.n595 0.00962857
R58323 DVSS.n22760 DVSS.n593 0.00962857
R58324 DVSS.n22765 DVSS.n593 0.00962857
R58325 DVSS.n22765 DVSS.n591 0.00962857
R58326 DVSS.n22769 DVSS.n591 0.00962857
R58327 DVSS.n22771 DVSS.n22769 0.00962857
R58328 DVSS.n22771 DVSS.n589 0.00962857
R58329 DVSS.n22776 DVSS.n589 0.00962857
R58330 DVSS.n22778 DVSS.n22776 0.00962857
R58331 DVSS.n22780 DVSS.n22778 0.00962857
R58332 DVSS.n22780 DVSS.n586 0.00962857
R58333 DVSS.n22785 DVSS.n586 0.00962857
R58334 DVSS.n22787 DVSS.n22785 0.00962857
R58335 DVSS.n22789 DVSS.n22787 0.00962857
R58336 DVSS.n22789 DVSS.n583 0.00962857
R58337 DVSS.n22793 DVSS.n583 0.00962857
R58338 DVSS.n22793 DVSS.n546 0.00962857
R58339 DVSS.n22800 DVSS.n546 0.00962857
R58340 DVSS.n22800 DVSS.n544 0.00962857
R58341 DVSS.n22805 DVSS.n544 0.00962857
R58342 DVSS.n22805 DVSS.n541 0.00962857
R58343 DVSS.n22809 DVSS.n541 0.00962857
R58344 DVSS.n22811 DVSS.n22809 0.00962857
R58345 DVSS.n22813 DVSS.n22811 0.00962857
R58346 DVSS.n22813 DVSS.n539 0.00962857
R58347 DVSS.n22818 DVSS.n539 0.00962857
R58348 DVSS.n22820 DVSS.n22818 0.00962857
R58349 DVSS.n22822 DVSS.n22820 0.00962857
R58350 DVSS.n22822 DVSS.n536 0.00962857
R58351 DVSS.n22827 DVSS.n536 0.00962857
R58352 DVSS.n22829 DVSS.n22827 0.00962857
R58353 DVSS.n22831 DVSS.n22829 0.00962857
R58354 DVSS.n22831 DVSS.n533 0.00962857
R58355 DVSS.n22835 DVSS.n533 0.00962857
R58356 DVSS.n22835 DVSS.n495 0.00962857
R58357 DVSS.n22841 DVSS.n495 0.00962857
R58358 DVSS.n22841 DVSS.n493 0.00962857
R58359 DVSS.n22846 DVSS.n493 0.00962857
R58360 DVSS.n22846 DVSS.n491 0.00962857
R58361 DVSS.n22850 DVSS.n491 0.00962857
R58362 DVSS.n22852 DVSS.n22850 0.00962857
R58363 DVSS.n22852 DVSS.n489 0.00962857
R58364 DVSS.n22857 DVSS.n489 0.00962857
R58365 DVSS.n22859 DVSS.n22857 0.00962857
R58366 DVSS.n22861 DVSS.n22859 0.00962857
R58367 DVSS.n22861 DVSS.n486 0.00962857
R58368 DVSS.n22866 DVSS.n486 0.00962857
R58369 DVSS.n22868 DVSS.n22866 0.00962857
R58370 DVSS.n22869 DVSS.n22868 0.00962857
R58371 DVSS.n22872 DVSS.n457 0.00962857
R58372 DVSS.n22881 DVSS.n457 0.00962857
R58373 DVSS.n22881 DVSS.n455 0.00962857
R58374 DVSS.n16571 DVSS.n16569 0.00962857
R58375 DVSS.n16571 DVSS.n16566 0.00962857
R58376 DVSS.n16576 DVSS.n16566 0.00962857
R58377 DVSS.n16578 DVSS.n16576 0.00962857
R58378 DVSS.n16580 DVSS.n16578 0.00962857
R58379 DVSS.n16580 DVSS.n16563 0.00962857
R58380 DVSS.n16585 DVSS.n16563 0.00962857
R58381 DVSS.n16587 DVSS.n16585 0.00962857
R58382 DVSS.n16589 DVSS.n16587 0.00962857
R58383 DVSS.n16589 DVSS.n16560 0.00962857
R58384 DVSS.n16593 DVSS.n16560 0.00962857
R58385 DVSS.n16593 DVSS.n16333 0.00962857
R58386 DVSS.n16599 DVSS.n16333 0.00962857
R58387 DVSS.n16599 DVSS.n16331 0.00962857
R58388 DVSS.n16604 DVSS.n16331 0.00962857
R58389 DVSS.n16604 DVSS.n16329 0.00962857
R58390 DVSS.n16608 DVSS.n16329 0.00962857
R58391 DVSS.n16610 DVSS.n16608 0.00962857
R58392 DVSS.n16610 DVSS.n16327 0.00962857
R58393 DVSS.n16615 DVSS.n16327 0.00962857
R58394 DVSS.n16617 DVSS.n16615 0.00962857
R58395 DVSS.n16619 DVSS.n16617 0.00962857
R58396 DVSS.n16619 DVSS.n16324 0.00962857
R58397 DVSS.n16624 DVSS.n16324 0.00962857
R58398 DVSS.n16626 DVSS.n16624 0.00962857
R58399 DVSS.n16628 DVSS.n16626 0.00962857
R58400 DVSS.n16628 DVSS.n16321 0.00962857
R58401 DVSS.n16632 DVSS.n16321 0.00962857
R58402 DVSS.n16632 DVSS.n16291 0.00962857
R58403 DVSS.n16641 DVSS.n16291 0.00962857
R58404 DVSS.n16641 DVSS.n16289 0.00962857
R58405 DVSS.n16646 DVSS.n16289 0.00962857
R58406 DVSS.n16646 DVSS.n16286 0.00962857
R58407 DVSS.n16650 DVSS.n16286 0.00962857
R58408 DVSS.n16652 DVSS.n16650 0.00962857
R58409 DVSS.n16654 DVSS.n16652 0.00962857
R58410 DVSS.n16654 DVSS.n16284 0.00962857
R58411 DVSS.n16659 DVSS.n16284 0.00962857
R58412 DVSS.n16661 DVSS.n16659 0.00962857
R58413 DVSS.n16663 DVSS.n16661 0.00962857
R58414 DVSS.n16663 DVSS.n16281 0.00962857
R58415 DVSS.n16668 DVSS.n16281 0.00962857
R58416 DVSS.n16670 DVSS.n16668 0.00962857
R58417 DVSS.n16672 DVSS.n16670 0.00962857
R58418 DVSS.n16672 DVSS.n16277 0.00962857
R58419 DVSS.n16677 DVSS.n16277 0.00962857
R58420 DVSS.n16677 DVSS.n16278 0.00962857
R58421 DVSS.n16278 DVSS.n16240 0.00962857
R58422 DVSS.n16684 DVSS.n16240 0.00962857
R58423 DVSS.n16684 DVSS.n16238 0.00962857
R58424 DVSS.n16688 DVSS.n16238 0.00962857
R58425 DVSS.n16688 DVSS.n16236 0.00962857
R58426 DVSS.n16692 DVSS.n16236 0.00962857
R58427 DVSS.n16692 DVSS.n16234 0.00962857
R58428 DVSS.n16697 DVSS.n16234 0.00962857
R58429 DVSS.n16699 DVSS.n16697 0.00962857
R58430 DVSS.n16701 DVSS.n16699 0.00962857
R58431 DVSS.n16701 DVSS.n16231 0.00962857
R58432 DVSS.n16706 DVSS.n16231 0.00962857
R58433 DVSS.n16708 DVSS.n16706 0.00962857
R58434 DVSS.n16710 DVSS.n16708 0.00962857
R58435 DVSS.n16710 DVSS.n16226 0.00962857
R58436 DVSS.n16820 DVSS.n16226 0.00962857
R58437 DVSS.n16820 DVSS.n16228 0.00962857
R58438 DVSS.n16816 DVSS.n16228 0.00962857
R58439 DVSS.n16816 DVSS.n16814 0.00962857
R58440 DVSS.n16814 DVSS.n16813 0.00962857
R58441 DVSS.n16813 DVSS.n16714 0.00962857
R58442 DVSS.n16809 DVSS.n16714 0.00962857
R58443 DVSS.n16809 DVSS.n16805 0.00962857
R58444 DVSS.n16805 DVSS.n16804 0.00962857
R58445 DVSS.n16804 DVSS.n16717 0.00962857
R58446 DVSS.n16799 DVSS.n16717 0.00962857
R58447 DVSS.n16799 DVSS.n16797 0.00962857
R58448 DVSS.n16797 DVSS.n16795 0.00962857
R58449 DVSS.n16795 DVSS.n16720 0.00962857
R58450 DVSS.n16790 DVSS.n16720 0.00962857
R58451 DVSS.n16790 DVSS.n16788 0.00962857
R58452 DVSS.n16788 DVSS.n16786 0.00962857
R58453 DVSS.n16786 DVSS.n16723 0.00962857
R58454 DVSS.n16781 DVSS.n16723 0.00962857
R58455 DVSS.n16781 DVSS.n16779 0.00962857
R58456 DVSS.n16779 DVSS.n16777 0.00962857
R58457 DVSS.n16777 DVSS.n16725 0.00962857
R58458 DVSS.n16773 DVSS.n16725 0.00962857
R58459 DVSS.n16773 DVSS.n16727 0.00962857
R58460 DVSS.n16769 DVSS.n16727 0.00962857
R58461 DVSS.n16769 DVSS.n16729 0.00962857
R58462 DVSS.n16765 DVSS.n16729 0.00962857
R58463 DVSS.n16765 DVSS.n16763 0.00962857
R58464 DVSS.n16763 DVSS.n16761 0.00962857
R58465 DVSS.n16761 DVSS.n16732 0.00962857
R58466 DVSS.n16756 DVSS.n16732 0.00962857
R58467 DVSS.n16756 DVSS.n16754 0.00962857
R58468 DVSS.n16754 DVSS.n16752 0.00962857
R58469 DVSS.n16752 DVSS.n16735 0.00962857
R58470 DVSS.n16747 DVSS.n16735 0.00962857
R58471 DVSS.n16745 DVSS.n16743 0.00962857
R58472 DVSS.n16743 DVSS.n16737 0.00962857
R58473 DVSS.n16738 DVSS.n16737 0.00962857
R58474 DVSS.n16568 DVSS.n15919 0.00962857
R58475 DVSS.n16598 DVSS.n16330 0.00962857
R58476 DVSS.n16605 DVSS.n16330 0.00962857
R58477 DVSS.n16606 DVSS.n16605 0.00962857
R58478 DVSS.n16607 DVSS.n16606 0.00962857
R58479 DVSS.n16647 DVSS.n16288 0.00962857
R58480 DVSS.n16648 DVSS.n16647 0.00962857
R58481 DVSS.n16649 DVSS.n16648 0.00962857
R58482 DVSS.n16683 DVSS.n16682 0.00962857
R58483 DVSS.n16683 DVSS.n16237 0.00962857
R58484 DVSS.n16689 DVSS.n16237 0.00962857
R58485 DVSS.n16690 DVSS.n16689 0.00962857
R58486 DVSS.n16691 DVSS.n16690 0.00962857
R58487 DVSS.n16806 DVSS.n16171 0.00962857
R58488 DVSS.n16808 DVSS.n16806 0.00962857
R58489 DVSS.n16808 DVSS.n16807 0.00962857
R58490 DVSS.n16772 DVSS.n15673 0.00962857
R58491 DVSS.n16772 DVSS.n16771 0.00962857
R58492 DVSS.n16771 DVSS.n16770 0.00962857
R58493 DVSS.n16770 DVSS.n16728 0.00962857
R58494 DVSS.n15613 DVSS.n15534 0.00962857
R58495 DVSS.n17781 DVSS.n15923 0.00962857
R58496 DVSS.n17781 DVSS.n15925 0.00962857
R58497 DVSS.n15971 DVSS.n15925 0.00962857
R58498 DVSS.n15973 DVSS.n15971 0.00962857
R58499 DVSS.n15973 DVSS.n15968 0.00962857
R58500 DVSS.n15978 DVSS.n15968 0.00962857
R58501 DVSS.n15980 DVSS.n15978 0.00962857
R58502 DVSS.n15982 DVSS.n15980 0.00962857
R58503 DVSS.n15982 DVSS.n15963 0.00962857
R58504 DVSS.n17671 DVSS.n15963 0.00962857
R58505 DVSS.n17671 DVSS.n15965 0.00962857
R58506 DVSS.n17667 DVSS.n15965 0.00962857
R58507 DVSS.n17667 DVSS.n17666 0.00962857
R58508 DVSS.n17666 DVSS.n17665 0.00962857
R58509 DVSS.n17665 DVSS.n15986 0.00962857
R58510 DVSS.n17661 DVSS.n15986 0.00962857
R58511 DVSS.n17661 DVSS.n15989 0.00962857
R58512 DVSS.n17657 DVSS.n15989 0.00962857
R58513 DVSS.n17657 DVSS.n15992 0.00962857
R58514 DVSS.n16042 DVSS.n15992 0.00962857
R58515 DVSS.n16044 DVSS.n16042 0.00962857
R58516 DVSS.n16044 DVSS.n16039 0.00962857
R58517 DVSS.n16049 DVSS.n16039 0.00962857
R58518 DVSS.n16051 DVSS.n16049 0.00962857
R58519 DVSS.n16053 DVSS.n16051 0.00962857
R58520 DVSS.n16053 DVSS.n16036 0.00962857
R58521 DVSS.n16058 DVSS.n16036 0.00962857
R58522 DVSS.n16060 DVSS.n16058 0.00962857
R58523 DVSS.n16062 DVSS.n16060 0.00962857
R58524 DVSS.n16062 DVSS.n16032 0.00962857
R58525 DVSS.n17651 DVSS.n16032 0.00962857
R58526 DVSS.n17651 DVSS.n16033 0.00962857
R58527 DVSS.n17647 DVSS.n16033 0.00962857
R58528 DVSS.n17647 DVSS.n16066 0.00962857
R58529 DVSS.n16112 DVSS.n16066 0.00962857
R58530 DVSS.n16116 DVSS.n16112 0.00962857
R58531 DVSS.n16118 DVSS.n16116 0.00962857
R58532 DVSS.n16120 DVSS.n16118 0.00962857
R58533 DVSS.n16120 DVSS.n16110 0.00962857
R58534 DVSS.n16125 DVSS.n16110 0.00962857
R58535 DVSS.n16127 DVSS.n16125 0.00962857
R58536 DVSS.n16129 DVSS.n16127 0.00962857
R58537 DVSS.n16129 DVSS.n16105 0.00962857
R58538 DVSS.n17638 DVSS.n16105 0.00962857
R58539 DVSS.n17638 DVSS.n16107 0.00962857
R58540 DVSS.n17634 DVSS.n16107 0.00962857
R58541 DVSS.n17634 DVSS.n17632 0.00962857
R58542 DVSS.n17632 DVSS.n17631 0.00962857
R58543 DVSS.n17631 DVSS.n16133 0.00962857
R58544 DVSS.n17627 DVSS.n16133 0.00962857
R58545 DVSS.n17627 DVSS.n16135 0.00962857
R58546 DVSS.n17623 DVSS.n16135 0.00962857
R58547 DVSS.n17623 DVSS.n16138 0.00962857
R58548 DVSS.n17619 DVSS.n16138 0.00962857
R58549 DVSS.n17619 DVSS.n16140 0.00962857
R58550 DVSS.n16864 DVSS.n16140 0.00962857
R58551 DVSS.n16866 DVSS.n16864 0.00962857
R58552 DVSS.n16866 DVSS.n16861 0.00962857
R58553 DVSS.n16871 DVSS.n16861 0.00962857
R58554 DVSS.n16873 DVSS.n16871 0.00962857
R58555 DVSS.n16875 DVSS.n16873 0.00962857
R58556 DVSS.n16875 DVSS.n16858 0.00962857
R58557 DVSS.n16880 DVSS.n16858 0.00962857
R58558 DVSS.n16882 DVSS.n16880 0.00962857
R58559 DVSS.n16884 DVSS.n16882 0.00962857
R58560 DVSS.n16884 DVSS.n16854 0.00962857
R58561 DVSS.n17613 DVSS.n16854 0.00962857
R58562 DVSS.n17613 DVSS.n16855 0.00962857
R58563 DVSS.n17609 DVSS.n16855 0.00962857
R58564 DVSS.n17609 DVSS.n16888 0.00962857
R58565 DVSS.n17547 DVSS.n16888 0.00962857
R58566 DVSS.n17602 DVSS.n17547 0.00962857
R58567 DVSS.n17602 DVSS.n17549 0.00962857
R58568 DVSS.n17598 DVSS.n17549 0.00962857
R58569 DVSS.n17598 DVSS.n17596 0.00962857
R58570 DVSS.n17596 DVSS.n17594 0.00962857
R58571 DVSS.n17594 DVSS.n17553 0.00962857
R58572 DVSS.n17589 DVSS.n17553 0.00962857
R58573 DVSS.n17589 DVSS.n17587 0.00962857
R58574 DVSS.n17587 DVSS.n17585 0.00962857
R58575 DVSS.n17585 DVSS.n17556 0.00962857
R58576 DVSS.n17580 DVSS.n17556 0.00962857
R58577 DVSS.n17580 DVSS.n17578 0.00962857
R58578 DVSS.n17578 DVSS.n17576 0.00962857
R58579 DVSS.n17576 DVSS.n17558 0.00962857
R58580 DVSS.n17572 DVSS.n17558 0.00962857
R58581 DVSS.n17572 DVSS.n17561 0.00962857
R58582 DVSS.n17568 DVSS.n17561 0.00962857
R58583 DVSS.n17568 DVSS.n17567 0.00962857
R58584 DVSS.n17567 DVSS.n17566 0.00962857
R58585 DVSS.n17566 DVSS.n15523 0.00962857
R58586 DVSS.n18196 DVSS.n15523 0.00962857
R58587 DVSS.n18196 DVSS.n15525 0.00962857
R58588 DVSS.n18192 DVSS.n15525 0.00962857
R58589 DVSS.n18192 DVSS.n18190 0.00962857
R58590 DVSS.n18190 DVSS.n18188 0.00962857
R58591 DVSS.n18188 DVSS.n15529 0.00962857
R58592 DVSS.n18183 DVSS.n18181 0.00962857
R58593 DVSS.n18181 DVSS.n15531 0.00962857
R58594 DVSS.n18176 DVSS.n15531 0.00962857
R58595 DVSS.n17784 DVSS.n15922 0.00962857
R58596 DVSS.n17664 DVSS.n15956 0.00962857
R58597 DVSS.n17664 DVSS.n17663 0.00962857
R58598 DVSS.n17663 DVSS.n17662 0.00962857
R58599 DVSS.n17662 DVSS.n15988 0.00962857
R58600 DVSS.n17652 DVSS.n16031 0.00962857
R58601 DVSS.n17646 DVSS.n16031 0.00962857
R58602 DVSS.n17646 DVSS.n17645 0.00962857
R58603 DVSS.n16136 DVSS.n16093 0.00962857
R58604 DVSS.n17626 DVSS.n16136 0.00962857
R58605 DVSS.n17626 DVSS.n17625 0.00962857
R58606 DVSS.n17625 DVSS.n17624 0.00962857
R58607 DVSS.n17624 DVSS.n16137 0.00962857
R58608 DVSS.n17614 DVSS.n16853 0.00962857
R58609 DVSS.n17608 DVSS.n16853 0.00962857
R58610 DVSS.n17608 DVSS.n17607 0.00962857
R58611 DVSS.n17575 DVSS.n17574 0.00962857
R58612 DVSS.n17574 DVSS.n17573 0.00962857
R58613 DVSS.n17573 DVSS.n17560 0.00962857
R58614 DVSS.n17560 DVSS.n15505 0.00962857
R58615 DVSS.n18175 DVSS.n18174 0.00962857
R58616 DVSS.n17721 DVSS.n17718 0.00962857
R58617 DVSS.n17726 DVSS.n17718 0.00962857
R58618 DVSS.n17728 DVSS.n17726 0.00962857
R58619 DVSS.n17730 DVSS.n17728 0.00962857
R58620 DVSS.n17730 DVSS.n17715 0.00962857
R58621 DVSS.n17735 DVSS.n17715 0.00962857
R58622 DVSS.n17737 DVSS.n17735 0.00962857
R58623 DVSS.n17739 DVSS.n17737 0.00962857
R58624 DVSS.n17739 DVSS.n17710 0.00962857
R58625 DVSS.n17769 DVSS.n17710 0.00962857
R58626 DVSS.n17769 DVSS.n17712 0.00962857
R58627 DVSS.n17765 DVSS.n17712 0.00962857
R58628 DVSS.n17765 DVSS.n17764 0.00962857
R58629 DVSS.n17764 DVSS.n17763 0.00962857
R58630 DVSS.n17763 DVSS.n17743 0.00962857
R58631 DVSS.n17759 DVSS.n17743 0.00962857
R58632 DVSS.n17759 DVSS.n17746 0.00962857
R58633 DVSS.n17755 DVSS.n17746 0.00962857
R58634 DVSS.n17755 DVSS.n17753 0.00962857
R58635 DVSS.n17753 DVSS.n17751 0.00962857
R58636 DVSS.n17751 DVSS.n15275 0.00962857
R58637 DVSS.n18376 DVSS.n15275 0.00962857
R58638 DVSS.n18376 DVSS.n15277 0.00962857
R58639 DVSS.n18372 DVSS.n15277 0.00962857
R58640 DVSS.n18372 DVSS.n18370 0.00962857
R58641 DVSS.n18370 DVSS.n18368 0.00962857
R58642 DVSS.n18368 DVSS.n15281 0.00962857
R58643 DVSS.n18363 DVSS.n15281 0.00962857
R58644 DVSS.n18363 DVSS.n18361 0.00962857
R58645 DVSS.n18361 DVSS.n18359 0.00962857
R58646 DVSS.n18359 DVSS.n15283 0.00962857
R58647 DVSS.n18355 DVSS.n15283 0.00962857
R58648 DVSS.n18355 DVSS.n15285 0.00962857
R58649 DVSS.n18351 DVSS.n15285 0.00962857
R58650 DVSS.n18351 DVSS.n15287 0.00962857
R58651 DVSS.n18347 DVSS.n15287 0.00962857
R58652 DVSS.n18347 DVSS.n15289 0.00962857
R58653 DVSS.n15335 DVSS.n15289 0.00962857
R58654 DVSS.n15335 DVSS.n15333 0.00962857
R58655 DVSS.n15340 DVSS.n15333 0.00962857
R58656 DVSS.n15342 DVSS.n15340 0.00962857
R58657 DVSS.n15344 DVSS.n15342 0.00962857
R58658 DVSS.n15344 DVSS.n15330 0.00962857
R58659 DVSS.n15349 DVSS.n15330 0.00962857
R58660 DVSS.n15351 DVSS.n15349 0.00962857
R58661 DVSS.n15353 DVSS.n15351 0.00962857
R58662 DVSS.n15353 DVSS.n15326 0.00962857
R58663 DVSS.n18341 DVSS.n15326 0.00962857
R58664 DVSS.n18341 DVSS.n15327 0.00962857
R58665 DVSS.n18337 DVSS.n15327 0.00962857
R58666 DVSS.n18337 DVSS.n15357 0.00962857
R58667 DVSS.n18333 DVSS.n15357 0.00962857
R58668 DVSS.n18333 DVSS.n15359 0.00962857
R58669 DVSS.n18329 DVSS.n15359 0.00962857
R58670 DVSS.n18329 DVSS.n15361 0.00962857
R58671 DVSS.n15408 DVSS.n15361 0.00962857
R58672 DVSS.n15410 DVSS.n15408 0.00962857
R58673 DVSS.n15410 DVSS.n15405 0.00962857
R58674 DVSS.n15415 DVSS.n15405 0.00962857
R58675 DVSS.n15417 DVSS.n15415 0.00962857
R58676 DVSS.n15419 DVSS.n15417 0.00962857
R58677 DVSS.n15419 DVSS.n15402 0.00962857
R58678 DVSS.n15424 DVSS.n15402 0.00962857
R58679 DVSS.n15426 DVSS.n15424 0.00962857
R58680 DVSS.n15428 DVSS.n15426 0.00962857
R58681 DVSS.n15428 DVSS.n15398 0.00962857
R58682 DVSS.n18323 DVSS.n15398 0.00962857
R58683 DVSS.n18323 DVSS.n15399 0.00962857
R58684 DVSS.n18319 DVSS.n15399 0.00962857
R58685 DVSS.n18319 DVSS.n15432 0.00962857
R58686 DVSS.n15467 DVSS.n15432 0.00962857
R58687 DVSS.n18312 DVSS.n15467 0.00962857
R58688 DVSS.n18312 DVSS.n15469 0.00962857
R58689 DVSS.n18308 DVSS.n15469 0.00962857
R58690 DVSS.n18308 DVSS.n18306 0.00962857
R58691 DVSS.n18306 DVSS.n18304 0.00962857
R58692 DVSS.n18304 DVSS.n15473 0.00962857
R58693 DVSS.n18299 DVSS.n15473 0.00962857
R58694 DVSS.n18299 DVSS.n18297 0.00962857
R58695 DVSS.n18297 DVSS.n18295 0.00962857
R58696 DVSS.n18295 DVSS.n15476 0.00962857
R58697 DVSS.n18290 DVSS.n15476 0.00962857
R58698 DVSS.n18290 DVSS.n18288 0.00962857
R58699 DVSS.n18288 DVSS.n18286 0.00962857
R58700 DVSS.n18286 DVSS.n15478 0.00962857
R58701 DVSS.n18282 DVSS.n15478 0.00962857
R58702 DVSS.n18282 DVSS.n15481 0.00962857
R58703 DVSS.n18278 DVSS.n15481 0.00962857
R58704 DVSS.n18278 DVSS.n15484 0.00962857
R58705 DVSS.n18238 DVSS.n15484 0.00962857
R58706 DVSS.n18272 DVSS.n18238 0.00962857
R58707 DVSS.n18272 DVSS.n18240 0.00962857
R58708 DVSS.n18268 DVSS.n18240 0.00962857
R58709 DVSS.n18268 DVSS.n18266 0.00962857
R58710 DVSS.n18266 DVSS.n18264 0.00962857
R58711 DVSS.n18264 DVSS.n18244 0.00962857
R58712 DVSS.n18259 DVSS.n18244 0.00962857
R58713 DVSS.n18257 DVSS.n18255 0.00962857
R58714 DVSS.n18255 DVSS.n18247 0.00962857
R58715 DVSS.n18250 DVSS.n18247 0.00962857
R58716 DVSS.n17720 DVSS.n17719 0.00962857
R58717 DVSS.n17762 DVSS.n17698 0.00962857
R58718 DVSS.n17762 DVSS.n17761 0.00962857
R58719 DVSS.n17761 DVSS.n17760 0.00962857
R58720 DVSS.n17760 DVSS.n17745 0.00962857
R58721 DVSS.n18354 DVSS.n15259 0.00962857
R58722 DVSS.n18354 DVSS.n18353 0.00962857
R58723 DVSS.n18353 DVSS.n18352 0.00962857
R58724 DVSS.n18342 DVSS.n15325 0.00962857
R58725 DVSS.n18336 DVSS.n15325 0.00962857
R58726 DVSS.n18336 DVSS.n18335 0.00962857
R58727 DVSS.n18335 DVSS.n18334 0.00962857
R58728 DVSS.n18334 DVSS.n15358 0.00962857
R58729 DVSS.n18324 DVSS.n15397 0.00962857
R58730 DVSS.n18318 DVSS.n15397 0.00962857
R58731 DVSS.n18318 DVSS.n18317 0.00962857
R58732 DVSS.n18285 DVSS.n18284 0.00962857
R58733 DVSS.n18284 DVSS.n18283 0.00962857
R58734 DVSS.n18283 DVSS.n15480 0.00962857
R58735 DVSS.n18277 DVSS.n15480 0.00962857
R58736 DVSS.n18249 DVSS.n18248 0.00962857
R58737 DVSS.n18494 DVSS.n15150 0.00962857
R58738 DVSS.n18494 DVSS.n15152 0.00962857
R58739 DVSS.n15195 DVSS.n15152 0.00962857
R58740 DVSS.n15195 DVSS.n15193 0.00962857
R58741 DVSS.n15200 DVSS.n15193 0.00962857
R58742 DVSS.n15202 DVSS.n15200 0.00962857
R58743 DVSS.n15204 DVSS.n15202 0.00962857
R58744 DVSS.n15204 DVSS.n15190 0.00962857
R58745 DVSS.n15208 DVSS.n15190 0.00962857
R58746 DVSS.n15216 DVSS.n15208 0.00962857
R58747 DVSS.n15218 DVSS.n15216 0.00962857
R58748 DVSS.n15218 DVSS.n15186 0.00962857
R58749 DVSS.n18488 DVSS.n15186 0.00962857
R58750 DVSS.n18488 DVSS.n15187 0.00962857
R58751 DVSS.n18484 DVSS.n15187 0.00962857
R58752 DVSS.n18484 DVSS.n15222 0.00962857
R58753 DVSS.n18480 DVSS.n15222 0.00962857
R58754 DVSS.n18480 DVSS.n15224 0.00962857
R58755 DVSS.n18476 DVSS.n15224 0.00962857
R58756 DVSS.n18476 DVSS.n15226 0.00962857
R58757 DVSS.n18411 DVSS.n15226 0.00962857
R58758 DVSS.n18411 DVSS.n18409 0.00962857
R58759 DVSS.n18416 DVSS.n18409 0.00962857
R58760 DVSS.n18418 DVSS.n18416 0.00962857
R58761 DVSS.n18420 DVSS.n18418 0.00962857
R58762 DVSS.n18420 DVSS.n18406 0.00962857
R58763 DVSS.n18425 DVSS.n18406 0.00962857
R58764 DVSS.n18426 DVSS.n18425 0.00962857
R58765 DVSS.n18435 DVSS.n18426 0.00962857
R58766 DVSS.n18435 DVSS.n18402 0.00962857
R58767 DVSS.n18470 DVSS.n18402 0.00962857
R58768 DVSS.n18470 DVSS.n18403 0.00962857
R58769 DVSS.n18466 DVSS.n18403 0.00962857
R58770 DVSS.n18466 DVSS.n18463 0.00962857
R58771 DVSS.n18463 DVSS.n18462 0.00962857
R58772 DVSS.n18462 DVSS.n18440 0.00962857
R58773 DVSS.n18457 DVSS.n18440 0.00962857
R58774 DVSS.n18457 DVSS.n18455 0.00962857
R58775 DVSS.n18455 DVSS.n18453 0.00962857
R58776 DVSS.n18453 DVSS.n18443 0.00962857
R58777 DVSS.n18448 DVSS.n18443 0.00962857
R58778 DVSS.n18448 DVSS.n18446 0.00962857
R58779 DVSS.n18446 DVSS.n14914 0.00962857
R58780 DVSS.n20004 DVSS.n14914 0.00962857
R58781 DVSS.n20004 DVSS.n14916 0.00962857
R58782 DVSS.n20000 DVSS.n14916 0.00962857
R58783 DVSS.n20000 DVSS.n19998 0.00962857
R58784 DVSS.n19998 DVSS.n19997 0.00962857
R58785 DVSS.n19997 DVSS.n14919 0.00962857
R58786 DVSS.n19993 DVSS.n14919 0.00962857
R58787 DVSS.n19993 DVSS.n14921 0.00962857
R58788 DVSS.n19989 DVSS.n14921 0.00962857
R58789 DVSS.n19989 DVSS.n14924 0.00962857
R58790 DVSS.n19985 DVSS.n14924 0.00962857
R58791 DVSS.n19985 DVSS.n14926 0.00962857
R58792 DVSS.n14970 DVSS.n14926 0.00962857
R58793 DVSS.n14972 DVSS.n14970 0.00962857
R58794 DVSS.n14972 DVSS.n14967 0.00962857
R58795 DVSS.n14977 DVSS.n14967 0.00962857
R58796 DVSS.n14979 DVSS.n14977 0.00962857
R58797 DVSS.n14981 DVSS.n14979 0.00962857
R58798 DVSS.n14981 DVSS.n14964 0.00962857
R58799 DVSS.n14986 DVSS.n14964 0.00962857
R58800 DVSS.n14994 DVSS.n14986 0.00962857
R58801 DVSS.n14996 DVSS.n14994 0.00962857
R58802 DVSS.n14996 DVSS.n14960 0.00962857
R58803 DVSS.n19979 DVSS.n14960 0.00962857
R58804 DVSS.n19979 DVSS.n14961 0.00962857
R58805 DVSS.n19975 DVSS.n14961 0.00962857
R58806 DVSS.n19975 DVSS.n15000 0.00962857
R58807 DVSS.n15044 DVSS.n15000 0.00962857
R58808 DVSS.n15048 DVSS.n15044 0.00962857
R58809 DVSS.n15050 DVSS.n15048 0.00962857
R58810 DVSS.n15052 DVSS.n15050 0.00962857
R58811 DVSS.n15052 DVSS.n15042 0.00962857
R58812 DVSS.n15057 DVSS.n15042 0.00962857
R58813 DVSS.n15059 DVSS.n15057 0.00962857
R58814 DVSS.n15061 DVSS.n15059 0.00962857
R58815 DVSS.n15061 DVSS.n15039 0.00962857
R58816 DVSS.n15065 DVSS.n15039 0.00962857
R58817 DVSS.n15073 DVSS.n15065 0.00962857
R58818 DVSS.n15075 DVSS.n15073 0.00962857
R58819 DVSS.n15075 DVSS.n15035 0.00962857
R58820 DVSS.n19968 DVSS.n15035 0.00962857
R58821 DVSS.n19968 DVSS.n15036 0.00962857
R58822 DVSS.n19964 DVSS.n15036 0.00962857
R58823 DVSS.n19964 DVSS.n15079 0.00962857
R58824 DVSS.n19960 DVSS.n15079 0.00962857
R58825 DVSS.n19960 DVSS.n15081 0.00962857
R58826 DVSS.n19956 DVSS.n15081 0.00962857
R58827 DVSS.n19956 DVSS.n15083 0.00962857
R58828 DVSS.n19949 DVSS.n15083 0.00962857
R58829 DVSS.n19949 DVSS.n15120 0.00962857
R58830 DVSS.n19945 DVSS.n15120 0.00962857
R58831 DVSS.n19945 DVSS.n19943 0.00962857
R58832 DVSS.n19943 DVSS.n19941 0.00962857
R58833 DVSS.n19941 DVSS.n15123 0.00962857
R58834 DVSS.n19936 DVSS.n19934 0.00962857
R58835 DVSS.n19934 DVSS.n15125 0.00962857
R58836 DVSS.n19929 DVSS.n15125 0.00962857
R58837 DVSS.n18497 DVSS.n15149 0.00962857
R58838 DVSS.n18489 DVSS.n15185 0.00962857
R58839 DVSS.n18483 DVSS.n15185 0.00962857
R58840 DVSS.n18483 DVSS.n18482 0.00962857
R58841 DVSS.n18482 DVSS.n18481 0.00962857
R58842 DVSS.n18471 DVSS.n18401 0.00962857
R58843 DVSS.n18465 DVSS.n18401 0.00962857
R58844 DVSS.n18465 DVSS.n18464 0.00962857
R58845 DVSS.n14922 DVSS.n14894 0.00962857
R58846 DVSS.n19992 DVSS.n14922 0.00962857
R58847 DVSS.n19992 DVSS.n19991 0.00962857
R58848 DVSS.n19991 DVSS.n19990 0.00962857
R58849 DVSS.n19990 DVSS.n14923 0.00962857
R58850 DVSS.n19980 DVSS.n14959 0.00962857
R58851 DVSS.n19974 DVSS.n14959 0.00962857
R58852 DVSS.n19974 DVSS.n19973 0.00962857
R58853 DVSS.n19969 DVSS.n15034 0.00962857
R58854 DVSS.n19963 DVSS.n15034 0.00962857
R58855 DVSS.n19963 DVSS.n19962 0.00962857
R58856 DVSS.n19962 DVSS.n19961 0.00962857
R58857 DVSS.n19928 DVSS.n19927 0.00962857
R58858 DVSS.n21149 DVSS.n13688 0.00962857
R58859 DVSS.n21149 DVSS.n13690 0.00962857
R58860 DVSS.n20745 DVSS.n13690 0.00962857
R58861 DVSS.n20747 DVSS.n20745 0.00962857
R58862 DVSS.n20749 DVSS.n20747 0.00962857
R58863 DVSS.n20749 DVSS.n20741 0.00962857
R58864 DVSS.n20754 DVSS.n20741 0.00962857
R58865 DVSS.n20756 DVSS.n20754 0.00962857
R58866 DVSS.n20758 DVSS.n20756 0.00962857
R58867 DVSS.n20758 DVSS.n20738 0.00962857
R58868 DVSS.n20763 DVSS.n20738 0.00962857
R58869 DVSS.n20764 DVSS.n20763 0.00962857
R58870 DVSS.n20765 DVSS.n20764 0.00962857
R58871 DVSS.n20765 DVSS.n20735 0.00962857
R58872 DVSS.n20770 DVSS.n20735 0.00962857
R58873 DVSS.n20770 DVSS.n20732 0.00962857
R58874 DVSS.n20774 DVSS.n20732 0.00962857
R58875 DVSS.n20776 DVSS.n20774 0.00962857
R58876 DVSS.n20778 DVSS.n20776 0.00962857
R58877 DVSS.n20778 DVSS.n20730 0.00962857
R58878 DVSS.n20783 DVSS.n20730 0.00962857
R58879 DVSS.n20785 DVSS.n20783 0.00962857
R58880 DVSS.n20787 DVSS.n20785 0.00962857
R58881 DVSS.n20787 DVSS.n20727 0.00962857
R58882 DVSS.n20792 DVSS.n20727 0.00962857
R58883 DVSS.n20794 DVSS.n20792 0.00962857
R58884 DVSS.n20796 DVSS.n20794 0.00962857
R58885 DVSS.n20796 DVSS.n20724 0.00962857
R58886 DVSS.n20800 DVSS.n20724 0.00962857
R58887 DVSS.n20800 DVSS.n14505 0.00962857
R58888 DVSS.n20807 DVSS.n14505 0.00962857
R58889 DVSS.n20807 DVSS.n14503 0.00962857
R58890 DVSS.n20812 DVSS.n14503 0.00962857
R58891 DVSS.n20812 DVSS.n14501 0.00962857
R58892 DVSS.n20820 DVSS.n14501 0.00962857
R58893 DVSS.n20822 DVSS.n20820 0.00962857
R58894 DVSS.n20822 DVSS.n14499 0.00962857
R58895 DVSS.n20827 DVSS.n14499 0.00962857
R58896 DVSS.n20829 DVSS.n20827 0.00962857
R58897 DVSS.n20831 DVSS.n20829 0.00962857
R58898 DVSS.n20831 DVSS.n14496 0.00962857
R58899 DVSS.n20836 DVSS.n14496 0.00962857
R58900 DVSS.n20838 DVSS.n20836 0.00962857
R58901 DVSS.n20840 DVSS.n20838 0.00962857
R58902 DVSS.n20840 DVSS.n14492 0.00962857
R58903 DVSS.n20845 DVSS.n14492 0.00962857
R58904 DVSS.n20845 DVSS.n14493 0.00962857
R58905 DVSS.n14493 DVSS.n14458 0.00962857
R58906 DVSS.n20852 DVSS.n14458 0.00962857
R58907 DVSS.n20852 DVSS.n14456 0.00962857
R58908 DVSS.n20857 DVSS.n14456 0.00962857
R58909 DVSS.n20857 DVSS.n14454 0.00962857
R58910 DVSS.n20861 DVSS.n14454 0.00962857
R58911 DVSS.n20863 DVSS.n20861 0.00962857
R58912 DVSS.n20863 DVSS.n14452 0.00962857
R58913 DVSS.n20868 DVSS.n14452 0.00962857
R58914 DVSS.n20870 DVSS.n20868 0.00962857
R58915 DVSS.n20872 DVSS.n20870 0.00962857
R58916 DVSS.n20872 DVSS.n14449 0.00962857
R58917 DVSS.n20877 DVSS.n14449 0.00962857
R58918 DVSS.n20879 DVSS.n20877 0.00962857
R58919 DVSS.n20881 DVSS.n20879 0.00962857
R58920 DVSS.n20881 DVSS.n14446 0.00962857
R58921 DVSS.n20885 DVSS.n14446 0.00962857
R58922 DVSS.n20885 DVSS.n14409 0.00962857
R58923 DVSS.n20892 DVSS.n14409 0.00962857
R58924 DVSS.n20892 DVSS.n14407 0.00962857
R58925 DVSS.n20897 DVSS.n14407 0.00962857
R58926 DVSS.n20897 DVSS.n14405 0.00962857
R58927 DVSS.n20901 DVSS.n14405 0.00962857
R58928 DVSS.n20903 DVSS.n20901 0.00962857
R58929 DVSS.n20903 DVSS.n14403 0.00962857
R58930 DVSS.n20908 DVSS.n14403 0.00962857
R58931 DVSS.n20910 DVSS.n20908 0.00962857
R58932 DVSS.n20912 DVSS.n20910 0.00962857
R58933 DVSS.n20912 DVSS.n14400 0.00962857
R58934 DVSS.n20917 DVSS.n14400 0.00962857
R58935 DVSS.n20919 DVSS.n20917 0.00962857
R58936 DVSS.n20921 DVSS.n20919 0.00962857
R58937 DVSS.n20921 DVSS.n14397 0.00962857
R58938 DVSS.n20925 DVSS.n14397 0.00962857
R58939 DVSS.n20925 DVSS.n14360 0.00962857
R58940 DVSS.n20932 DVSS.n14360 0.00962857
R58941 DVSS.n20932 DVSS.n14358 0.00962857
R58942 DVSS.n20936 DVSS.n14358 0.00962857
R58943 DVSS.n20936 DVSS.n14356 0.00962857
R58944 DVSS.n20940 DVSS.n14356 0.00962857
R58945 DVSS.n20940 DVSS.n14352 0.00962857
R58946 DVSS.n20974 DVSS.n14352 0.00962857
R58947 DVSS.n20974 DVSS.n14354 0.00962857
R58948 DVSS.n20970 DVSS.n14354 0.00962857
R58949 DVSS.n20970 DVSS.n20962 0.00962857
R58950 DVSS.n20962 DVSS.n20961 0.00962857
R58951 DVSS.n20961 DVSS.n20945 0.00962857
R58952 DVSS.n20956 DVSS.n20945 0.00962857
R58953 DVSS.n20956 DVSS.n20954 0.00962857
R58954 DVSS.n20954 DVSS.n20952 0.00962857
R58955 DVSS.n20948 DVSS.n14319 0.00962857
R58956 DVSS.n20980 DVSS.n14319 0.00962857
R58957 DVSS.n20980 DVSS.n14317 0.00962857
R58958 DVSS.n21152 DVSS.n13687 0.00962857
R58959 DVSS.n20734 DVSS.n13721 0.00962857
R58960 DVSS.n20771 DVSS.n20734 0.00962857
R58961 DVSS.n20772 DVSS.n20771 0.00962857
R58962 DVSS.n20773 DVSS.n20772 0.00962857
R58963 DVSS.n20806 DVSS.n14502 0.00962857
R58964 DVSS.n20813 DVSS.n14502 0.00962857
R58965 DVSS.n20814 DVSS.n20813 0.00962857
R58966 DVSS.n20851 DVSS.n20850 0.00962857
R58967 DVSS.n20851 DVSS.n14455 0.00962857
R58968 DVSS.n20858 DVSS.n14455 0.00962857
R58969 DVSS.n20859 DVSS.n20858 0.00962857
R58970 DVSS.n20860 DVSS.n20859 0.00962857
R58971 DVSS.n20898 DVSS.n14406 0.00962857
R58972 DVSS.n20899 DVSS.n20898 0.00962857
R58973 DVSS.n20900 DVSS.n20899 0.00962857
R58974 DVSS.n20937 DVSS.n14357 0.00962857
R58975 DVSS.n20938 DVSS.n20937 0.00962857
R58976 DVSS.n20939 DVSS.n20938 0.00962857
R58977 DVSS.n20939 DVSS.n14351 0.00962857
R58978 DVSS.n20983 DVSS.n14316 0.00962857
R58979 DVSS.n21184 DVSS.n21182 0.00962857
R58980 DVSS.n21184 DVSS.n13657 0.00962857
R58981 DVSS.n21189 DVSS.n13657 0.00962857
R58982 DVSS.n21191 DVSS.n21189 0.00962857
R58983 DVSS.n21193 DVSS.n21191 0.00962857
R58984 DVSS.n21193 DVSS.n13654 0.00962857
R58985 DVSS.n21198 DVSS.n13654 0.00962857
R58986 DVSS.n21200 DVSS.n21198 0.00962857
R58987 DVSS.n21207 DVSS.n21200 0.00962857
R58988 DVSS.n21207 DVSS.n13651 0.00962857
R58989 DVSS.n21211 DVSS.n13651 0.00962857
R58990 DVSS.n21211 DVSS.n13617 0.00962857
R58991 DVSS.n21217 DVSS.n13617 0.00962857
R58992 DVSS.n21217 DVSS.n13615 0.00962857
R58993 DVSS.n21222 DVSS.n13615 0.00962857
R58994 DVSS.n21222 DVSS.n13613 0.00962857
R58995 DVSS.n21226 DVSS.n13613 0.00962857
R58996 DVSS.n21228 DVSS.n21226 0.00962857
R58997 DVSS.n21228 DVSS.n13611 0.00962857
R58998 DVSS.n21233 DVSS.n13611 0.00962857
R58999 DVSS.n21235 DVSS.n21233 0.00962857
R59000 DVSS.n21237 DVSS.n21235 0.00962857
R59001 DVSS.n21237 DVSS.n13608 0.00962857
R59002 DVSS.n21242 DVSS.n13608 0.00962857
R59003 DVSS.n21244 DVSS.n21242 0.00962857
R59004 DVSS.n21246 DVSS.n21244 0.00962857
R59005 DVSS.n21246 DVSS.n13605 0.00962857
R59006 DVSS.n21250 DVSS.n13605 0.00962857
R59007 DVSS.n21250 DVSS.n13569 0.00962857
R59008 DVSS.n21259 DVSS.n13569 0.00962857
R59009 DVSS.n21259 DVSS.n13567 0.00962857
R59010 DVSS.n21264 DVSS.n13567 0.00962857
R59011 DVSS.n21264 DVSS.n13564 0.00962857
R59012 DVSS.n21268 DVSS.n13564 0.00962857
R59013 DVSS.n21270 DVSS.n21268 0.00962857
R59014 DVSS.n21272 DVSS.n21270 0.00962857
R59015 DVSS.n21272 DVSS.n13562 0.00962857
R59016 DVSS.n21277 DVSS.n13562 0.00962857
R59017 DVSS.n21279 DVSS.n21277 0.00962857
R59018 DVSS.n21281 DVSS.n21279 0.00962857
R59019 DVSS.n21281 DVSS.n13559 0.00962857
R59020 DVSS.n21286 DVSS.n13559 0.00962857
R59021 DVSS.n21288 DVSS.n21286 0.00962857
R59022 DVSS.n21290 DVSS.n21288 0.00962857
R59023 DVSS.n21290 DVSS.n13555 0.00962857
R59024 DVSS.n21295 DVSS.n13555 0.00962857
R59025 DVSS.n21295 DVSS.n13556 0.00962857
R59026 DVSS.n13556 DVSS.n13515 0.00962857
R59027 DVSS.n21302 DVSS.n13515 0.00962857
R59028 DVSS.n21302 DVSS.n13513 0.00962857
R59029 DVSS.n21307 DVSS.n13513 0.00962857
R59030 DVSS.n21307 DVSS.n13511 0.00962857
R59031 DVSS.n21311 DVSS.n13511 0.00962857
R59032 DVSS.n21313 DVSS.n21311 0.00962857
R59033 DVSS.n21313 DVSS.n13509 0.00962857
R59034 DVSS.n21318 DVSS.n13509 0.00962857
R59035 DVSS.n21320 DVSS.n21318 0.00962857
R59036 DVSS.n21322 DVSS.n21320 0.00962857
R59037 DVSS.n21322 DVSS.n13506 0.00962857
R59038 DVSS.n21327 DVSS.n13506 0.00962857
R59039 DVSS.n21329 DVSS.n21327 0.00962857
R59040 DVSS.n21331 DVSS.n21329 0.00962857
R59041 DVSS.n21331 DVSS.n13503 0.00962857
R59042 DVSS.n21335 DVSS.n13503 0.00962857
R59043 DVSS.n21335 DVSS.n13464 0.00962857
R59044 DVSS.n21342 DVSS.n13464 0.00962857
R59045 DVSS.n21342 DVSS.n13462 0.00962857
R59046 DVSS.n21347 DVSS.n13462 0.00962857
R59047 DVSS.n21347 DVSS.n13460 0.00962857
R59048 DVSS.n21351 DVSS.n13460 0.00962857
R59049 DVSS.n21353 DVSS.n21351 0.00962857
R59050 DVSS.n21353 DVSS.n13458 0.00962857
R59051 DVSS.n21358 DVSS.n13458 0.00962857
R59052 DVSS.n21360 DVSS.n21358 0.00962857
R59053 DVSS.n21362 DVSS.n21360 0.00962857
R59054 DVSS.n21362 DVSS.n13455 0.00962857
R59055 DVSS.n21367 DVSS.n13455 0.00962857
R59056 DVSS.n21369 DVSS.n21367 0.00962857
R59057 DVSS.n21371 DVSS.n21369 0.00962857
R59058 DVSS.n21371 DVSS.n13452 0.00962857
R59059 DVSS.n21375 DVSS.n13452 0.00962857
R59060 DVSS.n21375 DVSS.n13418 0.00962857
R59061 DVSS.n21386 DVSS.n13418 0.00962857
R59062 DVSS.n21386 DVSS.n13416 0.00962857
R59063 DVSS.n21390 DVSS.n13416 0.00962857
R59064 DVSS.n21390 DVSS.n13414 0.00962857
R59065 DVSS.n21394 DVSS.n13414 0.00962857
R59066 DVSS.n21394 DVSS.n13410 0.00962857
R59067 DVSS.n21428 DVSS.n13410 0.00962857
R59068 DVSS.n21428 DVSS.n13412 0.00962857
R59069 DVSS.n21424 DVSS.n13412 0.00962857
R59070 DVSS.n21424 DVSS.n21416 0.00962857
R59071 DVSS.n21416 DVSS.n21415 0.00962857
R59072 DVSS.n21415 DVSS.n21399 0.00962857
R59073 DVSS.n21410 DVSS.n21399 0.00962857
R59074 DVSS.n21410 DVSS.n21408 0.00962857
R59075 DVSS.n21408 DVSS.n21406 0.00962857
R59076 DVSS.n21402 DVSS.n13376 0.00962857
R59077 DVSS.n21434 DVSS.n13376 0.00962857
R59078 DVSS.n21434 DVSS.n13374 0.00962857
R59079 DVSS.n21181 DVSS.n21180 0.00962857
R59080 DVSS.n21216 DVSS.n13614 0.00962857
R59081 DVSS.n21223 DVSS.n13614 0.00962857
R59082 DVSS.n21224 DVSS.n21223 0.00962857
R59083 DVSS.n21225 DVSS.n21224 0.00962857
R59084 DVSS.n21265 DVSS.n13566 0.00962857
R59085 DVSS.n21266 DVSS.n21265 0.00962857
R59086 DVSS.n21267 DVSS.n21266 0.00962857
R59087 DVSS.n21301 DVSS.n21300 0.00962857
R59088 DVSS.n21301 DVSS.n13512 0.00962857
R59089 DVSS.n21308 DVSS.n13512 0.00962857
R59090 DVSS.n21309 DVSS.n21308 0.00962857
R59091 DVSS.n21310 DVSS.n21309 0.00962857
R59092 DVSS.n21348 DVSS.n13461 0.00962857
R59093 DVSS.n21349 DVSS.n21348 0.00962857
R59094 DVSS.n21350 DVSS.n21349 0.00962857
R59095 DVSS.n21391 DVSS.n13415 0.00962857
R59096 DVSS.n21392 DVSS.n21391 0.00962857
R59097 DVSS.n21393 DVSS.n21392 0.00962857
R59098 DVSS.n21393 DVSS.n13409 0.00962857
R59099 DVSS.n21437 DVSS.n13373 0.00962857
R59100 DVSS.n22638 DVSS.n729 0.00962857
R59101 DVSS.n22674 DVSS.n697 0.00962857
R59102 DVSS.n22681 DVSS.n697 0.00962857
R59103 DVSS.n22682 DVSS.n22681 0.00962857
R59104 DVSS.n22683 DVSS.n22682 0.00962857
R59105 DVSS.n22723 DVSS.n644 0.00962857
R59106 DVSS.n22724 DVSS.n22723 0.00962857
R59107 DVSS.n22725 DVSS.n22724 0.00962857
R59108 DVSS.n22759 DVSS.n22758 0.00962857
R59109 DVSS.n22759 DVSS.n592 0.00962857
R59110 DVSS.n22766 DVSS.n592 0.00962857
R59111 DVSS.n22767 DVSS.n22766 0.00962857
R59112 DVSS.n22768 DVSS.n22767 0.00962857
R59113 DVSS.n22806 DVSS.n543 0.00962857
R59114 DVSS.n22807 DVSS.n22806 0.00962857
R59115 DVSS.n22808 DVSS.n22807 0.00962857
R59116 DVSS.n22840 DVSS.n492 0.00962857
R59117 DVSS.n22847 DVSS.n492 0.00962857
R59118 DVSS.n22848 DVSS.n22847 0.00962857
R59119 DVSS.n22849 DVSS.n22848 0.00962857
R59120 DVSS.n22884 DVSS.n454 0.00962857
R59121 DVSS.n7110 DVSS.n7109 0.00956767
R59122 DVSS.n6249 DVSS.n6246 0.00937536
R59123 DVSS.n6666 DVSS.n6242 0.00937536
R59124 DVSS.n12774 DVSS.n12352 0.00937536
R59125 DVSS.n12775 DVSS.n12774 0.00937536
R59126 DVSS.n6250 DVSS.n6249 0.00937536
R59127 DVSS.n6250 DVSS.n6242 0.00937536
R59128 DVSS.n20160 DVSS.n20159 0.00934831
R59129 DVSS.n20272 DVSS.n20219 0.00934831
R59130 DVSS DVSS.n20224 0.00934831
R59131 DVSS.n10156 DVSS.n2071 0.00934279
R59132 DVSS.n10488 DVSS.n1621 0.00934279
R59133 DVSS.n10157 DVSS.n10155 0.00934279
R59134 DVSS.n10489 DVSS.n1622 0.00934279
R59135 DVSS.n18901 DVSS.n14555 0.00930435
R59136 DVSS.n18945 DVSS.n14554 0.00930435
R59137 DVSS.n20084 DVSS.n14591 0.00930435
R59138 DVSS.n20672 DVSS.n14602 0.00930435
R59139 DVSS.n20649 DVSS.n14630 0.00930435
R59140 DVSS.n20200 DVSS.n14635 0.00930435
R59141 DVSS.n20416 DVSS.n20359 0.00930435
R59142 DVSS.n20447 DVSS.n20446 0.00930435
R59143 DVSS.n18893 DVSS.n14524 0.00930435
R59144 DVSS.n18951 DVSS.n14521 0.00930435
R59145 DVSS.n20096 DVSS.n20016 0.00930435
R59146 DVSS.n20174 DVSS.n14874 0.00930435
R59147 DVSS.n20185 DVSS.n20184 0.00930435
R59148 DVSS.n20231 DVSS.n14867 0.00930435
R59149 DVSS.n20371 DVSS.n14858 0.00930435
R59150 DVSS.n20332 DVSS.n14855 0.00930435
R59151 DVSS.n9766 DVSS.n2713 0.00929699
R59152 DVSS.n8334 DVSS.n8333 0.00919799
R59153 DVSS.n12002 DVSS.n11996 0.00919799
R59154 DVSS.n8338 DVSS.n3844 0.00919799
R59155 DVSS.n12001 DVSS.n11998 0.00919799
R59156 DVSS.n8996 DVSS.n8995 0.00916165
R59157 DVSS.n11105 DVSS.n1506 0.00916165
R59158 DVSS.n21171 DVSS.n13367 0.00910927
R59159 DVSS.n19908 DVSS.n13367 0.00910927
R59160 DVSS.n21010 DVSS.n13368 0.00910927
R59161 DVSS.n14848 DVSS.n13368 0.00910927
R59162 DVSS.n15867 DVSS.n15862 0.00909155
R59163 DVSS.n17928 DVSS.n15766 0.00909155
R59164 DVSS.n18016 DVSS.n15558 0.00902113
R59165 DVSS.n17866 DVSS.n17865 0.0089507
R59166 DVSS.n17947 DVSS.n17945 0.0089507
R59167 DVSS.n8110 DVSS.n4023 0.00894978
R59168 DVSS.n12762 DVSS.n12458 0.00894978
R59169 DVSS.n8109 DVSS.n4024 0.00894978
R59170 DVSS.n12763 DVSS.n12554 0.00894978
R59171 DVSS.n22610 DVSS.n743 0.0089375
R59172 DVSS.n22911 DVSS.n443 0.0089375
R59173 DVSS.n16539 DVSS.n16478 0.00888983
R59174 DVSS.n18110 DVSS.n18109 0.00888983
R59175 DVSS.n18151 DVSS.n15563 0.00888028
R59176 DVSS.n22582 DVSS.n22581 0.00887209
R59177 DVSS.n22940 DVSS.n22939 0.00887209
R59178 DVSS.n20369 DVSS 0.0088427
R59179 DVSS.n17897 DVSS.n15802 0.00880986
R59180 DVSS.n18043 DVSS.n15693 0.00880986
R59181 DVSS.n17812 DVSS.n15905 0.00873944
R59182 DVSS.n5869 DVSS.n5530 0.00871477
R59183 DVSS.n7805 DVSS.n4819 0.00871477
R59184 DVSS.n5871 DVSS.n5529 0.00871477
R59185 DVSS.n7804 DVSS.n4820 0.00871477
R59186 DVSS.n12746 DVSS.n12554 0.0087125
R59187 DVSS.n12745 DVSS.n12458 0.0087125
R59188 DVSS.n6596 DVSS.n6235 0.0087125
R59189 DVSS.n6260 DVSS.n6236 0.0087125
R59190 DVSS.n15827 DVSS.n15806 0.00866901
R59191 DVSS.n17961 DVSS.n15697 0.00866901
R59192 DVSS.n8996 DVSS.n3040 0.0086203
R59193 DVSS.n13346 DVSS.n11105 0.0086203
R59194 DVSS.n17796 DVSS.n15900 0.00859859
R59195 DVSS.n15914 DVSS.n15897 0.00859859
R59196 DVSS.n18937 DVSS.n18877 0.00858989
R59197 DVSS.n20117 DVSS.n20057 0.00858989
R59198 DVSS.n20155 DVSS.n20154 0.00858989
R59199 DVSS.n20274 DVSS.n20218 0.00858989
R59200 DVSS.n20300 DVSS.n20299 0.00858989
R59201 DVSS.n20367 DVSS.n14688 0.00858989
R59202 DVSS.n18009 DVSS 0.00852817
R59203 DVSS.n17884 DVSS.n15816 0.00852817
R59204 DVSS.n17963 DVSS.n15698 0.00852817
R59205 DVSS.n9767 DVSS.n9766 0.00848496
R59206 DVSS.n17814 DVSS.n15893 0.00845775
R59207 DVSS.n17906 DVSS.n15821 0.00838732
R59208 DVSS.n18040 DVSS.n15701 0.00838732
R59209 DVSS.n12773 DVSS.n12772 0.008375
R59210 DVSS.n7811 DVSS.n7810 0.008375
R59211 DVSS.n6454 DVSS.n6453 0.008375
R59212 DVSS.n16323 DVSS.n16318 0.00834286
R59213 DVSS.n16700 DVSS.n16161 0.00834286
R59214 DVSS.n16048 DVSS.n16025 0.00834286
R59215 DVSS.n16865 DVSS.n16846 0.00834286
R59216 DVSS.n15276 DVSS.n15249 0.00834286
R59217 DVSS.n15409 DVSS.n15390 0.00834286
R59218 DVSS.n18415 DVSS.n18390 0.00834286
R59219 DVSS.n14971 DVSS.n14953 0.00834286
R59220 DVSS.n20786 DVSS.n20716 0.00834286
R59221 DVSS.n20869 DVSS.n14436 0.00834286
R59222 DVSS.n13607 DVSS.n13602 0.00834286
R59223 DVSS.n21319 DVSS.n13492 0.00834286
R59224 DVSS.n690 DVSS.n685 0.00834286
R59225 DVSS.n22777 DVSS.n577 0.00834286
R59226 DVSS.n18004 DVSS.n15549 0.0083169
R59227 DVSS.n16755 DVSS.n15601 0.00827857
R59228 DVSS.n15524 DVSS.n15502 0.00827857
R59229 DVSS.n18267 DVSS.n18229 0.00827857
R59230 DVSS.n15119 DVSS.n15113 0.00827857
R59231 DVSS.n20960 DVSS.n14347 0.00827857
R59232 DVSS.n21414 DVSS.n13405 0.00827857
R59233 DVSS.n22860 DVSS.n481 0.00827857
R59234 DVSS.n17861 DVSS.n15850 0.00824648
R59235 DVSS.n15771 DVSS.n15757 0.00824648
R59236 DVSS.n8993 DVSS.n2934 0.00823154
R59237 DVSS.n10767 DVSS.n1510 0.00823154
R59238 DVSS.n8994 DVSS.n8991 0.00823154
R59239 DVSS.n10769 DVSS.n1508 0.00823154
R59240 DVSS.n16640 DVSS.n16639 0.00821429
R59241 DVSS.n16227 DVSS.n16164 0.00821429
R59242 DVSS.n17653 DVSS.n16030 0.00821429
R59243 DVSS.n16881 DVSS.n16851 0.00821429
R59244 DVSS.n18380 DVSS.n15253 0.00821429
R59245 DVSS.n15425 DVSS.n15395 0.00821429
R59246 DVSS.n18472 DVSS.n18400 0.00821429
R59247 DVSS.n14993 DVSS.n14957 0.00821429
R59248 DVSS.n20805 DVSS.n14506 0.00821429
R59249 DVSS.n20888 DVSS.n20886 0.00821429
R59250 DVSS.n21258 DVSS.n21257 0.00821429
R59251 DVSS.n21338 DVSS.n21336 0.00821429
R59252 DVSS.n7448 DVSS.n7110 0.00821429
R59253 DVSS.n22716 DVSS.n22715 0.00821429
R59254 DVSS.n22796 DVSS.n22794 0.00821429
R59255 DVSS.n18761 DVSS.n18757 0.00819509
R59256 DVSS.n20471 DVSS.n14713 0.00819509
R59257 DVSS.n18757 DVSS.n18755 0.00819509
R59258 DVSS.n20612 DVSS.n14713 0.00819509
R59259 DVSS.n20558 DVSS.n20489 0.00817918
R59260 DVSS.n18018 DVSS.n15551 0.00817606
R59261 DVSS.n18119 DVSS.n15608 0.00815
R59262 DVSS.n15530 DVSS.n15498 0.00815
R59263 DVSS.n18246 DVSS.n18224 0.00815
R59264 DVSS.n15124 DVSS.n15108 0.00815
R59265 DVSS.n20979 DVSS.n20978 0.00815
R59266 DVSS.n21433 DVSS.n21432 0.00815
R59267 DVSS.n22880 DVSS.n22879 0.00815
R59268 DVSS.n17844 DVSS.n15854 0.00810563
R59269 DVSS.n17926 DVSS.n15761 0.00810563
R59270 DVSS.n18710 DVSS.n18708 0.00810135
R59271 DVSS.n16671 DVSS.n16257 0.00808571
R59272 DVSS.n16787 DVSS.n15656 0.00808571
R59273 DVSS.n17639 DVSS.n16076 0.00808571
R59274 DVSS.n17588 DVSS.n17543 0.00808571
R59275 DVSS.n15348 DVSS.n15311 0.00808571
R59276 DVSS.n18298 DVSS.n15463 0.00808571
R59277 DVSS.n20005 DVSS.n14877 0.00808571
R59278 DVSS.n15060 DVSS.n15020 0.00808571
R59279 DVSS.n20839 DVSS.n14477 0.00808571
R59280 DVSS.n20918 DVSS.n14379 0.00808571
R59281 DVSS.n21289 DVSS.n13535 0.00808571
R59282 DVSS.n21368 DVSS.n13438 0.00808571
R59283 DVSS.n22747 DVSS.n617 0.00808571
R59284 DVSS.n22826 DVSS.n518 0.00808571
R59285 DVSS.n18935 DVSS 0.00808427
R59286 DVSS.n18937 DVSS.n18912 0.00808427
R59287 DVSS.n20117 DVSS.n20056 0.00808427
R59288 DVSS.n20154 DVSS.n20040 0.00808427
R59289 DVSS.n20274 DVSS.n20222 0.00808427
R59290 DVSS.n20299 DVSS.n14660 0.00808427
R59291 DVSS.n20367 DVSS.n14683 0.00808427
R59292 DVSS.n7063 DVSS.n5528 0.00807895
R59293 DVSS.n7802 DVSS.n7801 0.00807895
R59294 DVSS.n16586 DVSS.n16556 0.00802143
R59295 DVSS.n15981 DVSS.n15952 0.00802143
R59296 DVSS.n17738 DVSS.n17687 0.00802143
R59297 DVSS.n15189 DVSS.n15180 0.00802143
R59298 DVSS.n20755 DVSS.n13717 0.00802143
R59299 DVSS.n21199 DVSS.n13647 0.00802143
R59300 DVSS.n22653 DVSS.n724 0.00802143
R59301 DVSS.n22623 DVSS.n22622 0.008
R59302 DVSS.n22899 DVSS.n22898 0.008
R59303 DVSS.n17833 DVSS.n15856 0.00796479
R59304 DVSS.n12349 DVSS.n12347 0.00796421
R59305 DVSS.n13104 DVSS.n12350 0.00796421
R59306 DVSS.n12755 DVSS.n12749 0.00796421
R59307 DVSS.n12753 DVSS.n12354 0.00796421
R59308 DVSS.n12769 DVSS.n12357 0.00796421
R59309 DVSS.n12363 DVSS.n12358 0.00796421
R59310 DVSS.n12505 DVSS.n12457 0.00796421
R59311 DVSS.n12507 DVSS.n12364 0.00796421
R59312 DVSS.n12504 DVSS.n12456 0.00796421
R59313 DVSS.n12508 DVSS.n12365 0.00796421
R59314 DVSS.n12503 DVSS.n12455 0.00796421
R59315 DVSS.n12509 DVSS.n12366 0.00796421
R59316 DVSS.n12502 DVSS.n12454 0.00796421
R59317 DVSS.n12510 DVSS.n12367 0.00796421
R59318 DVSS.n12501 DVSS.n12453 0.00796421
R59319 DVSS.n12511 DVSS.n12368 0.00796421
R59320 DVSS.n12500 DVSS.n12452 0.00796421
R59321 DVSS.n12512 DVSS.n12369 0.00796421
R59322 DVSS.n12499 DVSS.n12451 0.00796421
R59323 DVSS.n12513 DVSS.n12370 0.00796421
R59324 DVSS.n12498 DVSS.n12450 0.00796421
R59325 DVSS.n12514 DVSS.n12371 0.00796421
R59326 DVSS.n12497 DVSS.n12449 0.00796421
R59327 DVSS.n12515 DVSS.n12372 0.00796421
R59328 DVSS.n12496 DVSS.n12448 0.00796421
R59329 DVSS.n12516 DVSS.n12373 0.00796421
R59330 DVSS.n12495 DVSS.n12447 0.00796421
R59331 DVSS.n12517 DVSS.n12374 0.00796421
R59332 DVSS.n12494 DVSS.n12446 0.00796421
R59333 DVSS.n12518 DVSS.n12375 0.00796421
R59334 DVSS.n12493 DVSS.n12445 0.00796421
R59335 DVSS.n12519 DVSS.n12376 0.00796421
R59336 DVSS.n12492 DVSS.n12444 0.00796421
R59337 DVSS.n12520 DVSS.n12377 0.00796421
R59338 DVSS.n12491 DVSS.n12443 0.00796421
R59339 DVSS.n12521 DVSS.n12378 0.00796421
R59340 DVSS.n12490 DVSS.n12442 0.00796421
R59341 DVSS.n12522 DVSS.n12379 0.00796421
R59342 DVSS.n12489 DVSS.n12441 0.00796421
R59343 DVSS.n12523 DVSS.n12380 0.00796421
R59344 DVSS.n12488 DVSS.n12440 0.00796421
R59345 DVSS.n12524 DVSS.n12381 0.00796421
R59346 DVSS.n12487 DVSS.n12439 0.00796421
R59347 DVSS.n12525 DVSS.n12382 0.00796421
R59348 DVSS.n12486 DVSS.n12438 0.00796421
R59349 DVSS.n12526 DVSS.n12383 0.00796421
R59350 DVSS.n12485 DVSS.n12437 0.00796421
R59351 DVSS.n12527 DVSS.n12384 0.00796421
R59352 DVSS.n12484 DVSS.n12436 0.00796421
R59353 DVSS.n12528 DVSS.n12385 0.00796421
R59354 DVSS.n12483 DVSS.n12435 0.00796421
R59355 DVSS.n12529 DVSS.n12386 0.00796421
R59356 DVSS.n12482 DVSS.n12434 0.00796421
R59357 DVSS.n12530 DVSS.n12387 0.00796421
R59358 DVSS.n12481 DVSS.n12433 0.00796421
R59359 DVSS.n12531 DVSS.n12388 0.00796421
R59360 DVSS.n12480 DVSS.n12432 0.00796421
R59361 DVSS.n12532 DVSS.n12389 0.00796421
R59362 DVSS.n12479 DVSS.n12431 0.00796421
R59363 DVSS.n12533 DVSS.n12390 0.00796421
R59364 DVSS.n12478 DVSS.n12430 0.00796421
R59365 DVSS.n12534 DVSS.n12391 0.00796421
R59366 DVSS.n12477 DVSS.n12429 0.00796421
R59367 DVSS.n12535 DVSS.n12392 0.00796421
R59368 DVSS.n12476 DVSS.n12428 0.00796421
R59369 DVSS.n12536 DVSS.n12393 0.00796421
R59370 DVSS.n12475 DVSS.n12427 0.00796421
R59371 DVSS.n12537 DVSS.n12394 0.00796421
R59372 DVSS.n12474 DVSS.n12426 0.00796421
R59373 DVSS.n12538 DVSS.n12395 0.00796421
R59374 DVSS.n12473 DVSS.n12425 0.00796421
R59375 DVSS.n12539 DVSS.n12396 0.00796421
R59376 DVSS.n12472 DVSS.n12424 0.00796421
R59377 DVSS.n12540 DVSS.n12397 0.00796421
R59378 DVSS.n12471 DVSS.n12423 0.00796421
R59379 DVSS.n12541 DVSS.n12398 0.00796421
R59380 DVSS.n12470 DVSS.n12422 0.00796421
R59381 DVSS.n12542 DVSS.n12399 0.00796421
R59382 DVSS.n12469 DVSS.n12421 0.00796421
R59383 DVSS.n12543 DVSS.n12400 0.00796421
R59384 DVSS.n12468 DVSS.n12420 0.00796421
R59385 DVSS.n12544 DVSS.n12401 0.00796421
R59386 DVSS.n12467 DVSS.n12419 0.00796421
R59387 DVSS.n12545 DVSS.n12402 0.00796421
R59388 DVSS.n12466 DVSS.n12418 0.00796421
R59389 DVSS.n12546 DVSS.n12403 0.00796421
R59390 DVSS.n12465 DVSS.n12417 0.00796421
R59391 DVSS.n12547 DVSS.n12404 0.00796421
R59392 DVSS.n12464 DVSS.n12416 0.00796421
R59393 DVSS.n12548 DVSS.n12405 0.00796421
R59394 DVSS.n12463 DVSS.n12415 0.00796421
R59395 DVSS.n12549 DVSS.n12406 0.00796421
R59396 DVSS.n12462 DVSS.n12414 0.00796421
R59397 DVSS.n12550 DVSS.n12407 0.00796421
R59398 DVSS.n12461 DVSS.n12413 0.00796421
R59399 DVSS.n12551 DVSS.n12408 0.00796421
R59400 DVSS.n12460 DVSS.n12412 0.00796421
R59401 DVSS.n12552 DVSS.n12409 0.00796421
R59402 DVSS.n12459 DVSS.n12411 0.00796421
R59403 DVSS.n12743 DVSS.n12742 0.00796421
R59404 DVSS.n12745 DVSS.n12410 0.00796421
R59405 DVSS.n6663 DVSS.n6254 0.00796421
R59406 DVSS.n6665 DVSS.n6245 0.00796421
R59407 DVSS.n6662 DVSS.n6255 0.00796421
R59408 DVSS.n6658 DVSS.n6248 0.00796421
R59409 DVSS.n6650 DVSS.n6311 0.00796421
R59410 DVSS.n6310 DVSS.n6307 0.00796421
R59411 DVSS.n6649 DVSS.n6313 0.00796421
R59412 DVSS.n6312 DVSS.n6306 0.00796421
R59413 DVSS.n6648 DVSS.n6315 0.00796421
R59414 DVSS.n6314 DVSS.n6305 0.00796421
R59415 DVSS.n6647 DVSS.n6317 0.00796421
R59416 DVSS.n6316 DVSS.n6304 0.00796421
R59417 DVSS.n6646 DVSS.n6319 0.00796421
R59418 DVSS.n6318 DVSS.n6303 0.00796421
R59419 DVSS.n6645 DVSS.n6321 0.00796421
R59420 DVSS.n6320 DVSS.n6302 0.00796421
R59421 DVSS.n6644 DVSS.n6323 0.00796421
R59422 DVSS.n6322 DVSS.n6301 0.00796421
R59423 DVSS.n6643 DVSS.n6325 0.00796421
R59424 DVSS.n6324 DVSS.n6300 0.00796421
R59425 DVSS.n6642 DVSS.n6327 0.00796421
R59426 DVSS.n6326 DVSS.n6299 0.00796421
R59427 DVSS.n6641 DVSS.n6329 0.00796421
R59428 DVSS.n6328 DVSS.n6298 0.00796421
R59429 DVSS.n6640 DVSS.n6331 0.00796421
R59430 DVSS.n6330 DVSS.n6297 0.00796421
R59431 DVSS.n6639 DVSS.n6333 0.00796421
R59432 DVSS.n6332 DVSS.n6296 0.00796421
R59433 DVSS.n6638 DVSS.n6335 0.00796421
R59434 DVSS.n6334 DVSS.n6295 0.00796421
R59435 DVSS.n6637 DVSS.n6337 0.00796421
R59436 DVSS.n6336 DVSS.n6294 0.00796421
R59437 DVSS.n6636 DVSS.n6339 0.00796421
R59438 DVSS.n6338 DVSS.n6293 0.00796421
R59439 DVSS.n6635 DVSS.n6341 0.00796421
R59440 DVSS.n6340 DVSS.n6292 0.00796421
R59441 DVSS.n6634 DVSS.n6343 0.00796421
R59442 DVSS.n6342 DVSS.n6291 0.00796421
R59443 DVSS.n6633 DVSS.n6345 0.00796421
R59444 DVSS.n6344 DVSS.n6290 0.00796421
R59445 DVSS.n6632 DVSS.n6347 0.00796421
R59446 DVSS.n6346 DVSS.n6289 0.00796421
R59447 DVSS.n6631 DVSS.n6349 0.00796421
R59448 DVSS.n6348 DVSS.n6288 0.00796421
R59449 DVSS.n6630 DVSS.n6351 0.00796421
R59450 DVSS.n6350 DVSS.n6287 0.00796421
R59451 DVSS.n6629 DVSS.n6353 0.00796421
R59452 DVSS.n6352 DVSS.n6286 0.00796421
R59453 DVSS.n6628 DVSS.n6355 0.00796421
R59454 DVSS.n6354 DVSS.n6285 0.00796421
R59455 DVSS.n6627 DVSS.n6357 0.00796421
R59456 DVSS.n6356 DVSS.n6284 0.00796421
R59457 DVSS.n6626 DVSS.n6359 0.00796421
R59458 DVSS.n6358 DVSS.n6283 0.00796421
R59459 DVSS.n6625 DVSS.n6361 0.00796421
R59460 DVSS.n6360 DVSS.n6282 0.00796421
R59461 DVSS.n6624 DVSS.n6363 0.00796421
R59462 DVSS.n6362 DVSS.n6281 0.00796421
R59463 DVSS.n6623 DVSS.n6365 0.00796421
R59464 DVSS.n6364 DVSS.n6280 0.00796421
R59465 DVSS.n6622 DVSS.n6367 0.00796421
R59466 DVSS.n6366 DVSS.n6279 0.00796421
R59467 DVSS.n6621 DVSS.n6369 0.00796421
R59468 DVSS.n6368 DVSS.n6278 0.00796421
R59469 DVSS.n6620 DVSS.n6371 0.00796421
R59470 DVSS.n6370 DVSS.n6277 0.00796421
R59471 DVSS.n6619 DVSS.n6373 0.00796421
R59472 DVSS.n6372 DVSS.n6276 0.00796421
R59473 DVSS.n6618 DVSS.n6375 0.00796421
R59474 DVSS.n6374 DVSS.n6275 0.00796421
R59475 DVSS.n6617 DVSS.n6377 0.00796421
R59476 DVSS.n6376 DVSS.n6274 0.00796421
R59477 DVSS.n6616 DVSS.n6379 0.00796421
R59478 DVSS.n6378 DVSS.n6273 0.00796421
R59479 DVSS.n6615 DVSS.n6381 0.00796421
R59480 DVSS.n6380 DVSS.n6272 0.00796421
R59481 DVSS.n6614 DVSS.n6383 0.00796421
R59482 DVSS.n6382 DVSS.n6271 0.00796421
R59483 DVSS.n6613 DVSS.n6385 0.00796421
R59484 DVSS.n6384 DVSS.n6270 0.00796421
R59485 DVSS.n6612 DVSS.n6387 0.00796421
R59486 DVSS.n6386 DVSS.n6269 0.00796421
R59487 DVSS.n6611 DVSS.n6389 0.00796421
R59488 DVSS.n6388 DVSS.n6268 0.00796421
R59489 DVSS.n6610 DVSS.n6391 0.00796421
R59490 DVSS.n6390 DVSS.n6267 0.00796421
R59491 DVSS.n6609 DVSS.n6393 0.00796421
R59492 DVSS.n6392 DVSS.n6266 0.00796421
R59493 DVSS.n6608 DVSS.n6395 0.00796421
R59494 DVSS.n6394 DVSS.n6265 0.00796421
R59495 DVSS.n6607 DVSS.n6397 0.00796421
R59496 DVSS.n6396 DVSS.n6264 0.00796421
R59497 DVSS.n6606 DVSS.n6399 0.00796421
R59498 DVSS.n6398 DVSS.n6263 0.00796421
R59499 DVSS.n6605 DVSS.n6401 0.00796421
R59500 DVSS.n6400 DVSS.n6262 0.00796421
R59501 DVSS.n6604 DVSS.n6403 0.00796421
R59502 DVSS.n6402 DVSS.n6261 0.00796421
R59503 DVSS.n6603 DVSS.n6601 0.00796421
R59504 DVSS.n6404 DVSS.n6309 0.00796421
R59505 DVSS.n6651 DVSS.n6260 0.00796421
R59506 DVSS.n6651 DVSS.n6309 0.00796421
R59507 DVSS.n12743 DVSS.n12410 0.00796421
R59508 DVSS.n12742 DVSS.n12411 0.00796421
R59509 DVSS.n12459 DVSS.n12409 0.00796421
R59510 DVSS.n12552 DVSS.n12412 0.00796421
R59511 DVSS.n12460 DVSS.n12408 0.00796421
R59512 DVSS.n12551 DVSS.n12413 0.00796421
R59513 DVSS.n12461 DVSS.n12407 0.00796421
R59514 DVSS.n12550 DVSS.n12414 0.00796421
R59515 DVSS.n12462 DVSS.n12406 0.00796421
R59516 DVSS.n12549 DVSS.n12415 0.00796421
R59517 DVSS.n12463 DVSS.n12405 0.00796421
R59518 DVSS.n12548 DVSS.n12416 0.00796421
R59519 DVSS.n12464 DVSS.n12404 0.00796421
R59520 DVSS.n12547 DVSS.n12417 0.00796421
R59521 DVSS.n12465 DVSS.n12403 0.00796421
R59522 DVSS.n12546 DVSS.n12418 0.00796421
R59523 DVSS.n12466 DVSS.n12402 0.00796421
R59524 DVSS.n12545 DVSS.n12419 0.00796421
R59525 DVSS.n12467 DVSS.n12401 0.00796421
R59526 DVSS.n12544 DVSS.n12420 0.00796421
R59527 DVSS.n12468 DVSS.n12400 0.00796421
R59528 DVSS.n12543 DVSS.n12421 0.00796421
R59529 DVSS.n12469 DVSS.n12399 0.00796421
R59530 DVSS.n12542 DVSS.n12422 0.00796421
R59531 DVSS.n12470 DVSS.n12398 0.00796421
R59532 DVSS.n12541 DVSS.n12423 0.00796421
R59533 DVSS.n12471 DVSS.n12397 0.00796421
R59534 DVSS.n12540 DVSS.n12424 0.00796421
R59535 DVSS.n12472 DVSS.n12396 0.00796421
R59536 DVSS.n12539 DVSS.n12425 0.00796421
R59537 DVSS.n12473 DVSS.n12395 0.00796421
R59538 DVSS.n12538 DVSS.n12426 0.00796421
R59539 DVSS.n12474 DVSS.n12394 0.00796421
R59540 DVSS.n12537 DVSS.n12427 0.00796421
R59541 DVSS.n12475 DVSS.n12393 0.00796421
R59542 DVSS.n12536 DVSS.n12428 0.00796421
R59543 DVSS.n12476 DVSS.n12392 0.00796421
R59544 DVSS.n12535 DVSS.n12429 0.00796421
R59545 DVSS.n12477 DVSS.n12391 0.00796421
R59546 DVSS.n12534 DVSS.n12430 0.00796421
R59547 DVSS.n12478 DVSS.n12390 0.00796421
R59548 DVSS.n12533 DVSS.n12431 0.00796421
R59549 DVSS.n12479 DVSS.n12389 0.00796421
R59550 DVSS.n12532 DVSS.n12432 0.00796421
R59551 DVSS.n12480 DVSS.n12388 0.00796421
R59552 DVSS.n12531 DVSS.n12433 0.00796421
R59553 DVSS.n12481 DVSS.n12387 0.00796421
R59554 DVSS.n12530 DVSS.n12434 0.00796421
R59555 DVSS.n12482 DVSS.n12386 0.00796421
R59556 DVSS.n12529 DVSS.n12435 0.00796421
R59557 DVSS.n12483 DVSS.n12385 0.00796421
R59558 DVSS.n12528 DVSS.n12436 0.00796421
R59559 DVSS.n12484 DVSS.n12384 0.00796421
R59560 DVSS.n12527 DVSS.n12437 0.00796421
R59561 DVSS.n12485 DVSS.n12383 0.00796421
R59562 DVSS.n12526 DVSS.n12438 0.00796421
R59563 DVSS.n12486 DVSS.n12382 0.00796421
R59564 DVSS.n12525 DVSS.n12439 0.00796421
R59565 DVSS.n12487 DVSS.n12381 0.00796421
R59566 DVSS.n12524 DVSS.n12440 0.00796421
R59567 DVSS.n12488 DVSS.n12380 0.00796421
R59568 DVSS.n12523 DVSS.n12441 0.00796421
R59569 DVSS.n12489 DVSS.n12379 0.00796421
R59570 DVSS.n12522 DVSS.n12442 0.00796421
R59571 DVSS.n12490 DVSS.n12378 0.00796421
R59572 DVSS.n12521 DVSS.n12443 0.00796421
R59573 DVSS.n12491 DVSS.n12377 0.00796421
R59574 DVSS.n12520 DVSS.n12444 0.00796421
R59575 DVSS.n12492 DVSS.n12376 0.00796421
R59576 DVSS.n12519 DVSS.n12445 0.00796421
R59577 DVSS.n12493 DVSS.n12375 0.00796421
R59578 DVSS.n12518 DVSS.n12446 0.00796421
R59579 DVSS.n12494 DVSS.n12374 0.00796421
R59580 DVSS.n12517 DVSS.n12447 0.00796421
R59581 DVSS.n12495 DVSS.n12373 0.00796421
R59582 DVSS.n12516 DVSS.n12448 0.00796421
R59583 DVSS.n12496 DVSS.n12372 0.00796421
R59584 DVSS.n12515 DVSS.n12449 0.00796421
R59585 DVSS.n12497 DVSS.n12371 0.00796421
R59586 DVSS.n12514 DVSS.n12450 0.00796421
R59587 DVSS.n12498 DVSS.n12370 0.00796421
R59588 DVSS.n12513 DVSS.n12451 0.00796421
R59589 DVSS.n12499 DVSS.n12369 0.00796421
R59590 DVSS.n12512 DVSS.n12452 0.00796421
R59591 DVSS.n12500 DVSS.n12368 0.00796421
R59592 DVSS.n12511 DVSS.n12453 0.00796421
R59593 DVSS.n12501 DVSS.n12367 0.00796421
R59594 DVSS.n12510 DVSS.n12454 0.00796421
R59595 DVSS.n12502 DVSS.n12366 0.00796421
R59596 DVSS.n12509 DVSS.n12455 0.00796421
R59597 DVSS.n12503 DVSS.n12365 0.00796421
R59598 DVSS.n12508 DVSS.n12456 0.00796421
R59599 DVSS.n12504 DVSS.n12364 0.00796421
R59600 DVSS.n12507 DVSS.n12457 0.00796421
R59601 DVSS.n12505 DVSS.n12363 0.00796421
R59602 DVSS.n12769 DVSS.n12358 0.00796421
R59603 DVSS.n12362 DVSS.n12357 0.00796421
R59604 DVSS.n6659 DVSS.n6658 0.00796421
R59605 DVSS.n12753 DVSS.n12752 0.00796421
R59606 DVSS.n6660 DVSS.n6255 0.00796421
R59607 DVSS.n12759 DVSS.n12755 0.00796421
R59608 DVSS.n6650 DVSS.n6308 0.00796421
R59609 DVSS.n6311 DVSS.n6310 0.00796421
R59610 DVSS.n6649 DVSS.n6307 0.00796421
R59611 DVSS.n6313 DVSS.n6312 0.00796421
R59612 DVSS.n6648 DVSS.n6306 0.00796421
R59613 DVSS.n6315 DVSS.n6314 0.00796421
R59614 DVSS.n6647 DVSS.n6305 0.00796421
R59615 DVSS.n6317 DVSS.n6316 0.00796421
R59616 DVSS.n6646 DVSS.n6304 0.00796421
R59617 DVSS.n6319 DVSS.n6318 0.00796421
R59618 DVSS.n6645 DVSS.n6303 0.00796421
R59619 DVSS.n6321 DVSS.n6320 0.00796421
R59620 DVSS.n6644 DVSS.n6302 0.00796421
R59621 DVSS.n6323 DVSS.n6322 0.00796421
R59622 DVSS.n6643 DVSS.n6301 0.00796421
R59623 DVSS.n6325 DVSS.n6324 0.00796421
R59624 DVSS.n6642 DVSS.n6300 0.00796421
R59625 DVSS.n6327 DVSS.n6326 0.00796421
R59626 DVSS.n6641 DVSS.n6299 0.00796421
R59627 DVSS.n6329 DVSS.n6328 0.00796421
R59628 DVSS.n6640 DVSS.n6298 0.00796421
R59629 DVSS.n6331 DVSS.n6330 0.00796421
R59630 DVSS.n6639 DVSS.n6297 0.00796421
R59631 DVSS.n6333 DVSS.n6332 0.00796421
R59632 DVSS.n6638 DVSS.n6296 0.00796421
R59633 DVSS.n6335 DVSS.n6334 0.00796421
R59634 DVSS.n6637 DVSS.n6295 0.00796421
R59635 DVSS.n6337 DVSS.n6336 0.00796421
R59636 DVSS.n6636 DVSS.n6294 0.00796421
R59637 DVSS.n6339 DVSS.n6338 0.00796421
R59638 DVSS.n6635 DVSS.n6293 0.00796421
R59639 DVSS.n6341 DVSS.n6340 0.00796421
R59640 DVSS.n6634 DVSS.n6292 0.00796421
R59641 DVSS.n6343 DVSS.n6342 0.00796421
R59642 DVSS.n6633 DVSS.n6291 0.00796421
R59643 DVSS.n6345 DVSS.n6344 0.00796421
R59644 DVSS.n6632 DVSS.n6290 0.00796421
R59645 DVSS.n6347 DVSS.n6346 0.00796421
R59646 DVSS.n6631 DVSS.n6289 0.00796421
R59647 DVSS.n6349 DVSS.n6348 0.00796421
R59648 DVSS.n6630 DVSS.n6288 0.00796421
R59649 DVSS.n6351 DVSS.n6350 0.00796421
R59650 DVSS.n6629 DVSS.n6287 0.00796421
R59651 DVSS.n6353 DVSS.n6352 0.00796421
R59652 DVSS.n6628 DVSS.n6286 0.00796421
R59653 DVSS.n6355 DVSS.n6354 0.00796421
R59654 DVSS.n6627 DVSS.n6285 0.00796421
R59655 DVSS.n6357 DVSS.n6356 0.00796421
R59656 DVSS.n6626 DVSS.n6284 0.00796421
R59657 DVSS.n6359 DVSS.n6358 0.00796421
R59658 DVSS.n6625 DVSS.n6283 0.00796421
R59659 DVSS.n6361 DVSS.n6360 0.00796421
R59660 DVSS.n6624 DVSS.n6282 0.00796421
R59661 DVSS.n6363 DVSS.n6362 0.00796421
R59662 DVSS.n6623 DVSS.n6281 0.00796421
R59663 DVSS.n6365 DVSS.n6364 0.00796421
R59664 DVSS.n6622 DVSS.n6280 0.00796421
R59665 DVSS.n6367 DVSS.n6366 0.00796421
R59666 DVSS.n6621 DVSS.n6279 0.00796421
R59667 DVSS.n6369 DVSS.n6368 0.00796421
R59668 DVSS.n6620 DVSS.n6278 0.00796421
R59669 DVSS.n6371 DVSS.n6370 0.00796421
R59670 DVSS.n6619 DVSS.n6277 0.00796421
R59671 DVSS.n6373 DVSS.n6372 0.00796421
R59672 DVSS.n6618 DVSS.n6276 0.00796421
R59673 DVSS.n6375 DVSS.n6374 0.00796421
R59674 DVSS.n6617 DVSS.n6275 0.00796421
R59675 DVSS.n6377 DVSS.n6376 0.00796421
R59676 DVSS.n6616 DVSS.n6274 0.00796421
R59677 DVSS.n6379 DVSS.n6378 0.00796421
R59678 DVSS.n6615 DVSS.n6273 0.00796421
R59679 DVSS.n6381 DVSS.n6380 0.00796421
R59680 DVSS.n6614 DVSS.n6272 0.00796421
R59681 DVSS.n6383 DVSS.n6382 0.00796421
R59682 DVSS.n6613 DVSS.n6271 0.00796421
R59683 DVSS.n6385 DVSS.n6384 0.00796421
R59684 DVSS.n6612 DVSS.n6270 0.00796421
R59685 DVSS.n6387 DVSS.n6386 0.00796421
R59686 DVSS.n6611 DVSS.n6269 0.00796421
R59687 DVSS.n6389 DVSS.n6388 0.00796421
R59688 DVSS.n6610 DVSS.n6268 0.00796421
R59689 DVSS.n6391 DVSS.n6390 0.00796421
R59690 DVSS.n6609 DVSS.n6267 0.00796421
R59691 DVSS.n6393 DVSS.n6392 0.00796421
R59692 DVSS.n6608 DVSS.n6266 0.00796421
R59693 DVSS.n6395 DVSS.n6394 0.00796421
R59694 DVSS.n6607 DVSS.n6265 0.00796421
R59695 DVSS.n6397 DVSS.n6396 0.00796421
R59696 DVSS.n6606 DVSS.n6264 0.00796421
R59697 DVSS.n6399 DVSS.n6398 0.00796421
R59698 DVSS.n6605 DVSS.n6263 0.00796421
R59699 DVSS.n6401 DVSS.n6400 0.00796421
R59700 DVSS.n6604 DVSS.n6262 0.00796421
R59701 DVSS.n6403 DVSS.n6402 0.00796421
R59702 DVSS.n6603 DVSS.n6261 0.00796421
R59703 DVSS.n6601 DVSS.n6404 0.00796421
R59704 DVSS.n12347 DVSS.n12345 0.00796421
R59705 DVSS.n6254 DVSS.n6244 0.00796421
R59706 DVSS.n12350 DVSS.n12344 0.00796421
R59707 DVSS.n6245 DVSS.n6243 0.00796421
R59708 DVSS.n20665 DVSS 0.00795787
R59709 DVSS.n16283 DVSS.n16261 0.00795714
R59710 DVSS.n16803 DVSS.n15660 0.00795714
R59711 DVSS.n16117 DVSS.n16080 0.00795714
R59712 DVSS.n17606 DVSS.n16894 0.00795714
R59713 DVSS.n18345 DVSS.n15298 0.00795714
R59714 DVSS.n18316 DVSS.n15438 0.00795714
R59715 DVSS.n18456 DVSS.n14881 0.00795714
R59716 DVSS.n19972 DVSS.n15006 0.00795714
R59717 DVSS.n14498 DVSS.n14481 0.00795714
R59718 DVSS.n20902 DVSS.n14383 0.00795714
R59719 DVSS.n13561 DVSS.n13539 0.00795714
R59720 DVSS.n21352 DVSS.n13442 0.00795714
R59721 DVSS.n639 DVSS.n621 0.00795714
R59722 DVSS.n22810 DVSS.n522 0.00795714
R59723 DVSS.n9462 DVSS.n2725 0.007925
R59724 DVSS.n13332 DVSS.n11452 0.007925
R59725 DVSS.n16570 DVSS.n16551 0.00789286
R59726 DVSS.n16565 DVSS.n16352 0.00789286
R59727 DVSS.n17780 DVSS.n15926 0.00789286
R59728 DVSS.n15948 DVSS.n15947 0.00789286
R59729 DVSS.n17717 DVSS.n17682 0.00789286
R59730 DVSS.n17725 DVSS.n17680 0.00789286
R59731 DVSS.n18493 DVSS.n15153 0.00789286
R59732 DVSS.n15176 DVSS.n15175 0.00789286
R59733 DVSS.n21148 DVSS.n13691 0.00789286
R59734 DVSS.n13713 DVSS.n13712 0.00789286
R59735 DVSS.n21183 DVSS.n13642 0.00789286
R59736 DVSS.n13656 DVSS.n13640 0.00789286
R59737 DVSS.n22671 DVSS.n22670 0.00789286
R59738 DVSS.n731 DVSS.n714 0.00789286
R59739 DVSS.n13096 DVSS.n13095 0.00783696
R59740 DVSS.n22869 DVSS 0.00782857
R59741 DVSS.n16747 DVSS 0.00782857
R59742 DVSS.n16658 DVSS.n16271 0.00782857
R59743 DVSS.n16716 DVSS.n15662 0.00782857
R59744 DVSS DVSS.n15529 0.00782857
R59745 DVSS.n16119 DVSS.n16083 0.00782857
R59746 DVSS.n17603 DVSS.n16902 0.00782857
R59747 DVSS.n18259 DVSS 0.00782857
R59748 DVSS.n15334 DVSS.n15318 0.00782857
R59749 DVSS.n18313 DVSS.n15445 0.00782857
R59750 DVSS DVSS.n15123 0.00782857
R59751 DVSS.n18454 DVSS.n14884 0.00782857
R59752 DVSS.n15047 DVSS.n15026 0.00782857
R59753 DVSS.n20952 DVSS 0.00782857
R59754 DVSS.n20826 DVSS.n14486 0.00782857
R59755 DVSS.n14402 DVSS.n14386 0.00782857
R59756 DVSS.n21406 DVSS 0.00782857
R59757 DVSS.n21276 DVSS.n13544 0.00782857
R59758 DVSS.n13457 DVSS.n13445 0.00782857
R59759 DVSS.n22734 DVSS.n627 0.00782857
R59760 DVSS.n22812 DVSS.n526 0.00782857
R59761 DVSS.n17849 DVSS.n15852 0.00782394
R59762 DVSS.n17930 DVSS.n15759 0.00782394
R59763 DVSS.n16588 DVSS.n16348 0.00776429
R59764 DVSS.n17673 DVSS.n15958 0.00776429
R59765 DVSS.n17771 DVSS.n17706 0.00776429
R59766 DVSS.n15214 DVSS.n15209 0.00776429
R59767 DVSS.n20757 DVSS.n13727 0.00776429
R59768 DVSS.n21206 DVSS.n21205 0.00776429
R59769 DVSS.n22651 DVSS.n718 0.00776429
R59770 DVSS.n18014 DVSS.n15553 0.00775352
R59771 DVSS.n8989 DVSS.n2934 0.00774832
R59772 DVSS.n13348 DVSS.n10767 0.00774832
R59773 DVSS.n8991 DVSS.n8990 0.00774832
R59774 DVSS.n13347 DVSS.n10769 0.00774832
R59775 DVSS.n16679 DVSS.n16276 0.0077
R59776 DVSS.n16785 DVSS.n15666 0.0077
R59777 DVSS.n16106 DVSS.n16086 0.0077
R59778 DVSS.n17586 DVSS.n16906 0.0077
R59779 DVSS.n15350 DVSS.n15323 0.0077
R59780 DVSS.n18296 DVSS.n15449 0.0077
R59781 DVSS.n14915 DVSS.n14887 0.0077
R59782 DVSS.n15038 DVSS.n15031 0.0077
R59783 DVSS.n20847 DVSS.n14491 0.0077
R59784 DVSS.n20920 DVSS.n14391 0.0077
R59785 DVSS.n21297 DVSS.n13554 0.0077
R59786 DVSS.n21370 DVSS.n13450 0.0077
R59787 DVSS.n22755 DVSS.n632 0.0077
R59788 DVSS.n22828 DVSS.n531 0.0077
R59789 DVSS.n17946 DVSS.n15738 0.0076831
R59790 DVSS.n18046 DVSS.n15708 0.0076831
R59791 DVSS.n16742 DVSS.n15592 0.00763571
R59792 DVSS.n18180 DVSS.n15496 0.00763571
R59793 DVSS.n18254 DVSS.n18222 0.00763571
R59794 DVSS.n19933 DVSS.n15106 0.00763571
R59795 DVSS.n14342 DVSS.n14341 0.00763571
R59796 DVSS.n13400 DVSS.n13398 0.00763571
R59797 DVSS.n22875 DVSS.n470 0.00763571
R59798 DVSS.n16635 DVSS.n16306 0.00757143
R59799 DVSS.n16821 DVSS.n16154 0.00757143
R59800 DVSS.n16061 DVSS.n16015 0.00757143
R59801 DVSS.n16879 DVSS.n16838 0.00757143
R59802 DVSS.n18360 DVSS.n15240 0.00757143
R59803 DVSS.n15423 DVSS.n15382 0.00757143
R59804 DVSS.n18434 DVSS.n18432 0.00757143
R59805 DVSS.n14985 DVSS.n14946 0.00757143
R59806 DVSS.n20801 DVSS.n20722 0.00757143
R59807 DVSS.n14445 DVSS.n14427 0.00757143
R59808 DVSS.n21253 DVSS.n13584 0.00757143
R59809 DVSS.n13502 DVSS.n13483 0.00757143
R59810 DVSS.n22711 DVSS.n673 0.00757143
R59811 DVSS.n582 DVSS.n567 0.00757143
R59812 DVSS.n17895 DVSS.n15818 0.00754225
R59813 DVSS.n15726 DVSS.n15700 0.00754225
R59814 DVSS.n8336 DVSS.n3843 0.00753759
R59815 DVSS.n12342 DVSS.n12341 0.00753759
R59816 DVSS.n16731 DVSS.n15594 0.00750714
R59817 DVSS.n18201 DVSS.n18197 0.00750714
R59818 DVSS.n18239 DVSS.n18237 0.00750714
R59819 DVSS.n19950 DVSS.n15118 0.00750714
R59820 DVSS.n20968 DVSS.n20963 0.00750714
R59821 DVSS.n21422 DVSS.n21417 0.00750714
R59822 DVSS.n22858 DVSS.n474 0.00750714
R59823 DVSS.n8975 DVSS.n8974 0.007475
R59824 DVSS.n13116 DVSS.n13115 0.007475
R59825 DVSS.n17810 DVSS.n15895 0.00747183
R59826 DVSS.n16618 DVSS.n16310 0.00744286
R59827 DVSS.n16698 DVSS.n16158 0.00744286
R59828 DVSS.n16038 DVSS.n16019 0.00744286
R59829 DVSS.n16863 DVSS.n16842 0.00744286
R59830 DVSS.n18377 DVSS.n15244 0.00744286
R59831 DVSS.n15407 DVSS.n15386 0.00744286
R59832 DVSS.n18408 DVSS.n18386 0.00744286
R59833 DVSS.n14969 DVSS.n14950 0.00744286
R59834 DVSS.n20784 DVSS.n20709 0.00744286
R59835 DVSS.n20867 DVSS.n14431 0.00744286
R59836 DVSS.n21236 DVSS.n13591 0.00744286
R59837 DVSS.n21317 DVSS.n13487 0.00744286
R59838 DVSS.n22694 DVSS.n677 0.00744286
R59839 DVSS.n22775 DVSS.n571 0.00744286
R59840 DVSS.n17383 DVSS.n17382 0.00744149
R59841 DVSS.n17424 DVSS.n16933 0.00744149
R59842 DVSS.n17380 DVSS.n17310 0.00744149
R59843 DVSS.n17522 DVSS.n17521 0.00744149
R59844 DVSS.n17481 DVSS.n17118 0.00744149
R59845 DVSS.n17433 DVSS.n16924 0.00744149
R59846 DVSS.n13363 DVSS.n13362 0.00740226
R59847 DVSS.n17879 DVSS.n15813 0.00740141
R59848 DVSS.n7808 DVSS.n4812 0.00737773
R59849 DVSS.n7809 DVSS.n4813 0.00737773
R59850 DVSS.n17801 DVSS.n15903 0.00733099
R59851 DVSS.n18935 DVSS.n18912 0.00732584
R59852 DVSS.n20056 DVSS.n20055 0.00732584
R59853 DVSS.n20160 DVSS.n20040 0.00732584
R59854 DVSS.n14624 DVSS.n14623 0.00732584
R59855 DVSS.n20272 DVSS.n20222 0.00732584
R59856 DVSS.n20641 DVSS.n14660 0.00732584
R59857 DVSS.n20369 DVSS.n14683 0.00732584
R59858 DVSS.n16607 DVSS.n16312 0.00731429
R59859 DVSS.n15993 DVSS.n15988 0.00731429
R59860 DVSS.n17745 DVSS.n15246 0.00731429
R59861 DVSS.n18481 DVSS.n15223 0.00731429
R59862 DVSS.n20773 DVSS.n20711 0.00731429
R59863 DVSS.n21225 DVSS.n13593 0.00731429
R59864 DVSS.n22683 DVSS.n679 0.00731429
R59865 DVSS.n7061 DVSS.n5530 0.0072651
R59866 DVSS.n7799 DVSS.n4819 0.0072651
R59867 DVSS.n7062 DVSS.n5529 0.0072651
R59868 DVSS.n7800 DVSS.n4820 0.0072651
R59869 DVSS.n17886 DVSS.n15804 0.00726056
R59870 DVSS.n15729 DVSS.n15695 0.00726056
R59871 DVSS.n17821 DVSS.n15908 0.00719014
R59872 DVSS.n16623 DVSS.n16308 0.00718571
R59873 DVSS.n16230 DVSS.n16156 0.00718571
R59874 DVSS.n16050 DVSS.n16017 0.00718571
R59875 DVSS.n16860 DVSS.n16840 0.00718571
R59876 DVSS.n18371 DVSS.n15242 0.00718571
R59877 DVSS.n15404 DVSS.n15384 0.00718571
R59878 DVSS.n18417 DVSS.n18384 0.00718571
R59879 DVSS.n14966 DVSS.n14948 0.00718571
R59880 DVSS.n20726 DVSS.n20707 0.00718571
R59881 DVSS.n20871 DVSS.n14429 0.00718571
R59882 DVSS.n21241 DVSS.n13586 0.00718571
R59883 DVSS.n21321 DVSS.n13485 0.00718571
R59884 DVSS.n22699 DVSS.n675 0.00718571
R59885 DVSS.n22779 DVSS.n569 0.00718571
R59886 DVSS.n17799 DVSS.n17798 0.00716667
R59887 DVSS.n17800 DVSS.n17799 0.00716667
R59888 DVSS.n17800 DVSS.n15913 0.00716667
R59889 DVSS.n17807 DVSS.n15913 0.00716667
R59890 DVSS.n17808 DVSS.n17807 0.00716667
R59891 DVSS.n17809 DVSS.n17808 0.00716667
R59892 DVSS.n17809 DVSS.n15910 0.00716667
R59893 DVSS.n17816 DVSS.n15910 0.00716667
R59894 DVSS.n17817 DVSS.n17816 0.00716667
R59895 DVSS.n17818 DVSS.n17817 0.00716667
R59896 DVSS.n17818 DVSS.n15876 0.00716667
R59897 DVSS.n17826 DVSS.n15876 0.00716667
R59898 DVSS.n17827 DVSS.n17826 0.00716667
R59899 DVSS.n17829 DVSS.n17827 0.00716667
R59900 DVSS.n17829 DVSS.n17828 0.00716667
R59901 DVSS.n17828 DVSS.n15872 0.00716667
R59902 DVSS.n17837 DVSS.n15872 0.00716667
R59903 DVSS.n17838 DVSS.n17837 0.00716667
R59904 DVSS.n17839 DVSS.n17838 0.00716667
R59905 DVSS.n17839 DVSS.n15869 0.00716667
R59906 DVSS.n17846 DVSS.n15869 0.00716667
R59907 DVSS.n17847 DVSS.n17846 0.00716667
R59908 DVSS.n17848 DVSS.n17847 0.00716667
R59909 DVSS.n17848 DVSS.n15866 0.00716667
R59910 DVSS.n17855 DVSS.n15866 0.00716667
R59911 DVSS.n17856 DVSS.n17855 0.00716667
R59912 DVSS.n17857 DVSS.n17856 0.00716667
R59913 DVSS.n17857 DVSS.n15834 0.00716667
R59914 DVSS.n17868 DVSS.n15834 0.00716667
R59915 DVSS.n17869 DVSS.n17868 0.00716667
R59916 DVSS.n17871 DVSS.n17869 0.00716667
R59917 DVSS.n17871 DVSS.n17870 0.00716667
R59918 DVSS.n17870 DVSS.n15831 0.00716667
R59919 DVSS.n15831 DVSS.n15829 0.00716667
R59920 DVSS.n17881 DVSS.n15829 0.00716667
R59921 DVSS.n17882 DVSS.n17881 0.00716667
R59922 DVSS.n17883 DVSS.n17882 0.00716667
R59923 DVSS.n17883 DVSS.n15826 0.00716667
R59924 DVSS.n17890 DVSS.n15826 0.00716667
R59925 DVSS.n17891 DVSS.n17890 0.00716667
R59926 DVSS.n17892 DVSS.n17891 0.00716667
R59927 DVSS.n17892 DVSS.n15823 0.00716667
R59928 DVSS.n17899 DVSS.n15823 0.00716667
R59929 DVSS.n17900 DVSS.n17899 0.00716667
R59930 DVSS.n17901 DVSS.n17900 0.00716667
R59931 DVSS.n17902 DVSS.n17901 0.00716667
R59932 DVSS.n17902 DVSS.n15783 0.00716667
R59933 DVSS.n17912 DVSS.n15783 0.00716667
R59934 DVSS.n17913 DVSS.n17912 0.00716667
R59935 DVSS.n17915 DVSS.n17913 0.00716667
R59936 DVSS.n17915 DVSS.n17914 0.00716667
R59937 DVSS.n17914 DVSS.n15779 0.00716667
R59938 DVSS.n17923 DVSS.n15779 0.00716667
R59939 DVSS.n17924 DVSS.n17923 0.00716667
R59940 DVSS.n17925 DVSS.n17924 0.00716667
R59941 DVSS.n17925 DVSS.n15776 0.00716667
R59942 DVSS.n17932 DVSS.n15776 0.00716667
R59943 DVSS.n17933 DVSS.n17932 0.00716667
R59944 DVSS.n17934 DVSS.n17933 0.00716667
R59945 DVSS.n17934 DVSS.n15773 0.00716667
R59946 DVSS.n17941 DVSS.n15773 0.00716667
R59947 DVSS.n17942 DVSS.n17941 0.00716667
R59948 DVSS.n17943 DVSS.n17942 0.00716667
R59949 DVSS.n17943 DVSS.n15736 0.00716667
R59950 DVSS.n17952 DVSS.n15736 0.00716667
R59951 DVSS.n17953 DVSS.n17952 0.00716667
R59952 DVSS.n17955 DVSS.n17953 0.00716667
R59953 DVSS.n17955 DVSS.n17954 0.00716667
R59954 DVSS.n17954 DVSS.n15733 0.00716667
R59955 DVSS.n15733 DVSS.n15731 0.00716667
R59956 DVSS.n17965 DVSS.n15731 0.00716667
R59957 DVSS.n17966 DVSS.n17965 0.00716667
R59958 DVSS.n17967 DVSS.n17966 0.00716667
R59959 DVSS.n17967 DVSS.n15728 0.00716667
R59960 DVSS.n17974 DVSS.n15728 0.00716667
R59961 DVSS.n17975 DVSS.n17974 0.00716667
R59962 DVSS.n17976 DVSS.n17975 0.00716667
R59963 DVSS.n17977 DVSS.n17976 0.00716667
R59964 DVSS.n17978 DVSS.n17977 0.00716667
R59965 DVSS.n17979 DVSS.n17978 0.00716667
R59966 DVSS.n17980 DVSS.n17979 0.00716667
R59967 DVSS.n17981 DVSS.n17980 0.00716667
R59968 DVSS.n17982 DVSS.n17981 0.00716667
R59969 DVSS.n17983 DVSS.n17982 0.00716667
R59970 DVSS.n17986 DVSS.n17983 0.00716667
R59971 DVSS.n17987 DVSS.n17986 0.00716667
R59972 DVSS.n17988 DVSS.n17987 0.00716667
R59973 DVSS.n17989 DVSS.n17988 0.00716667
R59974 DVSS.n17990 DVSS.n17989 0.00716667
R59975 DVSS.n17991 DVSS.n17990 0.00716667
R59976 DVSS.n17992 DVSS.n17991 0.00716667
R59977 DVSS.n17993 DVSS.n17992 0.00716667
R59978 DVSS.n17994 DVSS.n17993 0.00716667
R59979 DVSS.n17995 DVSS.n17994 0.00716667
R59980 DVSS.n17996 DVSS.n17995 0.00716667
R59981 DVSS.n17997 DVSS.n17996 0.00716667
R59982 DVSS.n17998 DVSS.n17997 0.00716667
R59983 DVSS.n18000 DVSS.n17999 0.00716667
R59984 DVSS.n16753 DVSS.n15596 0.00712143
R59985 DVSS.n18191 DVSS.n15494 0.00712143
R59986 DVSS.n18265 DVSS.n18220 0.00712143
R59987 DVSS.n19944 DVSS.n15104 0.00712143
R59988 DVSS.n20944 DVSS.n14339 0.00712143
R59989 DVSS.n21398 DVSS.n13396 0.00712143
R59990 DVSS.n485 DVSS.n472 0.00712143
R59991 DVSS.n17905 DVSS.n15800 0.00711972
R59992 DVSS.n18038 DVSS.n15691 0.00711972
R59993 DVSS.n16815 DVSS.n16179 0.00705714
R59994 DVSS.n18079 DVSS.n15673 0.00705714
R59995 DVSS.n16883 DVSS.n16832 0.00705714
R59996 DVSS.n17575 DVSS.n16907 0.00705714
R59997 DVSS.n15427 DVSS.n15377 0.00705714
R59998 DVSS.n18285 DVSS.n15450 0.00705714
R59999 DVSS.n14995 DVSS.n14944 0.00705714
R60000 DVSS.n19970 DVSS.n19969 0.00705714
R60001 DVSS.n20887 DVSS.n14410 0.00705714
R60002 DVSS.n20930 DVSS.n14357 0.00705714
R60003 DVSS.n21337 DVSS.n13465 0.00705714
R60004 DVSS.n21384 DVSS.n13415 0.00705714
R60005 DVSS.n22795 DVSS.n547 0.00705714
R60006 DVSS.n22840 DVSS.n22839 0.00705714
R60007 DVSS.n21175 DVSS.n21174 0.00703846
R60008 DVSS.n6674 DVSS.n6234 0.007025
R60009 DVSS.n7075 DVSS.n7073 0.007025
R60010 DVSS.n10122 DVSS.n2367 0.00699624
R60011 DVSS.n10170 DVSS.n2024 0.00699624
R60012 DVSS.n9464 DVSS.n2727 0.00698472
R60013 DVSS.n11450 DVSS.n11199 0.00698472
R60014 DVSS.n9463 DVSS.n2726 0.00698472
R60015 DVSS.n13334 DVSS.n13333 0.00698472
R60016 DVSS.n17999 DVSS 0.00697887
R60017 DVSS.n17860 DVSS.n17859 0.00697887
R60018 DVSS.n17939 DVSS.n15768 0.00697887
R60019 DVSS.n16669 DVSS.n16273 0.00692857
R60020 DVSS.n16789 DVSS.n15664 0.00692857
R60021 DVSS.n16104 DVSS.n16085 0.00692857
R60022 DVSS.n17552 DVSS.n16904 0.00692857
R60023 DVSS.n15329 DVSS.n15320 0.00692857
R60024 DVSS.n15472 DVSS.n15447 0.00692857
R60025 DVSS.n14913 DVSS.n14886 0.00692857
R60026 DVSS.n15058 DVSS.n15028 0.00692857
R60027 DVSS.n20837 DVSS.n14488 0.00692857
R60028 DVSS.n20916 DVSS.n14388 0.00692857
R60029 DVSS.n21287 DVSS.n13546 0.00692857
R60030 DVSS.n21366 DVSS.n13447 0.00692857
R60031 DVSS.n22745 DVSS.n629 0.00692857
R60032 DVSS.n535 DVSS.n528 0.00692857
R60033 DVSS.n18020 DVSS.n15560 0.00690845
R60034 DVSS.n16584 DVSS.n16350 0.00686429
R60035 DVSS.n15979 DVSS.n15945 0.00686429
R60036 DVSS.n17736 DVSS.n17678 0.00686429
R60037 DVSS.n15203 DVSS.n15173 0.00686429
R60038 DVSS.n20753 DVSS.n13710 0.00686429
R60039 DVSS.n21197 DVSS.n13638 0.00686429
R60040 DVSS.n22655 DVSS.n716 0.00686429
R60041 DVSS.n19910 DVSS.n13672 0.00684146
R60042 DVSS.n17842 DVSS.n15859 0.00683803
R60043 DVSS.n15777 DVSS.n15763 0.00683803
R60044 DVSS.n18967 DVSS.n18877 0.00682022
R60045 DVSS.n20119 DVSS.n20057 0.00682022
R60046 DVSS.n20155 DVSS.n20153 0.00682022
R60047 DVSS.n20245 DVSS.n20218 0.00682022
R60048 DVSS.n20301 DVSS.n20300 0.00682022
R60049 DVSS.n20408 DVSS.n14688 0.00682022
R60050 DVSS.n16653 DVSS.n16268 0.0068
R60051 DVSS.n16115 DVSS.n16082 0.0068
R60052 DVSS.n18346 DVSS.n15291 0.0068
R60053 DVSS.n18439 DVSS.n14883 0.0068
R60054 DVSS.n20821 DVSS.n14483 0.0068
R60055 DVSS.n21271 DVSS.n13541 0.0068
R60056 DVSS.n22729 DVSS.n624 0.0068
R60057 DVSS.n8335 DVSS.n8334 0.00678188
R60058 DVSS.n12339 DVSS.n12002 0.00678188
R60059 DVSS.n8338 DVSS.n8337 0.00678188
R60060 DVSS.n12340 DVSS.n12001 0.00678188
R60061 DVSS.n19539 DVSS.n606 0.00677805
R60062 DVSS.n19544 DVSS.n561 0.00677805
R60063 DVSS.n19547 DVSS.n668 0.00677805
R60064 DVSS.n19543 DVSS.n506 0.00677805
R60065 DVSS.n16575 DVSS.n16554 0.00673571
R60066 DVSS.n15970 DVSS.n15950 0.00673571
R60067 DVSS.n17727 DVSS.n17685 0.00673571
R60068 DVSS.n15194 DVSS.n15178 0.00673571
R60069 DVSS.n20744 DVSS.n13715 0.00673571
R60070 DVSS.n21188 DVSS.n13645 0.00673571
R60071 DVSS.n22664 DVSS.n726 0.00673571
R60072 DVSS.n17835 DVSS.n15858 0.00669718
R60073 DVSS.n16660 DVSS.n16259 0.00667143
R60074 DVSS.n16798 DVSS.n15658 0.00667143
R60075 DVSS.n16109 DVSS.n16078 0.00667143
R60076 DVSS.n17548 DVSS.n17545 0.00667143
R60077 DVSS.n15332 DVSS.n15313 0.00667143
R60078 DVSS.n15468 DVSS.n15465 0.00667143
R60079 DVSS.n18452 DVSS.n14879 0.00667143
R60080 DVSS.n15049 DVSS.n15022 0.00667143
R60081 DVSS.n20828 DVSS.n14479 0.00667143
R60082 DVSS.n20907 DVSS.n14381 0.00667143
R60083 DVSS.n21278 DVSS.n13537 0.00667143
R60084 DVSS.n21357 DVSS.n13440 0.00667143
R60085 DVSS.n22736 DVSS.n619 0.00667143
R60086 DVSS.n538 DVSS.n520 0.00667143
R60087 DVSS.n17985 DVSS.n15561 0.00662676
R60088 DVSS.n16595 DVSS.n16559 0.00660714
R60089 DVSS.n17672 DVSS.n15954 0.00660714
R60090 DVSS.n17770 DVSS.n17690 0.00660714
R60091 DVSS.n15215 DVSS.n15183 0.00660714
R60092 DVSS.n20737 DVSS.n13719 0.00660714
R60093 DVSS.n21213 DVSS.n13650 0.00660714
R60094 DVSS.n22644 DVSS.n721 0.00660714
R60095 DVSS.n22603 DVSS.n745 0.00659375
R60096 DVSS.n22918 DVSS.n441 0.00659375
R60097 DVSS.n8977 DVSS.n3053 0.0065917
R60098 DVSS.n11992 DVSS.n11633 0.0065917
R60099 DVSS.n8976 DVSS.n3054 0.0065917
R60100 DVSS.n11990 DVSS.n11635 0.0065917
R60101 DVSS.n22668 DVSS.n22667 0.00658571
R60102 DVSS.n22667 DVSS.n22666 0.00658571
R60103 DVSS.n22666 DVSS.n22640 0.00658571
R60104 DVSS.n22659 DVSS.n22640 0.00658571
R60105 DVSS.n22659 DVSS.n22658 0.00658571
R60106 DVSS.n22658 DVSS.n22657 0.00658571
R60107 DVSS.n22657 DVSS.n22643 0.00658571
R60108 DVSS.n22650 DVSS.n22643 0.00658571
R60109 DVSS.n22650 DVSS.n22649 0.00658571
R60110 DVSS.n22649 DVSS.n22648 0.00658571
R60111 DVSS.n22648 DVSS.n699 0.00658571
R60112 DVSS.n22676 DVSS.n699 0.00658571
R60113 DVSS.n22677 DVSS.n22676 0.00658571
R60114 DVSS.n22679 DVSS.n22677 0.00658571
R60115 DVSS.n22679 DVSS.n22678 0.00658571
R60116 DVSS.n22678 DVSS.n695 0.00658571
R60117 DVSS.n22687 DVSS.n695 0.00658571
R60118 DVSS.n22688 DVSS.n22687 0.00658571
R60119 DVSS.n22689 DVSS.n22688 0.00658571
R60120 DVSS.n22689 DVSS.n692 0.00658571
R60121 DVSS.n22696 DVSS.n692 0.00658571
R60122 DVSS.n22697 DVSS.n22696 0.00658571
R60123 DVSS.n22698 DVSS.n22697 0.00658571
R60124 DVSS.n22698 DVSS.n689 0.00658571
R60125 DVSS.n22705 DVSS.n689 0.00658571
R60126 DVSS.n22706 DVSS.n22705 0.00658571
R60127 DVSS.n22707 DVSS.n22706 0.00658571
R60128 DVSS.n22707 DVSS.n646 0.00658571
R60129 DVSS.n22718 DVSS.n646 0.00658571
R60130 DVSS.n22719 DVSS.n22718 0.00658571
R60131 DVSS.n22721 DVSS.n22719 0.00658571
R60132 DVSS.n22721 DVSS.n22720 0.00658571
R60133 DVSS.n22720 DVSS.n643 0.00658571
R60134 DVSS.n643 DVSS.n641 0.00658571
R60135 DVSS.n22731 DVSS.n641 0.00658571
R60136 DVSS.n22732 DVSS.n22731 0.00658571
R60137 DVSS.n22733 DVSS.n22732 0.00658571
R60138 DVSS.n22733 DVSS.n638 0.00658571
R60139 DVSS.n22740 DVSS.n638 0.00658571
R60140 DVSS.n22741 DVSS.n22740 0.00658571
R60141 DVSS.n22742 DVSS.n22741 0.00658571
R60142 DVSS.n22742 DVSS.n635 0.00658571
R60143 DVSS.n22749 DVSS.n635 0.00658571
R60144 DVSS.n22750 DVSS.n22749 0.00658571
R60145 DVSS.n22752 DVSS.n22750 0.00658571
R60146 DVSS.n22752 DVSS.n22751 0.00658571
R60147 DVSS.n22751 DVSS.n594 0.00658571
R60148 DVSS.n22761 DVSS.n594 0.00658571
R60149 DVSS.n22762 DVSS.n22761 0.00658571
R60150 DVSS.n22764 DVSS.n22762 0.00658571
R60151 DVSS.n22764 DVSS.n22763 0.00658571
R60152 DVSS.n22763 DVSS.n590 0.00658571
R60153 DVSS.n22772 DVSS.n590 0.00658571
R60154 DVSS.n22773 DVSS.n22772 0.00658571
R60155 DVSS.n22774 DVSS.n22773 0.00658571
R60156 DVSS.n22774 DVSS.n587 0.00658571
R60157 DVSS.n22781 DVSS.n587 0.00658571
R60158 DVSS.n22782 DVSS.n22781 0.00658571
R60159 DVSS.n22783 DVSS.n22782 0.00658571
R60160 DVSS.n22783 DVSS.n584 0.00658571
R60161 DVSS.n22790 DVSS.n584 0.00658571
R60162 DVSS.n22791 DVSS.n22790 0.00658571
R60163 DVSS.n22792 DVSS.n22791 0.00658571
R60164 DVSS.n22792 DVSS.n545 0.00658571
R60165 DVSS.n22801 DVSS.n545 0.00658571
R60166 DVSS.n22802 DVSS.n22801 0.00658571
R60167 DVSS.n22804 DVSS.n22802 0.00658571
R60168 DVSS.n22804 DVSS.n22803 0.00658571
R60169 DVSS.n22803 DVSS.n542 0.00658571
R60170 DVSS.n542 DVSS.n540 0.00658571
R60171 DVSS.n22814 DVSS.n540 0.00658571
R60172 DVSS.n22815 DVSS.n22814 0.00658571
R60173 DVSS.n22816 DVSS.n22815 0.00658571
R60174 DVSS.n22816 DVSS.n537 0.00658571
R60175 DVSS.n22823 DVSS.n537 0.00658571
R60176 DVSS.n22824 DVSS.n22823 0.00658571
R60177 DVSS.n22825 DVSS.n22824 0.00658571
R60178 DVSS.n22825 DVSS.n534 0.00658571
R60179 DVSS.n22832 DVSS.n534 0.00658571
R60180 DVSS.n22833 DVSS.n22832 0.00658571
R60181 DVSS.n22834 DVSS.n22833 0.00658571
R60182 DVSS.n22834 DVSS.n494 0.00658571
R60183 DVSS.n22842 DVSS.n494 0.00658571
R60184 DVSS.n22843 DVSS.n22842 0.00658571
R60185 DVSS.n22845 DVSS.n22843 0.00658571
R60186 DVSS.n22845 DVSS.n22844 0.00658571
R60187 DVSS.n22844 DVSS.n490 0.00658571
R60188 DVSS.n22853 DVSS.n490 0.00658571
R60189 DVSS.n22854 DVSS.n22853 0.00658571
R60190 DVSS.n22855 DVSS.n22854 0.00658571
R60191 DVSS.n22855 DVSS.n487 0.00658571
R60192 DVSS.n22862 DVSS.n487 0.00658571
R60193 DVSS.n22863 DVSS.n22862 0.00658571
R60194 DVSS.n22864 DVSS.n22863 0.00658571
R60195 DVSS.n22864 DVSS.n484 0.00658571
R60196 DVSS.n22870 DVSS.n484 0.00658571
R60197 DVSS.n22871 DVSS.n22870 0.00658571
R60198 DVSS.n22882 DVSS.n456 0.00658571
R60199 DVSS.n16573 DVSS.n16572 0.00658571
R60200 DVSS.n16574 DVSS.n16573 0.00658571
R60201 DVSS.n16574 DVSS.n16564 0.00658571
R60202 DVSS.n16581 DVSS.n16564 0.00658571
R60203 DVSS.n16582 DVSS.n16581 0.00658571
R60204 DVSS.n16583 DVSS.n16582 0.00658571
R60205 DVSS.n16583 DVSS.n16561 0.00658571
R60206 DVSS.n16590 DVSS.n16561 0.00658571
R60207 DVSS.n16591 DVSS.n16590 0.00658571
R60208 DVSS.n16592 DVSS.n16591 0.00658571
R60209 DVSS.n16592 DVSS.n16332 0.00658571
R60210 DVSS.n16600 DVSS.n16332 0.00658571
R60211 DVSS.n16601 DVSS.n16600 0.00658571
R60212 DVSS.n16603 DVSS.n16601 0.00658571
R60213 DVSS.n16603 DVSS.n16602 0.00658571
R60214 DVSS.n16602 DVSS.n16328 0.00658571
R60215 DVSS.n16611 DVSS.n16328 0.00658571
R60216 DVSS.n16612 DVSS.n16611 0.00658571
R60217 DVSS.n16613 DVSS.n16612 0.00658571
R60218 DVSS.n16613 DVSS.n16325 0.00658571
R60219 DVSS.n16620 DVSS.n16325 0.00658571
R60220 DVSS.n16621 DVSS.n16620 0.00658571
R60221 DVSS.n16622 DVSS.n16621 0.00658571
R60222 DVSS.n16622 DVSS.n16322 0.00658571
R60223 DVSS.n16629 DVSS.n16322 0.00658571
R60224 DVSS.n16630 DVSS.n16629 0.00658571
R60225 DVSS.n16631 DVSS.n16630 0.00658571
R60226 DVSS.n16631 DVSS.n16290 0.00658571
R60227 DVSS.n16642 DVSS.n16290 0.00658571
R60228 DVSS.n16643 DVSS.n16642 0.00658571
R60229 DVSS.n16645 DVSS.n16643 0.00658571
R60230 DVSS.n16645 DVSS.n16644 0.00658571
R60231 DVSS.n16644 DVSS.n16287 0.00658571
R60232 DVSS.n16287 DVSS.n16285 0.00658571
R60233 DVSS.n16655 DVSS.n16285 0.00658571
R60234 DVSS.n16656 DVSS.n16655 0.00658571
R60235 DVSS.n16657 DVSS.n16656 0.00658571
R60236 DVSS.n16657 DVSS.n16282 0.00658571
R60237 DVSS.n16664 DVSS.n16282 0.00658571
R60238 DVSS.n16665 DVSS.n16664 0.00658571
R60239 DVSS.n16666 DVSS.n16665 0.00658571
R60240 DVSS.n16666 DVSS.n16279 0.00658571
R60241 DVSS.n16673 DVSS.n16279 0.00658571
R60242 DVSS.n16674 DVSS.n16673 0.00658571
R60243 DVSS.n16676 DVSS.n16674 0.00658571
R60244 DVSS.n16676 DVSS.n16675 0.00658571
R60245 DVSS.n16675 DVSS.n16239 0.00658571
R60246 DVSS.n16685 DVSS.n16239 0.00658571
R60247 DVSS.n16686 DVSS.n16685 0.00658571
R60248 DVSS.n16687 DVSS.n16686 0.00658571
R60249 DVSS.n16687 DVSS.n16235 0.00658571
R60250 DVSS.n16693 DVSS.n16235 0.00658571
R60251 DVSS.n16694 DVSS.n16693 0.00658571
R60252 DVSS.n16695 DVSS.n16694 0.00658571
R60253 DVSS.n16695 DVSS.n16232 0.00658571
R60254 DVSS.n16702 DVSS.n16232 0.00658571
R60255 DVSS.n16703 DVSS.n16702 0.00658571
R60256 DVSS.n16704 DVSS.n16703 0.00658571
R60257 DVSS.n16704 DVSS.n16229 0.00658571
R60258 DVSS.n16711 DVSS.n16229 0.00658571
R60259 DVSS.n16712 DVSS.n16711 0.00658571
R60260 DVSS.n16819 DVSS.n16712 0.00658571
R60261 DVSS.n16819 DVSS.n16818 0.00658571
R60262 DVSS.n16818 DVSS.n16817 0.00658571
R60263 DVSS.n16817 DVSS.n16713 0.00658571
R60264 DVSS.n16812 DVSS.n16713 0.00658571
R60265 DVSS.n16812 DVSS.n16811 0.00658571
R60266 DVSS.n16811 DVSS.n16810 0.00658571
R60267 DVSS.n16810 DVSS.n16715 0.00658571
R60268 DVSS.n16802 DVSS.n16715 0.00658571
R60269 DVSS.n16802 DVSS.n16801 0.00658571
R60270 DVSS.n16801 DVSS.n16800 0.00658571
R60271 DVSS.n16800 DVSS.n16718 0.00658571
R60272 DVSS.n16793 DVSS.n16718 0.00658571
R60273 DVSS.n16793 DVSS.n16792 0.00658571
R60274 DVSS.n16792 DVSS.n16791 0.00658571
R60275 DVSS.n16791 DVSS.n16721 0.00658571
R60276 DVSS.n16784 DVSS.n16721 0.00658571
R60277 DVSS.n16784 DVSS.n16783 0.00658571
R60278 DVSS.n16783 DVSS.n16782 0.00658571
R60279 DVSS.n16782 DVSS.n16724 0.00658571
R60280 DVSS.n16776 DVSS.n16724 0.00658571
R60281 DVSS.n16776 DVSS.n16775 0.00658571
R60282 DVSS.n16775 DVSS.n16774 0.00658571
R60283 DVSS.n16774 DVSS.n16726 0.00658571
R60284 DVSS.n16768 DVSS.n16726 0.00658571
R60285 DVSS.n16768 DVSS.n16767 0.00658571
R60286 DVSS.n16767 DVSS.n16766 0.00658571
R60287 DVSS.n16766 DVSS.n16730 0.00658571
R60288 DVSS.n16759 DVSS.n16730 0.00658571
R60289 DVSS.n16759 DVSS.n16758 0.00658571
R60290 DVSS.n16758 DVSS.n16757 0.00658571
R60291 DVSS.n16757 DVSS.n16733 0.00658571
R60292 DVSS.n16750 DVSS.n16733 0.00658571
R60293 DVSS.n16750 DVSS.n16749 0.00658571
R60294 DVSS.n16749 DVSS.n16748 0.00658571
R60295 DVSS.n16748 DVSS.n16736 0.00658571
R60296 DVSS.n16741 DVSS.n16740 0.00658571
R60297 DVSS.n17782 DVSS.n15924 0.00658571
R60298 DVSS.n15969 DVSS.n15924 0.00658571
R60299 DVSS.n15974 DVSS.n15969 0.00658571
R60300 DVSS.n15975 DVSS.n15974 0.00658571
R60301 DVSS.n15976 DVSS.n15975 0.00658571
R60302 DVSS.n15976 DVSS.n15966 0.00658571
R60303 DVSS.n15983 DVSS.n15966 0.00658571
R60304 DVSS.n15984 DVSS.n15983 0.00658571
R60305 DVSS.n17670 DVSS.n15984 0.00658571
R60306 DVSS.n17670 DVSS.n17669 0.00658571
R60307 DVSS.n17669 DVSS.n17668 0.00658571
R60308 DVSS.n17668 DVSS.n15985 0.00658571
R60309 DVSS.n15987 DVSS.n15985 0.00658571
R60310 DVSS.n15990 DVSS.n15987 0.00658571
R60311 DVSS.n17660 DVSS.n15990 0.00658571
R60312 DVSS.n17660 DVSS.n17659 0.00658571
R60313 DVSS.n17659 DVSS.n17658 0.00658571
R60314 DVSS.n17658 DVSS.n15991 0.00658571
R60315 DVSS.n16040 DVSS.n15991 0.00658571
R60316 DVSS.n16045 DVSS.n16040 0.00658571
R60317 DVSS.n16046 DVSS.n16045 0.00658571
R60318 DVSS.n16047 DVSS.n16046 0.00658571
R60319 DVSS.n16047 DVSS.n16037 0.00658571
R60320 DVSS.n16054 DVSS.n16037 0.00658571
R60321 DVSS.n16055 DVSS.n16054 0.00658571
R60322 DVSS.n16056 DVSS.n16055 0.00658571
R60323 DVSS.n16056 DVSS.n16034 0.00658571
R60324 DVSS.n16063 DVSS.n16034 0.00658571
R60325 DVSS.n16064 DVSS.n16063 0.00658571
R60326 DVSS.n17650 DVSS.n16064 0.00658571
R60327 DVSS.n17650 DVSS.n17649 0.00658571
R60328 DVSS.n17649 DVSS.n17648 0.00658571
R60329 DVSS.n17648 DVSS.n16065 0.00658571
R60330 DVSS.n16113 DVSS.n16065 0.00658571
R60331 DVSS.n16114 DVSS.n16113 0.00658571
R60332 DVSS.n16114 DVSS.n16111 0.00658571
R60333 DVSS.n16121 DVSS.n16111 0.00658571
R60334 DVSS.n16122 DVSS.n16121 0.00658571
R60335 DVSS.n16123 DVSS.n16122 0.00658571
R60336 DVSS.n16123 DVSS.n16108 0.00658571
R60337 DVSS.n16130 DVSS.n16108 0.00658571
R60338 DVSS.n16131 DVSS.n16130 0.00658571
R60339 DVSS.n17637 DVSS.n16131 0.00658571
R60340 DVSS.n17637 DVSS.n17636 0.00658571
R60341 DVSS.n17636 DVSS.n17635 0.00658571
R60342 DVSS.n17635 DVSS.n16132 0.00658571
R60343 DVSS.n17630 DVSS.n16132 0.00658571
R60344 DVSS.n17630 DVSS.n17629 0.00658571
R60345 DVSS.n17629 DVSS.n17628 0.00658571
R60346 DVSS.n17628 DVSS.n16134 0.00658571
R60347 DVSS.n17622 DVSS.n16134 0.00658571
R60348 DVSS.n17622 DVSS.n17621 0.00658571
R60349 DVSS.n17621 DVSS.n17620 0.00658571
R60350 DVSS.n17620 DVSS.n16139 0.00658571
R60351 DVSS.n16862 DVSS.n16139 0.00658571
R60352 DVSS.n16867 DVSS.n16862 0.00658571
R60353 DVSS.n16868 DVSS.n16867 0.00658571
R60354 DVSS.n16869 DVSS.n16868 0.00658571
R60355 DVSS.n16869 DVSS.n16859 0.00658571
R60356 DVSS.n16876 DVSS.n16859 0.00658571
R60357 DVSS.n16877 DVSS.n16876 0.00658571
R60358 DVSS.n16878 DVSS.n16877 0.00658571
R60359 DVSS.n16878 DVSS.n16856 0.00658571
R60360 DVSS.n16885 DVSS.n16856 0.00658571
R60361 DVSS.n16886 DVSS.n16885 0.00658571
R60362 DVSS.n17612 DVSS.n16886 0.00658571
R60363 DVSS.n17612 DVSS.n17611 0.00658571
R60364 DVSS.n17611 DVSS.n17610 0.00658571
R60365 DVSS.n17610 DVSS.n16887 0.00658571
R60366 DVSS.n17550 DVSS.n16887 0.00658571
R60367 DVSS.n17601 DVSS.n17550 0.00658571
R60368 DVSS.n17601 DVSS.n17600 0.00658571
R60369 DVSS.n17600 DVSS.n17599 0.00658571
R60370 DVSS.n17599 DVSS.n17551 0.00658571
R60371 DVSS.n17592 DVSS.n17551 0.00658571
R60372 DVSS.n17592 DVSS.n17591 0.00658571
R60373 DVSS.n17591 DVSS.n17590 0.00658571
R60374 DVSS.n17590 DVSS.n17554 0.00658571
R60375 DVSS.n17583 DVSS.n17554 0.00658571
R60376 DVSS.n17583 DVSS.n17582 0.00658571
R60377 DVSS.n17582 DVSS.n17581 0.00658571
R60378 DVSS.n17581 DVSS.n17557 0.00658571
R60379 DVSS.n17559 DVSS.n17557 0.00658571
R60380 DVSS.n17562 DVSS.n17559 0.00658571
R60381 DVSS.n17571 DVSS.n17562 0.00658571
R60382 DVSS.n17571 DVSS.n17570 0.00658571
R60383 DVSS.n17570 DVSS.n17569 0.00658571
R60384 DVSS.n17569 DVSS.n17563 0.00658571
R60385 DVSS.n17564 DVSS.n17563 0.00658571
R60386 DVSS.n17564 DVSS.n15526 0.00658571
R60387 DVSS.n18195 DVSS.n15526 0.00658571
R60388 DVSS.n18195 DVSS.n18194 0.00658571
R60389 DVSS.n18194 DVSS.n18193 0.00658571
R60390 DVSS.n18193 DVSS.n15527 0.00658571
R60391 DVSS.n18186 DVSS.n15527 0.00658571
R60392 DVSS.n18186 DVSS.n18185 0.00658571
R60393 DVSS.n18185 DVSS.n18184 0.00658571
R60394 DVSS.n18179 DVSS.n18178 0.00658571
R60395 DVSS.n17724 DVSS.n17723 0.00658571
R60396 DVSS.n17724 DVSS.n17716 0.00658571
R60397 DVSS.n17731 DVSS.n17716 0.00658571
R60398 DVSS.n17732 DVSS.n17731 0.00658571
R60399 DVSS.n17733 DVSS.n17732 0.00658571
R60400 DVSS.n17733 DVSS.n17713 0.00658571
R60401 DVSS.n17740 DVSS.n17713 0.00658571
R60402 DVSS.n17741 DVSS.n17740 0.00658571
R60403 DVSS.n17768 DVSS.n17741 0.00658571
R60404 DVSS.n17768 DVSS.n17767 0.00658571
R60405 DVSS.n17767 DVSS.n17766 0.00658571
R60406 DVSS.n17766 DVSS.n17742 0.00658571
R60407 DVSS.n17744 DVSS.n17742 0.00658571
R60408 DVSS.n17747 DVSS.n17744 0.00658571
R60409 DVSS.n17758 DVSS.n17747 0.00658571
R60410 DVSS.n17758 DVSS.n17757 0.00658571
R60411 DVSS.n17757 DVSS.n17756 0.00658571
R60412 DVSS.n17756 DVSS.n17748 0.00658571
R60413 DVSS.n17749 DVSS.n17748 0.00658571
R60414 DVSS.n17749 DVSS.n15278 0.00658571
R60415 DVSS.n18375 DVSS.n15278 0.00658571
R60416 DVSS.n18375 DVSS.n18374 0.00658571
R60417 DVSS.n18374 DVSS.n18373 0.00658571
R60418 DVSS.n18373 DVSS.n15279 0.00658571
R60419 DVSS.n18366 DVSS.n15279 0.00658571
R60420 DVSS.n18366 DVSS.n18365 0.00658571
R60421 DVSS.n18365 DVSS.n18364 0.00658571
R60422 DVSS.n18364 DVSS.n15282 0.00658571
R60423 DVSS.n18358 DVSS.n15282 0.00658571
R60424 DVSS.n18358 DVSS.n18357 0.00658571
R60425 DVSS.n18357 DVSS.n18356 0.00658571
R60426 DVSS.n18356 DVSS.n15284 0.00658571
R60427 DVSS.n18350 DVSS.n15284 0.00658571
R60428 DVSS.n18350 DVSS.n18349 0.00658571
R60429 DVSS.n18349 DVSS.n18348 0.00658571
R60430 DVSS.n18348 DVSS.n15288 0.00658571
R60431 DVSS.n15336 DVSS.n15288 0.00658571
R60432 DVSS.n15337 DVSS.n15336 0.00658571
R60433 DVSS.n15338 DVSS.n15337 0.00658571
R60434 DVSS.n15338 DVSS.n15331 0.00658571
R60435 DVSS.n15345 DVSS.n15331 0.00658571
R60436 DVSS.n15346 DVSS.n15345 0.00658571
R60437 DVSS.n15347 DVSS.n15346 0.00658571
R60438 DVSS.n15347 DVSS.n15328 0.00658571
R60439 DVSS.n15354 DVSS.n15328 0.00658571
R60440 DVSS.n15355 DVSS.n15354 0.00658571
R60441 DVSS.n18340 DVSS.n15355 0.00658571
R60442 DVSS.n18340 DVSS.n18339 0.00658571
R60443 DVSS.n18339 DVSS.n18338 0.00658571
R60444 DVSS.n18338 DVSS.n15356 0.00658571
R60445 DVSS.n18332 DVSS.n15356 0.00658571
R60446 DVSS.n18332 DVSS.n18331 0.00658571
R60447 DVSS.n18331 DVSS.n18330 0.00658571
R60448 DVSS.n18330 DVSS.n15360 0.00658571
R60449 DVSS.n15406 DVSS.n15360 0.00658571
R60450 DVSS.n15411 DVSS.n15406 0.00658571
R60451 DVSS.n15412 DVSS.n15411 0.00658571
R60452 DVSS.n15413 DVSS.n15412 0.00658571
R60453 DVSS.n15413 DVSS.n15403 0.00658571
R60454 DVSS.n15420 DVSS.n15403 0.00658571
R60455 DVSS.n15421 DVSS.n15420 0.00658571
R60456 DVSS.n15422 DVSS.n15421 0.00658571
R60457 DVSS.n15422 DVSS.n15400 0.00658571
R60458 DVSS.n15429 DVSS.n15400 0.00658571
R60459 DVSS.n15430 DVSS.n15429 0.00658571
R60460 DVSS.n18322 DVSS.n15430 0.00658571
R60461 DVSS.n18322 DVSS.n18321 0.00658571
R60462 DVSS.n18321 DVSS.n18320 0.00658571
R60463 DVSS.n18320 DVSS.n15431 0.00658571
R60464 DVSS.n15470 DVSS.n15431 0.00658571
R60465 DVSS.n18311 DVSS.n15470 0.00658571
R60466 DVSS.n18311 DVSS.n18310 0.00658571
R60467 DVSS.n18310 DVSS.n18309 0.00658571
R60468 DVSS.n18309 DVSS.n15471 0.00658571
R60469 DVSS.n18302 DVSS.n15471 0.00658571
R60470 DVSS.n18302 DVSS.n18301 0.00658571
R60471 DVSS.n18301 DVSS.n18300 0.00658571
R60472 DVSS.n18300 DVSS.n15474 0.00658571
R60473 DVSS.n18293 DVSS.n15474 0.00658571
R60474 DVSS.n18293 DVSS.n18292 0.00658571
R60475 DVSS.n18292 DVSS.n18291 0.00658571
R60476 DVSS.n18291 DVSS.n15477 0.00658571
R60477 DVSS.n15479 DVSS.n15477 0.00658571
R60478 DVSS.n15482 DVSS.n15479 0.00658571
R60479 DVSS.n18281 DVSS.n15482 0.00658571
R60480 DVSS.n18281 DVSS.n18280 0.00658571
R60481 DVSS.n18280 DVSS.n18279 0.00658571
R60482 DVSS.n18279 DVSS.n15483 0.00658571
R60483 DVSS.n18241 DVSS.n15483 0.00658571
R60484 DVSS.n18271 DVSS.n18241 0.00658571
R60485 DVSS.n18271 DVSS.n18270 0.00658571
R60486 DVSS.n18270 DVSS.n18269 0.00658571
R60487 DVSS.n18269 DVSS.n18242 0.00658571
R60488 DVSS.n18262 DVSS.n18242 0.00658571
R60489 DVSS.n18262 DVSS.n18261 0.00658571
R60490 DVSS.n18261 DVSS.n18260 0.00658571
R60491 DVSS.n18260 DVSS.n18245 0.00658571
R60492 DVSS.n18253 DVSS.n18252 0.00658571
R60493 DVSS.n18495 DVSS.n15151 0.00658571
R60494 DVSS.n15196 DVSS.n15151 0.00658571
R60495 DVSS.n15197 DVSS.n15196 0.00658571
R60496 DVSS.n15198 DVSS.n15197 0.00658571
R60497 DVSS.n15198 DVSS.n15191 0.00658571
R60498 DVSS.n15205 DVSS.n15191 0.00658571
R60499 DVSS.n15206 DVSS.n15205 0.00658571
R60500 DVSS.n15207 DVSS.n15206 0.00658571
R60501 DVSS.n15207 DVSS.n15188 0.00658571
R60502 DVSS.n15219 DVSS.n15188 0.00658571
R60503 DVSS.n15220 DVSS.n15219 0.00658571
R60504 DVSS.n18487 DVSS.n15220 0.00658571
R60505 DVSS.n18487 DVSS.n18486 0.00658571
R60506 DVSS.n18486 DVSS.n18485 0.00658571
R60507 DVSS.n18485 DVSS.n15221 0.00658571
R60508 DVSS.n18479 DVSS.n15221 0.00658571
R60509 DVSS.n18479 DVSS.n18478 0.00658571
R60510 DVSS.n18478 DVSS.n18477 0.00658571
R60511 DVSS.n18477 DVSS.n15225 0.00658571
R60512 DVSS.n18412 DVSS.n15225 0.00658571
R60513 DVSS.n18413 DVSS.n18412 0.00658571
R60514 DVSS.n18414 DVSS.n18413 0.00658571
R60515 DVSS.n18414 DVSS.n18407 0.00658571
R60516 DVSS.n18421 DVSS.n18407 0.00658571
R60517 DVSS.n18422 DVSS.n18421 0.00658571
R60518 DVSS.n18423 DVSS.n18422 0.00658571
R60519 DVSS.n18423 DVSS.n18404 0.00658571
R60520 DVSS.n18436 DVSS.n18404 0.00658571
R60521 DVSS.n18437 DVSS.n18436 0.00658571
R60522 DVSS.n18469 DVSS.n18437 0.00658571
R60523 DVSS.n18469 DVSS.n18468 0.00658571
R60524 DVSS.n18468 DVSS.n18467 0.00658571
R60525 DVSS.n18467 DVSS.n18438 0.00658571
R60526 DVSS.n18460 DVSS.n18438 0.00658571
R60527 DVSS.n18460 DVSS.n18459 0.00658571
R60528 DVSS.n18459 DVSS.n18458 0.00658571
R60529 DVSS.n18458 DVSS.n18441 0.00658571
R60530 DVSS.n18451 DVSS.n18441 0.00658571
R60531 DVSS.n18451 DVSS.n18450 0.00658571
R60532 DVSS.n18450 DVSS.n18449 0.00658571
R60533 DVSS.n18449 DVSS.n18444 0.00658571
R60534 DVSS.n18444 DVSS.n14917 0.00658571
R60535 DVSS.n20003 DVSS.n14917 0.00658571
R60536 DVSS.n20003 DVSS.n20002 0.00658571
R60537 DVSS.n20002 DVSS.n20001 0.00658571
R60538 DVSS.n20001 DVSS.n14918 0.00658571
R60539 DVSS.n19996 DVSS.n14918 0.00658571
R60540 DVSS.n19996 DVSS.n19995 0.00658571
R60541 DVSS.n19995 DVSS.n19994 0.00658571
R60542 DVSS.n19994 DVSS.n14920 0.00658571
R60543 DVSS.n19988 DVSS.n14920 0.00658571
R60544 DVSS.n19988 DVSS.n19987 0.00658571
R60545 DVSS.n19987 DVSS.n19986 0.00658571
R60546 DVSS.n19986 DVSS.n14925 0.00658571
R60547 DVSS.n14968 DVSS.n14925 0.00658571
R60548 DVSS.n14973 DVSS.n14968 0.00658571
R60549 DVSS.n14974 DVSS.n14973 0.00658571
R60550 DVSS.n14975 DVSS.n14974 0.00658571
R60551 DVSS.n14975 DVSS.n14965 0.00658571
R60552 DVSS.n14982 DVSS.n14965 0.00658571
R60553 DVSS.n14983 DVSS.n14982 0.00658571
R60554 DVSS.n14984 DVSS.n14983 0.00658571
R60555 DVSS.n14984 DVSS.n14962 0.00658571
R60556 DVSS.n14997 DVSS.n14962 0.00658571
R60557 DVSS.n14998 DVSS.n14997 0.00658571
R60558 DVSS.n19978 DVSS.n14998 0.00658571
R60559 DVSS.n19978 DVSS.n19977 0.00658571
R60560 DVSS.n19977 DVSS.n19976 0.00658571
R60561 DVSS.n19976 DVSS.n14999 0.00658571
R60562 DVSS.n15045 DVSS.n14999 0.00658571
R60563 DVSS.n15046 DVSS.n15045 0.00658571
R60564 DVSS.n15046 DVSS.n15043 0.00658571
R60565 DVSS.n15053 DVSS.n15043 0.00658571
R60566 DVSS.n15054 DVSS.n15053 0.00658571
R60567 DVSS.n15055 DVSS.n15054 0.00658571
R60568 DVSS.n15055 DVSS.n15040 0.00658571
R60569 DVSS.n15062 DVSS.n15040 0.00658571
R60570 DVSS.n15063 DVSS.n15062 0.00658571
R60571 DVSS.n15064 DVSS.n15063 0.00658571
R60572 DVSS.n15064 DVSS.n15037 0.00658571
R60573 DVSS.n15076 DVSS.n15037 0.00658571
R60574 DVSS.n15077 DVSS.n15076 0.00658571
R60575 DVSS.n19967 DVSS.n15077 0.00658571
R60576 DVSS.n19967 DVSS.n19966 0.00658571
R60577 DVSS.n19966 DVSS.n19965 0.00658571
R60578 DVSS.n19965 DVSS.n15078 0.00658571
R60579 DVSS.n19959 DVSS.n15078 0.00658571
R60580 DVSS.n19959 DVSS.n19958 0.00658571
R60581 DVSS.n19958 DVSS.n19957 0.00658571
R60582 DVSS.n19957 DVSS.n15082 0.00658571
R60583 DVSS.n19948 DVSS.n15082 0.00658571
R60584 DVSS.n19948 DVSS.n19947 0.00658571
R60585 DVSS.n19947 DVSS.n19946 0.00658571
R60586 DVSS.n19946 DVSS.n15121 0.00658571
R60587 DVSS.n19939 DVSS.n15121 0.00658571
R60588 DVSS.n19939 DVSS.n19938 0.00658571
R60589 DVSS.n19938 DVSS.n19937 0.00658571
R60590 DVSS.n19932 DVSS.n19931 0.00658571
R60591 DVSS.n21150 DVSS.n13689 0.00658571
R60592 DVSS.n20743 DVSS.n13689 0.00658571
R60593 DVSS.n20743 DVSS.n20742 0.00658571
R60594 DVSS.n20750 DVSS.n20742 0.00658571
R60595 DVSS.n20751 DVSS.n20750 0.00658571
R60596 DVSS.n20752 DVSS.n20751 0.00658571
R60597 DVSS.n20752 DVSS.n20739 0.00658571
R60598 DVSS.n20759 DVSS.n20739 0.00658571
R60599 DVSS.n20760 DVSS.n20759 0.00658571
R60600 DVSS.n20761 DVSS.n20760 0.00658571
R60601 DVSS.n20761 DVSS.n20736 0.00658571
R60602 DVSS.n20766 DVSS.n20736 0.00658571
R60603 DVSS.n20767 DVSS.n20766 0.00658571
R60604 DVSS.n20769 DVSS.n20767 0.00658571
R60605 DVSS.n20769 DVSS.n20768 0.00658571
R60606 DVSS.n20768 DVSS.n20733 0.00658571
R60607 DVSS.n20733 DVSS.n20731 0.00658571
R60608 DVSS.n20779 DVSS.n20731 0.00658571
R60609 DVSS.n20780 DVSS.n20779 0.00658571
R60610 DVSS.n20781 DVSS.n20780 0.00658571
R60611 DVSS.n20781 DVSS.n20728 0.00658571
R60612 DVSS.n20788 DVSS.n20728 0.00658571
R60613 DVSS.n20789 DVSS.n20788 0.00658571
R60614 DVSS.n20790 DVSS.n20789 0.00658571
R60615 DVSS.n20790 DVSS.n20725 0.00658571
R60616 DVSS.n20797 DVSS.n20725 0.00658571
R60617 DVSS.n20798 DVSS.n20797 0.00658571
R60618 DVSS.n20799 DVSS.n20798 0.00658571
R60619 DVSS.n20799 DVSS.n14504 0.00658571
R60620 DVSS.n20808 DVSS.n14504 0.00658571
R60621 DVSS.n20809 DVSS.n20808 0.00658571
R60622 DVSS.n20811 DVSS.n20809 0.00658571
R60623 DVSS.n20811 DVSS.n20810 0.00658571
R60624 DVSS.n20810 DVSS.n14500 0.00658571
R60625 DVSS.n20823 DVSS.n14500 0.00658571
R60626 DVSS.n20824 DVSS.n20823 0.00658571
R60627 DVSS.n20825 DVSS.n20824 0.00658571
R60628 DVSS.n20825 DVSS.n14497 0.00658571
R60629 DVSS.n20832 DVSS.n14497 0.00658571
R60630 DVSS.n20833 DVSS.n20832 0.00658571
R60631 DVSS.n20834 DVSS.n20833 0.00658571
R60632 DVSS.n20834 DVSS.n14494 0.00658571
R60633 DVSS.n20841 DVSS.n14494 0.00658571
R60634 DVSS.n20842 DVSS.n20841 0.00658571
R60635 DVSS.n20844 DVSS.n20842 0.00658571
R60636 DVSS.n20844 DVSS.n20843 0.00658571
R60637 DVSS.n20843 DVSS.n14457 0.00658571
R60638 DVSS.n20853 DVSS.n14457 0.00658571
R60639 DVSS.n20854 DVSS.n20853 0.00658571
R60640 DVSS.n20856 DVSS.n20854 0.00658571
R60641 DVSS.n20856 DVSS.n20855 0.00658571
R60642 DVSS.n20855 DVSS.n14453 0.00658571
R60643 DVSS.n20864 DVSS.n14453 0.00658571
R60644 DVSS.n20865 DVSS.n20864 0.00658571
R60645 DVSS.n20866 DVSS.n20865 0.00658571
R60646 DVSS.n20866 DVSS.n14450 0.00658571
R60647 DVSS.n20873 DVSS.n14450 0.00658571
R60648 DVSS.n20874 DVSS.n20873 0.00658571
R60649 DVSS.n20875 DVSS.n20874 0.00658571
R60650 DVSS.n20875 DVSS.n14447 0.00658571
R60651 DVSS.n20882 DVSS.n14447 0.00658571
R60652 DVSS.n20883 DVSS.n20882 0.00658571
R60653 DVSS.n20884 DVSS.n20883 0.00658571
R60654 DVSS.n20884 DVSS.n14408 0.00658571
R60655 DVSS.n20893 DVSS.n14408 0.00658571
R60656 DVSS.n20894 DVSS.n20893 0.00658571
R60657 DVSS.n20896 DVSS.n20894 0.00658571
R60658 DVSS.n20896 DVSS.n20895 0.00658571
R60659 DVSS.n20895 DVSS.n14404 0.00658571
R60660 DVSS.n20904 DVSS.n14404 0.00658571
R60661 DVSS.n20905 DVSS.n20904 0.00658571
R60662 DVSS.n20906 DVSS.n20905 0.00658571
R60663 DVSS.n20906 DVSS.n14401 0.00658571
R60664 DVSS.n20913 DVSS.n14401 0.00658571
R60665 DVSS.n20914 DVSS.n20913 0.00658571
R60666 DVSS.n20915 DVSS.n20914 0.00658571
R60667 DVSS.n20915 DVSS.n14398 0.00658571
R60668 DVSS.n20922 DVSS.n14398 0.00658571
R60669 DVSS.n20923 DVSS.n20922 0.00658571
R60670 DVSS.n20924 DVSS.n20923 0.00658571
R60671 DVSS.n20924 DVSS.n14359 0.00658571
R60672 DVSS.n20933 DVSS.n14359 0.00658571
R60673 DVSS.n20934 DVSS.n20933 0.00658571
R60674 DVSS.n20935 DVSS.n20934 0.00658571
R60675 DVSS.n20935 DVSS.n14355 0.00658571
R60676 DVSS.n20941 DVSS.n14355 0.00658571
R60677 DVSS.n20942 DVSS.n20941 0.00658571
R60678 DVSS.n20973 DVSS.n20942 0.00658571
R60679 DVSS.n20973 DVSS.n20972 0.00658571
R60680 DVSS.n20972 DVSS.n20971 0.00658571
R60681 DVSS.n20971 DVSS.n20943 0.00658571
R60682 DVSS.n20959 DVSS.n20943 0.00658571
R60683 DVSS.n20959 DVSS.n20958 0.00658571
R60684 DVSS.n20958 DVSS.n20957 0.00658571
R60685 DVSS.n20957 DVSS.n20946 0.00658571
R60686 DVSS.n20950 DVSS.n20946 0.00658571
R60687 DVSS.n20950 DVSS.n20949 0.00658571
R60688 DVSS.n20981 DVSS.n14318 0.00658571
R60689 DVSS.n21186 DVSS.n21185 0.00658571
R60690 DVSS.n21187 DVSS.n21186 0.00658571
R60691 DVSS.n21187 DVSS.n13655 0.00658571
R60692 DVSS.n21194 DVSS.n13655 0.00658571
R60693 DVSS.n21195 DVSS.n21194 0.00658571
R60694 DVSS.n21196 DVSS.n21195 0.00658571
R60695 DVSS.n21196 DVSS.n13652 0.00658571
R60696 DVSS.n21208 DVSS.n13652 0.00658571
R60697 DVSS.n21209 DVSS.n21208 0.00658571
R60698 DVSS.n21210 DVSS.n21209 0.00658571
R60699 DVSS.n21210 DVSS.n13616 0.00658571
R60700 DVSS.n21218 DVSS.n13616 0.00658571
R60701 DVSS.n21219 DVSS.n21218 0.00658571
R60702 DVSS.n21221 DVSS.n21219 0.00658571
R60703 DVSS.n21221 DVSS.n21220 0.00658571
R60704 DVSS.n21220 DVSS.n13612 0.00658571
R60705 DVSS.n21229 DVSS.n13612 0.00658571
R60706 DVSS.n21230 DVSS.n21229 0.00658571
R60707 DVSS.n21231 DVSS.n21230 0.00658571
R60708 DVSS.n21231 DVSS.n13609 0.00658571
R60709 DVSS.n21238 DVSS.n13609 0.00658571
R60710 DVSS.n21239 DVSS.n21238 0.00658571
R60711 DVSS.n21240 DVSS.n21239 0.00658571
R60712 DVSS.n21240 DVSS.n13606 0.00658571
R60713 DVSS.n21247 DVSS.n13606 0.00658571
R60714 DVSS.n21248 DVSS.n21247 0.00658571
R60715 DVSS.n21249 DVSS.n21248 0.00658571
R60716 DVSS.n21249 DVSS.n13568 0.00658571
R60717 DVSS.n21260 DVSS.n13568 0.00658571
R60718 DVSS.n21261 DVSS.n21260 0.00658571
R60719 DVSS.n21263 DVSS.n21261 0.00658571
R60720 DVSS.n21263 DVSS.n21262 0.00658571
R60721 DVSS.n21262 DVSS.n13565 0.00658571
R60722 DVSS.n13565 DVSS.n13563 0.00658571
R60723 DVSS.n21273 DVSS.n13563 0.00658571
R60724 DVSS.n21274 DVSS.n21273 0.00658571
R60725 DVSS.n21275 DVSS.n21274 0.00658571
R60726 DVSS.n21275 DVSS.n13560 0.00658571
R60727 DVSS.n21282 DVSS.n13560 0.00658571
R60728 DVSS.n21283 DVSS.n21282 0.00658571
R60729 DVSS.n21284 DVSS.n21283 0.00658571
R60730 DVSS.n21284 DVSS.n13557 0.00658571
R60731 DVSS.n21291 DVSS.n13557 0.00658571
R60732 DVSS.n21292 DVSS.n21291 0.00658571
R60733 DVSS.n21294 DVSS.n21292 0.00658571
R60734 DVSS.n21294 DVSS.n21293 0.00658571
R60735 DVSS.n21293 DVSS.n13514 0.00658571
R60736 DVSS.n21303 DVSS.n13514 0.00658571
R60737 DVSS.n21304 DVSS.n21303 0.00658571
R60738 DVSS.n21306 DVSS.n21304 0.00658571
R60739 DVSS.n21306 DVSS.n21305 0.00658571
R60740 DVSS.n21305 DVSS.n13510 0.00658571
R60741 DVSS.n21314 DVSS.n13510 0.00658571
R60742 DVSS.n21315 DVSS.n21314 0.00658571
R60743 DVSS.n21316 DVSS.n21315 0.00658571
R60744 DVSS.n21316 DVSS.n13507 0.00658571
R60745 DVSS.n21323 DVSS.n13507 0.00658571
R60746 DVSS.n21324 DVSS.n21323 0.00658571
R60747 DVSS.n21325 DVSS.n21324 0.00658571
R60748 DVSS.n21325 DVSS.n13504 0.00658571
R60749 DVSS.n21332 DVSS.n13504 0.00658571
R60750 DVSS.n21333 DVSS.n21332 0.00658571
R60751 DVSS.n21334 DVSS.n21333 0.00658571
R60752 DVSS.n21334 DVSS.n13463 0.00658571
R60753 DVSS.n21343 DVSS.n13463 0.00658571
R60754 DVSS.n21344 DVSS.n21343 0.00658571
R60755 DVSS.n21346 DVSS.n21344 0.00658571
R60756 DVSS.n21346 DVSS.n21345 0.00658571
R60757 DVSS.n21345 DVSS.n13459 0.00658571
R60758 DVSS.n21354 DVSS.n13459 0.00658571
R60759 DVSS.n21355 DVSS.n21354 0.00658571
R60760 DVSS.n21356 DVSS.n21355 0.00658571
R60761 DVSS.n21356 DVSS.n13456 0.00658571
R60762 DVSS.n21363 DVSS.n13456 0.00658571
R60763 DVSS.n21364 DVSS.n21363 0.00658571
R60764 DVSS.n21365 DVSS.n21364 0.00658571
R60765 DVSS.n21365 DVSS.n13453 0.00658571
R60766 DVSS.n21372 DVSS.n13453 0.00658571
R60767 DVSS.n21373 DVSS.n21372 0.00658571
R60768 DVSS.n21374 DVSS.n21373 0.00658571
R60769 DVSS.n21374 DVSS.n13417 0.00658571
R60770 DVSS.n21387 DVSS.n13417 0.00658571
R60771 DVSS.n21388 DVSS.n21387 0.00658571
R60772 DVSS.n21389 DVSS.n21388 0.00658571
R60773 DVSS.n21389 DVSS.n13413 0.00658571
R60774 DVSS.n21395 DVSS.n13413 0.00658571
R60775 DVSS.n21396 DVSS.n21395 0.00658571
R60776 DVSS.n21427 DVSS.n21396 0.00658571
R60777 DVSS.n21427 DVSS.n21426 0.00658571
R60778 DVSS.n21426 DVSS.n21425 0.00658571
R60779 DVSS.n21425 DVSS.n21397 0.00658571
R60780 DVSS.n21413 DVSS.n21397 0.00658571
R60781 DVSS.n21413 DVSS.n21412 0.00658571
R60782 DVSS.n21412 DVSS.n21411 0.00658571
R60783 DVSS.n21411 DVSS.n21400 0.00658571
R60784 DVSS.n21404 DVSS.n21400 0.00658571
R60785 DVSS.n21435 DVSS.n13375 0.00658571
R60786 DVSS.n17851 DVSS.n15863 0.00655634
R60787 DVSS.n15774 DVSS.n15767 0.00655634
R60788 DVSS.n16678 DVSS.n16255 0.00654286
R60789 DVSS.n16722 DVSS.n15654 0.00654286
R60790 DVSS.n17633 DVSS.n16099 0.00654286
R60791 DVSS.n17584 DVSS.n17540 0.00654286
R60792 DVSS.n15352 DVSS.n15309 0.00654286
R60793 DVSS.n18294 DVSS.n15460 0.00654286
R60794 DVSS.n19999 DVSS.n14908 0.00654286
R60795 DVSS.n15071 DVSS.n15066 0.00654286
R60796 DVSS.n20846 DVSS.n14475 0.00654286
R60797 DVSS.n14396 DVSS.n14395 0.00654286
R60798 DVSS.n21296 DVSS.n13533 0.00654286
R60799 DVSS.n13451 DVSS.n13436 0.00654286
R60800 DVSS.n22754 DVSS.n612 0.00654286
R60801 DVSS.n22830 DVSS.n516 0.00654286
R60802 DVSS.n6251 DVSS.n1501 0.00651579
R60803 DVSS.n13102 DVSS.n13101 0.00651579
R60804 DVSS.n22547 DVSS.n778 0.0065
R60805 DVSS.n23075 DVSS.n270 0.0065
R60806 DVSS.n22047 DVSS.n160 0.0065
R60807 DVSS.n22076 DVSS.n21556 0.0065
R60808 DVSS.n12974 DVSS.n160 0.0065
R60809 DVSS.n1486 DVSS.n1485 0.0065
R60810 DVSS.n21556 DVSS.n21555 0.0065
R60811 DVSS.n23190 DVSS.n54 0.0065
R60812 DVSS.n23190 DVSS.n55 0.0065
R60813 DVSS.n1485 DVSS.n1484 0.0065
R60814 DVSS.n22013 DVSS.n53 0.0065
R60815 DVSS.n23075 DVSS.n271 0.0065
R60816 DVSS.n22547 DVSS.n779 0.0065
R60817 DVSS.n23127 DVSS.n187 0.0065
R60818 DVSS.n23127 DVSS.n188 0.0065
R60819 DVSS.n22995 DVSS.n53 0.0065
R60820 DVSS.n18012 DVSS.n15557 0.00648592
R60821 DVSS.n8129 DVSS.n4008 0.00645489
R60822 DVSS.n17950 DVSS.n17949 0.00641549
R60823 DVSS.n15703 DVSS.n15690 0.00641549
R60824 DVSS DVSS.n456 0.00641429
R60825 DVSS.n16741 DVSS 0.00641429
R60826 DVSS.n16634 DVSS.n16633 0.00641429
R60827 DVSS.n16225 DVSS.n16163 0.00641429
R60828 DVSS.n18179 DVSS 0.00641429
R60829 DVSS.n16059 DVSS.n16027 0.00641429
R60830 DVSS.n16857 DVSS.n16848 0.00641429
R60831 DVSS.n18253 DVSS 0.00641429
R60832 DVSS.n18362 DVSS.n15251 0.00641429
R60833 DVSS.n15401 DVSS.n15392 0.00641429
R60834 DVSS.n19932 DVSS 0.00641429
R60835 DVSS.n18427 DVSS.n18392 0.00641429
R60836 DVSS.n14963 DVSS.n14955 0.00641429
R60837 DVSS DVSS.n14318 0.00641429
R60838 DVSS.n20723 DVSS.n20718 0.00641429
R60839 DVSS.n20880 DVSS.n14438 0.00641429
R60840 DVSS DVSS.n13375 0.00641429
R60841 DVSS.n21252 DVSS.n21251 0.00641429
R60842 DVSS.n21330 DVSS.n13494 0.00641429
R60843 DVSS.n22710 DVSS.n22709 0.00641429
R60844 DVSS.n22788 DVSS.n579 0.00641429
R60845 DVSS.n16504 DVSS.n16491 0.00637368
R60846 DVSS.n16508 DVSS.n16491 0.00637368
R60847 DVSS.n16509 DVSS.n16508 0.00637368
R60848 DVSS.n16510 DVSS.n16509 0.00637368
R60849 DVSS.n16510 DVSS.n16489 0.00637368
R60850 DVSS.n16514 DVSS.n16489 0.00637368
R60851 DVSS.n16515 DVSS.n16514 0.00637368
R60852 DVSS.n16515 DVSS.n16487 0.00637368
R60853 DVSS.n16519 DVSS.n16487 0.00637368
R60854 DVSS.n16520 DVSS.n16519 0.00637368
R60855 DVSS.n16521 DVSS.n16520 0.00637368
R60856 DVSS.n16521 DVSS.n16485 0.00637368
R60857 DVSS.n16525 DVSS.n16485 0.00637368
R60858 DVSS.n16526 DVSS.n16525 0.00637368
R60859 DVSS.n16527 DVSS.n16526 0.00637368
R60860 DVSS.n18147 DVSS.n15576 0.00637368
R60861 DVSS.n18143 DVSS.n15576 0.00637368
R60862 DVSS.n18143 DVSS.n18142 0.00637368
R60863 DVSS.n18142 DVSS.n18141 0.00637368
R60864 DVSS.n18141 DVSS.n15583 0.00637368
R60865 DVSS.n18137 DVSS.n15583 0.00637368
R60866 DVSS.n18137 DVSS.n18136 0.00637368
R60867 DVSS.n18136 DVSS.n15585 0.00637368
R60868 DVSS.n18132 DVSS.n15585 0.00637368
R60869 DVSS.n18132 DVSS.n18131 0.00637368
R60870 DVSS.n18131 DVSS.n18130 0.00637368
R60871 DVSS.n18130 DVSS.n15587 0.00637368
R60872 DVSS.n18126 DVSS.n15587 0.00637368
R60873 DVSS.n18126 DVSS.n18125 0.00637368
R60874 DVSS.n18125 DVSS.n18124 0.00637368
R60875 DVSS.n18903 DVSS.n14559 0.00636957
R60876 DVSS.n18943 DVSS.n14562 0.00636957
R60877 DVSS.n20675 DVSS.n20674 0.00636957
R60878 DVSS.n20125 DVSS.n14595 0.00636957
R60879 DVSS.n20202 DVSS.n14647 0.00636957
R60880 DVSS.n20646 DVSS.n20645 0.00636957
R60881 DVSS.n20429 DVSS.n20428 0.00636957
R60882 DVSS.n20445 DVSS.n20341 0.00636957
R60883 DVSS.n18888 DVSS.n14528 0.00636957
R60884 DVSS.n18947 DVSS.n14529 0.00636957
R60885 DVSS.n20107 DVSS.n20019 0.00636957
R60886 DVSS.n20098 DVSS.n20020 0.00636957
R60887 DVSS.n20204 DVSS.n20192 0.00636957
R60888 DVSS.n20318 DVSS.n20317 0.00636957
R60889 DVSS.n20365 DVSS.n20330 0.00636957
R60890 DVSS.n20344 DVSS.n20331 0.00636957
R60891 DVSS.n16760 DVSS.n15604 0.00635
R60892 DVSS.n15522 DVSS.n15504 0.00635
R60893 DVSS.n18274 DVSS.n18273 0.00635
R60894 DVSS.n19954 DVSS.n15091 0.00635
R60895 DVSS.n20969 DVSS.n14350 0.00635
R60896 DVSS.n21423 DVSS.n13408 0.00635
R60897 DVSS.n16404 DVSS.n16403 0.00635
R60898 DVSS.n18060 DVSS.n15684 0.00635
R60899 DVSS.n22856 DVSS.n478 0.00635
R60900 DVSS.n17824 DVSS.n17823 0.00634507
R60901 DVSS.n4010 DVSS.n4009 0.00631955
R60902 DVSS.n2709 DVSS.n2369 0.00629866
R60903 DVSS.n10168 DVSS.n2026 0.00629866
R60904 DVSS.n2711 DVSS.n2368 0.00629866
R60905 DVSS.n10169 DVSS.n2025 0.00629866
R60906 DVSS.n16616 DVSS.n16315 0.00628571
R60907 DVSS.n16696 DVSS.n16160 0.00628571
R60908 DVSS.n16043 DVSS.n16022 0.00628571
R60909 DVSS.n17617 DVSS.n16147 0.00628571
R60910 DVSS.n15274 DVSS.n15248 0.00628571
R60911 DVSS.n18327 DVSS.n15368 0.00628571
R60912 DVSS.n18410 DVSS.n18387 0.00628571
R60913 DVSS.n19983 DVSS.n14933 0.00628571
R60914 DVSS.n20782 DVSS.n20713 0.00628571
R60915 DVSS.n14451 DVSS.n14433 0.00628571
R60916 DVSS.n21234 DVSS.n13595 0.00628571
R60917 DVSS.n13508 DVSS.n13489 0.00628571
R60918 DVSS.n22692 DVSS.n682 0.00628571
R60919 DVSS.n588 DVSS.n574 0.00628571
R60920 DVSS.n17893 DVSS.n15803 0.00627465
R60921 DVSS.n17972 DVSS.n15694 0.00627465
R60922 DVSS.n12766 DVSS.n12554 0.0062375
R60923 DVSS.n12767 DVSS.n12458 0.0062375
R60924 DVSS.n6653 DVSS.n6235 0.0062375
R60925 DVSS.n6655 DVSS.n6236 0.0062375
R60926 DVSS.n15911 DVSS.n15904 0.00620423
R60927 DVSS.n6672 DVSS.n6236 0.00619869
R60928 DVSS.n7077 DVSS.n5185 0.00619869
R60929 DVSS.n6673 DVSS.n6235 0.00619869
R60930 DVSS.n7076 DVSS.n5186 0.00619869
R60931 DVSS.n16609 DVSS.n16314 0.00615714
R60932 DVSS.n17656 DVSS.n17655 0.00615714
R60933 DVSS.n17754 DVSS.n15247 0.00615714
R60934 DVSS.n15228 DVSS.n15227 0.00615714
R60935 DVSS.n20775 DVSS.n20712 0.00615714
R60936 DVSS.n21227 DVSS.n13594 0.00615714
R60937 DVSS.n22685 DVSS.n681 0.00615714
R60938 DVSS.n17822 DVSS.n15899 0.00613684
R60939 DVSS.n15564 DVSS.n15545 0.00613684
R60940 DVSS.n17877 DVSS.n15811 0.0061338
R60941 DVSS.n16405 DVSS 0.006125
R60942 DVSS DVSS.n18061 0.006125
R60943 DVSS.n21016 DVSS.n21015 0.006125
R60944 DVSS.n16728 DVSS.n15605 0.00609286
R60945 DVSS.n18205 DVSS.n15505 0.00609286
R60946 DVSS.n18277 DVSS.n18276 0.00609286
R60947 DVSS.n19961 DVSS.n15080 0.00609286
R60948 DVSS.n20976 DVSS.n14351 0.00609286
R60949 DVSS.n21430 DVSS.n13409 0.00609286
R60950 DVSS.n22849 DVSS.n475 0.00609286
R60951 DVSS.n4010 DVSS.n1503 0.00607561
R60952 DVSS.n9766 DVSS.n1504 0.00607561
R60953 DVSS.n7110 DVSS.n1502 0.00607561
R60954 DVSS.n13364 DVSS.n13363 0.00607561
R60955 DVSS.n17803 DVSS.n15896 0.00606338
R60956 DVSS.n18957 DVSS.n18878 0.0060618
R60957 DVSS.n20159 DVSS.n20044 0.0060618
R60958 DVSS.n20261 DVSS.n20219 0.0060618
R60959 DVSS.n20422 DVSS.n14689 0.0060618
R60960 DVSS.n16625 DVSS.n16319 0.00602857
R60961 DVSS.n16705 DVSS.n16162 0.00602857
R60962 DVSS.n16052 DVSS.n16026 0.00602857
R60963 DVSS.n16870 DVSS.n16847 0.00602857
R60964 DVSS.n18369 DVSS.n15250 0.00602857
R60965 DVSS.n15414 DVSS.n15391 0.00602857
R60966 DVSS.n18419 DVSS.n18391 0.00602857
R60967 DVSS.n14976 DVSS.n14954 0.00602857
R60968 DVSS.n20791 DVSS.n20717 0.00602857
R60969 DVSS.n14448 DVSS.n14437 0.00602857
R60970 DVSS.n21243 DVSS.n13603 0.00602857
R60971 DVSS.n13505 DVSS.n13493 0.00602857
R60972 DVSS.n22701 DVSS.n686 0.00602857
R60973 DVSS.n585 DVSS.n578 0.00602857
R60974 DVSS.n17888 DVSS.n15817 0.00599296
R60975 DVSS.n17968 DVSS.n15699 0.00599296
R60976 DVSS.n21590 DVSS.n21589 0.0059878
R60977 DVSS.n22339 DVSS.n1178 0.0059878
R60978 DVSS.n22458 DVSS.n870 0.0059878
R60979 DVSS.n22336 DVSS.n1199 0.0059878
R60980 DVSS.n16751 DVSS.n15600 0.00596429
R60981 DVSS.n18189 DVSS.n15501 0.00596429
R60982 DVSS.n18263 DVSS.n18228 0.00596429
R60983 DVSS.n19942 DVSS.n15112 0.00596429
R60984 DVSS.n20955 DVSS.n14346 0.00596429
R60985 DVSS.n21409 DVSS.n13404 0.00596429
R60986 DVSS.n22865 DVSS.n482 0.00596429
R60987 DVSS.n16394 DVSS.n16393 0.0059439
R60988 DVSS.n16395 DVSS.n16394 0.0059439
R60989 DVSS.n16395 DVSS.n16381 0.0059439
R60990 DVSS.n16399 DVSS.n16381 0.0059439
R60991 DVSS.n16400 DVSS.n16399 0.0059439
R60992 DVSS.n16401 DVSS.n16400 0.0059439
R60993 DVSS.n16401 DVSS.n16379 0.0059439
R60994 DVSS.n16406 DVSS.n16379 0.0059439
R60995 DVSS.n16407 DVSS.n16406 0.0059439
R60996 DVSS.n16408 DVSS.n16407 0.0059439
R60997 DVSS.n16408 DVSS.n16377 0.0059439
R60998 DVSS.n16412 DVSS.n16377 0.0059439
R60999 DVSS.n16413 DVSS.n16412 0.0059439
R61000 DVSS.n16414 DVSS.n16413 0.0059439
R61001 DVSS.n16414 DVSS.n16304 0.0059439
R61002 DVSS.n18048 DVSS.n15687 0.0059439
R61003 DVSS.n18052 DVSS.n15687 0.0059439
R61004 DVSS.n18053 DVSS.n18052 0.0059439
R61005 DVSS.n18054 DVSS.n18053 0.0059439
R61006 DVSS.n18054 DVSS.n15685 0.0059439
R61007 DVSS.n18058 DVSS.n15685 0.0059439
R61008 DVSS.n18059 DVSS.n18058 0.0059439
R61009 DVSS.n18059 DVSS.n15683 0.0059439
R61010 DVSS.n18063 DVSS.n15683 0.0059439
R61011 DVSS.n18064 DVSS.n18063 0.0059439
R61012 DVSS.n18065 DVSS.n18064 0.0059439
R61013 DVSS.n18065 DVSS.n15681 0.0059439
R61014 DVSS.n18069 DVSS.n15681 0.0059439
R61015 DVSS.n18070 DVSS.n18069 0.0059439
R61016 DVSS.n18071 DVSS.n18070 0.0059439
R61017 DVSS.n17820 DVSS.n15891 0.00592254
R61018 DVSS.n18002 DVSS.n18001 0.00591803
R61019 DVSS.n17795 DVSS.n15916 0.00591803
R61020 DVSS.n7038 DVSS.n7037 0.00591353
R61021 DVSS.n7823 DVSS.n7822 0.00591353
R61022 DVSS.n16824 DVSS.n16165 0.0059
R61023 DVSS.n15668 DVSS.n15653 0.0059
R61024 DVSS.n17615 DVSS.n16852 0.0059
R61025 DVSS.n17577 DVSS.n17535 0.0059
R61026 DVSS.n18325 DVSS.n15396 0.0059
R61027 DVSS.n18287 DVSS.n15456 0.0059
R61028 DVSS.n19981 DVSS.n14958 0.0059
R61029 DVSS.n15033 DVSS.n15017 0.0059
R61030 DVSS.n20891 DVSS.n20890 0.0059
R61031 DVSS.n20931 DVSS.n14361 0.0059
R61032 DVSS.n21341 DVSS.n21340 0.0059
R61033 DVSS.n21385 DVSS.n13419 0.0059
R61034 DVSS.n22799 DVSS.n22798 0.0059
R61035 DVSS.n512 DVSS.n496 0.0059
R61036 DVSS.n16550 DVSS.n16340 0.00585263
R61037 DVSS.n18116 DVSS.n18114 0.00585263
R61038 DVSS.n17908 DVSS.n15785 0.00585211
R61039 DVSS.n18036 DVSS.n15702 0.00585211
R61040 DVSS.n16598 DVSS.n16597 0.00583571
R61041 DVSS.n17777 DVSS.n15956 0.00583571
R61042 DVSS.n17774 DVSS.n17698 0.00583571
R61043 DVSS.n18490 DVSS.n18489 0.00583571
R61044 DVSS.n21145 DVSS.n13721 0.00583571
R61045 DVSS.n21216 DVSS.n21215 0.00583571
R61046 DVSS.n22674 DVSS.n22673 0.00583571
R61047 DVSS.n8122 DVSS.n3902 0.00581544
R61048 DVSS.n8124 DVSS.n8123 0.00581544
R61049 DVSS.n18008 DVSS.n15554 0.00578169
R61050 DVSS.n16667 DVSS.n16258 0.00577143
R61051 DVSS.n16719 DVSS.n15657 0.00577143
R61052 DVSS.n16128 DVSS.n16077 0.00577143
R61053 DVSS.n17593 DVSS.n17544 0.00577143
R61054 DVSS.n15343 DVSS.n15312 0.00577143
R61055 DVSS.n18303 DVSS.n15464 0.00577143
R61056 DVSS.n18445 DVSS.n14878 0.00577143
R61057 DVSS.n15056 DVSS.n15021 0.00577143
R61058 DVSS.n20835 DVSS.n14478 0.00577143
R61059 DVSS.n14399 DVSS.n14380 0.00577143
R61060 DVSS.n21285 DVSS.n13536 0.00577143
R61061 DVSS.n13454 DVSS.n13439 0.00577143
R61062 DVSS.n22743 DVSS.n618 0.00577143
R61063 DVSS.n22821 DVSS.n519 0.00577143
R61064 DVSS.n17907 DVSS.n15812 0.00572439
R61065 DVSS.n17948 DVSS.n15543 0.00572439
R61066 DVSS.n17864 DVSS.n15857 0.00572439
R61067 DVSS.n19002 DVSS.n13577 0.00572439
R61068 DVSS.n18045 DVSS.n15544 0.00572439
R61069 DVSS.n19181 DVSS.n13426 0.00572439
R61070 DVSS.n14795 DVSS.n14740 0.00572184
R61071 DVSS.n15864 DVSS.n15851 0.00571127
R61072 DVSS.n17937 DVSS.n15758 0.00571127
R61073 DVSS.n16562 DVSS.n16555 0.00570714
R61074 DVSS.n15977 DVSS.n15951 0.00570714
R61075 DVSS.n17734 DVSS.n17686 0.00570714
R61076 DVSS.n15201 DVSS.n15179 0.00570714
R61077 DVSS.n20740 DVSS.n13716 0.00570714
R61078 DVSS.n13653 DVSS.n13646 0.00570714
R61079 DVSS.n22641 DVSS.n725 0.00570714
R61080 DVSS.n7030 DVSS.n7029 0.005675
R61081 DVSS.n18822 DVSS.n18820 0.00566892
R61082 DVSS.n16651 DVSS.n16266 0.00564286
R61083 DVSS.n17644 DVSS.n16073 0.00564286
R61084 DVSS.n15290 DVSS.n15286 0.00564286
R61085 DVSS.n18461 DVSS.n14882 0.00564286
R61086 DVSS.n20819 DVSS.n20818 0.00564286
R61087 DVSS.n21269 DVSS.n13540 0.00564286
R61088 DVSS.n22727 DVSS.n622 0.00564286
R61089 DVSS.n18022 DVSS.n15550 0.00564085
R61090 DVSS.n19317 DVSS.n19307 0.00561579
R61091 DVSS.n19318 DVSS.n19317 0.00561579
R61092 DVSS.n19319 DVSS.n19318 0.00561579
R61093 DVSS.n19319 DVSS.n19305 0.00561579
R61094 DVSS.n19323 DVSS.n19305 0.00561579
R61095 DVSS.n19324 DVSS.n19323 0.00561579
R61096 DVSS.n19325 DVSS.n19324 0.00561579
R61097 DVSS.n19325 DVSS.n19303 0.00561579
R61098 DVSS.n19329 DVSS.n19303 0.00561579
R61099 DVSS.n19330 DVSS.n19329 0.00561579
R61100 DVSS.n19331 DVSS.n19330 0.00561579
R61101 DVSS.n19331 DVSS.n19301 0.00561579
R61102 DVSS.n19335 DVSS.n19301 0.00561579
R61103 DVSS.n19336 DVSS.n19335 0.00561579
R61104 DVSS.n19337 DVSS.n19336 0.00561579
R61105 DVSS.n19337 DVSS.n19299 0.00561579
R61106 DVSS.n19341 DVSS.n19299 0.00561579
R61107 DVSS.n19342 DVSS.n19341 0.00561579
R61108 DVSS.n19343 DVSS.n19342 0.00561579
R61109 DVSS.n19343 DVSS.n19297 0.00561579
R61110 DVSS.n19347 DVSS.n19297 0.00561579
R61111 DVSS.n19348 DVSS.n19347 0.00561579
R61112 DVSS.n19349 DVSS.n19348 0.00561579
R61113 DVSS.n19349 DVSS.n19295 0.00561579
R61114 DVSS.n19353 DVSS.n19295 0.00561579
R61115 DVSS.n19354 DVSS.n19353 0.00561579
R61116 DVSS.n19355 DVSS.n19354 0.00561579
R61117 DVSS.n19355 DVSS.n19293 0.00561579
R61118 DVSS.n19359 DVSS.n19293 0.00561579
R61119 DVSS.n19360 DVSS.n19359 0.00561579
R61120 DVSS.n19361 DVSS.n19360 0.00561579
R61121 DVSS.n19361 DVSS.n19291 0.00561579
R61122 DVSS.n19365 DVSS.n19291 0.00561579
R61123 DVSS.n19366 DVSS.n19365 0.00561579
R61124 DVSS.n19367 DVSS.n19366 0.00561579
R61125 DVSS.n19367 DVSS.n19289 0.00561579
R61126 DVSS.n19371 DVSS.n19289 0.00561579
R61127 DVSS.n19372 DVSS.n19371 0.00561579
R61128 DVSS.n19373 DVSS.n19372 0.00561579
R61129 DVSS.n19373 DVSS.n19287 0.00561579
R61130 DVSS.n19377 DVSS.n19287 0.00561579
R61131 DVSS.n19378 DVSS.n19377 0.00561579
R61132 DVSS.n19379 DVSS.n19378 0.00561579
R61133 DVSS.n19379 DVSS.n19285 0.00561579
R61134 DVSS.n19383 DVSS.n19285 0.00561579
R61135 DVSS.n19384 DVSS.n19383 0.00561579
R61136 DVSS.n19385 DVSS.n19384 0.00561579
R61137 DVSS.n19385 DVSS.n19283 0.00561579
R61138 DVSS.n19389 DVSS.n19283 0.00561579
R61139 DVSS.n19390 DVSS.n19389 0.00561579
R61140 DVSS.n19391 DVSS.n19390 0.00561579
R61141 DVSS.n19391 DVSS.n19281 0.00561579
R61142 DVSS.n19395 DVSS.n19281 0.00561579
R61143 DVSS.n19396 DVSS.n19395 0.00561579
R61144 DVSS.n19499 DVSS.n19396 0.00561579
R61145 DVSS.n19499 DVSS.n19498 0.00561579
R61146 DVSS.n19498 DVSS.n19497 0.00561579
R61147 DVSS.n19497 DVSS.n19397 0.00561579
R61148 DVSS.n19493 DVSS.n19397 0.00561579
R61149 DVSS.n19493 DVSS.n19492 0.00561579
R61150 DVSS.n19492 DVSS.n19491 0.00561579
R61151 DVSS.n19491 DVSS.n19399 0.00561579
R61152 DVSS.n19487 DVSS.n19399 0.00561579
R61153 DVSS.n19487 DVSS.n19486 0.00561579
R61154 DVSS.n19486 DVSS.n19485 0.00561579
R61155 DVSS.n19485 DVSS.n19401 0.00561579
R61156 DVSS.n19481 DVSS.n19401 0.00561579
R61157 DVSS.n19481 DVSS.n19480 0.00561579
R61158 DVSS.n19480 DVSS.n19479 0.00561579
R61159 DVSS.n19479 DVSS.n19403 0.00561579
R61160 DVSS.n19475 DVSS.n19403 0.00561579
R61161 DVSS.n19475 DVSS.n19474 0.00561579
R61162 DVSS.n19474 DVSS.n19473 0.00561579
R61163 DVSS.n19473 DVSS.n19405 0.00561579
R61164 DVSS.n19469 DVSS.n19405 0.00561579
R61165 DVSS.n19469 DVSS.n19468 0.00561579
R61166 DVSS.n19468 DVSS.n19467 0.00561579
R61167 DVSS.n19467 DVSS.n19407 0.00561579
R61168 DVSS.n19463 DVSS.n19407 0.00561579
R61169 DVSS.n19463 DVSS.n19462 0.00561579
R61170 DVSS.n19462 DVSS.n19461 0.00561579
R61171 DVSS.n19461 DVSS.n19409 0.00561579
R61172 DVSS.n19457 DVSS.n19409 0.00561579
R61173 DVSS.n19457 DVSS.n19456 0.00561579
R61174 DVSS.n19456 DVSS.n19455 0.00561579
R61175 DVSS.n19455 DVSS.n19411 0.00561579
R61176 DVSS.n19451 DVSS.n19411 0.00561579
R61177 DVSS.n19451 DVSS.n19450 0.00561579
R61178 DVSS.n19450 DVSS.n19449 0.00561579
R61179 DVSS.n19449 DVSS.n19413 0.00561579
R61180 DVSS.n19445 DVSS.n19413 0.00561579
R61181 DVSS.n19445 DVSS.n19444 0.00561579
R61182 DVSS.n19444 DVSS.n19443 0.00561579
R61183 DVSS.n19443 DVSS.n19415 0.00561579
R61184 DVSS.n19439 DVSS.n19415 0.00561579
R61185 DVSS.n19439 DVSS.n19438 0.00561579
R61186 DVSS.n19438 DVSS.n19437 0.00561579
R61187 DVSS.n19437 DVSS.n19417 0.00561579
R61188 DVSS.n19433 DVSS.n19417 0.00561579
R61189 DVSS.n19433 DVSS.n19432 0.00561579
R61190 DVSS.n19432 DVSS.n19431 0.00561579
R61191 DVSS.n19431 DVSS.n19419 0.00561579
R61192 DVSS.n19427 DVSS.n19419 0.00561579
R61193 DVSS.n19427 DVSS.n19426 0.00561579
R61194 DVSS.n19426 DVSS.n712 0.00561579
R61195 DVSS.n19421 DVSS.n19420 0.00561579
R61196 DVSS.n22217 DVSS.n22216 0.00561579
R61197 DVSS.n22211 DVSS.n22210 0.00561579
R61198 DVSS.n22210 DVSS.n22209 0.00561579
R61199 DVSS.n22209 DVSS.n1355 0.00561579
R61200 DVSS.n22205 DVSS.n1355 0.00561579
R61201 DVSS.n22205 DVSS.n22204 0.00561579
R61202 DVSS.n22204 DVSS.n22203 0.00561579
R61203 DVSS.n22203 DVSS.n1357 0.00561579
R61204 DVSS.n22199 DVSS.n1357 0.00561579
R61205 DVSS.n22199 DVSS.n22198 0.00561579
R61206 DVSS.n22198 DVSS.n22197 0.00561579
R61207 DVSS.n22197 DVSS.n1359 0.00561579
R61208 DVSS.n22193 DVSS.n1359 0.00561579
R61209 DVSS.n22193 DVSS.n22192 0.00561579
R61210 DVSS.n22192 DVSS.n22191 0.00561579
R61211 DVSS.n22191 DVSS.n1361 0.00561579
R61212 DVSS.n22187 DVSS.n1361 0.00561579
R61213 DVSS.n22187 DVSS.n22186 0.00561579
R61214 DVSS.n22177 DVSS.n22176 0.00561579
R61215 DVSS.n22161 DVSS.n22160 0.00561579
R61216 DVSS.n22145 DVSS.n22144 0.00561579
R61217 DVSS.n22133 DVSS.n881 0.00561579
R61218 DVSS.n22454 DVSS.n881 0.00561579
R61219 DVSS.n926 DVSS.n889 0.00561579
R61220 DVSS.n942 DVSS.n941 0.00561579
R61221 DVSS.n956 DVSS.n955 0.00561579
R61222 DVSS.n22450 DVSS.n925 0.00561579
R61223 DVSS.n22442 DVSS.n22441 0.00561579
R61224 DVSS.n22441 DVSS.n22440 0.00561579
R61225 DVSS.n22389 DVSS.n22388 0.00561579
R61226 DVSS.n22405 DVSS.n22404 0.00561579
R61227 DVSS.n22421 DVSS.n22420 0.00561579
R61228 DVSS.n19659 DVSS.n19138 0.00561579
R61229 DVSS.n19660 DVSS.n19659 0.00561579
R61230 DVSS.n19661 DVSS.n19660 0.00561579
R61231 DVSS.n19661 DVSS.n19136 0.00561579
R61232 DVSS.n19665 DVSS.n19136 0.00561579
R61233 DVSS.n19666 DVSS.n19665 0.00561579
R61234 DVSS.n19667 DVSS.n19666 0.00561579
R61235 DVSS.n19667 DVSS.n19134 0.00561579
R61236 DVSS.n19671 DVSS.n19134 0.00561579
R61237 DVSS.n19672 DVSS.n19671 0.00561579
R61238 DVSS.n19673 DVSS.n19672 0.00561579
R61239 DVSS.n19673 DVSS.n19132 0.00561579
R61240 DVSS.n19677 DVSS.n19132 0.00561579
R61241 DVSS.n19678 DVSS.n19677 0.00561579
R61242 DVSS.n19679 DVSS.n19678 0.00561579
R61243 DVSS.n19679 DVSS.n19130 0.00561579
R61244 DVSS.n19683 DVSS.n19130 0.00561579
R61245 DVSS.n19684 DVSS.n19683 0.00561579
R61246 DVSS.n19685 DVSS.n19684 0.00561579
R61247 DVSS.n19685 DVSS.n19128 0.00561579
R61248 DVSS.n19689 DVSS.n19128 0.00561579
R61249 DVSS.n19690 DVSS.n19689 0.00561579
R61250 DVSS.n19691 DVSS.n19690 0.00561579
R61251 DVSS.n19691 DVSS.n19126 0.00561579
R61252 DVSS.n19695 DVSS.n19126 0.00561579
R61253 DVSS.n19696 DVSS.n19695 0.00561579
R61254 DVSS.n19697 DVSS.n19696 0.00561579
R61255 DVSS.n19697 DVSS.n19124 0.00561579
R61256 DVSS.n19701 DVSS.n19124 0.00561579
R61257 DVSS.n19702 DVSS.n19701 0.00561579
R61258 DVSS.n19703 DVSS.n19702 0.00561579
R61259 DVSS.n19703 DVSS.n19122 0.00561579
R61260 DVSS.n19707 DVSS.n19122 0.00561579
R61261 DVSS.n19708 DVSS.n19707 0.00561579
R61262 DVSS.n19709 DVSS.n19708 0.00561579
R61263 DVSS.n19709 DVSS.n19120 0.00561579
R61264 DVSS.n19713 DVSS.n19120 0.00561579
R61265 DVSS.n19714 DVSS.n19713 0.00561579
R61266 DVSS.n19715 DVSS.n19714 0.00561579
R61267 DVSS.n19715 DVSS.n19118 0.00561579
R61268 DVSS.n19719 DVSS.n19118 0.00561579
R61269 DVSS.n19720 DVSS.n19719 0.00561579
R61270 DVSS.n19721 DVSS.n19720 0.00561579
R61271 DVSS.n19721 DVSS.n19116 0.00561579
R61272 DVSS.n19725 DVSS.n19116 0.00561579
R61273 DVSS.n19726 DVSS.n19725 0.00561579
R61274 DVSS.n19727 DVSS.n19726 0.00561579
R61275 DVSS.n19727 DVSS.n19114 0.00561579
R61276 DVSS.n19731 DVSS.n19114 0.00561579
R61277 DVSS.n19732 DVSS.n19731 0.00561579
R61278 DVSS.n19733 DVSS.n19732 0.00561579
R61279 DVSS.n19733 DVSS.n19112 0.00561579
R61280 DVSS.n19737 DVSS.n19112 0.00561579
R61281 DVSS.n19738 DVSS.n19737 0.00561579
R61282 DVSS.n19843 DVSS.n19738 0.00561579
R61283 DVSS.n19843 DVSS.n19842 0.00561579
R61284 DVSS.n19842 DVSS.n19841 0.00561579
R61285 DVSS.n19841 DVSS.n19739 0.00561579
R61286 DVSS.n19837 DVSS.n19739 0.00561579
R61287 DVSS.n19837 DVSS.n19836 0.00561579
R61288 DVSS.n19836 DVSS.n19835 0.00561579
R61289 DVSS.n19835 DVSS.n19741 0.00561579
R61290 DVSS.n19831 DVSS.n19741 0.00561579
R61291 DVSS.n19831 DVSS.n19830 0.00561579
R61292 DVSS.n19830 DVSS.n19829 0.00561579
R61293 DVSS.n19829 DVSS.n19743 0.00561579
R61294 DVSS.n19825 DVSS.n19743 0.00561579
R61295 DVSS.n19825 DVSS.n19824 0.00561579
R61296 DVSS.n19824 DVSS.n19823 0.00561579
R61297 DVSS.n19823 DVSS.n19745 0.00561579
R61298 DVSS.n19819 DVSS.n19745 0.00561579
R61299 DVSS.n19819 DVSS.n19818 0.00561579
R61300 DVSS.n19818 DVSS.n19817 0.00561579
R61301 DVSS.n19817 DVSS.n19747 0.00561579
R61302 DVSS.n19813 DVSS.n19747 0.00561579
R61303 DVSS.n19813 DVSS.n19812 0.00561579
R61304 DVSS.n19812 DVSS.n19811 0.00561579
R61305 DVSS.n19811 DVSS.n19749 0.00561579
R61306 DVSS.n19807 DVSS.n19749 0.00561579
R61307 DVSS.n19807 DVSS.n19806 0.00561579
R61308 DVSS.n19806 DVSS.n19805 0.00561579
R61309 DVSS.n19805 DVSS.n19751 0.00561579
R61310 DVSS.n19801 DVSS.n19751 0.00561579
R61311 DVSS.n19801 DVSS.n19800 0.00561579
R61312 DVSS.n19800 DVSS.n19799 0.00561579
R61313 DVSS.n19799 DVSS.n19753 0.00561579
R61314 DVSS.n19795 DVSS.n19753 0.00561579
R61315 DVSS.n19795 DVSS.n19794 0.00561579
R61316 DVSS.n19794 DVSS.n19793 0.00561579
R61317 DVSS.n19793 DVSS.n19755 0.00561579
R61318 DVSS.n19789 DVSS.n19755 0.00561579
R61319 DVSS.n19789 DVSS.n19788 0.00561579
R61320 DVSS.n19788 DVSS.n19787 0.00561579
R61321 DVSS.n19787 DVSS.n19757 0.00561579
R61322 DVSS.n19783 DVSS.n19757 0.00561579
R61323 DVSS.n19783 DVSS.n19782 0.00561579
R61324 DVSS.n19782 DVSS.n19781 0.00561579
R61325 DVSS.n19781 DVSS.n19759 0.00561579
R61326 DVSS.n19777 DVSS.n19759 0.00561579
R61327 DVSS.n19777 DVSS.n19776 0.00561579
R61328 DVSS.n19776 DVSS.n19775 0.00561579
R61329 DVSS.n19775 DVSS.n19761 0.00561579
R61330 DVSS.n19771 DVSS.n19761 0.00561579
R61331 DVSS.n19771 DVSS.n19770 0.00561579
R61332 DVSS.n19770 DVSS.n19769 0.00561579
R61333 DVSS.n19764 DVSS.n19763 0.00561579
R61334 DVSS.n22246 DVSS.n22245 0.00561579
R61335 DVSS.n22250 DVSS.n476 0.00561579
R61336 DVSS.n22250 DVSS.n1270 0.00561579
R61337 DVSS.n22254 DVSS.n1270 0.00561579
R61338 DVSS.n22255 DVSS.n22254 0.00561579
R61339 DVSS.n22256 DVSS.n22255 0.00561579
R61340 DVSS.n22256 DVSS.n1268 0.00561579
R61341 DVSS.n22260 DVSS.n1268 0.00561579
R61342 DVSS.n22261 DVSS.n22260 0.00561579
R61343 DVSS.n22262 DVSS.n22261 0.00561579
R61344 DVSS.n22262 DVSS.n1266 0.00561579
R61345 DVSS.n22266 DVSS.n1266 0.00561579
R61346 DVSS.n22267 DVSS.n22266 0.00561579
R61347 DVSS.n22268 DVSS.n22267 0.00561579
R61348 DVSS.n22268 DVSS.n1264 0.00561579
R61349 DVSS.n22272 DVSS.n1264 0.00561579
R61350 DVSS.n22273 DVSS.n22272 0.00561579
R61351 DVSS.n22274 DVSS.n22273 0.00561579
R61352 DVSS.n22286 DVSS.n22285 0.00561579
R61353 DVSS.n22302 DVSS.n22301 0.00561579
R61354 DVSS.n22318 DVSS.n22317 0.00561579
R61355 DVSS.n22331 DVSS.n22330 0.00561579
R61356 DVSS.n22332 DVSS.n22331 0.00561579
R61357 DVSS.n12821 DVSS.n12820 0.00561579
R61358 DVSS.n12837 DVSS.n12836 0.00561579
R61359 DVSS.n12851 DVSS.n12850 0.00561579
R61360 DVSS.n12867 DVSS.n12866 0.00561579
R61361 DVSS.n12874 DVSS.n36 0.00561579
R61362 DVSS.n12875 DVSS.n12874 0.00561579
R61363 DVSS.n12883 DVSS.n12882 0.00561579
R61364 DVSS.n12899 DVSS.n12898 0.00561579
R61365 DVSS.n12915 DVSS.n12914 0.00561579
R61366 DVSS.n16577 DVSS.n16351 0.00557857
R61367 DVSS.n15972 DVSS.n15946 0.00557857
R61368 DVSS.n17729 DVSS.n17679 0.00557857
R61369 DVSS.n15192 DVSS.n15174 0.00557857
R61370 DVSS.n20746 DVSS.n13711 0.00557857
R61371 DVSS.n21190 DVSS.n13639 0.00557857
R61372 DVSS.n22662 DVSS.n715 0.00557857
R61373 DVSS.n17840 DVSS.n15855 0.00557042
R61374 DVSS.n17921 DVSS.n15762 0.00557042
R61375 DVSS.n16529 DVSS.n16336 0.00556842
R61376 DVSS.n16531 DVSS.n16342 0.00556842
R61377 DVSS.n16533 DVSS.n16337 0.00556842
R61378 DVSS.n16535 DVSS.n16341 0.00556842
R61379 DVSS.n16537 DVSS.n16338 0.00556842
R61380 DVSS.n958 DVSS.n908 0.00556842
R61381 DVSS.n22391 DVSS.n1007 0.00556842
R61382 DVSS.n18121 DVSS.n15589 0.00556842
R61383 DVSS.n18120 DVSS.n15598 0.00556842
R61384 DVSS.n18096 DVSS.n15614 0.00556842
R61385 DVSS.n18098 DVSS.n15612 0.00556842
R61386 DVSS.n18100 DVSS.n15615 0.00556842
R61387 DVSS.n12853 DVSS.n9 0.00556842
R61388 DVSS.n12885 DVSS.n12810 0.00556842
R61389 DVSS.n18969 DVSS.n18913 0.00555618
R61390 DVSS.n20092 DVSS.n20054 0.00555618
R61391 DVSS.n20062 DVSS.n20050 0.00555618
R61392 DVSS.n20247 DVSS.n20223 0.00555618
R61393 DVSS.n20302 DVSS.n20210 0.00555618
R61394 DVSS.n20406 DVSS.n14684 0.00555618
R61395 DVSS.n21586 DVSS.n228 0.00554878
R61396 DVSS.n1197 DVSS.n148 0.00554878
R61397 DVSS.n22461 DVSS.n22460 0.00554878
R61398 DVSS.n1218 DVSS.n83 0.00554878
R61399 DVSS.n16662 DVSS.n16272 0.00551429
R61400 DVSS.n16796 DVSS.n15663 0.00551429
R61401 DVSS.n16124 DVSS.n16084 0.00551429
R61402 DVSS.n17597 DVSS.n16903 0.00551429
R61403 DVSS.n15339 DVSS.n15319 0.00551429
R61404 DVSS.n18307 DVSS.n15446 0.00551429
R61405 DVSS.n18442 DVSS.n14885 0.00551429
R61406 DVSS.n15051 DVSS.n15027 0.00551429
R61407 DVSS.n20830 DVSS.n14487 0.00551429
R61408 DVSS.n20909 DVSS.n14387 0.00551429
R61409 DVSS.n21280 DVSS.n13545 0.00551429
R61410 DVSS.n21359 DVSS.n13446 0.00551429
R61411 DVSS.n22738 DVSS.n628 0.00551429
R61412 DVSS.n22817 DVSS.n527 0.00551429
R61413 DVSS.n22883 DVSS.n455 0.00548841
R61414 DVSS.n22639 DVSS.n730 0.00548841
R61415 DVSS.n16739 DVSS.n16738 0.00548841
R61416 DVSS.n16569 DVSS.n16567 0.00548841
R61417 DVSS.n18177 DVSS.n18176 0.00548841
R61418 DVSS.n17783 DVSS.n15923 0.00548841
R61419 DVSS.n18251 DVSS.n18250 0.00548841
R61420 DVSS.n17722 DVSS.n17721 0.00548841
R61421 DVSS.n19930 DVSS.n19929 0.00548841
R61422 DVSS.n18496 DVSS.n15150 0.00548841
R61423 DVSS.n20982 DVSS.n14317 0.00548841
R61424 DVSS.n21151 DVSS.n13688 0.00548841
R61425 DVSS.n21436 DVSS.n13374 0.00548841
R61426 DVSS.n21182 DVSS.n13658 0.00548841
R61427 DVSS.n22229 DVSS.n711 0.00547368
R61428 DVSS.n22147 DVSS.n22122 0.00547368
R61429 DVSS.n938 DVSS.n921 0.00547368
R61430 DVSS.n22433 DVSS.n1000 0.00547368
R61431 DVSS.n22232 DVSS.n465 0.00547368
R61432 DVSS.n22314 DVSS.n1240 0.00547368
R61433 DVSS.n12833 DVSS.n20 0.00547368
R61434 DVSS.n13100 DVSS.n12776 0.00547368
R61435 DVSS.n16267 DVSS.n16247 0.00546098
R61436 DVSS.n16223 DVSS.n16172 0.00546098
R61437 DVSS.n16470 DVSS.n16300 0.00546098
R61438 DVSS.n18088 DVSS.n15635 0.00546098
R61439 DVSS.n16516 DVSS.n16488 0.00545763
R61440 DVSS.n18135 DVSS.n15584 0.00545763
R61441 DVSS.n16594 DVSS.n16346 0.00545
R61442 DVSS.n15964 DVSS.n15942 0.00545
R61443 DVSS.n17711 DVSS.n17675 0.00545
R61444 DVSS.n15217 DVSS.n15170 0.00545
R61445 DVSS.n20762 DVSS.n13707 0.00545
R61446 DVSS.n21212 DVSS.n13635 0.00545
R61447 DVSS.n22646 DVSS.n720 0.00545
R61448 DVSS.n15870 DVSS.n15855 0.00542958
R61449 DVSS.n17919 DVSS.n15762 0.00542958
R61450 DVSS.n16681 DVSS.n16241 0.00538571
R61451 DVSS.n16780 DVSS.n15667 0.00538571
R61452 DVSS.n17642 DVSS.n16087 0.00538571
R61453 DVSS.n17555 DVSS.n16908 0.00538571
R61454 DVSS.n18343 DVSS.n15324 0.00538571
R61455 DVSS.n15475 DVSS.n15451 0.00538571
R61456 DVSS.n20008 DVSS.n14888 0.00538571
R61457 DVSS.n15072 DVSS.n15032 0.00538571
R61458 DVSS.n20849 DVSS.n14459 0.00538571
R61459 DVSS.n20928 DVSS.n20926 0.00538571
R61460 DVSS.n21404 DVSS 0.00538571
R61461 DVSS.n21299 DVSS.n13516 0.00538571
R61462 DVSS.n21382 DVSS.n21376 0.00538571
R61463 DVSS.n22757 DVSS.n596 0.00538571
R61464 DVSS.n22837 DVSS.n532 0.00538571
R61465 DVSS.n22173 DVSS.n1381 0.00537895
R61466 DVSS.n22446 DVSS.n910 0.00537895
R61467 DVSS.n22407 DVSS.n1005 0.00537895
R61468 DVSS.n22288 DVSS.n1255 0.00537895
R61469 DVSS.n12869 DVSS.n27 0.00537895
R61470 DVSS.n12901 DVSS.n12801 0.00537895
R61471 DVSS.n9203 DVSS.n2875 0.00537218
R61472 DVSS.n10503 DVSS.n1612 0.00537218
R61473 DVSS.n15901 DVSS.n15898 0.00536196
R61474 DVSS.n15906 DVSS.n15894 0.00536196
R61475 DVSS.n15860 DVSS.n15853 0.00536196
R61476 DVSS.n17862 DVSS.n15836 0.00536196
R61477 DVSS.n15814 DVSS.n15805 0.00536196
R61478 DVSS.n15819 DVSS.n15801 0.00536196
R61479 DVSS.n15764 DVSS.n15760 0.00536196
R61480 DVSS.n15769 DVSS.n15756 0.00536196
R61481 DVSS.n15724 DVSS.n15696 0.00536196
R61482 DVSS.n15723 DVSS.n15692 0.00536196
R61483 DVSS.n15567 DVSS.n15552 0.00536196
R61484 DVSS.n15568 DVSS.n15548 0.00536196
R61485 DVSS.n15815 DVSS.n15814 0.00536196
R61486 DVSS.n15820 DVSS.n15819 0.00536196
R61487 DVSS.n15765 DVSS.n15764 0.00536196
R61488 DVSS.n15770 DVSS.n15769 0.00536196
R61489 DVSS.n15861 DVSS.n15860 0.00536196
R61490 DVSS.n17863 DVSS.n17862 0.00536196
R61491 DVSS.n15902 DVSS.n15901 0.00536196
R61492 DVSS.n15907 DVSS.n15906 0.00536196
R61493 DVSS.n15725 DVSS.n15696 0.00536196
R61494 DVSS.n18044 DVSS.n15692 0.00536196
R61495 DVSS.n15568 DVSS.n15562 0.00536196
R61496 DVSS.n15567 DVSS.n15559 0.00536196
R61497 DVSS.n18024 DVSS.n15550 0.00535915
R61498 DVSS.n7035 DVSS.n5877 0.00533221
R61499 DVSS.n7825 DVSS.n4472 0.00533221
R61500 DVSS.n7036 DVSS.n5875 0.00533221
R61501 DVSS.n7824 DVSS.n4473 0.00533221
R61502 DVSS.n16746 DVSS.n15597 0.00532143
R61503 DVSS.n15528 DVSS.n15495 0.00532143
R61504 DVSS.n18258 DVSS.n18221 0.00532143
R61505 DVSS.n15122 DVSS.n15105 0.00532143
R61506 DVSS.n20951 DVSS.n14340 0.00532143
R61507 DVSS.n21405 DVSS.n13397 0.00532143
R61508 DVSS.n483 DVSS.n471 0.00532143
R61509 DVSS.n17853 DVSS.n15851 0.00528873
R61510 DVSS.n17935 DVSS.n15758 0.00528873
R61511 DVSS.n22213 DVSS.n706 0.00528421
R61512 DVSS.n22163 DVSS.n1384 0.00528421
R61513 DVSS.n22454 DVSS.n22453 0.00528421
R61514 DVSS.n22417 DVSS.n989 0.00528421
R61515 DVSS.n469 DVSS.n459 0.00528421
R61516 DVSS.n22298 DVSS.n1258 0.00528421
R61517 DVSS.n22332 DVSS.n16 0.00528421
R61518 DVSS.n12911 DVSS.n12798 0.00528421
R61519 DVSS DVSS.n16517 0.00526695
R61520 DVSS.n18134 DVSS 0.00526695
R61521 DVSS.n16320 DVSS.n16307 0.00525714
R61522 DVSS.n16709 DVSS.n16155 0.00525714
R61523 DVSS.n16057 DVSS.n16016 0.00525714
R61524 DVSS.n16874 DVSS.n16839 0.00525714
R61525 DVSS.n15280 DVSS.n15241 0.00525714
R61526 DVSS.n15418 DVSS.n15383 0.00525714
R61527 DVSS.n18424 DVSS.n18383 0.00525714
R61528 DVSS.n14980 DVSS.n14947 0.00525714
R61529 DVSS.n20795 DVSS.n20706 0.00525714
R61530 DVSS.n20878 DVSS.n14428 0.00525714
R61531 DVSS.n13604 DVSS.n13585 0.00525714
R61532 DVSS.n21328 DVSS.n13484 0.00525714
R61533 DVSS.n687 DVSS.n674 0.00525714
R61534 DVSS.n22786 DVSS.n568 0.00525714
R61535 DVSS.n8596 DVSS.n8595 0.005225
R61536 DVSS.n18010 DVSS.n15554 0.00521831
R61537 DVSS.n16638 DVSS.n16313 0.00519756
R61538 DVSS.n16418 DVSS.n16293 0.00519756
R61539 DVSS.n16420 DVSS.n16303 0.00519756
R61540 DVSS.n16422 DVSS.n16294 0.00519756
R61541 DVSS.n16424 DVSS.n16302 0.00519756
R61542 DVSS.n15679 DVSS.n15669 0.00519756
R61543 DVSS.n18078 DVSS.n18077 0.00519756
R61544 DVSS.n18074 DVSS.n15670 0.00519756
R61545 DVSS.n15678 DVSS.n15652 0.00519756
R61546 DVSS.n18081 DVSS.n18080 0.00519756
R61547 DVSS.n16762 DVSS.n15593 0.00519286
R61548 DVSS.n17565 DVSS.n15492 0.00519286
R61549 DVSS.n18232 DVSS.n18218 0.00519286
R61550 DVSS.n19955 DVSS.n15085 0.00519286
R61551 DVSS.n14353 DVSS.n14337 0.00519286
R61552 DVSS.n13411 DVSS.n13394 0.00519286
R61553 DVSS.n488 DVSS.n477 0.00519286
R61554 DVSS.n22219 DVSS.n708 0.00518947
R61555 DVSS.n22157 DVSS.n22125 0.00518947
R61556 DVSS.n928 DVSS.n905 0.00518947
R61557 DVSS.n22423 DVSS.n1003 0.00518947
R61558 DVSS.n22242 DVSS.n468 0.00518947
R61559 DVSS.n22304 DVSS.n1243 0.00518947
R61560 DVSS.n12823 DVSS.n17 0.00518947
R61561 DVSS.n12917 DVSS.n12817 0.00518947
R61562 DVSS.n21458 DVSS.n21457 0.0051875
R61563 DVSS.n22954 DVSS.n428 0.0051875
R61564 DVSS.n17909 DVSS.n17908 0.00514789
R61565 DVSS.n18034 DVSS.n15702 0.00514789
R61566 DVSS.n16614 DVSS.n16311 0.00512857
R61567 DVSS.n16233 DVSS.n16159 0.00512857
R61568 DVSS.n16041 DVSS.n16020 0.00512857
R61569 DVSS.n17618 DVSS.n16141 0.00512857
R61570 DVSS.n17750 DVSS.n15245 0.00512857
R61571 DVSS.n18328 DVSS.n15362 0.00512857
R61572 DVSS.n18474 DVSS.n15234 0.00512857
R61573 DVSS.n19984 DVSS.n14927 0.00512857
R61574 DVSS.n20729 DVSS.n20710 0.00512857
R61575 DVSS.n20862 DVSS.n14432 0.00512857
R61576 DVSS.n21232 DVSS.n13592 0.00512857
R61577 DVSS.n21312 DVSS.n13488 0.00512857
R61578 DVSS.n22690 DVSS.n678 0.00512857
R61579 DVSS.n22770 DVSS.n572 0.00512857
R61580 DVSS.n662 DVSS.n604 0.00510976
R61581 DVSS.n660 DVSS.n558 0.00510976
R61582 DVSS.n665 DVSS.n664 0.00510976
R61583 DVSS.n659 DVSS.n504 0.00510976
R61584 DVSS.n22179 DVSS.n22129 0.00509474
R61585 DVSS.n22451 DVSS.n924 0.00509474
R61586 DVSS.n22401 DVSS.n1009 0.00509474
R61587 DVSS.n22282 DVSS.n1247 0.00509474
R61588 DVSS.n12863 DVSS.n6 0.00509474
R61589 DVSS.n12895 DVSS.n12813 0.00509474
R61590 DVSS.n15891 DVSS.n15878 0.00507746
R61591 DVSS DVSS.n15556 0.00507746
R61592 DVSS.n18985 DVSS.n18872 0.00505056
R61593 DVSS.n20625 DVSS.n14693 0.00505056
R61594 DVSS.n22372 DVSS.n1153 0.00502195
R61595 DVSS.n13088 DVSS.n13063 0.00502195
R61596 DVSS.n22385 DVSS.n1026 0.00502195
R61597 DVSS.n23003 DVSS.n369 0.00502195
R61598 DVSS.n7032 DVSS.n5882 0.00501965
R61599 DVSS.n7031 DVSS.n5884 0.00501965
R61600 DVSS.n15824 DVSS.n15817 0.00500704
R61601 DVSS.n17970 DVSS.n15699 0.00500704
R61602 DVSS.n16326 DVSS.n16311 0.005
R61603 DVSS.n16691 DVSS.n16159 0.005
R61604 DVSS.n16020 DVSS.n15999 0.005
R61605 DVSS.n16141 DVSS.n16137 0.005
R61606 DVSS.n17752 DVSS.n15245 0.005
R61607 DVSS.n15362 DVSS.n15358 0.005
R61608 DVSS.n18475 DVSS.n18474 0.005
R61609 DVSS.n14927 DVSS.n14923 0.005
R61610 DVSS.n20777 DVSS.n20710 0.005
R61611 DVSS.n20860 DVSS.n14432 0.005
R61612 DVSS.n13610 DVSS.n13592 0.005
R61613 DVSS.n21310 DVSS.n13488 0.005
R61614 DVSS.n719 DVSS.n702 0.005
R61615 DVSS.n22141 DVSS.n1388 0.005
R61616 DVSS.n944 DVSS.n918 0.005
R61617 DVSS.n19766 DVSS.n463 0.005
R61618 DVSS.n22320 DVSS.n1262 0.005
R61619 DVSS.n12839 DVSS.n12 0.005
R61620 DVSS.n693 DVSS.n678 0.005
R61621 DVSS.n22768 DVSS.n572 0.005
R61622 DVSS.n16552 DVSS.n16353 0.00498219
R61623 DVSS.n16557 DVSS.n16349 0.00498219
R61624 DVSS.n16316 DVSS.n16309 0.00498219
R61625 DVSS.n16636 DVSS.n16292 0.00498219
R61626 DVSS.n16269 DVSS.n16260 0.00498219
R61627 DVSS.n16274 DVSS.n16256 0.00498219
R61628 DVSS.n16185 DVSS.n16157 0.00498219
R61629 DVSS.n16184 DVSS.n16153 0.00498219
R61630 DVSS.n15676 DVSS.n15659 0.00498219
R61631 DVSS.n15675 DVSS.n15655 0.00498219
R61632 DVSS.n15602 DVSS.n15595 0.00498219
R61633 DVSS.n15606 DVSS.n15591 0.00498219
R61634 DVSS.n17779 DVSS.n15932 0.00498219
R61635 DVSS.n17674 DVSS.n15944 0.00498219
R61636 DVSS.n16023 DVSS.n16018 0.00498219
R61637 DVSS.n16028 DVSS.n16010 0.00498219
R61638 DVSS.n16102 DVSS.n16079 0.00498219
R61639 DVSS.n16101 DVSS.n16075 0.00498219
R61640 DVSS.n16844 DVSS.n16841 0.00498219
R61641 DVSS.n16849 DVSS.n16837 0.00498219
R61642 DVSS.n17604 DVSS.n17546 0.00498219
R61643 DVSS.n17542 DVSS.n17541 0.00498219
R61644 DVSS.n15513 DVSS.n15493 0.00498219
R61645 DVSS.n15514 DVSS.n15497 0.00498219
R61646 DVSS.n17683 DVSS.n17681 0.00498219
R61647 DVSS.n17688 DVSS.n17677 0.00498219
R61648 DVSS.n15272 DVSS.n15243 0.00498219
R61649 DVSS.n15271 DVSS.n15268 0.00498219
R61650 DVSS.n15316 DVSS.n15314 0.00498219
R61651 DVSS.n15321 DVSS.n15310 0.00498219
R61652 DVSS.n15388 DVSS.n15385 0.00498219
R61653 DVSS.n15393 DVSS.n15381 0.00498219
R61654 DVSS.n18314 DVSS.n15466 0.00498219
R61655 DVSS.n15462 DVSS.n15461 0.00498219
R61656 DVSS.n18230 DVSS.n18219 0.00498219
R61657 DVSS.n18225 DVSS.n18223 0.00498219
R61658 DVSS.n18492 DVSS.n15159 0.00498219
R61659 DVSS.n15181 DVSS.n15172 0.00498219
R61660 DVSS.n18388 DVSS.n18385 0.00498219
R61661 DVSS.n18433 DVSS.n18393 0.00498219
R61662 DVSS.n14910 DVSS.n14880 0.00498219
R61663 DVSS.n14909 DVSS.n14876 0.00498219
R61664 DVSS.n14951 DVSS.n14949 0.00498219
R61665 DVSS.n14992 DVSS.n14987 0.00498219
R61666 DVSS.n15024 DVSS.n15023 0.00498219
R61667 DVSS.n15029 DVSS.n15019 0.00498219
R61668 DVSS.n19951 DVSS.n15103 0.00498219
R61669 DVSS.n15109 DVSS.n15107 0.00498219
R61670 DVSS.n21147 DVSS.n13697 0.00498219
R61671 DVSS.n13728 DVSS.n13709 0.00498219
R61672 DVSS.n20714 DVSS.n20708 0.00498219
R61673 DVSS.n20802 DVSS.n20704 0.00498219
R61674 DVSS.n14484 DVSS.n14480 0.00498219
R61675 DVSS.n14489 DVSS.n14476 0.00498219
R61676 DVSS.n14434 DVSS.n14430 0.00498219
R61677 DVSS.n14444 DVSS.n14440 0.00498219
R61678 DVSS.n14384 DVSS.n14382 0.00498219
R61679 DVSS.n14389 DVSS.n14378 0.00498219
R61680 DVSS.n14348 DVSS.n14338 0.00498219
R61681 DVSS.n14343 DVSS.n14320 0.00498219
R61682 DVSS.n13643 DVSS.n13641 0.00498219
R61683 DVSS.n13648 DVSS.n13637 0.00498219
R61684 DVSS.n13596 DVSS.n13587 0.00498219
R61685 DVSS.n21254 DVSS.n13570 0.00498219
R61686 DVSS.n13542 DVSS.n13538 0.00498219
R61687 DVSS.n13553 DVSS.n13548 0.00498219
R61688 DVSS.n13490 DVSS.n13486 0.00498219
R61689 DVSS.n13501 DVSS.n13496 0.00498219
R61690 DVSS.n13443 DVSS.n13441 0.00498219
R61691 DVSS.n13448 DVSS.n13437 0.00498219
R61692 DVSS.n13406 DVSS.n13395 0.00498219
R61693 DVSS.n13401 DVSS.n13377 0.00498219
R61694 DVSS.n13543 DVSS.n13542 0.00498219
R61695 DVSS.n13548 DVSS.n13547 0.00498219
R61696 DVSS.n14485 DVSS.n14484 0.00498219
R61697 DVSS.n14490 DVSS.n14489 0.00498219
R61698 DVSS.n14912 DVSS.n14880 0.00498219
R61699 DVSS.n20006 DVSS.n14876 0.00498219
R61700 DVSS.n15317 DVSS.n15316 0.00498219
R61701 DVSS.n15322 DVSS.n15321 0.00498219
R61702 DVSS.n16103 DVSS.n16079 0.00498219
R61703 DVSS.n17640 DVSS.n16075 0.00498219
R61704 DVSS.n16270 DVSS.n16269 0.00498219
R61705 DVSS.n16275 DVSS.n16274 0.00498219
R61706 DVSS.n13491 DVSS.n13490 0.00498219
R61707 DVSS.n13496 DVSS.n13495 0.00498219
R61708 DVSS.n14435 DVSS.n14434 0.00498219
R61709 DVSS.n14440 DVSS.n14439 0.00498219
R61710 DVSS.n14952 DVSS.n14951 0.00498219
R61711 DVSS.n14987 DVSS.n14956 0.00498219
R61712 DVSS.n15389 DVSS.n15388 0.00498219
R61713 DVSS.n15394 DVSS.n15393 0.00498219
R61714 DVSS.n16845 DVSS.n16844 0.00498219
R61715 DVSS.n16850 DVSS.n16849 0.00498219
R61716 DVSS.n16224 DVSS.n16157 0.00498219
R61717 DVSS.n16822 DVSS.n16153 0.00498219
R61718 DVSS.n21255 DVSS.n21254 0.00498219
R61719 DVSS.n13601 DVSS.n13596 0.00498219
R61720 DVSS.n20715 DVSS.n20714 0.00498219
R61721 DVSS.n20803 DVSS.n20802 0.00498219
R61722 DVSS.n18389 DVSS.n18388 0.00498219
R61723 DVSS.n18399 DVSS.n18393 0.00498219
R61724 DVSS.n18378 DVSS.n15243 0.00498219
R61725 DVSS.n15268 DVSS.n15252 0.00498219
R61726 DVSS.n16024 DVSS.n16023 0.00498219
R61727 DVSS.n16029 DVSS.n16028 0.00498219
R61728 DVSS.n16317 DVSS.n16316 0.00498219
R61729 DVSS.n16637 DVSS.n16636 0.00498219
R61730 DVSS.n13644 DVSS.n13643 0.00498219
R61731 DVSS.n13649 DVSS.n13648 0.00498219
R61732 DVSS.n13714 DVSS.n13697 0.00498219
R61733 DVSS.n13728 DVSS.n13718 0.00498219
R61734 DVSS.n15177 DVSS.n15159 0.00498219
R61735 DVSS.n15182 DVSS.n15181 0.00498219
R61736 DVSS.n17684 DVSS.n17683 0.00498219
R61737 DVSS.n17689 DVSS.n17688 0.00498219
R61738 DVSS.n15949 DVSS.n15932 0.00498219
R61739 DVSS.n17674 DVSS.n15953 0.00498219
R61740 DVSS.n16553 DVSS.n16552 0.00498219
R61741 DVSS.n16558 DVSS.n16557 0.00498219
R61742 DVSS.n13444 DVSS.n13443 0.00498219
R61743 DVSS.n13449 DVSS.n13448 0.00498219
R61744 DVSS.n14385 DVSS.n14384 0.00498219
R61745 DVSS.n14390 DVSS.n14389 0.00498219
R61746 DVSS.n15025 DVSS.n15024 0.00498219
R61747 DVSS.n15030 DVSS.n15029 0.00498219
R61748 DVSS.n15466 DVSS.n15444 0.00498219
R61749 DVSS.n15461 DVSS.n15448 0.00498219
R61750 DVSS.n17546 DVSS.n16901 0.00498219
R61751 DVSS.n17541 DVSS.n16905 0.00498219
R61752 DVSS.n15676 DVSS.n15661 0.00498219
R61753 DVSS.n15675 DVSS.n15665 0.00498219
R61754 DVSS.n15603 DVSS.n15602 0.00498219
R61755 DVSS.n15607 DVSS.n15606 0.00498219
R61756 DVSS.n15514 DVSS.n15499 0.00498219
R61757 DVSS.n15513 DVSS.n15503 0.00498219
R61758 DVSS.n18226 DVSS.n18225 0.00498219
R61759 DVSS.n18231 DVSS.n18230 0.00498219
R61760 DVSS.n15110 DVSS.n15109 0.00498219
R61761 DVSS.n19952 DVSS.n19951 0.00498219
R61762 DVSS.n14344 DVSS.n14343 0.00498219
R61763 DVSS.n14349 DVSS.n14348 0.00498219
R61764 DVSS.n13402 DVSS.n13401 0.00498219
R61765 DVSS.n13407 DVSS.n13406 0.00498219
R61766 DVSS.n727 DVSS.n713 0.00498219
R61767 DVSS.n722 DVSS.n717 0.00498219
R61768 DVSS.n683 DVSS.n676 0.00498219
R61769 DVSS.n22712 DVSS.n648 0.00498219
R61770 DVSS.n625 DVSS.n620 0.00498219
R61771 DVSS.n630 DVSS.n616 0.00498219
R61772 DVSS.n575 DVSS.n570 0.00498219
R61773 DVSS.n580 DVSS.n566 0.00498219
R61774 DVSS.n524 DVSS.n521 0.00498219
R61775 DVSS.n529 DVSS.n517 0.00498219
R61776 DVSS.n480 DVSS.n479 0.00498219
R61777 DVSS.n22877 DVSS.n22876 0.00498219
R61778 DVSS.n22876 DVSS.n458 0.00498219
R61779 DVSS.n479 DVSS.n473 0.00498219
R61780 DVSS.n728 DVSS.n727 0.00498219
R61781 DVSS.n723 DVSS.n722 0.00498219
R61782 DVSS.n684 DVSS.n683 0.00498219
R61783 DVSS.n22713 DVSS.n22712 0.00498219
R61784 DVSS.n626 DVSS.n625 0.00498219
R61785 DVSS.n631 DVSS.n630 0.00498219
R61786 DVSS.n576 DVSS.n575 0.00498219
R61787 DVSS.n581 DVSS.n580 0.00498219
R61788 DVSS.n525 DVSS.n524 0.00498219
R61789 DVSS.n530 DVSS.n529 0.00498219
R61790 DVSS.n17805 DVSS.n15896 0.00493662
R61791 DVSS.n16764 DVSS.n15593 0.00493571
R61792 DVSS.n15511 DVSS.n15492 0.00493571
R61793 DVSS.n18218 DVSS.n15490 0.00493571
R61794 DVSS.n15085 DVSS.n15084 0.00493571
R61795 DVSS.n20975 DVSS.n14337 0.00493571
R61796 DVSS.n21429 DVSS.n13394 0.00493571
R61797 DVSS.n22851 DVSS.n477 0.00493571
R61798 DVSS.n22375 DVSS.n22374 0.00493415
R61799 DVSS.n13060 DVSS.n13001 0.00493415
R61800 DVSS.n22377 DVSS.n1078 0.00493415
R61801 DVSS.n13058 DVSS.n346 0.00493415
R61802 DVSS.n952 DVSS.n901 0.00490526
R61803 DVSS.n992 DVSS.n979 0.00490526
R61804 DVSS.n12847 DVSS.n23 0.00490526
R61805 DVSS.n12879 DVSS.n12805 0.00490526
R61806 DVSS.n17643 DVSS.n16081 0.00489024
R61807 DVSS.n17369 DVSS.n15293 0.00489024
R61808 DVSS.n17470 DVSS.n16148 0.00489024
R61809 DVSS.n17490 DVSS.n15364 0.00489024
R61810 DVSS.n17479 DVSS.n16000 0.00489024
R61811 DVSS.n17378 DVSS.n15255 0.00489024
R61812 DVSS.n17456 DVSS.n16895 0.00489024
R61813 DVSS.n17520 DVSS.n15434 0.00489024
R61814 DVSS.n16627 DVSS.n16307 0.00487143
R61815 DVSS.n16707 DVSS.n16155 0.00487143
R61816 DVSS.n16035 DVSS.n16016 0.00487143
R61817 DVSS.n16872 DVSS.n16839 0.00487143
R61818 DVSS.n18367 DVSS.n15241 0.00487143
R61819 DVSS.n15416 DVSS.n15383 0.00487143
R61820 DVSS.n18405 DVSS.n18383 0.00487143
R61821 DVSS.n14978 DVSS.n14947 0.00487143
R61822 DVSS.n20793 DVSS.n20706 0.00487143
R61823 DVSS.n20876 DVSS.n14428 0.00487143
R61824 DVSS.n21245 DVSS.n13585 0.00487143
R61825 DVSS.n21326 DVSS.n13484 0.00487143
R61826 DVSS.n22703 DVSS.n674 0.00487143
R61827 DVSS.n22784 DVSS.n568 0.00487143
R61828 DVSS.n17875 DVSS.n15811 0.0048662
R61829 DVSS.n9202 DVSS.n9201 0.00484899
R61830 DVSS.n1615 DVSS.n1614 0.00484899
R61831 DVSS.n9205 DVSS.n9204 0.00484899
R61832 DVSS.n10505 DVSS.n10504 0.00484899
R61833 DVSS.n17075 DVSS.n16095 0.00484634
R61834 DVSS.n16843 DVSS.n16150 0.00484634
R61835 DVSS.n16021 DVSS.n16002 0.00484634
R61836 DVSS.n17530 DVSS.n16897 0.00484634
R61837 DVSS.n8983 DVSS.n8982 0.00483083
R61838 DVSS.n11613 DVSS.n11106 0.00483083
R61839 DVSS.n960 DVSS.n916 0.00481053
R61840 DVSS.n22393 DVSS.n993 0.00481053
R61841 DVSS.n12855 DVSS.n24 0.00481053
R61842 DVSS.n12887 DVSS.n12804 0.00481053
R61843 DVSS.n16734 DVSS.n15597 0.00480714
R61844 DVSS.n18187 DVSS.n15495 0.00480714
R61845 DVSS.n18243 DVSS.n18221 0.00480714
R61846 DVSS.n19940 DVSS.n15105 0.00480714
R61847 DVSS.n20953 DVSS.n14340 0.00480714
R61848 DVSS.n21407 DVSS.n13397 0.00480714
R61849 DVSS.n22867 DVSS.n471 0.00480714
R61850 DVSS.n18955 DVSS.n18911 0.00479775
R61851 DVSS.n20156 DVSS.n20049 0.00479775
R61852 DVSS.n20221 DVSS.n20220 0.00479775
R61853 DVSS.n20424 DVSS.n14682 0.00479775
R61854 DVSS.n17805 DVSS.n15904 0.00479577
R61855 DVSS.n10134 DVSS.n10133 0.004775
R61856 DVSS.n10759 DVSS.n10758 0.004775
R61857 DVSS.n13792 DVSS.n13790 0.00476
R61858 DVSS.n13792 DVSS.n13786 0.00476
R61859 DVSS.n13797 DVSS.n13786 0.00476
R61860 DVSS.n13799 DVSS.n13797 0.00476
R61861 DVSS.n13801 DVSS.n13799 0.00476
R61862 DVSS.n13801 DVSS.n13783 0.00476
R61863 DVSS.n13806 DVSS.n13783 0.00476
R61864 DVSS.n13808 DVSS.n13806 0.00476
R61865 DVSS.n13810 DVSS.n13808 0.00476
R61866 DVSS.n13810 DVSS.n13780 0.00476
R61867 DVSS.n21127 DVSS.n13780 0.00476
R61868 DVSS.n21127 DVSS.n21126 0.00476
R61869 DVSS.n21126 DVSS.n21125 0.00476
R61870 DVSS.n21125 DVSS.n21124 0.00476
R61871 DVSS.n21124 DVSS.n13817 0.00476
R61872 DVSS.n21120 DVSS.n13817 0.00476
R61873 DVSS.n21120 DVSS.n21119 0.00476
R61874 DVSS.n21119 DVSS.n21118 0.00476
R61875 DVSS.n21118 DVSS.n13823 0.00476
R61876 DVSS.n13900 DVSS.n13823 0.00476
R61877 DVSS.n13902 DVSS.n13900 0.00476
R61878 DVSS.n13902 DVSS.n13896 0.00476
R61879 DVSS.n13907 DVSS.n13896 0.00476
R61880 DVSS.n13909 DVSS.n13907 0.00476
R61881 DVSS.n13911 DVSS.n13909 0.00476
R61882 DVSS.n13911 DVSS.n13893 0.00476
R61883 DVSS.n13916 DVSS.n13893 0.00476
R61884 DVSS.n13918 DVSS.n13916 0.00476
R61885 DVSS.n13920 DVSS.n13918 0.00476
R61886 DVSS.n13920 DVSS.n13890 0.00476
R61887 DVSS.n21112 DVSS.n13890 0.00476
R61888 DVSS.n21112 DVSS.n21111 0.00476
R61889 DVSS.n21111 DVSS.n21110 0.00476
R61890 DVSS.n21110 DVSS.n13926 0.00476
R61891 DVSS.n13986 DVSS.n13926 0.00476
R61892 DVSS.n13991 DVSS.n13986 0.00476
R61893 DVSS.n13993 DVSS.n13991 0.00476
R61894 DVSS.n13995 DVSS.n13993 0.00476
R61895 DVSS.n13995 DVSS.n13984 0.00476
R61896 DVSS.n14000 DVSS.n13984 0.00476
R61897 DVSS.n14002 DVSS.n14000 0.00476
R61898 DVSS.n14004 DVSS.n14002 0.00476
R61899 DVSS.n14004 DVSS.n13981 0.00476
R61900 DVSS.n21101 DVSS.n13981 0.00476
R61901 DVSS.n21101 DVSS.n21100 0.00476
R61902 DVSS.n21100 DVSS.n21098 0.00476
R61903 DVSS.n21098 DVSS.n21086 0.00476
R61904 DVSS.n21086 DVSS.n21085 0.00476
R61905 DVSS.n21085 DVSS.n21084 0.00476
R61906 DVSS.n21084 DVSS.n14013 0.00476
R61907 DVSS.n21080 DVSS.n14013 0.00476
R61908 DVSS.n21080 DVSS.n21079 0.00476
R61909 DVSS.n21079 DVSS.n21078 0.00476
R61910 DVSS.n21078 DVSS.n14019 0.00476
R61911 DVSS.n14097 DVSS.n14019 0.00476
R61912 DVSS.n14099 DVSS.n14097 0.00476
R61913 DVSS.n14101 DVSS.n14099 0.00476
R61914 DVSS.n14101 DVSS.n14092 0.00476
R61915 DVSS.n14106 DVSS.n14092 0.00476
R61916 DVSS.n14108 DVSS.n14106 0.00476
R61917 DVSS.n14110 DVSS.n14108 0.00476
R61918 DVSS.n14110 DVSS.n14089 0.00476
R61919 DVSS.n14115 DVSS.n14089 0.00476
R61920 DVSS.n14117 DVSS.n14115 0.00476
R61921 DVSS.n14119 DVSS.n14117 0.00476
R61922 DVSS.n14119 DVSS.n14086 0.00476
R61923 DVSS.n21072 DVSS.n14086 0.00476
R61924 DVSS.n21072 DVSS.n21071 0.00476
R61925 DVSS.n21071 DVSS.n21070 0.00476
R61926 DVSS.n21070 DVSS.n14125 0.00476
R61927 DVSS.n14200 DVSS.n14125 0.00476
R61928 DVSS.n14205 DVSS.n14200 0.00476
R61929 DVSS.n14207 DVSS.n14205 0.00476
R61930 DVSS.n14209 DVSS.n14207 0.00476
R61931 DVSS.n14209 DVSS.n14198 0.00476
R61932 DVSS.n14214 DVSS.n14198 0.00476
R61933 DVSS.n14216 DVSS.n14214 0.00476
R61934 DVSS.n14218 DVSS.n14216 0.00476
R61935 DVSS.n14218 DVSS.n14195 0.00476
R61936 DVSS.n14223 DVSS.n14195 0.00476
R61937 DVSS.n14225 DVSS.n14223 0.00476
R61938 DVSS.n14227 DVSS.n14225 0.00476
R61939 DVSS.n14227 DVSS.n14192 0.00476
R61940 DVSS.n21063 DVSS.n14192 0.00476
R61941 DVSS.n21063 DVSS.n21062 0.00476
R61942 DVSS.n21062 DVSS.n21061 0.00476
R61943 DVSS.n21061 DVSS.n14233 0.00476
R61944 DVSS.n21057 DVSS.n14233 0.00476
R61945 DVSS.n21057 DVSS.n21056 0.00476
R61946 DVSS.n21056 DVSS.n14238 0.00476
R61947 DVSS.n14296 DVSS.n14238 0.00476
R61948 DVSS.n21045 DVSS.n14296 0.00476
R61949 DVSS.n21045 DVSS.n21044 0.00476
R61950 DVSS.n21044 DVSS.n21042 0.00476
R61951 DVSS.n21042 DVSS.n21040 0.00476
R61952 DVSS.n21040 DVSS.n21038 0.00476
R61953 DVSS.n21038 DVSS.n21036 0.00476
R61954 DVSS.n21034 DVSS.n21032 0.00476
R61955 DVSS.n21032 DVSS.n21030 0.00476
R61956 DVSS.n21030 DVSS.n21028 0.00476
R61957 DVSS.n13789 DVSS.n13788 0.00476
R61958 DVSS.n21123 DVSS.n13757 0.00476
R61959 DVSS.n21123 DVSS.n21122 0.00476
R61960 DVSS.n21122 DVSS.n21121 0.00476
R61961 DVSS.n21121 DVSS.n13818 0.00476
R61962 DVSS.n21113 DVSS.n13889 0.00476
R61963 DVSS.n21109 DVSS.n13889 0.00476
R61964 DVSS.n21109 DVSS.n21108 0.00476
R61965 DVSS.n21083 DVSS.n13965 0.00476
R61966 DVSS.n21083 DVSS.n21082 0.00476
R61967 DVSS.n21082 DVSS.n21081 0.00476
R61968 DVSS.n21081 DVSS.n14014 0.00476
R61969 DVSS.n21077 DVSS.n14014 0.00476
R61970 DVSS.n21073 DVSS.n14085 0.00476
R61971 DVSS.n21069 DVSS.n14085 0.00476
R61972 DVSS.n21069 DVSS.n21068 0.00476
R61973 DVSS.n21064 DVSS.n14191 0.00476
R61974 DVSS.n21060 DVSS.n14191 0.00476
R61975 DVSS.n21060 DVSS.n21059 0.00476
R61976 DVSS.n21059 DVSS.n21058 0.00476
R61977 DVSS.n21027 DVSS.n21026 0.00476
R61978 DVSS.n21474 DVSS.n987 0.00476
R61979 DVSS.n21502 DVSS.n21501 0.00476
R61980 DVSS.n21510 DVSS.n21509 0.00476
R61981 DVSS.n21511 DVSS.n21510 0.00476
R61982 DVSS.n21543 DVSS.n1083 0.00476
R61983 DVSS.n21544 DVSS.n21543 0.00476
R61984 DVSS.n21545 DVSS.n21544 0.00476
R61985 DVSS.n291 DVSS.n290 0.00476
R61986 DVSS.n294 DVSS.n291 0.00476
R61987 DVSS.n295 DVSS.n294 0.00476
R61988 DVSS.n296 DVSS.n295 0.00476
R61989 DVSS.n297 DVSS.n296 0.00476
R61990 DVSS.n316 DVSS.n315 0.00476
R61991 DVSS.n317 DVSS.n316 0.00476
R61992 DVSS.n382 DVSS.n317 0.00476
R61993 DVSS.n23001 DVSS.n396 0.00476
R61994 DVSS.n402 DVSS.n396 0.00476
R61995 DVSS.n12794 DVSS.n403 0.00476
R61996 DVSS.n22972 DVSS.n421 0.00476
R61997 DVSS.n22570 DVSS.n758 0.00476
R61998 DVSS.n777 DVSS.n776 0.00476
R61999 DVSS.n784 DVSS.n780 0.00476
R62000 DVSS.n785 DVSS.n784 0.00476
R62001 DVSS.n22508 DVSS.n22505 0.00476
R62002 DVSS.n22509 DVSS.n22508 0.00476
R62003 DVSS.n22510 DVSS.n22509 0.00476
R62004 DVSS.n23096 DVSS.n201 0.00476
R62005 DVSS.n23102 DVSS.n201 0.00476
R62006 DVSS.n23103 DVSS.n23102 0.00476
R62007 DVSS.n23105 DVSS.n23103 0.00476
R62008 DVSS.n23105 DVSS.n23104 0.00476
R62009 DVSS.n23141 DVSS.n23139 0.00476
R62010 DVSS.n23141 DVSS.n23140 0.00476
R62011 DVSS.n23140 DVSS.n122 0.00476
R62012 DVSS.n23183 DVSS.n56 0.00476
R62013 DVSS.n23189 DVSS.n56 0.00476
R62014 DVSS.n23192 DVSS.n23191 0.00476
R62015 DVSS.n23222 DVSS.n3 0.00476
R62016 DVSS.n1408 DVSS.n1407 0.00476
R62017 DVSS.n22119 DVSS.n1393 0.00476
R62018 DVSS.n1436 DVSS.n1435 0.00476
R62019 DVSS.n1437 DVSS.n1436 0.00476
R62020 DVSS.n1456 DVSS.n1455 0.00476
R62021 DVSS.n1457 DVSS.n1456 0.00476
R62022 DVSS.n21627 DVSS.n1457 0.00476
R62023 DVSS.n22072 DVSS.n21639 0.00476
R62024 DVSS.n21667 DVSS.n21639 0.00476
R62025 DVSS.n21668 DVSS.n21667 0.00476
R62026 DVSS.n21669 DVSS.n21668 0.00476
R62027 DVSS.n21731 DVSS.n21669 0.00476
R62028 DVSS.n22044 DVSS.n21744 0.00476
R62029 DVSS.n21757 DVSS.n21744 0.00476
R62030 DVSS.n21758 DVSS.n21757 0.00476
R62031 DVSS.n21966 DVSS.n21965 0.00476
R62032 DVSS.n21967 DVSS.n21966 0.00476
R62033 DVSS.n21968 DVSS.n1238 0.00476
R62034 DVSS.n21989 DVSS.n21988 0.00476
R62035 DVSS.n1411 DVSS.n1405 0.00476
R62036 DVSS.n1413 DVSS.n1411 0.00476
R62037 DVSS.n1415 DVSS.n1413 0.00476
R62038 DVSS.n1415 DVSS.n1402 0.00476
R62039 DVSS.n1419 DVSS.n1402 0.00476
R62040 DVSS.n1421 DVSS.n1419 0.00476
R62041 DVSS.n1423 DVSS.n1421 0.00476
R62042 DVSS.n1423 DVSS.n1398 0.00476
R62043 DVSS.n1427 DVSS.n1398 0.00476
R62044 DVSS.n1429 DVSS.n1427 0.00476
R62045 DVSS.n1431 DVSS.n1429 0.00476
R62046 DVSS.n1431 DVSS.n1394 0.00476
R62047 DVSS.n22118 DVSS.n1394 0.00476
R62048 DVSS.n22118 DVSS.n1395 0.00476
R62049 DVSS.n22113 DVSS.n22112 0.00476
R62050 DVSS.n22112 DVSS.n22111 0.00476
R62051 DVSS.n22111 DVSS.n1438 0.00476
R62052 DVSS.n22107 DVSS.n1438 0.00476
R62053 DVSS.n22107 DVSS.n22106 0.00476
R62054 DVSS.n22106 DVSS.n22105 0.00476
R62055 DVSS.n22105 DVSS.n1443 0.00476
R62056 DVSS.n22101 DVSS.n1443 0.00476
R62057 DVSS.n22101 DVSS.n22100 0.00476
R62058 DVSS.n22100 DVSS.n22099 0.00476
R62059 DVSS.n22099 DVSS.n1448 0.00476
R62060 DVSS.n22095 DVSS.n1448 0.00476
R62061 DVSS.n22095 DVSS.n22094 0.00476
R62062 DVSS.n22094 DVSS.n22093 0.00476
R62063 DVSS.n22093 DVSS.n1453 0.00476
R62064 DVSS.n22089 DVSS.n1453 0.00476
R62065 DVSS.n22089 DVSS.n22088 0.00476
R62066 DVSS.n22088 DVSS.n22087 0.00476
R62067 DVSS.n22087 DVSS.n1458 0.00476
R62068 DVSS.n22083 DVSS.n1458 0.00476
R62069 DVSS.n22083 DVSS.n22082 0.00476
R62070 DVSS.n22082 DVSS.n22081 0.00476
R62071 DVSS.n22081 DVSS.n22078 0.00476
R62072 DVSS.n21651 DVSS.n21647 0.00476
R62073 DVSS.n21653 DVSS.n21651 0.00476
R62074 DVSS.n21655 DVSS.n21653 0.00476
R62075 DVSS.n21655 DVSS.n21644 0.00476
R62076 DVSS.n21659 DVSS.n21644 0.00476
R62077 DVSS.n21661 DVSS.n21659 0.00476
R62078 DVSS.n21663 DVSS.n21661 0.00476
R62079 DVSS.n21663 DVSS.n21640 0.00476
R62080 DVSS.n22071 DVSS.n21640 0.00476
R62081 DVSS.n22071 DVSS.n21641 0.00476
R62082 DVSS.n22067 DVSS.n21641 0.00476
R62083 DVSS.n22067 DVSS.n22066 0.00476
R62084 DVSS.n22066 DVSS.n22065 0.00476
R62085 DVSS.n22065 DVSS.n21670 0.00476
R62086 DVSS.n22061 DVSS.n21670 0.00476
R62087 DVSS.n22061 DVSS.n22060 0.00476
R62088 DVSS.n22060 DVSS.n22059 0.00476
R62089 DVSS.n22059 DVSS.n21675 0.00476
R62090 DVSS.n22055 DVSS.n21675 0.00476
R62091 DVSS.n22055 DVSS.n22054 0.00476
R62092 DVSS.n22054 DVSS.n22053 0.00476
R62093 DVSS.n22053 DVSS.n21680 0.00476
R62094 DVSS.n22049 DVSS.n21680 0.00476
R62095 DVSS.n21751 DVSS.n21749 0.00476
R62096 DVSS.n21753 DVSS.n21751 0.00476
R62097 DVSS.n21753 DVSS.n21745 0.00476
R62098 DVSS.n22043 DVSS.n21745 0.00476
R62099 DVSS.n22043 DVSS.n21746 0.00476
R62100 DVSS.n22039 DVSS.n21746 0.00476
R62101 DVSS.n22039 DVSS.n22038 0.00476
R62102 DVSS.n22038 DVSS.n22037 0.00476
R62103 DVSS.n22037 DVSS.n21760 0.00476
R62104 DVSS.n22033 DVSS.n21760 0.00476
R62105 DVSS.n22033 DVSS.n22032 0.00476
R62106 DVSS.n22032 DVSS.n22031 0.00476
R62107 DVSS.n22031 DVSS.n21765 0.00476
R62108 DVSS.n22027 DVSS.n21765 0.00476
R62109 DVSS.n22027 DVSS.n22026 0.00476
R62110 DVSS.n22026 DVSS.n22025 0.00476
R62111 DVSS.n22025 DVSS.n21770 0.00476
R62112 DVSS.n22021 DVSS.n21770 0.00476
R62113 DVSS.n22021 DVSS.n22020 0.00476
R62114 DVSS.n22020 DVSS.n22019 0.00476
R62115 DVSS.n22019 DVSS.n21775 0.00476
R62116 DVSS.n22015 DVSS.n21775 0.00476
R62117 DVSS.n22015 DVSS.n22014 0.00476
R62118 DVSS.n22012 DVSS.n21969 0.00476
R62119 DVSS.n22008 DVSS.n21969 0.00476
R62120 DVSS.n22008 DVSS.n22007 0.00476
R62121 DVSS.n22007 DVSS.n22006 0.00476
R62122 DVSS.n22006 DVSS.n21975 0.00476
R62123 DVSS.n22002 DVSS.n21975 0.00476
R62124 DVSS.n22002 DVSS.n22001 0.00476
R62125 DVSS.n22001 DVSS.n22000 0.00476
R62126 DVSS.n22000 DVSS.n21981 0.00476
R62127 DVSS.n21996 DVSS.n21981 0.00476
R62128 DVSS.n21995 DVSS.n21994 0.00476
R62129 DVSS.n21994 DVSS.n21987 0.00476
R62130 DVSS.n21990 DVSS.n21987 0.00476
R62131 DVSS.n22567 DVSS.n759 0.00476
R62132 DVSS.n22567 DVSS.n22566 0.00476
R62133 DVSS.n22566 DVSS.n22565 0.00476
R62134 DVSS.n22565 DVSS.n764 0.00476
R62135 DVSS.n22561 DVSS.n764 0.00476
R62136 DVSS.n22561 DVSS.n22560 0.00476
R62137 DVSS.n22560 DVSS.n22559 0.00476
R62138 DVSS.n22559 DVSS.n769 0.00476
R62139 DVSS.n22555 DVSS.n769 0.00476
R62140 DVSS.n22555 DVSS.n22554 0.00476
R62141 DVSS.n22554 DVSS.n22553 0.00476
R62142 DVSS.n22553 DVSS.n774 0.00476
R62143 DVSS.n22549 DVSS.n774 0.00476
R62144 DVSS.n22549 DVSS.n22548 0.00476
R62145 DVSS.n22546 DVSS.n781 0.00476
R62146 DVSS.n22542 DVSS.n781 0.00476
R62147 DVSS.n22542 DVSS.n22541 0.00476
R62148 DVSS.n22541 DVSS.n22540 0.00476
R62149 DVSS.n22540 DVSS.n788 0.00476
R62150 DVSS.n22536 DVSS.n788 0.00476
R62151 DVSS.n22536 DVSS.n22535 0.00476
R62152 DVSS.n22535 DVSS.n22534 0.00476
R62153 DVSS.n22534 DVSS.n793 0.00476
R62154 DVSS.n22530 DVSS.n793 0.00476
R62155 DVSS.n22530 DVSS.n22529 0.00476
R62156 DVSS.n22529 DVSS.n22528 0.00476
R62157 DVSS.n22528 DVSS.n798 0.00476
R62158 DVSS.n22524 DVSS.n798 0.00476
R62159 DVSS.n22524 DVSS.n22523 0.00476
R62160 DVSS.n22523 DVSS.n22522 0.00476
R62161 DVSS.n22522 DVSS.n22506 0.00476
R62162 DVSS.n22518 DVSS.n22506 0.00476
R62163 DVSS.n22518 DVSS.n22517 0.00476
R62164 DVSS.n22517 DVSS.n22516 0.00476
R62165 DVSS.n22516 DVSS.n22513 0.00476
R62166 DVSS.n22513 DVSS.n273 0.00476
R62167 DVSS.n23074 DVSS.n273 0.00476
R62168 DVSS.n23079 DVSS.n23077 0.00476
R62169 DVSS.n23079 DVSS.n267 0.00476
R62170 DVSS.n23083 DVSS.n267 0.00476
R62171 DVSS.n23085 DVSS.n23083 0.00476
R62172 DVSS.n23087 DVSS.n23085 0.00476
R62173 DVSS.n23087 DVSS.n264 0.00476
R62174 DVSS.n23091 DVSS.n264 0.00476
R62175 DVSS.n23091 DVSS.n204 0.00476
R62176 DVSS.n23097 DVSS.n204 0.00476
R62177 DVSS.n23097 DVSS.n202 0.00476
R62178 DVSS.n23101 DVSS.n202 0.00476
R62179 DVSS.n23101 DVSS.n200 0.00476
R62180 DVSS.n23106 DVSS.n200 0.00476
R62181 DVSS.n23106 DVSS.n197 0.00476
R62182 DVSS.n23110 DVSS.n197 0.00476
R62183 DVSS.n23112 DVSS.n23110 0.00476
R62184 DVSS.n23114 DVSS.n23112 0.00476
R62185 DVSS.n23114 DVSS.n194 0.00476
R62186 DVSS.n23118 DVSS.n194 0.00476
R62187 DVSS.n23120 DVSS.n23118 0.00476
R62188 DVSS.n23122 DVSS.n23120 0.00476
R62189 DVSS.n23122 DVSS.n190 0.00476
R62190 DVSS.n23126 DVSS.n190 0.00476
R62191 DVSS.n23129 DVSS.n184 0.00476
R62192 DVSS.n23134 DVSS.n184 0.00476
R62193 DVSS.n23134 DVSS.n185 0.00476
R62194 DVSS.n185 DVSS.n124 0.00476
R62195 DVSS.n23142 DVSS.n124 0.00476
R62196 DVSS.n23142 DVSS.n121 0.00476
R62197 DVSS.n23146 DVSS.n121 0.00476
R62198 DVSS.n23148 DVSS.n23146 0.00476
R62199 DVSS.n23150 DVSS.n23148 0.00476
R62200 DVSS.n23150 DVSS.n118 0.00476
R62201 DVSS.n23154 DVSS.n118 0.00476
R62202 DVSS.n23156 DVSS.n23154 0.00476
R62203 DVSS.n23158 DVSS.n23156 0.00476
R62204 DVSS.n23158 DVSS.n114 0.00476
R62205 DVSS.n23162 DVSS.n114 0.00476
R62206 DVSS.n23164 DVSS.n23162 0.00476
R62207 DVSS.n23174 DVSS.n23164 0.00476
R62208 DVSS.n23174 DVSS.n111 0.00476
R62209 DVSS.n23178 DVSS.n111 0.00476
R62210 DVSS.n23178 DVSS.n59 0.00476
R62211 DVSS.n23184 DVSS.n59 0.00476
R62212 DVSS.n23184 DVSS.n57 0.00476
R62213 DVSS.n23188 DVSS.n57 0.00476
R62214 DVSS.n23193 DVSS.n50 0.00476
R62215 DVSS.n23197 DVSS.n50 0.00476
R62216 DVSS.n23199 DVSS.n23197 0.00476
R62217 DVSS.n23201 DVSS.n23199 0.00476
R62218 DVSS.n23201 DVSS.n47 0.00476
R62219 DVSS.n23205 DVSS.n47 0.00476
R62220 DVSS.n23207 DVSS.n23205 0.00476
R62221 DVSS.n23209 DVSS.n23207 0.00476
R62222 DVSS.n23209 DVSS.n44 0.00476
R62223 DVSS.n23214 DVSS.n44 0.00476
R62224 DVSS.n23214 DVSS.n0 0.00476
R62225 DVSS.n23227 DVSS.n2 0.00476
R62226 DVSS.n23223 DVSS.n2 0.00476
R62227 DVSS.n21477 DVSS.n21476 0.00476
R62228 DVSS.n21479 DVSS.n21477 0.00476
R62229 DVSS.n21479 DVSS.n1497 0.00476
R62230 DVSS.n21483 DVSS.n1497 0.00476
R62231 DVSS.n21485 DVSS.n21483 0.00476
R62232 DVSS.n21487 DVSS.n21485 0.00476
R62233 DVSS.n21487 DVSS.n1493 0.00476
R62234 DVSS.n21491 DVSS.n1493 0.00476
R62235 DVSS.n21493 DVSS.n21491 0.00476
R62236 DVSS.n21495 DVSS.n21493 0.00476
R62237 DVSS.n21495 DVSS.n1489 0.00476
R62238 DVSS.n21499 DVSS.n1489 0.00476
R62239 DVSS.n21500 DVSS.n21499 0.00476
R62240 DVSS.n21503 DVSS.n21500 0.00476
R62241 DVSS.n21508 DVSS.n1483 0.00476
R62242 DVSS.n21512 DVSS.n1483 0.00476
R62243 DVSS.n21514 DVSS.n21512 0.00476
R62244 DVSS.n21514 DVSS.n1480 0.00476
R62245 DVSS.n21518 DVSS.n1480 0.00476
R62246 DVSS.n21520 DVSS.n21518 0.00476
R62247 DVSS.n21522 DVSS.n21520 0.00476
R62248 DVSS.n21522 DVSS.n1476 0.00476
R62249 DVSS.n21526 DVSS.n1476 0.00476
R62250 DVSS.n21528 DVSS.n21526 0.00476
R62251 DVSS.n21530 DVSS.n21528 0.00476
R62252 DVSS.n21530 DVSS.n1472 0.00476
R62253 DVSS.n21534 DVSS.n1472 0.00476
R62254 DVSS.n21536 DVSS.n21534 0.00476
R62255 DVSS.n21537 DVSS.n21536 0.00476
R62256 DVSS.n21537 DVSS.n1469 0.00476
R62257 DVSS.n21542 DVSS.n1469 0.00476
R62258 DVSS.n21542 DVSS.n1468 0.00476
R62259 DVSS.n21546 DVSS.n1468 0.00476
R62260 DVSS.n21548 DVSS.n21546 0.00476
R62261 DVSS.n21548 DVSS.n1465 0.00476
R62262 DVSS.n21552 DVSS.n1465 0.00476
R62263 DVSS.n21553 DVSS.n21552 0.00476
R62264 DVSS.n23069 DVSS.n23068 0.00476
R62265 DVSS.n23068 DVSS.n23067 0.00476
R62266 DVSS.n23067 DVSS.n282 0.00476
R62267 DVSS.n23063 DVSS.n282 0.00476
R62268 DVSS.n23063 DVSS.n23062 0.00476
R62269 DVSS.n23062 DVSS.n23061 0.00476
R62270 DVSS.n23061 DVSS.n287 0.00476
R62271 DVSS.n23057 DVSS.n287 0.00476
R62272 DVSS.n23057 DVSS.n23056 0.00476
R62273 DVSS.n23056 DVSS.n23055 0.00476
R62274 DVSS.n23055 DVSS.n292 0.00476
R62275 DVSS.n23051 DVSS.n292 0.00476
R62276 DVSS.n23051 DVSS.n23050 0.00476
R62277 DVSS.n23050 DVSS.n23049 0.00476
R62278 DVSS.n23049 DVSS.n298 0.00476
R62279 DVSS.n23045 DVSS.n298 0.00476
R62280 DVSS.n23045 DVSS.n23044 0.00476
R62281 DVSS.n23044 DVSS.n23043 0.00476
R62282 DVSS.n23043 DVSS.n303 0.00476
R62283 DVSS.n23039 DVSS.n303 0.00476
R62284 DVSS.n23039 DVSS.n23038 0.00476
R62285 DVSS.n23038 DVSS.n23037 0.00476
R62286 DVSS.n23037 DVSS.n308 0.00476
R62287 DVSS.n23032 DVSS.n23031 0.00476
R62288 DVSS.n23031 DVSS.n23030 0.00476
R62289 DVSS.n23030 DVSS.n313 0.00476
R62290 DVSS.n23026 DVSS.n313 0.00476
R62291 DVSS.n23026 DVSS.n23025 0.00476
R62292 DVSS.n23025 DVSS.n23024 0.00476
R62293 DVSS.n23024 DVSS.n318 0.00476
R62294 DVSS.n23020 DVSS.n318 0.00476
R62295 DVSS.n23020 DVSS.n23019 0.00476
R62296 DVSS.n23019 DVSS.n23018 0.00476
R62297 DVSS.n23018 DVSS.n323 0.00476
R62298 DVSS.n23014 DVSS.n323 0.00476
R62299 DVSS.n23014 DVSS.n23013 0.00476
R62300 DVSS.n23013 DVSS.n23012 0.00476
R62301 DVSS.n23012 DVSS.n328 0.00476
R62302 DVSS.n23008 DVSS.n328 0.00476
R62303 DVSS.n23008 DVSS.n23007 0.00476
R62304 DVSS.n23007 DVSS.n23006 0.00476
R62305 DVSS.n23006 DVSS.n333 0.00476
R62306 DVSS.n397 DVSS.n333 0.00476
R62307 DVSS.n23000 DVSS.n397 0.00476
R62308 DVSS.n23000 DVSS.n398 0.00476
R62309 DVSS.n22996 DVSS.n398 0.00476
R62310 DVSS.n22994 DVSS.n404 0.00476
R62311 DVSS.n22990 DVSS.n404 0.00476
R62312 DVSS.n22990 DVSS.n22989 0.00476
R62313 DVSS.n22989 DVSS.n22988 0.00476
R62314 DVSS.n22988 DVSS.n409 0.00476
R62315 DVSS.n22984 DVSS.n409 0.00476
R62316 DVSS.n22984 DVSS.n22983 0.00476
R62317 DVSS.n22983 DVSS.n22982 0.00476
R62318 DVSS.n22982 DVSS.n414 0.00476
R62319 DVSS.n22978 DVSS.n414 0.00476
R62320 DVSS.n22977 DVSS.n22976 0.00476
R62321 DVSS.n22976 DVSS.n419 0.00476
R62322 DVSS.n420 DVSS.n419 0.00476
R62323 DVSS.n16680 DVSS.n16251 0.00475854
R62324 DVSS.n21827 DVSS.n602 0.00475854
R62325 DVSS.n16823 DVSS.n16176 0.00475854
R62326 DVSS.n21834 DVSS.n554 0.00475854
R62327 DVSS.n21830 DVSS.n655 0.00475854
R62328 DVSS.n21829 DVSS.n502 0.00475854
R62329 DVSS.n16682 DVSS.n16681 0.00474286
R62330 DVSS.n16778 DVSS.n15667 0.00474286
R62331 DVSS.n17642 DVSS.n16093 0.00474286
R62332 DVSS.n17579 DVSS.n16908 0.00474286
R62333 DVSS.n18343 DVSS.n18342 0.00474286
R62334 DVSS.n18289 DVSS.n15451 0.00474286
R62335 DVSS.n20008 DVSS.n14894 0.00474286
R62336 DVSS.n15074 DVSS.n15032 0.00474286
R62337 DVSS.n20850 DVSS.n20849 0.00474286
R62338 DVSS.n20928 DVSS.n20927 0.00474286
R62339 DVSS.n21300 DVSS.n21299 0.00474286
R62340 DVSS.n21382 DVSS.n21381 0.00474286
R62341 DVSS.n22758 DVSS.n22757 0.00474286
R62342 DVSS.n22837 DVSS.n22836 0.00474286
R62343 DVSS.n15824 DVSS.n15803 0.00472535
R62344 DVSS.n17970 DVSS.n15694 0.00472535
R62345 DVSS.n22227 DVSS.n703 0.00471579
R62346 DVSS.n22149 DVSS.n1387 0.00471579
R62347 DVSS.n936 DVSS.n903 0.00471579
R62348 DVSS.n22434 DVSS.n1012 0.00471579
R62349 DVSS.n22234 DVSS.n462 0.00471579
R62350 DVSS.n22312 DVSS.n1261 0.00471579
R62351 DVSS.n12831 DVSS.n13 0.00471579
R62352 DVSS.n13097 DVSS.n12795 0.00471579
R62353 DVSS.n21155 DVSS.n13684 0.00468605
R62354 DVSS.n16346 DVSS.n16334 0.00467857
R62355 DVSS DVSS.n15599 0.00467857
R62356 DVSS.n15955 DVSS.n15942 0.00467857
R62357 DVSS DVSS.n15500 0.00467857
R62358 DVSS.n17691 DVSS.n17675 0.00467857
R62359 DVSS DVSS.n18227 0.00467857
R62360 DVSS.n15184 DVSS.n15170 0.00467857
R62361 DVSS DVSS.n15111 0.00467857
R62362 DVSS.n13720 DVSS.n13707 0.00467857
R62363 DVSS DVSS.n14345 0.00467857
R62364 DVSS.n13635 DVSS.n13618 0.00467857
R62365 DVSS DVSS.n13403 0.00467857
R62366 DVSS.n720 DVSS.n701 0.00467857
R62367 DVSS.n22874 DVSS 0.00467857
R62368 DVSS.n22074 DVSS.n21629 0.00467073
R62369 DVSS.n22046 DVSS.n21733 0.00467073
R62370 DVSS.n21946 DVSS.n21850 0.00467073
R62371 DVSS.n21963 DVSS.n21950 0.00467073
R62372 DVSS.n17823 DVSS.n15878 0.00465493
R62373 DVSS.n14794 DVSS 0.00464676
R62374 DVSS.n3750 DVSS.n3502 0.00462664
R62375 DVSS.n8598 DVSS.n8597 0.00462664
R62376 DVSS.n22171 DVSS.n22128 0.00462105
R62377 DVSS.n22444 DVSS.n914 0.00462105
R62378 DVSS.n22409 DVSS.n995 0.00462105
R62379 DVSS.n22290 DVSS.n1246 0.00462105
R62380 DVSS.n28 DVSS.n5 0.00462105
R62381 DVSS.n12903 DVSS.n12814 0.00462105
R62382 DVSS.n16280 DVSS.n16272 0.00461429
R62383 DVSS.n16794 DVSS.n15663 0.00461429
R62384 DVSS.n16126 DVSS.n16084 0.00461429
R62385 DVSS.n17595 DVSS.n16903 0.00461429
R62386 DVSS.n15341 DVSS.n15319 0.00461429
R62387 DVSS.n18305 DVSS.n15446 0.00461429
R62388 DVSS.n18447 DVSS.n14885 0.00461429
R62389 DVSS.n15041 DVSS.n15027 0.00461429
R62390 DVSS.n14495 DVSS.n14487 0.00461429
R62391 DVSS.n20911 DVSS.n14387 0.00461429
R62392 DVSS.n13558 DVSS.n13545 0.00461429
R62393 DVSS.n21361 DVSS.n13446 0.00461429
R62394 DVSS.n636 DVSS.n628 0.00461429
R62395 DVSS.n22819 DVSS.n527 0.00461429
R62396 DVSS DVSS.n18824 0.00460473
R62397 DVSS.n17949 DVSS.n15734 0.00458451
R62398 DVSS.n18034 DVSS.n15690 0.00458451
R62399 DVSS.n13016 DVSS.n1143 0.00458293
R62400 DVSS.n13022 DVSS.n13020 0.00458293
R62401 DVSS.n13015 DVSS.n1088 0.00458293
R62402 DVSS.n13014 DVSS.n356 0.00458293
R62403 DVSS.n22978 DVSS 0.00458
R62404 DVSS.n16579 DVSS.n16351 0.00455
R62405 DVSS.n15967 DVSS.n15946 0.00455
R62406 DVSS.n17714 DVSS.n17679 0.00455
R62407 DVSS.n15199 DVSS.n15174 0.00455
R62408 DVSS.n20748 DVSS.n13711 0.00455
R62409 DVSS.n21192 DVSS.n13639 0.00455
R62410 DVSS.n22660 DVSS.n715 0.00455
R62411 DVSS.n22211 DVSS.n707 0.00452632
R62412 DVSS.n22165 DVSS.n22126 0.00452632
R62413 DVSS.n22415 DVSS.n1010 0.00452632
R62414 DVSS.n22878 DVSS.n476 0.00452632
R62415 DVSS.n22296 DVSS.n1244 0.00452632
R62416 DVSS.n12909 DVSS.n12816 0.00452632
R62417 DVSS.n18010 DVSS.n15557 0.00451408
R62418 DVSS.n23072 DVSS.n276 0.0045
R62419 DVSS.n21681 DVSS.n186 0.0045
R62420 DVSS.n21505 DVSS.n782 0.0045
R62421 DVSS.n23072 DVSS.n23071 0.0045
R62422 DVSS.n23034 DVSS.n186 0.0045
R62423 DVSS.n21970 DVSS.n52 0.0045
R62424 DVSS.n401 DVSS.n52 0.0045
R62425 DVSS.n22115 DVSS.n782 0.0045
R62426 DVSS.n16649 DVSS.n16266 0.00448571
R62427 DVSS.n17645 DVSS.n17644 0.00448571
R62428 DVSS.n18352 DVSS.n15286 0.00448571
R62429 DVSS.n18464 DVSS.n14882 0.00448571
R62430 DVSS.n20818 DVSS.n20814 0.00448571
R62431 DVSS.n21267 DVSS.n13540 0.00448571
R62432 DVSS.n22725 DVSS.n622 0.00448571
R62433 DVSS.n15132 DVSS.n15131 0.00448437
R62434 DVSS.n21005 DVSS.n21004 0.00448437
R62435 DVSS.n16494 DVSS.n15886 0.00447895
R62436 DVSS.n16496 DVSS.n15881 0.00447895
R62437 DVSS.n16498 DVSS.n15885 0.00447895
R62438 DVSS.n16500 DVSS.n15882 0.00447895
R62439 DVSS.n16502 DVSS.n15884 0.00447895
R62440 DVSS.n16504 DVSS.n15883 0.00447895
R62441 DVSS.n18153 DVSS.n15547 0.00447895
R62442 DVSS.n18152 DVSS.n15555 0.00447895
R62443 DVSS.n15577 DVSS.n15566 0.00447895
R62444 DVSS.n15579 DVSS.n15574 0.00447895
R62445 DVSS.n15575 DVSS.n15565 0.00447895
R62446 DVSS.n18148 DVSS.n18147 0.00447895
R62447 DVSS.n17853 DVSS.n15863 0.00444366
R62448 DVSS.n17935 DVSS.n15767 0.00444366
R62449 DVSS.n22221 DVSS.n705 0.00443158
R62450 DVSS.n22155 DVSS.n1385 0.00443158
R62451 DVSS.n930 DVSS.n919 0.00443158
R62452 DVSS.n22425 DVSS.n997 0.00443158
R62453 DVSS.n22240 DVSS.n460 0.00443158
R62454 DVSS.n22306 DVSS.n1259 0.00443158
R62455 DVSS.n12825 DVSS.n15 0.00443158
R62456 DVSS.n12919 DVSS.n12797 0.00443158
R62457 DVSS.n16579 DVSS.n16555 0.00442143
R62458 DVSS.n15967 DVSS.n15951 0.00442143
R62459 DVSS.n17714 DVSS.n17686 0.00442143
R62460 DVSS.n15199 DVSS.n15179 0.00442143
R62461 DVSS.n20748 DVSS.n13716 0.00442143
R62462 DVSS.n21192 DVSS.n13646 0.00442143
R62463 DVSS.n22660 DVSS.n725 0.00442143
R62464 DVSS.n15315 DVSS.n15297 0.00440732
R62465 DVSS.n623 DVSS.n605 0.00440732
R62466 DVSS.n15387 DVSS.n15367 0.00440732
R62467 DVSS.n573 DVSS.n559 0.00440732
R62468 DVSS.n15273 DVSS.n15258 0.00440732
R62469 DVSS.n680 DVSS.n666 0.00440732
R62470 DVSS.n15452 DVSS.n15437 0.00440732
R62471 DVSS.n523 DVSS.n505 0.00440732
R62472 DVSS.n18024 DVSS.n15561 0.00437324
R62473 DVSS.n8980 DVSS.n3044 0.00436577
R62474 DVSS.n11615 DVSS.n11108 0.00436577
R62475 DVSS.n8981 DVSS.n3047 0.00436577
R62476 DVSS.n11614 DVSS.n11107 0.00436577
R62477 DVSS.n16280 DVSS.n16258 0.00435714
R62478 DVSS.n16794 DVSS.n15657 0.00435714
R62479 DVSS.n16126 DVSS.n16077 0.00435714
R62480 DVSS.n17595 DVSS.n17544 0.00435714
R62481 DVSS.n15341 DVSS.n15312 0.00435714
R62482 DVSS.n18305 DVSS.n15464 0.00435714
R62483 DVSS.n18447 DVSS.n14878 0.00435714
R62484 DVSS.n15041 DVSS.n15021 0.00435714
R62485 DVSS.n14495 DVSS.n14478 0.00435714
R62486 DVSS.n20911 DVSS.n14380 0.00435714
R62487 DVSS.n13558 DVSS.n13536 0.00435714
R62488 DVSS.n21361 DVSS.n13439 0.00435714
R62489 DVSS.n636 DVSS.n618 0.00435714
R62490 DVSS.n22819 DVSS.n519 0.00435714
R62491 DVSS.n22182 DVSS.n1380 0.00433684
R62492 DVSS.n966 DVSS.n900 0.00433684
R62493 DVSS.n22399 DVSS.n991 0.00433684
R62494 DVSS.n22280 DVSS.n1254 0.00433684
R62495 DVSS.n12861 DVSS.n26 0.00433684
R62496 DVSS.n12893 DVSS.n12802 0.00433684
R62497 DVSS.n7837 DVSS.n4458 0.004325
R62498 DVSS.n21938 DVSS.n21601 0.00431951
R62499 DVSS.n21935 DVSS.n21704 0.00431951
R62500 DVSS.n21941 DVSS.n21940 0.00431951
R62501 DVSS.n21934 DVSS.n21797 0.00431951
R62502 DVSS.n15870 DVSS.n15858 0.00430282
R62503 DVSS.n16597 DVSS.n16334 0.00429286
R62504 DVSS.n17777 DVSS.n15955 0.00429286
R62505 DVSS.n17774 DVSS.n17691 0.00429286
R62506 DVSS.n18490 DVSS.n15184 0.00429286
R62507 DVSS.n21145 DVSS.n13720 0.00429286
R62508 DVSS.n21215 DVSS.n13618 0.00429286
R62509 DVSS.n22673 DVSS.n701 0.00429286
R62510 DVSS.n18914 DVSS.n18876 0.00429213
R62511 DVSS.n20094 DVSS.n20058 0.00429213
R62512 DVSS.n20143 DVSS.n20061 0.00429213
R62513 DVSS.n20284 DVSS.n20217 0.00429213
R62514 DVSS.n20306 DVSS.n20305 0.00429213
R62515 DVSS.n20385 DVSS.n14687 0.00429213
R62516 DVSS.n16548 DVSS.n16344 0.00428947
R62517 DVSS.n7082 DVSS.n5179 0.00428947
R62518 DVSS.n7448 DVSS.n7447 0.00428947
R62519 DVSS.n18112 DVSS.n18111 0.00428947
R62520 DVSS.n22672 DVSS.n712 0.00424211
R62521 DVSS.n22139 DVSS.n22121 0.00424211
R62522 DVSS.n946 DVSS.n907 0.00424211
R62523 DVSS.n19769 DVSS.n464 0.00424211
R62524 DVSS.n22323 DVSS.n1239 0.00424211
R62525 DVSS.n12841 DVSS.n21 0.00424211
R62526 DVSS.n10131 DVSS.n2413 0.00423362
R62527 DVSS.n10756 DVSS.n1522 0.00423362
R62528 DVSS.n10132 DVSS.n10130 0.00423362
R62529 DVSS.n10757 DVSS.n1520 0.00423362
R62530 DVSS.n246 DVSS.n217 0.00423171
R62531 DVSS.n13051 DVSS.n1131 0.00423171
R62532 DVSS.n166 DVSS.n137 0.00423171
R62533 DVSS.n13055 DVSS.n12997 0.00423171
R62534 DVSS.n22482 DVSS.n813 0.00423171
R62535 DVSS.n13050 DVSS.n1074 0.00423171
R62536 DVSS.n101 DVSS.n72 0.00423171
R62537 DVSS.n13049 DVSS.n342 0.00423171
R62538 DVSS.n16824 DVSS.n16171 0.00422857
R62539 DVSS.n16778 DVSS.n15653 0.00422857
R62540 DVSS.n17615 DVSS.n17614 0.00422857
R62541 DVSS.n17579 DVSS.n17535 0.00422857
R62542 DVSS.n18325 DVSS.n18324 0.00422857
R62543 DVSS.n18289 DVSS.n15456 0.00422857
R62544 DVSS.n19981 DVSS.n19980 0.00422857
R62545 DVSS.n15074 DVSS.n15017 0.00422857
R62546 DVSS.n20890 DVSS.n14406 0.00422857
R62547 DVSS.n20927 DVSS.n14361 0.00422857
R62548 DVSS.n21340 DVSS.n13461 0.00422857
R62549 DVSS.n21381 DVSS.n13419 0.00422857
R62550 DVSS.n22798 DVSS.n543 0.00422857
R62551 DVSS.n22836 DVSS.n512 0.00422857
R62552 DVSS.n20043 DVSS.n13927 0.00418781
R62553 DVSS.n21075 DVSS.n14074 0.00418781
R62554 DVSS.n16383 DVSS.n15845 0.00418781
R62555 DVSS.n16384 DVSS.n15839 0.00418781
R62556 DVSS.n16386 DVSS.n15843 0.00418781
R62557 DVSS.n16388 DVSS.n15840 0.00418781
R62558 DVSS.n16390 DVSS.n15842 0.00418781
R62559 DVSS.n16393 DVSS.n15841 0.00418781
R62560 DVSS.n21115 DVSS.n13879 0.00418781
R62561 DVSS.n15719 DVSS.n15718 0.00418781
R62562 DVSS.n15716 DVSS.n15706 0.00418781
R62563 DVSS.n15714 DVSS.n15710 0.00418781
R62564 DVSS.n15712 DVSS.n15707 0.00418781
R62565 DVSS.n15709 DVSS.n15689 0.00418781
R62566 DVSS.n18048 DVSS.n18047 0.00418781
R62567 DVSS.n21066 DVSS.n14180 0.00418781
R62568 DVSS.n16734 DVSS.n15600 0.00416429
R62569 DVSS.n18187 DVSS.n15501 0.00416429
R62570 DVSS.n18243 DVSS.n18228 0.00416429
R62571 DVSS.n19940 DVSS.n15112 0.00416429
R62572 DVSS.n20953 DVSS.n14346 0.00416429
R62573 DVSS.n21407 DVSS.n13404 0.00416429
R62574 DVSS.n22867 DVSS.n482 0.00416429
R62575 DVSS.n17840 DVSS.n15859 0.00416197
R62576 DVSS.n17921 DVSS.n15763 0.00416197
R62577 DVSS.n13906 DVSS.n13883 0.00416
R62578 DVSS.n14100 DVSS.n14078 0.00416
R62579 DVSS.n1475 DVSS.n1063 0.00416
R62580 DVSS.n12984 DVSS.n302 0.00416
R62581 DVSS.n22489 DVSS.n792 0.00416
R62582 DVSS.n193 DVSS.n170 0.00416
R62583 DVSS.n21865 DVSS.n1445 0.00416
R62584 DVSS.n21738 DVSS.n21737 0.00416
R62585 DVSS.n22135 DVSS.n1392 0.00414737
R62586 DVSS.n950 DVSS.n922 0.00414737
R62587 DVSS.n22437 DVSS.n22436 0.00414737
R62588 DVSS.n22327 DVSS.n1221 0.00414737
R62589 DVSS.n12845 DVSS.n10 0.00414737
R62590 DVSS.n12877 DVSS.n12809 0.00414737
R62591 DVSS.n17099 DVSS.n16067 0.0041439
R62592 DVSS.n17616 DVSS.n16827 0.0041439
R62593 DVSS.n17654 DVSS.n16005 0.0041439
R62594 DVSS.n17605 DVSS.n16900 0.0041439
R62595 DVSS.n21043 DVSS.n14262 0.00413
R62596 DVSS.n12790 DVSS.n411 0.00413
R62597 DVSS.n48 DVSS.n41 0.00413
R62598 DVSS.n21977 DVSS.n1235 0.00413
R62599 DVSS.n16627 DVSS.n16319 0.0041
R62600 DVSS.n16707 DVSS.n16162 0.0041
R62601 DVSS.n16035 DVSS.n16026 0.0041
R62602 DVSS.n16872 DVSS.n16847 0.0041
R62603 DVSS.n18367 DVSS.n15250 0.0041
R62604 DVSS.n15416 DVSS.n15391 0.0041
R62605 DVSS.n18405 DVSS.n18391 0.0041
R62606 DVSS.n14978 DVSS.n14954 0.0041
R62607 DVSS.n20793 DVSS.n20717 0.0041
R62608 DVSS.n20876 DVSS.n14437 0.0041
R62609 DVSS.n21114 DVSS.n13888 0.0041
R62610 DVSS.n14116 DVSS.n14083 0.0041
R62611 DVSS.n21245 DVSS.n13603 0.0041
R62612 DVSS.n21326 DVSS.n13493 0.0041
R62613 DVSS.n22703 DVSS.n686 0.0041
R62614 DVSS.n22784 DVSS.n578 0.0041
R62615 DVSS.n22379 DVSS.n1067 0.0041
R62616 DVSS.n12989 DVSS.n311 0.0041
R62617 DVSS.n22504 DVSS.n801 0.0041
R62618 DVSS.n23136 DVSS.n183 0.0041
R62619 DVSS.n21944 DVSS.n21870 0.0041
R62620 DVSS.n21750 DVSS.n21742 0.0041
R62621 DVSS.n18022 DVSS.n15560 0.00409155
R62622 DVSS.n21029 DVSS.n14258 0.00407
R62623 DVSS.n12785 DVSS.n12784 0.00407
R62624 DVSS.n23221 DVSS.n4 0.00407
R62625 DVSS.n21986 DVSS.n1231 0.00407
R62626 DVSS.n16426 DVSS.n16242 0.0040561
R62627 DVSS.n16220 DVSS.n16166 0.0040561
R62628 DVSS.n22185 DVSS.n1370 0.00405263
R62629 DVSS.n962 DVSS.n909 0.00405263
R62630 DVSS.n22395 DVSS.n1006 0.00405263
R62631 DVSS.n22276 DVSS.n1251 0.00405263
R62632 DVSS.n12857 DVSS.n8 0.00405263
R62633 DVSS.n12889 DVSS.n12811 0.00405263
R62634 DVSS.n21102 DVSS.n13942 0.00404
R62635 DVSS.n14217 DVSS.n14176 0.00404
R62636 DVSS.n1110 DVSS.n285 0.00404
R62637 DVSS.n391 DVSS.n378 0.00404
R62638 DVSS.n403 DVSS.n55 0.00404
R62639 DVSS.n23086 DVSS.n240 0.00404
R62640 DVSS.n115 DVSS.n96 0.00404
R62641 DVSS.n23192 DVSS.n23190 0.00404
R62642 DVSS.n21645 DVSS.n21623 0.00404
R62643 DVSS.n21820 DVSS.n21768 0.00404
R62644 DVSS.n21968 DVSS.n54 0.00404
R62645 DVSS.n22013 DVSS.n22012 0.00404
R62646 DVSS.n23193 DVSS.n53 0.00404
R62647 DVSS.n22995 DVSS.n22994 0.00404
R62648 DVSS.n16764 DVSS.n15605 0.00403571
R62649 DVSS.n18205 DVSS.n15511 0.00403571
R62650 DVSS.n18276 DVSS.n15490 0.00403571
R62651 DVSS.n15084 DVSS.n15080 0.00403571
R62652 DVSS.n20976 DVSS.n20975 0.00403571
R62653 DVSS.n21430 DVSS.n21429 0.00403571
R62654 DVSS.n22851 DVSS.n475 0.00403571
R62655 DVSS.n17860 DVSS.n15864 0.00402113
R62656 DVSS.n17937 DVSS.n15768 0.00402113
R62657 DVSS.n16463 DVSS.n16360 0.0040122
R62658 DVSS.n15644 DVSS.n15629 0.0040122
R62659 DVSS.n13807 DVSS.n13741 0.00401
R62660 DVSS.n1494 DVSS.n983 0.00401
R62661 DVSS.n895 DVSS.n894 0.00401
R62662 DVSS.n1397 DVSS.n1375 0.00401
R62663 DVSS.n13992 DVSS.n13946 0.00398
R62664 DVSS.n21067 DVSS.n14138 0.00398
R62665 DVSS.n1466 DVSS.n1114 0.00398
R62666 DVSS.n383 DVSS.n320 0.00398
R62667 DVSS.n272 DVSS.n244 0.00398
R62668 DVSS.n23147 DVSS.n100 0.00398
R62669 DVSS.n21626 DVSS.n1462 0.00398
R62670 DVSS.n21824 DVSS.n21759 0.00398
R62671 DVSS.n16326 DVSS.n16314 0.00397143
R62672 DVSS.n17655 DVSS.n15999 0.00397143
R62673 DVSS.n17752 DVSS.n15247 0.00397143
R62674 DVSS.n18475 DVSS.n15228 0.00397143
R62675 DVSS.n20777 DVSS.n20712 0.00397143
R62676 DVSS.n13610 DVSS.n13594 0.00397143
R62677 DVSS.n693 DVSS.n681 0.00397143
R62678 DVSS.n21916 DVSS.n21599 0.00396829
R62679 DVSS.n854 DVSS.n227 0.00396829
R62680 DVSS.n21913 DVSS.n21702 0.00396829
R62681 DVSS.n852 DVSS.n147 0.00396829
R62682 DVSS.n21919 DVSS.n21918 0.00396829
R62683 DVSS.n857 DVSS.n856 0.00396829
R62684 DVSS.n21912 DVSS.n21795 0.00396829
R62685 DVSS.n851 DVSS.n82 0.00396829
R62686 DVSS.n22225 DVSS.n710 0.00395789
R62687 DVSS.n22151 DVSS.n22123 0.00395789
R62688 DVSS.n934 DVSS.n920 0.00395789
R62689 DVSS.n22431 DVSS.n988 0.00395789
R62690 DVSS.n22236 DVSS.n466 0.00395789
R62691 DVSS.n22310 DVSS.n1241 0.00395789
R62692 DVSS.n12829 DVSS.n19 0.00395789
R62693 DVSS.n13098 DVSS.n12819 0.00395789
R62694 DVSS.n18008 DVSS.n15556 0.0039507
R62695 DVSS.n13791 DVSS.n13736 0.00395
R62696 DVSS.n13785 DVSS.n13734 0.00395
R62697 DVSS.n22435 DVSS.n1001 0.00395
R62698 DVSS.n21478 DVSS.n973 0.00395
R62699 DVSS.n22452 DVSS.n761 0.00395
R62700 DVSS.n883 DVSS.n762 0.00395
R62701 DVSS.n1406 DVSS.n1371 0.00395
R62702 DVSS.n1412 DVSS.n1368 0.00395
R62703 DVSS.n15890 DVSS.n15887 0.00393493
R62704 DVSS.n15892 DVSS.n15880 0.00393493
R62705 DVSS.n15889 DVSS.n15886 0.00393493
R62706 DVSS.n16347 DVSS.n16339 0.00393493
R62707 DVSS.n16345 DVSS.n15937 0.00393493
R62708 DVSS.n15943 DVSS.n15927 0.00393493
R62709 DVSS.n15941 DVSS.n15936 0.00393493
R62710 DVSS.n15959 DVSS.n15928 0.00393493
R62711 DVSS.n15940 DVSS.n15935 0.00393493
R62712 DVSS.n15960 DVSS.n15929 0.00393493
R62713 DVSS.n15939 DVSS.n15934 0.00393493
R62714 DVSS.n15961 DVSS.n15930 0.00393493
R62715 DVSS.n15938 DVSS.n15933 0.00393493
R62716 DVSS.n15962 DVSS.n15931 0.00393493
R62717 DVSS.n17776 DVSS.n15957 0.00393493
R62718 DVSS.n17692 DVSS.n17676 0.00393493
R62719 DVSS.n17773 DVSS.n17705 0.00393493
R62720 DVSS.n17772 DVSS.n17693 0.00393493
R62721 DVSS.n17704 DVSS.n17703 0.00393493
R62722 DVSS.n17707 DVSS.n17694 0.00393493
R62723 DVSS.n17702 DVSS.n17701 0.00393493
R62724 DVSS.n17708 DVSS.n17695 0.00393493
R62725 DVSS.n17700 DVSS.n17699 0.00393493
R62726 DVSS.n17709 DVSS.n17697 0.00393493
R62727 DVSS.n17696 DVSS.n15164 0.00393493
R62728 DVSS.n15171 DVSS.n15154 0.00393493
R62729 DVSS.n15169 DVSS.n15163 0.00393493
R62730 DVSS.n15210 DVSS.n15155 0.00393493
R62731 DVSS.n15168 DVSS.n15162 0.00393493
R62732 DVSS.n15211 DVSS.n15156 0.00393493
R62733 DVSS.n15167 DVSS.n15161 0.00393493
R62734 DVSS.n15212 DVSS.n15157 0.00393493
R62735 DVSS.n15166 DVSS.n15160 0.00393493
R62736 DVSS.n15213 DVSS.n15158 0.00393493
R62737 DVSS.n15165 DVSS.n13702 0.00393493
R62738 DVSS.n13708 DVSS.n13692 0.00393493
R62739 DVSS.n13706 DVSS.n13701 0.00393493
R62740 DVSS.n13723 DVSS.n13693 0.00393493
R62741 DVSS.n13705 DVSS.n13700 0.00393493
R62742 DVSS.n13724 DVSS.n13694 0.00393493
R62743 DVSS.n13704 DVSS.n13699 0.00393493
R62744 DVSS.n13725 DVSS.n13695 0.00393493
R62745 DVSS.n13703 DVSS.n13698 0.00393493
R62746 DVSS.n13726 DVSS.n13696 0.00393493
R62747 DVSS.n21144 DVSS.n13722 0.00393493
R62748 DVSS.n13746 DVSS.n13729 0.00393493
R62749 DVSS.n21141 DVSS.n13778 0.00393493
R62750 DVSS.n21140 DVSS.n13747 0.00393493
R62751 DVSS.n13777 DVSS.n13776 0.00393493
R62752 DVSS.n21129 DVSS.n13748 0.00393493
R62753 DVSS.n13775 DVSS.n13774 0.00393493
R62754 DVSS.n21130 DVSS.n13749 0.00393493
R62755 DVSS.n13773 DVSS.n13772 0.00393493
R62756 DVSS.n21131 DVSS.n13750 0.00393493
R62757 DVSS.n13771 DVSS.n13770 0.00393493
R62758 DVSS.n21132 DVSS.n13751 0.00393493
R62759 DVSS.n13769 DVSS.n13768 0.00393493
R62760 DVSS.n21133 DVSS.n13752 0.00393493
R62761 DVSS.n13767 DVSS.n13766 0.00393493
R62762 DVSS.n21134 DVSS.n13753 0.00393493
R62763 DVSS.n13765 DVSS.n13764 0.00393493
R62764 DVSS.n21135 DVSS.n13754 0.00393493
R62765 DVSS.n13763 DVSS.n13762 0.00393493
R62766 DVSS.n21136 DVSS.n13755 0.00393493
R62767 DVSS.n13761 DVSS.n13760 0.00393493
R62768 DVSS.n21137 DVSS.n13756 0.00393493
R62769 DVSS.n13759 DVSS.n13758 0.00393493
R62770 DVSS.n21138 DVSS.n13629 0.00393493
R62771 DVSS.n13636 DVSS.n13619 0.00393493
R62772 DVSS.n13634 DVSS.n13628 0.00393493
R62773 DVSS.n21201 DVSS.n13620 0.00393493
R62774 DVSS.n13633 DVSS.n13627 0.00393493
R62775 DVSS.n21202 DVSS.n13621 0.00393493
R62776 DVSS.n13632 DVSS.n13626 0.00393493
R62777 DVSS.n21203 DVSS.n13622 0.00393493
R62778 DVSS.n13631 DVSS.n13625 0.00393493
R62779 DVSS.n21204 DVSS.n13623 0.00393493
R62780 DVSS.n13630 DVSS.n13624 0.00393493
R62781 DVSS.n13630 DVSS.n13623 0.00393493
R62782 DVSS.n21204 DVSS.n13625 0.00393493
R62783 DVSS.n13631 DVSS.n13622 0.00393493
R62784 DVSS.n21203 DVSS.n13626 0.00393493
R62785 DVSS.n13632 DVSS.n13621 0.00393493
R62786 DVSS.n21202 DVSS.n13627 0.00393493
R62787 DVSS.n13633 DVSS.n13620 0.00393493
R62788 DVSS.n21201 DVSS.n13628 0.00393493
R62789 DVSS.n13634 DVSS.n13619 0.00393493
R62790 DVSS.n21214 DVSS.n13636 0.00393493
R62791 DVSS.n21138 DVSS.n13759 0.00393493
R62792 DVSS.n13758 DVSS.n13756 0.00393493
R62793 DVSS.n21137 DVSS.n13761 0.00393493
R62794 DVSS.n13760 DVSS.n13755 0.00393493
R62795 DVSS.n21136 DVSS.n13763 0.00393493
R62796 DVSS.n13762 DVSS.n13754 0.00393493
R62797 DVSS.n21135 DVSS.n13765 0.00393493
R62798 DVSS.n13764 DVSS.n13753 0.00393493
R62799 DVSS.n21134 DVSS.n13767 0.00393493
R62800 DVSS.n13766 DVSS.n13752 0.00393493
R62801 DVSS.n21133 DVSS.n13769 0.00393493
R62802 DVSS.n13768 DVSS.n13751 0.00393493
R62803 DVSS.n21132 DVSS.n13771 0.00393493
R62804 DVSS.n13770 DVSS.n13750 0.00393493
R62805 DVSS.n21131 DVSS.n13773 0.00393493
R62806 DVSS.n13772 DVSS.n13749 0.00393493
R62807 DVSS.n21130 DVSS.n13775 0.00393493
R62808 DVSS.n13774 DVSS.n13748 0.00393493
R62809 DVSS.n21129 DVSS.n13777 0.00393493
R62810 DVSS.n13776 DVSS.n13747 0.00393493
R62811 DVSS.n21141 DVSS.n21140 0.00393493
R62812 DVSS.n13778 DVSS.n13746 0.00393493
R62813 DVSS.n21143 DVSS.n13729 0.00393493
R62814 DVSS.n13722 DVSS.n13696 0.00393493
R62815 DVSS.n13726 DVSS.n13698 0.00393493
R62816 DVSS.n13703 DVSS.n13695 0.00393493
R62817 DVSS.n13725 DVSS.n13699 0.00393493
R62818 DVSS.n13704 DVSS.n13694 0.00393493
R62819 DVSS.n13724 DVSS.n13700 0.00393493
R62820 DVSS.n13705 DVSS.n13693 0.00393493
R62821 DVSS.n13723 DVSS.n13701 0.00393493
R62822 DVSS.n13706 DVSS.n13692 0.00393493
R62823 DVSS.n21146 DVSS.n13708 0.00393493
R62824 DVSS.n15165 DVSS.n15158 0.00393493
R62825 DVSS.n15213 DVSS.n15160 0.00393493
R62826 DVSS.n15166 DVSS.n15157 0.00393493
R62827 DVSS.n15212 DVSS.n15161 0.00393493
R62828 DVSS.n15167 DVSS.n15156 0.00393493
R62829 DVSS.n15211 DVSS.n15162 0.00393493
R62830 DVSS.n15168 DVSS.n15155 0.00393493
R62831 DVSS.n15210 DVSS.n15163 0.00393493
R62832 DVSS.n15169 DVSS.n15154 0.00393493
R62833 DVSS.n18491 DVSS.n15171 0.00393493
R62834 DVSS.n17697 DVSS.n17696 0.00393493
R62835 DVSS.n17709 DVSS.n17700 0.00393493
R62836 DVSS.n17699 DVSS.n17695 0.00393493
R62837 DVSS.n17708 DVSS.n17702 0.00393493
R62838 DVSS.n17701 DVSS.n17694 0.00393493
R62839 DVSS.n17707 DVSS.n17704 0.00393493
R62840 DVSS.n17703 DVSS.n17693 0.00393493
R62841 DVSS.n17773 DVSS.n17772 0.00393493
R62842 DVSS.n17705 DVSS.n17692 0.00393493
R62843 DVSS.n17775 DVSS.n17676 0.00393493
R62844 DVSS.n15957 DVSS.n15931 0.00393493
R62845 DVSS.n15962 DVSS.n15933 0.00393493
R62846 DVSS.n15938 DVSS.n15930 0.00393493
R62847 DVSS.n15961 DVSS.n15934 0.00393493
R62848 DVSS.n15939 DVSS.n15929 0.00393493
R62849 DVSS.n15960 DVSS.n15935 0.00393493
R62850 DVSS.n15940 DVSS.n15928 0.00393493
R62851 DVSS.n15959 DVSS.n15936 0.00393493
R62852 DVSS.n15941 DVSS.n15927 0.00393493
R62853 DVSS.n17778 DVSS.n15943 0.00393493
R62854 DVSS.n16345 DVSS.n16339 0.00393493
R62855 DVSS.n16347 DVSS.n16340 0.00393493
R62856 DVSS.n15889 DVSS.n15880 0.00393493
R62857 DVSS.n15892 DVSS.n15887 0.00393493
R62858 DVSS.n15890 DVSS.n15879 0.00393493
R62859 DVSS.n18149 DVSS.n15569 0.00393493
R62860 DVSS.n15573 DVSS.n15571 0.00393493
R62861 DVSS.n15572 DVSS.n15547 0.00393493
R62862 DVSS.n18115 DVSS.n15609 0.00393493
R62863 DVSS.n18118 DVSS.n18117 0.00393493
R62864 DVSS.n15512 DVSS.n15510 0.00393493
R62865 DVSS.n18198 DVSS.n15517 0.00393493
R62866 DVSS.n15516 DVSS.n15509 0.00393493
R62867 DVSS.n18199 DVSS.n15519 0.00393493
R62868 DVSS.n15518 DVSS.n15508 0.00393493
R62869 DVSS.n18200 DVSS.n15521 0.00393493
R62870 DVSS.n15520 DVSS.n15507 0.00393493
R62871 DVSS.n18204 DVSS.n18202 0.00393493
R62872 DVSS.n18203 DVSS.n15506 0.00393493
R62873 DVSS.n18206 DVSS.n15491 0.00393493
R62874 DVSS.n18217 DVSS.n15489 0.00393493
R62875 DVSS.n18233 DVSS.n18208 0.00393493
R62876 DVSS.n18216 DVSS.n15488 0.00393493
R62877 DVSS.n18234 DVSS.n18209 0.00393493
R62878 DVSS.n18215 DVSS.n15487 0.00393493
R62879 DVSS.n18235 DVSS.n18210 0.00393493
R62880 DVSS.n18214 DVSS.n15486 0.00393493
R62881 DVSS.n18236 DVSS.n18211 0.00393493
R62882 DVSS.n18213 DVSS.n15485 0.00393493
R62883 DVSS.n18275 DVSS.n18212 0.00393493
R62884 DVSS.n15092 DVSS.n15090 0.00393493
R62885 DVSS.n15114 DVSS.n15095 0.00393493
R62886 DVSS.n15094 DVSS.n15089 0.00393493
R62887 DVSS.n15115 DVSS.n15097 0.00393493
R62888 DVSS.n15096 DVSS.n15088 0.00393493
R62889 DVSS.n15116 DVSS.n15099 0.00393493
R62890 DVSS.n15098 DVSS.n15087 0.00393493
R62891 DVSS.n15117 DVSS.n15101 0.00393493
R62892 DVSS.n15100 DVSS.n15086 0.00393493
R62893 DVSS.n19953 DVSS.n15102 0.00393493
R62894 DVSS.n14336 DVSS.n14325 0.00393493
R62895 DVSS.n20964 DVSS.n14327 0.00393493
R62896 DVSS.n14335 DVSS.n14324 0.00393493
R62897 DVSS.n20965 DVSS.n14328 0.00393493
R62898 DVSS.n14334 DVSS.n14323 0.00393493
R62899 DVSS.n20966 DVSS.n14329 0.00393493
R62900 DVSS.n14333 DVSS.n14322 0.00393493
R62901 DVSS.n20967 DVSS.n14330 0.00393493
R62902 DVSS.n14332 DVSS.n14321 0.00393493
R62903 DVSS.n20977 DVSS.n14331 0.00393493
R62904 DVSS.n14278 DVSS.n14240 0.00393493
R62905 DVSS.n14295 DVSS.n14273 0.00393493
R62906 DVSS.n14279 DVSS.n14241 0.00393493
R62907 DVSS.n14294 DVSS.n14272 0.00393493
R62908 DVSS.n14280 DVSS.n14242 0.00393493
R62909 DVSS.n14293 DVSS.n14271 0.00393493
R62910 DVSS.n14281 DVSS.n14243 0.00393493
R62911 DVSS.n14292 DVSS.n14270 0.00393493
R62912 DVSS.n14282 DVSS.n14244 0.00393493
R62913 DVSS.n14291 DVSS.n14269 0.00393493
R62914 DVSS.n14283 DVSS.n14245 0.00393493
R62915 DVSS.n14290 DVSS.n14268 0.00393493
R62916 DVSS.n14284 DVSS.n14246 0.00393493
R62917 DVSS.n14289 DVSS.n14267 0.00393493
R62918 DVSS.n14285 DVSS.n14247 0.00393493
R62919 DVSS.n14288 DVSS.n14266 0.00393493
R62920 DVSS.n14286 DVSS.n14248 0.00393493
R62921 DVSS.n14287 DVSS.n14265 0.00393493
R62922 DVSS.n21049 DVSS.n14249 0.00393493
R62923 DVSS.n21048 DVSS.n14264 0.00393493
R62924 DVSS.n21050 DVSS.n14250 0.00393493
R62925 DVSS.n21052 DVSS.n14252 0.00393493
R62926 DVSS.n21053 DVSS.n14251 0.00393493
R62927 DVSS.n13393 DVSS.n13382 0.00393493
R62928 DVSS.n21418 DVSS.n13384 0.00393493
R62929 DVSS.n13392 DVSS.n13381 0.00393493
R62930 DVSS.n21419 DVSS.n13385 0.00393493
R62931 DVSS.n13391 DVSS.n13380 0.00393493
R62932 DVSS.n21420 DVSS.n13386 0.00393493
R62933 DVSS.n13390 DVSS.n13379 0.00393493
R62934 DVSS.n21421 DVSS.n13387 0.00393493
R62935 DVSS.n13389 DVSS.n13378 0.00393493
R62936 DVSS.n21431 DVSS.n13388 0.00393493
R62937 DVSS.n15571 DVSS.n15569 0.00393493
R62938 DVSS.n15573 DVSS.n15572 0.00393493
R62939 DVSS.n18116 DVSS.n18115 0.00393493
R62940 DVSS.n18117 DVSS.n15609 0.00393493
R62941 DVSS.n15515 DVSS.n15512 0.00393493
R62942 DVSS.n18198 DVSS.n15510 0.00393493
R62943 DVSS.n15517 DVSS.n15516 0.00393493
R62944 DVSS.n18199 DVSS.n15509 0.00393493
R62945 DVSS.n15519 DVSS.n15518 0.00393493
R62946 DVSS.n18200 DVSS.n15508 0.00393493
R62947 DVSS.n15521 DVSS.n15520 0.00393493
R62948 DVSS.n18202 DVSS.n15507 0.00393493
R62949 DVSS.n18204 DVSS.n18203 0.00393493
R62950 DVSS.n15506 DVSS.n15491 0.00393493
R62951 DVSS.n18217 DVSS.n18207 0.00393493
R62952 DVSS.n18233 DVSS.n15489 0.00393493
R62953 DVSS.n18216 DVSS.n18208 0.00393493
R62954 DVSS.n18234 DVSS.n15488 0.00393493
R62955 DVSS.n18215 DVSS.n18209 0.00393493
R62956 DVSS.n18235 DVSS.n15487 0.00393493
R62957 DVSS.n18214 DVSS.n18210 0.00393493
R62958 DVSS.n18236 DVSS.n15486 0.00393493
R62959 DVSS.n18213 DVSS.n18211 0.00393493
R62960 DVSS.n18212 DVSS.n15485 0.00393493
R62961 DVSS.n15093 DVSS.n15092 0.00393493
R62962 DVSS.n15114 DVSS.n15090 0.00393493
R62963 DVSS.n15095 DVSS.n15094 0.00393493
R62964 DVSS.n15115 DVSS.n15089 0.00393493
R62965 DVSS.n15097 DVSS.n15096 0.00393493
R62966 DVSS.n15116 DVSS.n15088 0.00393493
R62967 DVSS.n15099 DVSS.n15098 0.00393493
R62968 DVSS.n15117 DVSS.n15087 0.00393493
R62969 DVSS.n15101 DVSS.n15100 0.00393493
R62970 DVSS.n15102 DVSS.n15086 0.00393493
R62971 DVSS.n14336 DVSS.n14326 0.00393493
R62972 DVSS.n20964 DVSS.n14325 0.00393493
R62973 DVSS.n14335 DVSS.n14327 0.00393493
R62974 DVSS.n20965 DVSS.n14324 0.00393493
R62975 DVSS.n14334 DVSS.n14328 0.00393493
R62976 DVSS.n20966 DVSS.n14323 0.00393493
R62977 DVSS.n14333 DVSS.n14329 0.00393493
R62978 DVSS.n20967 DVSS.n14322 0.00393493
R62979 DVSS.n14332 DVSS.n14330 0.00393493
R62980 DVSS.n14331 DVSS.n14321 0.00393493
R62981 DVSS.n14276 DVSS.n14240 0.00393493
R62982 DVSS.n14295 DVSS.n14278 0.00393493
R62983 DVSS.n14273 DVSS.n14241 0.00393493
R62984 DVSS.n14294 DVSS.n14279 0.00393493
R62985 DVSS.n14272 DVSS.n14242 0.00393493
R62986 DVSS.n14293 DVSS.n14280 0.00393493
R62987 DVSS.n14271 DVSS.n14243 0.00393493
R62988 DVSS.n14292 DVSS.n14281 0.00393493
R62989 DVSS.n14270 DVSS.n14244 0.00393493
R62990 DVSS.n14291 DVSS.n14282 0.00393493
R62991 DVSS.n14269 DVSS.n14245 0.00393493
R62992 DVSS.n14290 DVSS.n14283 0.00393493
R62993 DVSS.n14268 DVSS.n14246 0.00393493
R62994 DVSS.n14289 DVSS.n14284 0.00393493
R62995 DVSS.n14267 DVSS.n14247 0.00393493
R62996 DVSS.n14288 DVSS.n14285 0.00393493
R62997 DVSS.n14266 DVSS.n14248 0.00393493
R62998 DVSS.n14287 DVSS.n14286 0.00393493
R62999 DVSS.n14265 DVSS.n14249 0.00393493
R63000 DVSS.n21049 DVSS.n21048 0.00393493
R63001 DVSS.n14264 DVSS.n14250 0.00393493
R63002 DVSS.n21050 DVSS.n14252 0.00393493
R63003 DVSS.n21053 DVSS.n21052 0.00393493
R63004 DVSS.n13393 DVSS.n13383 0.00393493
R63005 DVSS.n21418 DVSS.n13382 0.00393493
R63006 DVSS.n13392 DVSS.n13384 0.00393493
R63007 DVSS.n21419 DVSS.n13381 0.00393493
R63008 DVSS.n13391 DVSS.n13385 0.00393493
R63009 DVSS.n21420 DVSS.n13380 0.00393493
R63010 DVSS.n13390 DVSS.n13386 0.00393493
R63011 DVSS.n21421 DVSS.n13379 0.00393493
R63012 DVSS.n13389 DVSS.n13387 0.00393493
R63013 DVSS.n13388 DVSS.n13378 0.00393493
R63014 DVSS.n18150 DVSS.n18149 0.00393493
R63015 DVSS.n21036 DVSS 0.00392
R63016 DVSS.n13994 DVSS.n13949 0.00392
R63017 DVSS.n14204 DVSS.n14183 0.00392
R63018 DVSS.n387 DVSS.n321 0.00392
R63019 DVSS.n23149 DVSS.n104 0.00392
R63020 DVSS.n21954 DVSS.n21953 0.00392
R63021 DVSS.n21996 DVSS 0.00392
R63022 DVSS.n13809 DVSS.n13730 0.00389
R63023 DVSS.n21492 DVSS.n977 0.00389
R63024 DVSS.n887 DVSS.n771 0.00389
R63025 DVSS.n1399 DVSS.n1364 0.00389
R63026 DVSS.n7080 DVSS.n5181 0.00388255
R63027 DVSS.n7450 DVSS.n4834 0.00388255
R63028 DVSS.n7081 DVSS.n5180 0.00388255
R63029 DVSS.n7449 DVSS.n4836 0.00388255
R63030 DVSS.n819 DVSS.n219 0.00388049
R63031 DVSS.n13030 DVSS.n1148 0.00388049
R63032 DVSS.n816 DVSS.n139 0.00388049
R63033 DVSS.n13036 DVSS.n13034 0.00388049
R63034 DVSS.n822 DVSS.n821 0.00388049
R63035 DVSS.n13029 DVSS.n1093 0.00388049
R63036 DVSS.n815 DVSS.n74 0.00388049
R63037 DVSS.n13028 DVSS.n361 0.00388049
R63038 DVSS.n15800 DVSS.n15785 0.00388028
R63039 DVSS.n18036 DVSS.n15691 0.00388028
R63040 DVSS.n22169 DVSS.n1382 0.00386316
R63041 DVSS.n22442 DVSS.n913 0.00386316
R63042 DVSS.n22411 DVSS.n1004 0.00386316
R63043 DVSS.n22292 DVSS.n1256 0.00386316
R63044 DVSS.n23220 DVSS.n36 0.00386316
R63045 DVSS.n12905 DVSS.n12800 0.00386316
R63046 DVSS.n21099 DVSS.n13952 0.00386
R63047 DVSS.n14194 DVSS.n14188 0.00386
R63048 DVSS.n1124 DVSS.n286 0.00386
R63049 DVSS.n394 DVSS.n330 0.00386
R63050 DVSS.n23093 DVSS.n263 0.00386
R63051 DVSS.n23163 DVSS.n109 0.00386
R63052 DVSS.n21660 DVSS.n21637 0.00386
R63053 DVSS.n21961 DVSS.n21769 0.00386
R63054 DVSS.n16614 DVSS.n16315 0.00384286
R63055 DVSS.n16233 DVSS.n16160 0.00384286
R63056 DVSS.n16041 DVSS.n16022 0.00384286
R63057 DVSS.n17618 DVSS.n17617 0.00384286
R63058 DVSS.n17750 DVSS.n15248 0.00384286
R63059 DVSS.n18328 DVSS.n18327 0.00384286
R63060 DVSS.n18387 DVSS.n15234 0.00384286
R63061 DVSS.n19984 DVSS.n19983 0.00384286
R63062 DVSS.n20729 DVSS.n20713 0.00384286
R63063 DVSS.n20862 DVSS.n14433 0.00384286
R63064 DVSS.n21232 DVSS.n13595 0.00384286
R63065 DVSS.n21312 DVSS.n13489 0.00384286
R63066 DVSS.n22690 DVSS.n682 0.00384286
R63067 DVSS.n22770 DVSS.n574 0.00384286
R63068 DVSS.n7840 DVSS.n7839 0.00384061
R63069 DVSS.n7838 DVSS.n4459 0.00384061
R63070 DVSS.n21031 DVSS.n14256 0.00383
R63071 DVSS.n12782 DVSS.n418 0.00383
R63072 DVSS.n21985 DVSS.n1229 0.00383
R63073 DVSS.n17821 DVSS.n17820 0.00380986
R63074 DVSS.n13919 DVSS.n13873 0.0038
R63075 DVSS.n14114 DVSS.n14069 0.0038
R63076 DVSS.n21535 DVSS.n1053 0.0038
R63077 DVSS.n12974 DVSS.n310 0.0038
R63078 DVSS.n22498 DVSS.n800 0.0038
R63079 DVSS.n23128 DVSS.n160 0.0038
R63080 DVSS.n21852 DVSS.n1452 0.0038
R63081 DVSS.n22047 DVSS.n21694 0.0038
R63082 DVSS.n21749 DVSS.n187 0.0038
R63083 DVSS.n23129 DVSS.n23127 0.0038
R63084 DVSS.n23032 DVSS.n188 0.0038
R63085 DVSS.n18897 DVSS.n18882 0.00378652
R63086 DVSS.n20338 DVSS.n20337 0.00378652
R63087 DVSS.n16762 DVSS.n15604 0.00377857
R63088 DVSS.n17565 DVSS.n15504 0.00377857
R63089 DVSS.n18274 DVSS.n18232 0.00377857
R63090 DVSS.n19955 DVSS.n19954 0.00377857
R63091 DVSS.n14353 DVSS.n14350 0.00377857
R63092 DVSS.n13411 DVSS.n13408 0.00377857
R63093 DVSS.n488 DVSS.n478 0.00377857
R63094 DVSS.n21047 DVSS.n21046 0.00377
R63095 DVSS.n12791 DVSS.n12778 0.00377
R63096 DVSS.n46 DVSS.n34 0.00377
R63097 DVSS.n21974 DVSS.n1225 0.00377
R63098 DVSS.n22167 DVSS.n1383 0.00376842
R63099 DVSS.n22413 DVSS.n990 0.00376842
R63100 DVSS.n22294 DVSS.n1257 0.00376842
R63101 DVSS.n12907 DVSS.n12799 0.00376842
R63102 DVSS.n8610 DVSS.n8609 0.00374812
R63103 DVSS.n13127 DVSS.n13126 0.00374812
R63104 DVSS.n13103 DVSS.n13102 0.00374812
R63105 DVSS.n13895 DVSS.n13877 0.00374
R63106 DVSS.n14098 DVSS.n14073 0.00374
R63107 DVSS.n21521 DVSS.n1057 0.00374
R63108 DVSS.n12978 DVSS.n301 0.00374
R63109 DVSS.n22476 DVSS.n791 0.00374
R63110 DVSS.n23113 DVSS.n164 0.00374
R63111 DVSS.n21862 DVSS.n21856 0.00374
R63112 DVSS.n21730 DVSS.n21674 0.00374
R63113 DVSS.n17888 DVSS.n15804 0.00373944
R63114 DVSS.n17968 DVSS.n15695 0.00373944
R63115 DVSS.n15796 DVSS.n15787 0.00372031
R63116 DVSS.n15797 DVSS.n15788 0.00372031
R63117 DVSS.n15798 DVSS.n15789 0.00372031
R63118 DVSS.n15799 DVSS.n15790 0.00372031
R63119 DVSS.n16252 DVSS.n16244 0.00372031
R63120 DVSS.n16253 DVSS.n16245 0.00372031
R63121 DVSS.n16254 DVSS.n16096 0.00372031
R63122 DVSS.n16100 DVSS.n16070 0.00372031
R63123 DVSS.n16097 DVSS.n16090 0.00372031
R63124 DVSS.n16098 DVSS.n16094 0.00372031
R63125 DVSS.n17643 DVSS.n16074 0.00372031
R63126 DVSS.n15308 DVSS.n15302 0.00372031
R63127 DVSS.n15307 DVSS.n15300 0.00372031
R63128 DVSS.n14907 DVSS.n14902 0.00372031
R63129 DVSS.n14906 DVSS.n14900 0.00372031
R63130 DVSS.n14905 DVSS.n14898 0.00372031
R63131 DVSS.n14904 DVSS.n14896 0.00372031
R63132 DVSS.n20009 DVSS.n14875 0.00372031
R63133 DVSS.n14474 DVSS.n14469 0.00372031
R63134 DVSS.n14473 DVSS.n14468 0.00372031
R63135 DVSS.n14472 DVSS.n14467 0.00372031
R63136 DVSS.n14471 DVSS.n14466 0.00372031
R63137 DVSS.n20048 DVSS.n20041 0.00372031
R63138 DVSS.n20158 DVSS.n20047 0.00372031
R63139 DVSS.n13976 DVSS.n13955 0.00372031
R63140 DVSS.n21087 DVSS.n13956 0.00372031
R63141 DVSS.n21088 DVSS.n13957 0.00372031
R63142 DVSS.n21089 DVSS.n13958 0.00372031
R63143 DVSS.n21090 DVSS.n13959 0.00372031
R63144 DVSS.n21091 DVSS.n13960 0.00372031
R63145 DVSS.n21092 DVSS.n13961 0.00372031
R63146 DVSS.n21093 DVSS.n13962 0.00372031
R63147 DVSS.n21094 DVSS.n13963 0.00372031
R63148 DVSS.n21095 DVSS.n13964 0.00372031
R63149 DVSS.n21106 DVSS.n13940 0.00372031
R63150 DVSS.n13534 DVSS.n13517 0.00372031
R63151 DVSS.n13532 DVSS.n13526 0.00372031
R63152 DVSS.n13549 DVSS.n13518 0.00372031
R63153 DVSS.n13531 DVSS.n13525 0.00372031
R63154 DVSS.n13550 DVSS.n13519 0.00372031
R63155 DVSS.n13530 DVSS.n13524 0.00372031
R63156 DVSS.n13551 DVSS.n13520 0.00372031
R63157 DVSS.n13529 DVSS.n13523 0.00372031
R63158 DVSS.n13552 DVSS.n13521 0.00372031
R63159 DVSS.n13528 DVSS.n13522 0.00372031
R63160 DVSS.n608 DVSS.n598 0.00372031
R63161 DVSS.n613 DVSS.n597 0.00372031
R63162 DVSS.n614 DVSS.n599 0.00372031
R63163 DVSS.n611 DVSS.n604 0.00372031
R63164 DVSS.n610 DVSS.n603 0.00372031
R63165 DVSS.n615 DVSS.n601 0.00372031
R63166 DVSS.n609 DVSS.n602 0.00372031
R63167 DVSS.n21614 DVSS.n21602 0.00372031
R63168 DVSS.n21616 DVSS.n21558 0.00372031
R63169 DVSS.n21613 DVSS.n21601 0.00372031
R63170 DVSS.n21612 DVSS.n21600 0.00372031
R63171 DVSS.n21617 DVSS.n21560 0.00372031
R63172 DVSS.n21611 DVSS.n21599 0.00372031
R63173 DVSS.n21610 DVSS.n21598 0.00372031
R63174 DVSS.n21618 DVSS.n21562 0.00372031
R63175 DVSS.n21609 DVSS.n21597 0.00372031
R63176 DVSS.n21608 DVSS.n21596 0.00372031
R63177 DVSS.n21619 DVSS.n21564 0.00372031
R63178 DVSS.n21607 DVSS.n21595 0.00372031
R63179 DVSS.n21606 DVSS.n21594 0.00372031
R63180 DVSS.n21620 DVSS.n21566 0.00372031
R63181 DVSS.n21605 DVSS.n21593 0.00372031
R63182 DVSS.n21621 DVSS.n21592 0.00372031
R63183 DVSS.n21604 DVSS.n21590 0.00372031
R63184 DVSS.n256 DVSS.n207 0.00372031
R63185 DVSS.n238 DVSS.n227 0.00372031
R63186 DVSS.n237 DVSS.n226 0.00372031
R63187 DVSS.n257 DVSS.n209 0.00372031
R63188 DVSS.n236 DVSS.n225 0.00372031
R63189 DVSS.n235 DVSS.n224 0.00372031
R63190 DVSS.n258 DVSS.n211 0.00372031
R63191 DVSS.n234 DVSS.n223 0.00372031
R63192 DVSS.n233 DVSS.n222 0.00372031
R63193 DVSS.n259 DVSS.n213 0.00372031
R63194 DVSS.n232 DVSS.n221 0.00372031
R63195 DVSS.n261 DVSS.n220 0.00372031
R63196 DVSS.n230 DVSS.n215 0.00372031
R63197 DVSS.n255 DVSS.n206 0.00372031
R63198 DVSS.n260 DVSS.n216 0.00372031
R63199 DVSS.n231 DVSS.n218 0.00372031
R63200 DVSS.n23094 DVSS.n229 0.00372031
R63201 DVSS.n1161 DVSS.n1150 0.00372031
R63202 DVSS.n1149 DVSS.n1129 0.00372031
R63203 DVSS.n1157 DVSS.n1127 0.00372031
R63204 DVSS.n1158 DVSS.n1130 0.00372031
R63205 DVSS.n1147 DVSS.n1146 0.00372031
R63206 DVSS.n1162 DVSS.n1152 0.00372031
R63207 DVSS.n1160 DVSS.n1145 0.00372031
R63208 DVSS.n1144 DVSS.n1132 0.00372031
R63209 DVSS.n1156 DVSS.n1126 0.00372031
R63210 DVSS.n1159 DVSS.n1133 0.00372031
R63211 DVSS.n1142 DVSS.n1141 0.00372031
R63212 DVSS.n1163 DVSS.n1107 0.00372031
R63213 DVSS.n1140 DVSS.n1109 0.00372031
R63214 DVSS.n1139 DVSS.n1134 0.00372031
R63215 DVSS.n1155 DVSS.n1125 0.00372031
R63216 DVSS.n1137 DVSS.n1136 0.00372031
R63217 DVSS.n20048 DVSS.n20046 0.00372031
R63218 DVSS.n20047 DVSS.n20041 0.00372031
R63219 DVSS.n13528 DVSS.n13521 0.00372031
R63220 DVSS.n13552 DVSS.n13523 0.00372031
R63221 DVSS.n13529 DVSS.n13520 0.00372031
R63222 DVSS.n13551 DVSS.n13524 0.00372031
R63223 DVSS.n13530 DVSS.n13519 0.00372031
R63224 DVSS.n13550 DVSS.n13525 0.00372031
R63225 DVSS.n13531 DVSS.n13518 0.00372031
R63226 DVSS.n13549 DVSS.n13526 0.00372031
R63227 DVSS.n13532 DVSS.n13517 0.00372031
R63228 DVSS.n21298 DVSS.n13534 0.00372031
R63229 DVSS.n13966 DVSS.n13940 0.00372031
R63230 DVSS.n21095 DVSS.n13967 0.00372031
R63231 DVSS.n21094 DVSS.n13968 0.00372031
R63232 DVSS.n21093 DVSS.n13969 0.00372031
R63233 DVSS.n21092 DVSS.n13970 0.00372031
R63234 DVSS.n21091 DVSS.n13971 0.00372031
R63235 DVSS.n21090 DVSS.n13972 0.00372031
R63236 DVSS.n21089 DVSS.n13973 0.00372031
R63237 DVSS.n21088 DVSS.n13974 0.00372031
R63238 DVSS.n21087 DVSS.n13975 0.00372031
R63239 DVSS.n21104 DVSS.n13976 0.00372031
R63240 DVSS.n14471 DVSS.n14463 0.00372031
R63241 DVSS.n14472 DVSS.n14462 0.00372031
R63242 DVSS.n14473 DVSS.n14461 0.00372031
R63243 DVSS.n14474 DVSS.n14460 0.00372031
R63244 DVSS.n14893 DVSS.n14875 0.00372031
R63245 DVSS.n14904 DVSS.n14892 0.00372031
R63246 DVSS.n14905 DVSS.n14891 0.00372031
R63247 DVSS.n14906 DVSS.n14890 0.00372031
R63248 DVSS.n14907 DVSS.n14889 0.00372031
R63249 DVSS.n15307 DVSS.n15295 0.00372031
R63250 DVSS.n15308 DVSS.n15294 0.00372031
R63251 DVSS.n16092 DVSS.n16074 0.00372031
R63252 DVSS.n16098 DVSS.n16091 0.00372031
R63253 DVSS.n16097 DVSS.n16070 0.00372031
R63254 DVSS.n16100 DVSS.n16089 0.00372031
R63255 DVSS.n16254 DVSS.n16246 0.00372031
R63256 DVSS.n16253 DVSS.n16248 0.00372031
R63257 DVSS.n16252 DVSS.n16249 0.00372031
R63258 DVSS.n15799 DVSS.n15791 0.00372031
R63259 DVSS.n15798 DVSS.n15792 0.00372031
R63260 DVSS.n15797 DVSS.n15793 0.00372031
R63261 DVSS.n15796 DVSS.n15794 0.00372031
R63262 DVSS.n15755 DVSS.n15751 0.00372031
R63263 DVSS.n15750 DVSS.n15740 0.00372031
R63264 DVSS.n15754 DVSS.n15749 0.00372031
R63265 DVSS.n15748 DVSS.n15741 0.00372031
R63266 DVSS.n15753 DVSS.n15747 0.00372031
R63267 DVSS.n15746 DVSS.n15742 0.00372031
R63268 DVSS.n15752 DVSS.n15745 0.00372031
R63269 DVSS.n15744 DVSS.n15743 0.00372031
R63270 DVSS.n16182 DVSS.n16174 0.00372031
R63271 DVSS.n16177 DVSS.n16168 0.00372031
R63272 DVSS.n16181 DVSS.n16173 0.00372031
R63273 DVSS.n16178 DVSS.n16169 0.00372031
R63274 DVSS.n16183 DVSS.n16175 0.00372031
R63275 DVSS.n16180 DVSS.n16170 0.00372031
R63276 DVSS.n16825 DVSS.n16152 0.00372031
R63277 DVSS.n16828 DVSS.n16143 0.00372031
R63278 DVSS.n16836 DVSS.n16151 0.00372031
R63279 DVSS.n16829 DVSS.n16144 0.00372031
R63280 DVSS.n16833 DVSS.n16142 0.00372031
R63281 DVSS.n16834 DVSS.n16145 0.00372031
R63282 DVSS.n16831 DVSS.n16149 0.00372031
R63283 DVSS.n16835 DVSS.n16146 0.00372031
R63284 DVSS.n16830 DVSS.n16148 0.00372031
R63285 DVSS.n15379 DVSS.n15365 0.00372031
R63286 DVSS.n15376 DVSS.n15370 0.00372031
R63287 DVSS.n15380 DVSS.n15366 0.00372031
R63288 DVSS.n15375 DVSS.n15369 0.00372031
R63289 DVSS.n15378 DVSS.n15363 0.00372031
R63290 DVSS.n15374 DVSS.n14938 0.00372031
R63291 DVSS.n14945 DVSS.n14928 0.00372031
R63292 DVSS.n14943 DVSS.n14937 0.00372031
R63293 DVSS.n14988 DVSS.n14929 0.00372031
R63294 DVSS.n14942 DVSS.n14936 0.00372031
R63295 DVSS.n14989 DVSS.n14930 0.00372031
R63296 DVSS.n14941 DVSS.n14935 0.00372031
R63297 DVSS.n14990 DVSS.n14931 0.00372031
R63298 DVSS.n14940 DVSS.n14934 0.00372031
R63299 DVSS.n14991 DVSS.n14932 0.00372031
R63300 DVSS.n14939 DVSS.n14864 0.00372031
R63301 DVSS.n14426 DVSS.n14411 0.00372031
R63302 DVSS.n14424 DVSS.n14423 0.00372031
R63303 DVSS.n14441 DVSS.n14412 0.00372031
R63304 DVSS.n14422 DVSS.n14421 0.00372031
R63305 DVSS.n14442 DVSS.n14413 0.00372031
R63306 DVSS.n14420 DVSS.n14419 0.00372031
R63307 DVSS.n14443 DVSS.n14414 0.00372031
R63308 DVSS.n14418 DVSS.n14417 0.00372031
R63309 DVSS.n20303 DVSS.n20213 0.00372031
R63310 DVSS.n20304 DVSS.n14044 0.00372031
R63311 DVSS.n14067 DVSS.n14043 0.00372031
R63312 DVSS.n14045 DVSS.n14021 0.00372031
R63313 DVSS.n14066 DVSS.n14042 0.00372031
R63314 DVSS.n14046 DVSS.n14022 0.00372031
R63315 DVSS.n14065 DVSS.n14041 0.00372031
R63316 DVSS.n14047 DVSS.n14023 0.00372031
R63317 DVSS.n14064 DVSS.n14040 0.00372031
R63318 DVSS.n14048 DVSS.n14024 0.00372031
R63319 DVSS.n14063 DVSS.n14039 0.00372031
R63320 DVSS.n14049 DVSS.n14025 0.00372031
R63321 DVSS.n14062 DVSS.n14038 0.00372031
R63322 DVSS.n14050 DVSS.n14026 0.00372031
R63323 DVSS.n14061 DVSS.n14037 0.00372031
R63324 DVSS.n14051 DVSS.n14027 0.00372031
R63325 DVSS.n14060 DVSS.n14036 0.00372031
R63326 DVSS.n14052 DVSS.n14028 0.00372031
R63327 DVSS.n14059 DVSS.n14035 0.00372031
R63328 DVSS.n14053 DVSS.n14029 0.00372031
R63329 DVSS.n14058 DVSS.n14034 0.00372031
R63330 DVSS.n14054 DVSS.n14030 0.00372031
R63331 DVSS.n14057 DVSS.n14033 0.00372031
R63332 DVSS.n14055 DVSS.n14031 0.00372031
R63333 DVSS.n13482 DVSS.n13466 0.00372031
R63334 DVSS.n13480 DVSS.n13479 0.00372031
R63335 DVSS.n13497 DVSS.n13467 0.00372031
R63336 DVSS.n13478 DVSS.n13477 0.00372031
R63337 DVSS.n13498 DVSS.n13468 0.00372031
R63338 DVSS.n13476 DVSS.n13475 0.00372031
R63339 DVSS.n13499 DVSS.n13469 0.00372031
R63340 DVSS.n13474 DVSS.n13473 0.00372031
R63341 DVSS.n13500 DVSS.n13470 0.00372031
R63342 DVSS.n13472 DVSS.n13471 0.00372031
R63343 DVSS.n560 DVSS.n549 0.00372031
R63344 DVSS.n563 DVSS.n548 0.00372031
R63345 DVSS.n564 DVSS.n550 0.00372031
R63346 DVSS.n558 DVSS.n557 0.00372031
R63347 DVSS.n556 DVSS.n555 0.00372031
R63348 DVSS.n565 DVSS.n552 0.00372031
R63349 DVSS.n554 DVSS.n553 0.00372031
R63350 DVSS.n21717 DVSS.n21705 0.00372031
R63351 DVSS.n21719 DVSS.n21684 0.00372031
R63352 DVSS.n21716 DVSS.n21704 0.00372031
R63353 DVSS.n21715 DVSS.n21703 0.00372031
R63354 DVSS.n21720 DVSS.n21686 0.00372031
R63355 DVSS.n21714 DVSS.n21702 0.00372031
R63356 DVSS.n21713 DVSS.n21701 0.00372031
R63357 DVSS.n21721 DVSS.n21688 0.00372031
R63358 DVSS.n21712 DVSS.n21700 0.00372031
R63359 DVSS.n21711 DVSS.n21699 0.00372031
R63360 DVSS.n21722 DVSS.n21690 0.00372031
R63361 DVSS.n21710 DVSS.n21698 0.00372031
R63362 DVSS.n21709 DVSS.n21697 0.00372031
R63363 DVSS.n21723 DVSS.n21692 0.00372031
R63364 DVSS.n21708 DVSS.n21696 0.00372031
R63365 DVSS.n21724 DVSS.n21695 0.00372031
R63366 DVSS.n21707 DVSS.n1178 0.00372031
R63367 DVSS.n176 DVSS.n127 0.00372031
R63368 DVSS.n158 DVSS.n147 0.00372031
R63369 DVSS.n157 DVSS.n146 0.00372031
R63370 DVSS.n177 DVSS.n129 0.00372031
R63371 DVSS.n156 DVSS.n145 0.00372031
R63372 DVSS.n155 DVSS.n144 0.00372031
R63373 DVSS.n178 DVSS.n131 0.00372031
R63374 DVSS.n154 DVSS.n143 0.00372031
R63375 DVSS.n153 DVSS.n142 0.00372031
R63376 DVSS.n179 DVSS.n133 0.00372031
R63377 DVSS.n152 DVSS.n141 0.00372031
R63378 DVSS.n181 DVSS.n140 0.00372031
R63379 DVSS.n150 DVSS.n135 0.00372031
R63380 DVSS.n175 DVSS.n126 0.00372031
R63381 DVSS.n180 DVSS.n136 0.00372031
R63382 DVSS.n151 DVSS.n138 0.00372031
R63383 DVSS.n23137 DVSS.n149 0.00372031
R63384 DVSS.n13039 DVSS.n13037 0.00372031
R63385 DVSS.n13038 DVSS.n12995 0.00372031
R63386 DVSS.n12994 DVSS.n12992 0.00372031
R63387 DVSS.n13035 DVSS.n12996 0.00372031
R63388 DVSS.n13027 DVSS.n13026 0.00372031
R63389 DVSS.n13056 DVSS.n13048 0.00372031
R63390 DVSS.n13025 DVSS.n13023 0.00372031
R63391 DVSS.n13024 DVSS.n12999 0.00372031
R63392 DVSS.n12998 DVSS.n12991 0.00372031
R63393 DVSS.n13021 DVSS.n13000 0.00372031
R63394 DVSS.n13013 DVSS.n13012 0.00372031
R63395 DVSS.n13061 DVSS.n13057 0.00372031
R63396 DVSS.n13011 DVSS.n13009 0.00372031
R63397 DVSS.n13010 DVSS.n13003 0.00372031
R63398 DVSS.n13002 DVSS.n12962 0.00372031
R63399 DVSS.n13007 DVSS.n13006 0.00372031
R63400 DVSS.n20213 DVSS.n20212 0.00372031
R63401 DVSS.n20304 DVSS.n20303 0.00372031
R63402 DVSS.n13471 DVSS.n13470 0.00372031
R63403 DVSS.n13500 DVSS.n13474 0.00372031
R63404 DVSS.n13473 DVSS.n13469 0.00372031
R63405 DVSS.n13499 DVSS.n13476 0.00372031
R63406 DVSS.n13475 DVSS.n13468 0.00372031
R63407 DVSS.n13498 DVSS.n13478 0.00372031
R63408 DVSS.n13477 DVSS.n13467 0.00372031
R63409 DVSS.n13497 DVSS.n13480 0.00372031
R63410 DVSS.n13479 DVSS.n13466 0.00372031
R63411 DVSS.n21339 DVSS.n13482 0.00372031
R63412 DVSS.n14055 DVSS.n14033 0.00372031
R63413 DVSS.n14057 DVSS.n14030 0.00372031
R63414 DVSS.n14054 DVSS.n14034 0.00372031
R63415 DVSS.n14058 DVSS.n14029 0.00372031
R63416 DVSS.n14053 DVSS.n14035 0.00372031
R63417 DVSS.n14059 DVSS.n14028 0.00372031
R63418 DVSS.n14052 DVSS.n14036 0.00372031
R63419 DVSS.n14060 DVSS.n14027 0.00372031
R63420 DVSS.n14051 DVSS.n14037 0.00372031
R63421 DVSS.n14061 DVSS.n14026 0.00372031
R63422 DVSS.n14050 DVSS.n14038 0.00372031
R63423 DVSS.n14062 DVSS.n14025 0.00372031
R63424 DVSS.n14049 DVSS.n14039 0.00372031
R63425 DVSS.n14063 DVSS.n14024 0.00372031
R63426 DVSS.n14048 DVSS.n14040 0.00372031
R63427 DVSS.n14064 DVSS.n14023 0.00372031
R63428 DVSS.n14047 DVSS.n14041 0.00372031
R63429 DVSS.n14065 DVSS.n14022 0.00372031
R63430 DVSS.n14046 DVSS.n14042 0.00372031
R63431 DVSS.n14066 DVSS.n14021 0.00372031
R63432 DVSS.n14045 DVSS.n14043 0.00372031
R63433 DVSS.n14067 DVSS.n14020 0.00372031
R63434 DVSS.n14417 DVSS.n14414 0.00372031
R63435 DVSS.n14443 DVSS.n14420 0.00372031
R63436 DVSS.n14419 DVSS.n14413 0.00372031
R63437 DVSS.n14442 DVSS.n14422 0.00372031
R63438 DVSS.n14421 DVSS.n14412 0.00372031
R63439 DVSS.n14441 DVSS.n14424 0.00372031
R63440 DVSS.n14423 DVSS.n14411 0.00372031
R63441 DVSS.n20889 DVSS.n14426 0.00372031
R63442 DVSS.n14939 DVSS.n14932 0.00372031
R63443 DVSS.n14991 DVSS.n14934 0.00372031
R63444 DVSS.n14940 DVSS.n14931 0.00372031
R63445 DVSS.n14990 DVSS.n14935 0.00372031
R63446 DVSS.n14941 DVSS.n14930 0.00372031
R63447 DVSS.n14989 DVSS.n14936 0.00372031
R63448 DVSS.n14942 DVSS.n14929 0.00372031
R63449 DVSS.n14988 DVSS.n14937 0.00372031
R63450 DVSS.n14943 DVSS.n14928 0.00372031
R63451 DVSS.n19982 DVSS.n14945 0.00372031
R63452 DVSS.n15374 DVSS.n15367 0.00372031
R63453 DVSS.n15378 DVSS.n15369 0.00372031
R63454 DVSS.n15375 DVSS.n15366 0.00372031
R63455 DVSS.n15380 DVSS.n15370 0.00372031
R63456 DVSS.n15376 DVSS.n15365 0.00372031
R63457 DVSS.n15379 DVSS.n15371 0.00372031
R63458 DVSS.n16830 DVSS.n16146 0.00372031
R63459 DVSS.n16835 DVSS.n16149 0.00372031
R63460 DVSS.n16831 DVSS.n16145 0.00372031
R63461 DVSS.n16834 DVSS.n16150 0.00372031
R63462 DVSS.n16833 DVSS.n16144 0.00372031
R63463 DVSS.n16829 DVSS.n16151 0.00372031
R63464 DVSS.n16836 DVSS.n16143 0.00372031
R63465 DVSS.n16828 DVSS.n16826 0.00372031
R63466 DVSS.n16170 DVSS.n16152 0.00372031
R63467 DVSS.n16180 DVSS.n16172 0.00372031
R63468 DVSS.n16183 DVSS.n16169 0.00372031
R63469 DVSS.n16178 DVSS.n16173 0.00372031
R63470 DVSS.n16181 DVSS.n16168 0.00372031
R63471 DVSS.n16177 DVSS.n16174 0.00372031
R63472 DVSS.n16182 DVSS.n16167 0.00372031
R63473 DVSS.n15745 DVSS.n15744 0.00372031
R63474 DVSS.n15752 DVSS.n15742 0.00372031
R63475 DVSS.n15747 DVSS.n15746 0.00372031
R63476 DVSS.n15753 DVSS.n15741 0.00372031
R63477 DVSS.n15749 DVSS.n15748 0.00372031
R63478 DVSS.n15754 DVSS.n15740 0.00372031
R63479 DVSS.n15751 DVSS.n15750 0.00372031
R63480 DVSS.n15755 DVSS.n15739 0.00372031
R63481 DVSS.n15847 DVSS.n15846 0.00372031
R63482 DVSS.n15849 DVSS.n15838 0.00372031
R63483 DVSS.n15845 DVSS.n15844 0.00372031
R63484 DVSS.n16305 DVSS.n16297 0.00372031
R63485 DVSS.n16299 DVSS.n16298 0.00372031
R63486 DVSS.n16006 DVSS.n15995 0.00372031
R63487 DVSS.n16014 DVSS.n16003 0.00372031
R63488 DVSS.n16007 DVSS.n15996 0.00372031
R63489 DVSS.n16011 DVSS.n15994 0.00372031
R63490 DVSS.n16012 DVSS.n15997 0.00372031
R63491 DVSS.n16009 DVSS.n16001 0.00372031
R63492 DVSS.n16013 DVSS.n15998 0.00372031
R63493 DVSS.n16008 DVSS.n16000 0.00372031
R63494 DVSS.n15264 DVSS.n15256 0.00372031
R63495 DVSS.n15270 DVSS.n15263 0.00372031
R63496 DVSS.n15262 DVSS.n15257 0.00372031
R63497 DVSS.n15269 DVSS.n15261 0.00372031
R63498 DVSS.n15260 DVSS.n15254 0.00372031
R63499 DVSS.n18381 DVSS.n15239 0.00372031
R63500 DVSS.n18382 DVSS.n15229 0.00372031
R63501 DVSS.n18398 DVSS.n15238 0.00372031
R63502 DVSS.n18428 DVSS.n15230 0.00372031
R63503 DVSS.n18397 DVSS.n15237 0.00372031
R63504 DVSS.n18429 DVSS.n15231 0.00372031
R63505 DVSS.n18396 DVSS.n15236 0.00372031
R63506 DVSS.n18430 DVSS.n15232 0.00372031
R63507 DVSS.n18395 DVSS.n15235 0.00372031
R63508 DVSS.n18431 DVSS.n15233 0.00372031
R63509 DVSS.n18394 DVSS.n14536 0.00372031
R63510 DVSS.n20705 DVSS.n14507 0.00372031
R63511 DVSS.n20703 DVSS.n14516 0.00372031
R63512 DVSS.n20719 DVSS.n14508 0.00372031
R63513 DVSS.n20702 DVSS.n14515 0.00372031
R63514 DVSS.n20720 DVSS.n14509 0.00372031
R63515 DVSS.n20701 DVSS.n14514 0.00372031
R63516 DVSS.n20721 DVSS.n14510 0.00372031
R63517 DVSS.n20700 DVSS.n14513 0.00372031
R63518 DVSS.n18874 DVSS.n18870 0.00372031
R63519 DVSS.n18875 DVSS.n13849 0.00372031
R63520 DVSS.n13872 DVSS.n13848 0.00372031
R63521 DVSS.n13850 DVSS.n13826 0.00372031
R63522 DVSS.n13871 DVSS.n13847 0.00372031
R63523 DVSS.n13851 DVSS.n13827 0.00372031
R63524 DVSS.n13870 DVSS.n13846 0.00372031
R63525 DVSS.n13852 DVSS.n13828 0.00372031
R63526 DVSS.n13869 DVSS.n13845 0.00372031
R63527 DVSS.n13853 DVSS.n13829 0.00372031
R63528 DVSS.n13868 DVSS.n13844 0.00372031
R63529 DVSS.n13854 DVSS.n13830 0.00372031
R63530 DVSS.n13867 DVSS.n13843 0.00372031
R63531 DVSS.n13855 DVSS.n13831 0.00372031
R63532 DVSS.n13866 DVSS.n13842 0.00372031
R63533 DVSS.n13856 DVSS.n13832 0.00372031
R63534 DVSS.n13865 DVSS.n13841 0.00372031
R63535 DVSS.n13857 DVSS.n13833 0.00372031
R63536 DVSS.n13864 DVSS.n13840 0.00372031
R63537 DVSS.n13858 DVSS.n13834 0.00372031
R63538 DVSS.n13863 DVSS.n13839 0.00372031
R63539 DVSS.n13859 DVSS.n13835 0.00372031
R63540 DVSS.n13862 DVSS.n13838 0.00372031
R63541 DVSS.n13860 DVSS.n13836 0.00372031
R63542 DVSS.n13582 DVSS.n13571 0.00372031
R63543 DVSS.n13583 DVSS.n13580 0.00372031
R63544 DVSS.n667 DVSS.n650 0.00372031
R63545 DVSS.n670 DVSS.n649 0.00372031
R63546 DVSS.n671 DVSS.n651 0.00372031
R63547 DVSS.n665 DVSS.n658 0.00372031
R63548 DVSS.n657 DVSS.n656 0.00372031
R63549 DVSS.n672 DVSS.n653 0.00372031
R63550 DVSS.n655 DVSS.n654 0.00372031
R63551 DVSS.n21943 DVSS.n21851 0.00372031
R63552 DVSS.n21942 DVSS.n21871 0.00372031
R63553 DVSS.n21941 DVSS.n21933 0.00372031
R63554 DVSS.n21931 DVSS.n21921 0.00372031
R63555 DVSS.n21920 DVSS.n21873 0.00372031
R63556 DVSS.n21930 DVSS.n21919 0.00372031
R63557 DVSS.n21929 DVSS.n21911 0.00372031
R63558 DVSS.n21910 DVSS.n21875 0.00372031
R63559 DVSS.n21928 DVSS.n21909 0.00372031
R63560 DVSS.n21927 DVSS.n21901 0.00372031
R63561 DVSS.n21900 DVSS.n21877 0.00372031
R63562 DVSS.n21926 DVSS.n21899 0.00372031
R63563 DVSS.n21925 DVSS.n21891 0.00372031
R63564 DVSS.n21890 DVSS.n21879 0.00372031
R63565 DVSS.n21924 DVSS.n21889 0.00372031
R63566 DVSS.n21882 DVSS.n21881 0.00372031
R63567 DVSS.n21923 DVSS.n870 0.00372031
R63568 DVSS.n22492 DVSS.n803 0.00372031
R63569 DVSS.n22471 DVSS.n857 0.00372031
R63570 DVSS.n22470 DVSS.n850 0.00372031
R63571 DVSS.n22493 DVSS.n805 0.00372031
R63572 DVSS.n22469 DVSS.n849 0.00372031
R63573 DVSS.n22468 DVSS.n841 0.00372031
R63574 DVSS.n22494 DVSS.n807 0.00372031
R63575 DVSS.n22467 DVSS.n840 0.00372031
R63576 DVSS.n22466 DVSS.n832 0.00372031
R63577 DVSS.n22495 DVSS.n809 0.00372031
R63578 DVSS.n22465 DVSS.n831 0.00372031
R63579 DVSS.n22497 DVSS.n823 0.00372031
R63580 DVSS.n22463 DVSS.n811 0.00372031
R63581 DVSS.n22491 DVSS.n802 0.00372031
R63582 DVSS.n22496 DVSS.n812 0.00372031
R63583 DVSS.n22464 DVSS.n814 0.00372031
R63584 DVSS.n22503 DVSS.n22462 0.00372031
R63585 DVSS.n1095 DVSS.n1094 0.00372031
R63586 DVSS.n1101 DVSS.n1072 0.00372031
R63587 DVSS.n1071 DVSS.n1069 0.00372031
R63588 DVSS.n1092 DVSS.n1073 0.00372031
R63589 DVSS.n1105 DVSS.n1091 0.00372031
R63590 DVSS.n1098 DVSS.n1097 0.00372031
R63591 DVSS.n1090 DVSS.n1089 0.00372031
R63592 DVSS.n1102 DVSS.n1076 0.00372031
R63593 DVSS.n1075 DVSS.n1068 0.00372031
R63594 DVSS.n1087 DVSS.n1077 0.00372031
R63595 DVSS.n1104 DVSS.n1086 0.00372031
R63596 DVSS.n22378 DVSS.n1099 0.00372031
R63597 DVSS.n1085 DVSS.n1084 0.00372031
R63598 DVSS.n1103 DVSS.n1080 0.00372031
R63599 DVSS.n1079 DVSS.n1017 0.00372031
R63600 DVSS.n1082 DVSS.n1052 0.00372031
R63601 DVSS.n18984 DVSS.n18874 0.00372031
R63602 DVSS.n18875 DVSS.n18870 0.00372031
R63603 DVSS.n13583 DVSS.n13571 0.00372031
R63604 DVSS.n21256 DVSS.n13582 0.00372031
R63605 DVSS.n13860 DVSS.n13838 0.00372031
R63606 DVSS.n13862 DVSS.n13835 0.00372031
R63607 DVSS.n13859 DVSS.n13839 0.00372031
R63608 DVSS.n13863 DVSS.n13834 0.00372031
R63609 DVSS.n13858 DVSS.n13840 0.00372031
R63610 DVSS.n13864 DVSS.n13833 0.00372031
R63611 DVSS.n13857 DVSS.n13841 0.00372031
R63612 DVSS.n13865 DVSS.n13832 0.00372031
R63613 DVSS.n13856 DVSS.n13842 0.00372031
R63614 DVSS.n13866 DVSS.n13831 0.00372031
R63615 DVSS.n13855 DVSS.n13843 0.00372031
R63616 DVSS.n13867 DVSS.n13830 0.00372031
R63617 DVSS.n13854 DVSS.n13844 0.00372031
R63618 DVSS.n13868 DVSS.n13829 0.00372031
R63619 DVSS.n13853 DVSS.n13845 0.00372031
R63620 DVSS.n13869 DVSS.n13828 0.00372031
R63621 DVSS.n13852 DVSS.n13846 0.00372031
R63622 DVSS.n13870 DVSS.n13827 0.00372031
R63623 DVSS.n13851 DVSS.n13847 0.00372031
R63624 DVSS.n13871 DVSS.n13826 0.00372031
R63625 DVSS.n13850 DVSS.n13848 0.00372031
R63626 DVSS.n13872 DVSS.n13825 0.00372031
R63627 DVSS.n20700 DVSS.n14510 0.00372031
R63628 DVSS.n20721 DVSS.n14514 0.00372031
R63629 DVSS.n20701 DVSS.n14509 0.00372031
R63630 DVSS.n20720 DVSS.n14515 0.00372031
R63631 DVSS.n20702 DVSS.n14508 0.00372031
R63632 DVSS.n20719 DVSS.n14516 0.00372031
R63633 DVSS.n20703 DVSS.n14507 0.00372031
R63634 DVSS.n20804 DVSS.n20705 0.00372031
R63635 DVSS.n18394 DVSS.n15233 0.00372031
R63636 DVSS.n18431 DVSS.n15235 0.00372031
R63637 DVSS.n18395 DVSS.n15232 0.00372031
R63638 DVSS.n18430 DVSS.n15236 0.00372031
R63639 DVSS.n18396 DVSS.n15231 0.00372031
R63640 DVSS.n18429 DVSS.n15237 0.00372031
R63641 DVSS.n18397 DVSS.n15230 0.00372031
R63642 DVSS.n18428 DVSS.n15238 0.00372031
R63643 DVSS.n18398 DVSS.n15229 0.00372031
R63644 DVSS.n18473 DVSS.n18382 0.00372031
R63645 DVSS.n15258 DVSS.n15239 0.00372031
R63646 DVSS.n15261 DVSS.n15260 0.00372031
R63647 DVSS.n15269 DVSS.n15257 0.00372031
R63648 DVSS.n15263 DVSS.n15262 0.00372031
R63649 DVSS.n15270 DVSS.n15256 0.00372031
R63650 DVSS.n15265 DVSS.n15264 0.00372031
R63651 DVSS.n16008 DVSS.n15998 0.00372031
R63652 DVSS.n16013 DVSS.n16001 0.00372031
R63653 DVSS.n16009 DVSS.n15997 0.00372031
R63654 DVSS.n16012 DVSS.n16002 0.00372031
R63655 DVSS.n16011 DVSS.n15996 0.00372031
R63656 DVSS.n16007 DVSS.n16003 0.00372031
R63657 DVSS.n16014 DVSS.n15995 0.00372031
R63658 DVSS.n16006 DVSS.n16004 0.00372031
R63659 DVSS.n16298 DVSS.n16297 0.00372031
R63660 DVSS.n16305 DVSS.n16300 0.00372031
R63661 DVSS.n15844 DVSS.n15838 0.00372031
R63662 DVSS.n15849 DVSS.n15847 0.00372031
R63663 DVSS.n15846 DVSS.n15837 0.00372031
R63664 DVSS.n15722 DVSS.n15720 0.00372031
R63665 DVSS.n15721 DVSS.n15705 0.00372031
R63666 DVSS.n15719 DVSS.n15711 0.00372031
R63667 DVSS.n15672 DVSS.n15671 0.00372031
R63668 DVSS.n15677 DVSS.n15674 0.00372031
R63669 DVSS.n17531 DVSS.n16890 0.00372031
R63670 DVSS.n17539 DVSS.n16898 0.00372031
R63671 DVSS.n17532 DVSS.n16891 0.00372031
R63672 DVSS.n17536 DVSS.n16889 0.00372031
R63673 DVSS.n17537 DVSS.n16892 0.00372031
R63674 DVSS.n17534 DVSS.n16896 0.00372031
R63675 DVSS.n17538 DVSS.n16893 0.00372031
R63676 DVSS.n17533 DVSS.n16895 0.00372031
R63677 DVSS.n15458 DVSS.n15435 0.00372031
R63678 DVSS.n15455 DVSS.n15440 0.00372031
R63679 DVSS.n15459 DVSS.n15436 0.00372031
R63680 DVSS.n15454 DVSS.n15439 0.00372031
R63681 DVSS.n15457 DVSS.n15433 0.00372031
R63682 DVSS.n15453 DVSS.n15011 0.00372031
R63683 DVSS.n15018 DVSS.n15001 0.00372031
R63684 DVSS.n15016 DVSS.n15010 0.00372031
R63685 DVSS.n15067 DVSS.n15002 0.00372031
R63686 DVSS.n15015 DVSS.n15009 0.00372031
R63687 DVSS.n15068 DVSS.n15003 0.00372031
R63688 DVSS.n15014 DVSS.n15008 0.00372031
R63689 DVSS.n15069 DVSS.n15004 0.00372031
R63690 DVSS.n15013 DVSS.n15007 0.00372031
R63691 DVSS.n15070 DVSS.n15005 0.00372031
R63692 DVSS.n15012 DVSS.n14853 0.00372031
R63693 DVSS.n14377 DVSS.n14362 0.00372031
R63694 DVSS.n14375 DVSS.n14374 0.00372031
R63695 DVSS.n14392 DVSS.n14363 0.00372031
R63696 DVSS.n14373 DVSS.n14372 0.00372031
R63697 DVSS.n14393 DVSS.n14364 0.00372031
R63698 DVSS.n14371 DVSS.n14370 0.00372031
R63699 DVSS.n14394 DVSS.n14365 0.00372031
R63700 DVSS.n14369 DVSS.n14368 0.00372031
R63701 DVSS.n14678 DVSS.n14674 0.00372031
R63702 DVSS.n14679 DVSS.n14150 0.00372031
R63703 DVSS.n14173 DVSS.n14149 0.00372031
R63704 DVSS.n14151 DVSS.n14127 0.00372031
R63705 DVSS.n14172 DVSS.n14148 0.00372031
R63706 DVSS.n14152 DVSS.n14128 0.00372031
R63707 DVSS.n14171 DVSS.n14147 0.00372031
R63708 DVSS.n14153 DVSS.n14129 0.00372031
R63709 DVSS.n14170 DVSS.n14146 0.00372031
R63710 DVSS.n14154 DVSS.n14130 0.00372031
R63711 DVSS.n14169 DVSS.n14145 0.00372031
R63712 DVSS.n14155 DVSS.n14131 0.00372031
R63713 DVSS.n14168 DVSS.n14144 0.00372031
R63714 DVSS.n14156 DVSS.n14132 0.00372031
R63715 DVSS.n14167 DVSS.n14143 0.00372031
R63716 DVSS.n14157 DVSS.n14133 0.00372031
R63717 DVSS.n14166 DVSS.n14142 0.00372031
R63718 DVSS.n14158 DVSS.n14134 0.00372031
R63719 DVSS.n14165 DVSS.n14141 0.00372031
R63720 DVSS.n14159 DVSS.n14135 0.00372031
R63721 DVSS.n14164 DVSS.n14140 0.00372031
R63722 DVSS.n14160 DVSS.n14136 0.00372031
R63723 DVSS.n14163 DVSS.n14139 0.00372031
R63724 DVSS.n14161 DVSS.n14137 0.00372031
R63725 DVSS.n13431 DVSS.n13420 0.00372031
R63726 DVSS.n13435 DVSS.n13429 0.00372031
R63727 DVSS.n508 DVSS.n498 0.00372031
R63728 DVSS.n513 DVSS.n497 0.00372031
R63729 DVSS.n514 DVSS.n499 0.00372031
R63730 DVSS.n511 DVSS.n504 0.00372031
R63731 DVSS.n510 DVSS.n503 0.00372031
R63732 DVSS.n515 DVSS.n501 0.00372031
R63733 DVSS.n509 DVSS.n502 0.00372031
R63734 DVSS.n21810 DVSS.n21798 0.00372031
R63735 DVSS.n21812 DVSS.n21778 0.00372031
R63736 DVSS.n21809 DVSS.n21797 0.00372031
R63737 DVSS.n21808 DVSS.n21796 0.00372031
R63738 DVSS.n21813 DVSS.n21780 0.00372031
R63739 DVSS.n21807 DVSS.n21795 0.00372031
R63740 DVSS.n21806 DVSS.n21794 0.00372031
R63741 DVSS.n21814 DVSS.n21782 0.00372031
R63742 DVSS.n21805 DVSS.n21793 0.00372031
R63743 DVSS.n21804 DVSS.n21792 0.00372031
R63744 DVSS.n21815 DVSS.n21784 0.00372031
R63745 DVSS.n21803 DVSS.n21791 0.00372031
R63746 DVSS.n21802 DVSS.n21790 0.00372031
R63747 DVSS.n21816 DVSS.n21786 0.00372031
R63748 DVSS.n21801 DVSS.n21789 0.00372031
R63749 DVSS.n21817 DVSS.n21788 0.00372031
R63750 DVSS.n21800 DVSS.n1199 0.00372031
R63751 DVSS.n23166 DVSS.n62 0.00372031
R63752 DVSS.n93 DVSS.n82 0.00372031
R63753 DVSS.n92 DVSS.n81 0.00372031
R63754 DVSS.n23167 DVSS.n64 0.00372031
R63755 DVSS.n91 DVSS.n80 0.00372031
R63756 DVSS.n90 DVSS.n79 0.00372031
R63757 DVSS.n23168 DVSS.n66 0.00372031
R63758 DVSS.n89 DVSS.n78 0.00372031
R63759 DVSS.n88 DVSS.n77 0.00372031
R63760 DVSS.n23169 DVSS.n68 0.00372031
R63761 DVSS.n87 DVSS.n76 0.00372031
R63762 DVSS.n23171 DVSS.n75 0.00372031
R63763 DVSS.n85 DVSS.n70 0.00372031
R63764 DVSS.n23165 DVSS.n61 0.00372031
R63765 DVSS.n23170 DVSS.n71 0.00372031
R63766 DVSS.n86 DVSS.n73 0.00372031
R63767 DVSS.n23181 DVSS.n84 0.00372031
R63768 DVSS.n363 DVSS.n362 0.00372031
R63769 DVSS.n370 DVSS.n340 0.00372031
R63770 DVSS.n339 DVSS.n337 0.00372031
R63771 DVSS.n360 DVSS.n341 0.00372031
R63772 DVSS.n375 DVSS.n359 0.00372031
R63773 DVSS.n366 DVSS.n365 0.00372031
R63774 DVSS.n358 DVSS.n357 0.00372031
R63775 DVSS.n371 DVSS.n344 0.00372031
R63776 DVSS.n343 DVSS.n336 0.00372031
R63777 DVSS.n355 DVSS.n345 0.00372031
R63778 DVSS.n374 DVSS.n354 0.00372031
R63779 DVSS.n368 DVSS.n367 0.00372031
R63780 DVSS.n353 DVSS.n352 0.00372031
R63781 DVSS.n372 DVSS.n348 0.00372031
R63782 DVSS.n347 DVSS.n335 0.00372031
R63783 DVSS.n373 DVSS.n349 0.00372031
R63784 DVSS.n20626 DVSS.n14678 0.00372031
R63785 DVSS.n14679 DVSS.n14674 0.00372031
R63786 DVSS.n13435 DVSS.n13420 0.00372031
R63787 DVSS.n21383 DVSS.n13431 0.00372031
R63788 DVSS.n14161 DVSS.n14139 0.00372031
R63789 DVSS.n14163 DVSS.n14136 0.00372031
R63790 DVSS.n14160 DVSS.n14140 0.00372031
R63791 DVSS.n14164 DVSS.n14135 0.00372031
R63792 DVSS.n14159 DVSS.n14141 0.00372031
R63793 DVSS.n14165 DVSS.n14134 0.00372031
R63794 DVSS.n14158 DVSS.n14142 0.00372031
R63795 DVSS.n14166 DVSS.n14133 0.00372031
R63796 DVSS.n14157 DVSS.n14143 0.00372031
R63797 DVSS.n14167 DVSS.n14132 0.00372031
R63798 DVSS.n14156 DVSS.n14144 0.00372031
R63799 DVSS.n14168 DVSS.n14131 0.00372031
R63800 DVSS.n14155 DVSS.n14145 0.00372031
R63801 DVSS.n14169 DVSS.n14130 0.00372031
R63802 DVSS.n14154 DVSS.n14146 0.00372031
R63803 DVSS.n14170 DVSS.n14129 0.00372031
R63804 DVSS.n14153 DVSS.n14147 0.00372031
R63805 DVSS.n14171 DVSS.n14128 0.00372031
R63806 DVSS.n14152 DVSS.n14148 0.00372031
R63807 DVSS.n14172 DVSS.n14127 0.00372031
R63808 DVSS.n14151 DVSS.n14149 0.00372031
R63809 DVSS.n14173 DVSS.n14126 0.00372031
R63810 DVSS.n14368 DVSS.n14365 0.00372031
R63811 DVSS.n14394 DVSS.n14371 0.00372031
R63812 DVSS.n14370 DVSS.n14364 0.00372031
R63813 DVSS.n14393 DVSS.n14373 0.00372031
R63814 DVSS.n14372 DVSS.n14363 0.00372031
R63815 DVSS.n14392 DVSS.n14375 0.00372031
R63816 DVSS.n14374 DVSS.n14362 0.00372031
R63817 DVSS.n20929 DVSS.n14377 0.00372031
R63818 DVSS.n15012 DVSS.n15005 0.00372031
R63819 DVSS.n15070 DVSS.n15007 0.00372031
R63820 DVSS.n15013 DVSS.n15004 0.00372031
R63821 DVSS.n15069 DVSS.n15008 0.00372031
R63822 DVSS.n15014 DVSS.n15003 0.00372031
R63823 DVSS.n15068 DVSS.n15009 0.00372031
R63824 DVSS.n15015 DVSS.n15002 0.00372031
R63825 DVSS.n15067 DVSS.n15010 0.00372031
R63826 DVSS.n15016 DVSS.n15001 0.00372031
R63827 DVSS.n19971 DVSS.n15018 0.00372031
R63828 DVSS.n15453 DVSS.n15437 0.00372031
R63829 DVSS.n15457 DVSS.n15439 0.00372031
R63830 DVSS.n15454 DVSS.n15436 0.00372031
R63831 DVSS.n15459 DVSS.n15440 0.00372031
R63832 DVSS.n15455 DVSS.n15435 0.00372031
R63833 DVSS.n15458 DVSS.n15441 0.00372031
R63834 DVSS.n17533 DVSS.n16893 0.00372031
R63835 DVSS.n17538 DVSS.n16896 0.00372031
R63836 DVSS.n17534 DVSS.n16892 0.00372031
R63837 DVSS.n17537 DVSS.n16897 0.00372031
R63838 DVSS.n17536 DVSS.n16891 0.00372031
R63839 DVSS.n17532 DVSS.n16898 0.00372031
R63840 DVSS.n17539 DVSS.n16890 0.00372031
R63841 DVSS.n17531 DVSS.n16899 0.00372031
R63842 DVSS.n15674 DVSS.n15672 0.00372031
R63843 DVSS.n15671 DVSS.n15635 0.00372031
R63844 DVSS.n15711 DVSS.n15705 0.00372031
R63845 DVSS.n15722 DVSS.n15721 0.00372031
R63846 DVSS.n15720 DVSS.n15704 0.00372031
R63847 DVSS.n654 DVSS.n653 0.00372031
R63848 DVSS.n672 DVSS.n657 0.00372031
R63849 DVSS.n656 DVSS.n652 0.00372031
R63850 DVSS.n658 DVSS.n651 0.00372031
R63851 DVSS.n671 DVSS.n666 0.00372031
R63852 DVSS.n670 DVSS.n650 0.00372031
R63853 DVSS.n668 DVSS.n667 0.00372031
R63854 DVSS.n609 DVSS.n601 0.00372031
R63855 DVSS.n615 DVSS.n603 0.00372031
R63856 DVSS.n610 DVSS.n600 0.00372031
R63857 DVSS.n611 DVSS.n599 0.00372031
R63858 DVSS.n614 DVSS.n605 0.00372031
R63859 DVSS.n613 DVSS.n598 0.00372031
R63860 DVSS.n608 DVSS.n606 0.00372031
R63861 DVSS.n553 DVSS.n552 0.00372031
R63862 DVSS.n565 DVSS.n556 0.00372031
R63863 DVSS.n555 DVSS.n551 0.00372031
R63864 DVSS.n557 DVSS.n550 0.00372031
R63865 DVSS.n564 DVSS.n559 0.00372031
R63866 DVSS.n563 DVSS.n549 0.00372031
R63867 DVSS.n561 DVSS.n560 0.00372031
R63868 DVSS.n509 DVSS.n501 0.00372031
R63869 DVSS.n515 DVSS.n503 0.00372031
R63870 DVSS.n510 DVSS.n500 0.00372031
R63871 DVSS.n511 DVSS.n499 0.00372031
R63872 DVSS.n514 DVSS.n505 0.00372031
R63873 DVSS.n513 DVSS.n498 0.00372031
R63874 DVSS.n508 DVSS.n506 0.00372031
R63875 DVSS.n22380 DVSS.n1052 0.00372031
R63876 DVSS.n1080 DVSS.n1079 0.00372031
R63877 DVSS.n1103 DVSS.n1085 0.00372031
R63878 DVSS.n1084 DVSS.n1078 0.00372031
R63879 DVSS.n1099 DVSS.n1086 0.00372031
R63880 DVSS.n1104 DVSS.n1077 0.00372031
R63881 DVSS.n1088 DVSS.n1087 0.00372031
R63882 DVSS.n1076 DVSS.n1075 0.00372031
R63883 DVSS.n1102 DVSS.n1090 0.00372031
R63884 DVSS.n1089 DVSS.n1074 0.00372031
R63885 DVSS.n1097 DVSS.n1091 0.00372031
R63886 DVSS.n1105 DVSS.n1073 0.00372031
R63887 DVSS.n1093 DVSS.n1092 0.00372031
R63888 DVSS.n1072 DVSS.n1071 0.00372031
R63889 DVSS.n1101 DVSS.n1095 0.00372031
R63890 DVSS.n1094 DVSS.n1070 0.00372031
R63891 DVSS.n1138 DVSS.n1137 0.00372031
R63892 DVSS.n1155 DVSS.n1134 0.00372031
R63893 DVSS.n1140 DVSS.n1139 0.00372031
R63894 DVSS.n22374 DVSS.n1109 0.00372031
R63895 DVSS.n1163 DVSS.n1142 0.00372031
R63896 DVSS.n1141 DVSS.n1133 0.00372031
R63897 DVSS.n1159 DVSS.n1143 0.00372031
R63898 DVSS.n1156 DVSS.n1132 0.00372031
R63899 DVSS.n1145 DVSS.n1144 0.00372031
R63900 DVSS.n1160 DVSS.n1131 0.00372031
R63901 DVSS.n1162 DVSS.n1147 0.00372031
R63902 DVSS.n1146 DVSS.n1130 0.00372031
R63903 DVSS.n1158 DVSS.n1148 0.00372031
R63904 DVSS.n1157 DVSS.n1129 0.00372031
R63905 DVSS.n1150 DVSS.n1149 0.00372031
R63906 DVSS.n1161 DVSS.n1128 0.00372031
R63907 DVSS.n13008 DVSS.n13007 0.00372031
R63908 DVSS.n13003 DVSS.n13002 0.00372031
R63909 DVSS.n13011 DVSS.n13010 0.00372031
R63910 DVSS.n13009 DVSS.n13001 0.00372031
R63911 DVSS.n13057 DVSS.n13013 0.00372031
R63912 DVSS.n13012 DVSS.n13000 0.00372031
R63913 DVSS.n13022 DVSS.n13021 0.00372031
R63914 DVSS.n12999 DVSS.n12998 0.00372031
R63915 DVSS.n13025 DVSS.n13024 0.00372031
R63916 DVSS.n13023 DVSS.n12997 0.00372031
R63917 DVSS.n13048 DVSS.n13027 0.00372031
R63918 DVSS.n13026 DVSS.n12996 0.00372031
R63919 DVSS.n13036 DVSS.n13035 0.00372031
R63920 DVSS.n12995 DVSS.n12994 0.00372031
R63921 DVSS.n13039 DVSS.n13038 0.00372031
R63922 DVSS.n13037 DVSS.n12993 0.00372031
R63923 DVSS.n373 DVSS.n351 0.00372031
R63924 DVSS.n348 DVSS.n347 0.00372031
R63925 DVSS.n372 DVSS.n353 0.00372031
R63926 DVSS.n352 DVSS.n346 0.00372031
R63927 DVSS.n367 DVSS.n354 0.00372031
R63928 DVSS.n374 DVSS.n345 0.00372031
R63929 DVSS.n356 DVSS.n355 0.00372031
R63930 DVSS.n344 DVSS.n343 0.00372031
R63931 DVSS.n371 DVSS.n358 0.00372031
R63932 DVSS.n357 DVSS.n342 0.00372031
R63933 DVSS.n365 DVSS.n359 0.00372031
R63934 DVSS.n375 DVSS.n341 0.00372031
R63935 DVSS.n361 DVSS.n360 0.00372031
R63936 DVSS.n340 DVSS.n339 0.00372031
R63937 DVSS.n370 DVSS.n363 0.00372031
R63938 DVSS.n362 DVSS.n338 0.00372031
R63939 DVSS.n22462 DVSS.n814 0.00372031
R63940 DVSS.n22464 DVSS.n812 0.00372031
R63941 DVSS.n22496 DVSS.n822 0.00372031
R63942 DVSS.n22491 DVSS.n811 0.00372031
R63943 DVSS.n22463 DVSS.n823 0.00372031
R63944 DVSS.n22497 DVSS.n810 0.00372031
R63945 DVSS.n22465 DVSS.n809 0.00372031
R63946 DVSS.n22495 DVSS.n832 0.00372031
R63947 DVSS.n22466 DVSS.n808 0.00372031
R63948 DVSS.n22467 DVSS.n807 0.00372031
R63949 DVSS.n22494 DVSS.n841 0.00372031
R63950 DVSS.n22468 DVSS.n806 0.00372031
R63951 DVSS.n22469 DVSS.n805 0.00372031
R63952 DVSS.n22493 DVSS.n850 0.00372031
R63953 DVSS.n22470 DVSS.n804 0.00372031
R63954 DVSS.n22471 DVSS.n803 0.00372031
R63955 DVSS.n22492 DVSS.n22461 0.00372031
R63956 DVSS.n229 DVSS.n218 0.00372031
R63957 DVSS.n231 DVSS.n216 0.00372031
R63958 DVSS.n260 DVSS.n219 0.00372031
R63959 DVSS.n255 DVSS.n215 0.00372031
R63960 DVSS.n230 DVSS.n220 0.00372031
R63961 DVSS.n261 DVSS.n214 0.00372031
R63962 DVSS.n232 DVSS.n213 0.00372031
R63963 DVSS.n259 DVSS.n222 0.00372031
R63964 DVSS.n233 DVSS.n212 0.00372031
R63965 DVSS.n234 DVSS.n211 0.00372031
R63966 DVSS.n258 DVSS.n224 0.00372031
R63967 DVSS.n235 DVSS.n210 0.00372031
R63968 DVSS.n236 DVSS.n209 0.00372031
R63969 DVSS.n257 DVSS.n226 0.00372031
R63970 DVSS.n237 DVSS.n208 0.00372031
R63971 DVSS.n238 DVSS.n207 0.00372031
R63972 DVSS.n256 DVSS.n228 0.00372031
R63973 DVSS.n149 DVSS.n138 0.00372031
R63974 DVSS.n151 DVSS.n136 0.00372031
R63975 DVSS.n180 DVSS.n139 0.00372031
R63976 DVSS.n175 DVSS.n135 0.00372031
R63977 DVSS.n150 DVSS.n140 0.00372031
R63978 DVSS.n181 DVSS.n134 0.00372031
R63979 DVSS.n152 DVSS.n133 0.00372031
R63980 DVSS.n179 DVSS.n142 0.00372031
R63981 DVSS.n153 DVSS.n132 0.00372031
R63982 DVSS.n154 DVSS.n131 0.00372031
R63983 DVSS.n178 DVSS.n144 0.00372031
R63984 DVSS.n155 DVSS.n130 0.00372031
R63985 DVSS.n156 DVSS.n129 0.00372031
R63986 DVSS.n177 DVSS.n146 0.00372031
R63987 DVSS.n157 DVSS.n128 0.00372031
R63988 DVSS.n158 DVSS.n127 0.00372031
R63989 DVSS.n176 DVSS.n148 0.00372031
R63990 DVSS.n84 DVSS.n73 0.00372031
R63991 DVSS.n86 DVSS.n71 0.00372031
R63992 DVSS.n23170 DVSS.n74 0.00372031
R63993 DVSS.n23165 DVSS.n70 0.00372031
R63994 DVSS.n85 DVSS.n75 0.00372031
R63995 DVSS.n23171 DVSS.n69 0.00372031
R63996 DVSS.n87 DVSS.n68 0.00372031
R63997 DVSS.n23169 DVSS.n77 0.00372031
R63998 DVSS.n88 DVSS.n67 0.00372031
R63999 DVSS.n89 DVSS.n66 0.00372031
R64000 DVSS.n23168 DVSS.n79 0.00372031
R64001 DVSS.n90 DVSS.n65 0.00372031
R64002 DVSS.n91 DVSS.n64 0.00372031
R64003 DVSS.n23167 DVSS.n81 0.00372031
R64004 DVSS.n92 DVSS.n63 0.00372031
R64005 DVSS.n93 DVSS.n62 0.00372031
R64006 DVSS.n23166 DVSS.n83 0.00372031
R64007 DVSS.n21923 DVSS.n21882 0.00372031
R64008 DVSS.n21881 DVSS.n21880 0.00372031
R64009 DVSS.n21924 DVSS.n21879 0.00372031
R64010 DVSS.n21891 DVSS.n21890 0.00372031
R64011 DVSS.n21925 DVSS.n21878 0.00372031
R64012 DVSS.n21926 DVSS.n21877 0.00372031
R64013 DVSS.n21901 DVSS.n21900 0.00372031
R64014 DVSS.n21927 DVSS.n21876 0.00372031
R64015 DVSS.n21928 DVSS.n21875 0.00372031
R64016 DVSS.n21911 DVSS.n21910 0.00372031
R64017 DVSS.n21929 DVSS.n21874 0.00372031
R64018 DVSS.n21930 DVSS.n21873 0.00372031
R64019 DVSS.n21921 DVSS.n21920 0.00372031
R64020 DVSS.n21931 DVSS.n21872 0.00372031
R64021 DVSS.n21933 DVSS.n21871 0.00372031
R64022 DVSS.n21943 DVSS.n21942 0.00372031
R64023 DVSS.n21945 DVSS.n21851 0.00372031
R64024 DVSS.n21604 DVSS.n21592 0.00372031
R64025 DVSS.n21621 DVSS.n21567 0.00372031
R64026 DVSS.n21605 DVSS.n21566 0.00372031
R64027 DVSS.n21620 DVSS.n21594 0.00372031
R64028 DVSS.n21606 DVSS.n21565 0.00372031
R64029 DVSS.n21607 DVSS.n21564 0.00372031
R64030 DVSS.n21619 DVSS.n21596 0.00372031
R64031 DVSS.n21608 DVSS.n21563 0.00372031
R64032 DVSS.n21609 DVSS.n21562 0.00372031
R64033 DVSS.n21618 DVSS.n21598 0.00372031
R64034 DVSS.n21610 DVSS.n21561 0.00372031
R64035 DVSS.n21611 DVSS.n21560 0.00372031
R64036 DVSS.n21617 DVSS.n21600 0.00372031
R64037 DVSS.n21612 DVSS.n21559 0.00372031
R64038 DVSS.n21613 DVSS.n21558 0.00372031
R64039 DVSS.n21616 DVSS.n21602 0.00372031
R64040 DVSS.n21614 DVSS.n21557 0.00372031
R64041 DVSS.n21707 DVSS.n21695 0.00372031
R64042 DVSS.n21724 DVSS.n21693 0.00372031
R64043 DVSS.n21708 DVSS.n21692 0.00372031
R64044 DVSS.n21723 DVSS.n21697 0.00372031
R64045 DVSS.n21709 DVSS.n21691 0.00372031
R64046 DVSS.n21710 DVSS.n21690 0.00372031
R64047 DVSS.n21722 DVSS.n21699 0.00372031
R64048 DVSS.n21711 DVSS.n21689 0.00372031
R64049 DVSS.n21712 DVSS.n21688 0.00372031
R64050 DVSS.n21721 DVSS.n21701 0.00372031
R64051 DVSS.n21713 DVSS.n21687 0.00372031
R64052 DVSS.n21714 DVSS.n21686 0.00372031
R64053 DVSS.n21720 DVSS.n21703 0.00372031
R64054 DVSS.n21715 DVSS.n21685 0.00372031
R64055 DVSS.n21716 DVSS.n21684 0.00372031
R64056 DVSS.n21719 DVSS.n21705 0.00372031
R64057 DVSS.n21717 DVSS.n21683 0.00372031
R64058 DVSS.n21800 DVSS.n21788 0.00372031
R64059 DVSS.n21817 DVSS.n21787 0.00372031
R64060 DVSS.n21801 DVSS.n21786 0.00372031
R64061 DVSS.n21816 DVSS.n21790 0.00372031
R64062 DVSS.n21802 DVSS.n21785 0.00372031
R64063 DVSS.n21803 DVSS.n21784 0.00372031
R64064 DVSS.n21815 DVSS.n21792 0.00372031
R64065 DVSS.n21804 DVSS.n21783 0.00372031
R64066 DVSS.n21805 DVSS.n21782 0.00372031
R64067 DVSS.n21814 DVSS.n21794 0.00372031
R64068 DVSS.n21806 DVSS.n21781 0.00372031
R64069 DVSS.n21807 DVSS.n21780 0.00372031
R64070 DVSS.n21813 DVSS.n21796 0.00372031
R64071 DVSS.n21808 DVSS.n21779 0.00372031
R64072 DVSS.n21809 DVSS.n21778 0.00372031
R64073 DVSS.n21812 DVSS.n21798 0.00372031
R64074 DVSS.n21810 DVSS.n21777 0.00372031
R64075 DVSS.n15807 DVSS.n15786 0.00372031
R64076 DVSS.n15808 DVSS.n15787 0.00372031
R64077 DVSS.n15809 DVSS.n15788 0.00372031
R64078 DVSS.n15810 DVSS.n15789 0.00372031
R64079 DVSS.n16263 DVSS.n16243 0.00372031
R64080 DVSS.n16264 DVSS.n16244 0.00372031
R64081 DVSS.n16262 DVSS.n16250 0.00372031
R64082 DVSS.n16265 DVSS.n16247 0.00372031
R64083 DVSS.n17641 DVSS.n16069 0.00372031
R64084 DVSS.n16088 DVSS.n16068 0.00372031
R64085 DVSS.n16095 DVSS.n16071 0.00372031
R64086 DVSS.n16094 DVSS.n16072 0.00372031
R64087 DVSS.n15304 DVSS.n15303 0.00372031
R64088 DVSS.n15302 DVSS.n15301 0.00372031
R64089 DVSS.n15299 DVSS.n15292 0.00372031
R64090 DVSS.n15297 DVSS.n15296 0.00372031
R64091 DVSS.n20007 DVSS.n14911 0.00372031
R64092 DVSS.n14902 DVSS.n14901 0.00372031
R64093 DVSS.n14900 DVSS.n14899 0.00372031
R64094 DVSS.n14898 DVSS.n14897 0.00372031
R64095 DVSS.n14896 DVSS.n14895 0.00372031
R64096 DVSS.n20848 DVSS.n14482 0.00372031
R64097 DVSS.n20815 DVSS.n14469 0.00372031
R64098 DVSS.n20816 DVSS.n14468 0.00372031
R64099 DVSS.n20817 DVSS.n14467 0.00372031
R64100 DVSS.n13954 DVSS.n13928 0.00372031
R64101 DVSS.n13955 DVSS.n13929 0.00372031
R64102 DVSS.n13956 DVSS.n13930 0.00372031
R64103 DVSS.n13957 DVSS.n13931 0.00372031
R64104 DVSS.n13958 DVSS.n13932 0.00372031
R64105 DVSS.n13959 DVSS.n13933 0.00372031
R64106 DVSS.n13960 DVSS.n13934 0.00372031
R64107 DVSS.n13961 DVSS.n13935 0.00372031
R64108 DVSS.n13962 DVSS.n13936 0.00372031
R64109 DVSS.n13963 DVSS.n13937 0.00372031
R64110 DVSS.n13964 DVSS.n13938 0.00372031
R64111 DVSS.n13966 DVSS.n13938 0.00372031
R64112 DVSS.n13967 DVSS.n13937 0.00372031
R64113 DVSS.n13968 DVSS.n13936 0.00372031
R64114 DVSS.n13969 DVSS.n13935 0.00372031
R64115 DVSS.n13970 DVSS.n13934 0.00372031
R64116 DVSS.n13971 DVSS.n13933 0.00372031
R64117 DVSS.n13972 DVSS.n13932 0.00372031
R64118 DVSS.n13973 DVSS.n13931 0.00372031
R64119 DVSS.n13974 DVSS.n13930 0.00372031
R64120 DVSS.n13975 DVSS.n13929 0.00372031
R64121 DVSS.n21104 DVSS.n13928 0.00372031
R64122 DVSS.n20817 DVSS.n14463 0.00372031
R64123 DVSS.n20816 DVSS.n14462 0.00372031
R64124 DVSS.n20815 DVSS.n14461 0.00372031
R64125 DVSS.n14482 DVSS.n14460 0.00372031
R64126 DVSS.n14895 DVSS.n14893 0.00372031
R64127 DVSS.n14897 DVSS.n14892 0.00372031
R64128 DVSS.n14899 DVSS.n14891 0.00372031
R64129 DVSS.n14901 DVSS.n14890 0.00372031
R64130 DVSS.n14911 DVSS.n14889 0.00372031
R64131 DVSS.n15296 DVSS.n14903 0.00372031
R64132 DVSS.n15300 DVSS.n15299 0.00372031
R64133 DVSS.n15301 DVSS.n15295 0.00372031
R64134 DVSS.n15303 DVSS.n15294 0.00372031
R64135 DVSS.n16092 DVSS.n16072 0.00372031
R64136 DVSS.n16091 DVSS.n16071 0.00372031
R64137 DVSS.n16090 DVSS.n16068 0.00372031
R64138 DVSS.n16089 DVSS.n16069 0.00372031
R64139 DVSS.n16265 DVSS.n16246 0.00372031
R64140 DVSS.n16262 DVSS.n16245 0.00372031
R64141 DVSS.n16264 DVSS.n16248 0.00372031
R64142 DVSS.n16263 DVSS.n16249 0.00372031
R64143 DVSS.n15810 DVSS.n15791 0.00372031
R64144 DVSS.n15809 DVSS.n15792 0.00372031
R64145 DVSS.n15808 DVSS.n15793 0.00372031
R64146 DVSS.n15807 DVSS.n15794 0.00372031
R64147 DVSS.n13597 DVSS.n13572 0.00372031
R64148 DVSS.n13588 DVSS.n13572 0.00372031
R64149 DVSS.n13598 DVSS.n13573 0.00372031
R64150 DVSS.n13589 DVSS.n13573 0.00372031
R64151 DVSS.n13599 DVSS.n13574 0.00372031
R64152 DVSS.n13600 DVSS.n13575 0.00372031
R64153 DVSS.n13590 DVSS.n13575 0.00372031
R64154 DVSS.n13590 DVSS.n13576 0.00372031
R64155 DVSS.n13600 DVSS.n13577 0.00372031
R64156 DVSS.n13589 DVSS.n13578 0.00372031
R64157 DVSS.n13599 DVSS.n13578 0.00372031
R64158 DVSS.n13588 DVSS.n13579 0.00372031
R64159 DVSS.n13598 DVSS.n13579 0.00372031
R64160 DVSS.n13597 DVSS.n13580 0.00372031
R64161 DVSS.n21377 DVSS.n13421 0.00372031
R64162 DVSS.n13432 DVSS.n13421 0.00372031
R64163 DVSS.n21378 DVSS.n13422 0.00372031
R64164 DVSS.n13433 DVSS.n13422 0.00372031
R64165 DVSS.n21379 DVSS.n13423 0.00372031
R64166 DVSS.n21380 DVSS.n13424 0.00372031
R64167 DVSS.n13434 DVSS.n13424 0.00372031
R64168 DVSS.n13434 DVSS.n13425 0.00372031
R64169 DVSS.n21380 DVSS.n13426 0.00372031
R64170 DVSS.n13433 DVSS.n13427 0.00372031
R64171 DVSS.n21379 DVSS.n13427 0.00372031
R64172 DVSS.n13432 DVSS.n13428 0.00372031
R64173 DVSS.n21378 DVSS.n13428 0.00372031
R64174 DVSS.n21377 DVSS.n13429 0.00372031
R64175 DVSS.n16634 DVSS.n16320 0.00371429
R64176 DVSS.n16709 DVSS.n16163 0.00371429
R64177 DVSS.n16057 DVSS.n16027 0.00371429
R64178 DVSS.n16874 DVSS.n16848 0.00371429
R64179 DVSS.n15280 DVSS.n15251 0.00371429
R64180 DVSS.n15418 DVSS.n15392 0.00371429
R64181 DVSS.n18424 DVSS.n18392 0.00371429
R64182 DVSS.n14980 DVSS.n14955 0.00371429
R64183 DVSS.n20795 DVSS.n20718 0.00371429
R64184 DVSS.n20878 DVSS.n14438 0.00371429
R64185 DVSS.n21252 DVSS.n13604 0.00371429
R64186 DVSS.n21328 DVSS.n13494 0.00371429
R64187 DVSS.n22710 DVSS.n687 0.00371429
R64188 DVSS.n22786 DVSS.n579 0.00371429
R64189 DVSS.n18344 DVSS.n15306 0.00370488
R64190 DVSS.n22756 DVSS.n607 0.00370488
R64191 DVSS.n18326 DVSS.n15373 0.00370488
R64192 DVSS.n22797 DVSS.n562 0.00370488
R64193 DVSS.n18379 DVSS.n15267 0.00370488
R64194 DVSS.n22714 DVSS.n669 0.00370488
R64195 DVSS.n18315 DVSS.n15443 0.00370488
R64196 DVSS.n22838 DVSS.n507 0.00370488
R64197 DVSS.n13824 DVSS.n13818 0.00368
R64198 DVSS.n21511 DVSS.n1059 0.00368
R64199 DVSS.n22478 DVSS.n785 0.00368
R64200 DVSS.n21858 DVSS.n1437 0.00368
R64201 DVSS.n22223 DVSS.n709 0.00367368
R64202 DVSS.n22153 DVSS.n22124 0.00367368
R64203 DVSS.n932 DVSS.n906 0.00367368
R64204 DVSS.n22427 DVSS.n1002 0.00367368
R64205 DVSS.n22238 DVSS.n467 0.00367368
R64206 DVSS.n22308 DVSS.n1242 0.00367368
R64207 DVSS.n12827 DVSS.n18 0.00367368
R64208 DVSS.n12921 DVSS.n12818 0.00367368
R64209 DVSS.n17803 DVSS.n15903 0.00366901
R64210 DVSS.n16746 DVSS.n15599 0.00365
R64211 DVSS.n15528 DVSS.n15500 0.00365
R64212 DVSS.n18258 DVSS.n18227 0.00365
R64213 DVSS.n15122 DVSS.n15111 0.00365
R64214 DVSS.n20951 DVSS.n14345 0.00365
R64215 DVSS.n21405 DVSS.n13403 0.00365
R64216 DVSS.n22874 DVSS.n483 0.00365
R64217 DVSS.n13908 DVSS.n13875 0.00362
R64218 DVSS.n14091 DVSS.n14071 0.00362
R64219 DVSS.n1477 DVSS.n1055 0.00362
R64220 DVSS.n12983 DVSS.n12976 0.00362
R64221 DVSS.n22488 DVSS.n22474 0.00362
R64222 DVSS.n195 DVSS.n162 0.00362
R64223 DVSS.n21854 DVSS.n1446 0.00362
R64224 DVSS.n21728 DVSS.n21677 0.00362
R64225 DVSS.n21906 DVSS.n21597 0.00361707
R64226 DVSS.n846 DVSS.n225 0.00361707
R64227 DVSS.n21903 DVSS.n21700 0.00361707
R64228 DVSS.n843 DVSS.n145 0.00361707
R64229 DVSS.n21909 DVSS.n21908 0.00361707
R64230 DVSS.n849 DVSS.n848 0.00361707
R64231 DVSS.n21902 DVSS.n21793 0.00361707
R64232 DVSS.n842 DVSS.n80 0.00361707
R64233 DVSS.n17877 DVSS.n15813 0.00359859
R64234 DVSS.n21041 DVSS.n14254 0.00359
R64235 DVSS.n12780 DVSS.n412 0.00359
R64236 DVSS.n23206 DVSS.n32 0.00359
R64237 DVSS.n21978 DVSS.n1227 0.00359
R64238 DVSS.n16255 DVSS.n16241 0.00358571
R64239 DVSS.n16780 DVSS.n15654 0.00358571
R64240 DVSS.n16099 DVSS.n16087 0.00358571
R64241 DVSS.n17555 DVSS.n17540 0.00358571
R64242 DVSS.n15324 DVSS.n15309 0.00358571
R64243 DVSS.n15475 DVSS.n15460 0.00358571
R64244 DVSS.n14908 DVSS.n14888 0.00358571
R64245 DVSS.n15072 DVSS.n15071 0.00358571
R64246 DVSS.n14475 DVSS.n14459 0.00358571
R64247 DVSS.n20926 DVSS.n14395 0.00358571
R64248 DVSS.n13533 DVSS.n13516 0.00358571
R64249 DVSS.n21376 DVSS.n13436 0.00358571
R64250 DVSS.n612 DVSS.n596 0.00358571
R64251 DVSS.n532 DVSS.n516 0.00358571
R64252 DVSS.n22183 DVSS.n22130 0.00357895
R64253 DVSS.n964 DVSS.n923 0.00357895
R64254 DVSS.n22397 DVSS.n1008 0.00357895
R64255 DVSS.n22278 DVSS.n1248 0.00357895
R64256 DVSS.n12859 DVSS.n7 0.00357895
R64257 DVSS.n12891 DVSS.n12812 0.00357895
R64258 DVSS.n14118 DVSS.n14056 0.00356
R64259 DVSS.n21065 DVSS.n21064 0.00356
R64260 DVSS.n12972 DVSS.n312 0.00356
R64261 DVSS.n23002 DVSS.n23001 0.00356
R64262 DVSS.n23135 DVSS.n159 0.00356
R64263 DVSS.n23183 DVSS.n23182 0.00356
R64264 DVSS.n21752 DVSS.n21718 0.00356
R64265 DVSS.n21965 DVSS.n21964 0.00356
R64266 DVSS.n21647 DVSS.n271 0.00356
R64267 DVSS.n23077 DVSS.n23075 0.00356
R64268 DVSS.n23069 DVSS.n270 0.00356
R64269 DVSS.n19311 DVSS.n19309 0.00355644
R64270 DVSS.n19310 DVSS.n19307 0.00355644
R64271 DVSS.n19311 DVSS.n19310 0.00355644
R64272 DVSS.n19313 DVSS.n19309 0.00355644
R64273 DVSS.n19655 DVSS.n19654 0.00355644
R64274 DVSS.n19655 DVSS.n13399 0.00355644
R64275 DVSS.n19654 DVSS.n19140 0.00355644
R64276 DVSS.n19140 DVSS.n19138 0.00355644
R64277 DVSS.n18953 DVSS.n18879 0.00353371
R64278 DVSS.n20157 DVSS.n14611 0.00353371
R64279 DVSS.n20653 DVSS.n14625 0.00353371
R64280 DVSS.n20284 DVSS 0.00353371
R64281 DVSS.n20346 DVSS.n14690 0.00353371
R64282 DVSS.n16541 DVSS.n16540 0.00353158
R64283 DVSS.n18108 DVSS.n18107 0.00353158
R64284 DVSS DVSS.n1 0.00353
R64285 DVSS DVSS.n23227 0.00353
R64286 DVSS.n21886 DVSS.n21567 0.00352927
R64287 DVSS.n828 DVSS.n214 0.00352927
R64288 DVSS.n13042 DVSS.n1128 0.00352927
R64289 DVSS.n21884 DVSS.n21693 0.00352927
R64290 DVSS.n825 DVSS.n134 0.00352927
R64291 DVSS.n13046 DVSS.n12993 0.00352927
R64292 DVSS.n21888 DVSS.n21880 0.00352927
R64293 DVSS.n830 DVSS.n810 0.00352927
R64294 DVSS.n13041 DVSS.n1070 0.00352927
R64295 DVSS.n21883 DVSS.n21787 0.00352927
R64296 DVSS.n824 DVSS.n69 0.00352927
R64297 DVSS.n13040 DVSS.n338 0.00352927
R64298 DVSS.n15911 DVSS.n15895 0.00352817
R64299 DVSS.n16595 DVSS.n16594 0.00352143
R64300 DVSS.n15964 DVSS.n15954 0.00352143
R64301 DVSS.n17711 DVSS.n17690 0.00352143
R64302 DVSS.n15217 DVSS.n15183 0.00352143
R64303 DVSS.n20762 DVSS.n13719 0.00352143
R64304 DVSS.n21213 DVSS.n21212 0.00352143
R64305 DVSS.n22646 DVSS.n721 0.00352143
R64306 DVSS.n13980 DVSS.n13951 0.0035
R64307 DVSS.n14215 DVSS.n14185 0.0035
R64308 DVSS.n1121 DVSS.n284 0.0035
R64309 DVSS.n390 DVSS.n327 0.0035
R64310 DVSS.n23084 DVSS.n252 0.0035
R64311 DVSS.n113 DVSS.n106 0.0035
R64312 DVSS.n21643 DVSS.n21634 0.0035
R64313 DVSS.n21957 DVSS.n21767 0.0035
R64314 DVSS.n22137 DVSS.n1391 0.00348421
R64315 DVSS.n948 DVSS.n917 0.00348421
R64316 DVSS.n22324 DVSS.n1223 0.00348421
R64317 DVSS.n12843 DVSS.n11 0.00348421
R64318 DVSS.n12773 DVSS.n12351 0.00347744
R64319 DVSS.n13805 DVSS.n13732 0.00347
R64320 DVSS.n1492 DVSS.n975 0.00347
R64321 DVSS.n885 DVSS.n768 0.00347
R64322 DVSS.n1422 DVSS.n1366 0.00347
R64323 DVSS.n17893 DVSS.n15818 0.00345775
R64324 DVSS.n17972 DVSS.n15700 0.00345775
R64325 DVSS.n16662 DVSS.n16259 0.00345714
R64326 DVSS.n16796 DVSS.n15658 0.00345714
R64327 DVSS.n16124 DVSS.n16078 0.00345714
R64328 DVSS.n17597 DVSS.n17545 0.00345714
R64329 DVSS.n15339 DVSS.n15313 0.00345714
R64330 DVSS.n18307 DVSS.n15465 0.00345714
R64331 DVSS.n18442 DVSS.n14879 0.00345714
R64332 DVSS.n15051 DVSS.n15022 0.00345714
R64333 DVSS.n20830 DVSS.n14479 0.00345714
R64334 DVSS.n20909 DVSS.n14381 0.00345714
R64335 DVSS.n21280 DVSS.n13537 0.00345714
R64336 DVSS.n21359 DVSS.n13440 0.00345714
R64337 DVSS.n22738 DVSS.n619 0.00345714
R64338 DVSS.n22817 DVSS.n520 0.00345714
R64339 DVSS.n13990 DVSS.n13948 0.00344
R64340 DVSS.n1464 DVSS.n1116 0.00344
R64341 DVSS.n22512 DVSS.n247 0.00344
R64342 DVSS.n21630 DVSS.n1461 0.00344
R64343 DVSS.n20689 DVSS.n14549 0.00343478
R64344 DVSS.n14561 DVSS.n14560 0.00343478
R64345 DVSS.n14593 DVSS.n14584 0.00343478
R64346 DVSS.n20123 DVSS.n14592 0.00343478
R64347 DVSS.n20310 DVSS.n14634 0.00343478
R64348 DVSS.n14651 DVSS.n14650 0.00343478
R64349 DVSS.n20431 DVSS.n20430 0.00343478
R64350 DVSS.n20357 DVSS.n20356 0.00343478
R64351 DVSS.n14538 DVSS.n14523 0.00343478
R64352 DVSS.n14540 DVSS.n14537 0.00343478
R64353 DVSS.n20110 DVSS.n20109 0.00343478
R64354 DVSS.n20112 DVSS.n20017 0.00343478
R64355 DVSS.n20195 DVSS.n14866 0.00343478
R64356 DVSS.n20194 DVSS.n14863 0.00343478
R64357 DVSS.n20363 DVSS.n20362 0.00343478
R64358 DVSS.n20350 DVSS.n14856 0.00343478
R64359 DVSS.n13796 DVSS.n13739 0.00341
R64360 DVSS.n1496 DVSS.n985 0.00341
R64361 DVSS.n898 DVSS.n763 0.00341
R64362 DVSS.n1414 DVSS.n1373 0.00341
R64363 DVSS.n3414 DVSS.n3407 0.00339933
R64364 DVSS.n11628 DVSS.n11621 0.00339933
R64365 DVSS.n3412 DVSS.n3408 0.00339933
R64366 DVSS.n11626 DVSS.n11623 0.00339933
R64367 DVSS.n20042 DVSS.n14466 0.00339756
R64368 DVSS.n20045 DVSS.n14464 0.00339756
R64369 DVSS.n20046 DVSS.n14465 0.00339756
R64370 DVSS.n20209 DVSS.n14418 0.00339756
R64371 DVSS.n20211 DVSS.n14415 0.00339756
R64372 DVSS.n20212 DVSS.n14416 0.00339756
R64373 DVSS.n18871 DVSS.n14513 0.00339756
R64374 DVSS.n18873 DVSS.n14511 0.00339756
R64375 DVSS.n18984 DVSS.n14512 0.00339756
R64376 DVSS.n14675 DVSS.n14369 0.00339756
R64377 DVSS.n14677 DVSS.n14366 0.00339756
R64378 DVSS.n20626 DVSS.n14367 0.00339756
R64379 DVSS.n16577 DVSS.n16554 0.00339286
R64380 DVSS.n15972 DVSS.n15950 0.00339286
R64381 DVSS.n17729 DVSS.n17685 0.00339286
R64382 DVSS.n15192 DVSS.n15178 0.00339286
R64383 DVSS.n20746 DVSS.n13715 0.00339286
R64384 DVSS.n21190 DVSS.n13645 0.00339286
R64385 DVSS.n22662 DVSS.n726 0.00339286
R64386 DVSS.n22137 DVSS.n22120 0.00338947
R64387 DVSS.n948 DVSS.n902 0.00338947
R64388 DVSS.n22440 DVSS.n970 0.00338947
R64389 DVSS.n22326 DVSS.n1223 0.00338947
R64390 DVSS.n12843 DVSS.n22 0.00338947
R64391 DVSS.n12875 DVSS.n12808 0.00338947
R64392 DVSS.n13983 DVSS.n13944 0.00338
R64393 DVSS.n14206 DVSS.n14178 0.00338
R64394 DVSS.n1112 DVSS.n279 0.00338
R64395 DVSS.n380 DVSS.n322 0.00338
R64396 DVSS.n23076 DVSS.n242 0.00338
R64397 DVSS.n117 DVSS.n98 0.00338
R64398 DVSS.n21625 DVSS.n21591 0.00338
R64399 DVSS.n21822 DVSS.n21762 0.00338
R64400 DVSS.n17456 DVSS.n17434 0.00336948
R64401 DVSS.n17423 DVSS.n17199 0.00336948
R64402 DVSS.n16937 DVSS.n16936 0.00336948
R64403 DVSS.n13092 DVSS.n384 0.00336948
R64404 DVSS.n13093 DVSS.n13092 0.00336948
R64405 DVSS.n16938 DVSS.n16937 0.00336948
R64406 DVSS.n17425 DVSS.n17199 0.00336948
R64407 DVSS.n17452 DVSS.n17434 0.00336948
R64408 DVSS.n17475 DVSS.n17140 0.00336948
R64409 DVSS.n17141 DVSS.n17138 0.00336948
R64410 DVSS.n17408 DVSS.n17260 0.00336948
R64411 DVSS.n17406 DVSS.n17261 0.00336948
R64412 DVSS.n17366 DVSS.n17359 0.00336948
R64413 DVSS.n20010 DVSS.n14470 0.00336948
R64414 DVSS.n20673 DVSS.n14585 0.00336948
R64415 DVSS.n19216 DVSS.n19171 0.00336948
R64416 DVSS.n19170 DVSS.n19041 0.00336948
R64417 DVSS.n19592 DVSS.n19252 0.00336948
R64418 DVSS.n21586 DVSS.n21568 0.00336948
R64419 DVSS.n22369 DVSS.n1165 0.00336948
R64420 DVSS.n21589 DVSS.n21568 0.00336948
R64421 DVSS.n14585 DVSS.n13947 0.00336948
R64422 DVSS.n20173 DVSS.n20010 0.00336948
R64423 DVSS.n17359 DVSS.n17332 0.00336948
R64424 DVSS.n17408 DVSS.n17261 0.00336948
R64425 DVSS.n17260 DVSS.n17259 0.00336948
R64426 DVSS.n17475 DVSS.n17141 0.00336948
R64427 DVSS.n17140 DVSS.n16081 0.00336948
R64428 DVSS.n17468 DVSS.n17175 0.00336948
R64429 DVSS.n17459 DVSS.n17173 0.00336948
R64430 DVSS.n17416 DVSS.n17225 0.00336948
R64431 DVSS.n17414 DVSS.n17226 0.00336948
R64432 DVSS.n17492 DVSS.n16941 0.00336948
R64433 DVSS.n14865 DVSS.n14425 0.00336948
R64434 DVSS.n20647 DVSS.n14633 0.00336948
R64435 DVSS.n19161 DVSS.n19157 0.00336948
R64436 DVSS.n19159 DVSS.n19158 0.00336948
R64437 DVSS.n19089 DVSS.n19069 0.00336948
R64438 DVSS.n1197 DVSS.n1179 0.00336948
R64439 DVSS.n12961 DVSS.n12960 0.00336948
R64440 DVSS.n22339 DVSS.n1179 0.00336948
R64441 DVSS.n14633 DVSS.n14631 0.00336948
R64442 DVSS.n20316 DVSS.n14865 0.00336948
R64443 DVSS.n16941 DVSS.n16940 0.00336948
R64444 DVSS.n17416 DVSS.n17226 0.00336948
R64445 DVSS.n17225 DVSS.n17224 0.00336948
R64446 DVSS.n17468 DVSS.n17459 0.00336948
R64447 DVSS.n17470 DVSS.n17175 0.00336948
R64448 DVSS.n17121 DVSS.n17119 0.00336948
R64449 DVSS.n17301 DVSS.n17295 0.00336948
R64450 DVSS.n17403 DVSS.n17303 0.00336948
R64451 DVSS.n17401 DVSS.n17304 0.00336948
R64452 DVSS.n17327 DVSS.n17312 0.00336948
R64453 DVSS.n20699 DVSS.n14517 0.00336948
R64454 DVSS.n14550 DVSS.n14548 0.00336948
R64455 DVSS.n19029 DVSS.n19004 0.00336948
R64456 DVSS.n19899 DVSS.n19031 0.00336948
R64457 DVSS.n19515 DVSS.n19269 0.00336948
R64458 DVSS.n22460 DVSS.n858 0.00336948
R64459 DVSS.n22383 DVSS.n1044 0.00336948
R64460 DVSS.n22458 DVSS.n858 0.00336948
R64461 DVSS.n20688 DVSS.n14550 0.00336948
R64462 DVSS.n20697 DVSS.n14517 0.00336948
R64463 DVSS.n17372 DVSS.n17327 0.00336948
R64464 DVSS.n17403 DVSS.n17304 0.00336948
R64465 DVSS.n17303 DVSS.n17302 0.00336948
R64466 DVSS.n17295 DVSS.n17119 0.00336948
R64467 DVSS.n17479 DVSS.n17121 0.00336948
R64468 DVSS.n19512 DVSS.n19269 0.00336948
R64469 DVSS.n19252 DVSS.n19065 0.00336948
R64470 DVSS.n19850 DVSS.n19069 0.00336948
R64471 DVSS.n19031 DVSS.n19029 0.00336948
R64472 DVSS.n19171 DVSS.n19170 0.00336948
R64473 DVSS.n19158 DVSS.n19157 0.00336948
R64474 DVSS.n19901 DVSS.n19004 0.00336948
R64475 DVSS.n19249 DVSS.n19216 0.00336948
R64476 DVSS.n19623 DVSS.n19161 0.00336948
R64477 DVSS.n1044 DVSS.n1015 0.00336948
R64478 DVSS.n22371 DVSS.n1165 0.00336948
R64479 DVSS.n12960 DVSS.n12959 0.00336948
R64480 DVSS.n17445 DVSS.n17426 0.00336948
R64481 DVSS.n17210 DVSS.n17209 0.00336948
R64482 DVSS.n14854 DVSS.n14376 0.00336948
R64483 DVSS.n20450 DVSS.n13430 0.00336948
R64484 DVSS.n19148 DVSS.n19142 0.00336948
R64485 DVSS.n19146 DVSS.n19143 0.00336948
R64486 DVSS.n19109 DVSS.n19091 0.00336948
R64487 DVSS.n1218 DVSS.n1200 0.00336948
R64488 DVSS.n19143 DVSS.n19142 0.00336948
R64489 DVSS.n19651 DVSS.n19148 0.00336948
R64490 DVSS.n19847 DVSS.n19091 0.00336948
R64491 DVSS.n22336 DVSS.n1200 0.00336948
R64492 DVSS.n20450 DVSS.n14668 0.00336948
R64493 DVSS.n20458 DVSS.n14854 0.00336948
R64494 DVSS.n17423 DVSS.n17210 0.00336948
R64495 DVSS.n17452 DVSS.n17445 0.00336948
R64496 DVSS.n13779 DVSS.n13744 0.00335
R64497 DVSS.n21494 DVSS.n981 0.00335
R64498 DVSS.n892 DVSS.n772 0.00335
R64499 DVSS.n1428 DVSS.n1377 0.00335
R64500 DVSS.n1409 DVSS.n1405 0.00334793
R64501 DVSS.n22569 DVSS.n759 0.00334793
R64502 DVSS.n21476 DVSS.n21475 0.00334793
R64503 DVSS.n21480 DVSS.n1499 0.00334
R64504 DVSS.n21481 DVSS.n21480 0.00334
R64505 DVSS.n21482 DVSS.n21481 0.00334
R64506 DVSS.n21482 DVSS.n1495 0.00334
R64507 DVSS.n21488 DVSS.n1495 0.00334
R64508 DVSS.n21489 DVSS.n21488 0.00334
R64509 DVSS.n21490 DVSS.n21489 0.00334
R64510 DVSS.n21490 DVSS.n1491 0.00334
R64511 DVSS.n21496 DVSS.n1491 0.00334
R64512 DVSS.n21497 DVSS.n21496 0.00334
R64513 DVSS.n21498 DVSS.n21497 0.00334
R64514 DVSS.n21498 DVSS.n1487 0.00334
R64515 DVSS.n21504 DVSS.n1487 0.00334
R64516 DVSS.n21507 DVSS.n21506 0.00334
R64517 DVSS.n21506 DVSS.n1482 0.00334
R64518 DVSS.n21515 DVSS.n1482 0.00334
R64519 DVSS.n21516 DVSS.n21515 0.00334
R64520 DVSS.n21517 DVSS.n21516 0.00334
R64521 DVSS.n21517 DVSS.n1478 0.00334
R64522 DVSS.n21523 DVSS.n1478 0.00334
R64523 DVSS.n21524 DVSS.n21523 0.00334
R64524 DVSS.n21525 DVSS.n21524 0.00334
R64525 DVSS.n21525 DVSS.n1474 0.00334
R64526 DVSS.n21531 DVSS.n1474 0.00334
R64527 DVSS.n21532 DVSS.n21531 0.00334
R64528 DVSS.n21533 DVSS.n21532 0.00334
R64529 DVSS.n21533 DVSS.n1470 0.00334
R64530 DVSS.n21538 DVSS.n1470 0.00334
R64531 DVSS.n21539 DVSS.n21538 0.00334
R64532 DVSS.n21541 DVSS.n21539 0.00334
R64533 DVSS.n21541 DVSS.n21540 0.00334
R64534 DVSS.n21540 DVSS.n1467 0.00334
R64535 DVSS.n21549 DVSS.n1467 0.00334
R64536 DVSS.n21550 DVSS.n21549 0.00334
R64537 DVSS.n21551 DVSS.n21550 0.00334
R64538 DVSS.n21551 DVSS.n277 0.00334
R64539 DVSS.n23070 DVSS.n278 0.00334
R64540 DVSS.n23066 DVSS.n278 0.00334
R64541 DVSS.n23066 DVSS.n23065 0.00334
R64542 DVSS.n23065 DVSS.n23064 0.00334
R64543 DVSS.n23064 DVSS.n283 0.00334
R64544 DVSS.n23060 DVSS.n283 0.00334
R64545 DVSS.n23060 DVSS.n23059 0.00334
R64546 DVSS.n23059 DVSS.n23058 0.00334
R64547 DVSS.n23058 DVSS.n288 0.00334
R64548 DVSS.n23054 DVSS.n288 0.00334
R64549 DVSS.n23054 DVSS.n23053 0.00334
R64550 DVSS.n23053 DVSS.n23052 0.00334
R64551 DVSS.n23052 DVSS.n293 0.00334
R64552 DVSS.n23048 DVSS.n293 0.00334
R64553 DVSS.n23048 DVSS.n23047 0.00334
R64554 DVSS.n23047 DVSS.n23046 0.00334
R64555 DVSS.n23046 DVSS.n299 0.00334
R64556 DVSS.n23042 DVSS.n299 0.00334
R64557 DVSS.n23042 DVSS.n23041 0.00334
R64558 DVSS.n23041 DVSS.n23040 0.00334
R64559 DVSS.n23040 DVSS.n304 0.00334
R64560 DVSS.n23036 DVSS.n304 0.00334
R64561 DVSS.n23036 DVSS.n23035 0.00334
R64562 DVSS.n23033 DVSS.n309 0.00334
R64563 DVSS.n23029 DVSS.n309 0.00334
R64564 DVSS.n23029 DVSS.n23028 0.00334
R64565 DVSS.n23028 DVSS.n23027 0.00334
R64566 DVSS.n23027 DVSS.n314 0.00334
R64567 DVSS.n23023 DVSS.n314 0.00334
R64568 DVSS.n23023 DVSS.n23022 0.00334
R64569 DVSS.n23022 DVSS.n23021 0.00334
R64570 DVSS.n23021 DVSS.n319 0.00334
R64571 DVSS.n23017 DVSS.n319 0.00334
R64572 DVSS.n23017 DVSS.n23016 0.00334
R64573 DVSS.n23016 DVSS.n23015 0.00334
R64574 DVSS.n23015 DVSS.n324 0.00334
R64575 DVSS.n23011 DVSS.n324 0.00334
R64576 DVSS.n23011 DVSS.n23010 0.00334
R64577 DVSS.n23010 DVSS.n23009 0.00334
R64578 DVSS.n23009 DVSS.n329 0.00334
R64579 DVSS.n332 DVSS.n329 0.00334
R64580 DVSS.n399 DVSS.n332 0.00334
R64581 DVSS.n400 DVSS.n399 0.00334
R64582 DVSS.n22999 DVSS.n400 0.00334
R64583 DVSS.n22999 DVSS.n22998 0.00334
R64584 DVSS.n22998 DVSS.n22997 0.00334
R64585 DVSS.n22993 DVSS.n22992 0.00334
R64586 DVSS.n22992 DVSS.n22991 0.00334
R64587 DVSS.n22991 DVSS.n405 0.00334
R64588 DVSS.n22987 DVSS.n405 0.00334
R64589 DVSS.n22987 DVSS.n22986 0.00334
R64590 DVSS.n22986 DVSS.n22985 0.00334
R64591 DVSS.n22985 DVSS.n410 0.00334
R64592 DVSS.n22981 DVSS.n410 0.00334
R64593 DVSS.n22981 DVSS.n22980 0.00334
R64594 DVSS.n22980 DVSS.n22979 0.00334
R64595 DVSS.n22979 DVSS.n415 0.00334
R64596 DVSS.n22975 DVSS.n22974 0.00334
R64597 DVSS.n22568 DVSS.n760 0.00334
R64598 DVSS.n22564 DVSS.n760 0.00334
R64599 DVSS.n22564 DVSS.n22563 0.00334
R64600 DVSS.n22563 DVSS.n22562 0.00334
R64601 DVSS.n22562 DVSS.n765 0.00334
R64602 DVSS.n22558 DVSS.n765 0.00334
R64603 DVSS.n22558 DVSS.n22557 0.00334
R64604 DVSS.n22557 DVSS.n22556 0.00334
R64605 DVSS.n22556 DVSS.n770 0.00334
R64606 DVSS.n22552 DVSS.n770 0.00334
R64607 DVSS.n22552 DVSS.n22551 0.00334
R64608 DVSS.n22551 DVSS.n22550 0.00334
R64609 DVSS.n22550 DVSS.n775 0.00334
R64610 DVSS.n22545 DVSS.n22544 0.00334
R64611 DVSS.n22544 DVSS.n22543 0.00334
R64612 DVSS.n22543 DVSS.n783 0.00334
R64613 DVSS.n22539 DVSS.n783 0.00334
R64614 DVSS.n22539 DVSS.n22538 0.00334
R64615 DVSS.n22538 DVSS.n22537 0.00334
R64616 DVSS.n22537 DVSS.n789 0.00334
R64617 DVSS.n22533 DVSS.n789 0.00334
R64618 DVSS.n22533 DVSS.n22532 0.00334
R64619 DVSS.n22532 DVSS.n22531 0.00334
R64620 DVSS.n22531 DVSS.n794 0.00334
R64621 DVSS.n22527 DVSS.n794 0.00334
R64622 DVSS.n22527 DVSS.n22526 0.00334
R64623 DVSS.n22526 DVSS.n22525 0.00334
R64624 DVSS.n22525 DVSS.n799 0.00334
R64625 DVSS.n22521 DVSS.n799 0.00334
R64626 DVSS.n22521 DVSS.n22520 0.00334
R64627 DVSS.n22520 DVSS.n22519 0.00334
R64628 DVSS.n22519 DVSS.n22507 0.00334
R64629 DVSS.n22515 DVSS.n22507 0.00334
R64630 DVSS.n22515 DVSS.n22514 0.00334
R64631 DVSS.n22514 DVSS.n275 0.00334
R64632 DVSS.n23073 DVSS.n275 0.00334
R64633 DVSS.n23080 DVSS.n269 0.00334
R64634 DVSS.n23081 DVSS.n23080 0.00334
R64635 DVSS.n23082 DVSS.n23081 0.00334
R64636 DVSS.n23082 DVSS.n265 0.00334
R64637 DVSS.n23088 DVSS.n265 0.00334
R64638 DVSS.n23089 DVSS.n23088 0.00334
R64639 DVSS.n23090 DVSS.n23089 0.00334
R64640 DVSS.n23090 DVSS.n203 0.00334
R64641 DVSS.n23098 DVSS.n203 0.00334
R64642 DVSS.n23099 DVSS.n23098 0.00334
R64643 DVSS.n23100 DVSS.n23099 0.00334
R64644 DVSS.n23100 DVSS.n199 0.00334
R64645 DVSS.n23107 DVSS.n199 0.00334
R64646 DVSS.n23108 DVSS.n23107 0.00334
R64647 DVSS.n23109 DVSS.n23108 0.00334
R64648 DVSS.n23109 DVSS.n196 0.00334
R64649 DVSS.n23115 DVSS.n196 0.00334
R64650 DVSS.n23116 DVSS.n23115 0.00334
R64651 DVSS.n23117 DVSS.n23116 0.00334
R64652 DVSS.n23117 DVSS.n192 0.00334
R64653 DVSS.n23123 DVSS.n192 0.00334
R64654 DVSS.n23124 DVSS.n23123 0.00334
R64655 DVSS.n23125 DVSS.n23124 0.00334
R64656 DVSS.n23131 DVSS.n23130 0.00334
R64657 DVSS.n23133 DVSS.n23131 0.00334
R64658 DVSS.n23133 DVSS.n23132 0.00334
R64659 DVSS.n23132 DVSS.n123 0.00334
R64660 DVSS.n23143 DVSS.n123 0.00334
R64661 DVSS.n23144 DVSS.n23143 0.00334
R64662 DVSS.n23145 DVSS.n23144 0.00334
R64663 DVSS.n23145 DVSS.n120 0.00334
R64664 DVSS.n23151 DVSS.n120 0.00334
R64665 DVSS.n23152 DVSS.n23151 0.00334
R64666 DVSS.n23153 DVSS.n23152 0.00334
R64667 DVSS.n23153 DVSS.n116 0.00334
R64668 DVSS.n23159 DVSS.n116 0.00334
R64669 DVSS.n23160 DVSS.n23159 0.00334
R64670 DVSS.n23161 DVSS.n23160 0.00334
R64671 DVSS.n23161 DVSS.n112 0.00334
R64672 DVSS.n23175 DVSS.n112 0.00334
R64673 DVSS.n23176 DVSS.n23175 0.00334
R64674 DVSS.n23177 DVSS.n23176 0.00334
R64675 DVSS.n23177 DVSS.n58 0.00334
R64676 DVSS.n23185 DVSS.n58 0.00334
R64677 DVSS.n23186 DVSS.n23185 0.00334
R64678 DVSS.n23187 DVSS.n23186 0.00334
R64679 DVSS.n23195 DVSS.n23194 0.00334
R64680 DVSS.n23196 DVSS.n23195 0.00334
R64681 DVSS.n23196 DVSS.n49 0.00334
R64682 DVSS.n23202 DVSS.n49 0.00334
R64683 DVSS.n23203 DVSS.n23202 0.00334
R64684 DVSS.n23204 DVSS.n23203 0.00334
R64685 DVSS.n23204 DVSS.n45 0.00334
R64686 DVSS.n23210 DVSS.n45 0.00334
R64687 DVSS.n23211 DVSS.n23210 0.00334
R64688 DVSS.n23213 DVSS.n23211 0.00334
R64689 DVSS.n23213 DVSS.n23212 0.00334
R64690 DVSS.n23226 DVSS.n23225 0.00334
R64691 DVSS.n1410 DVSS.n1404 0.00334
R64692 DVSS.n1416 DVSS.n1404 0.00334
R64693 DVSS.n1417 DVSS.n1416 0.00334
R64694 DVSS.n1418 DVSS.n1417 0.00334
R64695 DVSS.n1418 DVSS.n1400 0.00334
R64696 DVSS.n1424 DVSS.n1400 0.00334
R64697 DVSS.n1425 DVSS.n1424 0.00334
R64698 DVSS.n1426 DVSS.n1425 0.00334
R64699 DVSS.n1426 DVSS.n1396 0.00334
R64700 DVSS.n1432 DVSS.n1396 0.00334
R64701 DVSS.n1433 DVSS.n1432 0.00334
R64702 DVSS.n22117 DVSS.n1433 0.00334
R64703 DVSS.n22117 DVSS.n22116 0.00334
R64704 DVSS.n22114 DVSS.n1434 0.00334
R64705 DVSS.n22110 DVSS.n1434 0.00334
R64706 DVSS.n22110 DVSS.n22109 0.00334
R64707 DVSS.n22109 DVSS.n22108 0.00334
R64708 DVSS.n22108 DVSS.n1439 0.00334
R64709 DVSS.n22104 DVSS.n1439 0.00334
R64710 DVSS.n22104 DVSS.n22103 0.00334
R64711 DVSS.n22103 DVSS.n22102 0.00334
R64712 DVSS.n22102 DVSS.n1444 0.00334
R64713 DVSS.n22098 DVSS.n1444 0.00334
R64714 DVSS.n22098 DVSS.n22097 0.00334
R64715 DVSS.n22097 DVSS.n22096 0.00334
R64716 DVSS.n22096 DVSS.n1449 0.00334
R64717 DVSS.n22092 DVSS.n1449 0.00334
R64718 DVSS.n22092 DVSS.n22091 0.00334
R64719 DVSS.n22091 DVSS.n22090 0.00334
R64720 DVSS.n22090 DVSS.n1454 0.00334
R64721 DVSS.n22086 DVSS.n1454 0.00334
R64722 DVSS.n22086 DVSS.n22085 0.00334
R64723 DVSS.n22085 DVSS.n22084 0.00334
R64724 DVSS.n22084 DVSS.n1459 0.00334
R64725 DVSS.n22080 DVSS.n1459 0.00334
R64726 DVSS.n22080 DVSS.n22079 0.00334
R64727 DVSS.n21650 DVSS.n21649 0.00334
R64728 DVSS.n21650 DVSS.n21646 0.00334
R64729 DVSS.n21656 DVSS.n21646 0.00334
R64730 DVSS.n21657 DVSS.n21656 0.00334
R64731 DVSS.n21658 DVSS.n21657 0.00334
R64732 DVSS.n21658 DVSS.n21642 0.00334
R64733 DVSS.n21664 DVSS.n21642 0.00334
R64734 DVSS.n21665 DVSS.n21664 0.00334
R64735 DVSS.n22070 DVSS.n21665 0.00334
R64736 DVSS.n22070 DVSS.n22069 0.00334
R64737 DVSS.n22069 DVSS.n22068 0.00334
R64738 DVSS.n22068 DVSS.n21666 0.00334
R64739 DVSS.n22064 DVSS.n21666 0.00334
R64740 DVSS.n22064 DVSS.n22063 0.00334
R64741 DVSS.n22063 DVSS.n22062 0.00334
R64742 DVSS.n22062 DVSS.n21671 0.00334
R64743 DVSS.n22058 DVSS.n21671 0.00334
R64744 DVSS.n22058 DVSS.n22057 0.00334
R64745 DVSS.n22057 DVSS.n22056 0.00334
R64746 DVSS.n22056 DVSS.n21676 0.00334
R64747 DVSS.n22052 DVSS.n21676 0.00334
R64748 DVSS.n22052 DVSS.n22051 0.00334
R64749 DVSS.n22051 DVSS.n22050 0.00334
R64750 DVSS.n21748 DVSS.n21747 0.00334
R64751 DVSS.n21754 DVSS.n21747 0.00334
R64752 DVSS.n21755 DVSS.n21754 0.00334
R64753 DVSS.n22042 DVSS.n21755 0.00334
R64754 DVSS.n22042 DVSS.n22041 0.00334
R64755 DVSS.n22041 DVSS.n22040 0.00334
R64756 DVSS.n22040 DVSS.n21756 0.00334
R64757 DVSS.n22036 DVSS.n21756 0.00334
R64758 DVSS.n22036 DVSS.n22035 0.00334
R64759 DVSS.n22035 DVSS.n22034 0.00334
R64760 DVSS.n22034 DVSS.n21761 0.00334
R64761 DVSS.n22030 DVSS.n21761 0.00334
R64762 DVSS.n22030 DVSS.n22029 0.00334
R64763 DVSS.n22029 DVSS.n22028 0.00334
R64764 DVSS.n22028 DVSS.n21766 0.00334
R64765 DVSS.n22024 DVSS.n21766 0.00334
R64766 DVSS.n22024 DVSS.n22023 0.00334
R64767 DVSS.n22023 DVSS.n22022 0.00334
R64768 DVSS.n22022 DVSS.n21771 0.00334
R64769 DVSS.n22018 DVSS.n21771 0.00334
R64770 DVSS.n22018 DVSS.n22017 0.00334
R64771 DVSS.n22017 DVSS.n22016 0.00334
R64772 DVSS.n22016 DVSS.n21776 0.00334
R64773 DVSS.n22011 DVSS.n22010 0.00334
R64774 DVSS.n22010 DVSS.n22009 0.00334
R64775 DVSS.n22009 DVSS.n21971 0.00334
R64776 DVSS.n22005 DVSS.n21971 0.00334
R64777 DVSS.n22005 DVSS.n22004 0.00334
R64778 DVSS.n22004 DVSS.n22003 0.00334
R64779 DVSS.n22003 DVSS.n21976 0.00334
R64780 DVSS.n21999 DVSS.n21976 0.00334
R64781 DVSS.n21999 DVSS.n21998 0.00334
R64782 DVSS.n21998 DVSS.n21997 0.00334
R64783 DVSS.n21997 DVSS.n21982 0.00334
R64784 DVSS.n21993 DVSS.n21992 0.00334
R64785 DVSS.n13794 DVSS.n13793 0.00334
R64786 DVSS.n13795 DVSS.n13794 0.00334
R64787 DVSS.n13795 DVSS.n13784 0.00334
R64788 DVSS.n13802 DVSS.n13784 0.00334
R64789 DVSS.n13803 DVSS.n13802 0.00334
R64790 DVSS.n13804 DVSS.n13803 0.00334
R64791 DVSS.n13804 DVSS.n13781 0.00334
R64792 DVSS.n13811 DVSS.n13781 0.00334
R64793 DVSS.n13812 DVSS.n13811 0.00334
R64794 DVSS.n13813 DVSS.n13812 0.00334
R64795 DVSS.n13814 DVSS.n13813 0.00334
R64796 DVSS.n13815 DVSS.n13814 0.00334
R64797 DVSS.n13816 DVSS.n13815 0.00334
R64798 DVSS.n13819 DVSS.n13816 0.00334
R64799 DVSS.n13820 DVSS.n13819 0.00334
R64800 DVSS.n13821 DVSS.n13820 0.00334
R64801 DVSS.n13822 DVSS.n13821 0.00334
R64802 DVSS.n13897 DVSS.n13822 0.00334
R64803 DVSS.n13898 DVSS.n13897 0.00334
R64804 DVSS.n13903 DVSS.n13898 0.00334
R64805 DVSS.n13904 DVSS.n13903 0.00334
R64806 DVSS.n13905 DVSS.n13904 0.00334
R64807 DVSS.n13905 DVSS.n13894 0.00334
R64808 DVSS.n13912 DVSS.n13894 0.00334
R64809 DVSS.n13913 DVSS.n13912 0.00334
R64810 DVSS.n13914 DVSS.n13913 0.00334
R64811 DVSS.n13914 DVSS.n13891 0.00334
R64812 DVSS.n13921 DVSS.n13891 0.00334
R64813 DVSS.n13922 DVSS.n13921 0.00334
R64814 DVSS.n13923 DVSS.n13922 0.00334
R64815 DVSS.n13924 DVSS.n13923 0.00334
R64816 DVSS.n13925 DVSS.n13924 0.00334
R64817 DVSS.n13987 DVSS.n13925 0.00334
R64818 DVSS.n13988 DVSS.n13987 0.00334
R64819 DVSS.n13989 DVSS.n13988 0.00334
R64820 DVSS.n13989 DVSS.n13985 0.00334
R64821 DVSS.n13996 DVSS.n13985 0.00334
R64822 DVSS.n13997 DVSS.n13996 0.00334
R64823 DVSS.n13998 DVSS.n13997 0.00334
R64824 DVSS.n13998 DVSS.n13982 0.00334
R64825 DVSS.n14005 DVSS.n13982 0.00334
R64826 DVSS.n14006 DVSS.n14005 0.00334
R64827 DVSS.n14007 DVSS.n14006 0.00334
R64828 DVSS.n14008 DVSS.n14007 0.00334
R64829 DVSS.n14009 DVSS.n14008 0.00334
R64830 DVSS.n14010 DVSS.n14009 0.00334
R64831 DVSS.n14011 DVSS.n14010 0.00334
R64832 DVSS.n14012 DVSS.n14011 0.00334
R64833 DVSS.n14015 DVSS.n14012 0.00334
R64834 DVSS.n14016 DVSS.n14015 0.00334
R64835 DVSS.n14017 DVSS.n14016 0.00334
R64836 DVSS.n14018 DVSS.n14017 0.00334
R64837 DVSS.n14094 DVSS.n14018 0.00334
R64838 DVSS.n14095 DVSS.n14094 0.00334
R64839 DVSS.n14095 DVSS.n14093 0.00334
R64840 DVSS.n14102 DVSS.n14093 0.00334
R64841 DVSS.n14103 DVSS.n14102 0.00334
R64842 DVSS.n14104 DVSS.n14103 0.00334
R64843 DVSS.n14104 DVSS.n14090 0.00334
R64844 DVSS.n14111 DVSS.n14090 0.00334
R64845 DVSS.n14112 DVSS.n14111 0.00334
R64846 DVSS.n14113 DVSS.n14112 0.00334
R64847 DVSS.n14113 DVSS.n14087 0.00334
R64848 DVSS.n14120 DVSS.n14087 0.00334
R64849 DVSS.n14121 DVSS.n14120 0.00334
R64850 DVSS.n14122 DVSS.n14121 0.00334
R64851 DVSS.n14123 DVSS.n14122 0.00334
R64852 DVSS.n14124 DVSS.n14123 0.00334
R64853 DVSS.n14201 DVSS.n14124 0.00334
R64854 DVSS.n14202 DVSS.n14201 0.00334
R64855 DVSS.n14203 DVSS.n14202 0.00334
R64856 DVSS.n14203 DVSS.n14199 0.00334
R64857 DVSS.n14210 DVSS.n14199 0.00334
R64858 DVSS.n14211 DVSS.n14210 0.00334
R64859 DVSS.n14212 DVSS.n14211 0.00334
R64860 DVSS.n14212 DVSS.n14196 0.00334
R64861 DVSS.n14219 DVSS.n14196 0.00334
R64862 DVSS.n14220 DVSS.n14219 0.00334
R64863 DVSS.n14221 DVSS.n14220 0.00334
R64864 DVSS.n14221 DVSS.n14193 0.00334
R64865 DVSS.n14228 DVSS.n14193 0.00334
R64866 DVSS.n14229 DVSS.n14228 0.00334
R64867 DVSS.n14230 DVSS.n14229 0.00334
R64868 DVSS.n14231 DVSS.n14230 0.00334
R64869 DVSS.n14232 DVSS.n14231 0.00334
R64870 DVSS.n14235 DVSS.n14232 0.00334
R64871 DVSS.n14236 DVSS.n14235 0.00334
R64872 DVSS.n14237 DVSS.n14236 0.00334
R64873 DVSS.n14297 DVSS.n14237 0.00334
R64874 DVSS.n14298 DVSS.n14297 0.00334
R64875 DVSS.n14299 DVSS.n14298 0.00334
R64876 DVSS.n14300 DVSS.n14299 0.00334
R64877 DVSS.n14301 DVSS.n14300 0.00334
R64878 DVSS.n14302 DVSS.n14301 0.00334
R64879 DVSS.n14303 DVSS.n14302 0.00334
R64880 DVSS.n14304 DVSS.n14303 0.00334
R64881 DVSS.n14307 DVSS.n14306 0.00334
R64882 DVSS.n16651 DVSS.n16268 0.00332857
R64883 DVSS.n16082 DVSS.n16073 0.00332857
R64884 DVSS.n15291 DVSS.n15290 0.00332857
R64885 DVSS.n18461 DVSS.n14883 0.00332857
R64886 DVSS.n20819 DVSS.n14483 0.00332857
R64887 DVSS.n21269 DVSS.n13541 0.00332857
R64888 DVSS.n22727 DVSS.n624 0.00332857
R64889 DVSS.n21097 DVSS.n21096 0.00332
R64890 DVSS.n14222 DVSS.n14174 0.00332
R64891 DVSS.n21509 DVSS.n1486 0.00332
R64892 DVSS.n1123 DVSS.n1108 0.00332
R64893 DVSS.n334 DVSS.n331 0.00332
R64894 DVSS.n1485 DVSS.n780 0.00332
R64895 DVSS.n23092 DVSS.n239 0.00332
R64896 DVSS.n23173 DVSS.n23172 0.00332
R64897 DVSS.n1484 DVSS.n1435 0.00332
R64898 DVSS.n21662 DVSS.n21615 0.00332
R64899 DVSS.n21960 DVSS.n21818 0.00332
R64900 DVSS.n22113 DVSS.n779 0.00332
R64901 DVSS.n22547 DVSS.n22546 0.00332
R64902 DVSS.n21508 DVSS.n778 0.00332
R64903 DVSS.n17950 DVSS.n15738 0.0033169
R64904 DVSS.n18046 DVSS.n15703 0.0033169
R64905 DVSS.n16467 DVSS.n16466 0.00330976
R64906 DVSS.n18085 DVSS.n18084 0.00330976
R64907 DVSS.n22130 DVSS.n1379 0.00329474
R64908 DVSS.n964 DVSS.n915 0.00329474
R64909 DVSS.n22397 DVSS.n994 0.00329474
R64910 DVSS.n22278 DVSS.n1253 0.00329474
R64911 DVSS.n12859 DVSS.n25 0.00329474
R64912 DVSS.n12891 DVSS.n12803 0.00329474
R64913 DVSS.n21464 DVSS.n21450 0.0032907
R64914 DVSS.n22962 DVSS.n426 0.0032907
R64915 DVSS.n23217 DVSS.n23216 0.00329
R64916 DVSS.n21896 DVSS.n21595 0.00326585
R64917 DVSS.n837 DVSS.n223 0.00326585
R64918 DVSS.n21893 DVSS.n21698 0.00326585
R64919 DVSS.n834 DVSS.n143 0.00326585
R64920 DVSS.n21899 DVSS.n21898 0.00326585
R64921 DVSS.n840 DVSS.n839 0.00326585
R64922 DVSS.n21892 DVSS.n21791 0.00326585
R64923 DVSS.n833 DVSS.n78 0.00326585
R64924 DVSS.n16562 DVSS.n16350 0.00326429
R64925 DVSS.n15977 DVSS.n15945 0.00326429
R64926 DVSS.n17734 DVSS.n17678 0.00326429
R64927 DVSS.n15201 DVSS.n15173 0.00326429
R64928 DVSS.n20740 DVSS.n13710 0.00326429
R64929 DVSS.n13653 DVSS.n13638 0.00326429
R64930 DVSS.n22641 DVSS.n716 0.00326429
R64931 DVSS.n21993 DVSS 0.00326
R64932 DVSS.n14306 DVSS 0.00326
R64933 DVSS.n13917 DVSS.n13885 0.00326
R64934 DVSS.n14088 DVSS.n14080 0.00326
R64935 DVSS.n1473 DVSS.n1065 0.00326
R64936 DVSS.n12987 DVSS.n12986 0.00326
R64937 DVSS.n22500 DVSS.n22499 0.00326
R64938 DVSS.n191 DVSS.n172 0.00326
R64939 DVSS.n21868 DVSS.n1451 0.00326
R64940 DVSS.n22048 DVSS.n21682 0.00326
R64941 DVSS.n18012 DVSS.n15553 0.00324648
R64942 DVSS.n21051 DVSS.n14277 0.00323
R64943 DVSS.n12793 DVSS.n408 0.00323
R64944 DVSS.n23200 DVSS.n38 0.00323
R64945 DVSS.n21973 DVSS.n1237 0.00323
R64946 DVSS.n10120 DVSS.n10119 0.00320677
R64947 DVSS.n10456 DVSS.n1964 0.00320677
R64948 DVSS.n16667 DVSS.n16273 0.0032
R64949 DVSS.n16719 DVSS.n15664 0.0032
R64950 DVSS.n16128 DVSS.n16085 0.0032
R64951 DVSS.n17593 DVSS.n16904 0.0032
R64952 DVSS.n15343 DVSS.n15320 0.0032
R64953 DVSS.n18303 DVSS.n15447 0.0032
R64954 DVSS.n18445 DVSS.n14886 0.0032
R64955 DVSS.n15056 DVSS.n15028 0.0032
R64956 DVSS.n20835 DVSS.n14488 0.0032
R64957 DVSS.n14399 DVSS.n14388 0.0032
R64958 DVSS.n13901 DVSS.n13880 0.0032
R64959 DVSS.n14096 DVSS.n14075 0.0032
R64960 DVSS.n21285 DVSS.n13546 0.0032
R64961 DVSS.n13454 DVSS.n13447 0.0032
R64962 DVSS.n22223 DVSS.n704 0.0032
R64963 DVSS.n22153 DVSS.n1386 0.0032
R64964 DVSS.n932 DVSS.n904 0.0032
R64965 DVSS.n22427 DVSS.n1011 0.0032
R64966 DVSS.n22238 DVSS.n461 0.0032
R64967 DVSS.n22308 DVSS.n1260 0.0032
R64968 DVSS.n12827 DVSS.n14 0.0032
R64969 DVSS.n12921 DVSS.n12796 0.0032
R64970 DVSS.n22743 DVSS.n629 0.0032
R64971 DVSS.n22821 DVSS.n528 0.0032
R64972 DVSS.n21519 DVSS.n1061 0.0032
R64973 DVSS.n12981 DVSS.n300 0.0032
R64974 DVSS.n22485 DVSS.n790 0.0032
R64975 DVSS.n23111 DVSS.n167 0.0032
R64976 DVSS.n21861 DVSS.n1442 0.0032
R64977 DVSS.n21734 DVSS.n21673 0.0032
R64978 DVSS.n21896 DVSS.n21565 0.00317805
R64979 DVSS.n837 DVSS.n212 0.00317805
R64980 DVSS.n21893 DVSS.n21691 0.00317805
R64981 DVSS.n834 DVSS.n132 0.00317805
R64982 DVSS.n21898 DVSS.n21878 0.00317805
R64983 DVSS.n839 DVSS.n808 0.00317805
R64984 DVSS.n21892 DVSS.n21785 0.00317805
R64985 DVSS.n833 DVSS.n67 0.00317805
R64986 DVSS.n17851 DVSS.n15852 0.00317606
R64987 DVSS.n15774 DVSS.n15759 0.00317606
R64988 DVSS.n21117 DVSS.n21116 0.00314
R64989 DVSS.n21513 DVSS.n1060 0.00314
R64990 DVSS.n22483 DVSS.n786 0.00314
R64991 DVSS.n21860 DVSS.n21859 0.00314
R64992 DVSS.n21058 DVSS.n14234 0.00311
R64993 DVSS.n13099 DVSS.n12794 0.00311
R64994 DVSS.n12787 DVSS 0.00311
R64995 DVSS.n23191 DVSS.n35 0.00311
R64996 DVSS.n22325 DVSS.n1238 0.00311
R64997 DVSS.n22167 DVSS.n22127 0.00310526
R64998 DVSS.n22413 DVSS.n996 0.00310526
R64999 DVSS.n22294 DVSS.n1245 0.00310526
R65000 DVSS.n12907 DVSS.n12815 0.00310526
R65001 DVSS.n21028 DVSS.n14308 0.00309529
R65002 DVSS.n13790 DVSS.n13787 0.00309529
R65003 DVSS.n21991 DVSS.n21990 0.00309529
R65004 DVSS.n23224 DVSS.n23223 0.00309529
R65005 DVSS.n13910 DVSS.n13884 0.00308
R65006 DVSS.n14105 DVSS.n14079 0.00308
R65007 DVSS.n21527 DVSS.n1064 0.00308
R65008 DVSS.n12985 DVSS.n305 0.00308
R65009 DVSS.n22490 DVSS.n795 0.00308
R65010 DVSS.n23119 DVSS.n171 0.00308
R65011 DVSS.n21867 DVSS.n1447 0.00308
R65012 DVSS.n21739 DVSS.n21678 0.00308
R65013 DVSS.n16179 DVSS.n16165 0.00307143
R65014 DVSS.n18079 DVSS.n15668 0.00307143
R65015 DVSS.n16852 DVSS.n16832 0.00307143
R65016 DVSS.n17577 DVSS.n16907 0.00307143
R65017 DVSS.n15396 DVSS.n15377 0.00307143
R65018 DVSS.n18287 DVSS.n15450 0.00307143
R65019 DVSS.n14958 DVSS.n14944 0.00307143
R65020 DVSS.n19970 DVSS.n15033 0.00307143
R65021 DVSS.n20891 DVSS.n14410 0.00307143
R65022 DVSS.n20931 DVSS.n20930 0.00307143
R65023 DVSS.n21341 DVSS.n13465 0.00307143
R65024 DVSS.n21385 DVSS.n21384 0.00307143
R65025 DVSS.n22799 DVSS.n547 0.00307143
R65026 DVSS.n22839 DVSS.n496 0.00307143
R65027 DVSS.n21039 DVSS.n14261 0.00305
R65028 DVSS.n12789 DVSS.n413 0.00305
R65029 DVSS.n23208 DVSS.n42 0.00305
R65030 DVSS.n21979 DVSS.n1234 0.00305
R65031 DVSS.n20042 DVSS.n14464 0.00304634
R65032 DVSS.n20045 DVSS.n14465 0.00304634
R65033 DVSS.n20209 DVSS.n14415 0.00304634
R65034 DVSS.n20211 DVSS.n14416 0.00304634
R65035 DVSS.n18871 DVSS.n14511 0.00304634
R65036 DVSS.n18873 DVSS.n14512 0.00304634
R65037 DVSS.n14675 DVSS.n14366 0.00304634
R65038 DVSS.n14677 DVSS.n14367 0.00304634
R65039 DVSS.n17835 DVSS.n15856 0.00303521
R65040 DVSS.n18983 DVSS.n18982 0.00302809
R65041 DVSS.n20129 DVSS.n20053 0.00302809
R65042 DVSS.n20141 DVSS.n20051 0.00302809
R65043 DVSS.n20286 DVSS.n20224 0.00302809
R65044 DVSS.n20214 DVSS.n20208 0.00302809
R65045 DVSS.n20383 DVSS.n14685 0.00302809
R65046 DVSS.n21074 DVSS.n14084 0.00302
R65047 DVSS.n14190 DVSS.n14162 0.00302
R65048 DVSS.n13062 DVSS.n12990 0.00302
R65049 DVSS.n395 DVSS.n376 0.00302
R65050 DVSS.n23138 DVSS.n125 0.00302
R65051 DVSS.n94 DVSS.n60 0.00302
R65052 DVSS.n22045 DVSS.n21743 0.00302
R65053 DVSS.n21811 DVSS.n21774 0.00302
R65054 DVSS.n22169 DVSS.n22127 0.00301053
R65055 DVSS.n22411 DVSS.n996 0.00301053
R65056 DVSS.n22292 DVSS.n1245 0.00301053
R65057 DVSS.n12905 DVSS.n12815 0.00301053
R65058 DVSS.n16751 DVSS.n15596 0.00300714
R65059 DVSS.n18189 DVSS.n15494 0.00300714
R65060 DVSS.n18263 DVSS.n18220 0.00300714
R65061 DVSS.n19942 DVSS.n15104 0.00300714
R65062 DVSS.n20955 DVSS.n14339 0.00300714
R65063 DVSS.n21409 DVSS.n13396 0.00300714
R65064 DVSS.n22865 DVSS.n472 0.00300714
R65065 DVSS.n21142 DVSS.n13757 0.00299
R65066 DVSS.n21501 DVSS.n978 0.00299
R65067 DVSS.n888 DVSS.n776 0.00299
R65068 DVSS.n22184 DVSS.n22119 0.00299
R65069 DVSS.n14003 DVSS.n13943 0.00296
R65070 DVSS.n14213 DVSS.n14177 0.00296
R65071 DVSS.n1120 DVSS.n1111 0.00296
R65072 DVSS.n379 DVSS.n326 0.00296
R65073 DVSS.n268 DVSS.n241 0.00296
R65074 DVSS.n23157 DVSS.n97 0.00296
R65075 DVSS.n21654 DVSS.n21624 0.00296
R65076 DVSS.n21956 DVSS.n21821 0.00296
R65077 DVSS.n16625 DVSS.n16308 0.00294286
R65078 DVSS.n16705 DVSS.n16156 0.00294286
R65079 DVSS.n16052 DVSS.n16017 0.00294286
R65080 DVSS.n16870 DVSS.n16840 0.00294286
R65081 DVSS.n18369 DVSS.n15242 0.00294286
R65082 DVSS.n15414 DVSS.n15384 0.00294286
R65083 DVSS.n18419 DVSS.n18384 0.00294286
R65084 DVSS.n14976 DVSS.n14948 0.00294286
R65085 DVSS.n20791 DVSS.n20707 0.00294286
R65086 DVSS.n14448 DVSS.n14429 0.00294286
R65087 DVSS.n21243 DVSS.n13586 0.00294286
R65088 DVSS.n13505 DVSS.n13485 0.00294286
R65089 DVSS.n22701 DVSS.n675 0.00294286
R65090 DVSS.n585 DVSS.n569 0.00294286
R65091 DVSS.n13782 DVSS.n13740 0.00293
R65092 DVSS.n21486 DVSS.n984 0.00293
R65093 DVSS.n896 DVSS.n767 0.00293
R65094 DVSS.n1420 DVSS.n1374 0.00293
R65095 DVSS.n10117 DVSS.n2717 0.00291611
R65096 DVSS.n2021 DVSS.n1966 0.00291611
R65097 DVSS.n10118 DVSS.n2715 0.00291611
R65098 DVSS.n2023 DVSS.n1965 0.00291611
R65099 DVSS.n22225 DVSS.n704 0.00291579
R65100 DVSS.n22151 DVSS.n1386 0.00291579
R65101 DVSS.n934 DVSS.n904 0.00291579
R65102 DVSS.n22431 DVSS.n1011 0.00291579
R65103 DVSS.n22236 DVSS.n461 0.00291579
R65104 DVSS.n22310 DVSS.n1260 0.00291579
R65105 DVSS.n12829 DVSS.n14 0.00291579
R65106 DVSS.n12819 DVSS.n12796 0.00291579
R65107 DVSS.n21886 DVSS.n21593 0.00291463
R65108 DVSS.n828 DVSS.n221 0.00291463
R65109 DVSS.n13042 DVSS.n1151 0.00291463
R65110 DVSS.n21884 DVSS.n21696 0.00291463
R65111 DVSS.n825 DVSS.n141 0.00291463
R65112 DVSS.n13047 DVSS.n13046 0.00291463
R65113 DVSS.n21889 DVSS.n21888 0.00291463
R65114 DVSS.n831 DVSS.n830 0.00291463
R65115 DVSS.n13041 DVSS.n1096 0.00291463
R65116 DVSS.n21883 DVSS.n21789 0.00291463
R65117 DVSS.n824 DVSS.n76 0.00291463
R65118 DVSS.n13040 DVSS.n364 0.00291463
R65119 DVSS.n21107 DVSS.n13939 0.0029
R65120 DVSS.n21547 DVSS.n1115 0.0029
R65121 DVSS.n22511 DVSS.n245 0.0029
R65122 DVSS.n21628 DVSS.n1460 0.0029
R65123 DVSS.n17842 DVSS.n15854 0.00289437
R65124 DVSS.n15777 DVSS.n15761 0.00289437
R65125 DVSS.n13798 DVSS.n13733 0.00287
R65126 DVSS.n1498 DVSS.n974 0.00287
R65127 DVSS.n897 DVSS.n884 0.00287
R65128 DVSS.n1401 DVSS.n1367 0.00287
R65129 DVSS.n22993 DVSS.n401 0.00286
R65130 DVSS.n23194 DVSS.n52 0.00286
R65131 DVSS.n22011 DVSS.n21970 0.00286
R65132 DVSS.n13737 DVSS.n13735 0.00285923
R65133 DVSS.n13742 DVSS.n13731 0.00285923
R65134 DVSS.n13881 DVSS.n13876 0.00285923
R65135 DVSS.n13886 DVSS.n13861 0.00285923
R65136 DVSS.n13978 DVSS.n13945 0.00285923
R65137 DVSS.n13977 DVSS.n13941 0.00285923
R65138 DVSS.n14076 DVSS.n14072 0.00285923
R65139 DVSS.n14081 DVSS.n14068 0.00285923
R65140 DVSS.n14181 DVSS.n14179 0.00285923
R65141 DVSS.n14186 DVSS.n14175 0.00285923
R65142 DVSS.n14274 DVSS.n14253 0.00285923
R65143 DVSS.n14275 DVSS.n14257 0.00285923
R65144 DVSS.n13979 DVSS.n13945 0.00285923
R65145 DVSS.n21103 DVSS.n13941 0.00285923
R65146 DVSS.n14077 DVSS.n14076 0.00285923
R65147 DVSS.n14082 DVSS.n14081 0.00285923
R65148 DVSS.n13882 DVSS.n13881 0.00285923
R65149 DVSS.n13887 DVSS.n13886 0.00285923
R65150 DVSS.n13738 DVSS.n13737 0.00285923
R65151 DVSS.n13743 DVSS.n13742 0.00285923
R65152 DVSS.n14182 DVSS.n14181 0.00285923
R65153 DVSS.n14187 DVSS.n14186 0.00285923
R65154 DVSS.n14275 DVSS.n14259 0.00285923
R65155 DVSS.n14274 DVSS.n14263 0.00285923
R65156 DVSS.n999 DVSS.n972 0.00285923
R65157 DVSS.n998 DVSS.n976 0.00285923
R65158 DVSS.n1081 DVSS.n1056 0.00285923
R65159 DVSS.n1106 DVSS.n1100 0.00285923
R65160 DVSS.n1135 DVSS.n1113 0.00285923
R65161 DVSS.n1164 DVSS.n1154 0.00285923
R65162 DVSS.n13005 DVSS.n12977 0.00285923
R65163 DVSS.n13004 DVSS.n12973 0.00285923
R65164 DVSS.n385 DVSS.n381 0.00285923
R65165 DVSS.n392 DVSS.n377 0.00285923
R65166 DVSS.n12806 DVSS.n12779 0.00285923
R65167 DVSS.n12807 DVSS.n12783 0.00285923
R65168 DVSS.n12807 DVSS.n12786 0.00285923
R65169 DVSS.n12806 DVSS.n12792 0.00285923
R65170 DVSS.n999 DVSS.n986 0.00285923
R65171 DVSS.n998 DVSS.n982 0.00285923
R65172 DVSS.n1081 DVSS.n1062 0.00285923
R65173 DVSS.n1100 DVSS.n1066 0.00285923
R65174 DVSS.n1135 DVSS.n1117 0.00285923
R65175 DVSS.n1154 DVSS.n1122 0.00285923
R65176 DVSS.n13005 DVSS.n12982 0.00285923
R65177 DVSS.n13004 DVSS.n12988 0.00285923
R65178 DVSS.n386 DVSS.n385 0.00285923
R65179 DVSS.n393 DVSS.n392 0.00285923
R65180 DVSS.n912 DVSS.n882 0.00285923
R65181 DVSS.n911 DVSS.n886 0.00285923
R65182 DVSS.n22486 DVSS.n22475 0.00285923
R65183 DVSS.n22501 DVSS.n22472 0.00285923
R65184 DVSS.n248 DVSS.n243 0.00285923
R65185 DVSS.n262 DVSS.n254 0.00285923
R65186 DVSS.n168 DVSS.n163 0.00285923
R65187 DVSS.n182 DVSS.n174 0.00285923
R65188 DVSS.n102 DVSS.n99 0.00285923
R65189 DVSS.n107 DVSS.n95 0.00285923
R65190 DVSS.n39 DVSS.n33 0.00285923
R65191 DVSS.n23218 DVSS.n29 0.00285923
R65192 DVSS.n23219 DVSS.n23218 0.00285923
R65193 DVSS.n40 DVSS.n39 0.00285923
R65194 DVSS.n912 DVSS.n899 0.00285923
R65195 DVSS.n911 DVSS.n893 0.00285923
R65196 DVSS.n22487 DVSS.n22486 0.00285923
R65197 DVSS.n22502 DVSS.n22501 0.00285923
R65198 DVSS.n249 DVSS.n248 0.00285923
R65199 DVSS.n254 DVSS.n253 0.00285923
R65200 DVSS.n169 DVSS.n168 0.00285923
R65201 DVSS.n174 DVSS.n173 0.00285923
R65202 DVSS.n103 DVSS.n102 0.00285923
R65203 DVSS.n108 DVSS.n107 0.00285923
R65204 DVSS.n1390 DVSS.n1369 0.00285923
R65205 DVSS.n1389 DVSS.n1365 0.00285923
R65206 DVSS.n21863 DVSS.n21855 0.00285923
R65207 DVSS.n21932 DVSS.n21922 0.00285923
R65208 DVSS.n21631 DVSS.n1463 0.00285923
R65209 DVSS.n21635 DVSS.n21622 0.00285923
R65210 DVSS.n21735 DVSS.n21729 0.00285923
R65211 DVSS.n21740 DVSS.n21725 0.00285923
R65212 DVSS.n21951 DVSS.n21823 0.00285923
R65213 DVSS.n21958 DVSS.n21819 0.00285923
R65214 DVSS.n1250 DVSS.n1226 0.00285923
R65215 DVSS.n1249 DVSS.n1230 0.00285923
R65216 DVSS.n1250 DVSS.n1236 0.00285923
R65217 DVSS.n1249 DVSS.n1232 0.00285923
R65218 DVSS.n1390 DVSS.n1372 0.00285923
R65219 DVSS.n1389 DVSS.n1376 0.00285923
R65220 DVSS.n21864 DVSS.n21863 0.00285923
R65221 DVSS.n21922 DVSS.n21869 0.00285923
R65222 DVSS.n21632 DVSS.n21631 0.00285923
R65223 DVSS.n21636 DVSS.n21635 0.00285923
R65224 DVSS.n21736 DVSS.n21735 0.00285923
R65225 DVSS.n21741 DVSS.n21740 0.00285923
R65226 DVSS.n21952 DVSS.n21951 0.00285923
R65227 DVSS.n21959 DVSS.n21958 0.00285923
R65228 DVSS.n21465 DVSS.n21448 0.00284375
R65229 DVSS.n22963 DVSS.n424 0.00284375
R65230 DVSS.n13999 DVSS.n13950 0.00284
R65231 DVSS.n14208 DVSS.n14184 0.00284
R65232 DVSS.n13677 DVSS.n13673 0.00284
R65233 DVSS.n21162 DVSS.n13675 0.00284
R65234 DVSS.n21157 DVSS.n21156 0.00284
R65235 DVSS.n13685 DVSS.n13684 0.00284
R65236 DVSS.n18510 DVSS.n18509 0.00284
R65237 DVSS.n1119 DVSS.n280 0.00284
R65238 DVSS.n389 DVSS.n388 0.00284
R65239 DVSS.n23078 DVSS.n251 0.00284
R65240 DVSS.n119 DVSS.n105 0.00284
R65241 DVSS.n21648 DVSS.n21633 0.00284
R65242 DVSS.n21955 DVSS.n21763 0.00284
R65243 DVSS.n21906 DVSS.n21563 0.00282683
R65244 DVSS.n846 DVSS.n210 0.00282683
R65245 DVSS.n21903 DVSS.n21689 0.00282683
R65246 DVSS.n843 DVSS.n130 0.00282683
R65247 DVSS.n21908 DVSS.n21876 0.00282683
R65248 DVSS.n848 DVSS.n806 0.00282683
R65249 DVSS.n21902 DVSS.n21783 0.00282683
R65250 DVSS.n842 DVSS.n65 0.00282683
R65251 DVSS.n18020 DVSS.n15551 0.00282394
R65252 DVSS.n1379 DVSS.n1370 0.00282105
R65253 DVSS.n962 DVSS.n915 0.00282105
R65254 DVSS.n22395 DVSS.n994 0.00282105
R65255 DVSS.n22276 DVSS.n1253 0.00282105
R65256 DVSS.n12857 DVSS.n25 0.00282105
R65257 DVSS.n12889 DVSS.n12803 0.00282105
R65258 DVSS.n22975 DVSS 0.00282
R65259 DVSS.n16609 DVSS.n16312 0.00281429
R65260 DVSS.n17656 DVSS.n15993 0.00281429
R65261 DVSS.n17754 DVSS.n15246 0.00281429
R65262 DVSS.n15227 DVSS.n15223 0.00281429
R65263 DVSS.n20775 DVSS.n20711 0.00281429
R65264 DVSS.n21227 DVSS.n13593 0.00281429
R65265 DVSS.n22685 DVSS.n679 0.00281429
R65266 DVSS.n21139 DVSS.n21128 0.00281
R65267 DVSS.n1488 DVSS.n980 0.00281
R65268 DVSS.n891 DVSS.n773 0.00281
R65269 DVSS.n1430 DVSS.n1363 0.00281
R65270 DVSS DVSS.n14304 0.00278
R65271 DVSS.n21105 DVSS.n13953 0.00278
R65272 DVSS.n14224 DVSS.n14189 0.00278
R65273 DVSS.n22373 DVSS.n289 0.00278
R65274 DVSS.n23005 DVSS.n23004 0.00278
R65275 DVSS.n23095 DVSS.n205 0.00278
R65276 DVSS.n23180 DVSS.n110 0.00278
R65277 DVSS.n22073 DVSS.n21638 0.00278
R65278 DVSS.n21962 DVSS.n21772 0.00278
R65279 DVSS.n20680 DVSS.n14579 0.00277528
R65280 DVSS.n20143 DVSS 0.00277528
R65281 DVSS.n17859 DVSS.n15850 0.00275352
R65282 DVSS.n17939 DVSS.n15757 0.00275352
R65283 DVSS.n21035 DVSS.n14255 0.00275
R65284 DVSS.n12781 DVSS.n416 0.00275
R65285 DVSS.n23215 DVSS.n31 0.00275
R65286 DVSS.n21983 DVSS.n1228 0.00275
R65287 DVSS.n15306 DVSS.n15292 0.00273902
R65288 DVSS.n607 DVSS.n597 0.00273902
R65289 DVSS.n15373 DVSS.n15363 0.00273902
R65290 DVSS.n562 DVSS.n548 0.00273902
R65291 DVSS.n15267 DVSS.n15254 0.00273902
R65292 DVSS.n669 DVSS.n649 0.00273902
R65293 DVSS.n15443 DVSS.n15433 0.00273902
R65294 DVSS.n507 DVSS.n497 0.00273902
R65295 DVSS.n22135 DVSS.n22120 0.00272632
R65296 DVSS.n950 DVSS.n902 0.00272632
R65297 DVSS.n22437 DVSS.n970 0.00272632
R65298 DVSS.n22327 DVSS.n22326 0.00272632
R65299 DVSS.n12845 DVSS.n22 0.00272632
R65300 DVSS.n12877 DVSS.n12808 0.00272632
R65301 DVSS.n13915 DVSS.n13874 0.00272
R65302 DVSS.n14109 DVSS.n14070 0.00272
R65303 DVSS.n1471 DVSS.n1054 0.00272
R65304 DVSS.n21555 DVSS.n1118 0.00272
R65305 DVSS.n12975 DVSS.n307 0.00272
R65306 DVSS.n22473 DVSS.n797 0.00272
R65307 DVSS.n21556 DVSS.n250 0.00272
R65308 DVSS.n189 DVSS.n161 0.00272
R65309 DVSS.n21853 DVSS.n1450 0.00272
R65310 DVSS.n22076 DVSS.n22075 0.00272
R65311 DVSS.n21727 DVSS.n21726 0.00272
R65312 DVSS.n23034 DVSS.n23033 0.0027
R65313 DVSS.n23130 DVSS.n186 0.0027
R65314 DVSS.n21748 DVSS.n21681 0.0027
R65315 DVSS.n21054 DVSS.n14239 0.00269
R65316 DVSS.n12777 DVSS.n407 0.00269
R65317 DVSS.n23198 DVSS.n37 0.00269
R65318 DVSS.n21972 DVSS.n1224 0.00269
R65319 DVSS.n16616 DVSS.n16310 0.00268571
R65320 DVSS.n16696 DVSS.n16158 0.00268571
R65321 DVSS.n16043 DVSS.n16019 0.00268571
R65322 DVSS.n16842 DVSS.n16147 0.00268571
R65323 DVSS.n15274 DVSS.n15244 0.00268571
R65324 DVSS.n15386 DVSS.n15368 0.00268571
R65325 DVSS.n18410 DVSS.n18386 0.00268571
R65326 DVSS.n14950 DVSS.n14933 0.00268571
R65327 DVSS.n20782 DVSS.n20709 0.00268571
R65328 DVSS.n14451 DVSS.n14431 0.00268571
R65329 DVSS.n21234 DVSS.n13591 0.00268571
R65330 DVSS.n13508 DVSS.n13487 0.00268571
R65331 DVSS.n22692 DVSS.n677 0.00268571
R65332 DVSS.n588 DVSS.n571 0.00268571
R65333 DVSS.n18006 DVSS.n15549 0.0026831
R65334 DVSS.n8116 DVSS.n8115 0.00266541
R65335 DVSS.n13899 DVSS.n13878 0.00266
R65336 DVSS.n21076 DVSS.n14032 0.00266
R65337 DVSS.n1481 DVSS.n1058 0.00266
R65338 DVSS.n12980 DVSS.n12979 0.00266
R65339 DVSS.n22484 DVSS.n22477 0.00266
R65340 DVSS.n198 DVSS.n165 0.00266
R65341 DVSS.n21857 DVSS.n1441 0.00266
R65342 DVSS.n21732 DVSS.n21672 0.00266
R65343 DVSS.n12348 DVSS.n12344 0.0026375
R65344 DVSS.n12752 DVSS.n12751 0.0026375
R65345 DVSS.n6243 DVSS.n6241 0.0026375
R65346 DVSS.n6659 DVSS.n6240 0.0026375
R65347 DVSS.n22139 DVSS.n1391 0.00263158
R65348 DVSS.n946 DVSS.n917 0.00263158
R65349 DVSS.n22324 DVSS.n22323 0.00263158
R65350 DVSS.n12841 DVSS.n11 0.00263158
R65351 DVSS.n16760 DVSS.n15594 0.00262143
R65352 DVSS.n18201 DVSS.n15522 0.00262143
R65353 DVSS.n18273 DVSS.n18237 0.00262143
R65354 DVSS.n15118 DVSS.n15091 0.00262143
R65355 DVSS.n20969 DVSS.n20968 0.00262143
R65356 DVSS.n21423 DVSS.n21422 0.00262143
R65357 DVSS.n22856 DVSS.n474 0.00262143
R65358 DVSS.n17906 DVSS.n17905 0.00261268
R65359 DVSS.n18038 DVSS.n15701 0.00261268
R65360 DVSS.n13878 DVSS.n13837 0.0026
R65361 DVSS.n21077 DVSS.n21076 0.0026
R65362 DVSS.n1479 DVSS.n1058 0.0026
R65363 DVSS.n12979 DVSS.n297 0.0026
R65364 DVSS.n22477 DVSS.n787 0.0026
R65365 DVSS.n23104 DVSS.n165 0.0026
R65366 DVSS.n21857 DVSS.n1440 0.0026
R65367 DVSS.n21732 DVSS.n21731 0.0026
R65368 DVSS.n21055 DVSS.n21054 0.00257
R65369 DVSS.n12777 DVSS.n406 0.00257
R65370 DVSS.n51 DVSS.n37 0.00257
R65371 DVSS.n1252 DVSS.n1224 0.00257
R65372 DVSS.n819 DVSS.n206 0.00256341
R65373 DVSS.n13030 DVSS.n1127 0.00256341
R65374 DVSS.n816 DVSS.n126 0.00256341
R65375 DVSS.n13034 DVSS.n12992 0.00256341
R65376 DVSS.n821 DVSS.n802 0.00256341
R65377 DVSS.n13029 DVSS.n1069 0.00256341
R65378 DVSS.n815 DVSS.n61 0.00256341
R65379 DVSS.n13028 DVSS.n337 0.00256341
R65380 DVSS.n16633 DVSS.n16306 0.00255714
R65381 DVSS.n16225 DVSS.n16154 0.00255714
R65382 DVSS.n16059 DVSS.n16015 0.00255714
R65383 DVSS.n16857 DVSS.n16838 0.00255714
R65384 DVSS.n18362 DVSS.n15240 0.00255714
R65385 DVSS.n15401 DVSS.n15382 0.00255714
R65386 DVSS.n18432 DVSS.n18427 0.00255714
R65387 DVSS.n14963 DVSS.n14946 0.00255714
R65388 DVSS.n20723 DVSS.n20722 0.00255714
R65389 DVSS.n20880 DVSS.n14427 0.00255714
R65390 DVSS.n21251 DVSS.n13584 0.00255714
R65391 DVSS.n21330 DVSS.n13483 0.00255714
R65392 DVSS.n22709 DVSS.n673 0.00255714
R65393 DVSS.n22788 DVSS.n567 0.00255714
R65394 DVSS.n15908 DVSS.n15893 0.00254225
R65395 DVSS.n23071 DVSS.n23070 0.00254
R65396 DVSS.n23072 DVSS.n269 0.00254
R65397 DVSS.n21649 DVSS.n276 0.00254
R65398 DVSS.n13892 DVSS.n13874 0.00254
R65399 DVSS.n14107 DVSS.n14070 0.00254
R65400 DVSS.n21529 DVSS.n1054 0.00254
R65401 DVSS.n12975 DVSS.n306 0.00254
R65402 DVSS.n22473 DVSS.n796 0.00254
R65403 DVSS.n23121 DVSS.n161 0.00254
R65404 DVSS.n21866 DVSS.n21853 0.00254
R65405 DVSS.n21727 DVSS.n21679 0.00254
R65406 DVSS.n16541 DVSS.n16343 0.00253684
R65407 DVSS.n22183 DVSS.n22182 0.00253684
R65408 DVSS.n966 DVSS.n923 0.00253684
R65409 DVSS.n22399 DVSS.n1008 0.00253684
R65410 DVSS.n18107 DVSS.n15611 0.00253684
R65411 DVSS.n22280 DVSS.n1248 0.00253684
R65412 DVSS.n12861 DVSS.n7 0.00253684
R65413 DVSS.n12893 DVSS.n12812 0.00253684
R65414 DVSS.n7831 DVSS.n7830 0.002525
R65415 DVSS.n18883 DVSS.n18881 0.00252247
R65416 DVSS.n20438 DVSS.n14692 0.00252247
R65417 DVSS.n21037 DVSS.n14255 0.00251
R65418 DVSS.n12788 DVSS.n12781 0.00251
R65419 DVSS.n43 DVSS.n31 0.00251
R65420 DVSS.n21980 DVSS.n1228 0.00251
R65421 DVSS.n16744 DVSS.n15592 0.00249286
R65422 DVSS.n18182 DVSS.n15496 0.00249286
R65423 DVSS.n18256 DVSS.n18222 0.00249286
R65424 DVSS.n19935 DVSS.n15106 0.00249286
R65425 DVSS.n20947 DVSS.n14341 0.00249286
R65426 DVSS.n21401 DVSS.n13398 0.00249286
R65427 DVSS.n22873 DVSS.n470 0.00249286
R65428 DVSS.n21105 DVSS.n13965 0.00248
R65429 DVSS.n14226 DVSS.n14189 0.00248
R65430 DVSS.n22373 DVSS.n290 0.00248
R65431 DVSS.n23004 DVSS.n350 0.00248
R65432 DVSS.n23096 DVSS.n23095 0.00248
R65433 DVSS.n23180 DVSS.n23179 0.00248
R65434 DVSS.n22073 DVSS.n22072 0.00248
R65435 DVSS.n21962 DVSS.n21773 0.00248
R65436 DVSS.n21916 DVSS.n21561 0.00247561
R65437 DVSS.n854 DVSS.n208 0.00247561
R65438 DVSS.n21913 DVSS.n21687 0.00247561
R65439 DVSS.n852 DVSS.n128 0.00247561
R65440 DVSS.n21918 DVSS.n21874 0.00247561
R65441 DVSS.n856 DVSS.n804 0.00247561
R65442 DVSS.n21912 DVSS.n21781 0.00247561
R65443 DVSS.n851 DVSS.n63 0.00247561
R65444 DVSS DVSS.n18007 0.00247183
R65445 DVSS.n17886 DVSS.n15816 0.00247183
R65446 DVSS.n15729 DVSS.n15698 0.00247183
R65447 DVSS.n18006 DVSS 0.00247183
R65448 DVSS.n21139 DVSS.n13745 0.00245
R65449 DVSS DVSS.n14260 0.00245
R65450 DVSS.n1490 DVSS.n980 0.00245
R65451 DVSS.n891 DVSS.n890 0.00245
R65452 DVSS.n1378 DVSS.n1363 0.00245
R65453 DVSS DVSS.n1233 0.00245
R65454 DVSS.n22221 DVSS.n709 0.00244211
R65455 DVSS.n22155 DVSS.n22124 0.00244211
R65456 DVSS.n930 DVSS.n906 0.00244211
R65457 DVSS.n22425 DVSS.n1002 0.00244211
R65458 DVSS.n22240 DVSS.n467 0.00244211
R65459 DVSS.n22306 DVSS.n1242 0.00244211
R65460 DVSS.n12825 DVSS.n18 0.00244211
R65461 DVSS.n12919 DVSS.n12818 0.00244211
R65462 DVSS.n8113 DVSS.n4013 0.00243289
R65463 DVSS.n8114 DVSS.n4016 0.00243289
R65464 DVSS.n16679 DVSS.n16678 0.00242857
R65465 DVSS.n16722 DVSS.n15666 0.00242857
R65466 DVSS.n17633 DVSS.n16086 0.00242857
R65467 DVSS.n17584 DVSS.n16906 0.00242857
R65468 DVSS.n15352 DVSS.n15323 0.00242857
R65469 DVSS.n18294 DVSS.n15449 0.00242857
R65470 DVSS.n19999 DVSS.n14887 0.00242857
R65471 DVSS.n15066 DVSS.n15031 0.00242857
R65472 DVSS.n20847 DVSS.n20846 0.00242857
R65473 DVSS.n14396 DVSS.n14391 0.00242857
R65474 DVSS.n21297 DVSS.n21296 0.00242857
R65475 DVSS.n13451 DVSS.n13450 0.00242857
R65476 DVSS.n22755 DVSS.n22754 0.00242857
R65477 DVSS.n22830 DVSS.n531 0.00242857
R65478 DVSS.n14001 DVSS.n13950 0.00242
R65479 DVSS.n14197 DVSS.n14184 0.00242
R65480 DVSS.n1119 DVSS.n281 0.00242
R65481 DVSS.n389 DVSS.n325 0.00242
R65482 DVSS.n266 DVSS.n251 0.00242
R65483 DVSS.n23155 DVSS.n105 0.00242
R65484 DVSS.n21652 DVSS.n21633 0.00242
R65485 DVSS.n21955 DVSS.n21764 0.00242
R65486 DVSS.n17794 DVSS.n15900 0.00240141
R65487 DVSS.n17801 DVSS.n15897 0.00240141
R65488 DVSS.n16494 DVSS.n15881 0.00239474
R65489 DVSS.n16496 DVSS.n15885 0.00239474
R65490 DVSS.n16498 DVSS.n15882 0.00239474
R65491 DVSS.n16500 DVSS.n15884 0.00239474
R65492 DVSS.n16502 DVSS.n15883 0.00239474
R65493 DVSS.n18153 DVSS.n18152 0.00239474
R65494 DVSS.n15566 DVSS.n15555 0.00239474
R65495 DVSS.n15577 DVSS.n15574 0.00239474
R65496 DVSS.n15579 DVSS.n15565 0.00239474
R65497 DVSS.n18148 DVSS.n15575 0.00239474
R65498 DVSS.n13800 DVSS.n13733 0.00239
R65499 DVSS.n21484 DVSS.n974 0.00239
R65500 DVSS.n884 DVSS.n766 0.00239
R65501 DVSS.n1403 DVSS.n1367 0.00239
R65502 DVSS.n16426 DVSS.n16250 0.0023878
R65503 DVSS.n16220 DVSS.n16175 0.0023878
R65504 DVSS.n16467 DVSS.n16295 0.0023878
R65505 DVSS.n18085 DVSS.n15646 0.0023878
R65506 DVSS.n21507 DVSS.n21505 0.00238
R65507 DVSS.n22545 DVSS.n782 0.00238
R65508 DVSS.n22115 DVSS.n22114 0.00238
R65509 DVSS.n16559 DVSS.n16348 0.00236429
R65510 DVSS.n17673 DVSS.n17672 0.00236429
R65511 DVSS.n17771 DVSS.n17770 0.00236429
R65512 DVSS.n15215 DVSS.n15214 0.00236429
R65513 DVSS.n20737 DVSS.n13727 0.00236429
R65514 DVSS.n21205 DVSS.n13650 0.00236429
R65515 DVSS.n22644 DVSS.n718 0.00236429
R65516 DVSS.n21108 DVSS.n21107 0.00236
R65517 DVSS.n21545 DVSS.n1115 0.00236
R65518 DVSS.n22510 DVSS.n245 0.00236
R65519 DVSS.n21628 DVSS.n21627 0.00236
R65520 DVSS.n22165 DVSS.n1383 0.00234737
R65521 DVSS.n22415 DVSS.n990 0.00234737
R65522 DVSS.n22296 DVSS.n1257 0.00234737
R65523 DVSS.n12909 DVSS.n12799 0.00234737
R65524 DVSS.n17879 DVSS.n15806 0.00233099
R65525 DVSS.n17959 DVSS.n15697 0.00233099
R65526 DVSS.n13800 DVSS.n13740 0.00233
R65527 DVSS.n21484 DVSS.n984 0.00233
R65528 DVSS.n896 DVSS.n766 0.00233
R65529 DVSS.n1403 DVSS.n1374 0.00233
R65530 DVSS.n22872 DVSS 0.0023
R65531 DVSS DVSS.n16745 0.0023
R65532 DVSS.n16660 DVSS.n16271 0.0023
R65533 DVSS.n16798 DVSS.n15662 0.0023
R65534 DVSS.n16744 DVSS 0.0023
R65535 DVSS.n18183 DVSS 0.0023
R65536 DVSS.n16109 DVSS.n16083 0.0023
R65537 DVSS.n17548 DVSS.n16902 0.0023
R65538 DVSS.n18182 DVSS 0.0023
R65539 DVSS DVSS.n18257 0.0023
R65540 DVSS.n15332 DVSS.n15318 0.0023
R65541 DVSS.n15468 DVSS.n15445 0.0023
R65542 DVSS.n18256 DVSS 0.0023
R65543 DVSS.n19936 DVSS 0.0023
R65544 DVSS.n18452 DVSS.n14884 0.0023
R65545 DVSS.n15049 DVSS.n15026 0.0023
R65546 DVSS.n19935 DVSS 0.0023
R65547 DVSS.n20948 DVSS 0.0023
R65548 DVSS.n20828 DVSS.n14486 0.0023
R65549 DVSS.n20907 DVSS.n14386 0.0023
R65550 DVSS.n20947 DVSS 0.0023
R65551 DVSS.n14001 DVSS.n13943 0.0023
R65552 DVSS.n14197 DVSS.n14177 0.0023
R65553 DVSS.n21402 DVSS 0.0023
R65554 DVSS.n21278 DVSS.n13544 0.0023
R65555 DVSS.n21357 DVSS.n13445 0.0023
R65556 DVSS.n21401 DVSS 0.0023
R65557 DVSS.n17099 DVSS.n16088 0.0023
R65558 DVSS.n16827 DVSS.n16142 0.0023
R65559 DVSS.n16005 DVSS.n15994 0.0023
R65560 DVSS.n16900 DVSS.n16889 0.0023
R65561 DVSS.n22736 DVSS.n627 0.0023
R65562 DVSS.n538 DVSS.n526 0.0023
R65563 DVSS DVSS.n22873 0.0023
R65564 DVSS.n18519 DVSS.n15145 0.0023
R65565 DVSS.n17788 DVSS.n15920 0.0023
R65566 DVSS.n18170 DVSS.n15533 0.0023
R65567 DVSS.n19923 DVSS.n15137 0.0023
R65568 DVSS.n1111 DVSS.n281 0.0023
R65569 DVSS.n379 DVSS.n325 0.0023
R65570 DVSS.n266 DVSS.n241 0.0023
R65571 DVSS.n23155 DVSS.n97 0.0023
R65572 DVSS.n21652 DVSS.n21624 0.0023
R65573 DVSS.n21821 DVSS.n21764 0.0023
R65574 DVSS.n21142 DVSS.n13745 0.00227
R65575 DVSS.n1490 DVSS.n978 0.00227
R65576 DVSS.n890 DVSS.n888 0.00227
R65577 DVSS.n22184 DVSS.n1378 0.00227
R65578 DVSS.n18910 DVSS.n18909 0.00226966
R65579 DVSS.n20348 DVSS.n14681 0.00226966
R65580 DVSS.n7828 DVSS.n4467 0.00226856
R65581 DVSS.n7829 DVSS.n4465 0.00226856
R65582 DVSS.n17810 DVSS.n15905 0.00226056
R65583 DVSS.n20158 DVSS.n13927 0.0022561
R65584 DVSS.n20043 DVSS.n13954 0.0022561
R65585 DVSS.n21075 DVSS.n14044 0.0022561
R65586 DVSS.n14074 DVSS.n14020 0.0022561
R65587 DVSS.n16383 DVSS.n15839 0.0022561
R65588 DVSS.n16384 DVSS.n15843 0.0022561
R65589 DVSS.n16386 DVSS.n15840 0.0022561
R65590 DVSS.n16388 DVSS.n15842 0.0022561
R65591 DVSS.n16390 DVSS.n15841 0.0022561
R65592 DVSS.n21115 DVSS.n13849 0.0022561
R65593 DVSS.n13879 DVSS.n13825 0.0022561
R65594 DVSS.n15718 DVSS.n15706 0.0022561
R65595 DVSS.n15716 DVSS.n15710 0.0022561
R65596 DVSS.n15714 DVSS.n15707 0.0022561
R65597 DVSS.n15712 DVSS.n15709 0.0022561
R65598 DVSS.n18047 DVSS.n15689 0.0022561
R65599 DVSS.n21066 DVSS.n14150 0.0022561
R65600 DVSS.n14180 DVSS.n14126 0.0022561
R65601 DVSS.n22171 DVSS.n1382 0.00225263
R65602 DVSS.n22444 DVSS.n913 0.00225263
R65603 DVSS.n22409 DVSS.n1004 0.00225263
R65604 DVSS.n22290 DVSS.n1256 0.00225263
R65605 DVSS.n23220 DVSS.n28 0.00225263
R65606 DVSS.n12903 DVSS.n12800 0.00225263
R65607 DVSS.n21074 DVSS.n21073 0.00224
R65608 DVSS.n14226 DVSS.n14162 0.00224
R65609 DVSS.n13062 DVSS.n315 0.00224
R65610 DVSS.n376 DVSS.n350 0.00224
R65611 DVSS.n23139 DVSS.n23138 0.00224
R65612 DVSS.n23179 DVSS.n94 0.00224
R65613 DVSS.n22045 DVSS.n22044 0.00224
R65614 DVSS.n21811 DVSS.n21773 0.00224
R65615 DVSS.n16568 DVSS.n16551 0.00223571
R65616 DVSS.n16575 DVSS.n16352 0.00223571
R65617 DVSS.n15926 DVSS.n15922 0.00223571
R65618 DVSS.n15970 DVSS.n15947 0.00223571
R65619 DVSS.n17720 DVSS.n17682 0.00223571
R65620 DVSS.n17727 DVSS.n17680 0.00223571
R65621 DVSS.n15153 DVSS.n15149 0.00223571
R65622 DVSS.n15194 DVSS.n15175 0.00223571
R65623 DVSS.n13691 DVSS.n13687 0.00223571
R65624 DVSS.n20744 DVSS.n13712 0.00223571
R65625 DVSS.n21181 DVSS.n13642 0.00223571
R65626 DVSS.n21188 DVSS.n13640 0.00223571
R65627 DVSS.n22671 DVSS.n729 0.00223571
R65628 DVSS.n22664 DVSS.n714 0.00223571
R65629 DVSS.n23094 DVSS.n246 0.0022122
R65630 DVSS.n13051 DVSS.n1152 0.0022122
R65631 DVSS.n23137 DVSS.n166 0.0022122
R65632 DVSS.n13056 DVSS.n13055 0.0022122
R65633 DVSS.n22503 DVSS.n22482 0.0022122
R65634 DVSS.n13050 DVSS.n1098 0.0022122
R65635 DVSS.n23181 DVSS.n101 0.0022122
R65636 DVSS.n13049 DVSS.n366 0.0022122
R65637 DVSS.n21037 DVSS.n14261 0.00221
R65638 DVSS.n12789 DVSS.n12788 0.00221
R65639 DVSS.n43 DVSS.n42 0.00221
R65640 DVSS.n21980 DVSS.n1234 0.00221
R65641 DVSS.n17895 DVSS.n15802 0.00219014
R65642 DVSS.n15726 DVSS.n15693 0.00219014
R65643 DVSS.n20559 DVSS 0.00218942
R65644 DVSS.n13892 DVSS.n13884 0.00218
R65645 DVSS.n14107 DVSS.n14079 0.00218
R65646 DVSS.n21529 DVSS.n1064 0.00218
R65647 DVSS.n12985 DVSS.n306 0.00218
R65648 DVSS.n22490 DVSS.n796 0.00218
R65649 DVSS.n23121 DVSS.n171 0.00218
R65650 DVSS.n21867 DVSS.n21866 0.00218
R65651 DVSS.n21739 DVSS.n21679 0.00218
R65652 DVSS DVSS.n18712 0.0021723
R65653 DVSS.n16653 DVSS.n16261 0.00217143
R65654 DVSS.n16807 DVSS.n15660 0.00217143
R65655 DVSS.n16115 DVSS.n16080 0.00217143
R65656 DVSS.n17607 DVSS.n17606 0.00217143
R65657 DVSS.n18346 DVSS.n18345 0.00217143
R65658 DVSS.n18317 DVSS.n18316 0.00217143
R65659 DVSS.n18439 DVSS.n14881 0.00217143
R65660 DVSS.n19973 DVSS.n19972 0.00217143
R65661 DVSS.n20821 DVSS.n14481 0.00217143
R65662 DVSS.n20900 DVSS.n14383 0.00217143
R65663 DVSS.n21271 DVSS.n13539 0.00217143
R65664 DVSS.n21350 DVSS.n13442 0.00217143
R65665 DVSS.n22729 DVSS.n621 0.00217143
R65666 DVSS.n22808 DVSS.n522 0.00217143
R65667 DVSS.n22227 DVSS.n710 0.00215789
R65668 DVSS.n22149 DVSS.n22123 0.00215789
R65669 DVSS.n936 DVSS.n920 0.00215789
R65670 DVSS.n1012 DVSS.n988 0.00215789
R65671 DVSS.n22234 DVSS.n466 0.00215789
R65672 DVSS.n22312 DVSS.n1241 0.00215789
R65673 DVSS.n12831 DVSS.n19 0.00215789
R65674 DVSS.n13098 DVSS.n13097 0.00215789
R65675 DVSS.n21055 DVSS.n14234 0.00215
R65676 DVSS.n13099 DVSS.n406 0.00215
R65677 DVSS.n51 DVSS.n35 0.00215
R65678 DVSS.n22325 DVSS.n1252 0.00215
R65679 DVSS.n21938 DVSS.n21559 0.00212439
R65680 DVSS.n21935 DVSS.n21685 0.00212439
R65681 DVSS.n21940 DVSS.n21872 0.00212439
R65682 DVSS.n21934 DVSS.n21779 0.00212439
R65683 DVSS.n6684 DVSS.n6683 0.00212406
R65684 DVSS.n8096 DVSS.n8095 0.00212406
R65685 DVSS.n21116 DVSS.n13837 0.00212
R65686 DVSS.n1479 DVSS.n1060 0.00212
R65687 DVSS.n22483 DVSS.n787 0.00212
R65688 DVSS.n21860 DVSS.n1440 0.00212
R65689 DVSS.n18151 DVSS.n15570 0.00211972
R65690 DVSS.n16584 DVSS.n16556 0.00210714
R65691 DVSS.n15979 DVSS.n15952 0.00210714
R65692 DVSS.n17736 DVSS.n17687 0.00210714
R65693 DVSS.n15203 DVSS.n15180 0.00210714
R65694 DVSS.n20753 DVSS.n13717 0.00210714
R65695 DVSS.n21197 DVSS.n13647 0.00210714
R65696 DVSS.n22655 DVSS.n724 0.00210714
R65697 DVSS.n10112 DVSS.n10111 0.002075
R65698 DVSS.n13354 DVSS.n13353 0.002075
R65699 DVSS.n22186 DVSS.n22185 0.00206316
R65700 DVSS.n960 DVSS.n909 0.00206316
R65701 DVSS.n22393 DVSS.n1006 0.00206316
R65702 DVSS.n22274 DVSS.n1251 0.00206316
R65703 DVSS.n12855 DVSS.n8 0.00206316
R65704 DVSS.n12887 DVSS.n12811 0.00206316
R65705 DVSS.n13899 DVSS.n13880 0.00206
R65706 DVSS.n14075 DVSS.n14032 0.00206
R65707 DVSS.n1481 DVSS.n1061 0.00206
R65708 DVSS.n12981 DVSS.n12980 0.00206
R65709 DVSS.n22485 DVSS.n22484 0.00206
R65710 DVSS.n198 DVSS.n167 0.00206
R65711 DVSS.n21861 DVSS.n1441 0.00206
R65712 DVSS.n21734 DVSS.n21672 0.00206
R65713 DVSS.n17865 DVSS.n15832 0.0020493
R65714 DVSS.n17947 DVSS.n17946 0.0020493
R65715 DVSS.n16669 DVSS.n16257 0.00204286
R65716 DVSS.n16789 DVSS.n15656 0.00204286
R65717 DVSS.n16104 DVSS.n16076 0.00204286
R65718 DVSS.n17552 DVSS.n17543 0.00204286
R65719 DVSS.n15329 DVSS.n15311 0.00204286
R65720 DVSS.n15472 DVSS.n15463 0.00204286
R65721 DVSS.n14913 DVSS.n14877 0.00204286
R65722 DVSS.n15058 DVSS.n15020 0.00204286
R65723 DVSS.n20837 DVSS.n14477 0.00204286
R65724 DVSS.n20916 DVSS.n14379 0.00204286
R65725 DVSS.n21287 DVSS.n13535 0.00204286
R65726 DVSS.n21366 DVSS.n13438 0.00204286
R65727 DVSS.n22745 DVSS.n617 0.00204286
R65728 DVSS.n535 DVSS.n518 0.00204286
R65729 DVSS.n18344 DVSS.n15315 0.00203659
R65730 DVSS.n22756 DVSS.n623 0.00203659
R65731 DVSS.n18326 DVSS.n15387 0.00203659
R65732 DVSS.n22797 DVSS.n573 0.00203659
R65733 DVSS.n18379 DVSS.n15273 0.00203659
R65734 DVSS.n22714 DVSS.n680 0.00203659
R65735 DVSS.n18315 DVSS.n15452 0.00203659
R65736 DVSS.n22838 DVSS.n523 0.00203659
R65737 DVSS.n21051 DVSS.n14239 0.00203
R65738 DVSS.n12793 DVSS.n407 0.00203
R65739 DVSS.n23198 DVSS.n38 0.00203
R65740 DVSS.n21972 DVSS.n1237 0.00203
R65741 DVSS.n20640 DVSS.n20639 0.00201685
R65742 DVSS.n13915 DVSS.n13885 0.002
R65743 DVSS.n14109 DVSS.n14080 0.002
R65744 DVSS.n1471 DVSS.n1065 0.002
R65745 DVSS.n12987 DVSS.n307 0.002
R65746 DVSS.n22500 DVSS.n797 0.002
R65747 DVSS.n189 DVSS.n172 0.002
R65748 DVSS.n21868 DVSS.n1450 0.002
R65749 DVSS.n21726 DVSS.n21682 0.002
R65750 DVSS.n18014 DVSS.n15558 0.00197887
R65751 DVSS.n18119 DVSS.n15613 0.00197857
R65752 DVSS.n18175 DVSS.n15498 0.00197857
R65753 DVSS.n18249 DVSS.n18224 0.00197857
R65754 DVSS.n19928 DVSS.n15108 0.00197857
R65755 DVSS.n20978 DVSS.n14316 0.00197857
R65756 DVSS.n21432 DVSS.n13373 0.00197857
R65757 DVSS.n22879 DVSS.n454 0.00197857
R65758 DVSS.n21035 DVSS.n14260 0.00197
R65759 DVSS.n12787 DVSS.n416 0.00197
R65760 DVSS.n23217 DVSS.n23215 0.00197
R65761 DVSS.n21983 DVSS.n1233 0.00197
R65762 DVSS.n22133 DVSS.n1392 0.00196842
R65763 DVSS.n952 DVSS.n922 0.00196842
R65764 DVSS.n22436 DVSS.n979 0.00196842
R65765 DVSS.n22330 DVSS.n1221 0.00196842
R65766 DVSS.n12847 DVSS.n10 0.00196842
R65767 DVSS.n12879 DVSS.n12809 0.00196842
R65768 DVSS.n23212 DVSS 0.00196
R65769 DVSS.n6681 DVSS.n5891 0.00194966
R65770 DVSS.n4370 DVSS.n4363 0.00194966
R65771 DVSS.n6682 DVSS.n5892 0.00194966
R65772 DVSS.n4368 DVSS.n4364 0.00194966
R65773 DVSS.n21096 DVSS.n13953 0.00194
R65774 DVSS.n14224 DVSS.n14174 0.00194
R65775 DVSS.n21502 DVSS.n1486 0.00194
R65776 DVSS.n1108 DVSS.n289 0.00194
R65777 DVSS.n23005 DVSS.n334 0.00194
R65778 DVSS.n1485 DVSS.n777 0.00194
R65779 DVSS.n239 DVSS.n205 0.00194
R65780 DVSS.n23172 DVSS.n110 0.00194
R65781 DVSS.n1484 DVSS.n1393 0.00194
R65782 DVSS.n21638 DVSS.n21615 0.00194
R65783 DVSS.n21818 DVSS.n21772 0.00194
R65784 DVSS.n1395 DVSS.n779 0.00194
R65785 DVSS.n22548 DVSS.n22547 0.00194
R65786 DVSS.n21503 DVSS.n778 0.00194
R65787 DVSS.n16639 DVSS.n16288 0.00191429
R65788 DVSS.n16815 DVSS.n16164 0.00191429
R65789 DVSS.n17653 DVSS.n17652 0.00191429
R65790 DVSS.n16883 DVSS.n16851 0.00191429
R65791 DVSS.n18380 DVSS.n15259 0.00191429
R65792 DVSS.n15427 DVSS.n15395 0.00191429
R65793 DVSS.n18472 DVSS.n18471 0.00191429
R65794 DVSS.n14995 DVSS.n14957 0.00191429
R65795 DVSS.n20806 DVSS.n20805 0.00191429
R65796 DVSS.n20888 DVSS.n20887 0.00191429
R65797 DVSS.n21257 DVSS.n13566 0.00191429
R65798 DVSS.n21338 DVSS.n21337 0.00191429
R65799 DVSS.n22715 DVSS.n644 0.00191429
R65800 DVSS.n22796 DVSS.n22795 0.00191429
R65801 DVSS.n21128 DVSS.n13744 0.00191
R65802 DVSS.n1488 DVSS.n981 0.00191
R65803 DVSS.n892 DVSS.n773 0.00191
R65804 DVSS.n1430 DVSS.n1377 0.00191
R65805 DVSS.n17849 DVSS.n15862 0.00190845
R65806 DVSS.n17930 DVSS.n15766 0.00190845
R65807 DVSS.n23226 DVSS 0.00188
R65808 DVSS.n13999 DVSS.n13944 0.00188
R65809 DVSS.n14208 DVSS.n14178 0.00188
R65810 DVSS.n1112 DVSS.n280 0.00188
R65811 DVSS.n388 DVSS.n380 0.00188
R65812 DVSS.n23078 DVSS.n242 0.00188
R65813 DVSS.n119 DVSS.n98 0.00188
R65814 DVSS.n21648 DVSS.n21625 0.00188
R65815 DVSS.n21822 DVSS.n21763 0.00188
R65816 DVSS.n10114 DVSS.n2722 0.00187555
R65817 DVSS.n13351 DVSS.n1514 0.00187555
R65818 DVSS.n10113 DVSS.n2724 0.00187555
R65819 DVSS.n13352 DVSS.n1516 0.00187555
R65820 DVSS.n22672 DVSS.n719 0.00187368
R65821 DVSS.n22141 DVSS.n22121 0.00187368
R65822 DVSS.n944 DVSS.n907 0.00187368
R65823 DVSS.n19766 DVSS.n464 0.00187368
R65824 DVSS.n22320 DVSS.n1239 0.00187368
R65825 DVSS.n12839 DVSS.n21 0.00187368
R65826 DVSS.n13016 DVSS.n1126 0.00186098
R65827 DVSS.n13020 DVSS.n12991 0.00186098
R65828 DVSS.n13015 DVSS.n1068 0.00186098
R65829 DVSS.n13014 DVSS.n336 0.00186098
R65830 DVSS.n16753 DVSS.n15601 0.00185
R65831 DVSS.n18191 DVSS.n15502 0.00185
R65832 DVSS.n18265 DVSS.n18229 0.00185
R65833 DVSS.n19944 DVSS.n15113 0.00185
R65834 DVSS.n20944 DVSS.n14347 0.00185
R65835 DVSS.n13798 DVSS.n13739 0.00185
R65836 DVSS.n21398 DVSS.n13405 0.00185
R65837 DVSS.n485 DVSS.n481 0.00185
R65838 DVSS.n1498 DVSS.n985 0.00185
R65839 DVSS.n898 DVSS.n897 0.00185
R65840 DVSS.n1401 DVSS.n1373 0.00185
R65841 DVSS.n13948 DVSS.n13939 0.00182
R65842 DVSS.n21547 DVSS.n1116 0.00182
R65843 DVSS.n22511 DVSS.n247 0.00182
R65844 DVSS.n21630 DVSS.n1460 0.00182
R65845 DVSS.n13782 DVSS.n13732 0.00179
R65846 DVSS.n21486 DVSS.n975 0.00179
R65847 DVSS.n885 DVSS.n767 0.00179
R65848 DVSS.n1420 DVSS.n1366 0.00179
R65849 DVSS.n16623 DVSS.n16318 0.00178571
R65850 DVSS.n16230 DVSS.n16161 0.00178571
R65851 DVSS.n16050 DVSS.n16025 0.00178571
R65852 DVSS.n16860 DVSS.n16846 0.00178571
R65853 DVSS.n18371 DVSS.n15249 0.00178571
R65854 DVSS.n15404 DVSS.n15390 0.00178571
R65855 DVSS.n18417 DVSS.n18390 0.00178571
R65856 DVSS.n14966 DVSS.n14953 0.00178571
R65857 DVSS.n20726 DVSS.n20716 0.00178571
R65858 DVSS.n20871 DVSS.n14436 0.00178571
R65859 DVSS.n21241 DVSS.n13602 0.00178571
R65860 DVSS.n21321 DVSS.n13492 0.00178571
R65861 DVSS.n22699 DVSS.n685 0.00178571
R65862 DVSS.n22779 DVSS.n577 0.00178571
R65863 DVSS.n16548 DVSS.n16335 0.00177895
R65864 DVSS.n22179 DVSS.n1380 0.00177895
R65865 DVSS.n924 DVSS.n900 0.00177895
R65866 DVSS.n22401 DVSS.n991 0.00177895
R65867 DVSS.n18112 DVSS.n15616 0.00177895
R65868 DVSS.n22282 DVSS.n1254 0.00177895
R65869 DVSS.n12863 DVSS.n26 0.00177895
R65870 DVSS.n12895 DVSS.n12802 0.00177895
R65871 DVSS.n21629 DVSS.n21557 0.00177317
R65872 DVSS.n21733 DVSS.n21683 0.00177317
R65873 DVSS.n21946 DVSS.n21945 0.00177317
R65874 DVSS.n21950 DVSS.n21777 0.00177317
R65875 DVSS DVSS.n18878 0.00176405
R65876 DVSS.n18917 DVSS.n18915 0.00176405
R65877 DVSS.n20131 DVSS.n20059 0.00176405
R65878 DVSS.n20078 DVSS.n20060 0.00176405
R65879 DVSS.n20225 DVSS.n20216 0.00176405
R65880 DVSS.n20226 DVSS.n20215 0.00176405
R65881 DVSS.n14686 DVSS.n14676 0.00176405
R65882 DVSS.n14003 DVSS.n13951 0.00176
R65883 DVSS.n14213 DVSS.n14185 0.00176
R65884 DVSS.n1121 DVSS.n1120 0.00176
R65885 DVSS.n390 DVSS.n326 0.00176
R65886 DVSS.n268 DVSS.n252 0.00176
R65887 DVSS.n23157 DVSS.n106 0.00176
R65888 DVSS.n21654 DVSS.n21634 0.00176
R65889 DVSS.n21957 DVSS.n21956 0.00176
R65890 DVSS DVSS.n0 0.00173
R65891 DVSS.n21298 DVSS.n13527 0.00172927
R65892 DVSS.n21339 DVSS.n13481 0.00172927
R65893 DVSS.n21256 DVSS.n13581 0.00172927
R65894 DVSS.n14084 DVSS.n14056 0.0017
R65895 DVSS.n21065 DVSS.n14190 0.0017
R65896 DVSS DVSS.n21403 0.0017
R65897 DVSS.n21555 DVSS.n21554 0.0017
R65898 DVSS.n12990 DVSS.n12972 0.0017
R65899 DVSS.n23002 DVSS.n395 0.0017
R65900 DVSS.n21556 DVSS.n274 0.0017
R65901 DVSS.n159 DVSS.n125 0.0017
R65902 DVSS.n23182 DVSS.n60 0.0017
R65903 DVSS.n22077 DVSS.n22076 0.0017
R65904 DVSS.n21743 DVSS.n21718 0.0017
R65905 DVSS.n21964 DVSS.n21774 0.0017
R65906 DVSS.n22078 DVSS.n271 0.0017
R65907 DVSS.n23075 DVSS.n23074 0.0017
R65908 DVSS.n21553 DVSS.n270 0.0017
R65909 DVSS.n16251 DVSS.n16242 0.00168537
R65910 DVSS.n16176 DVSS.n16166 0.00168537
R65911 DVSS.n16360 DVSS.n16301 0.00168537
R65912 DVSS.n15650 DVSS.n15629 0.00168537
R65913 DVSS.n19212 DVSS.n19172 0.00168421
R65914 DVSS.n19208 DVSS.n19207 0.00168421
R65915 DVSS.n22219 DVSS.n705 0.00168421
R65916 DVSS.n22157 DVSS.n1385 0.00168421
R65917 DVSS.n928 DVSS.n919 0.00168421
R65918 DVSS.n22423 DVSS.n997 0.00168421
R65919 DVSS.n22242 DVSS.n460 0.00168421
R65920 DVSS.n22304 DVSS.n1259 0.00168421
R65921 DVSS.n12823 DVSS.n15 0.00168421
R65922 DVSS.n12917 DVSS.n12797 0.00168421
R65923 DVSS.n21039 DVSS.n14254 0.00167
R65924 DVSS.n12780 DVSS.n413 0.00167
R65925 DVSS.n23208 DVSS.n32 0.00167
R65926 DVSS.n21979 DVSS.n1227 0.00167
R65927 DVSS.n13910 DVSS.n13875 0.00164
R65928 DVSS.n14105 DVSS.n14071 0.00164
R65929 DVSS.n21527 DVSS.n1055 0.00164
R65930 DVSS.n12976 DVSS.n305 0.00164
R65931 DVSS.n22474 DVSS.n795 0.00164
R65932 DVSS.n23119 DVSS.n162 0.00164
R65933 DVSS.n21854 DVSS.n1447 0.00164
R65934 DVSS.n21728 DVSS.n21678 0.00164
R65935 DVSS.n20614 DVSS.n20613 0.00163764
R65936 DVSS.n17844 DVSS.n15861 0.00162676
R65937 DVSS.n17926 DVSS.n15765 0.00162676
R65938 DVSS.n8621 DVSS.n8620 0.001625
R65939 DVSS.n17075 DVSS.n16067 0.00159756
R65940 DVSS.n17616 DVSS.n16843 0.00159756
R65941 DVSS.n17654 DVSS.n16021 0.00159756
R65942 DVSS.n17605 DVSS.n17530 0.00159756
R65943 DVSS.n22213 DVSS.n707 0.00158947
R65944 DVSS.n22163 DVSS.n22126 0.00158947
R65945 DVSS.n22417 DVSS.n1010 0.00158947
R65946 DVSS.n22878 DVSS.n469 0.00158947
R65947 DVSS.n22298 DVSS.n1244 0.00158947
R65948 DVSS.n12911 DVSS.n12816 0.00158947
R65949 DVSS.n6251 DVSS.n6246 0.00158271
R65950 DVSS.n9765 DVSS.n9764 0.00158271
R65951 DVSS.n10483 DVSS.n1616 0.00158271
R65952 DVSS.n21117 DVSS.n13824 0.00158
R65953 DVSS.n21513 DVSS.n1059 0.00158
R65954 DVSS.n22478 DVSS.n786 0.00158
R65955 DVSS.n21859 DVSS.n21858 0.00158
R65956 DVSS.n18018 DVSS.n15559 0.00155634
R65957 DVSS.n17369 DVSS.n15304 0.00155366
R65958 DVSS.n17490 DVSS.n15371 0.00155366
R65959 DVSS.n17378 DVSS.n15265 0.00155366
R65960 DVSS.n17520 DVSS.n15441 0.00155366
R65961 DVSS.n16618 DVSS.n16317 0.00152857
R65962 DVSS.n16698 DVSS.n16224 0.00152857
R65963 DVSS.n16038 DVSS.n16024 0.00152857
R65964 DVSS.n16863 DVSS.n16845 0.00152857
R65965 DVSS.n18378 DVSS.n18377 0.00152857
R65966 DVSS.n15407 DVSS.n15389 0.00152857
R65967 DVSS.n18408 DVSS.n18389 0.00152857
R65968 DVSS.n14969 DVSS.n14952 0.00152857
R65969 DVSS.n20784 DVSS.n20715 0.00152857
R65970 DVSS.n20867 DVSS.n14435 0.00152857
R65971 DVSS.n21236 DVSS.n13601 0.00152857
R65972 DVSS.n21317 DVSS.n13491 0.00152857
R65973 DVSS.n22694 DVSS.n684 0.00152857
R65974 DVSS.n22775 DVSS.n576 0.00152857
R65975 DVSS.n13901 DVSS.n13877 0.00152
R65976 DVSS.n14096 DVSS.n14073 0.00152
R65977 DVSS.n21519 DVSS.n1057 0.00152
R65978 DVSS.n12978 DVSS.n300 0.00152
R65979 DVSS.n22476 DVSS.n790 0.00152
R65980 DVSS.n23111 DVSS.n164 0.00152
R65981 DVSS.n21856 DVSS.n1442 0.00152
R65982 DVSS.n21730 DVSS.n21673 0.00152
R65983 DVSS.n22375 DVSS.n1107 0.00150976
R65984 DVSS.n13061 DVSS.n13060 0.00150976
R65985 DVSS.n22378 DVSS.n22377 0.00150976
R65986 DVSS.n13058 DVSS.n368 0.00150976
R65987 DVSS.n15888 DVSS 0.00149474
R65988 DVSS.n22173 DVSS.n22128 0.00149474
R65989 DVSS.n22446 DVSS.n914 0.00149474
R65990 DVSS.n22407 DVSS.n995 0.00149474
R65991 DVSS.n15536 DVSS 0.00149474
R65992 DVSS.n22288 DVSS.n1246 0.00149474
R65993 DVSS.n12869 DVSS.n5 0.00149474
R65994 DVSS.n12901 DVSS.n12814 0.00149474
R65995 DVSS.n21047 DVSS.n14277 0.00149
R65996 DVSS.n12778 DVSS.n408 0.00149
R65997 DVSS.n23200 DVSS.n34 0.00149
R65998 DVSS.n21973 DVSS.n1225 0.00149
R65999 DVSS.n17863 DVSS.n17861 0.00148592
R66000 DVSS.n15771 DVSS.n15770 0.00148592
R66001 DVSS.n8623 DVSS.n3067 0.00148253
R66002 DVSS.n8622 DVSS.n3068 0.00148253
R66003 DVSS.n2738 DVSS.n2731 0.00146644
R66004 DVSS.n10485 DVSS.n1618 0.00146644
R66005 DVSS.n2736 DVSS.n2732 0.00146644
R66006 DVSS.n10484 DVSS.n1617 0.00146644
R66007 DVSS.n16731 DVSS.n15603 0.00146429
R66008 DVSS.n18197 DVSS.n15503 0.00146429
R66009 DVSS.n18239 DVSS.n18231 0.00146429
R66010 DVSS.n19952 DVSS.n19950 0.00146429
R66011 DVSS.n20963 DVSS.n14349 0.00146429
R66012 DVSS.n21417 DVSS.n13407 0.00146429
R66013 DVSS.n22858 DVSS.n480 0.00146429
R66014 DVSS.n21505 DVSS.n21504 0.00146
R66015 DVSS.n782 DVSS.n775 0.00146
R66016 DVSS.n22116 DVSS.n22115 0.00146
R66017 DVSS.n13917 DVSS.n13873 0.00146
R66018 DVSS.n14088 DVSS.n14069 0.00146
R66019 DVSS.n1473 DVSS.n1053 0.00146
R66020 DVSS.n12986 DVSS.n12974 0.00146
R66021 DVSS.n22499 DVSS.n22498 0.00146
R66022 DVSS.n191 DVSS.n160 0.00146
R66023 DVSS.n21852 DVSS.n1451 0.00146
R66024 DVSS.n22048 DVSS.n22047 0.00146
R66025 DVSS.n22049 DVSS.n187 0.00146
R66026 DVSS.n23127 DVSS.n23126 0.00146
R66027 DVSS.n308 DVSS.n188 0.00146
R66028 DVSS.n21033 DVSS.n14256 0.00143
R66029 DVSS.n12782 DVSS.n417 0.00143
R66030 DVSS.n23216 DVSS.n30 0.00143
R66031 DVSS.n21984 DVSS.n1229 0.00143
R66032 DVSS.n15795 DVSS 0.00142195
R66033 DVSS.n1153 DVSS.n1125 0.00142195
R66034 DVSS.n15538 DVSS 0.00142195
R66035 DVSS.n13088 DVSS.n12962 0.00142195
R66036 DVSS.n15848 DVSS 0.00142195
R66037 DVSS.n22385 DVSS.n1017 0.00142195
R66038 DVSS.n15537 DVSS 0.00142195
R66039 DVSS.n369 DVSS.n335 0.00142195
R66040 DVSS.n18004 DVSS.n15562 0.00141549
R66041 DVSS.n16637 DVSS.n16635 0.0014
R66042 DVSS.n16822 DVSS.n16821 0.0014
R66043 DVSS.n16061 DVSS.n16029 0.0014
R66044 DVSS.n16879 DVSS.n16850 0.0014
R66045 DVSS.n18360 DVSS.n15252 0.0014
R66046 DVSS.n15423 DVSS.n15394 0.0014
R66047 DVSS.n18434 DVSS.n18433 0.0014
R66048 DVSS.n14985 DVSS.n14956 0.0014
R66049 DVSS.n20803 DVSS.n20801 0.0014
R66050 DVSS.n14445 DVSS.n14439 0.0014
R66051 DVSS.n21097 DVSS.n13952 0.0014
R66052 DVSS.n14222 DVSS.n14188 0.0014
R66053 DVSS.n21255 DVSS.n21253 0.0014
R66054 DVSS.n13502 DVSS.n13495 0.0014
R66055 DVSS.n22229 DVSS.n703 0.0014
R66056 DVSS.n22147 DVSS.n1387 0.0014
R66057 DVSS.n938 DVSS.n903 0.0014
R66058 DVSS.n22434 DVSS.n22433 0.0014
R66059 DVSS.n22232 DVSS.n462 0.0014
R66060 DVSS.n22314 DVSS.n1261 0.0014
R66061 DVSS.n12833 DVSS.n13 0.0014
R66062 DVSS.n12795 DVSS.n12776 0.0014
R66063 DVSS.n22713 DVSS.n22711 0.0014
R66064 DVSS.n582 DVSS.n581 0.0014
R66065 DVSS.n1124 DVSS.n1123 0.0014
R66066 DVSS.n394 DVSS.n331 0.0014
R66067 DVSS.n23093 DVSS.n23092 0.0014
R66068 DVSS.n23173 DVSS.n109 0.0014
R66069 DVSS.n21662 DVSS.n21637 0.0014
R66070 DVSS.n21961 DVSS.n21960 0.0014
R66071 DVSS.n13779 DVSS.n13730 0.00137
R66072 DVSS.n21494 DVSS.n977 0.00137
R66073 DVSS.n887 DVSS.n772 0.00137
R66074 DVSS.n1428 DVSS.n1364 0.00137
R66075 DVSS.n15821 DVSS.n15801 0.00134507
R66076 DVSS.n18040 DVSS.n15723 0.00134507
R66077 DVSS DVSS.n21034 0.00134
R66078 DVSS.n13983 DVSS.n13949 0.00134
R66079 DVSS.n14206 DVSS.n14183 0.00134
R66080 DVSS.n21033 DVSS 0.00134
R66081 DVSS.n1118 DVSS.n279 0.00134
R66082 DVSS.n387 DVSS.n322 0.00134
R66083 DVSS.n23076 DVSS.n250 0.00134
R66084 DVSS.n117 DVSS.n104 0.00134
R66085 DVSS.n22075 DVSS.n21591 0.00134
R66086 DVSS.n21954 DVSS.n21762 0.00134
R66087 DVSS.n21984 DVSS 0.00134
R66088 DVSS DVSS.n21995 0.00134
R66089 DVSS.n16742 DVSS.n15607 0.00133571
R66090 DVSS.n18180 DVSS.n15499 0.00133571
R66091 DVSS.n18254 DVSS.n18226 0.00133571
R66092 DVSS.n19933 DVSS.n15110 0.00133571
R66093 DVSS.n14344 DVSS.n14342 0.00133571
R66094 DVSS.n13402 DVSS.n13400 0.00133571
R66095 DVSS.n22877 DVSS.n22875 0.00133571
R66096 DVSS.n662 DVSS.n600 0.00133415
R66097 DVSS.n660 DVSS.n551 0.00133415
R66098 DVSS.n664 DVSS.n652 0.00133415
R66099 DVSS.n659 DVSS.n500 0.00133415
R66100 DVSS.n6453 DVSS.n6252 0.00131203
R66101 DVSS.n13789 DVSS.n13736 0.00131
R66102 DVSS.n13796 DVSS.n13734 0.00131
R66103 DVSS.n22435 DVSS.n987 0.00131
R66104 DVSS.n1496 DVSS.n973 0.00131
R66105 DVSS.n22452 DVSS.n758 0.00131
R66106 DVSS.n883 DVSS.n763 0.00131
R66107 DVSS.n1407 DVSS.n1371 0.00131
R66108 DVSS.n1414 DVSS.n1368 0.00131
R66109 DVSS.n16527 DVSS.n16336 0.00130526
R66110 DVSS.n16529 DVSS.n16342 0.00130526
R66111 DVSS.n16531 DVSS.n16337 0.00130526
R66112 DVSS.n16533 DVSS.n16341 0.00130526
R66113 DVSS.n16535 DVSS.n16338 0.00130526
R66114 DVSS.n16537 DVSS.n16343 0.00130526
R66115 DVSS.n16540 DVSS.n16335 0.00130526
R66116 DVSS.n16596 DVSS.n16344 0.00130526
R66117 DVSS.n958 DVSS.n916 0.00130526
R66118 DVSS.n22391 DVSS.n993 0.00130526
R66119 DVSS.n18124 DVSS.n15589 0.00130526
R66120 DVSS.n18121 DVSS.n18120 0.00130526
R66121 DVSS.n15614 DVSS.n15598 0.00130526
R66122 DVSS.n18096 DVSS.n15612 0.00130526
R66123 DVSS.n18098 DVSS.n15615 0.00130526
R66124 DVSS.n18100 DVSS.n15611 0.00130526
R66125 DVSS.n18108 DVSS.n15616 0.00130526
R66126 DVSS.n18111 DVSS.n15610 0.00130526
R66127 DVSS.n12853 DVSS.n24 0.00130526
R66128 DVSS.n12885 DVSS.n12804 0.00130526
R66129 DVSS.n23071 DVSS.n277 0.0013
R66130 DVSS.n23073 DVSS.n23072 0.0013
R66131 DVSS.n22079 DVSS.n276 0.0013
R66132 DVSS.n12760 DVSS.n12750 0.00128471
R66133 DVSS.n12757 DVSS.n12750 0.00128471
R66134 DVSS.n13990 DVSS.n13946 0.00128
R66135 DVSS.n21068 DVSS.n21067 0.00128
R66136 DVSS.n1464 DVSS.n1114 0.00128
R66137 DVSS.n383 DVSS.n382 0.00128
R66138 DVSS.n22512 DVSS.n244 0.00128
R66139 DVSS.n122 DVSS.n100 0.00128
R66140 DVSS.n21626 DVSS.n1461 0.00128
R66141 DVSS.n21824 DVSS.n21758 0.00128
R66142 DVSS.n17814 DVSS.n15907 0.00127465
R66143 DVSS.n16276 DVSS.n16256 0.00127143
R66144 DVSS.n16785 DVSS.n15655 0.00127143
R66145 DVSS.n16106 DVSS.n16101 0.00127143
R66146 DVSS.n17586 DVSS.n17542 0.00127143
R66147 DVSS.n15350 DVSS.n15310 0.00127143
R66148 DVSS.n18296 DVSS.n15462 0.00127143
R66149 DVSS.n14915 DVSS.n14909 0.00127143
R66150 DVSS.n15038 DVSS.n15019 0.00127143
R66151 DVSS.n14491 DVSS.n14476 0.00127143
R66152 DVSS.n20920 DVSS.n14378 0.00127143
R66153 DVSS.n13554 DVSS.n13553 0.00127143
R66154 DVSS.n21370 DVSS.n13437 0.00127143
R66155 DVSS.n632 DVSS.n616 0.00127143
R66156 DVSS.n22828 DVSS.n517 0.00127143
R66157 DVSS.n18868 DVSS.n18867 0.00125843
R66158 DVSS.n18908 DVSS.n18907 0.00125843
R66159 DVSS.n20441 DVSS.n14680 0.00125843
R66160 DVSS.n13805 DVSS.n13741 0.00125
R66161 DVSS.n1492 DVSS.n983 0.00125
R66162 DVSS.n895 DVSS.n768 0.00125
R66163 DVSS.n1422 DVSS.n1375 0.00125
R66164 DVSS.n16638 DVSS.n16304 0.00124634
R66165 DVSS.n16313 DVSS.n16293 0.00124634
R66166 DVSS.n16418 DVSS.n16303 0.00124634
R66167 DVSS.n16420 DVSS.n16294 0.00124634
R66168 DVSS.n16422 DVSS.n16302 0.00124634
R66169 DVSS.n16424 DVSS.n16295 0.00124634
R66170 DVSS.n16466 DVSS.n16301 0.00124634
R66171 DVSS.n16463 DVSS.n16296 0.00124634
R66172 DVSS.n18071 DVSS.n15669 0.00124634
R66173 DVSS.n18078 DVSS.n15679 0.00124634
R66174 DVSS.n18077 DVSS.n15670 0.00124634
R66175 DVSS.n18074 DVSS.n15678 0.00124634
R66176 DVSS.n18080 DVSS.n15652 0.00124634
R66177 DVSS.n18081 DVSS.n15646 0.00124634
R66178 DVSS.n18084 DVSS.n15650 0.00124634
R66179 DVSS.n15644 DVSS.n15630 0.00124634
R66180 DVSS.n13980 DVSS.n13942 0.00122
R66181 DVSS.n14215 DVSS.n14176 0.00122
R66182 DVSS.n1110 DVSS.n284 0.00122
R66183 DVSS.n378 DVSS.n327 0.00122
R66184 DVSS.n402 DVSS.n55 0.00122
R66185 DVSS.n23084 DVSS.n240 0.00122
R66186 DVSS.n113 DVSS.n96 0.00122
R66187 DVSS.n23190 DVSS.n23189 0.00122
R66188 DVSS.n21643 DVSS.n21623 0.00122
R66189 DVSS.n21820 DVSS.n21767 0.00122
R66190 DVSS.n21967 DVSS.n54 0.00122
R66191 DVSS.n22014 DVSS.n22013 0.00122
R66192 DVSS.n23188 DVSS.n53 0.00122
R66193 DVSS.n22996 DVSS.n22995 0.00122
R66194 DVSS.n955 DVSS.n901 0.00121053
R66195 DVSS.n22388 DVSS.n992 0.00121053
R66196 DVSS.n12850 DVSS.n23 0.00121053
R66197 DVSS.n12882 DVSS.n12805 0.00121053
R66198 DVSS.n16588 DVSS.n16558 0.00120714
R66199 DVSS.n15958 DVSS.n15953 0.00120714
R66200 DVSS.n17706 DVSS.n17689 0.00120714
R66201 DVSS.n15209 DVSS.n15182 0.00120714
R66202 DVSS.n20757 DVSS.n13718 0.00120714
R66203 DVSS.n21206 DVSS.n13649 0.00120714
R66204 DVSS.n22651 DVSS.n723 0.00120714
R66205 DVSS.n17884 DVSS.n15805 0.00120422
R66206 DVSS.n17963 DVSS.n15724 0.00120422
R66207 DVSS.n21027 DVSS.n14258 0.00119
R66208 DVSS.n12785 DVSS.n421 0.00119
R66209 DVSS.n23222 DVSS.n23221 0.00119
R66210 DVSS.n21989 DVSS.n1231 0.00119
R66211 DVSS.n7052 DVSS.n7051 0.001175
R66212 DVSS.n21114 DVSS.n21113 0.00116
R66213 DVSS.n14118 DVSS.n14083 0.00116
R66214 DVSS.n22379 DVSS.n1083 0.00116
R66215 DVSS.n12989 DVSS.n312 0.00116
R66216 DVSS.n22505 DVSS.n22504 0.00116
R66217 DVSS.n23136 DVSS.n23135 0.00116
R66218 DVSS.n21944 DVSS.n1455 0.00116
R66219 DVSS.n21752 DVSS.n21742 0.00116
R66220 DVSS.n16658 DVSS.n16260 0.00114286
R66221 DVSS.n16716 DVSS.n15659 0.00114286
R66222 DVSS.n16119 DVSS.n16102 0.00114286
R66223 DVSS.n17604 DVSS.n17603 0.00114286
R66224 DVSS.n15334 DVSS.n15314 0.00114286
R66225 DVSS.n18314 DVSS.n18313 0.00114286
R66226 DVSS.n18454 DVSS.n14910 0.00114286
R66227 DVSS.n15047 DVSS.n15023 0.00114286
R66228 DVSS.n20826 DVSS.n14480 0.00114286
R66229 DVSS.n14402 DVSS.n14382 0.00114286
R66230 DVSS.n21276 DVSS.n13538 0.00114286
R66231 DVSS.n13457 DVSS.n13441 0.00114286
R66232 DVSS.n22734 DVSS.n620 0.00114286
R66233 DVSS.n22812 DVSS.n521 0.00114286
R66234 DVSS.n23035 DVSS.n23034 0.00114
R66235 DVSS.n23125 DVSS.n186 0.00114
R66236 DVSS.n22050 DVSS.n21681 0.00114
R66237 DVSS.n17796 DVSS.n15898 0.0011338
R66238 DVSS.n15914 DVSS.n15902 0.0011338
R66239 DVSS.n21041 DVSS.n14262 0.00113
R66240 DVSS.n12790 DVSS.n412 0.00113
R66241 DVSS.n23206 DVSS.n41 0.00113
R66242 DVSS.n21978 DVSS.n1235 0.00113
R66243 DVSS.n19421 DVSS.n702 0.00111579
R66244 DVSS.n22144 DVSS.n1388 0.00111579
R66245 DVSS.n942 DVSS.n918 0.00111579
R66246 DVSS.n19764 DVSS.n463 0.00111579
R66247 DVSS.n22318 DVSS.n1262 0.00111579
R66248 DVSS.n12837 DVSS.n12 0.00111579
R66249 DVSS.n13908 DVSS.n13883 0.0011
R66250 DVSS.n14091 DVSS.n14078 0.0011
R66251 DVSS.n1477 DVSS.n1063 0.0011
R66252 DVSS.n12984 DVSS.n12983 0.0011
R66253 DVSS.n22489 DVSS.n22488 0.0011
R66254 DVSS.n195 DVSS.n170 0.0011
R66255 DVSS.n21865 DVSS.n1446 0.0011
R66256 DVSS.n21738 DVSS.n21677 0.0011
R66257 DVSS.n7049 DVSS.n5575 0.00108952
R66258 DVSS.n7050 DVSS.n7048 0.00108952
R66259 DVSS.n16570 DVSS.n16353 0.00107857
R66260 DVSS.n16565 DVSS.n16553 0.00107857
R66261 DVSS.n17780 DVSS.n17779 0.00107857
R66262 DVSS.n15949 DVSS.n15948 0.00107857
R66263 DVSS.n17717 DVSS.n17681 0.00107857
R66264 DVSS.n17725 DVSS.n17684 0.00107857
R66265 DVSS.n18493 DVSS.n18492 0.00107857
R66266 DVSS.n15177 DVSS.n15176 0.00107857
R66267 DVSS.n21148 DVSS.n21147 0.00107857
R66268 DVSS.n13714 DVSS.n13713 0.00107857
R66269 DVSS.n21183 DVSS.n13641 0.00107857
R66270 DVSS.n13656 DVSS.n13644 0.00107857
R66271 DVSS.n22670 DVSS.n713 0.00107857
R66272 DVSS.n731 DVSS.n728 0.00107857
R66273 DVSS.n6657 DVSS.n6237 0.00106946
R66274 DVSS.n7797 DVSS.n7461 0.00106946
R66275 DVSS.n3946 DVSS.n3846 0.00106946
R66276 DVSS.n13122 DVSS.n13121 0.00106946
R66277 DVSS.n6688 DVSS.n5890 0.00106487
R66278 DVSS.n10498 DVSS.n10497 0.00106487
R66279 DVSS.n15827 DVSS.n15815 0.00106338
R66280 DVSS.n17961 DVSS.n15725 0.00106338
R66281 DVSS.n14305 DVSS 0.00106
R66282 DVSS.n9770 DVSS.n2730 0.0010465
R66283 DVSS.n8629 DVSS.n8628 0.00104135
R66284 DVSS.n13135 DVSS.n13134 0.00104135
R66285 DVSS.n8332 DVSS.n8331 0.00103731
R66286 DVSS.n2936 DVSS.n2932 0.00103731
R66287 DVSS.n6652 DVSS.n6257 0.00103272
R66288 DVSS.n6602 DVSS.n6258 0.00103272
R66289 DVSS.n6259 DVSS.n6256 0.00103272
R66290 DVSS.n6661 DVSS.n6656 0.00103272
R66291 DVSS.n8616 DVSS.n8614 0.00102813
R66292 DVSS.n9184 DVSS.n2878 0.00102813
R66293 DVSS.n16596 DVSS.n16550 0.00102105
R66294 DVSS.n22177 DVSS.n22129 0.00102105
R66295 DVSS.n22451 DVSS.n22450 0.00102105
R66296 DVSS.n22404 DVSS.n1009 0.00102105
R66297 DVSS.n18114 DVSS.n15610 0.00102105
R66298 DVSS.n22285 DVSS.n1247 0.00102105
R66299 DVSS.n12866 DVSS.n6 0.00102105
R66300 DVSS.n12898 DVSS.n12813 0.00102105
R66301 DVSS DVSS.n415 0.00102
R66302 DVSS.n3904 DVSS.n3900 0.00101894
R66303 DVSS.n9199 DVSS.n9198 0.00101894
R66304 DVSS.n16283 DVSS.n16270 0.00101429
R66305 DVSS.n16803 DVSS.n15661 0.00101429
R66306 DVSS.n16117 DVSS.n16103 0.00101429
R66307 DVSS.n16901 DVSS.n16894 0.00101429
R66308 DVSS.n15317 DVSS.n15298 0.00101429
R66309 DVSS.n15444 DVSS.n15438 0.00101429
R66310 DVSS.n18456 DVSS.n14912 0.00101429
R66311 DVSS.n15025 DVSS.n15006 0.00101429
R66312 DVSS.n14498 DVSS.n14485 0.00101429
R66313 DVSS.n20902 DVSS.n14385 0.00101429
R66314 DVSS.n13561 DVSS.n13543 0.00101429
R66315 DVSS.n21352 DVSS.n13444 0.00101429
R66316 DVSS.n639 DVSS.n626 0.00101429
R66317 DVSS.n22810 DVSS.n525 0.00101429
R66318 DVSS.n4469 DVSS.n4371 0.00100976
R66319 DVSS.n18884 DVSS.n18880 0.00100562
R66320 DVSS DVSS.n14689 0.00100562
R66321 DVSS.n20440 DVSS.n14691 0.00100562
R66322 DVSS.n2073 DVSS.n2027 0.00100517
R66323 DVSS.n10460 DVSS.n2019 0.00100057
R66324 DVSS.n17812 DVSS.n15894 0.000992958
R66325 DVSS.n7069 DVSS.n5525 0.000991389
R66326 DVSS.n7796 DVSS.n7795 0.000991389
R66327 DVSS.n11111 DVSS.n11110 0.000991389
R66328 DVSS.n19316 DVSS.n19315 0.00098913
R66329 DVSS.n22429 DVSS.n22428 0.00098913
R66330 DVSS.n19658 DVSS.n19657 0.00098913
R66331 DVSS.n8626 DVSS.n3060 0.000983221
R66332 DVSS.n13132 DVSS.n11502 0.000983221
R66333 DVSS.n8627 DVSS.n3061 0.000983221
R66334 DVSS.n13133 DVSS.n11619 0.000983221
R66335 DVSS.n16680 DVSS.n16267 0.000982927
R66336 DVSS.n22369 DVSS.n1138 0.000982927
R66337 DVSS.n16823 DVSS.n16223 0.000982927
R66338 DVSS.n13008 DVSS.n12961 0.000982927
R66339 DVSS.n16470 DVSS.n16296 0.000982927
R66340 DVSS.n22383 DVSS.n22380 0.000982927
R66341 DVSS.n18088 DVSS.n15630 0.000982927
R66342 DVSS.n13093 DVSS.n351 0.000982927
R66343 DVSS.n7087 DVSS.n5176 0.000982204
R66344 DVSS.n11458 DVSS.n11457 0.000982204
R66345 DVSS.n22997 DVSS.n401 0.00098
R66346 DVSS.n23187 DVSS.n52 0.00098
R66347 DVSS.n21970 DVSS.n21776 0.00098
R66348 DVSS.n13895 DVSS.n13882 0.00098
R66349 DVSS.n14098 DVSS.n14077 0.00098
R66350 DVSS.n21521 DVSS.n1062 0.00098
R66351 DVSS.n12982 DVSS.n301 0.00098
R66352 DVSS.n22487 DVSS.n791 0.00098
R66353 DVSS.n23113 DVSS.n169 0.00098
R66354 DVSS.n21864 DVSS.n21862 0.00098
R66355 DVSS.n21736 DVSS.n21674 0.00098
R66356 DVSS.n7451 DVSS.n4825 0.000977612
R66357 DVSS.n7807 DVSS.n7806 0.00097302
R66358 DVSS.n10152 DVSS.n2364 0.00097302
R66359 DVSS.n13340 DVSS.n11153 0.00097302
R66360 DVSS.n8102 DVSS.n8101 0.000963835
R66361 DVSS.n13120 DVSS.n11631 0.000959242
R66362 DVSS.n12337 DVSS.n12336 0.000959242
R66363 DVSS.n3848 DVSS.n3755 0.00095465
R66364 DVSS.n9188 DVSS.n2890 0.00095465
R66365 DVSS.n16586 DVSS.n16349 0.00095
R66366 DVSS.n15981 DVSS.n15944 0.00095
R66367 DVSS.n17738 DVSS.n17677 0.00095
R66368 DVSS.n15189 DVSS.n15172 0.00095
R66369 DVSS.n20755 DVSS.n13709 0.00095
R66370 DVSS.n21046 DVSS.n14263 0.00095
R66371 DVSS.n21199 DVSS.n13637 0.00095
R66372 DVSS.n22653 DVSS.n717 0.00095
R66373 DVSS.n12792 DVSS.n12791 0.00095
R66374 DVSS.n46 DVSS.n40 0.00095
R66375 DVSS.n21974 DVSS.n1236 0.00095
R66376 DVSS.n7033 DVSS.n5880 0.000945465
R66377 DVSS.n8635 DVSS.n8634 0.000945465
R66378 DVSS.n5889 DVSS.n5878 0.000940873
R66379 DVSS.n8321 DVSS.n3858 0.00093628
R66380 DVSS.n2880 DVSS.n2787 0.00093628
R66381 DVSS.n10166 DVSS.n2070 0.00093628
R66382 DVSS.n10126 DVSS.n2706 0.000927095
R66383 DVSS.n22217 DVSS.n708 0.000926316
R66384 DVSS.n22160 DVSS.n22125 0.000926316
R66385 DVSS.n926 DVSS.n905 0.000926316
R66386 DVSS.n22421 DVSS.n1003 0.000926316
R66387 DVSS.n22245 DVSS.n468 0.000926316
R66388 DVSS.n22302 DVSS.n1243 0.000926316
R66389 DVSS.n12821 DVSS.n17 0.000926316
R66390 DVSS.n12915 DVSS.n12817 0.000926316
R66391 DVSS.n17897 DVSS.n15820 0.000922535
R66392 DVSS.n18044 DVSS.n18043 0.000922535
R66393 DVSS.n11981 DVSS.n11980 0.000922503
R66394 DVSS.n12756 DVSS.n12359 0.000922503
R66395 DVSS.n12758 DVSS.n12506 0.000922503
R66396 DVSS.n12754 DVSS.n12360 0.000922503
R66397 DVSS.n12553 DVSS.n12361 0.000922503
R66398 DVSS.n13919 DVSS.n13887 0.00092
R66399 DVSS.n14114 DVSS.n14082 0.00092
R66400 DVSS.n21535 DVSS.n1066 0.00092
R66401 DVSS.n12988 DVSS.n310 0.00092
R66402 DVSS.n22502 DVSS.n800 0.00092
R66403 DVSS.n23128 DVSS.n173 0.00092
R66404 DVSS.n21869 DVSS.n1452 0.00092
R66405 DVSS.n21741 DVSS.n21694 0.00092
R66406 DVSS.n7079 DVSS.n5182 0.00091791
R66407 DVSS.n7044 DVSS.n5867 0.000908726
R66408 DVSS.n10755 DVSS.n10754 0.000908726
R66409 DVSS.n13359 DVSS.n1511 0.000908726
R66410 DVSS.n2013 DVSS.n2012 0.000904133
R66411 DVSS.n10496 DVSS.n1568 0.000904133
R66412 DVSS.n7103 DVSS.n4832 0.000894948
R66413 DVSS.n7816 DVSS.n7815 0.000890356
R66414 DVSS.n10143 DVSS.n10142 0.000890356
R66415 DVSS.n13337 DVSS.n11198 0.000890356
R66416 DVSS.n13111 DVSS.n13110 0.000890356
R66417 DVSS.n21031 DVSS.n14259 0.00089
R66418 DVSS.n12786 DVSS.n418 0.00089
R66419 DVSS.n23219 DVSS.n1 0.00089
R66420 DVSS.n21985 DVSS.n1232 0.00089
R66421 DVSS.n16671 DVSS.n16275 0.000885714
R66422 DVSS.n16787 DVSS.n15665 0.000885714
R66423 DVSS.n17640 DVSS.n17639 0.000885714
R66424 DVSS.n17588 DVSS.n16905 0.000885714
R66425 DVSS.n15348 DVSS.n15322 0.000885714
R66426 DVSS.n18298 DVSS.n15448 0.000885714
R66427 DVSS.n20006 DVSS.n20005 0.000885714
R66428 DVSS.n15060 DVSS.n15030 0.000885714
R66429 DVSS.n20839 DVSS.n14490 0.000885714
R66430 DVSS.n20918 DVSS.n14390 0.000885714
R66431 DVSS.n21289 DVSS.n13547 0.000885714
R66432 DVSS.n21368 DVSS.n13449 0.000885714
R66433 DVSS.n22747 DVSS.n631 0.000885714
R66434 DVSS.n22826 DVSS.n530 0.000885714
R66435 DVSS.n10486 DVSS.n1620 0.000876579
R66436 DVSS.n6680 DVSS.n5888 0.000871986
R66437 DVSS.n8090 DVSS.n4413 0.000871986
R66438 DVSS.n8590 DVSS.n8589 0.000871986
R66439 DVSS.n3046 DVSS.n3045 0.000871986
R66440 DVSS.n10115 DVSS.n2720 0.000862801
R66441 DVSS.n21099 DVSS.n13977 0.00086
R66442 DVSS.n14194 DVSS.n14175 0.00086
R66443 DVSS.n1164 DVSS.n286 0.00086
R66444 DVSS.n377 DVSS.n330 0.00086
R66445 DVSS.n263 DVSS.n262 0.00086
R66446 DVSS.n23163 DVSS.n95 0.00086
R66447 DVSS.n21660 DVSS.n21622 0.00086
R66448 DVSS.n21819 DVSS.n21769 0.00086
R66449 DVSS.n13326 DVSS.n11500 0.000858209
R66450 DVSS.n4015 DVSS.n4014 0.000853617
R66451 DVSS.n9457 DVSS.n9456 0.000853617
R66452 DVSS.n15563 DVSS.n15548 0.000852113
R66453 DVSS.n17332 DVSS.n15305 0.000851219
R66454 DVSS.n17366 DVSS.n15293 0.000851219
R66455 DVSS.n16940 DVSS.n15372 0.000851219
R66456 DVSS.n17492 DVSS.n15364 0.000851219
R66457 DVSS.n17372 DVSS.n15266 0.000851219
R66458 DVSS.n17312 DVSS.n15255 0.000851219
R66459 DVSS.n16938 DVSS.n15442 0.000851219
R66460 DVSS.n16936 DVSS.n15434 0.000851219
R66461 DVSS.n11109 DVSS.n10766 0.000844432
R66462 DVSS.n12761 DVSS.n12748 0.000844432
R66463 DVSS.n2729 DVSS.n2718 0.000839839
R66464 DVSS.n11646 DVSS.n11622 0.000839839
R66465 DVSS.n6671 DVSS.n6670 0.000835247
R66466 DVSS.n5184 DVSS.n5183 0.000835247
R66467 DVSS.n7105 DVSS.n7104 0.000835247
R66468 DVSS.n11643 DVSS.n11546 0.000835247
R66469 DVSS.n22216 DVSS.n706 0.000831579
R66470 DVSS.n22161 DVSS.n1384 0.000831579
R66471 DVSS.n22453 DVSS.n889 0.000831579
R66472 DVSS.n22420 DVSS.n989 0.000831579
R66473 DVSS.n22246 DVSS.n459 0.000831579
R66474 DVSS.n22301 DVSS.n1258 0.000831579
R66475 DVSS.n12820 DVSS.n16 0.000831579
R66476 DVSS.n12914 DVSS.n12798 0.000831579
R66477 DVSS.n13809 DVSS.n13743 0.00083
R66478 DVSS.n21492 DVSS.n982 0.00083
R66479 DVSS.n893 DVSS.n771 0.00083
R66480 DVSS.n1399 DVSS.n1376 0.00083
R66481 DVSS.n7045 DVSS.n5577 0.000826062
R66482 DVSS.n5577 DVSS.n5531 0.000826062
R66483 DVSS.n7059 DVSS.n5574 0.000826062
R66484 DVSS.n13350 DVSS.n10765 0.000826062
R66485 DVSS.n8625 DVSS.n3066 0.00082147
R66486 DVSS.n10478 DVSS.n10475 0.00082147
R66487 DVSS.n15608 DVSS.n15591 0.000821429
R66488 DVSS.n15530 DVSS.n15497 0.000821429
R66489 DVSS.n18246 DVSS.n18223 0.000821429
R66490 DVSS.n15124 DVSS.n15107 0.000821429
R66491 DVSS.n20979 DVSS.n14320 0.000821429
R66492 DVSS.n21433 DVSS.n13377 0.000821429
R66493 DVSS.n22880 DVSS.n458 0.000821429
R66494 DVSS.n6670 DVSS.n6239 0.000816877
R66495 DVSS.n10478 DVSS.n10477 0.000816877
R66496 DVSS.n7818 DVSS.n7817 0.000807692
R66497 DVSS.n2708 DVSS.n2370 0.000807692
R66498 DVSS.n13358 DVSS.n1512 0.000807692
R66499 DVSS.n12748 DVSS.n11995 0.000807692
R66500 DVSS.n4886 DVSS.n4885 0.0008031
R66501 DVSS.n13994 DVSS.n13978 0.0008
R66502 DVSS.n14204 DVSS.n14179 0.0008
R66503 DVSS.n21554 DVSS.n1113 0.0008
R66504 DVSS.n381 DVSS.n321 0.0008
R66505 DVSS.n274 DVSS.n243 0.0008
R66506 DVSS.n23149 DVSS.n99 0.0008
R66507 DVSS.n30 DVSS 0.0008
R66508 DVSS.n22077 DVSS.n1463 0.0008
R66509 DVSS.n21953 DVSS.n21823 0.0008
R66510 DVSS.n9456 DVSS.n2739 0.000798507
R66511 DVSS.n10476 DVSS.n1961 0.000793915
R66512 DVSS.n6238 DVSS.n6231 0.000789323
R66513 DVSS.n8100 DVSS.n4362 0.000789323
R66514 DVSS.n8605 DVSS.n3415 0.000789323
R66515 DVSS.n8624 DVSS.n3059 0.000789323
R66516 DVSS.n8979 DVSS.n8978 0.000789323
R66517 DVSS.n17866 DVSS.n15836 0.00078169
R66518 DVSS.n17945 DVSS.n15756 0.00078169
R66519 DVSS.n8589 DVSS.n3415 0.000780138
R66520 DVSS.n13323 DVSS.n11546 0.000775545
R66521 DVSS.n8112 DVSS.n8111 0.000770953
R66522 DVSS.n9760 DVSS.n2739 0.000770953
R66523 DVSS.n2781 DVSS.n2728 0.000770953
R66524 DVSS.n13791 DVSS.n13735 0.00077
R66525 DVSS.n13785 DVSS.n13738 0.00077
R66526 DVSS.n1001 DVSS.n972 0.00077
R66527 DVSS.n21478 DVSS.n986 0.00077
R66528 DVSS.n882 DVSS.n761 0.00077
R66529 DVSS.n899 DVSS.n762 0.00077
R66530 DVSS.n1406 DVSS.n1369 0.00077
R66531 DVSS.n1412 DVSS.n1372 0.00077
R66532 DVSS.n7817 DVSS.n7816 0.000761768
R66533 DVSS.n7827 DVSS.n4468 0.000761768
R66534 DVSS.n4471 DVSS.n4470 0.000761768
R66535 DVSS.n13110 DVSS.n11995 0.000761768
R66536 DVSS.n7836 DVSS.n4362 0.000757176
R66537 DVSS.n8112 DVSS.n4021 0.000757176
R66538 DVSS.n8604 DVSS.n3457 0.000757176
R66539 DVSS.n8601 DVSS.n3406 0.000757176
R66540 DVSS.n16640 DVSS.n16292 0.000757143
R66541 DVSS.n16227 DVSS.n16184 0.000757143
R66542 DVSS.n16030 DVSS.n16010 0.000757143
R66543 DVSS.n16881 DVSS.n16837 0.000757143
R66544 DVSS.n15271 DVSS.n15253 0.000757143
R66545 DVSS.n15425 DVSS.n15381 0.000757143
R66546 DVSS.n18400 DVSS.n18399 0.000757143
R66547 DVSS.n14993 DVSS.n14992 0.000757143
R66548 DVSS.n20704 DVSS.n14506 0.000757143
R66549 DVSS.n20886 DVSS.n14444 0.000757143
R66550 DVSS.n21258 DVSS.n13570 0.000757143
R66551 DVSS.n21336 DVSS.n13501 0.000757143
R66552 DVSS.n22716 DVSS.n648 0.000757143
R66553 DVSS.n22794 DVSS.n566 0.000757143
R66554 DVSS.n6239 DVSS.n6238 0.000752583
R66555 DVSS.n4885 DVSS.n4840 0.000752583
R66556 DVSS.n10477 DVSS.n10476 0.000752583
R66557 DVSS.n11504 DVSS.n11500 0.000752583
R66558 DVSS.n8615 DVSS.n3066 0.000747991
R66559 DVSS.n7045 DVSS.n7044 0.000743398
R66560 DVSS.n7060 DVSS.n5531 0.000743398
R66561 DVSS.n10127 DVSS.n2415 0.000743398
R66562 DVSS.n10141 DVSS.n2370 0.000743398
R66563 DVSS.n13359 DVSS.n13358 0.000743398
R66564 DVSS.n13350 DVSS.n13349 0.000743398
R66565 DVSS.n13992 DVSS.n13979 0.00074
R66566 DVSS.n14182 DVSS.n14138 0.00074
R66567 DVSS.n1466 DVSS.n1117 0.00074
R66568 DVSS.n386 DVSS.n320 0.00074
R66569 DVSS.n272 DVSS.n249 0.00074
R66570 DVSS.n23147 DVSS.n103 0.00074
R66571 DVSS.n21632 DVSS.n1462 0.00074
R66572 DVSS.n21952 DVSS.n21759 0.00074
R66573 DVSS.n8633 DVSS.n3059 0.000738806
R66574 DVSS.n15899 DVSS.n15879 0.000736842
R66575 DVSS.n22176 DVSS.n1381 0.000736842
R66576 DVSS.n925 DVSS.n910 0.000736842
R66577 DVSS.n22405 DVSS.n1005 0.000736842
R66578 DVSS.n18150 DVSS.n15545 0.000736842
R66579 DVSS.n22286 DVSS.n1255 0.000736842
R66580 DVSS.n12867 DVSS.n27 0.000736842
R66581 DVSS.n12899 DVSS.n12801 0.000736842
R66582 DVSS.n6671 DVSS.n6237 0.000734214
R66583 DVSS.n7104 DVSS.n7103 0.000734214
R66584 DVSS.n2012 DVSS.n1967 0.000734214
R66585 DVSS.n11643 DVSS.n11622 0.000734214
R66586 DVSS.n7078 DVSS.n5184 0.000729621
R66587 DVSS.n10116 DVSS.n2718 0.000729621
R66588 DVSS.n7827 DVSS.n7826 0.000725029
R66589 DVSS.n10127 DVSS.n10126 0.000725029
R66590 DVSS.n12761 DVSS.n12760 0.000725029
R66591 DVSS.n7105 DVSS.n7102 0.000720436
R66592 DVSS.n15812 DVSS.n15786 0.000719512
R66593 DVSS.n22372 DVSS.n22371 0.000719512
R66594 DVSS.n15739 DVSS.n15543 0.000719512
R66595 DVSS.n13063 DVSS.n12959 0.000719512
R66596 DVSS.n15857 DVSS.n15837 0.000719512
R66597 DVSS.n19002 DVSS.n13574 0.000719512
R66598 DVSS.n1026 DVSS.n1015 0.000719512
R66599 DVSS.n15704 DVSS.n15544 0.000719512
R66600 DVSS.n19181 DVSS.n13423 0.000719512
R66601 DVSS.n23003 DVSS.n384 0.000719512
R66602 DVSS.n4014 DVSS.n3858 0.000715844
R66603 DVSS.n18016 DVSS.n15552 0.000711268
R66604 DVSS.n13807 DVSS.n13731 0.00071
R66605 DVSS.n1494 DVSS.n976 0.00071
R66606 DVSS.n894 DVSS.n886 0.00071
R66607 DVSS.n1397 DVSS.n1365 0.00071
R66608 DVSS.n3460 DVSS.n3457 0.000706659
R66609 DVSS.n8970 DVSS.n8635 0.000706659
R66610 DVSS.n8091 DVSS.n8090 0.000697474
R66611 DVSS.n3045 DVSS.n2890 0.000697474
R66612 DVSS.n9759 DVSS.n9465 0.000692882
R66613 DVSS.n9771 DVSS.n2728 0.000692882
R66614 DVSS.n16755 DVSS.n15595 0.000692857
R66615 DVSS.n15524 DVSS.n15493 0.000692857
R66616 DVSS.n18267 DVSS.n18219 0.000692857
R66617 DVSS.n15119 DVSS.n15103 0.000692857
R66618 DVSS.n20960 DVSS.n14338 0.000692857
R66619 DVSS.n21414 DVSS.n13395 0.000692857
R66620 DVSS.n22860 DVSS.n473 0.000692857
R66621 DVSS.n8103 DVSS.n8102 0.000688289
R66622 DVSS.n8601 DVSS.n3460 0.000688289
R66623 DVSS.n9760 DVSS.n9759 0.000688289
R66624 DVSS.n9465 DVSS.n2781 0.000688289
R66625 DVSS DVSS.n17998 0.000687793
R66626 DVSS.n21103 DVSS.n21102 0.00068
R66627 DVSS.n14217 DVSS.n14187 0.00068
R66628 DVSS.n1122 DVSS.n285 0.00068
R66629 DVSS.n393 DVSS.n391 0.00068
R66630 DVSS DVSS.n417 0.00068
R66631 DVSS.n23086 DVSS.n253 0.00068
R66632 DVSS.n115 DVSS.n108 0.00068
R66633 DVSS.n21645 DVSS.n21636 0.00068
R66634 DVSS.n21959 DVSS.n21768 0.00068
R66635 DVSS DVSS.n22977 0.00068
R66636 DVSS.n8970 DVSS.n8969 0.000679104
R66637 DVSS.n8978 DVSS.n3052 0.000679104
R66638 DVSS.n10142 DVSS.n2364 0.000679104
R66639 DVSS.n13111 DVSS.n11994 0.000679104
R66640 DVSS.n4022 DVSS.n4015 0.000674512
R66641 DVSS.n13337 DVSS.n11156 0.000674512
R66642 DVSS.n22871 DVSS 0.000671429
R66643 DVSS DVSS.n16736 0.000671429
R66644 DVSS.n18184 DVSS 0.000671429
R66645 DVSS DVSS.n18245 0.000671429
R66646 DVSS.n19937 DVSS 0.000671429
R66647 DVSS.n20949 DVSS 0.000671429
R66648 DVSS.n21403 DVSS 0.000671429
R66649 DVSS.n6680 DVSS.n6679 0.00066992
R66650 DVSS.n7088 DVSS.n7087 0.00066992
R66651 DVSS.n10487 DVSS.n10486 0.00066992
R66652 DVSS.n13327 DVSS.n11458 0.00066992
R66653 DVSS.n7826 DVSS.n4471 0.000665327
R66654 DVSS.n1568 DVSS.n1523 0.000665327
R66655 DVSS.n5879 DVSS.n5867 0.000660735
R66656 DVSS.n5574 DVSS.n5525 0.000660735
R66657 DVSS.n7815 DVSS.n4811 0.000660735
R66658 DVSS.n1566 DVSS.n1511 0.000660735
R66659 DVSS.n11110 DVSS.n11109 0.000660735
R66660 DVSS.n9455 DVSS.n2787 0.000656142
R66661 DVSS.n7068 DVSS.n5182 0.00065155
R66662 DVSS.n7452 DVSS.n7451 0.00065155
R66663 DVSS.n10461 DVSS.n10460 0.00065155
R66664 DVSS.n11982 DVSS.n11981 0.00065155
R66665 DVSS.n21029 DVSS.n14257 0.00065
R66666 DVSS.n12784 DVSS.n12783 0.00065
R66667 DVSS.n29 DVSS.n4 0.00065
R66668 DVSS.n21986 DVSS.n1230 0.00065
R66669 DVSS.n2720 DVSS.n2719 0.000646958
R66670 DVSS.n12757 DVSS.n12359 0.000646958
R66671 DVSS.n12756 DVSS.n12506 0.000646958
R66672 DVSS.n12758 DVSS.n12360 0.000646958
R66673 DVSS.n12754 DVSS.n12553 0.000646958
R66674 DVSS.n12768 DVSS.n12361 0.000646958
R66675 DVSS.n4470 DVSS.n4469 0.000642365
R66676 DVSS.n2719 DVSS.n2706 0.000642365
R66677 DVSS.n19420 DVSS.n711 0.000642105
R66678 DVSS.n22145 DVSS.n22122 0.000642105
R66679 DVSS.n941 DVSS.n921 0.000642105
R66680 DVSS.n19763 DVSS.n465 0.000642105
R66681 DVSS.n22317 DVSS.n1240 0.000642105
R66682 DVSS.n12836 DVSS.n20 0.000642105
R66683 DVSS.n15867 DVSS.n15853 0.000640845
R66684 DVSS.n17928 DVSS.n15760 0.000640845
R66685 DVSS.n10167 DVSS.n10166 0.00063318
R66686 DVSS.n7034 DVSS.n5878 0.000628588
R66687 DVSS.n8320 DVSS.n3900 0.000628588
R66688 DVSS.n16323 DVSS.n16309 0.000628571
R66689 DVSS.n16700 DVSS.n16185 0.000628571
R66690 DVSS.n16048 DVSS.n16018 0.000628571
R66691 DVSS.n16865 DVSS.n16841 0.000628571
R66692 DVSS.n15276 DVSS.n15272 0.000628571
R66693 DVSS.n15409 DVSS.n15385 0.000628571
R66694 DVSS.n18415 DVSS.n18385 0.000628571
R66695 DVSS.n14971 DVSS.n14949 0.000628571
R66696 DVSS.n20786 DVSS.n20708 0.000628571
R66697 DVSS.n20869 DVSS.n14430 0.000628571
R66698 DVSS.n13607 DVSS.n13587 0.000628571
R66699 DVSS.n21319 DVSS.n13486 0.000628571
R66700 DVSS.n690 DVSS.n676 0.000628571
R66701 DVSS.n22777 DVSS.n570 0.000628571
R66702 DVSS.n14623 DVSS 0.000626404
R66703 DVSS.n8103 DVSS.n4021 0.000623995
R66704 DVSS.n8111 DVSS.n4022 0.000623995
R66705 DVSS.n8614 DVSS.n3406 0.000623995
R66706 DVSS.n8634 DVSS.n8633 0.000623995
R66707 DVSS.n8979 DVSS 0.000623995
R66708 DVSS.n13888 DVSS.n13861 0.00062
R66709 DVSS.n14116 DVSS.n14068 0.00062
R66710 DVSS.n1106 DVSS.n1067 0.00062
R66711 DVSS.n12973 DVSS.n311 0.00062
R66712 DVSS.n22472 DVSS.n801 0.00062
R66713 DVSS.n183 DVSS.n182 0.00062
R66714 DVSS.n21932 DVSS.n21870 0.00062
R66715 DVSS.n21750 DVSS.n21725 0.00062
R66716 DVSS.n6679 DVSS.n6231 0.000610218
R66717 DVSS.n6689 DVSS.n5888 0.000610218
R66718 DVSS.n3848 DVSS.n3799 0.000610218
R66719 DVSS.n8590 DVSS.n8588 0.000610218
R66720 DVSS.n8101 DVSS.n8100 0.000605626
R66721 DVSS.n8605 DVSS.n8604 0.000605626
R66722 DVSS.n9771 DVSS.n9770 0.000605626
R66723 DVSS.n10487 DVSS.n1961 0.000605626
R66724 DVSS.n10495 DVSS.n1620 0.000605626
R66725 DVSS.n3052 DVSS.n3046 0.000601033
R66726 DVSS.n2708 DVSS.n2415 0.000601033
R66727 DVSS.n7088 DVSS.n4886 0.000596441
R66728 DVSS.n7102 DVSS.n4840 0.000596441
R66729 DVSS.n7807 DVSS.n4818 0.000596441
R66730 DVSS.n10152 DVSS.n10151 0.000596441
R66731 DVSS.n13341 DVSS.n13340 0.000596441
R66732 DVSS.n12338 DVSS.n11631 0.000596441
R66733 DVSS.n12338 DVSS.n12337 0.000596441
R66734 DVSS.n21043 DVSS.n14253 0.00059
R66735 DVSS.n12779 DVSS.n411 0.00059
R66736 DVSS.n48 DVSS.n33 0.00059
R66737 DVSS.n21977 DVSS.n1226 0.00059
R66738 DVSS.n6689 DVSS.n6688 0.000587256
R66739 DVSS.n5183 DVSS.n5176 0.000587256
R66740 DVSS.n8588 DVSS.n3755 0.000587256
R66741 DVSS.n10498 DVSS.n10495 0.000587256
R66742 DVSS.n11457 DVSS.n11198 0.000587256
R66743 DVSS.n7060 DVSS.n7059 0.000582664
R66744 DVSS.n7818 DVSS.n4468 0.000582664
R66745 DVSS.n10754 DVSS.n1566 0.000582664
R66746 DVSS DVSS.n21982 0.00058
R66747 DVSS DVSS.n14305 0.00058
R66748 DVSS.n7034 DVSS.n7033 0.000578071
R66749 DVSS.n7069 DVSS.n7068 0.000578071
R66750 DVSS.n10755 DVSS.n1523 0.000578071
R66751 DVSS.n13341 DVSS.n11111 0.000578071
R66752 DVSS.n11982 DVSS.n11646 0.000578071
R66753 DVSS.n11980 DVSS.n11630 0.000578071
R66754 DVSS.n9188 DVSS.n9187 0.000573479
R66755 DVSS.n9199 DVSS.n2831 0.000573479
R66756 DVSS.n7461 DVSS.n7460 0.000568886
R66757 DVSS.n2070 DVSS.n2019 0.000568886
R66758 DVSS.n13122 DVSS.n11630 0.000568886
R66759 DVSS.n7795 DVSS.n4818 0.000564294
R66760 DVSS.n13349 DVSS.n10766 0.000564294
R66761 DVSS.n13906 DVSS.n13876 0.00056
R66762 DVSS.n14100 DVSS.n14072 0.00056
R66763 DVSS.n1475 DVSS.n1056 0.00056
R66764 DVSS.n12977 DVSS.n302 0.00056
R66765 DVSS.n22475 DVSS.n792 0.00056
R66766 DVSS.n193 DVSS.n163 0.00056
R66767 DVSS.n21855 DVSS.n1445 0.00056
R66768 DVSS.n21737 DVSS.n21729 0.00056
R66769 DVSS.n8091 DVSS.n4371 0.000559702
R66770 DVSS.n8969 DVSS 0.000559702
R66771 DVSS.n2880 DVSS.n2831 0.000559702
R66772 DVSS.n9457 DVSS.n9455 0.000559702
R66773 DVSS.n10116 DVSS.n10115 0.000559702
R66774 DVSS.n9198 DVSS.n2878 0.000550517
R66775 DVSS.n10151 DVSS.n2073 0.000550517
R66776 DVSS.n956 DVSS.n908 0.000547368
R66777 DVSS.n22389 DVSS.n1007 0.000547368
R66778 DVSS.n12851 DVSS.n9 0.000547368
R66779 DVSS.n12883 DVSS.n12810 0.000547368
R66780 DVSS.n5880 DVSS.n5879 0.000545924
R66781 DVSS.n8317 DVSS.n3946 0.000545924
R66782 DVSS.n8616 DVSS.n8615 0.000541332
R66783 DVSS.n8625 DVSS.n8624 0.000541332
R66784 DVSS.n9187 DVSS.n2932 0.000541332
R66785 DVSS.n9184 DVSS.n2937 0.000541332
R66786 DVSS.n13327 DVSS.n13326 0.000541332
R66787 DVSS.n13323 DVSS.n11504 0.000541332
R66788 DVSS.n6654 DVSS.n6257 0.000536739
R66789 DVSS.n6652 DVSS.n6258 0.000536739
R66790 DVSS.n6602 DVSS.n6256 0.000536739
R66791 DVSS.n6661 DVSS.n6259 0.000536739
R66792 DVSS.n6657 DVSS.n6656 0.000536739
R66793 DVSS.n8331 DVSS.n3846 0.000532147
R66794 DVSS.n2937 DVSS.n2936 0.000532147
R66795 DVSS.n7452 DVSS.n4832 0.000522962
R66796 DVSS.n7460 DVSS.n4825 0.000522962
R66797 DVSS.n7836 DVSS.n4413 0.000522962
R66798 DVSS.n2730 DVSS.n2729 0.000522962
R66799 DVSS.n7806 DVSS.n4811 0.00051837
R66800 DVSS.n10143 DVSS.n10141 0.00051837
R66801 DVSS.n10765 DVSS.n1512 0.00051837
R66802 DVSS.n7797 DVSS.n7796 0.000513777
R66803 DVSS.n10167 DVSS.n2027 0.000513777
R66804 DVSS.n10461 DVSS.n2013 0.000513777
R66805 DVSS.n10475 DVSS.n1967 0.000513777
R66806 DVSS.n13121 DVSS.n13120 0.000513777
R66807 DVSS.n12336 DVSS.n11994 0.000513777
R66808 DVSS.n5890 DVSS.n5889 0.000504592
R66809 DVSS.n7079 DVSS.n7078 0.000504592
R66810 DVSS.n8321 DVSS.n8320 0.000504592
R66811 DVSS.n8317 DVSS.n3904 0.000504592
R66812 DVSS.n8332 DVSS.n3799 0.000504592
R66813 DVSS.n10497 DVSS.n10496 0.000504592
R66814 DVSS.n11156 DVSS.n11153 0.000504592
R66815 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_1.D.n17 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_1.D.t12 47.1029
R66816 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_1.D.n6 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_1.D.t31 47.1029
R66817 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_1.D.n4 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_1.D.t15 47.1029
R66818 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_1.D.n2 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_1.D.t26 47.1029
R66819 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_1.D.n17 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_1.D.t11 38.0648
R66820 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_1.D.n18 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_1.D.t20 38.0648
R66821 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_1.D.n19 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_1.D.t9 38.0648
R66822 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_1.D.n20 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_1.D.t32 38.0648
R66823 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_1.D.n21 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_1.D.t24 38.0648
R66824 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_1.D.n22 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_1.D.t18 38.0648
R66825 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_1.D.n23 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_1.D.t30 38.0648
R66826 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_1.D.n24 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_1.D.t29 38.0648
R66827 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_1.D.n25 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_1.D.t10 38.0648
R66828 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_1.D.n26 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_1.D.t6 38.0648
R66829 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_1.D.n27 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_1.D.t27 38.0648
R66830 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_1.D.n6 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_1.D.t16 38.0648
R66831 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_1.D.n7 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_1.D.t25 38.0648
R66832 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_1.D.n8 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_1.D.t33 38.0648
R66833 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_1.D.n9 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_1.D.t13 38.0648
R66834 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_1.D.n10 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_1.D.t19 38.0648
R66835 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_1.D.n11 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_1.D.t28 38.0648
R66836 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_1.D.n12 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_1.D.t5 38.0648
R66837 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_1.D.n13 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_1.D.t17 38.0648
R66838 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_1.D.n14 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_1.D.t21 38.0648
R66839 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_1.D.n15 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_1.D.t7 38.0648
R66840 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_1.D.n16 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_1.D.t8 38.0648
R66841 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_1.D.n4 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_1.D.t14 38.0648
R66842 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_1.D.n5 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_1.D.t23 38.0648
R66843 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_1.D.n2 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_1.D.t4 38.0648
R66844 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_1.D.n3 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_1.D.t22 38.0648
R66845 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_1.D.n18 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_1.D.n17 9.0386
R66846 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_1.D.n19 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_1.D.n18 9.0386
R66847 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_1.D.n20 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_1.D.n19 9.0386
R66848 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_1.D.n21 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_1.D.n20 9.0386
R66849 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_1.D.n22 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_1.D.n21 9.0386
R66850 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_1.D.n23 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_1.D.n22 9.0386
R66851 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_1.D.n24 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_1.D.n23 9.0386
R66852 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_1.D.n25 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_1.D.n24 9.0386
R66853 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_1.D.n26 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_1.D.n25 9.0386
R66854 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_1.D.n27 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_1.D.n26 9.0386
R66855 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_1.D.n7 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_1.D.n6 9.0386
R66856 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_1.D.n8 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_1.D.n7 9.0386
R66857 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_1.D.n9 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_1.D.n8 9.0386
R66858 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_1.D.n10 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_1.D.n9 9.0386
R66859 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_1.D.n11 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_1.D.n10 9.0386
R66860 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_1.D.n12 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_1.D.n11 9.0386
R66861 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_1.D.n13 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_1.D.n12 9.0386
R66862 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_1.D.n14 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_1.D.n13 9.0386
R66863 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_1.D.n15 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_1.D.n14 9.0386
R66864 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_1.D.n16 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_1.D.n15 9.0386
R66865 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_1.D.n5 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_1.D.n4 9.0386
R66866 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_1.D.n3 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_1.D.n2 9.0386
R66867 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_1.D.n1 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_1.D.n16 4.51955
R66868 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_1.D.n1 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_1.D.n27 4.51955
R66869 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_1.D.n0 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_1.D.n3 4.51955
R66870 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_1.D.n0 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_1.D.n5 4.51955
R66871 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_1.D.n1 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_1.D.t3 2.87695
R66872 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_1.D.n1 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_1.D.n0 2.37212
R66873 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_1.D.t0 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_1.D.t1 1.95734
R66874 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_1.D.t3 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_1.D.t2 1.87633
R66875 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_1.D.t0 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_1.D.n1 1.56603
R66876 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531459_0.D.n3 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531459_0.D.t4 47.1029
R66877 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531459_0.D.n1 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531459_0.D.t9 47.1029
R66878 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531459_0.D.n6 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531459_0.D.t7 47.1029
R66879 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531459_0.D.n6 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531459_0.D.t11 47.1029
R66880 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531459_0.D.n3 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531459_0.D.t3 38.0648
R66881 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531459_0.D.n4 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531459_0.D.t8 38.0648
R66882 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531459_0.D.n1 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531459_0.D.t10 38.0648
R66883 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531459_0.D.n2 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531459_0.D.t5 38.0648
R66884 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531459_0.D.n6 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531459_0.D.t6 38.0648
R66885 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531459_0.D.n4 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531459_0.D.n3 9.0386
R66886 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531459_0.D.n2 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531459_0.D.n1 9.0386
R66887 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531459_0.D.n5 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531459_0.D.n2 4.51955
R66888 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531459_0.D.n5 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531459_0.D.n4 4.51955
R66889 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531459_0.D.n0 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531459_0.D.t2 2.8466
R66890 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531459_0.D.n0 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531459_0.D.n5 2.40746
R66891 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531459_0.D.n0 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531459_0.D.t0 1.87633
R66892 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531459_0.D.n0 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531459_0.D.n6 1.76725
R66893 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531459_0.D.n0 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531459_0.D.t1 1.65385
R66894 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/comp018green_esd_rc_v5p0_0.ppolyf_u_CDNS_406619531453_2.MINUS GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/comp018green_esd_rc_v5p0_0.ppolyf_u_CDNS_406619531453_2.MINUS.t0 11.0117
R66895 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/comp018green_esd_rc_v5p0_0.ppolyf_u_CDNS_406619531453_2.MINUS GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/comp018green_esd_rc_v5p0_0.ppolyf_u_CDNS_406619531453_2.MINUS.t1 11.0117
R66896 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/comp018green_esd_rc_v5p0_0.ppolyf_u_CDNS_406619531453_2.PLUS.t0 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/comp018green_esd_rc_v5p0_0.ppolyf_u_CDNS_406619531453_2.PLUS.t1 22.3936
R66897 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/comp018green_esd_rc_v5p0_0.VRC GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/comp018green_esd_rc_v5p0_0.VRC.t0 11.0117
R66898 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/comp018green_esd_rc_v5p0_0.VRC GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/comp018green_esd_rc_v5p0_0.VRC.n12 0.6125
R66899 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/comp018green_esd_rc_v5p0_0.VRC.n12 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/comp018green_esd_rc_v5p0_0.VRC.n18 1.2266
R66900 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/comp018green_esd_rc_v5p0_0.VRC.n19 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/comp018green_esd_rc_v5p0_0.VRC 0.225727
R66901 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/comp018green_esd_rc_v5p0_0.VRC GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/comp018green_esd_rc_v5p0_0.VRC.n18 0.00644
R66902 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/comp018green_esd_rc_v5p0_0.VRC.t9 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/comp018green_esd_rc_v5p0_0.VRC.n19 4.75334
R66903 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/comp018green_esd_rc_v5p0_0.VRC GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/comp018green_esd_rc_v5p0_0.VRC.n19 0.225727
R66904 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/comp018green_esd_rc_v5p0_0.VRC.n18 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/comp018green_esd_rc_v5p0_0.VRC.n16 0.767246
R66905 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/comp018green_esd_rc_v5p0_0.VRC.n17 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/comp018green_esd_rc_v5p0_0.VRC 0.225727
R66906 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/comp018green_esd_rc_v5p0_0.VRC GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/comp018green_esd_rc_v5p0_0.VRC.n16 0.00644
R66907 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/comp018green_esd_rc_v5p0_0.VRC.t8 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/comp018green_esd_rc_v5p0_0.VRC.n17 4.75334
R66908 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/comp018green_esd_rc_v5p0_0.VRC GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/comp018green_esd_rc_v5p0_0.VRC.n17 0.225727
R66909 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/comp018green_esd_rc_v5p0_0.VRC.n16 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/comp018green_esd_rc_v5p0_0.VRC.n14 0.767246
R66910 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/comp018green_esd_rc_v5p0_0.VRC.n15 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/comp018green_esd_rc_v5p0_0.VRC 0.225727
R66911 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/comp018green_esd_rc_v5p0_0.VRC GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/comp018green_esd_rc_v5p0_0.VRC.n14 0.00644
R66912 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/comp018green_esd_rc_v5p0_0.VRC.t13 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/comp018green_esd_rc_v5p0_0.VRC.n15 4.75334
R66913 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/comp018green_esd_rc_v5p0_0.VRC GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/comp018green_esd_rc_v5p0_0.VRC.n15 0.225727
R66914 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/comp018green_esd_rc_v5p0_0.VRC.n13 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/comp018green_esd_rc_v5p0_0.VRC 0.225727
R66915 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/comp018green_esd_rc_v5p0_0.VRC GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/comp018green_esd_rc_v5p0_0.VRC.n14 0.773185
R66916 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/comp018green_esd_rc_v5p0_0.VRC.t10 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/comp018green_esd_rc_v5p0_0.VRC.n13 4.75334
R66917 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/comp018green_esd_rc_v5p0_0.VRC GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/comp018green_esd_rc_v5p0_0.VRC.n13 0.225727
R66918 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/comp018green_esd_rc_v5p0_0.VRC.n12 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/comp018green_esd_rc_v5p0_0.VRC.n4 6.26225
R66919 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/comp018green_esd_rc_v5p0_0.VRC.n4 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/comp018green_esd_rc_v5p0_0.VRC 0.332722
R66920 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/comp018green_esd_rc_v5p0_0.VRC GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/comp018green_esd_rc_v5p0_0.VRC.n10 0.894378
R66921 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/comp018green_esd_rc_v5p0_0.VRC.n10 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/comp018green_esd_rc_v5p0_0.VRC 0.00644
R66922 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/comp018green_esd_rc_v5p0_0.VRC.n11 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/comp018green_esd_rc_v5p0_0.VRC 0.225727
R66923 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/comp018green_esd_rc_v5p0_0.VRC.t5 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/comp018green_esd_rc_v5p0_0.VRC.n11 4.75334
R66924 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/comp018green_esd_rc_v5p0_0.VRC GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/comp018green_esd_rc_v5p0_0.VRC.n11 0.225727
R66925 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/comp018green_esd_rc_v5p0_0.VRC.n10 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/comp018green_esd_rc_v5p0_0.VRC.n8 0.767246
R66926 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/comp018green_esd_rc_v5p0_0.VRC.n8 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/comp018green_esd_rc_v5p0_0.VRC 0.00644
R66927 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/comp018green_esd_rc_v5p0_0.VRC.n9 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/comp018green_esd_rc_v5p0_0.VRC 0.225727
R66928 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/comp018green_esd_rc_v5p0_0.VRC.t4 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/comp018green_esd_rc_v5p0_0.VRC.n9 4.75334
R66929 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/comp018green_esd_rc_v5p0_0.VRC GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/comp018green_esd_rc_v5p0_0.VRC.n9 0.225727
R66930 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/comp018green_esd_rc_v5p0_0.VRC.n8 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/comp018green_esd_rc_v5p0_0.VRC.n6 0.767246
R66931 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/comp018green_esd_rc_v5p0_0.VRC.n6 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/comp018green_esd_rc_v5p0_0.VRC 0.00644
R66932 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/comp018green_esd_rc_v5p0_0.VRC.n7 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/comp018green_esd_rc_v5p0_0.VRC 0.225727
R66933 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/comp018green_esd_rc_v5p0_0.VRC.t7 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/comp018green_esd_rc_v5p0_0.VRC.n7 4.75334
R66934 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/comp018green_esd_rc_v5p0_0.VRC GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/comp018green_esd_rc_v5p0_0.VRC.n7 0.225727
R66935 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/comp018green_esd_rc_v5p0_0.VRC.n6 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/comp018green_esd_rc_v5p0_0.VRC 0.773185
R66936 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/comp018green_esd_rc_v5p0_0.VRC.n5 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/comp018green_esd_rc_v5p0_0.VRC 0.225727
R66937 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/comp018green_esd_rc_v5p0_0.VRC.t6 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/comp018green_esd_rc_v5p0_0.VRC.n5 4.75334
R66938 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/comp018green_esd_rc_v5p0_0.VRC GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/comp018green_esd_rc_v5p0_0.VRC.n5 0.225727
R66939 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/comp018green_esd_rc_v5p0_0.VRC.n3 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/comp018green_esd_rc_v5p0_0.VRC.n2 1.0005
R66940 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/comp018green_esd_rc_v5p0_0.VRC.n4 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/comp018green_esd_rc_v5p0_0.VRC.n3 2.62726
R66941 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/comp018green_esd_rc_v5p0_0.VRC.n3 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/comp018green_esd_rc_v5p0_0.VRC.t3 36.8287
R66942 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/comp018green_esd_rc_v5p0_0.VRC.n2 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/comp018green_esd_rc_v5p0_0.VRC.n0 4.51955
R66943 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/comp018green_esd_rc_v5p0_0.VRC.n2 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/comp018green_esd_rc_v5p0_0.VRC.n1 4.51955
R66944 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/comp018green_esd_rc_v5p0_0.VRC.n1 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/comp018green_esd_rc_v5p0_0.VRC.t2 38.0648
R66945 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/comp018green_esd_rc_v5p0_0.VRC.n1 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/comp018green_esd_rc_v5p0_0.VRC.t1 47.1029
R66946 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/comp018green_esd_rc_v5p0_0.VRC.n0 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/comp018green_esd_rc_v5p0_0.VRC.t11 38.0648
R66947 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/comp018green_esd_rc_v5p0_0.VRC.n0 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/comp018green_esd_rc_v5p0_0.VRC.t12 47.1029
R66948 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/comp018green_esd_rc_v5p0_0.ppolyf_u_CDNS_406619531453_4.PLUS.t0 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/comp018green_esd_rc_v5p0_0.ppolyf_u_CDNS_406619531453_4.PLUS.t1 22.3936
R66949 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/comp018green_esd_rc_v5p0_0.ppolyf_u_CDNS_406619531453_1.MINUS.t0 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/comp018green_esd_rc_v5p0_0.ppolyf_u_CDNS_406619531453_1.MINUS.t1 22.3936
R66950 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/comp018green_esd_rc_v5p0_0.ppolyf_u_CDNS_406619531453_0.PLUS.t0 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/comp018green_esd_rc_v5p0_0.ppolyf_u_CDNS_406619531453_0.PLUS 11.0117
R66951 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/comp018green_esd_rc_v5p0_0.ppolyf_u_CDNS_406619531453_0.PLUS GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/comp018green_esd_rc_v5p0_0.ppolyf_u_CDNS_406619531453_0.PLUS.t1 11.0117
R66952 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/comp018green_esd_rc_v5p0_0.ppolyf_u_CDNS_406619531453_3.PLUS.t0 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/comp018green_esd_rc_v5p0_0.ppolyf_u_CDNS_406619531453_3.PLUS 11.0117
R66953 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/comp018green_esd_rc_v5p0_0.ppolyf_u_CDNS_406619531453_3.PLUS GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/comp018green_esd_rc_v5p0_0.ppolyf_u_CDNS_406619531453_3.PLUS.t1 11.0117
R66954 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/comp018green_esd_rc_v5p0_0.ppolyf_u_CDNS_406619531453_3.MINUS GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/comp018green_esd_rc_v5p0_0.ppolyf_u_CDNS_406619531453_3.MINUS.t0 11.0117
R66955 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/comp018green_esd_rc_v5p0_0.ppolyf_u_CDNS_406619531453_3.MINUS GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/comp018green_esd_rc_v5p0_0.ppolyf_u_CDNS_406619531453_3.MINUS.t1 11.0117
R66956 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/comp018green_esd_rc_v5p0_0.ppolyf_u_CDNS_406619531453_4.MINUS GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/comp018green_esd_rc_v5p0_0.ppolyf_u_CDNS_406619531453_4.MINUS.t0 11.0117
R66957 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/comp018green_esd_rc_v5p0_0.ppolyf_u_CDNS_406619531453_4.MINUS GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/comp018green_esd_rc_v5p0_0.ppolyf_u_CDNS_406619531453_4.MINUS.t1 11.0117
R66958 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/comp018green_esd_rc_v5p0_0.ppolyf_u_CDNS_406619531453_1.PLUS.t0 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/comp018green_esd_rc_v5p0_0.ppolyf_u_CDNS_406619531453_1.PLUS.t1 22.3936
R66959 VDD.n48 VDD.n47 13.4781
R66960 VDD.n44 VDD.n13 0.4505
R66961 VDD.n43 VDD.n15 0.4505
R66962 VDD.n18 VDD.n14 0.4505
R66963 VDD.n39 VDD.n38 0.4505
R66964 VDD.n37 VDD.n17 0.4505
R66965 VDD.n36 VDD.n35 0.4505
R66966 VDD.n20 VDD.n19 0.4505
R66967 VDD.n31 VDD.n30 0.4505
R66968 VDD.n29 VDD.n22 0.4505
R66969 VDD.n28 VDD.n27 0.4505
R66970 VDD.n24 VDD.n23 0.4505
R66971 VDD.n52 VDD.n51 0.4505
R66972 VDD.n53 VDD.n8 0.4505
R66973 VDD.n55 VDD.n54 0.4505
R66974 VDD.n6 VDD.n5 0.4505
R66975 VDD.n60 VDD.n59 0.4505
R66976 VDD.n61 VDD.n4 0.4505
R66977 VDD.n64 VDD.n63 0.4505
R66978 VDD.n62 VDD.n2 0.4505
R66979 VDD.n68 VDD.n1 0.4505
R66980 VDD.n70 VDD.n69 0.4505
R66981 VDD.n72 VDD.n71 0.4505
R66982 VDD.n51 VDD.n50 0.4505
R66983 VDD.n8 VDD.n7 0.4505
R66984 VDD.n56 VDD.n55 0.4505
R66985 VDD.n57 VDD.n6 0.4505
R66986 VDD.n59 VDD.n58 0.4505
R66987 VDD.n4 VDD.n3 0.4505
R66988 VDD.n65 VDD.n64 0.4505
R66989 VDD.n66 VDD.n2 0.4505
R66990 VDD.n68 VDD.n67 0.4505
R66991 VDD.n69 VDD.n0 0.4505
R66992 VDD.n49 VDD.n10 0.4505
R66993 VDD.n44 VDD.n12 0.4505
R66994 VDD.n43 VDD.n42 0.4505
R66995 VDD.n41 VDD.n14 0.4505
R66996 VDD.n40 VDD.n39 0.4505
R66997 VDD.n17 VDD.n16 0.4505
R66998 VDD.n35 VDD.n34 0.4505
R66999 VDD.n33 VDD.n20 0.4505
R67000 VDD.n32 VDD.n31 0.4505
R67001 VDD.n22 VDD.n21 0.4505
R67002 VDD.n27 VDD.n26 0.4505
R67003 VDD.n46 VDD.n45 0.4505
R67004 VDD.n73 VDD 0.130161
R67005 VDD.n25 VDD 0.130161
R67006 VDD VDD.n73 0.101206
R67007 VDD VDD.n25 0.101206
R67008 VDD.n48 VDD.n9 0.0737595
R67009 VDD.n47 VDD.n11 0.0737595
R67010 VDD.n13 VDD.n11 0.0585093
R67011 VDD.n52 VDD.n9 0.0585093
R67012 VDD.n45 VDD.n11 0.0267299
R67013 VDD.n10 VDD.n9 0.0267299
R67014 VDD.n25 VDD.n24 0.0142814
R67015 VDD.n73 VDD.n72 0.0142814
R67016 VDD.n45 VDD.n44 0.00962857
R67017 VDD.n44 VDD.n43 0.00962857
R67018 VDD.n43 VDD.n14 0.00962857
R67019 VDD.n39 VDD.n14 0.00962857
R67020 VDD.n39 VDD.n17 0.00962857
R67021 VDD.n35 VDD.n17 0.00962857
R67022 VDD.n35 VDD.n20 0.00962857
R67023 VDD.n31 VDD.n20 0.00962857
R67024 VDD.n31 VDD.n22 0.00962857
R67025 VDD.n27 VDD.n22 0.00962857
R67026 VDD.n51 VDD.n10 0.00962857
R67027 VDD.n51 VDD.n8 0.00962857
R67028 VDD.n55 VDD.n8 0.00962857
R67029 VDD.n55 VDD.n6 0.00962857
R67030 VDD.n59 VDD.n6 0.00962857
R67031 VDD.n59 VDD.n4 0.00962857
R67032 VDD.n64 VDD.n4 0.00962857
R67033 VDD.n64 VDD.n2 0.00962857
R67034 VDD.n68 VDD.n2 0.00962857
R67035 VDD.n69 VDD.n68 0.00962857
R67036 VDD.n50 VDD.n49 0.00962857
R67037 VDD.n50 VDD.n7 0.00962857
R67038 VDD.n56 VDD.n7 0.00962857
R67039 VDD.n57 VDD.n56 0.00962857
R67040 VDD.n58 VDD.n57 0.00962857
R67041 VDD.n58 VDD.n3 0.00962857
R67042 VDD.n65 VDD.n3 0.00962857
R67043 VDD.n66 VDD.n65 0.00962857
R67044 VDD.n67 VDD.n66 0.00962857
R67045 VDD.n67 VDD.n0 0.00962857
R67046 VDD.n46 VDD.n12 0.00962857
R67047 VDD.n42 VDD.n12 0.00962857
R67048 VDD.n42 VDD.n41 0.00962857
R67049 VDD.n41 VDD.n40 0.00962857
R67050 VDD.n40 VDD.n16 0.00962857
R67051 VDD.n34 VDD.n16 0.00962857
R67052 VDD.n34 VDD.n33 0.00962857
R67053 VDD.n33 VDD.n32 0.00962857
R67054 VDD.n32 VDD.n21 0.00962857
R67055 VDD.n26 VDD.n21 0.00962857
R67056 VDD.n27 VDD 0.00782857
R67057 VDD.n69 VDD 0.00782857
R67058 VDD VDD.n0 0.00782857
R67059 VDD.n26 VDD 0.00782857
R67060 VDD.n15 VDD.n13 0.00658571
R67061 VDD.n18 VDD.n15 0.00658571
R67062 VDD.n38 VDD.n18 0.00658571
R67063 VDD.n38 VDD.n37 0.00658571
R67064 VDD.n37 VDD.n36 0.00658571
R67065 VDD.n36 VDD.n19 0.00658571
R67066 VDD.n30 VDD.n19 0.00658571
R67067 VDD.n30 VDD.n29 0.00658571
R67068 VDD.n29 VDD.n28 0.00658571
R67069 VDD.n28 VDD.n23 0.00658571
R67070 VDD.n53 VDD.n52 0.00658571
R67071 VDD.n54 VDD.n53 0.00658571
R67072 VDD.n54 VDD.n5 0.00658571
R67073 VDD.n60 VDD.n5 0.00658571
R67074 VDD.n61 VDD.n60 0.00658571
R67075 VDD.n63 VDD.n61 0.00658571
R67076 VDD.n63 VDD.n62 0.00658571
R67077 VDD.n62 VDD.n1 0.00658571
R67078 VDD.n70 VDD.n1 0.00658571
R67079 VDD VDD.n70 0.00538571
R67080 VDD.n24 VDD 0.0023
R67081 VDD.n72 VDD 0.0023
R67082 VDD.n49 VDD.n48 0.00191429
R67083 VDD.n47 VDD.n46 0.00191429
R67084 VDD.n71 VDD 0.0017
R67085 VDD VDD.n23 0.000671429
R67086 VDD.n71 VDD 0.000671429
C0 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/comp018green_esd_rc_v5p0_0.ppolyf_u_CDNS_406619531453_2.MINUS GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/comp018green_esd_rc_v5p0_0.ppolyf_u_CDNS_406619531453_4.MINUS 0.034604f
C1 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/comp018green_esd_rc_v5p0_0.ppolyf_u_CDNS_406619531453_4.MINUS DVDD 0.365886f
C2 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/comp018green_esd_rc_v5p0_0.ppolyf_u_CDNS_406619531453_4.MINUS VDD 3.57e-19
C3 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/comp018green_esd_rc_v5p0_0.ppolyf_u_CDNS_406619531453_5.MINUS GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/comp018green_esd_rc_v5p0_0.VRC 1.19e-19
C4 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/comp018green_esd_rc_v5p0_0.ppolyf_u_CDNS_406619531453_5.MINUS DVDD 0.365689f
C5 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/comp018green_esd_rc_v5p0_0.ppolyf_u_CDNS_406619531453_0.PLUS DVDD 0.39484f
C6 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/comp018green_esd_rc_v5p0_0.ppolyf_u_CDNS_406619531453_5.MINUS VDD 3.57e-19
C7 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/comp018green_esd_rc_v5p0_0.ppolyf_u_CDNS_406619531453_4.MINUS GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/comp018green_esd_rc_v5p0_0.ppolyf_u_CDNS_406619531453_5.MINUS 0.034604f
C8 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/comp018green_esd_rc_v5p0_0.ppolyf_u_CDNS_406619531453_3.MINUS GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/comp018green_esd_rc_v5p0_0.VRC 3.97e-19
C9 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/comp018green_esd_rc_v5p0_0.ppolyf_u_CDNS_406619531453_3.MINUS DVDD 0.367095f
C10 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/comp018green_esd_rc_v5p0_0.ppolyf_u_CDNS_406619531453_3.MINUS VDD 3.57e-19
C11 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/comp018green_esd_rc_v5p0_0.VRC GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D 0.003635f
C12 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D DVDD 0.140423p
C13 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/comp018green_esd_rc_v5p0_0.ppolyf_u_CDNS_406619531453_5.MINUS GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/comp018green_esd_rc_v5p0_0.ppolyf_u_CDNS_406619531453_3.MINUS 0.034604f
C14 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/comp018green_esd_rc_v5p0_0.ppolyf_u_CDNS_406619531453_2.MINUS DVDD 0.401222f
C15 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/comp018green_esd_rc_v5p0_0.ppolyf_u_CDNS_406619531453_3.PLUS DVDD 0.367212f
C16 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/comp018green_esd_rc_v5p0_0.ppolyf_u_CDNS_406619531453_2.MINUS VDD 3.57e-19
C17 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/comp018green_esd_rc_v5p0_0.VRC DVDD 5.07478f
C18 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/comp018green_esd_rc_v5p0_0.VRC VDD 0.186557f
C19 DVDD VDD 29.6195f
C20 VDD DVSS 0.120571p
C21 DVDD DVSS 2.019451p
C22 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D DVSS 0.371754p
C23 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/comp018green_esd_rc_v5p0_0.VRC DVSS 0.197185p
C24 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/comp018green_esd_rc_v5p0_0.ppolyf_u_CDNS_406619531453_0.PLUS DVSS 0.335584f
C25 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/comp018green_esd_rc_v5p0_0.ppolyf_u_CDNS_406619531453_3.MINUS DVSS 0.327749f
C26 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/comp018green_esd_rc_v5p0_0.ppolyf_u_CDNS_406619531453_3.PLUS DVSS 0.328934f
C27 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/comp018green_esd_rc_v5p0_0.ppolyf_u_CDNS_406619531453_5.MINUS DVSS 0.330163f
C28 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/comp018green_esd_rc_v5p0_0.ppolyf_u_CDNS_406619531453_4.MINUS DVSS 0.330163f
C29 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/comp018green_esd_rc_v5p0_0.ppolyf_u_CDNS_406619531453_2.MINUS DVSS 0.328845f
C30 VDD.n0 DVSS 0.04178f
C31 VDD.n1 DVSS 0.04635f
C32 VDD.n2 DVSS 0.04635f
C33 VDD.n3 DVSS 0.04635f
C34 VDD.n4 DVSS 0.04635f
C35 VDD.n5 DVSS 0.04635f
C36 VDD.n6 DVSS 0.04635f
C37 VDD.n7 DVSS 0.04635f
C38 VDD.n8 DVSS 0.04635f
C39 VDD.n9 DVSS 6.10826f
C40 VDD.n10 DVSS 0.157676f
C41 VDD.n11 DVSS 6.10826f
C42 VDD.n12 DVSS 0.04635f
C43 VDD.n13 DVSS 3.50137f
C44 VDD.n14 DVSS 0.04635f
C45 VDD.n15 DVSS 0.04635f
C46 VDD.n16 DVSS 0.04635f
C47 VDD.n17 DVSS 0.04635f
C48 VDD.n18 DVSS 0.04635f
C49 VDD.n19 DVSS 0.04635f
C50 VDD.n20 DVSS 0.04635f
C51 VDD.n21 DVSS 0.04635f
C52 VDD.n22 DVSS 0.04635f
C53 VDD.n23 DVSS 0.023828f
C54 VDD.n24 DVSS 0.061015f
C55 VDD.n25 DVSS 0.223333f
C56 VDD.n26 DVSS 0.04178f
C57 VDD.n27 DVSS 0.04178f
C58 VDD.n28 DVSS 0.04635f
C59 VDD.n29 DVSS 0.04635f
C60 VDD.n30 DVSS 0.04635f
C61 VDD.n31 DVSS 0.04635f
C62 VDD.n32 DVSS 0.04635f
C63 VDD.n33 DVSS 0.04635f
C64 VDD.n34 DVSS 0.04635f
C65 VDD.n35 DVSS 0.04635f
C66 VDD.n36 DVSS 0.04635f
C67 VDD.n37 DVSS 0.04635f
C68 VDD.n38 DVSS 0.04635f
C69 VDD.n39 DVSS 0.04635f
C70 VDD.n40 DVSS 0.04635f
C71 VDD.n41 DVSS 0.04635f
C72 VDD.n42 DVSS 0.04635f
C73 VDD.n43 DVSS 0.04635f
C74 VDD.n44 DVSS 0.04635f
C75 VDD.n45 DVSS 0.157676f
C76 VDD.n46 DVSS 0.026765f
C77 VDD.n47 DVSS 2.85102f
C78 VDD.n48 DVSS 2.85093f
C79 VDD.n49 DVSS 0.026765f
C80 VDD.n50 DVSS 0.04635f
C81 VDD.n51 DVSS 0.04635f
C82 VDD.n52 DVSS 3.50137f
C83 VDD.n53 DVSS 0.04635f
C84 VDD.n54 DVSS 0.04635f
C85 VDD.n55 DVSS 0.04635f
C86 VDD.n56 DVSS 0.04635f
C87 VDD.n57 DVSS 0.04635f
C88 VDD.n58 DVSS 0.04635f
C89 VDD.n59 DVSS 0.04635f
C90 VDD.n60 DVSS 0.04635f
C91 VDD.n61 DVSS 0.04635f
C92 VDD.n62 DVSS 0.04635f
C93 VDD.n63 DVSS 0.04635f
C94 VDD.n64 DVSS 0.04635f
C95 VDD.n65 DVSS 0.04635f
C96 VDD.n66 DVSS 0.04635f
C97 VDD.n67 DVSS 0.04635f
C98 VDD.n68 DVSS 0.04635f
C99 VDD.n69 DVSS 0.04178f
C100 VDD.n70 DVSS 0.04178f
C101 VDD.n71 DVSS 0.005223f
C102 VDD.n72 DVSS 0.061015f
C103 VDD.n73 DVSS 0.223333f
C104 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/comp018green_esd_rc_v5p0_0.VRC.t0 DVSS 7.51e-19
C105 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/comp018green_esd_rc_v5p0_0.VRC.t12 DVSS 0.007154f
C106 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/comp018green_esd_rc_v5p0_0.VRC.n0 DVSS 0.006386f
C107 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/comp018green_esd_rc_v5p0_0.VRC.t11 DVSS 0.006489f
C108 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/comp018green_esd_rc_v5p0_0.VRC.t1 DVSS 0.007154f
C109 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/comp018green_esd_rc_v5p0_0.VRC.n1 DVSS 0.006386f
C110 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/comp018green_esd_rc_v5p0_0.VRC.t2 DVSS 0.006489f
C111 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/comp018green_esd_rc_v5p0_0.VRC.n2 DVSS 2.47e-19
C112 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/comp018green_esd_rc_v5p0_0.VRC.n3 DVSS 0.041889f
C113 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/comp018green_esd_rc_v5p0_0.VRC.t3 DVSS 0.006457f
C114 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/comp018green_esd_rc_v5p0_0.VRC.n4 DVSS 0.078598f
C115 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/comp018green_esd_rc_v5p0_0.VRC.t6 DVSS 0.30082f
C116 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/comp018green_esd_rc_v5p0_0.VRC.n6 DVSS 0.0218f
C117 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/comp018green_esd_rc_v5p0_0.VRC.t7 DVSS 0.30082f
C118 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/comp018green_esd_rc_v5p0_0.VRC.n8 DVSS 0.021728f
C119 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/comp018green_esd_rc_v5p0_0.VRC.t4 DVSS 0.30082f
C120 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/comp018green_esd_rc_v5p0_0.VRC.n10 DVSS 0.02355f
C121 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/comp018green_esd_rc_v5p0_0.VRC.t5 DVSS 0.30082f
C122 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/comp018green_esd_rc_v5p0_0.VRC.n12 DVSS 0.066169f
C123 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/comp018green_esd_rc_v5p0_0.VRC.t10 DVSS 0.30082f
C124 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/comp018green_esd_rc_v5p0_0.VRC.n14 DVSS 0.0218f
C125 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/comp018green_esd_rc_v5p0_0.VRC.t13 DVSS 0.30082f
C126 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/comp018green_esd_rc_v5p0_0.VRC.n16 DVSS 0.021728f
C127 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/comp018green_esd_rc_v5p0_0.VRC.t8 DVSS 0.30082f
C128 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/comp018green_esd_rc_v5p0_0.VRC.n18 DVSS 0.02634f
C129 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/comp018green_esd_rc_v5p0_0.VRC.t9 DVSS 0.30082f
C130 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531459_0.D.t0 DVSS 0.428625f
C131 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531459_0.D.t2 DVSS 0.326607f
C132 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531459_0.D.n0 DVSS 1.49938f
C133 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531459_0.D.t1 DVSS 0.332988f
C134 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531459_0.D.t9 DVSS 0.396162f
C135 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531459_0.D.t10 DVSS 0.359359f
C136 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531459_0.D.n1 DVSS 0.36046f
C137 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531459_0.D.t5 DVSS 0.359359f
C138 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531459_0.D.n2 DVSS 0.198632f
C139 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531459_0.D.t4 DVSS 0.396162f
C140 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531459_0.D.t3 DVSS 0.359359f
C141 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531459_0.D.n3 DVSS 0.36046f
C142 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531459_0.D.t8 DVSS 0.359359f
C143 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531459_0.D.n4 DVSS 0.198632f
C144 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531459_0.D.n5 DVSS 0.270963f
C145 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531459_0.D.t11 DVSS 0.396162f
C146 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531459_0.D.t7 DVSS 0.396162f
C147 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531459_0.D.t6 DVSS 0.359359f
C148 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531459_0.D.n6 DVSS 0.541808f
C149 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_1.D.n0 DVSS 0.139192f
C150 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_1.D.n1 DVSS 1.54267f
C151 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_1.D.t1 DVSS 0.45513f
C152 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_1.D.t0 DVSS 1.68789f
C153 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_1.D.t2 DVSS 0.453717f
C154 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_1.D.t3 DVSS 1.1716f
C155 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_1.D.t26 DVSS 0.419355f
C156 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_1.D.t4 DVSS 0.380396f
C157 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_1.D.n2 DVSS 0.381563f
C158 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_1.D.t22 DVSS 0.380396f
C159 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_1.D.n3 DVSS 0.21026f
C160 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_1.D.t15 DVSS 0.419355f
C161 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_1.D.t14 DVSS 0.380396f
C162 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_1.D.n4 DVSS 0.381563f
C163 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_1.D.t23 DVSS 0.380396f
C164 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_1.D.n5 DVSS 0.21026f
C165 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_1.D.t31 DVSS 0.419355f
C166 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_1.D.t16 DVSS 0.380396f
C167 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_1.D.n6 DVSS 0.381563f
C168 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_1.D.t25 DVSS 0.380396f
C169 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_1.D.n7 DVSS 0.217488f
C170 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_1.D.t33 DVSS 0.380396f
C171 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_1.D.n8 DVSS 0.217488f
C172 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_1.D.t13 DVSS 0.380396f
C173 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_1.D.n9 DVSS 0.217488f
C174 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_1.D.t19 DVSS 0.380396f
C175 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_1.D.n10 DVSS 0.217488f
C176 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_1.D.t28 DVSS 0.380396f
C177 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_1.D.n11 DVSS 0.217488f
C178 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_1.D.t5 DVSS 0.380396f
C179 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_1.D.n12 DVSS 0.217488f
C180 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_1.D.t17 DVSS 0.380396f
C181 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_1.D.n13 DVSS 0.217488f
C182 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_1.D.t21 DVSS 0.380396f
C183 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_1.D.n14 DVSS 0.217488f
C184 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_1.D.t7 DVSS 0.380396f
C185 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_1.D.n15 DVSS 0.217488f
C186 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_1.D.t8 DVSS 0.380396f
C187 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_1.D.n16 DVSS 0.21026f
C188 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_1.D.t12 DVSS 0.419355f
C189 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_1.D.t11 DVSS 0.380396f
C190 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_1.D.n17 DVSS 0.381563f
C191 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_1.D.t20 DVSS 0.380396f
C192 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_1.D.n18 DVSS 0.217488f
C193 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_1.D.t9 DVSS 0.380396f
C194 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_1.D.n19 DVSS 0.217488f
C195 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_1.D.t32 DVSS 0.380396f
C196 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_1.D.n20 DVSS 0.217488f
C197 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_1.D.t24 DVSS 0.380396f
C198 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_1.D.n21 DVSS 0.217488f
C199 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_1.D.t18 DVSS 0.380396f
C200 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_1.D.n22 DVSS 0.217488f
C201 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_1.D.t30 DVSS 0.380396f
C202 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_1.D.n23 DVSS 0.217488f
C203 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_1.D.t29 DVSS 0.380396f
C204 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_1.D.n24 DVSS 0.217488f
C205 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_1.D.t10 DVSS 0.380396f
C206 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_1.D.n25 DVSS 0.217488f
C207 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_1.D.t6 DVSS 0.380396f
C208 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_1.D.n26 DVSS 0.217488f
C209 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_1.D.t27 DVSS 0.380396f
C210 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_1.D.n27 DVSS 0.21026f
C211 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n0 DVSS 1.8071f
C212 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n1 DVSS 1.36365f
C213 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n2 DVSS 1.08485f
C214 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n3 DVSS 1.32384f
C215 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n4 DVSS 1.33565f
C216 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n5 DVSS 1.08373f
C217 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n6 DVSS 1.31923f
C218 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n7 DVSS 3.83312f
C219 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n8 DVSS 1.12015f
C220 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n9 DVSS 1.32384f
C221 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n10 DVSS 0.164547f
C222 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n11 DVSS 0.132556f
C223 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n12 DVSS 1.09441f
C224 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n13 DVSS 0.148653f
C225 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n14 DVSS 0.202716f
C226 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n15 DVSS 0.195803f
C227 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n16 DVSS 0.148653f
C228 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n17 DVSS 1.89711f
C229 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n18 DVSS 0.135251f
C230 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n19 DVSS 0.080926f
C231 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n20 DVSS 0.067727f
C232 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n21 DVSS 0.080926f
C233 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n22 DVSS 0.080926f
C234 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n23 DVSS 0.080926f
C235 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n24 DVSS 0.080926f
C236 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n25 DVSS 0.080926f
C237 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n26 DVSS 0.080926f
C238 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n27 DVSS 0.080926f
C239 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n28 DVSS 0.060915f
C240 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n29 DVSS 0.080926f
C241 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n30 DVSS 0.047375f
C242 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n31 DVSS 0.080926f
C243 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n32 DVSS 0.080926f
C244 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n33 DVSS 0.080926f
C245 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n34 DVSS 0.080926f
C246 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n35 DVSS 0.080926f
C247 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n36 DVSS 0.080926f
C248 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n37 DVSS 0.080926f
C249 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n38 DVSS 0.074432f
C250 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n39 DVSS 0.155483f
C251 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n40 DVSS 1.1182f
C252 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n41 DVSS 0.080926f
C253 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n42 DVSS 0.080926f
C254 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n43 DVSS 0.067727f
C255 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n44 DVSS 0.080926f
C256 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n45 DVSS 0.080926f
C257 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n46 DVSS 0.080926f
C258 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n47 DVSS 0.080926f
C259 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n48 DVSS 0.080926f
C260 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n49 DVSS 0.080926f
C261 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n50 DVSS 0.080926f
C262 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n51 DVSS 0.060915f
C263 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n52 DVSS 0.080926f
C264 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n53 DVSS 0.047375f
C265 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n54 DVSS 0.080926f
C266 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n55 DVSS 0.080926f
C267 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n56 DVSS 0.080926f
C268 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n57 DVSS 0.080926f
C269 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n58 DVSS 0.080926f
C270 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n59 DVSS 0.080926f
C271 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n60 DVSS 0.155483f
C272 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n61 DVSS 0.074432f
C273 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n62 DVSS 1.12226f
C274 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n63 DVSS 0.135251f
C275 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n64 DVSS 0.080926f
C276 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n65 DVSS 0.067727f
C277 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n66 DVSS 0.080926f
C278 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n67 DVSS 0.080926f
C279 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n68 DVSS 0.080926f
C280 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n69 DVSS 0.080926f
C281 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n70 DVSS 0.080926f
C282 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n71 DVSS 0.080926f
C283 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n72 DVSS 0.080926f
C284 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n73 DVSS 0.060915f
C285 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n74 DVSS 0.080926f
C286 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n75 DVSS 0.047375f
C287 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n76 DVSS 0.080926f
C288 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n77 DVSS 0.080926f
C289 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n78 DVSS 0.080926f
C290 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n79 DVSS 0.080926f
C291 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n80 DVSS 0.080926f
C292 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n81 DVSS 0.080926f
C293 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n82 DVSS 0.080926f
C294 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n83 DVSS 0.074432f
C295 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n84 DVSS 0.657969f
C296 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n85 DVSS 1.11876f
C297 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n86 DVSS 1.16277f
C298 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n87 DVSS 0.135251f
C299 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n88 DVSS 1.16826f
C300 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n89 DVSS 1.16277f
C301 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.t3 DVSS 0.099757f
C302 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n90 DVSS 0.107847f
C303 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n91 DVSS 0.219556f
C304 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.t11 DVSS 0.099757f
C305 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n92 DVSS 0.107847f
C306 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.t5 DVSS 0.099757f
C307 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n93 DVSS 0.078524f
C308 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.t7 DVSS 0.099757f
C309 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n94 DVSS 0.107847f
C310 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n95 DVSS 0.107847f
C311 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.t10 DVSS 0.099757f
C312 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n96 DVSS 0.107847f
C313 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.t9 DVSS 0.099757f
C314 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n97 DVSS 0.107847f
C315 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.t1 DVSS 0.099757f
C316 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n98 DVSS 0.107847f
C317 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.t2 DVSS 0.099757f
C318 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n99 DVSS 0.107847f
C319 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.t14 DVSS 0.099757f
C320 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.t12 DVSS 0.272103f
C321 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.t4 DVSS 0.128443f
C322 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.t15 DVSS 0.024353f
C323 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.t0 DVSS 0.024353f
C324 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n100 DVSS 0.080376f
C325 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.t13 DVSS 0.075054f
C326 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n101 DVSS 0.039523f
C327 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n102 DVSS 0.068017f
C328 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.t16 DVSS 0.024353f
C329 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n103 DVSS 0.021026f
C330 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.t41 DVSS 0.663518f
C331 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.t26 DVSS 0.663518f
C332 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.t47 DVSS 0.663518f
C333 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.t90 DVSS 0.663518f
C334 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.t61 DVSS 0.663518f
C335 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.t21 DVSS 0.663518f
C336 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.t85 DVSS 0.663518f
C337 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.t27 DVSS 0.663518f
C338 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.t72 DVSS 0.663518f
C339 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n104 DVSS 0.363297f
C340 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n105 DVSS 0.37381f
C341 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n106 DVSS 0.37381f
C342 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n107 DVSS 0.37381f
C343 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n108 DVSS 0.37381f
C344 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n109 DVSS 0.37381f
C345 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n110 DVSS 0.37381f
C346 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n111 DVSS 0.37381f
C347 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n112 DVSS 0.725746f
C348 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.t37 DVSS 0.689343f
C349 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n113 DVSS 0.725746f
C350 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n114 DVSS 0.37381f
C351 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n115 DVSS 0.37381f
C352 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n116 DVSS 0.37381f
C353 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n117 DVSS 0.37381f
C354 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n118 DVSS 0.37381f
C355 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n119 DVSS 0.37381f
C356 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n120 DVSS 0.37381f
C357 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n121 DVSS 0.363297f
C358 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.t96 DVSS 0.663518f
C359 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.t31 DVSS 0.663518f
C360 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.t89 DVSS 0.663518f
C361 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.t46 DVSS 0.663518f
C362 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.t59 DVSS 0.663518f
C363 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.t36 DVSS 0.663518f
C364 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.t53 DVSS 0.663518f
C365 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.t30 DVSS 0.663518f
C366 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.t69 DVSS 0.663518f
C367 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n122 DVSS 0.363297f
C368 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n123 DVSS 0.37381f
C369 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n124 DVSS 0.37381f
C370 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n125 DVSS 0.37381f
C371 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n126 DVSS 0.37381f
C372 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n127 DVSS 0.37381f
C373 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n128 DVSS 0.37381f
C374 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n129 DVSS 0.37381f
C375 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n130 DVSS 0.725746f
C376 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.t19 DVSS 0.689343f
C377 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n131 DVSS 0.725746f
C378 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n132 DVSS 0.37381f
C379 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n133 DVSS 0.37381f
C380 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n134 DVSS 0.37381f
C381 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n135 DVSS 0.37381f
C382 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n136 DVSS 0.37381f
C383 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n137 DVSS 0.37381f
C384 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n138 DVSS 0.37381f
C385 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n139 DVSS 0.363297f
C386 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n140 DVSS 0.172297f
C387 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n141 DVSS 0.146915f
C388 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.t25 DVSS 0.663518f
C389 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.t68 DVSS 0.663518f
C390 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.t29 DVSS 0.663518f
C391 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.t76 DVSS 0.663518f
C392 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.t84 DVSS 0.663518f
C393 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.t43 DVSS 0.663518f
C394 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.t70 DVSS 0.663518f
C395 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.t52 DVSS 0.663518f
C396 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.t80 DVSS 0.663518f
C397 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n142 DVSS 0.363297f
C398 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n143 DVSS 0.37381f
C399 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n144 DVSS 0.37381f
C400 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n145 DVSS 0.37381f
C401 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n146 DVSS 0.37381f
C402 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n147 DVSS 0.37381f
C403 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n148 DVSS 0.37381f
C404 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n149 DVSS 0.37381f
C405 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n150 DVSS 0.725746f
C406 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.t67 DVSS 0.689343f
C407 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n151 DVSS 0.725746f
C408 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n152 DVSS 0.37381f
C409 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n153 DVSS 0.37381f
C410 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n154 DVSS 0.37381f
C411 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n155 DVSS 0.37381f
C412 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n156 DVSS 0.37381f
C413 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n157 DVSS 0.37381f
C414 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n158 DVSS 0.37381f
C415 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n159 DVSS 0.363297f
C416 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.t58 DVSS 0.663518f
C417 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.t94 DVSS 0.663518f
C418 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.t51 DVSS 0.663518f
C419 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.t86 DVSS 0.663518f
C420 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.t39 DVSS 0.663518f
C421 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.t18 DVSS 0.663518f
C422 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.t34 DVSS 0.663518f
C423 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.t78 DVSS 0.663518f
C424 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.t24 DVSS 0.663518f
C425 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n160 DVSS 0.363297f
C426 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n161 DVSS 0.37381f
C427 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n162 DVSS 0.37381f
C428 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n163 DVSS 0.37381f
C429 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n164 DVSS 0.37381f
C430 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n165 DVSS 0.37381f
C431 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n166 DVSS 0.37381f
C432 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n167 DVSS 0.37381f
C433 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n168 DVSS 0.725746f
C434 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.t64 DVSS 0.689343f
C435 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n169 DVSS 0.725746f
C436 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n170 DVSS 0.37381f
C437 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n171 DVSS 0.37381f
C438 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n172 DVSS 0.37381f
C439 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n173 DVSS 0.37381f
C440 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n174 DVSS 0.37381f
C441 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n175 DVSS 0.37381f
C442 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n176 DVSS 0.37381f
C443 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n177 DVSS 0.363297f
C444 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n178 DVSS 0.021026f
C445 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n179 DVSS 0.053562f
C446 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n180 DVSS 0.021026f
C447 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.t44 DVSS 0.663518f
C448 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.t75 DVSS 0.663518f
C449 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.t54 DVSS 0.663518f
C450 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.t83 DVSS 0.663518f
C451 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.t40 DVSS 0.663518f
C452 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.t88 DVSS 0.663518f
C453 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.t45 DVSS 0.663518f
C454 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.t32 DVSS 0.663518f
C455 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.t60 DVSS 0.663518f
C456 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n181 DVSS 0.363297f
C457 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n182 DVSS 0.37381f
C458 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n183 DVSS 0.37381f
C459 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n184 DVSS 0.37381f
C460 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n185 DVSS 0.37381f
C461 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n186 DVSS 0.37381f
C462 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n187 DVSS 0.37381f
C463 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n188 DVSS 0.37381f
C464 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n189 DVSS 0.725746f
C465 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.t20 DVSS 0.689343f
C466 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n190 DVSS 0.725746f
C467 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n191 DVSS 0.37381f
C468 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n192 DVSS 0.37381f
C469 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n193 DVSS 0.37381f
C470 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n194 DVSS 0.37381f
C471 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n195 DVSS 0.37381f
C472 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n196 DVSS 0.37381f
C473 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n197 DVSS 0.37381f
C474 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n198 DVSS 0.363297f
C475 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.t66 DVSS 0.663518f
C476 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.t35 DVSS 0.663518f
C477 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.t79 DVSS 0.663518f
C478 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.t92 DVSS 0.663518f
C479 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.t74 DVSS 0.663518f
C480 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.t82 DVSS 0.663518f
C481 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.t57 DVSS 0.663518f
C482 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.t17 DVSS 0.663518f
C483 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.t50 DVSS 0.663518f
C484 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n199 DVSS 0.363297f
C485 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n200 DVSS 0.37381f
C486 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n201 DVSS 0.37381f
C487 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n202 DVSS 0.37381f
C488 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n203 DVSS 0.37381f
C489 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n204 DVSS 0.37381f
C490 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n205 DVSS 0.37381f
C491 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n206 DVSS 0.37381f
C492 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n207 DVSS 0.725746f
C493 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.t87 DVSS 0.689343f
C494 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n208 DVSS 0.725746f
C495 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n209 DVSS 0.37381f
C496 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n210 DVSS 0.37381f
C497 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n211 DVSS 0.37381f
C498 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n212 DVSS 0.37381f
C499 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n213 DVSS 0.37381f
C500 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n214 DVSS 0.37381f
C501 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n215 DVSS 0.37381f
C502 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n216 DVSS 0.363297f
C503 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n217 DVSS 0.172297f
C504 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n218 DVSS 0.363297f
C505 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.t42 DVSS 0.663518f
C506 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.t81 DVSS 0.663518f
C507 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.t33 DVSS 0.663518f
C508 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.t77 DVSS 0.663518f
C509 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.t48 DVSS 0.663518f
C510 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.t62 DVSS 0.663518f
C511 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.t22 DVSS 0.663518f
C512 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.t55 DVSS 0.663518f
C513 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.t95 DVSS 0.663518f
C514 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.t91 DVSS 0.663518f
C515 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.t49 DVSS 0.663518f
C516 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.t93 DVSS 0.663518f
C517 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.t63 DVSS 0.663518f
C518 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.t23 DVSS 0.663518f
C519 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.t73 DVSS 0.663518f
C520 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.t28 DVSS 0.663518f
C521 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.t56 DVSS 0.663518f
C522 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.t38 DVSS 0.663518f
C523 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n219 DVSS 0.37381f
C524 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n220 DVSS 0.37381f
C525 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n221 DVSS 0.37381f
C526 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n222 DVSS 0.37381f
C527 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n223 DVSS 0.37381f
C528 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n224 DVSS 0.37381f
C529 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n225 DVSS 0.37381f
C530 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n226 DVSS 0.725746f
C531 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.t65 DVSS 0.689343f
C532 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n227 DVSS 0.725746f
C533 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n228 DVSS 0.37381f
C534 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n229 DVSS 0.37381f
C535 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n230 DVSS 0.37381f
C536 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n231 DVSS 0.37381f
C537 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n232 DVSS 0.37381f
C538 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n233 DVSS 0.37381f
C539 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n234 DVSS 0.37381f
C540 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n235 DVSS 0.363297f
C541 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n236 DVSS 0.021026f
C542 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n237 DVSS 0.363297f
C543 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n238 DVSS 0.37381f
C544 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n239 DVSS 0.37381f
C545 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n240 DVSS 0.37381f
C546 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n241 DVSS 0.37381f
C547 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n242 DVSS 0.37381f
C548 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n243 DVSS 0.37381f
C549 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n244 DVSS 0.37381f
C550 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n245 DVSS 0.725746f
C551 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.t71 DVSS 0.689343f
C552 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n246 DVSS 0.725746f
C553 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n247 DVSS 0.37381f
C554 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n248 DVSS 0.37381f
C555 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n249 DVSS 0.37381f
C556 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n250 DVSS 0.37381f
C557 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n251 DVSS 0.37381f
C558 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n252 DVSS 0.37381f
C559 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n253 DVSS 0.37381f
C560 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n254 DVSS 0.363297f
C561 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n255 DVSS 0.053562f
C562 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n256 DVSS 0.053562f
C563 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n257 DVSS 1.52893f
C564 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.t6 DVSS 0.024353f
C565 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n258 DVSS 0.048705f
C566 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n259 DVSS 0.073677f
C567 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n260 DVSS 0.15975f
C568 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.t8 DVSS 0.075054f
C569 GF_NI_DVSS_BASE_0.comp018green_esd_clamp_v5p0_DVSS_0/nmos_6p0_CDNS_406619531458_0.D.n261 DVSS 0.039523f
C570 DVDD.n0 DVSS 0.02223f
C571 DVDD.n1 DVSS 0.024661f
C572 DVDD.n2 DVSS 0.024661f
C573 DVDD.n3 DVSS 0.024661f
C574 DVDD.n4 DVSS 0.024661f
C575 DVDD.n5 DVSS 0.024661f
C576 DVDD.n6 DVSS 0.024661f
C577 DVDD.n7 DVSS 0.024661f
C578 DVDD.n8 DVSS 0.024661f
C579 DVDD.n9 DVSS 0.024661f
C580 DVDD.n10 DVSS 0.024661f
C581 DVDD.n11 DVSS 0.01233f
C582 DVDD.n12 DVSS 0.024661f
C583 DVDD.n13 DVSS 0.024661f
C584 DVDD.n14 DVSS 0.024661f
C585 DVDD.n15 DVSS 0.024661f
C586 DVDD.n16 DVSS 0.00226f
C587 DVDD.n17 DVSS 0.010767f
C588 DVDD.n18 DVSS 0.001538f
C589 DVDD.n19 DVSS 0.003076f
C590 DVDD.n20 DVSS 0.003076f
C591 DVDD.n21 DVSS 0.001538f
C592 DVDD.n22 DVSS 0.002928f
C593 DVDD.n23 DVSS 0.003076f
C594 DVDD.n24 DVSS 0.003076f
C595 DVDD.n25 DVSS 0.001538f
C596 DVDD.n26 DVSS 0.003052f
C597 DVDD.n27 DVSS 4.9e-19
C598 DVDD.n28 DVSS 5.09e-19
C599 DVDD.n29 DVSS 9.8e-19
C600 DVDD.n30 DVSS 0.001161f
C601 DVDD.n31 DVSS 0.350325f
C602 DVDD.n32 DVSS 9.8e-19
C603 DVDD.n33 DVSS 0.001161f
C604 DVDD.n34 DVSS 9.8e-19
C605 DVDD.n36 DVSS 0.001161f
C606 DVDD.n37 DVSS 9.8e-19
C607 DVDD.n39 DVSS 0.001161f
C608 DVDD.t5 DVSS 0.00165f
C609 DVDD.n41 DVSS 0.002127f
C610 DVDD.n42 DVSS 0.001161f
C611 DVDD.n43 DVSS 8.77e-19
C612 DVDD.n44 DVSS 0.001161f
C613 DVDD.n45 DVSS 0.150384f
C614 DVDD.n46 DVSS 0.001161f
C615 DVDD.n47 DVSS 0.0013f
C616 DVDD.n48 DVSS 8.77e-19
C617 DVDD.n49 DVSS 0.001161f
C618 DVDD.t4 DVSS 0.088863f
C619 DVDD.n50 DVSS 0.001161f
C620 DVDD.n51 DVSS 0.001161f
C621 DVDD.n52 DVSS 0.001161f
C622 DVDD.t70 DVSS 0.088863f
C623 DVDD.n53 DVSS 0.001161f
C624 DVDD.n54 DVSS 8.77e-19
C625 DVDD.n55 DVSS 0.001161f
C626 DVDD.n56 DVSS 0.143548f
C627 DVDD.n57 DVSS 0.001161f
C628 DVDD.n58 DVSS 0.001161f
C629 DVDD.n59 DVSS 0.001161f
C630 DVDD.n60 DVSS 0.157219f
C631 DVDD.n61 DVSS 0.001161f
C632 DVDD.n62 DVSS 8.77e-19
C633 DVDD.n63 DVSS 0.001161f
C634 DVDD.t71 DVSS 0.088863f
C635 DVDD.n64 DVSS 0.001161f
C636 DVDD.n65 DVSS 0.001161f
C637 DVDD.n66 DVSS 0.001161f
C638 DVDD.t6 DVSS 0.088863f
C639 DVDD.n67 DVSS 0.001161f
C640 DVDD.n68 DVSS 8.77e-19
C641 DVDD.n69 DVSS 0.001161f
C642 DVDD.n70 DVSS 0.136712f
C643 DVDD.n71 DVSS 0.001161f
C644 DVDD.n72 DVSS 0.001161f
C645 DVDD.n73 DVSS 0.001161f
C646 DVDD.n74 DVSS 0.164055f
C647 DVDD.n75 DVSS 0.001161f
C648 DVDD.n76 DVSS 8.77e-19
C649 DVDD.n77 DVSS 0.001161f
C650 DVDD.t52 DVSS 0.088863f
C651 DVDD.n78 DVSS 0.001161f
C652 DVDD.n79 DVSS 0.001161f
C653 DVDD.n80 DVSS 0.001161f
C654 DVDD.t9 DVSS 0.088863f
C655 DVDD.n81 DVSS 0.001161f
C656 DVDD.n82 DVSS 8.77e-19
C657 DVDD.n83 DVSS 0.001161f
C658 DVDD.n84 DVSS 0.129877f
C659 DVDD.n85 DVSS 0.001161f
C660 DVDD.n86 DVSS 0.001161f
C661 DVDD.n87 DVSS 0.001161f
C662 DVDD.n88 DVSS 0.17089f
C663 DVDD.n89 DVSS 0.001161f
C664 DVDD.n90 DVSS 8.77e-19
C665 DVDD.n91 DVSS 0.001161f
C666 DVDD.t12 DVSS 0.088863f
C667 DVDD.n92 DVSS 0.001161f
C668 DVDD.n93 DVSS 0.001161f
C669 DVDD.n94 DVSS 0.001161f
C670 DVDD.t27 DVSS 0.088863f
C671 DVDD.n95 DVSS 0.001161f
C672 DVDD.n96 DVSS 8.77e-19
C673 DVDD.n97 DVSS 0.001161f
C674 DVDD.n98 DVSS 0.123041f
C675 DVDD.n99 DVSS 0.001161f
C676 DVDD.n100 DVSS 0.001161f
C677 DVDD.n101 DVSS 0.001161f
C678 DVDD.n102 DVSS 0.220449f
C679 DVDD.n103 DVSS 0.001189f
C680 DVDD.n104 DVSS 9.8e-19
C681 DVDD.n105 DVSS 0.001161f
C682 DVDD.n167 DVSS 0.001161f
C683 DVDD.n169 DVSS 5.09e-19
C684 DVDD.n170 DVSS 0.002059f
C685 DVDD.n171 DVSS 0.005483f
C686 DVDD.n172 DVSS 4.9e-19
C687 DVDD.n173 DVSS 9.24e-19
C688 DVDD.n174 DVSS 0.002059f
C689 DVDD.n175 DVSS 0.003076f
C690 DVDD.n176 DVSS 0.064196f
C691 DVDD.n177 DVSS 0.023631f
C692 DVDD.n178 DVSS 0.011968f
C693 DVDD.n179 DVSS 0.008245f
C694 DVDD.n180 DVSS 0.007156f
C695 DVDD.n181 DVSS 0.003523f
C696 DVDD.n182 DVSS 0.003076f
C697 DVDD.n183 DVSS 0.007046f
C698 DVDD.n184 DVSS 0.465466f
C699 DVDD.n185 DVSS 0.003076f
C700 DVDD.n186 DVSS 0.065183f
C701 DVDD.n187 DVSS 0.065324f
C702 DVDD.n188 DVSS 0.031815f
C703 DVDD.n189 DVSS 0.040378f
C704 DVDD.n190 DVSS 0.03889f
C705 DVDD.n191 DVSS 0.031918f
C706 DVDD.n192 DVSS 0.040378f
C707 DVDD.n193 DVSS 0.03889f
C708 DVDD.n194 DVSS 0.007613f
C709 DVDD.n195 DVSS 0.071557f
C710 DVDD.n196 DVSS 0.031918f
C711 DVDD.n197 DVSS 0.031815f
C712 DVDD.n198 DVSS 0.040378f
C713 DVDD.n199 DVSS 0.03889f
C714 DVDD.n200 DVSS 0.005384f
C715 DVDD.n201 DVSS 0.03889f
C716 DVDD.n202 DVSS 0.023073f
C717 DVDD.n203 DVSS 0.052845f
C718 DVDD.n204 DVSS 0.052845f
C719 DVDD.n205 DVSS 0.023073f
C720 DVDD.n206 DVSS 0.023073f
C721 DVDD.n207 DVSS 0.062707f
C722 DVDD.n208 DVSS 0.08485f
C723 DVDD.n209 DVSS 0.052845f
C724 DVDD.n210 DVSS 0.023073f
C725 DVDD.n211 DVSS 0.023073f
C726 DVDD.n212 DVSS 0.023073f
C727 DVDD.n213 DVSS 0.040378f
C728 DVDD.n214 DVSS 0.071557f
C729 DVDD.n215 DVSS 0.031917f
C730 DVDD.n216 DVSS 0.03889f
C731 DVDD.n217 DVSS 0.040378f
C732 DVDD.n218 DVSS 0.031815f
C733 DVDD.n219 DVSS 0.040378f
C734 DVDD.n220 DVSS 0.03889f
C735 DVDD.n221 DVSS 0.031917f
C736 DVDD.n222 DVSS 0.005185f
C737 DVDD.n223 DVSS 0.005384f
C738 DVDD.n224 DVSS 0.03889f
C739 DVDD.n225 DVSS 0.031815f
C740 DVDD.n226 DVSS 0.065321f
C741 DVDD.n227 DVSS 0.065181f
C742 DVDD.n228 DVSS 0.040378f
C743 DVDD.n229 DVSS 0.052845f
C744 DVDD.n230 DVSS 0.20396f
C745 DVDD.n231 DVSS 0.052845f
C746 DVDD.n232 DVSS 0.066256f
C747 DVDD.n233 DVSS 0.447728f
C748 DVDD.n234 DVSS 0.023073f
C749 DVDD.n235 DVSS 0.003076f
C750 DVDD.n236 DVSS 0.003076f
C751 DVDD.n237 DVSS 0.026423f
C752 DVDD.n238 DVSS 0.152989f
C753 DVDD.n239 DVSS 0.053362f
C754 DVDD.n240 DVSS 0.053408f
C755 DVDD.n241 DVSS 0.001538f
C756 DVDD.n242 DVSS 0.031074f
C757 DVDD.n243 DVSS 0.023073f
C758 DVDD.n244 DVSS 0.003076f
C759 DVDD.n245 DVSS 0.003076f
C760 DVDD.n246 DVSS 0.003076f
C761 DVDD.n247 DVSS 0.003076f
C762 DVDD.n248 DVSS 0.003076f
C763 DVDD.n249 DVSS 0.003076f
C764 DVDD.n250 DVSS 0.003076f
C765 DVDD.n251 DVSS 0.003076f
C766 DVDD.n252 DVSS 0.003076f
C767 DVDD.n253 DVSS 0.003076f
C768 DVDD.n254 DVSS 0.003076f
C769 DVDD.n255 DVSS 0.001538f
C770 DVDD.n256 DVSS 0.003163f
C771 DVDD.t17 DVSS 0.065353f
C772 DVDD.t18 DVSS 0.013249f
C773 DVDD.t24 DVSS 0.003225f
C774 DVDD.t58 DVSS 0.003225f
C775 DVDD.n257 DVSS 0.011936f
C776 DVDD.t33 DVSS 0.003225f
C777 DVDD.t22 DVSS 0.003225f
C778 DVDD.n258 DVSS 0.011936f
C779 DVDD.t43 DVSS 0.003225f
C780 DVDD.t69 DVSS 0.003225f
C781 DVDD.n259 DVSS 0.011663f
C782 DVDD.n260 DVSS 0.008739f
C783 DVDD.n261 DVSS 0.004305f
C784 DVDD.n262 DVSS 0.001538f
C785 DVDD.n263 DVSS 0.01697f
C786 DVDD.n264 DVSS 0.001538f
C787 DVDD.n265 DVSS 0.003076f
C788 DVDD.n266 DVSS 0.003076f
C789 DVDD.n267 DVSS 0.003076f
C790 DVDD.n268 DVSS 0.003076f
C791 DVDD.n269 DVSS 0.003076f
C792 DVDD.n270 DVSS 0.003076f
C793 DVDD.n271 DVSS 0.003076f
C794 DVDD.n272 DVSS 0.003076f
C795 DVDD.n273 DVSS 0.014092f
C796 DVDD.n274 DVSS 0.028184f
C797 DVDD.n275 DVSS 0.028184f
C798 DVDD.n276 DVSS 0.028184f
C799 DVDD.n277 DVSS 0.028184f
C800 DVDD.n278 DVSS 0.028184f
C801 DVDD.n279 DVSS 0.027092f
C802 DVDD.n280 DVSS 0.018062f
C803 DVDD.n281 DVSS 0.018062f
C804 DVDD.n282 DVSS 0.033866f
C805 DVDD.n283 DVSS 0.045402f
C806 DVDD.n284 DVSS 0.028184f
C807 DVDD.n285 DVSS 0.040514f
C808 DVDD.n286 DVSS 0.028184f
C809 DVDD.n287 DVSS 0.040514f
C810 DVDD.n288 DVSS 0.028184f
C811 DVDD.n289 DVSS 0.028184f
C812 DVDD.n290 DVSS 0.028184f
C813 DVDD.n291 DVSS 0.028184f
C814 DVDD.n292 DVSS 0.028184f
C815 DVDD.n293 DVSS 0.028184f
C816 DVDD.n294 DVSS 0.026001f
C817 DVDD.n295 DVSS 0.026001f
C818 DVDD.n296 DVSS 0.004764f
C819 DVDD.n297 DVSS 0.003076f
C820 DVDD.n298 DVSS 0.003076f
C821 DVDD.n301 DVSS 0.003523f
C822 DVDD.n302 DVSS 0.005384f
C823 DVDD.n303 DVSS 0.007046f
C824 DVDD.n304 DVSS 0.005384f
C825 DVDD.n305 DVSS 0.00698f
C826 DVDD.n306 DVSS 0.003076f
C827 DVDD.n307 DVSS 0.003399f
C828 DVDD.n308 DVSS 0.008245f
C829 DVDD.n309 DVSS 0.008245f
C830 DVDD.n312 DVSS 0.026423f
C831 DVDD.n313 DVSS 0.024376f
C832 DVDD.n314 DVSS 0.031819f
C833 DVDD.n315 DVSS 0.006948f
C834 DVDD.n316 DVSS 0.008245f
C835 DVDD.n317 DVSS 0.006682f
C836 DVDD.n318 DVSS 0.008245f
C837 DVDD.n319 DVSS 0.008245f
C838 DVDD.n320 DVSS 0.008245f
C839 DVDD.n321 DVSS 0.008245f
C840 DVDD.n322 DVSS 0.008245f
C841 DVDD.n323 DVSS 0.00359f
C842 DVDD.n324 DVSS 0.007613f
C843 DVDD.n325 DVSS 0.008245f
C844 DVDD.n326 DVSS 0.023073f
C845 DVDD.n328 DVSS 0.008245f
C846 DVDD.n330 DVSS 0.008245f
C847 DVDD.n331 DVSS 0.00359f
C848 DVDD.n333 DVSS 0.005818f
C849 DVDD.n335 DVSS 0.008245f
C850 DVDD.n337 DVSS 0.008245f
C851 DVDD.n339 DVSS 0.008245f
C852 DVDD.n341 DVSS 0.008245f
C853 DVDD.n342 DVSS 0.005685f
C854 DVDD.n344 DVSS 0.008245f
C855 DVDD.n345 DVSS 0.005419f
C856 DVDD.n355 DVSS 0.02512f
C857 DVDD.n357 DVSS 0.006416f
C858 DVDD.n358 DVSS 0.01188f
C859 DVDD.n359 DVSS 0.01104f
C860 DVDD.n360 DVSS 0.004999f
C861 DVDD.n361 DVSS 0.001538f
C862 DVDD.n362 DVSS 0.051543f
C863 DVDD.n363 DVSS 0.00289f
C864 DVDD.n364 DVSS 0.002791f
C865 DVDD.n365 DVSS 0.002692f
C866 DVDD.n366 DVSS 0.002593f
C867 DVDD.n367 DVSS 0.002493f
C868 DVDD.n368 DVSS 0.023073f
C869 DVDD.n369 DVSS 0.003076f
C870 DVDD.n370 DVSS 0.002121f
C871 DVDD.n371 DVSS 0.003076f
C872 DVDD.n372 DVSS 0.002022f
C873 DVDD.n373 DVSS 0.003076f
C874 DVDD.n374 DVSS 0.001923f
C875 DVDD.n375 DVSS 0.003076f
C876 DVDD.n376 DVSS 0.001824f
C877 DVDD.n377 DVSS 0.003076f
C878 DVDD.n378 DVSS 0.001724f
C879 DVDD.n379 DVSS 0.003076f
C880 DVDD.n380 DVSS 0.001538f
C881 DVDD.n381 DVSS 0.027944f
C882 DVDD.n383 DVSS 0.051543f
C883 DVDD.n384 DVSS 0.001538f
C884 DVDD.n385 DVSS 0.00299f
C885 DVDD.n386 DVSS 0.00289f
C886 DVDD.n387 DVSS 0.002791f
C887 DVDD.n388 DVSS 0.023073f
C888 DVDD.n389 DVSS 0.001824f
C889 DVDD.n390 DVSS 0.003076f
C890 DVDD.n391 DVSS 0.003076f
C891 DVDD.n392 DVSS 0.003076f
C892 DVDD.n393 DVSS 0.003076f
C893 DVDD.n394 DVSS 0.003076f
C894 DVDD.n395 DVSS 0.001724f
C895 DVDD.n396 DVSS 0.003076f
C896 DVDD.n397 DVSS 0.001625f
C897 DVDD.n398 DVSS 0.001538f
C898 DVDD.n399 DVSS 0.001538f
C899 DVDD.n400 DVSS 0.003064f
C900 DVDD.n401 DVSS 0.031074f
C901 DVDD.n402 DVSS 0.001538f
C902 DVDD.n403 DVSS 0.003076f
C903 DVDD.n404 DVSS 0.003076f
C904 DVDD.n405 DVSS 0.003076f
C905 DVDD.n406 DVSS 0.003076f
C906 DVDD.n407 DVSS 0.001538f
C907 DVDD.n408 DVSS 0.001538f
C908 DVDD.n409 DVSS 0.001538f
C909 DVDD.n410 DVSS 0.001538f
C910 DVDD.n411 DVSS 0.027944f
C911 DVDD.n412 DVSS 0.001538f
C912 DVDD.n413 DVSS 0.051543f
C913 DVDD.n414 DVSS 0.001538f
C914 DVDD.n415 DVSS 0.001538f
C915 DVDD.n416 DVSS 0.001538f
C916 DVDD.n417 DVSS 0.002965f
C917 DVDD.n418 DVSS 0.003076f
C918 DVDD.n419 DVSS 0.00299f
C919 DVDD.n420 DVSS 0.023073f
C920 DVDD.n421 DVSS 0.003076f
C921 DVDD.n422 DVSS 0.001625f
C922 DVDD.n423 DVSS 0.001538f
C923 DVDD.n424 DVSS 0.001551f
C924 DVDD.n425 DVSS 0.001538f
C925 DVDD.n426 DVSS 0.001538f
C926 DVDD.n427 DVSS 0.001538f
C927 DVDD.n428 DVSS 0.001538f
C928 DVDD.n429 DVSS 0.024004f
C929 DVDD.n430 DVSS 0.002667f
C930 DVDD.n431 DVSS 0.002766f
C931 DVDD.n432 DVSS 0.002866f
C932 DVDD.n433 DVSS 0.001538f
C933 DVDD.n434 DVSS 0.001538f
C934 DVDD.n435 DVSS 0.003064f
C935 DVDD.n436 DVSS 0.031074f
C936 DVDD.n437 DVSS 0.001538f
C937 DVDD.n438 DVSS 0.001538f
C938 DVDD.n439 DVSS 0.00165f
C939 DVDD.n440 DVSS 0.003076f
C940 DVDD.n441 DVSS 0.001749f
C941 DVDD.n442 DVSS 0.003076f
C942 DVDD.n443 DVSS 0.008261f
C943 DVDD.n444 DVSS 0.004122f
C944 DVDD.n445 DVSS 0.001538f
C945 DVDD.n446 DVSS 0.002766f
C946 DVDD.n447 DVSS 0.001538f
C947 DVDD.n448 DVSS 0.023073f
C948 DVDD.n449 DVSS 0.002667f
C949 DVDD.n450 DVSS 0.002866f
C950 DVDD.n451 DVSS 0.001538f
C951 DVDD.n452 DVSS 0.001538f
C952 DVDD.n453 DVSS 0.003064f
C953 DVDD.n454 DVSS 0.042611f
C954 DVDD.n455 DVSS 0.001538f
C955 DVDD.n456 DVSS 0.001538f
C956 DVDD.n457 DVSS 0.001538f
C957 DVDD.n458 DVSS 0.00165f
C958 DVDD.n459 DVSS 0.003076f
C959 DVDD.n460 DVSS 0.001749f
C960 DVDD.n461 DVSS 0.003076f
C961 DVDD.n462 DVSS 0.003076f
C962 DVDD.n463 DVSS 0.008262f
C963 DVDD.n464 DVSS 0.001538f
C964 DVDD.n465 DVSS 0.001538f
C965 DVDD.n466 DVSS 0.003076f
C966 DVDD.n467 DVSS 0.003076f
C967 DVDD.n468 DVSS 0.001538f
C968 DVDD.n469 DVSS 0.001538f
C969 DVDD.n470 DVSS 0.001538f
C970 DVDD.n471 DVSS 0.001538f
C971 DVDD.n472 DVSS 0.026423f
C972 DVDD.n473 DVSS 0.013013f
C973 DVDD.n474 DVSS 0.01188f
C974 DVDD.n475 DVSS 0.018359f
C975 DVDD.n476 DVSS 0.027687f
C976 DVDD.n477 DVSS 0.001538f
C977 DVDD.n478 DVSS 0.010767f
C978 DVDD.n479 DVSS 0.002642f
C979 DVDD.n480 DVSS 0.002741f
C980 DVDD.n481 DVSS 0.023706f
C981 DVDD.n482 DVSS 0.003076f
C982 DVDD.n483 DVSS 0.001873f
C983 DVDD.n484 DVSS 0.003076f
C984 DVDD.n485 DVSS 0.001972f
C985 DVDD.n486 DVSS 0.004081f
C986 DVDD.n487 DVSS 0.024661f
C987 DVDD.n488 DVSS 0.024661f
C988 DVDD.n489 DVSS 0.024661f
C989 DVDD.n490 DVSS 0.024661f
C990 DVDD.n491 DVSS 0.024661f
C991 DVDD.n492 DVSS 0.024661f
C992 DVDD.n493 DVSS 0.024661f
C993 DVDD.n494 DVSS 0.024661f
C994 DVDD.n495 DVSS 0.024661f
C995 DVDD.n496 DVSS 0.024661f
C996 DVDD.n497 DVSS 0.024661f
C997 DVDD.n498 DVSS 0.024661f
C998 DVDD.n499 DVSS 0.024661f
C999 DVDD.n500 DVSS 0.024661f
C1000 DVDD.n501 DVSS 0.024661f
C1001 DVDD.n502 DVSS 0.024661f
C1002 DVDD.n503 DVSS 0.024661f
C1003 DVDD.n504 DVSS 0.024661f
C1004 DVDD.n505 DVSS 0.024661f
C1005 DVDD.n506 DVSS 0.01233f
C1006 DVDD.n507 DVSS 0.024661f
C1007 DVDD.n508 DVSS 0.024661f
C1008 DVDD.n509 DVSS 0.024661f
C1009 DVDD.n510 DVSS 0.011375f
C1010 DVDD.n511 DVSS 0.008245f
C1011 DVDD.n513 DVSS 0.008245f
C1012 DVDD.n515 DVSS 0.008245f
C1013 DVDD.n516 DVSS 0.014501f
C1014 DVDD.n518 DVSS 0.004754f
C1015 DVDD.n520 DVSS 0.00502f
C1016 DVDD.n522 DVSS 0.005286f
C1017 DVDD.n524 DVSS 0.032447f
C1018 DVDD.n525 DVSS 0.01188f
C1019 DVDD.n526 DVSS 0.015319f
C1020 DVDD.n527 DVSS 0.004081f
C1021 DVDD.n528 DVSS 0.027944f
C1022 DVDD.n529 DVSS 0.027944f
C1023 DVDD.n530 DVSS 0.027944f
C1024 DVDD.n531 DVSS 0.027944f
C1025 DVDD.n532 DVSS 0.027944f
C1026 DVDD.n533 DVSS 0.027944f
C1027 DVDD.n534 DVSS 0.027944f
C1028 DVDD.n535 DVSS 0.027944f
C1029 DVDD.n536 DVSS 0.027944f
C1030 DVDD.n537 DVSS 0.027944f
C1031 DVDD.n538 DVSS 0.027944f
C1032 DVDD.n539 DVSS 0.027944f
C1033 DVDD.n540 DVSS 0.027944f
C1034 DVDD.n541 DVSS 0.027944f
C1035 DVDD.n542 DVSS 0.027944f
C1036 DVDD.n543 DVSS 0.055632f
C1037 DVDD.n544 DVSS 0.319527f
C1038 DVDD.n545 DVSS 1.00617f
C1039 DVDD.n546 DVSS 0.672128f
C1040 DVDD.n547 DVSS 0.00493f
C1041 DVDD.n549 DVSS 0.008644f
C1042 DVDD.n551 DVSS 0.00493f
C1043 DVDD.n553 DVSS 0.117609f
C1044 DVDD.n555 DVSS 0.032447f
C1045 DVDD.n556 DVSS 0.035866f
C1046 DVDD.n557 DVSS 0.018831f
C1047 DVDD.n558 DVSS 0.001538f
C1048 DVDD.n560 DVSS 0.002841f
C1049 DVDD.n561 DVSS 0.00134f
C1050 DVDD.n562 DVSS 0.001538f
C1051 DVDD.n564 DVSS 0.002841f
C1052 DVDD.n565 DVSS 0.00134f
C1053 DVDD.n566 DVSS 0.004122f
C1054 DVDD.n568 DVSS 0.00493f
C1055 DVDD.n569 DVSS 0.00493f
C1056 DVDD.n571 DVSS -0.285103f
C1057 DVDD.n573 DVSS 0.001538f
C1058 DVDD.n575 DVSS 0.002841f
C1059 DVDD.n576 DVSS 0.00134f
C1060 DVDD.n577 DVSS 0.001538f
C1061 DVDD.n579 DVSS 0.002841f
C1062 DVDD.n580 DVSS 0.026423f
C1063 DVDD.n581 DVSS 0.023073f
C1064 DVDD.n582 DVSS 0.004999f
C1065 DVDD.n584 DVSS 0.001538f
C1066 DVDD.n585 DVSS 0.003076f
C1067 DVDD.n586 DVSS 0.001538f
C1068 DVDD.n587 DVSS 0.001538f
C1069 DVDD.n588 DVSS 0.003076f
C1070 DVDD.n589 DVSS 0.003076f
C1071 DVDD.n590 DVSS 0.003076f
C1072 DVDD.n591 DVSS 0.003076f
C1073 DVDD.n592 DVSS 0.003076f
C1074 DVDD.n593 DVSS 0.003076f
C1075 DVDD.n594 DVSS 0.003076f
C1076 DVDD.n595 DVSS 0.003076f
C1077 DVDD.n596 DVSS 0.001538f
C1078 DVDD.n597 DVSS 0.002171f
C1079 DVDD.n598 DVSS 0.001538f
C1080 DVDD.n599 DVSS 0.00134f
C1081 DVDD.n600 DVSS 0.001538f
C1082 DVDD.n601 DVSS 0.003076f
C1083 DVDD.n602 DVSS 0.003076f
C1084 DVDD.n603 DVSS 0.017305f
C1085 DVDD.n604 DVSS 0.014092f
C1086 DVDD.n605 DVSS 0.014092f
C1087 DVDD.n606 DVSS 0.004305f
C1088 DVDD.t3 DVSS 0.013249f
C1089 DVDD.n607 DVSS 0.012648f
C1090 DVDD.t23 DVSS 0.046552f
C1091 DVDD.t57 DVSS 0.046552f
C1092 DVDD.t32 DVSS 0.046552f
C1093 DVDD.t21 DVSS 0.046552f
C1094 DVDD.t42 DVSS 0.046552f
C1095 DVDD.t68 DVSS 0.046552f
C1096 DVDD.t10 DVSS 0.046552f
C1097 DVDD.t25 DVSS 0.046552f
C1098 DVDD.t59 DVSS 0.046552f
C1099 DVDD.t30 DVSS 0.046552f
C1100 DVDD.t53 DVSS 0.046552f
C1101 DVDD.t66 DVSS 0.046552f
C1102 DVDD.t28 DVSS 0.046552f
C1103 DVDD.t50 DVSS 0.046552f
C1104 DVDD.t13 DVSS 0.03148f
C1105 DVDD.t11 DVSS 0.003225f
C1106 DVDD.t26 DVSS 0.003225f
C1107 DVDD.n608 DVSS 0.011936f
C1108 DVDD.n609 DVSS 0.010223f
C1109 DVDD.t60 DVSS 0.003225f
C1110 DVDD.t31 DVSS 0.003225f
C1111 DVDD.n610 DVSS 0.011936f
C1112 DVDD.n611 DVSS 0.010076f
C1113 DVDD.t54 DVSS 0.003225f
C1114 DVDD.t67 DVSS 0.003225f
C1115 DVDD.n612 DVSS 0.011936f
C1116 DVDD.n613 DVSS 0.010076f
C1117 DVDD.t29 DVSS 0.003225f
C1118 DVDD.t51 DVSS 0.003225f
C1119 DVDD.n614 DVSS 0.011936f
C1120 DVDD.n615 DVSS 0.010107f
C1121 DVDD.n616 DVSS 0.011769f
C1122 DVDD.t14 DVSS 0.003225f
C1123 DVDD.t16 DVSS 0.003225f
C1124 DVDD.n617 DVSS 0.011663f
C1125 DVDD.t41 DVSS 0.003225f
C1126 DVDD.t56 DVSS 0.003225f
C1127 DVDD.n618 DVSS 0.011936f
C1128 DVDD.t74 DVSS 0.003225f
C1129 DVDD.t49 DVSS 0.003225f
C1130 DVDD.n619 DVSS 0.011936f
C1131 DVDD.t35 DVSS 0.003225f
C1132 DVDD.t45 DVSS 0.003225f
C1133 DVDD.n620 DVSS 0.011936f
C1134 DVDD.t20 DVSS 0.013249f
C1135 DVDD.t65 DVSS 0.003225f
C1136 DVDD.t37 DVSS 0.003225f
C1137 DVDD.n621 DVSS 0.011663f
C1138 DVDD.t39 DVSS 0.003225f
C1139 DVDD.t47 DVSS 0.003225f
C1140 DVDD.n622 DVSS 0.011936f
C1141 DVDD.t63 DVSS 0.003225f
C1142 DVDD.t1 DVSS 0.003225f
C1143 DVDD.n623 DVSS 0.011936f
C1144 DVDD.n624 DVSS 0.010076f
C1145 DVDD.n625 DVSS 0.009654f
C1146 DVDD.n626 DVSS 0.004305f
C1147 DVDD.n627 DVSS 0.001538f
C1148 DVDD.n628 DVSS 0.027489f
C1149 DVDD.n629 DVSS 0.001538f
C1150 DVDD.n630 DVSS 0.003076f
C1151 DVDD.n631 DVSS 0.003076f
C1152 DVDD.n632 DVSS 0.003076f
C1153 DVDD.n633 DVSS 0.003076f
C1154 DVDD.n634 DVSS 0.003076f
C1155 DVDD.n635 DVSS 0.003076f
C1156 DVDD.n636 DVSS 0.003076f
C1157 DVDD.n637 DVSS 0.003076f
C1158 DVDD.n638 DVSS 0.014092f
C1159 DVDD.n639 DVSS 0.028184f
C1160 DVDD.n640 DVSS 0.028184f
C1161 DVDD.n641 DVSS 0.028184f
C1162 DVDD.n642 DVSS 0.028184f
C1163 DVDD.n643 DVSS 0.028184f
C1164 DVDD.n644 DVSS 0.016573f
C1165 DVDD.n645 DVSS 0.078941f
C1166 DVDD.n646 DVSS 0.033611f
C1167 DVDD.n647 DVSS 0.028184f
C1168 DVDD.n648 DVSS 0.028184f
C1169 DVDD.n649 DVSS 0.028184f
C1170 DVDD.n650 DVSS 0.028184f
C1171 DVDD.n651 DVSS 0.028184f
C1172 DVDD.n652 DVSS 0.028184f
C1173 DVDD.n653 DVSS 0.028184f
C1174 DVDD.n654 DVSS 0.028184f
C1175 DVDD.n655 DVSS 0.028184f
C1176 DVDD.n656 DVSS 0.040514f
C1177 DVDD.n657 DVSS 0.009229f
C1178 DVDD.n658 DVSS 0.025802f
C1179 DVDD.n659 DVSS 0.030888f
C1180 DVDD.n660 DVSS 0.052845f
C1181 DVDD.n661 DVSS 0.052845f
C1182 DVDD.n662 DVSS 0.028184f
C1183 DVDD.n663 DVSS 0.028184f
C1184 DVDD.n664 DVSS 0.028184f
C1185 DVDD.n665 DVSS 0.028184f
C1186 DVDD.n666 DVSS 0.028184f
C1187 DVDD.n667 DVSS 0.028184f
C1188 DVDD.n668 DVSS 0.028184f
C1189 DVDD.n669 DVSS 0.028184f
C1190 DVDD.n670 DVSS 0.028184f
C1191 DVDD.n671 DVSS 0.085347f
C1192 DVDD.n672 DVSS 0.03166f
C1193 DVDD.n673 DVSS 0.071557f
C1194 DVDD.n674 DVSS 0.06984f
C1195 DVDD.n675 DVSS 0.088583f
C1196 DVDD.n676 DVSS 0.024413f
C1197 DVDD.n677 DVSS 0.024413f
C1198 DVDD.n678 DVSS 0.024413f
C1199 DVDD.n679 DVSS 0.028184f
C1200 DVDD.n680 DVSS 0.028184f
C1201 DVDD.n681 DVSS 0.028184f
C1202 DVDD.n682 DVSS 0.028184f
C1203 DVDD.n683 DVSS 0.028184f
C1204 DVDD.n684 DVSS 0.028184f
C1205 DVDD.n685 DVSS 0.028184f
C1206 DVDD.n686 DVSS 0.028184f
C1207 DVDD.n687 DVSS 0.028184f
C1208 DVDD.n688 DVSS 0.028184f
C1209 DVDD.n689 DVSS 0.028184f
C1210 DVDD.n690 DVSS 0.028184f
C1211 DVDD.n691 DVSS 0.028184f
C1212 DVDD.n692 DVSS 0.028184f
C1213 DVDD.n693 DVSS 0.028184f
C1214 DVDD.n694 DVSS 0.025802f
C1215 DVDD.n695 DVSS 0.025802f
C1216 DVDD.n696 DVSS 0.026423f
C1217 DVDD.n697 DVSS 0.052845f
C1218 DVDD.n698 DVSS 0.052845f
C1219 DVDD.n699 DVSS 0.043355f
C1220 DVDD.n700 DVSS 0.003076f
C1221 DVDD.n701 DVSS 0.023631f
C1222 DVDD.n702 DVSS 0.052845f
C1223 DVDD.n703 DVSS 0.052845f
C1224 DVDD.n704 DVSS 0.052845f
C1225 DVDD.n705 DVSS 0.026423f
C1226 DVDD.n706 DVSS 0.023073f
C1227 DVDD.n707 DVSS 0.003076f
C1228 DVDD.n708 DVSS 0.023073f
C1229 DVDD.n709 DVSS 0.052845f
C1230 DVDD.n710 DVSS 0.08485f
C1231 DVDD.n711 DVSS 0.08485f
C1232 DVDD.n712 DVSS 0.026423f
C1233 DVDD.n713 DVSS 0.026423f
C1234 DVDD.n714 DVSS 0.023073f
C1235 DVDD.n715 DVSS 0.025492f
C1236 DVDD.n716 DVSS 0.003076f
C1237 DVDD.n717 DVSS 0.023073f
C1238 DVDD.n718 DVSS 0.062707f
C1239 DVDD.n719 DVSS 0.052845f
C1240 DVDD.n720 DVSS 0.040378f
C1241 DVDD.n721 DVSS 0.052845f
C1242 DVDD.n722 DVSS 0.052845f
C1243 DVDD.n723 DVSS 0.026423f
C1244 DVDD.n724 DVSS 0.024004f
C1245 DVDD.n725 DVSS 0.003076f
C1246 DVDD.n726 DVSS 0.023073f
C1247 DVDD.n727 DVSS 0.003076f
C1248 DVDD.n728 DVSS 0.023073f
C1249 DVDD.n729 DVSS 0.007613f
C1250 DVDD.n730 DVSS 0.05553f
C1251 DVDD.n731 DVSS 0.007613f
C1252 DVDD.n732 DVSS 0.023073f
C1253 DVDD.n733 DVSS 0.003076f
C1254 DVDD.n734 DVSS 0.023073f
C1255 DVDD.n735 DVSS 0.003076f
C1256 DVDD.n736 DVSS 0.023073f
C1257 DVDD.n737 DVSS 0.026423f
C1258 DVDD.n738 DVSS 0.03889f
C1259 DVDD.n739 DVSS 0.052845f
C1260 DVDD.n740 DVSS 0.053408f
C1261 DVDD.n741 DVSS 0.023073f
C1262 DVDD.n742 DVSS 0.026423f
C1263 DVDD.n743 DVSS 0.003076f
C1264 DVDD.n744 DVSS 0.001538f
C1265 DVDD.n745 DVSS 0.031819f
C1266 DVDD.n746 DVSS 0.023073f
C1267 DVDD.n747 DVSS 0.003076f
C1268 DVDD.n748 DVSS 0.003076f
C1269 DVDD.n749 DVSS 0.003076f
C1270 DVDD.n750 DVSS 0.003076f
C1271 DVDD.n751 DVSS 0.003076f
C1272 DVDD.n752 DVSS 0.003076f
C1273 DVDD.n753 DVSS 0.003076f
C1274 DVDD.n754 DVSS 0.003076f
C1275 DVDD.n755 DVSS 0.003076f
C1276 DVDD.n756 DVSS 0.003076f
C1277 DVDD.n757 DVSS 0.001538f
C1278 DVDD.n758 DVSS 0.052845f
C1279 DVDD.n759 DVSS 0.052845f
C1280 DVDD.n760 DVSS 0.052845f
C1281 DVDD.n761 DVSS 0.052845f
C1282 DVDD.n762 DVSS 0.052845f
C1283 DVDD.n763 DVSS 0.052845f
C1284 DVDD.n764 DVSS 0.052845f
C1285 DVDD.n765 DVSS 0.052845f
C1286 DVDD.n766 DVSS 0.052845f
C1287 DVDD.n767 DVSS 0.052845f
C1288 DVDD.n768 DVSS 0.052845f
C1289 DVDD.n769 DVSS 0.052845f
C1290 DVDD.n770 DVSS 0.052845f
C1291 DVDD.n771 DVSS 0.052845f
C1292 DVDD.n772 DVSS 0.052845f
C1293 DVDD.n773 DVSS 0.052845f
C1294 DVDD.n774 DVSS 0.003076f
C1295 DVDD.n775 DVSS 0.003076f
C1296 DVDD.n776 DVSS 0.003076f
C1297 DVDD.n777 DVSS 0.003076f
C1298 DVDD.n778 DVSS 0.003076f
C1299 DVDD.n779 DVSS 0.003076f
C1300 DVDD.n780 DVSS 0.003076f
C1301 DVDD.n781 DVSS 0.003076f
C1302 DVDD.n782 DVSS 0.003076f
C1303 DVDD.n783 DVSS 0.003076f
C1304 DVDD.n784 DVSS 0.026423f
C1305 DVDD.n785 DVSS 0.052845f
C1306 DVDD.n786 DVSS 0.880191f
C1307 DVDD.n787 DVSS 0.9643f
C1308 DVDD.n788 DVSS 0.018855f
C1309 DVDD.n789 DVSS 0.028184f
C1310 DVDD.n790 DVSS 0.02342f
C1311 DVDD.n791 DVSS 0.028184f
C1312 DVDD.n792 DVSS 0.028184f
C1313 DVDD.n793 DVSS 0.028184f
C1314 DVDD.n794 DVSS 0.028184f
C1315 DVDD.n795 DVSS 0.028184f
C1316 DVDD.n796 DVSS 0.028184f
C1317 DVDD.n797 DVSS 0.028184f
C1318 DVDD.n798 DVSS 0.028184f
C1319 DVDD.n799 DVSS 0.017268f
C1320 DVDD.n800 DVSS 0.017268f
C1321 DVDD.n801 DVSS 0.065184f
C1322 DVDD.n802 DVSS 0.140744f
C1323 DVDD.n803 DVSS 0.041426f
C1324 DVDD.n804 DVSS 0.065325f
C1325 DVDD.n805 DVSS 0.146476f
C1326 DVDD.n806 DVSS 0.017268f
C1327 DVDD.n807 DVSS 0.028184f
C1328 DVDD.n808 DVSS 0.028184f
C1329 DVDD.n809 DVSS 0.028184f
C1330 DVDD.n810 DVSS 0.028184f
C1331 DVDD.n811 DVSS 0.028184f
C1332 DVDD.n812 DVSS 0.028184f
C1333 DVDD.n813 DVSS 0.028184f
C1334 DVDD.n814 DVSS 0.028184f
C1335 DVDD.n815 DVSS 0.028184f
C1336 DVDD.n816 DVSS 0.028184f
C1337 DVDD.n817 DVSS 0.028184f
C1338 DVDD.n818 DVSS 0.028184f
C1339 DVDD.n819 DVSS 0.028184f
C1340 DVDD.n820 DVSS 0.028184f
C1341 DVDD.n821 DVSS 0.028184f
C1342 DVDD.n822 DVSS 0.028184f
C1343 DVDD.n823 DVSS 0.018855f
C1344 DVDD.n824 DVSS 0.028184f
C1345 DVDD.n825 DVSS 0.028184f
C1346 DVDD.n826 DVSS 0.028184f
C1347 DVDD.n827 DVSS 0.018855f
C1348 DVDD.n828 DVSS 0.706057f
C1349 DVDD.n829 DVSS 0.001538f
C1350 DVDD.n830 DVSS 0.003076f
C1351 DVDD.n831 DVSS 0.003076f
C1352 DVDD.n832 DVSS 0.003076f
C1353 DVDD.n833 DVSS 0.003076f
C1354 DVDD.n834 DVSS 0.003076f
C1355 DVDD.n835 DVSS 0.003076f
C1356 DVDD.n836 DVSS 0.003076f
C1357 DVDD.n837 DVSS 0.003076f
C1358 DVDD.n838 DVSS 0.001538f
C1359 DVDD.n839 DVSS 0.028184f
C1360 DVDD.n840 DVSS 0.028184f
C1361 DVDD.n841 DVSS 0.028184f
C1362 DVDD.n842 DVSS 0.028184f
C1363 DVDD.n843 DVSS 0.028184f
C1364 DVDD.n844 DVSS 0.028184f
C1365 DVDD.n845 DVSS 0.028184f
C1366 DVDD.n846 DVSS 0.026795f
C1367 DVDD.n847 DVSS 0.026795f
C1368 DVDD.n848 DVSS 0.018062f
C1369 DVDD.n849 DVSS 0.031815f
C1370 DVDD.n850 DVSS 0.033611f
C1371 DVDD.n851 DVSS 0.028184f
C1372 DVDD.n852 DVSS 0.028184f
C1373 DVDD.n853 DVSS 0.028184f
C1374 DVDD.n854 DVSS 0.028184f
C1375 DVDD.n855 DVSS 0.028184f
C1376 DVDD.n856 DVSS 0.028184f
C1377 DVDD.n857 DVSS 0.028184f
C1378 DVDD.n858 DVSS 0.028184f
C1379 DVDD.n859 DVSS 0.028184f
C1380 DVDD.n860 DVSS 0.018062f
C1381 DVDD.n861 DVSS 0.018062f
C1382 DVDD.n862 DVSS 0.082136f
C1383 DVDD.n863 DVSS 0.031917f
C1384 DVDD.n864 DVSS 0.078941f
C1385 DVDD.n865 DVSS 0.026795f
C1386 DVDD.n866 DVSS 0.028184f
C1387 DVDD.n867 DVSS 0.028184f
C1388 DVDD.n868 DVSS 0.028184f
C1389 DVDD.n869 DVSS 0.028184f
C1390 DVDD.n870 DVSS 0.028184f
C1391 DVDD.n871 DVSS 0.028184f
C1392 DVDD.n872 DVSS 0.028184f
C1393 DVDD.n873 DVSS 0.028184f
C1394 DVDD.n874 DVSS 0.028184f
C1395 DVDD.n875 DVSS 0.028184f
C1396 DVDD.n876 DVSS 0.028184f
C1397 DVDD.n877 DVSS 0.028184f
C1398 DVDD.n878 DVSS 0.028184f
C1399 DVDD.n879 DVSS 0.028184f
C1400 DVDD.n880 DVSS 0.022726f
C1401 DVDD.n881 DVSS 0.001538f
C1402 DVDD.n882 DVSS 0.031074f
C1403 DVDD.n883 DVSS 0.002593f
C1404 DVDD.n884 DVSS 0.002493f
C1405 DVDD.n885 DVSS 0.001538f
C1406 DVDD.n886 DVSS 0.00134f
C1407 DVDD.n887 DVSS 0.023073f
C1408 DVDD.n888 DVSS 0.003076f
C1409 DVDD.n889 DVSS 0.001538f
C1410 DVDD.n890 DVSS 0.003076f
C1411 DVDD.n891 DVSS 0.003076f
C1412 DVDD.n892 DVSS 0.003076f
C1413 DVDD.n893 DVSS 0.003076f
C1414 DVDD.n894 DVSS 0.002121f
C1415 DVDD.n895 DVSS 0.003076f
C1416 DVDD.n896 DVSS 0.002022f
C1417 DVDD.n898 DVSS 0.002394f
C1418 DVDD.n899 DVSS 0.004999f
C1419 DVDD.n900 DVSS 0.001538f
C1420 DVDD.n901 DVSS 0.031819f
C1421 DVDD.n902 DVSS 0.00289f
C1422 DVDD.n903 DVSS 0.002791f
C1423 DVDD.n904 DVSS 0.002692f
C1424 DVDD.n905 DVSS 0.002593f
C1425 DVDD.n906 DVSS 0.002493f
C1426 DVDD.n907 DVSS 0.023073f
C1427 DVDD.n908 DVSS 0.003076f
C1428 DVDD.n909 DVSS 0.002121f
C1429 DVDD.n910 DVSS 0.003076f
C1430 DVDD.n911 DVSS 0.002022f
C1431 DVDD.n912 DVSS 0.003076f
C1432 DVDD.n913 DVSS 0.001923f
C1433 DVDD.n914 DVSS 0.003076f
C1434 DVDD.n915 DVSS 0.001824f
C1435 DVDD.n916 DVSS 0.003076f
C1436 DVDD.n917 DVSS 0.001724f
C1437 DVDD.n918 DVSS 0.003076f
C1438 DVDD.n919 DVSS 0.001538f
C1439 DVDD.n920 DVSS 0.027687f
C1440 DVDD.n922 DVSS 0.031819f
C1441 DVDD.n923 DVSS 0.001538f
C1442 DVDD.n924 DVSS 0.00299f
C1443 DVDD.n925 DVSS 0.00289f
C1444 DVDD.n926 DVSS 0.002791f
C1445 DVDD.n927 DVSS 0.023073f
C1446 DVDD.n928 DVSS 0.001824f
C1447 DVDD.n929 DVSS 0.003076f
C1448 DVDD.n930 DVSS 0.003076f
C1449 DVDD.n931 DVSS 0.003076f
C1450 DVDD.n932 DVSS 0.003076f
C1451 DVDD.n933 DVSS 0.003076f
C1452 DVDD.n934 DVSS 0.001724f
C1453 DVDD.n935 DVSS 0.003076f
C1454 DVDD.n936 DVSS 0.001625f
C1455 DVDD.n937 DVSS 0.001538f
C1456 DVDD.n938 DVSS 0.001538f
C1457 DVDD.n939 DVSS 0.003064f
C1458 DVDD.n940 DVSS 0.050798f
C1459 DVDD.n941 DVSS 0.001538f
C1460 DVDD.n942 DVSS 0.003076f
C1461 DVDD.n943 DVSS 0.003076f
C1462 DVDD.n944 DVSS 0.003076f
C1463 DVDD.n945 DVSS 0.003076f
C1464 DVDD.n946 DVSS 0.001538f
C1465 DVDD.n947 DVSS 0.001538f
C1466 DVDD.n948 DVSS 0.001538f
C1467 DVDD.n949 DVSS 0.001538f
C1468 DVDD.n950 DVSS 0.027687f
C1469 DVDD.n951 DVSS 0.001538f
C1470 DVDD.n952 DVSS 0.031819f
C1471 DVDD.n953 DVSS 0.001538f
C1472 DVDD.n954 DVSS 0.001538f
C1473 DVDD.n955 DVSS 0.001538f
C1474 DVDD.n956 DVSS 0.002965f
C1475 DVDD.n957 DVSS 0.003076f
C1476 DVDD.n958 DVSS 0.00299f
C1477 DVDD.n959 DVSS 0.023073f
C1478 DVDD.n960 DVSS 0.003076f
C1479 DVDD.n961 DVSS 0.001625f
C1480 DVDD.n962 DVSS 0.001538f
C1481 DVDD.n963 DVSS 0.001551f
C1482 DVDD.n964 DVSS 0.001538f
C1483 DVDD.n965 DVSS 0.001538f
C1484 DVDD.n966 DVSS 0.002667f
C1485 DVDD.n967 DVSS 0.002766f
C1486 DVDD.n968 DVSS 0.002866f
C1487 DVDD.n969 DVSS 0.001538f
C1488 DVDD.n970 DVSS 0.001538f
C1489 DVDD.n971 DVSS 0.003064f
C1490 DVDD.n972 DVSS 0.050798f
C1491 DVDD.n973 DVSS 0.001538f
C1492 DVDD.n974 DVSS 0.001538f
C1493 DVDD.n975 DVSS 0.00165f
C1494 DVDD.n976 DVSS 0.003076f
C1495 DVDD.t131 DVSS 0.032253f
C1496 DVDD.t141 DVSS 0.032253f
C1497 DVDD.n977 DVSS 0.064506f
C1498 DVDD.n978 DVSS 0.00768f
C1499 DVDD.n979 DVSS 0.004688f
C1500 DVDD.n980 DVSS 0.002866f
C1501 DVDD.n981 DVSS 0.001538f
C1502 DVDD.n982 DVSS 0.023073f
C1503 DVDD.n983 DVSS 0.002667f
C1504 DVDD.n984 DVSS 0.002766f
C1505 DVDD.n985 DVSS 0.001538f
C1506 DVDD.n986 DVSS 0.001538f
C1507 DVDD.n987 DVSS 0.003064f
C1508 DVDD.n988 DVSS 0.017305f
C1509 DVDD.n989 DVSS 0.001538f
C1510 DVDD.n990 DVSS 0.001538f
C1511 DVDD.n991 DVSS 0.001538f
C1512 DVDD.n992 DVSS 0.00165f
C1513 DVDD.n993 DVSS 0.003076f
C1514 DVDD.n994 DVSS 0.003076f
C1515 DVDD.n995 DVSS 0.001848f
C1516 DVDD.n996 DVSS 0.003076f
C1517 DVDD.n997 DVSS 0.008261f
C1518 DVDD.n998 DVSS 0.001538f
C1519 DVDD.n999 DVSS 0.001538f
C1520 DVDD.n1000 DVSS 0.003076f
C1521 DVDD.n1001 DVSS 0.003076f
C1522 DVDD.n1002 DVSS 0.001538f
C1523 DVDD.n1003 DVSS 0.001538f
C1524 DVDD.n1004 DVSS 0.001538f
C1525 DVDD.n1005 DVSS 0.001538f
C1526 DVDD.n1006 DVSS 0.026423f
C1527 DVDD.n1007 DVSS 0.027944f
C1528 DVDD.n1008 DVSS 0.001538f
C1529 DVDD.n1009 DVSS 0.027687f
C1530 DVDD.n1010 DVSS 0.01188f
C1531 DVDD.n1011 DVSS 0.027944f
C1532 DVDD.t143 DVSS 0.032253f
C1533 DVDD.t86 DVSS 0.032253f
C1534 DVDD.n1012 DVSS 0.064506f
C1535 DVDD.n1013 DVSS 0.011628f
C1536 DVDD.n1014 DVSS 0.004122f
C1537 DVDD.n1015 DVSS 0.024376f
C1538 DVDD.n1016 DVSS 0.026423f
C1539 DVDD.n1017 DVSS 0.02512f
C1540 DVDD.n1018 DVSS 0.023073f
C1541 DVDD.n1019 DVSS 0.007148f
C1542 DVDD.n1021 DVSS 0.008245f
C1543 DVDD.n1023 DVSS 0.008245f
C1544 DVDD.n1024 DVSS 0.007414f
C1545 DVDD.n1027 DVSS 0.008245f
C1546 DVDD.n1029 DVSS 0.008245f
C1547 DVDD.n1031 DVSS 0.008245f
C1548 DVDD.n1033 DVSS 0.008245f
C1549 DVDD.n1034 DVSS 0.007946f
C1550 DVDD.n1036 DVSS 0.008245f
C1551 DVDD.n1038 DVSS 0.008012f
C1552 DVDD.n1040 DVSS 0.008245f
C1553 DVDD.n1042 DVSS 0.007746f
C1554 DVDD.n1043 DVSS 0.052845f
C1555 DVDD.n1044 DVSS 0.052845f
C1556 DVDD.n1045 DVSS 0.052845f
C1557 DVDD.n1046 DVSS 0.052845f
C1558 DVDD.n1047 DVSS 0.052845f
C1559 DVDD.n1048 DVSS 0.052845f
C1560 DVDD.n1049 DVSS 0.052845f
C1561 DVDD.n1050 DVSS 0.052845f
C1562 DVDD.n1051 DVSS 0.052845f
C1563 DVDD.n1052 DVSS 0.052845f
C1564 DVDD.n1053 DVSS 0.052845f
C1565 DVDD.n1054 DVSS 0.052845f
C1566 DVDD.n1055 DVSS 0.052845f
C1567 DVDD.n1056 DVSS 0.052845f
C1568 DVDD.n1057 DVSS 0.052845f
C1569 DVDD.n1058 DVSS 0.052845f
C1570 DVDD.n1059 DVSS 0.032377f
C1571 DVDD.n1060 DVSS 0.063637f
C1572 DVDD.n1061 DVSS 0.046891f
C1573 DVDD.n1062 DVSS 0.100852f
C1574 DVDD.n1063 DVSS 0.032377f
C1575 DVDD.n1064 DVSS 0.052845f
C1576 DVDD.n1065 DVSS 0.100852f
C1577 DVDD.n1066 DVSS 0.046891f
C1578 DVDD.n1067 DVSS 0.052845f
C1579 DVDD.n1068 DVSS 0.052845f
C1580 DVDD.n1069 DVSS 0.052845f
C1581 DVDD.n1070 DVSS 0.052845f
C1582 DVDD.n1071 DVSS 0.052845f
C1583 DVDD.n1072 DVSS 0.052845f
C1584 DVDD.n1073 DVSS 0.052845f
C1585 DVDD.n1074 DVSS 0.052845f
C1586 DVDD.n1075 DVSS 0.052845f
C1587 DVDD.n1076 DVSS 0.052845f
C1588 DVDD.n1077 DVSS 0.052845f
C1589 DVDD.n1078 DVSS 0.052845f
C1590 DVDD.n1079 DVSS 0.052845f
C1591 DVDD.n1080 DVSS 0.052845f
C1592 DVDD.n1081 DVSS 0.052845f
C1593 DVDD.n1082 DVSS 0.052845f
C1594 DVDD.n1083 DVSS 0.052845f
C1595 DVDD.n1084 DVSS 0.052845f
C1596 DVDD.n1085 DVSS 0.052845f
C1597 DVDD.n1086 DVSS 0.052845f
C1598 DVDD.n1087 DVSS 0.052845f
C1599 DVDD.n1088 DVSS 0.052845f
C1600 DVDD.n1089 DVSS 0.052845f
C1601 DVDD.n1090 DVSS 0.052845f
C1602 DVDD.n1091 DVSS 0.052845f
C1603 DVDD.n1092 DVSS 0.052845f
C1604 DVDD.n1093 DVSS 0.026423f
C1605 DVDD.n1094 DVSS 0.052845f
C1606 DVDD.n1095 DVSS 0.052845f
C1607 DVDD.n1096 DVSS 0.052845f
C1608 DVDD.n1097 DVSS 0.030888f
C1609 DVDD.n1098 DVSS 0.001538f
C1610 DVDD.n1099 DVSS 0.003064f
C1611 DVDD.n1100 DVSS 0.017305f
C1612 DVDD.n1102 DVSS 0.001538f
C1613 DVDD.n1103 DVSS 0.003076f
C1614 DVDD.n1104 DVSS 0.003076f
C1615 DVDD.n1105 DVSS 0.003076f
C1616 DVDD.n1106 DVSS 0.003076f
C1617 DVDD.n1107 DVSS 0.003076f
C1618 DVDD.n1108 DVSS 0.003076f
C1619 DVDD.n1109 DVSS 0.003076f
C1620 DVDD.n1110 DVSS 0.003076f
C1621 DVDD.n1111 DVSS 0.003076f
C1622 DVDD.n1112 DVSS 0.001538f
C1623 DVDD.n1113 DVSS 0.001538f
C1624 DVDD.n1114 DVSS 0.003076f
C1625 DVDD.n1115 DVSS 0.001538f
C1626 DVDD.n1116 DVSS 0.001538f
C1627 DVDD.n1117 DVSS 0.001625f
C1628 DVDD.n1118 DVSS 0.001538f
C1629 DVDD.n1119 DVSS 0.004122f
C1630 DVDD.n1120 DVSS 0.001538f
C1631 DVDD.n1121 DVSS 0.001625f
C1632 DVDD.n1122 DVSS 0.001538f
C1633 DVDD.n1123 DVSS 0.031074f
C1634 DVDD.n1124 DVSS 0.001538f
C1635 DVDD.n1125 DVSS 0.00289f
C1636 DVDD.n1126 DVSS 0.002791f
C1637 DVDD.n1127 DVSS 0.005768f
C1638 DVDD.n1128 DVSS 0.023073f
C1639 DVDD.n1129 DVSS 0.001824f
C1640 DVDD.n1130 DVSS 0.003076f
C1641 DVDD.n1131 DVSS 0.003076f
C1642 DVDD.n1132 DVSS 0.003076f
C1643 DVDD.n1133 DVSS 0.003076f
C1644 DVDD.n1134 DVSS 0.003076f
C1645 DVDD.n1135 DVSS 0.001724f
C1646 DVDD.n1136 DVSS 0.003076f
C1647 DVDD.n1137 DVSS 0.001538f
C1648 DVDD.n1138 DVSS 0.008262f
C1649 DVDD.n1139 DVSS 0.003064f
C1650 DVDD.n1140 DVSS 0.052845f
C1651 DVDD.n1141 DVSS 0.052845f
C1652 DVDD.n1142 DVSS 0.052845f
C1653 DVDD.n1143 DVSS 0.052845f
C1654 DVDD.n1144 DVSS 0.052845f
C1655 DVDD.n1145 DVSS 0.052845f
C1656 DVDD.n1146 DVSS 0.052845f
C1657 DVDD.n1147 DVSS 0.052845f
C1658 DVDD.n1148 DVSS 0.052845f
C1659 DVDD.n1149 DVSS 0.052845f
C1660 DVDD.n1150 DVSS 0.052845f
C1661 DVDD.n1151 DVSS 0.052845f
C1662 DVDD.n1152 DVSS 0.052845f
C1663 DVDD.n1153 DVSS 0.052845f
C1664 DVDD.n1154 DVSS 0.052845f
C1665 DVDD.n1155 DVSS 0.052845f
C1666 DVDD.n1156 DVSS 0.052845f
C1667 DVDD.n1157 DVSS 0.052845f
C1668 DVDD.n1158 DVSS 0.052845f
C1669 DVDD.n1159 DVSS 0.052845f
C1670 DVDD.n1160 DVSS 0.052845f
C1671 DVDD.n1161 DVSS 0.052845f
C1672 DVDD.n1162 DVSS 0.052845f
C1673 DVDD.n1163 DVSS 0.052845f
C1674 DVDD.n1164 DVSS 0.052845f
C1675 DVDD.n1165 DVSS 0.052845f
C1676 DVDD.n1166 DVSS 0.052845f
C1677 DVDD.n1167 DVSS 0.052845f
C1678 DVDD.n1168 DVSS 0.033866f
C1679 DVDD.n1169 DVSS 0.052845f
C1680 DVDD.n1170 DVSS 0.052845f
C1681 DVDD.n1171 DVSS 0.033866f
C1682 DVDD.n1172 DVSS 0.063637f
C1683 DVDD.n1173 DVSS 0.100852f
C1684 DVDD.n1174 DVSS 0.045402f
C1685 DVDD.n1175 DVSS 0.052845f
C1686 DVDD.n1176 DVSS 0.100852f
C1687 DVDD.n1177 DVSS 0.052845f
C1688 DVDD.n1178 DVSS 0.052845f
C1689 DVDD.n1179 DVSS 0.052845f
C1690 DVDD.n1180 DVSS 0.052845f
C1691 DVDD.n1181 DVSS 0.052845f
C1692 DVDD.n1182 DVSS 0.052845f
C1693 DVDD.n1183 DVSS 0.052845f
C1694 DVDD.n1184 DVSS 0.052845f
C1695 DVDD.n1185 DVSS 0.052845f
C1696 DVDD.n1186 DVSS 0.052845f
C1697 DVDD.n1187 DVSS 0.052845f
C1698 DVDD.n1188 DVSS 0.052845f
C1699 DVDD.n1189 DVSS 0.026423f
C1700 DVDD.n1190 DVSS 0.052845f
C1701 DVDD.n1191 DVSS 0.052845f
C1702 DVDD.n1192 DVSS 0.052845f
C1703 DVDD.n1193 DVSS 0.052845f
C1704 DVDD.n1207 DVSS 0.01188f
C1705 DVDD.t119 DVSS 0.032253f
C1706 DVDD.t151 DVSS 0.032253f
C1707 DVDD.n1208 DVSS 0.064506f
C1708 DVDD.n1209 DVSS 0.011628f
C1709 DVDD.n1210 DVSS 0.011569f
C1710 DVDD.n1211 DVSS 0.008245f
C1711 DVDD.n1212 DVSS 0.008012f
C1712 DVDD.n1213 DVSS 0.008245f
C1713 DVDD.n1214 DVSS 0.007746f
C1714 DVDD.n1215 DVSS 0.008245f
C1715 DVDD.n1216 DVSS 0.008245f
C1716 DVDD.n1217 DVSS 0.008245f
C1717 DVDD.n1218 DVSS 0.008245f
C1718 DVDD.n1219 DVSS 0.008245f
C1719 DVDD.n1220 DVSS 0.00748f
C1720 DVDD.n1221 DVSS 0.015459f
C1721 DVDD.n1222 DVSS 0.023073f
C1722 DVDD.n1223 DVSS 0.001538f
C1723 DVDD.n1224 DVSS 0.008262f
C1724 DVDD.n1225 DVSS 0.027687f
C1725 DVDD.n1226 DVSS 0.01188f
C1726 DVDD.n1227 DVSS 0.001824f
C1727 DVDD.n1228 DVSS 0.002791f
C1728 DVDD.n1229 DVSS 0.008261f
C1729 DVDD.n1230 DVSS 0.001538f
C1730 DVDD.n1231 DVSS 0.027944f
C1731 DVDD.t112 DVSS 0.032253f
C1732 DVDD.t132 DVSS 0.032253f
C1733 DVDD.n1232 DVSS 0.064506f
C1734 DVDD.n1233 DVSS 0.011628f
C1735 DVDD.n1234 DVSS 0.004122f
C1736 DVDD.n1235 DVSS 0.004887f
C1737 DVDD.n1236 DVSS 0.008245f
C1738 DVDD.n1237 DVSS 0.008245f
C1739 DVDD.n1238 DVSS 0.008245f
C1740 DVDD.n1239 DVSS 0.008245f
C1741 DVDD.n1240 DVSS 0.008245f
C1742 DVDD.n1241 DVSS 0.001538f
C1743 DVDD.n1242 DVSS 0.008262f
C1744 DVDD.n1243 DVSS 0.027687f
C1745 DVDD.n1244 DVSS 0.01188f
C1746 DVDD.n1245 DVSS 0.001724f
C1747 DVDD.n1246 DVSS 0.00289f
C1748 DVDD.n1247 DVSS 0.008261f
C1749 DVDD.n1248 DVSS 0.001538f
C1750 DVDD.n1249 DVSS 0.027944f
C1751 DVDD.t126 DVSS 0.032253f
C1752 DVDD.t78 DVSS 0.032253f
C1753 DVDD.n1250 DVSS 0.064506f
C1754 DVDD.n1251 DVSS 0.011628f
C1755 DVDD.n1252 DVSS 0.004122f
C1756 DVDD.n1253 DVSS 0.004621f
C1757 DVDD.n1254 DVSS 0.008245f
C1758 DVDD.n1255 DVSS 0.004355f
C1759 DVDD.n1256 DVSS 0.008245f
C1760 DVDD.n1257 DVSS 0.027687f
C1761 DVDD.n1258 DVSS 0.01188f
C1762 DVDD.n1259 DVSS 0.001551f
C1763 DVDD.n1260 DVSS 0.008261f
C1764 DVDD.n1261 DVSS 0.027944f
C1765 DVDD.t76 DVSS 0.032253f
C1766 DVDD.t90 DVSS 0.032253f
C1767 DVDD.n1262 DVSS 0.064506f
C1768 DVDD.n1263 DVSS 0.011628f
C1769 DVDD.n1264 DVSS 0.004122f
C1770 DVDD.n1265 DVSS 0.008212f
C1771 DVDD.n1273 DVSS 0.052845f
C1772 DVDD.n1274 DVSS 0.052845f
C1773 DVDD.n1275 DVSS 0.052845f
C1774 DVDD.n1276 DVSS 0.052845f
C1775 DVDD.n1277 DVSS 0.052845f
C1776 DVDD.n1278 DVSS 0.052845f
C1777 DVDD.n1279 DVSS 0.052845f
C1778 DVDD.n1280 DVSS 0.052845f
C1779 DVDD.n1281 DVSS 0.052845f
C1780 DVDD.n1282 DVSS 0.052845f
C1781 DVDD.n1283 DVSS 0.052845f
C1782 DVDD.n1284 DVSS 0.052845f
C1783 DVDD.n1285 DVSS 0.052845f
C1784 DVDD.n1286 DVSS 0.052845f
C1785 DVDD.n1287 DVSS 0.052845f
C1786 DVDD.n1288 DVSS 0.052845f
C1787 DVDD.n1289 DVSS 0.100852f
C1788 DVDD.n1290 DVSS 0.052845f
C1789 DVDD.n1291 DVSS 0.052845f
C1790 DVDD.n1292 DVSS 0.052845f
C1791 DVDD.n1293 DVSS 0.052845f
C1792 DVDD.n1294 DVSS 0.052845f
C1793 DVDD.n1295 DVSS 0.052845f
C1794 DVDD.n1296 DVSS 0.052845f
C1795 DVDD.n1297 DVSS 0.052845f
C1796 DVDD.n1298 DVSS 0.052845f
C1797 DVDD.n1299 DVSS 0.052845f
C1798 DVDD.n1300 DVSS 0.052845f
C1799 DVDD.n1301 DVSS 0.052845f
C1800 DVDD.n1302 DVSS 0.052845f
C1801 DVDD.n1303 DVSS 0.052845f
C1802 DVDD.n1304 DVSS 0.052845f
C1803 DVDD.n1305 DVSS 0.052845f
C1804 DVDD.n1306 DVSS 0.052845f
C1805 DVDD.n1307 DVSS 0.052845f
C1806 DVDD.n1308 DVSS 0.052845f
C1807 DVDD.n1309 DVSS 0.052845f
C1808 DVDD.n1310 DVSS 0.052845f
C1809 DVDD.n1311 DVSS 0.052845f
C1810 DVDD.n1312 DVSS 0.052845f
C1811 DVDD.n1313 DVSS 0.052845f
C1812 DVDD.n1314 DVSS 0.052845f
C1813 DVDD.n1315 DVSS 0.052845f
C1814 DVDD.n1316 DVSS 0.052845f
C1815 DVDD.n1317 DVSS 0.052845f
C1816 DVDD.n1318 DVSS 0.052845f
C1817 DVDD.n1319 DVSS 0.052845f
C1818 DVDD.n1320 DVSS 0.030888f
C1819 DVDD.n1321 DVSS 0.100852f
C1820 DVDD.n1322 DVSS 0.048379f
C1821 DVDD.n1323 DVSS 0.052845f
C1822 DVDD.n1324 DVSS 0.048379f
C1823 DVDD.n1325 DVSS 0.063637f
C1824 DVDD.n1326 DVSS 0.017305f
C1825 DVDD.n1327 DVSS 0.052845f
C1826 DVDD.n1328 DVSS 0.100852f
C1827 DVDD.n1329 DVSS 0.063637f
C1828 DVDD.n1330 DVSS 0.063637f
C1829 DVDD.n1331 DVSS 0.030888f
C1830 DVDD.n1332 DVSS 0.052845f
C1831 DVDD.n1333 DVSS 0.052845f
C1832 DVDD.n1334 DVSS 0.052845f
C1833 DVDD.n1335 DVSS 0.052845f
C1834 DVDD.n1336 DVSS 0.052845f
C1835 DVDD.n1337 DVSS 0.052845f
C1836 DVDD.n1338 DVSS 0.052845f
C1837 DVDD.n1339 DVSS 0.052845f
C1838 DVDD.n1340 DVSS 0.052845f
C1839 DVDD.n1341 DVSS 0.052845f
C1840 DVDD.n1342 DVSS 0.052845f
C1841 DVDD.n1343 DVSS 0.052845f
C1842 DVDD.n1344 DVSS 0.052845f
C1843 DVDD.n1345 DVSS 0.047635f
C1844 DVDD.n1346 DVSS 0.047635f
C1845 DVDD.n1347 DVSS 0.005954f
C1846 DVDD.n1348 DVSS 0.075079f
C1847 DVDD.n1349 DVSS 0.243482f
C1848 DVDD.n1350 DVSS 0.047635f
C1849 DVDD.n1351 DVSS 0.052845f
C1850 DVDD.n1352 DVSS 0.052845f
C1851 DVDD.n1353 DVSS 0.052845f
C1852 DVDD.n1354 DVSS 0.052845f
C1853 DVDD.n1355 DVSS 0.052845f
C1854 DVDD.n1356 DVSS 0.052845f
C1855 DVDD.n1357 DVSS 0.052845f
C1856 DVDD.n1358 DVSS 0.052845f
C1857 DVDD.n1359 DVSS 0.052845f
C1858 DVDD.n1360 DVSS 0.052845f
C1859 DVDD.n1361 DVSS 0.052845f
C1860 DVDD.n1362 DVSS 0.052845f
C1861 DVDD.n1363 DVSS 0.052845f
C1862 DVDD.n1364 DVSS 0.052845f
C1863 DVDD.n1365 DVSS 0.048379f
C1864 DVDD.n1366 DVSS 0.048379f
C1865 DVDD.n1367 DVSS 0.100852f
C1866 DVDD.n1368 DVSS 0.052845f
C1867 DVDD.n1369 DVSS 0.052845f
C1868 DVDD.n1370 DVSS 0.026423f
C1869 DVDD.n1371 DVSS 0.002394f
C1870 DVDD.n1372 DVSS 0.001538f
C1871 DVDD.n1373 DVSS 0.003076f
C1872 DVDD.n1374 DVSS 0.001538f
C1873 DVDD.n1375 DVSS 0.001538f
C1874 DVDD.n1376 DVSS 0.003076f
C1875 DVDD.n1377 DVSS 0.001538f
C1876 DVDD.n1378 DVSS 0.001538f
C1877 DVDD.n1379 DVSS 0.003076f
C1878 DVDD.n1380 DVSS 0.001538f
C1879 DVDD.n1381 DVSS 0.001538f
C1880 DVDD.n1382 DVSS 0.003076f
C1881 DVDD.n1383 DVSS 0.001538f
C1882 DVDD.n1384 DVSS 0.001538f
C1883 DVDD.n1385 DVSS 0.003076f
C1884 DVDD.n1386 DVSS 0.001538f
C1885 DVDD.n1387 DVSS 0.001724f
C1886 DVDD.n1388 DVSS 0.001538f
C1887 DVDD.n1389 DVSS 0.004122f
C1888 DVDD.n1390 DVSS 0.001538f
C1889 DVDD.n1391 DVSS 0.001724f
C1890 DVDD.n1392 DVSS 0.001538f
C1891 DVDD.n1393 DVSS 0.031074f
C1892 DVDD.n1394 DVSS 0.002791f
C1893 DVDD.n1395 DVSS 0.002692f
C1894 DVDD.n1396 DVSS 0.002593f
C1895 DVDD.n1397 DVSS 0.002493f
C1896 DVDD.n1398 DVSS 0.023073f
C1897 DVDD.n1399 DVSS 0.003076f
C1898 DVDD.n1400 DVSS 0.002121f
C1899 DVDD.n1401 DVSS 0.003076f
C1900 DVDD.n1402 DVSS 0.002022f
C1901 DVDD.n1403 DVSS 0.003076f
C1902 DVDD.n1404 DVSS 0.001923f
C1903 DVDD.n1405 DVSS 0.003076f
C1904 DVDD.n1406 DVSS 0.001824f
C1905 DVDD.n1407 DVSS 0.003076f
C1906 DVDD.n1408 DVSS 0.003076f
C1907 DVDD.n1409 DVSS 0.052845f
C1908 DVDD.n1410 DVSS 0.052845f
C1909 DVDD.n1411 DVSS 0.052845f
C1910 DVDD.n1412 DVSS 0.052845f
C1911 DVDD.n1413 DVSS 0.052845f
C1912 DVDD.n1414 DVSS 0.052845f
C1913 DVDD.n1415 DVSS 0.052845f
C1914 DVDD.n1416 DVSS 0.052845f
C1915 DVDD.n1417 DVSS 0.052845f
C1916 DVDD.n1418 DVSS 0.052845f
C1917 DVDD.n1419 DVSS 0.052845f
C1918 DVDD.n1420 DVSS 0.052845f
C1919 DVDD.n1421 DVSS 0.052845f
C1920 DVDD.n1422 DVSS 0.052845f
C1921 DVDD.n1423 DVSS 0.052845f
C1922 DVDD.n1424 DVSS 0.052845f
C1923 DVDD.n1425 DVSS 0.052845f
C1924 DVDD.n1426 DVSS 0.052845f
C1925 DVDD.n1427 DVSS 0.052845f
C1926 DVDD.n1428 DVSS 0.052845f
C1927 DVDD.n1429 DVSS 0.052845f
C1928 DVDD.n1430 DVSS 0.052845f
C1929 DVDD.n1431 DVSS 0.052845f
C1930 DVDD.n1432 DVSS 0.052845f
C1931 DVDD.n1433 DVSS 0.052845f
C1932 DVDD.n1434 DVSS 0.052845f
C1933 DVDD.n1435 DVSS 0.052845f
C1934 DVDD.n1436 DVSS 0.001538f
C1935 DVDD.n1437 DVSS 0.001538f
C1936 DVDD.n1438 DVSS 0.001538f
C1937 DVDD.n1439 DVSS 0.001538f
C1938 DVDD.n1440 DVSS 0.001538f
C1939 DVDD.n1441 DVSS 0.001538f
C1940 DVDD.n1442 DVSS 0.001538f
C1941 DVDD.n1443 DVSS 0.001538f
C1942 DVDD.n1444 DVSS 0.001538f
C1943 DVDD.n1445 DVSS 0.001538f
C1944 DVDD.n1446 DVSS 0.026423f
C1945 DVDD.n1447 DVSS 0.052845f
C1946 DVDD.n1448 DVSS 0.052845f
C1947 DVDD.n1449 DVSS 0.052845f
C1948 DVDD.n1450 DVSS 0.052845f
C1949 DVDD.n1451 DVSS 0.033866f
C1950 DVDD.n1452 DVSS 0.063637f
C1951 DVDD.n1453 DVSS 0.052845f
C1952 DVDD.n1454 DVSS 0.045402f
C1953 DVDD.n1455 DVSS 0.052845f
C1954 DVDD.n1456 DVSS 0.052845f
C1955 DVDD.n1457 DVSS 0.052845f
C1956 DVDD.n1458 DVSS 0.052845f
C1957 DVDD.n1459 DVSS 0.052845f
C1958 DVDD.n1460 DVSS 0.052845f
C1959 DVDD.n1461 DVSS 0.052845f
C1960 DVDD.n1462 DVSS 0.052845f
C1961 DVDD.n1463 DVSS 0.052845f
C1962 DVDD.n1464 DVSS 0.052845f
C1963 DVDD.n1465 DVSS 0.052845f
C1964 DVDD.n1466 DVSS 0.052845f
C1965 DVDD.n1467 DVSS 0.052845f
C1966 DVDD.n1468 DVSS 0.052845f
C1967 DVDD.n1469 DVSS 0.052845f
C1968 DVDD.n1470 DVSS 0.008245f
C1969 DVDD.n1471 DVSS 0.007746f
C1970 DVDD.n1472 DVSS 0.008245f
C1971 DVDD.n1473 DVSS 0.00748f
C1972 DVDD.n1474 DVSS 0.008245f
C1973 DVDD.n1475 DVSS 0.007214f
C1974 DVDD.n1476 DVSS 0.008245f
C1975 DVDD.n1477 DVSS 0.006948f
C1976 DVDD.n1478 DVSS 0.008245f
C1977 DVDD.n1479 DVSS 0.006682f
C1978 DVDD.n1480 DVSS 0.008245f
C1979 DVDD.n1481 DVSS 0.023073f
C1980 DVDD.n1482 DVSS 0.008245f
C1981 DVDD.n1483 DVSS 0.001538f
C1982 DVDD.n1484 DVSS 0.008262f
C1983 DVDD.n1485 DVSS 0.027687f
C1984 DVDD.n1486 DVSS 0.01188f
C1985 DVDD.n1487 DVSS 0.002121f
C1986 DVDD.n1488 DVSS 0.002493f
C1987 DVDD.n1489 DVSS 0.008261f
C1988 DVDD.n1490 DVSS 0.001538f
C1989 DVDD.n1491 DVSS 0.027944f
C1990 DVDD.t89 DVSS 0.032253f
C1991 DVDD.t77 DVSS 0.032253f
C1992 DVDD.n1492 DVSS 0.064506f
C1993 DVDD.n1493 DVSS 0.011628f
C1994 DVDD.n1494 DVSS 0.004122f
C1995 DVDD.n1495 DVSS 0.005685f
C1996 DVDD.n1496 DVSS 0.008245f
C1997 DVDD.n1497 DVSS 0.001538f
C1998 DVDD.n1498 DVSS 0.008262f
C1999 DVDD.n1499 DVSS 0.027687f
C2000 DVDD.n1500 DVSS 0.01188f
C2001 DVDD.n1501 DVSS 0.002022f
C2002 DVDD.n1502 DVSS 0.002593f
C2003 DVDD.n1503 DVSS 0.008261f
C2004 DVDD.n1504 DVSS 0.001538f
C2005 DVDD.n1505 DVSS 0.027944f
C2006 DVDD.t136 DVSS 0.032253f
C2007 DVDD.t92 DVSS 0.032253f
C2008 DVDD.n1506 DVSS 0.064506f
C2009 DVDD.n1507 DVSS 0.011628f
C2010 DVDD.n1508 DVSS 0.004122f
C2011 DVDD.n1509 DVSS 0.005419f
C2012 DVDD.n1510 DVSS 0.008245f
C2013 DVDD.n1511 DVSS 0.001538f
C2014 DVDD.n1512 DVSS 0.008262f
C2015 DVDD.n1513 DVSS 0.027687f
C2016 DVDD.n1514 DVSS 0.01188f
C2017 DVDD.n1515 DVSS 0.001923f
C2018 DVDD.n1516 DVSS 0.002692f
C2019 DVDD.n1517 DVSS 0.008261f
C2020 DVDD.n1518 DVSS 0.001538f
C2021 DVDD.n1519 DVSS 0.027944f
C2022 DVDD.t146 DVSS 0.032253f
C2023 DVDD.t145 DVSS 0.032253f
C2024 DVDD.n1520 DVSS 0.064506f
C2025 DVDD.n1521 DVSS 0.011628f
C2026 DVDD.n1522 DVSS 0.004122f
C2027 DVDD.n1523 DVSS 0.005153f
C2028 DVDD.n1524 DVSS 0.008245f
C2029 DVDD.n1525 DVSS 0.001538f
C2030 DVDD.n1526 DVSS 0.008262f
C2031 DVDD.n1527 DVSS 0.027687f
C2032 DVDD.n1528 DVSS 0.01188f
C2033 DVDD.n1529 DVSS 0.001824f
C2034 DVDD.n1530 DVSS 0.002791f
C2035 DVDD.n1531 DVSS 0.008261f
C2036 DVDD.n1532 DVSS 0.001538f
C2037 DVDD.n1533 DVSS 0.027944f
C2038 DVDD.t135 DVSS 0.032253f
C2039 DVDD.t104 DVSS 0.032253f
C2040 DVDD.n1534 DVSS 0.064506f
C2041 DVDD.n1535 DVSS 0.011628f
C2042 DVDD.n1536 DVSS 0.004122f
C2043 DVDD.n1537 DVSS 0.004887f
C2044 DVDD.n1538 DVSS 0.008245f
C2045 DVDD.n1539 DVSS 0.004621f
C2046 DVDD.n1540 DVSS 0.008245f
C2047 DVDD.n1548 DVSS 0.026423f
C2048 DVDD.n1549 DVSS 0.01188f
C2049 DVDD.t100 DVSS 0.032253f
C2050 DVDD.t144 DVSS 0.032253f
C2051 DVDD.n1550 DVSS 0.064506f
C2052 DVDD.n1551 DVSS 0.011628f
C2053 DVDD.n1552 DVSS 0.011569f
C2054 DVDD.n1564 DVSS 0.02512f
C2055 DVDD.n1565 DVSS 0.052845f
C2056 DVDD.n1566 DVSS 0.052845f
C2057 DVDD.n1567 DVSS 0.052845f
C2058 DVDD.n1568 DVSS 0.052845f
C2059 DVDD.n1569 DVSS 0.052845f
C2060 DVDD.n1570 DVSS 0.052845f
C2061 DVDD.n1571 DVSS 0.052845f
C2062 DVDD.n1572 DVSS 0.052845f
C2063 DVDD.n1573 DVSS 0.052845f
C2064 DVDD.n1574 DVSS 0.052845f
C2065 DVDD.n1575 DVSS 0.052845f
C2066 DVDD.n1576 DVSS 0.052845f
C2067 DVDD.n1577 DVSS 0.052845f
C2068 DVDD.n1578 DVSS 0.052845f
C2069 DVDD.n1579 DVSS 0.052845f
C2070 DVDD.n1580 DVSS 0.052845f
C2071 DVDD.n1581 DVSS 0.052845f
C2072 DVDD.n1582 DVSS 0.032377f
C2073 DVDD.n1583 DVSS 0.032377f
C2074 DVDD.n1584 DVSS 0.046891f
C2075 DVDD.n1585 DVSS 0.052845f
C2076 DVDD.n1586 DVSS 0.063637f
C2077 DVDD.n1587 DVSS 0.052845f
C2078 DVDD.n1588 DVSS 0.052845f
C2079 DVDD.n1589 DVSS 0.052845f
C2080 DVDD.n1590 DVSS 0.052845f
C2081 DVDD.n1591 DVSS 0.052845f
C2082 DVDD.n1592 DVSS 0.052845f
C2083 DVDD.n1593 DVSS 0.002593f
C2084 DVDD.n1594 DVSS 0.002493f
C2085 DVDD.n1595 DVSS 0.001538f
C2086 DVDD.n1596 DVSS 0.00134f
C2087 DVDD.n1597 DVSS 0.025778f
C2088 DVDD.n1598 DVSS 0.025778f
C2089 DVDD.n1599 DVSS 0.023073f
C2090 DVDD.n1600 DVSS 0.003076f
C2091 DVDD.n1601 DVSS 0.001538f
C2092 DVDD.n1602 DVSS 0.003076f
C2093 DVDD.n1603 DVSS 0.003076f
C2094 DVDD.n1604 DVSS 0.003076f
C2095 DVDD.n1605 DVSS 0.003076f
C2096 DVDD.n1606 DVSS 0.002121f
C2097 DVDD.n1607 DVSS 0.003076f
C2098 DVDD.n1608 DVSS 0.052845f
C2099 DVDD.n1609 DVSS 0.052845f
C2100 DVDD.n1610 DVSS 0.052845f
C2101 DVDD.n1611 DVSS 0.052845f
C2102 DVDD.n1612 DVSS 0.052845f
C2103 DVDD.n1613 DVSS 0.052845f
C2104 DVDD.n1614 DVSS 0.052845f
C2105 DVDD.n1615 DVSS 0.052845f
C2106 DVDD.n1616 DVSS 0.052845f
C2107 DVDD.n1617 DVSS 0.052845f
C2108 DVDD.n1618 DVSS 0.052845f
C2109 DVDD.n1619 DVSS 0.052845f
C2110 DVDD.n1620 DVSS 0.052845f
C2111 DVDD.n1621 DVSS 0.052845f
C2112 DVDD.n1622 DVSS 0.052845f
C2113 DVDD.n1623 DVSS 0.052845f
C2114 DVDD.n1624 DVSS 0.052845f
C2115 DVDD.n1625 DVSS 0.052845f
C2116 DVDD.n1626 DVSS 0.052845f
C2117 DVDD.n1627 DVSS 0.052845f
C2118 DVDD.n1628 DVSS 0.052845f
C2119 DVDD.n1629 DVSS 0.052845f
C2120 DVDD.n1630 DVSS 0.052845f
C2121 DVDD.n1631 DVSS 0.052845f
C2122 DVDD.n1632 DVSS 0.052845f
C2123 DVDD.n1633 DVSS 0.030888f
C2124 DVDD.n1634 DVSS 0.048379f
C2125 DVDD.n1635 DVSS 0.052845f
C2126 DVDD.n1636 DVSS 0.052845f
C2127 DVDD.n1637 DVSS 0.052845f
C2128 DVDD.n1638 DVSS 0.052845f
C2129 DVDD.n1639 DVSS 0.052845f
C2130 DVDD.n1640 DVSS 0.052845f
C2131 DVDD.n1641 DVSS 0.052845f
C2132 DVDD.n1642 DVSS 0.052845f
C2133 DVDD.n1643 DVSS 0.052845f
C2134 DVDD.n1644 DVSS 0.052845f
C2135 DVDD.n1645 DVSS 0.052845f
C2136 DVDD.n1646 DVSS 0.052845f
C2137 DVDD.n1647 DVSS 0.052845f
C2138 DVDD.n1648 DVSS 0.052845f
C2139 DVDD.n1649 DVSS 0.047635f
C2140 DVDD.n1650 DVSS 0.005954f
C2141 DVDD.n1651 DVSS 0.243482f
C2142 DVDD.n1652 DVSS 0.075079f
C2143 DVDD.n1653 DVSS 0.047635f
C2144 DVDD.n1654 DVSS 0.047635f
C2145 DVDD.n1655 DVSS 0.052845f
C2146 DVDD.n1656 DVSS 0.052845f
C2147 DVDD.n1657 DVSS 0.052845f
C2148 DVDD.n1658 DVSS 0.052845f
C2149 DVDD.n1659 DVSS 0.052845f
C2150 DVDD.n1660 DVSS 0.052845f
C2151 DVDD.n1661 DVSS 0.052845f
C2152 DVDD.n1662 DVSS 0.052845f
C2153 DVDD.n1663 DVSS 0.052845f
C2154 DVDD.n1664 DVSS 0.052845f
C2155 DVDD.n1665 DVSS 0.052845f
C2156 DVDD.n1666 DVSS 0.052845f
C2157 DVDD.n1667 DVSS 0.052845f
C2158 DVDD.n1668 DVSS 0.048379f
C2159 DVDD.n1669 DVSS 0.048379f
C2160 DVDD.n1670 DVSS 0.063637f
C2161 DVDD.n1671 DVSS 0.030888f
C2162 DVDD.n1672 DVSS 0.052845f
C2163 DVDD.n1673 DVSS 0.052845f
C2164 DVDD.n1674 DVSS 0.043355f
C2165 DVDD.n1675 DVSS 0.052845f
C2166 DVDD.n1676 DVSS 0.052845f
C2167 DVDD.n1677 DVSS 0.052845f
C2168 DVDD.n1678 DVSS 0.052845f
C2169 DVDD.n1679 DVSS 0.052845f
C2170 DVDD.n1680 DVSS 0.052845f
C2171 DVDD.n1681 DVSS 0.052845f
C2172 DVDD.n1682 DVSS 0.052845f
C2173 DVDD.n1683 DVSS 0.052845f
C2174 DVDD.n1684 DVSS 0.052845f
C2175 DVDD.n1685 DVSS 0.052845f
C2176 DVDD.n1686 DVSS 0.052845f
C2177 DVDD.n1687 DVSS 0.052845f
C2178 DVDD.n1688 DVSS 0.052845f
C2179 DVDD.n1689 DVSS 0.052845f
C2180 DVDD.n1690 DVSS 0.052845f
C2181 DVDD.n1691 DVSS 0.052845f
C2182 DVDD.n1692 DVSS 0.052845f
C2183 DVDD.n1693 DVSS 0.052845f
C2184 DVDD.n1694 DVSS 0.052845f
C2185 DVDD.n1695 DVSS 0.052845f
C2186 DVDD.n1696 DVSS 0.052845f
C2187 DVDD.n1697 DVSS 0.031074f
C2188 DVDD.n1698 DVSS 0.001538f
C2189 DVDD.n1699 DVSS 0.003076f
C2190 DVDD.n1700 DVSS 0.001538f
C2191 DVDD.n1701 DVSS 0.002171f
C2192 DVDD.n1702 DVSS 0.003076f
C2193 DVDD.n1703 DVSS 0.003076f
C2194 DVDD.n1704 DVSS 0.003076f
C2195 DVDD.n1705 DVSS 0.003076f
C2196 DVDD.n1706 DVSS 0.001538f
C2197 DVDD.n1707 DVSS 0.001538f
C2198 DVDD.n1709 DVSS 0.026423f
C2199 DVDD.n1710 DVSS 0.001538f
C2200 DVDD.n1711 DVSS 0.002022f
C2201 DVDD.n1712 DVSS 0.002593f
C2202 DVDD.n1713 DVSS 0.008261f
C2203 DVDD.n1714 DVSS 0.004122f
C2204 DVDD.n1715 DVSS 0.002022f
C2205 DVDD.n1717 DVSS 0.031819f
C2206 DVDD.n1718 DVSS 0.002493f
C2207 DVDD.n1719 DVSS 0.001538f
C2208 DVDD.n1720 DVSS 0.00134f
C2209 DVDD.n1721 DVSS 0.025778f
C2210 DVDD.n1722 DVSS 0.025778f
C2211 DVDD.n1723 DVSS 0.023073f
C2212 DVDD.n1724 DVSS 0.003076f
C2213 DVDD.n1725 DVSS 0.001538f
C2214 DVDD.n1726 DVSS 0.003076f
C2215 DVDD.n1727 DVSS 0.003076f
C2216 DVDD.n1728 DVSS 0.003076f
C2217 DVDD.n1729 DVSS 0.003076f
C2218 DVDD.t153 DVSS 0.032253f
C2219 DVDD.t99 DVSS 0.032253f
C2220 DVDD.n1730 DVSS 0.064506f
C2221 DVDD.n1731 DVSS 0.002121f
C2222 DVDD.n1732 DVSS 0.002493f
C2223 DVDD.n1733 DVSS 0.008261f
C2224 DVDD.n1734 DVSS 0.001538f
C2225 DVDD.n1735 DVSS 0.027944f
C2226 DVDD.n1736 DVSS 0.011628f
C2227 DVDD.n1737 DVSS 0.004122f
C2228 DVDD.n1738 DVSS 0.01188f
C2229 DVDD.n1739 DVSS 0.008262f
C2230 DVDD.n1740 DVSS 0.027687f
C2231 DVDD.n1741 DVSS 0.001538f
C2232 DVDD.n1742 DVSS 0.002121f
C2233 DVDD.n1743 DVSS 0.001538f
C2234 DVDD.n1744 DVSS 0.052845f
C2235 DVDD.n1745 DVSS 0.052845f
C2236 DVDD.n1746 DVSS 0.052845f
C2237 DVDD.n1747 DVSS 0.052845f
C2238 DVDD.n1748 DVSS 0.052845f
C2239 DVDD.n1749 DVSS 0.052845f
C2240 DVDD.n1750 DVSS 0.052845f
C2241 DVDD.n1751 DVSS 0.033866f
C2242 DVDD.n1752 DVSS 0.033866f
C2243 DVDD.n1753 DVSS 0.052845f
C2244 DVDD.n1754 DVSS 0.052845f
C2245 DVDD.n1755 DVSS 0.052845f
C2246 DVDD.n1756 DVSS 0.052845f
C2247 DVDD.n1757 DVSS 0.052845f
C2248 DVDD.n1758 DVSS 0.052845f
C2249 DVDD.n1759 DVSS 0.052845f
C2250 DVDD.n1760 DVSS 0.052845f
C2251 DVDD.n1761 DVSS 0.052845f
C2252 DVDD.n1762 DVSS 0.052845f
C2253 DVDD.n1763 DVSS 0.052845f
C2254 DVDD.n1764 DVSS 0.052845f
C2255 DVDD.n1765 DVSS 0.052845f
C2256 DVDD.n1766 DVSS 0.052845f
C2257 DVDD.n1767 DVSS 0.052845f
C2258 DVDD.n1768 DVSS 0.052845f
C2259 DVDD.n1769 DVSS 0.052845f
C2260 DVDD.n1770 DVSS 0.052845f
C2261 DVDD.n1771 DVSS 0.052845f
C2262 DVDD.n1772 DVSS 0.052845f
C2263 DVDD.n1773 DVSS 0.908729f
C2264 DVDD.n1774 DVSS 0.20542f
C2265 DVDD.n1775 DVSS 0.766395f
C2266 DVDD.n1776 DVSS 0.242697f
C2267 DVDD.n1777 DVSS 0.9643f
C2268 DVDD.n1778 DVSS 0.052845f
C2269 DVDD.n1779 DVSS 0.043914f
C2270 DVDD.n1780 DVSS 0.72918f
C2271 DVDD.n1781 DVSS 0.9643f
C2272 DVDD.n1782 DVSS 0.052845f
C2273 DVDD.n1783 DVSS 0.043914f
C2274 DVDD.n1784 DVSS 0.242697f
C2275 DVDD.n1785 DVSS 0.205482f
C2276 DVDD.n1786 DVSS 0.052845f
C2277 DVDD.n1787 DVSS 0.052845f
C2278 DVDD.n1788 DVSS 0.003076f
C2279 DVDD.n1789 DVSS 0.001538f
C2280 DVDD.n1790 DVSS 0.002171f
C2281 DVDD.n1791 DVSS 0.003076f
C2282 DVDD.n1792 DVSS 0.003076f
C2283 DVDD.n1793 DVSS 0.003076f
C2284 DVDD.n1794 DVSS 0.003076f
C2285 DVDD.n1795 DVSS 0.001538f
C2286 DVDD.n1796 DVSS 0.001538f
C2287 DVDD.n1797 DVSS 0.001538f
C2288 DVDD.n1798 DVSS 0.026423f
C2289 DVDD.n1799 DVSS 0.052845f
C2290 DVDD.n1800 DVSS 0.052845f
C2291 DVDD.n1801 DVSS 0.052845f
C2292 DVDD.n1802 DVSS 0.052845f
C2293 DVDD.n1803 DVSS 0.052845f
C2294 DVDD.n1804 DVSS 0.052845f
C2295 DVDD.n1805 DVSS 0.052845f
C2296 DVDD.n1806 DVSS 0.052845f
C2297 DVDD.n1807 DVSS 0.052845f
C2298 DVDD.n1808 DVSS 0.052845f
C2299 DVDD.n1809 DVSS 0.052845f
C2300 DVDD.n1810 DVSS 0.052845f
C2301 DVDD.n1811 DVSS 0.052845f
C2302 DVDD.n1812 DVSS 0.052845f
C2303 DVDD.n1813 DVSS 0.052845f
C2304 DVDD.n1814 DVSS 0.052845f
C2305 DVDD.n1815 DVSS 0.052845f
C2306 DVDD.n1816 DVSS 0.052845f
C2307 DVDD.n1817 DVSS 0.052845f
C2308 DVDD.n1818 DVSS 0.052845f
C2309 DVDD.n1819 DVSS 0.052845f
C2310 DVDD.n1820 DVSS 0.052845f
C2311 DVDD.n1821 DVSS 0.052845f
C2312 DVDD.n1822 DVSS 0.052845f
C2313 DVDD.n1823 DVSS 0.052845f
C2314 DVDD.n1824 DVSS 0.052845f
C2315 DVDD.n1825 DVSS 0.052845f
C2316 DVDD.n1826 DVSS 0.052845f
C2317 DVDD.n1827 DVSS 0.052845f
C2318 DVDD.n1828 DVSS 0.052845f
C2319 DVDD.n1829 DVSS 0.052845f
C2320 DVDD.n1830 DVSS 0.052845f
C2321 DVDD.n1831 DVSS 0.052845f
C2322 DVDD.n1832 DVSS 0.052845f
C2323 DVDD.n1833 DVSS 0.052845f
C2324 DVDD.n1834 DVSS 0.052845f
C2325 DVDD.n1835 DVSS 0.052845f
C2326 DVDD.n1836 DVSS 0.052845f
C2327 DVDD.n1837 DVSS 0.052845f
C2328 DVDD.n1838 DVSS 0.052845f
C2329 DVDD.n1839 DVSS 0.052845f
C2330 DVDD.n1840 DVSS 0.052845f
C2331 DVDD.n1841 DVSS 0.052845f
C2332 DVDD.n1842 DVSS 0.052845f
C2333 DVDD.n1843 DVSS 0.042611f
C2334 DVDD.n1844 DVSS 0.052845f
C2335 DVDD.n1845 DVSS 0.052845f
C2336 DVDD.n1846 DVSS 0.043914f
C2337 DVDD.n1847 DVSS 0.043914f
C2338 DVDD.n1848 DVSS 0.903314f
C2339 DVDD.n1849 DVSS 0.940529f
C2340 DVDD.n1850 DVSS 0.052845f
C2341 DVDD.n1851 DVSS 0.043914f
C2342 DVDD.n1852 DVSS 0.043914f
C2343 DVDD.n1853 DVSS 0.940529f
C2344 DVDD.n1854 DVSS 0.9643f
C2345 DVDD.n1855 DVSS 0.766395f
C2346 DVDD.n1856 DVSS 0.964426f
C2347 DVDD.n1857 DVSS 0.723701f
C2348 DVDD.n1858 DVSS 0.031074f
C2349 DVDD.n1859 DVSS 0.043914f
C2350 DVDD.n1860 DVSS 0.043914f
C2351 DVDD.n1861 DVSS 0.052845f
C2352 DVDD.n1862 DVSS 0.052845f
C2353 DVDD.n1863 DVSS 0.052845f
C2354 DVDD.n1864 DVSS 0.052845f
C2355 DVDD.n1865 DVSS 0.052845f
C2356 DVDD.n1866 DVSS 0.052845f
C2357 DVDD.n1867 DVSS 0.052845f
C2358 DVDD.n1868 DVSS 0.052845f
C2359 DVDD.n1869 DVSS 0.052845f
C2360 DVDD.n1870 DVSS 0.052845f
C2361 DVDD.n1871 DVSS 0.052845f
C2362 DVDD.n1872 DVSS 0.052845f
C2363 DVDD.n1873 DVSS 0.052845f
C2364 DVDD.n1874 DVSS 0.052845f
C2365 DVDD.n1875 DVSS 0.052845f
C2366 DVDD.n1876 DVSS 0.052845f
C2367 DVDD.n1877 DVSS 0.052845f
C2368 DVDD.n1878 DVSS 0.052845f
C2369 DVDD.n1879 DVSS 0.052845f
C2370 DVDD.n1880 DVSS 0.052845f
C2371 DVDD.n1881 DVSS 0.052845f
C2372 DVDD.n1882 DVSS 0.052845f
C2373 DVDD.n1883 DVSS 0.052845f
C2374 DVDD.n1884 DVSS 0.052845f
C2375 DVDD.n1885 DVSS 0.052845f
C2376 DVDD.n1886 DVSS 0.052845f
C2377 DVDD.n1887 DVSS 0.052845f
C2378 DVDD.n1888 DVSS 0.052845f
C2379 DVDD.n1889 DVSS 0.052845f
C2380 DVDD.n1890 DVSS 0.052845f
C2381 DVDD.n1891 DVSS 0.052845f
C2382 DVDD.n1892 DVSS 0.052845f
C2383 DVDD.n1893 DVSS 0.052845f
C2384 DVDD.n1894 DVSS 0.052845f
C2385 DVDD.n1895 DVSS 0.052845f
C2386 DVDD.n1896 DVSS 0.052845f
C2387 DVDD.n1897 DVSS 0.052845f
C2388 DVDD.n1898 DVSS 0.052845f
C2389 DVDD.n1899 DVSS 0.052845f
C2390 DVDD.n1900 DVSS 0.052845f
C2391 DVDD.n1901 DVSS 0.052845f
C2392 DVDD.n1902 DVSS 0.052845f
C2393 DVDD.n1903 DVSS 0.052845f
C2394 DVDD.n1904 DVSS 0.033866f
C2395 DVDD.n1905 DVSS 0.033866f
C2396 DVDD.n1906 DVSS 0.063637f
C2397 DVDD.n1907 DVSS 0.052845f
C2398 DVDD.n1908 DVSS 0.052845f
C2399 DVDD.n1909 DVSS 0.052845f
C2400 DVDD.n1910 DVSS 0.052845f
C2401 DVDD.n1911 DVSS 0.052845f
C2402 DVDD.n1912 DVSS 0.052845f
C2403 DVDD.n1913 DVSS 0.052845f
C2404 DVDD.n1914 DVSS 0.052845f
C2405 DVDD.n1915 DVSS 0.052845f
C2406 DVDD.n1916 DVSS 0.052845f
C2407 DVDD.n1917 DVSS 0.052845f
C2408 DVDD.n1918 DVSS 0.052845f
C2409 DVDD.n1919 DVSS 0.052845f
C2410 DVDD.n1920 DVSS 0.052845f
C2411 DVDD.n1921 DVSS 0.052845f
C2412 DVDD.n1922 DVSS 0.023073f
C2413 DVDD.n1923 DVSS 0.052845f
C2414 DVDD.n1924 DVSS 0.052845f
C2415 DVDD.n1925 DVSS 0.031819f
C2416 DVDD.n1926 DVSS 0.052845f
C2417 DVDD.n1927 DVSS 0.052845f
C2418 DVDD.n1928 DVSS 0.052845f
C2419 DVDD.n1929 DVSS 0.052845f
C2420 DVDD.n1930 DVSS 0.052845f
C2421 DVDD.n1931 DVSS 0.052845f
C2422 DVDD.n1932 DVSS 0.052845f
C2423 DVDD.n1933 DVSS 0.052845f
C2424 DVDD.n1934 DVSS 0.052845f
C2425 DVDD.n1935 DVSS 0.052845f
C2426 DVDD.n1936 DVSS 0.052845f
C2427 DVDD.n1937 DVSS 0.052845f
C2428 DVDD.n1938 DVSS 0.052845f
C2429 DVDD.n1939 DVSS 0.045402f
C2430 DVDD.n1940 DVSS 0.045402f
C2431 DVDD.n1941 DVSS 0.045402f
C2432 DVDD.n1942 DVSS 0.063637f
C2433 DVDD.n1943 DVSS 0.100852f
C2434 DVDD.n1944 DVSS 0.100852f
C2435 DVDD.n1945 DVSS 0.063637f
C2436 DVDD.n1946 DVSS 0.045402f
C2437 DVDD.n1947 DVSS 0.052845f
C2438 DVDD.n1948 DVSS 0.052845f
C2439 DVDD.n1949 DVSS 0.052845f
C2440 DVDD.n1950 DVSS 0.052845f
C2441 DVDD.n1951 DVSS 0.052845f
C2442 DVDD.n1952 DVSS 0.052845f
C2443 DVDD.n1953 DVSS 0.052845f
C2444 DVDD.n1954 DVSS 0.052845f
C2445 DVDD.n1955 DVSS 0.052845f
C2446 DVDD.n1956 DVSS 0.052845f
C2447 DVDD.n1957 DVSS 0.052845f
C2448 DVDD.n1958 DVSS 0.052845f
C2449 DVDD.n1959 DVSS 0.052845f
C2450 DVDD.n1960 DVSS 0.052845f
C2451 DVDD.n1961 DVSS 0.052845f
C2452 DVDD.n1962 DVSS 0.052845f
C2453 DVDD.n1963 DVSS 0.052845f
C2454 DVDD.n1964 DVSS 0.052845f
C2455 DVDD.n1965 DVSS 0.052845f
C2456 DVDD.n1966 DVSS 0.052845f
C2457 DVDD.n1967 DVSS 0.052845f
C2458 DVDD.n1968 DVSS 0.052845f
C2459 DVDD.n1969 DVSS 0.052845f
C2460 DVDD.n1970 DVSS 0.052845f
C2461 DVDD.n1971 DVSS 0.052845f
C2462 DVDD.n1972 DVSS 0.052845f
C2463 DVDD.n1973 DVSS 0.052845f
C2464 DVDD.n1974 DVSS 0.052845f
C2465 DVDD.n1975 DVSS 0.052845f
C2466 DVDD.n1976 DVSS 0.063637f
C2467 DVDD.n1977 DVSS 0.032377f
C2468 DVDD.n1978 DVSS 0.052845f
C2469 DVDD.n1979 DVSS 0.052845f
C2470 DVDD.n1980 DVSS 0.032377f
C2471 DVDD.n1981 DVSS 0.052845f
C2472 DVDD.n1982 DVSS 0.052845f
C2473 DVDD.n1983 DVSS 0.052845f
C2474 DVDD.n1984 DVSS 0.052845f
C2475 DVDD.n1985 DVSS 0.052845f
C2476 DVDD.n1986 DVSS 0.052845f
C2477 DVDD.n1987 DVSS 0.052845f
C2478 DVDD.n1988 DVSS 0.052845f
C2479 DVDD.n1989 DVSS 0.052845f
C2480 DVDD.n1990 DVSS 0.052845f
C2481 DVDD.n1991 DVSS 0.052845f
C2482 DVDD.n1992 DVSS 0.052845f
C2483 DVDD.n1993 DVSS 0.052845f
C2484 DVDD.n1994 DVSS 0.031074f
C2485 DVDD.n1995 DVSS 0.052845f
C2486 DVDD.n1996 DVSS 0.023073f
C2487 DVDD.n1997 DVSS 0.052845f
C2488 DVDD.n1998 DVSS 0.052845f
C2489 DVDD.n1999 DVSS 0.052845f
C2490 DVDD.n2000 DVSS 0.052845f
C2491 DVDD.n2001 DVSS 0.052845f
C2492 DVDD.n2002 DVSS 0.052845f
C2493 DVDD.n2003 DVSS 0.052845f
C2494 DVDD.n2004 DVSS 0.052845f
C2495 DVDD.n2005 DVSS 0.052845f
C2496 DVDD.n2006 DVSS 0.052845f
C2497 DVDD.n2007 DVSS 0.052845f
C2498 DVDD.n2008 DVSS 0.052845f
C2499 DVDD.n2009 DVSS 0.052845f
C2500 DVDD.n2010 DVSS 0.052845f
C2501 DVDD.n2011 DVSS 0.052845f
C2502 DVDD.n2012 DVSS 0.052845f
C2503 DVDD.n2013 DVSS 0.052845f
C2504 DVDD.n2014 DVSS 0.045402f
C2505 DVDD.n2015 DVSS 0.045402f
C2506 DVDD.n2016 DVSS 0.063637f
C2507 DVDD.n2017 DVSS 0.033866f
C2508 DVDD.n2018 DVSS 0.033866f
C2509 DVDD.n2019 DVSS 0.052845f
C2510 DVDD.n2020 DVSS 0.052845f
C2511 DVDD.n2021 DVSS 0.052845f
C2512 DVDD.n2022 DVSS 0.052845f
C2513 DVDD.n2023 DVSS 0.052845f
C2514 DVDD.n2024 DVSS 0.050798f
C2515 DVDD.n2025 DVSS 0.001538f
C2516 DVDD.n2026 DVSS 0.003076f
C2517 DVDD.n2027 DVSS 0.001538f
C2518 DVDD.n2028 DVSS 0.002171f
C2519 DVDD.n2029 DVSS 0.003076f
C2520 DVDD.n2030 DVSS 0.003076f
C2521 DVDD.n2031 DVSS 0.003076f
C2522 DVDD.n2032 DVSS 0.003076f
C2523 DVDD.n2033 DVSS 0.001538f
C2524 DVDD.n2034 DVSS 0.026423f
C2525 DVDD.n2035 DVSS 0.001538f
C2526 DVDD.n2036 DVSS 0.003076f
C2527 DVDD.n2037 DVSS 0.026423f
C2528 DVDD.n2038 DVSS 0.002593f
C2529 DVDD.n2039 DVSS 0.001538f
C2530 DVDD.n2040 DVSS 0.008262f
C2531 DVDD.n2041 DVSS 0.027687f
C2532 DVDD.n2042 DVSS 0.01188f
C2533 DVDD.t150 DVSS 0.032253f
C2534 DVDD.t106 DVSS 0.032253f
C2535 DVDD.n2043 DVSS 0.064506f
C2536 DVDD.n2044 DVSS 0.011628f
C2537 DVDD.n2045 DVSS 0.027944f
C2538 DVDD.n2046 DVSS 0.001538f
C2539 DVDD.n2047 DVSS 0.002022f
C2540 DVDD.n2048 DVSS 0.026423f
C2541 DVDD.n2049 DVSS 0.051543f
C2542 DVDD.n2050 DVSS 0.052845f
C2543 DVDD.n2051 DVSS 0.052845f
C2544 DVDD.n2052 DVSS 0.052845f
C2545 DVDD.n2053 DVSS 0.052845f
C2546 DVDD.n2054 DVSS 0.052845f
C2547 DVDD.n2055 DVSS 0.046891f
C2548 DVDD.n2056 DVSS 0.046891f
C2549 DVDD.n2057 DVSS 0.063637f
C2550 DVDD.n2058 DVSS 0.046891f
C2551 DVDD.n2059 DVSS 0.052845f
C2552 DVDD.n2060 DVSS 0.052845f
C2553 DVDD.n2061 DVSS 0.052845f
C2554 DVDD.n2062 DVSS 0.052845f
C2555 DVDD.n2063 DVSS 0.052845f
C2556 DVDD.n2064 DVSS 0.052845f
C2557 DVDD.n2065 DVSS 0.052845f
C2558 DVDD.n2066 DVSS 0.052845f
C2559 DVDD.n2067 DVSS 0.052845f
C2560 DVDD.n2068 DVSS 0.001538f
C2561 DVDD.n2069 DVSS 0.001538f
C2562 DVDD.n2070 DVSS 0.001538f
C2563 DVDD.n2071 DVSS 0.001538f
C2564 DVDD.n2072 DVSS 0.001538f
C2565 DVDD.n2073 DVSS 0.001538f
C2566 DVDD.n2074 DVSS 0.001538f
C2567 DVDD.n2075 DVSS 0.001538f
C2568 DVDD.n2076 DVSS 0.001538f
C2569 DVDD.n2077 DVSS 0.001538f
C2570 DVDD.n2078 DVSS 0.026423f
C2571 DVDD.n2079 DVSS 0.052845f
C2572 DVDD.n2080 DVSS 0.052845f
C2573 DVDD.n2081 DVSS 0.052845f
C2574 DVDD.n2082 DVSS 0.052845f
C2575 DVDD.n2083 DVSS 0.052845f
C2576 DVDD.n2084 DVSS 0.052845f
C2577 DVDD.n2085 DVSS 0.052845f
C2578 DVDD.n2086 DVSS 0.052845f
C2579 DVDD.n2087 DVSS 0.052845f
C2580 DVDD.n2088 DVSS 0.052845f
C2581 DVDD.n2089 DVSS 0.052845f
C2582 DVDD.n2090 DVSS 0.052845f
C2583 DVDD.n2091 DVSS 0.052845f
C2584 DVDD.n2092 DVSS 0.052845f
C2585 DVDD.n2093 DVSS 0.052845f
C2586 DVDD.n2094 DVSS 0.052845f
C2587 DVDD.n2095 DVSS 0.052845f
C2588 DVDD.n2096 DVSS 0.052845f
C2589 DVDD.n2097 DVSS 0.043355f
C2590 DVDD.n2098 DVSS 0.052845f
C2591 DVDD.n2099 DVSS 0.052845f
C2592 DVDD.n2100 DVSS 0.052845f
C2593 DVDD.n2101 DVSS 0.052845f
C2594 DVDD.n2102 DVSS 0.052845f
C2595 DVDD.n2103 DVSS 0.052845f
C2596 DVDD.n2104 DVSS 0.052845f
C2597 DVDD.n2105 DVSS 0.052845f
C2598 DVDD.n2106 DVSS 0.052845f
C2599 DVDD.n2107 DVSS 0.052845f
C2600 DVDD.n2108 DVSS 0.052845f
C2601 DVDD.n2109 DVSS 0.052845f
C2602 DVDD.n2110 DVSS 0.052845f
C2603 DVDD.n2111 DVSS 0.052845f
C2604 DVDD.n2112 DVSS 0.052845f
C2605 DVDD.n2113 DVSS 0.052845f
C2606 DVDD.n2114 DVSS 0.052845f
C2607 DVDD.n2115 DVSS 0.052845f
C2608 DVDD.n2116 DVSS 0.052845f
C2609 DVDD.n2117 DVSS 0.052845f
C2610 DVDD.n2118 DVSS 0.052845f
C2611 DVDD.n2119 DVSS 0.052845f
C2612 DVDD.n2120 DVSS 0.052845f
C2613 DVDD.n2121 DVSS 0.052845f
C2614 DVDD.n2122 DVSS 0.031074f
C2615 DVDD.n2123 DVSS 0.052845f
C2616 DVDD.n2124 DVSS 0.052845f
C2617 DVDD.n2125 DVSS 0.052845f
C2618 DVDD.n2126 DVSS 0.052845f
C2619 DVDD.n2127 DVSS 0.052845f
C2620 DVDD.n2128 DVSS 0.052845f
C2621 DVDD.n2129 DVSS 0.052845f
C2622 DVDD.n2130 DVSS 0.046891f
C2623 DVDD.n2131 DVSS 0.046891f
C2624 DVDD.n2132 DVSS 0.100852f
C2625 DVDD.n2133 DVSS 0.032377f
C2626 DVDD.n2134 DVSS 0.032377f
C2627 DVDD.n2135 DVSS 0.052845f
C2628 DVDD.n2136 DVSS 0.052845f
C2629 DVDD.n2137 DVSS 0.052845f
C2630 DVDD.n2138 DVSS 0.052845f
C2631 DVDD.n2139 DVSS 0.052845f
C2632 DVDD.n2140 DVSS 0.052845f
C2633 DVDD.n2141 DVSS 0.052845f
C2634 DVDD.n2142 DVSS 0.052845f
C2635 DVDD.n2143 DVSS 0.052845f
C2636 DVDD.n2144 DVSS 0.052845f
C2637 DVDD.n2145 DVSS 0.052845f
C2638 DVDD.n2146 DVSS 0.052845f
C2639 DVDD.n2147 DVSS 0.052845f
C2640 DVDD.n2148 DVSS 0.031074f
C2641 DVDD.n2149 DVSS 0.052845f
C2642 DVDD.n2150 DVSS 0.052845f
C2643 DVDD.n2151 DVSS 0.023073f
C2644 DVDD.n2152 DVSS 0.024376f
C2645 DVDD.n2153 DVSS 0.004355f
C2646 DVDD.n2154 DVSS 0.026423f
C2647 DVDD.n2155 DVSS 0.031819f
C2648 DVDD.n2156 DVSS 0.052845f
C2649 DVDD.n2157 DVSS 0.052845f
C2650 DVDD.n2158 DVSS 0.052845f
C2651 DVDD.n2159 DVSS 0.052845f
C2652 DVDD.n2160 DVSS 0.052845f
C2653 DVDD.n2161 DVSS 0.052845f
C2654 DVDD.n2162 DVSS 0.052845f
C2655 DVDD.n2163 DVSS 0.052845f
C2656 DVDD.n2164 DVSS 0.052845f
C2657 DVDD.n2165 DVSS 0.052845f
C2658 DVDD.n2166 DVSS 0.052845f
C2659 DVDD.n2167 DVSS 0.052845f
C2660 DVDD.n2168 DVSS 0.052845f
C2661 DVDD.n2169 DVSS 0.052845f
C2662 DVDD.n2170 DVSS 0.045402f
C2663 DVDD.n2171 DVSS 0.045402f
C2664 DVDD.n2172 DVSS 0.100852f
C2665 DVDD.n2173 DVSS 0.033866f
C2666 DVDD.n2174 DVSS 0.033866f
C2667 DVDD.n2175 DVSS 0.052845f
C2668 DVDD.n2176 DVSS 0.052845f
C2669 DVDD.n2177 DVSS 0.052845f
C2670 DVDD.n2178 DVSS 0.052845f
C2671 DVDD.n2179 DVSS 0.050798f
C2672 DVDD.n2180 DVSS 0.052845f
C2673 DVDD.n2181 DVSS 0.052845f
C2674 DVDD.n2182 DVSS 0.052845f
C2675 DVDD.n2183 DVSS 0.052845f
C2676 DVDD.n2184 DVSS 0.052845f
C2677 DVDD.n2185 DVSS 0.052845f
C2678 DVDD.n2186 DVSS 0.052845f
C2679 DVDD.n2187 DVSS 0.052845f
C2680 DVDD.n2188 DVSS 0.052845f
C2681 DVDD.n2189 DVSS 0.052845f
C2682 DVDD.n2190 DVSS 0.052845f
C2683 DVDD.n2191 DVSS 0.052845f
C2684 DVDD.n2192 DVSS 0.052845f
C2685 DVDD.n2193 DVSS 0.052845f
C2686 DVDD.n2194 DVSS 0.052845f
C2687 DVDD.n2195 DVSS 0.052845f
C2688 DVDD.n2196 DVSS 0.052845f
C2689 DVDD.n2197 DVSS 0.052845f
C2690 DVDD.n2198 DVSS 0.052845f
C2691 DVDD.n2199 DVSS 0.052845f
C2692 DVDD.n2200 DVSS 0.052845f
C2693 DVDD.n2201 DVSS 0.052845f
C2694 DVDD.n2202 DVSS 0.052845f
C2695 DVDD.n2203 DVSS 0.052845f
C2696 DVDD.n2204 DVSS 0.052845f
C2697 DVDD.n2205 DVSS 0.042611f
C2698 DVDD.n2206 DVSS 0.001538f
C2699 DVDD.n2207 DVSS 0.001538f
C2700 DVDD.n2208 DVSS 0.001538f
C2701 DVDD.n2209 DVSS 0.001538f
C2702 DVDD.n2210 DVSS 0.001538f
C2703 DVDD.n2211 DVSS 0.001538f
C2704 DVDD.n2212 DVSS 0.001538f
C2705 DVDD.n2213 DVSS 0.001538f
C2706 DVDD.n2214 DVSS 0.001538f
C2707 DVDD.n2215 DVSS 0.001538f
C2708 DVDD.n2216 DVSS 0.026423f
C2709 DVDD.n2217 DVSS 0.001538f
C2710 DVDD.n2218 DVSS 0.011041f
C2711 DVDD.n2219 DVSS 0.001625f
C2712 DVDD.n2220 DVSS 0.026423f
C2713 DVDD.n2221 DVSS 0.00289f
C2714 DVDD.n2222 DVSS 0.008262f
C2715 DVDD.n2223 DVSS 0.027687f
C2716 DVDD.n2224 DVSS 0.01188f
C2717 DVDD.t130 DVSS 0.032253f
C2718 DVDD.t147 DVSS 0.032253f
C2719 DVDD.n2225 DVSS 0.064506f
C2720 DVDD.n2226 DVSS 0.011628f
C2721 DVDD.n2227 DVSS 0.027944f
C2722 DVDD.n2228 DVSS 0.008261f
C2723 DVDD.n2229 DVSS 0.00289f
C2724 DVDD.n2230 DVSS 0.001538f
C2725 DVDD.n2231 DVSS 0.005768f
C2726 DVDD.n2232 DVSS 0.01104f
C2727 DVDD.n2233 DVSS 0.001625f
C2728 DVDD.n2234 DVSS 0.003076f
C2729 DVDD.n2235 DVSS 0.001538f
C2730 DVDD.n2236 DVSS 0.026423f
C2731 DVDD.n2237 DVSS 0.023073f
C2732 DVDD.n2238 DVSS 0.052845f
C2733 DVDD.n2239 DVSS 0.030888f
C2734 DVDD.n2240 DVSS 0.030888f
C2735 DVDD.n2241 DVSS 0.100852f
C2736 DVDD.n2242 DVSS 0.048379f
C2737 DVDD.n2243 DVSS 0.052845f
C2738 DVDD.n2244 DVSS 0.052845f
C2739 DVDD.n2245 DVSS 0.052845f
C2740 DVDD.n2246 DVSS 0.052845f
C2741 DVDD.n2247 DVSS 0.052845f
C2742 DVDD.n2248 DVSS 0.052845f
C2743 DVDD.n2249 DVSS 0.052845f
C2744 DVDD.n2250 DVSS 0.052845f
C2745 DVDD.n2251 DVSS 0.052845f
C2746 DVDD.n2252 DVSS 0.052845f
C2747 DVDD.n2253 DVSS 0.052845f
C2748 DVDD.n2254 DVSS 0.052845f
C2749 DVDD.n2255 DVSS 0.052845f
C2750 DVDD.n2256 DVSS 0.052845f
C2751 DVDD.n2257 DVSS 0.027167f
C2752 DVDD.n2258 DVSS 0.075079f
C2753 DVDD.n2259 DVSS 0.243482f
C2754 DVDD.n2260 DVSS 0.047635f
C2755 DVDD.n2261 DVSS 0.047635f
C2756 DVDD.n2262 DVSS 0.052845f
C2757 DVDD.n2263 DVSS 0.052845f
C2758 DVDD.n2264 DVSS 0.052845f
C2759 DVDD.n2265 DVSS 0.052845f
C2760 DVDD.n2266 DVSS 0.052845f
C2761 DVDD.n2267 DVSS 0.052845f
C2762 DVDD.n2268 DVSS 0.052845f
C2763 DVDD.n2269 DVSS 0.052845f
C2764 DVDD.n2270 DVSS 0.052845f
C2765 DVDD.n2271 DVSS 0.052845f
C2766 DVDD.n2272 DVSS 0.052845f
C2767 DVDD.n2273 DVSS 0.052845f
C2768 DVDD.n2274 DVSS 0.052845f
C2769 DVDD.n2275 DVSS 0.048379f
C2770 DVDD.n2276 DVSS 0.048379f
C2771 DVDD.n2277 DVSS 0.100852f
C2772 DVDD.n2278 DVSS 0.100852f
C2773 DVDD.n2279 DVSS 0.063637f
C2774 DVDD.n2280 DVSS 0.052845f
C2775 DVDD.n2281 DVSS 0.052845f
C2776 DVDD.n2282 DVSS 0.052845f
C2777 DVDD.n2283 DVSS 0.052845f
C2778 DVDD.n2284 DVSS 0.052845f
C2779 DVDD.n2285 DVSS 0.052845f
C2780 DVDD.n2286 DVSS 0.052845f
C2781 DVDD.n2287 DVSS 0.052845f
C2782 DVDD.n2288 DVSS 0.052845f
C2783 DVDD.n2289 DVSS 0.052845f
C2784 DVDD.n2290 DVSS 0.052845f
C2785 DVDD.n2291 DVSS 0.052845f
C2786 DVDD.n2292 DVSS 0.052845f
C2787 DVDD.n2293 DVSS 0.047635f
C2788 DVDD.n2294 DVSS 0.005954f
C2789 DVDD.n2295 DVSS 0.243482f
C2790 DVDD.n2296 DVSS 0.075079f
C2791 DVDD.n2297 DVSS 0.047635f
C2792 DVDD.n2298 DVSS 0.047635f
C2793 DVDD.n2299 DVSS 0.052845f
C2794 DVDD.n2300 DVSS 0.052845f
C2795 DVDD.n2301 DVSS 0.052845f
C2796 DVDD.n2302 DVSS 0.052845f
C2797 DVDD.n2303 DVSS 0.052845f
C2798 DVDD.n2304 DVSS 0.052845f
C2799 DVDD.n2305 DVSS 0.052845f
C2800 DVDD.n2306 DVSS 0.052845f
C2801 DVDD.n2307 DVSS 0.052845f
C2802 DVDD.n2308 DVSS 0.052845f
C2803 DVDD.n2309 DVSS 0.052845f
C2804 DVDD.n2310 DVSS 0.052845f
C2805 DVDD.n2311 DVSS 0.052845f
C2806 DVDD.n2312 DVSS 0.048379f
C2807 DVDD.n2313 DVSS 0.048379f
C2808 DVDD.n2314 DVSS 0.063637f
C2809 DVDD.n2315 DVSS 0.030888f
C2810 DVDD.n2316 DVSS 0.052845f
C2811 DVDD.n2317 DVSS 0.052845f
C2812 DVDD.n2318 DVSS 0.043355f
C2813 DVDD.n2319 DVSS 0.052845f
C2814 DVDD.n2320 DVSS 0.052845f
C2815 DVDD.n2321 DVSS 0.052845f
C2816 DVDD.n2322 DVSS 0.052845f
C2817 DVDD.n2323 DVSS 0.052845f
C2818 DVDD.n2324 DVSS 0.052845f
C2819 DVDD.n2325 DVSS 0.052845f
C2820 DVDD.n2326 DVSS 0.052845f
C2821 DVDD.n2327 DVSS 0.052845f
C2822 DVDD.n2328 DVSS 0.052845f
C2823 DVDD.n2329 DVSS 0.052845f
C2824 DVDD.n2330 DVSS 0.052845f
C2825 DVDD.n2331 DVSS 0.052845f
C2826 DVDD.n2332 DVSS 0.052845f
C2827 DVDD.n2333 DVSS 0.052845f
C2828 DVDD.n2334 DVSS 0.052845f
C2829 DVDD.n2335 DVSS 0.052845f
C2830 DVDD.n2336 DVSS 0.052845f
C2831 DVDD.n2337 DVSS 0.052845f
C2832 DVDD.n2338 DVSS 0.052845f
C2833 DVDD.n2339 DVSS 0.052845f
C2834 DVDD.n2340 DVSS 0.052845f
C2835 DVDD.n2341 DVSS 0.052845f
C2836 DVDD.n2342 DVSS 0.052845f
C2837 DVDD.n2343 DVSS 0.052845f
C2838 DVDD.n2344 DVSS 0.052845f
C2839 DVDD.n2345 DVSS 0.052845f
C2840 DVDD.n2346 DVSS 0.052845f
C2841 DVDD.n2347 DVSS 0.052845f
C2842 DVDD.n2348 DVSS 0.046891f
C2843 DVDD.n2349 DVSS 0.046891f
C2844 DVDD.n2350 DVSS 0.063637f
C2845 DVDD.n2351 DVSS 0.100852f
C2846 DVDD.n2352 DVSS 0.032377f
C2847 DVDD.n2353 DVSS 0.032377f
C2848 DVDD.n2354 DVSS 0.052845f
C2849 DVDD.n2355 DVSS 0.052845f
C2850 DVDD.n2356 DVSS 0.052845f
C2851 DVDD.n2357 DVSS 0.052845f
C2852 DVDD.n2358 DVSS 0.052845f
C2853 DVDD.n2359 DVSS 0.052845f
C2854 DVDD.n2360 DVSS 0.052845f
C2855 DVDD.n2361 DVSS 0.052845f
C2856 DVDD.n2362 DVSS 0.052845f
C2857 DVDD.n2363 DVSS 0.052845f
C2858 DVDD.n2364 DVSS 0.052845f
C2859 DVDD.n2365 DVSS 0.052845f
C2860 DVDD.n2366 DVSS 0.052845f
C2861 DVDD.n2367 DVSS 0.052845f
C2862 DVDD.n2368 DVSS 0.031074f
C2863 DVDD.n2369 DVSS 0.026423f
C2864 DVDD.n2370 DVSS 0.004156f
C2865 DVDD.n2371 DVSS 0.024376f
C2866 DVDD.n2372 DVSS 0.012068f
C2867 DVDD.n2373 DVSS 0.02512f
C2868 DVDD.n2374 DVSS 0.023073f
C2869 DVDD.n2375 DVSS 0.052845f
C2870 DVDD.n2376 DVSS 0.052845f
C2871 DVDD.n2377 DVSS 0.031819f
C2872 DVDD.n2378 DVSS 0.052845f
C2873 DVDD.n2379 DVSS 0.052845f
C2874 DVDD.n2380 DVSS 0.052845f
C2875 DVDD.n2381 DVSS 0.052845f
C2876 DVDD.n2382 DVSS 0.052845f
C2877 DVDD.n2383 DVSS 0.052845f
C2878 DVDD.n2384 DVSS 0.052845f
C2879 DVDD.n2385 DVSS 0.052845f
C2880 DVDD.n2386 DVSS 0.052845f
C2881 DVDD.n2387 DVSS 0.052845f
C2882 DVDD.n2388 DVSS 0.052845f
C2883 DVDD.n2389 DVSS 0.052845f
C2884 DVDD.n2390 DVSS 0.052845f
C2885 DVDD.n2391 DVSS 0.045402f
C2886 DVDD.n2392 DVSS 0.045402f
C2887 DVDD.n2393 DVSS 0.100852f
C2888 DVDD.n2394 DVSS 0.033866f
C2889 DVDD.n2395 DVSS 0.052845f
C2890 DVDD.n2396 DVSS 0.052845f
C2891 DVDD.n2397 DVSS 0.052845f
C2892 DVDD.n2398 DVSS 0.052845f
C2893 DVDD.n2399 DVSS 0.052845f
C2894 DVDD.n2400 DVSS 0.052845f
C2895 DVDD.n2401 DVSS 0.052845f
C2896 DVDD.n2402 DVSS 0.052845f
C2897 DVDD.n2403 DVSS 0.052845f
C2898 DVDD.n2404 DVSS 0.052845f
C2899 DVDD.n2405 DVSS 0.052845f
C2900 DVDD.n2406 DVSS 0.052845f
C2901 DVDD.n2407 DVSS 0.052845f
C2902 DVDD.n2408 DVSS 0.052845f
C2903 DVDD.n2409 DVSS 0.052845f
C2904 DVDD.n2410 DVSS 0.052845f
C2905 DVDD.n2411 DVSS 0.052845f
C2906 DVDD.n2412 DVSS 0.052845f
C2907 DVDD.n2413 DVSS 0.052845f
C2908 DVDD.n2414 DVSS 0.052845f
C2909 DVDD.n2415 DVSS 0.052845f
C2910 DVDD.n2416 DVSS 0.052845f
C2911 DVDD.n2417 DVSS 0.052845f
C2912 DVDD.n2418 DVSS 0.052845f
C2913 DVDD.n2419 DVSS 0.052845f
C2914 DVDD.n2420 DVSS 0.052845f
C2915 DVDD.n2421 DVSS 0.052845f
C2916 DVDD.n2422 DVSS 0.052845f
C2917 DVDD.n2423 DVSS 0.052845f
C2918 DVDD.n2424 DVSS 0.052845f
C2919 DVDD.n2425 DVSS 0.042611f
C2920 DVDD.n2427 DVSS 0.001538f
C2921 DVDD.n2428 DVSS 0.003076f
C2922 DVDD.n2429 DVSS 0.003076f
C2923 DVDD.n2430 DVSS 0.003076f
C2924 DVDD.n2431 DVSS 0.003076f
C2925 DVDD.n2432 DVSS 0.001538f
C2926 DVDD.n2433 DVSS 0.001538f
C2927 DVDD.n2434 DVSS 0.001538f
C2928 DVDD.n2435 DVSS 0.00289f
C2929 DVDD.n2436 DVSS 0.011041f
C2930 DVDD.n2437 DVSS 0.004503f
C2931 DVDD.n2438 DVSS 0.026423f
C2932 DVDD.n2439 DVSS 0.001538f
C2933 DVDD.n2440 DVSS 0.001551f
C2934 DVDD.n2441 DVSS 0.026423f
C2935 DVDD.n2442 DVSS 0.00299f
C2936 DVDD.n2443 DVSS 0.008262f
C2937 DVDD.n2444 DVSS 0.027687f
C2938 DVDD.n2445 DVSS 0.01188f
C2939 DVDD.t98 DVSS 0.032253f
C2940 DVDD.t111 DVSS 0.032253f
C2941 DVDD.n2446 DVSS 0.064506f
C2942 DVDD.n2447 DVSS 0.011628f
C2943 DVDD.n2448 DVSS 0.027944f
C2944 DVDD.n2449 DVSS 0.008261f
C2945 DVDD.n2450 DVSS 0.00299f
C2946 DVDD.n2451 DVSS 0.001538f
C2947 DVDD.n2452 DVSS 0.00289f
C2948 DVDD.n2453 DVSS 0.01104f
C2949 DVDD.n2454 DVSS 0.001538f
C2950 DVDD.n2455 DVSS 0.004503f
C2951 DVDD.n2456 DVSS 0.026423f
C2952 DVDD.n2457 DVSS 0.023073f
C2953 DVDD.n2458 DVSS 0.052845f
C2954 DVDD.n2459 DVSS 0.052845f
C2955 DVDD.n2460 DVSS 0.043355f
C2956 DVDD.n2461 DVSS 0.052845f
C2957 DVDD.n2462 DVSS 0.052845f
C2958 DVDD.n2463 DVSS 0.052845f
C2959 DVDD.n2464 DVSS 0.052845f
C2960 DVDD.n2465 DVSS 0.052845f
C2961 DVDD.n2466 DVSS 0.052845f
C2962 DVDD.n2467 DVSS 0.052845f
C2963 DVDD.n2468 DVSS 0.052845f
C2964 DVDD.n2469 DVSS 0.052845f
C2965 DVDD.n2470 DVSS 0.052845f
C2966 DVDD.n2471 DVSS 0.052845f
C2967 DVDD.n2472 DVSS 0.052845f
C2968 DVDD.n2473 DVSS 0.052845f
C2969 DVDD.n2474 DVSS 0.052845f
C2970 DVDD.n2475 DVSS 0.052845f
C2971 DVDD.n2476 DVSS 0.052845f
C2972 DVDD.n2477 DVSS 0.052845f
C2973 DVDD.n2478 DVSS 0.052845f
C2974 DVDD.n2479 DVSS 0.052845f
C2975 DVDD.n2480 DVSS 0.052845f
C2976 DVDD.n2481 DVSS 0.052845f
C2977 DVDD.n2482 DVSS 0.052845f
C2978 DVDD.n2483 DVSS 0.052845f
C2979 DVDD.n2484 DVSS 0.052845f
C2980 DVDD.n2485 DVSS 0.052845f
C2981 DVDD.n2486 DVSS 0.052845f
C2982 DVDD.n2487 DVSS 0.052845f
C2983 DVDD.n2488 DVSS 0.052845f
C2984 DVDD.n2489 DVSS 0.052845f
C2985 DVDD.n2490 DVSS 0.046891f
C2986 DVDD.n2491 DVSS 0.046891f
C2987 DVDD.n2492 DVSS 0.100852f
C2988 DVDD.n2493 DVSS 0.063637f
C2989 DVDD.n2494 DVSS 0.032377f
C2990 DVDD.n2495 DVSS 0.032377f
C2991 DVDD.n2496 DVSS 0.052845f
C2992 DVDD.n2497 DVSS 0.052845f
C2993 DVDD.n2498 DVSS 0.052845f
C2994 DVDD.n2499 DVSS 0.052845f
C2995 DVDD.n2500 DVSS 0.052845f
C2996 DVDD.n2501 DVSS 0.052845f
C2997 DVDD.n2502 DVSS 0.052845f
C2998 DVDD.n2503 DVSS 0.052845f
C2999 DVDD.n2504 DVSS 0.052845f
C3000 DVDD.n2505 DVSS 0.052845f
C3001 DVDD.n2506 DVSS 0.052845f
C3002 DVDD.n2507 DVSS 0.052845f
C3003 DVDD.n2508 DVSS 0.052845f
C3004 DVDD.n2509 DVSS 0.052845f
C3005 DVDD.n2510 DVSS 0.031074f
C3006 DVDD.n2511 DVSS 0.008245f
C3007 DVDD.n2513 DVSS 0.001538f
C3008 DVDD.n2514 DVSS 0.001625f
C3009 DVDD.n2515 DVSS 0.00299f
C3010 DVDD.n2516 DVSS 0.008262f
C3011 DVDD.n2517 DVSS 0.027687f
C3012 DVDD.n2518 DVSS 0.01188f
C3013 DVDD.n2519 DVSS 0.001625f
C3014 DVDD.n2520 DVSS 0.00299f
C3015 DVDD.n2521 DVSS 0.008261f
C3016 DVDD.n2522 DVSS 0.001538f
C3017 DVDD.n2523 DVSS 0.027944f
C3018 DVDD.t96 DVSS 0.032253f
C3019 DVDD.t140 DVSS 0.032253f
C3020 DVDD.n2524 DVSS 0.064506f
C3021 DVDD.n2525 DVSS 0.011628f
C3022 DVDD.n2526 DVSS 0.004122f
C3023 DVDD.n2527 DVSS 0.004355f
C3024 DVDD.n2529 DVSS 0.008212f
C3025 DVDD.n2530 DVSS 0.001538f
C3026 DVDD.n2531 DVSS 0.001551f
C3027 DVDD.n2532 DVSS 0.008262f
C3028 DVDD.n2533 DVSS 0.027687f
C3029 DVDD.n2534 DVSS 0.01188f
C3030 DVDD.n2535 DVSS 0.001551f
C3031 DVDD.n2536 DVSS 0.008261f
C3032 DVDD.n2537 DVSS 0.001538f
C3033 DVDD.n2538 DVSS 0.027944f
C3034 DVDD.t109 DVSS 0.032253f
C3035 DVDD.t83 DVSS 0.032253f
C3036 DVDD.n2539 DVSS 0.064506f
C3037 DVDD.n2540 DVSS 0.011628f
C3038 DVDD.n2541 DVSS 0.004122f
C3039 DVDD.n2542 DVSS 0.004156f
C3040 DVDD.n2544 DVSS 0.008245f
C3041 DVDD.n2546 DVSS 0.008245f
C3042 DVDD.n2548 DVSS 0.001538f
C3043 DVDD.n2549 DVSS 0.002965f
C3044 DVDD.n2550 DVSS 0.008262f
C3045 DVDD.n2551 DVSS 0.027687f
C3046 DVDD.n2552 DVSS 0.01188f
C3047 DVDD.n2553 DVSS 0.002965f
C3048 DVDD.n2554 DVSS 0.008261f
C3049 DVDD.n2555 DVSS 0.001538f
C3050 DVDD.n2556 DVSS 0.027944f
C3051 DVDD.t97 DVSS 0.032253f
C3052 DVDD.t107 DVSS 0.032253f
C3053 DVDD.n2557 DVSS 0.064506f
C3054 DVDD.n2558 DVSS 0.011628f
C3055 DVDD.n2559 DVSS 0.004122f
C3056 DVDD.n2561 DVSS 0.004422f
C3057 DVDD.n2563 DVSS 0.004954f
C3058 DVDD.n2564 DVSS 0.026423f
C3059 DVDD.n2565 DVSS 0.049203f
C3060 DVDD.t142 DVSS 0.032253f
C3061 DVDD.t124 DVSS 0.032253f
C3062 DVDD.n2566 DVSS 0.064506f
C3063 DVDD.n2567 DVSS 0.011628f
C3064 DVDD.n2568 DVSS 0.064329f
C3065 DVDD.n2569 DVSS 0.016855f
C3066 DVDD.n2570 DVSS 0.01188f
C3067 DVDD.t133 DVSS 0.032253f
C3068 DVDD.t85 DVSS 0.032253f
C3069 DVDD.n2571 DVSS 0.064506f
C3070 DVDD.n2572 DVSS 0.011628f
C3071 DVDD.n2573 DVSS 0.027944f
C3072 DVDD.n2574 DVSS 0.001538f
C3073 DVDD.n2575 DVSS 0.010767f
C3074 DVDD.n2576 DVSS 0.002642f
C3075 DVDD.n2577 DVSS 0.002741f
C3076 DVDD.n2578 DVSS 0.018322f
C3077 DVDD.n2579 DVSS 0.003076f
C3078 DVDD.n2580 DVSS 0.001873f
C3079 DVDD.n2581 DVSS 0.003076f
C3080 DVDD.n2582 DVSS 0.001538f
C3081 DVDD.n2583 DVSS 0.020233f
C3082 DVDD.n2584 DVSS 0.001538f
C3083 DVDD.n2585 DVSS 0.004122f
C3084 DVDD.n2586 DVSS 0.001538f
C3085 DVDD.n2587 DVSS 0.002642f
C3086 DVDD.n2588 DVSS 0.001538f
C3087 DVDD.n2589 DVSS 0.010767f
C3088 DVDD.n2590 DVSS 0.002741f
C3089 DVDD.n2591 DVSS 0.019885f
C3090 DVDD.n2592 DVSS 0.001774f
C3091 DVDD.n2593 DVSS 0.003076f
C3092 DVDD.t103 DVSS 0.032253f
C3093 DVDD.t87 DVSS 0.032253f
C3094 DVDD.n2594 DVSS 0.064506f
C3095 DVDD.n2595 DVSS 0.010767f
C3096 DVDD.n2596 DVSS 0.007081f
C3097 DVDD.n2597 DVSS 0.008245f
C3098 DVDD.n2599 DVSS 0.008245f
C3099 DVDD.n2601 DVSS 0.011723f
C3100 DVDD.n2603 DVSS 0.007347f
C3101 DVDD.n2604 DVSS 0.008261f
C3102 DVDD.n2605 DVSS 0.002741f
C3103 DVDD.n2606 DVSS 0.001538f
C3104 DVDD.n2607 DVSS 0.010767f
C3105 DVDD.n2608 DVSS 0.002642f
C3106 DVDD.n2609 DVSS 0.014501f
C3107 DVDD.n2610 DVSS 0.006289f
C3108 DVDD.n2611 DVSS 0.001774f
C3109 DVDD.n2612 DVSS 0.003076f
C3110 DVDD.n2613 DVSS 0.003076f
C3111 DVDD.n2614 DVSS 0.001972f
C3112 DVDD.n2615 DVSS 0.024661f
C3113 DVDD.n2616 DVSS 0.024661f
C3114 DVDD.n2617 DVSS 0.024661f
C3115 DVDD.n2618 DVSS 0.024661f
C3116 DVDD.n2619 DVSS 0.024661f
C3117 DVDD.n2620 DVSS 0.024661f
C3118 DVDD.n2621 DVSS 0.024661f
C3119 DVDD.n2622 DVSS 0.024661f
C3120 DVDD.n2623 DVSS 0.024661f
C3121 DVDD.n2624 DVSS 0.024661f
C3122 DVDD.n2625 DVSS 0.024661f
C3123 DVDD.n2626 DVSS 0.024661f
C3124 DVDD.n2627 DVSS 0.024661f
C3125 DVDD.n2628 DVSS 0.024661f
C3126 DVDD.n2629 DVSS 0.024661f
C3127 DVDD.n2630 DVSS 0.024661f
C3128 DVDD.n2631 DVSS 0.024661f
C3129 DVDD.n2632 DVSS 0.024661f
C3130 DVDD.n2633 DVSS 0.024661f
C3131 DVDD.n2634 DVSS 0.024661f
C3132 DVDD.n2635 DVSS 0.024661f
C3133 DVDD.n2636 DVSS 0.024661f
C3134 DVDD.n2637 DVSS 0.024661f
C3135 DVDD.n2638 DVSS 0.024661f
C3136 DVDD.n2639 DVSS 0.024661f
C3137 DVDD.n2640 DVSS 0.024661f
C3138 DVDD.n2641 DVSS 0.024661f
C3139 DVDD.n2642 DVSS 0.024661f
C3140 DVDD.n2643 DVSS 0.024661f
C3141 DVDD.n2644 DVSS 0.024661f
C3142 DVDD.n2645 DVSS 0.024661f
C3143 DVDD.n2646 DVSS 0.024661f
C3144 DVDD.n2647 DVSS 0.024661f
C3145 DVDD.n2648 DVSS 0.024661f
C3146 DVDD.n2649 DVSS 0.024661f
C3147 DVDD.n2650 DVSS 0.024661f
C3148 DVDD.n2651 DVSS 0.024661f
C3149 DVDD.n2652 DVSS 0.024661f
C3150 DVDD.n2653 DVSS 0.024661f
C3151 DVDD.n2654 DVSS 0.024661f
C3152 DVDD.n2655 DVSS 0.024661f
C3153 DVDD.n2656 DVSS 0.024661f
C3154 DVDD.n2657 DVSS 0.024661f
C3155 DVDD.n2658 DVSS 0.024661f
C3156 DVDD.n2659 DVSS 0.024661f
C3157 DVDD.n2660 DVSS 0.024661f
C3158 DVDD.n2661 DVSS 0.024661f
C3159 DVDD.n2662 DVSS 0.024661f
C3160 DVDD.n2663 DVSS 0.024661f
C3161 DVDD.n2664 DVSS 0.024661f
C3162 DVDD.n2665 DVSS 0.024661f
C3163 DVDD.n2666 DVSS 0.024661f
C3164 DVDD.n2667 DVSS 0.024661f
C3165 DVDD.n2668 DVSS 0.024661f
C3166 DVDD.n2669 DVSS 0.024661f
C3167 DVDD.n2670 DVSS 0.024661f
C3168 DVDD.n2671 DVSS 0.024661f
C3169 DVDD.n2672 DVSS 0.024661f
C3170 DVDD.n2673 DVSS 0.024661f
C3171 DVDD.n2674 DVSS 0.024661f
C3172 DVDD.n2675 DVSS 0.024661f
C3173 DVDD.n2676 DVSS 0.024661f
C3174 DVDD.n2677 DVSS 0.024661f
C3175 DVDD.n2678 DVSS 0.024661f
C3176 DVDD.n2679 DVSS 0.024661f
C3177 DVDD.n2680 DVSS 0.024661f
C3178 DVDD.n2681 DVSS 0.024661f
C3179 DVDD.n2682 DVSS 0.024661f
C3180 DVDD.n2683 DVSS 0.024661f
C3181 DVDD.n2684 DVSS 0.118858f
C3182 DVDD.n2685 DVSS 0.032461f
C3183 DVDD.n2686 DVSS 0.002779f
C3184 DVDD.n2687 DVSS 0.02223f
C3185 DVDD.n2688 DVSS 0.02223f
C3186 DVDD.n2689 DVSS 0.02223f
C3187 DVDD.n2690 DVSS 0.024661f
C3188 DVDD.n2691 DVSS 0.024661f
C3189 DVDD.n2692 DVSS 0.024661f
C3190 DVDD.n2693 DVSS 0.024661f
C3191 DVDD.n2694 DVSS 0.024661f
C3192 DVDD.n2695 DVSS 0.024661f
C3193 DVDD.n2696 DVSS 0.024661f
C3194 DVDD.n2697 DVSS 0.024661f
C3195 DVDD.n2698 DVSS 0.024661f
C3196 DVDD.n2699 DVSS 0.024661f
C3197 DVDD.n2700 DVSS 0.024661f
C3198 DVDD.n2701 DVSS 0.024661f
C3199 DVDD.n2702 DVSS 0.024661f
C3200 DVDD.n2703 DVSS 0.024661f
C3201 DVDD.n2704 DVSS 0.024661f
C3202 DVDD.n2705 DVSS 0.024661f
C3203 DVDD.n2706 DVSS 0.024661f
C3204 DVDD.n2707 DVSS 0.024661f
C3205 DVDD.n2708 DVSS 0.024661f
C3206 DVDD.n2709 DVSS 0.024661f
C3207 DVDD.n2710 DVSS 0.024661f
C3208 DVDD.n2711 DVSS 0.024661f
C3209 DVDD.n2712 DVSS 0.024661f
C3210 DVDD.n2713 DVSS 0.024661f
C3211 DVDD.n2714 DVSS 0.024661f
C3212 DVDD.n2715 DVSS 0.024661f
C3213 DVDD.n2716 DVSS 0.024661f
C3214 DVDD.n2717 DVSS 0.024661f
C3215 DVDD.n2718 DVSS 0.024661f
C3216 DVDD.n2719 DVSS 0.024661f
C3217 DVDD.n2720 DVSS 0.024661f
C3218 DVDD.n2721 DVSS 0.024661f
C3219 DVDD.n2722 DVSS 0.024661f
C3220 DVDD.n2723 DVSS 0.024661f
C3221 DVDD.n2724 DVSS 0.024661f
C3222 DVDD.n2725 DVSS 0.024661f
C3223 DVDD.n2726 DVSS 0.024661f
C3224 DVDD.n2727 DVSS 0.024661f
C3225 DVDD.n2728 DVSS 0.024661f
C3226 DVDD.n2729 DVSS 0.024661f
C3227 DVDD.n2730 DVSS 0.024661f
C3228 DVDD.n2731 DVSS 0.024661f
C3229 DVDD.n2732 DVSS 0.024661f
C3230 DVDD.n2733 DVSS 0.024661f
C3231 DVDD.n2734 DVSS 0.024661f
C3232 DVDD.n2735 DVSS 0.024661f
C3233 DVDD.n2736 DVSS 0.024661f
C3234 DVDD.n2737 DVSS 0.024661f
C3235 DVDD.n2738 DVSS 0.024661f
C3236 DVDD.n2739 DVSS 0.024661f
C3237 DVDD.n2740 DVSS 0.024661f
C3238 DVDD.n2741 DVSS 0.024661f
C3239 DVDD.n2742 DVSS 0.024661f
C3240 DVDD.n2743 DVSS 0.024661f
C3241 DVDD.n2744 DVSS 0.024661f
C3242 DVDD.n2745 DVSS 0.024661f
C3243 DVDD.n2746 DVSS 0.024661f
C3244 DVDD.n2747 DVSS 0.024053f
C3245 DVDD.n2748 DVSS 0.001538f
C3246 DVDD.n2749 DVSS 0.001538f
C3247 DVDD.n2750 DVSS 0.001538f
C3248 DVDD.n2751 DVSS 0.01233f
C3249 DVDD.n2752 DVSS 0.001538f
C3250 DVDD.n2753 DVSS 0.001538f
C3251 DVDD.n2754 DVSS 0.01233f
C3252 DVDD.n2755 DVSS 0.001873f
C3253 DVDD.n2756 DVSS 0.001538f
C3254 DVDD.n2757 DVSS 0.027944f
C3255 DVDD.n2758 DVSS 0.011628f
C3256 DVDD.n2759 DVSS 0.004122f
C3257 DVDD.n2760 DVSS 0.01188f
C3258 DVDD.n2761 DVSS 0.001538f
C3259 DVDD.n2762 DVSS 0.027687f
C3260 DVDD.n2763 DVSS 0.008262f
C3261 DVDD.n2764 DVSS 0.001873f
C3262 DVDD.n2765 DVSS 0.003076f
C3263 DVDD.n2766 DVSS 0.018831f
C3264 DVDD.t79 DVSS 0.032253f
C3265 DVDD.t94 DVSS 0.032253f
C3266 DVDD.n2767 DVSS 0.064506f
C3267 DVDD.n2768 DVSS 0.011628f
C3268 DVDD.n2769 DVSS 0.01188f
C3269 DVDD.n2770 DVSS 0.027687f
C3270 DVDD.n2771 DVSS 0.027687f
C3271 DVDD.n2772 DVSS 0.027687f
C3272 DVDD.n2773 DVSS 0.027687f
C3273 DVDD.n2774 DVSS 0.027687f
C3274 DVDD.n2775 DVSS 0.027687f
C3275 DVDD.n2776 DVSS 0.027687f
C3276 DVDD.n2777 DVSS 0.027687f
C3277 DVDD.n2778 DVSS 0.027687f
C3278 DVDD.n2779 DVSS 0.027687f
C3279 DVDD.n2780 DVSS 0.027687f
C3280 DVDD.n2781 DVSS 0.027687f
C3281 DVDD.t75 DVSS 0.032253f
C3282 DVDD.t129 DVSS 0.032253f
C3283 DVDD.n2782 DVSS 0.064506f
C3284 DVDD.n2783 DVSS 0.01188f
C3285 DVDD.t122 DVSS 0.032253f
C3286 DVDD.t105 DVSS 0.032253f
C3287 DVDD.n2784 DVSS 0.064506f
C3288 DVDD.n2785 DVSS 0.011628f
C3289 DVDD.n2786 DVSS 0.032447f
C3290 DVDD.n2787 DVSS 0.01188f
C3291 DVDD.t101 DVSS 0.032253f
C3292 DVDD.t102 DVSS 0.032253f
C3293 DVDD.n2788 DVSS 0.064506f
C3294 DVDD.n2789 DVSS 0.011628f
C3295 DVDD.n2790 DVSS 0.032447f
C3296 DVDD.n2791 DVSS 0.01188f
C3297 DVDD.t93 DVSS 0.032253f
C3298 DVDD.t148 DVSS 0.032253f
C3299 DVDD.n2792 DVSS 0.064506f
C3300 DVDD.n2793 DVSS 0.011628f
C3301 DVDD.n2794 DVSS 0.032447f
C3302 DVDD.n2795 DVSS 0.01188f
C3303 DVDD.t82 DVSS 0.032253f
C3304 DVDD.t114 DVSS 0.032253f
C3305 DVDD.n2796 DVSS 0.064506f
C3306 DVDD.n2797 DVSS 0.011628f
C3307 DVDD.n2798 DVSS 0.065427f
C3308 DVDD.n2799 DVSS 0.01188f
C3309 DVDD.t121 DVSS 0.032253f
C3310 DVDD.t152 DVSS 0.032253f
C3311 DVDD.n2800 DVSS 0.064506f
C3312 DVDD.n2801 DVSS 0.011628f
C3313 DVDD.n2802 DVSS 0.065427f
C3314 DVDD.n2803 DVSS 0.01188f
C3315 DVDD.t125 DVSS 0.032253f
C3316 DVDD.t154 DVSS 0.032253f
C3317 DVDD.n2804 DVSS 0.064506f
C3318 DVDD.n2805 DVSS 0.011628f
C3319 DVDD.n2806 DVSS 0.032447f
C3320 DVDD.n2807 DVSS 0.01188f
C3321 DVDD.t116 DVSS 0.032253f
C3322 DVDD.t134 DVSS 0.032253f
C3323 DVDD.n2808 DVSS 0.064506f
C3324 DVDD.n2809 DVSS 0.011628f
C3325 DVDD.n2810 DVSS 0.032447f
C3326 DVDD.n2811 DVSS 0.01188f
C3327 DVDD.t127 DVSS 0.032253f
C3328 DVDD.t149 DVSS 0.032253f
C3329 DVDD.n2812 DVSS 0.064506f
C3330 DVDD.n2813 DVSS 0.011628f
C3331 DVDD.n2814 DVSS 0.032447f
C3332 DVDD.n2815 DVSS 0.01188f
C3333 DVDD.t115 DVSS 0.032253f
C3334 DVDD.t138 DVSS 0.032253f
C3335 DVDD.n2816 DVSS 0.064506f
C3336 DVDD.n2817 DVSS 0.011628f
C3337 DVDD.n2818 DVSS 0.032447f
C3338 DVDD.n2819 DVSS 0.01188f
C3339 DVDD.t84 DVSS 0.032253f
C3340 DVDD.t81 DVSS 0.032253f
C3341 DVDD.n2820 DVSS 0.064506f
C3342 DVDD.n2821 DVSS 0.011628f
C3343 DVDD.n2822 DVSS 0.032447f
C3344 DVDD.n2823 DVSS 0.01188f
C3345 DVDD.t88 DVSS 0.032253f
C3346 DVDD.t123 DVSS 0.032253f
C3347 DVDD.n2824 DVSS 0.064506f
C3348 DVDD.n2825 DVSS 0.011628f
C3349 DVDD.n2826 DVSS 0.032447f
C3350 DVDD.n2827 DVSS 0.011628f
C3351 DVDD.n2828 DVSS 0.032447f
C3352 DVDD.n2829 DVSS 0.01188f
C3353 DVDD.n2830 DVSS 0.018831f
C3354 DVDD.n2831 DVSS 0.018831f
C3355 DVDD.n2832 DVSS 0.018831f
C3356 DVDD.n2833 DVSS 0.031137f
C3357 DVDD.n2834 DVSS 0.031137f
C3358 DVDD.n2835 DVSS 0.018831f
C3359 DVDD.n2836 DVSS 0.018831f
C3360 DVDD.n2837 DVSS 0.018831f
C3361 DVDD.n2838 DVSS 0.018831f
C3362 DVDD.n2839 DVSS 0.018831f
C3363 DVDD.n2840 DVSS 0.018831f
C3364 DVDD.n2841 DVSS 0.018831f
C3365 DVDD.n2842 DVSS 0.027687f
C3366 DVDD.t137 DVSS 0.032253f
C3367 DVDD.t108 DVSS 0.032253f
C3368 DVDD.n2843 DVSS 0.064506f
C3369 DVDD.n2844 DVSS 0.011628f
C3370 DVDD.n2845 DVSS 0.01188f
C3371 DVDD.n2846 DVSS 0.027687f
C3372 DVDD.n2847 DVSS 0.012107f
C3373 DVDD.n2848 DVSS 0.012107f
C3374 DVDD.n2849 DVSS 0.012107f
C3375 DVDD.n2850 DVSS 0.012107f
C3376 DVDD.n2851 DVSS 0.012107f
C3377 DVDD.n2852 DVSS 0.012107f
C3378 DVDD.n2853 DVSS 0.012107f
C3379 DVDD.n2854 DVSS 0.012107f
C3380 DVDD.n2855 DVSS 0.024413f
C3381 DVDD.n2856 DVSS 0.024413f
C3382 DVDD.n2857 DVSS 0.012107f
C3383 DVDD.n2858 DVSS 0.012107f
C3384 DVDD.n2859 DVSS 0.012107f
C3385 DVDD.n2860 DVSS 0.012107f
C3386 DVDD.n2861 DVSS 0.008597f
C3387 DVDD.n2862 DVSS 0.027687f
C3388 DVDD.n2863 DVSS 0.015321f
C3389 DVDD.n2864 DVSS 0.385829f
C3390 DVDD.n2865 DVSS 0.024661f
C3391 DVDD.n2866 DVSS 0.024661f
C3392 DVDD.n2867 DVSS 0.024661f
C3393 DVDD.n2868 DVSS 0.024661f
C3394 DVDD.n2869 DVSS 0.024661f
C3395 DVDD.n2870 DVSS 0.024661f
C3396 DVDD.n2871 DVSS 0.024661f
C3397 DVDD.n2872 DVSS 0.024661f
C3398 DVDD.n2873 DVSS 0.024661f
C3399 DVDD.n2874 DVSS 0.024661f
C3400 DVDD.n2875 DVSS 0.024661f
C3401 DVDD.n2876 DVSS 0.024661f
C3402 DVDD.n2877 DVSS 0.024661f
C3403 DVDD.n2878 DVSS 0.024661f
C3404 DVDD.n2879 DVSS 0.024661f
C3405 DVDD.n2880 DVSS 0.024661f
C3406 DVDD.n2881 DVSS 0.024661f
C3407 DVDD.n2882 DVSS 0.024661f
C3408 DVDD.n2883 DVSS 0.024661f
C3409 DVDD.n2884 DVSS 0.024661f
C3410 DVDD.n2885 DVSS 0.024661f
C3411 DVDD.n2886 DVSS 0.024661f
C3412 DVDD.n2887 DVSS 0.024661f
C3413 DVDD.n2888 DVSS 0.024661f
C3414 DVDD.n2889 DVSS 0.024661f
C3415 DVDD.n2890 DVSS 0.024661f
C3416 DVDD.n2891 DVSS 0.024661f
C3417 DVDD.n2892 DVSS 0.024661f
C3418 DVDD.n2893 DVSS 0.024661f
C3419 DVDD.n2894 DVSS 0.024661f
C3420 DVDD.n2895 DVSS 0.024661f
C3421 DVDD.n2896 DVSS 0.024661f
C3422 DVDD.n2897 DVSS 0.024661f
C3423 DVDD.n2898 DVSS 0.024661f
C3424 DVDD.n2899 DVSS 0.024661f
C3425 DVDD.n2900 DVSS 0.024661f
C3426 DVDD.n2901 DVSS 0.024661f
C3427 DVDD.n2902 DVSS 0.024661f
C3428 DVDD.n2903 DVSS 0.024661f
C3429 DVDD.n2904 DVSS 0.024661f
C3430 DVDD.n2905 DVSS 0.080215f
C3431 DVDD.n2906 DVSS 0.588441f
C3432 DVDD.n2907 DVSS 0.001538f
C3433 DVDD.n2908 DVSS 0.001538f
C3434 DVDD.n2909 DVSS 0.001538f
C3435 DVDD.n2910 DVSS 0.001538f
C3436 DVDD.n2911 DVSS 0.342943f
C3437 DVDD.n2912 DVSS 0.004081f
C3438 DVDD.n2913 DVSS 0.001538f
C3439 DVDD.n2914 DVSS 0.01233f
C3440 DVDD.n2915 DVSS 0.001972f
C3441 DVDD.n2916 DVSS 0.008262f
C3442 DVDD.n2917 DVSS 0.027687f
C3443 DVDD.n2918 DVSS 0.01188f
C3444 DVDD.t80 DVSS 0.032253f
C3445 DVDD.t91 DVSS 0.032253f
C3446 DVDD.n2919 DVSS 0.064506f
C3447 DVDD.n2920 DVSS 0.011628f
C3448 DVDD.n2921 DVSS 0.027944f
C3449 DVDD.n2922 DVSS 0.008261f
C3450 DVDD.n2923 DVSS 0.001972f
C3451 DVDD.n2924 DVSS 0.001538f
C3452 DVDD.n2925 DVSS 0.001538f
C3453 DVDD.n2926 DVSS 0.001538f
C3454 DVDD.n2927 DVSS 0.01233f
C3455 DVDD.n2928 DVSS 0.001538f
C3456 DVDD.n2929 DVSS 0.004081f
C3457 DVDD.n2930 DVSS 0.01233f
C3458 DVDD.n2931 DVSS 0.001774f
C3459 DVDD.n2932 DVSS 0.013012f
C3460 DVDD.n2933 DVSS 0.030726f
C3461 DVDD.n2934 DVSS 0.018359f
C3462 DVDD.n2935 DVSS 0.026423f
C3463 DVDD.n2936 DVSS 0.001749f
C3464 DVDD.n2937 DVSS 0.008261f
C3465 DVDD.n2938 DVSS 0.001538f
C3466 DVDD.n2939 DVSS 0.027944f
C3467 DVDD.n2940 DVSS 0.011628f
C3468 DVDD.n2941 DVSS 0.004122f
C3469 DVDD.n2942 DVSS 0.01188f
C3470 DVDD.n2943 DVSS 0.008262f
C3471 DVDD.n2944 DVSS 0.027687f
C3472 DVDD.n2945 DVSS 0.001538f
C3473 DVDD.n2946 DVSS 0.001749f
C3474 DVDD.n2947 DVSS 0.003076f
C3475 DVDD.n2948 DVSS 0.001848f
C3476 DVDD.n2949 DVSS 0.026423f
C3477 DVDD.n2950 DVSS 0.003076f
C3478 DVDD.n2951 DVSS 0.001538f
C3479 DVDD.n2952 DVSS 0.026423f
C3480 DVDD.n2953 DVSS 0.00289f
C3481 DVDD.n2954 DVSS 0.004317f
C3482 DVDD.n2955 DVSS 0.004503f
C3483 DVDD.n2956 DVSS 0.026423f
C3484 DVDD.n2957 DVSS 0.001538f
C3485 DVDD.n2958 DVSS 0.001551f
C3486 DVDD.n2959 DVSS 0.026423f
C3487 DVDD.n2960 DVSS 0.005768f
C3488 DVDD.n2961 DVSS 0.004317f
C3489 DVDD.n2962 DVSS 0.001625f
C3490 DVDD.n2963 DVSS 0.026423f
C3491 DVDD.n2964 DVSS 0.002394f
C3492 DVDD.n2965 DVSS 0.004317f
C3493 DVDD.n2966 DVSS 0.027687f
C3494 DVDD.n2967 DVSS 0.011041f
C3495 DVDD.n2968 DVSS 0.004999f
C3496 DVDD.n2969 DVSS 0.026423f
C3497 DVDD.n2970 DVSS 0.025778f
C3498 DVDD.n2971 DVSS 0.025778f
C3499 DVDD.n2972 DVSS 0.014092f
C3500 DVDD.n2973 DVSS 0.012306f
C3501 DVDD.n2974 DVSS 0.014092f
C3502 DVDD.n2975 DVSS 0.016573f
C3503 DVDD.n2976 DVSS 0.02342f
C3504 DVDD.n2977 DVSS 0.182359f
C3505 DVDD.n2978 DVSS 0.043914f
C3506 DVDD.n2979 DVSS 0.043914f
C3507 DVDD.n2980 DVSS 0.052845f
C3508 DVDD.n2981 DVSS 0.052845f
C3509 DVDD.n2982 DVSS 0.052845f
C3510 DVDD.n2983 DVSS 0.042611f
C3511 DVDD.n2984 DVSS 0.052845f
C3512 DVDD.n2985 DVSS 0.052845f
C3513 DVDD.n2986 DVSS 0.052845f
C3514 DVDD.n2987 DVSS 0.052845f
C3515 DVDD.n2988 DVSS 0.052845f
C3516 DVDD.n2989 DVSS 0.052845f
C3517 DVDD.n2990 DVSS 0.052845f
C3518 DVDD.n2991 DVSS 0.052845f
C3519 DVDD.n2992 DVSS 0.052845f
C3520 DVDD.n2993 DVSS 0.052845f
C3521 DVDD.n2994 DVSS 0.052845f
C3522 DVDD.n2995 DVSS 0.052845f
C3523 DVDD.n2996 DVSS 0.052845f
C3524 DVDD.n2997 DVSS 0.052845f
C3525 DVDD.n2998 DVSS 0.052845f
C3526 DVDD.n2999 DVSS 0.052845f
C3527 DVDD.n3000 DVSS 0.052845f
C3528 DVDD.n3001 DVSS 0.052845f
C3529 DVDD.n3002 DVSS 0.052845f
C3530 DVDD.n3003 DVSS 0.052845f
C3531 DVDD.n3004 DVSS 0.052845f
C3532 DVDD.n3005 DVSS 0.052845f
C3533 DVDD.n3006 DVSS 0.052845f
C3534 DVDD.n3007 DVSS 0.052845f
C3535 DVDD.n3008 DVSS 0.052845f
C3536 DVDD.n3009 DVSS 0.052845f
C3537 DVDD.n3010 DVSS 0.052845f
C3538 DVDD.n3011 DVSS 0.052845f
C3539 DVDD.n3012 DVSS 0.052845f
C3540 DVDD.n3013 DVSS 0.052845f
C3541 DVDD.n3014 DVSS 0.052845f
C3542 DVDD.n3015 DVSS 0.052845f
C3543 DVDD.n3016 DVSS 0.052845f
C3544 DVDD.n3017 DVSS 0.052845f
C3545 DVDD.n3018 DVSS 0.052845f
C3546 DVDD.n3019 DVSS 0.052845f
C3547 DVDD.n3020 DVSS 0.033866f
C3548 DVDD.n3021 DVSS 0.033866f
C3549 DVDD.n3022 DVSS 0.052845f
C3550 DVDD.n3023 DVSS 0.052845f
C3551 DVDD.n3024 DVSS 0.052845f
C3552 DVDD.n3025 DVSS 0.052845f
C3553 DVDD.n3026 DVSS 0.052845f
C3554 DVDD.n3027 DVSS 0.050798f
C3555 DVDD.n3028 DVSS 0.003076f
C3556 DVDD.n3029 DVSS 0.003076f
C3557 DVDD.n3030 DVSS 0.003076f
C3558 DVDD.n3031 DVSS 0.003076f
C3559 DVDD.n3032 DVSS 0.003076f
C3560 DVDD.n3033 DVSS 0.003076f
C3561 DVDD.n3034 DVSS 0.003076f
C3562 DVDD.n3035 DVSS 0.003076f
C3563 DVDD.n3036 DVSS 0.003076f
C3564 DVDD.n3037 DVSS 0.026423f
C3565 DVDD.n3038 DVSS 0.003076f
C3566 DVDD.n3039 DVSS 0.003076f
C3567 DVDD.n3040 DVSS 0.026423f
C3568 DVDD.n3041 DVSS 0.085321f
C3569 DVDD.n3042 DVSS 0.085321f
C3570 DVDD.n3043 DVSS 0.003076f
C3571 DVDD.n3044 DVSS 0.023631f
C3572 DVDD.n3045 DVSS 0.023073f
C3573 DVDD.n3046 DVSS 0.052845f
C3574 DVDD.n3047 DVSS 0.053362f
C3575 DVDD.n3048 DVSS 0.152989f
C3576 DVDD.n3049 DVSS 0.052845f
C3577 DVDD.n3050 DVSS 0.052845f
C3578 DVDD.n3051 DVSS 0.023073f
C3579 DVDD.n3052 DVSS 0.026423f
C3580 DVDD.n3053 DVSS 0.003076f
C3581 DVDD.n3054 DVSS 0.003076f
C3582 DVDD.n3055 DVSS 0.023073f
C3583 DVDD.n3056 DVSS 0.026423f
C3584 DVDD.n3057 DVSS 0.003076f
C3585 DVDD.n3058 DVSS 0.026423f
C3586 DVDD.n3059 DVSS 0.003076f
C3587 DVDD.n3060 DVSS 0.003076f
C3588 DVDD.n3061 DVSS 0.025492f
C3589 DVDD.n3062 DVSS 0.024004f
C3590 DVDD.n3063 DVSS 0.003076f
C3591 DVDD.n3064 DVSS 0.062707f
C3592 DVDD.n3065 DVSS 0.026423f
C3593 DVDD.n3066 DVSS 0.006004f
C3594 DVDD.n3067 DVSS 0.026423f
C3595 DVDD.n3068 DVSS 0.006004f
C3596 DVDD.n3069 DVSS 0.003076f
C3597 DVDD.n3070 DVSS 0.024004f
C3598 DVDD.n3071 DVSS 0.025492f
C3599 DVDD.n3072 DVSS 0.003076f
C3600 DVDD.n3073 DVSS 0.003076f
C3601 DVDD.n3074 DVSS 0.026423f
C3602 DVDD.n3075 DVSS 0.023073f
C3603 DVDD.n3076 DVSS 0.026423f
C3604 DVDD.n3077 DVSS 0.003076f
C3605 DVDD.n3078 DVSS 0.003076f
C3606 DVDD.n3079 DVSS 0.023073f
C3607 DVDD.n3080 DVSS 0.023073f
C3608 DVDD.n3081 DVSS 0.003076f
C3609 DVDD.n3082 DVSS 0.026423f
C3610 DVDD.n3083 DVSS 0.040378f
C3611 DVDD.n3084 DVSS 0.052845f
C3612 DVDD.n3085 DVSS 0.052845f
C3613 DVDD.n3086 DVSS 0.052845f
C3614 DVDD.n3087 DVSS 0.024004f
C3615 DVDD.n3088 DVSS 0.006004f
C3616 DVDD.n3089 DVSS 0.023073f
C3617 DVDD.n3090 DVSS 0.062707f
C3618 DVDD.n3091 DVSS 0.052845f
C3619 DVDD.n3092 DVSS 0.08485f
C3620 DVDD.n3093 DVSS 0.08485f
C3621 DVDD.n3094 DVSS 0.052845f
C3622 DVDD.n3095 DVSS 0.052845f
C3623 DVDD.n3096 DVSS 0.026423f
C3624 DVDD.n3097 DVSS 0.025492f
C3625 DVDD.n3098 DVSS 0.003076f
C3626 DVDD.n3099 DVSS 0.023073f
C3627 DVDD.n3100 DVSS 0.026423f
C3628 DVDD.n3101 DVSS 0.052845f
C3629 DVDD.n3102 DVSS 0.052845f
C3630 DVDD.n3103 DVSS 0.023073f
C3631 DVDD.n3104 DVSS 0.040378f
C3632 DVDD.n3105 DVSS 0.052845f
C3633 DVDD.n3106 DVSS 0.023073f
C3634 DVDD.n3107 DVSS 0.026423f
C3635 DVDD.n3108 DVSS 0.003076f
C3636 DVDD.n3109 DVSS 0.003076f
C3637 DVDD.n3110 DVSS 0.003076f
C3638 DVDD.n3111 DVSS 0.024004f
C3639 DVDD.n3112 DVSS 0.023073f
C3640 DVDD.n3113 DVSS 0.052845f
C3641 DVDD.n3114 DVSS 0.08485f
C3642 DVDD.n3115 DVSS 0.08485f
C3643 DVDD.n3116 DVSS 0.062707f
C3644 DVDD.n3117 DVSS 0.026423f
C3645 DVDD.n3118 DVSS 0.006004f
C3646 DVDD.n3119 DVSS 0.003076f
C3647 DVDD.n3120 DVSS 0.003076f
C3648 DVDD.n3121 DVSS 0.025492f
C3649 DVDD.n3122 DVSS 0.023073f
C3650 DVDD.n3123 DVSS 0.052845f
C3651 DVDD.n3124 DVSS 0.052845f
C3652 DVDD.n3125 DVSS 0.023073f
C3653 DVDD.n3126 DVSS 0.026423f
C3654 DVDD.n3127 DVSS 0.003076f
C3655 DVDD.n3128 DVSS 0.003076f
C3656 DVDD.n3129 DVSS 0.008245f
C3657 DVDD.n3130 DVSS 0.023073f
C3658 DVDD.n3131 DVSS 0.003076f
C3659 DVDD.n3132 DVSS 0.008245f
C3660 DVDD.n3133 DVSS 0.026423f
C3661 DVDD.n3134 DVSS 0.023073f
C3662 DVDD.n3135 DVSS 0.052845f
C3663 DVDD.n3136 DVSS 0.052845f
C3664 DVDD.n3137 DVSS 0.087827f
C3665 DVDD.n3138 DVSS 0.052845f
C3666 DVDD.n3139 DVSS 0.023631f
C3667 DVDD.n3140 DVSS 0.008245f
C3668 DVDD.n3141 DVSS 0.003151f
C3669 DVDD.n3142 DVSS 0.007046f
C3670 DVDD.n3143 DVSS 0.007046f
C3671 DVDD.n3144 DVSS 0.007046f
C3672 DVDD.n3145 DVSS 0.003523f
C3673 DVDD.n3146 DVSS 0.003076f
C3674 DVDD.n3147 DVSS 0.008245f
C3675 DVDD.n3148 DVSS 0.023073f
C3676 DVDD.n3149 DVSS 0.003076f
C3677 DVDD.n3150 DVSS 0.026423f
C3678 DVDD.n3151 DVSS 0.03889f
C3679 DVDD.n3152 DVSS 0.052845f
C3680 DVDD.n3153 DVSS 0.065321f
C3681 DVDD.n3154 DVSS 0.064737f
C3682 DVDD.n3155 DVSS 0.040378f
C3683 DVDD.n3156 DVSS 0.040378f
C3684 DVDD.n3157 DVSS 0.005185f
C3685 DVDD.n3158 DVSS 0.005384f
C3686 DVDD.n3159 DVSS 0.031765f
C3687 DVDD.n3160 DVSS 0.040378f
C3688 DVDD.n3161 DVSS 0.03889f
C3689 DVDD.n3162 DVSS 0.070897f
C3690 DVDD.n3163 DVSS 0.031917f
C3691 DVDD.n3164 DVSS 0.03889f
C3692 DVDD.n3165 DVSS 0.040378f
C3693 DVDD.n3166 DVSS 0.03889f
C3694 DVDD.n3167 DVSS 0.031917f
C3695 DVDD.n3168 DVSS 0.023073f
C3696 DVDD.n3169 DVSS 0.447695f
C3697 DVDD.n3170 DVSS 0.005185f
C3698 DVDD.n3171 DVSS 0.005384f
C3699 DVDD.n3172 DVSS 0.03889f
C3700 DVDD.n3173 DVSS 0.040378f
C3701 DVDD.n3174 DVSS 0.066256f
C3702 DVDD.n3175 DVSS 0.040378f
C3703 DVDD.n3176 DVSS 0.052845f
C3704 DVDD.n3177 DVSS 0.023073f
C3705 DVDD.n3178 DVSS 0.003076f
C3706 DVDD.n3179 DVSS 0.026423f
C3707 DVDD.n3180 DVSS 0.052845f
C3708 DVDD.n3181 DVSS 0.052416f
C3709 DVDD.n3182 DVSS 0.023073f
C3710 DVDD.n3183 DVSS 0.025492f
C3711 DVDD.n3184 DVSS 0.025852f
C3712 DVDD.n3185 DVSS 0.025852f
C3713 DVDD.n3186 DVSS 0.003076f
C3714 DVDD.n3187 DVSS 0.003076f
C3715 DVDD.n3188 DVSS 0.024004f
C3716 DVDD.n3189 DVSS 0.023073f
C3717 DVDD.n3190 DVSS 0.052845f
C3718 DVDD.n3191 DVSS 0.050332f
C3719 DVDD.n3192 DVSS 0.150127f
C3720 DVDD.n3193 DVSS 0.052845f
C3721 DVDD.n3194 DVSS 0.052845f
C3722 DVDD.n3195 DVSS 0.023073f
C3723 DVDD.n3196 DVSS 0.023073f
C3724 DVDD.n3197 DVSS 0.026423f
C3725 DVDD.n3198 DVSS 0.003076f
C3726 DVDD.n3199 DVSS 0.003076f
C3727 DVDD.n3200 DVSS 0.003076f
C3728 DVDD.n3201 DVSS 0.026423f
C3729 DVDD.n3202 DVSS 0.052845f
C3730 DVDD.n3203 DVSS 0.052845f
C3731 DVDD.n3204 DVSS 0.052845f
C3732 DVDD.n3205 DVSS 0.087827f
C3733 DVDD.n3206 DVSS 0.025864f
C3734 DVDD.n3207 DVSS 0.087827f
C3735 DVDD.n3208 DVSS 0.087827f
C3736 DVDD.n3209 DVSS 0.052845f
C3737 DVDD.n3210 DVSS 0.052845f
C3738 DVDD.n3211 DVSS 0.023631f
C3739 DVDD.n3212 DVSS 0.023073f
C3740 DVDD.n3213 DVSS 0.003076f
C3741 DVDD.n3214 DVSS 0.003076f
C3742 DVDD.n3215 DVSS 0.026423f
C3743 DVDD.n3216 DVSS 0.052845f
C3744 DVDD.n3217 DVSS 0.03889f
C3745 DVDD.n3218 DVSS 0.052845f
C3746 DVDD.n3219 DVSS 0.052845f
C3747 DVDD.n3220 DVSS 0.023073f
C3748 DVDD.n3221 DVSS 0.026423f
C3749 DVDD.n3222 DVSS 0.003076f
C3750 DVDD.n3223 DVSS 0.003076f
C3751 DVDD.n3224 DVSS 0.026423f
C3752 DVDD.n3225 DVSS 0.023073f
C3753 DVDD.n3226 DVSS 0.052845f
C3754 DVDD.n3227 DVSS 0.087827f
C3755 DVDD.n3228 DVSS 0.064196f
C3756 DVDD.n3229 DVSS 0.064196f
C3757 DVDD.n3230 DVSS 0.025864f
C3758 DVDD.n3231 DVSS 0.003076f
C3759 DVDD.n3232 DVSS 0.023631f
C3760 DVDD.n3233 DVSS 0.023073f
C3761 DVDD.n3234 DVSS 0.052845f
C3762 DVDD.n3235 DVSS 0.052845f
C3763 DVDD.n3236 DVSS 0.023073f
C3764 DVDD.n3237 DVSS 0.026423f
C3765 DVDD.n3238 DVSS 0.003076f
C3766 DVDD.n3239 DVSS 0.003076f
C3767 DVDD.n3240 DVSS 0.026423f
C3768 DVDD.n3241 DVSS 0.023073f
C3769 DVDD.n3242 DVSS 0.03889f
C3770 DVDD.n3243 DVSS 0.040378f
C3771 DVDD.n3244 DVSS 0.040378f
C3772 DVDD.n3245 DVSS 0.052845f
C3773 DVDD.n3246 DVSS 0.023073f
C3774 DVDD.n3247 DVSS 0.003076f
C3775 DVDD.n3248 DVSS 0.003076f
C3776 DVDD.n3249 DVSS 0.026423f
C3777 DVDD.n3250 DVSS 0.052845f
C3778 DVDD.n3251 DVSS 0.052845f
C3779 DVDD.n3252 DVSS 0.052845f
C3780 DVDD.n3253 DVSS 0.087827f
C3781 DVDD.n3254 DVSS 0.025864f
C3782 DVDD.n3255 DVSS 5.09e-19
C3783 DVDD.n3256 DVSS 0.002059f
C3784 DVDD.n3257 DVSS 4.9e-19
C3785 DVDD.n3258 DVSS 0.001161f
C3786 DVDD.n3259 DVSS 4.9e-19
C3787 DVDD.n3260 DVSS 0.001161f
C3788 DVDD.n3261 DVSS 0.001161f
C3789 DVDD.n3262 DVSS 9.8e-19
C3790 DVDD.n3263 DVSS 9.8e-19
C3791 DVDD.n3264 DVSS 0.001161f
C3792 DVDD.n3265 DVSS 0.001161f
C3793 DVDD.n3266 DVSS 9.8e-19
C3794 DVDD.n3267 DVSS 9.8e-19
C3795 DVDD.n3268 DVSS 0.001161f
C3796 DVDD.n3269 DVSS 0.001161f
C3797 DVDD.n3270 DVSS 9.8e-19
C3798 DVDD.n3271 DVSS 9.8e-19
C3799 DVDD.n3272 DVSS 0.001161f
C3800 DVDD.n3273 DVSS 0.001161f
C3801 DVDD.n3274 DVSS 9.8e-19
C3802 DVDD.n3275 DVSS 9.8e-19
C3803 DVDD.n3276 DVSS 0.001161f
C3804 DVDD.n3277 DVSS 0.001161f
C3805 DVDD.n3278 DVSS 9.8e-19
C3806 DVDD.n3279 DVSS 9.8e-19
C3807 DVDD.n3280 DVSS 0.001161f
C3808 DVDD.n3281 DVSS 0.001161f
C3809 DVDD.n3282 DVSS 9.8e-19
C3810 DVDD.n3283 DVSS 9.8e-19
C3811 DVDD.n3284 DVSS 0.001161f
C3812 DVDD.n3285 DVSS 0.001161f
C3813 DVDD.n3286 DVSS 9.8e-19
C3814 DVDD.n3287 DVSS 9.8e-19
C3815 DVDD.n3288 DVSS 0.001161f
C3816 DVDD.n3289 DVSS 0.001161f
C3817 DVDD.n3290 DVSS 9.8e-19
C3818 DVDD.n3291 DVSS 9.8e-19
C3819 DVDD.n3292 DVSS 0.001161f
C3820 DVDD.n3293 DVSS 0.001161f
C3821 DVDD.n3294 DVSS 9.8e-19
C3822 DVDD.n3295 DVSS 9.8e-19
C3823 DVDD.n3296 DVSS 0.001161f
C3824 DVDD.n3297 DVSS 0.001161f
C3825 DVDD.n3298 DVSS 9.8e-19
C3826 DVDD.n3299 DVSS 9.43e-19
C3827 DVDD.n3300 DVSS 0.001161f
C3828 DVDD.n3301 DVSS 0.001161f
C3829 DVDD.n3302 DVSS 5.09e-19
C3830 DVDD.n3303 DVSS 4.9e-19
C3831 DVDD.n3304 DVSS 0.001161f
C3832 DVDD.n3305 DVSS 5.09e-19
C3833 DVDD.n3306 DVSS 9.8e-19
C3834 DVDD.n3307 DVSS 5.09e-19
C3835 DVDD.n3308 DVSS 0.001161f
C3836 DVDD.n3309 DVSS 0.001161f
C3837 DVDD.n3310 DVSS 5.09e-19
C3838 DVDD.n3311 DVSS 4.9e-19
C3839 DVDD.n3312 DVSS 9.43e-19
C3840 DVDD.n3313 DVSS 0.001161f
C3841 DVDD.n3314 DVSS 0.001161f
C3842 DVDD.n3315 DVSS 9.8e-19
C3843 DVDD.n3316 DVSS 9.8e-19
C3844 DVDD.n3317 DVSS 0.001161f
C3845 DVDD.n3318 DVSS 0.001161f
C3846 DVDD.n3319 DVSS 9.8e-19
C3847 DVDD.n3320 DVSS 9.8e-19
C3848 DVDD.n3321 DVSS 0.001161f
C3849 DVDD.n3322 DVSS 0.001161f
C3850 DVDD.n3323 DVSS 9.8e-19
C3851 DVDD.n3324 DVSS 9.8e-19
C3852 DVDD.n3325 DVSS 0.001161f
C3853 DVDD.n3326 DVSS 0.001161f
C3854 DVDD.n3327 DVSS 9.8e-19
C3855 DVDD.n3328 DVSS 9.8e-19
C3856 DVDD.n3329 DVSS 0.001161f
C3857 DVDD.n3330 DVSS 0.001161f
C3858 DVDD.n3331 DVSS 9.8e-19
C3859 DVDD.n3332 DVSS 9.8e-19
C3860 DVDD.n3333 DVSS 0.001161f
C3861 DVDD.n3334 DVSS 0.001161f
C3862 DVDD.n3335 DVSS 9.8e-19
C3863 DVDD.n3336 DVSS 9.8e-19
C3864 DVDD.n3337 DVSS 0.001161f
C3865 DVDD.n3338 DVSS 0.001161f
C3866 DVDD.n3339 DVSS 9.8e-19
C3867 DVDD.n3340 DVSS 9.8e-19
C3868 DVDD.n3341 DVSS 0.001161f
C3869 DVDD.n3342 DVSS 0.001161f
C3870 DVDD.n3343 DVSS 9.8e-19
C3871 DVDD.n3344 DVSS 9.8e-19
C3872 DVDD.n3345 DVSS 0.001161f
C3873 DVDD.n3346 DVSS 0.001161f
C3874 DVDD.n3347 DVSS 9.8e-19
C3875 DVDD.n3348 DVSS 9.8e-19
C3876 DVDD.n3349 DVSS 0.001161f
C3877 DVDD.n3350 DVSS 0.001161f
C3878 DVDD.n3351 DVSS 9.8e-19
C3879 DVDD.n3352 DVSS 0.001161f
C3880 DVDD.n3353 DVSS 0.001161f
C3881 DVDD.n3354 DVSS 9.24e-19
C3882 DVDD.n3355 DVSS 4.9e-19
C3883 DVDD.n3356 DVSS 0.003076f
C3884 DVDD.n3357 DVSS 0.064196f
C3885 DVDD.n3358 DVSS 0.026423f
C3886 DVDD.n3359 DVSS 0.087827f
C3887 DVDD.n3360 DVSS 0.052845f
C3888 DVDD.n3361 DVSS 0.052845f
C3889 DVDD.n3362 DVSS 0.052845f
C3890 DVDD.n3363 DVSS 0.023073f
C3891 DVDD.n3364 DVSS 0.003076f
C3892 DVDD.n3365 DVSS 0.026423f
C3893 DVDD.n3366 DVSS 0.023073f
C3894 DVDD.n3367 DVSS 0.003076f
C3895 DVDD.n3368 DVSS 0.026423f
C3896 DVDD.n3369 DVSS 0.052845f
C3897 DVDD.n3370 DVSS 0.052416f
C3898 DVDD.n3371 DVSS 0.023073f
C3899 DVDD.n3372 DVSS 0.025492f
C3900 DVDD.n3373 DVSS 0.01233f
C3901 DVDD.n3374 DVSS 0.01233f
C3902 DVDD.n3375 DVSS 0.003052f
C3903 DVDD.n3376 DVSS 4.9e-19
C3904 DVDD.n3377 DVSS 5.09e-19
C3905 DVDD.n3378 DVSS 9.8e-19
C3906 DVDD.n3380 DVSS 0.001161f
C3907 DVDD.n3381 DVSS 9.8e-19
C3908 DVDD.n3383 DVSS 0.001161f
C3909 DVDD.n3384 DVSS 9.8e-19
C3910 DVDD.n3386 DVSS 0.001161f
C3911 DVDD.n3387 DVSS 9.8e-19
C3912 DVDD.n3389 DVSS 0.001161f
C3913 DVDD.n3390 DVSS 9.8e-19
C3914 DVDD.n3392 DVSS 0.001161f
C3915 DVDD.n3393 DVSS 4.9e-19
C3916 DVDD.n3395 DVSS 5.09e-19
C3917 DVDD.n3396 DVSS 0.001161f
C3918 DVDD.n3397 DVSS 4.9e-19
C3919 DVDD.n3398 DVSS 5.09e-19
C3920 DVDD.n3399 DVSS 0.008178f
C3921 DVDD.n3400 DVSS 4.9e-19
C3922 DVDD.n3401 DVSS 0.004189f
C3923 DVDD.n3402 DVSS 5.09e-19
C3924 DVDD.n3403 DVSS 9.8e-19
C3925 DVDD.n3405 DVSS 0.001161f
C3926 DVDD.n3406 DVSS 0.001161f
C3927 DVDD.n3408 DVSS 0.001161f
C3928 DVDD.n3409 DVSS 9.8e-19
C3929 DVDD.n3411 DVSS 0.001161f
C3930 DVDD.n3412 DVSS 9.8e-19
C3931 DVDD.n3414 DVSS 0.001161f
C3932 DVDD.n3415 DVSS 9.8e-19
C3933 DVDD.n3417 DVSS 0.001161f
C3934 DVDD.n3418 DVSS 9.8e-19
C3935 DVDD.n3420 DVSS 0.001161f
C3936 DVDD.n3421 DVSS 4.9e-19
C3937 DVDD.n3423 DVSS 5.09e-19
C3938 DVDD.n3424 DVSS 0.001161f
C3939 DVDD.n3425 DVSS 0.003052f
C3940 DVDD.n3426 DVSS 0.01233f
C3941 DVDD.n3427 DVSS 0.01233f
C3942 DVDD.n3428 DVSS 0.003076f
C3943 DVDD.n3429 DVSS 0.050332f
C3944 DVDD.n3430 DVSS 0.023073f
C3945 DVDD.n3433 DVSS 0.014849f
C3946 DVDD.n3434 DVSS 0.008245f
C3947 DVDD.n3435 DVSS 0.004455f
C3948 DVDD.n3438 DVSS 0.010767f
C3949 DVDD.n3439 DVSS 0.008245f
C3950 DVDD.n3441 DVSS 0.010767f
C3951 DVDD.n3445 DVSS 0.011723f
C3952 DVDD.n3446 DVSS 0.008245f
C3953 DVDD.n3447 DVSS 0.008245f
C3954 DVDD.n3448 DVSS 0.024661f
C3955 DVDD.n3449 DVSS 0.024661f
C3956 DVDD.n3450 DVSS 0.024661f
C3957 DVDD.n3451 DVSS 0.024661f
C3958 DVDD.n3452 DVSS 0.024661f
C3959 DVDD.n3453 DVSS 0.024661f
C3960 DVDD.n3454 DVSS 0.024661f
C3961 DVDD.n3455 DVSS 0.024661f
C3962 DVDD.n3456 DVSS 0.024661f
C3963 DVDD.n3457 DVSS 0.024661f
C3964 DVDD.n3458 DVSS 0.024661f
C3965 DVDD.n3459 DVSS 0.024661f
C3966 DVDD.n3460 DVSS 0.024661f
C3967 DVDD.n3461 DVSS 0.024661f
C3968 DVDD.n3462 DVSS 0.024661f
C3969 DVDD.n3463 DVSS 0.024661f
C3970 DVDD.n3464 DVSS 0.024661f
C3971 DVDD.n3465 DVSS 0.024661f
C3972 DVDD.n3466 DVSS 0.024661f
C3973 DVDD.n3467 DVSS 0.024661f
C3974 DVDD.n3468 DVSS 0.014849f
C3975 DVDD.n3469 DVSS 0.024661f
C3976 DVDD.n3470 DVSS 0.024661f
C3977 DVDD.n3471 DVSS 0.024661f
C3978 DVDD.n3472 DVSS 0.024661f
C3979 DVDD.n3473 DVSS 0.024661f
C3980 DVDD.n3474 DVSS 0.024661f
C3981 DVDD.n3475 DVSS 0.024661f
C3982 DVDD.n3476 DVSS 0.024661f
C3983 DVDD.n3477 DVSS 0.024661f
C3984 DVDD.n3478 DVSS 0.024661f
C3985 DVDD.n3479 DVSS 0.024661f
C3986 DVDD.n3480 DVSS 0.024661f
C3987 DVDD.n3481 DVSS 0.385637f
C3988 DVDD.n3482 DVSS 0.024661f
C3989 DVDD.n3483 DVSS 0.010767f
C3990 DVDD.n3484 DVSS 0.003076f
C3991 DVDD.n3485 DVSS 0.050332f
C3992 DVDD.n3486 DVSS 0.024004f
C3993 DVDD.n3487 DVSS 0.150127f
C3994 DVDD.n3488 DVSS 0.052845f
C3995 DVDD.n3489 DVSS 0.052845f
C3996 DVDD.n3490 DVSS 0.025492f
C3997 DVDD.n3491 DVSS 0.023073f
C3998 DVDD.n3492 DVSS 0.003076f
C3999 DVDD.n3493 DVSS 0.023073f
C4000 DVDD.n3494 DVSS 0.026423f
C4001 DVDD.n3495 DVSS 0.003076f
C4002 DVDD.n3496 DVSS 0.003076f
C4003 DVDD.n3497 DVSS 0.026423f
C4004 DVDD.n3498 DVSS 0.023073f
C4005 DVDD.n3499 DVSS 0.052845f
C4006 DVDD.n3500 DVSS 0.052845f
C4007 DVDD.n3501 DVSS 0.023073f
C4008 DVDD.n3502 DVSS 0.052416f
C4009 DVDD.n3503 DVSS 0.025852f
C4010 DVDD.n3504 DVSS 0.025852f
C4011 DVDD.n3505 DVSS 0.00226f
C4012 DVDD.n3506 DVSS 0.001538f
C4013 DVDD.n3507 DVSS 0.003076f
C4014 DVDD.n3508 DVSS 0.003388f
C4015 DVDD.n3509 DVSS 0.002693f
C4016 DVDD.n3510 DVSS 0.054232f
C4017 DVDD.n3511 DVSS 0.001538f
C4018 DVDD.n3512 DVSS 0.003076f
C4019 DVDD.n3513 DVSS 0.003076f
C4020 DVDD.n3514 DVSS 0.003076f
C4021 DVDD.n3515 DVSS 0.001538f
C4022 DVDD.n3516 DVSS 0.001662f
C4023 DVDD.n3517 DVSS 0.001464f
C4024 DVDD.n3518 DVSS 0.00134f
C4025 DVDD.n3519 DVSS 0.054841f
C4026 DVDD.n3520 DVSS 0.00134f
C4027 DVDD.n3522 DVSS 0.00134f
C4028 DVDD.n3523 DVSS 0.028092f
C4029 DVDD.n3524 DVSS 0.002679f
C4030 DVDD.t160 DVSS 0.198479f
C4031 DVDD.n3525 DVSS 0.031051f
C4032 DVDD.n3526 DVSS 0.054842f
C4033 DVDD.n3527 DVSS 0.054232f
C4034 DVDD.n3528 DVSS 0.002693f
C4035 DVDD.n3529 DVSS 0.002679f
C4036 DVDD.n3530 DVSS 0.00493f
C4037 DVDD.n3531 DVSS 0.002679f
C4038 DVDD.n3532 DVSS 0.00493f
C4039 DVDD.n3533 DVSS 0.002679f
C4040 DVDD.n3534 DVSS 0.00493f
C4041 DVDD.n3535 DVSS 0.002679f
C4042 DVDD.n3536 DVSS 0.00493f
C4043 DVDD.n3537 DVSS 0.002679f
C4044 DVDD.n3538 DVSS -0.118241f
C4045 DVDD.n3539 DVSS 0.002679f
C4046 DVDD.n3540 DVSS 0.00493f
C4047 DVDD.n3541 DVSS 0.002679f
C4048 DVDD.n3542 DVSS 0.00493f
C4049 DVDD.n3543 DVSS 0.002679f
C4050 DVDD.n3544 DVSS 0.00493f
C4051 DVDD.n3545 DVSS 0.002679f
C4052 DVDD.n3546 DVSS 0.00493f
C4053 DVDD.n3547 DVSS 0.002679f
C4054 DVDD.n3548 DVSS 0.002693f
C4055 DVDD.n3549 DVSS 0.057866f
C4056 DVDD.n3550 DVSS 0.012517f
C4057 DVDD.n3551 DVSS 0.001538f
C4058 DVDD.n3552 DVSS 0.010767f
C4059 DVDD.n3553 DVSS 0.018322f
C4060 DVDD.n3554 DVSS 0.001538f
C4061 DVDD.n3555 DVSS 0.003076f
C4062 DVDD.n3556 DVSS 0.003076f
C4063 DVDD.n3557 DVSS 0.003076f
C4064 DVDD.n3558 DVSS 0.024661f
C4065 DVDD.n3559 DVSS 0.024661f
C4066 DVDD.n3560 DVSS 0.024661f
C4067 DVDD.n3561 DVSS 0.024661f
C4068 DVDD.n3562 DVSS 0.024661f
C4069 DVDD.n3563 DVSS 0.024661f
C4070 DVDD.n3564 DVSS 0.024661f
C4071 DVDD.n3565 DVSS 0.024661f
C4072 DVDD.n3566 DVSS 0.024661f
C4073 DVDD.n3567 DVSS 0.024661f
C4074 DVDD.n3568 DVSS 0.024661f
C4075 DVDD.n3569 DVSS 0.024661f
C4076 DVDD.n3570 DVSS 0.024661f
C4077 DVDD.n3571 DVSS 0.024661f
C4078 DVDD.n3572 DVSS 0.024661f
C4079 DVDD.n3573 DVSS 0.024661f
C4080 DVDD.n3574 DVSS 0.024661f
C4081 DVDD.n3575 DVSS 0.010767f
C4082 DVDD.n3576 DVSS 0.00134f
C4083 DVDD.n3577 DVSS 0.00134f
C4084 DVDD.n3578 DVSS 0.00134f
C4085 DVDD.n3579 DVSS 0.00134f
C4086 DVDD.n3580 DVSS 0.00134f
C4087 DVDD.n3581 DVSS 0.00134f
C4088 DVDD.n3582 DVSS 0.00134f
C4089 DVDD.n3583 DVSS 0.00134f
C4090 DVDD.n3584 DVSS 0.00134f
C4091 DVDD.n3585 DVSS 0.00134f
C4092 DVDD.n3586 DVSS 0.10316f
C4093 DVDD.n3587 DVSS 0.001538f
C4094 DVDD.n3588 DVSS 0.024661f
C4095 DVDD.n3589 DVSS 0.024661f
C4096 DVDD.n3590 DVSS 0.024661f
C4097 DVDD.n3591 DVSS 0.024661f
C4098 DVDD.n3592 DVSS 0.024661f
C4099 DVDD.n3593 DVSS 0.024661f
C4100 DVDD.n3594 DVSS 0.024661f
C4101 DVDD.n3595 DVSS 0.024661f
C4102 DVDD.n3596 DVSS 0.024661f
C4103 DVDD.n3597 DVSS 0.024661f
C4104 DVDD.n3598 DVSS 0.024661f
C4105 DVDD.n3599 DVSS 0.024661f
C4106 DVDD.n3600 DVSS 0.024661f
C4107 DVDD.n3601 DVSS 0.024661f
C4108 DVDD.n3602 DVSS 0.024661f
C4109 DVDD.n3603 DVSS 0.024661f
C4110 DVDD.n3604 DVSS 0.024661f
C4111 DVDD.n3605 DVSS 0.010767f
C4112 DVDD.n3606 DVSS 0.008245f
C4113 DVDD.n3607 DVSS 0.008245f
C4114 DVDD.n3608 DVSS 0.008245f
C4115 DVDD.n3609 DVSS 0.008245f
C4116 DVDD.n3610 DVSS 0.008245f
C4117 DVDD.n3611 DVSS 0.068419f
C4118 DVDD.n3612 DVSS 0.008245f
C4119 DVDD.n3613 DVSS 0.008245f
C4120 DVDD.n3614 DVSS 0.008245f
C4121 DVDD.n3615 DVSS 0.008245f
C4122 DVDD.n3622 DVSS 0.011375f
C4123 DVDD.n3627 DVSS 0.01233f
C4124 DVDD.n3628 DVSS 0.024661f
C4125 DVDD.n3629 DVSS 0.024661f
C4126 DVDD.n3630 DVSS 0.024661f
C4127 DVDD.n3631 DVSS 0.024661f
C4128 DVDD.n3632 DVSS 0.024661f
C4129 DVDD.n3633 DVSS 0.024661f
C4130 DVDD.n3634 DVSS 0.024661f
C4131 DVDD.n3635 DVSS 0.024661f
C4132 DVDD.n3636 DVSS 0.024661f
C4133 DVDD.n3637 DVSS 0.024661f
C4134 DVDD.n3638 DVSS 0.024661f
C4135 DVDD.n3639 DVSS 0.024661f
C4136 DVDD.n3640 DVSS 0.024661f
C4137 DVDD.n3641 DVSS 0.024661f
C4138 DVDD.n3642 DVSS 0.024661f
C4139 DVDD.n3643 DVSS 0.024661f
C4140 DVDD.n3644 DVSS 0.01233f
C4141 DVDD.n3645 DVSS 0.024661f
C4142 DVDD.n3646 DVSS 0.024661f
C4143 DVDD.n3647 DVSS 0.024661f
C4144 DVDD.n3648 DVSS 0.024661f
C4145 DVDD.n3649 DVSS 0.00134f
C4146 DVDD.n3650 DVSS 0.00134f
C4147 DVDD.n3651 DVSS 0.022707f
C4148 DVDD.n3652 DVSS 0.00134f
C4149 DVDD.n3653 DVSS 0.00134f
C4150 DVDD.n3654 DVSS 0.010767f
C4151 DVDD.n3655 DVSS 0.00134f
C4152 DVDD.n3656 DVSS 0.00134f
C4153 DVDD.n3657 DVSS 0.00134f
C4154 DVDD.n3658 DVSS 0.00134f
C4155 DVDD.n3659 DVSS 0.00134f
C4156 DVDD.n3660 DVSS 0.001538f
C4157 DVDD.n3661 DVSS 0.001476f
C4158 DVDD.n3662 DVSS 0.013397f
C4159 DVDD.n3663 DVSS 0.013397f
C4160 DVDD.n3664 DVSS 0.002679f
C4161 DVDD.n3665 DVSS 0.013397f
C4162 DVDD.n3666 DVSS 0.051813f
C4163 DVDD.n3667 DVSS 0.054232f
C4164 DVDD.n3668 DVSS 0.063552f
C4165 DVDD.n3669 DVSS 0.00134f
C4166 DVDD.n3671 DVSS 0.00134f
C4167 DVDD.n3673 DVSS 0.00134f
C4168 DVDD.t159 DVSS 0.198479f
C4169 DVDD.n3674 DVSS 0.002679f
C4170 DVDD.n3675 DVSS 0.00134f
C4171 DVDD.n3676 DVSS 0.063552f
C4172 DVDD.n3677 DVSS 0.031051f
C4173 DVDD.n3678 DVSS 0.063551f
C4174 DVDD.n3679 DVSS 0.031051f
C4175 DVDD.n3680 DVSS 0.002679f
C4176 DVDD.t156 DVSS 0.198479f
C4177 DVDD.n3681 DVSS 0.031051f
C4178 DVDD.n3682 DVSS 0.011228f
C4179 DVDD.n3683 DVSS 0.002679f
C4180 DVDD.n3686 DVSS 0.003698f
C4181 DVDD.n3687 DVSS 0.00493f
C4182 DVDD.n3688 DVSS 0.002679f
C4183 DVDD.n3689 DVSS 0.00493f
C4184 DVDD.n3690 DVSS 0.002679f
C4185 DVDD.n3691 DVSS 0.00493f
C4186 DVDD.n3692 DVSS 0.002679f
C4187 DVDD.n3693 DVSS 0.00493f
C4188 DVDD.n3694 DVSS 0.002679f
C4189 DVDD.n3695 DVSS 0.00493f
C4190 DVDD.n3696 DVSS 0.002679f
C4191 DVDD.n3697 DVSS 0.057866f
C4192 DVDD.n3698 DVSS 0.012517f
C4193 DVDD.n3699 DVSS 0.342976f
C4194 DVDD.n3700 DVSS 0.010767f
C4195 DVDD.n3701 DVSS 0.024661f
C4196 DVDD.n3702 DVSS 0.080216f
C4197 DVDD.n3703 DVSS 0.024661f
C4198 DVDD.n3704 DVSS 0.588581f
C4199 DVDD.n3705 DVSS 0.024661f
C4200 DVDD.n3706 DVSS 0.024661f
C4201 DVDD.n3707 DVSS 0.024661f
C4202 DVDD.n3708 DVSS 0.024661f
C4203 DVDD.n3709 DVSS 0.024661f
C4204 DVDD.n3710 DVSS 0.024661f
C4205 DVDD.n3711 DVSS 0.024661f
C4206 DVDD.n3712 DVSS 0.024661f
C4207 DVDD.n3713 DVSS 0.024661f
C4208 DVDD.n3714 DVSS 0.024661f
C4209 DVDD.n3715 DVSS 0.024661f
C4210 DVDD.n3716 DVSS 0.024661f
C4211 DVDD.n3717 DVSS 0.024661f
C4212 DVDD.n3718 DVSS 0.024661f
C4213 DVDD.n3719 DVSS 0.024661f
C4214 DVDD.n3720 DVSS 0.024661f
C4215 DVDD.n3721 DVSS 0.024661f
C4216 DVDD.n3722 DVSS 0.024661f
C4217 DVDD.n3723 DVSS 0.024661f
C4218 DVDD.n3724 DVSS 0.024661f
C4219 DVDD.n3725 DVSS 0.024661f
C4220 DVDD.n3726 DVSS 0.024661f
C4221 DVDD.n3727 DVSS 0.024661f
C4222 DVDD.n3728 DVSS 0.024661f
C4223 DVDD.n3729 DVSS 0.024661f
C4224 DVDD.n3730 DVSS 0.024661f
C4225 DVDD.n3731 DVSS 0.024661f
C4226 DVDD.n3732 DVSS 0.024661f
C4227 DVDD.n3733 DVSS 0.024661f
C4228 DVDD.n3734 DVSS 0.024661f
C4229 DVDD.n3735 DVSS 0.024661f
C4230 DVDD.n3736 DVSS 0.024661f
C4231 DVDD.n3737 DVSS 0.024661f
C4232 DVDD.n3738 DVSS 0.024661f
C4233 DVDD.n3739 DVSS 0.024661f
C4234 DVDD.n3740 DVSS 0.024661f
C4235 DVDD.n3741 DVSS 0.024661f
C4236 DVDD.n3742 DVSS 0.385657f
C4237 DVDD.n3743 DVSS 0.024661f
C4238 DVDD.n3744 DVSS 0.019885f
C4239 DVDD.n3745 DVSS 0.01233f
C4240 DVDD.n3746 DVSS 0.001538f
C4241 DVDD.n3747 DVSS 0.003076f
C4242 DVDD.n3748 DVSS 0.003076f
C4243 DVDD.n3749 DVSS 0.003076f
C4244 DVDD.n3750 DVSS 0.003076f
C4245 DVDD.n3751 DVSS 0.003076f
C4246 DVDD.n3752 DVSS 0.003076f
C4247 DVDD.n3753 DVSS 0.003076f
C4248 DVDD.n3754 DVSS 0.003076f
C4249 DVDD.n3755 DVSS 0.001538f
C4250 DVDD.n3756 DVSS 0.035774f
C4251 DVDD.n3757 DVSS 0.204625f
C4252 DVDD.t155 DVSS 0.617722f
C4253 DVDD.n3759 DVSS 0.200207f
C4254 DVDD.n3760 DVSS 0.025152f
C4255 DVDD.n3761 DVSS 0.016319f
C4256 DVDD.n3762 DVSS 0.004474f
C4257 DVDD.n3763 DVSS 0.002693f
C4258 DVDD.n3764 DVSS 0.00493f
C4259 DVDD.n3765 DVSS 0.00493f
C4260 DVDD.n3766 DVSS 0.002679f
C4261 DVDD.n3767 DVSS 0.002679f
C4262 DVDD.n3768 DVSS 0.002679f
C4263 DVDD.n3769 DVSS 0.00493f
C4264 DVDD.n3770 DVSS 0.00493f
C4265 DVDD.n3771 DVSS 0.00493f
C4266 DVDD.n3772 DVSS 0.002679f
C4267 DVDD.n3773 DVSS 0.002679f
C4268 DVDD.n3774 DVSS 0.002679f
C4269 DVDD.n3775 DVSS 0.00493f
C4270 DVDD.n3776 DVSS 0.00493f
C4271 DVDD.n3777 DVSS 0.00493f
C4272 DVDD.n3778 DVSS 0.002679f
C4273 DVDD.n3779 DVSS 0.002679f
C4274 DVDD.n3780 DVSS 0.002679f
C4275 DVDD.n3781 DVSS 0.00493f
C4276 DVDD.n3782 DVSS 0.00493f
C4277 DVDD.n3783 DVSS 0.00493f
C4278 DVDD.n3784 DVSS 0.002679f
C4279 DVDD.n3785 DVSS 0.002679f
C4280 DVDD.n3786 DVSS 0.002679f
C4281 DVDD.n3787 DVSS 0.00493f
C4282 DVDD.n3788 DVSS 0.00493f
C4283 DVDD.n3789 DVSS 0.00493f
C4284 DVDD.n3790 DVSS 0.002679f
C4285 DVDD.n3791 DVSS 0.002679f
C4286 DVDD.n3792 DVSS 0.002679f
C4287 DVDD.n3793 DVSS 0.00493f
C4288 DVDD.n3794 DVSS 0.002679f
C4289 DVDD.n3795 DVSS 0.00493f
C4290 DVDD.n3796 DVSS 0.002679f
C4291 DVDD.n3797 DVSS 0.00493f
C4292 DVDD.n3798 DVSS 0.002679f
C4293 DVDD.n3799 DVSS 0.00493f
C4294 DVDD.n3800 DVSS 0.003582f
C4295 DVDD.n3801 DVSS 0.00493f
C4296 DVDD.n3802 DVSS 0.002679f
C4297 DVDD.n3803 DVSS 0.002679f
C4298 DVDD.n3804 DVSS 0.002679f
C4299 DVDD.n3805 DVSS 0.00493f
C4300 DVDD.n3806 DVSS 0.00493f
C4301 DVDD.n3807 DVSS 0.00493f
C4302 DVDD.n3808 DVSS 0.002679f
C4303 DVDD.n3809 DVSS 0.002679f
C4304 DVDD.n3810 DVSS 0.002679f
C4305 DVDD.n3811 DVSS 0.00493f
C4306 DVDD.n3812 DVSS 0.00493f
C4307 DVDD.n3813 DVSS 0.00493f
C4308 DVDD.n3814 DVSS 0.002679f
C4309 DVDD.n3815 DVSS 0.002679f
C4310 DVDD.n3816 DVSS 0.002679f
C4311 DVDD.n3817 DVSS 0.00493f
C4312 DVDD.n3818 DVSS 0.00493f
C4313 DVDD.n3819 DVSS 0.00493f
C4314 DVDD.n3820 DVSS 0.002679f
C4315 DVDD.n3821 DVSS 0.002679f
C4316 DVDD.n3822 DVSS 0.002679f
C4317 DVDD.n3823 DVSS 0.00493f
C4318 DVDD.n3824 DVSS 0.00493f
C4319 DVDD.n3825 DVSS 0.00493f
C4320 DVDD.n3826 DVSS 0.002679f
C4321 DVDD.n3827 DVSS 0.002679f
C4322 DVDD.n3828 DVSS 0.002679f
C4323 DVDD.n3829 DVSS 0.003698f
C4324 DVDD.n3830 DVSS -0.118241f
C4325 DVDD.n3831 DVSS 0.373549f
C4326 DVDD.n3835 DVSS 0.00493f
C4327 DVDD.n3837 DVSS 0.00493f
C4328 DVDD.n3838 DVSS 0.054232f
C4329 DVDD.n3840 DVSS 0.007181f
C4330 DVDD.n3841 DVSS 0.054232f
C4331 DVDD.n3842 DVSS 0.003923f
C4332 DVDD.n3843 DVSS -0.212535f
C4333 DVDD.n3844 DVSS 0.261329f
C4334 DVDD.n3845 DVSS 0.373549f
C4335 DVDD.n3846 DVSS 0.261329f
C4336 DVDD.n3847 DVSS -0.212535f
C4337 DVDD.n3848 DVSS 0.00493f
C4338 DVDD.n3849 DVSS 0.007181f
C4339 DVDD.n3850 DVSS 0.00134f
C4340 DVDD.n3851 DVSS 0.00134f
C4341 DVDD.n3852 DVSS 0.002679f
C4342 DVDD.n3853 DVSS 0.013397f
C4343 DVDD.n3854 DVSS 0.002679f
C4344 DVDD.n3855 DVSS 0.047684f
C4345 DVDD.n3856 DVSS 0.013397f
C4346 DVDD.n3857 DVSS 0.001451f
C4347 DVDD.n3858 DVSS 0.001427f
C4348 DVDD.n3859 DVSS 0.013397f
C4349 DVDD.n3860 DVSS 0.001538f
C4350 DVDD.n3861 DVSS 0.013397f
C4351 DVDD.n3862 DVSS 0.001538f
C4352 DVDD.n3863 DVSS 0.013397f
C4353 DVDD.n3864 DVSS 0.001538f
C4354 DVDD.n3865 DVSS 0.013397f
C4355 DVDD.n3866 DVSS 0.001538f
C4356 DVDD.n3867 DVSS 0.013397f
C4357 DVDD.n3868 DVSS 0.001538f
C4358 DVDD.n3869 DVSS 0.013397f
C4359 DVDD.n3870 DVSS 0.001538f
C4360 DVDD.n3871 DVSS 0.013397f
C4361 DVDD.n3872 DVSS 0.013397f
C4362 DVDD.n3873 DVSS 0.001402f
C4363 DVDD.n3874 DVSS 0.001476f
C4364 DVDD.n3875 DVSS 0.013397f
C4365 DVDD.n3876 DVSS 0.001538f
C4366 DVDD.n3877 DVSS 0.013397f
C4367 DVDD.n3878 DVSS 0.013397f
C4368 DVDD.n3879 DVSS 0.002345f
C4369 DVDD.n3880 DVSS 0.002679f
C4370 DVDD.n3881 DVSS 0.013397f
C4371 DVDD.n3882 DVSS 0.013397f
C4372 DVDD.n3883 DVSS 0.013397f
C4373 DVDD.n3884 DVSS 0.002679f
C4374 DVDD.n3885 DVSS 0.002679f
C4375 DVDD.n3886 DVSS 0.002679f
C4376 DVDD.n3887 DVSS 0.013397f
C4377 DVDD.n3888 DVSS 0.013397f
C4378 DVDD.t161 DVSS 0.617722f
C4379 DVDD.n3890 DVSS 0.018249f
C4380 DVDD.n3891 DVSS 0.014948f
C4381 DVDD.n3892 DVSS 0.014948f
C4382 DVDD.n3893 DVSS 0.051813f
C4383 DVDD.n3894 DVSS 0.054232f
C4384 DVDD.n3895 DVSS 0.00493f
C4385 DVDD.n3897 DVSS 0.054232f
C4386 DVDD.n3899 DVSS 0.067887f
C4387 DVDD.n3900 DVSS 0.054232f
C4388 DVDD.n3901 DVSS 0.028092f
C4389 DVDD.n3902 DVSS 0.028092f
C4390 DVDD.t162 DVSS 0.198479f
C4391 DVDD.n3904 DVSS 0.00134f
C4392 DVDD.n3905 DVSS 0.00134f
C4393 DVDD.n3906 DVSS 0.031051f
C4394 DVDD.n3907 DVSS 0.063551f
C4395 DVDD.n3908 DVSS 0.052984f
C4396 DVDD.n3909 DVSS 0.054842f
C4397 DVDD.n3910 DVSS 0.063551f
C4398 DVDD.n3911 DVSS 0.031051f
C4399 DVDD.n3912 DVSS 0.063552f
C4400 DVDD.n3913 DVSS 0.054841f
C4401 DVDD.n3914 DVSS 0.052977f
C4402 DVDD.n3915 DVSS 0.011249f
C4403 DVDD.n3916 DVSS 0.00134f
C4404 DVDD.n3917 DVSS 0.00134f
C4405 DVDD.n3918 DVSS 0.014948f
C4406 DVDD.n3919 DVSS 0.014948f
C4407 DVDD.n3920 DVSS 0.001538f
C4408 DVDD.n3921 DVSS 0.013397f
C4409 DVDD.n3922 DVSS 0.001538f
C4410 DVDD.n3923 DVSS 0.013397f
C4411 DVDD.n3924 DVSS 0.001538f
C4412 DVDD.n3925 DVSS 0.013397f
C4413 DVDD.n3926 DVSS 0.001538f
C4414 DVDD.n3927 DVSS 0.013397f
C4415 DVDD.n3928 DVSS 0.001538f
C4416 DVDD.n3929 DVSS 0.013397f
C4417 DVDD.n3930 DVSS 0.013397f
C4418 DVDD.n3931 DVSS 0.001427f
C4419 DVDD.n3932 DVSS 0.001451f
C4420 DVDD.n3933 DVSS 0.013397f
C4421 DVDD.n3934 DVSS 0.001538f
C4422 DVDD.n3935 DVSS 0.047788f
C4423 DVDD.n3936 DVSS 0.103037f
C4424 DVDD.t157 DVSS 0.617722f
C4425 DVDD.n3938 DVSS 0.018249f
C4426 DVDD.n3939 DVSS 0.013397f
C4427 DVDD.n3940 DVSS 0.002679f
C4428 DVDD.n3941 DVSS 0.002679f
C4429 DVDD.n3942 DVSS 0.002679f
C4430 DVDD.n3943 DVSS 0.013397f
C4431 DVDD.n3944 DVSS 0.013397f
C4432 DVDD.n3945 DVSS 0.013397f
C4433 DVDD.n3946 DVSS 0.002679f
C4434 DVDD.n3947 DVSS 0.002679f
C4435 DVDD.n3948 DVSS 0.002345f
C4436 DVDD.n3949 DVSS 0.013397f
C4437 DVDD.n3950 DVSS 0.001538f
C4438 DVDD.n3951 DVSS 0.013397f
C4439 DVDD.n3952 DVSS 0.013397f
C4440 DVDD.n3953 DVSS 0.013397f
C4441 DVDD.n3954 DVSS 0.001402f
C4442 DVDD.n3955 DVSS 0.00134f
C4443 DVDD.n3956 DVSS 0.01233f
C4444 DVDD.n3957 DVSS 0.014849f
C4445 DVDD.n3958 DVSS 0.024661f
C4446 DVDD.n3959 DVSS 0.024661f
C4447 DVDD.n3960 DVSS 0.024661f
C4448 DVDD.n3961 DVSS 0.024661f
C4449 DVDD.n3962 DVSS 0.024661f
C4450 DVDD.n3963 DVSS 0.023706f
C4451 DVDD.n3964 DVSS 0.024661f
C4452 DVDD.n3965 DVSS 0.024661f
C4453 DVDD.n3966 DVSS 0.024661f
C4454 DVDD.n3967 DVSS 0.024661f
C4455 DVDD.n3968 DVSS 0.024661f
C4456 DVDD.n3969 DVSS 0.024661f
C4457 DVDD.n3970 DVSS 0.024661f
C4458 DVDD.n3971 DVSS 0.024661f
C4459 DVDD.n3972 DVSS 0.024661f
C4460 DVDD.n3973 DVSS 0.024661f
C4461 DVDD.n3974 DVSS 0.024661f
C4462 DVDD.n3975 DVSS 0.024661f
C4463 DVDD.n3976 DVSS 0.024661f
C4464 DVDD.n3977 DVSS 0.024661f
C4465 DVDD.n3978 DVSS 0.024661f
C4466 DVDD.n3979 DVSS 0.024661f
C4467 DVDD.n3980 DVSS 0.024661f
C4468 DVDD.n3981 DVSS 0.024661f
C4469 DVDD.n3982 DVSS 0.024661f
C4470 DVDD.n3983 DVSS 0.024661f
C4471 DVDD.n3984 DVSS 0.024661f
C4472 DVDD.n3985 DVSS 0.024661f
C4473 DVDD.n3986 DVSS 0.024661f
C4474 DVDD.n3987 DVSS 0.024661f
C4475 DVDD.n3988 DVSS 0.024661f
C4476 DVDD.n3989 DVSS 0.014849f
C4477 DVDD.n3990 DVSS 0.024661f
C4478 DVDD.n3991 DVSS 0.024661f
C4479 DVDD.n3992 DVSS 0.024661f
C4480 DVDD.n3993 DVSS 0.024661f
C4481 DVDD.n3994 DVSS 0.024661f
C4482 DVDD.n3995 DVSS 0.024661f
C4483 DVDD.n3996 DVSS 0.024661f
C4484 DVDD.n3997 DVSS 0.010767f
C4485 DVDD.n3998 DVSS 0.011723f
C4486 DVDD.n4000 DVSS 0.107715f
C4487 DVDD.n4001 DVSS 0.01233f
C4488 DVDD.n4002 DVSS 0.014501f
C4489 DVDD.n4003 DVSS 0.024661f
C4490 DVDD.n4004 DVSS 0.024661f
C4491 DVDD.n4005 DVSS 0.024661f
C4492 DVDD.n4006 DVSS 0.024661f
C4493 DVDD.n4007 DVSS 0.024661f
C4494 DVDD.n4008 DVSS 0.024661f
C4495 DVDD.n4009 DVSS 0.024661f
C4496 DVDD.n4010 DVSS 0.024661f
C4497 DVDD.n4011 DVSS 0.024661f
C4498 DVDD.n4012 DVSS 0.024661f
C4499 DVDD.n4013 DVSS 0.024661f
C4500 DVDD.n4014 DVSS 0.024661f
C4501 DVDD.n4015 DVSS 0.024661f
C4502 DVDD.n4016 DVSS 0.024661f
C4503 DVDD.n4017 DVSS 0.024661f
C4504 DVDD.n4018 DVSS 0.024661f
C4505 DVDD.n4019 DVSS 0.024661f
C4506 DVDD.n4020 DVSS 0.024661f
C4507 DVDD.n4021 DVSS 0.024661f
C4508 DVDD.n4022 DVSS 0.024661f
C4509 DVDD.n4023 DVSS 0.024661f
C4510 DVDD.n4024 DVSS 0.024661f
C4511 DVDD.n4025 DVSS 0.024661f
C4512 DVDD.n4026 DVSS 0.024661f
C4513 DVDD.n4027 DVSS 0.024661f
C4514 DVDD.n4028 DVSS 0.024661f
C4515 DVDD.n4029 DVSS 0.024661f
C4516 DVDD.n4030 DVSS 0.024661f
C4517 DVDD.n4031 DVSS 0.024661f
C4518 DVDD.n4032 DVSS 0.024661f
C4519 DVDD.n4033 DVSS 0.024661f
C4520 DVDD.n4034 DVSS 0.024053f
C4521 DVDD.n4035 DVSS 0.01233f
C4522 DVDD.n4036 DVSS 0.022708f
C4523 DVDD.n4037 DVSS 0.01233f
C4524 DVDD.n4038 DVSS 0.014501f
C4525 DVDD.n4039 DVSS 0.024661f
C4526 DVDD.n4040 DVSS 0.024661f
C4527 DVDD.n4041 DVSS 0.024661f
C4528 DVDD.n4042 DVSS 0.024661f
C4529 DVDD.n4043 DVSS 0.024661f
C4530 DVDD.n4044 DVSS 0.024661f
C4531 DVDD.n4045 DVSS 0.024661f
C4532 DVDD.n4046 DVSS 0.024661f
C4533 DVDD.n4047 DVSS 0.024661f
C4534 DVDD.n4048 DVSS 0.024661f
C4535 DVDD.n4049 DVSS 0.024661f
C4536 DVDD.n4050 DVSS 0.024661f
C4537 DVDD.n4051 DVSS 0.024661f
C4538 DVDD.n4052 DVSS 0.024661f
C4539 DVDD.n4053 DVSS 0.024661f
C4540 DVDD.n4054 DVSS 0.024661f
C4541 DVDD.n4055 DVSS 0.024661f
C4542 DVDD.n4056 DVSS 0.024661f
C4543 DVDD.n4057 DVSS 0.024661f
C4544 DVDD.n4058 DVSS 0.024661f
C4545 DVDD.n4059 DVSS 0.024661f
C4546 DVDD.n4060 DVSS 0.024661f
C4547 DVDD.n4061 DVSS 0.024661f
C4548 DVDD.n4062 DVSS 0.024661f
C4549 DVDD.n4063 DVSS 0.024661f
C4550 DVDD.n4064 DVSS 0.024661f
C4551 DVDD.n4065 DVSS 0.024661f
C4552 DVDD.n4066 DVSS 0.024661f
C4553 DVDD.n4067 DVSS 0.024661f
C4554 DVDD.n4068 DVSS 0.024661f
C4555 DVDD.n4069 DVSS 0.024661f
C4556 DVDD.n4070 DVSS 0.024661f
C4557 DVDD.n4071 DVSS 0.024661f
C4558 DVDD.n4072 DVSS 0.024661f
C4559 DVDD.n4073 DVSS 0.024661f
C4560 DVDD.n4074 DVSS 0.024661f
C4561 DVDD.n4075 DVSS 0.024661f
C4562 DVDD.n4076 DVSS 0.024661f
C4563 DVDD.n4077 DVSS 0.024661f
C4564 DVDD.n4078 DVSS 0.118858f
C4565 DVDD.n4079 DVSS 0.032461f
C4566 DVDD.n4080 DVSS 0.012678f
C4567 DVDD.n4081 DVSS 0.024661f
C4568 DVDD.n4082 DVSS 0.02223f
C4569 DVDD.n4083 DVSS 0.02223f
C4570 DVDD.n4084 DVSS 0.024661f
C4571 DVDD.n4085 DVSS 0.024661f
C4572 DVDD.n4086 DVSS 0.024661f
C4573 DVDD.n4087 DVSS 0.024661f
C4574 DVDD.n4088 DVSS 0.024661f
C4575 DVDD.n4089 DVSS 0.024661f
C4576 DVDD.n4090 DVSS 0.024661f
C4577 DVDD.n4091 DVSS 0.024661f
C4578 DVDD.n4092 DVSS 0.024661f
C4579 DVDD.n4093 DVSS 0.024661f
C4580 DVDD.n4094 DVSS 0.024661f
C4581 DVDD.n4095 DVSS 0.024661f
C4582 DVDD.n4096 DVSS 0.024661f
C4583 DVDD.n4097 DVSS 0.024661f
C4584 DVDD.n4098 DVSS 0.024661f
C4585 DVDD.n4099 DVSS 0.024661f
C4586 DVDD.n4100 DVSS 0.024661f
C4587 DVDD.n4101 DVSS 0.024661f
C4588 DVDD.n4102 DVSS 0.024661f
C4589 DVDD.n4103 DVSS 0.024661f
C4590 DVDD.n4104 DVSS 0.024661f
C4591 DVDD.n4105 DVSS 0.024661f
C4592 DVDD.n4106 DVSS 0.024661f
C4593 DVDD.n4107 DVSS 0.024661f
C4594 DVDD.n4108 DVSS 0.020233f
C4595 DVDD.n4109 DVSS 0.003076f
C4596 DVDD.n4110 DVSS 0.003076f
C4597 DVDD.n4111 DVSS 0.003076f
C4598 DVDD.n4112 DVSS 0.01233f
C4599 DVDD.n4113 DVSS 0.003076f
C4600 DVDD.n4114 DVSS 0.003076f
C4601 DVDD.n4115 DVSS 0.01233f
C4602 DVDD.n4116 DVSS 0.035774f
C4603 DVDD.t158 DVSS 0.617722f
C4604 DVDD.n4118 DVSS 0.204625f
C4605 DVDD.n4119 DVSS 0.200207f
C4606 DVDD.n4120 DVSS 0.025152f
C4607 DVDD.n4121 DVSS 0.016319f
C4608 DVDD.n4122 DVSS 0.004474f
C4609 DVDD.n4123 DVSS 0.002679f
C4610 DVDD.n4124 DVSS 0.00493f
C4611 DVDD.n4125 DVSS 0.00493f
C4612 DVDD.n4126 DVSS 0.00493f
C4613 DVDD.n4127 DVSS 0.002679f
C4614 DVDD.n4128 DVSS 0.002679f
C4615 DVDD.n4129 DVSS 0.002679f
C4616 DVDD.n4130 DVSS 0.00493f
C4617 DVDD.n4131 DVSS 0.00493f
C4618 DVDD.n4132 DVSS 0.00493f
C4619 DVDD.n4133 DVSS 0.002679f
C4620 DVDD.n4134 DVSS 0.002679f
C4621 DVDD.n4135 DVSS 0.002679f
C4622 DVDD.n4136 DVSS 0.00493f
C4623 DVDD.n4137 DVSS 0.00493f
C4624 DVDD.n4138 DVSS 0.00493f
C4625 DVDD.n4139 DVSS 0.002679f
C4626 DVDD.n4140 DVSS 0.002679f
C4627 DVDD.n4141 DVSS 0.002679f
C4628 DVDD.n4142 DVSS 0.00493f
C4629 DVDD.n4143 DVSS 0.00493f
C4630 DVDD.n4144 DVSS 0.00493f
C4631 DVDD.n4145 DVSS 0.002679f
C4632 DVDD.n4146 DVSS 0.002679f
C4633 DVDD.n4147 DVSS 0.002679f
C4634 DVDD.n4148 DVSS 0.00493f
C4635 DVDD.n4149 DVSS 0.00493f
C4636 DVDD.n4150 DVSS 0.003698f
C4637 DVDD.n4151 DVSS 0.002679f
C4638 DVDD.n4152 DVSS 0.002679f
C4639 DVDD.n4153 DVSS 0.003698f
C4640 DVDD.n4154 DVSS 0.00493f
C4641 DVDD.n4155 DVSS 0.00493f
C4642 DVDD.n4156 DVSS 0.002679f
C4643 DVDD.n4157 DVSS 0.002679f
C4644 DVDD.n4158 DVSS 0.002679f
C4645 DVDD.n4159 DVSS 0.00493f
C4646 DVDD.n4160 DVSS 0.00493f
C4647 DVDD.n4161 DVSS 0.00493f
C4648 DVDD.n4162 DVSS 0.002679f
C4649 DVDD.n4163 DVSS 0.002679f
C4650 DVDD.n4164 DVSS 0.002679f
C4651 DVDD.n4165 DVSS 0.00493f
C4652 DVDD.n4166 DVSS 0.00493f
C4653 DVDD.n4167 DVSS 0.00493f
C4654 DVDD.n4168 DVSS 0.002679f
C4655 DVDD.n4169 DVSS 0.002679f
C4656 DVDD.n4170 DVSS 0.002679f
C4657 DVDD.n4171 DVSS 0.00493f
C4658 DVDD.n4172 DVSS 0.00493f
C4659 DVDD.n4173 DVSS 0.00493f
C4660 DVDD.n4174 DVSS 0.002679f
C4661 DVDD.n4175 DVSS 0.002679f
C4662 DVDD.n4176 DVSS 0.002679f
C4663 DVDD.n4177 DVSS 0.00493f
C4664 DVDD.n4178 DVSS 0.00493f
C4665 DVDD.n4179 DVSS 0.00493f
C4666 DVDD.n4180 DVSS 0.002679f
C4667 DVDD.n4181 DVSS 0.003582f
C4668 DVDD.n4182 DVSS 0.003388f
C4669 DVDD.n4183 DVSS 0.001538f
C4670 DVDD.n4184 DVSS 0.005683f
C4671 DVDD.n4185 DVSS 0.052292f
C4672 DVDD.n4186 DVSS 0.051813f
C4673 DVDD.n4187 DVSS 0.001538f
C4674 DVDD.n4188 DVSS 0.003076f
C4675 DVDD.n4189 DVSS 0.003076f
C4676 DVDD.n4190 DVSS 0.003076f
C4677 DVDD.n4191 DVSS 0.001538f
C4678 DVDD.n4192 DVSS 0.001662f
C4679 DVDD.n4193 DVSS 0.001464f
C4680 DVDD.n4194 DVSS 0.00134f
C4681 DVDD.n4195 DVSS 0.00134f
C4682 DVDD.n4196 DVSS 0.011236f
C4683 DVDD.n4197 DVSS 0.052992f
C4684 DVDD.n4198 DVSS 0.063551f
C4685 DVDD.n4199 DVSS 0.028092f
C4686 DVDD.n4200 DVSS 0.063552f
C4687 DVDD.n4201 DVSS 0.05297f
C4688 DVDD.n4202 DVSS 0.00134f
C4689 DVDD.n4203 DVSS 0.011242f
C4690 DVDD.n4204 DVSS 0.051813f
C4691 DVDD.n4205 DVSS 0.052292f
C4692 DVDD.n4206 DVSS 0.005683f
C4693 DVDD.n4207 DVSS 0.001538f
C4694 DVDD.n4208 DVSS 0.002928f
C4695 DVDD.n4209 DVSS 0.001538f
C4696 DVDD.n4210 DVSS 0.001538f
C4697 DVDD.n4211 DVSS 0.080216f
C4698 DVDD.n4212 DVSS 0.588581f
C4699 DVDD.n4213 DVSS 0.001538f
C4700 DVDD.n4214 DVSS 0.003076f
C4701 DVDD.n4215 DVSS 0.003052f
C4702 DVDD.n4216 DVSS 4.9e-19
C4703 DVDD.n4217 DVSS 6.32e-19
C4704 DVDD.n4219 DVSS 9.8e-19
C4705 DVDD.n4220 DVSS 0.001161f
C4706 DVDD.n4221 DVSS 9.8e-19
C4707 DVDD.n4222 DVSS 0.001161f
C4708 DVDD.n4223 DVSS 9.8e-19
C4709 DVDD.n4224 DVSS 0.001161f
C4710 DVDD.n4225 DVSS 9.8e-19
C4711 DVDD.n4226 DVSS 0.001083f
C4712 DVDD.n4227 DVSS 9.8e-19
C4713 DVDD.n4228 DVSS 0.001161f
C4714 DVDD.n4230 DVSS 0.001161f
C4715 DVDD.n4232 DVSS 0.001161f
C4716 DVDD.n4233 DVSS 9.8e-19
C4717 DVDD.n4234 DVSS 9.8e-19
C4718 DVDD.n4235 DVSS 9.8e-19
C4719 DVDD.n4236 DVSS 0.001161f
C4720 DVDD.n4238 DVSS 0.001161f
C4721 DVDD.n4240 DVSS 0.001161f
C4722 DVDD.n4241 DVSS 9.8e-19
C4723 DVDD.n4242 DVSS 9.8e-19
C4724 DVDD.n4243 DVSS 9.8e-19
C4725 DVDD.n4244 DVSS 0.001161f
C4726 DVDD.n4246 DVSS 0.001161f
C4727 DVDD.n4248 DVSS 0.001161f
C4728 DVDD.n4249 DVSS 9.8e-19
C4729 DVDD.n4250 DVSS 9.8e-19
C4730 DVDD.n4251 DVSS 9.8e-19
C4731 DVDD.n4252 DVSS 0.001161f
C4732 DVDD.n4254 DVSS 0.001161f
C4733 DVDD.n4255 DVSS 0.001161f
C4734 DVDD.n4256 DVSS 9.8e-19
C4735 DVDD.n4257 DVSS 9.8e-19
C4736 DVDD.n4258 DVSS 0.001161f
C4737 DVDD.n4259 DVSS 0.001161f
C4738 DVDD.n4261 DVSS 8.2e-19
C4739 DVDD.n4262 DVSS 0.001161f
C4740 DVDD.n4263 DVSS 9.8e-19
C4741 DVDD.n4265 DVSS 0.001161f
C4742 DVDD.n4266 DVSS 9.8e-19
C4743 DVDD.n4268 DVSS 0.001161f
C4744 DVDD.n4269 DVSS 9.8e-19
C4745 DVDD.n4271 DVSS 0.001161f
C4746 DVDD.n4272 DVSS 9.8e-19
C4747 DVDD.n4274 DVSS 0.001161f
C4748 DVDD.n4275 DVSS 9.8e-19
C4749 DVDD.n4277 DVSS 0.001161f
C4750 DVDD.n4278 DVSS 5.28e-19
C4751 DVDD.n4279 DVSS 0.001161f
C4752 DVDD.n4281 DVSS 0.001161f
C4753 DVDD.n4282 DVSS 0.001161f
C4754 DVDD.n4283 DVSS 9.8e-19
C4755 DVDD.n4284 DVSS 9.8e-19
C4756 DVDD.n4285 DVSS 9.8e-19
C4757 DVDD.n4286 DVSS 0.001161f
C4758 DVDD.n4288 DVSS 0.001161f
C4759 DVDD.n4289 DVSS 0.001161f
C4760 DVDD.n4290 DVSS 9.8e-19
C4761 DVDD.n4291 DVSS 9.8e-19
C4762 DVDD.n4292 DVSS 9.8e-19
C4763 DVDD.n4293 DVSS 0.001161f
C4764 DVDD.n4295 DVSS 0.001161f
C4765 DVDD.n4296 DVSS 0.001161f
C4766 DVDD.n4297 DVSS 9.8e-19
C4767 DVDD.n4298 DVSS 9.8e-19
C4768 DVDD.n4299 DVSS 9.8e-19
C4769 DVDD.n4300 DVSS 0.001161f
C4770 DVDD.n4302 DVSS 0.001161f
C4771 DVDD.n4303 DVSS 0.001161f
C4772 DVDD.n4304 DVSS 9.8e-19
C4773 DVDD.n4305 DVSS 9.8e-19
C4774 DVDD.n4306 DVSS 9.8e-19
C4775 DVDD.n4307 DVSS 0.001161f
C4776 DVDD.n4309 DVSS 0.001161f
C4777 DVDD.n4310 DVSS 0.001161f
C4778 DVDD.n4311 DVSS 9.8e-19
C4779 DVDD.n4312 DVSS 9.8e-19
C4780 DVDD.n4313 DVSS 9.8e-19
C4781 DVDD.n4314 DVSS 0.001161f
C4782 DVDD.n4316 DVSS 0.001161f
C4783 DVDD.n4317 DVSS 0.001161f
C4784 DVDD.n4318 DVSS 5.09e-19
C4785 DVDD.n4319 DVSS 4.9e-19
C4786 DVDD.n4320 DVSS 0.001538f
C4787 DVDD.n4321 DVSS 0.001563f
C4788 DVDD.n4322 DVSS 0.342994f
C4789 DVDD.n4323 DVSS 0.003076f
C4790 DVDD.n4324 DVSS 0.003076f
C4791 DVDD.n4325 DVSS 0.01233f
C4792 DVDD.n4326 DVSS 0.019885f
C4793 DVDD.n4327 DVSS 0.024661f
C4794 DVDD.n4328 DVSS 0.024661f
C4795 DVDD.n4329 DVSS 0.024661f
C4796 DVDD.n4330 DVSS 0.024661f
C4797 DVDD.n4331 DVSS 0.024661f
C4798 DVDD.n4332 DVSS 0.024661f
C4799 DVDD.n4333 DVSS 0.024661f
C4800 DVDD.n4334 DVSS 0.024661f
C4801 DVDD.n4335 DVSS 0.024661f
C4802 DVDD.n4336 DVSS 0.024661f
C4803 DVDD.n4337 DVSS 0.024661f
C4804 DVDD.n4338 DVSS 0.024661f
C4805 DVDD.n4339 DVSS 0.024661f
C4806 DVDD.n4340 DVSS 0.024661f
C4807 DVDD.n4341 DVSS 0.024661f
C4808 DVDD.n4342 DVSS 0.024661f
C4809 DVDD.n4343 DVSS 0.024661f
C4810 DVDD.n4344 DVSS 0.024661f
C4811 DVDD.n4345 DVSS 0.024661f
C4812 DVDD.n4346 DVSS 0.024661f
C4813 DVDD.n4347 DVSS 0.024661f
C4814 DVDD.n4348 DVSS 0.024661f
C4815 DVDD.n4349 DVSS 0.024661f
C4816 DVDD.n4350 DVSS 0.024661f
C4817 DVDD.n4351 DVSS 0.024661f
C4818 DVDD.n4352 DVSS 0.024661f
C4819 DVDD.n4353 DVSS 0.024661f
C4820 DVDD.n4354 DVSS 0.024661f
C4821 DVDD.n4355 DVSS 0.024661f
C4822 DVDD.n4356 DVSS 0.024661f
C4823 DVDD.n4357 DVSS 0.024661f
C4824 DVDD.n4358 DVSS 0.010767f
C4825 DVDD.n4359 DVSS 0.024661f
C4826 DVDD.n4360 DVSS 0.023706f
C4827 DVDD.n4361 DVSS 0.024661f
C4828 DVDD.n4362 DVSS 0.024661f
C4829 DVDD.n4363 DVSS 0.024661f
C4830 DVDD.n4364 DVSS 0.024661f
C4831 DVDD.n4365 DVSS 0.024661f
C4832 DVDD.n4366 DVSS 0.024661f
C4833 DVDD.n4367 DVSS 0.024661f
C4834 DVDD.n4368 DVSS 0.024661f
C4835 DVDD.n4369 DVSS 0.024661f
C4836 DVDD.n4370 DVSS 0.024661f
C4837 DVDD.n4371 DVSS 0.024661f
C4838 DVDD.n4372 DVSS 0.024661f
C4839 DVDD.n4373 DVSS 0.024661f
C4840 DVDD.n4374 DVSS 0.024661f
C4841 DVDD.n4375 DVSS 0.024661f
C4842 DVDD.n4376 DVSS 0.024661f
C4843 DVDD.n4377 DVSS 0.024661f
C4844 DVDD.n4378 DVSS 0.024661f
C4845 DVDD.n4379 DVSS 0.024661f
C4846 DVDD.n4380 DVSS 0.024661f
C4847 DVDD.n4381 DVSS 0.024661f
C4848 DVDD.n4382 DVSS 0.024661f
C4849 DVDD.n4383 DVSS 0.024661f
C4850 DVDD.n4384 DVSS 0.024661f
C4851 DVDD.n4385 DVSS 0.024661f
C4852 DVDD.n4386 DVSS 0.024661f
C4853 DVDD.n4387 DVSS 0.024661f
C4854 DVDD.n4388 DVSS 0.024661f
C4855 DVDD.n4389 DVSS 0.024661f
C4856 DVDD.n4390 DVSS 0.024661f
C4857 DVDD.n4391 DVSS 0.024661f
C4858 DVDD.n4392 DVSS 0.024661f
C4859 DVDD.n4393 DVSS 0.024661f
C4860 DVDD.n4394 DVSS 0.024661f
C4861 DVDD.n4395 DVSS 0.024661f
C4862 DVDD.n4396 DVSS 0.024661f
C4863 DVDD.n4397 DVSS 0.024661f
C4864 DVDD.n4398 DVSS 0.024661f
C4865 DVDD.n4399 DVSS 0.024661f
C4866 DVDD.n4400 DVSS 0.024661f
C4867 DVDD.n4401 DVSS 0.024661f
C4868 DVDD.n4402 DVSS 0.024661f
C4869 DVDD.n4403 DVSS 0.024661f
C4870 DVDD.n4404 DVSS 0.024661f
C4871 DVDD.n4405 DVSS 0.024661f
C4872 DVDD.n4406 DVSS 0.024661f
C4873 DVDD.n4407 DVSS 0.024661f
C4874 DVDD.n4408 DVSS 0.024661f
C4875 DVDD.n4409 DVSS 0.010767f
C4876 DVDD.n4410 DVSS 0.024661f
C4877 DVDD.n4411 DVSS 0.024661f
C4878 DVDD.n4412 DVSS 0.014501f
C4879 DVDD.n4413 DVSS 0.024661f
C4880 DVDD.n4414 DVSS 0.024661f
C4881 DVDD.n4415 DVSS 0.024661f
C4882 DVDD.n4416 DVSS 0.024661f
C4883 DVDD.n4417 DVSS 0.024661f
C4884 DVDD.n4418 DVSS 0.024661f
C4885 DVDD.n4419 DVSS 0.024661f
C4886 DVDD.n4420 DVSS 0.024661f
C4887 DVDD.n4421 DVSS 0.024661f
C4888 DVDD.n4422 DVSS 0.024661f
C4889 DVDD.n4423 DVSS 0.024661f
C4890 DVDD.n4424 DVSS 0.024661f
C4891 DVDD.n4425 DVSS 0.024661f
C4892 DVDD.n4426 DVSS 0.024661f
C4893 DVDD.n4427 DVSS 0.024661f
C4894 DVDD.n4428 DVSS 0.024661f
C4895 DVDD.n4429 DVSS 0.024661f
C4896 DVDD.n4430 DVSS 0.024661f
C4897 DVDD.n4431 DVSS 0.024661f
C4898 DVDD.n4432 DVSS 0.024661f
C4899 DVDD.n4433 DVSS 0.024661f
C4900 DVDD.n4434 DVSS 0.024661f
C4901 DVDD.n4435 DVSS 0.024661f
C4902 DVDD.n4436 DVSS 0.024661f
C4903 DVDD.n4437 DVSS 0.024661f
C4904 DVDD.n4438 DVSS 0.024661f
C4905 DVDD.n4439 DVSS 0.024661f
C4906 DVDD.n4440 DVSS 0.024661f
C4907 DVDD.n4441 DVSS 0.024661f
C4908 DVDD.n4442 DVSS 0.024661f
C4909 DVDD.n4443 DVSS 0.024661f
C4910 DVDD.n4444 DVSS 0.024661f
C4911 DVDD.n4445 DVSS 0.024661f
C4912 DVDD.n4446 DVSS 0.024661f
C4913 DVDD.n4447 DVSS 0.024661f
C4914 DVDD.n4448 DVSS 0.024661f
C4915 DVDD.n4449 DVSS 0.024661f
C4916 DVDD.n4450 DVSS 0.024661f
C4917 DVDD.n4451 DVSS 0.024661f
C4918 DVDD.n4452 DVSS 0.024661f
C4919 DVDD.n4453 DVSS 0.024661f
C4920 DVDD.n4454 DVSS 0.024053f
C4921 DVDD.n4455 DVSS 0.024661f
C4922 DVDD.n4456 DVSS 0.024661f
C4923 DVDD.n4457 DVSS 0.024661f
C4924 DVDD.n4458 DVSS 0.024661f
C4925 DVDD.n4459 DVSS 0.024661f
C4926 DVDD.n4460 DVSS 0.024661f
C4927 DVDD.n4461 DVSS 0.024661f
C4928 DVDD.n4462 DVSS 0.024661f
C4929 DVDD.n4463 DVSS 0.024661f
C4930 DVDD.n4464 DVSS 0.024661f
C4931 DVDD.n4465 DVSS 0.024661f
C4932 DVDD.n4466 DVSS 0.024661f
C4933 DVDD.n4467 DVSS 0.024661f
C4934 DVDD.n4468 DVSS 0.024661f
C4935 DVDD.n4469 DVSS 0.024661f
C4936 DVDD.n4470 DVSS 0.024661f
C4937 DVDD.n4471 DVSS 0.024661f
C4938 DVDD.n4472 DVSS 0.024661f
C4939 DVDD.n4473 DVSS 0.024661f
C4940 DVDD.n4474 DVSS 0.024661f
C4941 DVDD.n4475 DVSS 0.024661f
C4942 DVDD.n4476 DVSS 0.024661f
C4943 DVDD.n4477 DVSS 0.024661f
C4944 DVDD.n4478 DVSS 0.024661f
C4945 DVDD.n4479 DVSS 0.024661f
C4946 DVDD.n4480 DVSS 0.024661f
C4947 DVDD.n4481 DVSS 0.024661f
C4948 DVDD.n4482 DVSS 0.024661f
C4949 DVDD.n4483 DVSS 0.024661f
C4950 DVDD.n4484 DVSS 0.024661f
C4951 DVDD.n4485 DVSS 0.014501f
C4952 DVDD.n4486 DVSS 0.008245f
C4953 DVDD.n4488 DVSS 0.01233f
C4954 DVDD.n4489 DVSS 0.008245f
C4955 DVDD.n4491 DVSS 0.011375f
C4956 DVDD.n4492 DVSS 0.008245f
C4957 DVDD.n4493 DVSS 0.01233f
C4958 DVDD.n4494 DVSS 0.069283f
C4959 DVDD.n4495 DVSS 0.008245f
C4960 DVDD.n4496 DVSS 0.006751f
C4961 DVDD.n4497 DVSS 0.0032f
C4962 DVDD.n4498 DVSS 0.003076f
C4963 DVDD.n4499 DVSS 0.003523f
C4964 DVDD.n4500 DVSS 0.003076f
C4965 DVDD.n4501 DVSS 0.008245f
C4966 DVDD.n4502 DVSS 0.023073f
C4967 DVDD.n4503 DVSS 0.003076f
C4968 DVDD.n4504 DVSS 0.024004f
C4969 DVDD.n4505 DVSS 0.003399f
C4970 DVDD.n4506 DVSS 0.008245f
C4971 DVDD.n4507 DVSS 0.025492f
C4972 DVDD.n4508 DVSS 0.052845f
C4973 DVDD.n4509 DVSS 0.052845f
C4974 DVDD.n4510 DVSS 0.052845f
C4975 DVDD.n4511 DVSS 0.150127f
C4976 DVDD.n4512 DVSS 0.052845f
C4977 DVDD.n4513 DVSS 0.023073f
C4978 DVDD.n4514 DVSS 0.026423f
C4979 DVDD.n4515 DVSS 0.003076f
C4980 DVDD.n4516 DVSS 0.003076f
C4981 DVDD.n4517 DVSS 0.003076f
C4982 DVDD.n4518 DVSS 0.023073f
C4983 DVDD.n4519 DVSS 0.026423f
C4984 DVDD.n4520 DVSS 0.003076f
C4985 DVDD.n4521 DVSS 0.003076f
C4986 DVDD.n4522 DVSS 0.003523f
C4987 DVDD.n4523 DVSS 0.008245f
C4988 DVDD.n4524 DVSS 0.008245f
C4989 DVDD.n4525 DVSS 0.008245f
C4990 DVDD.n4526 DVSS 0.003523f
C4991 DVDD.n4527 DVSS 0.003076f
C4992 DVDD.n4528 DVSS 0.007046f
C4993 DVDD.n4529 DVSS 0.007046f
C4994 DVDD.n4530 DVSS 0.019986f
C4995 DVDD.n4531 DVSS 0.007046f
C4996 DVDD.n4532 DVSS 0.007046f
C4997 DVDD.n4533 DVSS 0.003076f
C4998 DVDD.n4534 DVSS 0.00698f
C4999 DVDD.n4535 DVSS 0.069283f
C5000 DVDD.n4536 DVSS 0.052416f
C5001 DVDD.n4537 DVSS 0.025852f
C5002 DVDD.n4538 DVSS 0.025852f
C5003 DVDD.n4539 DVSS 0.001538f
C5004 DVDD.n4540 DVSS 0.003076f
C5005 DVDD.n4541 DVSS 0.003076f
C5006 DVDD.n4542 DVSS 0.001538f
C5007 DVDD.n4543 DVSS 0.001563f
C5008 DVDD.n4544 DVSS 0.001538f
C5009 DVDD.n4545 DVSS 4.9e-19
C5010 DVDD.n4546 DVSS 9.8e-19
C5011 DVDD.n4548 DVSS 0.001161f
C5012 DVDD.n4549 DVSS 9.8e-19
C5013 DVDD.n4551 DVSS 0.001161f
C5014 DVDD.n4552 DVSS 9.8e-19
C5015 DVDD.n4554 DVSS 0.001161f
C5016 DVDD.n4555 DVSS 9.8e-19
C5017 DVDD.n4557 DVSS 0.001161f
C5018 DVDD.n4558 DVSS 9.8e-19
C5019 DVDD.n4561 DVSS 0.001161f
C5020 DVDD.n4562 DVSS 8.2e-19
C5021 DVDD.n4563 DVSS 9.8e-19
C5022 DVDD.n4564 DVSS 0.001161f
C5023 DVDD.n4566 DVSS 0.001161f
C5024 DVDD.n4567 DVSS 0.001161f
C5025 DVDD.n4568 DVSS 9.8e-19
C5026 DVDD.n4569 DVSS 9.8e-19
C5027 DVDD.n4570 DVSS 9.8e-19
C5028 DVDD.n4571 DVSS 0.001161f
C5029 DVDD.n4573 DVSS 0.001161f
C5030 DVDD.n4574 DVSS 0.001161f
C5031 DVDD.n4575 DVSS 9.8e-19
C5032 DVDD.n4576 DVSS 9.8e-19
C5033 DVDD.n4577 DVSS 9.8e-19
C5034 DVDD.n4578 DVSS 0.001161f
C5035 DVDD.n4580 DVSS 0.001161f
C5036 DVDD.n4581 DVSS 0.001161f
C5037 DVDD.n4582 DVSS 9.8e-19
C5038 DVDD.n4583 DVSS 9.8e-19
C5039 DVDD.n4584 DVSS 9.8e-19
C5040 DVDD.n4585 DVSS 0.001161f
C5041 DVDD.n4587 DVSS 0.001161f
C5042 DVDD.n4588 DVSS 0.001161f
C5043 DVDD.n4589 DVSS 9.8e-19
C5044 DVDD.n4590 DVSS 9.8e-19
C5045 DVDD.n4591 DVSS 9.8e-19
C5046 DVDD.n4592 DVSS 0.001161f
C5047 DVDD.n4594 DVSS 0.001161f
C5048 DVDD.n4595 DVSS 0.001161f
C5049 DVDD.n4596 DVSS 9.8e-19
C5050 DVDD.n4597 DVSS 9.8e-19
C5051 DVDD.n4598 DVSS 5.28e-19
C5052 DVDD.n4599 DVSS 0.001161f
C5053 DVDD.n4601 DVSS 0.001161f
C5054 DVDD.n4602 DVSS 0.001161f
C5055 DVDD.n4603 DVSS 9.24e-19
C5056 DVDD.n4604 DVSS 9.8e-19
C5057 DVDD.n4605 DVSS 9.8e-19
C5058 DVDD.n4606 DVSS 0.001161f
C5059 DVDD.n4608 DVSS 0.001161f
C5060 DVDD.n4609 DVSS 0.001161f
C5061 DVDD.n4610 DVSS 9.8e-19
C5062 DVDD.n4611 DVSS 9.8e-19
C5063 DVDD.n4612 DVSS 9.8e-19
C5064 DVDD.n4613 DVSS 0.001161f
C5065 DVDD.n4615 DVSS 0.001161f
C5066 DVDD.n4616 DVSS 0.001161f
C5067 DVDD.n4617 DVSS 9.8e-19
C5068 DVDD.n4618 DVSS 9.8e-19
C5069 DVDD.n4619 DVSS 9.8e-19
C5070 DVDD.n4620 DVSS 0.001161f
C5071 DVDD.n4622 DVSS 0.001161f
C5072 DVDD.n4623 DVSS 0.001161f
C5073 DVDD.n4624 DVSS 9.8e-19
C5074 DVDD.n4625 DVSS 9.8e-19
C5075 DVDD.n4626 DVSS 9.8e-19
C5076 DVDD.n4627 DVSS 0.001161f
C5077 DVDD.n4629 DVSS 0.001161f
C5078 DVDD.n4630 DVSS 0.001161f
C5079 DVDD.n4631 DVSS 9.8e-19
C5080 DVDD.n4632 DVSS 9.8e-19
C5081 DVDD.n4633 DVSS 9.8e-19
C5082 DVDD.n4634 DVSS 0.001161f
C5083 DVDD.n4636 DVSS 0.001161f
C5084 DVDD.n4637 DVSS 0.001161f
C5085 DVDD.n4638 DVSS 9.43e-19
C5086 DVDD.n4639 DVSS 4.9e-19
C5087 DVDD.n4640 DVSS 0.004122f
C5088 DVDD.n4641 DVSS 9.8e-19
C5089 DVDD.n4642 DVSS 5.09e-19
C5090 DVDD.n4643 DVSS 0.001161f
C5091 DVDD.n4645 DVSS 0.001161f
C5092 DVDD.n4646 DVSS 0.001161f
C5093 DVDD.n4647 DVSS 9.43e-19
C5094 DVDD.n4648 DVSS 9.8e-19
C5095 DVDD.n4649 DVSS 9.8e-19
C5096 DVDD.n4650 DVSS 0.001161f
C5097 DVDD.n4652 DVSS 0.001161f
C5098 DVDD.n4653 DVSS 0.001161f
C5099 DVDD.n4654 DVSS 9.8e-19
C5100 DVDD.n4655 DVSS 9.8e-19
C5101 DVDD.n4656 DVSS 9.8e-19
C5102 DVDD.n4657 DVSS 0.001161f
C5103 DVDD.n4659 DVSS 0.001161f
C5104 DVDD.n4660 DVSS 0.001161f
C5105 DVDD.n4661 DVSS 9.8e-19
C5106 DVDD.n4662 DVSS 9.8e-19
C5107 DVDD.n4663 DVSS 9.8e-19
C5108 DVDD.n4664 DVSS 0.001161f
C5109 DVDD.n4666 DVSS 0.001161f
C5110 DVDD.n4667 DVSS 0.001161f
C5111 DVDD.n4668 DVSS 9.8e-19
C5112 DVDD.n4669 DVSS 9.8e-19
C5113 DVDD.n4670 DVSS 9.8e-19
C5114 DVDD.n4671 DVSS 0.001161f
C5115 DVDD.n4673 DVSS 0.001161f
C5116 DVDD.n4674 DVSS 0.001161f
C5117 DVDD.n4675 DVSS 9.8e-19
C5118 DVDD.n4676 DVSS 9.8e-19
C5119 DVDD.n4677 DVSS 9.8e-19
C5120 DVDD.n4678 DVSS 0.001161f
C5121 DVDD.n4680 DVSS 0.001161f
C5122 DVDD.n4681 DVSS 0.001161f
C5123 DVDD.n4682 DVSS 9.24e-19
C5124 DVDD.n4683 DVSS 4.9e-19
C5125 DVDD.n4684 DVSS 0.001538f
C5126 DVDD.n4685 DVSS 0.001563f
C5127 DVDD.n4686 DVSS 0.001538f
C5128 DVDD.n4687 DVSS 0.003076f
C5129 DVDD.n4688 DVSS 0.003076f
C5130 DVDD.n4689 DVSS 0.001538f
C5131 DVDD.n4690 DVSS 0.025852f
C5132 DVDD.n4691 DVSS 0.025852f
C5133 DVDD.n4692 DVSS 0.003076f
C5134 DVDD.n4693 DVSS 0.003076f
C5135 DVDD.n4694 DVSS 0.024004f
C5136 DVDD.n4695 DVSS 0.023073f
C5137 DVDD.n4696 DVSS 0.052845f
C5138 DVDD.n4697 DVSS 0.050332f
C5139 DVDD.n4698 DVSS 0.150127f
C5140 DVDD.n4699 DVSS 0.052845f
C5141 DVDD.n4700 DVSS 0.052845f
C5142 DVDD.n4701 DVSS 0.023073f
C5143 DVDD.n4702 DVSS 0.023073f
C5144 DVDD.n4703 DVSS 0.026423f
C5145 DVDD.n4704 DVSS 0.003076f
C5146 DVDD.n4705 DVSS 0.003076f
C5147 DVDD.n4706 DVSS 0.003076f
C5148 DVDD.n4707 DVSS 0.026423f
C5149 DVDD.n4708 DVSS 0.023073f
C5150 DVDD.n4709 DVSS 0.052845f
C5151 DVDD.n4710 DVSS 0.052845f
C5152 DVDD.n4711 DVSS 0.052845f
C5153 DVDD.n4712 DVSS 0.052845f
C5154 DVDD.n4713 DVSS 0.023073f
C5155 DVDD.n4714 DVSS 0.026423f
C5156 DVDD.n4715 DVSS 0.003076f
C5157 DVDD.n4716 DVSS 0.003076f
C5158 DVDD.n4717 DVSS 0.023631f
C5159 DVDD.n4718 DVSS 0.025864f
C5160 DVDD.n4719 DVSS 0.064196f
C5161 DVDD.n4720 DVSS 0.087827f
C5162 DVDD.n4721 DVSS 0.087827f
C5163 DVDD.n4722 DVSS 0.087827f
C5164 DVDD.n4723 DVSS 0.03889f
C5165 DVDD.n4724 DVSS 0.023073f
C5166 DVDD.n4725 DVSS 0.026423f
C5167 DVDD.n4726 DVSS 0.003076f
C5168 DVDD.n4727 DVSS 0.003076f
C5169 DVDD.n4728 DVSS 0.003076f
C5170 DVDD.n4729 DVSS 0.026423f
C5171 DVDD.n4730 DVSS 0.023073f
C5172 DVDD.n4731 DVSS 0.052845f
C5173 DVDD.n4732 DVSS 0.052845f
C5174 DVDD.n4733 DVSS 0.052845f
C5175 DVDD.n4734 DVSS 0.052845f
C5176 DVDD.n4735 DVSS 0.052845f
C5177 DVDD.n4736 DVSS 0.023073f
C5178 DVDD.n4737 DVSS 0.023631f
C5179 DVDD.n4738 DVSS 0.025864f
C5180 DVDD.n4739 DVSS 0.005483f
C5181 DVDD.n4740 DVSS 0.004466f
C5182 DVDD.n4741 DVSS 4.9e-19
C5183 DVDD.n4742 DVSS 5.28e-19
C5184 DVDD.n4743 DVSS 0.001161f
C5185 DVDD.n4744 DVSS 0.001161f
C5186 DVDD.n4745 DVSS 9.8e-19
C5187 DVDD.n4746 DVSS 9.8e-19
C5188 DVDD.n4747 DVSS 0.001161f
C5189 DVDD.n4748 DVSS 0.001161f
C5190 DVDD.n4749 DVSS 9.8e-19
C5191 DVDD.n4750 DVSS 9.8e-19
C5192 DVDD.n4751 DVSS 0.001161f
C5193 DVDD.n4752 DVSS 0.001161f
C5194 DVDD.n4753 DVSS 9.8e-19
C5195 DVDD.n4754 DVSS 9.8e-19
C5196 DVDD.n4755 DVSS 0.001161f
C5197 DVDD.n4756 DVSS 0.001161f
C5198 DVDD.n4757 DVSS 9.8e-19
C5199 DVDD.n4758 DVSS 9.8e-19
C5200 DVDD.n4759 DVSS 0.001161f
C5201 DVDD.n4760 DVSS 0.001161f
C5202 DVDD.n4761 DVSS 9.8e-19
C5203 DVDD.n4762 DVSS 9.8e-19
C5204 DVDD.n4763 DVSS 0.001161f
C5205 DVDD.n4764 DVSS 0.001161f
C5206 DVDD.n4765 DVSS 9.8e-19
C5207 DVDD.n4766 DVSS 9.8e-19
C5208 DVDD.n4767 DVSS 0.001161f
C5209 DVDD.n4768 DVSS 0.001161f
C5210 DVDD.n4769 DVSS 9.8e-19
C5211 DVDD.n4770 DVSS 9.8e-19
C5212 DVDD.n4771 DVSS 0.001161f
C5213 DVDD.n4772 DVSS 0.001161f
C5214 DVDD.n4773 DVSS 9.8e-19
C5215 DVDD.n4774 DVSS 9.8e-19
C5216 DVDD.n4775 DVSS 0.001161f
C5217 DVDD.n4776 DVSS 0.001161f
C5218 DVDD.n4777 DVSS 9.8e-19
C5219 DVDD.n4778 DVSS 9.8e-19
C5220 DVDD.n4779 DVSS 0.001161f
C5221 DVDD.n4780 DVSS 0.001161f
C5222 DVDD.n4781 DVSS 9.8e-19
C5223 DVDD.n4782 DVSS 9.8e-19
C5224 DVDD.n4783 DVSS 0.001161f
C5225 DVDD.n4784 DVSS 0.001161f
C5226 DVDD.n4785 DVSS 8.2e-19
C5227 DVDD.n4786 DVSS 4.9e-19
C5228 DVDD.n4787 DVSS 0.003076f
C5229 DVDD.n4788 DVSS 0.064196f
C5230 DVDD.n4789 DVSS 0.064196f
C5231 DVDD.n4790 DVSS 0.026423f
C5232 DVDD.n4791 DVSS 0.087827f
C5233 DVDD.n4792 DVSS 0.087827f
C5234 DVDD.n4793 DVSS 0.087827f
C5235 DVDD.n4794 DVSS 0.052845f
C5236 DVDD.n4795 DVSS 0.052845f
C5237 DVDD.n4796 DVSS 0.03889f
C5238 DVDD.n4797 DVSS 0.052845f
C5239 DVDD.n4798 DVSS 0.052845f
C5240 DVDD.n4799 DVSS 0.023073f
C5241 DVDD.n4800 DVSS 0.003076f
C5242 DVDD.n4801 DVSS 0.026423f
C5243 DVDD.n4802 DVSS 0.003076f
C5244 DVDD.n4803 DVSS 0.003076f
C5245 DVDD.n4804 DVSS 0.026423f
C5246 DVDD.n4805 DVSS 0.023073f
C5247 DVDD.n4806 DVSS 0.052845f
C5248 DVDD.n4807 DVSS 0.052845f
C5249 DVDD.n4808 DVSS 0.023073f
C5250 DVDD.n4809 DVSS 0.023631f
C5251 DVDD.n4810 DVSS 0.025864f
C5252 DVDD.n4811 DVSS 0.005483f
C5253 DVDD.n4812 DVSS 0.001161f
C5254 DVDD.n4813 DVSS 9.8e-19
C5255 DVDD.n4814 DVSS 9.8e-19
C5256 DVDD.n4815 DVSS 0.001161f
C5257 DVDD.n4816 DVSS 0.001161f
C5258 DVDD.n4817 DVSS 9.8e-19
C5259 DVDD.n4818 DVSS 9.8e-19
C5260 DVDD.n4819 DVSS 0.001161f
C5261 DVDD.n4820 DVSS 0.001161f
C5262 DVDD.n4821 DVSS 9.8e-19
C5263 DVDD.n4822 DVSS 9.8e-19
C5264 DVDD.n4823 DVSS 0.001161f
C5265 DVDD.n4824 DVSS 0.001161f
C5266 DVDD.n4825 DVSS 9.8e-19
C5267 DVDD.n4826 DVSS 9.8e-19
C5268 DVDD.n4827 DVSS 0.001161f
C5269 DVDD.n4828 DVSS 0.001161f
C5270 DVDD.n4829 DVSS 9.8e-19
C5271 DVDD.n4830 DVSS 9.8e-19
C5272 DVDD.n4831 DVSS 0.001161f
C5273 DVDD.n4832 DVSS 0.001161f
C5274 DVDD.n4833 DVSS 9.8e-19
C5275 DVDD.n4834 DVSS 9.8e-19
C5276 DVDD.n4835 DVSS 0.001161f
C5277 DVDD.n4836 DVSS 0.001161f
C5278 DVDD.n4837 DVSS 9.8e-19
C5279 DVDD.n4838 DVSS 9.8e-19
C5280 DVDD.n4839 DVSS 0.001161f
C5281 DVDD.n4840 DVSS 0.001161f
C5282 DVDD.n4841 DVSS 9.8e-19
C5283 DVDD.n4842 DVSS 6.32e-19
C5284 DVDD.n4843 DVSS 0.001161f
C5285 DVDD.n4844 DVSS 0.001161f
C5286 DVDD.n4845 DVSS 5.09e-19
C5287 DVDD.n4846 DVSS 4.9e-19
C5288 DVDD.n4847 DVSS 0.004466f
C5289 DVDD.n4848 DVSS 0.002059f
C5290 DVDD.n4849 DVSS 0.003076f
C5291 DVDD.n4850 DVSS 0.023631f
C5292 DVDD.n4851 DVSS 0.023073f
C5293 DVDD.n4852 DVSS 0.052845f
C5294 DVDD.n4853 DVSS 0.052845f
C5295 DVDD.n4854 DVSS 0.023073f
C5296 DVDD.n4855 DVSS 0.026423f
C5297 DVDD.n4856 DVSS 0.003076f
C5298 DVDD.n4857 DVSS 0.003076f
C5299 DVDD.n4858 DVSS 0.026423f
C5300 DVDD.n4859 DVSS 0.023073f
C5301 DVDD.n4860 DVSS 0.03889f
C5302 DVDD.n4861 DVSS 0.204821f
C5303 DVDD.n4862 DVSS 0.031765f
C5304 DVDD.n4863 DVSS 0.463259f
C5305 DVDD.n4864 DVSS 0.03889f
C5306 DVDD.n4865 DVSS 0.052845f
C5307 DVDD.n4866 DVSS 0.052845f
C5308 DVDD.n4867 DVSS 0.052845f
C5309 DVDD.n4868 DVSS 0.052845f
C5310 DVDD.n4869 DVSS 0.023073f
C5311 DVDD.n4870 DVSS 0.026423f
C5312 DVDD.n4871 DVSS 0.003076f
C5313 DVDD.n4872 DVSS 0.003076f
C5314 DVDD.n4873 DVSS 0.003076f
C5315 DVDD.n4874 DVSS 0.023073f
C5316 DVDD.n4875 DVSS 0.026423f
C5317 DVDD.n4876 DVSS 0.008245f
C5318 DVDD.n4877 DVSS 0.003523f
C5319 DVDD.n4878 DVSS 0.003076f
C5320 DVDD.n4879 DVSS 0.007046f
C5321 DVDD.n4880 DVSS 0.020366f
C5322 DVDD.n4881 DVSS 0.007156f
C5323 DVDD.n4882 DVSS 0.007112f
C5324 DVDD.n4883 DVSS 0.005519f
C5325 DVDD.n4884 DVSS 0.025864f
C5326 DVDD.n4885 DVSS 0.064196f
C5327 DVDD.n4886 DVSS 0.087827f
C5328 DVDD.n4887 DVSS 0.087827f
C5329 DVDD.n4888 DVSS 0.087827f
C5330 DVDD.n4889 DVSS 0.052845f
C5331 DVDD.n4890 DVSS 0.03889f
C5332 DVDD.n4891 DVSS 0.052845f
C5333 DVDD.n4892 DVSS 0.052845f
C5334 DVDD.n4893 DVSS 0.052845f
C5335 DVDD.n4894 DVSS 0.023073f
C5336 DVDD.n4895 DVSS 0.026423f
C5337 DVDD.n4896 DVSS 0.003076f
C5338 DVDD.n4897 DVSS 0.003076f
C5339 DVDD.n4898 DVSS 0.026423f
C5340 DVDD.n4899 DVSS 0.003523f
C5341 DVDD.n4900 DVSS 0.003076f
C5342 DVDD.n4901 DVSS 0.003523f
C5343 DVDD.n4902 DVSS 0.008245f
C5344 DVDD.n4903 DVSS 0.026423f
C5345 DVDD.n4904 DVSS 0.008245f
C5346 DVDD.n4905 DVSS 0.003523f
C5347 DVDD.n4906 DVSS 0.007046f
C5348 DVDD.n4907 DVSS 0.005384f
C5349 DVDD.n4908 DVSS 0.00698f
C5350 DVDD.n4909 DVSS 0.003076f
C5351 DVDD.n4910 DVSS 0.003399f
C5352 DVDD.n4911 DVSS 0.008245f
C5353 DVDD.n4912 DVSS 0.024004f
C5354 DVDD.n4913 DVSS 0.026423f
C5355 DVDD.n4914 DVSS 0.026423f
C5356 DVDD.n4915 DVSS 0.008245f
C5357 DVDD.n4916 DVSS 0.006751f
C5358 DVDD.n4917 DVSS 0.0032f
C5359 DVDD.n4918 DVSS 0.003076f
C5360 DVDD.n4919 DVSS 0.003076f
C5361 DVDD.n4920 DVSS 0.003523f
C5362 DVDD.n4921 DVSS 0.008245f
C5363 DVDD.n4922 DVSS 0.026423f
C5364 DVDD.n4923 DVSS 0.026423f
C5365 DVDD.n4924 DVSS 0.008245f
C5366 DVDD.n4925 DVSS 0.003076f
C5367 DVDD.n4926 DVSS 0.003523f
C5368 DVDD.n4927 DVSS 0.005185f
C5369 DVDD.n4928 DVSS 0.007046f
C5370 DVDD.n4929 DVSS 0.007112f
C5371 DVDD.n4930 DVSS 0.003076f
C5372 DVDD.n4931 DVSS 0.003523f
C5373 DVDD.n4932 DVSS 0.008245f
C5374 DVDD.n4933 DVSS 0.023631f
C5375 DVDD.n4934 DVSS 0.053408f
C5376 DVDD.n4936 DVSS 0.026423f
C5377 DVDD.n4937 DVSS 0.024376f
C5378 DVDD.n4938 DVSS 0.031819f
C5379 DVDD.n4939 DVSS 0.008245f
C5380 DVDD.n4940 DVSS 0.008245f
C5381 DVDD.n4941 DVSS 0.008245f
C5382 DVDD.n4942 DVSS 0.008245f
C5383 DVDD.n4943 DVSS 0.008245f
C5384 DVDD.n4944 DVSS 0.008245f
C5385 DVDD.n4945 DVSS 0.008245f
C5386 DVDD.n4946 DVSS 0.008245f
C5387 DVDD.n4947 DVSS 0.008245f
C5388 DVDD.n4948 DVSS 0.008245f
C5389 DVDD.n4949 DVSS 0.008245f
C5390 DVDD.n4950 DVSS 0.052845f
C5391 DVDD.n4951 DVSS 0.052845f
C5392 DVDD.n4952 DVSS 0.052845f
C5393 DVDD.n4953 DVSS 0.052845f
C5394 DVDD.n4954 DVSS 0.052845f
C5395 DVDD.n4955 DVSS 0.052845f
C5396 DVDD.n4956 DVSS 0.052845f
C5397 DVDD.n4957 DVSS 0.052845f
C5398 DVDD.n4958 DVSS 0.052845f
C5399 DVDD.n4959 DVSS 0.045402f
C5400 DVDD.n4960 DVSS 0.045402f
C5401 DVDD.n4961 DVSS 0.052845f
C5402 DVDD.n4962 DVSS 0.052845f
C5403 DVDD.n4963 DVSS 0.052845f
C5404 DVDD.n4964 DVSS 0.052845f
C5405 DVDD.n4965 DVSS 0.052845f
C5406 DVDD.n4966 DVSS 0.052845f
C5407 DVDD.n4967 DVSS 0.052845f
C5408 DVDD.n4968 DVSS 0.052845f
C5409 DVDD.n4969 DVSS 0.052845f
C5410 DVDD.n4970 DVSS 0.052845f
C5411 DVDD.n4971 DVSS 0.052845f
C5412 DVDD.n4972 DVSS 0.052845f
C5413 DVDD.n4973 DVSS 0.052845f
C5414 DVDD.n4974 DVSS 0.052845f
C5415 DVDD.n4975 DVSS 0.052845f
C5416 DVDD.n4976 DVSS 0.052845f
C5417 DVDD.n4977 DVSS 0.052845f
C5418 DVDD.n4978 DVSS 0.052845f
C5419 DVDD.n4979 DVSS 0.052845f
C5420 DVDD.n4980 DVSS 0.052845f
C5421 DVDD.n4981 DVSS 0.052845f
C5422 DVDD.n4982 DVSS 0.052845f
C5423 DVDD.n4983 DVSS 0.052845f
C5424 DVDD.n4984 DVSS 0.052845f
C5425 DVDD.n4985 DVSS 0.052845f
C5426 DVDD.n4986 DVSS 0.052845f
C5427 DVDD.n4987 DVSS 0.052845f
C5428 DVDD.n4988 DVSS 0.052845f
C5429 DVDD.n4989 DVSS 0.052845f
C5430 DVDD.n4990 DVSS 0.052845f
C5431 DVDD.n4991 DVSS 0.052845f
C5432 DVDD.n4992 DVSS 0.052845f
C5433 DVDD.n4993 DVSS 0.052845f
C5434 DVDD.n4994 DVSS 0.052845f
C5435 DVDD.n4995 DVSS 0.052845f
C5436 DVDD.n4996 DVSS 0.052845f
C5437 DVDD.n4997 DVSS 0.040514f
C5438 DVDD.n4998 DVSS 0.052845f
C5439 DVDD.n4999 DVSS 0.032377f
C5440 DVDD.n5000 DVSS 0.017268f
C5441 DVDD.n5001 DVSS 0.025008f
C5442 DVDD.n5002 DVSS 0.028184f
C5443 DVDD.n5003 DVSS 0.028184f
C5444 DVDD.n5004 DVSS 0.028184f
C5445 DVDD.n5005 DVSS 0.028184f
C5446 DVDD.n5006 DVSS 0.028184f
C5447 DVDD.n5007 DVSS 0.028184f
C5448 DVDD.n5008 DVSS 0.028184f
C5449 DVDD.n5009 DVSS 0.028184f
C5450 DVDD.n5010 DVSS 0.018855f
C5451 DVDD.n5011 DVSS 0.007046f
C5452 DVDD.n5012 DVSS 0.007156f
C5453 DVDD.n5013 DVSS 0.007046f
C5454 DVDD.n5014 DVSS 0.003523f
C5455 DVDD.n5015 DVSS 0.003076f
C5456 DVDD.n5017 DVSS 0.008478f
C5457 DVDD.n5018 DVSS 0.007112f
C5458 DVDD.n5019 DVSS 0.003076f
C5459 DVDD.n5020 DVSS 0.003151f
C5460 DVDD.n5021 DVSS 0.008245f
C5461 DVDD.n5022 DVSS 0.008245f
C5462 DVDD.n5024 DVSS 0.003523f
C5463 DVDD.n5025 DVSS 0.008245f
C5464 DVDD.n5026 DVSS 0.008245f
C5465 DVDD.n5027 DVSS 0.003523f
C5466 DVDD.n5028 DVSS 0.003076f
C5467 DVDD.n5029 DVSS 0.007046f
C5468 DVDD.n5030 DVSS 0.020366f
C5469 DVDD.n5031 DVSS 0.007046f
C5470 DVDD.n5032 DVSS 0.020195f
C5471 DVDD.n5033 DVSS 0.005185f
C5472 DVDD.n5034 DVSS 0.005185f
C5473 DVDD.n5035 DVSS 0.020195f
C5474 DVDD.n5036 DVSS 0.018855f
C5475 DVDD.n5037 DVSS 0.016573f
C5476 DVDD.n5038 DVSS 0.028184f
C5477 DVDD.n5039 DVSS 0.028184f
C5478 DVDD.n5040 DVSS 0.028184f
C5479 DVDD.n5041 DVSS 0.028184f
C5480 DVDD.n5042 DVSS 0.028184f
C5481 DVDD.n5043 DVSS 0.028184f
C5482 DVDD.n5044 DVSS 0.028184f
C5483 DVDD.n5045 DVSS 0.028184f
C5484 DVDD.n5046 DVSS 0.028184f
C5485 DVDD.n5047 DVSS 0.028184f
C5486 DVDD.n5048 DVSS 0.028184f
C5487 DVDD.n5049 DVSS 0.028184f
C5488 DVDD.n5050 DVSS 0.028184f
C5489 DVDD.n5051 DVSS 0.028184f
C5490 DVDD.n5052 DVSS 0.028184f
C5491 DVDD.n5053 DVSS 0.028184f
C5492 DVDD.n5054 DVSS 0.017268f
C5493 DVDD.n5055 DVSS 0.028184f
C5494 DVDD.n5056 DVSS 0.028184f
C5495 DVDD.n5057 DVSS 0.028184f
C5496 DVDD.n5058 DVSS 0.017268f
C5497 DVDD.n5059 DVSS 0.028184f
C5498 DVDD.n5060 DVSS 0.028184f
C5499 DVDD.n5061 DVSS 0.025008f
C5500 DVDD.n5062 DVSS 0.028184f
C5501 DVDD.n5063 DVSS 0.028184f
C5502 DVDD.n5064 DVSS 0.028184f
C5503 DVDD.n5065 DVSS 0.028184f
C5504 DVDD.n5066 DVSS 0.028184f
C5505 DVDD.n5067 DVSS 0.028184f
C5506 DVDD.n5068 DVSS 0.028184f
C5507 DVDD.n5069 DVSS 0.025008f
C5508 DVDD.n5070 DVSS 0.040514f
C5509 DVDD.n5071 DVSS 0.046891f
C5510 DVDD.n5072 DVSS 0.052845f
C5511 DVDD.n5073 DVSS 0.052845f
C5512 DVDD.n5074 DVSS 0.052845f
C5513 DVDD.n5075 DVSS 0.052845f
C5514 DVDD.n5076 DVSS 0.052845f
C5515 DVDD.n5077 DVSS 0.052845f
C5516 DVDD.n5078 DVSS 0.052845f
C5517 DVDD.n5079 DVSS 0.003076f
C5518 DVDD.n5080 DVSS 0.023073f
C5519 DVDD.n5081 DVSS 0.052845f
C5520 DVDD.n5082 DVSS 0.023073f
C5521 DVDD.n5083 DVSS 0.040378f
C5522 DVDD.n5084 DVSS 0.08485f
C5523 DVDD.n5085 DVSS 0.08485f
C5524 DVDD.n5086 DVSS 0.003076f
C5525 DVDD.n5087 DVSS 0.003076f
C5526 DVDD.n5088 DVSS 0.026423f
C5527 DVDD.n5089 DVSS 0.023073f
C5528 DVDD.n5090 DVSS 0.052845f
C5529 DVDD.n5091 DVSS 0.023073f
C5530 DVDD.n5092 DVSS 0.052845f
C5531 DVDD.n5093 DVSS 0.040378f
C5532 DVDD.n5094 DVSS 0.052845f
C5533 DVDD.n5095 DVSS 0.062707f
C5534 DVDD.n5096 DVSS 0.062707f
C5535 DVDD.n5097 DVSS 0.08485f
C5536 DVDD.n5098 DVSS 0.08485f
C5537 DVDD.n5099 DVSS 0.052845f
C5538 DVDD.n5100 DVSS 0.052845f
C5539 DVDD.n5101 DVSS 0.052845f
C5540 DVDD.n5102 DVSS 0.023073f
C5541 DVDD.n5103 DVSS 0.025492f
C5542 DVDD.n5104 DVSS 0.003076f
C5543 DVDD.n5105 DVSS 0.003076f
C5544 DVDD.n5106 DVSS 0.006004f
C5545 DVDD.n5107 DVSS 0.006004f
C5546 DVDD.n5108 DVSS 0.003076f
C5547 DVDD.n5109 DVSS 0.003399f
C5548 DVDD.n5110 DVSS 0.008245f
C5549 DVDD.n5111 DVSS 0.025492f
C5550 DVDD.n5112 DVSS 0.024004f
C5551 DVDD.n5113 DVSS 0.023073f
C5552 DVDD.n5114 DVSS 0.052845f
C5553 DVDD.n5115 DVSS 0.052845f
C5554 DVDD.n5116 DVSS 0.052845f
C5555 DVDD.n5117 DVSS 0.052845f
C5556 DVDD.n5118 DVSS 0.052845f
C5557 DVDD.n5119 DVSS 0.023073f
C5558 DVDD.n5120 DVSS 0.026423f
C5559 DVDD.n5121 DVSS 0.003076f
C5560 DVDD.n5122 DVSS 0.003076f
C5561 DVDD.n5123 DVSS 0.003076f
C5562 DVDD.n5124 DVSS 0.003076f
C5563 DVDD.n5125 DVSS 0.003076f
C5564 DVDD.n5126 DVSS 0.023073f
C5565 DVDD.n5127 DVSS 0.052845f
C5566 DVDD.n5128 DVSS 0.023073f
C5567 DVDD.n5129 DVSS 0.03889f
C5568 DVDD.n5130 DVSS 0.026423f
C5569 DVDD.n5131 DVSS 0.023073f
C5570 DVDD.n5132 DVSS 0.052845f
C5571 DVDD.n5133 DVSS 0.052845f
C5572 DVDD.n5134 DVSS 0.152989f
C5573 DVDD.n5135 DVSS 0.053362f
C5574 DVDD.n5136 DVSS 0.052845f
C5575 DVDD.n5137 DVSS 0.023073f
C5576 DVDD.n5138 DVSS 0.026423f
C5577 DVDD.n5139 DVSS 0.003076f
C5578 DVDD.n5140 DVSS 0.003076f
C5579 DVDD.n5141 DVSS 0.085321f
C5580 DVDD.n5142 DVSS 0.085321f
C5581 DVDD.n5143 DVSS 0.023073f
C5582 DVDD.n5144 DVSS 0.003076f
C5583 DVDD.n5145 DVSS 0.003076f
C5584 DVDD.n5146 DVSS 0.003076f
C5585 DVDD.n5147 DVSS 0.003076f
C5586 DVDD.n5148 DVSS 0.003076f
C5587 DVDD.n5149 DVSS 0.003076f
C5588 DVDD.n5150 DVSS 0.003076f
C5589 DVDD.n5151 DVSS 0.003076f
C5590 DVDD.n5152 DVSS 0.003076f
C5591 DVDD.n5153 DVSS 0.003076f
C5592 DVDD.n5154 DVSS 0.001538f
C5593 DVDD.n5155 DVSS 0.052845f
C5594 DVDD.n5156 DVSS 0.052845f
C5595 DVDD.n5157 DVSS 0.052845f
C5596 DVDD.n5158 DVSS 0.052845f
C5597 DVDD.n5159 DVSS 0.052845f
C5598 DVDD.n5160 DVSS 0.052845f
C5599 DVDD.n5161 DVSS 0.052845f
C5600 DVDD.n5162 DVSS 0.052845f
C5601 DVDD.n5163 DVSS 0.052845f
C5602 DVDD.n5164 DVSS 0.052845f
C5603 DVDD.n5165 DVSS 0.052845f
C5604 DVDD.n5166 DVSS 0.052845f
C5605 DVDD.n5167 DVSS 0.052845f
C5606 DVDD.n5168 DVSS 0.052845f
C5607 DVDD.n5169 DVSS 0.052845f
C5608 DVDD.n5170 DVSS 0.052845f
C5609 DVDD.n5171 DVSS 0.052845f
C5610 DVDD.n5172 DVSS 0.052845f
C5611 DVDD.n5173 DVSS 0.052845f
C5612 DVDD.n5174 DVSS 0.052845f
C5613 DVDD.n5175 DVSS 0.052845f
C5614 DVDD.n5176 DVSS 0.052845f
C5615 DVDD.n5177 DVSS 0.052845f
C5616 DVDD.n5178 DVSS 0.052845f
C5617 DVDD.n5179 DVSS 0.052845f
C5618 DVDD.n5180 DVSS 0.052845f
C5619 DVDD.n5181 DVSS 0.052845f
C5620 DVDD.n5182 DVSS 0.052845f
C5621 DVDD.n5183 DVSS 0.052845f
C5622 DVDD.n5184 DVSS 0.052845f
C5623 DVDD.n5185 DVSS 0.052845f
C5624 DVDD.n5186 DVSS 0.052845f
C5625 DVDD.n5187 DVSS 0.052845f
C5626 DVDD.n5188 DVSS 0.052845f
C5627 DVDD.n5189 DVSS 0.052845f
C5628 DVDD.n5190 DVSS 0.052845f
C5629 DVDD.n5191 DVSS 0.052845f
C5630 DVDD.n5192 DVSS 0.052845f
C5631 DVDD.n5193 DVSS 0.052845f
C5632 DVDD.n5194 DVSS 0.052845f
C5633 DVDD.n5195 DVSS 0.052845f
C5634 DVDD.n5196 DVSS 0.052845f
C5635 DVDD.n5197 DVSS 0.052845f
C5636 DVDD.n5198 DVSS 0.052845f
C5637 DVDD.n5199 DVSS 0.052845f
C5638 DVDD.n5200 DVSS 0.052845f
C5639 DVDD.n5201 DVSS 0.031074f
C5640 DVDD.n5202 DVSS 0.001538f
C5641 DVDD.n5203 DVSS 0.003076f
C5642 DVDD.n5204 DVSS 0.003076f
C5643 DVDD.n5205 DVSS 0.003076f
C5644 DVDD.n5206 DVSS 0.003076f
C5645 DVDD.n5207 DVSS 0.003076f
C5646 DVDD.n5208 DVSS 0.003076f
C5647 DVDD.n5209 DVSS 0.003076f
C5648 DVDD.n5210 DVSS 0.003076f
C5649 DVDD.n5211 DVSS 0.003076f
C5650 DVDD.n5212 DVSS 0.026423f
C5651 DVDD.n5213 DVSS 0.003076f
C5652 DVDD.n5214 DVSS 0.003076f
C5653 DVDD.n5215 DVSS 0.026423f
C5654 DVDD.n5216 DVSS 0.051543f
C5655 DVDD.n5217 DVSS 0.052845f
C5656 DVDD.n5218 DVSS 0.052845f
C5657 DVDD.n5219 DVSS 0.052845f
C5658 DVDD.n5220 DVSS 0.052845f
C5659 DVDD.n5221 DVSS 0.052845f
C5660 DVDD.n5222 DVSS 0.046891f
C5661 DVDD.n5223 DVSS 0.046891f
C5662 DVDD.n5224 DVSS 0.040514f
C5663 DVDD.n5225 DVSS 0.032377f
C5664 DVDD.n5226 DVSS 0.032377f
C5665 DVDD.n5227 DVSS 0.052845f
C5666 DVDD.n5228 DVSS 0.052845f
C5667 DVDD.n5229 DVSS 0.052845f
C5668 DVDD.n5230 DVSS 0.052845f
C5669 DVDD.n5231 DVSS 0.052845f
C5670 DVDD.n5232 DVSS 0.052845f
C5671 DVDD.n5233 DVSS 0.052845f
C5672 DVDD.n5234 DVSS 0.052845f
C5673 DVDD.n5235 DVSS 0.052845f
C5674 DVDD.n5236 DVSS 0.052845f
C5675 DVDD.n5237 DVSS 0.052845f
C5676 DVDD.n5238 DVSS 0.052845f
C5677 DVDD.n5239 DVSS 0.052845f
C5678 DVDD.n5240 DVSS 0.031074f
C5679 DVDD.n5241 DVSS 0.052845f
C5680 DVDD.n5242 DVSS 0.023073f
C5681 DVDD.n5243 DVSS 0.052845f
C5682 DVDD.n5244 DVSS 0.052845f
C5683 DVDD.n5245 DVSS 0.023073f
C5684 DVDD.n5247 DVSS 0.008245f
C5685 DVDD.n5249 DVSS 0.008245f
C5686 DVDD.n5251 DVSS 0.008245f
C5687 DVDD.n5253 DVSS 0.008245f
C5688 DVDD.n5255 DVSS 0.008245f
C5689 DVDD.n5257 DVSS 0.008245f
C5690 DVDD.n5259 DVSS 0.008245f
C5691 DVDD.n5261 DVSS 0.008245f
C5692 DVDD.n5263 DVSS 0.008245f
C5693 DVDD.n5265 DVSS 0.008245f
C5694 DVDD.n5267 DVSS 0.008245f
C5695 DVDD.n5278 DVSS 0.02512f
C5696 DVDD.n5280 DVSS 0.011536f
C5697 DVDD.n5281 DVSS 0.026423f
C5698 DVDD.n5282 DVSS 0.228661f
C5699 DVDD.n5283 DVSS 0.228661f
C5700 DVDD.n5284 DVSS 0.008245f
C5701 DVDD.n5285 DVSS 0.003151f
C5702 DVDD.n5286 DVSS 0.003076f
C5703 DVDD.n5287 DVSS 0.007046f
C5704 DVDD.n5288 DVSS 0.007156f
C5705 DVDD.n5289 DVSS 0.020366f
C5706 DVDD.n5290 DVSS 0.007046f
C5707 DVDD.n5291 DVSS 0.007046f
C5708 DVDD.n5292 DVSS 0.003076f
C5709 DVDD.n5293 DVSS 0.003523f
C5710 DVDD.n5294 DVSS 0.008245f
C5711 DVDD.n5295 DVSS 0.008245f
C5712 DVDD.n5296 DVSS 0.008245f
C5713 DVDD.n5297 DVSS 0.003523f
C5714 DVDD.n5298 DVSS 0.003076f
C5715 DVDD.n5299 DVSS 0.005384f
C5716 DVDD.n5300 DVSS 0.007046f
C5717 DVDD.n5301 DVSS 0.007046f
C5718 DVDD.n5302 DVSS 0.019986f
C5719 DVDD.n5303 DVSS 0.007046f
C5720 DVDD.n5304 DVSS 0.007046f
C5721 DVDD.n5305 DVSS 0.003076f
C5722 DVDD.n5306 DVSS 0.00698f
C5723 DVDD.n5307 DVSS 0.016091f
C5724 DVDD.n5308 DVSS 0.016091f
C5725 DVDD.n5309 DVSS 0.008245f
C5726 DVDD.n5310 DVSS 0.0032f
C5727 DVDD.n5311 DVSS 0.003076f
C5728 DVDD.n5312 DVSS 0.007046f
C5729 DVDD.n5313 DVSS 0.006751f
C5730 DVDD.n5314 DVSS 0.019986f
C5731 DVDD.n5315 DVSS 0.007046f
C5732 DVDD.n5316 DVSS 0.007046f
C5733 DVDD.n5317 DVSS 0.003076f
C5734 DVDD.n5318 DVSS 0.003523f
C5735 DVDD.n5319 DVSS 0.008245f
C5736 DVDD.n5320 DVSS 0.008245f
C5737 DVDD.n5321 DVSS 0.449908f
C5738 DVDD.n5322 DVSS 0.023073f
C5739 DVDD.n5323 DVSS 0.023073f
C5740 DVDD.n5324 DVSS 0.026423f
C5741 DVDD.n5325 DVSS 0.003076f
C5742 DVDD.n5326 DVSS 0.003076f
C5743 DVDD.n5327 DVSS 0.003076f
C5744 DVDD.n5328 DVSS 0.025492f
C5745 DVDD.n5329 DVSS 0.023073f
C5746 DVDD.n5330 DVSS 0.052845f
C5747 DVDD.n5331 DVSS 0.052845f
C5748 DVDD.n5332 DVSS 0.052845f
C5749 DVDD.n5333 DVSS 0.08485f
C5750 DVDD.n5334 DVSS 0.08485f
C5751 DVDD.n5335 DVSS 0.062707f
C5752 DVDD.n5336 DVSS 0.026423f
C5753 DVDD.n5337 DVSS 0.006004f
C5754 DVDD.n5338 DVSS 0.006004f
C5755 DVDD.n5339 DVSS 0.003076f
C5756 DVDD.n5340 DVSS 0.003076f
C5757 DVDD.n5341 DVSS 0.024004f
C5758 DVDD.n5342 DVSS 0.023073f
C5759 DVDD.n5343 DVSS 0.052845f
C5760 DVDD.n5344 DVSS 0.052845f
C5761 DVDD.n5345 DVSS 0.052845f
C5762 DVDD.n5346 DVSS 0.052845f
C5763 DVDD.n5347 DVSS 0.052845f
C5764 DVDD.n5348 DVSS 0.040378f
C5765 DVDD.n5349 DVSS 0.023073f
C5766 DVDD.n5350 DVSS 0.026423f
C5767 DVDD.n5351 DVSS 0.003076f
C5768 DVDD.n5352 DVSS 0.003076f
C5769 DVDD.n5353 DVSS 0.03889f
C5770 DVDD.n5354 DVSS 0.023073f
C5771 DVDD.n5355 DVSS 0.023073f
C5772 DVDD.n5356 DVSS 0.026423f
C5773 DVDD.n5357 DVSS 0.003076f
C5774 DVDD.n5358 DVSS 0.003076f
C5775 DVDD.n5359 DVSS 0.003076f
C5776 DVDD.n5360 DVSS 0.026423f
C5777 DVDD.n5361 DVSS 0.023073f
C5778 DVDD.n5362 DVSS 0.052845f
C5779 DVDD.n5363 DVSS 0.152989f
C5780 DVDD.n5364 DVSS 0.053362f
C5781 DVDD.n5365 DVSS 0.053408f
C5782 DVDD.n5366 DVSS 0.085321f
C5783 DVDD.n5367 DVSS 0.085321f
C5784 DVDD.n5368 DVSS 0.001538f
C5785 DVDD.n5369 DVSS 0.003076f
C5786 DVDD.n5370 DVSS 0.003076f
C5787 DVDD.n5371 DVSS 0.003076f
C5788 DVDD.n5372 DVSS 0.003076f
C5789 DVDD.n5373 DVSS 0.003076f
C5790 DVDD.n5374 DVSS 0.003076f
C5791 DVDD.n5375 DVSS 0.003076f
C5792 DVDD.n5376 DVSS 0.003076f
C5793 DVDD.n5377 DVSS 0.003076f
C5794 DVDD.n5378 DVSS 0.003076f
C5795 DVDD.n5379 DVSS 0.003076f
C5796 DVDD.n5380 DVSS 0.003076f
C5797 DVDD.n5381 DVSS 0.003076f
C5798 DVDD.n5382 DVSS 0.003076f
C5799 DVDD.n5383 DVSS 0.003076f
C5800 DVDD.n5384 DVSS 0.003076f
C5801 DVDD.n5385 DVSS 0.003076f
C5802 DVDD.n5386 DVSS 0.003076f
C5803 DVDD.n5387 DVSS 0.003076f
C5804 DVDD.n5388 DVSS 0.001538f
C5805 DVDD.n5389 DVSS 0.003076f
C5806 DVDD.n5390 DVSS 0.003076f
C5807 DVDD.n5391 DVSS 0.026423f
C5808 DVDD.n5392 DVSS 0.023073f
C5809 DVDD.n5393 DVSS 0.052845f
C5810 DVDD.n5394 DVSS 0.030888f
C5811 DVDD.n5395 DVSS 0.017305f
C5812 DVDD.n5396 DVSS 0.040514f
C5813 DVDD.n5397 DVSS 0.052845f
C5814 DVDD.n5398 DVSS 0.052845f
C5815 DVDD.n5399 DVSS 0.052845f
C5816 DVDD.n5400 DVSS 0.052845f
C5817 DVDD.n5401 DVSS 0.052845f
C5818 DVDD.n5402 DVSS 0.052845f
C5819 DVDD.n5403 DVSS 0.052845f
C5820 DVDD.n5404 DVSS 0.052845f
C5821 DVDD.n5405 DVSS 0.052845f
C5822 DVDD.n5406 DVSS 0.052845f
C5823 DVDD.n5407 DVSS 0.052845f
C5824 DVDD.n5408 DVSS 0.052845f
C5825 DVDD.n5409 DVSS 0.047635f
C5826 DVDD.n5410 DVSS 0.005954f
C5827 DVDD.n5411 DVSS 0.243482f
C5828 DVDD.n5412 DVSS 0.075079f
C5829 DVDD.n5413 DVSS 0.047635f
C5830 DVDD.n5414 DVSS 0.047635f
C5831 DVDD.n5415 DVSS 0.052845f
C5832 DVDD.n5416 DVSS 0.052845f
C5833 DVDD.n5417 DVSS 0.052845f
C5834 DVDD.n5418 DVSS 0.052845f
C5835 DVDD.n5419 DVSS 0.052845f
C5836 DVDD.n5420 DVSS 0.052845f
C5837 DVDD.n5421 DVSS 0.052845f
C5838 DVDD.n5422 DVSS 0.052845f
C5839 DVDD.n5423 DVSS 0.052845f
C5840 DVDD.n5424 DVSS 0.052845f
C5841 DVDD.n5425 DVSS 0.052845f
C5842 DVDD.n5426 DVSS 0.052845f
C5843 DVDD.n5427 DVSS 0.052845f
C5844 DVDD.n5428 DVSS 0.048379f
C5845 DVDD.n5429 DVSS 0.048379f
C5846 DVDD.n5430 DVSS 0.048379f
C5847 DVDD.n5431 DVSS 0.040514f
C5848 DVDD.n5432 DVSS 0.016474f
C5849 DVDD.n5433 DVSS 0.016474f
C5850 DVDD.n5434 DVSS 0.012306f
C5851 DVDD.n5435 DVSS 0.028184f
C5852 DVDD.n5436 DVSS 0.023123f
C5853 DVDD.n5437 DVSS 0.028184f
C5854 DVDD.n5438 DVSS 0.028184f
C5855 DVDD.n5439 DVSS 0.028184f
C5856 DVDD.n5440 DVSS 0.028184f
C5857 DVDD.n5441 DVSS 0.028184f
C5858 DVDD.n5442 DVSS 0.028184f
C5859 DVDD.n5443 DVSS 0.028184f
C5860 DVDD.n5444 DVSS 0.028184f
C5861 DVDD.n5445 DVSS 0.028184f
C5862 DVDD.n5446 DVSS 0.028184f
C5863 DVDD.n5447 DVSS 0.028184f
C5864 DVDD.n5448 DVSS 0.028184f
C5865 DVDD.n5449 DVSS 0.028184f
C5866 DVDD.n5450 DVSS 0.028184f
C5867 DVDD.n5451 DVSS 0.028184f
C5868 DVDD.n5452 DVSS 0.019649f
C5869 DVDD.n5453 DVSS 0.019649f
C5870 DVDD.n5454 DVSS 0.019649f
C5871 DVDD.n5455 DVSS 0.031815f
C5872 DVDD.n5456 DVSS 0.031917f
C5873 DVDD.n5457 DVSS 0.082136f
C5874 DVDD.n5458 DVSS 0.025207f
C5875 DVDD.n5459 DVSS 0.025207f
C5876 DVDD.n5460 DVSS 0.025207f
C5877 DVDD.n5461 DVSS 0.028184f
C5878 DVDD.n5462 DVSS 0.028184f
C5879 DVDD.n5463 DVSS 0.028184f
C5880 DVDD.n5464 DVSS 0.028184f
C5881 DVDD.n5465 DVSS 0.028184f
C5882 DVDD.n5466 DVSS 0.028184f
C5883 DVDD.n5467 DVSS 0.028184f
C5884 DVDD.n5468 DVSS 0.012306f
C5885 DVDD.n5469 DVSS 0.014092f
C5886 DVDD.n5470 DVSS 0.003163f
C5887 DVDD.n5471 DVSS 0.004391f
C5888 DVDD.n5472 DVSS 0.002071f
C5889 DVDD.n5473 DVSS 0.008435f
C5890 DVDD.n5474 DVSS 0.013072f
C5891 DVDD.n5475 DVSS 0.010076f
C5892 DVDD.n5476 DVSS 0.010076f
C5893 DVDD.n5477 DVSS 0.01023f
C5894 DVDD.n5478 DVSS 0.00844f
C5895 DVDD.n5479 DVSS -0.045065f
C5896 DVDD.n5480 DVSS -0.023927f
C5897 DVDD.t15 DVSS 0.038348f
C5898 DVDD.t40 DVSS 0.046552f
C5899 DVDD.t55 DVSS 0.046552f
C5900 DVDD.t73 DVSS 0.046552f
C5901 DVDD.t48 DVSS 0.046552f
C5902 DVDD.t34 DVSS 0.046552f
C5903 DVDD.t44 DVSS 0.046552f
C5904 DVDD.t19 DVSS 0.06296f
C5905 DVDD.t64 DVSS 0.06296f
C5906 DVDD.t36 DVSS 0.046552f
C5907 DVDD.t38 DVSS 0.046552f
C5908 DVDD.t46 DVSS 0.046552f
C5909 DVDD.t62 DVSS 0.046552f
C5910 DVDD.t0 DVSS 0.046552f
C5911 DVDD.t2 DVSS 0.065353f
C5912 DVDD.n5481 DVSS 0.070654f
C5913 DVDD.n5482 DVSS 0.005596f
C5914 DVDD.n5483 DVSS 0.003163f
C5915 DVDD.n5484 DVSS 0.001538f
C5916 DVDD.n5485 DVSS 0.003076f
C5917 DVDD.n5486 DVSS 0.003076f
C5918 DVDD.n5487 DVSS 0.003076f
C5919 DVDD.n5488 DVSS 0.003076f
C5920 DVDD.n5489 DVSS 0.003076f
C5921 DVDD.n5490 DVSS 0.003076f
C5922 DVDD.n5491 DVSS 0.003076f
C5923 DVDD.n5492 DVSS 0.003076f
C5924 DVDD.n5493 DVSS 0.001538f
C5925 DVDD.n5494 DVSS 0.025778f
C5926 DVDD.n5495 DVSS 0.001538f
C5927 DVDD.n5496 DVSS 0.025778f
C5928 DVDD.n5497 DVSS 0.026423f
C5929 DVDD.n5498 DVSS 0.00134f
C5930 DVDD.n5499 DVSS 0.001538f
C5931 DVDD.n5500 DVSS 0.054096f
C5932 DVDD.n5501 DVSS 0.054096f
C5933 DVDD.n5502 DVSS 0.001538f
C5934 DVDD.n5503 DVSS 0.054232f
C5935 DVDD.n5505 DVSS 0.004122f
C5936 DVDD.n5506 DVSS 0.054232f
C5937 DVDD.n5507 DVSS 0.004122f
C5938 DVDD.n5508 DVSS 0.054232f
C5939 DVDD.n5509 DVSS 0.054232f
C5940 DVDD.n5510 DVSS 0.001538f
C5941 DVDD.n5511 DVSS 0.054096f
C5942 DVDD.n5512 DVSS 0.054096f
C5943 DVDD.n5513 DVSS 0.001538f
C5944 DVDD.n5514 DVSS 0.319527f
C5945 DVDD.n5515 DVSS 0.010218f
C5946 DVDD.n5516 DVSS 0.382769f
C5947 DVDD.n5517 DVSS 0.042587f
C5948 DVDD.n5518 DVSS 0.027687f
C5949 DVDD.n5519 DVSS 0.01188f
C5950 DVDD.t113 DVSS 0.032253f
C5951 DVDD.t110 DVSS 0.032253f
C5952 DVDD.n5520 DVSS 0.064506f
C5953 DVDD.n5521 DVSS 0.011628f
C5954 DVDD.n5522 DVSS 0.060706f
C5955 DVDD.n5523 DVSS 0.048073f
C5956 DVDD.n5524 DVSS 0.055616f
C5957 DVDD.n5525 DVSS 0.007181f
C5958 DVDD.n5526 DVSS -0.285103f
C5959 DVDD.n5527 DVSS 1.00617f
C5960 DVDD.n5528 DVSS 0.672128f
C5961 DVDD.n5529 DVSS 0.010161f
C5962 DVDD.n5530 DVSS 0.01883f
C5963 DVDD.n5531 DVSS 0.01883f
C5964 DVDD.n5532 DVSS 0.01883f
C5965 DVDD.n5533 DVSS 0.01883f
C5966 DVDD.n5534 DVSS 0.031135f
C5967 DVDD.n5535 DVSS 0.031135f
C5968 DVDD.n5536 DVSS 0.01883f
C5969 DVDD.n5537 DVSS 0.01883f
C5970 DVDD.n5538 DVSS 0.01883f
C5971 DVDD.n5539 DVSS 0.01883f
C5972 DVDD.n5540 DVSS 0.01883f
C5973 DVDD.n5541 DVSS 0.01883f
C5974 DVDD.n5542 DVSS 0.01883f
C5975 DVDD.n5543 DVSS 0.01883f
C5976 DVDD.n5544 DVSS 0.042589f
C5977 DVDD.n5545 DVSS 0.382842f
C5978 DVDD.n5546 DVSS 0.117573f
C5979 DVDD.n5547 DVSS 0.035866f
C5980 DVDD.n5548 DVSS 0.012107f
C5981 DVDD.n5549 DVSS 0.012107f
C5982 DVDD.n5550 DVSS 0.012107f
C5983 DVDD.n5551 DVSS 0.012107f
C5984 DVDD.n5552 DVSS 0.012107f
C5985 DVDD.n5553 DVSS 0.012107f
C5986 DVDD.n5554 DVSS 0.012107f
C5987 DVDD.n5555 DVSS 0.012107f
C5988 DVDD.n5556 DVSS 0.024413f
C5989 DVDD.n5557 DVSS 0.024413f
C5990 DVDD.n5558 DVSS 0.012107f
C5991 DVDD.n5559 DVSS 0.012107f
C5992 DVDD.n5560 DVSS 0.012107f
C5993 DVDD.n5561 DVSS 0.012107f
C5994 DVDD.n5562 DVSS 0.008597f
C5995 DVDD.n5563 DVSS 0.027944f
C5996 DVDD.t120 DVSS 0.032253f
C5997 DVDD.t95 DVSS 0.032253f
C5998 DVDD.n5564 DVSS 0.064506f
C5999 DVDD.n5565 DVSS 0.011628f
C6000 DVDD.n5566 DVSS 0.023039f
C6001 DVDD.n5567 DVSS 0.010938f
C6002 DVDD.n5568 DVSS 0.01233f
C6003 DVDD.n5569 DVSS 0.010767f
C6004 DVDD.n5570 DVSS 0.024661f
C6005 DVDD.n5571 DVSS 0.024661f
C6006 DVDD.n5572 DVSS 0.024661f
C6007 DVDD.n5573 DVSS 0.024661f
C6008 DVDD.n5574 DVSS 0.024661f
C6009 DVDD.n5575 DVSS 0.014849f
C6010 DVDD.n5576 DVSS 0.024661f
C6011 DVDD.n5577 DVSS 0.024661f
C6012 DVDD.n5578 DVSS 0.024661f
C6013 DVDD.n5579 DVSS 0.024661f
C6014 DVDD.n5580 DVSS 0.024661f
C6015 DVDD.n5581 DVSS 0.024661f
C6016 DVDD.n5582 DVSS 0.024661f
C6017 DVDD.n5583 DVSS 0.024661f
C6018 DVDD.n5584 DVSS 0.024661f
C6019 DVDD.n5585 DVSS 0.024661f
C6020 DVDD.n5586 DVSS 0.024661f
C6021 DVDD.n5587 DVSS 0.024661f
C6022 DVDD.n5588 DVSS 0.024661f
C6023 DVDD.n5589 DVSS 0.024661f
C6024 DVDD.n5590 DVSS 0.024661f
C6025 DVDD.n5591 DVSS 0.024661f
C6026 DVDD.n5592 DVSS 0.024661f
C6027 DVDD.n5593 DVSS 0.024661f
C6028 DVDD.n5594 DVSS 0.024661f
C6029 DVDD.n5595 DVSS 0.024661f
C6030 DVDD.n5596 DVSS 0.024661f
C6031 DVDD.n5597 DVSS 0.024661f
C6032 DVDD.n5598 DVSS 0.024661f
C6033 DVDD.n5599 DVSS 0.024661f
C6034 DVDD.n5600 DVSS 0.024661f
C6035 DVDD.n5601 DVSS 0.024661f
C6036 DVDD.n5602 DVSS 0.024661f
C6037 DVDD.n5603 DVSS 0.024661f
C6038 DVDD.n5604 DVSS 0.024661f
C6039 DVDD.n5605 DVSS 0.024661f
C6040 DVDD.n5606 DVSS 0.024661f
C6041 DVDD.n5607 DVSS 0.024661f
C6042 DVDD.n5608 DVSS 0.014849f
C6043 DVDD.n5609 DVSS 0.001538f
C6044 DVDD.n5610 DVSS 0.001538f
C6045 DVDD.n5611 DVSS 0.001538f
C6046 DVDD.n5612 DVSS 0.01233f
C6047 DVDD.n5613 DVSS 0.001538f
C6048 DVDD.n5614 DVSS 0.001538f
C6049 DVDD.n5615 DVSS 0.01233f
C6050 DVDD.n5616 DVSS 0.001774f
C6051 DVDD.n5617 DVSS 0.006289f
C6052 DVDD.n5618 DVSS 0.024004f
C6053 DVDD.n5619 DVSS 0.027687f
C6054 DVDD.n5620 DVSS 0.030727f
C6055 DVDD.n5621 DVSS 0.018359f
C6056 DVDD.n5622 DVSS 0.026423f
C6057 DVDD.n5623 DVSS 0.001848f
C6058 DVDD.n5624 DVSS 0.008262f
C6059 DVDD.n5625 DVSS 0.027687f
C6060 DVDD.n5626 DVSS 0.01188f
C6061 DVDD.t117 DVSS 0.032253f
C6062 DVDD.t118 DVSS 0.032253f
C6063 DVDD.n5627 DVSS 0.064506f
C6064 DVDD.n5628 DVSS 0.011628f
C6065 DVDD.n5629 DVSS 0.027944f
C6066 DVDD.n5630 DVSS 0.001538f
C6067 DVDD.n5631 DVSS 0.001848f
C6068 DVDD.n5632 DVSS 0.003076f
C6069 DVDD.n5633 DVSS 0.026423f
C6070 DVDD.n5634 DVSS 0.018359f
C6071 DVDD.n5635 DVSS 0.026423f
C6072 DVDD.n5636 DVSS 0.00289f
C6073 DVDD.n5637 DVSS 0.004317f
C6074 DVDD.n5638 DVSS 0.004503f
C6075 DVDD.n5639 DVSS 0.026423f
C6076 DVDD.n5640 DVSS 0.001538f
C6077 DVDD.n5641 DVSS 0.001551f
C6078 DVDD.n5642 DVSS 0.026423f
C6079 DVDD.n5643 DVSS 0.005768f
C6080 DVDD.n5644 DVSS 0.004317f
C6081 DVDD.n5645 DVSS 0.001625f
C6082 DVDD.n5646 DVSS 0.026423f
C6083 DVDD.n5647 DVSS 0.002394f
C6084 DVDD.n5648 DVSS 0.004317f
C6085 DVDD.n5649 DVSS 0.027944f
C6086 DVDD.t139 DVSS 0.032253f
C6087 DVDD.t128 DVSS 0.032253f
C6088 DVDD.n5650 DVSS 0.064506f
C6089 DVDD.n5651 DVSS 0.011628f
C6090 DVDD.n5652 DVSS 0.011569f
C6091 DVDD.n5653 DVSS 0.013398f
C6092 DVDD.n5654 DVSS 0.026423f
C6093 DVDD.n5655 DVSS 0.069084f
C6094 DVDD.n5656 DVSS 0.069084f
C6095 DVDD.n5657 DVSS 0.008245f
C6096 DVDD.n5658 DVSS 0.0032f
C6097 DVDD.n5659 DVSS 0.003076f
C6098 DVDD.n5660 DVSS 0.007046f
C6099 DVDD.n5661 DVSS 0.006751f
C6100 DVDD.n5662 DVSS 0.019986f
C6101 DVDD.n5663 DVSS 0.007046f
C6102 DVDD.n5664 DVSS 0.007046f
C6103 DVDD.n5665 DVSS 0.003076f
C6104 DVDD.n5666 DVSS 0.003523f
C6105 DVDD.n5667 DVSS 0.008245f
C6106 DVDD.n5668 DVSS 0.008245f
C6107 DVDD.n5669 DVSS 0.017714f
C6108 DVDD.n5670 DVSS 0.026001f
C6109 DVDD.n5671 DVSS 0.028184f
C6110 DVDD.n5672 DVSS 0.028184f
C6111 DVDD.n5673 DVSS 0.028184f
C6112 DVDD.n5674 DVSS 0.028184f
C6113 DVDD.n5675 DVSS 0.028184f
C6114 DVDD.n5676 DVSS 0.028184f
C6115 DVDD.n5677 DVSS 0.028184f
C6116 DVDD.n5678 DVSS 0.028184f
C6117 DVDD.n5679 DVSS 0.028184f
C6118 DVDD.n5680 DVSS 0.028184f
C6119 DVDD.n5681 DVSS 0.028184f
C6120 DVDD.n5682 DVSS 0.028184f
C6121 DVDD.n5683 DVSS 0.028184f
C6122 DVDD.n5684 DVSS 0.028184f
C6123 DVDD.n5685 DVSS 0.028184f
C6124 DVDD.n5686 DVSS 0.028184f
C6125 DVDD.n5687 DVSS 0.024214f
C6126 DVDD.n5688 DVSS 0.024214f
C6127 DVDD.n5689 DVSS 0.024214f
C6128 DVDD.n5690 DVSS 0.040514f
C6129 DVDD.n5691 DVSS 0.018062f
C6130 DVDD.n5692 DVSS 0.028184f
C6131 DVDD.n5693 DVSS 0.028184f
C6132 DVDD.n5694 DVSS 0.028184f
C6133 DVDD.n5695 DVSS 0.028184f
C6134 DVDD.n5696 DVSS 0.028184f
C6135 DVDD.n5697 DVSS 0.028184f
C6136 DVDD.n5698 DVSS 0.028184f
C6137 DVDD.n5699 DVSS 0.028184f
C6138 DVDD.n5700 DVSS 0.028184f
C6139 DVDD.n5701 DVSS 0.028184f
C6140 DVDD.n5702 DVSS 0.012306f
C6141 DVDD.n5703 DVSS 0.014092f
C6142 DVDD.n5704 DVSS 0.003163f
C6143 DVDD.n5705 DVSS 0.004391f
C6144 DVDD.n5706 DVSS 0.002071f
C6145 DVDD.n5707 DVSS 0.009654f
C6146 DVDD.n5708 DVSS 0.010076f
C6147 DVDD.n5709 DVSS 0.012648f
C6148 DVDD.n5710 DVSS 0.070654f
C6149 DVDD.n5711 DVSS 0.005596f
C6150 DVDD.n5712 DVSS 0.004305f
C6151 DVDD.n5713 DVSS 0.026423f
C6152 DVDD.n5714 DVSS 0.085321f
C6153 DVDD.n5715 DVSS 0.085321f
C6154 DVDD.n5716 DVSS 0.003076f
C6155 DVDD.n5717 DVSS 0.023631f
C6156 DVDD.n5718 DVSS 0.023073f
C6157 DVDD.n5719 DVSS 0.052845f
C6158 DVDD.n5720 DVSS 0.052845f
C6159 DVDD.n5721 DVSS 0.023073f
C6160 DVDD.n5722 DVSS 0.026423f
C6161 DVDD.n5723 DVSS 0.003076f
C6162 DVDD.n5724 DVSS 0.003076f
C6163 DVDD.n5725 DVSS 0.026423f
C6164 DVDD.n5726 DVSS 0.023073f
C6165 DVDD.n5727 DVSS 0.03889f
C6166 DVDD.n5728 DVSS 0.03889f
C6167 DVDD.n5729 DVSS 0.462884f
C6168 DVDD.n5730 DVSS 0.040378f
C6169 DVDD.n5731 DVSS 0.052845f
C6170 DVDD.n5732 DVSS 0.052845f
C6171 DVDD.n5733 DVSS 0.052845f
C6172 DVDD.n5734 DVSS 0.052845f
C6173 DVDD.n5735 DVSS 0.052845f
C6174 DVDD.n5736 DVSS 0.08485f
C6175 DVDD.n5737 DVSS 0.08485f
C6176 DVDD.n5738 DVSS 0.08485f
C6177 DVDD.n5739 DVSS 0.052845f
C6178 DVDD.n5740 DVSS 0.052845f
C6179 DVDD.n5741 DVSS 0.052845f
C6180 DVDD.n5742 DVSS 0.052845f
C6181 DVDD.n5743 DVSS 0.040378f
C6182 DVDD.n5744 DVSS 0.040378f
C6183 DVDD.n5745 DVSS 0.206339f
C6184 DVDD.n5746 DVSS 0.005185f
C6185 DVDD.n5747 DVSS 0.005185f
C6186 DVDD.n5748 DVSS 0.007046f
C6187 DVDD.n5749 DVSS 0.020366f
C6188 DVDD.n5750 DVSS 0.007046f
C6189 DVDD.n5751 DVSS 0.007046f
C6190 DVDD.n5752 DVSS 0.003076f
C6191 DVDD.n5753 DVSS 0.003151f
C6192 DVDD.n5754 DVSS 0.007112f
C6193 DVDD.n5755 DVSS 0.014694f
C6194 DVDD.n5756 DVSS 0.025864f
C6195 DVDD.n5757 DVSS 0.005483f
C6196 DVDD.n5758 DVSS 0.004466f
C6197 DVDD.n5759 DVSS 4.9e-19
C6198 DVDD.n5760 DVSS 5.09e-19
C6199 DVDD.n5761 DVSS 0.001161f
C6200 DVDD.n5762 DVSS 0.001161f
C6201 DVDD.n5763 DVSS 5.28e-19
C6202 DVDD.n5764 DVSS 9.8e-19
C6203 DVDD.n5765 DVSS 0.001161f
C6204 DVDD.n5766 DVSS 0.001161f
C6205 DVDD.n5767 DVSS 9.8e-19
C6206 DVDD.n5768 DVSS 9.8e-19
C6207 DVDD.n5769 DVSS 0.001161f
C6208 DVDD.n5770 DVSS 0.001161f
C6209 DVDD.n5771 DVSS 9.8e-19
C6210 DVDD.n5772 DVSS 9.8e-19
C6211 DVDD.n5773 DVSS 0.001161f
C6212 DVDD.n5774 DVSS 0.001161f
C6213 DVDD.n5775 DVSS 9.8e-19
C6214 DVDD.n5776 DVSS 9.8e-19
C6215 DVDD.n5777 DVSS 0.001161f
C6216 DVDD.n5778 DVSS 0.001161f
C6217 DVDD.n5779 DVSS 9.8e-19
C6218 DVDD.n5780 DVSS 9.8e-19
C6219 DVDD.n5781 DVSS 0.001161f
C6220 DVDD.n5782 DVSS 0.001161f
C6221 DVDD.n5783 DVSS 9.8e-19
C6222 DVDD.n5784 DVSS 9.8e-19
C6223 DVDD.n5785 DVSS 0.001161f
C6224 DVDD.n5786 DVSS 0.001161f
C6225 DVDD.n5787 DVSS 9.8e-19
C6226 DVDD.n5788 DVSS 9.8e-19
C6227 DVDD.n5789 DVSS 0.001161f
C6228 DVDD.n5790 DVSS 0.001161f
C6229 DVDD.n5791 DVSS 9.8e-19
C6230 DVDD.n5792 DVSS 9.8e-19
C6231 DVDD.n5793 DVSS 0.001161f
C6232 DVDD.n5794 DVSS 0.001161f
C6233 DVDD.n5795 DVSS 9.8e-19
C6234 DVDD.n5796 DVSS 9.8e-19
C6235 DVDD.n5797 DVSS 0.001161f
C6236 DVDD.n5798 DVSS 0.001161f
C6237 DVDD.n5799 DVSS 9.8e-19
C6238 DVDD.n5800 DVSS 9.8e-19
C6239 DVDD.n5801 DVSS 0.001161f
C6240 DVDD.n5802 DVSS 0.001161f
C6241 DVDD.n5803 DVSS 9.8e-19
C6242 DVDD.n5804 DVSS 0.001161f
C6243 DVDD.n5805 DVSS 0.001161f
C6244 DVDD.n5806 DVSS 8.2e-19
C6245 DVDD.n5807 DVSS 4.9e-19
C6246 DVDD.n5808 DVSS 0.004466f
C6247 DVDD.n5809 DVSS 4.9e-19
C6248 DVDD.n5810 DVSS 6.32e-19
C6249 DVDD.n5811 DVSS 0.001161f
C6250 DVDD.n5812 DVSS 0.001161f
C6251 DVDD.n5813 DVSS 9.8e-19
C6252 DVDD.n5814 DVSS 9.8e-19
C6253 DVDD.n5815 DVSS 0.001161f
C6254 DVDD.n5816 DVSS 0.001161f
C6255 DVDD.n5817 DVSS 9.8e-19
C6256 DVDD.n5818 DVSS 9.8e-19
C6257 DVDD.n5819 DVSS 0.001161f
C6258 DVDD.n5820 DVSS 0.001161f
C6259 DVDD.n5821 DVSS 9.8e-19
C6260 DVDD.n5822 DVSS 9.8e-19
C6261 DVDD.n5823 DVSS 0.001161f
C6262 DVDD.n5824 DVSS 0.001161f
C6263 DVDD.n5825 DVSS 9.8e-19
C6264 DVDD.n5826 DVSS 9.8e-19
C6265 DVDD.n5827 DVSS 0.001161f
C6266 DVDD.n5828 DVSS 0.001161f
C6267 DVDD.n5829 DVSS 9.8e-19
C6268 DVDD.n5830 DVSS 0.001161f
C6269 DVDD.n5831 DVSS 0.002855f
C6270 DVDD.n5832 DVSS 1.14e-19
C6271 DVDD.n5833 DVSS 0.001691f
C6272 DVDD.n5834 DVSS 8.77e-19
C6273 DVDD.n5835 DVSS 8.77e-19
C6274 DVDD.n5836 DVSS 8.77e-19
C6275 DVDD.n5837 DVSS 0.001161f
C6276 DVDD.n5838 DVSS 8.77e-19
C6277 DVDD.n5839 DVSS 8.77e-19
C6278 DVDD.n5840 DVSS 8.77e-19
C6279 DVDD.n5841 DVSS 8.77e-19
C6280 DVDD.n5842 DVSS 0.001161f
C6281 DVDD.n5843 DVSS 8.77e-19
C6282 DVDD.n5844 DVSS 8.77e-19
C6283 DVDD.n5845 DVSS 8.77e-19
C6284 DVDD.n5846 DVSS 8.77e-19
C6285 DVDD.n5847 DVSS 0.001161f
C6286 DVDD.n5848 DVSS 8.77e-19
C6287 DVDD.n5849 DVSS 8.77e-19
C6288 DVDD.n5850 DVSS 8.77e-19
C6289 DVDD.n5851 DVSS 8.77e-19
C6290 DVDD.n5852 DVSS 0.001161f
C6291 DVDD.n5853 DVSS 8.77e-19
C6292 DVDD.n5854 DVSS 8.77e-19
C6293 DVDD.n5855 DVSS 8.77e-19
C6294 DVDD.n5856 DVSS 8.77e-19
C6295 DVDD.n5857 DVSS 0.001161f
C6296 DVDD.n5858 DVSS 8.77e-19
C6297 DVDD.n5859 DVSS 8.77e-19
C6298 DVDD.n5860 DVSS 8.77e-19
C6299 DVDD.n5861 DVSS 8.77e-19
C6300 DVDD.n5862 DVSS 0.001161f
C6301 DVDD.n5863 DVSS 8.77e-19
C6302 DVDD.n5864 DVSS 8.77e-19
C6303 DVDD.n5865 DVSS 8.77e-19
C6304 DVDD.n5866 DVSS 8.77e-19
C6305 DVDD.n5867 DVSS 0.001161f
C6306 DVDD.n5868 DVSS 8.77e-19
C6307 DVDD.n5869 DVSS 8.77e-19
C6308 DVDD.n5870 DVSS 8.77e-19
C6309 DVDD.n5871 DVSS 8.77e-19
C6310 DVDD.n5872 DVSS 0.001189f
C6311 DVDD.n5873 DVSS 9.45e-19
C6312 DVDD.n5874 DVSS 0.00209f
C6313 DVDD.n5875 DVSS 0.002922f
C6314 DVDD.n5876 DVSS 0.002922f
C6315 DVDD.n5877 DVSS 0.350325f
C6316 DVDD.n5879 DVSS 0.001691f
C6317 DVDD.n5880 DVSS 0.0013f
C6318 DVDD.n5881 DVSS 9.28e-19
C6319 DVDD.n5882 DVSS 8.77e-19
C6320 DVDD.n5883 DVSS 0.001161f
C6321 DVDD.n5884 DVSS 0.150384f
C6322 DVDD.t7 DVSS 0.088863f
C6323 DVDD.n5885 DVSS 0.116206f
C6324 DVDD.n5886 DVSS 0.177726f
C6325 DVDD.n5887 DVSS 0.001161f
C6326 DVDD.n5888 DVSS 8.77e-19
C6327 DVDD.n5889 DVSS 8.77e-19
C6328 DVDD.n5890 DVSS 8.77e-19
C6329 DVDD.n5891 DVSS 0.001161f
C6330 DVDD.n5892 DVSS 0.143548f
C6331 DVDD.n5893 DVSS 0.177726f
C6332 DVDD.n5894 DVSS 0.095699f
C6333 DVDD.n5895 DVSS 0.001161f
C6334 DVDD.n5896 DVSS 8.77e-19
C6335 DVDD.n5897 DVSS 8.77e-19
C6336 DVDD.n5898 DVSS 8.77e-19
C6337 DVDD.n5899 DVSS 0.001161f
C6338 DVDD.n5900 DVSS 0.157219f
C6339 DVDD.t8 DVSS 0.088863f
C6340 DVDD.n5901 DVSS 0.10937f
C6341 DVDD.n5902 DVSS 0.177726f
C6342 DVDD.n5903 DVSS 0.001161f
C6343 DVDD.n5904 DVSS 8.77e-19
C6344 DVDD.n5905 DVSS 8.77e-19
C6345 DVDD.n5906 DVSS 8.77e-19
C6346 DVDD.n5907 DVSS 0.001161f
C6347 DVDD.n5908 DVSS 0.136712f
C6348 DVDD.n5909 DVSS 0.177726f
C6349 DVDD.n5910 DVSS 0.102534f
C6350 DVDD.n5911 DVSS 0.001161f
C6351 DVDD.n5912 DVSS 8.77e-19
C6352 DVDD.n5913 DVSS 8.77e-19
C6353 DVDD.n5914 DVSS 8.77e-19
C6354 DVDD.n5915 DVSS 0.001161f
C6355 DVDD.n5916 DVSS 0.164055f
C6356 DVDD.t72 DVSS 0.088863f
C6357 DVDD.n5917 DVSS 0.102534f
C6358 DVDD.n5918 DVSS 0.177726f
C6359 DVDD.n5919 DVSS 0.001161f
C6360 DVDD.n5920 DVSS 8.77e-19
C6361 DVDD.n5921 DVSS 8.77e-19
C6362 DVDD.n5922 DVSS 8.77e-19
C6363 DVDD.n5923 DVSS 0.001161f
C6364 DVDD.n5924 DVSS 0.129877f
C6365 DVDD.n5925 DVSS 0.177726f
C6366 DVDD.n5926 DVSS 0.10937f
C6367 DVDD.n5927 DVSS 0.001161f
C6368 DVDD.n5928 DVSS 8.77e-19
C6369 DVDD.n5929 DVSS 8.77e-19
C6370 DVDD.n5930 DVSS 8.77e-19
C6371 DVDD.n5931 DVSS 0.001161f
C6372 DVDD.n5932 DVSS 0.17089f
C6373 DVDD.t61 DVSS 0.088863f
C6374 DVDD.n5933 DVSS 0.095699f
C6375 DVDD.n5934 DVSS 0.177726f
C6376 DVDD.n5935 DVSS 0.001161f
C6377 DVDD.n5936 DVSS 8.77e-19
C6378 DVDD.n5937 DVSS 8.77e-19
C6379 DVDD.n5938 DVSS 8.77e-19
C6380 DVDD.n5939 DVSS 0.001161f
C6381 DVDD.n5940 DVSS 0.123041f
C6382 DVDD.n5941 DVSS 0.177726f
C6383 DVDD.n5942 DVSS 0.116206f
C6384 DVDD.n5943 DVSS 0.001161f
C6385 DVDD.n5944 DVSS 8.77e-19
C6386 DVDD.n5945 DVSS 8.77e-19
C6387 DVDD.n5946 DVSS 9.28e-19
C6388 DVDD.n5947 DVSS 0.001083f
C6389 DVDD.n5948 DVSS 0.220449f
C6390 DVDD.n5949 DVSS 0.001083f
C6391 DVDD.n5950 DVSS 9.28e-19
C6392 DVDD.n5951 DVSS 7.93e-19
C6393 DVDD.n5952 DVSS 0.00159f
C6394 DVDD.n5953 DVSS 9.8e-19
C6395 DVDD.n5954 DVSS 9.8e-19
C6396 DVDD.n5955 DVSS 0.001161f
C6397 DVDD.n5957 DVSS 0.001161f
C6398 DVDD.n5958 DVSS 0.001161f
C6399 DVDD.n5959 DVSS 5.75e-19
C6400 DVDD.n5960 DVSS 9.8e-19
C6401 DVDD.n5961 DVSS 9.8e-19
C6402 DVDD.n5962 DVSS 0.001161f
C6403 DVDD.n5964 DVSS 0.001161f
C6404 DVDD.n5965 DVSS 0.001161f
C6405 DVDD.n5966 DVSS 9.8e-19
C6406 DVDD.n5967 DVSS 9.8e-19
C6407 DVDD.n5968 DVSS 9.8e-19
C6408 DVDD.n5969 DVSS 0.001161f
C6409 DVDD.n5971 DVSS 0.001161f
C6410 DVDD.n5972 DVSS 0.001161f
C6411 DVDD.n5973 DVSS 9.8e-19
C6412 DVDD.n5974 DVSS 9.8e-19
C6413 DVDD.n5975 DVSS 9.8e-19
C6414 DVDD.n5976 DVSS 0.001161f
C6415 DVDD.n5978 DVSS 0.001161f
C6416 DVDD.n5979 DVSS 0.001161f
C6417 DVDD.n5981 DVSS 0.001161f
C6418 DVDD.n5982 DVSS 6.32e-19
C6419 DVDD.n5983 DVSS 4.9e-19
C6420 DVDD.n5984 DVSS 0.001538f
C6421 DVDD.n5985 DVSS 0.001538f
C6422 DVDD.n5986 DVSS 0.001563f
C6423 DVDD.n5987 DVSS 0.01233f
C6424 DVDD.n5988 DVSS 0.020233f
C6425 DVDD.n5989 DVSS 0.024661f
C6426 DVDD.n5990 DVSS 0.024661f
C6427 DVDD.n5991 DVSS 0.024661f
C6428 DVDD.n5992 DVSS 0.024661f
C6429 DVDD.n5993 DVSS 0.024661f
C6430 DVDD.n5994 DVSS 0.018322f
C6431 DVDD.n5995 DVSS 0.024661f
C6432 DVDD.n5996 DVSS 0.024661f
C6433 DVDD.n5997 DVSS 0.024661f
C6434 DVDD.n5998 DVSS 0.024661f
C6435 DVDD.n5999 DVSS 0.024661f
C6436 DVDD.n6000 DVSS 0.024661f
C6437 DVDD.n6001 DVSS 0.024661f
C6438 DVDD.n6002 DVSS 0.024661f
C6439 DVDD.n6003 DVSS 0.024661f
C6440 DVDD.n6004 DVSS 0.024661f
C6441 DVDD.n6005 DVSS 0.024661f
C6442 DVDD.n6006 DVSS 0.024661f
C6443 DVDD.n6007 DVSS 0.024661f
C6444 DVDD.n6008 DVSS 0.024661f
C6445 DVDD.n6009 DVSS 0.024661f
C6446 DVDD.n6010 DVSS 0.024661f
C6447 DVDD.n6011 DVSS 0.024661f
C6448 DVDD.n6012 DVSS 0.024661f
C6449 DVDD.n6013 DVSS 0.024661f
C6450 DVDD.n6014 DVSS 0.024661f
C6451 DVDD.n6015 DVSS 0.02223f
C6452 DVDD.n6016 DVSS 0.024661f
C6453 DVDD.n6017 DVSS 0.012678f
C6454 DVDD.n6018 DVSS 0.032464f
C6455 DVDD.n6019 DVSS 0.118823f
.ends

