* NGSPICE file created from gf180mcu_fd_io__dvdd_pex.ext - technology: gf180mcuD

.subckt gf180mcu_fd_io__dvdd_pex VSS DVSS DVDD
X0 DVDD.t61 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_1.D.t4 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.t6 DVDD.t60 pfet_06v0 ad=1.3p pd=5.52u as=1.3p ps=5.52u w=5u l=0.7u
X1 DVDD.t152 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.t17 DVSS.t188 DVSS.t187 nfet_06v0 ad=12.999999p pd=50.52u as=12.999999p ps=50.52u w=50u l=0.7u
X2 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.t9 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_1.D.t5 DVDD.t59 DVDD.t58 pfet_06v0 ad=1.3p pd=5.52u as=1.3p ps=5.52u w=5u l=0.7u
X3 DVDD.t151 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.t18 DVSS.t186 DVSS.t185 nfet_06v0 ad=12.999999p pd=50.52u as=12.999999p ps=50.52u w=50u l=0.7u
X4 DVDD.t150 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.t19 DVSS.t184 DVSS.t183 nfet_06v0 ad=12.999999p pd=50.52u as=12.999999p ps=50.52u w=50u l=0.7u
X5 DVDD.t57 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_1.D.t6 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.t7 DVDD.t56 pfet_06v0 ad=1.3p pd=5.52u as=1.3p ps=5.52u w=5u l=0.7u
X6 DVDD.t55 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_1.D.t7 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.t14 DVDD.t54 pfet_06v0 ad=2.2p pd=10.879999u as=1.3p ps=5.52u w=5u l=0.7u
X7 DVSS.t182 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.t20 DVDD.t149 DVSS.t181 nfet_06v0 ad=12.999999p pd=50.52u as=12.999999p ps=50.52u w=50u l=0.7u
X8 DVSS.t180 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.t21 DVDD.t148 DVSS.t179 nfet_06v0 ad=12.999999p pd=50.52u as=12.999999p ps=50.52u w=50u l=0.7u
X9 DVSS.t178 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.t22 DVDD.t147 DVSS.t177 nfet_06v0 ad=12.999999p pd=50.52u as=12.999999p ps=50.52u w=50u l=0.7u
X10 DVSS.t176 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.t23 DVDD.t146 DVSS.t175 nfet_06v0 ad=12.999999p pd=50.52u as=12.999999p ps=50.52u w=50u l=0.7u
X11 DVSS.t174 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.t24 DVDD.t145 DVSS.t173 nfet_06v0 ad=12.999999p pd=50.52u as=12.999999p ps=50.52u w=50u l=0.7u
X12 DVDD.t155 DVSS.t28 cap_nmos_06v0 c_width=15u c_length=15u
X13 DVDD.t144 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.t25 DVSS.t172 DVSS.t171 nfet_06v0 ad=12.999999p pd=50.52u as=12.999999p ps=50.52u w=50u l=0.7u
X14 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_1.D.t3 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531459_0.D.t3 DVDD.t154 DVDD.t153 pfet_06v0 ad=2.2p pd=10.879999u as=1.3p ps=5.52u w=5u l=0.7u
X15 DVDD.t143 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.t26 DVSS.t170 DVSS.t169 nfet_06v0 ad=12.999999p pd=50.52u as=12.999999p ps=50.52u w=50u l=0.7u
X16 DVDD.t142 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.t27 DVSS.t168 DVSS.t167 nfet_06v0 ad=12.999999p pd=50.52u as=12.999999p ps=50.52u w=50u l=0.7u
X17 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.t13 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_1.D.t8 DVDD.t53 DVDD.t52 pfet_06v0 ad=1.3p pd=5.52u as=1.3p ps=5.52u w=5u l=0.7u
X18 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.t10 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_1.D.t9 DVDD.t51 DVDD.t50 pfet_06v0 ad=1.3p pd=5.52u as=1.3p ps=5.52u w=5u l=0.7u
X19 DVSS.t166 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.t28 DVDD.t141 DVSS.t165 nfet_06v0 ad=12.999999p pd=50.52u as=12.999999p ps=50.52u w=50u l=0.7u
X20 DVSS.t164 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.t29 DVDD.t140 DVSS.t163 nfet_06v0 ad=12.999999p pd=50.52u as=12.999999p ps=50.52u w=50u l=0.7u
X21 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/comp018green_esd_rc_v5p0_0.ppolyf_u_CDNS_406619531453_1.MINUS.t1 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/comp018green_esd_rc_v5p0_0.ppolyf_u_CDNS_406619531453_0.PLUS.t1 DVDD.t69 ppolyf_u r_width=0.8u r_length=63.854996u
X22 DVDD.t139 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.t30 DVSS.t162 DVSS.t161 nfet_06v0 ad=21.999998p pd=0.10088m as=12.999999p ps=50.52u w=50u l=0.7u
X23 DVDD.t5 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/comp018green_esd_rc_v5p0_0.VRC.t1 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531459_0.D.t1 DVDD.t4 pfet_06v0 ad=1.3p pd=5.52u as=1.3p ps=5.52u w=5u l=0.7u
X24 DVDD.t138 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.t31 DVSS.t160 DVSS.t159 nfet_06v0 ad=12.999999p pd=50.52u as=12.999999p ps=50.52u w=50u l=0.7u
D0 DVSS.t24 DVDD.t156 diode_nd2ps_06v0 pj=82u area=40p
X25 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531459_0.D.t1 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/comp018green_esd_rc_v5p0_0.VRC.t2 DVDD.t3 DVDD.t2 pfet_06v0 ad=1.3p pd=5.52u as=1.3p ps=5.52u w=5u l=0.7u
X26 DVSS.t158 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.t32 DVDD.t137 DVSS.t157 nfet_06v0 ad=12.999999p pd=50.52u as=12.999999p ps=50.52u w=50u l=0.7u
X27 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/comp018green_esd_rc_v5p0_0.ppolyf_u_CDNS_406619531453_5.MINUS.t0 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/comp018green_esd_rc_v5p0_0.ppolyf_u_CDNS_406619531453_3.PLUS.t0 DVDD.t13 ppolyf_u r_width=0.8u r_length=63.854996u
X28 DVSS.t156 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.t33 DVDD.t136 DVSS.t155 nfet_06v0 ad=12.999999p pd=50.52u as=12.999999p ps=50.52u w=50u l=0.7u
X29 DVDD.t157 DVSS.t27 cap_nmos_06v0 c_width=15u c_length=15u
X30 DVDD.t158 DVSS.t26 cap_nmos_06v0 c_width=15u c_length=15u
X31 DVSS.t23 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_1.D.t10 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.t3 DVSS.t22 nfet_06v0 ad=1.3p pd=5.52u as=1.3p ps=5.52u w=5u l=0.7u
X32 DVDD.t135 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.t34 DVSS.t154 DVSS.t153 nfet_06v0 ad=12.999999p pd=50.52u as=12.999999p ps=50.52u w=50u l=0.7u
X33 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.t2 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_1.D.t11 DVSS.t21 DVSS.t20 nfet_06v0 ad=1.3p pd=5.52u as=1.3p ps=5.52u w=5u l=0.7u
X34 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/comp018green_esd_rc_v5p0_0.ppolyf_u_CDNS_406619531453_2.MINUS.t1 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/comp018green_esd_rc_v5p0_0.ppolyf_u_CDNS_406619531453_4.PLUS.t0 DVDD.t68 ppolyf_u r_width=0.8u r_length=63.854996u
X35 DVDD.t134 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.t35 DVSS.t152 DVSS.t151 nfet_06v0 ad=12.999999p pd=50.52u as=12.999999p ps=50.52u w=50u l=0.7u
X36 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.t4 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_1.D.t12 DVDD.t49 DVDD.t48 pfet_06v0 ad=1.3p pd=5.52u as=1.3p ps=5.52u w=5u l=0.7u
X37 DVDD.t133 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.t36 DVSS.t150 DVSS.t149 nfet_06v0 ad=12.999999p pd=50.52u as=12.999999p ps=50.52u w=50u l=0.7u
X38 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531459_0.D.t2 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/comp018green_esd_rc_v5p0_0.VRC.t3 DVSS.t7 DVSS.t6 nfet_06v0 ad=2.2p pd=10.879999u as=2.2p ps=10.879999u w=5u l=0.7u
X39 DVSS.t148 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.t37 DVDD.t132 DVSS.t147 nfet_06v0 ad=12.999999p pd=50.52u as=21.999998p ps=0.10088m w=50u l=0.7u
X40 DVSS.t146 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.t38 DVDD.t131 DVSS.t145 nfet_06v0 ad=12.999999p pd=50.52u as=12.999999p ps=50.52u w=50u l=0.7u
X41 DVSS.t144 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.t39 DVDD.t130 DVSS.t143 nfet_06v0 ad=12.999999p pd=50.52u as=12.999999p ps=50.52u w=50u l=0.7u
X42 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_1.D.t0 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531459_0.D.t4 DVSS.t11 DVSS.t10 nfet_06v0 ad=1.3p pd=5.52u as=2.2p ps=10.879999u w=5u l=0.7u
X43 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.t8 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_1.D.t13 DVDD.t47 DVDD.t46 pfet_06v0 ad=1.3p pd=5.52u as=1.3p ps=5.52u w=5u l=0.7u
X44 DVSS.t142 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.t40 DVDD.t129 DVSS.t141 nfet_06v0 ad=12.999999p pd=50.52u as=12.999999p ps=50.52u w=50u l=0.7u
X45 DVSS.t192 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531459_0.D.t5 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_1.D.t2 DVSS.t191 nfet_06v0 ad=1.3p pd=5.52u as=1.3p ps=5.52u w=5u l=0.7u
X46 DVDD.t128 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.t41 DVSS.t140 DVSS.t139 nfet_06v0 ad=12.999999p pd=50.52u as=12.999999p ps=50.52u w=50u l=0.7u
X47 DVDD.t45 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_1.D.t14 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.t15 DVDD.t44 pfet_06v0 ad=1.3p pd=5.52u as=1.3p ps=5.52u w=5u l=0.7u
X48 DVDD.t127 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.t42 DVSS.t138 DVSS.t137 nfet_06v0 ad=12.999999p pd=50.52u as=12.999999p ps=50.52u w=50u l=0.7u
X49 DVDD.t126 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.t43 DVSS.t136 DVSS.t135 nfet_06v0 ad=12.999999p pd=50.52u as=12.999999p ps=50.52u w=50u l=0.7u
X50 DVDD.t125 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.t44 DVSS.t134 DVSS.t133 nfet_06v0 ad=12.999999p pd=50.52u as=12.999999p ps=50.52u w=50u l=0.7u
X51 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.t15 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_1.D.t15 DVDD.t43 DVDD.t42 pfet_06v0 ad=1.3p pd=5.52u as=1.3p ps=5.52u w=5u l=0.7u
X52 DVDD.t124 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.t45 DVSS.t132 DVSS.t131 nfet_06v0 ad=12.999999p pd=50.52u as=12.999999p ps=50.52u w=50u l=0.7u
X53 DVDD.t41 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_1.D.t16 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.t5 DVDD.t40 pfet_06v0 ad=1.3p pd=5.52u as=1.3p ps=5.52u w=5u l=0.7u
X54 DVSS.t130 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.t46 DVDD.t123 DVSS.t129 nfet_06v0 ad=12.999999p pd=50.52u as=12.999999p ps=50.52u w=50u l=0.7u
X55 DVDD.t122 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.t47 DVSS.t128 DVSS.t127 nfet_06v0 ad=21.999998p pd=0.10088m as=12.999999p ps=50.52u w=50u l=0.7u
X56 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/comp018green_esd_rc_v5p0_0.VRC.t4 DVSS.t4 cap_nmos_06v0 c_width=25u c_length=10u
X57 DVDD.t121 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.t48 DVSS.t126 DVSS.t125 nfet_06v0 ad=12.999999p pd=50.52u as=12.999999p ps=50.52u w=50u l=0.7u
X58 DVDD.t39 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_1.D.t17 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.t9 DVDD.t38 pfet_06v0 ad=1.3p pd=5.52u as=1.3p ps=5.52u w=5u l=0.7u
X59 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/comp018green_esd_rc_v5p0_0.VRC.t0 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/comp018green_esd_rc_v5p0_0.ppolyf_u_CDNS_406619531453_0.PLUS.t0 DVDD.t65 ppolyf_u r_width=0.8u r_length=63.854996u
X60 DVDD.t120 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.t49 DVSS.t124 DVSS.t123 nfet_06v0 ad=12.999999p pd=50.52u as=12.999999p ps=50.52u w=50u l=0.7u
X61 DVDD.t37 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_1.D.t18 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.t11 DVDD.t36 pfet_06v0 ad=1.3p pd=5.52u as=1.3p ps=5.52u w=5u l=0.7u
X62 DVDD.t119 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.t50 DVSS.t122 DVSS.t121 nfet_06v0 ad=12.999999p pd=50.52u as=12.999999p ps=50.52u w=50u l=0.7u
X63 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/comp018green_esd_rc_v5p0_0.VRC.t5 DVSS.t5 cap_nmos_06v0 c_width=25u c_length=10u
X64 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.t11 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_1.D.t19 DVDD.t35 DVDD.t34 pfet_06v0 ad=1.3p pd=5.52u as=2.2p ps=10.879999u w=5u l=0.7u
X65 DVSS.t120 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.t51 DVDD.t118 DVSS.t119 nfet_06v0 ad=12.999999p pd=50.52u as=12.999999p ps=50.52u w=50u l=0.7u
X66 DVSS.t118 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.t52 DVDD.t117 DVSS.t117 nfet_06v0 ad=12.999999p pd=50.52u as=12.999999p ps=50.52u w=50u l=0.7u
X67 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/comp018green_esd_rc_v5p0_0.VRC.t6 DVSS.t9 cap_nmos_06v0 c_width=25u c_length=10u
X68 DVDD.t33 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_1.D.t20 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.t12 DVDD.t32 pfet_06v0 ad=1.3p pd=5.52u as=1.3p ps=5.52u w=5u l=0.7u
X69 DVDD.t116 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.t53 DVSS.t116 DVSS.t115 nfet_06v0 ad=12.999999p pd=50.52u as=12.999999p ps=50.52u w=50u l=0.7u
X70 DVDD.t115 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.t54 DVSS.t114 DVSS.t113 nfet_06v0 ad=12.999999p pd=50.52u as=12.999999p ps=50.52u w=50u l=0.7u
X71 DVDD.t114 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.t55 DVSS.t112 DVSS.t111 nfet_06v0 ad=12.999999p pd=50.52u as=12.999999p ps=50.52u w=50u l=0.7u
X72 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.t14 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_1.D.t21 DVDD.t31 DVDD.t30 pfet_06v0 ad=1.3p pd=5.52u as=1.3p ps=5.52u w=5u l=0.7u
X73 DVSS.t19 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_1.D.t22 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.t1 DVSS.t18 nfet_06v0 ad=1.3p pd=5.52u as=1.3p ps=5.52u w=5u l=0.7u
X74 DVSS.t110 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.t56 DVDD.t113 DVSS.t109 nfet_06v0 ad=12.999999p pd=50.52u as=12.999999p ps=50.52u w=50u l=0.7u
X75 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.t1 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_1.D.t23 DVSS.t17 DVSS.t16 nfet_06v0 ad=1.3p pd=5.52u as=1.3p ps=5.52u w=5u l=0.7u
X76 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/comp018green_esd_rc_v5p0_0.ppolyf_u_CDNS_406619531453_3.MINUS.t0 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/comp018green_esd_rc_v5p0_0.ppolyf_u_CDNS_406619531453_3.PLUS.t1 DVDD.t66 ppolyf_u r_width=0.8u r_length=63.854996u
X77 DVSS.t108 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.t57 DVDD.t112 DVSS.t107 nfet_06v0 ad=12.999999p pd=50.52u as=12.999999p ps=50.52u w=50u l=0.7u
X78 DVDD.t111 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.t58 DVSS.t106 DVSS.t105 nfet_06v0 ad=12.999999p pd=50.52u as=12.999999p ps=50.52u w=50u l=0.7u
X79 DVSS.t15 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_1.D.t24 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.t0 DVSS.t14 nfet_06v0 ad=2.2p pd=10.879999u as=1.3p ps=5.52u w=5u l=0.7u
X80 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/comp018green_esd_rc_v5p0_0.ppolyf_u_CDNS_406619531453_4.MINUS.t1 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/comp018green_esd_rc_v5p0_0.ppolyf_u_CDNS_406619531453_4.PLUS.t1 DVDD.t70 ppolyf_u r_width=0.8u r_length=63.854996u
X81 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/comp018green_esd_rc_v5p0_0.VRC.t7 DVSS.t1 cap_nmos_06v0 c_width=25u c_length=10u
X82 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/comp018green_esd_rc_v5p0_0.VRC.t8 DVSS.t2 cap_nmos_06v0 c_width=25u c_length=10u
X83 DVDD.t11 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531459_0.D.t6 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_1.D.t1 DVDD.t10 pfet_06v0 ad=1.3p pd=5.52u as=1.3p ps=5.52u w=5u l=0.7u
X84 DVDD.t110 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.t59 DVSS.t104 DVSS.t103 nfet_06v0 ad=12.999999p pd=50.52u as=12.999999p ps=50.52u w=50u l=0.7u
X85 DVDD.t109 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.t60 DVSS.t102 DVSS.t101 nfet_06v0 ad=12.999999p pd=50.52u as=12.999999p ps=50.52u w=50u l=0.7u
X86 DVDD.t108 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.t61 DVSS.t100 DVSS.t99 nfet_06v0 ad=12.999999p pd=50.52u as=12.999999p ps=50.52u w=50u l=0.7u
X87 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/comp018green_esd_rc_v5p0_0.ppolyf_u_CDNS_406619531453_4.MINUS.t0 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/comp018green_esd_rc_v5p0_0.ppolyf_u_CDNS_406619531453_5.PLUS.t0 DVDD.t67 ppolyf_u r_width=0.8u r_length=63.854996u
X88 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_1.D.t1 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531459_0.D.t7 DVDD.t9 DVDD.t8 pfet_06v0 ad=1.3p pd=5.52u as=1.3p ps=5.52u w=5u l=0.7u
X89 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_1.D.t2 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531459_0.D.t8 DVSS.t190 DVSS.t189 nfet_06v0 ad=1.3p pd=5.52u as=1.3p ps=5.52u w=5u l=0.7u
X90 DVSS.t98 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.t62 DVDD.t107 DVSS.t97 nfet_06v0 ad=12.999999p pd=50.52u as=12.999999p ps=50.52u w=50u l=0.7u
X91 DVSS.t198 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531459_0.D.t9 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_1.D.t2 DVSS.t197 nfet_06v0 ad=1.3p pd=5.52u as=1.3p ps=5.52u w=5u l=0.7u
X92 DVDD.t29 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_1.D.t25 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.t16 DVDD.t28 pfet_06v0 ad=1.3p pd=5.52u as=1.3p ps=5.52u w=5u l=0.7u
X93 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/comp018green_esd_rc_v5p0_0.VRC.t9 DVSS.t8 cap_nmos_06v0 c_width=25u c_length=10u
X94 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/comp018green_esd_rc_v5p0_0.VRC.t10 DVSS.t3 cap_nmos_06v0 c_width=25u c_length=10u
X95 DVDD.t106 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.t63 DVSS.t96 DVSS.t95 nfet_06v0 ad=12.999999p pd=50.52u as=12.999999p ps=50.52u w=50u l=0.7u
X96 DVSS.t94 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.t64 DVDD.t105 DVSS.t93 nfet_06v0 ad=12.999999p pd=50.52u as=12.999999p ps=50.52u w=50u l=0.7u
X97 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.t7 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_1.D.t26 DVDD.t27 DVDD.t26 pfet_06v0 ad=1.3p pd=5.52u as=1.3p ps=5.52u w=5u l=0.7u
X98 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.t12 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_1.D.t27 DVDD.t25 DVDD.t24 pfet_06v0 ad=1.3p pd=5.52u as=1.3p ps=5.52u w=5u l=0.7u
X99 DVDD.t104 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.t65 DVSS.t92 DVSS.t91 nfet_06v0 ad=12.999999p pd=50.52u as=12.999999p ps=50.52u w=50u l=0.7u
X100 DVSS.t90 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.t66 DVDD.t103 DVSS.t89 nfet_06v0 ad=12.999999p pd=50.52u as=12.999999p ps=50.52u w=50u l=0.7u
X101 DVSS.t88 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.t67 DVDD.t102 DVSS.t87 nfet_06v0 ad=12.999999p pd=50.52u as=12.999999p ps=50.52u w=50u l=0.7u
X102 DVDD.t64 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/comp018green_esd_rc_v5p0_0.ppolyf_u_CDNS_406619531453_2.PLUS.t1 DVDD.t63 ppolyf_u r_width=0.8u r_length=63.854996u
X103 DVSS.t86 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.t68 DVDD.t101 DVSS.t85 nfet_06v0 ad=12.999999p pd=50.52u as=12.999999p ps=50.52u w=50u l=0.7u
X104 DVSS.t84 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.t69 DVDD.t100 DVSS.t83 nfet_06v0 ad=12.999999p pd=50.52u as=21.999998p ps=0.10088m w=50u l=0.7u
X105 DVDD.t99 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.t70 DVSS.t82 DVSS.t81 nfet_06v0 ad=21.999998p pd=0.10088m as=12.999999p ps=50.52u w=50u l=0.7u
X106 DVDD.t98 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.t71 DVSS.t80 DVSS.t79 nfet_06v0 ad=12.999999p pd=50.52u as=12.999999p ps=50.52u w=50u l=0.7u
D1 DVSS.t24 DVDD.t159 diode_nd2ps_06v0 pj=82u area=40p
X107 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/comp018green_esd_rc_v5p0_0.VRC.t11 DVSS.t0 cap_nmos_06v0 c_width=25u c_length=10u
X108 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.t5 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_1.D.t28 DVDD.t23 DVDD.t22 pfet_06v0 ad=1.3p pd=5.52u as=1.3p ps=5.52u w=5u l=0.7u
X109 DVDD.t97 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.t72 DVSS.t78 DVSS.t77 nfet_06v0 ad=12.999999p pd=50.52u as=12.999999p ps=50.52u w=50u l=0.7u
X110 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.t16 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_1.D.t29 DVDD.t21 DVDD.t20 pfet_06v0 ad=1.3p pd=5.52u as=1.3p ps=5.52u w=5u l=0.7u
X111 DVSS.t76 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.t73 DVDD.t96 DVSS.t75 nfet_06v0 ad=12.999999p pd=50.52u as=12.999999p ps=50.52u w=50u l=0.7u
X112 DVSS.t74 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.t74 DVDD.t95 DVSS.t73 nfet_06v0 ad=12.999999p pd=50.52u as=12.999999p ps=50.52u w=50u l=0.7u
D2 DVSS.t24 DVDD.t160 diode_nd2ps_06v0 pj=82u area=40p
X113 DVDD.t19 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_1.D.t30 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.t13 DVDD.t18 pfet_06v0 ad=1.3p pd=5.52u as=1.3p ps=5.52u w=5u l=0.7u
X114 DVSS.t72 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.t75 DVDD.t94 DVSS.t71 nfet_06v0 ad=12.999999p pd=50.52u as=21.999998p ps=0.10088m w=50u l=0.7u
X115 DVSS.t70 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.t76 DVDD.t93 DVSS.t69 nfet_06v0 ad=12.999999p pd=50.52u as=12.999999p ps=50.52u w=50u l=0.7u
X116 DVDD.t17 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_1.D.t31 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.t10 DVDD.t16 pfet_06v0 ad=1.3p pd=5.52u as=1.3p ps=5.52u w=5u l=0.7u
X117 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/comp018green_esd_rc_v5p0_0.ppolyf_u_CDNS_406619531453_3.MINUS.t1 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/comp018green_esd_rc_v5p0_0.ppolyf_u_CDNS_406619531453_1.PLUS.t1 DVDD.t71 ppolyf_u r_width=0.8u r_length=63.854996u
X118 DVDD.t92 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.t77 DVSS.t68 DVSS.t67 nfet_06v0 ad=12.999999p pd=50.52u as=12.999999p ps=50.52u w=50u l=0.7u
X119 DVDD.t91 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.t78 DVSS.t66 DVSS.t65 nfet_06v0 ad=12.999999p pd=50.52u as=12.999999p ps=50.52u w=50u l=0.7u
X120 DVDD.t90 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.t79 DVSS.t64 DVSS.t63 nfet_06v0 ad=12.999999p pd=50.52u as=12.999999p ps=50.52u w=50u l=0.7u
X121 DVDD.t161 DVSS.t25 cap_nmos_06v0 c_width=15u c_length=15u
X122 DVSS.t62 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.t80 DVDD.t89 DVSS.t61 nfet_06v0 ad=12.999999p pd=50.52u as=12.999999p ps=50.52u w=50u l=0.7u
X123 DVSS.t60 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.t81 DVDD.t88 DVSS.t59 nfet_06v0 ad=12.999999p pd=50.52u as=12.999999p ps=50.52u w=50u l=0.7u
X124 DVSS.t58 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.t82 DVDD.t87 DVSS.t57 nfet_06v0 ad=12.999999p pd=50.52u as=12.999999p ps=50.52u w=50u l=0.7u
X125 DVSS.t56 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.t83 DVDD.t86 DVSS.t55 nfet_06v0 ad=12.999999p pd=50.52u as=12.999999p ps=50.52u w=50u l=0.7u
X126 DVSS.t54 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.t84 DVDD.t85 DVSS.t53 nfet_06v0 ad=12.999999p pd=50.52u as=12.999999p ps=50.52u w=50u l=0.7u
X127 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/comp018green_esd_rc_v5p0_0.ppolyf_u_CDNS_406619531453_1.MINUS.t0 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/comp018green_esd_rc_v5p0_0.ppolyf_u_CDNS_406619531453_1.PLUS.t0 DVDD.t12 ppolyf_u r_width=0.8u r_length=63.854996u
X128 DVDD.t84 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.t85 DVSS.t52 DVSS.t51 nfet_06v0 ad=12.999999p pd=50.52u as=12.999999p ps=50.52u w=50u l=0.7u
X129 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_1.D.t2 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531459_0.D.t10 DVSS.t196 DVSS.t195 nfet_06v0 ad=1.3p pd=5.52u as=1.3p ps=5.52u w=5u l=0.7u
X130 DVDD.t83 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.t86 DVSS.t50 DVSS.t49 nfet_06v0 ad=12.999999p pd=50.52u as=12.999999p ps=50.52u w=50u l=0.7u
X131 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/comp018green_esd_rc_v5p0_0.ppolyf_u_CDNS_406619531453_5.MINUS.t1 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/comp018green_esd_rc_v5p0_0.ppolyf_u_CDNS_406619531453_5.PLUS.t1 DVDD.t72 ppolyf_u r_width=0.8u r_length=63.854996u
X132 DVSS.t48 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.t87 DVDD.t82 DVSS.t47 nfet_06v0 ad=12.999999p pd=50.52u as=12.999999p ps=50.52u w=50u l=0.7u
D3 DVSS.t24 DVDD.t162 diode_nd2ps_06v0 pj=82u area=40p
X133 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.t0 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_1.D.t32 DVSS.t13 DVSS.t12 nfet_06v0 ad=1.3p pd=5.52u as=1.3p ps=5.52u w=5u l=0.7u
X134 DVDD.t7 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/comp018green_esd_rc_v5p0_0.VRC.t12 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531459_0.D.t0 DVDD.t6 pfet_06v0 ad=1.3p pd=5.52u as=1.3p ps=5.52u w=5u l=0.7u
X135 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531459_0.D.t0 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/comp018green_esd_rc_v5p0_0.VRC.t13 DVDD.t1 DVDD.t0 pfet_06v0 ad=1.3p pd=5.52u as=2.2p ps=10.879999u w=5u l=0.7u
X136 DVSS.t46 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.t88 DVDD.t81 DVSS.t45 nfet_06v0 ad=12.999999p pd=50.52u as=12.999999p ps=50.52u w=50u l=0.7u
X137 DVSS.t44 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.t89 DVDD.t80 DVSS.t43 nfet_06v0 ad=12.999999p pd=50.52u as=12.999999p ps=50.52u w=50u l=0.7u
X138 DVSS.t42 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.t90 DVDD.t79 DVSS.t41 nfet_06v0 ad=12.999999p pd=50.52u as=21.999998p ps=0.10088m w=50u l=0.7u
X139 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/comp018green_esd_rc_v5p0_0.ppolyf_u_CDNS_406619531453_2.MINUS.t0 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/comp018green_esd_rc_v5p0_0.ppolyf_u_CDNS_406619531453_2.PLUS.t0 DVDD.t62 ppolyf_u r_width=0.8u r_length=63.854996u
X140 DVDD.t78 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.t91 DVSS.t40 DVSS.t39 nfet_06v0 ad=12.999999p pd=50.52u as=12.999999p ps=50.52u w=50u l=0.7u
X141 DVSS.t194 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531459_0.D.t11 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_1.D.t0 DVSS.t193 nfet_06v0 ad=1.3p pd=5.52u as=1.3p ps=5.52u w=5u l=0.7u
X142 DVDD.t77 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.t92 DVSS.t38 DVSS.t37 nfet_06v0 ad=21.999998p pd=0.10088m as=12.999999p ps=50.52u w=50u l=0.7u
X143 DVDD.t76 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.t93 DVSS.t36 DVSS.t35 nfet_06v0 ad=12.999999p pd=50.52u as=12.999999p ps=50.52u w=50u l=0.7u
X144 DVDD.t15 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_1.D.t33 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.t8 DVDD.t14 pfet_06v0 ad=1.3p pd=5.52u as=1.3p ps=5.52u w=5u l=0.7u
X145 DVSS.t34 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.t94 DVDD.t75 DVSS.t33 nfet_06v0 ad=12.999999p pd=50.52u as=12.999999p ps=50.52u w=50u l=0.7u
X146 DVSS.t32 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.t95 DVDD.t74 DVSS.t31 nfet_06v0 ad=12.999999p pd=50.52u as=12.999999p ps=50.52u w=50u l=0.7u
X147 DVSS.t30 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.t96 DVDD.t73 DVSS.t29 nfet_06v0 ad=12.999999p pd=50.52u as=12.999999p ps=50.52u w=50u l=0.7u
R0 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_1.D.n17 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_1.D.t19 47.1029
R1 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_1.D.n6 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_1.D.t7 47.1029
R2 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_1.D.n4 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_1.D.t11 47.1029
R3 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_1.D.n2 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_1.D.t24 47.1029
R4 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_1.D.n17 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_1.D.t18 38.0648
R5 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_1.D.n18 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_1.D.t28 38.0648
R6 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_1.D.n19 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_1.D.t16 38.0648
R7 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_1.D.n20 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_1.D.t8 38.0648
R8 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_1.D.n21 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_1.D.t30 38.0648
R9 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_1.D.n22 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_1.D.t26 38.0648
R10 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_1.D.n23 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_1.D.t6 38.0648
R11 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_1.D.n24 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_1.D.t5 38.0648
R12 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_1.D.n25 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_1.D.t17 38.0648
R13 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_1.D.n26 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_1.D.t13 38.0648
R14 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_1.D.n27 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_1.D.t33 38.0648
R15 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_1.D.n6 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_1.D.t21 38.0648
R16 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_1.D.n7 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_1.D.t31 38.0648
R17 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_1.D.n8 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_1.D.t9 38.0648
R18 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_1.D.n9 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_1.D.t20 38.0648
R19 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_1.D.n10 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_1.D.t27 38.0648
R20 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_1.D.n11 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_1.D.t4 38.0648
R21 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_1.D.n12 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_1.D.t12 38.0648
R22 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_1.D.n13 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_1.D.t25 38.0648
R23 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_1.D.n14 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_1.D.t29 38.0648
R24 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_1.D.n15 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_1.D.t14 38.0648
R25 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_1.D.n16 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_1.D.t15 38.0648
R26 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_1.D.n4 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_1.D.t10 38.0648
R27 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_1.D.n5 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_1.D.t23 38.0648
R28 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_1.D.n2 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_1.D.t32 38.0648
R29 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_1.D.n3 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_1.D.t22 38.0648
R30 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_1.D.n18 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_1.D.n17 9.0386
R31 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_1.D.n19 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_1.D.n18 9.0386
R32 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_1.D.n20 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_1.D.n19 9.0386
R33 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_1.D.n21 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_1.D.n20 9.0386
R34 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_1.D.n22 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_1.D.n21 9.0386
R35 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_1.D.n23 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_1.D.n22 9.0386
R36 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_1.D.n24 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_1.D.n23 9.0386
R37 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_1.D.n25 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_1.D.n24 9.0386
R38 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_1.D.n26 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_1.D.n25 9.0386
R39 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_1.D.n27 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_1.D.n26 9.0386
R40 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_1.D.n7 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_1.D.n6 9.0386
R41 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_1.D.n8 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_1.D.n7 9.0386
R42 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_1.D.n9 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_1.D.n8 9.0386
R43 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_1.D.n10 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_1.D.n9 9.0386
R44 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_1.D.n11 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_1.D.n10 9.0386
R45 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_1.D.n12 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_1.D.n11 9.0386
R46 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_1.D.n13 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_1.D.n12 9.0386
R47 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_1.D.n14 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_1.D.n13 9.0386
R48 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_1.D.n15 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_1.D.n14 9.0386
R49 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_1.D.n16 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_1.D.n15 9.0386
R50 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_1.D.n5 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_1.D.n4 9.0386
R51 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_1.D.n3 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_1.D.n2 9.0386
R52 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_1.D.n1 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_1.D.n16 4.51955
R53 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_1.D.n1 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_1.D.n27 4.51955
R54 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_1.D.n0 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_1.D.n3 4.51955
R55 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_1.D.n0 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_1.D.n5 4.51955
R56 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_1.D.n1 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_1.D.t3 2.87695
R57 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_1.D.n1 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_1.D.n0 2.37212
R58 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_1.D.t2 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_1.D.t0 1.95734
R59 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_1.D.t3 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_1.D.t1 1.87633
R60 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_1.D.t2 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_1.D.n1 1.56603
R61 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n246 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.t37 273.524
R62 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.t37 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n245 273.524
R63 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n227 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.t70 273.524
R64 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.t70 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n226 273.524
R65 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.t47 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n112 273.524
R66 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n113 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.t47 273.524
R67 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n131 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.t90 273.524
R68 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.t90 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n130 273.524
R69 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n151 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.t30 273.524
R70 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.t30 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n150 273.524
R71 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.t69 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n168 273.524
R72 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n169 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.t69 273.524
R73 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.t92 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n189 273.524
R74 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n190 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.t92 273.524
R75 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n208 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.t75 273.524
R76 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.t75 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n207 273.524
R77 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n226 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.t32 263.844
R78 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n227 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.t32 263.844
R79 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n225 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.t63 263.844
R80 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n228 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.t63 263.844
R81 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n224 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.t20 263.844
R82 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n229 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.t20 263.844
R83 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n223 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.t54 263.844
R84 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n230 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.t54 263.844
R85 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n222 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.t94 263.844
R86 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n231 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.t94 263.844
R87 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n221 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.t53 263.844
R88 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n232 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.t53 263.844
R89 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n220 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.t82 263.844
R90 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n233 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.t82 263.844
R91 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n219 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.t41 263.844
R92 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n234 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.t41 263.844
R93 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.t73 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n218 263.844
R94 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n235 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.t73 263.844
R95 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n254 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.t34 263.844
R96 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n237 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.t34 263.844
R97 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n253 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.t88 263.844
R98 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n238 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.t88 263.844
R99 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n252 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.t26 263.844
R100 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n239 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.t26 263.844
R101 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n251 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.t80 263.844
R102 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n240 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.t80 263.844
R103 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n250 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.t18 263.844
R104 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n241 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.t18 263.844
R105 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n249 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.t56 263.844
R106 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n242 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.t56 263.844
R107 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n248 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.t31 263.844
R108 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n243 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.t31 263.844
R109 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n247 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.t46 263.844
R110 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n244 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.t46 263.844
R111 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n246 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.t25 263.844
R112 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n245 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.t25 263.844
R113 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n130 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.t50 263.844
R114 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n131 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.t50 263.844
R115 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n129 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.t24 263.844
R116 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n132 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.t24 263.844
R117 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n128 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.t61 263.844
R118 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n133 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.t61 263.844
R119 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n127 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.t29 263.844
R120 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n134 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.t29 263.844
R121 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n126 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.t65 263.844
R122 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n135 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.t65 263.844
R123 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n125 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.t96 263.844
R124 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n136 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.t96 263.844
R125 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n124 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.t78 263.844
R126 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n137 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.t78 263.844
R127 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n123 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.t40 263.844
R128 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n138 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.t40 263.844
R129 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n122 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.t86 263.844
R130 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n139 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.t86 263.844
R131 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n104 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.t51 263.844
R132 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n121 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.t51 263.844
R133 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n105 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.t72 263.844
R134 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n120 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.t72 263.844
R135 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n106 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.t57 263.844
R136 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n119 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.t57 263.844
R137 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n107 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.t79 263.844
R138 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n118 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.t79 263.844
R139 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n108 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.t67 263.844
R140 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n117 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.t67 263.844
R141 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n109 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.t93 263.844
R142 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n116 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.t93 263.844
R143 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n110 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.t52 263.844
R144 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n115 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.t52 263.844
R145 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n111 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.t36 263.844
R146 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n114 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.t36 263.844
R147 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n112 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.t62 263.844
R148 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n113 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.t62 263.844
R149 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n169 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.t19 263.844
R150 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n168 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.t19 263.844
R151 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n170 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.t81 263.844
R152 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n167 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.t81 263.844
R153 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n171 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.t27 263.844
R154 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n166 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.t27 263.844
R155 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n172 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.t64 263.844
R156 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n165 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.t64 263.844
R157 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n173 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.t49 263.844
R158 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n164 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.t49 263.844
R159 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n174 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.t74 263.844
R160 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n163 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.t74 263.844
R161 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n175 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.t59 263.844
R162 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n162 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.t59 263.844
R163 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n176 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.t84 263.844
R164 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n161 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.t84 263.844
R165 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n177 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.t45 263.844
R166 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n160 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.t45 263.844
R167 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n159 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.t95 263.844
R168 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n142 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.t95 263.844
R169 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n158 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.t55 263.844
R170 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n143 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.t55 263.844
R171 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n157 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.t22 263.844
R172 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n144 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.t22 263.844
R173 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n156 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.t60 263.844
R174 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n145 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.t60 263.844
R175 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n155 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.t68 263.844
R176 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n146 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.t68 263.844
R177 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n154 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.t35 263.844
R178 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n147 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.t35 263.844
R179 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n153 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.t76 263.844
R180 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n148 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.t76 263.844
R181 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n152 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.t44 263.844
R182 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n149 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.t44 263.844
R183 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n151 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.t87 263.844
R184 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n150 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.t87 263.844
R185 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n207 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.t42 263.844
R186 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n208 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.t42 263.844
R187 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n206 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.t83 263.844
R188 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n209 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.t83 263.844
R189 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n205 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.t48 263.844
R190 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n210 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.t48 263.844
R191 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n204 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.t89 263.844
R192 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n211 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.t89 263.844
R193 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n203 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.t58 263.844
R194 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n212 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.t58 263.844
R195 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n202 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.t21 263.844
R196 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n213 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.t21 263.844
R197 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n201 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.t43 263.844
R198 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n214 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.t43 263.844
R199 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n200 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.t28 263.844
R200 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n215 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.t28 263.844
R201 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n199 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.t71 263.844
R202 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n216 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.t71 263.844
R203 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n181 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.t38 263.844
R204 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n198 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.t38 263.844
R205 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n182 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.t77 263.844
R206 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n197 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.t77 263.844
R207 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n183 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.t23 263.844
R208 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n196 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.t23 263.844
R209 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n184 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.t91 263.844
R210 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n195 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.t91 263.844
R211 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n185 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.t33 263.844
R212 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n194 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.t33 263.844
R213 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n186 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.t17 263.844
R214 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n193 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.t17 263.844
R215 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n187 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.t39 263.844
R216 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n192 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.t39 263.844
R217 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n188 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.t85 263.844
R218 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n191 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.t85 263.844
R219 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n189 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.t66 263.844
R220 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n190 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.t66 263.844
R221 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n228 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n227 9.68093
R222 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n229 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n228 9.68093
R223 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n230 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n229 9.68093
R224 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n231 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n230 9.68093
R225 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n232 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n231 9.68093
R226 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n233 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n232 9.68093
R227 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n234 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n233 9.68093
R228 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n235 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n234 9.68093
R229 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n238 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n237 9.68093
R230 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n239 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n238 9.68093
R231 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n240 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n239 9.68093
R232 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n241 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n240 9.68093
R233 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n242 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n241 9.68093
R234 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n243 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n242 9.68093
R235 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n244 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n243 9.68093
R236 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n245 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n244 9.68093
R237 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n226 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n225 9.68093
R238 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n225 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n224 9.68093
R239 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n224 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n223 9.68093
R240 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n223 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n222 9.68093
R241 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n222 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n221 9.68093
R242 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n221 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n220 9.68093
R243 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n220 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n219 9.68093
R244 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n219 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n218 9.68093
R245 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n254 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n253 9.68093
R246 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n253 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n252 9.68093
R247 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n252 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n251 9.68093
R248 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n251 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n250 9.68093
R249 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n250 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n249 9.68093
R250 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n249 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n248 9.68093
R251 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n248 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n247 9.68093
R252 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n247 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n246 9.68093
R253 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n114 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n113 9.68093
R254 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n115 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n114 9.68093
R255 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n116 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n115 9.68093
R256 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n117 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n116 9.68093
R257 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n118 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n117 9.68093
R258 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n119 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n118 9.68093
R259 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n120 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n119 9.68093
R260 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n121 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n120 9.68093
R261 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n139 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n138 9.68093
R262 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n138 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n137 9.68093
R263 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n137 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n136 9.68093
R264 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n136 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n135 9.68093
R265 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n135 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n134 9.68093
R266 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n134 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n133 9.68093
R267 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n133 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n132 9.68093
R268 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n132 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n131 9.68093
R269 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n112 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n111 9.68093
R270 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n111 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n110 9.68093
R271 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n110 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n109 9.68093
R272 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n109 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n108 9.68093
R273 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n108 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n107 9.68093
R274 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n107 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n106 9.68093
R275 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n106 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n105 9.68093
R276 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n105 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n104 9.68093
R277 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n123 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n122 9.68093
R278 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n124 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n123 9.68093
R279 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n125 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n124 9.68093
R280 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n126 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n125 9.68093
R281 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n127 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n126 9.68093
R282 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n128 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n127 9.68093
R283 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n129 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n128 9.68093
R284 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n130 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n129 9.68093
R285 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n150 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n149 9.68093
R286 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n149 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n148 9.68093
R287 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n148 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n147 9.68093
R288 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n147 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n146 9.68093
R289 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n146 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n145 9.68093
R290 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n145 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n144 9.68093
R291 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n144 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n143 9.68093
R292 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n143 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n142 9.68093
R293 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n161 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n160 9.68093
R294 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n162 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n161 9.68093
R295 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n163 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n162 9.68093
R296 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n164 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n163 9.68093
R297 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n165 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n164 9.68093
R298 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n166 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n165 9.68093
R299 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n167 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n166 9.68093
R300 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n168 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n167 9.68093
R301 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n152 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n151 9.68093
R302 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n153 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n152 9.68093
R303 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n154 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n153 9.68093
R304 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n155 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n154 9.68093
R305 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n156 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n155 9.68093
R306 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n157 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n156 9.68093
R307 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n158 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n157 9.68093
R308 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n159 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n158 9.68093
R309 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n177 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n176 9.68093
R310 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n176 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n175 9.68093
R311 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n175 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n174 9.68093
R312 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n174 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n173 9.68093
R313 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n173 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n172 9.68093
R314 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n172 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n171 9.68093
R315 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n171 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n170 9.68093
R316 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n170 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n169 9.68093
R317 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n191 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n190 9.68093
R318 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n192 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n191 9.68093
R319 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n193 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n192 9.68093
R320 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n194 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n193 9.68093
R321 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n195 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n194 9.68093
R322 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n196 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n195 9.68093
R323 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n197 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n196 9.68093
R324 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n198 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n197 9.68093
R325 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n216 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n215 9.68093
R326 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n215 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n214 9.68093
R327 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n214 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n213 9.68093
R328 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n213 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n212 9.68093
R329 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n212 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n211 9.68093
R330 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n211 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n210 9.68093
R331 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n210 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n209 9.68093
R332 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n209 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n208 9.68093
R333 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n189 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n188 9.68093
R334 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n188 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n187 9.68093
R335 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n187 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n186 9.68093
R336 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n186 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n185 9.68093
R337 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n185 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n184 9.68093
R338 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n184 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n183 9.68093
R339 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n183 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n182 9.68093
R340 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n182 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n181 9.68093
R341 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n200 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n199 9.68093
R342 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n201 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n200 9.68093
R343 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n202 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n201 9.68093
R344 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n203 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n202 9.68093
R345 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n204 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n203 9.68093
R346 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n205 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n204 9.68093
R347 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n206 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n205 9.68093
R348 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n207 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n206 9.68093
R349 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n236 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n235 4.84072
R350 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n237 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n236 4.84072
R351 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n7 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n218 4.84072
R352 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n7 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n254 4.84072
R353 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n140 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n121 4.84072
R354 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n140 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n139 4.84072
R355 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n104 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n103 4.84072
R356 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n122 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n103 4.84072
R357 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n142 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n141 4.84072
R358 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n160 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n141 4.84072
R359 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n178 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n159 4.84072
R360 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n178 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n177 4.84072
R361 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n217 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n198 4.84072
R362 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n217 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n216 4.84072
R363 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n181 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n180 4.84072
R364 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n199 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n180 4.84072
R365 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n85 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n0 5.09602
R366 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n1 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n62 5.10883
R367 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n40 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n4 5.09332
R368 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n7 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n12 4.98233
R369 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n257 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n84 4.33869
R370 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n260 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n91 4.14642
R371 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n257 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n0 4.13574
R372 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n17 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n15 0.10684
R373 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n16 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n14 0.226809
R374 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n13 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n11 0.226809
R375 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n12 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n10 1.11398
R376 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n18 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n89 1.11398
R377 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n19 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n20 0.534346
R378 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n21 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n22 0.534346
R379 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n23 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n24 0.534346
R380 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n25 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n26 0.534346
R381 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n27 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n28 0.534346
R382 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n29 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n30 0.534346
R383 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n31 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n32 0.534346
R384 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n33 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n34 0.534346
R385 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n35 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n36 0.534346
R386 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n37 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n38 0.534346
R387 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n39 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n40 0.73001
R388 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n88 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n87 1.11398
R389 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n43 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n42 0.534346
R390 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n45 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n41 0.534346
R391 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n47 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n44 0.534346
R392 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n49 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n46 0.534346
R393 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n51 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n48 0.534346
R394 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n53 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n50 0.534346
R395 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n55 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n52 0.534346
R396 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n57 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n54 0.534346
R397 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n59 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n56 0.534346
R398 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n61 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n58 0.534346
R399 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n62 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n60 0.73001
R400 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n63 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n86 1.11398
R401 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n64 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n65 0.534346
R402 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n66 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n67 0.534346
R403 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n68 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n69 0.534346
R404 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n70 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n71 0.534346
R405 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n72 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n73 0.534346
R406 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n74 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n75 0.534346
R407 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n76 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n77 0.534346
R408 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n78 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n79 0.534346
R409 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n80 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n81 0.534346
R410 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n82 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n83 0.534346
R411 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n84 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n85 0.73001
R412 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.t5 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.t11 1.8765
R413 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n91 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.t14 1.29859
R414 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n90 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.t10 1.29859
R415 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n92 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.t12 1.29859
R416 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n95 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.t16 1.29859
R417 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n94 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.t15 1.29859
R418 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n96 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.t8 1.29859
R419 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n97 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.t9 1.29859
R420 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n98 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.t7 1.29859
R421 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n99 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.t13 1.29859
R422 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n259 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n102 1.16318
R423 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n102 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n257 0.97572
R424 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n93 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n100 0.931354
R425 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n101 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.t1 0.912457
R426 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n261 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.t0 0.912457
R427 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n260 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n259 0.578395
R428 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n91 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n90 0.578395
R429 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n90 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n92 0.578395
R430 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n92 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n93 0.578395
R431 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n93 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n95 0.578395
R432 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n95 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n94 0.578395
R433 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n94 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n96 0.578395
R434 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n96 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n97 0.578395
R435 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n97 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n98 0.578395
R436 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n98 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n99 0.578395
R437 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n99 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.t5 0.578395
R438 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n2 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n1 0.620373
R439 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n5 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n4 0.630944
R440 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n63 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n60 0.5045
R441 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n87 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n39 0.5045
R442 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n18 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n10 0.5045
R443 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n259 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n101 0.467486
R444 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n261 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n260 0.467486
R445 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n102 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n258 0.467055
R446 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n100 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.t6 0.3645
R447 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n100 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.t4 0.3645
R448 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n258 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.t3 0.3281
R449 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n258 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.t2 0.3281
R450 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n17 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n7 6.11209
R451 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n101 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D 0.149031
R452 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n261 0.149031
R453 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n11 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n10 0.229028
R454 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n256 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n103 0.0821327
R455 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n179 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n178 0.0821327
R456 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n255 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n180 0.0821327
R457 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n83 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n85 0.169667
R458 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n81 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n83 0.192757
R459 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n79 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n81 0.192757
R460 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n77 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n79 0.192757
R461 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n75 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n77 0.192757
R462 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n75 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n256 0.0723285
R463 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n73 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n256 0.120928
R464 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n71 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n73 0.192757
R465 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n69 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n71 0.192757
R466 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n67 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n69 0.192757
R467 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n65 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n67 0.192757
R468 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n65 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n86 0.145469
R469 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n2 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n0 0.188574
R470 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n3 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n2 0.150067
R471 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n3 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n140 0.191209
R472 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n86 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n3 5.29016
R473 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n61 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n62 0.169667
R474 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n59 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n61 0.192757
R475 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n57 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n59 0.192757
R476 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n55 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n57 0.192757
R477 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n53 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n55 0.192757
R478 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n179 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n53 0.0723285
R479 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n51 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n179 0.120928
R480 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n49 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n51 0.192757
R481 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n47 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n49 0.192757
R482 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n45 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n47 0.192757
R483 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n43 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n45 0.192757
R484 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n88 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n43 0.145469
R485 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n5 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n1 0.221781
R486 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n6 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n5 0.102099
R487 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n6 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n141 0.168375
R488 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n88 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n6 5.31608
R489 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n38 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n40 0.169667
R490 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n36 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n38 0.192757
R491 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n34 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n36 0.192757
R492 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n32 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n34 0.192757
R493 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n30 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n32 0.192757
R494 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n30 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n255 0.0723285
R495 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n28 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n255 0.120928
R496 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n26 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n28 0.192757
R497 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n24 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n26 0.192757
R498 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n22 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n24 0.192757
R499 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n20 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n22 0.192757
R500 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n20 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n89 0.145469
R501 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n8 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n7 1.04643
R502 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n16 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n13 0.385014
R503 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n16 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n15 0.24315
R504 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n84 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n82 0.1949
R505 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n82 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n80 0.1949
R506 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n80 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n78 0.1949
R507 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n78 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n76 0.1949
R508 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n76 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n74 0.1949
R509 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n74 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n72 0.1949
R510 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n72 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n70 0.1949
R511 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n70 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n68 0.1949
R512 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n68 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n66 0.1949
R513 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n66 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n64 0.1949
R514 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n64 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n63 0.1949
R515 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n58 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n60 0.1949
R516 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n56 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n58 0.1949
R517 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n54 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n56 0.1949
R518 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n52 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n54 0.1949
R519 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n50 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n52 0.1949
R520 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n48 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n50 0.1949
R521 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n46 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n48 0.1949
R522 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n44 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n46 0.1949
R523 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n41 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n44 0.1949
R524 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n42 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n41 0.1949
R525 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n87 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n42 0.1949
R526 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n39 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n37 0.1949
R527 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n37 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n35 0.1949
R528 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n35 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n33 0.1949
R529 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n33 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n31 0.1949
R530 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n31 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n29 0.1949
R531 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n29 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n27 0.1949
R532 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n27 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n25 0.1949
R533 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n25 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n23 0.1949
R534 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n23 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n21 0.1949
R535 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n21 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n19 0.1949
R536 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n19 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n18 0.1949
R537 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n14 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n11 0.360357
R538 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n17 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n14 0.482631
R539 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n13 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n12 0.337726
R540 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n236 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n15 0.155273
R541 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n8 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n4 0.188574
R542 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n9 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n8 0.150067
R543 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n9 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n217 0.191209
R544 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n89 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n9 5.29016
R545 DVDD.n16402 DVDD.n16401 33140.3
R546 DVDD.n16403 DVDD.n16402 33140.3
R547 DVDD.n16403 DVDD.n2292 33140.3
R548 DVDD.n16401 DVDD.n2292 33140.3
R549 DVDD.n21015 DVDD.n18821 12187
R550 DVDD.n21017 DVDD.n18821 12187
R551 DVDD.n21017 DVDD.n21016 12187
R552 DVDD.n21016 DVDD.n21015 12187
R553 DVDD.n4372 DVDD.t54 285.2
R554 DVDD.t0 DVDD.n4353 285.18
R555 DVDD.t34 DVDD.t153 270.481
R556 DVDD.t54 DVDD.t30 158.649
R557 DVDD.t30 DVDD.t16 158.649
R558 DVDD.t16 DVDD.t50 158.649
R559 DVDD.t50 DVDD.t32 158.649
R560 DVDD.t32 DVDD.t24 158.649
R561 DVDD.t24 DVDD.t60 158.649
R562 DVDD.t60 DVDD.t48 158.649
R563 DVDD.t48 DVDD.t28 158.649
R564 DVDD.t28 DVDD.t20 158.649
R565 DVDD.t20 DVDD.t44 158.649
R566 DVDD.t44 DVDD.t42 158.649
R567 DVDD.t42 DVDD.t14 158.649
R568 DVDD.t14 DVDD.t46 158.649
R569 DVDD.t46 DVDD.t38 158.649
R570 DVDD.t38 DVDD.t58 158.649
R571 DVDD.t56 DVDD.t26 158.649
R572 DVDD.t26 DVDD.t18 158.649
R573 DVDD.t18 DVDD.t52 158.649
R574 DVDD.t52 DVDD.t40 158.649
R575 DVDD.t40 DVDD.t22 158.649
R576 DVDD.t22 DVDD.t36 158.649
R577 DVDD.t36 DVDD.t34 158.649
R578 DVDD.t153 DVDD.t10 158.649
R579 DVDD.t10 DVDD.t8 158.649
R580 DVDD.t8 DVDD.t4 158.649
R581 DVDD.t4 DVDD.t2 158.649
R582 DVDD.t2 DVDD.t6 158.649
R583 DVDD.t6 DVDD.t0 158.649
R584 DVDD.n4354 DVDD.t56 102.731
R585 DVDD.t58 DVDD.n4354 55.9173
R586 DVDD.n21502 DVDD.n21501 29.1205
R587 DVDD.n19409 DVDD.n19218 11.1794
R588 DVDD.n21497 DVDD.n18560 11.1794
R589 DVDD DVDD.t64 11.0117
R590 DVDD.n19413 DVDD.n19412 8.60804
R591 DVDD.n21496 DVDD.n18621 7.6305
R592 DVDD.n21499 DVDD.n21498 7.6305
R593 DVDD.n19409 DVDD.n19408 7.54986
R594 DVDD.n19402 DVDD.n19338 7.54986
R595 DVDD.n19402 DVDD.n19401 7.54986
R596 DVDD.n19400 DVDD.n19342 7.54986
R597 DVDD.n19394 DVDD.n19342 7.54986
R598 DVDD.n19393 DVDD.n19392 7.54986
R599 DVDD.n19386 DVDD.n19352 7.54986
R600 DVDD.n19386 DVDD.n19385 7.54986
R601 DVDD.n19384 DVDD.n19356 7.54986
R602 DVDD.n19378 DVDD.n19356 7.54986
R603 DVDD.n21276 DVDD.n18650 7.54986
R604 DVDD.n21283 DVDD.n18646 7.54986
R605 DVDD.n21283 DVDD.n21282 7.54986
R606 DVDD.n21289 DVDD.n18639 7.54986
R607 DVDD.n21295 DVDD.n18639 7.54986
R608 DVDD.n21301 DVDD.n18635 7.54986
R609 DVDD.n21308 DVDD.n18631 7.54986
R610 DVDD.n21308 DVDD.n21307 7.54986
R611 DVDD.n21314 DVDD.n18624 7.54986
R612 DVDD.n21321 DVDD.n18624 7.54986
R613 DVDD.n21497 DVDD.n18619 7.54986
R614 DVDD.n19333 DVDD.n19332 7.2805
R615 DVDD.n19330 DVDD.n19318 7.2805
R616 DVDD.n19326 DVDD.n19325 7.2805
R617 DVDD.n19323 DVDD.n19321 7.2805
R618 DVDD.n19630 DVDD.n19629 7.2805
R619 DVDD.n19627 DVDD.n19219 7.2805
R620 DVDD.n19623 DVDD.n19622 7.2805
R621 DVDD.n19620 DVDD.n19222 7.2805
R622 DVDD.n19616 DVDD.n19615 7.2805
R623 DVDD.n19613 DVDD.n19225 7.2805
R624 DVDD.n19609 DVDD.n19608 7.2805
R625 DVDD.n19606 DVDD.n19228 7.2805
R626 DVDD.n19602 DVDD.n19601 7.2805
R627 DVDD.n19599 DVDD.n19231 7.2805
R628 DVDD.n19595 DVDD.n19594 7.2805
R629 DVDD.n19592 DVDD.n19234 7.2805
R630 DVDD.n19588 DVDD.n19587 7.2805
R631 DVDD.n19585 DVDD.n19239 7.2805
R632 DVDD.n19581 DVDD.n19580 7.2805
R633 DVDD.n19578 DVDD.n19242 7.2805
R634 DVDD.n19574 DVDD.n19573 7.2805
R635 DVDD.n19571 DVDD.n19245 7.2805
R636 DVDD.n19567 DVDD.n19566 7.2805
R637 DVDD.n19564 DVDD.n19248 7.2805
R638 DVDD.n19560 DVDD.n19559 7.2805
R639 DVDD.n19557 DVDD.n19251 7.2805
R640 DVDD.n19551 DVDD.n19550 7.2805
R641 DVDD.n19548 DVDD.n19254 7.2805
R642 DVDD.n19544 DVDD.n19543 7.2805
R643 DVDD.n19541 DVDD.n19257 7.2805
R644 DVDD.n19537 DVDD.n19536 7.2805
R645 DVDD.n19534 DVDD.n19260 7.2805
R646 DVDD.n19530 DVDD.n19529 7.2805
R647 DVDD.n19527 DVDD.n19263 7.2805
R648 DVDD.n19523 DVDD.n19522 7.2805
R649 DVDD.n19520 DVDD.n19266 7.2805
R650 DVDD.n19516 DVDD.n19515 7.2805
R651 DVDD.n19513 DVDD.n19269 7.2805
R652 DVDD.n19509 DVDD.n19508 7.2805
R653 DVDD.n19506 DVDD.n19272 7.2805
R654 DVDD.n19500 DVDD.n19499 7.2805
R655 DVDD.n19497 DVDD.n19275 7.2805
R656 DVDD.n19493 DVDD.n19492 7.2805
R657 DVDD.n19490 DVDD.n19278 7.2805
R658 DVDD.n19486 DVDD.n19485 7.2805
R659 DVDD.n19483 DVDD.n19281 7.2805
R660 DVDD.n19479 DVDD.n19478 7.2805
R661 DVDD.n19476 DVDD.n19284 7.2805
R662 DVDD.n19472 DVDD.n19471 7.2805
R663 DVDD.n19469 DVDD.n19287 7.2805
R664 DVDD.n19465 DVDD.n19464 7.2805
R665 DVDD.n19462 DVDD.n19292 7.2805
R666 DVDD.n19458 DVDD.n19457 7.2805
R667 DVDD.n19455 DVDD.n19295 7.2805
R668 DVDD.n19451 DVDD.n19450 7.2805
R669 DVDD.n19448 DVDD.n19298 7.2805
R670 DVDD.n19444 DVDD.n19443 7.2805
R671 DVDD.n19441 DVDD.n19301 7.2805
R672 DVDD.n19437 DVDD.n19436 7.2805
R673 DVDD.n19434 DVDD.n19304 7.2805
R674 DVDD.n19430 DVDD.n19429 7.2805
R675 DVDD.n19427 DVDD.n19307 7.2805
R676 DVDD.n19422 DVDD.n19421 7.2805
R677 DVDD.n19419 DVDD.n19310 7.2805
R678 DVDD.n19415 DVDD.n19414 7.2805
R679 DVDD.n19407 DVDD.n19315 7.2805
R680 DVDD.n19407 DVDD.n19316 7.2805
R681 DVDD.n19403 DVDD.n19316 7.2805
R682 DVDD.n19403 DVDD.n19337 7.2805
R683 DVDD.n19399 DVDD.n19337 7.2805
R684 DVDD.n19399 DVDD.n19343 7.2805
R685 DVDD.n19395 DVDD.n19343 7.2805
R686 DVDD.n19395 DVDD.n19345 7.2805
R687 DVDD.n19391 DVDD.n19345 7.2805
R688 DVDD.n19391 DVDD.n19349 7.2805
R689 DVDD.n19387 DVDD.n19349 7.2805
R690 DVDD.n19387 DVDD.n19351 7.2805
R691 DVDD.n19383 DVDD.n19351 7.2805
R692 DVDD.n19383 DVDD.n19357 7.2805
R693 DVDD.n19379 DVDD.n19357 7.2805
R694 DVDD.n19379 DVDD.n18651 7.2805
R695 DVDD.n21275 DVDD.n18651 7.2805
R696 DVDD.n21275 DVDD.n18645 7.2805
R697 DVDD.n21284 DVDD.n18645 7.2805
R698 DVDD.n21284 DVDD.n18643 7.2805
R699 DVDD.n21288 DVDD.n18643 7.2805
R700 DVDD.n21288 DVDD.n18638 7.2805
R701 DVDD.n21296 DVDD.n18638 7.2805
R702 DVDD.n21296 DVDD.n18636 7.2805
R703 DVDD.n21300 DVDD.n18636 7.2805
R704 DVDD.n21300 DVDD.n18630 7.2805
R705 DVDD.n21309 DVDD.n18630 7.2805
R706 DVDD.n21309 DVDD.n18628 7.2805
R707 DVDD.n21313 DVDD.n18628 7.2805
R708 DVDD.n21313 DVDD.n18623 7.2805
R709 DVDD.n21322 DVDD.n18623 7.2805
R710 DVDD.n21322 DVDD.n18620 7.2805
R711 DVDD.n21496 DVDD.n18620 7.2805
R712 DVDD.n19410 DVDD.n19314 7.2805
R713 DVDD.n19359 DVDD.n19314 7.2805
R714 DVDD.n19359 DVDD.n19339 7.2805
R715 DVDD.n19340 DVDD.n19339 7.2805
R716 DVDD.n19341 DVDD.n19340 7.2805
R717 DVDD.n19364 DVDD.n19341 7.2805
R718 DVDD.n19364 DVDD.n19346 7.2805
R719 DVDD.n19347 DVDD.n19346 7.2805
R720 DVDD.n19348 DVDD.n19347 7.2805
R721 DVDD.n19369 DVDD.n19348 7.2805
R722 DVDD.n19369 DVDD.n19353 7.2805
R723 DVDD.n19354 DVDD.n19353 7.2805
R724 DVDD.n19355 DVDD.n19354 7.2805
R725 DVDD.n19358 DVDD.n19355 7.2805
R726 DVDD.n19377 DVDD.n19358 7.2805
R727 DVDD.n19377 DVDD.n18649 7.2805
R728 DVDD.n21277 DVDD.n18649 7.2805
R729 DVDD.n21277 DVDD.n18647 7.2805
R730 DVDD.n21281 DVDD.n18647 7.2805
R731 DVDD.n21281 DVDD.n18642 7.2805
R732 DVDD.n21290 DVDD.n18642 7.2805
R733 DVDD.n21290 DVDD.n18640 7.2805
R734 DVDD.n21294 DVDD.n18640 7.2805
R735 DVDD.n21294 DVDD.n18634 7.2805
R736 DVDD.n21302 DVDD.n18634 7.2805
R737 DVDD.n21302 DVDD.n18632 7.2805
R738 DVDD.n21306 DVDD.n18632 7.2805
R739 DVDD.n21306 DVDD.n18627 7.2805
R740 DVDD.n21315 DVDD.n18627 7.2805
R741 DVDD.n21315 DVDD.n18625 7.2805
R742 DVDD.n21320 DVDD.n18625 7.2805
R743 DVDD.n21320 DVDD.n18617 7.2805
R744 DVDD.n21498 DVDD.n18617 7.2805
R745 DVDD.n21492 DVDD.n18621 7.2805
R746 DVDD.n21490 DVDD.n21489 7.2805
R747 DVDD.n21487 DVDD.n21327 7.2805
R748 DVDD.n21483 DVDD.n21482 7.2805
R749 DVDD.n21480 DVDD.n21330 7.2805
R750 DVDD.n21476 DVDD.n21475 7.2805
R751 DVDD.n21473 DVDD.n21374 7.2805
R752 DVDD.n21469 DVDD.n21468 7.2805
R753 DVDD.n21466 DVDD.n21377 7.2805
R754 DVDD.n21462 DVDD.n21461 7.2805
R755 DVDD.n21459 DVDD.n21380 7.2805
R756 DVDD.n21455 DVDD.n21454 7.2805
R757 DVDD.n21452 DVDD.n21383 7.2805
R758 DVDD.n21448 DVDD.n21447 7.2805
R759 DVDD.n21445 DVDD.n21386 7.2805
R760 DVDD.n21439 DVDD.n21438 7.2805
R761 DVDD.n21436 DVDD.n21389 7.2805
R762 DVDD.n21432 DVDD.n21431 7.2805
R763 DVDD.n21429 DVDD.n21392 7.2805
R764 DVDD.n21425 DVDD.n21424 7.2805
R765 DVDD.n21422 DVDD.n21395 7.2805
R766 DVDD.n21418 DVDD.n21417 7.2805
R767 DVDD.n21415 DVDD.n21398 7.2805
R768 DVDD.n21411 DVDD.n21410 7.2805
R769 DVDD.n21408 DVDD.n21401 7.2805
R770 DVDD.n21404 DVDD.n21403 7.2805
R771 DVDD.n21643 DVDD.n21642 7.2805
R772 DVDD.n21640 DVDD.n18561 7.2805
R773 DVDD.n21636 DVDD.n21635 7.2805
R774 DVDD.n21633 DVDD.n18564 7.2805
R775 DVDD.n21629 DVDD.n21628 7.2805
R776 DVDD.n21626 DVDD.n18567 7.2805
R777 DVDD.n21622 DVDD.n21621 7.2805
R778 DVDD.n21619 DVDD.n18570 7.2805
R779 DVDD.n21615 DVDD.n21614 7.2805
R780 DVDD.n21612 DVDD.n18573 7.2805
R781 DVDD.n21608 DVDD.n21607 7.2805
R782 DVDD.n21605 DVDD.n18576 7.2805
R783 DVDD.n21601 DVDD.n21600 7.2805
R784 DVDD.n21598 DVDD.n18579 7.2805
R785 DVDD.n21579 DVDD.n21578 7.2805
R786 DVDD.n21576 DVDD.n18582 7.2805
R787 DVDD.n21572 DVDD.n21571 7.2805
R788 DVDD.n21569 DVDD.n18585 7.2805
R789 DVDD.n21565 DVDD.n21564 7.2805
R790 DVDD.n21562 DVDD.n18588 7.2805
R791 DVDD.n21558 DVDD.n21557 7.2805
R792 DVDD.n21555 DVDD.n18591 7.2805
R793 DVDD.n21551 DVDD.n21550 7.2805
R794 DVDD.n21548 DVDD.n18594 7.2805
R795 DVDD.n21544 DVDD.n21543 7.2805
R796 DVDD.n21541 DVDD.n18598 7.2805
R797 DVDD.n21537 DVDD.n21536 7.2805
R798 DVDD.n21534 DVDD.n18601 7.2805
R799 DVDD.n21530 DVDD.n21529 7.2805
R800 DVDD.n21527 DVDD.n18604 7.2805
R801 DVDD.n21523 DVDD.n21522 7.2805
R802 DVDD.n21520 DVDD.n18607 7.2805
R803 DVDD.n21516 DVDD.n21515 7.2805
R804 DVDD.n21513 DVDD.n18610 7.2805
R805 DVDD.n21509 DVDD.n21508 7.2805
R806 DVDD.n21506 DVDD.n18613 7.2805
R807 DVDD.t68 DVDD.n19393 6.96914
R808 DVDD.n21301 DVDD.t12 6.96914
R809 DVDD.n21501 DVDD.n18616 6.39315
R810 DVDD.t72 DVDD.n18650 6.38842
R811 DVDD.n21276 DVDD.t13 6.38842
R812 DVDD.n19411 DVDD.n19410 6.3005
R813 DVDD.n19410 DVDD.n19409 6.3005
R814 DVDD.n19314 DVDD.n19313 6.3005
R815 DVDD.n19408 DVDD.n19314 6.3005
R816 DVDD.n19360 DVDD.n19359 6.3005
R817 DVDD.n19359 DVDD.n19338 6.3005
R818 DVDD.n19361 DVDD.n19339 6.3005
R819 DVDD.n19402 DVDD.n19339 6.3005
R820 DVDD.n19362 DVDD.n19340 6.3005
R821 DVDD.n19401 DVDD.n19340 6.3005
R822 DVDD.n19363 DVDD.n19341 6.3005
R823 DVDD.n19400 DVDD.n19341 6.3005
R824 DVDD.n19365 DVDD.n19364 6.3005
R825 DVDD.n19364 DVDD.n19342 6.3005
R826 DVDD.n19366 DVDD.n19346 6.3005
R827 DVDD.n19394 DVDD.n19346 6.3005
R828 DVDD.n19367 DVDD.n19347 6.3005
R829 DVDD.n19393 DVDD.n19347 6.3005
R830 DVDD.n19368 DVDD.n19348 6.3005
R831 DVDD.n19392 DVDD.n19348 6.3005
R832 DVDD.n19370 DVDD.n19369 6.3005
R833 DVDD.n19369 DVDD.n19352 6.3005
R834 DVDD.n19371 DVDD.n19353 6.3005
R835 DVDD.n19386 DVDD.n19353 6.3005
R836 DVDD.n19372 DVDD.n19354 6.3005
R837 DVDD.n19385 DVDD.n19354 6.3005
R838 DVDD.n19373 DVDD.n19355 6.3005
R839 DVDD.n19384 DVDD.n19355 6.3005
R840 DVDD.n19374 DVDD.n19358 6.3005
R841 DVDD.n19358 DVDD.n19356 6.3005
R842 DVDD.n19377 DVDD.n19376 6.3005
R843 DVDD.n19378 DVDD.n19377 6.3005
R844 DVDD.n19375 DVDD.n18649 6.3005
R845 DVDD.n18650 DVDD.n18649 6.3005
R846 DVDD.n21278 DVDD.n21277 6.3005
R847 DVDD.n21277 DVDD.n21276 6.3005
R848 DVDD.n21279 DVDD.n18647 6.3005
R849 DVDD.n18647 DVDD.n18646 6.3005
R850 DVDD.n21281 DVDD.n21280 6.3005
R851 DVDD.n21283 DVDD.n21281 6.3005
R852 DVDD.n18642 DVDD.n18641 6.3005
R853 DVDD.n21282 DVDD.n18642 6.3005
R854 DVDD.n21291 DVDD.n21290 6.3005
R855 DVDD.n21290 DVDD.n21289 6.3005
R856 DVDD.n21292 DVDD.n18640 6.3005
R857 DVDD.n18640 DVDD.n18639 6.3005
R858 DVDD.n21294 DVDD.n21293 6.3005
R859 DVDD.n21295 DVDD.n21294 6.3005
R860 DVDD.n18634 DVDD.n18633 6.3005
R861 DVDD.n18635 DVDD.n18634 6.3005
R862 DVDD.n21303 DVDD.n21302 6.3005
R863 DVDD.n21302 DVDD.n21301 6.3005
R864 DVDD.n21304 DVDD.n18632 6.3005
R865 DVDD.n18632 DVDD.n18631 6.3005
R866 DVDD.n21306 DVDD.n21305 6.3005
R867 DVDD.n21308 DVDD.n21306 6.3005
R868 DVDD.n18627 DVDD.n18626 6.3005
R869 DVDD.n21307 DVDD.n18627 6.3005
R870 DVDD.n21316 DVDD.n21315 6.3005
R871 DVDD.n21315 DVDD.n21314 6.3005
R872 DVDD.n21317 DVDD.n18625 6.3005
R873 DVDD.n18625 DVDD.n18624 6.3005
R874 DVDD.n21320 DVDD.n21319 6.3005
R875 DVDD.n21321 DVDD.n21320 6.3005
R876 DVDD.n21318 DVDD.n18617 6.3005
R877 DVDD.n18619 DVDD.n18617 6.3005
R878 DVDD.n21498 DVDD.n18618 6.3005
R879 DVDD.n21498 DVDD.n21497 6.3005
R880 DVDD.n21499 DVDD.n18616 6.3005
R881 DVDD.n21502 DVDD.n18560 6.3005
R882 DVDD.n21504 DVDD.n18613 6.3005
R883 DVDD.n21506 DVDD.n21505 6.3005
R884 DVDD.n21508 DVDD.n18611 6.3005
R885 DVDD.n21510 DVDD.n21509 6.3005
R886 DVDD.n21511 DVDD.n18610 6.3005
R887 DVDD.n21513 DVDD.n21512 6.3005
R888 DVDD.n21515 DVDD.n18608 6.3005
R889 DVDD.n21517 DVDD.n21516 6.3005
R890 DVDD.n21518 DVDD.n18607 6.3005
R891 DVDD.n21520 DVDD.n21519 6.3005
R892 DVDD.n21522 DVDD.n18605 6.3005
R893 DVDD.n21524 DVDD.n21523 6.3005
R894 DVDD.n21525 DVDD.n18604 6.3005
R895 DVDD.n21527 DVDD.n21526 6.3005
R896 DVDD.n21529 DVDD.n18602 6.3005
R897 DVDD.n21531 DVDD.n21530 6.3005
R898 DVDD.n21532 DVDD.n18601 6.3005
R899 DVDD.n21534 DVDD.n21533 6.3005
R900 DVDD.n21536 DVDD.n18599 6.3005
R901 DVDD.n21538 DVDD.n21537 6.3005
R902 DVDD.n21539 DVDD.n18598 6.3005
R903 DVDD.n21541 DVDD.n21540 6.3005
R904 DVDD.n21543 DVDD.n18597 6.3005
R905 DVDD.n21545 DVDD.n21544 6.3005
R906 DVDD.n21546 DVDD.n18594 6.3005
R907 DVDD.n21548 DVDD.n21547 6.3005
R908 DVDD.n21550 DVDD.n18592 6.3005
R909 DVDD.n21552 DVDD.n21551 6.3005
R910 DVDD.n21553 DVDD.n18591 6.3005
R911 DVDD.n21555 DVDD.n21554 6.3005
R912 DVDD.n21557 DVDD.n18589 6.3005
R913 DVDD.n21559 DVDD.n21558 6.3005
R914 DVDD.n21560 DVDD.n18588 6.3005
R915 DVDD.n21562 DVDD.n21561 6.3005
R916 DVDD.n21564 DVDD.n18586 6.3005
R917 DVDD.n21566 DVDD.n21565 6.3005
R918 DVDD.n21567 DVDD.n18585 6.3005
R919 DVDD.n21569 DVDD.n21568 6.3005
R920 DVDD.n21571 DVDD.n18583 6.3005
R921 DVDD.n21573 DVDD.n21572 6.3005
R922 DVDD.n21574 DVDD.n18582 6.3005
R923 DVDD.n21576 DVDD.n21575 6.3005
R924 DVDD.n21578 DVDD.n18580 6.3005
R925 DVDD.n21580 DVDD.n21579 6.3005
R926 DVDD.n21581 DVDD.n18579 6.3005
R927 DVDD.n21598 DVDD.n21597 6.3005
R928 DVDD.n21600 DVDD.n18577 6.3005
R929 DVDD.n21602 DVDD.n21601 6.3005
R930 DVDD.n21603 DVDD.n18576 6.3005
R931 DVDD.n21605 DVDD.n21604 6.3005
R932 DVDD.n21607 DVDD.n18574 6.3005
R933 DVDD.n21609 DVDD.n21608 6.3005
R934 DVDD.n21610 DVDD.n18573 6.3005
R935 DVDD.n21612 DVDD.n21611 6.3005
R936 DVDD.n21614 DVDD.n18571 6.3005
R937 DVDD.n21616 DVDD.n21615 6.3005
R938 DVDD.n21617 DVDD.n18570 6.3005
R939 DVDD.n21619 DVDD.n21618 6.3005
R940 DVDD.n21621 DVDD.n18568 6.3005
R941 DVDD.n21623 DVDD.n21622 6.3005
R942 DVDD.n21624 DVDD.n18567 6.3005
R943 DVDD.n21626 DVDD.n21625 6.3005
R944 DVDD.n21628 DVDD.n18565 6.3005
R945 DVDD.n21630 DVDD.n21629 6.3005
R946 DVDD.n21631 DVDD.n18564 6.3005
R947 DVDD.n21633 DVDD.n21632 6.3005
R948 DVDD.n21635 DVDD.n18562 6.3005
R949 DVDD.n21637 DVDD.n21636 6.3005
R950 DVDD.n21638 DVDD.n18561 6.3005
R951 DVDD.n21640 DVDD.n21639 6.3005
R952 DVDD.n21642 DVDD.n18558 6.3005
R953 DVDD.n21644 DVDD.n21643 6.3005
R954 DVDD.n21403 DVDD.n18557 6.3005
R955 DVDD.n21405 DVDD.n21404 6.3005
R956 DVDD.n21406 DVDD.n21401 6.3005
R957 DVDD.n21408 DVDD.n21407 6.3005
R958 DVDD.n21410 DVDD.n21399 6.3005
R959 DVDD.n21412 DVDD.n21411 6.3005
R960 DVDD.n21413 DVDD.n21398 6.3005
R961 DVDD.n21415 DVDD.n21414 6.3005
R962 DVDD.n21417 DVDD.n21396 6.3005
R963 DVDD.n21419 DVDD.n21418 6.3005
R964 DVDD.n21420 DVDD.n21395 6.3005
R965 DVDD.n21422 DVDD.n21421 6.3005
R966 DVDD.n21424 DVDD.n21393 6.3005
R967 DVDD.n21426 DVDD.n21425 6.3005
R968 DVDD.n21427 DVDD.n21392 6.3005
R969 DVDD.n21429 DVDD.n21428 6.3005
R970 DVDD.n21431 DVDD.n21390 6.3005
R971 DVDD.n21433 DVDD.n21432 6.3005
R972 DVDD.n21434 DVDD.n21389 6.3005
R973 DVDD.n21436 DVDD.n21435 6.3005
R974 DVDD.n21438 DVDD.n21387 6.3005
R975 DVDD.n21440 DVDD.n21439 6.3005
R976 DVDD.n21443 DVDD.n21386 6.3005
R977 DVDD.n21445 DVDD.n21444 6.3005
R978 DVDD.n21447 DVDD.n21384 6.3005
R979 DVDD.n21449 DVDD.n21448 6.3005
R980 DVDD.n21450 DVDD.n21383 6.3005
R981 DVDD.n21452 DVDD.n21451 6.3005
R982 DVDD.n21454 DVDD.n21381 6.3005
R983 DVDD.n21456 DVDD.n21455 6.3005
R984 DVDD.n21457 DVDD.n21380 6.3005
R985 DVDD.n21459 DVDD.n21458 6.3005
R986 DVDD.n21461 DVDD.n21378 6.3005
R987 DVDD.n21463 DVDD.n21462 6.3005
R988 DVDD.n21464 DVDD.n21377 6.3005
R989 DVDD.n21466 DVDD.n21465 6.3005
R990 DVDD.n21468 DVDD.n21375 6.3005
R991 DVDD.n21470 DVDD.n21469 6.3005
R992 DVDD.n21471 DVDD.n21374 6.3005
R993 DVDD.n21473 DVDD.n21472 6.3005
R994 DVDD.n21475 DVDD.n21372 6.3005
R995 DVDD.n21477 DVDD.n21476 6.3005
R996 DVDD.n21478 DVDD.n21330 6.3005
R997 DVDD.n21480 DVDD.n21479 6.3005
R998 DVDD.n21482 DVDD.n21328 6.3005
R999 DVDD.n21484 DVDD.n21483 6.3005
R1000 DVDD.n21485 DVDD.n21327 6.3005
R1001 DVDD.n21487 DVDD.n21486 6.3005
R1002 DVDD.n21489 DVDD.n21326 6.3005
R1003 DVDD.n21490 DVDD.n21325 6.3005
R1004 DVDD.n21493 DVDD.n21492 6.3005
R1005 DVDD.n21494 DVDD.n18621 6.3005
R1006 DVDD.n18621 DVDD.n18560 6.3005
R1007 DVDD.n21496 DVDD.n21495 6.3005
R1008 DVDD.n21497 DVDD.n21496 6.3005
R1009 DVDD.n21324 DVDD.n18620 6.3005
R1010 DVDD.n18620 DVDD.n18619 6.3005
R1011 DVDD.n21323 DVDD.n21322 6.3005
R1012 DVDD.n21322 DVDD.n21321 6.3005
R1013 DVDD.n18623 DVDD.n18622 6.3005
R1014 DVDD.n18624 DVDD.n18623 6.3005
R1015 DVDD.n21313 DVDD.n21312 6.3005
R1016 DVDD.n21314 DVDD.n21313 6.3005
R1017 DVDD.n21311 DVDD.n18628 6.3005
R1018 DVDD.n21307 DVDD.n18628 6.3005
R1019 DVDD.n21310 DVDD.n21309 6.3005
R1020 DVDD.n21309 DVDD.n21308 6.3005
R1021 DVDD.n18630 DVDD.n18629 6.3005
R1022 DVDD.n18631 DVDD.n18630 6.3005
R1023 DVDD.n21300 DVDD.n21299 6.3005
R1024 DVDD.n21301 DVDD.n21300 6.3005
R1025 DVDD.n21298 DVDD.n18636 6.3005
R1026 DVDD.n18636 DVDD.n18635 6.3005
R1027 DVDD.n21297 DVDD.n21296 6.3005
R1028 DVDD.n21296 DVDD.n21295 6.3005
R1029 DVDD.n18638 DVDD.n18637 6.3005
R1030 DVDD.n18639 DVDD.n18638 6.3005
R1031 DVDD.n21288 DVDD.n21287 6.3005
R1032 DVDD.n21289 DVDD.n21288 6.3005
R1033 DVDD.n21286 DVDD.n18643 6.3005
R1034 DVDD.n21282 DVDD.n18643 6.3005
R1035 DVDD.n21285 DVDD.n21284 6.3005
R1036 DVDD.n21284 DVDD.n21283 6.3005
R1037 DVDD.n18645 DVDD.n18644 6.3005
R1038 DVDD.n18646 DVDD.n18645 6.3005
R1039 DVDD.n21275 DVDD.n21274 6.3005
R1040 DVDD.n21276 DVDD.n21275 6.3005
R1041 DVDD.n18652 DVDD.n18651 6.3005
R1042 DVDD.n18651 DVDD.n18650 6.3005
R1043 DVDD.n19380 DVDD.n19379 6.3005
R1044 DVDD.n19379 DVDD.n19378 6.3005
R1045 DVDD.n19381 DVDD.n19357 6.3005
R1046 DVDD.n19357 DVDD.n19356 6.3005
R1047 DVDD.n19383 DVDD.n19382 6.3005
R1048 DVDD.n19384 DVDD.n19383 6.3005
R1049 DVDD.n19351 DVDD.n19350 6.3005
R1050 DVDD.n19385 DVDD.n19351 6.3005
R1051 DVDD.n19388 DVDD.n19387 6.3005
R1052 DVDD.n19387 DVDD.n19386 6.3005
R1053 DVDD.n19389 DVDD.n19349 6.3005
R1054 DVDD.n19352 DVDD.n19349 6.3005
R1055 DVDD.n19391 DVDD.n19390 6.3005
R1056 DVDD.n19392 DVDD.n19391 6.3005
R1057 DVDD.n19345 DVDD.n19344 6.3005
R1058 DVDD.n19393 DVDD.n19345 6.3005
R1059 DVDD.n19396 DVDD.n19395 6.3005
R1060 DVDD.n19395 DVDD.n19394 6.3005
R1061 DVDD.n19397 DVDD.n19343 6.3005
R1062 DVDD.n19343 DVDD.n19342 6.3005
R1063 DVDD.n19399 DVDD.n19398 6.3005
R1064 DVDD.n19400 DVDD.n19399 6.3005
R1065 DVDD.n19337 DVDD.n19336 6.3005
R1066 DVDD.n19401 DVDD.n19337 6.3005
R1067 DVDD.n19404 DVDD.n19403 6.3005
R1068 DVDD.n19403 DVDD.n19402 6.3005
R1069 DVDD.n19405 DVDD.n19316 6.3005
R1070 DVDD.n19338 DVDD.n19316 6.3005
R1071 DVDD.n19407 DVDD.n19406 6.3005
R1072 DVDD.n19408 DVDD.n19407 6.3005
R1073 DVDD.n19335 DVDD.n19315 6.3005
R1074 DVDD.n19409 DVDD.n19315 6.3005
R1075 DVDD.n19414 DVDD.n19311 6.3005
R1076 DVDD.n19416 DVDD.n19415 6.3005
R1077 DVDD.n19417 DVDD.n19310 6.3005
R1078 DVDD.n19419 DVDD.n19418 6.3005
R1079 DVDD.n19421 DVDD.n19308 6.3005
R1080 DVDD.n19423 DVDD.n19422 6.3005
R1081 DVDD.n19424 DVDD.n19307 6.3005
R1082 DVDD.n19427 DVDD.n19426 6.3005
R1083 DVDD.n19429 DVDD.n19305 6.3005
R1084 DVDD.n19431 DVDD.n19430 6.3005
R1085 DVDD.n19432 DVDD.n19304 6.3005
R1086 DVDD.n19434 DVDD.n19433 6.3005
R1087 DVDD.n19436 DVDD.n19302 6.3005
R1088 DVDD.n19438 DVDD.n19437 6.3005
R1089 DVDD.n19439 DVDD.n19301 6.3005
R1090 DVDD.n19441 DVDD.n19440 6.3005
R1091 DVDD.n19443 DVDD.n19299 6.3005
R1092 DVDD.n19445 DVDD.n19444 6.3005
R1093 DVDD.n19446 DVDD.n19298 6.3005
R1094 DVDD.n19448 DVDD.n19447 6.3005
R1095 DVDD.n19450 DVDD.n19296 6.3005
R1096 DVDD.n19452 DVDD.n19451 6.3005
R1097 DVDD.n19453 DVDD.n19295 6.3005
R1098 DVDD.n19455 DVDD.n19454 6.3005
R1099 DVDD.n19457 DVDD.n19293 6.3005
R1100 DVDD.n19459 DVDD.n19458 6.3005
R1101 DVDD.n19460 DVDD.n19292 6.3005
R1102 DVDD.n19462 DVDD.n19461 6.3005
R1103 DVDD.n19464 DVDD.n19291 6.3005
R1104 DVDD.n19466 DVDD.n19465 6.3005
R1105 DVDD.n19467 DVDD.n19287 6.3005
R1106 DVDD.n19469 DVDD.n19468 6.3005
R1107 DVDD.n19471 DVDD.n19285 6.3005
R1108 DVDD.n19473 DVDD.n19472 6.3005
R1109 DVDD.n19474 DVDD.n19284 6.3005
R1110 DVDD.n19476 DVDD.n19475 6.3005
R1111 DVDD.n19478 DVDD.n19282 6.3005
R1112 DVDD.n19480 DVDD.n19479 6.3005
R1113 DVDD.n19481 DVDD.n19281 6.3005
R1114 DVDD.n19483 DVDD.n19482 6.3005
R1115 DVDD.n19485 DVDD.n19279 6.3005
R1116 DVDD.n19487 DVDD.n19486 6.3005
R1117 DVDD.n19488 DVDD.n19278 6.3005
R1118 DVDD.n19490 DVDD.n19489 6.3005
R1119 DVDD.n19492 DVDD.n19276 6.3005
R1120 DVDD.n19494 DVDD.n19493 6.3005
R1121 DVDD.n19495 DVDD.n19275 6.3005
R1122 DVDD.n19497 DVDD.n19496 6.3005
R1123 DVDD.n19499 DVDD.n19273 6.3005
R1124 DVDD.n19501 DVDD.n19500 6.3005
R1125 DVDD.n19502 DVDD.n19272 6.3005
R1126 DVDD.n19506 DVDD.n19505 6.3005
R1127 DVDD.n19508 DVDD.n19270 6.3005
R1128 DVDD.n19510 DVDD.n19509 6.3005
R1129 DVDD.n19511 DVDD.n19269 6.3005
R1130 DVDD.n19513 DVDD.n19512 6.3005
R1131 DVDD.n19515 DVDD.n19267 6.3005
R1132 DVDD.n19517 DVDD.n19516 6.3005
R1133 DVDD.n19518 DVDD.n19266 6.3005
R1134 DVDD.n19520 DVDD.n19519 6.3005
R1135 DVDD.n19522 DVDD.n19264 6.3005
R1136 DVDD.n19524 DVDD.n19523 6.3005
R1137 DVDD.n19525 DVDD.n19263 6.3005
R1138 DVDD.n19527 DVDD.n19526 6.3005
R1139 DVDD.n19529 DVDD.n19261 6.3005
R1140 DVDD.n19531 DVDD.n19530 6.3005
R1141 DVDD.n19532 DVDD.n19260 6.3005
R1142 DVDD.n19534 DVDD.n19533 6.3005
R1143 DVDD.n19536 DVDD.n19258 6.3005
R1144 DVDD.n19538 DVDD.n19537 6.3005
R1145 DVDD.n19539 DVDD.n19257 6.3005
R1146 DVDD.n19541 DVDD.n19540 6.3005
R1147 DVDD.n19543 DVDD.n19255 6.3005
R1148 DVDD.n19545 DVDD.n19544 6.3005
R1149 DVDD.n19546 DVDD.n19254 6.3005
R1150 DVDD.n19548 DVDD.n19547 6.3005
R1151 DVDD.n19550 DVDD.n19252 6.3005
R1152 DVDD.n19552 DVDD.n19551 6.3005
R1153 DVDD.n19555 DVDD.n19251 6.3005
R1154 DVDD.n19557 DVDD.n19556 6.3005
R1155 DVDD.n19559 DVDD.n19249 6.3005
R1156 DVDD.n19561 DVDD.n19560 6.3005
R1157 DVDD.n19562 DVDD.n19248 6.3005
R1158 DVDD.n19564 DVDD.n19563 6.3005
R1159 DVDD.n19566 DVDD.n19246 6.3005
R1160 DVDD.n19568 DVDD.n19567 6.3005
R1161 DVDD.n19569 DVDD.n19245 6.3005
R1162 DVDD.n19571 DVDD.n19570 6.3005
R1163 DVDD.n19573 DVDD.n19243 6.3005
R1164 DVDD.n19575 DVDD.n19574 6.3005
R1165 DVDD.n19576 DVDD.n19242 6.3005
R1166 DVDD.n19578 DVDD.n19577 6.3005
R1167 DVDD.n19580 DVDD.n19240 6.3005
R1168 DVDD.n19582 DVDD.n19581 6.3005
R1169 DVDD.n19583 DVDD.n19239 6.3005
R1170 DVDD.n19585 DVDD.n19584 6.3005
R1171 DVDD.n19587 DVDD.n19237 6.3005
R1172 DVDD.n19589 DVDD.n19588 6.3005
R1173 DVDD.n19590 DVDD.n19234 6.3005
R1174 DVDD.n19592 DVDD.n19591 6.3005
R1175 DVDD.n19594 DVDD.n19232 6.3005
R1176 DVDD.n19596 DVDD.n19595 6.3005
R1177 DVDD.n19597 DVDD.n19231 6.3005
R1178 DVDD.n19599 DVDD.n19598 6.3005
R1179 DVDD.n19601 DVDD.n19229 6.3005
R1180 DVDD.n19603 DVDD.n19602 6.3005
R1181 DVDD.n19604 DVDD.n19228 6.3005
R1182 DVDD.n19606 DVDD.n19605 6.3005
R1183 DVDD.n19608 DVDD.n19226 6.3005
R1184 DVDD.n19610 DVDD.n19609 6.3005
R1185 DVDD.n19611 DVDD.n19225 6.3005
R1186 DVDD.n19613 DVDD.n19612 6.3005
R1187 DVDD.n19615 DVDD.n19223 6.3005
R1188 DVDD.n19617 DVDD.n19616 6.3005
R1189 DVDD.n19618 DVDD.n19222 6.3005
R1190 DVDD.n19620 DVDD.n19619 6.3005
R1191 DVDD.n19622 DVDD.n19220 6.3005
R1192 DVDD.n19624 DVDD.n19623 6.3005
R1193 DVDD.n19625 DVDD.n19219 6.3005
R1194 DVDD.n19627 DVDD.n19626 6.3005
R1195 DVDD.n19629 DVDD.n19216 6.3005
R1196 DVDD.n19631 DVDD.n19630 6.3005
R1197 DVDD.n19321 DVDD.n19215 6.3005
R1198 DVDD.n19323 DVDD.n19322 6.3005
R1199 DVDD.n19325 DVDD.n19319 6.3005
R1200 DVDD.n19327 DVDD.n19326 6.3005
R1201 DVDD.n19328 DVDD.n19318 6.3005
R1202 DVDD.n19330 DVDD.n19329 6.3005
R1203 DVDD.n19332 DVDD.n19317 6.3005
R1204 DVDD.n19334 DVDD.n19333 6.3005
R1205 DVDD.n19333 DVDD.n19218 6.3005
R1206 DVDD.n19392 DVDD.t70 5.8077
R1207 DVDD.t71 DVDD.n18635 5.8077
R1208 DVDD.n19408 DVDD.t63 5.22698
R1209 DVDD.t65 DVDD.n18619 5.22698
R1210 DVDD.t62 DVDD.n19400 4.64626
R1211 DVDD.n21307 DVDD.t69 4.64626
R1212 DVDD.n21503 DVDD.n18615 4.60138
R1213 DVDD.n18797 DVDD.n104 4.5005
R1214 DVDD.n21050 DVDD.n104 4.5005
R1215 DVDD.n18794 DVDD.n97 4.5005
R1216 DVDD.n21051 DVDD.n18801 4.5005
R1217 DVDD.n21051 DVDD.n18792 4.5005
R1218 DVDD.n21051 DVDD.n18804 4.5005
R1219 DVDD.n21051 DVDD.n18791 4.5005
R1220 DVDD.n21051 DVDD.n18807 4.5005
R1221 DVDD.n21051 DVDD.n18790 4.5005
R1222 DVDD.n21051 DVDD.n18810 4.5005
R1223 DVDD.n21051 DVDD.n18789 4.5005
R1224 DVDD.n21051 DVDD.n18813 4.5005
R1225 DVDD.n21051 DVDD.n18788 4.5005
R1226 DVDD.n21051 DVDD.n18816 4.5005
R1227 DVDD.n21051 DVDD.n18787 4.5005
R1228 DVDD.n21051 DVDD.n21050 4.5005
R1229 DVDD.n19098 DVDD.n18770 4.5005
R1230 DVDD.n18773 DVDD.n18770 4.5005
R1231 DVDD.n21053 DVDD.n18770 4.5005
R1232 DVDD.n21053 DVDD.n21052 4.5005
R1233 DVDD.n19105 DVDD.n19094 4.5005
R1234 DVDD.n19121 DVDD.n19094 4.5005
R1235 DVDD.n20933 DVDD.n18868 4.5005
R1236 DVDD.n20949 DVDD.n18868 4.5005
R1237 DVDD.n20465 DVDD.n18907 4.5005
R1238 DVDD.n20479 DVDD.n20465 4.5005
R1239 DVDD.n20482 DVDD.n20465 4.5005
R1240 DVDD.n20482 DVDD.n19033 4.5005
R1241 DVDD.n20464 DVDD.n19817 4.5005
R1242 DVDD.n20464 DVDD.n19818 4.5005
R1243 DVDD.n20464 DVDD.n20463 4.5005
R1244 DVDD.n19820 DVDD.n19818 4.5005
R1245 DVDD.n20463 DVDD.n19820 4.5005
R1246 DVDD.n20462 DVDD.n19817 4.5005
R1247 DVDD.n20462 DVDD.n20450 4.5005
R1248 DVDD.n20462 DVDD.n20448 4.5005
R1249 DVDD.n20462 DVDD.n20452 4.5005
R1250 DVDD.n20462 DVDD.n20447 4.5005
R1251 DVDD.n20462 DVDD.n20454 4.5005
R1252 DVDD.n20462 DVDD.n20446 4.5005
R1253 DVDD.n20462 DVDD.n20456 4.5005
R1254 DVDD.n20462 DVDD.n20445 4.5005
R1255 DVDD.n20462 DVDD.n20458 4.5005
R1256 DVDD.n20462 DVDD.n20444 4.5005
R1257 DVDD.n20462 DVDD.n20460 4.5005
R1258 DVDD.n20463 DVDD.n20462 4.5005
R1259 DVDD.n9668 DVDD.n9661 4.5005
R1260 DVDD.n10068 DVDD.n9668 4.5005
R1261 DVDD.n9686 DVDD.n9668 4.5005
R1262 DVDD.n9690 DVDD.n9668 4.5005
R1263 DVDD.n9684 DVDD.n9668 4.5005
R1264 DVDD.n9691 DVDD.n9668 4.5005
R1265 DVDD.n9683 DVDD.n9668 4.5005
R1266 DVDD.n9692 DVDD.n9668 4.5005
R1267 DVDD.n9682 DVDD.n9668 4.5005
R1268 DVDD.n9695 DVDD.n9668 4.5005
R1269 DVDD.n9680 DVDD.n9668 4.5005
R1270 DVDD.n10066 DVDD.n9668 4.5005
R1271 DVDD.n10068 DVDD.n9666 4.5005
R1272 DVDD.n9686 DVDD.n9666 4.5005
R1273 DVDD.n9689 DVDD.n9666 4.5005
R1274 DVDD.n9685 DVDD.n9666 4.5005
R1275 DVDD.n9690 DVDD.n9666 4.5005
R1276 DVDD.n9684 DVDD.n9666 4.5005
R1277 DVDD.n9691 DVDD.n9666 4.5005
R1278 DVDD.n9683 DVDD.n9666 4.5005
R1279 DVDD.n9692 DVDD.n9666 4.5005
R1280 DVDD.n9682 DVDD.n9666 4.5005
R1281 DVDD.n9694 DVDD.n9666 4.5005
R1282 DVDD.n9681 DVDD.n9666 4.5005
R1283 DVDD.n9695 DVDD.n9666 4.5005
R1284 DVDD.n10066 DVDD.n9666 4.5005
R1285 DVDD.n10068 DVDD.n9670 4.5005
R1286 DVDD.n9686 DVDD.n9670 4.5005
R1287 DVDD.n9689 DVDD.n9670 4.5005
R1288 DVDD.n9685 DVDD.n9670 4.5005
R1289 DVDD.n9690 DVDD.n9670 4.5005
R1290 DVDD.n9684 DVDD.n9670 4.5005
R1291 DVDD.n9691 DVDD.n9670 4.5005
R1292 DVDD.n9683 DVDD.n9670 4.5005
R1293 DVDD.n9692 DVDD.n9670 4.5005
R1294 DVDD.n9682 DVDD.n9670 4.5005
R1295 DVDD.n9694 DVDD.n9670 4.5005
R1296 DVDD.n9681 DVDD.n9670 4.5005
R1297 DVDD.n9695 DVDD.n9670 4.5005
R1298 DVDD.n10066 DVDD.n9670 4.5005
R1299 DVDD.n10068 DVDD.n9665 4.5005
R1300 DVDD.n9686 DVDD.n9665 4.5005
R1301 DVDD.n9689 DVDD.n9665 4.5005
R1302 DVDD.n9685 DVDD.n9665 4.5005
R1303 DVDD.n9690 DVDD.n9665 4.5005
R1304 DVDD.n9684 DVDD.n9665 4.5005
R1305 DVDD.n9691 DVDD.n9665 4.5005
R1306 DVDD.n9683 DVDD.n9665 4.5005
R1307 DVDD.n9692 DVDD.n9665 4.5005
R1308 DVDD.n9682 DVDD.n9665 4.5005
R1309 DVDD.n9694 DVDD.n9665 4.5005
R1310 DVDD.n9681 DVDD.n9665 4.5005
R1311 DVDD.n9695 DVDD.n9665 4.5005
R1312 DVDD.n9680 DVDD.n9665 4.5005
R1313 DVDD.n10066 DVDD.n9665 4.5005
R1314 DVDD.n10068 DVDD.n9672 4.5005
R1315 DVDD.n9686 DVDD.n9672 4.5005
R1316 DVDD.n9689 DVDD.n9672 4.5005
R1317 DVDD.n9685 DVDD.n9672 4.5005
R1318 DVDD.n9690 DVDD.n9672 4.5005
R1319 DVDD.n9684 DVDD.n9672 4.5005
R1320 DVDD.n9691 DVDD.n9672 4.5005
R1321 DVDD.n9683 DVDD.n9672 4.5005
R1322 DVDD.n9692 DVDD.n9672 4.5005
R1323 DVDD.n9682 DVDD.n9672 4.5005
R1324 DVDD.n9694 DVDD.n9672 4.5005
R1325 DVDD.n9681 DVDD.n9672 4.5005
R1326 DVDD.n9695 DVDD.n9672 4.5005
R1327 DVDD.n10066 DVDD.n9672 4.5005
R1328 DVDD.n10068 DVDD.n9664 4.5005
R1329 DVDD.n9686 DVDD.n9664 4.5005
R1330 DVDD.n9689 DVDD.n9664 4.5005
R1331 DVDD.n9685 DVDD.n9664 4.5005
R1332 DVDD.n9690 DVDD.n9664 4.5005
R1333 DVDD.n9684 DVDD.n9664 4.5005
R1334 DVDD.n9691 DVDD.n9664 4.5005
R1335 DVDD.n9683 DVDD.n9664 4.5005
R1336 DVDD.n9692 DVDD.n9664 4.5005
R1337 DVDD.n9682 DVDD.n9664 4.5005
R1338 DVDD.n9694 DVDD.n9664 4.5005
R1339 DVDD.n9681 DVDD.n9664 4.5005
R1340 DVDD.n9695 DVDD.n9664 4.5005
R1341 DVDD.n10066 DVDD.n9664 4.5005
R1342 DVDD.n10068 DVDD.n9674 4.5005
R1343 DVDD.n9686 DVDD.n9674 4.5005
R1344 DVDD.n9689 DVDD.n9674 4.5005
R1345 DVDD.n9685 DVDD.n9674 4.5005
R1346 DVDD.n9690 DVDD.n9674 4.5005
R1347 DVDD.n9684 DVDD.n9674 4.5005
R1348 DVDD.n9691 DVDD.n9674 4.5005
R1349 DVDD.n9683 DVDD.n9674 4.5005
R1350 DVDD.n9692 DVDD.n9674 4.5005
R1351 DVDD.n9682 DVDD.n9674 4.5005
R1352 DVDD.n9694 DVDD.n9674 4.5005
R1353 DVDD.n9681 DVDD.n9674 4.5005
R1354 DVDD.n9695 DVDD.n9674 4.5005
R1355 DVDD.n9680 DVDD.n9674 4.5005
R1356 DVDD.n10066 DVDD.n9674 4.5005
R1357 DVDD.n10068 DVDD.n9663 4.5005
R1358 DVDD.n9686 DVDD.n9663 4.5005
R1359 DVDD.n9689 DVDD.n9663 4.5005
R1360 DVDD.n9685 DVDD.n9663 4.5005
R1361 DVDD.n9690 DVDD.n9663 4.5005
R1362 DVDD.n9684 DVDD.n9663 4.5005
R1363 DVDD.n9691 DVDD.n9663 4.5005
R1364 DVDD.n9683 DVDD.n9663 4.5005
R1365 DVDD.n9692 DVDD.n9663 4.5005
R1366 DVDD.n9682 DVDD.n9663 4.5005
R1367 DVDD.n9694 DVDD.n9663 4.5005
R1368 DVDD.n9681 DVDD.n9663 4.5005
R1369 DVDD.n9695 DVDD.n9663 4.5005
R1370 DVDD.n9680 DVDD.n9663 4.5005
R1371 DVDD.n10066 DVDD.n9663 4.5005
R1372 DVDD.n16113 DVDD.n3007 4.5005
R1373 DVDD.n3033 DVDD.n3007 4.5005
R1374 DVDD.n3031 DVDD.n3007 4.5005
R1375 DVDD.n3036 DVDD.n3007 4.5005
R1376 DVDD.n3029 DVDD.n3007 4.5005
R1377 DVDD.n3037 DVDD.n3007 4.5005
R1378 DVDD.n3028 DVDD.n3007 4.5005
R1379 DVDD.n3038 DVDD.n3007 4.5005
R1380 DVDD.n3027 DVDD.n3007 4.5005
R1381 DVDD.n16142 DVDD.n3007 4.5005
R1382 DVDD.n16144 DVDD.n3007 4.5005
R1383 DVDD.n3033 DVDD.n3009 4.5005
R1384 DVDD.n3031 DVDD.n3009 4.5005
R1385 DVDD.n3035 DVDD.n3009 4.5005
R1386 DVDD.n3030 DVDD.n3009 4.5005
R1387 DVDD.n3036 DVDD.n3009 4.5005
R1388 DVDD.n3029 DVDD.n3009 4.5005
R1389 DVDD.n3037 DVDD.n3009 4.5005
R1390 DVDD.n3028 DVDD.n3009 4.5005
R1391 DVDD.n3038 DVDD.n3009 4.5005
R1392 DVDD.n3027 DVDD.n3009 4.5005
R1393 DVDD.n3040 DVDD.n3009 4.5005
R1394 DVDD.n3026 DVDD.n3009 4.5005
R1395 DVDD.n16142 DVDD.n3009 4.5005
R1396 DVDD.n16144 DVDD.n3009 4.5005
R1397 DVDD.n3033 DVDD.n3006 4.5005
R1398 DVDD.n3031 DVDD.n3006 4.5005
R1399 DVDD.n3035 DVDD.n3006 4.5005
R1400 DVDD.n3030 DVDD.n3006 4.5005
R1401 DVDD.n3036 DVDD.n3006 4.5005
R1402 DVDD.n3029 DVDD.n3006 4.5005
R1403 DVDD.n3037 DVDD.n3006 4.5005
R1404 DVDD.n3028 DVDD.n3006 4.5005
R1405 DVDD.n3038 DVDD.n3006 4.5005
R1406 DVDD.n3027 DVDD.n3006 4.5005
R1407 DVDD.n3040 DVDD.n3006 4.5005
R1408 DVDD.n3026 DVDD.n3006 4.5005
R1409 DVDD.n16142 DVDD.n3006 4.5005
R1410 DVDD.n3006 DVDD.n2995 4.5005
R1411 DVDD.n16144 DVDD.n3006 4.5005
R1412 DVDD.n3033 DVDD.n3011 4.5005
R1413 DVDD.n3031 DVDD.n3011 4.5005
R1414 DVDD.n3035 DVDD.n3011 4.5005
R1415 DVDD.n3030 DVDD.n3011 4.5005
R1416 DVDD.n3036 DVDD.n3011 4.5005
R1417 DVDD.n3029 DVDD.n3011 4.5005
R1418 DVDD.n3037 DVDD.n3011 4.5005
R1419 DVDD.n3028 DVDD.n3011 4.5005
R1420 DVDD.n3038 DVDD.n3011 4.5005
R1421 DVDD.n3027 DVDD.n3011 4.5005
R1422 DVDD.n3040 DVDD.n3011 4.5005
R1423 DVDD.n3026 DVDD.n3011 4.5005
R1424 DVDD.n16142 DVDD.n3011 4.5005
R1425 DVDD.n16144 DVDD.n3011 4.5005
R1426 DVDD.n3033 DVDD.n3005 4.5005
R1427 DVDD.n3031 DVDD.n3005 4.5005
R1428 DVDD.n3035 DVDD.n3005 4.5005
R1429 DVDD.n3030 DVDD.n3005 4.5005
R1430 DVDD.n3036 DVDD.n3005 4.5005
R1431 DVDD.n3029 DVDD.n3005 4.5005
R1432 DVDD.n3037 DVDD.n3005 4.5005
R1433 DVDD.n3028 DVDD.n3005 4.5005
R1434 DVDD.n3038 DVDD.n3005 4.5005
R1435 DVDD.n3027 DVDD.n3005 4.5005
R1436 DVDD.n3040 DVDD.n3005 4.5005
R1437 DVDD.n3026 DVDD.n3005 4.5005
R1438 DVDD.n16142 DVDD.n3005 4.5005
R1439 DVDD.n16144 DVDD.n3005 4.5005
R1440 DVDD.n3033 DVDD.n3012 4.5005
R1441 DVDD.n3031 DVDD.n3012 4.5005
R1442 DVDD.n3035 DVDD.n3012 4.5005
R1443 DVDD.n3030 DVDD.n3012 4.5005
R1444 DVDD.n3036 DVDD.n3012 4.5005
R1445 DVDD.n3029 DVDD.n3012 4.5005
R1446 DVDD.n3037 DVDD.n3012 4.5005
R1447 DVDD.n3028 DVDD.n3012 4.5005
R1448 DVDD.n3038 DVDD.n3012 4.5005
R1449 DVDD.n3027 DVDD.n3012 4.5005
R1450 DVDD.n3040 DVDD.n3012 4.5005
R1451 DVDD.n3026 DVDD.n3012 4.5005
R1452 DVDD.n16142 DVDD.n3012 4.5005
R1453 DVDD.n3012 DVDD.n2995 4.5005
R1454 DVDD.n16144 DVDD.n3012 4.5005
R1455 DVDD.n3033 DVDD.n3004 4.5005
R1456 DVDD.n3031 DVDD.n3004 4.5005
R1457 DVDD.n3035 DVDD.n3004 4.5005
R1458 DVDD.n3030 DVDD.n3004 4.5005
R1459 DVDD.n3036 DVDD.n3004 4.5005
R1460 DVDD.n3029 DVDD.n3004 4.5005
R1461 DVDD.n3037 DVDD.n3004 4.5005
R1462 DVDD.n3028 DVDD.n3004 4.5005
R1463 DVDD.n3038 DVDD.n3004 4.5005
R1464 DVDD.n3027 DVDD.n3004 4.5005
R1465 DVDD.n3040 DVDD.n3004 4.5005
R1466 DVDD.n3026 DVDD.n3004 4.5005
R1467 DVDD.n16142 DVDD.n3004 4.5005
R1468 DVDD.n16144 DVDD.n3004 4.5005
R1469 DVDD.n3033 DVDD.n3014 4.5005
R1470 DVDD.n3031 DVDD.n3014 4.5005
R1471 DVDD.n3035 DVDD.n3014 4.5005
R1472 DVDD.n3030 DVDD.n3014 4.5005
R1473 DVDD.n3036 DVDD.n3014 4.5005
R1474 DVDD.n3029 DVDD.n3014 4.5005
R1475 DVDD.n3037 DVDD.n3014 4.5005
R1476 DVDD.n3028 DVDD.n3014 4.5005
R1477 DVDD.n3038 DVDD.n3014 4.5005
R1478 DVDD.n3027 DVDD.n3014 4.5005
R1479 DVDD.n3040 DVDD.n3014 4.5005
R1480 DVDD.n3026 DVDD.n3014 4.5005
R1481 DVDD.n16142 DVDD.n3014 4.5005
R1482 DVDD.n16144 DVDD.n3014 4.5005
R1483 DVDD.n3033 DVDD.n3003 4.5005
R1484 DVDD.n3031 DVDD.n3003 4.5005
R1485 DVDD.n3035 DVDD.n3003 4.5005
R1486 DVDD.n3030 DVDD.n3003 4.5005
R1487 DVDD.n3036 DVDD.n3003 4.5005
R1488 DVDD.n3029 DVDD.n3003 4.5005
R1489 DVDD.n3037 DVDD.n3003 4.5005
R1490 DVDD.n3028 DVDD.n3003 4.5005
R1491 DVDD.n3038 DVDD.n3003 4.5005
R1492 DVDD.n3027 DVDD.n3003 4.5005
R1493 DVDD.n3040 DVDD.n3003 4.5005
R1494 DVDD.n3026 DVDD.n3003 4.5005
R1495 DVDD.n16142 DVDD.n3003 4.5005
R1496 DVDD.n3003 DVDD.n2995 4.5005
R1497 DVDD.n16144 DVDD.n3003 4.5005
R1498 DVDD.n3033 DVDD.n3016 4.5005
R1499 DVDD.n3031 DVDD.n3016 4.5005
R1500 DVDD.n3035 DVDD.n3016 4.5005
R1501 DVDD.n3030 DVDD.n3016 4.5005
R1502 DVDD.n3036 DVDD.n3016 4.5005
R1503 DVDD.n3029 DVDD.n3016 4.5005
R1504 DVDD.n3037 DVDD.n3016 4.5005
R1505 DVDD.n3028 DVDD.n3016 4.5005
R1506 DVDD.n3038 DVDD.n3016 4.5005
R1507 DVDD.n3027 DVDD.n3016 4.5005
R1508 DVDD.n3040 DVDD.n3016 4.5005
R1509 DVDD.n3026 DVDD.n3016 4.5005
R1510 DVDD.n16142 DVDD.n3016 4.5005
R1511 DVDD.n16144 DVDD.n3016 4.5005
R1512 DVDD.n3033 DVDD.n3002 4.5005
R1513 DVDD.n3031 DVDD.n3002 4.5005
R1514 DVDD.n3035 DVDD.n3002 4.5005
R1515 DVDD.n3030 DVDD.n3002 4.5005
R1516 DVDD.n3036 DVDD.n3002 4.5005
R1517 DVDD.n3029 DVDD.n3002 4.5005
R1518 DVDD.n3037 DVDD.n3002 4.5005
R1519 DVDD.n3028 DVDD.n3002 4.5005
R1520 DVDD.n3038 DVDD.n3002 4.5005
R1521 DVDD.n3027 DVDD.n3002 4.5005
R1522 DVDD.n3040 DVDD.n3002 4.5005
R1523 DVDD.n3026 DVDD.n3002 4.5005
R1524 DVDD.n16142 DVDD.n3002 4.5005
R1525 DVDD.n16144 DVDD.n3002 4.5005
R1526 DVDD.n3033 DVDD.n3017 4.5005
R1527 DVDD.n3031 DVDD.n3017 4.5005
R1528 DVDD.n3035 DVDD.n3017 4.5005
R1529 DVDD.n3030 DVDD.n3017 4.5005
R1530 DVDD.n3036 DVDD.n3017 4.5005
R1531 DVDD.n3029 DVDD.n3017 4.5005
R1532 DVDD.n3037 DVDD.n3017 4.5005
R1533 DVDD.n3028 DVDD.n3017 4.5005
R1534 DVDD.n3038 DVDD.n3017 4.5005
R1535 DVDD.n3027 DVDD.n3017 4.5005
R1536 DVDD.n3040 DVDD.n3017 4.5005
R1537 DVDD.n3026 DVDD.n3017 4.5005
R1538 DVDD.n16142 DVDD.n3017 4.5005
R1539 DVDD.n3017 DVDD.n2995 4.5005
R1540 DVDD.n16144 DVDD.n3017 4.5005
R1541 DVDD.n3033 DVDD.n3001 4.5005
R1542 DVDD.n3031 DVDD.n3001 4.5005
R1543 DVDD.n3035 DVDD.n3001 4.5005
R1544 DVDD.n3030 DVDD.n3001 4.5005
R1545 DVDD.n3036 DVDD.n3001 4.5005
R1546 DVDD.n3029 DVDD.n3001 4.5005
R1547 DVDD.n3037 DVDD.n3001 4.5005
R1548 DVDD.n3028 DVDD.n3001 4.5005
R1549 DVDD.n3038 DVDD.n3001 4.5005
R1550 DVDD.n3027 DVDD.n3001 4.5005
R1551 DVDD.n3040 DVDD.n3001 4.5005
R1552 DVDD.n3026 DVDD.n3001 4.5005
R1553 DVDD.n16142 DVDD.n3001 4.5005
R1554 DVDD.n3001 DVDD.n2995 4.5005
R1555 DVDD.n16144 DVDD.n3001 4.5005
R1556 DVDD.n3033 DVDD.n3019 4.5005
R1557 DVDD.n3031 DVDD.n3019 4.5005
R1558 DVDD.n3035 DVDD.n3019 4.5005
R1559 DVDD.n3030 DVDD.n3019 4.5005
R1560 DVDD.n3036 DVDD.n3019 4.5005
R1561 DVDD.n3029 DVDD.n3019 4.5005
R1562 DVDD.n3037 DVDD.n3019 4.5005
R1563 DVDD.n3028 DVDD.n3019 4.5005
R1564 DVDD.n3038 DVDD.n3019 4.5005
R1565 DVDD.n3027 DVDD.n3019 4.5005
R1566 DVDD.n3040 DVDD.n3019 4.5005
R1567 DVDD.n3026 DVDD.n3019 4.5005
R1568 DVDD.n16142 DVDD.n3019 4.5005
R1569 DVDD.n16144 DVDD.n3019 4.5005
R1570 DVDD.n3033 DVDD.n3000 4.5005
R1571 DVDD.n3031 DVDD.n3000 4.5005
R1572 DVDD.n3035 DVDD.n3000 4.5005
R1573 DVDD.n3030 DVDD.n3000 4.5005
R1574 DVDD.n3036 DVDD.n3000 4.5005
R1575 DVDD.n3029 DVDD.n3000 4.5005
R1576 DVDD.n3037 DVDD.n3000 4.5005
R1577 DVDD.n3028 DVDD.n3000 4.5005
R1578 DVDD.n3038 DVDD.n3000 4.5005
R1579 DVDD.n3027 DVDD.n3000 4.5005
R1580 DVDD.n3040 DVDD.n3000 4.5005
R1581 DVDD.n3026 DVDD.n3000 4.5005
R1582 DVDD.n16142 DVDD.n3000 4.5005
R1583 DVDD.n16144 DVDD.n3000 4.5005
R1584 DVDD.n3033 DVDD.n3020 4.5005
R1585 DVDD.n3031 DVDD.n3020 4.5005
R1586 DVDD.n3035 DVDD.n3020 4.5005
R1587 DVDD.n3030 DVDD.n3020 4.5005
R1588 DVDD.n3036 DVDD.n3020 4.5005
R1589 DVDD.n3029 DVDD.n3020 4.5005
R1590 DVDD.n3037 DVDD.n3020 4.5005
R1591 DVDD.n3028 DVDD.n3020 4.5005
R1592 DVDD.n3038 DVDD.n3020 4.5005
R1593 DVDD.n3027 DVDD.n3020 4.5005
R1594 DVDD.n3040 DVDD.n3020 4.5005
R1595 DVDD.n3026 DVDD.n3020 4.5005
R1596 DVDD.n16142 DVDD.n3020 4.5005
R1597 DVDD.n3020 DVDD.n2995 4.5005
R1598 DVDD.n16144 DVDD.n3020 4.5005
R1599 DVDD.n3033 DVDD.n2999 4.5005
R1600 DVDD.n3031 DVDD.n2999 4.5005
R1601 DVDD.n3035 DVDD.n2999 4.5005
R1602 DVDD.n3030 DVDD.n2999 4.5005
R1603 DVDD.n3036 DVDD.n2999 4.5005
R1604 DVDD.n3029 DVDD.n2999 4.5005
R1605 DVDD.n3037 DVDD.n2999 4.5005
R1606 DVDD.n3028 DVDD.n2999 4.5005
R1607 DVDD.n3038 DVDD.n2999 4.5005
R1608 DVDD.n3027 DVDD.n2999 4.5005
R1609 DVDD.n3040 DVDD.n2999 4.5005
R1610 DVDD.n3026 DVDD.n2999 4.5005
R1611 DVDD.n16142 DVDD.n2999 4.5005
R1612 DVDD.n2999 DVDD.n2995 4.5005
R1613 DVDD.n16144 DVDD.n2999 4.5005
R1614 DVDD.n3033 DVDD.n3022 4.5005
R1615 DVDD.n3031 DVDD.n3022 4.5005
R1616 DVDD.n3035 DVDD.n3022 4.5005
R1617 DVDD.n3030 DVDD.n3022 4.5005
R1618 DVDD.n3036 DVDD.n3022 4.5005
R1619 DVDD.n3029 DVDD.n3022 4.5005
R1620 DVDD.n3037 DVDD.n3022 4.5005
R1621 DVDD.n3028 DVDD.n3022 4.5005
R1622 DVDD.n3038 DVDD.n3022 4.5005
R1623 DVDD.n3027 DVDD.n3022 4.5005
R1624 DVDD.n3040 DVDD.n3022 4.5005
R1625 DVDD.n3026 DVDD.n3022 4.5005
R1626 DVDD.n16142 DVDD.n3022 4.5005
R1627 DVDD.n16144 DVDD.n3022 4.5005
R1628 DVDD.n3033 DVDD.n2998 4.5005
R1629 DVDD.n3031 DVDD.n2998 4.5005
R1630 DVDD.n3035 DVDD.n2998 4.5005
R1631 DVDD.n3030 DVDD.n2998 4.5005
R1632 DVDD.n3036 DVDD.n2998 4.5005
R1633 DVDD.n3029 DVDD.n2998 4.5005
R1634 DVDD.n3037 DVDD.n2998 4.5005
R1635 DVDD.n3028 DVDD.n2998 4.5005
R1636 DVDD.n3038 DVDD.n2998 4.5005
R1637 DVDD.n3027 DVDD.n2998 4.5005
R1638 DVDD.n3040 DVDD.n2998 4.5005
R1639 DVDD.n3026 DVDD.n2998 4.5005
R1640 DVDD.n16142 DVDD.n2998 4.5005
R1641 DVDD.n16144 DVDD.n2998 4.5005
R1642 DVDD.n3033 DVDD.n3023 4.5005
R1643 DVDD.n3031 DVDD.n3023 4.5005
R1644 DVDD.n3035 DVDD.n3023 4.5005
R1645 DVDD.n3030 DVDD.n3023 4.5005
R1646 DVDD.n3036 DVDD.n3023 4.5005
R1647 DVDD.n3029 DVDD.n3023 4.5005
R1648 DVDD.n3037 DVDD.n3023 4.5005
R1649 DVDD.n3028 DVDD.n3023 4.5005
R1650 DVDD.n3038 DVDD.n3023 4.5005
R1651 DVDD.n3027 DVDD.n3023 4.5005
R1652 DVDD.n3040 DVDD.n3023 4.5005
R1653 DVDD.n3026 DVDD.n3023 4.5005
R1654 DVDD.n16142 DVDD.n3023 4.5005
R1655 DVDD.n3023 DVDD.n2995 4.5005
R1656 DVDD.n16144 DVDD.n3023 4.5005
R1657 DVDD.n16113 DVDD.n2997 4.5005
R1658 DVDD.n3033 DVDD.n2997 4.5005
R1659 DVDD.n3031 DVDD.n2997 4.5005
R1660 DVDD.n3035 DVDD.n2997 4.5005
R1661 DVDD.n3030 DVDD.n2997 4.5005
R1662 DVDD.n3036 DVDD.n2997 4.5005
R1663 DVDD.n3029 DVDD.n2997 4.5005
R1664 DVDD.n3037 DVDD.n2997 4.5005
R1665 DVDD.n3028 DVDD.n2997 4.5005
R1666 DVDD.n3038 DVDD.n2997 4.5005
R1667 DVDD.n3027 DVDD.n2997 4.5005
R1668 DVDD.n3040 DVDD.n2997 4.5005
R1669 DVDD.n3026 DVDD.n2997 4.5005
R1670 DVDD.n16142 DVDD.n2997 4.5005
R1671 DVDD.n2997 DVDD.n2995 4.5005
R1672 DVDD.n16144 DVDD.n2997 4.5005
R1673 DVDD.n2769 DVDD.n2752 4.5005
R1674 DVDD.n2769 DVDD.n2753 4.5005
R1675 DVDD.n2769 DVDD.n2751 4.5005
R1676 DVDD.n2769 DVDD.n2755 4.5005
R1677 DVDD.n2769 DVDD.n2749 4.5005
R1678 DVDD.n2769 DVDD.n2756 4.5005
R1679 DVDD.n2769 DVDD.n2748 4.5005
R1680 DVDD.n2769 DVDD.n2757 4.5005
R1681 DVDD.n2769 DVDD.n2710 4.5005
R1682 DVDD.n2769 DVDD.n2766 4.5005
R1683 DVDD.n2769 DVDD.n2746 4.5005
R1684 DVDD.n16255 DVDD.n2769 4.5005
R1685 DVDD.n2752 DVDD.n2723 4.5005
R1686 DVDD.n2753 DVDD.n2723 4.5005
R1687 DVDD.n2751 DVDD.n2723 4.5005
R1688 DVDD.n2754 DVDD.n2723 4.5005
R1689 DVDD.n2750 DVDD.n2723 4.5005
R1690 DVDD.n2755 DVDD.n2723 4.5005
R1691 DVDD.n2749 DVDD.n2723 4.5005
R1692 DVDD.n2756 DVDD.n2723 4.5005
R1693 DVDD.n2748 DVDD.n2723 4.5005
R1694 DVDD.n2757 DVDD.n2723 4.5005
R1695 DVDD.n2723 DVDD.n2710 4.5005
R1696 DVDD.n16257 DVDD.n2723 4.5005
R1697 DVDD.n2764 DVDD.n2723 4.5005
R1698 DVDD.n2766 DVDD.n2723 4.5005
R1699 DVDD.n16255 DVDD.n2723 4.5005
R1700 DVDD.n2752 DVDD.n2721 4.5005
R1701 DVDD.n2753 DVDD.n2721 4.5005
R1702 DVDD.n2751 DVDD.n2721 4.5005
R1703 DVDD.n2754 DVDD.n2721 4.5005
R1704 DVDD.n2750 DVDD.n2721 4.5005
R1705 DVDD.n2755 DVDD.n2721 4.5005
R1706 DVDD.n2749 DVDD.n2721 4.5005
R1707 DVDD.n2756 DVDD.n2721 4.5005
R1708 DVDD.n2748 DVDD.n2721 4.5005
R1709 DVDD.n2757 DVDD.n2721 4.5005
R1710 DVDD.n2721 DVDD.n2710 4.5005
R1711 DVDD.n16257 DVDD.n2721 4.5005
R1712 DVDD.n2766 DVDD.n2721 4.5005
R1713 DVDD.n16255 DVDD.n2721 4.5005
R1714 DVDD.n2752 DVDD.n2724 4.5005
R1715 DVDD.n2753 DVDD.n2724 4.5005
R1716 DVDD.n2751 DVDD.n2724 4.5005
R1717 DVDD.n2754 DVDD.n2724 4.5005
R1718 DVDD.n2750 DVDD.n2724 4.5005
R1719 DVDD.n2755 DVDD.n2724 4.5005
R1720 DVDD.n2749 DVDD.n2724 4.5005
R1721 DVDD.n2756 DVDD.n2724 4.5005
R1722 DVDD.n2748 DVDD.n2724 4.5005
R1723 DVDD.n2757 DVDD.n2724 4.5005
R1724 DVDD.n2724 DVDD.n2710 4.5005
R1725 DVDD.n16257 DVDD.n2724 4.5005
R1726 DVDD.n2766 DVDD.n2724 4.5005
R1727 DVDD.n16255 DVDD.n2724 4.5005
R1728 DVDD.n2752 DVDD.n2720 4.5005
R1729 DVDD.n2753 DVDD.n2720 4.5005
R1730 DVDD.n2751 DVDD.n2720 4.5005
R1731 DVDD.n2754 DVDD.n2720 4.5005
R1732 DVDD.n2750 DVDD.n2720 4.5005
R1733 DVDD.n2755 DVDD.n2720 4.5005
R1734 DVDD.n2749 DVDD.n2720 4.5005
R1735 DVDD.n2756 DVDD.n2720 4.5005
R1736 DVDD.n2748 DVDD.n2720 4.5005
R1737 DVDD.n2757 DVDD.n2720 4.5005
R1738 DVDD.n2720 DVDD.n2710 4.5005
R1739 DVDD.n16257 DVDD.n2720 4.5005
R1740 DVDD.n2764 DVDD.n2720 4.5005
R1741 DVDD.n2766 DVDD.n2720 4.5005
R1742 DVDD.n16255 DVDD.n2720 4.5005
R1743 DVDD.n2752 DVDD.n2725 4.5005
R1744 DVDD.n2753 DVDD.n2725 4.5005
R1745 DVDD.n2751 DVDD.n2725 4.5005
R1746 DVDD.n2754 DVDD.n2725 4.5005
R1747 DVDD.n2750 DVDD.n2725 4.5005
R1748 DVDD.n2755 DVDD.n2725 4.5005
R1749 DVDD.n2749 DVDD.n2725 4.5005
R1750 DVDD.n2756 DVDD.n2725 4.5005
R1751 DVDD.n2748 DVDD.n2725 4.5005
R1752 DVDD.n2757 DVDD.n2725 4.5005
R1753 DVDD.n2725 DVDD.n2710 4.5005
R1754 DVDD.n16257 DVDD.n2725 4.5005
R1755 DVDD.n2764 DVDD.n2725 4.5005
R1756 DVDD.n2766 DVDD.n2725 4.5005
R1757 DVDD.n16255 DVDD.n2725 4.5005
R1758 DVDD.n2752 DVDD.n2719 4.5005
R1759 DVDD.n2753 DVDD.n2719 4.5005
R1760 DVDD.n2751 DVDD.n2719 4.5005
R1761 DVDD.n2754 DVDD.n2719 4.5005
R1762 DVDD.n2750 DVDD.n2719 4.5005
R1763 DVDD.n2755 DVDD.n2719 4.5005
R1764 DVDD.n2749 DVDD.n2719 4.5005
R1765 DVDD.n2756 DVDD.n2719 4.5005
R1766 DVDD.n2748 DVDD.n2719 4.5005
R1767 DVDD.n2757 DVDD.n2719 4.5005
R1768 DVDD.n2719 DVDD.n2710 4.5005
R1769 DVDD.n16257 DVDD.n2719 4.5005
R1770 DVDD.n2766 DVDD.n2719 4.5005
R1771 DVDD.n16255 DVDD.n2719 4.5005
R1772 DVDD.n2752 DVDD.n2726 4.5005
R1773 DVDD.n2753 DVDD.n2726 4.5005
R1774 DVDD.n2751 DVDD.n2726 4.5005
R1775 DVDD.n2754 DVDD.n2726 4.5005
R1776 DVDD.n2750 DVDD.n2726 4.5005
R1777 DVDD.n2755 DVDD.n2726 4.5005
R1778 DVDD.n2749 DVDD.n2726 4.5005
R1779 DVDD.n2756 DVDD.n2726 4.5005
R1780 DVDD.n2748 DVDD.n2726 4.5005
R1781 DVDD.n2757 DVDD.n2726 4.5005
R1782 DVDD.n2726 DVDD.n2710 4.5005
R1783 DVDD.n16257 DVDD.n2726 4.5005
R1784 DVDD.n2766 DVDD.n2726 4.5005
R1785 DVDD.n16255 DVDD.n2726 4.5005
R1786 DVDD.n2752 DVDD.n2718 4.5005
R1787 DVDD.n2753 DVDD.n2718 4.5005
R1788 DVDD.n2751 DVDD.n2718 4.5005
R1789 DVDD.n2754 DVDD.n2718 4.5005
R1790 DVDD.n2750 DVDD.n2718 4.5005
R1791 DVDD.n2755 DVDD.n2718 4.5005
R1792 DVDD.n2749 DVDD.n2718 4.5005
R1793 DVDD.n2756 DVDD.n2718 4.5005
R1794 DVDD.n2748 DVDD.n2718 4.5005
R1795 DVDD.n2757 DVDD.n2718 4.5005
R1796 DVDD.n2718 DVDD.n2710 4.5005
R1797 DVDD.n16257 DVDD.n2718 4.5005
R1798 DVDD.n2764 DVDD.n2718 4.5005
R1799 DVDD.n2766 DVDD.n2718 4.5005
R1800 DVDD.n16255 DVDD.n2718 4.5005
R1801 DVDD.n2752 DVDD.n2727 4.5005
R1802 DVDD.n2753 DVDD.n2727 4.5005
R1803 DVDD.n2751 DVDD.n2727 4.5005
R1804 DVDD.n2754 DVDD.n2727 4.5005
R1805 DVDD.n2750 DVDD.n2727 4.5005
R1806 DVDD.n2755 DVDD.n2727 4.5005
R1807 DVDD.n2749 DVDD.n2727 4.5005
R1808 DVDD.n2756 DVDD.n2727 4.5005
R1809 DVDD.n2748 DVDD.n2727 4.5005
R1810 DVDD.n2757 DVDD.n2727 4.5005
R1811 DVDD.n2727 DVDD.n2710 4.5005
R1812 DVDD.n16257 DVDD.n2727 4.5005
R1813 DVDD.n2764 DVDD.n2727 4.5005
R1814 DVDD.n2766 DVDD.n2727 4.5005
R1815 DVDD.n16255 DVDD.n2727 4.5005
R1816 DVDD.n2752 DVDD.n2717 4.5005
R1817 DVDD.n2753 DVDD.n2717 4.5005
R1818 DVDD.n2751 DVDD.n2717 4.5005
R1819 DVDD.n2754 DVDD.n2717 4.5005
R1820 DVDD.n2750 DVDD.n2717 4.5005
R1821 DVDD.n2755 DVDD.n2717 4.5005
R1822 DVDD.n2749 DVDD.n2717 4.5005
R1823 DVDD.n2756 DVDD.n2717 4.5005
R1824 DVDD.n2748 DVDD.n2717 4.5005
R1825 DVDD.n2757 DVDD.n2717 4.5005
R1826 DVDD.n2717 DVDD.n2710 4.5005
R1827 DVDD.n16257 DVDD.n2717 4.5005
R1828 DVDD.n2766 DVDD.n2717 4.5005
R1829 DVDD.n16255 DVDD.n2717 4.5005
R1830 DVDD.n2752 DVDD.n2728 4.5005
R1831 DVDD.n2753 DVDD.n2728 4.5005
R1832 DVDD.n2751 DVDD.n2728 4.5005
R1833 DVDD.n2754 DVDD.n2728 4.5005
R1834 DVDD.n2750 DVDD.n2728 4.5005
R1835 DVDD.n2755 DVDD.n2728 4.5005
R1836 DVDD.n2749 DVDD.n2728 4.5005
R1837 DVDD.n2756 DVDD.n2728 4.5005
R1838 DVDD.n2748 DVDD.n2728 4.5005
R1839 DVDD.n2757 DVDD.n2728 4.5005
R1840 DVDD.n2728 DVDD.n2710 4.5005
R1841 DVDD.n16257 DVDD.n2728 4.5005
R1842 DVDD.n2766 DVDD.n2728 4.5005
R1843 DVDD.n16255 DVDD.n2728 4.5005
R1844 DVDD.n2752 DVDD.n2716 4.5005
R1845 DVDD.n2753 DVDD.n2716 4.5005
R1846 DVDD.n2751 DVDD.n2716 4.5005
R1847 DVDD.n2754 DVDD.n2716 4.5005
R1848 DVDD.n2750 DVDD.n2716 4.5005
R1849 DVDD.n2755 DVDD.n2716 4.5005
R1850 DVDD.n2749 DVDD.n2716 4.5005
R1851 DVDD.n2756 DVDD.n2716 4.5005
R1852 DVDD.n2748 DVDD.n2716 4.5005
R1853 DVDD.n2757 DVDD.n2716 4.5005
R1854 DVDD.n2716 DVDD.n2710 4.5005
R1855 DVDD.n16257 DVDD.n2716 4.5005
R1856 DVDD.n2764 DVDD.n2716 4.5005
R1857 DVDD.n2766 DVDD.n2716 4.5005
R1858 DVDD.n16255 DVDD.n2716 4.5005
R1859 DVDD.n2752 DVDD.n2729 4.5005
R1860 DVDD.n2753 DVDD.n2729 4.5005
R1861 DVDD.n2751 DVDD.n2729 4.5005
R1862 DVDD.n2754 DVDD.n2729 4.5005
R1863 DVDD.n2750 DVDD.n2729 4.5005
R1864 DVDD.n2755 DVDD.n2729 4.5005
R1865 DVDD.n2749 DVDD.n2729 4.5005
R1866 DVDD.n2756 DVDD.n2729 4.5005
R1867 DVDD.n2748 DVDD.n2729 4.5005
R1868 DVDD.n2757 DVDD.n2729 4.5005
R1869 DVDD.n2729 DVDD.n2710 4.5005
R1870 DVDD.n16257 DVDD.n2729 4.5005
R1871 DVDD.n2764 DVDD.n2729 4.5005
R1872 DVDD.n2766 DVDD.n2729 4.5005
R1873 DVDD.n16255 DVDD.n2729 4.5005
R1874 DVDD.n2752 DVDD.n2715 4.5005
R1875 DVDD.n2753 DVDD.n2715 4.5005
R1876 DVDD.n2751 DVDD.n2715 4.5005
R1877 DVDD.n2754 DVDD.n2715 4.5005
R1878 DVDD.n2750 DVDD.n2715 4.5005
R1879 DVDD.n2755 DVDD.n2715 4.5005
R1880 DVDD.n2749 DVDD.n2715 4.5005
R1881 DVDD.n2756 DVDD.n2715 4.5005
R1882 DVDD.n2748 DVDD.n2715 4.5005
R1883 DVDD.n2757 DVDD.n2715 4.5005
R1884 DVDD.n2715 DVDD.n2710 4.5005
R1885 DVDD.n16257 DVDD.n2715 4.5005
R1886 DVDD.n2766 DVDD.n2715 4.5005
R1887 DVDD.n16255 DVDD.n2715 4.5005
R1888 DVDD.n2752 DVDD.n2730 4.5005
R1889 DVDD.n2753 DVDD.n2730 4.5005
R1890 DVDD.n2751 DVDD.n2730 4.5005
R1891 DVDD.n2754 DVDD.n2730 4.5005
R1892 DVDD.n2750 DVDD.n2730 4.5005
R1893 DVDD.n2755 DVDD.n2730 4.5005
R1894 DVDD.n2749 DVDD.n2730 4.5005
R1895 DVDD.n2756 DVDD.n2730 4.5005
R1896 DVDD.n2748 DVDD.n2730 4.5005
R1897 DVDD.n2757 DVDD.n2730 4.5005
R1898 DVDD.n2730 DVDD.n2710 4.5005
R1899 DVDD.n16257 DVDD.n2730 4.5005
R1900 DVDD.n2766 DVDD.n2730 4.5005
R1901 DVDD.n16255 DVDD.n2730 4.5005
R1902 DVDD.n2752 DVDD.n2714 4.5005
R1903 DVDD.n2753 DVDD.n2714 4.5005
R1904 DVDD.n2751 DVDD.n2714 4.5005
R1905 DVDD.n2754 DVDD.n2714 4.5005
R1906 DVDD.n2750 DVDD.n2714 4.5005
R1907 DVDD.n2755 DVDD.n2714 4.5005
R1908 DVDD.n2749 DVDD.n2714 4.5005
R1909 DVDD.n2756 DVDD.n2714 4.5005
R1910 DVDD.n2748 DVDD.n2714 4.5005
R1911 DVDD.n2757 DVDD.n2714 4.5005
R1912 DVDD.n2714 DVDD.n2710 4.5005
R1913 DVDD.n16257 DVDD.n2714 4.5005
R1914 DVDD.n2766 DVDD.n2714 4.5005
R1915 DVDD.n16255 DVDD.n2714 4.5005
R1916 DVDD.n2752 DVDD.n2731 4.5005
R1917 DVDD.n2753 DVDD.n2731 4.5005
R1918 DVDD.n2751 DVDD.n2731 4.5005
R1919 DVDD.n2754 DVDD.n2731 4.5005
R1920 DVDD.n2750 DVDD.n2731 4.5005
R1921 DVDD.n2755 DVDD.n2731 4.5005
R1922 DVDD.n2749 DVDD.n2731 4.5005
R1923 DVDD.n2756 DVDD.n2731 4.5005
R1924 DVDD.n2748 DVDD.n2731 4.5005
R1925 DVDD.n2757 DVDD.n2731 4.5005
R1926 DVDD.n2731 DVDD.n2710 4.5005
R1927 DVDD.n16257 DVDD.n2731 4.5005
R1928 DVDD.n2766 DVDD.n2731 4.5005
R1929 DVDD.n16255 DVDD.n2731 4.5005
R1930 DVDD.n2752 DVDD.n2713 4.5005
R1931 DVDD.n2753 DVDD.n2713 4.5005
R1932 DVDD.n2751 DVDD.n2713 4.5005
R1933 DVDD.n2754 DVDD.n2713 4.5005
R1934 DVDD.n2750 DVDD.n2713 4.5005
R1935 DVDD.n2755 DVDD.n2713 4.5005
R1936 DVDD.n2749 DVDD.n2713 4.5005
R1937 DVDD.n2756 DVDD.n2713 4.5005
R1938 DVDD.n2748 DVDD.n2713 4.5005
R1939 DVDD.n2757 DVDD.n2713 4.5005
R1940 DVDD.n2713 DVDD.n2710 4.5005
R1941 DVDD.n16257 DVDD.n2713 4.5005
R1942 DVDD.n2766 DVDD.n2713 4.5005
R1943 DVDD.n16255 DVDD.n2713 4.5005
R1944 DVDD.n2752 DVDD.n2732 4.5005
R1945 DVDD.n2753 DVDD.n2732 4.5005
R1946 DVDD.n2751 DVDD.n2732 4.5005
R1947 DVDD.n2754 DVDD.n2732 4.5005
R1948 DVDD.n2750 DVDD.n2732 4.5005
R1949 DVDD.n2755 DVDD.n2732 4.5005
R1950 DVDD.n2749 DVDD.n2732 4.5005
R1951 DVDD.n2756 DVDD.n2732 4.5005
R1952 DVDD.n2748 DVDD.n2732 4.5005
R1953 DVDD.n2757 DVDD.n2732 4.5005
R1954 DVDD.n2732 DVDD.n2710 4.5005
R1955 DVDD.n16257 DVDD.n2732 4.5005
R1956 DVDD.n2766 DVDD.n2732 4.5005
R1957 DVDD.n16255 DVDD.n2732 4.5005
R1958 DVDD.n2752 DVDD.n2712 4.5005
R1959 DVDD.n2753 DVDD.n2712 4.5005
R1960 DVDD.n2751 DVDD.n2712 4.5005
R1961 DVDD.n2754 DVDD.n2712 4.5005
R1962 DVDD.n2750 DVDD.n2712 4.5005
R1963 DVDD.n2755 DVDD.n2712 4.5005
R1964 DVDD.n2749 DVDD.n2712 4.5005
R1965 DVDD.n2756 DVDD.n2712 4.5005
R1966 DVDD.n2748 DVDD.n2712 4.5005
R1967 DVDD.n2757 DVDD.n2712 4.5005
R1968 DVDD.n2712 DVDD.n2710 4.5005
R1969 DVDD.n16257 DVDD.n2712 4.5005
R1970 DVDD.n2764 DVDD.n2712 4.5005
R1971 DVDD.n2766 DVDD.n2712 4.5005
R1972 DVDD.n16255 DVDD.n2712 4.5005
R1973 DVDD.n2752 DVDD.n2733 4.5005
R1974 DVDD.n2753 DVDD.n2733 4.5005
R1975 DVDD.n2751 DVDD.n2733 4.5005
R1976 DVDD.n2754 DVDD.n2733 4.5005
R1977 DVDD.n2750 DVDD.n2733 4.5005
R1978 DVDD.n2755 DVDD.n2733 4.5005
R1979 DVDD.n2749 DVDD.n2733 4.5005
R1980 DVDD.n2756 DVDD.n2733 4.5005
R1981 DVDD.n2748 DVDD.n2733 4.5005
R1982 DVDD.n2757 DVDD.n2733 4.5005
R1983 DVDD.n2733 DVDD.n2710 4.5005
R1984 DVDD.n16257 DVDD.n2733 4.5005
R1985 DVDD.n2764 DVDD.n2733 4.5005
R1986 DVDD.n2766 DVDD.n2733 4.5005
R1987 DVDD.n16255 DVDD.n2733 4.5005
R1988 DVDD.n2752 DVDD.n2711 4.5005
R1989 DVDD.n2753 DVDD.n2711 4.5005
R1990 DVDD.n2751 DVDD.n2711 4.5005
R1991 DVDD.n2754 DVDD.n2711 4.5005
R1992 DVDD.n2750 DVDD.n2711 4.5005
R1993 DVDD.n2755 DVDD.n2711 4.5005
R1994 DVDD.n2749 DVDD.n2711 4.5005
R1995 DVDD.n2756 DVDD.n2711 4.5005
R1996 DVDD.n2748 DVDD.n2711 4.5005
R1997 DVDD.n2757 DVDD.n2711 4.5005
R1998 DVDD.n2711 DVDD.n2710 4.5005
R1999 DVDD.n16257 DVDD.n2711 4.5005
R2000 DVDD.n2766 DVDD.n2711 4.5005
R2001 DVDD.n16255 DVDD.n2711 4.5005
R2002 DVDD.n16256 DVDD.n2752 4.5005
R2003 DVDD.n16256 DVDD.n2753 4.5005
R2004 DVDD.n16256 DVDD.n2751 4.5005
R2005 DVDD.n16256 DVDD.n2754 4.5005
R2006 DVDD.n16256 DVDD.n2750 4.5005
R2007 DVDD.n16256 DVDD.n2755 4.5005
R2008 DVDD.n16256 DVDD.n2749 4.5005
R2009 DVDD.n16256 DVDD.n2756 4.5005
R2010 DVDD.n16256 DVDD.n2748 4.5005
R2011 DVDD.n16256 DVDD.n2757 4.5005
R2012 DVDD.n16256 DVDD.n2710 4.5005
R2013 DVDD.n16257 DVDD.n16256 4.5005
R2014 DVDD.n16256 DVDD.n2766 4.5005
R2015 DVDD.n16256 DVDD.n2746 4.5005
R2016 DVDD.n16256 DVDD.n16255 4.5005
R2017 DVDD.n2691 DVDD.n2656 4.5005
R2018 DVDD.n2693 DVDD.n2656 4.5005
R2019 DVDD.n2690 DVDD.n2656 4.5005
R2020 DVDD.n2696 DVDD.n2656 4.5005
R2021 DVDD.n2688 DVDD.n2656 4.5005
R2022 DVDD.n2697 DVDD.n2656 4.5005
R2023 DVDD.n2687 DVDD.n2656 4.5005
R2024 DVDD.n2698 DVDD.n2656 4.5005
R2025 DVDD.n2686 DVDD.n2656 4.5005
R2026 DVDD.n16268 DVDD.n2656 4.5005
R2027 DVDD.n16270 DVDD.n2656 4.5005
R2028 DVDD.n2691 DVDD.n2658 4.5005
R2029 DVDD.n2693 DVDD.n2658 4.5005
R2030 DVDD.n2690 DVDD.n2658 4.5005
R2031 DVDD.n2695 DVDD.n2658 4.5005
R2032 DVDD.n2689 DVDD.n2658 4.5005
R2033 DVDD.n2696 DVDD.n2658 4.5005
R2034 DVDD.n2688 DVDD.n2658 4.5005
R2035 DVDD.n2697 DVDD.n2658 4.5005
R2036 DVDD.n2687 DVDD.n2658 4.5005
R2037 DVDD.n2698 DVDD.n2658 4.5005
R2038 DVDD.n2686 DVDD.n2658 4.5005
R2039 DVDD.n2700 DVDD.n2658 4.5005
R2040 DVDD.n16268 DVDD.n2658 4.5005
R2041 DVDD.n16270 DVDD.n2658 4.5005
R2042 DVDD.n2691 DVDD.n2655 4.5005
R2043 DVDD.n2693 DVDD.n2655 4.5005
R2044 DVDD.n2690 DVDD.n2655 4.5005
R2045 DVDD.n2695 DVDD.n2655 4.5005
R2046 DVDD.n2689 DVDD.n2655 4.5005
R2047 DVDD.n2696 DVDD.n2655 4.5005
R2048 DVDD.n2688 DVDD.n2655 4.5005
R2049 DVDD.n2697 DVDD.n2655 4.5005
R2050 DVDD.n2687 DVDD.n2655 4.5005
R2051 DVDD.n2698 DVDD.n2655 4.5005
R2052 DVDD.n2686 DVDD.n2655 4.5005
R2053 DVDD.n2700 DVDD.n2655 4.5005
R2054 DVDD.n16268 DVDD.n2655 4.5005
R2055 DVDD.n2655 DVDD.n2644 4.5005
R2056 DVDD.n16270 DVDD.n2655 4.5005
R2057 DVDD.n2691 DVDD.n2660 4.5005
R2058 DVDD.n2693 DVDD.n2660 4.5005
R2059 DVDD.n2690 DVDD.n2660 4.5005
R2060 DVDD.n2695 DVDD.n2660 4.5005
R2061 DVDD.n2689 DVDD.n2660 4.5005
R2062 DVDD.n2696 DVDD.n2660 4.5005
R2063 DVDD.n2688 DVDD.n2660 4.5005
R2064 DVDD.n2697 DVDD.n2660 4.5005
R2065 DVDD.n2687 DVDD.n2660 4.5005
R2066 DVDD.n2698 DVDD.n2660 4.5005
R2067 DVDD.n2686 DVDD.n2660 4.5005
R2068 DVDD.n2700 DVDD.n2660 4.5005
R2069 DVDD.n2685 DVDD.n2660 4.5005
R2070 DVDD.n16268 DVDD.n2660 4.5005
R2071 DVDD.n16270 DVDD.n2660 4.5005
R2072 DVDD.n2691 DVDD.n2654 4.5005
R2073 DVDD.n2693 DVDD.n2654 4.5005
R2074 DVDD.n2690 DVDD.n2654 4.5005
R2075 DVDD.n2695 DVDD.n2654 4.5005
R2076 DVDD.n2689 DVDD.n2654 4.5005
R2077 DVDD.n2696 DVDD.n2654 4.5005
R2078 DVDD.n2688 DVDD.n2654 4.5005
R2079 DVDD.n2697 DVDD.n2654 4.5005
R2080 DVDD.n2687 DVDD.n2654 4.5005
R2081 DVDD.n2698 DVDD.n2654 4.5005
R2082 DVDD.n2686 DVDD.n2654 4.5005
R2083 DVDD.n2700 DVDD.n2654 4.5005
R2084 DVDD.n16268 DVDD.n2654 4.5005
R2085 DVDD.n16270 DVDD.n2654 4.5005
R2086 DVDD.n2691 DVDD.n2662 4.5005
R2087 DVDD.n2693 DVDD.n2662 4.5005
R2088 DVDD.n2690 DVDD.n2662 4.5005
R2089 DVDD.n2695 DVDD.n2662 4.5005
R2090 DVDD.n2689 DVDD.n2662 4.5005
R2091 DVDD.n2696 DVDD.n2662 4.5005
R2092 DVDD.n2688 DVDD.n2662 4.5005
R2093 DVDD.n2697 DVDD.n2662 4.5005
R2094 DVDD.n2687 DVDD.n2662 4.5005
R2095 DVDD.n2698 DVDD.n2662 4.5005
R2096 DVDD.n2686 DVDD.n2662 4.5005
R2097 DVDD.n2700 DVDD.n2662 4.5005
R2098 DVDD.n16268 DVDD.n2662 4.5005
R2099 DVDD.n16270 DVDD.n2662 4.5005
R2100 DVDD.n2691 DVDD.n2653 4.5005
R2101 DVDD.n2693 DVDD.n2653 4.5005
R2102 DVDD.n2690 DVDD.n2653 4.5005
R2103 DVDD.n2695 DVDD.n2653 4.5005
R2104 DVDD.n2689 DVDD.n2653 4.5005
R2105 DVDD.n2696 DVDD.n2653 4.5005
R2106 DVDD.n2688 DVDD.n2653 4.5005
R2107 DVDD.n2697 DVDD.n2653 4.5005
R2108 DVDD.n2687 DVDD.n2653 4.5005
R2109 DVDD.n2698 DVDD.n2653 4.5005
R2110 DVDD.n2686 DVDD.n2653 4.5005
R2111 DVDD.n2700 DVDD.n2653 4.5005
R2112 DVDD.n2685 DVDD.n2653 4.5005
R2113 DVDD.n16268 DVDD.n2653 4.5005
R2114 DVDD.n16270 DVDD.n2653 4.5005
R2115 DVDD.n2691 DVDD.n2664 4.5005
R2116 DVDD.n2693 DVDD.n2664 4.5005
R2117 DVDD.n2690 DVDD.n2664 4.5005
R2118 DVDD.n2695 DVDD.n2664 4.5005
R2119 DVDD.n2689 DVDD.n2664 4.5005
R2120 DVDD.n2696 DVDD.n2664 4.5005
R2121 DVDD.n2688 DVDD.n2664 4.5005
R2122 DVDD.n2697 DVDD.n2664 4.5005
R2123 DVDD.n2687 DVDD.n2664 4.5005
R2124 DVDD.n2698 DVDD.n2664 4.5005
R2125 DVDD.n2686 DVDD.n2664 4.5005
R2126 DVDD.n2700 DVDD.n2664 4.5005
R2127 DVDD.n2685 DVDD.n2664 4.5005
R2128 DVDD.n16268 DVDD.n2664 4.5005
R2129 DVDD.n16270 DVDD.n2664 4.5005
R2130 DVDD.n2691 DVDD.n2652 4.5005
R2131 DVDD.n2693 DVDD.n2652 4.5005
R2132 DVDD.n2690 DVDD.n2652 4.5005
R2133 DVDD.n2695 DVDD.n2652 4.5005
R2134 DVDD.n2689 DVDD.n2652 4.5005
R2135 DVDD.n2696 DVDD.n2652 4.5005
R2136 DVDD.n2688 DVDD.n2652 4.5005
R2137 DVDD.n2697 DVDD.n2652 4.5005
R2138 DVDD.n2687 DVDD.n2652 4.5005
R2139 DVDD.n2698 DVDD.n2652 4.5005
R2140 DVDD.n2686 DVDD.n2652 4.5005
R2141 DVDD.n2700 DVDD.n2652 4.5005
R2142 DVDD.n16268 DVDD.n2652 4.5005
R2143 DVDD.n16270 DVDD.n2652 4.5005
R2144 DVDD.n2691 DVDD.n2666 4.5005
R2145 DVDD.n2693 DVDD.n2666 4.5005
R2146 DVDD.n2690 DVDD.n2666 4.5005
R2147 DVDD.n2695 DVDD.n2666 4.5005
R2148 DVDD.n2689 DVDD.n2666 4.5005
R2149 DVDD.n2696 DVDD.n2666 4.5005
R2150 DVDD.n2688 DVDD.n2666 4.5005
R2151 DVDD.n2697 DVDD.n2666 4.5005
R2152 DVDD.n2687 DVDD.n2666 4.5005
R2153 DVDD.n2698 DVDD.n2666 4.5005
R2154 DVDD.n2686 DVDD.n2666 4.5005
R2155 DVDD.n2700 DVDD.n2666 4.5005
R2156 DVDD.n16268 DVDD.n2666 4.5005
R2157 DVDD.n16270 DVDD.n2666 4.5005
R2158 DVDD.n2691 DVDD.n2651 4.5005
R2159 DVDD.n2693 DVDD.n2651 4.5005
R2160 DVDD.n2690 DVDD.n2651 4.5005
R2161 DVDD.n2695 DVDD.n2651 4.5005
R2162 DVDD.n2689 DVDD.n2651 4.5005
R2163 DVDD.n2696 DVDD.n2651 4.5005
R2164 DVDD.n2688 DVDD.n2651 4.5005
R2165 DVDD.n2697 DVDD.n2651 4.5005
R2166 DVDD.n2687 DVDD.n2651 4.5005
R2167 DVDD.n2698 DVDD.n2651 4.5005
R2168 DVDD.n2686 DVDD.n2651 4.5005
R2169 DVDD.n2700 DVDD.n2651 4.5005
R2170 DVDD.n2685 DVDD.n2651 4.5005
R2171 DVDD.n16268 DVDD.n2651 4.5005
R2172 DVDD.n16270 DVDD.n2651 4.5005
R2173 DVDD.n2691 DVDD.n2668 4.5005
R2174 DVDD.n2693 DVDD.n2668 4.5005
R2175 DVDD.n2690 DVDD.n2668 4.5005
R2176 DVDD.n2695 DVDD.n2668 4.5005
R2177 DVDD.n2689 DVDD.n2668 4.5005
R2178 DVDD.n2696 DVDD.n2668 4.5005
R2179 DVDD.n2688 DVDD.n2668 4.5005
R2180 DVDD.n2697 DVDD.n2668 4.5005
R2181 DVDD.n2687 DVDD.n2668 4.5005
R2182 DVDD.n2698 DVDD.n2668 4.5005
R2183 DVDD.n2686 DVDD.n2668 4.5005
R2184 DVDD.n2700 DVDD.n2668 4.5005
R2185 DVDD.n2685 DVDD.n2668 4.5005
R2186 DVDD.n16268 DVDD.n2668 4.5005
R2187 DVDD.n16270 DVDD.n2668 4.5005
R2188 DVDD.n2691 DVDD.n2650 4.5005
R2189 DVDD.n2693 DVDD.n2650 4.5005
R2190 DVDD.n2690 DVDD.n2650 4.5005
R2191 DVDD.n2695 DVDD.n2650 4.5005
R2192 DVDD.n2689 DVDD.n2650 4.5005
R2193 DVDD.n2696 DVDD.n2650 4.5005
R2194 DVDD.n2688 DVDD.n2650 4.5005
R2195 DVDD.n2697 DVDD.n2650 4.5005
R2196 DVDD.n2687 DVDD.n2650 4.5005
R2197 DVDD.n2698 DVDD.n2650 4.5005
R2198 DVDD.n2686 DVDD.n2650 4.5005
R2199 DVDD.n2700 DVDD.n2650 4.5005
R2200 DVDD.n16268 DVDD.n2650 4.5005
R2201 DVDD.n16270 DVDD.n2650 4.5005
R2202 DVDD.n2691 DVDD.n2670 4.5005
R2203 DVDD.n2693 DVDD.n2670 4.5005
R2204 DVDD.n2690 DVDD.n2670 4.5005
R2205 DVDD.n2695 DVDD.n2670 4.5005
R2206 DVDD.n2689 DVDD.n2670 4.5005
R2207 DVDD.n2696 DVDD.n2670 4.5005
R2208 DVDD.n2688 DVDD.n2670 4.5005
R2209 DVDD.n2697 DVDD.n2670 4.5005
R2210 DVDD.n2687 DVDD.n2670 4.5005
R2211 DVDD.n2698 DVDD.n2670 4.5005
R2212 DVDD.n2686 DVDD.n2670 4.5005
R2213 DVDD.n2700 DVDD.n2670 4.5005
R2214 DVDD.n16268 DVDD.n2670 4.5005
R2215 DVDD.n16270 DVDD.n2670 4.5005
R2216 DVDD.n2691 DVDD.n2649 4.5005
R2217 DVDD.n2693 DVDD.n2649 4.5005
R2218 DVDD.n2690 DVDD.n2649 4.5005
R2219 DVDD.n2695 DVDD.n2649 4.5005
R2220 DVDD.n2689 DVDD.n2649 4.5005
R2221 DVDD.n2696 DVDD.n2649 4.5005
R2222 DVDD.n2688 DVDD.n2649 4.5005
R2223 DVDD.n2697 DVDD.n2649 4.5005
R2224 DVDD.n2687 DVDD.n2649 4.5005
R2225 DVDD.n2698 DVDD.n2649 4.5005
R2226 DVDD.n2686 DVDD.n2649 4.5005
R2227 DVDD.n2700 DVDD.n2649 4.5005
R2228 DVDD.n2685 DVDD.n2649 4.5005
R2229 DVDD.n16268 DVDD.n2649 4.5005
R2230 DVDD.n16270 DVDD.n2649 4.5005
R2231 DVDD.n2691 DVDD.n2672 4.5005
R2232 DVDD.n2693 DVDD.n2672 4.5005
R2233 DVDD.n2690 DVDD.n2672 4.5005
R2234 DVDD.n2695 DVDD.n2672 4.5005
R2235 DVDD.n2689 DVDD.n2672 4.5005
R2236 DVDD.n2696 DVDD.n2672 4.5005
R2237 DVDD.n2688 DVDD.n2672 4.5005
R2238 DVDD.n2697 DVDD.n2672 4.5005
R2239 DVDD.n2687 DVDD.n2672 4.5005
R2240 DVDD.n2698 DVDD.n2672 4.5005
R2241 DVDD.n2686 DVDD.n2672 4.5005
R2242 DVDD.n2700 DVDD.n2672 4.5005
R2243 DVDD.n2685 DVDD.n2672 4.5005
R2244 DVDD.n16268 DVDD.n2672 4.5005
R2245 DVDD.n16270 DVDD.n2672 4.5005
R2246 DVDD.n2691 DVDD.n2648 4.5005
R2247 DVDD.n2693 DVDD.n2648 4.5005
R2248 DVDD.n2690 DVDD.n2648 4.5005
R2249 DVDD.n2695 DVDD.n2648 4.5005
R2250 DVDD.n2689 DVDD.n2648 4.5005
R2251 DVDD.n2696 DVDD.n2648 4.5005
R2252 DVDD.n2688 DVDD.n2648 4.5005
R2253 DVDD.n2697 DVDD.n2648 4.5005
R2254 DVDD.n2687 DVDD.n2648 4.5005
R2255 DVDD.n2698 DVDD.n2648 4.5005
R2256 DVDD.n2686 DVDD.n2648 4.5005
R2257 DVDD.n2700 DVDD.n2648 4.5005
R2258 DVDD.n16268 DVDD.n2648 4.5005
R2259 DVDD.n16270 DVDD.n2648 4.5005
R2260 DVDD.n2691 DVDD.n2674 4.5005
R2261 DVDD.n2693 DVDD.n2674 4.5005
R2262 DVDD.n2690 DVDD.n2674 4.5005
R2263 DVDD.n2695 DVDD.n2674 4.5005
R2264 DVDD.n2689 DVDD.n2674 4.5005
R2265 DVDD.n2696 DVDD.n2674 4.5005
R2266 DVDD.n2688 DVDD.n2674 4.5005
R2267 DVDD.n2697 DVDD.n2674 4.5005
R2268 DVDD.n2687 DVDD.n2674 4.5005
R2269 DVDD.n2698 DVDD.n2674 4.5005
R2270 DVDD.n2686 DVDD.n2674 4.5005
R2271 DVDD.n2700 DVDD.n2674 4.5005
R2272 DVDD.n16268 DVDD.n2674 4.5005
R2273 DVDD.n16270 DVDD.n2674 4.5005
R2274 DVDD.n2691 DVDD.n2647 4.5005
R2275 DVDD.n2693 DVDD.n2647 4.5005
R2276 DVDD.n2690 DVDD.n2647 4.5005
R2277 DVDD.n2695 DVDD.n2647 4.5005
R2278 DVDD.n2689 DVDD.n2647 4.5005
R2279 DVDD.n2696 DVDD.n2647 4.5005
R2280 DVDD.n2688 DVDD.n2647 4.5005
R2281 DVDD.n2697 DVDD.n2647 4.5005
R2282 DVDD.n2687 DVDD.n2647 4.5005
R2283 DVDD.n2698 DVDD.n2647 4.5005
R2284 DVDD.n2686 DVDD.n2647 4.5005
R2285 DVDD.n2700 DVDD.n2647 4.5005
R2286 DVDD.n2685 DVDD.n2647 4.5005
R2287 DVDD.n16268 DVDD.n2647 4.5005
R2288 DVDD.n16270 DVDD.n2647 4.5005
R2289 DVDD.n2691 DVDD.n2676 4.5005
R2290 DVDD.n2693 DVDD.n2676 4.5005
R2291 DVDD.n2690 DVDD.n2676 4.5005
R2292 DVDD.n2695 DVDD.n2676 4.5005
R2293 DVDD.n2689 DVDD.n2676 4.5005
R2294 DVDD.n2696 DVDD.n2676 4.5005
R2295 DVDD.n2688 DVDD.n2676 4.5005
R2296 DVDD.n2697 DVDD.n2676 4.5005
R2297 DVDD.n2687 DVDD.n2676 4.5005
R2298 DVDD.n2698 DVDD.n2676 4.5005
R2299 DVDD.n2686 DVDD.n2676 4.5005
R2300 DVDD.n2700 DVDD.n2676 4.5005
R2301 DVDD.n2685 DVDD.n2676 4.5005
R2302 DVDD.n16268 DVDD.n2676 4.5005
R2303 DVDD.n16270 DVDD.n2676 4.5005
R2304 DVDD.n2691 DVDD.n2646 4.5005
R2305 DVDD.n2693 DVDD.n2646 4.5005
R2306 DVDD.n2690 DVDD.n2646 4.5005
R2307 DVDD.n2695 DVDD.n2646 4.5005
R2308 DVDD.n2689 DVDD.n2646 4.5005
R2309 DVDD.n2696 DVDD.n2646 4.5005
R2310 DVDD.n2688 DVDD.n2646 4.5005
R2311 DVDD.n2697 DVDD.n2646 4.5005
R2312 DVDD.n2687 DVDD.n2646 4.5005
R2313 DVDD.n2698 DVDD.n2646 4.5005
R2314 DVDD.n2686 DVDD.n2646 4.5005
R2315 DVDD.n2700 DVDD.n2646 4.5005
R2316 DVDD.n16268 DVDD.n2646 4.5005
R2317 DVDD.n16270 DVDD.n2646 4.5005
R2318 DVDD.n2691 DVDD.n2678 4.5005
R2319 DVDD.n2693 DVDD.n2678 4.5005
R2320 DVDD.n2690 DVDD.n2678 4.5005
R2321 DVDD.n2695 DVDD.n2678 4.5005
R2322 DVDD.n2689 DVDD.n2678 4.5005
R2323 DVDD.n2696 DVDD.n2678 4.5005
R2324 DVDD.n2688 DVDD.n2678 4.5005
R2325 DVDD.n2697 DVDD.n2678 4.5005
R2326 DVDD.n2687 DVDD.n2678 4.5005
R2327 DVDD.n2698 DVDD.n2678 4.5005
R2328 DVDD.n2686 DVDD.n2678 4.5005
R2329 DVDD.n2700 DVDD.n2678 4.5005
R2330 DVDD.n16268 DVDD.n2678 4.5005
R2331 DVDD.n16270 DVDD.n2678 4.5005
R2332 DVDD.n2691 DVDD.n2645 4.5005
R2333 DVDD.n2693 DVDD.n2645 4.5005
R2334 DVDD.n2690 DVDD.n2645 4.5005
R2335 DVDD.n2695 DVDD.n2645 4.5005
R2336 DVDD.n2689 DVDD.n2645 4.5005
R2337 DVDD.n2696 DVDD.n2645 4.5005
R2338 DVDD.n2688 DVDD.n2645 4.5005
R2339 DVDD.n2697 DVDD.n2645 4.5005
R2340 DVDD.n2687 DVDD.n2645 4.5005
R2341 DVDD.n2698 DVDD.n2645 4.5005
R2342 DVDD.n2686 DVDD.n2645 4.5005
R2343 DVDD.n2700 DVDD.n2645 4.5005
R2344 DVDD.n2685 DVDD.n2645 4.5005
R2345 DVDD.n16268 DVDD.n2645 4.5005
R2346 DVDD.n16270 DVDD.n2645 4.5005
R2347 DVDD.n16269 DVDD.n2691 4.5005
R2348 DVDD.n16269 DVDD.n2693 4.5005
R2349 DVDD.n16269 DVDD.n2690 4.5005
R2350 DVDD.n16269 DVDD.n2695 4.5005
R2351 DVDD.n16269 DVDD.n2689 4.5005
R2352 DVDD.n16269 DVDD.n2696 4.5005
R2353 DVDD.n16269 DVDD.n2688 4.5005
R2354 DVDD.n16269 DVDD.n2697 4.5005
R2355 DVDD.n16269 DVDD.n2687 4.5005
R2356 DVDD.n16269 DVDD.n2698 4.5005
R2357 DVDD.n16269 DVDD.n2686 4.5005
R2358 DVDD.n16269 DVDD.n2700 4.5005
R2359 DVDD.n16269 DVDD.n2685 4.5005
R2360 DVDD.n16269 DVDD.n16268 4.5005
R2361 DVDD.n16269 DVDD.n2644 4.5005
R2362 DVDD.n16270 DVDD.n16269 4.5005
R2363 DVDD.n2361 DVDD.n2341 4.5005
R2364 DVDD.n2361 DVDD.n2342 4.5005
R2365 DVDD.n2361 DVDD.n2340 4.5005
R2366 DVDD.n2361 DVDD.n2344 4.5005
R2367 DVDD.n2361 DVDD.n2338 4.5005
R2368 DVDD.n2361 DVDD.n2345 4.5005
R2369 DVDD.n2361 DVDD.n2337 4.5005
R2370 DVDD.n2361 DVDD.n2346 4.5005
R2371 DVDD.n2361 DVDD.n2336 4.5005
R2372 DVDD.n2361 DVDD.n2348 4.5005
R2373 DVDD.n16390 DVDD.n2361 4.5005
R2374 DVDD.n16394 DVDD.n2361 4.5005
R2375 DVDD.n2363 DVDD.n2341 4.5005
R2376 DVDD.n2363 DVDD.n2342 4.5005
R2377 DVDD.n2363 DVDD.n2340 4.5005
R2378 DVDD.n2363 DVDD.n2343 4.5005
R2379 DVDD.n2363 DVDD.n2339 4.5005
R2380 DVDD.n2363 DVDD.n2344 4.5005
R2381 DVDD.n2363 DVDD.n2338 4.5005
R2382 DVDD.n2363 DVDD.n2345 4.5005
R2383 DVDD.n2363 DVDD.n2337 4.5005
R2384 DVDD.n2363 DVDD.n2346 4.5005
R2385 DVDD.n2363 DVDD.n2336 4.5005
R2386 DVDD.n2363 DVDD.n2347 4.5005
R2387 DVDD.n2363 DVDD.n2335 4.5005
R2388 DVDD.n2363 DVDD.n2348 4.5005
R2389 DVDD.n16394 DVDD.n2363 4.5005
R2390 DVDD.n2358 DVDD.n2341 4.5005
R2391 DVDD.n2358 DVDD.n2342 4.5005
R2392 DVDD.n2358 DVDD.n2340 4.5005
R2393 DVDD.n2358 DVDD.n2343 4.5005
R2394 DVDD.n2358 DVDD.n2339 4.5005
R2395 DVDD.n2358 DVDD.n2344 4.5005
R2396 DVDD.n2358 DVDD.n2338 4.5005
R2397 DVDD.n2358 DVDD.n2345 4.5005
R2398 DVDD.n2358 DVDD.n2337 4.5005
R2399 DVDD.n2358 DVDD.n2346 4.5005
R2400 DVDD.n2358 DVDD.n2336 4.5005
R2401 DVDD.n2358 DVDD.n2347 4.5005
R2402 DVDD.n2358 DVDD.n2348 4.5005
R2403 DVDD.n16394 DVDD.n2358 4.5005
R2404 DVDD.n2365 DVDD.n2341 4.5005
R2405 DVDD.n2365 DVDD.n2342 4.5005
R2406 DVDD.n2365 DVDD.n2340 4.5005
R2407 DVDD.n2365 DVDD.n2343 4.5005
R2408 DVDD.n2365 DVDD.n2339 4.5005
R2409 DVDD.n2365 DVDD.n2344 4.5005
R2410 DVDD.n2365 DVDD.n2338 4.5005
R2411 DVDD.n2365 DVDD.n2345 4.5005
R2412 DVDD.n2365 DVDD.n2337 4.5005
R2413 DVDD.n2365 DVDD.n2346 4.5005
R2414 DVDD.n2365 DVDD.n2336 4.5005
R2415 DVDD.n2365 DVDD.n2347 4.5005
R2416 DVDD.n2365 DVDD.n2348 4.5005
R2417 DVDD.n16394 DVDD.n2365 4.5005
R2418 DVDD.n2357 DVDD.n2341 4.5005
R2419 DVDD.n2357 DVDD.n2342 4.5005
R2420 DVDD.n2357 DVDD.n2340 4.5005
R2421 DVDD.n2357 DVDD.n2343 4.5005
R2422 DVDD.n2357 DVDD.n2339 4.5005
R2423 DVDD.n2357 DVDD.n2344 4.5005
R2424 DVDD.n2357 DVDD.n2338 4.5005
R2425 DVDD.n2357 DVDD.n2345 4.5005
R2426 DVDD.n2357 DVDD.n2337 4.5005
R2427 DVDD.n2357 DVDD.n2346 4.5005
R2428 DVDD.n2357 DVDD.n2336 4.5005
R2429 DVDD.n2357 DVDD.n2347 4.5005
R2430 DVDD.n2357 DVDD.n2335 4.5005
R2431 DVDD.n2357 DVDD.n2348 4.5005
R2432 DVDD.n16394 DVDD.n2357 4.5005
R2433 DVDD.n2366 DVDD.n2341 4.5005
R2434 DVDD.n2366 DVDD.n2342 4.5005
R2435 DVDD.n2366 DVDD.n2340 4.5005
R2436 DVDD.n2366 DVDD.n2343 4.5005
R2437 DVDD.n2366 DVDD.n2339 4.5005
R2438 DVDD.n2366 DVDD.n2344 4.5005
R2439 DVDD.n2366 DVDD.n2338 4.5005
R2440 DVDD.n2366 DVDD.n2345 4.5005
R2441 DVDD.n2366 DVDD.n2337 4.5005
R2442 DVDD.n2366 DVDD.n2346 4.5005
R2443 DVDD.n2366 DVDD.n2336 4.5005
R2444 DVDD.n2366 DVDD.n2347 4.5005
R2445 DVDD.n2366 DVDD.n2335 4.5005
R2446 DVDD.n2366 DVDD.n2348 4.5005
R2447 DVDD.n16394 DVDD.n2366 4.5005
R2448 DVDD.n2356 DVDD.n2341 4.5005
R2449 DVDD.n2356 DVDD.n2342 4.5005
R2450 DVDD.n2356 DVDD.n2340 4.5005
R2451 DVDD.n2356 DVDD.n2343 4.5005
R2452 DVDD.n2356 DVDD.n2339 4.5005
R2453 DVDD.n2356 DVDD.n2344 4.5005
R2454 DVDD.n2356 DVDD.n2338 4.5005
R2455 DVDD.n2356 DVDD.n2345 4.5005
R2456 DVDD.n2356 DVDD.n2337 4.5005
R2457 DVDD.n2356 DVDD.n2346 4.5005
R2458 DVDD.n2356 DVDD.n2336 4.5005
R2459 DVDD.n2356 DVDD.n2347 4.5005
R2460 DVDD.n2356 DVDD.n2348 4.5005
R2461 DVDD.n16394 DVDD.n2356 4.5005
R2462 DVDD.n2368 DVDD.n2341 4.5005
R2463 DVDD.n2368 DVDD.n2342 4.5005
R2464 DVDD.n2368 DVDD.n2340 4.5005
R2465 DVDD.n2368 DVDD.n2343 4.5005
R2466 DVDD.n2368 DVDD.n2339 4.5005
R2467 DVDD.n2368 DVDD.n2344 4.5005
R2468 DVDD.n2368 DVDD.n2338 4.5005
R2469 DVDD.n2368 DVDD.n2345 4.5005
R2470 DVDD.n2368 DVDD.n2337 4.5005
R2471 DVDD.n2368 DVDD.n2346 4.5005
R2472 DVDD.n2368 DVDD.n2336 4.5005
R2473 DVDD.n2368 DVDD.n2347 4.5005
R2474 DVDD.n2368 DVDD.n2348 4.5005
R2475 DVDD.n16394 DVDD.n2368 4.5005
R2476 DVDD.n2355 DVDD.n2341 4.5005
R2477 DVDD.n2355 DVDD.n2342 4.5005
R2478 DVDD.n2355 DVDD.n2340 4.5005
R2479 DVDD.n2355 DVDD.n2343 4.5005
R2480 DVDD.n2355 DVDD.n2339 4.5005
R2481 DVDD.n2355 DVDD.n2344 4.5005
R2482 DVDD.n2355 DVDD.n2338 4.5005
R2483 DVDD.n2355 DVDD.n2345 4.5005
R2484 DVDD.n2355 DVDD.n2337 4.5005
R2485 DVDD.n2355 DVDD.n2346 4.5005
R2486 DVDD.n2355 DVDD.n2336 4.5005
R2487 DVDD.n2355 DVDD.n2347 4.5005
R2488 DVDD.n2355 DVDD.n2335 4.5005
R2489 DVDD.n2355 DVDD.n2348 4.5005
R2490 DVDD.n16394 DVDD.n2355 4.5005
R2491 DVDD.n2369 DVDD.n2341 4.5005
R2492 DVDD.n2369 DVDD.n2342 4.5005
R2493 DVDD.n2369 DVDD.n2340 4.5005
R2494 DVDD.n2369 DVDD.n2343 4.5005
R2495 DVDD.n2369 DVDD.n2339 4.5005
R2496 DVDD.n2369 DVDD.n2344 4.5005
R2497 DVDD.n2369 DVDD.n2338 4.5005
R2498 DVDD.n2369 DVDD.n2345 4.5005
R2499 DVDD.n2369 DVDD.n2337 4.5005
R2500 DVDD.n2369 DVDD.n2346 4.5005
R2501 DVDD.n2369 DVDD.n2336 4.5005
R2502 DVDD.n2369 DVDD.n2347 4.5005
R2503 DVDD.n2369 DVDD.n2335 4.5005
R2504 DVDD.n2369 DVDD.n2348 4.5005
R2505 DVDD.n16394 DVDD.n2369 4.5005
R2506 DVDD.n2354 DVDD.n2341 4.5005
R2507 DVDD.n2354 DVDD.n2342 4.5005
R2508 DVDD.n2354 DVDD.n2340 4.5005
R2509 DVDD.n2354 DVDD.n2343 4.5005
R2510 DVDD.n2354 DVDD.n2339 4.5005
R2511 DVDD.n2354 DVDD.n2344 4.5005
R2512 DVDD.n2354 DVDD.n2338 4.5005
R2513 DVDD.n2354 DVDD.n2345 4.5005
R2514 DVDD.n2354 DVDD.n2337 4.5005
R2515 DVDD.n2354 DVDD.n2346 4.5005
R2516 DVDD.n2354 DVDD.n2336 4.5005
R2517 DVDD.n2354 DVDD.n2347 4.5005
R2518 DVDD.n2354 DVDD.n2348 4.5005
R2519 DVDD.n16394 DVDD.n2354 4.5005
R2520 DVDD.n2371 DVDD.n2341 4.5005
R2521 DVDD.n2371 DVDD.n2342 4.5005
R2522 DVDD.n2371 DVDD.n2340 4.5005
R2523 DVDD.n2371 DVDD.n2343 4.5005
R2524 DVDD.n2371 DVDD.n2339 4.5005
R2525 DVDD.n2371 DVDD.n2344 4.5005
R2526 DVDD.n2371 DVDD.n2338 4.5005
R2527 DVDD.n2371 DVDD.n2345 4.5005
R2528 DVDD.n2371 DVDD.n2337 4.5005
R2529 DVDD.n2371 DVDD.n2346 4.5005
R2530 DVDD.n2371 DVDD.n2336 4.5005
R2531 DVDD.n2371 DVDD.n2347 4.5005
R2532 DVDD.n2371 DVDD.n2348 4.5005
R2533 DVDD.n16394 DVDD.n2371 4.5005
R2534 DVDD.n2353 DVDD.n2341 4.5005
R2535 DVDD.n2353 DVDD.n2342 4.5005
R2536 DVDD.n2353 DVDD.n2340 4.5005
R2537 DVDD.n2353 DVDD.n2343 4.5005
R2538 DVDD.n2353 DVDD.n2339 4.5005
R2539 DVDD.n2353 DVDD.n2344 4.5005
R2540 DVDD.n2353 DVDD.n2338 4.5005
R2541 DVDD.n2353 DVDD.n2345 4.5005
R2542 DVDD.n2353 DVDD.n2337 4.5005
R2543 DVDD.n2353 DVDD.n2346 4.5005
R2544 DVDD.n2353 DVDD.n2336 4.5005
R2545 DVDD.n2353 DVDD.n2347 4.5005
R2546 DVDD.n2353 DVDD.n2348 4.5005
R2547 DVDD.n16394 DVDD.n2353 4.5005
R2548 DVDD.n2373 DVDD.n2341 4.5005
R2549 DVDD.n2373 DVDD.n2342 4.5005
R2550 DVDD.n2373 DVDD.n2340 4.5005
R2551 DVDD.n2373 DVDD.n2343 4.5005
R2552 DVDD.n2373 DVDD.n2339 4.5005
R2553 DVDD.n2373 DVDD.n2344 4.5005
R2554 DVDD.n2373 DVDD.n2338 4.5005
R2555 DVDD.n2373 DVDD.n2345 4.5005
R2556 DVDD.n2373 DVDD.n2337 4.5005
R2557 DVDD.n2373 DVDD.n2346 4.5005
R2558 DVDD.n2373 DVDD.n2336 4.5005
R2559 DVDD.n2373 DVDD.n2347 4.5005
R2560 DVDD.n2373 DVDD.n2348 4.5005
R2561 DVDD.n16394 DVDD.n2373 4.5005
R2562 DVDD.n2352 DVDD.n2341 4.5005
R2563 DVDD.n2352 DVDD.n2342 4.5005
R2564 DVDD.n2352 DVDD.n2340 4.5005
R2565 DVDD.n2352 DVDD.n2343 4.5005
R2566 DVDD.n2352 DVDD.n2339 4.5005
R2567 DVDD.n2352 DVDD.n2344 4.5005
R2568 DVDD.n2352 DVDD.n2338 4.5005
R2569 DVDD.n2352 DVDD.n2345 4.5005
R2570 DVDD.n2352 DVDD.n2337 4.5005
R2571 DVDD.n2352 DVDD.n2346 4.5005
R2572 DVDD.n2352 DVDD.n2336 4.5005
R2573 DVDD.n2352 DVDD.n2347 4.5005
R2574 DVDD.n2352 DVDD.n2348 4.5005
R2575 DVDD.n16394 DVDD.n2352 4.5005
R2576 DVDD.n2375 DVDD.n2341 4.5005
R2577 DVDD.n2375 DVDD.n2342 4.5005
R2578 DVDD.n2375 DVDD.n2340 4.5005
R2579 DVDD.n2375 DVDD.n2343 4.5005
R2580 DVDD.n2375 DVDD.n2339 4.5005
R2581 DVDD.n2375 DVDD.n2344 4.5005
R2582 DVDD.n2375 DVDD.n2338 4.5005
R2583 DVDD.n2375 DVDD.n2345 4.5005
R2584 DVDD.n2375 DVDD.n2337 4.5005
R2585 DVDD.n2375 DVDD.n2346 4.5005
R2586 DVDD.n2375 DVDD.n2336 4.5005
R2587 DVDD.n2375 DVDD.n2347 4.5005
R2588 DVDD.n2375 DVDD.n2348 4.5005
R2589 DVDD.n16394 DVDD.n2375 4.5005
R2590 DVDD.n16395 DVDD.n2341 4.5005
R2591 DVDD.n16395 DVDD.n2342 4.5005
R2592 DVDD.n16395 DVDD.n2340 4.5005
R2593 DVDD.n16395 DVDD.n2343 4.5005
R2594 DVDD.n16395 DVDD.n2339 4.5005
R2595 DVDD.n16395 DVDD.n2344 4.5005
R2596 DVDD.n16395 DVDD.n2338 4.5005
R2597 DVDD.n16395 DVDD.n2345 4.5005
R2598 DVDD.n16395 DVDD.n2337 4.5005
R2599 DVDD.n16395 DVDD.n2346 4.5005
R2600 DVDD.n16395 DVDD.n2336 4.5005
R2601 DVDD.n16395 DVDD.n2347 4.5005
R2602 DVDD.n16395 DVDD.n2335 4.5005
R2603 DVDD.n16395 DVDD.n2348 4.5005
R2604 DVDD.n16395 DVDD.n16394 4.5005
R2605 DVDD.n2377 DVDD.n2341 4.5005
R2606 DVDD.n2377 DVDD.n2342 4.5005
R2607 DVDD.n2377 DVDD.n2340 4.5005
R2608 DVDD.n2377 DVDD.n2343 4.5005
R2609 DVDD.n2377 DVDD.n2339 4.5005
R2610 DVDD.n2377 DVDD.n2344 4.5005
R2611 DVDD.n2377 DVDD.n2338 4.5005
R2612 DVDD.n2377 DVDD.n2345 4.5005
R2613 DVDD.n2377 DVDD.n2337 4.5005
R2614 DVDD.n2377 DVDD.n2346 4.5005
R2615 DVDD.n2377 DVDD.n2336 4.5005
R2616 DVDD.n2377 DVDD.n2347 4.5005
R2617 DVDD.n2377 DVDD.n2348 4.5005
R2618 DVDD.n16394 DVDD.n2377 4.5005
R2619 DVDD.n2351 DVDD.n2341 4.5005
R2620 DVDD.n2351 DVDD.n2342 4.5005
R2621 DVDD.n2351 DVDD.n2340 4.5005
R2622 DVDD.n2351 DVDD.n2343 4.5005
R2623 DVDD.n2351 DVDD.n2339 4.5005
R2624 DVDD.n2351 DVDD.n2344 4.5005
R2625 DVDD.n2351 DVDD.n2338 4.5005
R2626 DVDD.n2351 DVDD.n2345 4.5005
R2627 DVDD.n2351 DVDD.n2337 4.5005
R2628 DVDD.n2351 DVDD.n2346 4.5005
R2629 DVDD.n2351 DVDD.n2336 4.5005
R2630 DVDD.n2351 DVDD.n2347 4.5005
R2631 DVDD.n2351 DVDD.n2348 4.5005
R2632 DVDD.n16394 DVDD.n2351 4.5005
R2633 DVDD.n16393 DVDD.n2341 4.5005
R2634 DVDD.n16393 DVDD.n2342 4.5005
R2635 DVDD.n16393 DVDD.n2340 4.5005
R2636 DVDD.n16393 DVDD.n2343 4.5005
R2637 DVDD.n16393 DVDD.n2339 4.5005
R2638 DVDD.n16393 DVDD.n2344 4.5005
R2639 DVDD.n16393 DVDD.n2338 4.5005
R2640 DVDD.n16393 DVDD.n2345 4.5005
R2641 DVDD.n16393 DVDD.n2337 4.5005
R2642 DVDD.n16393 DVDD.n2346 4.5005
R2643 DVDD.n16393 DVDD.n2336 4.5005
R2644 DVDD.n16393 DVDD.n2347 4.5005
R2645 DVDD.n16393 DVDD.n2348 4.5005
R2646 DVDD.n16394 DVDD.n16393 4.5005
R2647 DVDD.n2350 DVDD.n2341 4.5005
R2648 DVDD.n2350 DVDD.n2342 4.5005
R2649 DVDD.n2350 DVDD.n2340 4.5005
R2650 DVDD.n2350 DVDD.n2343 4.5005
R2651 DVDD.n2350 DVDD.n2339 4.5005
R2652 DVDD.n2350 DVDD.n2344 4.5005
R2653 DVDD.n2350 DVDD.n2338 4.5005
R2654 DVDD.n2350 DVDD.n2345 4.5005
R2655 DVDD.n2350 DVDD.n2337 4.5005
R2656 DVDD.n2350 DVDD.n2346 4.5005
R2657 DVDD.n2350 DVDD.n2336 4.5005
R2658 DVDD.n2350 DVDD.n2347 4.5005
R2659 DVDD.n2350 DVDD.n2335 4.5005
R2660 DVDD.n2350 DVDD.n2348 4.5005
R2661 DVDD.n16394 DVDD.n2350 4.5005
R2662 DVDD.n4389 DVDD.n4329 4.5005
R2663 DVDD.n4406 DVDD.n4329 4.5005
R2664 DVDD.n4391 DVDD.n4329 4.5005
R2665 DVDD.n4403 DVDD.n4329 4.5005
R2666 DVDD.n4392 DVDD.n4329 4.5005
R2667 DVDD.n4402 DVDD.n4329 4.5005
R2668 DVDD.n4393 DVDD.n4329 4.5005
R2669 DVDD.n4534 DVDD.n4329 4.5005
R2670 DVDD.n4399 DVDD.n4329 4.5005
R2671 DVDD.n4329 DVDD.n4323 4.5005
R2672 DVDD.n4558 DVDD.n4329 4.5005
R2673 DVDD.n4389 DVDD.n4328 4.5005
R2674 DVDD.n4406 DVDD.n4328 4.5005
R2675 DVDD.n4390 DVDD.n4328 4.5005
R2676 DVDD.n4405 DVDD.n4328 4.5005
R2677 DVDD.n4391 DVDD.n4328 4.5005
R2678 DVDD.n4403 DVDD.n4328 4.5005
R2679 DVDD.n4392 DVDD.n4328 4.5005
R2680 DVDD.n4402 DVDD.n4328 4.5005
R2681 DVDD.n4393 DVDD.n4328 4.5005
R2682 DVDD.n4534 DVDD.n4328 4.5005
R2683 DVDD.n4394 DVDD.n4328 4.5005
R2684 DVDD.n4401 DVDD.n4328 4.5005
R2685 DVDD.n4399 DVDD.n4328 4.5005
R2686 DVDD.n4558 DVDD.n4328 4.5005
R2687 DVDD.n4399 DVDD.n4331 4.5005
R2688 DVDD.n4558 DVDD.n4331 4.5005
R2689 DVDD.n4327 DVDD.n4323 4.5005
R2690 DVDD.n4558 DVDD.n4327 4.5005
R2691 DVDD.n4332 DVDD.n4323 4.5005
R2692 DVDD.n4558 DVDD.n4332 4.5005
R2693 DVDD.n4326 DVDD.n4323 4.5005
R2694 DVDD.n4558 DVDD.n4326 4.5005
R2695 DVDD.n4386 DVDD.n4323 4.5005
R2696 DVDD.n4558 DVDD.n4386 4.5005
R2697 DVDD.n4399 DVDD.n4325 4.5005
R2698 DVDD.n4325 DVDD.n4323 4.5005
R2699 DVDD.n4558 DVDD.n4325 4.5005
R2700 DVDD.n4387 DVDD.n4323 4.5005
R2701 DVDD.n4558 DVDD.n4387 4.5005
R2702 DVDD.n4324 DVDD.n4323 4.5005
R2703 DVDD.n4558 DVDD.n4324 4.5005
R2704 DVDD.n4557 DVDD.n4399 4.5005
R2705 DVDD.n4557 DVDD.n4323 4.5005
R2706 DVDD.n4558 DVDD.n4557 4.5005
R2707 DVDD.n4531 DVDD.n4495 4.5005
R2708 DVDD.n4531 DVDD.n4497 4.5005
R2709 DVDD.n4531 DVDD.n4494 4.5005
R2710 DVDD.n4531 DVDD.n4500 4.5005
R2711 DVDD.n4531 DVDD.n4492 4.5005
R2712 DVDD.n4531 DVDD.n4501 4.5005
R2713 DVDD.n4531 DVDD.n4491 4.5005
R2714 DVDD.n4531 DVDD.n4502 4.5005
R2715 DVDD.n4531 DVDD.n4504 4.5005
R2716 DVDD.n4532 DVDD.n4531 4.5005
R2717 DVDD.n4495 DVDD.n4479 4.5005
R2718 DVDD.n4497 DVDD.n4479 4.5005
R2719 DVDD.n4494 DVDD.n4479 4.5005
R2720 DVDD.n4498 DVDD.n4479 4.5005
R2721 DVDD.n4493 DVDD.n4479 4.5005
R2722 DVDD.n4500 DVDD.n4479 4.5005
R2723 DVDD.n4492 DVDD.n4479 4.5005
R2724 DVDD.n4501 DVDD.n4479 4.5005
R2725 DVDD.n4491 DVDD.n4479 4.5005
R2726 DVDD.n4502 DVDD.n4479 4.5005
R2727 DVDD.n4534 DVDD.n4479 4.5005
R2728 DVDD.n4503 DVDD.n4479 4.5005
R2729 DVDD.n4504 DVDD.n4479 4.5005
R2730 DVDD.n4532 DVDD.n4479 4.5005
R2731 DVDD.n4495 DVDD.n4473 4.5005
R2732 DVDD.n4497 DVDD.n4473 4.5005
R2733 DVDD.n4494 DVDD.n4473 4.5005
R2734 DVDD.n4498 DVDD.n4473 4.5005
R2735 DVDD.n4493 DVDD.n4473 4.5005
R2736 DVDD.n4500 DVDD.n4473 4.5005
R2737 DVDD.n4492 DVDD.n4473 4.5005
R2738 DVDD.n4501 DVDD.n4473 4.5005
R2739 DVDD.n4491 DVDD.n4473 4.5005
R2740 DVDD.n4502 DVDD.n4473 4.5005
R2741 DVDD.n4534 DVDD.n4473 4.5005
R2742 DVDD.n4503 DVDD.n4473 4.5005
R2743 DVDD.n4504 DVDD.n4473 4.5005
R2744 DVDD.n4532 DVDD.n4473 4.5005
R2745 DVDD.n4495 DVDD.n4480 4.5005
R2746 DVDD.n4497 DVDD.n4480 4.5005
R2747 DVDD.n4494 DVDD.n4480 4.5005
R2748 DVDD.n4498 DVDD.n4480 4.5005
R2749 DVDD.n4493 DVDD.n4480 4.5005
R2750 DVDD.n4500 DVDD.n4480 4.5005
R2751 DVDD.n4492 DVDD.n4480 4.5005
R2752 DVDD.n4501 DVDD.n4480 4.5005
R2753 DVDD.n4491 DVDD.n4480 4.5005
R2754 DVDD.n4502 DVDD.n4480 4.5005
R2755 DVDD.n4534 DVDD.n4480 4.5005
R2756 DVDD.n4503 DVDD.n4480 4.5005
R2757 DVDD.n4504 DVDD.n4480 4.5005
R2758 DVDD.n4532 DVDD.n4480 4.5005
R2759 DVDD.n4495 DVDD.n4472 4.5005
R2760 DVDD.n4497 DVDD.n4472 4.5005
R2761 DVDD.n4494 DVDD.n4472 4.5005
R2762 DVDD.n4498 DVDD.n4472 4.5005
R2763 DVDD.n4493 DVDD.n4472 4.5005
R2764 DVDD.n4500 DVDD.n4472 4.5005
R2765 DVDD.n4492 DVDD.n4472 4.5005
R2766 DVDD.n4501 DVDD.n4472 4.5005
R2767 DVDD.n4491 DVDD.n4472 4.5005
R2768 DVDD.n4502 DVDD.n4472 4.5005
R2769 DVDD.n4534 DVDD.n4472 4.5005
R2770 DVDD.n4503 DVDD.n4472 4.5005
R2771 DVDD.n4504 DVDD.n4472 4.5005
R2772 DVDD.n4532 DVDD.n4472 4.5005
R2773 DVDD.n4495 DVDD.n4481 4.5005
R2774 DVDD.n4497 DVDD.n4481 4.5005
R2775 DVDD.n4494 DVDD.n4481 4.5005
R2776 DVDD.n4498 DVDD.n4481 4.5005
R2777 DVDD.n4493 DVDD.n4481 4.5005
R2778 DVDD.n4500 DVDD.n4481 4.5005
R2779 DVDD.n4492 DVDD.n4481 4.5005
R2780 DVDD.n4501 DVDD.n4481 4.5005
R2781 DVDD.n4491 DVDD.n4481 4.5005
R2782 DVDD.n4502 DVDD.n4481 4.5005
R2783 DVDD.n4534 DVDD.n4481 4.5005
R2784 DVDD.n4503 DVDD.n4481 4.5005
R2785 DVDD.n4504 DVDD.n4481 4.5005
R2786 DVDD.n4532 DVDD.n4481 4.5005
R2787 DVDD.n4495 DVDD.n4471 4.5005
R2788 DVDD.n4497 DVDD.n4471 4.5005
R2789 DVDD.n4494 DVDD.n4471 4.5005
R2790 DVDD.n4498 DVDD.n4471 4.5005
R2791 DVDD.n4493 DVDD.n4471 4.5005
R2792 DVDD.n4500 DVDD.n4471 4.5005
R2793 DVDD.n4492 DVDD.n4471 4.5005
R2794 DVDD.n4501 DVDD.n4471 4.5005
R2795 DVDD.n4491 DVDD.n4471 4.5005
R2796 DVDD.n4502 DVDD.n4471 4.5005
R2797 DVDD.n4534 DVDD.n4471 4.5005
R2798 DVDD.n4503 DVDD.n4471 4.5005
R2799 DVDD.n4504 DVDD.n4471 4.5005
R2800 DVDD.n4532 DVDD.n4471 4.5005
R2801 DVDD.n4495 DVDD.n4482 4.5005
R2802 DVDD.n4497 DVDD.n4482 4.5005
R2803 DVDD.n4494 DVDD.n4482 4.5005
R2804 DVDD.n4498 DVDD.n4482 4.5005
R2805 DVDD.n4493 DVDD.n4482 4.5005
R2806 DVDD.n4500 DVDD.n4482 4.5005
R2807 DVDD.n4492 DVDD.n4482 4.5005
R2808 DVDD.n4501 DVDD.n4482 4.5005
R2809 DVDD.n4491 DVDD.n4482 4.5005
R2810 DVDD.n4502 DVDD.n4482 4.5005
R2811 DVDD.n4534 DVDD.n4482 4.5005
R2812 DVDD.n4503 DVDD.n4482 4.5005
R2813 DVDD.n4504 DVDD.n4482 4.5005
R2814 DVDD.n4532 DVDD.n4482 4.5005
R2815 DVDD.n4495 DVDD.n4470 4.5005
R2816 DVDD.n4497 DVDD.n4470 4.5005
R2817 DVDD.n4494 DVDD.n4470 4.5005
R2818 DVDD.n4498 DVDD.n4470 4.5005
R2819 DVDD.n4493 DVDD.n4470 4.5005
R2820 DVDD.n4500 DVDD.n4470 4.5005
R2821 DVDD.n4492 DVDD.n4470 4.5005
R2822 DVDD.n4501 DVDD.n4470 4.5005
R2823 DVDD.n4491 DVDD.n4470 4.5005
R2824 DVDD.n4502 DVDD.n4470 4.5005
R2825 DVDD.n4534 DVDD.n4470 4.5005
R2826 DVDD.n4503 DVDD.n4470 4.5005
R2827 DVDD.n4504 DVDD.n4470 4.5005
R2828 DVDD.n4532 DVDD.n4470 4.5005
R2829 DVDD.n4495 DVDD.n4483 4.5005
R2830 DVDD.n4497 DVDD.n4483 4.5005
R2831 DVDD.n4494 DVDD.n4483 4.5005
R2832 DVDD.n4498 DVDD.n4483 4.5005
R2833 DVDD.n4493 DVDD.n4483 4.5005
R2834 DVDD.n4500 DVDD.n4483 4.5005
R2835 DVDD.n4492 DVDD.n4483 4.5005
R2836 DVDD.n4501 DVDD.n4483 4.5005
R2837 DVDD.n4491 DVDD.n4483 4.5005
R2838 DVDD.n4502 DVDD.n4483 4.5005
R2839 DVDD.n4534 DVDD.n4483 4.5005
R2840 DVDD.n4503 DVDD.n4483 4.5005
R2841 DVDD.n4504 DVDD.n4483 4.5005
R2842 DVDD.n4532 DVDD.n4483 4.5005
R2843 DVDD.n4495 DVDD.n4469 4.5005
R2844 DVDD.n4497 DVDD.n4469 4.5005
R2845 DVDD.n4494 DVDD.n4469 4.5005
R2846 DVDD.n4498 DVDD.n4469 4.5005
R2847 DVDD.n4493 DVDD.n4469 4.5005
R2848 DVDD.n4500 DVDD.n4469 4.5005
R2849 DVDD.n4492 DVDD.n4469 4.5005
R2850 DVDD.n4501 DVDD.n4469 4.5005
R2851 DVDD.n4491 DVDD.n4469 4.5005
R2852 DVDD.n4502 DVDD.n4469 4.5005
R2853 DVDD.n4534 DVDD.n4469 4.5005
R2854 DVDD.n4503 DVDD.n4469 4.5005
R2855 DVDD.n4504 DVDD.n4469 4.5005
R2856 DVDD.n4532 DVDD.n4469 4.5005
R2857 DVDD.n4495 DVDD.n4484 4.5005
R2858 DVDD.n4497 DVDD.n4484 4.5005
R2859 DVDD.n4494 DVDD.n4484 4.5005
R2860 DVDD.n4498 DVDD.n4484 4.5005
R2861 DVDD.n4493 DVDD.n4484 4.5005
R2862 DVDD.n4500 DVDD.n4484 4.5005
R2863 DVDD.n4492 DVDD.n4484 4.5005
R2864 DVDD.n4501 DVDD.n4484 4.5005
R2865 DVDD.n4491 DVDD.n4484 4.5005
R2866 DVDD.n4502 DVDD.n4484 4.5005
R2867 DVDD.n4534 DVDD.n4484 4.5005
R2868 DVDD.n4503 DVDD.n4484 4.5005
R2869 DVDD.n4504 DVDD.n4484 4.5005
R2870 DVDD.n4532 DVDD.n4484 4.5005
R2871 DVDD.n4495 DVDD.n4468 4.5005
R2872 DVDD.n4497 DVDD.n4468 4.5005
R2873 DVDD.n4494 DVDD.n4468 4.5005
R2874 DVDD.n4498 DVDD.n4468 4.5005
R2875 DVDD.n4493 DVDD.n4468 4.5005
R2876 DVDD.n4500 DVDD.n4468 4.5005
R2877 DVDD.n4492 DVDD.n4468 4.5005
R2878 DVDD.n4501 DVDD.n4468 4.5005
R2879 DVDD.n4491 DVDD.n4468 4.5005
R2880 DVDD.n4502 DVDD.n4468 4.5005
R2881 DVDD.n4534 DVDD.n4468 4.5005
R2882 DVDD.n4503 DVDD.n4468 4.5005
R2883 DVDD.n4504 DVDD.n4468 4.5005
R2884 DVDD.n4532 DVDD.n4468 4.5005
R2885 DVDD.n4495 DVDD.n4485 4.5005
R2886 DVDD.n4497 DVDD.n4485 4.5005
R2887 DVDD.n4494 DVDD.n4485 4.5005
R2888 DVDD.n4498 DVDD.n4485 4.5005
R2889 DVDD.n4493 DVDD.n4485 4.5005
R2890 DVDD.n4500 DVDD.n4485 4.5005
R2891 DVDD.n4492 DVDD.n4485 4.5005
R2892 DVDD.n4501 DVDD.n4485 4.5005
R2893 DVDD.n4491 DVDD.n4485 4.5005
R2894 DVDD.n4502 DVDD.n4485 4.5005
R2895 DVDD.n4534 DVDD.n4485 4.5005
R2896 DVDD.n4503 DVDD.n4485 4.5005
R2897 DVDD.n4504 DVDD.n4485 4.5005
R2898 DVDD.n4532 DVDD.n4485 4.5005
R2899 DVDD.n4495 DVDD.n4467 4.5005
R2900 DVDD.n4497 DVDD.n4467 4.5005
R2901 DVDD.n4494 DVDD.n4467 4.5005
R2902 DVDD.n4498 DVDD.n4467 4.5005
R2903 DVDD.n4493 DVDD.n4467 4.5005
R2904 DVDD.n4500 DVDD.n4467 4.5005
R2905 DVDD.n4492 DVDD.n4467 4.5005
R2906 DVDD.n4501 DVDD.n4467 4.5005
R2907 DVDD.n4491 DVDD.n4467 4.5005
R2908 DVDD.n4502 DVDD.n4467 4.5005
R2909 DVDD.n4534 DVDD.n4467 4.5005
R2910 DVDD.n4503 DVDD.n4467 4.5005
R2911 DVDD.n4504 DVDD.n4467 4.5005
R2912 DVDD.n4532 DVDD.n4467 4.5005
R2913 DVDD.n4495 DVDD.n4486 4.5005
R2914 DVDD.n4497 DVDD.n4486 4.5005
R2915 DVDD.n4494 DVDD.n4486 4.5005
R2916 DVDD.n4498 DVDD.n4486 4.5005
R2917 DVDD.n4493 DVDD.n4486 4.5005
R2918 DVDD.n4500 DVDD.n4486 4.5005
R2919 DVDD.n4492 DVDD.n4486 4.5005
R2920 DVDD.n4501 DVDD.n4486 4.5005
R2921 DVDD.n4491 DVDD.n4486 4.5005
R2922 DVDD.n4502 DVDD.n4486 4.5005
R2923 DVDD.n4534 DVDD.n4486 4.5005
R2924 DVDD.n4503 DVDD.n4486 4.5005
R2925 DVDD.n4504 DVDD.n4486 4.5005
R2926 DVDD.n4532 DVDD.n4486 4.5005
R2927 DVDD.n4495 DVDD.n4466 4.5005
R2928 DVDD.n4497 DVDD.n4466 4.5005
R2929 DVDD.n4494 DVDD.n4466 4.5005
R2930 DVDD.n4498 DVDD.n4466 4.5005
R2931 DVDD.n4493 DVDD.n4466 4.5005
R2932 DVDD.n4500 DVDD.n4466 4.5005
R2933 DVDD.n4492 DVDD.n4466 4.5005
R2934 DVDD.n4501 DVDD.n4466 4.5005
R2935 DVDD.n4491 DVDD.n4466 4.5005
R2936 DVDD.n4502 DVDD.n4466 4.5005
R2937 DVDD.n4534 DVDD.n4466 4.5005
R2938 DVDD.n4503 DVDD.n4466 4.5005
R2939 DVDD.n4504 DVDD.n4466 4.5005
R2940 DVDD.n4532 DVDD.n4466 4.5005
R2941 DVDD.n4495 DVDD.n4487 4.5005
R2942 DVDD.n4497 DVDD.n4487 4.5005
R2943 DVDD.n4494 DVDD.n4487 4.5005
R2944 DVDD.n4498 DVDD.n4487 4.5005
R2945 DVDD.n4493 DVDD.n4487 4.5005
R2946 DVDD.n4500 DVDD.n4487 4.5005
R2947 DVDD.n4492 DVDD.n4487 4.5005
R2948 DVDD.n4501 DVDD.n4487 4.5005
R2949 DVDD.n4491 DVDD.n4487 4.5005
R2950 DVDD.n4502 DVDD.n4487 4.5005
R2951 DVDD.n4534 DVDD.n4487 4.5005
R2952 DVDD.n4503 DVDD.n4487 4.5005
R2953 DVDD.n4504 DVDD.n4487 4.5005
R2954 DVDD.n4532 DVDD.n4487 4.5005
R2955 DVDD.n4495 DVDD.n4465 4.5005
R2956 DVDD.n4497 DVDD.n4465 4.5005
R2957 DVDD.n4494 DVDD.n4465 4.5005
R2958 DVDD.n4498 DVDD.n4465 4.5005
R2959 DVDD.n4493 DVDD.n4465 4.5005
R2960 DVDD.n4500 DVDD.n4465 4.5005
R2961 DVDD.n4492 DVDD.n4465 4.5005
R2962 DVDD.n4501 DVDD.n4465 4.5005
R2963 DVDD.n4491 DVDD.n4465 4.5005
R2964 DVDD.n4502 DVDD.n4465 4.5005
R2965 DVDD.n4534 DVDD.n4465 4.5005
R2966 DVDD.n4503 DVDD.n4465 4.5005
R2967 DVDD.n4504 DVDD.n4465 4.5005
R2968 DVDD.n4532 DVDD.n4465 4.5005
R2969 DVDD.n4495 DVDD.n4488 4.5005
R2970 DVDD.n4497 DVDD.n4488 4.5005
R2971 DVDD.n4494 DVDD.n4488 4.5005
R2972 DVDD.n4498 DVDD.n4488 4.5005
R2973 DVDD.n4493 DVDD.n4488 4.5005
R2974 DVDD.n4500 DVDD.n4488 4.5005
R2975 DVDD.n4492 DVDD.n4488 4.5005
R2976 DVDD.n4501 DVDD.n4488 4.5005
R2977 DVDD.n4491 DVDD.n4488 4.5005
R2978 DVDD.n4502 DVDD.n4488 4.5005
R2979 DVDD.n4534 DVDD.n4488 4.5005
R2980 DVDD.n4503 DVDD.n4488 4.5005
R2981 DVDD.n4504 DVDD.n4488 4.5005
R2982 DVDD.n4532 DVDD.n4488 4.5005
R2983 DVDD.n4495 DVDD.n4464 4.5005
R2984 DVDD.n4497 DVDD.n4464 4.5005
R2985 DVDD.n4494 DVDD.n4464 4.5005
R2986 DVDD.n4498 DVDD.n4464 4.5005
R2987 DVDD.n4493 DVDD.n4464 4.5005
R2988 DVDD.n4500 DVDD.n4464 4.5005
R2989 DVDD.n4492 DVDD.n4464 4.5005
R2990 DVDD.n4501 DVDD.n4464 4.5005
R2991 DVDD.n4491 DVDD.n4464 4.5005
R2992 DVDD.n4502 DVDD.n4464 4.5005
R2993 DVDD.n4534 DVDD.n4464 4.5005
R2994 DVDD.n4503 DVDD.n4464 4.5005
R2995 DVDD.n4504 DVDD.n4464 4.5005
R2996 DVDD.n4532 DVDD.n4464 4.5005
R2997 DVDD.n4533 DVDD.n4495 4.5005
R2998 DVDD.n4533 DVDD.n4497 4.5005
R2999 DVDD.n4533 DVDD.n4494 4.5005
R3000 DVDD.n4533 DVDD.n4498 4.5005
R3001 DVDD.n4533 DVDD.n4493 4.5005
R3002 DVDD.n4533 DVDD.n4500 4.5005
R3003 DVDD.n4533 DVDD.n4492 4.5005
R3004 DVDD.n4533 DVDD.n4501 4.5005
R3005 DVDD.n4533 DVDD.n4491 4.5005
R3006 DVDD.n4533 DVDD.n4502 4.5005
R3007 DVDD.n4534 DVDD.n4533 4.5005
R3008 DVDD.n4533 DVDD.n4503 4.5005
R3009 DVDD.n4533 DVDD.n4504 4.5005
R3010 DVDD.n4533 DVDD.n4532 4.5005
R3011 DVDD.n4495 DVDD.n4463 4.5005
R3012 DVDD.n4497 DVDD.n4463 4.5005
R3013 DVDD.n4494 DVDD.n4463 4.5005
R3014 DVDD.n4498 DVDD.n4463 4.5005
R3015 DVDD.n4493 DVDD.n4463 4.5005
R3016 DVDD.n4500 DVDD.n4463 4.5005
R3017 DVDD.n4492 DVDD.n4463 4.5005
R3018 DVDD.n4501 DVDD.n4463 4.5005
R3019 DVDD.n4491 DVDD.n4463 4.5005
R3020 DVDD.n4502 DVDD.n4463 4.5005
R3021 DVDD.n4534 DVDD.n4463 4.5005
R3022 DVDD.n4503 DVDD.n4463 4.5005
R3023 DVDD.n4504 DVDD.n4463 4.5005
R3024 DVDD.n4532 DVDD.n4463 4.5005
R3025 DVDD.n4495 DVDD.n298 4.5005
R3026 DVDD.n4497 DVDD.n298 4.5005
R3027 DVDD.n4494 DVDD.n298 4.5005
R3028 DVDD.n4498 DVDD.n298 4.5005
R3029 DVDD.n4493 DVDD.n298 4.5005
R3030 DVDD.n4500 DVDD.n298 4.5005
R3031 DVDD.n4492 DVDD.n298 4.5005
R3032 DVDD.n4501 DVDD.n298 4.5005
R3033 DVDD.n4491 DVDD.n298 4.5005
R3034 DVDD.n4502 DVDD.n298 4.5005
R3035 DVDD.n4534 DVDD.n298 4.5005
R3036 DVDD.n4503 DVDD.n298 4.5005
R3037 DVDD.n4528 DVDD.n298 4.5005
R3038 DVDD.n4504 DVDD.n298 4.5005
R3039 DVDD.n4532 DVDD.n298 4.5005
R3040 DVDD.n22160 DVDD.n22159 4.5005
R3041 DVDD.n22159 DVDD.n299 4.5005
R3042 DVDD.n22159 DVDD.n297 4.5005
R3043 DVDD.n22159 DVDD.n300 4.5005
R3044 DVDD.n22159 DVDD.n295 4.5005
R3045 DVDD.n22159 DVDD.n301 4.5005
R3046 DVDD.n22159 DVDD.n294 4.5005
R3047 DVDD.n22159 DVDD.n302 4.5005
R3048 DVDD.n22159 DVDD.n293 4.5005
R3049 DVDD.n22159 DVDD.n303 4.5005
R3050 DVDD.n22159 DVDD.n22158 4.5005
R3051 DVDD.n309 DVDD.n299 4.5005
R3052 DVDD.n309 DVDD.n297 4.5005
R3053 DVDD.n323 DVDD.n309 4.5005
R3054 DVDD.n322 DVDD.n309 4.5005
R3055 DVDD.n309 DVDD.n300 4.5005
R3056 DVDD.n309 DVDD.n295 4.5005
R3057 DVDD.n309 DVDD.n301 4.5005
R3058 DVDD.n309 DVDD.n294 4.5005
R3059 DVDD.n309 DVDD.n302 4.5005
R3060 DVDD.n309 DVDD.n293 4.5005
R3061 DVDD.n22156 DVDD.n309 4.5005
R3062 DVDD.n321 DVDD.n309 4.5005
R3063 DVDD.n309 DVDD.n303 4.5005
R3064 DVDD.n22158 DVDD.n309 4.5005
R3065 DVDD.n311 DVDD.n299 4.5005
R3066 DVDD.n311 DVDD.n297 4.5005
R3067 DVDD.n323 DVDD.n311 4.5005
R3068 DVDD.n322 DVDD.n311 4.5005
R3069 DVDD.n311 DVDD.n300 4.5005
R3070 DVDD.n311 DVDD.n295 4.5005
R3071 DVDD.n311 DVDD.n301 4.5005
R3072 DVDD.n311 DVDD.n294 4.5005
R3073 DVDD.n311 DVDD.n302 4.5005
R3074 DVDD.n311 DVDD.n293 4.5005
R3075 DVDD.n22156 DVDD.n311 4.5005
R3076 DVDD.n321 DVDD.n311 4.5005
R3077 DVDD.n311 DVDD.n303 4.5005
R3078 DVDD.n22158 DVDD.n311 4.5005
R3079 DVDD.n308 DVDD.n299 4.5005
R3080 DVDD.n308 DVDD.n297 4.5005
R3081 DVDD.n323 DVDD.n308 4.5005
R3082 DVDD.n322 DVDD.n308 4.5005
R3083 DVDD.n308 DVDD.n300 4.5005
R3084 DVDD.n308 DVDD.n295 4.5005
R3085 DVDD.n308 DVDD.n301 4.5005
R3086 DVDD.n308 DVDD.n294 4.5005
R3087 DVDD.n308 DVDD.n302 4.5005
R3088 DVDD.n308 DVDD.n293 4.5005
R3089 DVDD.n22156 DVDD.n308 4.5005
R3090 DVDD.n321 DVDD.n308 4.5005
R3091 DVDD.n308 DVDD.n303 4.5005
R3092 DVDD.n22158 DVDD.n308 4.5005
R3093 DVDD.n312 DVDD.n299 4.5005
R3094 DVDD.n312 DVDD.n297 4.5005
R3095 DVDD.n323 DVDD.n312 4.5005
R3096 DVDD.n322 DVDD.n312 4.5005
R3097 DVDD.n312 DVDD.n300 4.5005
R3098 DVDD.n312 DVDD.n295 4.5005
R3099 DVDD.n312 DVDD.n301 4.5005
R3100 DVDD.n312 DVDD.n294 4.5005
R3101 DVDD.n312 DVDD.n302 4.5005
R3102 DVDD.n312 DVDD.n293 4.5005
R3103 DVDD.n22156 DVDD.n312 4.5005
R3104 DVDD.n321 DVDD.n312 4.5005
R3105 DVDD.n312 DVDD.n303 4.5005
R3106 DVDD.n22158 DVDD.n312 4.5005
R3107 DVDD.n307 DVDD.n299 4.5005
R3108 DVDD.n307 DVDD.n297 4.5005
R3109 DVDD.n323 DVDD.n307 4.5005
R3110 DVDD.n322 DVDD.n307 4.5005
R3111 DVDD.n307 DVDD.n300 4.5005
R3112 DVDD.n307 DVDD.n295 4.5005
R3113 DVDD.n307 DVDD.n301 4.5005
R3114 DVDD.n307 DVDD.n294 4.5005
R3115 DVDD.n307 DVDD.n302 4.5005
R3116 DVDD.n307 DVDD.n293 4.5005
R3117 DVDD.n22156 DVDD.n307 4.5005
R3118 DVDD.n321 DVDD.n307 4.5005
R3119 DVDD.n307 DVDD.n303 4.5005
R3120 DVDD.n22158 DVDD.n307 4.5005
R3121 DVDD.n313 DVDD.n299 4.5005
R3122 DVDD.n313 DVDD.n297 4.5005
R3123 DVDD.n323 DVDD.n313 4.5005
R3124 DVDD.n322 DVDD.n313 4.5005
R3125 DVDD.n313 DVDD.n300 4.5005
R3126 DVDD.n313 DVDD.n295 4.5005
R3127 DVDD.n313 DVDD.n301 4.5005
R3128 DVDD.n313 DVDD.n294 4.5005
R3129 DVDD.n313 DVDD.n302 4.5005
R3130 DVDD.n313 DVDD.n293 4.5005
R3131 DVDD.n22156 DVDD.n313 4.5005
R3132 DVDD.n321 DVDD.n313 4.5005
R3133 DVDD.n313 DVDD.n303 4.5005
R3134 DVDD.n22158 DVDD.n313 4.5005
R3135 DVDD.n306 DVDD.n299 4.5005
R3136 DVDD.n306 DVDD.n297 4.5005
R3137 DVDD.n323 DVDD.n306 4.5005
R3138 DVDD.n322 DVDD.n306 4.5005
R3139 DVDD.n306 DVDD.n300 4.5005
R3140 DVDD.n306 DVDD.n295 4.5005
R3141 DVDD.n306 DVDD.n301 4.5005
R3142 DVDD.n306 DVDD.n294 4.5005
R3143 DVDD.n306 DVDD.n302 4.5005
R3144 DVDD.n306 DVDD.n293 4.5005
R3145 DVDD.n22156 DVDD.n306 4.5005
R3146 DVDD.n321 DVDD.n306 4.5005
R3147 DVDD.n306 DVDD.n303 4.5005
R3148 DVDD.n22158 DVDD.n306 4.5005
R3149 DVDD.n314 DVDD.n299 4.5005
R3150 DVDD.n314 DVDD.n297 4.5005
R3151 DVDD.n323 DVDD.n314 4.5005
R3152 DVDD.n322 DVDD.n314 4.5005
R3153 DVDD.n314 DVDD.n300 4.5005
R3154 DVDD.n314 DVDD.n295 4.5005
R3155 DVDD.n314 DVDD.n301 4.5005
R3156 DVDD.n314 DVDD.n294 4.5005
R3157 DVDD.n314 DVDD.n302 4.5005
R3158 DVDD.n314 DVDD.n293 4.5005
R3159 DVDD.n22156 DVDD.n314 4.5005
R3160 DVDD.n321 DVDD.n314 4.5005
R3161 DVDD.n314 DVDD.n303 4.5005
R3162 DVDD.n22158 DVDD.n314 4.5005
R3163 DVDD.n305 DVDD.n299 4.5005
R3164 DVDD.n305 DVDD.n297 4.5005
R3165 DVDD.n323 DVDD.n305 4.5005
R3166 DVDD.n322 DVDD.n305 4.5005
R3167 DVDD.n305 DVDD.n300 4.5005
R3168 DVDD.n305 DVDD.n295 4.5005
R3169 DVDD.n305 DVDD.n301 4.5005
R3170 DVDD.n305 DVDD.n294 4.5005
R3171 DVDD.n305 DVDD.n302 4.5005
R3172 DVDD.n305 DVDD.n293 4.5005
R3173 DVDD.n22156 DVDD.n305 4.5005
R3174 DVDD.n321 DVDD.n305 4.5005
R3175 DVDD.n305 DVDD.n303 4.5005
R3176 DVDD.n22158 DVDD.n305 4.5005
R3177 DVDD.n22157 DVDD.n299 4.5005
R3178 DVDD.n22157 DVDD.n297 4.5005
R3179 DVDD.n22157 DVDD.n323 4.5005
R3180 DVDD.n22157 DVDD.n322 4.5005
R3181 DVDD.n22157 DVDD.n300 4.5005
R3182 DVDD.n22157 DVDD.n295 4.5005
R3183 DVDD.n22157 DVDD.n301 4.5005
R3184 DVDD.n22157 DVDD.n294 4.5005
R3185 DVDD.n22157 DVDD.n302 4.5005
R3186 DVDD.n22157 DVDD.n293 4.5005
R3187 DVDD.n22157 DVDD.n22156 4.5005
R3188 DVDD.n22157 DVDD.n321 4.5005
R3189 DVDD.n22157 DVDD.n303 4.5005
R3190 DVDD.n22157 DVDD.n320 4.5005
R3191 DVDD.n22158 DVDD.n22157 4.5005
R3192 DVDD.n19045 DVDD.n19028 4.5005
R3193 DVDD.n19046 DVDD.n19028 4.5005
R3194 DVDD.n19040 DVDD.n19028 4.5005
R3195 DVDD.n19049 DVDD.n19028 4.5005
R3196 DVDD.n19038 DVDD.n19028 4.5005
R3197 DVDD.n19050 DVDD.n19028 4.5005
R3198 DVDD.n19037 DVDD.n19028 4.5005
R3199 DVDD.n19051 DVDD.n19028 4.5005
R3200 DVDD.n19036 DVDD.n19028 4.5005
R3201 DVDD.n20777 DVDD.n19028 4.5005
R3202 DVDD.n19057 DVDD.n19028 4.5005
R3203 DVDD.n20779 DVDD.n19028 4.5005
R3204 DVDD.n19046 DVDD.n19027 4.5005
R3205 DVDD.n19040 DVDD.n19027 4.5005
R3206 DVDD.n19048 DVDD.n19027 4.5005
R3207 DVDD.n19039 DVDD.n19027 4.5005
R3208 DVDD.n19049 DVDD.n19027 4.5005
R3209 DVDD.n19038 DVDD.n19027 4.5005
R3210 DVDD.n19050 DVDD.n19027 4.5005
R3211 DVDD.n19037 DVDD.n19027 4.5005
R3212 DVDD.n19051 DVDD.n19027 4.5005
R3213 DVDD.n19036 DVDD.n19027 4.5005
R3214 DVDD.n19053 DVDD.n19027 4.5005
R3215 DVDD.n19035 DVDD.n19027 4.5005
R3216 DVDD.n20777 DVDD.n19027 4.5005
R3217 DVDD.n19057 DVDD.n19027 4.5005
R3218 DVDD.n20779 DVDD.n19027 4.5005
R3219 DVDD.n19046 DVDD.n19029 4.5005
R3220 DVDD.n19040 DVDD.n19029 4.5005
R3221 DVDD.n19048 DVDD.n19029 4.5005
R3222 DVDD.n19039 DVDD.n19029 4.5005
R3223 DVDD.n19049 DVDD.n19029 4.5005
R3224 DVDD.n19038 DVDD.n19029 4.5005
R3225 DVDD.n19050 DVDD.n19029 4.5005
R3226 DVDD.n19037 DVDD.n19029 4.5005
R3227 DVDD.n19051 DVDD.n19029 4.5005
R3228 DVDD.n19036 DVDD.n19029 4.5005
R3229 DVDD.n19053 DVDD.n19029 4.5005
R3230 DVDD.n19035 DVDD.n19029 4.5005
R3231 DVDD.n20777 DVDD.n19029 4.5005
R3232 DVDD.n20779 DVDD.n19029 4.5005
R3233 DVDD.n19046 DVDD.n19026 4.5005
R3234 DVDD.n19040 DVDD.n19026 4.5005
R3235 DVDD.n19048 DVDD.n19026 4.5005
R3236 DVDD.n19039 DVDD.n19026 4.5005
R3237 DVDD.n19049 DVDD.n19026 4.5005
R3238 DVDD.n19038 DVDD.n19026 4.5005
R3239 DVDD.n19050 DVDD.n19026 4.5005
R3240 DVDD.n19037 DVDD.n19026 4.5005
R3241 DVDD.n19051 DVDD.n19026 4.5005
R3242 DVDD.n19036 DVDD.n19026 4.5005
R3243 DVDD.n19053 DVDD.n19026 4.5005
R3244 DVDD.n19035 DVDD.n19026 4.5005
R3245 DVDD.n20777 DVDD.n19026 4.5005
R3246 DVDD.n20779 DVDD.n19026 4.5005
R3247 DVDD.n19046 DVDD.n19030 4.5005
R3248 DVDD.n19040 DVDD.n19030 4.5005
R3249 DVDD.n19048 DVDD.n19030 4.5005
R3250 DVDD.n19039 DVDD.n19030 4.5005
R3251 DVDD.n19049 DVDD.n19030 4.5005
R3252 DVDD.n19038 DVDD.n19030 4.5005
R3253 DVDD.n19050 DVDD.n19030 4.5005
R3254 DVDD.n19037 DVDD.n19030 4.5005
R3255 DVDD.n19051 DVDD.n19030 4.5005
R3256 DVDD.n19036 DVDD.n19030 4.5005
R3257 DVDD.n19053 DVDD.n19030 4.5005
R3258 DVDD.n19035 DVDD.n19030 4.5005
R3259 DVDD.n20777 DVDD.n19030 4.5005
R3260 DVDD.n20779 DVDD.n19030 4.5005
R3261 DVDD.n19046 DVDD.n19025 4.5005
R3262 DVDD.n19040 DVDD.n19025 4.5005
R3263 DVDD.n19048 DVDD.n19025 4.5005
R3264 DVDD.n19039 DVDD.n19025 4.5005
R3265 DVDD.n19049 DVDD.n19025 4.5005
R3266 DVDD.n19038 DVDD.n19025 4.5005
R3267 DVDD.n19050 DVDD.n19025 4.5005
R3268 DVDD.n19037 DVDD.n19025 4.5005
R3269 DVDD.n19051 DVDD.n19025 4.5005
R3270 DVDD.n19036 DVDD.n19025 4.5005
R3271 DVDD.n19053 DVDD.n19025 4.5005
R3272 DVDD.n19035 DVDD.n19025 4.5005
R3273 DVDD.n20777 DVDD.n19025 4.5005
R3274 DVDD.n20779 DVDD.n19025 4.5005
R3275 DVDD.n19046 DVDD.n19031 4.5005
R3276 DVDD.n19040 DVDD.n19031 4.5005
R3277 DVDD.n19048 DVDD.n19031 4.5005
R3278 DVDD.n19039 DVDD.n19031 4.5005
R3279 DVDD.n19049 DVDD.n19031 4.5005
R3280 DVDD.n19038 DVDD.n19031 4.5005
R3281 DVDD.n19050 DVDD.n19031 4.5005
R3282 DVDD.n19037 DVDD.n19031 4.5005
R3283 DVDD.n19051 DVDD.n19031 4.5005
R3284 DVDD.n19036 DVDD.n19031 4.5005
R3285 DVDD.n19053 DVDD.n19031 4.5005
R3286 DVDD.n19035 DVDD.n19031 4.5005
R3287 DVDD.n20777 DVDD.n19031 4.5005
R3288 DVDD.n19057 DVDD.n19031 4.5005
R3289 DVDD.n20779 DVDD.n19031 4.5005
R3290 DVDD.n20779 DVDD.n19024 4.5005
R3291 DVDD.n20779 DVDD.n19032 4.5005
R3292 DVDD.n19046 DVDD.n19023 4.5005
R3293 DVDD.n19040 DVDD.n19023 4.5005
R3294 DVDD.n19048 DVDD.n19023 4.5005
R3295 DVDD.n19039 DVDD.n19023 4.5005
R3296 DVDD.n19049 DVDD.n19023 4.5005
R3297 DVDD.n19038 DVDD.n19023 4.5005
R3298 DVDD.n19050 DVDD.n19023 4.5005
R3299 DVDD.n19037 DVDD.n19023 4.5005
R3300 DVDD.n19051 DVDD.n19023 4.5005
R3301 DVDD.n19036 DVDD.n19023 4.5005
R3302 DVDD.n19053 DVDD.n19023 4.5005
R3303 DVDD.n19035 DVDD.n19023 4.5005
R3304 DVDD.n20777 DVDD.n19023 4.5005
R3305 DVDD.n20779 DVDD.n19023 4.5005
R3306 DVDD.n20778 DVDD.n19045 4.5005
R3307 DVDD.n20778 DVDD.n19046 4.5005
R3308 DVDD.n20778 DVDD.n19040 4.5005
R3309 DVDD.n20778 DVDD.n19048 4.5005
R3310 DVDD.n20778 DVDD.n19039 4.5005
R3311 DVDD.n20778 DVDD.n19049 4.5005
R3312 DVDD.n20778 DVDD.n19038 4.5005
R3313 DVDD.n20778 DVDD.n19050 4.5005
R3314 DVDD.n20778 DVDD.n19037 4.5005
R3315 DVDD.n20778 DVDD.n19051 4.5005
R3316 DVDD.n20778 DVDD.n19036 4.5005
R3317 DVDD.n20778 DVDD.n19053 4.5005
R3318 DVDD.n20778 DVDD.n19035 4.5005
R3319 DVDD.n20778 DVDD.n20777 4.5005
R3320 DVDD.n20779 DVDD.n20778 4.5005
R3321 DVDD.n19891 DVDD.n19879 4.5005
R3322 DVDD.n19936 DVDD.n19879 4.5005
R3323 DVDD.n19890 DVDD.n19879 4.5005
R3324 DVDD.n19939 DVDD.n19879 4.5005
R3325 DVDD.n19888 DVDD.n19879 4.5005
R3326 DVDD.n19940 DVDD.n19879 4.5005
R3327 DVDD.n19887 DVDD.n19879 4.5005
R3328 DVDD.n19941 DVDD.n19879 4.5005
R3329 DVDD.n19886 DVDD.n19879 4.5005
R3330 DVDD.n20283 DVDD.n19879 4.5005
R3331 DVDD.n19879 DVDD.n19873 4.5005
R3332 DVDD.n20285 DVDD.n19879 4.5005
R3333 DVDD.n19891 DVDD.n19878 4.5005
R3334 DVDD.n19936 DVDD.n19878 4.5005
R3335 DVDD.n19890 DVDD.n19878 4.5005
R3336 DVDD.n19938 DVDD.n19878 4.5005
R3337 DVDD.n19889 DVDD.n19878 4.5005
R3338 DVDD.n19939 DVDD.n19878 4.5005
R3339 DVDD.n19888 DVDD.n19878 4.5005
R3340 DVDD.n19940 DVDD.n19878 4.5005
R3341 DVDD.n19887 DVDD.n19878 4.5005
R3342 DVDD.n19941 DVDD.n19878 4.5005
R3343 DVDD.n19886 DVDD.n19878 4.5005
R3344 DVDD.n19943 DVDD.n19878 4.5005
R3345 DVDD.n19885 DVDD.n19878 4.5005
R3346 DVDD.n20283 DVDD.n19878 4.5005
R3347 DVDD.n19878 DVDD.n19873 4.5005
R3348 DVDD.n20285 DVDD.n19878 4.5005
R3349 DVDD.n19891 DVDD.n19880 4.5005
R3350 DVDD.n19936 DVDD.n19880 4.5005
R3351 DVDD.n19890 DVDD.n19880 4.5005
R3352 DVDD.n19938 DVDD.n19880 4.5005
R3353 DVDD.n19889 DVDD.n19880 4.5005
R3354 DVDD.n19939 DVDD.n19880 4.5005
R3355 DVDD.n19888 DVDD.n19880 4.5005
R3356 DVDD.n19940 DVDD.n19880 4.5005
R3357 DVDD.n19887 DVDD.n19880 4.5005
R3358 DVDD.n19941 DVDD.n19880 4.5005
R3359 DVDD.n19886 DVDD.n19880 4.5005
R3360 DVDD.n19943 DVDD.n19880 4.5005
R3361 DVDD.n19885 DVDD.n19880 4.5005
R3362 DVDD.n20283 DVDD.n19880 4.5005
R3363 DVDD.n19880 DVDD.n19873 4.5005
R3364 DVDD.n20285 DVDD.n19880 4.5005
R3365 DVDD.n19891 DVDD.n19877 4.5005
R3366 DVDD.n19936 DVDD.n19877 4.5005
R3367 DVDD.n19890 DVDD.n19877 4.5005
R3368 DVDD.n19938 DVDD.n19877 4.5005
R3369 DVDD.n19889 DVDD.n19877 4.5005
R3370 DVDD.n19939 DVDD.n19877 4.5005
R3371 DVDD.n19888 DVDD.n19877 4.5005
R3372 DVDD.n19940 DVDD.n19877 4.5005
R3373 DVDD.n19887 DVDD.n19877 4.5005
R3374 DVDD.n19941 DVDD.n19877 4.5005
R3375 DVDD.n19886 DVDD.n19877 4.5005
R3376 DVDD.n19943 DVDD.n19877 4.5005
R3377 DVDD.n19885 DVDD.n19877 4.5005
R3378 DVDD.n20283 DVDD.n19877 4.5005
R3379 DVDD.n19877 DVDD.n19873 4.5005
R3380 DVDD.n20285 DVDD.n19877 4.5005
R3381 DVDD.n19891 DVDD.n19881 4.5005
R3382 DVDD.n19936 DVDD.n19881 4.5005
R3383 DVDD.n19890 DVDD.n19881 4.5005
R3384 DVDD.n19938 DVDD.n19881 4.5005
R3385 DVDD.n19889 DVDD.n19881 4.5005
R3386 DVDD.n19939 DVDD.n19881 4.5005
R3387 DVDD.n19888 DVDD.n19881 4.5005
R3388 DVDD.n19940 DVDD.n19881 4.5005
R3389 DVDD.n19887 DVDD.n19881 4.5005
R3390 DVDD.n19941 DVDD.n19881 4.5005
R3391 DVDD.n19886 DVDD.n19881 4.5005
R3392 DVDD.n19943 DVDD.n19881 4.5005
R3393 DVDD.n19885 DVDD.n19881 4.5005
R3394 DVDD.n20283 DVDD.n19881 4.5005
R3395 DVDD.n19881 DVDD.n19873 4.5005
R3396 DVDD.n20285 DVDD.n19881 4.5005
R3397 DVDD.n19891 DVDD.n19876 4.5005
R3398 DVDD.n19936 DVDD.n19876 4.5005
R3399 DVDD.n19890 DVDD.n19876 4.5005
R3400 DVDD.n19938 DVDD.n19876 4.5005
R3401 DVDD.n19889 DVDD.n19876 4.5005
R3402 DVDD.n19939 DVDD.n19876 4.5005
R3403 DVDD.n19888 DVDD.n19876 4.5005
R3404 DVDD.n19940 DVDD.n19876 4.5005
R3405 DVDD.n19887 DVDD.n19876 4.5005
R3406 DVDD.n19941 DVDD.n19876 4.5005
R3407 DVDD.n19886 DVDD.n19876 4.5005
R3408 DVDD.n19943 DVDD.n19876 4.5005
R3409 DVDD.n19885 DVDD.n19876 4.5005
R3410 DVDD.n20283 DVDD.n19876 4.5005
R3411 DVDD.n19876 DVDD.n19873 4.5005
R3412 DVDD.n20285 DVDD.n19876 4.5005
R3413 DVDD.n19891 DVDD.n19882 4.5005
R3414 DVDD.n19936 DVDD.n19882 4.5005
R3415 DVDD.n19890 DVDD.n19882 4.5005
R3416 DVDD.n19938 DVDD.n19882 4.5005
R3417 DVDD.n19889 DVDD.n19882 4.5005
R3418 DVDD.n19939 DVDD.n19882 4.5005
R3419 DVDD.n19888 DVDD.n19882 4.5005
R3420 DVDD.n19940 DVDD.n19882 4.5005
R3421 DVDD.n19887 DVDD.n19882 4.5005
R3422 DVDD.n19941 DVDD.n19882 4.5005
R3423 DVDD.n19886 DVDD.n19882 4.5005
R3424 DVDD.n19943 DVDD.n19882 4.5005
R3425 DVDD.n19885 DVDD.n19882 4.5005
R3426 DVDD.n20283 DVDD.n19882 4.5005
R3427 DVDD.n19882 DVDD.n19873 4.5005
R3428 DVDD.n20285 DVDD.n19882 4.5005
R3429 DVDD.n19891 DVDD.n19875 4.5005
R3430 DVDD.n19936 DVDD.n19875 4.5005
R3431 DVDD.n19890 DVDD.n19875 4.5005
R3432 DVDD.n19938 DVDD.n19875 4.5005
R3433 DVDD.n19889 DVDD.n19875 4.5005
R3434 DVDD.n19939 DVDD.n19875 4.5005
R3435 DVDD.n19888 DVDD.n19875 4.5005
R3436 DVDD.n19940 DVDD.n19875 4.5005
R3437 DVDD.n19887 DVDD.n19875 4.5005
R3438 DVDD.n19941 DVDD.n19875 4.5005
R3439 DVDD.n19886 DVDD.n19875 4.5005
R3440 DVDD.n19943 DVDD.n19875 4.5005
R3441 DVDD.n19885 DVDD.n19875 4.5005
R3442 DVDD.n20283 DVDD.n19875 4.5005
R3443 DVDD.n19875 DVDD.n19873 4.5005
R3444 DVDD.n20285 DVDD.n19875 4.5005
R3445 DVDD.n19891 DVDD.n19883 4.5005
R3446 DVDD.n19936 DVDD.n19883 4.5005
R3447 DVDD.n19890 DVDD.n19883 4.5005
R3448 DVDD.n19938 DVDD.n19883 4.5005
R3449 DVDD.n19889 DVDD.n19883 4.5005
R3450 DVDD.n19939 DVDD.n19883 4.5005
R3451 DVDD.n19888 DVDD.n19883 4.5005
R3452 DVDD.n19940 DVDD.n19883 4.5005
R3453 DVDD.n19887 DVDD.n19883 4.5005
R3454 DVDD.n19941 DVDD.n19883 4.5005
R3455 DVDD.n19886 DVDD.n19883 4.5005
R3456 DVDD.n19943 DVDD.n19883 4.5005
R3457 DVDD.n19885 DVDD.n19883 4.5005
R3458 DVDD.n20283 DVDD.n19883 4.5005
R3459 DVDD.n19883 DVDD.n19873 4.5005
R3460 DVDD.n20285 DVDD.n19883 4.5005
R3461 DVDD.n19891 DVDD.n19874 4.5005
R3462 DVDD.n19936 DVDD.n19874 4.5005
R3463 DVDD.n19890 DVDD.n19874 4.5005
R3464 DVDD.n19938 DVDD.n19874 4.5005
R3465 DVDD.n19889 DVDD.n19874 4.5005
R3466 DVDD.n19939 DVDD.n19874 4.5005
R3467 DVDD.n19888 DVDD.n19874 4.5005
R3468 DVDD.n19940 DVDD.n19874 4.5005
R3469 DVDD.n19887 DVDD.n19874 4.5005
R3470 DVDD.n19941 DVDD.n19874 4.5005
R3471 DVDD.n19886 DVDD.n19874 4.5005
R3472 DVDD.n19943 DVDD.n19874 4.5005
R3473 DVDD.n19885 DVDD.n19874 4.5005
R3474 DVDD.n20283 DVDD.n19874 4.5005
R3475 DVDD.n19874 DVDD.n19873 4.5005
R3476 DVDD.n20285 DVDD.n19874 4.5005
R3477 DVDD.n20284 DVDD.n19891 4.5005
R3478 DVDD.n20284 DVDD.n19936 4.5005
R3479 DVDD.n20284 DVDD.n19890 4.5005
R3480 DVDD.n20284 DVDD.n19938 4.5005
R3481 DVDD.n20284 DVDD.n19889 4.5005
R3482 DVDD.n20284 DVDD.n19939 4.5005
R3483 DVDD.n20284 DVDD.n19888 4.5005
R3484 DVDD.n20284 DVDD.n19940 4.5005
R3485 DVDD.n20284 DVDD.n19887 4.5005
R3486 DVDD.n20284 DVDD.n19941 4.5005
R3487 DVDD.n20284 DVDD.n19886 4.5005
R3488 DVDD.n20284 DVDD.n19943 4.5005
R3489 DVDD.n20284 DVDD.n19885 4.5005
R3490 DVDD.n20284 DVDD.n20283 4.5005
R3491 DVDD.n20284 DVDD.n19873 4.5005
R3492 DVDD.n20285 DVDD.n20284 4.5005
R3493 DVDD.n19057 DVDD.n19032 4.5005
R3494 DVDD.n20777 DVDD.n19032 4.5005
R3495 DVDD.n19035 DVDD.n19032 4.5005
R3496 DVDD.n19053 DVDD.n19032 4.5005
R3497 DVDD.n19036 DVDD.n19032 4.5005
R3498 DVDD.n19051 DVDD.n19032 4.5005
R3499 DVDD.n19037 DVDD.n19032 4.5005
R3500 DVDD.n19050 DVDD.n19032 4.5005
R3501 DVDD.n19038 DVDD.n19032 4.5005
R3502 DVDD.n19049 DVDD.n19032 4.5005
R3503 DVDD.n19039 DVDD.n19032 4.5005
R3504 DVDD.n19048 DVDD.n19032 4.5005
R3505 DVDD.n19040 DVDD.n19032 4.5005
R3506 DVDD.n19046 DVDD.n19032 4.5005
R3507 DVDD.n19057 DVDD.n19024 4.5005
R3508 DVDD.n20777 DVDD.n19024 4.5005
R3509 DVDD.n19035 DVDD.n19024 4.5005
R3510 DVDD.n19053 DVDD.n19024 4.5005
R3511 DVDD.n19036 DVDD.n19024 4.5005
R3512 DVDD.n19051 DVDD.n19024 4.5005
R3513 DVDD.n19037 DVDD.n19024 4.5005
R3514 DVDD.n19050 DVDD.n19024 4.5005
R3515 DVDD.n19038 DVDD.n19024 4.5005
R3516 DVDD.n19049 DVDD.n19024 4.5005
R3517 DVDD.n19039 DVDD.n19024 4.5005
R3518 DVDD.n19048 DVDD.n19024 4.5005
R3519 DVDD.n19040 DVDD.n19024 4.5005
R3520 DVDD.n19046 DVDD.n19024 4.5005
R3521 DVDD.n19045 DVDD.n19024 4.5005
R3522 DVDD.n4557 DVDD.n4401 4.5005
R3523 DVDD.n4557 DVDD.n4394 4.5005
R3524 DVDD.n4401 DVDD.n4324 4.5005
R3525 DVDD.n4394 DVDD.n4324 4.5005
R3526 DVDD.n4534 DVDD.n4324 4.5005
R3527 DVDD.n4401 DVDD.n4387 4.5005
R3528 DVDD.n4394 DVDD.n4387 4.5005
R3529 DVDD.n4534 DVDD.n4387 4.5005
R3530 DVDD.n4401 DVDD.n4325 4.5005
R3531 DVDD.n4394 DVDD.n4325 4.5005
R3532 DVDD.n4534 DVDD.n4325 4.5005
R3533 DVDD.n4401 DVDD.n4386 4.5005
R3534 DVDD.n4394 DVDD.n4386 4.5005
R3535 DVDD.n4534 DVDD.n4386 4.5005
R3536 DVDD.n4401 DVDD.n4326 4.5005
R3537 DVDD.n4394 DVDD.n4326 4.5005
R3538 DVDD.n4534 DVDD.n4326 4.5005
R3539 DVDD.n4401 DVDD.n4332 4.5005
R3540 DVDD.n4394 DVDD.n4332 4.5005
R3541 DVDD.n4534 DVDD.n4332 4.5005
R3542 DVDD.n4401 DVDD.n4327 4.5005
R3543 DVDD.n4394 DVDD.n4327 4.5005
R3544 DVDD.n4534 DVDD.n4327 4.5005
R3545 DVDD.n4401 DVDD.n4331 4.5005
R3546 DVDD.n4394 DVDD.n4331 4.5005
R3547 DVDD.n4534 DVDD.n4331 4.5005
R3548 DVDD.n4393 DVDD.n4331 4.5005
R3549 DVDD.n4393 DVDD.n4327 4.5005
R3550 DVDD.n4393 DVDD.n4332 4.5005
R3551 DVDD.n4393 DVDD.n4326 4.5005
R3552 DVDD.n4393 DVDD.n4386 4.5005
R3553 DVDD.n4393 DVDD.n4325 4.5005
R3554 DVDD.n4393 DVDD.n4387 4.5005
R3555 DVDD.n4393 DVDD.n4324 4.5005
R3556 DVDD.n4557 DVDD.n4393 4.5005
R3557 DVDD.n4557 DVDD.n4402 4.5005
R3558 DVDD.n4557 DVDD.n4392 4.5005
R3559 DVDD.n4557 DVDD.n4403 4.5005
R3560 DVDD.n4402 DVDD.n4324 4.5005
R3561 DVDD.n4392 DVDD.n4324 4.5005
R3562 DVDD.n4403 DVDD.n4324 4.5005
R3563 DVDD.n4402 DVDD.n4387 4.5005
R3564 DVDD.n4392 DVDD.n4387 4.5005
R3565 DVDD.n4403 DVDD.n4387 4.5005
R3566 DVDD.n4402 DVDD.n4325 4.5005
R3567 DVDD.n4392 DVDD.n4325 4.5005
R3568 DVDD.n4403 DVDD.n4325 4.5005
R3569 DVDD.n4402 DVDD.n4386 4.5005
R3570 DVDD.n4392 DVDD.n4386 4.5005
R3571 DVDD.n4403 DVDD.n4386 4.5005
R3572 DVDD.n4402 DVDD.n4326 4.5005
R3573 DVDD.n4392 DVDD.n4326 4.5005
R3574 DVDD.n4403 DVDD.n4326 4.5005
R3575 DVDD.n4402 DVDD.n4332 4.5005
R3576 DVDD.n4392 DVDD.n4332 4.5005
R3577 DVDD.n4403 DVDD.n4332 4.5005
R3578 DVDD.n4402 DVDD.n4327 4.5005
R3579 DVDD.n4392 DVDD.n4327 4.5005
R3580 DVDD.n4403 DVDD.n4327 4.5005
R3581 DVDD.n4402 DVDD.n4331 4.5005
R3582 DVDD.n4392 DVDD.n4331 4.5005
R3583 DVDD.n4403 DVDD.n4331 4.5005
R3584 DVDD.n4391 DVDD.n4331 4.5005
R3585 DVDD.n4391 DVDD.n4327 4.5005
R3586 DVDD.n4391 DVDD.n4332 4.5005
R3587 DVDD.n4391 DVDD.n4326 4.5005
R3588 DVDD.n4391 DVDD.n4386 4.5005
R3589 DVDD.n4391 DVDD.n4325 4.5005
R3590 DVDD.n4391 DVDD.n4387 4.5005
R3591 DVDD.n4391 DVDD.n4324 4.5005
R3592 DVDD.n4557 DVDD.n4391 4.5005
R3593 DVDD.n4557 DVDD.n4405 4.5005
R3594 DVDD.n4557 DVDD.n4390 4.5005
R3595 DVDD.n4557 DVDD.n4406 4.5005
R3596 DVDD.n4405 DVDD.n4324 4.5005
R3597 DVDD.n4390 DVDD.n4324 4.5005
R3598 DVDD.n4406 DVDD.n4324 4.5005
R3599 DVDD.n4405 DVDD.n4387 4.5005
R3600 DVDD.n4390 DVDD.n4387 4.5005
R3601 DVDD.n4406 DVDD.n4387 4.5005
R3602 DVDD.n4405 DVDD.n4325 4.5005
R3603 DVDD.n4390 DVDD.n4325 4.5005
R3604 DVDD.n4406 DVDD.n4325 4.5005
R3605 DVDD.n4405 DVDD.n4386 4.5005
R3606 DVDD.n4390 DVDD.n4386 4.5005
R3607 DVDD.n4406 DVDD.n4386 4.5005
R3608 DVDD.n4405 DVDD.n4326 4.5005
R3609 DVDD.n4390 DVDD.n4326 4.5005
R3610 DVDD.n4406 DVDD.n4326 4.5005
R3611 DVDD.n4405 DVDD.n4332 4.5005
R3612 DVDD.n4390 DVDD.n4332 4.5005
R3613 DVDD.n4406 DVDD.n4332 4.5005
R3614 DVDD.n4405 DVDD.n4327 4.5005
R3615 DVDD.n4390 DVDD.n4327 4.5005
R3616 DVDD.n4406 DVDD.n4327 4.5005
R3617 DVDD.n4405 DVDD.n4331 4.5005
R3618 DVDD.n4390 DVDD.n4331 4.5005
R3619 DVDD.n4406 DVDD.n4331 4.5005
R3620 DVDD.n4389 DVDD.n4331 4.5005
R3621 DVDD.n4389 DVDD.n4327 4.5005
R3622 DVDD.n4389 DVDD.n4332 4.5005
R3623 DVDD.n4389 DVDD.n4326 4.5005
R3624 DVDD.n4389 DVDD.n4386 4.5005
R3625 DVDD.n4389 DVDD.n4325 4.5005
R3626 DVDD.n4389 DVDD.n4387 4.5005
R3627 DVDD.n4389 DVDD.n4324 4.5005
R3628 DVDD.n4557 DVDD.n4389 4.5005
R3629 DVDD.n4555 DVDD.n4386 4.5005
R3630 DVDD.n2341 DVDD.n2296 4.5005
R3631 DVDD.n2342 DVDD.n2296 4.5005
R3632 DVDD.n2340 DVDD.n2296 4.5005
R3633 DVDD.n2343 DVDD.n2296 4.5005
R3634 DVDD.n2339 DVDD.n2296 4.5005
R3635 DVDD.n2344 DVDD.n2296 4.5005
R3636 DVDD.n2338 DVDD.n2296 4.5005
R3637 DVDD.n2345 DVDD.n2296 4.5005
R3638 DVDD.n2337 DVDD.n2296 4.5005
R3639 DVDD.n2346 DVDD.n2296 4.5005
R3640 DVDD.n2336 DVDD.n2296 4.5005
R3641 DVDD.n2347 DVDD.n2296 4.5005
R3642 DVDD.n2348 DVDD.n2296 4.5005
R3643 DVDD.n16390 DVDD.n2296 4.5005
R3644 DVDD.n16394 DVDD.n2296 4.5005
R3645 DVDD.n2341 DVDD.n2306 4.5005
R3646 DVDD.n2342 DVDD.n2306 4.5005
R3647 DVDD.n2340 DVDD.n2306 4.5005
R3648 DVDD.n2343 DVDD.n2306 4.5005
R3649 DVDD.n2339 DVDD.n2306 4.5005
R3650 DVDD.n2344 DVDD.n2306 4.5005
R3651 DVDD.n2338 DVDD.n2306 4.5005
R3652 DVDD.n2345 DVDD.n2306 4.5005
R3653 DVDD.n2337 DVDD.n2306 4.5005
R3654 DVDD.n2346 DVDD.n2306 4.5005
R3655 DVDD.n2336 DVDD.n2306 4.5005
R3656 DVDD.n2347 DVDD.n2306 4.5005
R3657 DVDD.n2335 DVDD.n2306 4.5005
R3658 DVDD.n2348 DVDD.n2306 4.5005
R3659 DVDD.n16390 DVDD.n2306 4.5005
R3660 DVDD.n16394 DVDD.n2306 4.5005
R3661 DVDD.n2341 DVDD.n2325 4.5005
R3662 DVDD.n2342 DVDD.n2325 4.5005
R3663 DVDD.n2340 DVDD.n2325 4.5005
R3664 DVDD.n2343 DVDD.n2325 4.5005
R3665 DVDD.n2339 DVDD.n2325 4.5005
R3666 DVDD.n2344 DVDD.n2325 4.5005
R3667 DVDD.n2338 DVDD.n2325 4.5005
R3668 DVDD.n2345 DVDD.n2325 4.5005
R3669 DVDD.n2337 DVDD.n2325 4.5005
R3670 DVDD.n2346 DVDD.n2325 4.5005
R3671 DVDD.n2336 DVDD.n2325 4.5005
R3672 DVDD.n2347 DVDD.n2325 4.5005
R3673 DVDD.n2335 DVDD.n2325 4.5005
R3674 DVDD.n2348 DVDD.n2325 4.5005
R3675 DVDD.n16390 DVDD.n2325 4.5005
R3676 DVDD.n16394 DVDD.n2325 4.5005
R3677 DVDD.n3033 DVDD.n3024 4.5005
R3678 DVDD.n3031 DVDD.n3024 4.5005
R3679 DVDD.n3035 DVDD.n3024 4.5005
R3680 DVDD.n3030 DVDD.n3024 4.5005
R3681 DVDD.n3036 DVDD.n3024 4.5005
R3682 DVDD.n3029 DVDD.n3024 4.5005
R3683 DVDD.n3037 DVDD.n3024 4.5005
R3684 DVDD.n3028 DVDD.n3024 4.5005
R3685 DVDD.n3038 DVDD.n3024 4.5005
R3686 DVDD.n3027 DVDD.n3024 4.5005
R3687 DVDD.n3040 DVDD.n3024 4.5005
R3688 DVDD.n3026 DVDD.n3024 4.5005
R3689 DVDD.n16142 DVDD.n3024 4.5005
R3690 DVDD.n3024 DVDD.n2995 4.5005
R3691 DVDD.n16144 DVDD.n3024 4.5005
R3692 DVDD.n3033 DVDD.n2996 4.5005
R3693 DVDD.n3031 DVDD.n2996 4.5005
R3694 DVDD.n3035 DVDD.n2996 4.5005
R3695 DVDD.n3030 DVDD.n2996 4.5005
R3696 DVDD.n3036 DVDD.n2996 4.5005
R3697 DVDD.n3029 DVDD.n2996 4.5005
R3698 DVDD.n3037 DVDD.n2996 4.5005
R3699 DVDD.n3028 DVDD.n2996 4.5005
R3700 DVDD.n3038 DVDD.n2996 4.5005
R3701 DVDD.n3027 DVDD.n2996 4.5005
R3702 DVDD.n3040 DVDD.n2996 4.5005
R3703 DVDD.n3026 DVDD.n2996 4.5005
R3704 DVDD.n16142 DVDD.n2996 4.5005
R3705 DVDD.n2996 DVDD.n2995 4.5005
R3706 DVDD.n16144 DVDD.n2996 4.5005
R3707 DVDD.n16143 DVDD.n3033 4.5005
R3708 DVDD.n16143 DVDD.n3031 4.5005
R3709 DVDD.n16143 DVDD.n3035 4.5005
R3710 DVDD.n16143 DVDD.n3030 4.5005
R3711 DVDD.n16143 DVDD.n3036 4.5005
R3712 DVDD.n16143 DVDD.n3029 4.5005
R3713 DVDD.n16143 DVDD.n3037 4.5005
R3714 DVDD.n16143 DVDD.n3028 4.5005
R3715 DVDD.n16143 DVDD.n3038 4.5005
R3716 DVDD.n16143 DVDD.n3027 4.5005
R3717 DVDD.n16143 DVDD.n3040 4.5005
R3718 DVDD.n16143 DVDD.n3026 4.5005
R3719 DVDD.n16143 DVDD.n16142 4.5005
R3720 DVDD.n16143 DVDD.n2995 4.5005
R3721 DVDD.n16144 DVDD.n16143 4.5005
R3722 DVDD.n10068 DVDD.n9676 4.5005
R3723 DVDD.n9686 DVDD.n9676 4.5005
R3724 DVDD.n9689 DVDD.n9676 4.5005
R3725 DVDD.n9685 DVDD.n9676 4.5005
R3726 DVDD.n9690 DVDD.n9676 4.5005
R3727 DVDD.n9684 DVDD.n9676 4.5005
R3728 DVDD.n9691 DVDD.n9676 4.5005
R3729 DVDD.n9683 DVDD.n9676 4.5005
R3730 DVDD.n9692 DVDD.n9676 4.5005
R3731 DVDD.n9682 DVDD.n9676 4.5005
R3732 DVDD.n9694 DVDD.n9676 4.5005
R3733 DVDD.n9681 DVDD.n9676 4.5005
R3734 DVDD.n9695 DVDD.n9676 4.5005
R3735 DVDD.n9680 DVDD.n9676 4.5005
R3736 DVDD.n10066 DVDD.n9676 4.5005
R3737 DVDD.n10068 DVDD.n9662 4.5005
R3738 DVDD.n9686 DVDD.n9662 4.5005
R3739 DVDD.n9689 DVDD.n9662 4.5005
R3740 DVDD.n9685 DVDD.n9662 4.5005
R3741 DVDD.n9690 DVDD.n9662 4.5005
R3742 DVDD.n9684 DVDD.n9662 4.5005
R3743 DVDD.n9691 DVDD.n9662 4.5005
R3744 DVDD.n9683 DVDD.n9662 4.5005
R3745 DVDD.n9692 DVDD.n9662 4.5005
R3746 DVDD.n9682 DVDD.n9662 4.5005
R3747 DVDD.n9694 DVDD.n9662 4.5005
R3748 DVDD.n9681 DVDD.n9662 4.5005
R3749 DVDD.n9695 DVDD.n9662 4.5005
R3750 DVDD.n9680 DVDD.n9662 4.5005
R3751 DVDD.n10066 DVDD.n9662 4.5005
R3752 DVDD.n10068 DVDD.n10067 4.5005
R3753 DVDD.n10067 DVDD.n9686 4.5005
R3754 DVDD.n10067 DVDD.n9689 4.5005
R3755 DVDD.n10067 DVDD.n9685 4.5005
R3756 DVDD.n10067 DVDD.n9690 4.5005
R3757 DVDD.n10067 DVDD.n9684 4.5005
R3758 DVDD.n10067 DVDD.n9691 4.5005
R3759 DVDD.n10067 DVDD.n9683 4.5005
R3760 DVDD.n10067 DVDD.n9692 4.5005
R3761 DVDD.n10067 DVDD.n9682 4.5005
R3762 DVDD.n10067 DVDD.n9694 4.5005
R3763 DVDD.n10067 DVDD.n9681 4.5005
R3764 DVDD.n10067 DVDD.n9695 4.5005
R3765 DVDD.n10067 DVDD.n9680 4.5005
R3766 DVDD.n10067 DVDD.n10066 4.5005
R3767 DVDD.n21049 DVDD.n66 4.5005
R3768 DVDD.n21019 DVDD.n66 4.5005
R3769 DVDD.n21049 DVDD.n21048 4.5005
R3770 DVDD.n21048 DVDD.n21027 4.5005
R3771 DVDD.n21048 DVDD.n21025 4.5005
R3772 DVDD.n21048 DVDD.n21030 4.5005
R3773 DVDD.n21048 DVDD.n21024 4.5005
R3774 DVDD.n21048 DVDD.n21033 4.5005
R3775 DVDD.n21048 DVDD.n21023 4.5005
R3776 DVDD.n21048 DVDD.n21036 4.5005
R3777 DVDD.n21048 DVDD.n21022 4.5005
R3778 DVDD.n21048 DVDD.n21039 4.5005
R3779 DVDD.n21048 DVDD.n21021 4.5005
R3780 DVDD.n21048 DVDD.n21042 4.5005
R3781 DVDD.n21048 DVDD.n21020 4.5005
R3782 DVDD.n21048 DVDD.n21044 4.5005
R3783 DVDD.n21048 DVDD.n21019 4.5005
R3784 DVDD.n19101 DVDD.n19100 4.5005
R3785 DVDD.n19100 DVDD.n18819 4.5005
R3786 DVDD.n20925 DVDD.n20923 4.5005
R3787 DVDD.n20926 DVDD.n20925 4.5005
R3788 DVDD.n20922 DVDD.n18909 4.5005
R3789 DVDD.n20922 DVDD.n18820 4.5005
R3790 DVDD.n20919 DVDD.n18909 4.5005
R3791 DVDD.n20919 DVDD.n20908 4.5005
R3792 DVDD.n20919 DVDD.n20906 4.5005
R3793 DVDD.n20919 DVDD.n20910 4.5005
R3794 DVDD.n20919 DVDD.n20905 4.5005
R3795 DVDD.n20919 DVDD.n20912 4.5005
R3796 DVDD.n20919 DVDD.n20904 4.5005
R3797 DVDD.n20919 DVDD.n20914 4.5005
R3798 DVDD.n20919 DVDD.n20903 4.5005
R3799 DVDD.n20919 DVDD.n20916 4.5005
R3800 DVDD.n20919 DVDD.n20902 4.5005
R3801 DVDD.n20919 DVDD.n20918 4.5005
R3802 DVDD.n20919 DVDD.n20901 4.5005
R3803 DVDD.n20920 DVDD.n20919 4.5005
R3804 DVDD.n20919 DVDD.n18820 4.5005
R3805 DVDD.n21048 DVDD.n21047 4.5005
R3806 DVDD.n20919 DVDD.n18917 4.5005
R3807 DVDD.n10057 DVDD.n9741 4.5005
R3808 DVDD.n9957 DVDD.n9741 4.5005
R3809 DVDD.n9754 DVDD.n9741 4.5005
R3810 DVDD.n9958 DVDD.n9741 4.5005
R3811 DVDD.n9753 DVDD.n9741 4.5005
R3812 DVDD.n9959 DVDD.n9741 4.5005
R3813 DVDD.n9752 DVDD.n9741 4.5005
R3814 DVDD.n9962 DVDD.n9741 4.5005
R3815 DVDD.n10001 DVDD.n9741 4.5005
R3816 DVDD.n9963 DVDD.n9741 4.5005
R3817 DVDD.n9750 DVDD.n9741 4.5005
R3818 DVDD.n10055 DVDD.n9741 4.5005
R3819 DVDD.n10057 DVDD.n9737 4.5005
R3820 DVDD.n9956 DVDD.n9737 4.5005
R3821 DVDD.n9755 DVDD.n9737 4.5005
R3822 DVDD.n9957 DVDD.n9737 4.5005
R3823 DVDD.n9754 DVDD.n9737 4.5005
R3824 DVDD.n9958 DVDD.n9737 4.5005
R3825 DVDD.n9753 DVDD.n9737 4.5005
R3826 DVDD.n9959 DVDD.n9737 4.5005
R3827 DVDD.n9752 DVDD.n9737 4.5005
R3828 DVDD.n9961 DVDD.n9737 4.5005
R3829 DVDD.n9751 DVDD.n9737 4.5005
R3830 DVDD.n9962 DVDD.n9737 4.5005
R3831 DVDD.n9963 DVDD.n9737 4.5005
R3832 DVDD.n10055 DVDD.n9737 4.5005
R3833 DVDD.n10057 DVDD.n9742 4.5005
R3834 DVDD.n9956 DVDD.n9742 4.5005
R3835 DVDD.n9755 DVDD.n9742 4.5005
R3836 DVDD.n9957 DVDD.n9742 4.5005
R3837 DVDD.n9754 DVDD.n9742 4.5005
R3838 DVDD.n9958 DVDD.n9742 4.5005
R3839 DVDD.n9753 DVDD.n9742 4.5005
R3840 DVDD.n9959 DVDD.n9742 4.5005
R3841 DVDD.n9752 DVDD.n9742 4.5005
R3842 DVDD.n9961 DVDD.n9742 4.5005
R3843 DVDD.n9751 DVDD.n9742 4.5005
R3844 DVDD.n9962 DVDD.n9742 4.5005
R3845 DVDD.n9963 DVDD.n9742 4.5005
R3846 DVDD.n10055 DVDD.n9742 4.5005
R3847 DVDD.n10057 DVDD.n9736 4.5005
R3848 DVDD.n9956 DVDD.n9736 4.5005
R3849 DVDD.n9755 DVDD.n9736 4.5005
R3850 DVDD.n9957 DVDD.n9736 4.5005
R3851 DVDD.n9754 DVDD.n9736 4.5005
R3852 DVDD.n9958 DVDD.n9736 4.5005
R3853 DVDD.n9753 DVDD.n9736 4.5005
R3854 DVDD.n9959 DVDD.n9736 4.5005
R3855 DVDD.n9752 DVDD.n9736 4.5005
R3856 DVDD.n9961 DVDD.n9736 4.5005
R3857 DVDD.n9751 DVDD.n9736 4.5005
R3858 DVDD.n9962 DVDD.n9736 4.5005
R3859 DVDD.n9963 DVDD.n9736 4.5005
R3860 DVDD.n9750 DVDD.n9736 4.5005
R3861 DVDD.n10055 DVDD.n9736 4.5005
R3862 DVDD.n10057 DVDD.n9743 4.5005
R3863 DVDD.n9956 DVDD.n9743 4.5005
R3864 DVDD.n9755 DVDD.n9743 4.5005
R3865 DVDD.n9957 DVDD.n9743 4.5005
R3866 DVDD.n9754 DVDD.n9743 4.5005
R3867 DVDD.n9958 DVDD.n9743 4.5005
R3868 DVDD.n9753 DVDD.n9743 4.5005
R3869 DVDD.n9959 DVDD.n9743 4.5005
R3870 DVDD.n9752 DVDD.n9743 4.5005
R3871 DVDD.n9961 DVDD.n9743 4.5005
R3872 DVDD.n9751 DVDD.n9743 4.5005
R3873 DVDD.n9962 DVDD.n9743 4.5005
R3874 DVDD.n9963 DVDD.n9743 4.5005
R3875 DVDD.n10055 DVDD.n9743 4.5005
R3876 DVDD.n10057 DVDD.n9735 4.5005
R3877 DVDD.n9956 DVDD.n9735 4.5005
R3878 DVDD.n9755 DVDD.n9735 4.5005
R3879 DVDD.n9957 DVDD.n9735 4.5005
R3880 DVDD.n9754 DVDD.n9735 4.5005
R3881 DVDD.n9958 DVDD.n9735 4.5005
R3882 DVDD.n9753 DVDD.n9735 4.5005
R3883 DVDD.n9959 DVDD.n9735 4.5005
R3884 DVDD.n9752 DVDD.n9735 4.5005
R3885 DVDD.n9961 DVDD.n9735 4.5005
R3886 DVDD.n9751 DVDD.n9735 4.5005
R3887 DVDD.n9962 DVDD.n9735 4.5005
R3888 DVDD.n9963 DVDD.n9735 4.5005
R3889 DVDD.n10055 DVDD.n9735 4.5005
R3890 DVDD.n10057 DVDD.n9744 4.5005
R3891 DVDD.n9956 DVDD.n9744 4.5005
R3892 DVDD.n9755 DVDD.n9744 4.5005
R3893 DVDD.n9957 DVDD.n9744 4.5005
R3894 DVDD.n9754 DVDD.n9744 4.5005
R3895 DVDD.n9958 DVDD.n9744 4.5005
R3896 DVDD.n9753 DVDD.n9744 4.5005
R3897 DVDD.n9959 DVDD.n9744 4.5005
R3898 DVDD.n9752 DVDD.n9744 4.5005
R3899 DVDD.n9961 DVDD.n9744 4.5005
R3900 DVDD.n9751 DVDD.n9744 4.5005
R3901 DVDD.n9962 DVDD.n9744 4.5005
R3902 DVDD.n9963 DVDD.n9744 4.5005
R3903 DVDD.n9750 DVDD.n9744 4.5005
R3904 DVDD.n10055 DVDD.n9744 4.5005
R3905 DVDD.n10057 DVDD.n9734 4.5005
R3906 DVDD.n9956 DVDD.n9734 4.5005
R3907 DVDD.n9755 DVDD.n9734 4.5005
R3908 DVDD.n9957 DVDD.n9734 4.5005
R3909 DVDD.n9754 DVDD.n9734 4.5005
R3910 DVDD.n9958 DVDD.n9734 4.5005
R3911 DVDD.n9753 DVDD.n9734 4.5005
R3912 DVDD.n9959 DVDD.n9734 4.5005
R3913 DVDD.n9752 DVDD.n9734 4.5005
R3914 DVDD.n9961 DVDD.n9734 4.5005
R3915 DVDD.n9751 DVDD.n9734 4.5005
R3916 DVDD.n9962 DVDD.n9734 4.5005
R3917 DVDD.n10001 DVDD.n9734 4.5005
R3918 DVDD.n9963 DVDD.n9734 4.5005
R3919 DVDD.n10055 DVDD.n9734 4.5005
R3920 DVDD.n2962 DVDD.n2936 4.5005
R3921 DVDD.n2966 DVDD.n2936 4.5005
R3922 DVDD.n2960 DVDD.n2936 4.5005
R3923 DVDD.n2967 DVDD.n2936 4.5005
R3924 DVDD.n2959 DVDD.n2936 4.5005
R3925 DVDD.n2968 DVDD.n2936 4.5005
R3926 DVDD.n2958 DVDD.n2936 4.5005
R3927 DVDD.n2971 DVDD.n2936 4.5005
R3928 DVDD.n2980 DVDD.n2936 4.5005
R3929 DVDD.n16182 DVDD.n2936 4.5005
R3930 DVDD.n16184 DVDD.n2936 4.5005
R3931 DVDD.n2962 DVDD.n2938 4.5005
R3932 DVDD.n2965 DVDD.n2938 4.5005
R3933 DVDD.n2961 DVDD.n2938 4.5005
R3934 DVDD.n2966 DVDD.n2938 4.5005
R3935 DVDD.n2960 DVDD.n2938 4.5005
R3936 DVDD.n2967 DVDD.n2938 4.5005
R3937 DVDD.n2959 DVDD.n2938 4.5005
R3938 DVDD.n2968 DVDD.n2938 4.5005
R3939 DVDD.n2958 DVDD.n2938 4.5005
R3940 DVDD.n2970 DVDD.n2938 4.5005
R3941 DVDD.n2957 DVDD.n2938 4.5005
R3942 DVDD.n2971 DVDD.n2938 4.5005
R3943 DVDD.n16182 DVDD.n2938 4.5005
R3944 DVDD.n16184 DVDD.n2938 4.5005
R3945 DVDD.n2962 DVDD.n2935 4.5005
R3946 DVDD.n2965 DVDD.n2935 4.5005
R3947 DVDD.n2961 DVDD.n2935 4.5005
R3948 DVDD.n2966 DVDD.n2935 4.5005
R3949 DVDD.n2960 DVDD.n2935 4.5005
R3950 DVDD.n2967 DVDD.n2935 4.5005
R3951 DVDD.n2959 DVDD.n2935 4.5005
R3952 DVDD.n2968 DVDD.n2935 4.5005
R3953 DVDD.n2958 DVDD.n2935 4.5005
R3954 DVDD.n2970 DVDD.n2935 4.5005
R3955 DVDD.n2957 DVDD.n2935 4.5005
R3956 DVDD.n2971 DVDD.n2935 4.5005
R3957 DVDD.n16182 DVDD.n2935 4.5005
R3958 DVDD.n2935 DVDD.n2924 4.5005
R3959 DVDD.n16184 DVDD.n2935 4.5005
R3960 DVDD.n2962 DVDD.n2940 4.5005
R3961 DVDD.n2965 DVDD.n2940 4.5005
R3962 DVDD.n2961 DVDD.n2940 4.5005
R3963 DVDD.n2966 DVDD.n2940 4.5005
R3964 DVDD.n2960 DVDD.n2940 4.5005
R3965 DVDD.n2967 DVDD.n2940 4.5005
R3966 DVDD.n2959 DVDD.n2940 4.5005
R3967 DVDD.n2968 DVDD.n2940 4.5005
R3968 DVDD.n2958 DVDD.n2940 4.5005
R3969 DVDD.n2970 DVDD.n2940 4.5005
R3970 DVDD.n2957 DVDD.n2940 4.5005
R3971 DVDD.n2971 DVDD.n2940 4.5005
R3972 DVDD.n16182 DVDD.n2940 4.5005
R3973 DVDD.n16184 DVDD.n2940 4.5005
R3974 DVDD.n2962 DVDD.n2934 4.5005
R3975 DVDD.n2965 DVDD.n2934 4.5005
R3976 DVDD.n2961 DVDD.n2934 4.5005
R3977 DVDD.n2966 DVDD.n2934 4.5005
R3978 DVDD.n2960 DVDD.n2934 4.5005
R3979 DVDD.n2967 DVDD.n2934 4.5005
R3980 DVDD.n2959 DVDD.n2934 4.5005
R3981 DVDD.n2968 DVDD.n2934 4.5005
R3982 DVDD.n2958 DVDD.n2934 4.5005
R3983 DVDD.n2970 DVDD.n2934 4.5005
R3984 DVDD.n2957 DVDD.n2934 4.5005
R3985 DVDD.n2971 DVDD.n2934 4.5005
R3986 DVDD.n16182 DVDD.n2934 4.5005
R3987 DVDD.n16184 DVDD.n2934 4.5005
R3988 DVDD.n2962 DVDD.n2941 4.5005
R3989 DVDD.n2965 DVDD.n2941 4.5005
R3990 DVDD.n2961 DVDD.n2941 4.5005
R3991 DVDD.n2966 DVDD.n2941 4.5005
R3992 DVDD.n2960 DVDD.n2941 4.5005
R3993 DVDD.n2967 DVDD.n2941 4.5005
R3994 DVDD.n2959 DVDD.n2941 4.5005
R3995 DVDD.n2968 DVDD.n2941 4.5005
R3996 DVDD.n2958 DVDD.n2941 4.5005
R3997 DVDD.n2970 DVDD.n2941 4.5005
R3998 DVDD.n2957 DVDD.n2941 4.5005
R3999 DVDD.n2971 DVDD.n2941 4.5005
R4000 DVDD.n16182 DVDD.n2941 4.5005
R4001 DVDD.n2941 DVDD.n2924 4.5005
R4002 DVDD.n16184 DVDD.n2941 4.5005
R4003 DVDD.n2962 DVDD.n2933 4.5005
R4004 DVDD.n2965 DVDD.n2933 4.5005
R4005 DVDD.n2961 DVDD.n2933 4.5005
R4006 DVDD.n2966 DVDD.n2933 4.5005
R4007 DVDD.n2960 DVDD.n2933 4.5005
R4008 DVDD.n2967 DVDD.n2933 4.5005
R4009 DVDD.n2959 DVDD.n2933 4.5005
R4010 DVDD.n2968 DVDD.n2933 4.5005
R4011 DVDD.n2958 DVDD.n2933 4.5005
R4012 DVDD.n2970 DVDD.n2933 4.5005
R4013 DVDD.n2957 DVDD.n2933 4.5005
R4014 DVDD.n2971 DVDD.n2933 4.5005
R4015 DVDD.n16182 DVDD.n2933 4.5005
R4016 DVDD.n16184 DVDD.n2933 4.5005
R4017 DVDD.n2962 DVDD.n2943 4.5005
R4018 DVDD.n2965 DVDD.n2943 4.5005
R4019 DVDD.n2961 DVDD.n2943 4.5005
R4020 DVDD.n2966 DVDD.n2943 4.5005
R4021 DVDD.n2960 DVDD.n2943 4.5005
R4022 DVDD.n2967 DVDD.n2943 4.5005
R4023 DVDD.n2959 DVDD.n2943 4.5005
R4024 DVDD.n2968 DVDD.n2943 4.5005
R4025 DVDD.n2958 DVDD.n2943 4.5005
R4026 DVDD.n2970 DVDD.n2943 4.5005
R4027 DVDD.n2957 DVDD.n2943 4.5005
R4028 DVDD.n2971 DVDD.n2943 4.5005
R4029 DVDD.n16182 DVDD.n2943 4.5005
R4030 DVDD.n16184 DVDD.n2943 4.5005
R4031 DVDD.n2962 DVDD.n2932 4.5005
R4032 DVDD.n2965 DVDD.n2932 4.5005
R4033 DVDD.n2961 DVDD.n2932 4.5005
R4034 DVDD.n2966 DVDD.n2932 4.5005
R4035 DVDD.n2960 DVDD.n2932 4.5005
R4036 DVDD.n2967 DVDD.n2932 4.5005
R4037 DVDD.n2959 DVDD.n2932 4.5005
R4038 DVDD.n2968 DVDD.n2932 4.5005
R4039 DVDD.n2958 DVDD.n2932 4.5005
R4040 DVDD.n2970 DVDD.n2932 4.5005
R4041 DVDD.n2957 DVDD.n2932 4.5005
R4042 DVDD.n2971 DVDD.n2932 4.5005
R4043 DVDD.n16182 DVDD.n2932 4.5005
R4044 DVDD.n2932 DVDD.n2924 4.5005
R4045 DVDD.n16184 DVDD.n2932 4.5005
R4046 DVDD.n2962 DVDD.n2945 4.5005
R4047 DVDD.n2965 DVDD.n2945 4.5005
R4048 DVDD.n2961 DVDD.n2945 4.5005
R4049 DVDD.n2966 DVDD.n2945 4.5005
R4050 DVDD.n2960 DVDD.n2945 4.5005
R4051 DVDD.n2967 DVDD.n2945 4.5005
R4052 DVDD.n2959 DVDD.n2945 4.5005
R4053 DVDD.n2968 DVDD.n2945 4.5005
R4054 DVDD.n2958 DVDD.n2945 4.5005
R4055 DVDD.n2970 DVDD.n2945 4.5005
R4056 DVDD.n2957 DVDD.n2945 4.5005
R4057 DVDD.n2971 DVDD.n2945 4.5005
R4058 DVDD.n16182 DVDD.n2945 4.5005
R4059 DVDD.n16184 DVDD.n2945 4.5005
R4060 DVDD.n2962 DVDD.n2931 4.5005
R4061 DVDD.n2965 DVDD.n2931 4.5005
R4062 DVDD.n2961 DVDD.n2931 4.5005
R4063 DVDD.n2966 DVDD.n2931 4.5005
R4064 DVDD.n2960 DVDD.n2931 4.5005
R4065 DVDD.n2967 DVDD.n2931 4.5005
R4066 DVDD.n2959 DVDD.n2931 4.5005
R4067 DVDD.n2968 DVDD.n2931 4.5005
R4068 DVDD.n2958 DVDD.n2931 4.5005
R4069 DVDD.n2970 DVDD.n2931 4.5005
R4070 DVDD.n2957 DVDD.n2931 4.5005
R4071 DVDD.n2971 DVDD.n2931 4.5005
R4072 DVDD.n16182 DVDD.n2931 4.5005
R4073 DVDD.n16184 DVDD.n2931 4.5005
R4074 DVDD.n2962 DVDD.n2946 4.5005
R4075 DVDD.n2965 DVDD.n2946 4.5005
R4076 DVDD.n2961 DVDD.n2946 4.5005
R4077 DVDD.n2966 DVDD.n2946 4.5005
R4078 DVDD.n2960 DVDD.n2946 4.5005
R4079 DVDD.n2967 DVDD.n2946 4.5005
R4080 DVDD.n2959 DVDD.n2946 4.5005
R4081 DVDD.n2968 DVDD.n2946 4.5005
R4082 DVDD.n2958 DVDD.n2946 4.5005
R4083 DVDD.n2970 DVDD.n2946 4.5005
R4084 DVDD.n2957 DVDD.n2946 4.5005
R4085 DVDD.n2971 DVDD.n2946 4.5005
R4086 DVDD.n16182 DVDD.n2946 4.5005
R4087 DVDD.n2946 DVDD.n2924 4.5005
R4088 DVDD.n16184 DVDD.n2946 4.5005
R4089 DVDD.n2962 DVDD.n2930 4.5005
R4090 DVDD.n2965 DVDD.n2930 4.5005
R4091 DVDD.n2961 DVDD.n2930 4.5005
R4092 DVDD.n2966 DVDD.n2930 4.5005
R4093 DVDD.n2960 DVDD.n2930 4.5005
R4094 DVDD.n2967 DVDD.n2930 4.5005
R4095 DVDD.n2959 DVDD.n2930 4.5005
R4096 DVDD.n2968 DVDD.n2930 4.5005
R4097 DVDD.n2958 DVDD.n2930 4.5005
R4098 DVDD.n2970 DVDD.n2930 4.5005
R4099 DVDD.n2957 DVDD.n2930 4.5005
R4100 DVDD.n2971 DVDD.n2930 4.5005
R4101 DVDD.n2980 DVDD.n2930 4.5005
R4102 DVDD.n16182 DVDD.n2930 4.5005
R4103 DVDD.n16184 DVDD.n2930 4.5005
R4104 DVDD.n2962 DVDD.n2948 4.5005
R4105 DVDD.n2965 DVDD.n2948 4.5005
R4106 DVDD.n2961 DVDD.n2948 4.5005
R4107 DVDD.n2966 DVDD.n2948 4.5005
R4108 DVDD.n2960 DVDD.n2948 4.5005
R4109 DVDD.n2967 DVDD.n2948 4.5005
R4110 DVDD.n2959 DVDD.n2948 4.5005
R4111 DVDD.n2968 DVDD.n2948 4.5005
R4112 DVDD.n2958 DVDD.n2948 4.5005
R4113 DVDD.n2970 DVDD.n2948 4.5005
R4114 DVDD.n2957 DVDD.n2948 4.5005
R4115 DVDD.n2971 DVDD.n2948 4.5005
R4116 DVDD.n16182 DVDD.n2948 4.5005
R4117 DVDD.n16184 DVDD.n2948 4.5005
R4118 DVDD.n2962 DVDD.n2929 4.5005
R4119 DVDD.n2965 DVDD.n2929 4.5005
R4120 DVDD.n2961 DVDD.n2929 4.5005
R4121 DVDD.n2966 DVDD.n2929 4.5005
R4122 DVDD.n2960 DVDD.n2929 4.5005
R4123 DVDD.n2967 DVDD.n2929 4.5005
R4124 DVDD.n2959 DVDD.n2929 4.5005
R4125 DVDD.n2968 DVDD.n2929 4.5005
R4126 DVDD.n2958 DVDD.n2929 4.5005
R4127 DVDD.n2970 DVDD.n2929 4.5005
R4128 DVDD.n2957 DVDD.n2929 4.5005
R4129 DVDD.n2971 DVDD.n2929 4.5005
R4130 DVDD.n16182 DVDD.n2929 4.5005
R4131 DVDD.n16184 DVDD.n2929 4.5005
R4132 DVDD.n2962 DVDD.n2950 4.5005
R4133 DVDD.n2965 DVDD.n2950 4.5005
R4134 DVDD.n2961 DVDD.n2950 4.5005
R4135 DVDD.n2966 DVDD.n2950 4.5005
R4136 DVDD.n2960 DVDD.n2950 4.5005
R4137 DVDD.n2967 DVDD.n2950 4.5005
R4138 DVDD.n2959 DVDD.n2950 4.5005
R4139 DVDD.n2968 DVDD.n2950 4.5005
R4140 DVDD.n2958 DVDD.n2950 4.5005
R4141 DVDD.n2970 DVDD.n2950 4.5005
R4142 DVDD.n2957 DVDD.n2950 4.5005
R4143 DVDD.n2971 DVDD.n2950 4.5005
R4144 DVDD.n2980 DVDD.n2950 4.5005
R4145 DVDD.n16182 DVDD.n2950 4.5005
R4146 DVDD.n16184 DVDD.n2950 4.5005
R4147 DVDD.n2962 DVDD.n2928 4.5005
R4148 DVDD.n2965 DVDD.n2928 4.5005
R4149 DVDD.n2961 DVDD.n2928 4.5005
R4150 DVDD.n2966 DVDD.n2928 4.5005
R4151 DVDD.n2960 DVDD.n2928 4.5005
R4152 DVDD.n2967 DVDD.n2928 4.5005
R4153 DVDD.n2959 DVDD.n2928 4.5005
R4154 DVDD.n2968 DVDD.n2928 4.5005
R4155 DVDD.n2958 DVDD.n2928 4.5005
R4156 DVDD.n2970 DVDD.n2928 4.5005
R4157 DVDD.n2957 DVDD.n2928 4.5005
R4158 DVDD.n2971 DVDD.n2928 4.5005
R4159 DVDD.n2980 DVDD.n2928 4.5005
R4160 DVDD.n16182 DVDD.n2928 4.5005
R4161 DVDD.n16184 DVDD.n2928 4.5005
R4162 DVDD.n2962 DVDD.n2952 4.5005
R4163 DVDD.n2965 DVDD.n2952 4.5005
R4164 DVDD.n2961 DVDD.n2952 4.5005
R4165 DVDD.n2966 DVDD.n2952 4.5005
R4166 DVDD.n2960 DVDD.n2952 4.5005
R4167 DVDD.n2967 DVDD.n2952 4.5005
R4168 DVDD.n2959 DVDD.n2952 4.5005
R4169 DVDD.n2968 DVDD.n2952 4.5005
R4170 DVDD.n2958 DVDD.n2952 4.5005
R4171 DVDD.n2970 DVDD.n2952 4.5005
R4172 DVDD.n2957 DVDD.n2952 4.5005
R4173 DVDD.n2971 DVDD.n2952 4.5005
R4174 DVDD.n16182 DVDD.n2952 4.5005
R4175 DVDD.n16184 DVDD.n2952 4.5005
R4176 DVDD.n2962 DVDD.n2927 4.5005
R4177 DVDD.n2965 DVDD.n2927 4.5005
R4178 DVDD.n2961 DVDD.n2927 4.5005
R4179 DVDD.n2966 DVDD.n2927 4.5005
R4180 DVDD.n2960 DVDD.n2927 4.5005
R4181 DVDD.n2967 DVDD.n2927 4.5005
R4182 DVDD.n2959 DVDD.n2927 4.5005
R4183 DVDD.n2968 DVDD.n2927 4.5005
R4184 DVDD.n2958 DVDD.n2927 4.5005
R4185 DVDD.n2970 DVDD.n2927 4.5005
R4186 DVDD.n2957 DVDD.n2927 4.5005
R4187 DVDD.n2971 DVDD.n2927 4.5005
R4188 DVDD.n16182 DVDD.n2927 4.5005
R4189 DVDD.n16184 DVDD.n2927 4.5005
R4190 DVDD.n2962 DVDD.n2954 4.5005
R4191 DVDD.n2965 DVDD.n2954 4.5005
R4192 DVDD.n2961 DVDD.n2954 4.5005
R4193 DVDD.n2966 DVDD.n2954 4.5005
R4194 DVDD.n2960 DVDD.n2954 4.5005
R4195 DVDD.n2967 DVDD.n2954 4.5005
R4196 DVDD.n2959 DVDD.n2954 4.5005
R4197 DVDD.n2968 DVDD.n2954 4.5005
R4198 DVDD.n2958 DVDD.n2954 4.5005
R4199 DVDD.n2970 DVDD.n2954 4.5005
R4200 DVDD.n2957 DVDD.n2954 4.5005
R4201 DVDD.n2971 DVDD.n2954 4.5005
R4202 DVDD.n2980 DVDD.n2954 4.5005
R4203 DVDD.n16182 DVDD.n2954 4.5005
R4204 DVDD.n16184 DVDD.n2954 4.5005
R4205 DVDD.n2962 DVDD.n2926 4.5005
R4206 DVDD.n2965 DVDD.n2926 4.5005
R4207 DVDD.n2961 DVDD.n2926 4.5005
R4208 DVDD.n2966 DVDD.n2926 4.5005
R4209 DVDD.n2960 DVDD.n2926 4.5005
R4210 DVDD.n2967 DVDD.n2926 4.5005
R4211 DVDD.n2959 DVDD.n2926 4.5005
R4212 DVDD.n2968 DVDD.n2926 4.5005
R4213 DVDD.n2958 DVDD.n2926 4.5005
R4214 DVDD.n2970 DVDD.n2926 4.5005
R4215 DVDD.n2957 DVDD.n2926 4.5005
R4216 DVDD.n2971 DVDD.n2926 4.5005
R4217 DVDD.n2980 DVDD.n2926 4.5005
R4218 DVDD.n16182 DVDD.n2926 4.5005
R4219 DVDD.n2926 DVDD.n2924 4.5005
R4220 DVDD.n16184 DVDD.n2926 4.5005
R4221 DVDD.n16248 DVDD.n2791 4.5005
R4222 DVDD.n2825 DVDD.n2791 4.5005
R4223 DVDD.n2821 DVDD.n2791 4.5005
R4224 DVDD.n2826 DVDD.n2791 4.5005
R4225 DVDD.n2820 DVDD.n2791 4.5005
R4226 DVDD.n2827 DVDD.n2791 4.5005
R4227 DVDD.n2819 DVDD.n2791 4.5005
R4228 DVDD.n2830 DVDD.n2791 4.5005
R4229 DVDD.n2872 DVDD.n2791 4.5005
R4230 DVDD.n2831 DVDD.n2791 4.5005
R4231 DVDD.n2816 DVDD.n2791 4.5005
R4232 DVDD.n16246 DVDD.n2791 4.5005
R4233 DVDD.n16248 DVDD.n2793 4.5005
R4234 DVDD.n2824 DVDD.n2793 4.5005
R4235 DVDD.n2822 DVDD.n2793 4.5005
R4236 DVDD.n2825 DVDD.n2793 4.5005
R4237 DVDD.n2821 DVDD.n2793 4.5005
R4238 DVDD.n2826 DVDD.n2793 4.5005
R4239 DVDD.n2820 DVDD.n2793 4.5005
R4240 DVDD.n2827 DVDD.n2793 4.5005
R4241 DVDD.n2819 DVDD.n2793 4.5005
R4242 DVDD.n2829 DVDD.n2793 4.5005
R4243 DVDD.n2818 DVDD.n2793 4.5005
R4244 DVDD.n2830 DVDD.n2793 4.5005
R4245 DVDD.n2872 DVDD.n2793 4.5005
R4246 DVDD.n2831 DVDD.n2793 4.5005
R4247 DVDD.n16246 DVDD.n2793 4.5005
R4248 DVDD.n16248 DVDD.n2790 4.5005
R4249 DVDD.n2824 DVDD.n2790 4.5005
R4250 DVDD.n2822 DVDD.n2790 4.5005
R4251 DVDD.n2825 DVDD.n2790 4.5005
R4252 DVDD.n2821 DVDD.n2790 4.5005
R4253 DVDD.n2826 DVDD.n2790 4.5005
R4254 DVDD.n2820 DVDD.n2790 4.5005
R4255 DVDD.n2827 DVDD.n2790 4.5005
R4256 DVDD.n2819 DVDD.n2790 4.5005
R4257 DVDD.n2829 DVDD.n2790 4.5005
R4258 DVDD.n2818 DVDD.n2790 4.5005
R4259 DVDD.n2830 DVDD.n2790 4.5005
R4260 DVDD.n2831 DVDD.n2790 4.5005
R4261 DVDD.n16246 DVDD.n2790 4.5005
R4262 DVDD.n16248 DVDD.n2794 4.5005
R4263 DVDD.n2824 DVDD.n2794 4.5005
R4264 DVDD.n2822 DVDD.n2794 4.5005
R4265 DVDD.n2825 DVDD.n2794 4.5005
R4266 DVDD.n2821 DVDD.n2794 4.5005
R4267 DVDD.n2826 DVDD.n2794 4.5005
R4268 DVDD.n2820 DVDD.n2794 4.5005
R4269 DVDD.n2827 DVDD.n2794 4.5005
R4270 DVDD.n2819 DVDD.n2794 4.5005
R4271 DVDD.n2829 DVDD.n2794 4.5005
R4272 DVDD.n2818 DVDD.n2794 4.5005
R4273 DVDD.n2830 DVDD.n2794 4.5005
R4274 DVDD.n2831 DVDD.n2794 4.5005
R4275 DVDD.n16246 DVDD.n2794 4.5005
R4276 DVDD.n16248 DVDD.n2789 4.5005
R4277 DVDD.n2824 DVDD.n2789 4.5005
R4278 DVDD.n2822 DVDD.n2789 4.5005
R4279 DVDD.n2825 DVDD.n2789 4.5005
R4280 DVDD.n2821 DVDD.n2789 4.5005
R4281 DVDD.n2826 DVDD.n2789 4.5005
R4282 DVDD.n2820 DVDD.n2789 4.5005
R4283 DVDD.n2827 DVDD.n2789 4.5005
R4284 DVDD.n2819 DVDD.n2789 4.5005
R4285 DVDD.n2829 DVDD.n2789 4.5005
R4286 DVDD.n2818 DVDD.n2789 4.5005
R4287 DVDD.n2830 DVDD.n2789 4.5005
R4288 DVDD.n2872 DVDD.n2789 4.5005
R4289 DVDD.n2831 DVDD.n2789 4.5005
R4290 DVDD.n16246 DVDD.n2789 4.5005
R4291 DVDD.n16248 DVDD.n2795 4.5005
R4292 DVDD.n2824 DVDD.n2795 4.5005
R4293 DVDD.n2822 DVDD.n2795 4.5005
R4294 DVDD.n2825 DVDD.n2795 4.5005
R4295 DVDD.n2821 DVDD.n2795 4.5005
R4296 DVDD.n2826 DVDD.n2795 4.5005
R4297 DVDD.n2820 DVDD.n2795 4.5005
R4298 DVDD.n2827 DVDD.n2795 4.5005
R4299 DVDD.n2819 DVDD.n2795 4.5005
R4300 DVDD.n2829 DVDD.n2795 4.5005
R4301 DVDD.n2818 DVDD.n2795 4.5005
R4302 DVDD.n2830 DVDD.n2795 4.5005
R4303 DVDD.n2872 DVDD.n2795 4.5005
R4304 DVDD.n2831 DVDD.n2795 4.5005
R4305 DVDD.n16246 DVDD.n2795 4.5005
R4306 DVDD.n16248 DVDD.n2788 4.5005
R4307 DVDD.n2824 DVDD.n2788 4.5005
R4308 DVDD.n2822 DVDD.n2788 4.5005
R4309 DVDD.n2825 DVDD.n2788 4.5005
R4310 DVDD.n2821 DVDD.n2788 4.5005
R4311 DVDD.n2826 DVDD.n2788 4.5005
R4312 DVDD.n2820 DVDD.n2788 4.5005
R4313 DVDD.n2827 DVDD.n2788 4.5005
R4314 DVDD.n2819 DVDD.n2788 4.5005
R4315 DVDD.n2829 DVDD.n2788 4.5005
R4316 DVDD.n2818 DVDD.n2788 4.5005
R4317 DVDD.n2830 DVDD.n2788 4.5005
R4318 DVDD.n2831 DVDD.n2788 4.5005
R4319 DVDD.n16246 DVDD.n2788 4.5005
R4320 DVDD.n16248 DVDD.n2796 4.5005
R4321 DVDD.n2824 DVDD.n2796 4.5005
R4322 DVDD.n2822 DVDD.n2796 4.5005
R4323 DVDD.n2825 DVDD.n2796 4.5005
R4324 DVDD.n2821 DVDD.n2796 4.5005
R4325 DVDD.n2826 DVDD.n2796 4.5005
R4326 DVDD.n2820 DVDD.n2796 4.5005
R4327 DVDD.n2827 DVDD.n2796 4.5005
R4328 DVDD.n2819 DVDD.n2796 4.5005
R4329 DVDD.n2829 DVDD.n2796 4.5005
R4330 DVDD.n2818 DVDD.n2796 4.5005
R4331 DVDD.n2830 DVDD.n2796 4.5005
R4332 DVDD.n2831 DVDD.n2796 4.5005
R4333 DVDD.n16246 DVDD.n2796 4.5005
R4334 DVDD.n16248 DVDD.n2787 4.5005
R4335 DVDD.n2824 DVDD.n2787 4.5005
R4336 DVDD.n2822 DVDD.n2787 4.5005
R4337 DVDD.n2825 DVDD.n2787 4.5005
R4338 DVDD.n2821 DVDD.n2787 4.5005
R4339 DVDD.n2826 DVDD.n2787 4.5005
R4340 DVDD.n2820 DVDD.n2787 4.5005
R4341 DVDD.n2827 DVDD.n2787 4.5005
R4342 DVDD.n2819 DVDD.n2787 4.5005
R4343 DVDD.n2829 DVDD.n2787 4.5005
R4344 DVDD.n2818 DVDD.n2787 4.5005
R4345 DVDD.n2830 DVDD.n2787 4.5005
R4346 DVDD.n2872 DVDD.n2787 4.5005
R4347 DVDD.n2831 DVDD.n2787 4.5005
R4348 DVDD.n16246 DVDD.n2787 4.5005
R4349 DVDD.n16248 DVDD.n2797 4.5005
R4350 DVDD.n2824 DVDD.n2797 4.5005
R4351 DVDD.n2822 DVDD.n2797 4.5005
R4352 DVDD.n2825 DVDD.n2797 4.5005
R4353 DVDD.n2821 DVDD.n2797 4.5005
R4354 DVDD.n2826 DVDD.n2797 4.5005
R4355 DVDD.n2820 DVDD.n2797 4.5005
R4356 DVDD.n2827 DVDD.n2797 4.5005
R4357 DVDD.n2819 DVDD.n2797 4.5005
R4358 DVDD.n2829 DVDD.n2797 4.5005
R4359 DVDD.n2818 DVDD.n2797 4.5005
R4360 DVDD.n2830 DVDD.n2797 4.5005
R4361 DVDD.n2872 DVDD.n2797 4.5005
R4362 DVDD.n2831 DVDD.n2797 4.5005
R4363 DVDD.n16246 DVDD.n2797 4.5005
R4364 DVDD.n16248 DVDD.n2786 4.5005
R4365 DVDD.n2824 DVDD.n2786 4.5005
R4366 DVDD.n2822 DVDD.n2786 4.5005
R4367 DVDD.n2825 DVDD.n2786 4.5005
R4368 DVDD.n2821 DVDD.n2786 4.5005
R4369 DVDD.n2826 DVDD.n2786 4.5005
R4370 DVDD.n2820 DVDD.n2786 4.5005
R4371 DVDD.n2827 DVDD.n2786 4.5005
R4372 DVDD.n2819 DVDD.n2786 4.5005
R4373 DVDD.n2829 DVDD.n2786 4.5005
R4374 DVDD.n2818 DVDD.n2786 4.5005
R4375 DVDD.n2830 DVDD.n2786 4.5005
R4376 DVDD.n2831 DVDD.n2786 4.5005
R4377 DVDD.n16246 DVDD.n2786 4.5005
R4378 DVDD.n16248 DVDD.n2798 4.5005
R4379 DVDD.n2824 DVDD.n2798 4.5005
R4380 DVDD.n2822 DVDD.n2798 4.5005
R4381 DVDD.n2825 DVDD.n2798 4.5005
R4382 DVDD.n2821 DVDD.n2798 4.5005
R4383 DVDD.n2826 DVDD.n2798 4.5005
R4384 DVDD.n2820 DVDD.n2798 4.5005
R4385 DVDD.n2827 DVDD.n2798 4.5005
R4386 DVDD.n2819 DVDD.n2798 4.5005
R4387 DVDD.n2829 DVDD.n2798 4.5005
R4388 DVDD.n2818 DVDD.n2798 4.5005
R4389 DVDD.n2830 DVDD.n2798 4.5005
R4390 DVDD.n2831 DVDD.n2798 4.5005
R4391 DVDD.n16246 DVDD.n2798 4.5005
R4392 DVDD.n16248 DVDD.n2785 4.5005
R4393 DVDD.n2824 DVDD.n2785 4.5005
R4394 DVDD.n2822 DVDD.n2785 4.5005
R4395 DVDD.n2825 DVDD.n2785 4.5005
R4396 DVDD.n2821 DVDD.n2785 4.5005
R4397 DVDD.n2826 DVDD.n2785 4.5005
R4398 DVDD.n2820 DVDD.n2785 4.5005
R4399 DVDD.n2827 DVDD.n2785 4.5005
R4400 DVDD.n2819 DVDD.n2785 4.5005
R4401 DVDD.n2829 DVDD.n2785 4.5005
R4402 DVDD.n2818 DVDD.n2785 4.5005
R4403 DVDD.n2830 DVDD.n2785 4.5005
R4404 DVDD.n2872 DVDD.n2785 4.5005
R4405 DVDD.n2831 DVDD.n2785 4.5005
R4406 DVDD.n16246 DVDD.n2785 4.5005
R4407 DVDD.n16248 DVDD.n2799 4.5005
R4408 DVDD.n2824 DVDD.n2799 4.5005
R4409 DVDD.n2822 DVDD.n2799 4.5005
R4410 DVDD.n2825 DVDD.n2799 4.5005
R4411 DVDD.n2821 DVDD.n2799 4.5005
R4412 DVDD.n2826 DVDD.n2799 4.5005
R4413 DVDD.n2820 DVDD.n2799 4.5005
R4414 DVDD.n2827 DVDD.n2799 4.5005
R4415 DVDD.n2819 DVDD.n2799 4.5005
R4416 DVDD.n2829 DVDD.n2799 4.5005
R4417 DVDD.n2818 DVDD.n2799 4.5005
R4418 DVDD.n2830 DVDD.n2799 4.5005
R4419 DVDD.n2872 DVDD.n2799 4.5005
R4420 DVDD.n2831 DVDD.n2799 4.5005
R4421 DVDD.n16246 DVDD.n2799 4.5005
R4422 DVDD.n16248 DVDD.n2784 4.5005
R4423 DVDD.n2824 DVDD.n2784 4.5005
R4424 DVDD.n2822 DVDD.n2784 4.5005
R4425 DVDD.n2825 DVDD.n2784 4.5005
R4426 DVDD.n2821 DVDD.n2784 4.5005
R4427 DVDD.n2826 DVDD.n2784 4.5005
R4428 DVDD.n2820 DVDD.n2784 4.5005
R4429 DVDD.n2827 DVDD.n2784 4.5005
R4430 DVDD.n2819 DVDD.n2784 4.5005
R4431 DVDD.n2829 DVDD.n2784 4.5005
R4432 DVDD.n2818 DVDD.n2784 4.5005
R4433 DVDD.n2830 DVDD.n2784 4.5005
R4434 DVDD.n2831 DVDD.n2784 4.5005
R4435 DVDD.n16246 DVDD.n2784 4.5005
R4436 DVDD.n16248 DVDD.n2800 4.5005
R4437 DVDD.n2824 DVDD.n2800 4.5005
R4438 DVDD.n2822 DVDD.n2800 4.5005
R4439 DVDD.n2825 DVDD.n2800 4.5005
R4440 DVDD.n2821 DVDD.n2800 4.5005
R4441 DVDD.n2826 DVDD.n2800 4.5005
R4442 DVDD.n2820 DVDD.n2800 4.5005
R4443 DVDD.n2827 DVDD.n2800 4.5005
R4444 DVDD.n2819 DVDD.n2800 4.5005
R4445 DVDD.n2829 DVDD.n2800 4.5005
R4446 DVDD.n2818 DVDD.n2800 4.5005
R4447 DVDD.n2830 DVDD.n2800 4.5005
R4448 DVDD.n2831 DVDD.n2800 4.5005
R4449 DVDD.n16246 DVDD.n2800 4.5005
R4450 DVDD.n16248 DVDD.n2783 4.5005
R4451 DVDD.n2824 DVDD.n2783 4.5005
R4452 DVDD.n2822 DVDD.n2783 4.5005
R4453 DVDD.n2825 DVDD.n2783 4.5005
R4454 DVDD.n2821 DVDD.n2783 4.5005
R4455 DVDD.n2826 DVDD.n2783 4.5005
R4456 DVDD.n2820 DVDD.n2783 4.5005
R4457 DVDD.n2827 DVDD.n2783 4.5005
R4458 DVDD.n2819 DVDD.n2783 4.5005
R4459 DVDD.n2829 DVDD.n2783 4.5005
R4460 DVDD.n2818 DVDD.n2783 4.5005
R4461 DVDD.n2830 DVDD.n2783 4.5005
R4462 DVDD.n2831 DVDD.n2783 4.5005
R4463 DVDD.n16246 DVDD.n2783 4.5005
R4464 DVDD.n16248 DVDD.n2801 4.5005
R4465 DVDD.n2824 DVDD.n2801 4.5005
R4466 DVDD.n2822 DVDD.n2801 4.5005
R4467 DVDD.n2825 DVDD.n2801 4.5005
R4468 DVDD.n2821 DVDD.n2801 4.5005
R4469 DVDD.n2826 DVDD.n2801 4.5005
R4470 DVDD.n2820 DVDD.n2801 4.5005
R4471 DVDD.n2827 DVDD.n2801 4.5005
R4472 DVDD.n2819 DVDD.n2801 4.5005
R4473 DVDD.n2829 DVDD.n2801 4.5005
R4474 DVDD.n2818 DVDD.n2801 4.5005
R4475 DVDD.n2830 DVDD.n2801 4.5005
R4476 DVDD.n2831 DVDD.n2801 4.5005
R4477 DVDD.n16246 DVDD.n2801 4.5005
R4478 DVDD.n16248 DVDD.n2782 4.5005
R4479 DVDD.n2824 DVDD.n2782 4.5005
R4480 DVDD.n2822 DVDD.n2782 4.5005
R4481 DVDD.n2825 DVDD.n2782 4.5005
R4482 DVDD.n2821 DVDD.n2782 4.5005
R4483 DVDD.n2826 DVDD.n2782 4.5005
R4484 DVDD.n2820 DVDD.n2782 4.5005
R4485 DVDD.n2827 DVDD.n2782 4.5005
R4486 DVDD.n2819 DVDD.n2782 4.5005
R4487 DVDD.n2829 DVDD.n2782 4.5005
R4488 DVDD.n2818 DVDD.n2782 4.5005
R4489 DVDD.n2830 DVDD.n2782 4.5005
R4490 DVDD.n2831 DVDD.n2782 4.5005
R4491 DVDD.n16246 DVDD.n2782 4.5005
R4492 DVDD.n16248 DVDD.n2802 4.5005
R4493 DVDD.n2824 DVDD.n2802 4.5005
R4494 DVDD.n2822 DVDD.n2802 4.5005
R4495 DVDD.n2825 DVDD.n2802 4.5005
R4496 DVDD.n2821 DVDD.n2802 4.5005
R4497 DVDD.n2826 DVDD.n2802 4.5005
R4498 DVDD.n2820 DVDD.n2802 4.5005
R4499 DVDD.n2827 DVDD.n2802 4.5005
R4500 DVDD.n2819 DVDD.n2802 4.5005
R4501 DVDD.n2829 DVDD.n2802 4.5005
R4502 DVDD.n2818 DVDD.n2802 4.5005
R4503 DVDD.n2830 DVDD.n2802 4.5005
R4504 DVDD.n2831 DVDD.n2802 4.5005
R4505 DVDD.n16246 DVDD.n2802 4.5005
R4506 DVDD.n16248 DVDD.n2781 4.5005
R4507 DVDD.n2824 DVDD.n2781 4.5005
R4508 DVDD.n2822 DVDD.n2781 4.5005
R4509 DVDD.n2825 DVDD.n2781 4.5005
R4510 DVDD.n2821 DVDD.n2781 4.5005
R4511 DVDD.n2826 DVDD.n2781 4.5005
R4512 DVDD.n2820 DVDD.n2781 4.5005
R4513 DVDD.n2827 DVDD.n2781 4.5005
R4514 DVDD.n2819 DVDD.n2781 4.5005
R4515 DVDD.n2829 DVDD.n2781 4.5005
R4516 DVDD.n2818 DVDD.n2781 4.5005
R4517 DVDD.n2830 DVDD.n2781 4.5005
R4518 DVDD.n2872 DVDD.n2781 4.5005
R4519 DVDD.n2831 DVDD.n2781 4.5005
R4520 DVDD.n16246 DVDD.n2781 4.5005
R4521 DVDD.n16248 DVDD.n2803 4.5005
R4522 DVDD.n2824 DVDD.n2803 4.5005
R4523 DVDD.n2822 DVDD.n2803 4.5005
R4524 DVDD.n2825 DVDD.n2803 4.5005
R4525 DVDD.n2821 DVDD.n2803 4.5005
R4526 DVDD.n2826 DVDD.n2803 4.5005
R4527 DVDD.n2820 DVDD.n2803 4.5005
R4528 DVDD.n2827 DVDD.n2803 4.5005
R4529 DVDD.n2819 DVDD.n2803 4.5005
R4530 DVDD.n2829 DVDD.n2803 4.5005
R4531 DVDD.n2818 DVDD.n2803 4.5005
R4532 DVDD.n2830 DVDD.n2803 4.5005
R4533 DVDD.n2872 DVDD.n2803 4.5005
R4534 DVDD.n2831 DVDD.n2803 4.5005
R4535 DVDD.n16246 DVDD.n2803 4.5005
R4536 DVDD.n16248 DVDD.n2780 4.5005
R4537 DVDD.n2824 DVDD.n2780 4.5005
R4538 DVDD.n2822 DVDD.n2780 4.5005
R4539 DVDD.n2825 DVDD.n2780 4.5005
R4540 DVDD.n2821 DVDD.n2780 4.5005
R4541 DVDD.n2826 DVDD.n2780 4.5005
R4542 DVDD.n2820 DVDD.n2780 4.5005
R4543 DVDD.n2827 DVDD.n2780 4.5005
R4544 DVDD.n2819 DVDD.n2780 4.5005
R4545 DVDD.n2829 DVDD.n2780 4.5005
R4546 DVDD.n2818 DVDD.n2780 4.5005
R4547 DVDD.n2830 DVDD.n2780 4.5005
R4548 DVDD.n2831 DVDD.n2780 4.5005
R4549 DVDD.n16246 DVDD.n2780 4.5005
R4550 DVDD.n16248 DVDD.n16247 4.5005
R4551 DVDD.n16247 DVDD.n2824 4.5005
R4552 DVDD.n16247 DVDD.n2822 4.5005
R4553 DVDD.n16247 DVDD.n2825 4.5005
R4554 DVDD.n16247 DVDD.n2821 4.5005
R4555 DVDD.n16247 DVDD.n2826 4.5005
R4556 DVDD.n16247 DVDD.n2820 4.5005
R4557 DVDD.n16247 DVDD.n2827 4.5005
R4558 DVDD.n16247 DVDD.n2819 4.5005
R4559 DVDD.n16247 DVDD.n2829 4.5005
R4560 DVDD.n16247 DVDD.n2818 4.5005
R4561 DVDD.n16247 DVDD.n2830 4.5005
R4562 DVDD.n16247 DVDD.n2831 4.5005
R4563 DVDD.n16247 DVDD.n2816 4.5005
R4564 DVDD.n16247 DVDD.n16246 4.5005
R4565 DVDD.n2619 DVDD.n2583 4.5005
R4566 DVDD.n2623 DVDD.n2583 4.5005
R4567 DVDD.n2617 DVDD.n2583 4.5005
R4568 DVDD.n2624 DVDD.n2583 4.5005
R4569 DVDD.n2616 DVDD.n2583 4.5005
R4570 DVDD.n2625 DVDD.n2583 4.5005
R4571 DVDD.n2615 DVDD.n2583 4.5005
R4572 DVDD.n2628 DVDD.n2583 4.5005
R4573 DVDD.n2613 DVDD.n2583 4.5005
R4574 DVDD.n16312 DVDD.n2583 4.5005
R4575 DVDD.n16314 DVDD.n2583 4.5005
R4576 DVDD.n2619 DVDD.n2584 4.5005
R4577 DVDD.n2622 DVDD.n2584 4.5005
R4578 DVDD.n2618 DVDD.n2584 4.5005
R4579 DVDD.n2623 DVDD.n2584 4.5005
R4580 DVDD.n2617 DVDD.n2584 4.5005
R4581 DVDD.n2624 DVDD.n2584 4.5005
R4582 DVDD.n2616 DVDD.n2584 4.5005
R4583 DVDD.n2625 DVDD.n2584 4.5005
R4584 DVDD.n2615 DVDD.n2584 4.5005
R4585 DVDD.n2627 DVDD.n2584 4.5005
R4586 DVDD.n2614 DVDD.n2584 4.5005
R4587 DVDD.n2628 DVDD.n2584 4.5005
R4588 DVDD.n16312 DVDD.n2584 4.5005
R4589 DVDD.n16314 DVDD.n2584 4.5005
R4590 DVDD.n2619 DVDD.n2582 4.5005
R4591 DVDD.n2622 DVDD.n2582 4.5005
R4592 DVDD.n2618 DVDD.n2582 4.5005
R4593 DVDD.n2623 DVDD.n2582 4.5005
R4594 DVDD.n2617 DVDD.n2582 4.5005
R4595 DVDD.n2624 DVDD.n2582 4.5005
R4596 DVDD.n2616 DVDD.n2582 4.5005
R4597 DVDD.n2625 DVDD.n2582 4.5005
R4598 DVDD.n2615 DVDD.n2582 4.5005
R4599 DVDD.n2627 DVDD.n2582 4.5005
R4600 DVDD.n2614 DVDD.n2582 4.5005
R4601 DVDD.n2628 DVDD.n2582 4.5005
R4602 DVDD.n16312 DVDD.n2582 4.5005
R4603 DVDD.n2606 DVDD.n2582 4.5005
R4604 DVDD.n16314 DVDD.n2582 4.5005
R4605 DVDD.n2619 DVDD.n2585 4.5005
R4606 DVDD.n2622 DVDD.n2585 4.5005
R4607 DVDD.n2618 DVDD.n2585 4.5005
R4608 DVDD.n2623 DVDD.n2585 4.5005
R4609 DVDD.n2617 DVDD.n2585 4.5005
R4610 DVDD.n2624 DVDD.n2585 4.5005
R4611 DVDD.n2616 DVDD.n2585 4.5005
R4612 DVDD.n2625 DVDD.n2585 4.5005
R4613 DVDD.n2615 DVDD.n2585 4.5005
R4614 DVDD.n2627 DVDD.n2585 4.5005
R4615 DVDD.n2614 DVDD.n2585 4.5005
R4616 DVDD.n2628 DVDD.n2585 4.5005
R4617 DVDD.n2613 DVDD.n2585 4.5005
R4618 DVDD.n16312 DVDD.n2585 4.5005
R4619 DVDD.n16314 DVDD.n2585 4.5005
R4620 DVDD.n2619 DVDD.n2581 4.5005
R4621 DVDD.n2622 DVDD.n2581 4.5005
R4622 DVDD.n2618 DVDD.n2581 4.5005
R4623 DVDD.n2623 DVDD.n2581 4.5005
R4624 DVDD.n2617 DVDD.n2581 4.5005
R4625 DVDD.n2624 DVDD.n2581 4.5005
R4626 DVDD.n2616 DVDD.n2581 4.5005
R4627 DVDD.n2625 DVDD.n2581 4.5005
R4628 DVDD.n2615 DVDD.n2581 4.5005
R4629 DVDD.n2627 DVDD.n2581 4.5005
R4630 DVDD.n2614 DVDD.n2581 4.5005
R4631 DVDD.n2628 DVDD.n2581 4.5005
R4632 DVDD.n16312 DVDD.n2581 4.5005
R4633 DVDD.n16314 DVDD.n2581 4.5005
R4634 DVDD.n2619 DVDD.n2586 4.5005
R4635 DVDD.n2622 DVDD.n2586 4.5005
R4636 DVDD.n2618 DVDD.n2586 4.5005
R4637 DVDD.n2623 DVDD.n2586 4.5005
R4638 DVDD.n2617 DVDD.n2586 4.5005
R4639 DVDD.n2624 DVDD.n2586 4.5005
R4640 DVDD.n2616 DVDD.n2586 4.5005
R4641 DVDD.n2625 DVDD.n2586 4.5005
R4642 DVDD.n2615 DVDD.n2586 4.5005
R4643 DVDD.n2627 DVDD.n2586 4.5005
R4644 DVDD.n2614 DVDD.n2586 4.5005
R4645 DVDD.n2628 DVDD.n2586 4.5005
R4646 DVDD.n16312 DVDD.n2586 4.5005
R4647 DVDD.n16314 DVDD.n2586 4.5005
R4648 DVDD.n2619 DVDD.n2580 4.5005
R4649 DVDD.n2622 DVDD.n2580 4.5005
R4650 DVDD.n2618 DVDD.n2580 4.5005
R4651 DVDD.n2623 DVDD.n2580 4.5005
R4652 DVDD.n2617 DVDD.n2580 4.5005
R4653 DVDD.n2624 DVDD.n2580 4.5005
R4654 DVDD.n2616 DVDD.n2580 4.5005
R4655 DVDD.n2625 DVDD.n2580 4.5005
R4656 DVDD.n2615 DVDD.n2580 4.5005
R4657 DVDD.n2627 DVDD.n2580 4.5005
R4658 DVDD.n2614 DVDD.n2580 4.5005
R4659 DVDD.n2628 DVDD.n2580 4.5005
R4660 DVDD.n2613 DVDD.n2580 4.5005
R4661 DVDD.n16312 DVDD.n2580 4.5005
R4662 DVDD.n16314 DVDD.n2580 4.5005
R4663 DVDD.n2619 DVDD.n2587 4.5005
R4664 DVDD.n2622 DVDD.n2587 4.5005
R4665 DVDD.n2618 DVDD.n2587 4.5005
R4666 DVDD.n2623 DVDD.n2587 4.5005
R4667 DVDD.n2617 DVDD.n2587 4.5005
R4668 DVDD.n2624 DVDD.n2587 4.5005
R4669 DVDD.n2616 DVDD.n2587 4.5005
R4670 DVDD.n2625 DVDD.n2587 4.5005
R4671 DVDD.n2615 DVDD.n2587 4.5005
R4672 DVDD.n2627 DVDD.n2587 4.5005
R4673 DVDD.n2614 DVDD.n2587 4.5005
R4674 DVDD.n2628 DVDD.n2587 4.5005
R4675 DVDD.n2613 DVDD.n2587 4.5005
R4676 DVDD.n16312 DVDD.n2587 4.5005
R4677 DVDD.n16314 DVDD.n2587 4.5005
R4678 DVDD.n2619 DVDD.n2579 4.5005
R4679 DVDD.n2622 DVDD.n2579 4.5005
R4680 DVDD.n2618 DVDD.n2579 4.5005
R4681 DVDD.n2623 DVDD.n2579 4.5005
R4682 DVDD.n2617 DVDD.n2579 4.5005
R4683 DVDD.n2624 DVDD.n2579 4.5005
R4684 DVDD.n2616 DVDD.n2579 4.5005
R4685 DVDD.n2625 DVDD.n2579 4.5005
R4686 DVDD.n2615 DVDD.n2579 4.5005
R4687 DVDD.n2627 DVDD.n2579 4.5005
R4688 DVDD.n2614 DVDD.n2579 4.5005
R4689 DVDD.n2628 DVDD.n2579 4.5005
R4690 DVDD.n16312 DVDD.n2579 4.5005
R4691 DVDD.n16314 DVDD.n2579 4.5005
R4692 DVDD.n2619 DVDD.n2588 4.5005
R4693 DVDD.n2622 DVDD.n2588 4.5005
R4694 DVDD.n2618 DVDD.n2588 4.5005
R4695 DVDD.n2623 DVDD.n2588 4.5005
R4696 DVDD.n2617 DVDD.n2588 4.5005
R4697 DVDD.n2624 DVDD.n2588 4.5005
R4698 DVDD.n2616 DVDD.n2588 4.5005
R4699 DVDD.n2625 DVDD.n2588 4.5005
R4700 DVDD.n2615 DVDD.n2588 4.5005
R4701 DVDD.n2627 DVDD.n2588 4.5005
R4702 DVDD.n2614 DVDD.n2588 4.5005
R4703 DVDD.n2628 DVDD.n2588 4.5005
R4704 DVDD.n16312 DVDD.n2588 4.5005
R4705 DVDD.n16314 DVDD.n2588 4.5005
R4706 DVDD.n2619 DVDD.n2578 4.5005
R4707 DVDD.n2622 DVDD.n2578 4.5005
R4708 DVDD.n2618 DVDD.n2578 4.5005
R4709 DVDD.n2623 DVDD.n2578 4.5005
R4710 DVDD.n2617 DVDD.n2578 4.5005
R4711 DVDD.n2624 DVDD.n2578 4.5005
R4712 DVDD.n2616 DVDD.n2578 4.5005
R4713 DVDD.n2625 DVDD.n2578 4.5005
R4714 DVDD.n2615 DVDD.n2578 4.5005
R4715 DVDD.n2627 DVDD.n2578 4.5005
R4716 DVDD.n2614 DVDD.n2578 4.5005
R4717 DVDD.n2628 DVDD.n2578 4.5005
R4718 DVDD.n2613 DVDD.n2578 4.5005
R4719 DVDD.n16312 DVDD.n2578 4.5005
R4720 DVDD.n16314 DVDD.n2578 4.5005
R4721 DVDD.n2619 DVDD.n2589 4.5005
R4722 DVDD.n2622 DVDD.n2589 4.5005
R4723 DVDD.n2618 DVDD.n2589 4.5005
R4724 DVDD.n2623 DVDD.n2589 4.5005
R4725 DVDD.n2617 DVDD.n2589 4.5005
R4726 DVDD.n2624 DVDD.n2589 4.5005
R4727 DVDD.n2616 DVDD.n2589 4.5005
R4728 DVDD.n2625 DVDD.n2589 4.5005
R4729 DVDD.n2615 DVDD.n2589 4.5005
R4730 DVDD.n2627 DVDD.n2589 4.5005
R4731 DVDD.n2614 DVDD.n2589 4.5005
R4732 DVDD.n2628 DVDD.n2589 4.5005
R4733 DVDD.n2613 DVDD.n2589 4.5005
R4734 DVDD.n16312 DVDD.n2589 4.5005
R4735 DVDD.n16314 DVDD.n2589 4.5005
R4736 DVDD.n2619 DVDD.n2577 4.5005
R4737 DVDD.n2622 DVDD.n2577 4.5005
R4738 DVDD.n2618 DVDD.n2577 4.5005
R4739 DVDD.n2623 DVDD.n2577 4.5005
R4740 DVDD.n2617 DVDD.n2577 4.5005
R4741 DVDD.n2624 DVDD.n2577 4.5005
R4742 DVDD.n2616 DVDD.n2577 4.5005
R4743 DVDD.n2625 DVDD.n2577 4.5005
R4744 DVDD.n2615 DVDD.n2577 4.5005
R4745 DVDD.n2627 DVDD.n2577 4.5005
R4746 DVDD.n2614 DVDD.n2577 4.5005
R4747 DVDD.n2628 DVDD.n2577 4.5005
R4748 DVDD.n16312 DVDD.n2577 4.5005
R4749 DVDD.n16314 DVDD.n2577 4.5005
R4750 DVDD.n2619 DVDD.n2590 4.5005
R4751 DVDD.n2622 DVDD.n2590 4.5005
R4752 DVDD.n2618 DVDD.n2590 4.5005
R4753 DVDD.n2623 DVDD.n2590 4.5005
R4754 DVDD.n2617 DVDD.n2590 4.5005
R4755 DVDD.n2624 DVDD.n2590 4.5005
R4756 DVDD.n2616 DVDD.n2590 4.5005
R4757 DVDD.n2625 DVDD.n2590 4.5005
R4758 DVDD.n2615 DVDD.n2590 4.5005
R4759 DVDD.n2627 DVDD.n2590 4.5005
R4760 DVDD.n2614 DVDD.n2590 4.5005
R4761 DVDD.n2628 DVDD.n2590 4.5005
R4762 DVDD.n16312 DVDD.n2590 4.5005
R4763 DVDD.n16314 DVDD.n2590 4.5005
R4764 DVDD.n2619 DVDD.n2576 4.5005
R4765 DVDD.n2622 DVDD.n2576 4.5005
R4766 DVDD.n2618 DVDD.n2576 4.5005
R4767 DVDD.n2623 DVDD.n2576 4.5005
R4768 DVDD.n2617 DVDD.n2576 4.5005
R4769 DVDD.n2624 DVDD.n2576 4.5005
R4770 DVDD.n2616 DVDD.n2576 4.5005
R4771 DVDD.n2625 DVDD.n2576 4.5005
R4772 DVDD.n2615 DVDD.n2576 4.5005
R4773 DVDD.n2627 DVDD.n2576 4.5005
R4774 DVDD.n2614 DVDD.n2576 4.5005
R4775 DVDD.n2628 DVDD.n2576 4.5005
R4776 DVDD.n2613 DVDD.n2576 4.5005
R4777 DVDD.n16312 DVDD.n2576 4.5005
R4778 DVDD.n16314 DVDD.n2576 4.5005
R4779 DVDD.n2619 DVDD.n2591 4.5005
R4780 DVDD.n2622 DVDD.n2591 4.5005
R4781 DVDD.n2618 DVDD.n2591 4.5005
R4782 DVDD.n2623 DVDD.n2591 4.5005
R4783 DVDD.n2617 DVDD.n2591 4.5005
R4784 DVDD.n2624 DVDD.n2591 4.5005
R4785 DVDD.n2616 DVDD.n2591 4.5005
R4786 DVDD.n2625 DVDD.n2591 4.5005
R4787 DVDD.n2615 DVDD.n2591 4.5005
R4788 DVDD.n2627 DVDD.n2591 4.5005
R4789 DVDD.n2614 DVDD.n2591 4.5005
R4790 DVDD.n2628 DVDD.n2591 4.5005
R4791 DVDD.n2613 DVDD.n2591 4.5005
R4792 DVDD.n16312 DVDD.n2591 4.5005
R4793 DVDD.n16314 DVDD.n2591 4.5005
R4794 DVDD.n2619 DVDD.n2575 4.5005
R4795 DVDD.n2622 DVDD.n2575 4.5005
R4796 DVDD.n2618 DVDD.n2575 4.5005
R4797 DVDD.n2623 DVDD.n2575 4.5005
R4798 DVDD.n2617 DVDD.n2575 4.5005
R4799 DVDD.n2624 DVDD.n2575 4.5005
R4800 DVDD.n2616 DVDD.n2575 4.5005
R4801 DVDD.n2625 DVDD.n2575 4.5005
R4802 DVDD.n2615 DVDD.n2575 4.5005
R4803 DVDD.n2627 DVDD.n2575 4.5005
R4804 DVDD.n2614 DVDD.n2575 4.5005
R4805 DVDD.n2628 DVDD.n2575 4.5005
R4806 DVDD.n16312 DVDD.n2575 4.5005
R4807 DVDD.n16314 DVDD.n2575 4.5005
R4808 DVDD.n2619 DVDD.n2592 4.5005
R4809 DVDD.n2622 DVDD.n2592 4.5005
R4810 DVDD.n2618 DVDD.n2592 4.5005
R4811 DVDD.n2623 DVDD.n2592 4.5005
R4812 DVDD.n2617 DVDD.n2592 4.5005
R4813 DVDD.n2624 DVDD.n2592 4.5005
R4814 DVDD.n2616 DVDD.n2592 4.5005
R4815 DVDD.n2625 DVDD.n2592 4.5005
R4816 DVDD.n2615 DVDD.n2592 4.5005
R4817 DVDD.n2627 DVDD.n2592 4.5005
R4818 DVDD.n2614 DVDD.n2592 4.5005
R4819 DVDD.n2628 DVDD.n2592 4.5005
R4820 DVDD.n16312 DVDD.n2592 4.5005
R4821 DVDD.n16314 DVDD.n2592 4.5005
R4822 DVDD.n2619 DVDD.n2574 4.5005
R4823 DVDD.n2622 DVDD.n2574 4.5005
R4824 DVDD.n2618 DVDD.n2574 4.5005
R4825 DVDD.n2623 DVDD.n2574 4.5005
R4826 DVDD.n2617 DVDD.n2574 4.5005
R4827 DVDD.n2624 DVDD.n2574 4.5005
R4828 DVDD.n2616 DVDD.n2574 4.5005
R4829 DVDD.n2625 DVDD.n2574 4.5005
R4830 DVDD.n2615 DVDD.n2574 4.5005
R4831 DVDD.n2627 DVDD.n2574 4.5005
R4832 DVDD.n2614 DVDD.n2574 4.5005
R4833 DVDD.n2628 DVDD.n2574 4.5005
R4834 DVDD.n2613 DVDD.n2574 4.5005
R4835 DVDD.n16312 DVDD.n2574 4.5005
R4836 DVDD.n16314 DVDD.n2574 4.5005
R4837 DVDD.n2619 DVDD.n2593 4.5005
R4838 DVDD.n2622 DVDD.n2593 4.5005
R4839 DVDD.n2618 DVDD.n2593 4.5005
R4840 DVDD.n2623 DVDD.n2593 4.5005
R4841 DVDD.n2617 DVDD.n2593 4.5005
R4842 DVDD.n2624 DVDD.n2593 4.5005
R4843 DVDD.n2616 DVDD.n2593 4.5005
R4844 DVDD.n2625 DVDD.n2593 4.5005
R4845 DVDD.n2615 DVDD.n2593 4.5005
R4846 DVDD.n2627 DVDD.n2593 4.5005
R4847 DVDD.n2614 DVDD.n2593 4.5005
R4848 DVDD.n2628 DVDD.n2593 4.5005
R4849 DVDD.n2613 DVDD.n2593 4.5005
R4850 DVDD.n16312 DVDD.n2593 4.5005
R4851 DVDD.n16314 DVDD.n2593 4.5005
R4852 DVDD.n2619 DVDD.n2573 4.5005
R4853 DVDD.n2622 DVDD.n2573 4.5005
R4854 DVDD.n2618 DVDD.n2573 4.5005
R4855 DVDD.n2623 DVDD.n2573 4.5005
R4856 DVDD.n2617 DVDD.n2573 4.5005
R4857 DVDD.n2624 DVDD.n2573 4.5005
R4858 DVDD.n2616 DVDD.n2573 4.5005
R4859 DVDD.n2625 DVDD.n2573 4.5005
R4860 DVDD.n2615 DVDD.n2573 4.5005
R4861 DVDD.n2627 DVDD.n2573 4.5005
R4862 DVDD.n2614 DVDD.n2573 4.5005
R4863 DVDD.n2628 DVDD.n2573 4.5005
R4864 DVDD.n16312 DVDD.n2573 4.5005
R4865 DVDD.n16314 DVDD.n2573 4.5005
R4866 DVDD.n2619 DVDD.n2594 4.5005
R4867 DVDD.n2622 DVDD.n2594 4.5005
R4868 DVDD.n2618 DVDD.n2594 4.5005
R4869 DVDD.n2623 DVDD.n2594 4.5005
R4870 DVDD.n2617 DVDD.n2594 4.5005
R4871 DVDD.n2624 DVDD.n2594 4.5005
R4872 DVDD.n2616 DVDD.n2594 4.5005
R4873 DVDD.n2625 DVDD.n2594 4.5005
R4874 DVDD.n2615 DVDD.n2594 4.5005
R4875 DVDD.n2627 DVDD.n2594 4.5005
R4876 DVDD.n2614 DVDD.n2594 4.5005
R4877 DVDD.n2628 DVDD.n2594 4.5005
R4878 DVDD.n16312 DVDD.n2594 4.5005
R4879 DVDD.n16314 DVDD.n2594 4.5005
R4880 DVDD.n2619 DVDD.n2572 4.5005
R4881 DVDD.n2622 DVDD.n2572 4.5005
R4882 DVDD.n2618 DVDD.n2572 4.5005
R4883 DVDD.n2623 DVDD.n2572 4.5005
R4884 DVDD.n2617 DVDD.n2572 4.5005
R4885 DVDD.n2624 DVDD.n2572 4.5005
R4886 DVDD.n2616 DVDD.n2572 4.5005
R4887 DVDD.n2625 DVDD.n2572 4.5005
R4888 DVDD.n2615 DVDD.n2572 4.5005
R4889 DVDD.n2627 DVDD.n2572 4.5005
R4890 DVDD.n2614 DVDD.n2572 4.5005
R4891 DVDD.n2628 DVDD.n2572 4.5005
R4892 DVDD.n2613 DVDD.n2572 4.5005
R4893 DVDD.n16312 DVDD.n2572 4.5005
R4894 DVDD.n16314 DVDD.n2572 4.5005
R4895 DVDD.n16313 DVDD.n2619 4.5005
R4896 DVDD.n16313 DVDD.n2622 4.5005
R4897 DVDD.n16313 DVDD.n2618 4.5005
R4898 DVDD.n16313 DVDD.n2623 4.5005
R4899 DVDD.n16313 DVDD.n2617 4.5005
R4900 DVDD.n16313 DVDD.n2624 4.5005
R4901 DVDD.n16313 DVDD.n2616 4.5005
R4902 DVDD.n16313 DVDD.n2625 4.5005
R4903 DVDD.n16313 DVDD.n2615 4.5005
R4904 DVDD.n16313 DVDD.n2627 4.5005
R4905 DVDD.n16313 DVDD.n2614 4.5005
R4906 DVDD.n16313 DVDD.n2628 4.5005
R4907 DVDD.n16313 DVDD.n2613 4.5005
R4908 DVDD.n16313 DVDD.n16312 4.5005
R4909 DVDD.n16313 DVDD.n2606 4.5005
R4910 DVDD.n16314 DVDD.n16313 4.5005
R4911 DVDD.n2485 DVDD.n2385 4.5005
R4912 DVDD.n2485 DVDD.n2477 4.5005
R4913 DVDD.n2485 DVDD.n2436 4.5005
R4914 DVDD.n2485 DVDD.n2478 4.5005
R4915 DVDD.n2485 DVDD.n2435 4.5005
R4916 DVDD.n2485 DVDD.n2479 4.5005
R4917 DVDD.n2485 DVDD.n2434 4.5005
R4918 DVDD.n2485 DVDD.n2481 4.5005
R4919 DVDD.n2485 DVDD.n2432 4.5005
R4920 DVDD.n2485 DVDD.n2482 4.5005
R4921 DVDD.n2485 DVDD.n2424 4.5005
R4922 DVDD.n16368 DVDD.n2485 4.5005
R4923 DVDD.n2402 DVDD.n2385 4.5005
R4924 DVDD.n16370 DVDD.n2402 4.5005
R4925 DVDD.n2437 DVDD.n2402 4.5005
R4926 DVDD.n2477 DVDD.n2402 4.5005
R4927 DVDD.n2436 DVDD.n2402 4.5005
R4928 DVDD.n2478 DVDD.n2402 4.5005
R4929 DVDD.n2435 DVDD.n2402 4.5005
R4930 DVDD.n2479 DVDD.n2402 4.5005
R4931 DVDD.n2434 DVDD.n2402 4.5005
R4932 DVDD.n2480 DVDD.n2402 4.5005
R4933 DVDD.n2433 DVDD.n2402 4.5005
R4934 DVDD.n2481 DVDD.n2402 4.5005
R4935 DVDD.n2432 DVDD.n2402 4.5005
R4936 DVDD.n2482 DVDD.n2402 4.5005
R4937 DVDD.n16368 DVDD.n2402 4.5005
R4938 DVDD.n2400 DVDD.n2385 4.5005
R4939 DVDD.n16370 DVDD.n2400 4.5005
R4940 DVDD.n2437 DVDD.n2400 4.5005
R4941 DVDD.n2477 DVDD.n2400 4.5005
R4942 DVDD.n2436 DVDD.n2400 4.5005
R4943 DVDD.n2478 DVDD.n2400 4.5005
R4944 DVDD.n2435 DVDD.n2400 4.5005
R4945 DVDD.n2479 DVDD.n2400 4.5005
R4946 DVDD.n2434 DVDD.n2400 4.5005
R4947 DVDD.n2480 DVDD.n2400 4.5005
R4948 DVDD.n2433 DVDD.n2400 4.5005
R4949 DVDD.n2481 DVDD.n2400 4.5005
R4950 DVDD.n2482 DVDD.n2400 4.5005
R4951 DVDD.n16368 DVDD.n2400 4.5005
R4952 DVDD.n2403 DVDD.n2385 4.5005
R4953 DVDD.n16370 DVDD.n2403 4.5005
R4954 DVDD.n2437 DVDD.n2403 4.5005
R4955 DVDD.n2477 DVDD.n2403 4.5005
R4956 DVDD.n2436 DVDD.n2403 4.5005
R4957 DVDD.n2478 DVDD.n2403 4.5005
R4958 DVDD.n2435 DVDD.n2403 4.5005
R4959 DVDD.n2479 DVDD.n2403 4.5005
R4960 DVDD.n2434 DVDD.n2403 4.5005
R4961 DVDD.n2480 DVDD.n2403 4.5005
R4962 DVDD.n2433 DVDD.n2403 4.5005
R4963 DVDD.n2481 DVDD.n2403 4.5005
R4964 DVDD.n2482 DVDD.n2403 4.5005
R4965 DVDD.n16368 DVDD.n2403 4.5005
R4966 DVDD.n2399 DVDD.n2385 4.5005
R4967 DVDD.n16370 DVDD.n2399 4.5005
R4968 DVDD.n2437 DVDD.n2399 4.5005
R4969 DVDD.n2477 DVDD.n2399 4.5005
R4970 DVDD.n2436 DVDD.n2399 4.5005
R4971 DVDD.n2478 DVDD.n2399 4.5005
R4972 DVDD.n2435 DVDD.n2399 4.5005
R4973 DVDD.n2479 DVDD.n2399 4.5005
R4974 DVDD.n2434 DVDD.n2399 4.5005
R4975 DVDD.n2480 DVDD.n2399 4.5005
R4976 DVDD.n2433 DVDD.n2399 4.5005
R4977 DVDD.n2481 DVDD.n2399 4.5005
R4978 DVDD.n2432 DVDD.n2399 4.5005
R4979 DVDD.n2482 DVDD.n2399 4.5005
R4980 DVDD.n16368 DVDD.n2399 4.5005
R4981 DVDD.n2404 DVDD.n2385 4.5005
R4982 DVDD.n16370 DVDD.n2404 4.5005
R4983 DVDD.n2437 DVDD.n2404 4.5005
R4984 DVDD.n2477 DVDD.n2404 4.5005
R4985 DVDD.n2436 DVDD.n2404 4.5005
R4986 DVDD.n2478 DVDD.n2404 4.5005
R4987 DVDD.n2435 DVDD.n2404 4.5005
R4988 DVDD.n2479 DVDD.n2404 4.5005
R4989 DVDD.n2434 DVDD.n2404 4.5005
R4990 DVDD.n2480 DVDD.n2404 4.5005
R4991 DVDD.n2433 DVDD.n2404 4.5005
R4992 DVDD.n2481 DVDD.n2404 4.5005
R4993 DVDD.n2432 DVDD.n2404 4.5005
R4994 DVDD.n2482 DVDD.n2404 4.5005
R4995 DVDD.n16368 DVDD.n2404 4.5005
R4996 DVDD.n2398 DVDD.n2385 4.5005
R4997 DVDD.n16370 DVDD.n2398 4.5005
R4998 DVDD.n2437 DVDD.n2398 4.5005
R4999 DVDD.n2477 DVDD.n2398 4.5005
R5000 DVDD.n2436 DVDD.n2398 4.5005
R5001 DVDD.n2478 DVDD.n2398 4.5005
R5002 DVDD.n2435 DVDD.n2398 4.5005
R5003 DVDD.n2479 DVDD.n2398 4.5005
R5004 DVDD.n2434 DVDD.n2398 4.5005
R5005 DVDD.n2480 DVDD.n2398 4.5005
R5006 DVDD.n2433 DVDD.n2398 4.5005
R5007 DVDD.n2481 DVDD.n2398 4.5005
R5008 DVDD.n2482 DVDD.n2398 4.5005
R5009 DVDD.n16368 DVDD.n2398 4.5005
R5010 DVDD.n2405 DVDD.n2385 4.5005
R5011 DVDD.n16370 DVDD.n2405 4.5005
R5012 DVDD.n2437 DVDD.n2405 4.5005
R5013 DVDD.n2477 DVDD.n2405 4.5005
R5014 DVDD.n2436 DVDD.n2405 4.5005
R5015 DVDD.n2478 DVDD.n2405 4.5005
R5016 DVDD.n2435 DVDD.n2405 4.5005
R5017 DVDD.n2479 DVDD.n2405 4.5005
R5018 DVDD.n2434 DVDD.n2405 4.5005
R5019 DVDD.n2480 DVDD.n2405 4.5005
R5020 DVDD.n2433 DVDD.n2405 4.5005
R5021 DVDD.n2481 DVDD.n2405 4.5005
R5022 DVDD.n2482 DVDD.n2405 4.5005
R5023 DVDD.n16368 DVDD.n2405 4.5005
R5024 DVDD.n2397 DVDD.n2385 4.5005
R5025 DVDD.n16370 DVDD.n2397 4.5005
R5026 DVDD.n2437 DVDD.n2397 4.5005
R5027 DVDD.n2477 DVDD.n2397 4.5005
R5028 DVDD.n2436 DVDD.n2397 4.5005
R5029 DVDD.n2478 DVDD.n2397 4.5005
R5030 DVDD.n2435 DVDD.n2397 4.5005
R5031 DVDD.n2479 DVDD.n2397 4.5005
R5032 DVDD.n2434 DVDD.n2397 4.5005
R5033 DVDD.n2480 DVDD.n2397 4.5005
R5034 DVDD.n2433 DVDD.n2397 4.5005
R5035 DVDD.n2481 DVDD.n2397 4.5005
R5036 DVDD.n2432 DVDD.n2397 4.5005
R5037 DVDD.n2482 DVDD.n2397 4.5005
R5038 DVDD.n16368 DVDD.n2397 4.5005
R5039 DVDD.n2406 DVDD.n2385 4.5005
R5040 DVDD.n16370 DVDD.n2406 4.5005
R5041 DVDD.n2437 DVDD.n2406 4.5005
R5042 DVDD.n2477 DVDD.n2406 4.5005
R5043 DVDD.n2436 DVDD.n2406 4.5005
R5044 DVDD.n2478 DVDD.n2406 4.5005
R5045 DVDD.n2435 DVDD.n2406 4.5005
R5046 DVDD.n2479 DVDD.n2406 4.5005
R5047 DVDD.n2434 DVDD.n2406 4.5005
R5048 DVDD.n2480 DVDD.n2406 4.5005
R5049 DVDD.n2433 DVDD.n2406 4.5005
R5050 DVDD.n2481 DVDD.n2406 4.5005
R5051 DVDD.n2432 DVDD.n2406 4.5005
R5052 DVDD.n2482 DVDD.n2406 4.5005
R5053 DVDD.n16368 DVDD.n2406 4.5005
R5054 DVDD.n2396 DVDD.n2385 4.5005
R5055 DVDD.n16370 DVDD.n2396 4.5005
R5056 DVDD.n2437 DVDD.n2396 4.5005
R5057 DVDD.n2477 DVDD.n2396 4.5005
R5058 DVDD.n2436 DVDD.n2396 4.5005
R5059 DVDD.n2478 DVDD.n2396 4.5005
R5060 DVDD.n2435 DVDD.n2396 4.5005
R5061 DVDD.n2479 DVDD.n2396 4.5005
R5062 DVDD.n2434 DVDD.n2396 4.5005
R5063 DVDD.n2480 DVDD.n2396 4.5005
R5064 DVDD.n2433 DVDD.n2396 4.5005
R5065 DVDD.n2481 DVDD.n2396 4.5005
R5066 DVDD.n2482 DVDD.n2396 4.5005
R5067 DVDD.n16368 DVDD.n2396 4.5005
R5068 DVDD.n2407 DVDD.n2385 4.5005
R5069 DVDD.n16370 DVDD.n2407 4.5005
R5070 DVDD.n2437 DVDD.n2407 4.5005
R5071 DVDD.n2477 DVDD.n2407 4.5005
R5072 DVDD.n2436 DVDD.n2407 4.5005
R5073 DVDD.n2478 DVDD.n2407 4.5005
R5074 DVDD.n2435 DVDD.n2407 4.5005
R5075 DVDD.n2479 DVDD.n2407 4.5005
R5076 DVDD.n2434 DVDD.n2407 4.5005
R5077 DVDD.n2480 DVDD.n2407 4.5005
R5078 DVDD.n2433 DVDD.n2407 4.5005
R5079 DVDD.n2481 DVDD.n2407 4.5005
R5080 DVDD.n2482 DVDD.n2407 4.5005
R5081 DVDD.n16368 DVDD.n2407 4.5005
R5082 DVDD.n2395 DVDD.n2385 4.5005
R5083 DVDD.n16370 DVDD.n2395 4.5005
R5084 DVDD.n2437 DVDD.n2395 4.5005
R5085 DVDD.n2477 DVDD.n2395 4.5005
R5086 DVDD.n2436 DVDD.n2395 4.5005
R5087 DVDD.n2478 DVDD.n2395 4.5005
R5088 DVDD.n2435 DVDD.n2395 4.5005
R5089 DVDD.n2479 DVDD.n2395 4.5005
R5090 DVDD.n2434 DVDD.n2395 4.5005
R5091 DVDD.n2480 DVDD.n2395 4.5005
R5092 DVDD.n2433 DVDD.n2395 4.5005
R5093 DVDD.n2481 DVDD.n2395 4.5005
R5094 DVDD.n2482 DVDD.n2395 4.5005
R5095 DVDD.n16368 DVDD.n2395 4.5005
R5096 DVDD.n2408 DVDD.n2385 4.5005
R5097 DVDD.n16370 DVDD.n2408 4.5005
R5098 DVDD.n2437 DVDD.n2408 4.5005
R5099 DVDD.n2477 DVDD.n2408 4.5005
R5100 DVDD.n2436 DVDD.n2408 4.5005
R5101 DVDD.n2478 DVDD.n2408 4.5005
R5102 DVDD.n2435 DVDD.n2408 4.5005
R5103 DVDD.n2479 DVDD.n2408 4.5005
R5104 DVDD.n2434 DVDD.n2408 4.5005
R5105 DVDD.n2480 DVDD.n2408 4.5005
R5106 DVDD.n2433 DVDD.n2408 4.5005
R5107 DVDD.n2481 DVDD.n2408 4.5005
R5108 DVDD.n2482 DVDD.n2408 4.5005
R5109 DVDD.n16368 DVDD.n2408 4.5005
R5110 DVDD.n2394 DVDD.n2385 4.5005
R5111 DVDD.n16370 DVDD.n2394 4.5005
R5112 DVDD.n2437 DVDD.n2394 4.5005
R5113 DVDD.n2477 DVDD.n2394 4.5005
R5114 DVDD.n2436 DVDD.n2394 4.5005
R5115 DVDD.n2478 DVDD.n2394 4.5005
R5116 DVDD.n2435 DVDD.n2394 4.5005
R5117 DVDD.n2479 DVDD.n2394 4.5005
R5118 DVDD.n2434 DVDD.n2394 4.5005
R5119 DVDD.n2480 DVDD.n2394 4.5005
R5120 DVDD.n2433 DVDD.n2394 4.5005
R5121 DVDD.n2481 DVDD.n2394 4.5005
R5122 DVDD.n2482 DVDD.n2394 4.5005
R5123 DVDD.n16368 DVDD.n2394 4.5005
R5124 DVDD.n2409 DVDD.n2385 4.5005
R5125 DVDD.n16370 DVDD.n2409 4.5005
R5126 DVDD.n2437 DVDD.n2409 4.5005
R5127 DVDD.n2477 DVDD.n2409 4.5005
R5128 DVDD.n2436 DVDD.n2409 4.5005
R5129 DVDD.n2478 DVDD.n2409 4.5005
R5130 DVDD.n2435 DVDD.n2409 4.5005
R5131 DVDD.n2479 DVDD.n2409 4.5005
R5132 DVDD.n2434 DVDD.n2409 4.5005
R5133 DVDD.n2480 DVDD.n2409 4.5005
R5134 DVDD.n2433 DVDD.n2409 4.5005
R5135 DVDD.n2481 DVDD.n2409 4.5005
R5136 DVDD.n2482 DVDD.n2409 4.5005
R5137 DVDD.n16368 DVDD.n2409 4.5005
R5138 DVDD.n2393 DVDD.n2385 4.5005
R5139 DVDD.n16370 DVDD.n2393 4.5005
R5140 DVDD.n2437 DVDD.n2393 4.5005
R5141 DVDD.n2477 DVDD.n2393 4.5005
R5142 DVDD.n2436 DVDD.n2393 4.5005
R5143 DVDD.n2478 DVDD.n2393 4.5005
R5144 DVDD.n2435 DVDD.n2393 4.5005
R5145 DVDD.n2479 DVDD.n2393 4.5005
R5146 DVDD.n2434 DVDD.n2393 4.5005
R5147 DVDD.n2480 DVDD.n2393 4.5005
R5148 DVDD.n2433 DVDD.n2393 4.5005
R5149 DVDD.n2481 DVDD.n2393 4.5005
R5150 DVDD.n2432 DVDD.n2393 4.5005
R5151 DVDD.n2482 DVDD.n2393 4.5005
R5152 DVDD.n16368 DVDD.n2393 4.5005
R5153 DVDD.n2410 DVDD.n2385 4.5005
R5154 DVDD.n16370 DVDD.n2410 4.5005
R5155 DVDD.n2437 DVDD.n2410 4.5005
R5156 DVDD.n2477 DVDD.n2410 4.5005
R5157 DVDD.n2436 DVDD.n2410 4.5005
R5158 DVDD.n2478 DVDD.n2410 4.5005
R5159 DVDD.n2435 DVDD.n2410 4.5005
R5160 DVDD.n2479 DVDD.n2410 4.5005
R5161 DVDD.n2434 DVDD.n2410 4.5005
R5162 DVDD.n2480 DVDD.n2410 4.5005
R5163 DVDD.n2433 DVDD.n2410 4.5005
R5164 DVDD.n2481 DVDD.n2410 4.5005
R5165 DVDD.n2482 DVDD.n2410 4.5005
R5166 DVDD.n16368 DVDD.n2410 4.5005
R5167 DVDD.n2392 DVDD.n2385 4.5005
R5168 DVDD.n16370 DVDD.n2392 4.5005
R5169 DVDD.n2437 DVDD.n2392 4.5005
R5170 DVDD.n2477 DVDD.n2392 4.5005
R5171 DVDD.n2436 DVDD.n2392 4.5005
R5172 DVDD.n2478 DVDD.n2392 4.5005
R5173 DVDD.n2435 DVDD.n2392 4.5005
R5174 DVDD.n2479 DVDD.n2392 4.5005
R5175 DVDD.n2434 DVDD.n2392 4.5005
R5176 DVDD.n2480 DVDD.n2392 4.5005
R5177 DVDD.n2433 DVDD.n2392 4.5005
R5178 DVDD.n2481 DVDD.n2392 4.5005
R5179 DVDD.n2482 DVDD.n2392 4.5005
R5180 DVDD.n16368 DVDD.n2392 4.5005
R5181 DVDD.n2411 DVDD.n2385 4.5005
R5182 DVDD.n16370 DVDD.n2411 4.5005
R5183 DVDD.n2437 DVDD.n2411 4.5005
R5184 DVDD.n2477 DVDD.n2411 4.5005
R5185 DVDD.n2436 DVDD.n2411 4.5005
R5186 DVDD.n2478 DVDD.n2411 4.5005
R5187 DVDD.n2435 DVDD.n2411 4.5005
R5188 DVDD.n2479 DVDD.n2411 4.5005
R5189 DVDD.n2434 DVDD.n2411 4.5005
R5190 DVDD.n2480 DVDD.n2411 4.5005
R5191 DVDD.n2433 DVDD.n2411 4.5005
R5192 DVDD.n2481 DVDD.n2411 4.5005
R5193 DVDD.n2482 DVDD.n2411 4.5005
R5194 DVDD.n16368 DVDD.n2411 4.5005
R5195 DVDD.n2391 DVDD.n2385 4.5005
R5196 DVDD.n16370 DVDD.n2391 4.5005
R5197 DVDD.n2437 DVDD.n2391 4.5005
R5198 DVDD.n2477 DVDD.n2391 4.5005
R5199 DVDD.n2436 DVDD.n2391 4.5005
R5200 DVDD.n2478 DVDD.n2391 4.5005
R5201 DVDD.n2435 DVDD.n2391 4.5005
R5202 DVDD.n2479 DVDD.n2391 4.5005
R5203 DVDD.n2434 DVDD.n2391 4.5005
R5204 DVDD.n2480 DVDD.n2391 4.5005
R5205 DVDD.n2433 DVDD.n2391 4.5005
R5206 DVDD.n2481 DVDD.n2391 4.5005
R5207 DVDD.n2432 DVDD.n2391 4.5005
R5208 DVDD.n2482 DVDD.n2391 4.5005
R5209 DVDD.n16368 DVDD.n2391 4.5005
R5210 DVDD.n4262 DVDD.n4244 4.5005
R5211 DVDD.n4262 DVDD.n4250 4.5005
R5212 DVDD.n4262 DVDD.n4241 4.5005
R5213 DVDD.n4600 DVDD.n4262 4.5005
R5214 DVDD.n4262 DVDD.n4246 4.5005
R5215 DVDD.n4597 DVDD.n4262 4.5005
R5216 DVDD.n4262 DVDD.n4248 4.5005
R5217 DVDD.n4257 DVDD.n4244 4.5005
R5218 DVDD.n4257 DVDD.n4249 4.5005
R5219 DVDD.n4257 DVDD.n4243 4.5005
R5220 DVDD.n4257 DVDD.n4250 4.5005
R5221 DVDD.n4257 DVDD.n4241 4.5005
R5222 DVDD.n4257 DVDD.n4251 4.5005
R5223 DVDD.n4257 DVDD.n4240 4.5005
R5224 DVDD.n4600 DVDD.n4257 4.5005
R5225 DVDD.n4597 DVDD.n4257 4.5005
R5226 DVDD.n4257 DVDD.n4248 4.5005
R5227 DVDD.n4599 DVDD.n4245 4.5005
R5228 DVDD.n4599 DVDD.n4248 4.5005
R5229 DVDD.n4253 DVDD.n4246 4.5005
R5230 DVDD.n4253 DVDD.n4248 4.5005
R5231 DVDD.n4597 DVDD.n4268 4.5005
R5232 DVDD.n4268 DVDD.n4248 4.5005
R5233 DVDD.n4254 DVDD.n4245 4.5005
R5234 DVDD.n4254 DVDD.n4248 4.5005
R5235 DVDD.n4265 DVDD.n4246 4.5005
R5236 DVDD.n4265 DVDD.n4245 4.5005
R5237 DVDD.n4265 DVDD.n4248 4.5005
R5238 DVDD.n4255 DVDD.n4246 4.5005
R5239 DVDD.n4255 DVDD.n4245 4.5005
R5240 DVDD.n4255 DVDD.n4248 4.5005
R5241 DVDD.n4264 DVDD.n4245 4.5005
R5242 DVDD.n4264 DVDD.n4248 4.5005
R5243 DVDD.n4256 DVDD.n4245 4.5005
R5244 DVDD.n4256 DVDD.n4248 4.5005
R5245 DVDD.n4601 DVDD.n4246 4.5005
R5246 DVDD.n4601 DVDD.n4245 4.5005
R5247 DVDD.n4601 DVDD.n4248 4.5005
R5248 DVDD.n4633 DVDD.n4602 4.5005
R5249 DVDD.n4636 DVDD.n4602 4.5005
R5250 DVDD.n4630 DVDD.n4602 4.5005
R5251 DVDD.n4638 DVDD.n4602 4.5005
R5252 DVDD.n4629 DVDD.n4602 4.5005
R5253 DVDD.n4639 DVDD.n4602 4.5005
R5254 DVDD.n4628 DVDD.n4602 4.5005
R5255 DVDD.n4643 DVDD.n4602 4.5005
R5256 DVDD.n4626 DVDD.n4602 4.5005
R5257 DVDD.n4657 DVDD.n4602 4.5005
R5258 DVDD.n4659 DVDD.n4602 4.5005
R5259 DVDD.n4633 DVDD.n4603 4.5005
R5260 DVDD.n4635 DVDD.n4603 4.5005
R5261 DVDD.n4631 DVDD.n4603 4.5005
R5262 DVDD.n4636 DVDD.n4603 4.5005
R5263 DVDD.n4630 DVDD.n4603 4.5005
R5264 DVDD.n4638 DVDD.n4603 4.5005
R5265 DVDD.n4629 DVDD.n4603 4.5005
R5266 DVDD.n4639 DVDD.n4603 4.5005
R5267 DVDD.n4628 DVDD.n4603 4.5005
R5268 DVDD.n4642 DVDD.n4603 4.5005
R5269 DVDD.n4627 DVDD.n4603 4.5005
R5270 DVDD.n4643 DVDD.n4603 4.5005
R5271 DVDD.n4657 DVDD.n4603 4.5005
R5272 DVDD.n4659 DVDD.n4603 4.5005
R5273 DVDD.n4633 DVDD.n4239 4.5005
R5274 DVDD.n4635 DVDD.n4239 4.5005
R5275 DVDD.n4631 DVDD.n4239 4.5005
R5276 DVDD.n4636 DVDD.n4239 4.5005
R5277 DVDD.n4630 DVDD.n4239 4.5005
R5278 DVDD.n4638 DVDD.n4239 4.5005
R5279 DVDD.n4629 DVDD.n4239 4.5005
R5280 DVDD.n4639 DVDD.n4239 4.5005
R5281 DVDD.n4628 DVDD.n4239 4.5005
R5282 DVDD.n4642 DVDD.n4239 4.5005
R5283 DVDD.n4627 DVDD.n4239 4.5005
R5284 DVDD.n4643 DVDD.n4239 4.5005
R5285 DVDD.n4657 DVDD.n4239 4.5005
R5286 DVDD.n4659 DVDD.n4239 4.5005
R5287 DVDD.n4633 DVDD.n4604 4.5005
R5288 DVDD.n4635 DVDD.n4604 4.5005
R5289 DVDD.n4631 DVDD.n4604 4.5005
R5290 DVDD.n4636 DVDD.n4604 4.5005
R5291 DVDD.n4630 DVDD.n4604 4.5005
R5292 DVDD.n4638 DVDD.n4604 4.5005
R5293 DVDD.n4629 DVDD.n4604 4.5005
R5294 DVDD.n4639 DVDD.n4604 4.5005
R5295 DVDD.n4628 DVDD.n4604 4.5005
R5296 DVDD.n4642 DVDD.n4604 4.5005
R5297 DVDD.n4627 DVDD.n4604 4.5005
R5298 DVDD.n4643 DVDD.n4604 4.5005
R5299 DVDD.n4657 DVDD.n4604 4.5005
R5300 DVDD.n4659 DVDD.n4604 4.5005
R5301 DVDD.n4633 DVDD.n4238 4.5005
R5302 DVDD.n4635 DVDD.n4238 4.5005
R5303 DVDD.n4631 DVDD.n4238 4.5005
R5304 DVDD.n4636 DVDD.n4238 4.5005
R5305 DVDD.n4630 DVDD.n4238 4.5005
R5306 DVDD.n4638 DVDD.n4238 4.5005
R5307 DVDD.n4629 DVDD.n4238 4.5005
R5308 DVDD.n4639 DVDD.n4238 4.5005
R5309 DVDD.n4628 DVDD.n4238 4.5005
R5310 DVDD.n4642 DVDD.n4238 4.5005
R5311 DVDD.n4627 DVDD.n4238 4.5005
R5312 DVDD.n4643 DVDD.n4238 4.5005
R5313 DVDD.n4657 DVDD.n4238 4.5005
R5314 DVDD.n4659 DVDD.n4238 4.5005
R5315 DVDD.n4633 DVDD.n4605 4.5005
R5316 DVDD.n4635 DVDD.n4605 4.5005
R5317 DVDD.n4631 DVDD.n4605 4.5005
R5318 DVDD.n4636 DVDD.n4605 4.5005
R5319 DVDD.n4630 DVDD.n4605 4.5005
R5320 DVDD.n4638 DVDD.n4605 4.5005
R5321 DVDD.n4629 DVDD.n4605 4.5005
R5322 DVDD.n4639 DVDD.n4605 4.5005
R5323 DVDD.n4628 DVDD.n4605 4.5005
R5324 DVDD.n4642 DVDD.n4605 4.5005
R5325 DVDD.n4627 DVDD.n4605 4.5005
R5326 DVDD.n4643 DVDD.n4605 4.5005
R5327 DVDD.n4657 DVDD.n4605 4.5005
R5328 DVDD.n4659 DVDD.n4605 4.5005
R5329 DVDD.n4633 DVDD.n4237 4.5005
R5330 DVDD.n4635 DVDD.n4237 4.5005
R5331 DVDD.n4631 DVDD.n4237 4.5005
R5332 DVDD.n4636 DVDD.n4237 4.5005
R5333 DVDD.n4630 DVDD.n4237 4.5005
R5334 DVDD.n4638 DVDD.n4237 4.5005
R5335 DVDD.n4629 DVDD.n4237 4.5005
R5336 DVDD.n4639 DVDD.n4237 4.5005
R5337 DVDD.n4628 DVDD.n4237 4.5005
R5338 DVDD.n4642 DVDD.n4237 4.5005
R5339 DVDD.n4627 DVDD.n4237 4.5005
R5340 DVDD.n4643 DVDD.n4237 4.5005
R5341 DVDD.n4657 DVDD.n4237 4.5005
R5342 DVDD.n4659 DVDD.n4237 4.5005
R5343 DVDD.n4633 DVDD.n4606 4.5005
R5344 DVDD.n4635 DVDD.n4606 4.5005
R5345 DVDD.n4631 DVDD.n4606 4.5005
R5346 DVDD.n4636 DVDD.n4606 4.5005
R5347 DVDD.n4630 DVDD.n4606 4.5005
R5348 DVDD.n4638 DVDD.n4606 4.5005
R5349 DVDD.n4629 DVDD.n4606 4.5005
R5350 DVDD.n4639 DVDD.n4606 4.5005
R5351 DVDD.n4628 DVDD.n4606 4.5005
R5352 DVDD.n4642 DVDD.n4606 4.5005
R5353 DVDD.n4627 DVDD.n4606 4.5005
R5354 DVDD.n4643 DVDD.n4606 4.5005
R5355 DVDD.n4657 DVDD.n4606 4.5005
R5356 DVDD.n4659 DVDD.n4606 4.5005
R5357 DVDD.n4633 DVDD.n4236 4.5005
R5358 DVDD.n4635 DVDD.n4236 4.5005
R5359 DVDD.n4631 DVDD.n4236 4.5005
R5360 DVDD.n4636 DVDD.n4236 4.5005
R5361 DVDD.n4630 DVDD.n4236 4.5005
R5362 DVDD.n4638 DVDD.n4236 4.5005
R5363 DVDD.n4629 DVDD.n4236 4.5005
R5364 DVDD.n4639 DVDD.n4236 4.5005
R5365 DVDD.n4628 DVDD.n4236 4.5005
R5366 DVDD.n4642 DVDD.n4236 4.5005
R5367 DVDD.n4627 DVDD.n4236 4.5005
R5368 DVDD.n4643 DVDD.n4236 4.5005
R5369 DVDD.n4657 DVDD.n4236 4.5005
R5370 DVDD.n4659 DVDD.n4236 4.5005
R5371 DVDD.n4633 DVDD.n4607 4.5005
R5372 DVDD.n4635 DVDD.n4607 4.5005
R5373 DVDD.n4631 DVDD.n4607 4.5005
R5374 DVDD.n4636 DVDD.n4607 4.5005
R5375 DVDD.n4630 DVDD.n4607 4.5005
R5376 DVDD.n4638 DVDD.n4607 4.5005
R5377 DVDD.n4629 DVDD.n4607 4.5005
R5378 DVDD.n4639 DVDD.n4607 4.5005
R5379 DVDD.n4628 DVDD.n4607 4.5005
R5380 DVDD.n4642 DVDD.n4607 4.5005
R5381 DVDD.n4627 DVDD.n4607 4.5005
R5382 DVDD.n4643 DVDD.n4607 4.5005
R5383 DVDD.n4657 DVDD.n4607 4.5005
R5384 DVDD.n4659 DVDD.n4607 4.5005
R5385 DVDD.n4633 DVDD.n4235 4.5005
R5386 DVDD.n4635 DVDD.n4235 4.5005
R5387 DVDD.n4631 DVDD.n4235 4.5005
R5388 DVDD.n4636 DVDD.n4235 4.5005
R5389 DVDD.n4630 DVDD.n4235 4.5005
R5390 DVDD.n4638 DVDD.n4235 4.5005
R5391 DVDD.n4629 DVDD.n4235 4.5005
R5392 DVDD.n4639 DVDD.n4235 4.5005
R5393 DVDD.n4628 DVDD.n4235 4.5005
R5394 DVDD.n4642 DVDD.n4235 4.5005
R5395 DVDD.n4627 DVDD.n4235 4.5005
R5396 DVDD.n4643 DVDD.n4235 4.5005
R5397 DVDD.n4657 DVDD.n4235 4.5005
R5398 DVDD.n4659 DVDD.n4235 4.5005
R5399 DVDD.n4633 DVDD.n4608 4.5005
R5400 DVDD.n4635 DVDD.n4608 4.5005
R5401 DVDD.n4631 DVDD.n4608 4.5005
R5402 DVDD.n4636 DVDD.n4608 4.5005
R5403 DVDD.n4630 DVDD.n4608 4.5005
R5404 DVDD.n4638 DVDD.n4608 4.5005
R5405 DVDD.n4629 DVDD.n4608 4.5005
R5406 DVDD.n4639 DVDD.n4608 4.5005
R5407 DVDD.n4628 DVDD.n4608 4.5005
R5408 DVDD.n4642 DVDD.n4608 4.5005
R5409 DVDD.n4627 DVDD.n4608 4.5005
R5410 DVDD.n4643 DVDD.n4608 4.5005
R5411 DVDD.n4657 DVDD.n4608 4.5005
R5412 DVDD.n4659 DVDD.n4608 4.5005
R5413 DVDD.n4633 DVDD.n4234 4.5005
R5414 DVDD.n4635 DVDD.n4234 4.5005
R5415 DVDD.n4631 DVDD.n4234 4.5005
R5416 DVDD.n4636 DVDD.n4234 4.5005
R5417 DVDD.n4630 DVDD.n4234 4.5005
R5418 DVDD.n4638 DVDD.n4234 4.5005
R5419 DVDD.n4629 DVDD.n4234 4.5005
R5420 DVDD.n4639 DVDD.n4234 4.5005
R5421 DVDD.n4628 DVDD.n4234 4.5005
R5422 DVDD.n4642 DVDD.n4234 4.5005
R5423 DVDD.n4627 DVDD.n4234 4.5005
R5424 DVDD.n4643 DVDD.n4234 4.5005
R5425 DVDD.n4657 DVDD.n4234 4.5005
R5426 DVDD.n4659 DVDD.n4234 4.5005
R5427 DVDD.n4633 DVDD.n4609 4.5005
R5428 DVDD.n4635 DVDD.n4609 4.5005
R5429 DVDD.n4631 DVDD.n4609 4.5005
R5430 DVDD.n4636 DVDD.n4609 4.5005
R5431 DVDD.n4630 DVDD.n4609 4.5005
R5432 DVDD.n4638 DVDD.n4609 4.5005
R5433 DVDD.n4629 DVDD.n4609 4.5005
R5434 DVDD.n4639 DVDD.n4609 4.5005
R5435 DVDD.n4628 DVDD.n4609 4.5005
R5436 DVDD.n4642 DVDD.n4609 4.5005
R5437 DVDD.n4627 DVDD.n4609 4.5005
R5438 DVDD.n4643 DVDD.n4609 4.5005
R5439 DVDD.n4657 DVDD.n4609 4.5005
R5440 DVDD.n4659 DVDD.n4609 4.5005
R5441 DVDD.n4633 DVDD.n4233 4.5005
R5442 DVDD.n4635 DVDD.n4233 4.5005
R5443 DVDD.n4631 DVDD.n4233 4.5005
R5444 DVDD.n4636 DVDD.n4233 4.5005
R5445 DVDD.n4630 DVDD.n4233 4.5005
R5446 DVDD.n4638 DVDD.n4233 4.5005
R5447 DVDD.n4629 DVDD.n4233 4.5005
R5448 DVDD.n4639 DVDD.n4233 4.5005
R5449 DVDD.n4628 DVDD.n4233 4.5005
R5450 DVDD.n4642 DVDD.n4233 4.5005
R5451 DVDD.n4627 DVDD.n4233 4.5005
R5452 DVDD.n4643 DVDD.n4233 4.5005
R5453 DVDD.n4657 DVDD.n4233 4.5005
R5454 DVDD.n4659 DVDD.n4233 4.5005
R5455 DVDD.n4633 DVDD.n4610 4.5005
R5456 DVDD.n4635 DVDD.n4610 4.5005
R5457 DVDD.n4631 DVDD.n4610 4.5005
R5458 DVDD.n4636 DVDD.n4610 4.5005
R5459 DVDD.n4630 DVDD.n4610 4.5005
R5460 DVDD.n4638 DVDD.n4610 4.5005
R5461 DVDD.n4629 DVDD.n4610 4.5005
R5462 DVDD.n4639 DVDD.n4610 4.5005
R5463 DVDD.n4628 DVDD.n4610 4.5005
R5464 DVDD.n4642 DVDD.n4610 4.5005
R5465 DVDD.n4627 DVDD.n4610 4.5005
R5466 DVDD.n4643 DVDD.n4610 4.5005
R5467 DVDD.n4657 DVDD.n4610 4.5005
R5468 DVDD.n4659 DVDD.n4610 4.5005
R5469 DVDD.n4633 DVDD.n4232 4.5005
R5470 DVDD.n4635 DVDD.n4232 4.5005
R5471 DVDD.n4631 DVDD.n4232 4.5005
R5472 DVDD.n4636 DVDD.n4232 4.5005
R5473 DVDD.n4630 DVDD.n4232 4.5005
R5474 DVDD.n4638 DVDD.n4232 4.5005
R5475 DVDD.n4629 DVDD.n4232 4.5005
R5476 DVDD.n4639 DVDD.n4232 4.5005
R5477 DVDD.n4628 DVDD.n4232 4.5005
R5478 DVDD.n4642 DVDD.n4232 4.5005
R5479 DVDD.n4627 DVDD.n4232 4.5005
R5480 DVDD.n4643 DVDD.n4232 4.5005
R5481 DVDD.n4657 DVDD.n4232 4.5005
R5482 DVDD.n4659 DVDD.n4232 4.5005
R5483 DVDD.n4633 DVDD.n4611 4.5005
R5484 DVDD.n4635 DVDD.n4611 4.5005
R5485 DVDD.n4631 DVDD.n4611 4.5005
R5486 DVDD.n4636 DVDD.n4611 4.5005
R5487 DVDD.n4630 DVDD.n4611 4.5005
R5488 DVDD.n4638 DVDD.n4611 4.5005
R5489 DVDD.n4629 DVDD.n4611 4.5005
R5490 DVDD.n4639 DVDD.n4611 4.5005
R5491 DVDD.n4628 DVDD.n4611 4.5005
R5492 DVDD.n4642 DVDD.n4611 4.5005
R5493 DVDD.n4627 DVDD.n4611 4.5005
R5494 DVDD.n4643 DVDD.n4611 4.5005
R5495 DVDD.n4657 DVDD.n4611 4.5005
R5496 DVDD.n4659 DVDD.n4611 4.5005
R5497 DVDD.n4633 DVDD.n4231 4.5005
R5498 DVDD.n4635 DVDD.n4231 4.5005
R5499 DVDD.n4631 DVDD.n4231 4.5005
R5500 DVDD.n4636 DVDD.n4231 4.5005
R5501 DVDD.n4630 DVDD.n4231 4.5005
R5502 DVDD.n4638 DVDD.n4231 4.5005
R5503 DVDD.n4629 DVDD.n4231 4.5005
R5504 DVDD.n4639 DVDD.n4231 4.5005
R5505 DVDD.n4628 DVDD.n4231 4.5005
R5506 DVDD.n4642 DVDD.n4231 4.5005
R5507 DVDD.n4627 DVDD.n4231 4.5005
R5508 DVDD.n4643 DVDD.n4231 4.5005
R5509 DVDD.n4657 DVDD.n4231 4.5005
R5510 DVDD.n4659 DVDD.n4231 4.5005
R5511 DVDD.n4633 DVDD.n4612 4.5005
R5512 DVDD.n4635 DVDD.n4612 4.5005
R5513 DVDD.n4631 DVDD.n4612 4.5005
R5514 DVDD.n4636 DVDD.n4612 4.5005
R5515 DVDD.n4630 DVDD.n4612 4.5005
R5516 DVDD.n4638 DVDD.n4612 4.5005
R5517 DVDD.n4629 DVDD.n4612 4.5005
R5518 DVDD.n4639 DVDD.n4612 4.5005
R5519 DVDD.n4628 DVDD.n4612 4.5005
R5520 DVDD.n4642 DVDD.n4612 4.5005
R5521 DVDD.n4627 DVDD.n4612 4.5005
R5522 DVDD.n4643 DVDD.n4612 4.5005
R5523 DVDD.n4657 DVDD.n4612 4.5005
R5524 DVDD.n4659 DVDD.n4612 4.5005
R5525 DVDD.n4633 DVDD.n4230 4.5005
R5526 DVDD.n4635 DVDD.n4230 4.5005
R5527 DVDD.n4631 DVDD.n4230 4.5005
R5528 DVDD.n4636 DVDD.n4230 4.5005
R5529 DVDD.n4630 DVDD.n4230 4.5005
R5530 DVDD.n4638 DVDD.n4230 4.5005
R5531 DVDD.n4629 DVDD.n4230 4.5005
R5532 DVDD.n4639 DVDD.n4230 4.5005
R5533 DVDD.n4628 DVDD.n4230 4.5005
R5534 DVDD.n4642 DVDD.n4230 4.5005
R5535 DVDD.n4627 DVDD.n4230 4.5005
R5536 DVDD.n4643 DVDD.n4230 4.5005
R5537 DVDD.n4657 DVDD.n4230 4.5005
R5538 DVDD.n4659 DVDD.n4230 4.5005
R5539 DVDD.n4633 DVDD.n4613 4.5005
R5540 DVDD.n4635 DVDD.n4613 4.5005
R5541 DVDD.n4631 DVDD.n4613 4.5005
R5542 DVDD.n4636 DVDD.n4613 4.5005
R5543 DVDD.n4630 DVDD.n4613 4.5005
R5544 DVDD.n4638 DVDD.n4613 4.5005
R5545 DVDD.n4629 DVDD.n4613 4.5005
R5546 DVDD.n4639 DVDD.n4613 4.5005
R5547 DVDD.n4628 DVDD.n4613 4.5005
R5548 DVDD.n4642 DVDD.n4613 4.5005
R5549 DVDD.n4627 DVDD.n4613 4.5005
R5550 DVDD.n4643 DVDD.n4613 4.5005
R5551 DVDD.n4657 DVDD.n4613 4.5005
R5552 DVDD.n4659 DVDD.n4613 4.5005
R5553 DVDD.n4633 DVDD.n4229 4.5005
R5554 DVDD.n4635 DVDD.n4229 4.5005
R5555 DVDD.n4631 DVDD.n4229 4.5005
R5556 DVDD.n4636 DVDD.n4229 4.5005
R5557 DVDD.n4630 DVDD.n4229 4.5005
R5558 DVDD.n4638 DVDD.n4229 4.5005
R5559 DVDD.n4629 DVDD.n4229 4.5005
R5560 DVDD.n4639 DVDD.n4229 4.5005
R5561 DVDD.n4628 DVDD.n4229 4.5005
R5562 DVDD.n4642 DVDD.n4229 4.5005
R5563 DVDD.n4627 DVDD.n4229 4.5005
R5564 DVDD.n4643 DVDD.n4229 4.5005
R5565 DVDD.n4657 DVDD.n4229 4.5005
R5566 DVDD.n4659 DVDD.n4229 4.5005
R5567 DVDD.n4658 DVDD.n4633 4.5005
R5568 DVDD.n4658 DVDD.n4635 4.5005
R5569 DVDD.n4658 DVDD.n4631 4.5005
R5570 DVDD.n4658 DVDD.n4636 4.5005
R5571 DVDD.n4658 DVDD.n4630 4.5005
R5572 DVDD.n4658 DVDD.n4638 4.5005
R5573 DVDD.n4658 DVDD.n4629 4.5005
R5574 DVDD.n4658 DVDD.n4639 4.5005
R5575 DVDD.n4658 DVDD.n4628 4.5005
R5576 DVDD.n4658 DVDD.n4642 4.5005
R5577 DVDD.n4658 DVDD.n4627 4.5005
R5578 DVDD.n4658 DVDD.n4643 4.5005
R5579 DVDD.n4658 DVDD.n4626 4.5005
R5580 DVDD.n4658 DVDD.n4657 4.5005
R5581 DVDD.n4659 DVDD.n4658 4.5005
R5582 DVDD.n22140 DVDD.n361 4.5005
R5583 DVDD.n381 DVDD.n361 4.5005
R5584 DVDD.n377 DVDD.n361 4.5005
R5585 DVDD.n382 DVDD.n361 4.5005
R5586 DVDD.n376 DVDD.n361 4.5005
R5587 DVDD.n383 DVDD.n361 4.5005
R5588 DVDD.n375 DVDD.n361 4.5005
R5589 DVDD.n386 DVDD.n361 4.5005
R5590 DVDD.n426 DVDD.n361 4.5005
R5591 DVDD.n387 DVDD.n361 4.5005
R5592 DVDD.n22138 DVDD.n361 4.5005
R5593 DVDD.n22140 DVDD.n359 4.5005
R5594 DVDD.n380 DVDD.n359 4.5005
R5595 DVDD.n378 DVDD.n359 4.5005
R5596 DVDD.n381 DVDD.n359 4.5005
R5597 DVDD.n377 DVDD.n359 4.5005
R5598 DVDD.n382 DVDD.n359 4.5005
R5599 DVDD.n376 DVDD.n359 4.5005
R5600 DVDD.n383 DVDD.n359 4.5005
R5601 DVDD.n375 DVDD.n359 4.5005
R5602 DVDD.n385 DVDD.n359 4.5005
R5603 DVDD.n374 DVDD.n359 4.5005
R5604 DVDD.n386 DVDD.n359 4.5005
R5605 DVDD.n387 DVDD.n359 4.5005
R5606 DVDD.n22138 DVDD.n359 4.5005
R5607 DVDD.n22140 DVDD.n362 4.5005
R5608 DVDD.n380 DVDD.n362 4.5005
R5609 DVDD.n378 DVDD.n362 4.5005
R5610 DVDD.n381 DVDD.n362 4.5005
R5611 DVDD.n377 DVDD.n362 4.5005
R5612 DVDD.n382 DVDD.n362 4.5005
R5613 DVDD.n376 DVDD.n362 4.5005
R5614 DVDD.n383 DVDD.n362 4.5005
R5615 DVDD.n375 DVDD.n362 4.5005
R5616 DVDD.n385 DVDD.n362 4.5005
R5617 DVDD.n374 DVDD.n362 4.5005
R5618 DVDD.n386 DVDD.n362 4.5005
R5619 DVDD.n387 DVDD.n362 4.5005
R5620 DVDD.n22138 DVDD.n362 4.5005
R5621 DVDD.n22140 DVDD.n358 4.5005
R5622 DVDD.n380 DVDD.n358 4.5005
R5623 DVDD.n378 DVDD.n358 4.5005
R5624 DVDD.n381 DVDD.n358 4.5005
R5625 DVDD.n377 DVDD.n358 4.5005
R5626 DVDD.n382 DVDD.n358 4.5005
R5627 DVDD.n376 DVDD.n358 4.5005
R5628 DVDD.n383 DVDD.n358 4.5005
R5629 DVDD.n375 DVDD.n358 4.5005
R5630 DVDD.n385 DVDD.n358 4.5005
R5631 DVDD.n374 DVDD.n358 4.5005
R5632 DVDD.n386 DVDD.n358 4.5005
R5633 DVDD.n387 DVDD.n358 4.5005
R5634 DVDD.n22138 DVDD.n358 4.5005
R5635 DVDD.n22140 DVDD.n363 4.5005
R5636 DVDD.n380 DVDD.n363 4.5005
R5637 DVDD.n378 DVDD.n363 4.5005
R5638 DVDD.n381 DVDD.n363 4.5005
R5639 DVDD.n377 DVDD.n363 4.5005
R5640 DVDD.n382 DVDD.n363 4.5005
R5641 DVDD.n376 DVDD.n363 4.5005
R5642 DVDD.n383 DVDD.n363 4.5005
R5643 DVDD.n375 DVDD.n363 4.5005
R5644 DVDD.n385 DVDD.n363 4.5005
R5645 DVDD.n374 DVDD.n363 4.5005
R5646 DVDD.n386 DVDD.n363 4.5005
R5647 DVDD.n387 DVDD.n363 4.5005
R5648 DVDD.n22138 DVDD.n363 4.5005
R5649 DVDD.n22140 DVDD.n357 4.5005
R5650 DVDD.n380 DVDD.n357 4.5005
R5651 DVDD.n378 DVDD.n357 4.5005
R5652 DVDD.n381 DVDD.n357 4.5005
R5653 DVDD.n377 DVDD.n357 4.5005
R5654 DVDD.n382 DVDD.n357 4.5005
R5655 DVDD.n376 DVDD.n357 4.5005
R5656 DVDD.n383 DVDD.n357 4.5005
R5657 DVDD.n375 DVDD.n357 4.5005
R5658 DVDD.n385 DVDD.n357 4.5005
R5659 DVDD.n374 DVDD.n357 4.5005
R5660 DVDD.n386 DVDD.n357 4.5005
R5661 DVDD.n387 DVDD.n357 4.5005
R5662 DVDD.n22138 DVDD.n357 4.5005
R5663 DVDD.n22140 DVDD.n364 4.5005
R5664 DVDD.n380 DVDD.n364 4.5005
R5665 DVDD.n378 DVDD.n364 4.5005
R5666 DVDD.n381 DVDD.n364 4.5005
R5667 DVDD.n377 DVDD.n364 4.5005
R5668 DVDD.n382 DVDD.n364 4.5005
R5669 DVDD.n376 DVDD.n364 4.5005
R5670 DVDD.n383 DVDD.n364 4.5005
R5671 DVDD.n375 DVDD.n364 4.5005
R5672 DVDD.n385 DVDD.n364 4.5005
R5673 DVDD.n374 DVDD.n364 4.5005
R5674 DVDD.n386 DVDD.n364 4.5005
R5675 DVDD.n387 DVDD.n364 4.5005
R5676 DVDD.n22138 DVDD.n364 4.5005
R5677 DVDD.n22140 DVDD.n356 4.5005
R5678 DVDD.n380 DVDD.n356 4.5005
R5679 DVDD.n378 DVDD.n356 4.5005
R5680 DVDD.n381 DVDD.n356 4.5005
R5681 DVDD.n377 DVDD.n356 4.5005
R5682 DVDD.n382 DVDD.n356 4.5005
R5683 DVDD.n376 DVDD.n356 4.5005
R5684 DVDD.n383 DVDD.n356 4.5005
R5685 DVDD.n375 DVDD.n356 4.5005
R5686 DVDD.n385 DVDD.n356 4.5005
R5687 DVDD.n374 DVDD.n356 4.5005
R5688 DVDD.n386 DVDD.n356 4.5005
R5689 DVDD.n387 DVDD.n356 4.5005
R5690 DVDD.n22138 DVDD.n356 4.5005
R5691 DVDD.n22140 DVDD.n365 4.5005
R5692 DVDD.n380 DVDD.n365 4.5005
R5693 DVDD.n378 DVDD.n365 4.5005
R5694 DVDD.n381 DVDD.n365 4.5005
R5695 DVDD.n377 DVDD.n365 4.5005
R5696 DVDD.n382 DVDD.n365 4.5005
R5697 DVDD.n376 DVDD.n365 4.5005
R5698 DVDD.n383 DVDD.n365 4.5005
R5699 DVDD.n375 DVDD.n365 4.5005
R5700 DVDD.n385 DVDD.n365 4.5005
R5701 DVDD.n374 DVDD.n365 4.5005
R5702 DVDD.n386 DVDD.n365 4.5005
R5703 DVDD.n387 DVDD.n365 4.5005
R5704 DVDD.n22138 DVDD.n365 4.5005
R5705 DVDD.n22140 DVDD.n355 4.5005
R5706 DVDD.n380 DVDD.n355 4.5005
R5707 DVDD.n378 DVDD.n355 4.5005
R5708 DVDD.n381 DVDD.n355 4.5005
R5709 DVDD.n377 DVDD.n355 4.5005
R5710 DVDD.n382 DVDD.n355 4.5005
R5711 DVDD.n376 DVDD.n355 4.5005
R5712 DVDD.n383 DVDD.n355 4.5005
R5713 DVDD.n375 DVDD.n355 4.5005
R5714 DVDD.n385 DVDD.n355 4.5005
R5715 DVDD.n374 DVDD.n355 4.5005
R5716 DVDD.n386 DVDD.n355 4.5005
R5717 DVDD.n387 DVDD.n355 4.5005
R5718 DVDD.n22138 DVDD.n355 4.5005
R5719 DVDD.n22140 DVDD.n22139 4.5005
R5720 DVDD.n22139 DVDD.n380 4.5005
R5721 DVDD.n22139 DVDD.n378 4.5005
R5722 DVDD.n22139 DVDD.n381 4.5005
R5723 DVDD.n22139 DVDD.n377 4.5005
R5724 DVDD.n22139 DVDD.n382 4.5005
R5725 DVDD.n22139 DVDD.n376 4.5005
R5726 DVDD.n22139 DVDD.n383 4.5005
R5727 DVDD.n22139 DVDD.n375 4.5005
R5728 DVDD.n22139 DVDD.n385 4.5005
R5729 DVDD.n22139 DVDD.n374 4.5005
R5730 DVDD.n22139 DVDD.n386 4.5005
R5731 DVDD.n22139 DVDD.n387 4.5005
R5732 DVDD.n22139 DVDD.n372 4.5005
R5733 DVDD.n22139 DVDD.n22138 4.5005
R5734 DVDD.n20929 DVDD.n18896 4.5005
R5735 DVDD.n18896 DVDD.n18873 4.5005
R5736 DVDD.n18896 DVDD.n18885 4.5005
R5737 DVDD.n18896 DVDD.n18874 4.5005
R5738 DVDD.n18896 DVDD.n18884 4.5005
R5739 DVDD.n18896 DVDD.n18875 4.5005
R5740 DVDD.n18896 DVDD.n18883 4.5005
R5741 DVDD.n18896 DVDD.n18878 4.5005
R5742 DVDD.n18896 DVDD.n18881 4.5005
R5743 DVDD.n18896 DVDD.n18877 4.5005
R5744 DVDD.n18896 DVDD.n18882 4.5005
R5745 DVDD.n18896 DVDD.n18876 4.5005
R5746 DVDD.n20929 DVDD.n18892 4.5005
R5747 DVDD.n18892 DVDD.n18872 4.5005
R5748 DVDD.n18892 DVDD.n18886 4.5005
R5749 DVDD.n18892 DVDD.n18873 4.5005
R5750 DVDD.n18892 DVDD.n18885 4.5005
R5751 DVDD.n18892 DVDD.n18874 4.5005
R5752 DVDD.n18892 DVDD.n18884 4.5005
R5753 DVDD.n18892 DVDD.n18875 4.5005
R5754 DVDD.n18892 DVDD.n18883 4.5005
R5755 DVDD.n18892 DVDD.n18879 4.5005
R5756 DVDD.n18892 DVDD.n18880 4.5005
R5757 DVDD.n18892 DVDD.n18878 4.5005
R5758 DVDD.n18892 DVDD.n18881 4.5005
R5759 DVDD.n18892 DVDD.n18877 4.5005
R5760 DVDD.n18892 DVDD.n18876 4.5005
R5761 DVDD.n20929 DVDD.n18899 4.5005
R5762 DVDD.n18899 DVDD.n18872 4.5005
R5763 DVDD.n18899 DVDD.n18886 4.5005
R5764 DVDD.n18899 DVDD.n18873 4.5005
R5765 DVDD.n18899 DVDD.n18885 4.5005
R5766 DVDD.n18899 DVDD.n18874 4.5005
R5767 DVDD.n18899 DVDD.n18884 4.5005
R5768 DVDD.n18899 DVDD.n18875 4.5005
R5769 DVDD.n18899 DVDD.n18883 4.5005
R5770 DVDD.n18899 DVDD.n18879 4.5005
R5771 DVDD.n18899 DVDD.n18880 4.5005
R5772 DVDD.n18899 DVDD.n18878 4.5005
R5773 DVDD.n18899 DVDD.n18877 4.5005
R5774 DVDD.n18899 DVDD.n18876 4.5005
R5775 DVDD.n20929 DVDD.n18891 4.5005
R5776 DVDD.n18891 DVDD.n18872 4.5005
R5777 DVDD.n18891 DVDD.n18886 4.5005
R5778 DVDD.n18891 DVDD.n18873 4.5005
R5779 DVDD.n18891 DVDD.n18885 4.5005
R5780 DVDD.n18891 DVDD.n18874 4.5005
R5781 DVDD.n18891 DVDD.n18884 4.5005
R5782 DVDD.n18891 DVDD.n18875 4.5005
R5783 DVDD.n18891 DVDD.n18883 4.5005
R5784 DVDD.n18891 DVDD.n18879 4.5005
R5785 DVDD.n18891 DVDD.n18880 4.5005
R5786 DVDD.n18891 DVDD.n18878 4.5005
R5787 DVDD.n18891 DVDD.n18877 4.5005
R5788 DVDD.n18891 DVDD.n18876 4.5005
R5789 DVDD.n20929 DVDD.n18902 4.5005
R5790 DVDD.n18902 DVDD.n18872 4.5005
R5791 DVDD.n18902 DVDD.n18886 4.5005
R5792 DVDD.n18902 DVDD.n18873 4.5005
R5793 DVDD.n18902 DVDD.n18885 4.5005
R5794 DVDD.n18902 DVDD.n18874 4.5005
R5795 DVDD.n18902 DVDD.n18884 4.5005
R5796 DVDD.n18902 DVDD.n18875 4.5005
R5797 DVDD.n18902 DVDD.n18883 4.5005
R5798 DVDD.n18902 DVDD.n18879 4.5005
R5799 DVDD.n18902 DVDD.n18880 4.5005
R5800 DVDD.n18902 DVDD.n18878 4.5005
R5801 DVDD.n18902 DVDD.n18877 4.5005
R5802 DVDD.n18902 DVDD.n18876 4.5005
R5803 DVDD.n20929 DVDD.n18890 4.5005
R5804 DVDD.n18890 DVDD.n18872 4.5005
R5805 DVDD.n18890 DVDD.n18886 4.5005
R5806 DVDD.n18890 DVDD.n18873 4.5005
R5807 DVDD.n18890 DVDD.n18885 4.5005
R5808 DVDD.n18890 DVDD.n18874 4.5005
R5809 DVDD.n18890 DVDD.n18884 4.5005
R5810 DVDD.n18890 DVDD.n18875 4.5005
R5811 DVDD.n18890 DVDD.n18883 4.5005
R5812 DVDD.n18890 DVDD.n18879 4.5005
R5813 DVDD.n18890 DVDD.n18880 4.5005
R5814 DVDD.n18890 DVDD.n18878 4.5005
R5815 DVDD.n18890 DVDD.n18877 4.5005
R5816 DVDD.n18890 DVDD.n18876 4.5005
R5817 DVDD.n20929 DVDD.n18904 4.5005
R5818 DVDD.n18904 DVDD.n18872 4.5005
R5819 DVDD.n18904 DVDD.n18886 4.5005
R5820 DVDD.n18904 DVDD.n18873 4.5005
R5821 DVDD.n18904 DVDD.n18885 4.5005
R5822 DVDD.n18904 DVDD.n18874 4.5005
R5823 DVDD.n18904 DVDD.n18884 4.5005
R5824 DVDD.n18904 DVDD.n18875 4.5005
R5825 DVDD.n18904 DVDD.n18883 4.5005
R5826 DVDD.n18904 DVDD.n18879 4.5005
R5827 DVDD.n18904 DVDD.n18880 4.5005
R5828 DVDD.n18904 DVDD.n18878 4.5005
R5829 DVDD.n18904 DVDD.n18881 4.5005
R5830 DVDD.n18904 DVDD.n18877 4.5005
R5831 DVDD.n18904 DVDD.n18876 4.5005
R5832 DVDD.n20930 DVDD.n18879 4.5005
R5833 DVDD.n20930 DVDD.n18880 4.5005
R5834 DVDD.n20930 DVDD.n18878 4.5005
R5835 DVDD.n20930 DVDD.n18881 4.5005
R5836 DVDD.n20930 DVDD.n18877 4.5005
R5837 DVDD.n20930 DVDD.n18882 4.5005
R5838 DVDD.n20930 DVDD.n18876 4.5005
R5839 DVDD.n18879 DVDD.n18871 4.5005
R5840 DVDD.n18880 DVDD.n18871 4.5005
R5841 DVDD.n18878 DVDD.n18871 4.5005
R5842 DVDD.n18877 DVDD.n18871 4.5005
R5843 DVDD.n18882 DVDD.n18871 4.5005
R5844 DVDD.n18876 DVDD.n18871 4.5005
R5845 DVDD.n20929 DVDD.n18889 4.5005
R5846 DVDD.n18889 DVDD.n18872 4.5005
R5847 DVDD.n18889 DVDD.n18886 4.5005
R5848 DVDD.n18889 DVDD.n18873 4.5005
R5849 DVDD.n18889 DVDD.n18885 4.5005
R5850 DVDD.n18889 DVDD.n18874 4.5005
R5851 DVDD.n18889 DVDD.n18884 4.5005
R5852 DVDD.n18889 DVDD.n18875 4.5005
R5853 DVDD.n18889 DVDD.n18883 4.5005
R5854 DVDD.n18889 DVDD.n18879 4.5005
R5855 DVDD.n18889 DVDD.n18880 4.5005
R5856 DVDD.n18889 DVDD.n18878 4.5005
R5857 DVDD.n18889 DVDD.n18877 4.5005
R5858 DVDD.n18889 DVDD.n18876 4.5005
R5859 DVDD.n20929 DVDD.n20928 4.5005
R5860 DVDD.n20928 DVDD.n18872 4.5005
R5861 DVDD.n20928 DVDD.n18886 4.5005
R5862 DVDD.n20928 DVDD.n18873 4.5005
R5863 DVDD.n20928 DVDD.n18885 4.5005
R5864 DVDD.n20928 DVDD.n18874 4.5005
R5865 DVDD.n20928 DVDD.n18884 4.5005
R5866 DVDD.n20928 DVDD.n18875 4.5005
R5867 DVDD.n20928 DVDD.n18883 4.5005
R5868 DVDD.n20928 DVDD.n18879 4.5005
R5869 DVDD.n20928 DVDD.n18880 4.5005
R5870 DVDD.n20928 DVDD.n18878 4.5005
R5871 DVDD.n20928 DVDD.n18881 4.5005
R5872 DVDD.n20928 DVDD.n18877 4.5005
R5873 DVDD.n20928 DVDD.n18876 4.5005
R5874 DVDD.n20374 DVDD.n19841 4.5005
R5875 DVDD.n20374 DVDD.n19844 4.5005
R5876 DVDD.n20374 DVDD.n19839 4.5005
R5877 DVDD.n20374 DVDD.n19845 4.5005
R5878 DVDD.n20374 DVDD.n19838 4.5005
R5879 DVDD.n20374 DVDD.n19846 4.5005
R5880 DVDD.n20374 DVDD.n19837 4.5005
R5881 DVDD.n20374 DVDD.n19848 4.5005
R5882 DVDD.n20374 DVDD.n19835 4.5005
R5883 DVDD.n20374 DVDD.n19849 4.5005
R5884 DVDD.n20374 DVDD.n19834 4.5005
R5885 DVDD.n20420 DVDD.n20374 4.5005
R5886 DVDD.n19854 DVDD.n19841 4.5005
R5887 DVDD.n19854 DVDD.n19843 4.5005
R5888 DVDD.n19854 DVDD.n19840 4.5005
R5889 DVDD.n19854 DVDD.n19844 4.5005
R5890 DVDD.n19854 DVDD.n19839 4.5005
R5891 DVDD.n19854 DVDD.n19845 4.5005
R5892 DVDD.n19854 DVDD.n19838 4.5005
R5893 DVDD.n19854 DVDD.n19846 4.5005
R5894 DVDD.n19854 DVDD.n19837 4.5005
R5895 DVDD.n19854 DVDD.n19847 4.5005
R5896 DVDD.n19854 DVDD.n19836 4.5005
R5897 DVDD.n19854 DVDD.n19848 4.5005
R5898 DVDD.n19854 DVDD.n19835 4.5005
R5899 DVDD.n19854 DVDD.n19849 4.5005
R5900 DVDD.n19854 DVDD.n19834 4.5005
R5901 DVDD.n20420 DVDD.n19854 4.5005
R5902 DVDD.n20375 DVDD.n19841 4.5005
R5903 DVDD.n20375 DVDD.n19843 4.5005
R5904 DVDD.n20375 DVDD.n19840 4.5005
R5905 DVDD.n20375 DVDD.n19844 4.5005
R5906 DVDD.n20375 DVDD.n19839 4.5005
R5907 DVDD.n20375 DVDD.n19845 4.5005
R5908 DVDD.n20375 DVDD.n19838 4.5005
R5909 DVDD.n20375 DVDD.n19846 4.5005
R5910 DVDD.n20375 DVDD.n19837 4.5005
R5911 DVDD.n20375 DVDD.n19847 4.5005
R5912 DVDD.n20375 DVDD.n19836 4.5005
R5913 DVDD.n20375 DVDD.n19848 4.5005
R5914 DVDD.n20375 DVDD.n19835 4.5005
R5915 DVDD.n20375 DVDD.n19849 4.5005
R5916 DVDD.n20375 DVDD.n19834 4.5005
R5917 DVDD.n20420 DVDD.n20375 4.5005
R5918 DVDD.n19853 DVDD.n19841 4.5005
R5919 DVDD.n19853 DVDD.n19843 4.5005
R5920 DVDD.n19853 DVDD.n19840 4.5005
R5921 DVDD.n19853 DVDD.n19844 4.5005
R5922 DVDD.n19853 DVDD.n19839 4.5005
R5923 DVDD.n19853 DVDD.n19845 4.5005
R5924 DVDD.n19853 DVDD.n19838 4.5005
R5925 DVDD.n19853 DVDD.n19846 4.5005
R5926 DVDD.n19853 DVDD.n19837 4.5005
R5927 DVDD.n19853 DVDD.n19847 4.5005
R5928 DVDD.n19853 DVDD.n19836 4.5005
R5929 DVDD.n19853 DVDD.n19848 4.5005
R5930 DVDD.n19853 DVDD.n19835 4.5005
R5931 DVDD.n19853 DVDD.n19849 4.5005
R5932 DVDD.n19853 DVDD.n19834 4.5005
R5933 DVDD.n20420 DVDD.n19853 4.5005
R5934 DVDD.n20376 DVDD.n19841 4.5005
R5935 DVDD.n20376 DVDD.n19843 4.5005
R5936 DVDD.n20376 DVDD.n19840 4.5005
R5937 DVDD.n20376 DVDD.n19844 4.5005
R5938 DVDD.n20376 DVDD.n19839 4.5005
R5939 DVDD.n20376 DVDD.n19845 4.5005
R5940 DVDD.n20376 DVDD.n19838 4.5005
R5941 DVDD.n20376 DVDD.n19846 4.5005
R5942 DVDD.n20376 DVDD.n19837 4.5005
R5943 DVDD.n20376 DVDD.n19847 4.5005
R5944 DVDD.n20376 DVDD.n19836 4.5005
R5945 DVDD.n20376 DVDD.n19848 4.5005
R5946 DVDD.n20376 DVDD.n19835 4.5005
R5947 DVDD.n20376 DVDD.n19849 4.5005
R5948 DVDD.n20376 DVDD.n19834 4.5005
R5949 DVDD.n20420 DVDD.n20376 4.5005
R5950 DVDD.n19852 DVDD.n19841 4.5005
R5951 DVDD.n19852 DVDD.n19843 4.5005
R5952 DVDD.n19852 DVDD.n19840 4.5005
R5953 DVDD.n19852 DVDD.n19844 4.5005
R5954 DVDD.n19852 DVDD.n19839 4.5005
R5955 DVDD.n19852 DVDD.n19845 4.5005
R5956 DVDD.n19852 DVDD.n19838 4.5005
R5957 DVDD.n19852 DVDD.n19846 4.5005
R5958 DVDD.n19852 DVDD.n19837 4.5005
R5959 DVDD.n19852 DVDD.n19847 4.5005
R5960 DVDD.n19852 DVDD.n19836 4.5005
R5961 DVDD.n19852 DVDD.n19848 4.5005
R5962 DVDD.n19852 DVDD.n19835 4.5005
R5963 DVDD.n19852 DVDD.n19849 4.5005
R5964 DVDD.n19852 DVDD.n19834 4.5005
R5965 DVDD.n20420 DVDD.n19852 4.5005
R5966 DVDD.n20377 DVDD.n19841 4.5005
R5967 DVDD.n20377 DVDD.n19843 4.5005
R5968 DVDD.n20377 DVDD.n19840 4.5005
R5969 DVDD.n20377 DVDD.n19844 4.5005
R5970 DVDD.n20377 DVDD.n19839 4.5005
R5971 DVDD.n20377 DVDD.n19845 4.5005
R5972 DVDD.n20377 DVDD.n19838 4.5005
R5973 DVDD.n20377 DVDD.n19846 4.5005
R5974 DVDD.n20377 DVDD.n19837 4.5005
R5975 DVDD.n20377 DVDD.n19847 4.5005
R5976 DVDD.n20377 DVDD.n19836 4.5005
R5977 DVDD.n20377 DVDD.n19848 4.5005
R5978 DVDD.n20377 DVDD.n19835 4.5005
R5979 DVDD.n20377 DVDD.n19849 4.5005
R5980 DVDD.n20377 DVDD.n19834 4.5005
R5981 DVDD.n20420 DVDD.n20377 4.5005
R5982 DVDD.n19851 DVDD.n19841 4.5005
R5983 DVDD.n19851 DVDD.n19843 4.5005
R5984 DVDD.n19851 DVDD.n19840 4.5005
R5985 DVDD.n19851 DVDD.n19844 4.5005
R5986 DVDD.n19851 DVDD.n19839 4.5005
R5987 DVDD.n19851 DVDD.n19845 4.5005
R5988 DVDD.n19851 DVDD.n19838 4.5005
R5989 DVDD.n19851 DVDD.n19846 4.5005
R5990 DVDD.n19851 DVDD.n19837 4.5005
R5991 DVDD.n19851 DVDD.n19847 4.5005
R5992 DVDD.n19851 DVDD.n19836 4.5005
R5993 DVDD.n19851 DVDD.n19848 4.5005
R5994 DVDD.n19851 DVDD.n19835 4.5005
R5995 DVDD.n19851 DVDD.n19849 4.5005
R5996 DVDD.n19851 DVDD.n19834 4.5005
R5997 DVDD.n20420 DVDD.n19851 4.5005
R5998 DVDD.n20419 DVDD.n19841 4.5005
R5999 DVDD.n20419 DVDD.n19843 4.5005
R6000 DVDD.n20419 DVDD.n19840 4.5005
R6001 DVDD.n20419 DVDD.n19844 4.5005
R6002 DVDD.n20419 DVDD.n19839 4.5005
R6003 DVDD.n20419 DVDD.n19845 4.5005
R6004 DVDD.n20419 DVDD.n19838 4.5005
R6005 DVDD.n20419 DVDD.n19846 4.5005
R6006 DVDD.n20419 DVDD.n19837 4.5005
R6007 DVDD.n20419 DVDD.n19847 4.5005
R6008 DVDD.n20419 DVDD.n19836 4.5005
R6009 DVDD.n20419 DVDD.n19848 4.5005
R6010 DVDD.n20419 DVDD.n19835 4.5005
R6011 DVDD.n20419 DVDD.n19849 4.5005
R6012 DVDD.n20419 DVDD.n19834 4.5005
R6013 DVDD.n20420 DVDD.n20419 4.5005
R6014 DVDD.n20421 DVDD.n19841 4.5005
R6015 DVDD.n20421 DVDD.n19843 4.5005
R6016 DVDD.n20421 DVDD.n19840 4.5005
R6017 DVDD.n20421 DVDD.n19844 4.5005
R6018 DVDD.n20421 DVDD.n19839 4.5005
R6019 DVDD.n20421 DVDD.n19845 4.5005
R6020 DVDD.n20421 DVDD.n19838 4.5005
R6021 DVDD.n20421 DVDD.n19846 4.5005
R6022 DVDD.n20421 DVDD.n19837 4.5005
R6023 DVDD.n20421 DVDD.n19847 4.5005
R6024 DVDD.n20421 DVDD.n19836 4.5005
R6025 DVDD.n20421 DVDD.n19848 4.5005
R6026 DVDD.n20421 DVDD.n19835 4.5005
R6027 DVDD.n20421 DVDD.n19849 4.5005
R6028 DVDD.n20421 DVDD.n19834 4.5005
R6029 DVDD.n20421 DVDD.n20420 4.5005
R6030 DVDD.n19841 DVDD.n19832 4.5005
R6031 DVDD.n19843 DVDD.n19832 4.5005
R6032 DVDD.n19840 DVDD.n19832 4.5005
R6033 DVDD.n19844 DVDD.n19832 4.5005
R6034 DVDD.n19839 DVDD.n19832 4.5005
R6035 DVDD.n19845 DVDD.n19832 4.5005
R6036 DVDD.n19838 DVDD.n19832 4.5005
R6037 DVDD.n19846 DVDD.n19832 4.5005
R6038 DVDD.n19837 DVDD.n19832 4.5005
R6039 DVDD.n19847 DVDD.n19832 4.5005
R6040 DVDD.n19836 DVDD.n19832 4.5005
R6041 DVDD.n19848 DVDD.n19832 4.5005
R6042 DVDD.n19835 DVDD.n19832 4.5005
R6043 DVDD.n19849 DVDD.n19832 4.5005
R6044 DVDD.n19834 DVDD.n19832 4.5005
R6045 DVDD.n20420 DVDD.n19832 4.5005
R6046 DVDD.n18883 DVDD.n18871 4.5005
R6047 DVDD.n18875 DVDD.n18871 4.5005
R6048 DVDD.n18884 DVDD.n18871 4.5005
R6049 DVDD.n18874 DVDD.n18871 4.5005
R6050 DVDD.n18885 DVDD.n18871 4.5005
R6051 DVDD.n18873 DVDD.n18871 4.5005
R6052 DVDD.n18886 DVDD.n18871 4.5005
R6053 DVDD.n18872 DVDD.n18871 4.5005
R6054 DVDD.n20929 DVDD.n18871 4.5005
R6055 DVDD.n20930 DVDD.n18883 4.5005
R6056 DVDD.n20930 DVDD.n18875 4.5005
R6057 DVDD.n20930 DVDD.n18884 4.5005
R6058 DVDD.n20930 DVDD.n18874 4.5005
R6059 DVDD.n20930 DVDD.n18885 4.5005
R6060 DVDD.n20930 DVDD.n18873 4.5005
R6061 DVDD.n20930 DVDD.n18886 4.5005
R6062 DVDD.n20930 DVDD.n18872 4.5005
R6063 DVDD.n20930 DVDD.n20929 4.5005
R6064 DVDD.n4601 DVDD.n4244 4.5005
R6065 DVDD.n4256 DVDD.n4244 4.5005
R6066 DVDD.n4264 DVDD.n4244 4.5005
R6067 DVDD.n4255 DVDD.n4244 4.5005
R6068 DVDD.n4265 DVDD.n4244 4.5005
R6069 DVDD.n4254 DVDD.n4244 4.5005
R6070 DVDD.n4268 DVDD.n4244 4.5005
R6071 DVDD.n4253 DVDD.n4244 4.5005
R6072 DVDD.n4599 DVDD.n4244 4.5005
R6073 DVDD.n4599 DVDD.n4249 4.5005
R6074 DVDD.n4599 DVDD.n4243 4.5005
R6075 DVDD.n4253 DVDD.n4249 4.5005
R6076 DVDD.n4253 DVDD.n4243 4.5005
R6077 DVDD.n4268 DVDD.n4249 4.5005
R6078 DVDD.n4268 DVDD.n4243 4.5005
R6079 DVDD.n4254 DVDD.n4249 4.5005
R6080 DVDD.n4254 DVDD.n4243 4.5005
R6081 DVDD.n4265 DVDD.n4249 4.5005
R6082 DVDD.n4265 DVDD.n4243 4.5005
R6083 DVDD.n4255 DVDD.n4249 4.5005
R6084 DVDD.n4255 DVDD.n4243 4.5005
R6085 DVDD.n4264 DVDD.n4249 4.5005
R6086 DVDD.n4264 DVDD.n4243 4.5005
R6087 DVDD.n4256 DVDD.n4249 4.5005
R6088 DVDD.n4256 DVDD.n4243 4.5005
R6089 DVDD.n4601 DVDD.n4249 4.5005
R6090 DVDD.n4601 DVDD.n4243 4.5005
R6091 DVDD.n4599 DVDD.n4250 4.5005
R6092 DVDD.n4599 DVDD.n4241 4.5005
R6093 DVDD.n4253 DVDD.n4250 4.5005
R6094 DVDD.n4253 DVDD.n4241 4.5005
R6095 DVDD.n4268 DVDD.n4250 4.5005
R6096 DVDD.n4268 DVDD.n4241 4.5005
R6097 DVDD.n4254 DVDD.n4250 4.5005
R6098 DVDD.n4254 DVDD.n4241 4.5005
R6099 DVDD.n4265 DVDD.n4250 4.5005
R6100 DVDD.n4265 DVDD.n4241 4.5005
R6101 DVDD.n4255 DVDD.n4250 4.5005
R6102 DVDD.n4255 DVDD.n4241 4.5005
R6103 DVDD.n4264 DVDD.n4250 4.5005
R6104 DVDD.n4264 DVDD.n4241 4.5005
R6105 DVDD.n4256 DVDD.n4250 4.5005
R6106 DVDD.n4256 DVDD.n4241 4.5005
R6107 DVDD.n4601 DVDD.n4250 4.5005
R6108 DVDD.n4601 DVDD.n4241 4.5005
R6109 DVDD.n4599 DVDD.n4251 4.5005
R6110 DVDD.n4599 DVDD.n4240 4.5005
R6111 DVDD.n4253 DVDD.n4251 4.5005
R6112 DVDD.n4253 DVDD.n4240 4.5005
R6113 DVDD.n4268 DVDD.n4251 4.5005
R6114 DVDD.n4268 DVDD.n4240 4.5005
R6115 DVDD.n4254 DVDD.n4251 4.5005
R6116 DVDD.n4254 DVDD.n4240 4.5005
R6117 DVDD.n4265 DVDD.n4251 4.5005
R6118 DVDD.n4265 DVDD.n4240 4.5005
R6119 DVDD.n4255 DVDD.n4251 4.5005
R6120 DVDD.n4255 DVDD.n4240 4.5005
R6121 DVDD.n4264 DVDD.n4251 4.5005
R6122 DVDD.n4264 DVDD.n4240 4.5005
R6123 DVDD.n4256 DVDD.n4251 4.5005
R6124 DVDD.n4256 DVDD.n4240 4.5005
R6125 DVDD.n4601 DVDD.n4251 4.5005
R6126 DVDD.n4601 DVDD.n4240 4.5005
R6127 DVDD.n4601 DVDD.n4600 4.5005
R6128 DVDD.n4600 DVDD.n4256 4.5005
R6129 DVDD.n4600 DVDD.n4264 4.5005
R6130 DVDD.n4600 DVDD.n4255 4.5005
R6131 DVDD.n4600 DVDD.n4265 4.5005
R6132 DVDD.n4600 DVDD.n4254 4.5005
R6133 DVDD.n4600 DVDD.n4268 4.5005
R6134 DVDD.n4600 DVDD.n4253 4.5005
R6135 DVDD.n4600 DVDD.n4599 4.5005
R6136 DVDD.n2412 DVDD.n2385 4.5005
R6137 DVDD.n16370 DVDD.n2412 4.5005
R6138 DVDD.n2437 DVDD.n2412 4.5005
R6139 DVDD.n2477 DVDD.n2412 4.5005
R6140 DVDD.n2436 DVDD.n2412 4.5005
R6141 DVDD.n2478 DVDD.n2412 4.5005
R6142 DVDD.n2435 DVDD.n2412 4.5005
R6143 DVDD.n2479 DVDD.n2412 4.5005
R6144 DVDD.n2434 DVDD.n2412 4.5005
R6145 DVDD.n2480 DVDD.n2412 4.5005
R6146 DVDD.n2433 DVDD.n2412 4.5005
R6147 DVDD.n2481 DVDD.n2412 4.5005
R6148 DVDD.n2482 DVDD.n2412 4.5005
R6149 DVDD.n2424 DVDD.n2412 4.5005
R6150 DVDD.n16368 DVDD.n2412 4.5005
R6151 DVDD.n2390 DVDD.n2385 4.5005
R6152 DVDD.n16370 DVDD.n2390 4.5005
R6153 DVDD.n2437 DVDD.n2390 4.5005
R6154 DVDD.n2477 DVDD.n2390 4.5005
R6155 DVDD.n2436 DVDD.n2390 4.5005
R6156 DVDD.n2478 DVDD.n2390 4.5005
R6157 DVDD.n2435 DVDD.n2390 4.5005
R6158 DVDD.n2479 DVDD.n2390 4.5005
R6159 DVDD.n2434 DVDD.n2390 4.5005
R6160 DVDD.n2480 DVDD.n2390 4.5005
R6161 DVDD.n2433 DVDD.n2390 4.5005
R6162 DVDD.n2481 DVDD.n2390 4.5005
R6163 DVDD.n2432 DVDD.n2390 4.5005
R6164 DVDD.n2482 DVDD.n2390 4.5005
R6165 DVDD.n2424 DVDD.n2390 4.5005
R6166 DVDD.n16368 DVDD.n2390 4.5005
R6167 DVDD.n16369 DVDD.n2385 4.5005
R6168 DVDD.n16370 DVDD.n16369 4.5005
R6169 DVDD.n16369 DVDD.n2437 4.5005
R6170 DVDD.n16369 DVDD.n2477 4.5005
R6171 DVDD.n16369 DVDD.n2436 4.5005
R6172 DVDD.n16369 DVDD.n2478 4.5005
R6173 DVDD.n16369 DVDD.n2435 4.5005
R6174 DVDD.n16369 DVDD.n2479 4.5005
R6175 DVDD.n16369 DVDD.n2434 4.5005
R6176 DVDD.n16369 DVDD.n2480 4.5005
R6177 DVDD.n16369 DVDD.n2433 4.5005
R6178 DVDD.n16369 DVDD.n2481 4.5005
R6179 DVDD.n16369 DVDD.n2432 4.5005
R6180 DVDD.n16369 DVDD.n2482 4.5005
R6181 DVDD.n16369 DVDD.n2424 4.5005
R6182 DVDD.n16369 DVDD.n16368 4.5005
R6183 DVDD.n2962 DVDD.n2955 4.5005
R6184 DVDD.n2965 DVDD.n2955 4.5005
R6185 DVDD.n2961 DVDD.n2955 4.5005
R6186 DVDD.n2966 DVDD.n2955 4.5005
R6187 DVDD.n2960 DVDD.n2955 4.5005
R6188 DVDD.n2967 DVDD.n2955 4.5005
R6189 DVDD.n2959 DVDD.n2955 4.5005
R6190 DVDD.n2968 DVDD.n2955 4.5005
R6191 DVDD.n2958 DVDD.n2955 4.5005
R6192 DVDD.n2970 DVDD.n2955 4.5005
R6193 DVDD.n2957 DVDD.n2955 4.5005
R6194 DVDD.n2971 DVDD.n2955 4.5005
R6195 DVDD.n16182 DVDD.n2955 4.5005
R6196 DVDD.n2955 DVDD.n2924 4.5005
R6197 DVDD.n16184 DVDD.n2955 4.5005
R6198 DVDD.n2962 DVDD.n2925 4.5005
R6199 DVDD.n2965 DVDD.n2925 4.5005
R6200 DVDD.n2961 DVDD.n2925 4.5005
R6201 DVDD.n2966 DVDD.n2925 4.5005
R6202 DVDD.n2960 DVDD.n2925 4.5005
R6203 DVDD.n2967 DVDD.n2925 4.5005
R6204 DVDD.n2959 DVDD.n2925 4.5005
R6205 DVDD.n2968 DVDD.n2925 4.5005
R6206 DVDD.n2958 DVDD.n2925 4.5005
R6207 DVDD.n2970 DVDD.n2925 4.5005
R6208 DVDD.n2957 DVDD.n2925 4.5005
R6209 DVDD.n2971 DVDD.n2925 4.5005
R6210 DVDD.n16182 DVDD.n2925 4.5005
R6211 DVDD.n2925 DVDD.n2924 4.5005
R6212 DVDD.n16184 DVDD.n2925 4.5005
R6213 DVDD.n16183 DVDD.n2962 4.5005
R6214 DVDD.n16183 DVDD.n2965 4.5005
R6215 DVDD.n16183 DVDD.n2961 4.5005
R6216 DVDD.n16183 DVDD.n2966 4.5005
R6217 DVDD.n16183 DVDD.n2960 4.5005
R6218 DVDD.n16183 DVDD.n2967 4.5005
R6219 DVDD.n16183 DVDD.n2959 4.5005
R6220 DVDD.n16183 DVDD.n2968 4.5005
R6221 DVDD.n16183 DVDD.n2958 4.5005
R6222 DVDD.n16183 DVDD.n2970 4.5005
R6223 DVDD.n16183 DVDD.n2957 4.5005
R6224 DVDD.n16183 DVDD.n2971 4.5005
R6225 DVDD.n16183 DVDD.n16182 4.5005
R6226 DVDD.n16183 DVDD.n2924 4.5005
R6227 DVDD.n16184 DVDD.n16183 4.5005
R6228 DVDD.n10057 DVDD.n9745 4.5005
R6229 DVDD.n9956 DVDD.n9745 4.5005
R6230 DVDD.n9755 DVDD.n9745 4.5005
R6231 DVDD.n9957 DVDD.n9745 4.5005
R6232 DVDD.n9754 DVDD.n9745 4.5005
R6233 DVDD.n9958 DVDD.n9745 4.5005
R6234 DVDD.n9753 DVDD.n9745 4.5005
R6235 DVDD.n9959 DVDD.n9745 4.5005
R6236 DVDD.n9752 DVDD.n9745 4.5005
R6237 DVDD.n9961 DVDD.n9745 4.5005
R6238 DVDD.n9751 DVDD.n9745 4.5005
R6239 DVDD.n9962 DVDD.n9745 4.5005
R6240 DVDD.n10001 DVDD.n9745 4.5005
R6241 DVDD.n9963 DVDD.n9745 4.5005
R6242 DVDD.n10055 DVDD.n9745 4.5005
R6243 DVDD.n10057 DVDD.n9733 4.5005
R6244 DVDD.n9956 DVDD.n9733 4.5005
R6245 DVDD.n9755 DVDD.n9733 4.5005
R6246 DVDD.n9957 DVDD.n9733 4.5005
R6247 DVDD.n9754 DVDD.n9733 4.5005
R6248 DVDD.n9958 DVDD.n9733 4.5005
R6249 DVDD.n9753 DVDD.n9733 4.5005
R6250 DVDD.n9959 DVDD.n9733 4.5005
R6251 DVDD.n9752 DVDD.n9733 4.5005
R6252 DVDD.n9961 DVDD.n9733 4.5005
R6253 DVDD.n9751 DVDD.n9733 4.5005
R6254 DVDD.n9962 DVDD.n9733 4.5005
R6255 DVDD.n9963 DVDD.n9733 4.5005
R6256 DVDD.n9750 DVDD.n9733 4.5005
R6257 DVDD.n10055 DVDD.n9733 4.5005
R6258 DVDD.n10057 DVDD.n10056 4.5005
R6259 DVDD.n10056 DVDD.n9956 4.5005
R6260 DVDD.n10056 DVDD.n9755 4.5005
R6261 DVDD.n10056 DVDD.n9957 4.5005
R6262 DVDD.n10056 DVDD.n9754 4.5005
R6263 DVDD.n10056 DVDD.n9958 4.5005
R6264 DVDD.n10056 DVDD.n9753 4.5005
R6265 DVDD.n10056 DVDD.n9959 4.5005
R6266 DVDD.n10056 DVDD.n9752 4.5005
R6267 DVDD.n10056 DVDD.n9961 4.5005
R6268 DVDD.n10056 DVDD.n9751 4.5005
R6269 DVDD.n10056 DVDD.n9962 4.5005
R6270 DVDD.n10056 DVDD.n9963 4.5005
R6271 DVDD.n10056 DVDD.n9750 4.5005
R6272 DVDD.n10056 DVDD.n10055 4.5005
R6273 DVDD.n21083 DVDD.n18751 4.5005
R6274 DVDD.n21083 DVDD.n21082 4.5005
R6275 DVDD.n21082 DVDD.n18735 4.5005
R6276 DVDD.n21081 DVDD.n18751 4.5005
R6277 DVDD.n21081 DVDD.n21068 4.5005
R6278 DVDD.n21081 DVDD.n21066 4.5005
R6279 DVDD.n21081 DVDD.n21070 4.5005
R6280 DVDD.n21081 DVDD.n21065 4.5005
R6281 DVDD.n21081 DVDD.n21072 4.5005
R6282 DVDD.n21081 DVDD.n21064 4.5005
R6283 DVDD.n21081 DVDD.n21074 4.5005
R6284 DVDD.n21081 DVDD.n21063 4.5005
R6285 DVDD.n21081 DVDD.n21076 4.5005
R6286 DVDD.n21081 DVDD.n21062 4.5005
R6287 DVDD.n21081 DVDD.n21078 4.5005
R6288 DVDD.n21081 DVDD.n21061 4.5005
R6289 DVDD.n21081 DVDD.n21080 4.5005
R6290 DVDD.n21082 DVDD.n21081 4.5005
R6291 DVDD.n21055 DVDD.n21054 4.5005
R6292 DVDD.n21056 DVDD.n21055 4.5005
R6293 DVDD.n21058 DVDD.n21055 4.5005
R6294 DVDD.n21059 DVDD.n21058 4.5005
R6295 DVDD.n19123 DVDD.n19122 4.5005
R6296 DVDD.n19123 DVDD.n18830 4.5005
R6297 DVDD.n20950 DVDD.n18866 4.5005
R6298 DVDD.n20966 DVDD.n18866 4.5005
R6299 DVDD.n20535 DVDD.n20483 4.5005
R6300 DVDD.n20535 DVDD.n20485 4.5005
R6301 DVDD.n20535 DVDD.n20534 4.5005
R6302 DVDD.n20534 DVDD.n19129 4.5005
R6303 DVDD.n20538 DVDD.n19773 4.5005
R6304 DVDD.n20538 DVDD.n20537 4.5005
R6305 DVDD.n20539 DVDD.n20538 4.5005
R6306 DVDD.n20537 DVDD.n19788 4.5005
R6307 DVDD.n20539 DVDD.n19788 4.5005
R6308 DVDD.n20540 DVDD.n19773 4.5005
R6309 DVDD.n20540 DVDD.n19774 4.5005
R6310 DVDD.n20540 DVDD.n19772 4.5005
R6311 DVDD.n20540 DVDD.n19775 4.5005
R6312 DVDD.n20540 DVDD.n19771 4.5005
R6313 DVDD.n20540 DVDD.n19776 4.5005
R6314 DVDD.n20540 DVDD.n19770 4.5005
R6315 DVDD.n20540 DVDD.n19777 4.5005
R6316 DVDD.n20540 DVDD.n19769 4.5005
R6317 DVDD.n20540 DVDD.n19778 4.5005
R6318 DVDD.n20540 DVDD.n19768 4.5005
R6319 DVDD.n20540 DVDD.n19779 4.5005
R6320 DVDD.n20540 DVDD.n20539 4.5005
R6321 DVDD.n10094 DVDD.n9620 4.5005
R6322 DVDD.n10094 DVDD.n9621 4.5005
R6323 DVDD.n10094 DVDD.n9619 4.5005
R6324 DVDD.n10094 DVDD.n9622 4.5005
R6325 DVDD.n10094 DVDD.n9617 4.5005
R6326 DVDD.n10094 DVDD.n9623 4.5005
R6327 DVDD.n10094 DVDD.n9616 4.5005
R6328 DVDD.n10094 DVDD.n9624 4.5005
R6329 DVDD.n10094 DVDD.n9615 4.5005
R6330 DVDD.n10094 DVDD.n9625 4.5005
R6331 DVDD.n10094 DVDD.n9613 4.5005
R6332 DVDD.n10094 DVDD.n10093 4.5005
R6333 DVDD.n9631 DVDD.n9620 4.5005
R6334 DVDD.n9631 DVDD.n9621 4.5005
R6335 DVDD.n9631 DVDD.n9619 4.5005
R6336 DVDD.n9642 DVDD.n9631 4.5005
R6337 DVDD.n9641 DVDD.n9631 4.5005
R6338 DVDD.n9631 DVDD.n9622 4.5005
R6339 DVDD.n9631 DVDD.n9617 4.5005
R6340 DVDD.n9631 DVDD.n9623 4.5005
R6341 DVDD.n9631 DVDD.n9616 4.5005
R6342 DVDD.n9631 DVDD.n9624 4.5005
R6343 DVDD.n9631 DVDD.n9615 4.5005
R6344 DVDD.n10091 DVDD.n9631 4.5005
R6345 DVDD.n9631 DVDD.n9625 4.5005
R6346 DVDD.n10093 DVDD.n9631 4.5005
R6347 DVDD.n9634 DVDD.n9620 4.5005
R6348 DVDD.n9634 DVDD.n9621 4.5005
R6349 DVDD.n9634 DVDD.n9619 4.5005
R6350 DVDD.n9642 DVDD.n9634 4.5005
R6351 DVDD.n9641 DVDD.n9634 4.5005
R6352 DVDD.n9634 DVDD.n9622 4.5005
R6353 DVDD.n9634 DVDD.n9617 4.5005
R6354 DVDD.n9634 DVDD.n9623 4.5005
R6355 DVDD.n9634 DVDD.n9616 4.5005
R6356 DVDD.n9634 DVDD.n9624 4.5005
R6357 DVDD.n9634 DVDD.n9615 4.5005
R6358 DVDD.n10091 DVDD.n9634 4.5005
R6359 DVDD.n9634 DVDD.n9625 4.5005
R6360 DVDD.n10093 DVDD.n9634 4.5005
R6361 DVDD.n9630 DVDD.n9620 4.5005
R6362 DVDD.n9630 DVDD.n9621 4.5005
R6363 DVDD.n9630 DVDD.n9619 4.5005
R6364 DVDD.n9642 DVDD.n9630 4.5005
R6365 DVDD.n9641 DVDD.n9630 4.5005
R6366 DVDD.n9630 DVDD.n9622 4.5005
R6367 DVDD.n9630 DVDD.n9617 4.5005
R6368 DVDD.n9630 DVDD.n9623 4.5005
R6369 DVDD.n9630 DVDD.n9616 4.5005
R6370 DVDD.n9630 DVDD.n9624 4.5005
R6371 DVDD.n9630 DVDD.n9615 4.5005
R6372 DVDD.n10091 DVDD.n9630 4.5005
R6373 DVDD.n9630 DVDD.n9625 4.5005
R6374 DVDD.n9630 DVDD.n9613 4.5005
R6375 DVDD.n10093 DVDD.n9630 4.5005
R6376 DVDD.n9636 DVDD.n9620 4.5005
R6377 DVDD.n9636 DVDD.n9621 4.5005
R6378 DVDD.n9636 DVDD.n9619 4.5005
R6379 DVDD.n9642 DVDD.n9636 4.5005
R6380 DVDD.n9641 DVDD.n9636 4.5005
R6381 DVDD.n9636 DVDD.n9622 4.5005
R6382 DVDD.n9636 DVDD.n9617 4.5005
R6383 DVDD.n9636 DVDD.n9623 4.5005
R6384 DVDD.n9636 DVDD.n9616 4.5005
R6385 DVDD.n9636 DVDD.n9624 4.5005
R6386 DVDD.n9636 DVDD.n9615 4.5005
R6387 DVDD.n10091 DVDD.n9636 4.5005
R6388 DVDD.n9636 DVDD.n9625 4.5005
R6389 DVDD.n10093 DVDD.n9636 4.5005
R6390 DVDD.n9629 DVDD.n9620 4.5005
R6391 DVDD.n9629 DVDD.n9621 4.5005
R6392 DVDD.n9629 DVDD.n9619 4.5005
R6393 DVDD.n9642 DVDD.n9629 4.5005
R6394 DVDD.n9641 DVDD.n9629 4.5005
R6395 DVDD.n9629 DVDD.n9622 4.5005
R6396 DVDD.n9629 DVDD.n9617 4.5005
R6397 DVDD.n9629 DVDD.n9623 4.5005
R6398 DVDD.n9629 DVDD.n9616 4.5005
R6399 DVDD.n9629 DVDD.n9624 4.5005
R6400 DVDD.n9629 DVDD.n9615 4.5005
R6401 DVDD.n10091 DVDD.n9629 4.5005
R6402 DVDD.n9629 DVDD.n9625 4.5005
R6403 DVDD.n10093 DVDD.n9629 4.5005
R6404 DVDD.n9637 DVDD.n9620 4.5005
R6405 DVDD.n9637 DVDD.n9621 4.5005
R6406 DVDD.n9637 DVDD.n9619 4.5005
R6407 DVDD.n9642 DVDD.n9637 4.5005
R6408 DVDD.n9641 DVDD.n9637 4.5005
R6409 DVDD.n9637 DVDD.n9622 4.5005
R6410 DVDD.n9637 DVDD.n9617 4.5005
R6411 DVDD.n9637 DVDD.n9623 4.5005
R6412 DVDD.n9637 DVDD.n9616 4.5005
R6413 DVDD.n9637 DVDD.n9624 4.5005
R6414 DVDD.n9637 DVDD.n9615 4.5005
R6415 DVDD.n10091 DVDD.n9637 4.5005
R6416 DVDD.n9637 DVDD.n9625 4.5005
R6417 DVDD.n9637 DVDD.n9613 4.5005
R6418 DVDD.n10093 DVDD.n9637 4.5005
R6419 DVDD.n9628 DVDD.n9620 4.5005
R6420 DVDD.n9628 DVDD.n9621 4.5005
R6421 DVDD.n9628 DVDD.n9619 4.5005
R6422 DVDD.n9642 DVDD.n9628 4.5005
R6423 DVDD.n9641 DVDD.n9628 4.5005
R6424 DVDD.n9628 DVDD.n9622 4.5005
R6425 DVDD.n9628 DVDD.n9617 4.5005
R6426 DVDD.n9628 DVDD.n9623 4.5005
R6427 DVDD.n9628 DVDD.n9616 4.5005
R6428 DVDD.n9628 DVDD.n9624 4.5005
R6429 DVDD.n9628 DVDD.n9615 4.5005
R6430 DVDD.n10091 DVDD.n9628 4.5005
R6431 DVDD.n9648 DVDD.n9628 4.5005
R6432 DVDD.n9628 DVDD.n9625 4.5005
R6433 DVDD.n10093 DVDD.n9628 4.5005
R6434 DVDD.n9778 DVDD.n3080 4.5005
R6435 DVDD.n9778 DVDD.n3082 4.5005
R6436 DVDD.n9778 DVDD.n3079 4.5005
R6437 DVDD.n9778 DVDD.n3084 4.5005
R6438 DVDD.n9778 DVDD.n3077 4.5005
R6439 DVDD.n9778 DVDD.n3085 4.5005
R6440 DVDD.n9778 DVDD.n3076 4.5005
R6441 DVDD.n9778 DVDD.n3086 4.5005
R6442 DVDD.n9778 DVDD.n3075 4.5005
R6443 DVDD.n9778 DVDD.n3057 4.5005
R6444 DVDD.n9778 DVDD.n3053 4.5005
R6445 DVDD.n3096 DVDD.n3080 4.5005
R6446 DVDD.n3096 DVDD.n3082 4.5005
R6447 DVDD.n3096 DVDD.n3079 4.5005
R6448 DVDD.n3096 DVDD.n3083 4.5005
R6449 DVDD.n3096 DVDD.n3078 4.5005
R6450 DVDD.n3096 DVDD.n3084 4.5005
R6451 DVDD.n3096 DVDD.n3077 4.5005
R6452 DVDD.n3096 DVDD.n3085 4.5005
R6453 DVDD.n3096 DVDD.n3076 4.5005
R6454 DVDD.n3096 DVDD.n3086 4.5005
R6455 DVDD.n3096 DVDD.n3075 4.5005
R6456 DVDD.n16083 DVDD.n3096 4.5005
R6457 DVDD.n3096 DVDD.n3057 4.5005
R6458 DVDD.n3096 DVDD.n3053 4.5005
R6459 DVDD.n3080 DVDD.n3066 4.5005
R6460 DVDD.n3082 DVDD.n3066 4.5005
R6461 DVDD.n3079 DVDD.n3066 4.5005
R6462 DVDD.n3083 DVDD.n3066 4.5005
R6463 DVDD.n3078 DVDD.n3066 4.5005
R6464 DVDD.n3084 DVDD.n3066 4.5005
R6465 DVDD.n3077 DVDD.n3066 4.5005
R6466 DVDD.n3085 DVDD.n3066 4.5005
R6467 DVDD.n3076 DVDD.n3066 4.5005
R6468 DVDD.n3086 DVDD.n3066 4.5005
R6469 DVDD.n3075 DVDD.n3066 4.5005
R6470 DVDD.n16083 DVDD.n3066 4.5005
R6471 DVDD.n3066 DVDD.n3057 4.5005
R6472 DVDD.n16085 DVDD.n3066 4.5005
R6473 DVDD.n3066 DVDD.n3053 4.5005
R6474 DVDD.n3097 DVDD.n3080 4.5005
R6475 DVDD.n3097 DVDD.n3082 4.5005
R6476 DVDD.n3097 DVDD.n3079 4.5005
R6477 DVDD.n3097 DVDD.n3083 4.5005
R6478 DVDD.n3097 DVDD.n3078 4.5005
R6479 DVDD.n3097 DVDD.n3084 4.5005
R6480 DVDD.n3097 DVDD.n3077 4.5005
R6481 DVDD.n3097 DVDD.n3085 4.5005
R6482 DVDD.n3097 DVDD.n3076 4.5005
R6483 DVDD.n3097 DVDD.n3086 4.5005
R6484 DVDD.n3097 DVDD.n3075 4.5005
R6485 DVDD.n16083 DVDD.n3097 4.5005
R6486 DVDD.n3097 DVDD.n3057 4.5005
R6487 DVDD.n3097 DVDD.n3053 4.5005
R6488 DVDD.n3094 DVDD.n3080 4.5005
R6489 DVDD.n3094 DVDD.n3082 4.5005
R6490 DVDD.n3094 DVDD.n3079 4.5005
R6491 DVDD.n3094 DVDD.n3083 4.5005
R6492 DVDD.n3094 DVDD.n3078 4.5005
R6493 DVDD.n3094 DVDD.n3084 4.5005
R6494 DVDD.n3094 DVDD.n3077 4.5005
R6495 DVDD.n3094 DVDD.n3085 4.5005
R6496 DVDD.n3094 DVDD.n3076 4.5005
R6497 DVDD.n3094 DVDD.n3086 4.5005
R6498 DVDD.n3094 DVDD.n3075 4.5005
R6499 DVDD.n16083 DVDD.n3094 4.5005
R6500 DVDD.n3094 DVDD.n3057 4.5005
R6501 DVDD.n3094 DVDD.n3053 4.5005
R6502 DVDD.n3080 DVDD.n3070 4.5005
R6503 DVDD.n3082 DVDD.n3070 4.5005
R6504 DVDD.n3079 DVDD.n3070 4.5005
R6505 DVDD.n3083 DVDD.n3070 4.5005
R6506 DVDD.n3078 DVDD.n3070 4.5005
R6507 DVDD.n3084 DVDD.n3070 4.5005
R6508 DVDD.n3077 DVDD.n3070 4.5005
R6509 DVDD.n3085 DVDD.n3070 4.5005
R6510 DVDD.n3076 DVDD.n3070 4.5005
R6511 DVDD.n3086 DVDD.n3070 4.5005
R6512 DVDD.n3075 DVDD.n3070 4.5005
R6513 DVDD.n16083 DVDD.n3070 4.5005
R6514 DVDD.n3070 DVDD.n3057 4.5005
R6515 DVDD.n16085 DVDD.n3070 4.5005
R6516 DVDD.n3070 DVDD.n3053 4.5005
R6517 DVDD.n3093 DVDD.n3080 4.5005
R6518 DVDD.n3093 DVDD.n3082 4.5005
R6519 DVDD.n3093 DVDD.n3079 4.5005
R6520 DVDD.n3093 DVDD.n3083 4.5005
R6521 DVDD.n3093 DVDD.n3078 4.5005
R6522 DVDD.n3093 DVDD.n3084 4.5005
R6523 DVDD.n3093 DVDD.n3077 4.5005
R6524 DVDD.n3093 DVDD.n3085 4.5005
R6525 DVDD.n3093 DVDD.n3076 4.5005
R6526 DVDD.n3093 DVDD.n3086 4.5005
R6527 DVDD.n3093 DVDD.n3075 4.5005
R6528 DVDD.n16083 DVDD.n3093 4.5005
R6529 DVDD.n3093 DVDD.n3057 4.5005
R6530 DVDD.n3093 DVDD.n3053 4.5005
R6531 DVDD.n3098 DVDD.n3080 4.5005
R6532 DVDD.n3098 DVDD.n3082 4.5005
R6533 DVDD.n3098 DVDD.n3079 4.5005
R6534 DVDD.n3098 DVDD.n3083 4.5005
R6535 DVDD.n3098 DVDD.n3078 4.5005
R6536 DVDD.n3098 DVDD.n3084 4.5005
R6537 DVDD.n3098 DVDD.n3077 4.5005
R6538 DVDD.n3098 DVDD.n3085 4.5005
R6539 DVDD.n3098 DVDD.n3076 4.5005
R6540 DVDD.n3098 DVDD.n3086 4.5005
R6541 DVDD.n3098 DVDD.n3075 4.5005
R6542 DVDD.n16083 DVDD.n3098 4.5005
R6543 DVDD.n3098 DVDD.n3057 4.5005
R6544 DVDD.n3098 DVDD.n3053 4.5005
R6545 DVDD.n3080 DVDD.n3064 4.5005
R6546 DVDD.n3082 DVDD.n3064 4.5005
R6547 DVDD.n3079 DVDD.n3064 4.5005
R6548 DVDD.n3083 DVDD.n3064 4.5005
R6549 DVDD.n3078 DVDD.n3064 4.5005
R6550 DVDD.n3084 DVDD.n3064 4.5005
R6551 DVDD.n3077 DVDD.n3064 4.5005
R6552 DVDD.n3085 DVDD.n3064 4.5005
R6553 DVDD.n3076 DVDD.n3064 4.5005
R6554 DVDD.n3086 DVDD.n3064 4.5005
R6555 DVDD.n3075 DVDD.n3064 4.5005
R6556 DVDD.n16083 DVDD.n3064 4.5005
R6557 DVDD.n3064 DVDD.n3057 4.5005
R6558 DVDD.n16085 DVDD.n3064 4.5005
R6559 DVDD.n3064 DVDD.n3053 4.5005
R6560 DVDD.n3099 DVDD.n3080 4.5005
R6561 DVDD.n3099 DVDD.n3082 4.5005
R6562 DVDD.n3099 DVDD.n3079 4.5005
R6563 DVDD.n3099 DVDD.n3083 4.5005
R6564 DVDD.n3099 DVDD.n3078 4.5005
R6565 DVDD.n3099 DVDD.n3084 4.5005
R6566 DVDD.n3099 DVDD.n3077 4.5005
R6567 DVDD.n3099 DVDD.n3085 4.5005
R6568 DVDD.n3099 DVDD.n3076 4.5005
R6569 DVDD.n3099 DVDD.n3086 4.5005
R6570 DVDD.n3099 DVDD.n3075 4.5005
R6571 DVDD.n16083 DVDD.n3099 4.5005
R6572 DVDD.n3099 DVDD.n3057 4.5005
R6573 DVDD.n3099 DVDD.n3053 4.5005
R6574 DVDD.n3092 DVDD.n3080 4.5005
R6575 DVDD.n3092 DVDD.n3082 4.5005
R6576 DVDD.n3092 DVDD.n3079 4.5005
R6577 DVDD.n3092 DVDD.n3083 4.5005
R6578 DVDD.n3092 DVDD.n3078 4.5005
R6579 DVDD.n3092 DVDD.n3084 4.5005
R6580 DVDD.n3092 DVDD.n3077 4.5005
R6581 DVDD.n3092 DVDD.n3085 4.5005
R6582 DVDD.n3092 DVDD.n3076 4.5005
R6583 DVDD.n3092 DVDD.n3086 4.5005
R6584 DVDD.n3092 DVDD.n3075 4.5005
R6585 DVDD.n16083 DVDD.n3092 4.5005
R6586 DVDD.n3092 DVDD.n3057 4.5005
R6587 DVDD.n3092 DVDD.n3053 4.5005
R6588 DVDD.n3080 DVDD.n3072 4.5005
R6589 DVDD.n3082 DVDD.n3072 4.5005
R6590 DVDD.n3079 DVDD.n3072 4.5005
R6591 DVDD.n3083 DVDD.n3072 4.5005
R6592 DVDD.n3078 DVDD.n3072 4.5005
R6593 DVDD.n3084 DVDD.n3072 4.5005
R6594 DVDD.n3077 DVDD.n3072 4.5005
R6595 DVDD.n3085 DVDD.n3072 4.5005
R6596 DVDD.n3076 DVDD.n3072 4.5005
R6597 DVDD.n3086 DVDD.n3072 4.5005
R6598 DVDD.n3075 DVDD.n3072 4.5005
R6599 DVDD.n16083 DVDD.n3072 4.5005
R6600 DVDD.n3072 DVDD.n3057 4.5005
R6601 DVDD.n16085 DVDD.n3072 4.5005
R6602 DVDD.n3072 DVDD.n3053 4.5005
R6603 DVDD.n3091 DVDD.n3080 4.5005
R6604 DVDD.n3091 DVDD.n3082 4.5005
R6605 DVDD.n3091 DVDD.n3079 4.5005
R6606 DVDD.n3091 DVDD.n3083 4.5005
R6607 DVDD.n3091 DVDD.n3078 4.5005
R6608 DVDD.n3091 DVDD.n3084 4.5005
R6609 DVDD.n3091 DVDD.n3077 4.5005
R6610 DVDD.n3091 DVDD.n3085 4.5005
R6611 DVDD.n3091 DVDD.n3076 4.5005
R6612 DVDD.n3091 DVDD.n3086 4.5005
R6613 DVDD.n3091 DVDD.n3075 4.5005
R6614 DVDD.n16083 DVDD.n3091 4.5005
R6615 DVDD.n16081 DVDD.n3091 4.5005
R6616 DVDD.n3091 DVDD.n3057 4.5005
R6617 DVDD.n3091 DVDD.n3053 4.5005
R6618 DVDD.n3100 DVDD.n3080 4.5005
R6619 DVDD.n3100 DVDD.n3082 4.5005
R6620 DVDD.n3100 DVDD.n3079 4.5005
R6621 DVDD.n3100 DVDD.n3083 4.5005
R6622 DVDD.n3100 DVDD.n3078 4.5005
R6623 DVDD.n3100 DVDD.n3084 4.5005
R6624 DVDD.n3100 DVDD.n3077 4.5005
R6625 DVDD.n3100 DVDD.n3085 4.5005
R6626 DVDD.n3100 DVDD.n3076 4.5005
R6627 DVDD.n3100 DVDD.n3086 4.5005
R6628 DVDD.n3100 DVDD.n3075 4.5005
R6629 DVDD.n16083 DVDD.n3100 4.5005
R6630 DVDD.n3100 DVDD.n3057 4.5005
R6631 DVDD.n3100 DVDD.n3053 4.5005
R6632 DVDD.n3090 DVDD.n3080 4.5005
R6633 DVDD.n3090 DVDD.n3082 4.5005
R6634 DVDD.n3090 DVDD.n3079 4.5005
R6635 DVDD.n3090 DVDD.n3083 4.5005
R6636 DVDD.n3090 DVDD.n3078 4.5005
R6637 DVDD.n3090 DVDD.n3084 4.5005
R6638 DVDD.n3090 DVDD.n3077 4.5005
R6639 DVDD.n3090 DVDD.n3085 4.5005
R6640 DVDD.n3090 DVDD.n3076 4.5005
R6641 DVDD.n3090 DVDD.n3086 4.5005
R6642 DVDD.n3090 DVDD.n3075 4.5005
R6643 DVDD.n16083 DVDD.n3090 4.5005
R6644 DVDD.n3090 DVDD.n3057 4.5005
R6645 DVDD.n3090 DVDD.n3053 4.5005
R6646 DVDD.n3101 DVDD.n3080 4.5005
R6647 DVDD.n3101 DVDD.n3082 4.5005
R6648 DVDD.n3101 DVDD.n3079 4.5005
R6649 DVDD.n3101 DVDD.n3083 4.5005
R6650 DVDD.n3101 DVDD.n3078 4.5005
R6651 DVDD.n3101 DVDD.n3084 4.5005
R6652 DVDD.n3101 DVDD.n3077 4.5005
R6653 DVDD.n3101 DVDD.n3085 4.5005
R6654 DVDD.n3101 DVDD.n3076 4.5005
R6655 DVDD.n3101 DVDD.n3086 4.5005
R6656 DVDD.n3101 DVDD.n3075 4.5005
R6657 DVDD.n16083 DVDD.n3101 4.5005
R6658 DVDD.n16081 DVDD.n3101 4.5005
R6659 DVDD.n3101 DVDD.n3057 4.5005
R6660 DVDD.n3101 DVDD.n3053 4.5005
R6661 DVDD.n3089 DVDD.n3080 4.5005
R6662 DVDD.n3089 DVDD.n3082 4.5005
R6663 DVDD.n3089 DVDD.n3079 4.5005
R6664 DVDD.n3089 DVDD.n3083 4.5005
R6665 DVDD.n3089 DVDD.n3078 4.5005
R6666 DVDD.n3089 DVDD.n3084 4.5005
R6667 DVDD.n3089 DVDD.n3077 4.5005
R6668 DVDD.n3089 DVDD.n3085 4.5005
R6669 DVDD.n3089 DVDD.n3076 4.5005
R6670 DVDD.n3089 DVDD.n3086 4.5005
R6671 DVDD.n3089 DVDD.n3075 4.5005
R6672 DVDD.n16083 DVDD.n3089 4.5005
R6673 DVDD.n16081 DVDD.n3089 4.5005
R6674 DVDD.n3089 DVDD.n3057 4.5005
R6675 DVDD.n3089 DVDD.n3053 4.5005
R6676 DVDD.n3102 DVDD.n3080 4.5005
R6677 DVDD.n3102 DVDD.n3082 4.5005
R6678 DVDD.n3102 DVDD.n3079 4.5005
R6679 DVDD.n3102 DVDD.n3083 4.5005
R6680 DVDD.n3102 DVDD.n3078 4.5005
R6681 DVDD.n3102 DVDD.n3084 4.5005
R6682 DVDD.n3102 DVDD.n3077 4.5005
R6683 DVDD.n3102 DVDD.n3085 4.5005
R6684 DVDD.n3102 DVDD.n3076 4.5005
R6685 DVDD.n3102 DVDD.n3086 4.5005
R6686 DVDD.n3102 DVDD.n3075 4.5005
R6687 DVDD.n16083 DVDD.n3102 4.5005
R6688 DVDD.n3102 DVDD.n3057 4.5005
R6689 DVDD.n3102 DVDD.n3053 4.5005
R6690 DVDD.n3088 DVDD.n3080 4.5005
R6691 DVDD.n3088 DVDD.n3082 4.5005
R6692 DVDD.n3088 DVDD.n3079 4.5005
R6693 DVDD.n3088 DVDD.n3083 4.5005
R6694 DVDD.n3088 DVDD.n3078 4.5005
R6695 DVDD.n3088 DVDD.n3084 4.5005
R6696 DVDD.n3088 DVDD.n3077 4.5005
R6697 DVDD.n3088 DVDD.n3085 4.5005
R6698 DVDD.n3088 DVDD.n3076 4.5005
R6699 DVDD.n3088 DVDD.n3086 4.5005
R6700 DVDD.n3088 DVDD.n3075 4.5005
R6701 DVDD.n16083 DVDD.n3088 4.5005
R6702 DVDD.n3088 DVDD.n3057 4.5005
R6703 DVDD.n3088 DVDD.n3053 4.5005
R6704 DVDD.n16082 DVDD.n3080 4.5005
R6705 DVDD.n16082 DVDD.n3082 4.5005
R6706 DVDD.n16082 DVDD.n3079 4.5005
R6707 DVDD.n16082 DVDD.n3083 4.5005
R6708 DVDD.n16082 DVDD.n3078 4.5005
R6709 DVDD.n16082 DVDD.n3084 4.5005
R6710 DVDD.n16082 DVDD.n3077 4.5005
R6711 DVDD.n16082 DVDD.n3085 4.5005
R6712 DVDD.n16082 DVDD.n3076 4.5005
R6713 DVDD.n16082 DVDD.n3086 4.5005
R6714 DVDD.n16082 DVDD.n3075 4.5005
R6715 DVDD.n16083 DVDD.n16082 4.5005
R6716 DVDD.n16082 DVDD.n16081 4.5005
R6717 DVDD.n16082 DVDD.n3057 4.5005
R6718 DVDD.n16082 DVDD.n3053 4.5005
R6719 DVDD.n3080 DVDD.n3059 4.5005
R6720 DVDD.n3082 DVDD.n3059 4.5005
R6721 DVDD.n3079 DVDD.n3059 4.5005
R6722 DVDD.n3083 DVDD.n3059 4.5005
R6723 DVDD.n3078 DVDD.n3059 4.5005
R6724 DVDD.n3084 DVDD.n3059 4.5005
R6725 DVDD.n3077 DVDD.n3059 4.5005
R6726 DVDD.n3085 DVDD.n3059 4.5005
R6727 DVDD.n3076 DVDD.n3059 4.5005
R6728 DVDD.n3086 DVDD.n3059 4.5005
R6729 DVDD.n3075 DVDD.n3059 4.5005
R6730 DVDD.n16083 DVDD.n3059 4.5005
R6731 DVDD.n16081 DVDD.n3059 4.5005
R6732 DVDD.n3059 DVDD.n3057 4.5005
R6733 DVDD.n16085 DVDD.n3059 4.5005
R6734 DVDD.n3059 DVDD.n3053 4.5005
R6735 DVDD.n3193 DVDD.n3161 4.5005
R6736 DVDD.n3194 DVDD.n3161 4.5005
R6737 DVDD.n3192 DVDD.n3161 4.5005
R6738 DVDD.n15989 DVDD.n3161 4.5005
R6739 DVDD.n3190 DVDD.n3161 4.5005
R6740 DVDD.n3197 DVDD.n3161 4.5005
R6741 DVDD.n3189 DVDD.n3161 4.5005
R6742 DVDD.n3198 DVDD.n3161 4.5005
R6743 DVDD.n3188 DVDD.n3161 4.5005
R6744 DVDD.n3200 DVDD.n3161 4.5005
R6745 DVDD.n3186 DVDD.n3161 4.5005
R6746 DVDD.n15987 DVDD.n3161 4.5005
R6747 DVDD.n3193 DVDD.n3163 4.5005
R6748 DVDD.n3194 DVDD.n3163 4.5005
R6749 DVDD.n3192 DVDD.n3163 4.5005
R6750 DVDD.n3196 DVDD.n3163 4.5005
R6751 DVDD.n3191 DVDD.n3163 4.5005
R6752 DVDD.n15989 DVDD.n3163 4.5005
R6753 DVDD.n3190 DVDD.n3163 4.5005
R6754 DVDD.n3197 DVDD.n3163 4.5005
R6755 DVDD.n3189 DVDD.n3163 4.5005
R6756 DVDD.n3198 DVDD.n3163 4.5005
R6757 DVDD.n3188 DVDD.n3163 4.5005
R6758 DVDD.n3199 DVDD.n3163 4.5005
R6759 DVDD.n15937 DVDD.n3163 4.5005
R6760 DVDD.n3200 DVDD.n3163 4.5005
R6761 DVDD.n15987 DVDD.n3163 4.5005
R6762 DVDD.n3193 DVDD.n3160 4.5005
R6763 DVDD.n3194 DVDD.n3160 4.5005
R6764 DVDD.n3192 DVDD.n3160 4.5005
R6765 DVDD.n3196 DVDD.n3160 4.5005
R6766 DVDD.n3191 DVDD.n3160 4.5005
R6767 DVDD.n15989 DVDD.n3160 4.5005
R6768 DVDD.n3190 DVDD.n3160 4.5005
R6769 DVDD.n3197 DVDD.n3160 4.5005
R6770 DVDD.n3189 DVDD.n3160 4.5005
R6771 DVDD.n3198 DVDD.n3160 4.5005
R6772 DVDD.n3188 DVDD.n3160 4.5005
R6773 DVDD.n3199 DVDD.n3160 4.5005
R6774 DVDD.n3200 DVDD.n3160 4.5005
R6775 DVDD.n15987 DVDD.n3160 4.5005
R6776 DVDD.n3193 DVDD.n3164 4.5005
R6777 DVDD.n3194 DVDD.n3164 4.5005
R6778 DVDD.n3192 DVDD.n3164 4.5005
R6779 DVDD.n3196 DVDD.n3164 4.5005
R6780 DVDD.n3191 DVDD.n3164 4.5005
R6781 DVDD.n15989 DVDD.n3164 4.5005
R6782 DVDD.n3190 DVDD.n3164 4.5005
R6783 DVDD.n3197 DVDD.n3164 4.5005
R6784 DVDD.n3189 DVDD.n3164 4.5005
R6785 DVDD.n3198 DVDD.n3164 4.5005
R6786 DVDD.n3188 DVDD.n3164 4.5005
R6787 DVDD.n3199 DVDD.n3164 4.5005
R6788 DVDD.n3200 DVDD.n3164 4.5005
R6789 DVDD.n15987 DVDD.n3164 4.5005
R6790 DVDD.n3193 DVDD.n3159 4.5005
R6791 DVDD.n3194 DVDD.n3159 4.5005
R6792 DVDD.n3192 DVDD.n3159 4.5005
R6793 DVDD.n3196 DVDD.n3159 4.5005
R6794 DVDD.n3191 DVDD.n3159 4.5005
R6795 DVDD.n15989 DVDD.n3159 4.5005
R6796 DVDD.n3190 DVDD.n3159 4.5005
R6797 DVDD.n3197 DVDD.n3159 4.5005
R6798 DVDD.n3189 DVDD.n3159 4.5005
R6799 DVDD.n3198 DVDD.n3159 4.5005
R6800 DVDD.n3188 DVDD.n3159 4.5005
R6801 DVDD.n3199 DVDD.n3159 4.5005
R6802 DVDD.n15937 DVDD.n3159 4.5005
R6803 DVDD.n3200 DVDD.n3159 4.5005
R6804 DVDD.n15987 DVDD.n3159 4.5005
R6805 DVDD.n3193 DVDD.n3165 4.5005
R6806 DVDD.n3194 DVDD.n3165 4.5005
R6807 DVDD.n3192 DVDD.n3165 4.5005
R6808 DVDD.n3196 DVDD.n3165 4.5005
R6809 DVDD.n3191 DVDD.n3165 4.5005
R6810 DVDD.n15989 DVDD.n3165 4.5005
R6811 DVDD.n3190 DVDD.n3165 4.5005
R6812 DVDD.n3197 DVDD.n3165 4.5005
R6813 DVDD.n3189 DVDD.n3165 4.5005
R6814 DVDD.n3198 DVDD.n3165 4.5005
R6815 DVDD.n3188 DVDD.n3165 4.5005
R6816 DVDD.n3199 DVDD.n3165 4.5005
R6817 DVDD.n15937 DVDD.n3165 4.5005
R6818 DVDD.n3200 DVDD.n3165 4.5005
R6819 DVDD.n15987 DVDD.n3165 4.5005
R6820 DVDD.n3193 DVDD.n3158 4.5005
R6821 DVDD.n3194 DVDD.n3158 4.5005
R6822 DVDD.n3192 DVDD.n3158 4.5005
R6823 DVDD.n3196 DVDD.n3158 4.5005
R6824 DVDD.n3191 DVDD.n3158 4.5005
R6825 DVDD.n15989 DVDD.n3158 4.5005
R6826 DVDD.n3190 DVDD.n3158 4.5005
R6827 DVDD.n3197 DVDD.n3158 4.5005
R6828 DVDD.n3189 DVDD.n3158 4.5005
R6829 DVDD.n3198 DVDD.n3158 4.5005
R6830 DVDD.n3188 DVDD.n3158 4.5005
R6831 DVDD.n3199 DVDD.n3158 4.5005
R6832 DVDD.n3200 DVDD.n3158 4.5005
R6833 DVDD.n15987 DVDD.n3158 4.5005
R6834 DVDD.n3193 DVDD.n3166 4.5005
R6835 DVDD.n3194 DVDD.n3166 4.5005
R6836 DVDD.n3192 DVDD.n3166 4.5005
R6837 DVDD.n3196 DVDD.n3166 4.5005
R6838 DVDD.n3191 DVDD.n3166 4.5005
R6839 DVDD.n15989 DVDD.n3166 4.5005
R6840 DVDD.n3190 DVDD.n3166 4.5005
R6841 DVDD.n3197 DVDD.n3166 4.5005
R6842 DVDD.n3189 DVDD.n3166 4.5005
R6843 DVDD.n3198 DVDD.n3166 4.5005
R6844 DVDD.n3188 DVDD.n3166 4.5005
R6845 DVDD.n3199 DVDD.n3166 4.5005
R6846 DVDD.n3200 DVDD.n3166 4.5005
R6847 DVDD.n15987 DVDD.n3166 4.5005
R6848 DVDD.n3193 DVDD.n3157 4.5005
R6849 DVDD.n3194 DVDD.n3157 4.5005
R6850 DVDD.n3192 DVDD.n3157 4.5005
R6851 DVDD.n3196 DVDD.n3157 4.5005
R6852 DVDD.n3191 DVDD.n3157 4.5005
R6853 DVDD.n15989 DVDD.n3157 4.5005
R6854 DVDD.n3190 DVDD.n3157 4.5005
R6855 DVDD.n3197 DVDD.n3157 4.5005
R6856 DVDD.n3189 DVDD.n3157 4.5005
R6857 DVDD.n3198 DVDD.n3157 4.5005
R6858 DVDD.n3188 DVDD.n3157 4.5005
R6859 DVDD.n3199 DVDD.n3157 4.5005
R6860 DVDD.n15937 DVDD.n3157 4.5005
R6861 DVDD.n3200 DVDD.n3157 4.5005
R6862 DVDD.n15987 DVDD.n3157 4.5005
R6863 DVDD.n3193 DVDD.n3167 4.5005
R6864 DVDD.n3194 DVDD.n3167 4.5005
R6865 DVDD.n3192 DVDD.n3167 4.5005
R6866 DVDD.n3196 DVDD.n3167 4.5005
R6867 DVDD.n3191 DVDD.n3167 4.5005
R6868 DVDD.n15989 DVDD.n3167 4.5005
R6869 DVDD.n3190 DVDD.n3167 4.5005
R6870 DVDD.n3197 DVDD.n3167 4.5005
R6871 DVDD.n3189 DVDD.n3167 4.5005
R6872 DVDD.n3198 DVDD.n3167 4.5005
R6873 DVDD.n3188 DVDD.n3167 4.5005
R6874 DVDD.n3199 DVDD.n3167 4.5005
R6875 DVDD.n15937 DVDD.n3167 4.5005
R6876 DVDD.n3200 DVDD.n3167 4.5005
R6877 DVDD.n15987 DVDD.n3167 4.5005
R6878 DVDD.n3193 DVDD.n3156 4.5005
R6879 DVDD.n3194 DVDD.n3156 4.5005
R6880 DVDD.n3192 DVDD.n3156 4.5005
R6881 DVDD.n3196 DVDD.n3156 4.5005
R6882 DVDD.n3191 DVDD.n3156 4.5005
R6883 DVDD.n15989 DVDD.n3156 4.5005
R6884 DVDD.n3190 DVDD.n3156 4.5005
R6885 DVDD.n3197 DVDD.n3156 4.5005
R6886 DVDD.n3189 DVDD.n3156 4.5005
R6887 DVDD.n3198 DVDD.n3156 4.5005
R6888 DVDD.n3188 DVDD.n3156 4.5005
R6889 DVDD.n3199 DVDD.n3156 4.5005
R6890 DVDD.n3200 DVDD.n3156 4.5005
R6891 DVDD.n15987 DVDD.n3156 4.5005
R6892 DVDD.n3193 DVDD.n3168 4.5005
R6893 DVDD.n3194 DVDD.n3168 4.5005
R6894 DVDD.n3192 DVDD.n3168 4.5005
R6895 DVDD.n3196 DVDD.n3168 4.5005
R6896 DVDD.n3191 DVDD.n3168 4.5005
R6897 DVDD.n15989 DVDD.n3168 4.5005
R6898 DVDD.n3190 DVDD.n3168 4.5005
R6899 DVDD.n3197 DVDD.n3168 4.5005
R6900 DVDD.n3189 DVDD.n3168 4.5005
R6901 DVDD.n3198 DVDD.n3168 4.5005
R6902 DVDD.n3188 DVDD.n3168 4.5005
R6903 DVDD.n3199 DVDD.n3168 4.5005
R6904 DVDD.n3200 DVDD.n3168 4.5005
R6905 DVDD.n15987 DVDD.n3168 4.5005
R6906 DVDD.n3193 DVDD.n3155 4.5005
R6907 DVDD.n3194 DVDD.n3155 4.5005
R6908 DVDD.n3192 DVDD.n3155 4.5005
R6909 DVDD.n3196 DVDD.n3155 4.5005
R6910 DVDD.n3191 DVDD.n3155 4.5005
R6911 DVDD.n15989 DVDD.n3155 4.5005
R6912 DVDD.n3190 DVDD.n3155 4.5005
R6913 DVDD.n3197 DVDD.n3155 4.5005
R6914 DVDD.n3189 DVDD.n3155 4.5005
R6915 DVDD.n3198 DVDD.n3155 4.5005
R6916 DVDD.n3188 DVDD.n3155 4.5005
R6917 DVDD.n3199 DVDD.n3155 4.5005
R6918 DVDD.n15937 DVDD.n3155 4.5005
R6919 DVDD.n3200 DVDD.n3155 4.5005
R6920 DVDD.n15987 DVDD.n3155 4.5005
R6921 DVDD.n3193 DVDD.n3169 4.5005
R6922 DVDD.n3194 DVDD.n3169 4.5005
R6923 DVDD.n3192 DVDD.n3169 4.5005
R6924 DVDD.n3196 DVDD.n3169 4.5005
R6925 DVDD.n3191 DVDD.n3169 4.5005
R6926 DVDD.n15989 DVDD.n3169 4.5005
R6927 DVDD.n3190 DVDD.n3169 4.5005
R6928 DVDD.n3197 DVDD.n3169 4.5005
R6929 DVDD.n3189 DVDD.n3169 4.5005
R6930 DVDD.n3198 DVDD.n3169 4.5005
R6931 DVDD.n3188 DVDD.n3169 4.5005
R6932 DVDD.n3199 DVDD.n3169 4.5005
R6933 DVDD.n15937 DVDD.n3169 4.5005
R6934 DVDD.n3200 DVDD.n3169 4.5005
R6935 DVDD.n15987 DVDD.n3169 4.5005
R6936 DVDD.n3193 DVDD.n3154 4.5005
R6937 DVDD.n3194 DVDD.n3154 4.5005
R6938 DVDD.n3192 DVDD.n3154 4.5005
R6939 DVDD.n3196 DVDD.n3154 4.5005
R6940 DVDD.n3191 DVDD.n3154 4.5005
R6941 DVDD.n15989 DVDD.n3154 4.5005
R6942 DVDD.n3190 DVDD.n3154 4.5005
R6943 DVDD.n3197 DVDD.n3154 4.5005
R6944 DVDD.n3189 DVDD.n3154 4.5005
R6945 DVDD.n3198 DVDD.n3154 4.5005
R6946 DVDD.n3188 DVDD.n3154 4.5005
R6947 DVDD.n3199 DVDD.n3154 4.5005
R6948 DVDD.n3200 DVDD.n3154 4.5005
R6949 DVDD.n15987 DVDD.n3154 4.5005
R6950 DVDD.n3193 DVDD.n3170 4.5005
R6951 DVDD.n3194 DVDD.n3170 4.5005
R6952 DVDD.n3192 DVDD.n3170 4.5005
R6953 DVDD.n3196 DVDD.n3170 4.5005
R6954 DVDD.n3191 DVDD.n3170 4.5005
R6955 DVDD.n15989 DVDD.n3170 4.5005
R6956 DVDD.n3190 DVDD.n3170 4.5005
R6957 DVDD.n3197 DVDD.n3170 4.5005
R6958 DVDD.n3189 DVDD.n3170 4.5005
R6959 DVDD.n3198 DVDD.n3170 4.5005
R6960 DVDD.n3188 DVDD.n3170 4.5005
R6961 DVDD.n3199 DVDD.n3170 4.5005
R6962 DVDD.n3200 DVDD.n3170 4.5005
R6963 DVDD.n15987 DVDD.n3170 4.5005
R6964 DVDD.n3193 DVDD.n3153 4.5005
R6965 DVDD.n3194 DVDD.n3153 4.5005
R6966 DVDD.n3192 DVDD.n3153 4.5005
R6967 DVDD.n3196 DVDD.n3153 4.5005
R6968 DVDD.n3191 DVDD.n3153 4.5005
R6969 DVDD.n15989 DVDD.n3153 4.5005
R6970 DVDD.n3190 DVDD.n3153 4.5005
R6971 DVDD.n3197 DVDD.n3153 4.5005
R6972 DVDD.n3189 DVDD.n3153 4.5005
R6973 DVDD.n3198 DVDD.n3153 4.5005
R6974 DVDD.n3188 DVDD.n3153 4.5005
R6975 DVDD.n3199 DVDD.n3153 4.5005
R6976 DVDD.n3200 DVDD.n3153 4.5005
R6977 DVDD.n15987 DVDD.n3153 4.5005
R6978 DVDD.n3193 DVDD.n3171 4.5005
R6979 DVDD.n3194 DVDD.n3171 4.5005
R6980 DVDD.n3192 DVDD.n3171 4.5005
R6981 DVDD.n3196 DVDD.n3171 4.5005
R6982 DVDD.n3191 DVDD.n3171 4.5005
R6983 DVDD.n15989 DVDD.n3171 4.5005
R6984 DVDD.n3190 DVDD.n3171 4.5005
R6985 DVDD.n3197 DVDD.n3171 4.5005
R6986 DVDD.n3189 DVDD.n3171 4.5005
R6987 DVDD.n3198 DVDD.n3171 4.5005
R6988 DVDD.n3188 DVDD.n3171 4.5005
R6989 DVDD.n3199 DVDD.n3171 4.5005
R6990 DVDD.n3200 DVDD.n3171 4.5005
R6991 DVDD.n15987 DVDD.n3171 4.5005
R6992 DVDD.n3193 DVDD.n3152 4.5005
R6993 DVDD.n3194 DVDD.n3152 4.5005
R6994 DVDD.n3192 DVDD.n3152 4.5005
R6995 DVDD.n3196 DVDD.n3152 4.5005
R6996 DVDD.n3191 DVDD.n3152 4.5005
R6997 DVDD.n15989 DVDD.n3152 4.5005
R6998 DVDD.n3190 DVDD.n3152 4.5005
R6999 DVDD.n3197 DVDD.n3152 4.5005
R7000 DVDD.n3189 DVDD.n3152 4.5005
R7001 DVDD.n3198 DVDD.n3152 4.5005
R7002 DVDD.n3188 DVDD.n3152 4.5005
R7003 DVDD.n3199 DVDD.n3152 4.5005
R7004 DVDD.n3200 DVDD.n3152 4.5005
R7005 DVDD.n15987 DVDD.n3152 4.5005
R7006 DVDD.n3193 DVDD.n3172 4.5005
R7007 DVDD.n3194 DVDD.n3172 4.5005
R7008 DVDD.n3192 DVDD.n3172 4.5005
R7009 DVDD.n3196 DVDD.n3172 4.5005
R7010 DVDD.n3191 DVDD.n3172 4.5005
R7011 DVDD.n15989 DVDD.n3172 4.5005
R7012 DVDD.n3190 DVDD.n3172 4.5005
R7013 DVDD.n3197 DVDD.n3172 4.5005
R7014 DVDD.n3189 DVDD.n3172 4.5005
R7015 DVDD.n3198 DVDD.n3172 4.5005
R7016 DVDD.n3188 DVDD.n3172 4.5005
R7017 DVDD.n3199 DVDD.n3172 4.5005
R7018 DVDD.n3200 DVDD.n3172 4.5005
R7019 DVDD.n15987 DVDD.n3172 4.5005
R7020 DVDD.n3193 DVDD.n3151 4.5005
R7021 DVDD.n3194 DVDD.n3151 4.5005
R7022 DVDD.n3192 DVDD.n3151 4.5005
R7023 DVDD.n3196 DVDD.n3151 4.5005
R7024 DVDD.n3191 DVDD.n3151 4.5005
R7025 DVDD.n15989 DVDD.n3151 4.5005
R7026 DVDD.n3190 DVDD.n3151 4.5005
R7027 DVDD.n3197 DVDD.n3151 4.5005
R7028 DVDD.n3189 DVDD.n3151 4.5005
R7029 DVDD.n3198 DVDD.n3151 4.5005
R7030 DVDD.n3188 DVDD.n3151 4.5005
R7031 DVDD.n3199 DVDD.n3151 4.5005
R7032 DVDD.n15937 DVDD.n3151 4.5005
R7033 DVDD.n3200 DVDD.n3151 4.5005
R7034 DVDD.n15987 DVDD.n3151 4.5005
R7035 DVDD.n3193 DVDD.n3173 4.5005
R7036 DVDD.n3194 DVDD.n3173 4.5005
R7037 DVDD.n3192 DVDD.n3173 4.5005
R7038 DVDD.n3196 DVDD.n3173 4.5005
R7039 DVDD.n3191 DVDD.n3173 4.5005
R7040 DVDD.n15989 DVDD.n3173 4.5005
R7041 DVDD.n3190 DVDD.n3173 4.5005
R7042 DVDD.n3197 DVDD.n3173 4.5005
R7043 DVDD.n3189 DVDD.n3173 4.5005
R7044 DVDD.n3198 DVDD.n3173 4.5005
R7045 DVDD.n3188 DVDD.n3173 4.5005
R7046 DVDD.n3199 DVDD.n3173 4.5005
R7047 DVDD.n15937 DVDD.n3173 4.5005
R7048 DVDD.n3200 DVDD.n3173 4.5005
R7049 DVDD.n15987 DVDD.n3173 4.5005
R7050 DVDD.n3193 DVDD.n3150 4.5005
R7051 DVDD.n3194 DVDD.n3150 4.5005
R7052 DVDD.n3192 DVDD.n3150 4.5005
R7053 DVDD.n3196 DVDD.n3150 4.5005
R7054 DVDD.n3191 DVDD.n3150 4.5005
R7055 DVDD.n15989 DVDD.n3150 4.5005
R7056 DVDD.n3190 DVDD.n3150 4.5005
R7057 DVDD.n3197 DVDD.n3150 4.5005
R7058 DVDD.n3189 DVDD.n3150 4.5005
R7059 DVDD.n3198 DVDD.n3150 4.5005
R7060 DVDD.n3188 DVDD.n3150 4.5005
R7061 DVDD.n3199 DVDD.n3150 4.5005
R7062 DVDD.n3200 DVDD.n3150 4.5005
R7063 DVDD.n15987 DVDD.n3150 4.5005
R7064 DVDD.n15988 DVDD.n3193 4.5005
R7065 DVDD.n15988 DVDD.n3194 4.5005
R7066 DVDD.n15988 DVDD.n3192 4.5005
R7067 DVDD.n15988 DVDD.n3196 4.5005
R7068 DVDD.n15988 DVDD.n3191 4.5005
R7069 DVDD.n15989 DVDD.n15988 4.5005
R7070 DVDD.n15988 DVDD.n3190 4.5005
R7071 DVDD.n15988 DVDD.n3197 4.5005
R7072 DVDD.n15988 DVDD.n3189 4.5005
R7073 DVDD.n15988 DVDD.n3198 4.5005
R7074 DVDD.n15988 DVDD.n3188 4.5005
R7075 DVDD.n15988 DVDD.n3199 4.5005
R7076 DVDD.n15988 DVDD.n3200 4.5005
R7077 DVDD.n15988 DVDD.n3186 4.5005
R7078 DVDD.n15988 DVDD.n15987 4.5005
R7079 DVDD.n3285 DVDD.n3247 4.5005
R7080 DVDD.n3287 DVDD.n3247 4.5005
R7081 DVDD.n3284 DVDD.n3247 4.5005
R7082 DVDD.n3247 DVDD.n3235 4.5005
R7083 DVDD.n15909 DVDD.n3247 4.5005
R7084 DVDD.n3290 DVDD.n3247 4.5005
R7085 DVDD.n3281 DVDD.n3247 4.5005
R7086 DVDD.n3291 DVDD.n3247 4.5005
R7087 DVDD.n3280 DVDD.n3247 4.5005
R7088 DVDD.n3294 DVDD.n3247 4.5005
R7089 DVDD.n15907 DVDD.n3247 4.5005
R7090 DVDD.n3285 DVDD.n3249 4.5005
R7091 DVDD.n3287 DVDD.n3249 4.5005
R7092 DVDD.n3284 DVDD.n3249 4.5005
R7093 DVDD.n3289 DVDD.n3249 4.5005
R7094 DVDD.n3283 DVDD.n3249 4.5005
R7095 DVDD.n3249 DVDD.n3235 4.5005
R7096 DVDD.n15909 DVDD.n3249 4.5005
R7097 DVDD.n3290 DVDD.n3249 4.5005
R7098 DVDD.n3281 DVDD.n3249 4.5005
R7099 DVDD.n3291 DVDD.n3249 4.5005
R7100 DVDD.n3280 DVDD.n3249 4.5005
R7101 DVDD.n3293 DVDD.n3249 4.5005
R7102 DVDD.n3294 DVDD.n3249 4.5005
R7103 DVDD.n15907 DVDD.n3249 4.5005
R7104 DVDD.n3285 DVDD.n3246 4.5005
R7105 DVDD.n3287 DVDD.n3246 4.5005
R7106 DVDD.n3284 DVDD.n3246 4.5005
R7107 DVDD.n3289 DVDD.n3246 4.5005
R7108 DVDD.n3283 DVDD.n3246 4.5005
R7109 DVDD.n3246 DVDD.n3235 4.5005
R7110 DVDD.n15909 DVDD.n3246 4.5005
R7111 DVDD.n3290 DVDD.n3246 4.5005
R7112 DVDD.n3281 DVDD.n3246 4.5005
R7113 DVDD.n3291 DVDD.n3246 4.5005
R7114 DVDD.n3280 DVDD.n3246 4.5005
R7115 DVDD.n3293 DVDD.n3246 4.5005
R7116 DVDD.n3294 DVDD.n3246 4.5005
R7117 DVDD.n3272 DVDD.n3246 4.5005
R7118 DVDD.n15907 DVDD.n3246 4.5005
R7119 DVDD.n3285 DVDD.n3250 4.5005
R7120 DVDD.n3287 DVDD.n3250 4.5005
R7121 DVDD.n3284 DVDD.n3250 4.5005
R7122 DVDD.n3289 DVDD.n3250 4.5005
R7123 DVDD.n3283 DVDD.n3250 4.5005
R7124 DVDD.n3250 DVDD.n3235 4.5005
R7125 DVDD.n15909 DVDD.n3250 4.5005
R7126 DVDD.n3290 DVDD.n3250 4.5005
R7127 DVDD.n3281 DVDD.n3250 4.5005
R7128 DVDD.n3291 DVDD.n3250 4.5005
R7129 DVDD.n3280 DVDD.n3250 4.5005
R7130 DVDD.n3293 DVDD.n3250 4.5005
R7131 DVDD.n3279 DVDD.n3250 4.5005
R7132 DVDD.n3294 DVDD.n3250 4.5005
R7133 DVDD.n15907 DVDD.n3250 4.5005
R7134 DVDD.n3285 DVDD.n3245 4.5005
R7135 DVDD.n3287 DVDD.n3245 4.5005
R7136 DVDD.n3284 DVDD.n3245 4.5005
R7137 DVDD.n3289 DVDD.n3245 4.5005
R7138 DVDD.n3283 DVDD.n3245 4.5005
R7139 DVDD.n3245 DVDD.n3235 4.5005
R7140 DVDD.n15909 DVDD.n3245 4.5005
R7141 DVDD.n3290 DVDD.n3245 4.5005
R7142 DVDD.n3281 DVDD.n3245 4.5005
R7143 DVDD.n3291 DVDD.n3245 4.5005
R7144 DVDD.n3280 DVDD.n3245 4.5005
R7145 DVDD.n3293 DVDD.n3245 4.5005
R7146 DVDD.n3294 DVDD.n3245 4.5005
R7147 DVDD.n15907 DVDD.n3245 4.5005
R7148 DVDD.n3285 DVDD.n3251 4.5005
R7149 DVDD.n3287 DVDD.n3251 4.5005
R7150 DVDD.n3284 DVDD.n3251 4.5005
R7151 DVDD.n3289 DVDD.n3251 4.5005
R7152 DVDD.n3283 DVDD.n3251 4.5005
R7153 DVDD.n3251 DVDD.n3235 4.5005
R7154 DVDD.n15909 DVDD.n3251 4.5005
R7155 DVDD.n3290 DVDD.n3251 4.5005
R7156 DVDD.n3281 DVDD.n3251 4.5005
R7157 DVDD.n3291 DVDD.n3251 4.5005
R7158 DVDD.n3280 DVDD.n3251 4.5005
R7159 DVDD.n3293 DVDD.n3251 4.5005
R7160 DVDD.n3294 DVDD.n3251 4.5005
R7161 DVDD.n15907 DVDD.n3251 4.5005
R7162 DVDD.n3285 DVDD.n3244 4.5005
R7163 DVDD.n3287 DVDD.n3244 4.5005
R7164 DVDD.n3284 DVDD.n3244 4.5005
R7165 DVDD.n3289 DVDD.n3244 4.5005
R7166 DVDD.n3283 DVDD.n3244 4.5005
R7167 DVDD.n3244 DVDD.n3235 4.5005
R7168 DVDD.n15909 DVDD.n3244 4.5005
R7169 DVDD.n3290 DVDD.n3244 4.5005
R7170 DVDD.n3281 DVDD.n3244 4.5005
R7171 DVDD.n3291 DVDD.n3244 4.5005
R7172 DVDD.n3280 DVDD.n3244 4.5005
R7173 DVDD.n3293 DVDD.n3244 4.5005
R7174 DVDD.n3279 DVDD.n3244 4.5005
R7175 DVDD.n3294 DVDD.n3244 4.5005
R7176 DVDD.n15907 DVDD.n3244 4.5005
R7177 DVDD.n3285 DVDD.n3252 4.5005
R7178 DVDD.n3287 DVDD.n3252 4.5005
R7179 DVDD.n3284 DVDD.n3252 4.5005
R7180 DVDD.n3289 DVDD.n3252 4.5005
R7181 DVDD.n3283 DVDD.n3252 4.5005
R7182 DVDD.n3252 DVDD.n3235 4.5005
R7183 DVDD.n15909 DVDD.n3252 4.5005
R7184 DVDD.n3290 DVDD.n3252 4.5005
R7185 DVDD.n3281 DVDD.n3252 4.5005
R7186 DVDD.n3291 DVDD.n3252 4.5005
R7187 DVDD.n3280 DVDD.n3252 4.5005
R7188 DVDD.n3293 DVDD.n3252 4.5005
R7189 DVDD.n3279 DVDD.n3252 4.5005
R7190 DVDD.n3294 DVDD.n3252 4.5005
R7191 DVDD.n15907 DVDD.n3252 4.5005
R7192 DVDD.n3285 DVDD.n3243 4.5005
R7193 DVDD.n3287 DVDD.n3243 4.5005
R7194 DVDD.n3284 DVDD.n3243 4.5005
R7195 DVDD.n3289 DVDD.n3243 4.5005
R7196 DVDD.n3283 DVDD.n3243 4.5005
R7197 DVDD.n3243 DVDD.n3235 4.5005
R7198 DVDD.n15909 DVDD.n3243 4.5005
R7199 DVDD.n3290 DVDD.n3243 4.5005
R7200 DVDD.n3281 DVDD.n3243 4.5005
R7201 DVDD.n3291 DVDD.n3243 4.5005
R7202 DVDD.n3280 DVDD.n3243 4.5005
R7203 DVDD.n3293 DVDD.n3243 4.5005
R7204 DVDD.n3294 DVDD.n3243 4.5005
R7205 DVDD.n15907 DVDD.n3243 4.5005
R7206 DVDD.n3285 DVDD.n3253 4.5005
R7207 DVDD.n3287 DVDD.n3253 4.5005
R7208 DVDD.n3284 DVDD.n3253 4.5005
R7209 DVDD.n3289 DVDD.n3253 4.5005
R7210 DVDD.n3283 DVDD.n3253 4.5005
R7211 DVDD.n3253 DVDD.n3235 4.5005
R7212 DVDD.n15909 DVDD.n3253 4.5005
R7213 DVDD.n3290 DVDD.n3253 4.5005
R7214 DVDD.n3281 DVDD.n3253 4.5005
R7215 DVDD.n3291 DVDD.n3253 4.5005
R7216 DVDD.n3280 DVDD.n3253 4.5005
R7217 DVDD.n3293 DVDD.n3253 4.5005
R7218 DVDD.n3294 DVDD.n3253 4.5005
R7219 DVDD.n15907 DVDD.n3253 4.5005
R7220 DVDD.n3285 DVDD.n3242 4.5005
R7221 DVDD.n3287 DVDD.n3242 4.5005
R7222 DVDD.n3284 DVDD.n3242 4.5005
R7223 DVDD.n3289 DVDD.n3242 4.5005
R7224 DVDD.n3283 DVDD.n3242 4.5005
R7225 DVDD.n3242 DVDD.n3235 4.5005
R7226 DVDD.n15909 DVDD.n3242 4.5005
R7227 DVDD.n3290 DVDD.n3242 4.5005
R7228 DVDD.n3281 DVDD.n3242 4.5005
R7229 DVDD.n3291 DVDD.n3242 4.5005
R7230 DVDD.n3280 DVDD.n3242 4.5005
R7231 DVDD.n3293 DVDD.n3242 4.5005
R7232 DVDD.n3279 DVDD.n3242 4.5005
R7233 DVDD.n3294 DVDD.n3242 4.5005
R7234 DVDD.n15907 DVDD.n3242 4.5005
R7235 DVDD.n3285 DVDD.n3254 4.5005
R7236 DVDD.n3287 DVDD.n3254 4.5005
R7237 DVDD.n3284 DVDD.n3254 4.5005
R7238 DVDD.n3289 DVDD.n3254 4.5005
R7239 DVDD.n3283 DVDD.n3254 4.5005
R7240 DVDD.n3254 DVDD.n3235 4.5005
R7241 DVDD.n15909 DVDD.n3254 4.5005
R7242 DVDD.n3290 DVDD.n3254 4.5005
R7243 DVDD.n3281 DVDD.n3254 4.5005
R7244 DVDD.n3291 DVDD.n3254 4.5005
R7245 DVDD.n3280 DVDD.n3254 4.5005
R7246 DVDD.n3293 DVDD.n3254 4.5005
R7247 DVDD.n3279 DVDD.n3254 4.5005
R7248 DVDD.n3294 DVDD.n3254 4.5005
R7249 DVDD.n15907 DVDD.n3254 4.5005
R7250 DVDD.n3285 DVDD.n3241 4.5005
R7251 DVDD.n3287 DVDD.n3241 4.5005
R7252 DVDD.n3284 DVDD.n3241 4.5005
R7253 DVDD.n3289 DVDD.n3241 4.5005
R7254 DVDD.n3283 DVDD.n3241 4.5005
R7255 DVDD.n3241 DVDD.n3235 4.5005
R7256 DVDD.n15909 DVDD.n3241 4.5005
R7257 DVDD.n3290 DVDD.n3241 4.5005
R7258 DVDD.n3281 DVDD.n3241 4.5005
R7259 DVDD.n3291 DVDD.n3241 4.5005
R7260 DVDD.n3280 DVDD.n3241 4.5005
R7261 DVDD.n3293 DVDD.n3241 4.5005
R7262 DVDD.n3294 DVDD.n3241 4.5005
R7263 DVDD.n15907 DVDD.n3241 4.5005
R7264 DVDD.n3285 DVDD.n3255 4.5005
R7265 DVDD.n3287 DVDD.n3255 4.5005
R7266 DVDD.n3284 DVDD.n3255 4.5005
R7267 DVDD.n3289 DVDD.n3255 4.5005
R7268 DVDD.n3283 DVDD.n3255 4.5005
R7269 DVDD.n3255 DVDD.n3235 4.5005
R7270 DVDD.n15909 DVDD.n3255 4.5005
R7271 DVDD.n3290 DVDD.n3255 4.5005
R7272 DVDD.n3281 DVDD.n3255 4.5005
R7273 DVDD.n3291 DVDD.n3255 4.5005
R7274 DVDD.n3280 DVDD.n3255 4.5005
R7275 DVDD.n3293 DVDD.n3255 4.5005
R7276 DVDD.n3294 DVDD.n3255 4.5005
R7277 DVDD.n15907 DVDD.n3255 4.5005
R7278 DVDD.n3285 DVDD.n3240 4.5005
R7279 DVDD.n3287 DVDD.n3240 4.5005
R7280 DVDD.n3284 DVDD.n3240 4.5005
R7281 DVDD.n3289 DVDD.n3240 4.5005
R7282 DVDD.n3283 DVDD.n3240 4.5005
R7283 DVDD.n3240 DVDD.n3235 4.5005
R7284 DVDD.n15909 DVDD.n3240 4.5005
R7285 DVDD.n3290 DVDD.n3240 4.5005
R7286 DVDD.n3281 DVDD.n3240 4.5005
R7287 DVDD.n3291 DVDD.n3240 4.5005
R7288 DVDD.n3280 DVDD.n3240 4.5005
R7289 DVDD.n3293 DVDD.n3240 4.5005
R7290 DVDD.n3279 DVDD.n3240 4.5005
R7291 DVDD.n3294 DVDD.n3240 4.5005
R7292 DVDD.n15907 DVDD.n3240 4.5005
R7293 DVDD.n3285 DVDD.n3256 4.5005
R7294 DVDD.n3287 DVDD.n3256 4.5005
R7295 DVDD.n3284 DVDD.n3256 4.5005
R7296 DVDD.n3289 DVDD.n3256 4.5005
R7297 DVDD.n3283 DVDD.n3256 4.5005
R7298 DVDD.n3256 DVDD.n3235 4.5005
R7299 DVDD.n15909 DVDD.n3256 4.5005
R7300 DVDD.n3290 DVDD.n3256 4.5005
R7301 DVDD.n3281 DVDD.n3256 4.5005
R7302 DVDD.n3291 DVDD.n3256 4.5005
R7303 DVDD.n3280 DVDD.n3256 4.5005
R7304 DVDD.n3293 DVDD.n3256 4.5005
R7305 DVDD.n3279 DVDD.n3256 4.5005
R7306 DVDD.n3294 DVDD.n3256 4.5005
R7307 DVDD.n15907 DVDD.n3256 4.5005
R7308 DVDD.n3285 DVDD.n3239 4.5005
R7309 DVDD.n3287 DVDD.n3239 4.5005
R7310 DVDD.n3284 DVDD.n3239 4.5005
R7311 DVDD.n3289 DVDD.n3239 4.5005
R7312 DVDD.n3283 DVDD.n3239 4.5005
R7313 DVDD.n3239 DVDD.n3235 4.5005
R7314 DVDD.n15909 DVDD.n3239 4.5005
R7315 DVDD.n3290 DVDD.n3239 4.5005
R7316 DVDD.n3281 DVDD.n3239 4.5005
R7317 DVDD.n3291 DVDD.n3239 4.5005
R7318 DVDD.n3280 DVDD.n3239 4.5005
R7319 DVDD.n3293 DVDD.n3239 4.5005
R7320 DVDD.n3294 DVDD.n3239 4.5005
R7321 DVDD.n15907 DVDD.n3239 4.5005
R7322 DVDD.n3285 DVDD.n3257 4.5005
R7323 DVDD.n3287 DVDD.n3257 4.5005
R7324 DVDD.n3284 DVDD.n3257 4.5005
R7325 DVDD.n3289 DVDD.n3257 4.5005
R7326 DVDD.n3283 DVDD.n3257 4.5005
R7327 DVDD.n3257 DVDD.n3235 4.5005
R7328 DVDD.n15909 DVDD.n3257 4.5005
R7329 DVDD.n3290 DVDD.n3257 4.5005
R7330 DVDD.n3281 DVDD.n3257 4.5005
R7331 DVDD.n3291 DVDD.n3257 4.5005
R7332 DVDD.n3280 DVDD.n3257 4.5005
R7333 DVDD.n3293 DVDD.n3257 4.5005
R7334 DVDD.n3294 DVDD.n3257 4.5005
R7335 DVDD.n15907 DVDD.n3257 4.5005
R7336 DVDD.n3285 DVDD.n3238 4.5005
R7337 DVDD.n3287 DVDD.n3238 4.5005
R7338 DVDD.n3284 DVDD.n3238 4.5005
R7339 DVDD.n3289 DVDD.n3238 4.5005
R7340 DVDD.n3283 DVDD.n3238 4.5005
R7341 DVDD.n3238 DVDD.n3235 4.5005
R7342 DVDD.n15909 DVDD.n3238 4.5005
R7343 DVDD.n3290 DVDD.n3238 4.5005
R7344 DVDD.n3281 DVDD.n3238 4.5005
R7345 DVDD.n3291 DVDD.n3238 4.5005
R7346 DVDD.n3280 DVDD.n3238 4.5005
R7347 DVDD.n3293 DVDD.n3238 4.5005
R7348 DVDD.n3279 DVDD.n3238 4.5005
R7349 DVDD.n3294 DVDD.n3238 4.5005
R7350 DVDD.n15907 DVDD.n3238 4.5005
R7351 DVDD.n3285 DVDD.n3258 4.5005
R7352 DVDD.n3287 DVDD.n3258 4.5005
R7353 DVDD.n3284 DVDD.n3258 4.5005
R7354 DVDD.n3289 DVDD.n3258 4.5005
R7355 DVDD.n3283 DVDD.n3258 4.5005
R7356 DVDD.n3258 DVDD.n3235 4.5005
R7357 DVDD.n15909 DVDD.n3258 4.5005
R7358 DVDD.n3290 DVDD.n3258 4.5005
R7359 DVDD.n3281 DVDD.n3258 4.5005
R7360 DVDD.n3291 DVDD.n3258 4.5005
R7361 DVDD.n3280 DVDD.n3258 4.5005
R7362 DVDD.n3293 DVDD.n3258 4.5005
R7363 DVDD.n3279 DVDD.n3258 4.5005
R7364 DVDD.n3294 DVDD.n3258 4.5005
R7365 DVDD.n15907 DVDD.n3258 4.5005
R7366 DVDD.n3285 DVDD.n3237 4.5005
R7367 DVDD.n3287 DVDD.n3237 4.5005
R7368 DVDD.n3284 DVDD.n3237 4.5005
R7369 DVDD.n3289 DVDD.n3237 4.5005
R7370 DVDD.n3283 DVDD.n3237 4.5005
R7371 DVDD.n3237 DVDD.n3235 4.5005
R7372 DVDD.n15909 DVDD.n3237 4.5005
R7373 DVDD.n3290 DVDD.n3237 4.5005
R7374 DVDD.n3281 DVDD.n3237 4.5005
R7375 DVDD.n3291 DVDD.n3237 4.5005
R7376 DVDD.n3280 DVDD.n3237 4.5005
R7377 DVDD.n3293 DVDD.n3237 4.5005
R7378 DVDD.n3294 DVDD.n3237 4.5005
R7379 DVDD.n15907 DVDD.n3237 4.5005
R7380 DVDD.n3285 DVDD.n3259 4.5005
R7381 DVDD.n3287 DVDD.n3259 4.5005
R7382 DVDD.n3284 DVDD.n3259 4.5005
R7383 DVDD.n3289 DVDD.n3259 4.5005
R7384 DVDD.n3283 DVDD.n3259 4.5005
R7385 DVDD.n3259 DVDD.n3235 4.5005
R7386 DVDD.n15909 DVDD.n3259 4.5005
R7387 DVDD.n3290 DVDD.n3259 4.5005
R7388 DVDD.n3281 DVDD.n3259 4.5005
R7389 DVDD.n3291 DVDD.n3259 4.5005
R7390 DVDD.n3280 DVDD.n3259 4.5005
R7391 DVDD.n3293 DVDD.n3259 4.5005
R7392 DVDD.n3294 DVDD.n3259 4.5005
R7393 DVDD.n15907 DVDD.n3259 4.5005
R7394 DVDD.n3285 DVDD.n3236 4.5005
R7395 DVDD.n3287 DVDD.n3236 4.5005
R7396 DVDD.n3284 DVDD.n3236 4.5005
R7397 DVDD.n3289 DVDD.n3236 4.5005
R7398 DVDD.n3283 DVDD.n3236 4.5005
R7399 DVDD.n3236 DVDD.n3235 4.5005
R7400 DVDD.n15909 DVDD.n3236 4.5005
R7401 DVDD.n3290 DVDD.n3236 4.5005
R7402 DVDD.n3281 DVDD.n3236 4.5005
R7403 DVDD.n3291 DVDD.n3236 4.5005
R7404 DVDD.n3280 DVDD.n3236 4.5005
R7405 DVDD.n3293 DVDD.n3236 4.5005
R7406 DVDD.n3279 DVDD.n3236 4.5005
R7407 DVDD.n3294 DVDD.n3236 4.5005
R7408 DVDD.n15907 DVDD.n3236 4.5005
R7409 DVDD.n15908 DVDD.n3285 4.5005
R7410 DVDD.n15908 DVDD.n3287 4.5005
R7411 DVDD.n15908 DVDD.n3284 4.5005
R7412 DVDD.n15908 DVDD.n3289 4.5005
R7413 DVDD.n15908 DVDD.n3283 4.5005
R7414 DVDD.n15908 DVDD.n3235 4.5005
R7415 DVDD.n15909 DVDD.n15908 4.5005
R7416 DVDD.n15908 DVDD.n3290 4.5005
R7417 DVDD.n15908 DVDD.n3281 4.5005
R7418 DVDD.n15908 DVDD.n3291 4.5005
R7419 DVDD.n15908 DVDD.n3280 4.5005
R7420 DVDD.n15908 DVDD.n3293 4.5005
R7421 DVDD.n15908 DVDD.n3279 4.5005
R7422 DVDD.n15908 DVDD.n3294 4.5005
R7423 DVDD.n15908 DVDD.n3272 4.5005
R7424 DVDD.n15908 DVDD.n15907 4.5005
R7425 DVDD.n3395 DVDD.n3260 4.5005
R7426 DVDD.n3397 DVDD.n3260 4.5005
R7427 DVDD.n3394 DVDD.n3260 4.5005
R7428 DVDD.n3400 DVDD.n3260 4.5005
R7429 DVDD.n3392 DVDD.n3260 4.5005
R7430 DVDD.n3401 DVDD.n3260 4.5005
R7431 DVDD.n3391 DVDD.n3260 4.5005
R7432 DVDD.n3402 DVDD.n3260 4.5005
R7433 DVDD.n3390 DVDD.n3260 4.5005
R7434 DVDD.n15837 DVDD.n3260 4.5005
R7435 DVDD.n3381 DVDD.n3260 4.5005
R7436 DVDD.n15839 DVDD.n3260 4.5005
R7437 DVDD.n3395 DVDD.n3359 4.5005
R7438 DVDD.n3397 DVDD.n3359 4.5005
R7439 DVDD.n3394 DVDD.n3359 4.5005
R7440 DVDD.n3399 DVDD.n3359 4.5005
R7441 DVDD.n3393 DVDD.n3359 4.5005
R7442 DVDD.n3400 DVDD.n3359 4.5005
R7443 DVDD.n3392 DVDD.n3359 4.5005
R7444 DVDD.n3401 DVDD.n3359 4.5005
R7445 DVDD.n3391 DVDD.n3359 4.5005
R7446 DVDD.n3402 DVDD.n3359 4.5005
R7447 DVDD.n3390 DVDD.n3359 4.5005
R7448 DVDD.n3404 DVDD.n3359 4.5005
R7449 DVDD.n3389 DVDD.n3359 4.5005
R7450 DVDD.n15837 DVDD.n3359 4.5005
R7451 DVDD.n15839 DVDD.n3359 4.5005
R7452 DVDD.n3395 DVDD.n3358 4.5005
R7453 DVDD.n3397 DVDD.n3358 4.5005
R7454 DVDD.n3394 DVDD.n3358 4.5005
R7455 DVDD.n3399 DVDD.n3358 4.5005
R7456 DVDD.n3393 DVDD.n3358 4.5005
R7457 DVDD.n3400 DVDD.n3358 4.5005
R7458 DVDD.n3392 DVDD.n3358 4.5005
R7459 DVDD.n3401 DVDD.n3358 4.5005
R7460 DVDD.n3391 DVDD.n3358 4.5005
R7461 DVDD.n3402 DVDD.n3358 4.5005
R7462 DVDD.n3390 DVDD.n3358 4.5005
R7463 DVDD.n3404 DVDD.n3358 4.5005
R7464 DVDD.n15837 DVDD.n3358 4.5005
R7465 DVDD.n15839 DVDD.n3358 4.5005
R7466 DVDD.n3395 DVDD.n3360 4.5005
R7467 DVDD.n3397 DVDD.n3360 4.5005
R7468 DVDD.n3394 DVDD.n3360 4.5005
R7469 DVDD.n3399 DVDD.n3360 4.5005
R7470 DVDD.n3393 DVDD.n3360 4.5005
R7471 DVDD.n3400 DVDD.n3360 4.5005
R7472 DVDD.n3392 DVDD.n3360 4.5005
R7473 DVDD.n3401 DVDD.n3360 4.5005
R7474 DVDD.n3391 DVDD.n3360 4.5005
R7475 DVDD.n3402 DVDD.n3360 4.5005
R7476 DVDD.n3390 DVDD.n3360 4.5005
R7477 DVDD.n3404 DVDD.n3360 4.5005
R7478 DVDD.n15837 DVDD.n3360 4.5005
R7479 DVDD.n15839 DVDD.n3360 4.5005
R7480 DVDD.n3395 DVDD.n3357 4.5005
R7481 DVDD.n3397 DVDD.n3357 4.5005
R7482 DVDD.n3394 DVDD.n3357 4.5005
R7483 DVDD.n3399 DVDD.n3357 4.5005
R7484 DVDD.n3393 DVDD.n3357 4.5005
R7485 DVDD.n3400 DVDD.n3357 4.5005
R7486 DVDD.n3392 DVDD.n3357 4.5005
R7487 DVDD.n3401 DVDD.n3357 4.5005
R7488 DVDD.n3391 DVDD.n3357 4.5005
R7489 DVDD.n3402 DVDD.n3357 4.5005
R7490 DVDD.n3390 DVDD.n3357 4.5005
R7491 DVDD.n3404 DVDD.n3357 4.5005
R7492 DVDD.n3389 DVDD.n3357 4.5005
R7493 DVDD.n15837 DVDD.n3357 4.5005
R7494 DVDD.n15839 DVDD.n3357 4.5005
R7495 DVDD.n3395 DVDD.n3361 4.5005
R7496 DVDD.n3397 DVDD.n3361 4.5005
R7497 DVDD.n3394 DVDD.n3361 4.5005
R7498 DVDD.n3399 DVDD.n3361 4.5005
R7499 DVDD.n3393 DVDD.n3361 4.5005
R7500 DVDD.n3400 DVDD.n3361 4.5005
R7501 DVDD.n3392 DVDD.n3361 4.5005
R7502 DVDD.n3401 DVDD.n3361 4.5005
R7503 DVDD.n3391 DVDD.n3361 4.5005
R7504 DVDD.n3402 DVDD.n3361 4.5005
R7505 DVDD.n3390 DVDD.n3361 4.5005
R7506 DVDD.n3404 DVDD.n3361 4.5005
R7507 DVDD.n3389 DVDD.n3361 4.5005
R7508 DVDD.n15837 DVDD.n3361 4.5005
R7509 DVDD.n15839 DVDD.n3361 4.5005
R7510 DVDD.n3395 DVDD.n3356 4.5005
R7511 DVDD.n3397 DVDD.n3356 4.5005
R7512 DVDD.n3394 DVDD.n3356 4.5005
R7513 DVDD.n3399 DVDD.n3356 4.5005
R7514 DVDD.n3393 DVDD.n3356 4.5005
R7515 DVDD.n3400 DVDD.n3356 4.5005
R7516 DVDD.n3392 DVDD.n3356 4.5005
R7517 DVDD.n3401 DVDD.n3356 4.5005
R7518 DVDD.n3391 DVDD.n3356 4.5005
R7519 DVDD.n3402 DVDD.n3356 4.5005
R7520 DVDD.n3390 DVDD.n3356 4.5005
R7521 DVDD.n3404 DVDD.n3356 4.5005
R7522 DVDD.n15837 DVDD.n3356 4.5005
R7523 DVDD.n15839 DVDD.n3356 4.5005
R7524 DVDD.n3395 DVDD.n3362 4.5005
R7525 DVDD.n3397 DVDD.n3362 4.5005
R7526 DVDD.n3394 DVDD.n3362 4.5005
R7527 DVDD.n3399 DVDD.n3362 4.5005
R7528 DVDD.n3393 DVDD.n3362 4.5005
R7529 DVDD.n3400 DVDD.n3362 4.5005
R7530 DVDD.n3392 DVDD.n3362 4.5005
R7531 DVDD.n3401 DVDD.n3362 4.5005
R7532 DVDD.n3391 DVDD.n3362 4.5005
R7533 DVDD.n3402 DVDD.n3362 4.5005
R7534 DVDD.n3390 DVDD.n3362 4.5005
R7535 DVDD.n3404 DVDD.n3362 4.5005
R7536 DVDD.n15837 DVDD.n3362 4.5005
R7537 DVDD.n15839 DVDD.n3362 4.5005
R7538 DVDD.n3395 DVDD.n3355 4.5005
R7539 DVDD.n3397 DVDD.n3355 4.5005
R7540 DVDD.n3394 DVDD.n3355 4.5005
R7541 DVDD.n3399 DVDD.n3355 4.5005
R7542 DVDD.n3393 DVDD.n3355 4.5005
R7543 DVDD.n3400 DVDD.n3355 4.5005
R7544 DVDD.n3392 DVDD.n3355 4.5005
R7545 DVDD.n3401 DVDD.n3355 4.5005
R7546 DVDD.n3391 DVDD.n3355 4.5005
R7547 DVDD.n3402 DVDD.n3355 4.5005
R7548 DVDD.n3390 DVDD.n3355 4.5005
R7549 DVDD.n3404 DVDD.n3355 4.5005
R7550 DVDD.n3389 DVDD.n3355 4.5005
R7551 DVDD.n15837 DVDD.n3355 4.5005
R7552 DVDD.n15839 DVDD.n3355 4.5005
R7553 DVDD.n3395 DVDD.n3363 4.5005
R7554 DVDD.n3397 DVDD.n3363 4.5005
R7555 DVDD.n3394 DVDD.n3363 4.5005
R7556 DVDD.n3399 DVDD.n3363 4.5005
R7557 DVDD.n3393 DVDD.n3363 4.5005
R7558 DVDD.n3400 DVDD.n3363 4.5005
R7559 DVDD.n3392 DVDD.n3363 4.5005
R7560 DVDD.n3401 DVDD.n3363 4.5005
R7561 DVDD.n3391 DVDD.n3363 4.5005
R7562 DVDD.n3402 DVDD.n3363 4.5005
R7563 DVDD.n3390 DVDD.n3363 4.5005
R7564 DVDD.n3404 DVDD.n3363 4.5005
R7565 DVDD.n3389 DVDD.n3363 4.5005
R7566 DVDD.n15837 DVDD.n3363 4.5005
R7567 DVDD.n15839 DVDD.n3363 4.5005
R7568 DVDD.n3395 DVDD.n3354 4.5005
R7569 DVDD.n3397 DVDD.n3354 4.5005
R7570 DVDD.n3394 DVDD.n3354 4.5005
R7571 DVDD.n3399 DVDD.n3354 4.5005
R7572 DVDD.n3393 DVDD.n3354 4.5005
R7573 DVDD.n3400 DVDD.n3354 4.5005
R7574 DVDD.n3392 DVDD.n3354 4.5005
R7575 DVDD.n3401 DVDD.n3354 4.5005
R7576 DVDD.n3391 DVDD.n3354 4.5005
R7577 DVDD.n3402 DVDD.n3354 4.5005
R7578 DVDD.n3390 DVDD.n3354 4.5005
R7579 DVDD.n3404 DVDD.n3354 4.5005
R7580 DVDD.n15837 DVDD.n3354 4.5005
R7581 DVDD.n15839 DVDD.n3354 4.5005
R7582 DVDD.n3395 DVDD.n3364 4.5005
R7583 DVDD.n3397 DVDD.n3364 4.5005
R7584 DVDD.n3394 DVDD.n3364 4.5005
R7585 DVDD.n3399 DVDD.n3364 4.5005
R7586 DVDD.n3393 DVDD.n3364 4.5005
R7587 DVDD.n3400 DVDD.n3364 4.5005
R7588 DVDD.n3392 DVDD.n3364 4.5005
R7589 DVDD.n3401 DVDD.n3364 4.5005
R7590 DVDD.n3391 DVDD.n3364 4.5005
R7591 DVDD.n3402 DVDD.n3364 4.5005
R7592 DVDD.n3390 DVDD.n3364 4.5005
R7593 DVDD.n3404 DVDD.n3364 4.5005
R7594 DVDD.n15837 DVDD.n3364 4.5005
R7595 DVDD.n15839 DVDD.n3364 4.5005
R7596 DVDD.n3395 DVDD.n3353 4.5005
R7597 DVDD.n3397 DVDD.n3353 4.5005
R7598 DVDD.n3394 DVDD.n3353 4.5005
R7599 DVDD.n3399 DVDD.n3353 4.5005
R7600 DVDD.n3393 DVDD.n3353 4.5005
R7601 DVDD.n3400 DVDD.n3353 4.5005
R7602 DVDD.n3392 DVDD.n3353 4.5005
R7603 DVDD.n3401 DVDD.n3353 4.5005
R7604 DVDD.n3391 DVDD.n3353 4.5005
R7605 DVDD.n3402 DVDD.n3353 4.5005
R7606 DVDD.n3390 DVDD.n3353 4.5005
R7607 DVDD.n3404 DVDD.n3353 4.5005
R7608 DVDD.n15837 DVDD.n3353 4.5005
R7609 DVDD.n15839 DVDD.n3353 4.5005
R7610 DVDD.n3395 DVDD.n3365 4.5005
R7611 DVDD.n3397 DVDD.n3365 4.5005
R7612 DVDD.n3394 DVDD.n3365 4.5005
R7613 DVDD.n3399 DVDD.n3365 4.5005
R7614 DVDD.n3393 DVDD.n3365 4.5005
R7615 DVDD.n3400 DVDD.n3365 4.5005
R7616 DVDD.n3392 DVDD.n3365 4.5005
R7617 DVDD.n3401 DVDD.n3365 4.5005
R7618 DVDD.n3391 DVDD.n3365 4.5005
R7619 DVDD.n3402 DVDD.n3365 4.5005
R7620 DVDD.n3390 DVDD.n3365 4.5005
R7621 DVDD.n3404 DVDD.n3365 4.5005
R7622 DVDD.n15837 DVDD.n3365 4.5005
R7623 DVDD.n15839 DVDD.n3365 4.5005
R7624 DVDD.n3395 DVDD.n3352 4.5005
R7625 DVDD.n3397 DVDD.n3352 4.5005
R7626 DVDD.n3394 DVDD.n3352 4.5005
R7627 DVDD.n3399 DVDD.n3352 4.5005
R7628 DVDD.n3393 DVDD.n3352 4.5005
R7629 DVDD.n3400 DVDD.n3352 4.5005
R7630 DVDD.n3392 DVDD.n3352 4.5005
R7631 DVDD.n3401 DVDD.n3352 4.5005
R7632 DVDD.n3391 DVDD.n3352 4.5005
R7633 DVDD.n3402 DVDD.n3352 4.5005
R7634 DVDD.n3390 DVDD.n3352 4.5005
R7635 DVDD.n3404 DVDD.n3352 4.5005
R7636 DVDD.n15837 DVDD.n3352 4.5005
R7637 DVDD.n15839 DVDD.n3352 4.5005
R7638 DVDD.n3395 DVDD.n3366 4.5005
R7639 DVDD.n3397 DVDD.n3366 4.5005
R7640 DVDD.n3394 DVDD.n3366 4.5005
R7641 DVDD.n3399 DVDD.n3366 4.5005
R7642 DVDD.n3393 DVDD.n3366 4.5005
R7643 DVDD.n3400 DVDD.n3366 4.5005
R7644 DVDD.n3392 DVDD.n3366 4.5005
R7645 DVDD.n3401 DVDD.n3366 4.5005
R7646 DVDD.n3391 DVDD.n3366 4.5005
R7647 DVDD.n3402 DVDD.n3366 4.5005
R7648 DVDD.n3390 DVDD.n3366 4.5005
R7649 DVDD.n3404 DVDD.n3366 4.5005
R7650 DVDD.n15837 DVDD.n3366 4.5005
R7651 DVDD.n15839 DVDD.n3366 4.5005
R7652 DVDD.n3395 DVDD.n3351 4.5005
R7653 DVDD.n3397 DVDD.n3351 4.5005
R7654 DVDD.n3394 DVDD.n3351 4.5005
R7655 DVDD.n3399 DVDD.n3351 4.5005
R7656 DVDD.n3393 DVDD.n3351 4.5005
R7657 DVDD.n3400 DVDD.n3351 4.5005
R7658 DVDD.n3392 DVDD.n3351 4.5005
R7659 DVDD.n3401 DVDD.n3351 4.5005
R7660 DVDD.n3391 DVDD.n3351 4.5005
R7661 DVDD.n3402 DVDD.n3351 4.5005
R7662 DVDD.n3390 DVDD.n3351 4.5005
R7663 DVDD.n3404 DVDD.n3351 4.5005
R7664 DVDD.n3389 DVDD.n3351 4.5005
R7665 DVDD.n15837 DVDD.n3351 4.5005
R7666 DVDD.n15839 DVDD.n3351 4.5005
R7667 DVDD.n3395 DVDD.n3367 4.5005
R7668 DVDD.n3397 DVDD.n3367 4.5005
R7669 DVDD.n3394 DVDD.n3367 4.5005
R7670 DVDD.n3399 DVDD.n3367 4.5005
R7671 DVDD.n3393 DVDD.n3367 4.5005
R7672 DVDD.n3400 DVDD.n3367 4.5005
R7673 DVDD.n3392 DVDD.n3367 4.5005
R7674 DVDD.n3401 DVDD.n3367 4.5005
R7675 DVDD.n3391 DVDD.n3367 4.5005
R7676 DVDD.n3402 DVDD.n3367 4.5005
R7677 DVDD.n3390 DVDD.n3367 4.5005
R7678 DVDD.n3404 DVDD.n3367 4.5005
R7679 DVDD.n15837 DVDD.n3367 4.5005
R7680 DVDD.n15839 DVDD.n3367 4.5005
R7681 DVDD.n3395 DVDD.n3350 4.5005
R7682 DVDD.n3397 DVDD.n3350 4.5005
R7683 DVDD.n3394 DVDD.n3350 4.5005
R7684 DVDD.n3399 DVDD.n3350 4.5005
R7685 DVDD.n3393 DVDD.n3350 4.5005
R7686 DVDD.n3400 DVDD.n3350 4.5005
R7687 DVDD.n3392 DVDD.n3350 4.5005
R7688 DVDD.n3401 DVDD.n3350 4.5005
R7689 DVDD.n3391 DVDD.n3350 4.5005
R7690 DVDD.n3402 DVDD.n3350 4.5005
R7691 DVDD.n3390 DVDD.n3350 4.5005
R7692 DVDD.n3404 DVDD.n3350 4.5005
R7693 DVDD.n15837 DVDD.n3350 4.5005
R7694 DVDD.n15839 DVDD.n3350 4.5005
R7695 DVDD.n3395 DVDD.n3368 4.5005
R7696 DVDD.n3397 DVDD.n3368 4.5005
R7697 DVDD.n3394 DVDD.n3368 4.5005
R7698 DVDD.n3399 DVDD.n3368 4.5005
R7699 DVDD.n3393 DVDD.n3368 4.5005
R7700 DVDD.n3400 DVDD.n3368 4.5005
R7701 DVDD.n3392 DVDD.n3368 4.5005
R7702 DVDD.n3401 DVDD.n3368 4.5005
R7703 DVDD.n3391 DVDD.n3368 4.5005
R7704 DVDD.n3402 DVDD.n3368 4.5005
R7705 DVDD.n3390 DVDD.n3368 4.5005
R7706 DVDD.n3404 DVDD.n3368 4.5005
R7707 DVDD.n15837 DVDD.n3368 4.5005
R7708 DVDD.n15839 DVDD.n3368 4.5005
R7709 DVDD.n3395 DVDD.n3349 4.5005
R7710 DVDD.n3397 DVDD.n3349 4.5005
R7711 DVDD.n3394 DVDD.n3349 4.5005
R7712 DVDD.n3399 DVDD.n3349 4.5005
R7713 DVDD.n3393 DVDD.n3349 4.5005
R7714 DVDD.n3400 DVDD.n3349 4.5005
R7715 DVDD.n3392 DVDD.n3349 4.5005
R7716 DVDD.n3401 DVDD.n3349 4.5005
R7717 DVDD.n3391 DVDD.n3349 4.5005
R7718 DVDD.n3402 DVDD.n3349 4.5005
R7719 DVDD.n3390 DVDD.n3349 4.5005
R7720 DVDD.n3404 DVDD.n3349 4.5005
R7721 DVDD.n3389 DVDD.n3349 4.5005
R7722 DVDD.n15837 DVDD.n3349 4.5005
R7723 DVDD.n15839 DVDD.n3349 4.5005
R7724 DVDD.n4743 DVDD.n3728 4.5005
R7725 DVDD.n3733 DVDD.n3728 4.5005
R7726 DVDD.n4741 DVDD.n3728 4.5005
R7727 DVDD.n3735 DVDD.n3728 4.5005
R7728 DVDD.n3750 DVDD.n3728 4.5005
R7729 DVDD.n3736 DVDD.n3728 4.5005
R7730 DVDD.n3749 DVDD.n3728 4.5005
R7731 DVDD.n3737 DVDD.n3728 4.5005
R7732 DVDD.n3748 DVDD.n3728 4.5005
R7733 DVDD.n3739 DVDD.n3728 4.5005
R7734 DVDD.n4419 DVDD.n3728 4.5005
R7735 DVDD.n4743 DVDD.n3726 4.5005
R7736 DVDD.n3733 DVDD.n3726 4.5005
R7737 DVDD.n4741 DVDD.n3726 4.5005
R7738 DVDD.n3734 DVDD.n3726 4.5005
R7739 DVDD.n3752 DVDD.n3726 4.5005
R7740 DVDD.n3735 DVDD.n3726 4.5005
R7741 DVDD.n3750 DVDD.n3726 4.5005
R7742 DVDD.n3736 DVDD.n3726 4.5005
R7743 DVDD.n3749 DVDD.n3726 4.5005
R7744 DVDD.n3737 DVDD.n3726 4.5005
R7745 DVDD.n3748 DVDD.n3726 4.5005
R7746 DVDD.n3738 DVDD.n3726 4.5005
R7747 DVDD.n3739 DVDD.n3726 4.5005
R7748 DVDD.n4419 DVDD.n3726 4.5005
R7749 DVDD.n4419 DVDD.n3731 4.5005
R7750 DVDD.n4419 DVDD.n3724 4.5005
R7751 DVDD.n4419 DVDD.n3729 4.5005
R7752 DVDD.n3813 DVDD.n3783 4.5005
R7753 DVDD.n3814 DVDD.n3783 4.5005
R7754 DVDD.n3812 DVDD.n3783 4.5005
R7755 DVDD.n4158 DVDD.n3783 4.5005
R7756 DVDD.n3810 DVDD.n3783 4.5005
R7757 DVDD.n4159 DVDD.n3783 4.5005
R7758 DVDD.n3809 DVDD.n3783 4.5005
R7759 DVDD.n4161 DVDD.n3783 4.5005
R7760 DVDD.n3808 DVDD.n3783 4.5005
R7761 DVDD.n4177 DVDD.n3783 4.5005
R7762 DVDD.n4179 DVDD.n3783 4.5005
R7763 DVDD.n3813 DVDD.n3784 4.5005
R7764 DVDD.n3814 DVDD.n3784 4.5005
R7765 DVDD.n3812 DVDD.n3784 4.5005
R7766 DVDD.n3816 DVDD.n3784 4.5005
R7767 DVDD.n3811 DVDD.n3784 4.5005
R7768 DVDD.n4158 DVDD.n3784 4.5005
R7769 DVDD.n3810 DVDD.n3784 4.5005
R7770 DVDD.n4159 DVDD.n3784 4.5005
R7771 DVDD.n3809 DVDD.n3784 4.5005
R7772 DVDD.n4161 DVDD.n3784 4.5005
R7773 DVDD.n3808 DVDD.n3784 4.5005
R7774 DVDD.n4163 DVDD.n3784 4.5005
R7775 DVDD.n4177 DVDD.n3784 4.5005
R7776 DVDD.n4179 DVDD.n3784 4.5005
R7777 DVDD.n3813 DVDD.n3782 4.5005
R7778 DVDD.n3814 DVDD.n3782 4.5005
R7779 DVDD.n3812 DVDD.n3782 4.5005
R7780 DVDD.n3816 DVDD.n3782 4.5005
R7781 DVDD.n3811 DVDD.n3782 4.5005
R7782 DVDD.n4158 DVDD.n3782 4.5005
R7783 DVDD.n3810 DVDD.n3782 4.5005
R7784 DVDD.n4159 DVDD.n3782 4.5005
R7785 DVDD.n3809 DVDD.n3782 4.5005
R7786 DVDD.n4161 DVDD.n3782 4.5005
R7787 DVDD.n3808 DVDD.n3782 4.5005
R7788 DVDD.n4163 DVDD.n3782 4.5005
R7789 DVDD.n4177 DVDD.n3782 4.5005
R7790 DVDD.n4179 DVDD.n3782 4.5005
R7791 DVDD.n3813 DVDD.n3785 4.5005
R7792 DVDD.n3814 DVDD.n3785 4.5005
R7793 DVDD.n3812 DVDD.n3785 4.5005
R7794 DVDD.n3816 DVDD.n3785 4.5005
R7795 DVDD.n3811 DVDD.n3785 4.5005
R7796 DVDD.n4158 DVDD.n3785 4.5005
R7797 DVDD.n3810 DVDD.n3785 4.5005
R7798 DVDD.n4159 DVDD.n3785 4.5005
R7799 DVDD.n3809 DVDD.n3785 4.5005
R7800 DVDD.n4161 DVDD.n3785 4.5005
R7801 DVDD.n3808 DVDD.n3785 4.5005
R7802 DVDD.n4163 DVDD.n3785 4.5005
R7803 DVDD.n4177 DVDD.n3785 4.5005
R7804 DVDD.n4179 DVDD.n3785 4.5005
R7805 DVDD.n3813 DVDD.n3781 4.5005
R7806 DVDD.n3814 DVDD.n3781 4.5005
R7807 DVDD.n3812 DVDD.n3781 4.5005
R7808 DVDD.n3816 DVDD.n3781 4.5005
R7809 DVDD.n3811 DVDD.n3781 4.5005
R7810 DVDD.n4158 DVDD.n3781 4.5005
R7811 DVDD.n3810 DVDD.n3781 4.5005
R7812 DVDD.n4159 DVDD.n3781 4.5005
R7813 DVDD.n3809 DVDD.n3781 4.5005
R7814 DVDD.n4161 DVDD.n3781 4.5005
R7815 DVDD.n3808 DVDD.n3781 4.5005
R7816 DVDD.n4163 DVDD.n3781 4.5005
R7817 DVDD.n4177 DVDD.n3781 4.5005
R7818 DVDD.n4179 DVDD.n3781 4.5005
R7819 DVDD.n3813 DVDD.n3786 4.5005
R7820 DVDD.n3814 DVDD.n3786 4.5005
R7821 DVDD.n3812 DVDD.n3786 4.5005
R7822 DVDD.n3816 DVDD.n3786 4.5005
R7823 DVDD.n3811 DVDD.n3786 4.5005
R7824 DVDD.n4158 DVDD.n3786 4.5005
R7825 DVDD.n3810 DVDD.n3786 4.5005
R7826 DVDD.n4159 DVDD.n3786 4.5005
R7827 DVDD.n3809 DVDD.n3786 4.5005
R7828 DVDD.n4161 DVDD.n3786 4.5005
R7829 DVDD.n3808 DVDD.n3786 4.5005
R7830 DVDD.n4163 DVDD.n3786 4.5005
R7831 DVDD.n4177 DVDD.n3786 4.5005
R7832 DVDD.n4179 DVDD.n3786 4.5005
R7833 DVDD.n3813 DVDD.n3780 4.5005
R7834 DVDD.n3814 DVDD.n3780 4.5005
R7835 DVDD.n3812 DVDD.n3780 4.5005
R7836 DVDD.n3816 DVDD.n3780 4.5005
R7837 DVDD.n3811 DVDD.n3780 4.5005
R7838 DVDD.n4158 DVDD.n3780 4.5005
R7839 DVDD.n3810 DVDD.n3780 4.5005
R7840 DVDD.n4159 DVDD.n3780 4.5005
R7841 DVDD.n3809 DVDD.n3780 4.5005
R7842 DVDD.n4161 DVDD.n3780 4.5005
R7843 DVDD.n3808 DVDD.n3780 4.5005
R7844 DVDD.n4163 DVDD.n3780 4.5005
R7845 DVDD.n4177 DVDD.n3780 4.5005
R7846 DVDD.n4179 DVDD.n3780 4.5005
R7847 DVDD.n3813 DVDD.n3787 4.5005
R7848 DVDD.n3814 DVDD.n3787 4.5005
R7849 DVDD.n3812 DVDD.n3787 4.5005
R7850 DVDD.n3816 DVDD.n3787 4.5005
R7851 DVDD.n3811 DVDD.n3787 4.5005
R7852 DVDD.n4158 DVDD.n3787 4.5005
R7853 DVDD.n3810 DVDD.n3787 4.5005
R7854 DVDD.n4159 DVDD.n3787 4.5005
R7855 DVDD.n3809 DVDD.n3787 4.5005
R7856 DVDD.n4161 DVDD.n3787 4.5005
R7857 DVDD.n3808 DVDD.n3787 4.5005
R7858 DVDD.n4163 DVDD.n3787 4.5005
R7859 DVDD.n4177 DVDD.n3787 4.5005
R7860 DVDD.n4179 DVDD.n3787 4.5005
R7861 DVDD.n3813 DVDD.n3779 4.5005
R7862 DVDD.n3814 DVDD.n3779 4.5005
R7863 DVDD.n3812 DVDD.n3779 4.5005
R7864 DVDD.n3816 DVDD.n3779 4.5005
R7865 DVDD.n3811 DVDD.n3779 4.5005
R7866 DVDD.n4158 DVDD.n3779 4.5005
R7867 DVDD.n3810 DVDD.n3779 4.5005
R7868 DVDD.n4159 DVDD.n3779 4.5005
R7869 DVDD.n3809 DVDD.n3779 4.5005
R7870 DVDD.n4161 DVDD.n3779 4.5005
R7871 DVDD.n3808 DVDD.n3779 4.5005
R7872 DVDD.n4163 DVDD.n3779 4.5005
R7873 DVDD.n4177 DVDD.n3779 4.5005
R7874 DVDD.n4179 DVDD.n3779 4.5005
R7875 DVDD.n3813 DVDD.n3788 4.5005
R7876 DVDD.n3814 DVDD.n3788 4.5005
R7877 DVDD.n3812 DVDD.n3788 4.5005
R7878 DVDD.n3816 DVDD.n3788 4.5005
R7879 DVDD.n3811 DVDD.n3788 4.5005
R7880 DVDD.n4158 DVDD.n3788 4.5005
R7881 DVDD.n3810 DVDD.n3788 4.5005
R7882 DVDD.n4159 DVDD.n3788 4.5005
R7883 DVDD.n3809 DVDD.n3788 4.5005
R7884 DVDD.n4161 DVDD.n3788 4.5005
R7885 DVDD.n3808 DVDD.n3788 4.5005
R7886 DVDD.n4163 DVDD.n3788 4.5005
R7887 DVDD.n4177 DVDD.n3788 4.5005
R7888 DVDD.n4179 DVDD.n3788 4.5005
R7889 DVDD.n3813 DVDD.n3778 4.5005
R7890 DVDD.n3814 DVDD.n3778 4.5005
R7891 DVDD.n3812 DVDD.n3778 4.5005
R7892 DVDD.n3816 DVDD.n3778 4.5005
R7893 DVDD.n3811 DVDD.n3778 4.5005
R7894 DVDD.n4158 DVDD.n3778 4.5005
R7895 DVDD.n3810 DVDD.n3778 4.5005
R7896 DVDD.n4159 DVDD.n3778 4.5005
R7897 DVDD.n3809 DVDD.n3778 4.5005
R7898 DVDD.n4161 DVDD.n3778 4.5005
R7899 DVDD.n3808 DVDD.n3778 4.5005
R7900 DVDD.n4163 DVDD.n3778 4.5005
R7901 DVDD.n4177 DVDD.n3778 4.5005
R7902 DVDD.n4179 DVDD.n3778 4.5005
R7903 DVDD.n3813 DVDD.n3789 4.5005
R7904 DVDD.n3814 DVDD.n3789 4.5005
R7905 DVDD.n3812 DVDD.n3789 4.5005
R7906 DVDD.n3816 DVDD.n3789 4.5005
R7907 DVDD.n3811 DVDD.n3789 4.5005
R7908 DVDD.n4158 DVDD.n3789 4.5005
R7909 DVDD.n3810 DVDD.n3789 4.5005
R7910 DVDD.n4159 DVDD.n3789 4.5005
R7911 DVDD.n3809 DVDD.n3789 4.5005
R7912 DVDD.n4161 DVDD.n3789 4.5005
R7913 DVDD.n3808 DVDD.n3789 4.5005
R7914 DVDD.n4163 DVDD.n3789 4.5005
R7915 DVDD.n4177 DVDD.n3789 4.5005
R7916 DVDD.n4179 DVDD.n3789 4.5005
R7917 DVDD.n3813 DVDD.n3777 4.5005
R7918 DVDD.n3814 DVDD.n3777 4.5005
R7919 DVDD.n3812 DVDD.n3777 4.5005
R7920 DVDD.n3816 DVDD.n3777 4.5005
R7921 DVDD.n3811 DVDD.n3777 4.5005
R7922 DVDD.n4158 DVDD.n3777 4.5005
R7923 DVDD.n3810 DVDD.n3777 4.5005
R7924 DVDD.n4159 DVDD.n3777 4.5005
R7925 DVDD.n3809 DVDD.n3777 4.5005
R7926 DVDD.n4161 DVDD.n3777 4.5005
R7927 DVDD.n3808 DVDD.n3777 4.5005
R7928 DVDD.n4163 DVDD.n3777 4.5005
R7929 DVDD.n4177 DVDD.n3777 4.5005
R7930 DVDD.n4179 DVDD.n3777 4.5005
R7931 DVDD.n3813 DVDD.n3790 4.5005
R7932 DVDD.n3814 DVDD.n3790 4.5005
R7933 DVDD.n3812 DVDD.n3790 4.5005
R7934 DVDD.n3816 DVDD.n3790 4.5005
R7935 DVDD.n3811 DVDD.n3790 4.5005
R7936 DVDD.n4158 DVDD.n3790 4.5005
R7937 DVDD.n3810 DVDD.n3790 4.5005
R7938 DVDD.n4159 DVDD.n3790 4.5005
R7939 DVDD.n3809 DVDD.n3790 4.5005
R7940 DVDD.n4161 DVDD.n3790 4.5005
R7941 DVDD.n3808 DVDD.n3790 4.5005
R7942 DVDD.n4163 DVDD.n3790 4.5005
R7943 DVDD.n4177 DVDD.n3790 4.5005
R7944 DVDD.n4179 DVDD.n3790 4.5005
R7945 DVDD.n3813 DVDD.n3776 4.5005
R7946 DVDD.n3814 DVDD.n3776 4.5005
R7947 DVDD.n3812 DVDD.n3776 4.5005
R7948 DVDD.n3816 DVDD.n3776 4.5005
R7949 DVDD.n3811 DVDD.n3776 4.5005
R7950 DVDD.n4158 DVDD.n3776 4.5005
R7951 DVDD.n3810 DVDD.n3776 4.5005
R7952 DVDD.n4159 DVDD.n3776 4.5005
R7953 DVDD.n3809 DVDD.n3776 4.5005
R7954 DVDD.n4161 DVDD.n3776 4.5005
R7955 DVDD.n3808 DVDD.n3776 4.5005
R7956 DVDD.n4163 DVDD.n3776 4.5005
R7957 DVDD.n4177 DVDD.n3776 4.5005
R7958 DVDD.n4179 DVDD.n3776 4.5005
R7959 DVDD.n3813 DVDD.n3791 4.5005
R7960 DVDD.n3814 DVDD.n3791 4.5005
R7961 DVDD.n3812 DVDD.n3791 4.5005
R7962 DVDD.n3816 DVDD.n3791 4.5005
R7963 DVDD.n3811 DVDD.n3791 4.5005
R7964 DVDD.n4158 DVDD.n3791 4.5005
R7965 DVDD.n3810 DVDD.n3791 4.5005
R7966 DVDD.n4159 DVDD.n3791 4.5005
R7967 DVDD.n3809 DVDD.n3791 4.5005
R7968 DVDD.n4161 DVDD.n3791 4.5005
R7969 DVDD.n3808 DVDD.n3791 4.5005
R7970 DVDD.n4163 DVDD.n3791 4.5005
R7971 DVDD.n4177 DVDD.n3791 4.5005
R7972 DVDD.n4179 DVDD.n3791 4.5005
R7973 DVDD.n3813 DVDD.n3775 4.5005
R7974 DVDD.n3814 DVDD.n3775 4.5005
R7975 DVDD.n3812 DVDD.n3775 4.5005
R7976 DVDD.n3816 DVDD.n3775 4.5005
R7977 DVDD.n3811 DVDD.n3775 4.5005
R7978 DVDD.n4158 DVDD.n3775 4.5005
R7979 DVDD.n3810 DVDD.n3775 4.5005
R7980 DVDD.n4159 DVDD.n3775 4.5005
R7981 DVDD.n3809 DVDD.n3775 4.5005
R7982 DVDD.n4161 DVDD.n3775 4.5005
R7983 DVDD.n3808 DVDD.n3775 4.5005
R7984 DVDD.n4163 DVDD.n3775 4.5005
R7985 DVDD.n4177 DVDD.n3775 4.5005
R7986 DVDD.n4179 DVDD.n3775 4.5005
R7987 DVDD.n3813 DVDD.n3792 4.5005
R7988 DVDD.n3814 DVDD.n3792 4.5005
R7989 DVDD.n3812 DVDD.n3792 4.5005
R7990 DVDD.n3816 DVDD.n3792 4.5005
R7991 DVDD.n3811 DVDD.n3792 4.5005
R7992 DVDD.n4158 DVDD.n3792 4.5005
R7993 DVDD.n3810 DVDD.n3792 4.5005
R7994 DVDD.n4159 DVDD.n3792 4.5005
R7995 DVDD.n3809 DVDD.n3792 4.5005
R7996 DVDD.n4161 DVDD.n3792 4.5005
R7997 DVDD.n3808 DVDD.n3792 4.5005
R7998 DVDD.n4163 DVDD.n3792 4.5005
R7999 DVDD.n4177 DVDD.n3792 4.5005
R8000 DVDD.n4179 DVDD.n3792 4.5005
R8001 DVDD.n3813 DVDD.n3774 4.5005
R8002 DVDD.n3814 DVDD.n3774 4.5005
R8003 DVDD.n3812 DVDD.n3774 4.5005
R8004 DVDD.n3816 DVDD.n3774 4.5005
R8005 DVDD.n3811 DVDD.n3774 4.5005
R8006 DVDD.n4158 DVDD.n3774 4.5005
R8007 DVDD.n3810 DVDD.n3774 4.5005
R8008 DVDD.n4159 DVDD.n3774 4.5005
R8009 DVDD.n3809 DVDD.n3774 4.5005
R8010 DVDD.n4161 DVDD.n3774 4.5005
R8011 DVDD.n3808 DVDD.n3774 4.5005
R8012 DVDD.n4163 DVDD.n3774 4.5005
R8013 DVDD.n4177 DVDD.n3774 4.5005
R8014 DVDD.n4179 DVDD.n3774 4.5005
R8015 DVDD.n3813 DVDD.n3793 4.5005
R8016 DVDD.n3814 DVDD.n3793 4.5005
R8017 DVDD.n3812 DVDD.n3793 4.5005
R8018 DVDD.n3816 DVDD.n3793 4.5005
R8019 DVDD.n3811 DVDD.n3793 4.5005
R8020 DVDD.n4158 DVDD.n3793 4.5005
R8021 DVDD.n3810 DVDD.n3793 4.5005
R8022 DVDD.n4159 DVDD.n3793 4.5005
R8023 DVDD.n3809 DVDD.n3793 4.5005
R8024 DVDD.n4161 DVDD.n3793 4.5005
R8025 DVDD.n3808 DVDD.n3793 4.5005
R8026 DVDD.n4163 DVDD.n3793 4.5005
R8027 DVDD.n4177 DVDD.n3793 4.5005
R8028 DVDD.n4179 DVDD.n3793 4.5005
R8029 DVDD.n3813 DVDD.n3773 4.5005
R8030 DVDD.n3814 DVDD.n3773 4.5005
R8031 DVDD.n3812 DVDD.n3773 4.5005
R8032 DVDD.n3816 DVDD.n3773 4.5005
R8033 DVDD.n3811 DVDD.n3773 4.5005
R8034 DVDD.n4158 DVDD.n3773 4.5005
R8035 DVDD.n3810 DVDD.n3773 4.5005
R8036 DVDD.n4159 DVDD.n3773 4.5005
R8037 DVDD.n3809 DVDD.n3773 4.5005
R8038 DVDD.n4161 DVDD.n3773 4.5005
R8039 DVDD.n3808 DVDD.n3773 4.5005
R8040 DVDD.n4163 DVDD.n3773 4.5005
R8041 DVDD.n4177 DVDD.n3773 4.5005
R8042 DVDD.n4179 DVDD.n3773 4.5005
R8043 DVDD.n3813 DVDD.n3794 4.5005
R8044 DVDD.n3814 DVDD.n3794 4.5005
R8045 DVDD.n3812 DVDD.n3794 4.5005
R8046 DVDD.n3816 DVDD.n3794 4.5005
R8047 DVDD.n3811 DVDD.n3794 4.5005
R8048 DVDD.n4158 DVDD.n3794 4.5005
R8049 DVDD.n3810 DVDD.n3794 4.5005
R8050 DVDD.n4159 DVDD.n3794 4.5005
R8051 DVDD.n3809 DVDD.n3794 4.5005
R8052 DVDD.n4161 DVDD.n3794 4.5005
R8053 DVDD.n3808 DVDD.n3794 4.5005
R8054 DVDD.n4163 DVDD.n3794 4.5005
R8055 DVDD.n4177 DVDD.n3794 4.5005
R8056 DVDD.n4179 DVDD.n3794 4.5005
R8057 DVDD.n3813 DVDD.n3772 4.5005
R8058 DVDD.n3814 DVDD.n3772 4.5005
R8059 DVDD.n3812 DVDD.n3772 4.5005
R8060 DVDD.n3816 DVDD.n3772 4.5005
R8061 DVDD.n3811 DVDD.n3772 4.5005
R8062 DVDD.n4158 DVDD.n3772 4.5005
R8063 DVDD.n3810 DVDD.n3772 4.5005
R8064 DVDD.n4159 DVDD.n3772 4.5005
R8065 DVDD.n3809 DVDD.n3772 4.5005
R8066 DVDD.n4161 DVDD.n3772 4.5005
R8067 DVDD.n3808 DVDD.n3772 4.5005
R8068 DVDD.n4163 DVDD.n3772 4.5005
R8069 DVDD.n4177 DVDD.n3772 4.5005
R8070 DVDD.n4179 DVDD.n3772 4.5005
R8071 DVDD.n4178 DVDD.n3813 4.5005
R8072 DVDD.n4178 DVDD.n3814 4.5005
R8073 DVDD.n4178 DVDD.n3812 4.5005
R8074 DVDD.n4178 DVDD.n3816 4.5005
R8075 DVDD.n4178 DVDD.n3811 4.5005
R8076 DVDD.n4178 DVDD.n4158 4.5005
R8077 DVDD.n4178 DVDD.n3810 4.5005
R8078 DVDD.n4178 DVDD.n4159 4.5005
R8079 DVDD.n4178 DVDD.n3809 4.5005
R8080 DVDD.n4178 DVDD.n4161 4.5005
R8081 DVDD.n4178 DVDD.n3808 4.5005
R8082 DVDD.n4178 DVDD.n4163 4.5005
R8083 DVDD.n4178 DVDD.n3807 4.5005
R8084 DVDD.n4178 DVDD.n4177 4.5005
R8085 DVDD.n4179 DVDD.n4178 4.5005
R8086 DVDD.n260 DVDD.n243 4.5005
R8087 DVDD.n260 DVDD.n244 4.5005
R8088 DVDD.n260 DVDD.n242 4.5005
R8089 DVDD.n260 DVDD.n246 4.5005
R8090 DVDD.n260 DVDD.n240 4.5005
R8091 DVDD.n260 DVDD.n247 4.5005
R8092 DVDD.n260 DVDD.n239 4.5005
R8093 DVDD.n260 DVDD.n248 4.5005
R8094 DVDD.n260 DVDD.n238 4.5005
R8095 DVDD.n260 DVDD.n250 4.5005
R8096 DVDD.n22181 DVDD.n260 4.5005
R8097 DVDD.n256 DVDD.n243 4.5005
R8098 DVDD.n256 DVDD.n244 4.5005
R8099 DVDD.n256 DVDD.n242 4.5005
R8100 DVDD.n256 DVDD.n245 4.5005
R8101 DVDD.n256 DVDD.n241 4.5005
R8102 DVDD.n256 DVDD.n246 4.5005
R8103 DVDD.n256 DVDD.n240 4.5005
R8104 DVDD.n256 DVDD.n247 4.5005
R8105 DVDD.n256 DVDD.n239 4.5005
R8106 DVDD.n256 DVDD.n248 4.5005
R8107 DVDD.n256 DVDD.n238 4.5005
R8108 DVDD.n256 DVDD.n249 4.5005
R8109 DVDD.n256 DVDD.n250 4.5005
R8110 DVDD.n22181 DVDD.n256 4.5005
R8111 DVDD.n262 DVDD.n243 4.5005
R8112 DVDD.n262 DVDD.n244 4.5005
R8113 DVDD.n262 DVDD.n242 4.5005
R8114 DVDD.n262 DVDD.n245 4.5005
R8115 DVDD.n262 DVDD.n241 4.5005
R8116 DVDD.n262 DVDD.n246 4.5005
R8117 DVDD.n262 DVDD.n240 4.5005
R8118 DVDD.n262 DVDD.n247 4.5005
R8119 DVDD.n262 DVDD.n239 4.5005
R8120 DVDD.n262 DVDD.n248 4.5005
R8121 DVDD.n262 DVDD.n238 4.5005
R8122 DVDD.n262 DVDD.n249 4.5005
R8123 DVDD.n262 DVDD.n250 4.5005
R8124 DVDD.n22181 DVDD.n262 4.5005
R8125 DVDD.n255 DVDD.n243 4.5005
R8126 DVDD.n255 DVDD.n244 4.5005
R8127 DVDD.n255 DVDD.n242 4.5005
R8128 DVDD.n255 DVDD.n245 4.5005
R8129 DVDD.n255 DVDD.n241 4.5005
R8130 DVDD.n255 DVDD.n246 4.5005
R8131 DVDD.n255 DVDD.n240 4.5005
R8132 DVDD.n255 DVDD.n247 4.5005
R8133 DVDD.n255 DVDD.n239 4.5005
R8134 DVDD.n255 DVDD.n248 4.5005
R8135 DVDD.n255 DVDD.n238 4.5005
R8136 DVDD.n255 DVDD.n249 4.5005
R8137 DVDD.n255 DVDD.n250 4.5005
R8138 DVDD.n22181 DVDD.n255 4.5005
R8139 DVDD.n264 DVDD.n243 4.5005
R8140 DVDD.n264 DVDD.n244 4.5005
R8141 DVDD.n264 DVDD.n242 4.5005
R8142 DVDD.n264 DVDD.n245 4.5005
R8143 DVDD.n264 DVDD.n241 4.5005
R8144 DVDD.n264 DVDD.n246 4.5005
R8145 DVDD.n264 DVDD.n240 4.5005
R8146 DVDD.n264 DVDD.n247 4.5005
R8147 DVDD.n264 DVDD.n239 4.5005
R8148 DVDD.n264 DVDD.n248 4.5005
R8149 DVDD.n264 DVDD.n238 4.5005
R8150 DVDD.n264 DVDD.n249 4.5005
R8151 DVDD.n264 DVDD.n250 4.5005
R8152 DVDD.n22181 DVDD.n264 4.5005
R8153 DVDD.n254 DVDD.n243 4.5005
R8154 DVDD.n254 DVDD.n244 4.5005
R8155 DVDD.n254 DVDD.n242 4.5005
R8156 DVDD.n254 DVDD.n245 4.5005
R8157 DVDD.n254 DVDD.n241 4.5005
R8158 DVDD.n254 DVDD.n246 4.5005
R8159 DVDD.n254 DVDD.n240 4.5005
R8160 DVDD.n254 DVDD.n247 4.5005
R8161 DVDD.n254 DVDD.n239 4.5005
R8162 DVDD.n254 DVDD.n248 4.5005
R8163 DVDD.n254 DVDD.n238 4.5005
R8164 DVDD.n254 DVDD.n249 4.5005
R8165 DVDD.n254 DVDD.n250 4.5005
R8166 DVDD.n22181 DVDD.n254 4.5005
R8167 DVDD.n266 DVDD.n243 4.5005
R8168 DVDD.n266 DVDD.n244 4.5005
R8169 DVDD.n266 DVDD.n242 4.5005
R8170 DVDD.n266 DVDD.n245 4.5005
R8171 DVDD.n266 DVDD.n241 4.5005
R8172 DVDD.n266 DVDD.n246 4.5005
R8173 DVDD.n266 DVDD.n240 4.5005
R8174 DVDD.n266 DVDD.n247 4.5005
R8175 DVDD.n266 DVDD.n239 4.5005
R8176 DVDD.n266 DVDD.n248 4.5005
R8177 DVDD.n266 DVDD.n238 4.5005
R8178 DVDD.n266 DVDD.n249 4.5005
R8179 DVDD.n266 DVDD.n250 4.5005
R8180 DVDD.n22181 DVDD.n266 4.5005
R8181 DVDD.n253 DVDD.n243 4.5005
R8182 DVDD.n253 DVDD.n244 4.5005
R8183 DVDD.n253 DVDD.n242 4.5005
R8184 DVDD.n253 DVDD.n245 4.5005
R8185 DVDD.n253 DVDD.n241 4.5005
R8186 DVDD.n253 DVDD.n246 4.5005
R8187 DVDD.n253 DVDD.n240 4.5005
R8188 DVDD.n253 DVDD.n247 4.5005
R8189 DVDD.n253 DVDD.n239 4.5005
R8190 DVDD.n253 DVDD.n248 4.5005
R8191 DVDD.n253 DVDD.n238 4.5005
R8192 DVDD.n253 DVDD.n249 4.5005
R8193 DVDD.n253 DVDD.n250 4.5005
R8194 DVDD.n22181 DVDD.n253 4.5005
R8195 DVDD.n22180 DVDD.n243 4.5005
R8196 DVDD.n22180 DVDD.n244 4.5005
R8197 DVDD.n22180 DVDD.n242 4.5005
R8198 DVDD.n22180 DVDD.n245 4.5005
R8199 DVDD.n22180 DVDD.n241 4.5005
R8200 DVDD.n22180 DVDD.n246 4.5005
R8201 DVDD.n22180 DVDD.n240 4.5005
R8202 DVDD.n22180 DVDD.n247 4.5005
R8203 DVDD.n22180 DVDD.n239 4.5005
R8204 DVDD.n22180 DVDD.n248 4.5005
R8205 DVDD.n22180 DVDD.n238 4.5005
R8206 DVDD.n22180 DVDD.n249 4.5005
R8207 DVDD.n22180 DVDD.n250 4.5005
R8208 DVDD.n22181 DVDD.n22180 4.5005
R8209 DVDD.n252 DVDD.n243 4.5005
R8210 DVDD.n252 DVDD.n244 4.5005
R8211 DVDD.n252 DVDD.n242 4.5005
R8212 DVDD.n252 DVDD.n245 4.5005
R8213 DVDD.n252 DVDD.n241 4.5005
R8214 DVDD.n252 DVDD.n246 4.5005
R8215 DVDD.n252 DVDD.n240 4.5005
R8216 DVDD.n252 DVDD.n247 4.5005
R8217 DVDD.n252 DVDD.n239 4.5005
R8218 DVDD.n252 DVDD.n248 4.5005
R8219 DVDD.n252 DVDD.n238 4.5005
R8220 DVDD.n252 DVDD.n249 4.5005
R8221 DVDD.n252 DVDD.n250 4.5005
R8222 DVDD.n22181 DVDD.n252 4.5005
R8223 DVDD.n22182 DVDD.n243 4.5005
R8224 DVDD.n22182 DVDD.n244 4.5005
R8225 DVDD.n22182 DVDD.n242 4.5005
R8226 DVDD.n22182 DVDD.n245 4.5005
R8227 DVDD.n22182 DVDD.n241 4.5005
R8228 DVDD.n22182 DVDD.n246 4.5005
R8229 DVDD.n22182 DVDD.n240 4.5005
R8230 DVDD.n22182 DVDD.n247 4.5005
R8231 DVDD.n22182 DVDD.n239 4.5005
R8232 DVDD.n22182 DVDD.n248 4.5005
R8233 DVDD.n22182 DVDD.n238 4.5005
R8234 DVDD.n22182 DVDD.n249 4.5005
R8235 DVDD.n22182 DVDD.n250 4.5005
R8236 DVDD.n22182 DVDD.n236 4.5005
R8237 DVDD.n22182 DVDD.n22181 4.5005
R8238 DVDD.n19140 DVDD.n19124 4.5005
R8239 DVDD.n19141 DVDD.n19124 4.5005
R8240 DVDD.n19139 DVDD.n19124 4.5005
R8241 DVDD.n19144 DVDD.n19124 4.5005
R8242 DVDD.n19137 DVDD.n19124 4.5005
R8243 DVDD.n19145 DVDD.n19124 4.5005
R8244 DVDD.n19136 DVDD.n19124 4.5005
R8245 DVDD.n19146 DVDD.n19124 4.5005
R8246 DVDD.n19135 DVDD.n19124 4.5005
R8247 DVDD.n20734 DVDD.n19124 4.5005
R8248 DVDD.n19153 DVDD.n19124 4.5005
R8249 DVDD.n20736 DVDD.n19124 4.5005
R8250 DVDD.n19140 DVDD.n19078 4.5005
R8251 DVDD.n19141 DVDD.n19078 4.5005
R8252 DVDD.n19139 DVDD.n19078 4.5005
R8253 DVDD.n19143 DVDD.n19078 4.5005
R8254 DVDD.n19138 DVDD.n19078 4.5005
R8255 DVDD.n19144 DVDD.n19078 4.5005
R8256 DVDD.n19137 DVDD.n19078 4.5005
R8257 DVDD.n19145 DVDD.n19078 4.5005
R8258 DVDD.n19136 DVDD.n19078 4.5005
R8259 DVDD.n19146 DVDD.n19078 4.5005
R8260 DVDD.n19135 DVDD.n19078 4.5005
R8261 DVDD.n19148 DVDD.n19078 4.5005
R8262 DVDD.n19134 DVDD.n19078 4.5005
R8263 DVDD.n20734 DVDD.n19078 4.5005
R8264 DVDD.n20736 DVDD.n19078 4.5005
R8265 DVDD.n19140 DVDD.n19125 4.5005
R8266 DVDD.n19141 DVDD.n19125 4.5005
R8267 DVDD.n19139 DVDD.n19125 4.5005
R8268 DVDD.n19143 DVDD.n19125 4.5005
R8269 DVDD.n19138 DVDD.n19125 4.5005
R8270 DVDD.n19144 DVDD.n19125 4.5005
R8271 DVDD.n19137 DVDD.n19125 4.5005
R8272 DVDD.n19145 DVDD.n19125 4.5005
R8273 DVDD.n19136 DVDD.n19125 4.5005
R8274 DVDD.n19146 DVDD.n19125 4.5005
R8275 DVDD.n19135 DVDD.n19125 4.5005
R8276 DVDD.n19148 DVDD.n19125 4.5005
R8277 DVDD.n20734 DVDD.n19125 4.5005
R8278 DVDD.n20736 DVDD.n19125 4.5005
R8279 DVDD.n19140 DVDD.n19077 4.5005
R8280 DVDD.n19141 DVDD.n19077 4.5005
R8281 DVDD.n19139 DVDD.n19077 4.5005
R8282 DVDD.n19143 DVDD.n19077 4.5005
R8283 DVDD.n19138 DVDD.n19077 4.5005
R8284 DVDD.n19144 DVDD.n19077 4.5005
R8285 DVDD.n19137 DVDD.n19077 4.5005
R8286 DVDD.n19145 DVDD.n19077 4.5005
R8287 DVDD.n19136 DVDD.n19077 4.5005
R8288 DVDD.n19146 DVDD.n19077 4.5005
R8289 DVDD.n19135 DVDD.n19077 4.5005
R8290 DVDD.n19148 DVDD.n19077 4.5005
R8291 DVDD.n20734 DVDD.n19077 4.5005
R8292 DVDD.n20736 DVDD.n19077 4.5005
R8293 DVDD.n19140 DVDD.n19126 4.5005
R8294 DVDD.n19141 DVDD.n19126 4.5005
R8295 DVDD.n19139 DVDD.n19126 4.5005
R8296 DVDD.n19143 DVDD.n19126 4.5005
R8297 DVDD.n19138 DVDD.n19126 4.5005
R8298 DVDD.n19144 DVDD.n19126 4.5005
R8299 DVDD.n19137 DVDD.n19126 4.5005
R8300 DVDD.n19145 DVDD.n19126 4.5005
R8301 DVDD.n19136 DVDD.n19126 4.5005
R8302 DVDD.n19146 DVDD.n19126 4.5005
R8303 DVDD.n19135 DVDD.n19126 4.5005
R8304 DVDD.n19148 DVDD.n19126 4.5005
R8305 DVDD.n20734 DVDD.n19126 4.5005
R8306 DVDD.n20736 DVDD.n19126 4.5005
R8307 DVDD.n19140 DVDD.n19076 4.5005
R8308 DVDD.n19141 DVDD.n19076 4.5005
R8309 DVDD.n19139 DVDD.n19076 4.5005
R8310 DVDD.n19143 DVDD.n19076 4.5005
R8311 DVDD.n19138 DVDD.n19076 4.5005
R8312 DVDD.n19144 DVDD.n19076 4.5005
R8313 DVDD.n19137 DVDD.n19076 4.5005
R8314 DVDD.n19145 DVDD.n19076 4.5005
R8315 DVDD.n19136 DVDD.n19076 4.5005
R8316 DVDD.n19146 DVDD.n19076 4.5005
R8317 DVDD.n19135 DVDD.n19076 4.5005
R8318 DVDD.n19148 DVDD.n19076 4.5005
R8319 DVDD.n20734 DVDD.n19076 4.5005
R8320 DVDD.n20736 DVDD.n19076 4.5005
R8321 DVDD.n19140 DVDD.n19127 4.5005
R8322 DVDD.n19141 DVDD.n19127 4.5005
R8323 DVDD.n19139 DVDD.n19127 4.5005
R8324 DVDD.n19143 DVDD.n19127 4.5005
R8325 DVDD.n19138 DVDD.n19127 4.5005
R8326 DVDD.n19144 DVDD.n19127 4.5005
R8327 DVDD.n19137 DVDD.n19127 4.5005
R8328 DVDD.n19145 DVDD.n19127 4.5005
R8329 DVDD.n19136 DVDD.n19127 4.5005
R8330 DVDD.n19146 DVDD.n19127 4.5005
R8331 DVDD.n19135 DVDD.n19127 4.5005
R8332 DVDD.n19148 DVDD.n19127 4.5005
R8333 DVDD.n19134 DVDD.n19127 4.5005
R8334 DVDD.n20734 DVDD.n19127 4.5005
R8335 DVDD.n20736 DVDD.n19127 4.5005
R8336 DVDD.n20736 DVDD.n19075 4.5005
R8337 DVDD.n20736 DVDD.n19128 4.5005
R8338 DVDD.n19140 DVDD.n19074 4.5005
R8339 DVDD.n19141 DVDD.n19074 4.5005
R8340 DVDD.n19139 DVDD.n19074 4.5005
R8341 DVDD.n19143 DVDD.n19074 4.5005
R8342 DVDD.n19138 DVDD.n19074 4.5005
R8343 DVDD.n19144 DVDD.n19074 4.5005
R8344 DVDD.n19137 DVDD.n19074 4.5005
R8345 DVDD.n19145 DVDD.n19074 4.5005
R8346 DVDD.n19136 DVDD.n19074 4.5005
R8347 DVDD.n19146 DVDD.n19074 4.5005
R8348 DVDD.n19135 DVDD.n19074 4.5005
R8349 DVDD.n19148 DVDD.n19074 4.5005
R8350 DVDD.n20734 DVDD.n19074 4.5005
R8351 DVDD.n20736 DVDD.n19074 4.5005
R8352 DVDD.n20735 DVDD.n19140 4.5005
R8353 DVDD.n20735 DVDD.n19141 4.5005
R8354 DVDD.n20735 DVDD.n19139 4.5005
R8355 DVDD.n20735 DVDD.n19143 4.5005
R8356 DVDD.n20735 DVDD.n19138 4.5005
R8357 DVDD.n20735 DVDD.n19144 4.5005
R8358 DVDD.n20735 DVDD.n19137 4.5005
R8359 DVDD.n20735 DVDD.n19145 4.5005
R8360 DVDD.n20735 DVDD.n19136 4.5005
R8361 DVDD.n20735 DVDD.n19146 4.5005
R8362 DVDD.n20735 DVDD.n19135 4.5005
R8363 DVDD.n20735 DVDD.n19148 4.5005
R8364 DVDD.n20735 DVDD.n19134 4.5005
R8365 DVDD.n20735 DVDD.n20734 4.5005
R8366 DVDD.n20736 DVDD.n20735 4.5005
R8367 DVDD.n19977 DVDD.n19964 4.5005
R8368 DVDD.n20023 DVDD.n19964 4.5005
R8369 DVDD.n19976 DVDD.n19964 4.5005
R8370 DVDD.n20026 DVDD.n19964 4.5005
R8371 DVDD.n19974 DVDD.n19964 4.5005
R8372 DVDD.n20027 DVDD.n19964 4.5005
R8373 DVDD.n19973 DVDD.n19964 4.5005
R8374 DVDD.n20028 DVDD.n19964 4.5005
R8375 DVDD.n19972 DVDD.n19964 4.5005
R8376 DVDD.n20242 DVDD.n19964 4.5005
R8377 DVDD.n19970 DVDD.n19964 4.5005
R8378 DVDD.n20244 DVDD.n19964 4.5005
R8379 DVDD.n19977 DVDD.n19963 4.5005
R8380 DVDD.n20023 DVDD.n19963 4.5005
R8381 DVDD.n19976 DVDD.n19963 4.5005
R8382 DVDD.n20025 DVDD.n19963 4.5005
R8383 DVDD.n19975 DVDD.n19963 4.5005
R8384 DVDD.n20026 DVDD.n19963 4.5005
R8385 DVDD.n19974 DVDD.n19963 4.5005
R8386 DVDD.n20027 DVDD.n19963 4.5005
R8387 DVDD.n19973 DVDD.n19963 4.5005
R8388 DVDD.n20028 DVDD.n19963 4.5005
R8389 DVDD.n19972 DVDD.n19963 4.5005
R8390 DVDD.n20030 DVDD.n19963 4.5005
R8391 DVDD.n19971 DVDD.n19963 4.5005
R8392 DVDD.n20242 DVDD.n19963 4.5005
R8393 DVDD.n19970 DVDD.n19963 4.5005
R8394 DVDD.n20244 DVDD.n19963 4.5005
R8395 DVDD.n19977 DVDD.n19965 4.5005
R8396 DVDD.n20023 DVDD.n19965 4.5005
R8397 DVDD.n19976 DVDD.n19965 4.5005
R8398 DVDD.n20025 DVDD.n19965 4.5005
R8399 DVDD.n19975 DVDD.n19965 4.5005
R8400 DVDD.n20026 DVDD.n19965 4.5005
R8401 DVDD.n19974 DVDD.n19965 4.5005
R8402 DVDD.n20027 DVDD.n19965 4.5005
R8403 DVDD.n19973 DVDD.n19965 4.5005
R8404 DVDD.n20028 DVDD.n19965 4.5005
R8405 DVDD.n19972 DVDD.n19965 4.5005
R8406 DVDD.n20030 DVDD.n19965 4.5005
R8407 DVDD.n19971 DVDD.n19965 4.5005
R8408 DVDD.n20242 DVDD.n19965 4.5005
R8409 DVDD.n19970 DVDD.n19965 4.5005
R8410 DVDD.n20244 DVDD.n19965 4.5005
R8411 DVDD.n19977 DVDD.n19962 4.5005
R8412 DVDD.n20023 DVDD.n19962 4.5005
R8413 DVDD.n19976 DVDD.n19962 4.5005
R8414 DVDD.n20025 DVDD.n19962 4.5005
R8415 DVDD.n19975 DVDD.n19962 4.5005
R8416 DVDD.n20026 DVDD.n19962 4.5005
R8417 DVDD.n19974 DVDD.n19962 4.5005
R8418 DVDD.n20027 DVDD.n19962 4.5005
R8419 DVDD.n19973 DVDD.n19962 4.5005
R8420 DVDD.n20028 DVDD.n19962 4.5005
R8421 DVDD.n19972 DVDD.n19962 4.5005
R8422 DVDD.n20030 DVDD.n19962 4.5005
R8423 DVDD.n19971 DVDD.n19962 4.5005
R8424 DVDD.n20242 DVDD.n19962 4.5005
R8425 DVDD.n19970 DVDD.n19962 4.5005
R8426 DVDD.n20244 DVDD.n19962 4.5005
R8427 DVDD.n19977 DVDD.n19966 4.5005
R8428 DVDD.n20023 DVDD.n19966 4.5005
R8429 DVDD.n19976 DVDD.n19966 4.5005
R8430 DVDD.n20025 DVDD.n19966 4.5005
R8431 DVDD.n19975 DVDD.n19966 4.5005
R8432 DVDD.n20026 DVDD.n19966 4.5005
R8433 DVDD.n19974 DVDD.n19966 4.5005
R8434 DVDD.n20027 DVDD.n19966 4.5005
R8435 DVDD.n19973 DVDD.n19966 4.5005
R8436 DVDD.n20028 DVDD.n19966 4.5005
R8437 DVDD.n19972 DVDD.n19966 4.5005
R8438 DVDD.n20030 DVDD.n19966 4.5005
R8439 DVDD.n19971 DVDD.n19966 4.5005
R8440 DVDD.n20242 DVDD.n19966 4.5005
R8441 DVDD.n19970 DVDD.n19966 4.5005
R8442 DVDD.n20244 DVDD.n19966 4.5005
R8443 DVDD.n19977 DVDD.n19961 4.5005
R8444 DVDD.n20023 DVDD.n19961 4.5005
R8445 DVDD.n19976 DVDD.n19961 4.5005
R8446 DVDD.n20025 DVDD.n19961 4.5005
R8447 DVDD.n19975 DVDD.n19961 4.5005
R8448 DVDD.n20026 DVDD.n19961 4.5005
R8449 DVDD.n19974 DVDD.n19961 4.5005
R8450 DVDD.n20027 DVDD.n19961 4.5005
R8451 DVDD.n19973 DVDD.n19961 4.5005
R8452 DVDD.n20028 DVDD.n19961 4.5005
R8453 DVDD.n19972 DVDD.n19961 4.5005
R8454 DVDD.n20030 DVDD.n19961 4.5005
R8455 DVDD.n19971 DVDD.n19961 4.5005
R8456 DVDD.n20242 DVDD.n19961 4.5005
R8457 DVDD.n19970 DVDD.n19961 4.5005
R8458 DVDD.n20244 DVDD.n19961 4.5005
R8459 DVDD.n19977 DVDD.n19967 4.5005
R8460 DVDD.n20023 DVDD.n19967 4.5005
R8461 DVDD.n19976 DVDD.n19967 4.5005
R8462 DVDD.n20025 DVDD.n19967 4.5005
R8463 DVDD.n19975 DVDD.n19967 4.5005
R8464 DVDD.n20026 DVDD.n19967 4.5005
R8465 DVDD.n19974 DVDD.n19967 4.5005
R8466 DVDD.n20027 DVDD.n19967 4.5005
R8467 DVDD.n19973 DVDD.n19967 4.5005
R8468 DVDD.n20028 DVDD.n19967 4.5005
R8469 DVDD.n19972 DVDD.n19967 4.5005
R8470 DVDD.n20030 DVDD.n19967 4.5005
R8471 DVDD.n19971 DVDD.n19967 4.5005
R8472 DVDD.n20242 DVDD.n19967 4.5005
R8473 DVDD.n19970 DVDD.n19967 4.5005
R8474 DVDD.n20244 DVDD.n19967 4.5005
R8475 DVDD.n19977 DVDD.n19960 4.5005
R8476 DVDD.n20023 DVDD.n19960 4.5005
R8477 DVDD.n19976 DVDD.n19960 4.5005
R8478 DVDD.n20025 DVDD.n19960 4.5005
R8479 DVDD.n19975 DVDD.n19960 4.5005
R8480 DVDD.n20026 DVDD.n19960 4.5005
R8481 DVDD.n19974 DVDD.n19960 4.5005
R8482 DVDD.n20027 DVDD.n19960 4.5005
R8483 DVDD.n19973 DVDD.n19960 4.5005
R8484 DVDD.n20028 DVDD.n19960 4.5005
R8485 DVDD.n19972 DVDD.n19960 4.5005
R8486 DVDD.n20030 DVDD.n19960 4.5005
R8487 DVDD.n19971 DVDD.n19960 4.5005
R8488 DVDD.n20242 DVDD.n19960 4.5005
R8489 DVDD.n19970 DVDD.n19960 4.5005
R8490 DVDD.n20244 DVDD.n19960 4.5005
R8491 DVDD.n19977 DVDD.n19968 4.5005
R8492 DVDD.n20023 DVDD.n19968 4.5005
R8493 DVDD.n19976 DVDD.n19968 4.5005
R8494 DVDD.n20025 DVDD.n19968 4.5005
R8495 DVDD.n19975 DVDD.n19968 4.5005
R8496 DVDD.n20026 DVDD.n19968 4.5005
R8497 DVDD.n19974 DVDD.n19968 4.5005
R8498 DVDD.n20027 DVDD.n19968 4.5005
R8499 DVDD.n19973 DVDD.n19968 4.5005
R8500 DVDD.n20028 DVDD.n19968 4.5005
R8501 DVDD.n19972 DVDD.n19968 4.5005
R8502 DVDD.n20030 DVDD.n19968 4.5005
R8503 DVDD.n19971 DVDD.n19968 4.5005
R8504 DVDD.n20242 DVDD.n19968 4.5005
R8505 DVDD.n19970 DVDD.n19968 4.5005
R8506 DVDD.n20244 DVDD.n19968 4.5005
R8507 DVDD.n19977 DVDD.n19959 4.5005
R8508 DVDD.n20023 DVDD.n19959 4.5005
R8509 DVDD.n19976 DVDD.n19959 4.5005
R8510 DVDD.n20025 DVDD.n19959 4.5005
R8511 DVDD.n19975 DVDD.n19959 4.5005
R8512 DVDD.n20026 DVDD.n19959 4.5005
R8513 DVDD.n19974 DVDD.n19959 4.5005
R8514 DVDD.n20027 DVDD.n19959 4.5005
R8515 DVDD.n19973 DVDD.n19959 4.5005
R8516 DVDD.n20028 DVDD.n19959 4.5005
R8517 DVDD.n19972 DVDD.n19959 4.5005
R8518 DVDD.n20030 DVDD.n19959 4.5005
R8519 DVDD.n19971 DVDD.n19959 4.5005
R8520 DVDD.n20242 DVDD.n19959 4.5005
R8521 DVDD.n19970 DVDD.n19959 4.5005
R8522 DVDD.n20244 DVDD.n19959 4.5005
R8523 DVDD.n20243 DVDD.n19977 4.5005
R8524 DVDD.n20243 DVDD.n20023 4.5005
R8525 DVDD.n20243 DVDD.n19976 4.5005
R8526 DVDD.n20243 DVDD.n20025 4.5005
R8527 DVDD.n20243 DVDD.n19975 4.5005
R8528 DVDD.n20243 DVDD.n20026 4.5005
R8529 DVDD.n20243 DVDD.n19974 4.5005
R8530 DVDD.n20243 DVDD.n20027 4.5005
R8531 DVDD.n20243 DVDD.n19973 4.5005
R8532 DVDD.n20243 DVDD.n20028 4.5005
R8533 DVDD.n20243 DVDD.n19972 4.5005
R8534 DVDD.n20243 DVDD.n20030 4.5005
R8535 DVDD.n20243 DVDD.n19971 4.5005
R8536 DVDD.n20243 DVDD.n20242 4.5005
R8537 DVDD.n20243 DVDD.n19970 4.5005
R8538 DVDD.n20244 DVDD.n20243 4.5005
R8539 DVDD.n19153 DVDD.n19128 4.5005
R8540 DVDD.n20734 DVDD.n19128 4.5005
R8541 DVDD.n19148 DVDD.n19128 4.5005
R8542 DVDD.n19135 DVDD.n19128 4.5005
R8543 DVDD.n19146 DVDD.n19128 4.5005
R8544 DVDD.n19136 DVDD.n19128 4.5005
R8545 DVDD.n19145 DVDD.n19128 4.5005
R8546 DVDD.n19137 DVDD.n19128 4.5005
R8547 DVDD.n19144 DVDD.n19128 4.5005
R8548 DVDD.n19138 DVDD.n19128 4.5005
R8549 DVDD.n19143 DVDD.n19128 4.5005
R8550 DVDD.n19139 DVDD.n19128 4.5005
R8551 DVDD.n19141 DVDD.n19128 4.5005
R8552 DVDD.n19140 DVDD.n19128 4.5005
R8553 DVDD.n19153 DVDD.n19075 4.5005
R8554 DVDD.n20734 DVDD.n19075 4.5005
R8555 DVDD.n19134 DVDD.n19075 4.5005
R8556 DVDD.n19148 DVDD.n19075 4.5005
R8557 DVDD.n19135 DVDD.n19075 4.5005
R8558 DVDD.n19146 DVDD.n19075 4.5005
R8559 DVDD.n19136 DVDD.n19075 4.5005
R8560 DVDD.n19145 DVDD.n19075 4.5005
R8561 DVDD.n19137 DVDD.n19075 4.5005
R8562 DVDD.n19144 DVDD.n19075 4.5005
R8563 DVDD.n19138 DVDD.n19075 4.5005
R8564 DVDD.n19143 DVDD.n19075 4.5005
R8565 DVDD.n19139 DVDD.n19075 4.5005
R8566 DVDD.n19141 DVDD.n19075 4.5005
R8567 DVDD.n19140 DVDD.n19075 4.5005
R8568 DVDD.n3739 DVDD.n3729 4.5005
R8569 DVDD.n4441 DVDD.n3729 4.5005
R8570 DVDD.n3739 DVDD.n3725 4.5005
R8571 DVDD.n4441 DVDD.n3725 4.5005
R8572 DVDD.n3739 DVDD.n3730 4.5005
R8573 DVDD.n4441 DVDD.n3730 4.5005
R8574 DVDD.n3739 DVDD.n3724 4.5005
R8575 DVDD.n4441 DVDD.n3724 4.5005
R8576 DVDD.n3739 DVDD.n3731 4.5005
R8577 DVDD.n4441 DVDD.n3731 4.5005
R8578 DVDD.n3739 DVDD.n3723 4.5005
R8579 DVDD.n4441 DVDD.n3723 4.5005
R8580 DVDD.n3739 DVDD.n3732 4.5005
R8581 DVDD.n4441 DVDD.n3732 4.5005
R8582 DVDD.n3739 DVDD.n3722 4.5005
R8583 DVDD.n4441 DVDD.n3722 4.5005
R8584 DVDD.n4742 DVDD.n3746 4.5005
R8585 DVDD.n4742 DVDD.n3739 4.5005
R8586 DVDD.n4742 DVDD.n3738 4.5005
R8587 DVDD.n3738 DVDD.n3722 4.5005
R8588 DVDD.n3738 DVDD.n3732 4.5005
R8589 DVDD.n3738 DVDD.n3723 4.5005
R8590 DVDD.n3738 DVDD.n3731 4.5005
R8591 DVDD.n3738 DVDD.n3724 4.5005
R8592 DVDD.n3738 DVDD.n3730 4.5005
R8593 DVDD.n3738 DVDD.n3725 4.5005
R8594 DVDD.n3738 DVDD.n3729 4.5005
R8595 DVDD.n3748 DVDD.n3729 4.5005
R8596 DVDD.n3737 DVDD.n3729 4.5005
R8597 DVDD.n3749 DVDD.n3729 4.5005
R8598 DVDD.n3748 DVDD.n3725 4.5005
R8599 DVDD.n3737 DVDD.n3725 4.5005
R8600 DVDD.n3749 DVDD.n3725 4.5005
R8601 DVDD.n3748 DVDD.n3730 4.5005
R8602 DVDD.n3737 DVDD.n3730 4.5005
R8603 DVDD.n3749 DVDD.n3730 4.5005
R8604 DVDD.n3748 DVDD.n3724 4.5005
R8605 DVDD.n3737 DVDD.n3724 4.5005
R8606 DVDD.n3749 DVDD.n3724 4.5005
R8607 DVDD.n3748 DVDD.n3731 4.5005
R8608 DVDD.n3737 DVDD.n3731 4.5005
R8609 DVDD.n3749 DVDD.n3731 4.5005
R8610 DVDD.n3748 DVDD.n3723 4.5005
R8611 DVDD.n3737 DVDD.n3723 4.5005
R8612 DVDD.n3749 DVDD.n3723 4.5005
R8613 DVDD.n3748 DVDD.n3732 4.5005
R8614 DVDD.n3737 DVDD.n3732 4.5005
R8615 DVDD.n3749 DVDD.n3732 4.5005
R8616 DVDD.n3748 DVDD.n3722 4.5005
R8617 DVDD.n3737 DVDD.n3722 4.5005
R8618 DVDD.n3749 DVDD.n3722 4.5005
R8619 DVDD.n4742 DVDD.n3748 4.5005
R8620 DVDD.n4742 DVDD.n3737 4.5005
R8621 DVDD.n4742 DVDD.n3749 4.5005
R8622 DVDD.n4742 DVDD.n3736 4.5005
R8623 DVDD.n3736 DVDD.n3722 4.5005
R8624 DVDD.n3736 DVDD.n3732 4.5005
R8625 DVDD.n3736 DVDD.n3723 4.5005
R8626 DVDD.n3736 DVDD.n3731 4.5005
R8627 DVDD.n3736 DVDD.n3724 4.5005
R8628 DVDD.n3736 DVDD.n3730 4.5005
R8629 DVDD.n3736 DVDD.n3725 4.5005
R8630 DVDD.n3736 DVDD.n3729 4.5005
R8631 DVDD.n3750 DVDD.n3729 4.5005
R8632 DVDD.n3735 DVDD.n3729 4.5005
R8633 DVDD.n3752 DVDD.n3729 4.5005
R8634 DVDD.n3750 DVDD.n3725 4.5005
R8635 DVDD.n3735 DVDD.n3725 4.5005
R8636 DVDD.n3752 DVDD.n3725 4.5005
R8637 DVDD.n3750 DVDD.n3730 4.5005
R8638 DVDD.n3735 DVDD.n3730 4.5005
R8639 DVDD.n3752 DVDD.n3730 4.5005
R8640 DVDD.n3750 DVDD.n3724 4.5005
R8641 DVDD.n3735 DVDD.n3724 4.5005
R8642 DVDD.n3752 DVDD.n3724 4.5005
R8643 DVDD.n3750 DVDD.n3731 4.5005
R8644 DVDD.n3735 DVDD.n3731 4.5005
R8645 DVDD.n3752 DVDD.n3731 4.5005
R8646 DVDD.n3750 DVDD.n3723 4.5005
R8647 DVDD.n3735 DVDD.n3723 4.5005
R8648 DVDD.n3752 DVDD.n3723 4.5005
R8649 DVDD.n3750 DVDD.n3732 4.5005
R8650 DVDD.n3735 DVDD.n3732 4.5005
R8651 DVDD.n3752 DVDD.n3732 4.5005
R8652 DVDD.n3750 DVDD.n3722 4.5005
R8653 DVDD.n3735 DVDD.n3722 4.5005
R8654 DVDD.n3752 DVDD.n3722 4.5005
R8655 DVDD.n4742 DVDD.n3750 4.5005
R8656 DVDD.n4742 DVDD.n3735 4.5005
R8657 DVDD.n4742 DVDD.n3752 4.5005
R8658 DVDD.n4742 DVDD.n3734 4.5005
R8659 DVDD.n3734 DVDD.n3722 4.5005
R8660 DVDD.n3734 DVDD.n3732 4.5005
R8661 DVDD.n3734 DVDD.n3723 4.5005
R8662 DVDD.n3734 DVDD.n3731 4.5005
R8663 DVDD.n3734 DVDD.n3724 4.5005
R8664 DVDD.n3734 DVDD.n3730 4.5005
R8665 DVDD.n3734 DVDD.n3725 4.5005
R8666 DVDD.n3734 DVDD.n3729 4.5005
R8667 DVDD.n4741 DVDD.n3729 4.5005
R8668 DVDD.n3733 DVDD.n3729 4.5005
R8669 DVDD.n4743 DVDD.n3729 4.5005
R8670 DVDD.n4741 DVDD.n3725 4.5005
R8671 DVDD.n3733 DVDD.n3725 4.5005
R8672 DVDD.n4743 DVDD.n3725 4.5005
R8673 DVDD.n4741 DVDD.n3730 4.5005
R8674 DVDD.n3733 DVDD.n3730 4.5005
R8675 DVDD.n4743 DVDD.n3730 4.5005
R8676 DVDD.n4741 DVDD.n3724 4.5005
R8677 DVDD.n3733 DVDD.n3724 4.5005
R8678 DVDD.n4743 DVDD.n3724 4.5005
R8679 DVDD.n4741 DVDD.n3731 4.5005
R8680 DVDD.n3733 DVDD.n3731 4.5005
R8681 DVDD.n4743 DVDD.n3731 4.5005
R8682 DVDD.n4741 DVDD.n3723 4.5005
R8683 DVDD.n3733 DVDD.n3723 4.5005
R8684 DVDD.n4743 DVDD.n3723 4.5005
R8685 DVDD.n4741 DVDD.n3732 4.5005
R8686 DVDD.n3733 DVDD.n3732 4.5005
R8687 DVDD.n4743 DVDD.n3732 4.5005
R8688 DVDD.n4741 DVDD.n3722 4.5005
R8689 DVDD.n3733 DVDD.n3722 4.5005
R8690 DVDD.n4743 DVDD.n3722 4.5005
R8691 DVDD.n4742 DVDD.n4741 4.5005
R8692 DVDD.n4742 DVDD.n3733 4.5005
R8693 DVDD.n4743 DVDD.n4742 4.5005
R8694 DVDD.n3395 DVDD.n3369 4.5005
R8695 DVDD.n3397 DVDD.n3369 4.5005
R8696 DVDD.n3394 DVDD.n3369 4.5005
R8697 DVDD.n3399 DVDD.n3369 4.5005
R8698 DVDD.n3393 DVDD.n3369 4.5005
R8699 DVDD.n3400 DVDD.n3369 4.5005
R8700 DVDD.n3392 DVDD.n3369 4.5005
R8701 DVDD.n3401 DVDD.n3369 4.5005
R8702 DVDD.n3391 DVDD.n3369 4.5005
R8703 DVDD.n3402 DVDD.n3369 4.5005
R8704 DVDD.n3390 DVDD.n3369 4.5005
R8705 DVDD.n3404 DVDD.n3369 4.5005
R8706 DVDD.n15837 DVDD.n3369 4.5005
R8707 DVDD.n3381 DVDD.n3369 4.5005
R8708 DVDD.n15839 DVDD.n3369 4.5005
R8709 DVDD.n3395 DVDD.n3348 4.5005
R8710 DVDD.n3397 DVDD.n3348 4.5005
R8711 DVDD.n3394 DVDD.n3348 4.5005
R8712 DVDD.n3399 DVDD.n3348 4.5005
R8713 DVDD.n3393 DVDD.n3348 4.5005
R8714 DVDD.n3400 DVDD.n3348 4.5005
R8715 DVDD.n3392 DVDD.n3348 4.5005
R8716 DVDD.n3401 DVDD.n3348 4.5005
R8717 DVDD.n3391 DVDD.n3348 4.5005
R8718 DVDD.n3402 DVDD.n3348 4.5005
R8719 DVDD.n3390 DVDD.n3348 4.5005
R8720 DVDD.n3404 DVDD.n3348 4.5005
R8721 DVDD.n3389 DVDD.n3348 4.5005
R8722 DVDD.n15837 DVDD.n3348 4.5005
R8723 DVDD.n3381 DVDD.n3348 4.5005
R8724 DVDD.n15839 DVDD.n3348 4.5005
R8725 DVDD.n15838 DVDD.n3395 4.5005
R8726 DVDD.n15838 DVDD.n3397 4.5005
R8727 DVDD.n15838 DVDD.n3394 4.5005
R8728 DVDD.n15838 DVDD.n3399 4.5005
R8729 DVDD.n15838 DVDD.n3393 4.5005
R8730 DVDD.n15838 DVDD.n3400 4.5005
R8731 DVDD.n15838 DVDD.n3392 4.5005
R8732 DVDD.n15838 DVDD.n3401 4.5005
R8733 DVDD.n15838 DVDD.n3391 4.5005
R8734 DVDD.n15838 DVDD.n3402 4.5005
R8735 DVDD.n15838 DVDD.n3390 4.5005
R8736 DVDD.n15838 DVDD.n3404 4.5005
R8737 DVDD.n15838 DVDD.n3389 4.5005
R8738 DVDD.n15838 DVDD.n15837 4.5005
R8739 DVDD.n15838 DVDD.n3381 4.5005
R8740 DVDD.n15839 DVDD.n15838 4.5005
R8741 DVDD.n3080 DVDD.n3073 4.5005
R8742 DVDD.n3082 DVDD.n3073 4.5005
R8743 DVDD.n3079 DVDD.n3073 4.5005
R8744 DVDD.n3083 DVDD.n3073 4.5005
R8745 DVDD.n3078 DVDD.n3073 4.5005
R8746 DVDD.n3084 DVDD.n3073 4.5005
R8747 DVDD.n3077 DVDD.n3073 4.5005
R8748 DVDD.n3085 DVDD.n3073 4.5005
R8749 DVDD.n3076 DVDD.n3073 4.5005
R8750 DVDD.n3086 DVDD.n3073 4.5005
R8751 DVDD.n3075 DVDD.n3073 4.5005
R8752 DVDD.n16083 DVDD.n3073 4.5005
R8753 DVDD.n3073 DVDD.n3057 4.5005
R8754 DVDD.n16085 DVDD.n3073 4.5005
R8755 DVDD.n3073 DVDD.n3053 4.5005
R8756 DVDD.n3080 DVDD.n3058 4.5005
R8757 DVDD.n3082 DVDD.n3058 4.5005
R8758 DVDD.n3079 DVDD.n3058 4.5005
R8759 DVDD.n3083 DVDD.n3058 4.5005
R8760 DVDD.n3078 DVDD.n3058 4.5005
R8761 DVDD.n3084 DVDD.n3058 4.5005
R8762 DVDD.n3077 DVDD.n3058 4.5005
R8763 DVDD.n3085 DVDD.n3058 4.5005
R8764 DVDD.n3076 DVDD.n3058 4.5005
R8765 DVDD.n3086 DVDD.n3058 4.5005
R8766 DVDD.n3075 DVDD.n3058 4.5005
R8767 DVDD.n16083 DVDD.n3058 4.5005
R8768 DVDD.n3058 DVDD.n3057 4.5005
R8769 DVDD.n16085 DVDD.n3058 4.5005
R8770 DVDD.n3058 DVDD.n3053 4.5005
R8771 DVDD.n16084 DVDD.n3080 4.5005
R8772 DVDD.n16084 DVDD.n3082 4.5005
R8773 DVDD.n16084 DVDD.n3079 4.5005
R8774 DVDD.n16084 DVDD.n3083 4.5005
R8775 DVDD.n16084 DVDD.n3078 4.5005
R8776 DVDD.n16084 DVDD.n3084 4.5005
R8777 DVDD.n16084 DVDD.n3077 4.5005
R8778 DVDD.n16084 DVDD.n3085 4.5005
R8779 DVDD.n16084 DVDD.n3076 4.5005
R8780 DVDD.n16084 DVDD.n3086 4.5005
R8781 DVDD.n16084 DVDD.n3075 4.5005
R8782 DVDD.n16084 DVDD.n16083 4.5005
R8783 DVDD.n16084 DVDD.n3057 4.5005
R8784 DVDD.n16085 DVDD.n16084 4.5005
R8785 DVDD.n16084 DVDD.n3053 4.5005
R8786 DVDD.n9639 DVDD.n9620 4.5005
R8787 DVDD.n9639 DVDD.n9621 4.5005
R8788 DVDD.n9639 DVDD.n9619 4.5005
R8789 DVDD.n9642 DVDD.n9639 4.5005
R8790 DVDD.n9641 DVDD.n9639 4.5005
R8791 DVDD.n9639 DVDD.n9622 4.5005
R8792 DVDD.n9639 DVDD.n9617 4.5005
R8793 DVDD.n9639 DVDD.n9623 4.5005
R8794 DVDD.n9639 DVDD.n9616 4.5005
R8795 DVDD.n9639 DVDD.n9624 4.5005
R8796 DVDD.n9639 DVDD.n9615 4.5005
R8797 DVDD.n10091 DVDD.n9639 4.5005
R8798 DVDD.n9648 DVDD.n9639 4.5005
R8799 DVDD.n9639 DVDD.n9625 4.5005
R8800 DVDD.n10093 DVDD.n9639 4.5005
R8801 DVDD.n9627 DVDD.n9620 4.5005
R8802 DVDD.n9627 DVDD.n9621 4.5005
R8803 DVDD.n9627 DVDD.n9619 4.5005
R8804 DVDD.n9642 DVDD.n9627 4.5005
R8805 DVDD.n9641 DVDD.n9627 4.5005
R8806 DVDD.n9627 DVDD.n9622 4.5005
R8807 DVDD.n9627 DVDD.n9617 4.5005
R8808 DVDD.n9627 DVDD.n9623 4.5005
R8809 DVDD.n9627 DVDD.n9616 4.5005
R8810 DVDD.n9627 DVDD.n9624 4.5005
R8811 DVDD.n9627 DVDD.n9615 4.5005
R8812 DVDD.n10091 DVDD.n9627 4.5005
R8813 DVDD.n9627 DVDD.n9625 4.5005
R8814 DVDD.n9627 DVDD.n9613 4.5005
R8815 DVDD.n10093 DVDD.n9627 4.5005
R8816 DVDD.n10092 DVDD.n9620 4.5005
R8817 DVDD.n10092 DVDD.n9621 4.5005
R8818 DVDD.n10092 DVDD.n9619 4.5005
R8819 DVDD.n10092 DVDD.n9642 4.5005
R8820 DVDD.n10092 DVDD.n9641 4.5005
R8821 DVDD.n10092 DVDD.n9622 4.5005
R8822 DVDD.n10092 DVDD.n9617 4.5005
R8823 DVDD.n10092 DVDD.n9623 4.5005
R8824 DVDD.n10092 DVDD.n9616 4.5005
R8825 DVDD.n10092 DVDD.n9624 4.5005
R8826 DVDD.n10092 DVDD.n9615 4.5005
R8827 DVDD.n10092 DVDD.n10091 4.5005
R8828 DVDD.n10092 DVDD.n9625 4.5005
R8829 DVDD.n10092 DVDD.n9613 4.5005
R8830 DVDD.n10093 DVDD.n10092 4.5005
R8831 DVDD.n4978 DVDD.n3396 4.5005
R8832 DVDD.n16397 DVDD.n16396 4.5005
R8833 DVDD.n2475 DVDD.n2474 4.5005
R8834 DVDD.n3370 DVDD.n2293 4.5005
R8835 DVDD.n16399 DVDD.n2294 4.5005
R8836 DVDD.n2413 DVDD.n2324 4.5005
R8837 DVDD.n4978 DVDD.n4977 4.5005
R8838 DVDD.n4977 DVDD.n4952 4.5005
R8839 DVDD.n4977 DVDD.n4955 4.5005
R8840 DVDD.n4977 DVDD.n4951 4.5005
R8841 DVDD.n4977 DVDD.n4958 4.5005
R8842 DVDD.n4977 DVDD.n4950 4.5005
R8843 DVDD.n4977 DVDD.n4961 4.5005
R8844 DVDD.n4977 DVDD.n4949 4.5005
R8845 DVDD.n4977 DVDD.n4964 4.5005
R8846 DVDD.n4977 DVDD.n4948 4.5005
R8847 DVDD.n4977 DVDD.n4967 4.5005
R8848 DVDD.n4977 DVDD.n4947 4.5005
R8849 DVDD.n4977 DVDD.n4970 4.5005
R8850 DVDD.n4977 DVDD.n4946 4.5005
R8851 DVDD.n4977 DVDD.n4973 4.5005
R8852 DVDD.n4977 DVDD.n4945 4.5005
R8853 DVDD.n4977 DVDD.n4976 4.5005
R8854 DVDD.n4977 DVDD.n4944 4.5005
R8855 DVDD.n4977 DVDD.n2293 4.5005
R8856 DVDD.n16399 DVDD.n16398 4.5005
R8857 DVDD.n16398 DVDD.n2305 4.5005
R8858 DVDD.n16398 DVDD.n2308 4.5005
R8859 DVDD.n16398 DVDD.n2304 4.5005
R8860 DVDD.n16398 DVDD.n2310 4.5005
R8861 DVDD.n16398 DVDD.n2303 4.5005
R8862 DVDD.n16398 DVDD.n2312 4.5005
R8863 DVDD.n16398 DVDD.n2302 4.5005
R8864 DVDD.n16398 DVDD.n2314 4.5005
R8865 DVDD.n16398 DVDD.n2301 4.5005
R8866 DVDD.n16398 DVDD.n2316 4.5005
R8867 DVDD.n16398 DVDD.n2300 4.5005
R8868 DVDD.n16398 DVDD.n2318 4.5005
R8869 DVDD.n16398 DVDD.n2299 4.5005
R8870 DVDD.n16398 DVDD.n2320 4.5005
R8871 DVDD.n16398 DVDD.n2298 4.5005
R8872 DVDD.n16398 DVDD.n2322 4.5005
R8873 DVDD.n16398 DVDD.n2297 4.5005
R8874 DVDD.n16398 DVDD.n16397 4.5005
R8875 DVDD.n2473 DVDD.n2324 4.5005
R8876 DVDD.n2473 DVDD.n2456 4.5005
R8877 DVDD.n2473 DVDD.n2458 4.5005
R8878 DVDD.n2473 DVDD.n2455 4.5005
R8879 DVDD.n2473 DVDD.n2460 4.5005
R8880 DVDD.n2473 DVDD.n2454 4.5005
R8881 DVDD.n2473 DVDD.n2462 4.5005
R8882 DVDD.n2473 DVDD.n2453 4.5005
R8883 DVDD.n2473 DVDD.n2464 4.5005
R8884 DVDD.n2473 DVDD.n2452 4.5005
R8885 DVDD.n2473 DVDD.n2466 4.5005
R8886 DVDD.n2473 DVDD.n2451 4.5005
R8887 DVDD.n2473 DVDD.n2468 4.5005
R8888 DVDD.n2473 DVDD.n2450 4.5005
R8889 DVDD.n2473 DVDD.n2470 4.5005
R8890 DVDD.n2473 DVDD.n2449 4.5005
R8891 DVDD.n2473 DVDD.n2472 4.5005
R8892 DVDD.n2473 DVDD.n2448 4.5005
R8893 DVDD.n2474 DVDD.n2473 4.5005
R8894 DVDD.n4996 DVDD.n4995 4.5005
R8895 DVDD.n4996 DVDD.n4906 4.5005
R8896 DVDD.n4996 DVDD.n4985 4.5005
R8897 DVDD.n5002 DVDD.n4982 4.5005
R8898 DVDD.n4995 DVDD.n4992 4.5005
R8899 DVDD.n4987 DVDD.n4985 4.5005
R8900 DVDD.n5000 DVDD.n4989 4.5005
R8901 DVDD.n5000 DVDD.n4990 4.5005
R8902 DVDD.n5000 DVDD.n4988 4.5005
R8903 DVDD.n5000 DVDD.n4999 4.5005
R8904 DVDD.n5000 DVDD.n4982 4.5005
R8905 DVDD.n5001 DVDD.n5000 4.5005
R8906 DVDD.n5002 DVDD.n5001 4.5005
R8907 DVDD.n3978 DVDD.n3916 4.5005
R8908 DVDD.n3916 DVDD.n3910 4.5005
R8909 DVDD.n3927 DVDD.n3916 4.5005
R8910 DVDD.n3925 DVDD.n3916 4.5005
R8911 DVDD.n3930 DVDD.n3916 4.5005
R8912 DVDD.n3923 DVDD.n3916 4.5005
R8913 DVDD.n3931 DVDD.n3916 4.5005
R8914 DVDD.n3922 DVDD.n3916 4.5005
R8915 DVDD.n3932 DVDD.n3916 4.5005
R8916 DVDD.n3971 DVDD.n3916 4.5005
R8917 DVDD.n3965 DVDD.n3916 4.5005
R8918 DVDD.n3976 DVDD.n3916 4.5005
R8919 DVDD.n3978 DVDD.n3915 4.5005
R8920 DVDD.n3915 DVDD.n3910 4.5005
R8921 DVDD.n3927 DVDD.n3915 4.5005
R8922 DVDD.n3925 DVDD.n3915 4.5005
R8923 DVDD.n3929 DVDD.n3915 4.5005
R8924 DVDD.n3924 DVDD.n3915 4.5005
R8925 DVDD.n3930 DVDD.n3915 4.5005
R8926 DVDD.n3923 DVDD.n3915 4.5005
R8927 DVDD.n3931 DVDD.n3915 4.5005
R8928 DVDD.n3922 DVDD.n3915 4.5005
R8929 DVDD.n3932 DVDD.n3915 4.5005
R8930 DVDD.n3965 DVDD.n3915 4.5005
R8931 DVDD.n3976 DVDD.n3915 4.5005
R8932 DVDD.n3978 DVDD.n3917 4.5005
R8933 DVDD.n3917 DVDD.n3910 4.5005
R8934 DVDD.n3927 DVDD.n3917 4.5005
R8935 DVDD.n3925 DVDD.n3917 4.5005
R8936 DVDD.n3929 DVDD.n3917 4.5005
R8937 DVDD.n3924 DVDD.n3917 4.5005
R8938 DVDD.n3930 DVDD.n3917 4.5005
R8939 DVDD.n3923 DVDD.n3917 4.5005
R8940 DVDD.n3931 DVDD.n3917 4.5005
R8941 DVDD.n3922 DVDD.n3917 4.5005
R8942 DVDD.n3932 DVDD.n3917 4.5005
R8943 DVDD.n3965 DVDD.n3917 4.5005
R8944 DVDD.n3976 DVDD.n3917 4.5005
R8945 DVDD.n3978 DVDD.n3914 4.5005
R8946 DVDD.n3914 DVDD.n3910 4.5005
R8947 DVDD.n3927 DVDD.n3914 4.5005
R8948 DVDD.n3925 DVDD.n3914 4.5005
R8949 DVDD.n3929 DVDD.n3914 4.5005
R8950 DVDD.n3924 DVDD.n3914 4.5005
R8951 DVDD.n3930 DVDD.n3914 4.5005
R8952 DVDD.n3923 DVDD.n3914 4.5005
R8953 DVDD.n3931 DVDD.n3914 4.5005
R8954 DVDD.n3922 DVDD.n3914 4.5005
R8955 DVDD.n3932 DVDD.n3914 4.5005
R8956 DVDD.n3965 DVDD.n3914 4.5005
R8957 DVDD.n3976 DVDD.n3914 4.5005
R8958 DVDD.n3978 DVDD.n3918 4.5005
R8959 DVDD.n3918 DVDD.n3910 4.5005
R8960 DVDD.n3927 DVDD.n3918 4.5005
R8961 DVDD.n3925 DVDD.n3918 4.5005
R8962 DVDD.n3929 DVDD.n3918 4.5005
R8963 DVDD.n3924 DVDD.n3918 4.5005
R8964 DVDD.n3930 DVDD.n3918 4.5005
R8965 DVDD.n3923 DVDD.n3918 4.5005
R8966 DVDD.n3931 DVDD.n3918 4.5005
R8967 DVDD.n3922 DVDD.n3918 4.5005
R8968 DVDD.n3932 DVDD.n3918 4.5005
R8969 DVDD.n3965 DVDD.n3918 4.5005
R8970 DVDD.n3976 DVDD.n3918 4.5005
R8971 DVDD.n3978 DVDD.n3913 4.5005
R8972 DVDD.n3913 DVDD.n3910 4.5005
R8973 DVDD.n3927 DVDD.n3913 4.5005
R8974 DVDD.n3925 DVDD.n3913 4.5005
R8975 DVDD.n3929 DVDD.n3913 4.5005
R8976 DVDD.n3924 DVDD.n3913 4.5005
R8977 DVDD.n3930 DVDD.n3913 4.5005
R8978 DVDD.n3923 DVDD.n3913 4.5005
R8979 DVDD.n3931 DVDD.n3913 4.5005
R8980 DVDD.n3922 DVDD.n3913 4.5005
R8981 DVDD.n3932 DVDD.n3913 4.5005
R8982 DVDD.n3965 DVDD.n3913 4.5005
R8983 DVDD.n3976 DVDD.n3913 4.5005
R8984 DVDD.n3978 DVDD.n3919 4.5005
R8985 DVDD.n3919 DVDD.n3910 4.5005
R8986 DVDD.n3927 DVDD.n3919 4.5005
R8987 DVDD.n3925 DVDD.n3919 4.5005
R8988 DVDD.n3929 DVDD.n3919 4.5005
R8989 DVDD.n3924 DVDD.n3919 4.5005
R8990 DVDD.n3930 DVDD.n3919 4.5005
R8991 DVDD.n3923 DVDD.n3919 4.5005
R8992 DVDD.n3931 DVDD.n3919 4.5005
R8993 DVDD.n3922 DVDD.n3919 4.5005
R8994 DVDD.n3932 DVDD.n3919 4.5005
R8995 DVDD.n3965 DVDD.n3919 4.5005
R8996 DVDD.n3976 DVDD.n3919 4.5005
R8997 DVDD.n3978 DVDD.n3912 4.5005
R8998 DVDD.n3912 DVDD.n3910 4.5005
R8999 DVDD.n3927 DVDD.n3912 4.5005
R9000 DVDD.n3925 DVDD.n3912 4.5005
R9001 DVDD.n3929 DVDD.n3912 4.5005
R9002 DVDD.n3924 DVDD.n3912 4.5005
R9003 DVDD.n3930 DVDD.n3912 4.5005
R9004 DVDD.n3923 DVDD.n3912 4.5005
R9005 DVDD.n3931 DVDD.n3912 4.5005
R9006 DVDD.n3922 DVDD.n3912 4.5005
R9007 DVDD.n3932 DVDD.n3912 4.5005
R9008 DVDD.n3965 DVDD.n3912 4.5005
R9009 DVDD.n3976 DVDD.n3912 4.5005
R9010 DVDD.n3978 DVDD.n3920 4.5005
R9011 DVDD.n3920 DVDD.n3910 4.5005
R9012 DVDD.n3927 DVDD.n3920 4.5005
R9013 DVDD.n3925 DVDD.n3920 4.5005
R9014 DVDD.n3929 DVDD.n3920 4.5005
R9015 DVDD.n3924 DVDD.n3920 4.5005
R9016 DVDD.n3930 DVDD.n3920 4.5005
R9017 DVDD.n3923 DVDD.n3920 4.5005
R9018 DVDD.n3931 DVDD.n3920 4.5005
R9019 DVDD.n3922 DVDD.n3920 4.5005
R9020 DVDD.n3932 DVDD.n3920 4.5005
R9021 DVDD.n3965 DVDD.n3920 4.5005
R9022 DVDD.n3976 DVDD.n3920 4.5005
R9023 DVDD.n3978 DVDD.n3911 4.5005
R9024 DVDD.n3911 DVDD.n3910 4.5005
R9025 DVDD.n3927 DVDD.n3911 4.5005
R9026 DVDD.n3925 DVDD.n3911 4.5005
R9027 DVDD.n3929 DVDD.n3911 4.5005
R9028 DVDD.n3924 DVDD.n3911 4.5005
R9029 DVDD.n3930 DVDD.n3911 4.5005
R9030 DVDD.n3923 DVDD.n3911 4.5005
R9031 DVDD.n3931 DVDD.n3911 4.5005
R9032 DVDD.n3922 DVDD.n3911 4.5005
R9033 DVDD.n3932 DVDD.n3911 4.5005
R9034 DVDD.n3965 DVDD.n3911 4.5005
R9035 DVDD.n3976 DVDD.n3911 4.5005
R9036 DVDD.n3978 DVDD.n3977 4.5005
R9037 DVDD.n3977 DVDD.n3910 4.5005
R9038 DVDD.n3977 DVDD.n3927 4.5005
R9039 DVDD.n3977 DVDD.n3925 4.5005
R9040 DVDD.n3977 DVDD.n3929 4.5005
R9041 DVDD.n3977 DVDD.n3924 4.5005
R9042 DVDD.n3977 DVDD.n3930 4.5005
R9043 DVDD.n3977 DVDD.n3923 4.5005
R9044 DVDD.n3977 DVDD.n3931 4.5005
R9045 DVDD.n3977 DVDD.n3922 4.5005
R9046 DVDD.n3977 DVDD.n3932 4.5005
R9047 DVDD.n3977 DVDD.n3976 4.5005
R9048 DVDD.n3578 DVDD.n3558 4.5005
R9049 DVDD.n3578 DVDD.n3557 4.5005
R9050 DVDD.n3578 DVDD.n3559 4.5005
R9051 DVDD.n3578 DVDD.n3556 4.5005
R9052 DVDD.n3578 DVDD.n3561 4.5005
R9053 DVDD.n3578 DVDD.n3554 4.5005
R9054 DVDD.n3578 DVDD.n3562 4.5005
R9055 DVDD.n3578 DVDD.n3553 4.5005
R9056 DVDD.n3578 DVDD.n3563 4.5005
R9057 DVDD.n3578 DVDD.n3552 4.5005
R9058 DVDD.n3578 DVDD.n3564 4.5005
R9059 DVDD.n4838 DVDD.n3578 4.5005
R9060 DVDD.n4805 DVDD.n3558 4.5005
R9061 DVDD.n4805 DVDD.n3557 4.5005
R9062 DVDD.n4805 DVDD.n3559 4.5005
R9063 DVDD.n4805 DVDD.n3556 4.5005
R9064 DVDD.n4805 DVDD.n3560 4.5005
R9065 DVDD.n4805 DVDD.n3555 4.5005
R9066 DVDD.n4805 DVDD.n3561 4.5005
R9067 DVDD.n4805 DVDD.n3554 4.5005
R9068 DVDD.n4805 DVDD.n3562 4.5005
R9069 DVDD.n4805 DVDD.n3553 4.5005
R9070 DVDD.n4805 DVDD.n3563 4.5005
R9071 DVDD.n4805 DVDD.n3564 4.5005
R9072 DVDD.n4838 DVDD.n4805 4.5005
R9073 DVDD.n3576 DVDD.n3558 4.5005
R9074 DVDD.n3576 DVDD.n3557 4.5005
R9075 DVDD.n3576 DVDD.n3559 4.5005
R9076 DVDD.n3576 DVDD.n3556 4.5005
R9077 DVDD.n3576 DVDD.n3560 4.5005
R9078 DVDD.n3576 DVDD.n3555 4.5005
R9079 DVDD.n3576 DVDD.n3561 4.5005
R9080 DVDD.n3576 DVDD.n3554 4.5005
R9081 DVDD.n3576 DVDD.n3562 4.5005
R9082 DVDD.n3576 DVDD.n3553 4.5005
R9083 DVDD.n3576 DVDD.n3563 4.5005
R9084 DVDD.n3576 DVDD.n3564 4.5005
R9085 DVDD.n4838 DVDD.n3576 4.5005
R9086 DVDD.n4807 DVDD.n3558 4.5005
R9087 DVDD.n4807 DVDD.n3557 4.5005
R9088 DVDD.n4807 DVDD.n3559 4.5005
R9089 DVDD.n4807 DVDD.n3556 4.5005
R9090 DVDD.n4807 DVDD.n3560 4.5005
R9091 DVDD.n4807 DVDD.n3555 4.5005
R9092 DVDD.n4807 DVDD.n3561 4.5005
R9093 DVDD.n4807 DVDD.n3554 4.5005
R9094 DVDD.n4807 DVDD.n3562 4.5005
R9095 DVDD.n4807 DVDD.n3553 4.5005
R9096 DVDD.n4807 DVDD.n3563 4.5005
R9097 DVDD.n4807 DVDD.n3564 4.5005
R9098 DVDD.n4838 DVDD.n4807 4.5005
R9099 DVDD.n3575 DVDD.n3558 4.5005
R9100 DVDD.n3575 DVDD.n3557 4.5005
R9101 DVDD.n3575 DVDD.n3559 4.5005
R9102 DVDD.n3575 DVDD.n3556 4.5005
R9103 DVDD.n3575 DVDD.n3560 4.5005
R9104 DVDD.n3575 DVDD.n3555 4.5005
R9105 DVDD.n3575 DVDD.n3561 4.5005
R9106 DVDD.n3575 DVDD.n3554 4.5005
R9107 DVDD.n3575 DVDD.n3562 4.5005
R9108 DVDD.n3575 DVDD.n3553 4.5005
R9109 DVDD.n3575 DVDD.n3563 4.5005
R9110 DVDD.n3575 DVDD.n3564 4.5005
R9111 DVDD.n4838 DVDD.n3575 4.5005
R9112 DVDD.n4809 DVDD.n3558 4.5005
R9113 DVDD.n4809 DVDD.n3557 4.5005
R9114 DVDD.n4809 DVDD.n3559 4.5005
R9115 DVDD.n4809 DVDD.n3556 4.5005
R9116 DVDD.n4809 DVDD.n3560 4.5005
R9117 DVDD.n4809 DVDD.n3555 4.5005
R9118 DVDD.n4809 DVDD.n3561 4.5005
R9119 DVDD.n4809 DVDD.n3554 4.5005
R9120 DVDD.n4809 DVDD.n3562 4.5005
R9121 DVDD.n4809 DVDD.n3553 4.5005
R9122 DVDD.n4809 DVDD.n3563 4.5005
R9123 DVDD.n4809 DVDD.n3564 4.5005
R9124 DVDD.n4838 DVDD.n4809 4.5005
R9125 DVDD.n3574 DVDD.n3558 4.5005
R9126 DVDD.n3574 DVDD.n3557 4.5005
R9127 DVDD.n3574 DVDD.n3559 4.5005
R9128 DVDD.n3574 DVDD.n3556 4.5005
R9129 DVDD.n3574 DVDD.n3560 4.5005
R9130 DVDD.n3574 DVDD.n3555 4.5005
R9131 DVDD.n3574 DVDD.n3561 4.5005
R9132 DVDD.n3574 DVDD.n3554 4.5005
R9133 DVDD.n3574 DVDD.n3562 4.5005
R9134 DVDD.n3574 DVDD.n3553 4.5005
R9135 DVDD.n3574 DVDD.n3563 4.5005
R9136 DVDD.n3574 DVDD.n3564 4.5005
R9137 DVDD.n4838 DVDD.n3574 4.5005
R9138 DVDD.n4811 DVDD.n3558 4.5005
R9139 DVDD.n4811 DVDD.n3557 4.5005
R9140 DVDD.n4811 DVDD.n3559 4.5005
R9141 DVDD.n4811 DVDD.n3556 4.5005
R9142 DVDD.n4811 DVDD.n3560 4.5005
R9143 DVDD.n4811 DVDD.n3555 4.5005
R9144 DVDD.n4811 DVDD.n3561 4.5005
R9145 DVDD.n4811 DVDD.n3554 4.5005
R9146 DVDD.n4811 DVDD.n3562 4.5005
R9147 DVDD.n4811 DVDD.n3553 4.5005
R9148 DVDD.n4811 DVDD.n3563 4.5005
R9149 DVDD.n4811 DVDD.n3564 4.5005
R9150 DVDD.n4838 DVDD.n4811 4.5005
R9151 DVDD.n3573 DVDD.n3558 4.5005
R9152 DVDD.n3573 DVDD.n3557 4.5005
R9153 DVDD.n3573 DVDD.n3559 4.5005
R9154 DVDD.n3573 DVDD.n3556 4.5005
R9155 DVDD.n3573 DVDD.n3560 4.5005
R9156 DVDD.n3573 DVDD.n3555 4.5005
R9157 DVDD.n3573 DVDD.n3561 4.5005
R9158 DVDD.n3573 DVDD.n3554 4.5005
R9159 DVDD.n3573 DVDD.n3562 4.5005
R9160 DVDD.n3573 DVDD.n3553 4.5005
R9161 DVDD.n3573 DVDD.n3563 4.5005
R9162 DVDD.n3573 DVDD.n3564 4.5005
R9163 DVDD.n4838 DVDD.n3573 4.5005
R9164 DVDD.n4813 DVDD.n3558 4.5005
R9165 DVDD.n4813 DVDD.n3557 4.5005
R9166 DVDD.n4813 DVDD.n3559 4.5005
R9167 DVDD.n4813 DVDD.n3556 4.5005
R9168 DVDD.n4813 DVDD.n3560 4.5005
R9169 DVDD.n4813 DVDD.n3555 4.5005
R9170 DVDD.n4813 DVDD.n3561 4.5005
R9171 DVDD.n4813 DVDD.n3554 4.5005
R9172 DVDD.n4813 DVDD.n3562 4.5005
R9173 DVDD.n4813 DVDD.n3553 4.5005
R9174 DVDD.n4813 DVDD.n3563 4.5005
R9175 DVDD.n4813 DVDD.n3564 4.5005
R9176 DVDD.n4838 DVDD.n4813 4.5005
R9177 DVDD.n3572 DVDD.n3558 4.5005
R9178 DVDD.n3572 DVDD.n3557 4.5005
R9179 DVDD.n3572 DVDD.n3559 4.5005
R9180 DVDD.n3572 DVDD.n3556 4.5005
R9181 DVDD.n3572 DVDD.n3560 4.5005
R9182 DVDD.n3572 DVDD.n3555 4.5005
R9183 DVDD.n3572 DVDD.n3561 4.5005
R9184 DVDD.n3572 DVDD.n3554 4.5005
R9185 DVDD.n3572 DVDD.n3562 4.5005
R9186 DVDD.n3572 DVDD.n3553 4.5005
R9187 DVDD.n3572 DVDD.n3563 4.5005
R9188 DVDD.n3572 DVDD.n3564 4.5005
R9189 DVDD.n4838 DVDD.n3572 4.5005
R9190 DVDD.n4815 DVDD.n3558 4.5005
R9191 DVDD.n4815 DVDD.n3557 4.5005
R9192 DVDD.n4815 DVDD.n3559 4.5005
R9193 DVDD.n4815 DVDD.n3556 4.5005
R9194 DVDD.n4815 DVDD.n3560 4.5005
R9195 DVDD.n4815 DVDD.n3555 4.5005
R9196 DVDD.n4815 DVDD.n3561 4.5005
R9197 DVDD.n4815 DVDD.n3554 4.5005
R9198 DVDD.n4815 DVDD.n3562 4.5005
R9199 DVDD.n4815 DVDD.n3553 4.5005
R9200 DVDD.n4815 DVDD.n3563 4.5005
R9201 DVDD.n4815 DVDD.n3564 4.5005
R9202 DVDD.n4838 DVDD.n4815 4.5005
R9203 DVDD.n3571 DVDD.n3558 4.5005
R9204 DVDD.n3571 DVDD.n3557 4.5005
R9205 DVDD.n3571 DVDD.n3559 4.5005
R9206 DVDD.n3571 DVDD.n3556 4.5005
R9207 DVDD.n3571 DVDD.n3560 4.5005
R9208 DVDD.n3571 DVDD.n3555 4.5005
R9209 DVDD.n3571 DVDD.n3561 4.5005
R9210 DVDD.n3571 DVDD.n3554 4.5005
R9211 DVDD.n3571 DVDD.n3562 4.5005
R9212 DVDD.n3571 DVDD.n3553 4.5005
R9213 DVDD.n3571 DVDD.n3563 4.5005
R9214 DVDD.n3571 DVDD.n3564 4.5005
R9215 DVDD.n4838 DVDD.n3571 4.5005
R9216 DVDD.n4817 DVDD.n3558 4.5005
R9217 DVDD.n4817 DVDD.n3557 4.5005
R9218 DVDD.n4817 DVDD.n3559 4.5005
R9219 DVDD.n4817 DVDD.n3556 4.5005
R9220 DVDD.n4817 DVDD.n3560 4.5005
R9221 DVDD.n4817 DVDD.n3555 4.5005
R9222 DVDD.n4817 DVDD.n3561 4.5005
R9223 DVDD.n4817 DVDD.n3554 4.5005
R9224 DVDD.n4817 DVDD.n3562 4.5005
R9225 DVDD.n4817 DVDD.n3553 4.5005
R9226 DVDD.n4817 DVDD.n3563 4.5005
R9227 DVDD.n4817 DVDD.n3564 4.5005
R9228 DVDD.n4838 DVDD.n4817 4.5005
R9229 DVDD.n3570 DVDD.n3558 4.5005
R9230 DVDD.n3570 DVDD.n3557 4.5005
R9231 DVDD.n3570 DVDD.n3559 4.5005
R9232 DVDD.n3570 DVDD.n3556 4.5005
R9233 DVDD.n3570 DVDD.n3560 4.5005
R9234 DVDD.n3570 DVDD.n3555 4.5005
R9235 DVDD.n3570 DVDD.n3561 4.5005
R9236 DVDD.n3570 DVDD.n3554 4.5005
R9237 DVDD.n3570 DVDD.n3562 4.5005
R9238 DVDD.n3570 DVDD.n3553 4.5005
R9239 DVDD.n3570 DVDD.n3563 4.5005
R9240 DVDD.n3570 DVDD.n3564 4.5005
R9241 DVDD.n4838 DVDD.n3570 4.5005
R9242 DVDD.n4819 DVDD.n3558 4.5005
R9243 DVDD.n4819 DVDD.n3557 4.5005
R9244 DVDD.n4819 DVDD.n3559 4.5005
R9245 DVDD.n4819 DVDD.n3556 4.5005
R9246 DVDD.n4819 DVDD.n3560 4.5005
R9247 DVDD.n4819 DVDD.n3555 4.5005
R9248 DVDD.n4819 DVDD.n3561 4.5005
R9249 DVDD.n4819 DVDD.n3554 4.5005
R9250 DVDD.n4819 DVDD.n3562 4.5005
R9251 DVDD.n4819 DVDD.n3553 4.5005
R9252 DVDD.n4819 DVDD.n3563 4.5005
R9253 DVDD.n4819 DVDD.n3564 4.5005
R9254 DVDD.n4838 DVDD.n4819 4.5005
R9255 DVDD.n3569 DVDD.n3558 4.5005
R9256 DVDD.n3569 DVDD.n3557 4.5005
R9257 DVDD.n3569 DVDD.n3559 4.5005
R9258 DVDD.n3569 DVDD.n3556 4.5005
R9259 DVDD.n3569 DVDD.n3560 4.5005
R9260 DVDD.n3569 DVDD.n3555 4.5005
R9261 DVDD.n3569 DVDD.n3561 4.5005
R9262 DVDD.n3569 DVDD.n3554 4.5005
R9263 DVDD.n3569 DVDD.n3562 4.5005
R9264 DVDD.n3569 DVDD.n3553 4.5005
R9265 DVDD.n3569 DVDD.n3563 4.5005
R9266 DVDD.n3569 DVDD.n3564 4.5005
R9267 DVDD.n4838 DVDD.n3569 4.5005
R9268 DVDD.n4821 DVDD.n3558 4.5005
R9269 DVDD.n4821 DVDD.n3557 4.5005
R9270 DVDD.n4821 DVDD.n3559 4.5005
R9271 DVDD.n4821 DVDD.n3556 4.5005
R9272 DVDD.n4821 DVDD.n3560 4.5005
R9273 DVDD.n4821 DVDD.n3555 4.5005
R9274 DVDD.n4821 DVDD.n3561 4.5005
R9275 DVDD.n4821 DVDD.n3554 4.5005
R9276 DVDD.n4821 DVDD.n3562 4.5005
R9277 DVDD.n4821 DVDD.n3553 4.5005
R9278 DVDD.n4821 DVDD.n3563 4.5005
R9279 DVDD.n4821 DVDD.n3564 4.5005
R9280 DVDD.n4838 DVDD.n4821 4.5005
R9281 DVDD.n3568 DVDD.n3558 4.5005
R9282 DVDD.n3568 DVDD.n3557 4.5005
R9283 DVDD.n3568 DVDD.n3559 4.5005
R9284 DVDD.n3568 DVDD.n3556 4.5005
R9285 DVDD.n3568 DVDD.n3560 4.5005
R9286 DVDD.n3568 DVDD.n3555 4.5005
R9287 DVDD.n3568 DVDD.n3561 4.5005
R9288 DVDD.n3568 DVDD.n3554 4.5005
R9289 DVDD.n3568 DVDD.n3562 4.5005
R9290 DVDD.n3568 DVDD.n3553 4.5005
R9291 DVDD.n3568 DVDD.n3563 4.5005
R9292 DVDD.n3568 DVDD.n3564 4.5005
R9293 DVDD.n4838 DVDD.n3568 4.5005
R9294 DVDD.n4823 DVDD.n3558 4.5005
R9295 DVDD.n4823 DVDD.n3557 4.5005
R9296 DVDD.n4823 DVDD.n3559 4.5005
R9297 DVDD.n4823 DVDD.n3556 4.5005
R9298 DVDD.n4823 DVDD.n3560 4.5005
R9299 DVDD.n4823 DVDD.n3555 4.5005
R9300 DVDD.n4823 DVDD.n3561 4.5005
R9301 DVDD.n4823 DVDD.n3554 4.5005
R9302 DVDD.n4823 DVDD.n3562 4.5005
R9303 DVDD.n4823 DVDD.n3553 4.5005
R9304 DVDD.n4823 DVDD.n3563 4.5005
R9305 DVDD.n4823 DVDD.n3564 4.5005
R9306 DVDD.n4838 DVDD.n4823 4.5005
R9307 DVDD.n3567 DVDD.n3558 4.5005
R9308 DVDD.n3567 DVDD.n3557 4.5005
R9309 DVDD.n3567 DVDD.n3559 4.5005
R9310 DVDD.n3567 DVDD.n3556 4.5005
R9311 DVDD.n3567 DVDD.n3560 4.5005
R9312 DVDD.n3567 DVDD.n3555 4.5005
R9313 DVDD.n3567 DVDD.n3561 4.5005
R9314 DVDD.n3567 DVDD.n3554 4.5005
R9315 DVDD.n3567 DVDD.n3562 4.5005
R9316 DVDD.n3567 DVDD.n3553 4.5005
R9317 DVDD.n3567 DVDD.n3563 4.5005
R9318 DVDD.n3567 DVDD.n3564 4.5005
R9319 DVDD.n4838 DVDD.n3567 4.5005
R9320 DVDD.n4837 DVDD.n3558 4.5005
R9321 DVDD.n4837 DVDD.n3557 4.5005
R9322 DVDD.n4837 DVDD.n3559 4.5005
R9323 DVDD.n4837 DVDD.n3556 4.5005
R9324 DVDD.n4837 DVDD.n3560 4.5005
R9325 DVDD.n4837 DVDD.n3555 4.5005
R9326 DVDD.n4837 DVDD.n3561 4.5005
R9327 DVDD.n4837 DVDD.n3554 4.5005
R9328 DVDD.n4837 DVDD.n3562 4.5005
R9329 DVDD.n4837 DVDD.n3553 4.5005
R9330 DVDD.n4837 DVDD.n3563 4.5005
R9331 DVDD.n4837 DVDD.n3564 4.5005
R9332 DVDD.n4838 DVDD.n4837 4.5005
R9333 DVDD.n3566 DVDD.n3558 4.5005
R9334 DVDD.n3566 DVDD.n3557 4.5005
R9335 DVDD.n3566 DVDD.n3559 4.5005
R9336 DVDD.n3566 DVDD.n3556 4.5005
R9337 DVDD.n3566 DVDD.n3560 4.5005
R9338 DVDD.n3566 DVDD.n3555 4.5005
R9339 DVDD.n3566 DVDD.n3561 4.5005
R9340 DVDD.n3566 DVDD.n3554 4.5005
R9341 DVDD.n3566 DVDD.n3562 4.5005
R9342 DVDD.n3566 DVDD.n3553 4.5005
R9343 DVDD.n3566 DVDD.n3563 4.5005
R9344 DVDD.n3566 DVDD.n3564 4.5005
R9345 DVDD.n4838 DVDD.n3566 4.5005
R9346 DVDD.n4839 DVDD.n3558 4.5005
R9347 DVDD.n4839 DVDD.n3557 4.5005
R9348 DVDD.n4839 DVDD.n3559 4.5005
R9349 DVDD.n4839 DVDD.n3556 4.5005
R9350 DVDD.n4839 DVDD.n3560 4.5005
R9351 DVDD.n4839 DVDD.n3555 4.5005
R9352 DVDD.n4839 DVDD.n3561 4.5005
R9353 DVDD.n4839 DVDD.n3554 4.5005
R9354 DVDD.n4839 DVDD.n3562 4.5005
R9355 DVDD.n4839 DVDD.n3553 4.5005
R9356 DVDD.n4839 DVDD.n3563 4.5005
R9357 DVDD.n4839 DVDD.n3552 4.5005
R9358 DVDD.n4839 DVDD.n3564 4.5005
R9359 DVDD.n4839 DVDD.n4838 4.5005
R9360 DVDD.n4845 DVDD.n3527 4.5005
R9361 DVDD.n4845 DVDD.n3526 4.5005
R9362 DVDD.n4845 DVDD.n3528 4.5005
R9363 DVDD.n4845 DVDD.n3525 4.5005
R9364 DVDD.n4845 DVDD.n3530 4.5005
R9365 DVDD.n4845 DVDD.n3538 4.5005
R9366 DVDD.n4845 DVDD.n3531 4.5005
R9367 DVDD.n4842 DVDD.n3527 4.5005
R9368 DVDD.n4842 DVDD.n3526 4.5005
R9369 DVDD.n4842 DVDD.n3528 4.5005
R9370 DVDD.n4842 DVDD.n3525 4.5005
R9371 DVDD.n4842 DVDD.n3529 4.5005
R9372 DVDD.n4842 DVDD.n3524 4.5005
R9373 DVDD.n4842 DVDD.n3530 4.5005
R9374 DVDD.n4842 DVDD.n3531 4.5005
R9375 DVDD.n4840 DVDD.n3527 4.5005
R9376 DVDD.n4840 DVDD.n3526 4.5005
R9377 DVDD.n4840 DVDD.n3528 4.5005
R9378 DVDD.n4840 DVDD.n3525 4.5005
R9379 DVDD.n4840 DVDD.n3529 4.5005
R9380 DVDD.n4840 DVDD.n3524 4.5005
R9381 DVDD.n4840 DVDD.n3530 4.5005
R9382 DVDD.n4840 DVDD.n3531 4.5005
R9383 DVDD.n4852 DVDD.n3527 4.5005
R9384 DVDD.n4852 DVDD.n3526 4.5005
R9385 DVDD.n4852 DVDD.n3528 4.5005
R9386 DVDD.n4852 DVDD.n3525 4.5005
R9387 DVDD.n4852 DVDD.n3529 4.5005
R9388 DVDD.n4852 DVDD.n3524 4.5005
R9389 DVDD.n4852 DVDD.n3530 4.5005
R9390 DVDD.n4852 DVDD.n3531 4.5005
R9391 DVDD.n4856 DVDD.n3527 4.5005
R9392 DVDD.n4856 DVDD.n3526 4.5005
R9393 DVDD.n4856 DVDD.n3528 4.5005
R9394 DVDD.n4856 DVDD.n3525 4.5005
R9395 DVDD.n4856 DVDD.n3529 4.5005
R9396 DVDD.n4856 DVDD.n3524 4.5005
R9397 DVDD.n4856 DVDD.n3530 4.5005
R9398 DVDD.n4856 DVDD.n3531 4.5005
R9399 DVDD.n4854 DVDD.n3527 4.5005
R9400 DVDD.n4854 DVDD.n3526 4.5005
R9401 DVDD.n4854 DVDD.n3528 4.5005
R9402 DVDD.n4854 DVDD.n3525 4.5005
R9403 DVDD.n4854 DVDD.n3529 4.5005
R9404 DVDD.n4854 DVDD.n3524 4.5005
R9405 DVDD.n4854 DVDD.n3530 4.5005
R9406 DVDD.n4854 DVDD.n3531 4.5005
R9407 DVDD.n4867 DVDD.n3527 4.5005
R9408 DVDD.n4867 DVDD.n3526 4.5005
R9409 DVDD.n4867 DVDD.n3528 4.5005
R9410 DVDD.n4867 DVDD.n3525 4.5005
R9411 DVDD.n4867 DVDD.n3529 4.5005
R9412 DVDD.n4867 DVDD.n3524 4.5005
R9413 DVDD.n4867 DVDD.n3530 4.5005
R9414 DVDD.n4867 DVDD.n3531 4.5005
R9415 DVDD.n4869 DVDD.n3527 4.5005
R9416 DVDD.n4869 DVDD.n3526 4.5005
R9417 DVDD.n4869 DVDD.n3528 4.5005
R9418 DVDD.n4869 DVDD.n3525 4.5005
R9419 DVDD.n4869 DVDD.n3529 4.5005
R9420 DVDD.n4869 DVDD.n3524 4.5005
R9421 DVDD.n4869 DVDD.n3530 4.5005
R9422 DVDD.n4869 DVDD.n3531 4.5005
R9423 DVDD.n4873 DVDD.n3527 4.5005
R9424 DVDD.n4873 DVDD.n3526 4.5005
R9425 DVDD.n4873 DVDD.n3528 4.5005
R9426 DVDD.n4873 DVDD.n3525 4.5005
R9427 DVDD.n4873 DVDD.n3529 4.5005
R9428 DVDD.n4873 DVDD.n3524 4.5005
R9429 DVDD.n4873 DVDD.n3530 4.5005
R9430 DVDD.n4873 DVDD.n3531 4.5005
R9431 DVDD.n4871 DVDD.n3527 4.5005
R9432 DVDD.n4871 DVDD.n3526 4.5005
R9433 DVDD.n4871 DVDD.n3528 4.5005
R9434 DVDD.n4871 DVDD.n3525 4.5005
R9435 DVDD.n4871 DVDD.n3529 4.5005
R9436 DVDD.n4871 DVDD.n3524 4.5005
R9437 DVDD.n4871 DVDD.n3530 4.5005
R9438 DVDD.n4871 DVDD.n3531 4.5005
R9439 DVDD.n4880 DVDD.n3527 4.5005
R9440 DVDD.n4880 DVDD.n3526 4.5005
R9441 DVDD.n4880 DVDD.n3528 4.5005
R9442 DVDD.n4880 DVDD.n3525 4.5005
R9443 DVDD.n4880 DVDD.n3529 4.5005
R9444 DVDD.n4880 DVDD.n3524 4.5005
R9445 DVDD.n4880 DVDD.n3530 4.5005
R9446 DVDD.n4880 DVDD.n3531 4.5005
R9447 DVDD.n4880 DVDD.n3523 4.5005
R9448 DVDD.n15752 DVDD.n4881 4.5005
R9449 DVDD.n4904 DVDD.n4881 4.5005
R9450 DVDD.n15707 DVDD.n4881 4.5005
R9451 DVDD.n4903 DVDD.n4881 4.5005
R9452 DVDD.n15710 DVDD.n4881 4.5005
R9453 DVDD.n4901 DVDD.n4881 4.5005
R9454 DVDD.n15711 DVDD.n4881 4.5005
R9455 DVDD.n4900 DVDD.n4881 4.5005
R9456 DVDD.n15712 DVDD.n4881 4.5005
R9457 DVDD.n4899 DVDD.n4881 4.5005
R9458 DVDD.n15714 DVDD.n4881 4.5005
R9459 DVDD.n15750 DVDD.n4881 4.5005
R9460 DVDD.n15752 DVDD.n4882 4.5005
R9461 DVDD.n4904 DVDD.n4882 4.5005
R9462 DVDD.n15707 DVDD.n4882 4.5005
R9463 DVDD.n4903 DVDD.n4882 4.5005
R9464 DVDD.n15709 DVDD.n4882 4.5005
R9465 DVDD.n4902 DVDD.n4882 4.5005
R9466 DVDD.n15710 DVDD.n4882 4.5005
R9467 DVDD.n4901 DVDD.n4882 4.5005
R9468 DVDD.n15711 DVDD.n4882 4.5005
R9469 DVDD.n4900 DVDD.n4882 4.5005
R9470 DVDD.n15712 DVDD.n4882 4.5005
R9471 DVDD.n15714 DVDD.n4882 4.5005
R9472 DVDD.n15750 DVDD.n4882 4.5005
R9473 DVDD.n15752 DVDD.n3521 4.5005
R9474 DVDD.n4904 DVDD.n3521 4.5005
R9475 DVDD.n15707 DVDD.n3521 4.5005
R9476 DVDD.n4903 DVDD.n3521 4.5005
R9477 DVDD.n15709 DVDD.n3521 4.5005
R9478 DVDD.n4902 DVDD.n3521 4.5005
R9479 DVDD.n15710 DVDD.n3521 4.5005
R9480 DVDD.n4901 DVDD.n3521 4.5005
R9481 DVDD.n15711 DVDD.n3521 4.5005
R9482 DVDD.n4900 DVDD.n3521 4.5005
R9483 DVDD.n15712 DVDD.n3521 4.5005
R9484 DVDD.n15714 DVDD.n3521 4.5005
R9485 DVDD.n15750 DVDD.n3521 4.5005
R9486 DVDD.n15752 DVDD.n4883 4.5005
R9487 DVDD.n4904 DVDD.n4883 4.5005
R9488 DVDD.n15707 DVDD.n4883 4.5005
R9489 DVDD.n4903 DVDD.n4883 4.5005
R9490 DVDD.n15709 DVDD.n4883 4.5005
R9491 DVDD.n4902 DVDD.n4883 4.5005
R9492 DVDD.n15710 DVDD.n4883 4.5005
R9493 DVDD.n4901 DVDD.n4883 4.5005
R9494 DVDD.n15711 DVDD.n4883 4.5005
R9495 DVDD.n4900 DVDD.n4883 4.5005
R9496 DVDD.n15712 DVDD.n4883 4.5005
R9497 DVDD.n15714 DVDD.n4883 4.5005
R9498 DVDD.n15750 DVDD.n4883 4.5005
R9499 DVDD.n15752 DVDD.n3520 4.5005
R9500 DVDD.n4904 DVDD.n3520 4.5005
R9501 DVDD.n15707 DVDD.n3520 4.5005
R9502 DVDD.n4903 DVDD.n3520 4.5005
R9503 DVDD.n15709 DVDD.n3520 4.5005
R9504 DVDD.n4902 DVDD.n3520 4.5005
R9505 DVDD.n15710 DVDD.n3520 4.5005
R9506 DVDD.n4901 DVDD.n3520 4.5005
R9507 DVDD.n15711 DVDD.n3520 4.5005
R9508 DVDD.n4900 DVDD.n3520 4.5005
R9509 DVDD.n15712 DVDD.n3520 4.5005
R9510 DVDD.n15750 DVDD.n3520 4.5005
R9511 DVDD.n15752 DVDD.n4884 4.5005
R9512 DVDD.n4904 DVDD.n4884 4.5005
R9513 DVDD.n15707 DVDD.n4884 4.5005
R9514 DVDD.n4903 DVDD.n4884 4.5005
R9515 DVDD.n15709 DVDD.n4884 4.5005
R9516 DVDD.n4902 DVDD.n4884 4.5005
R9517 DVDD.n15710 DVDD.n4884 4.5005
R9518 DVDD.n4901 DVDD.n4884 4.5005
R9519 DVDD.n15711 DVDD.n4884 4.5005
R9520 DVDD.n4900 DVDD.n4884 4.5005
R9521 DVDD.n15712 DVDD.n4884 4.5005
R9522 DVDD.n4899 DVDD.n4884 4.5005
R9523 DVDD.n15714 DVDD.n4884 4.5005
R9524 DVDD.n4896 DVDD.n4884 4.5005
R9525 DVDD.n15750 DVDD.n4884 4.5005
R9526 DVDD.n15711 DVDD.n3519 4.5005
R9527 DVDD.n4900 DVDD.n3519 4.5005
R9528 DVDD.n15712 DVDD.n3519 4.5005
R9529 DVDD.n4899 DVDD.n3519 4.5005
R9530 DVDD.n15714 DVDD.n3519 4.5005
R9531 DVDD.n4896 DVDD.n3519 4.5005
R9532 DVDD.n15750 DVDD.n3519 4.5005
R9533 DVDD.n4901 DVDD.n3519 4.5005
R9534 DVDD.n15710 DVDD.n3519 4.5005
R9535 DVDD.n4902 DVDD.n3519 4.5005
R9536 DVDD.n15709 DVDD.n3519 4.5005
R9537 DVDD.n4903 DVDD.n3519 4.5005
R9538 DVDD.n15707 DVDD.n3519 4.5005
R9539 DVDD.n4904 DVDD.n3519 4.5005
R9540 DVDD.n15752 DVDD.n3519 4.5005
R9541 DVDD.n15711 DVDD.n4885 4.5005
R9542 DVDD.n4900 DVDD.n4885 4.5005
R9543 DVDD.n15712 DVDD.n4885 4.5005
R9544 DVDD.n4899 DVDD.n4885 4.5005
R9545 DVDD.n15714 DVDD.n4885 4.5005
R9546 DVDD.n4896 DVDD.n4885 4.5005
R9547 DVDD.n15750 DVDD.n4885 4.5005
R9548 DVDD.n4901 DVDD.n4885 4.5005
R9549 DVDD.n15710 DVDD.n4885 4.5005
R9550 DVDD.n4902 DVDD.n4885 4.5005
R9551 DVDD.n15709 DVDD.n4885 4.5005
R9552 DVDD.n4903 DVDD.n4885 4.5005
R9553 DVDD.n15707 DVDD.n4885 4.5005
R9554 DVDD.n4904 DVDD.n4885 4.5005
R9555 DVDD.n15752 DVDD.n4885 4.5005
R9556 DVDD.n15711 DVDD.n3518 4.5005
R9557 DVDD.n4900 DVDD.n3518 4.5005
R9558 DVDD.n15712 DVDD.n3518 4.5005
R9559 DVDD.n4899 DVDD.n3518 4.5005
R9560 DVDD.n15714 DVDD.n3518 4.5005
R9561 DVDD.n4896 DVDD.n3518 4.5005
R9562 DVDD.n15750 DVDD.n3518 4.5005
R9563 DVDD.n4901 DVDD.n3518 4.5005
R9564 DVDD.n15710 DVDD.n3518 4.5005
R9565 DVDD.n4902 DVDD.n3518 4.5005
R9566 DVDD.n15709 DVDD.n3518 4.5005
R9567 DVDD.n4903 DVDD.n3518 4.5005
R9568 DVDD.n15707 DVDD.n3518 4.5005
R9569 DVDD.n4904 DVDD.n3518 4.5005
R9570 DVDD.n15752 DVDD.n3518 4.5005
R9571 DVDD.n15752 DVDD.n4886 4.5005
R9572 DVDD.n4904 DVDD.n4886 4.5005
R9573 DVDD.n15707 DVDD.n4886 4.5005
R9574 DVDD.n4903 DVDD.n4886 4.5005
R9575 DVDD.n15709 DVDD.n4886 4.5005
R9576 DVDD.n4902 DVDD.n4886 4.5005
R9577 DVDD.n15710 DVDD.n4886 4.5005
R9578 DVDD.n4901 DVDD.n4886 4.5005
R9579 DVDD.n15711 DVDD.n4886 4.5005
R9580 DVDD.n4900 DVDD.n4886 4.5005
R9581 DVDD.n15712 DVDD.n4886 4.5005
R9582 DVDD.n4899 DVDD.n4886 4.5005
R9583 DVDD.n15714 DVDD.n4886 4.5005
R9584 DVDD.n4896 DVDD.n4886 4.5005
R9585 DVDD.n15750 DVDD.n4886 4.5005
R9586 DVDD.n15752 DVDD.n3517 4.5005
R9587 DVDD.n4904 DVDD.n3517 4.5005
R9588 DVDD.n15707 DVDD.n3517 4.5005
R9589 DVDD.n4903 DVDD.n3517 4.5005
R9590 DVDD.n15709 DVDD.n3517 4.5005
R9591 DVDD.n4902 DVDD.n3517 4.5005
R9592 DVDD.n15710 DVDD.n3517 4.5005
R9593 DVDD.n4901 DVDD.n3517 4.5005
R9594 DVDD.n15711 DVDD.n3517 4.5005
R9595 DVDD.n4900 DVDD.n3517 4.5005
R9596 DVDD.n15712 DVDD.n3517 4.5005
R9597 DVDD.n4899 DVDD.n3517 4.5005
R9598 DVDD.n15714 DVDD.n3517 4.5005
R9599 DVDD.n4896 DVDD.n3517 4.5005
R9600 DVDD.n15750 DVDD.n3517 4.5005
R9601 DVDD.n15752 DVDD.n4887 4.5005
R9602 DVDD.n4904 DVDD.n4887 4.5005
R9603 DVDD.n15707 DVDD.n4887 4.5005
R9604 DVDD.n4903 DVDD.n4887 4.5005
R9605 DVDD.n15709 DVDD.n4887 4.5005
R9606 DVDD.n4902 DVDD.n4887 4.5005
R9607 DVDD.n15710 DVDD.n4887 4.5005
R9608 DVDD.n4901 DVDD.n4887 4.5005
R9609 DVDD.n15711 DVDD.n4887 4.5005
R9610 DVDD.n4900 DVDD.n4887 4.5005
R9611 DVDD.n15712 DVDD.n4887 4.5005
R9612 DVDD.n4899 DVDD.n4887 4.5005
R9613 DVDD.n15714 DVDD.n4887 4.5005
R9614 DVDD.n4896 DVDD.n4887 4.5005
R9615 DVDD.n15750 DVDD.n4887 4.5005
R9616 DVDD.n15752 DVDD.n3516 4.5005
R9617 DVDD.n4904 DVDD.n3516 4.5005
R9618 DVDD.n15707 DVDD.n3516 4.5005
R9619 DVDD.n4903 DVDD.n3516 4.5005
R9620 DVDD.n15709 DVDD.n3516 4.5005
R9621 DVDD.n4902 DVDD.n3516 4.5005
R9622 DVDD.n15710 DVDD.n3516 4.5005
R9623 DVDD.n4901 DVDD.n3516 4.5005
R9624 DVDD.n15711 DVDD.n3516 4.5005
R9625 DVDD.n4900 DVDD.n3516 4.5005
R9626 DVDD.n15712 DVDD.n3516 4.5005
R9627 DVDD.n4899 DVDD.n3516 4.5005
R9628 DVDD.n15714 DVDD.n3516 4.5005
R9629 DVDD.n4896 DVDD.n3516 4.5005
R9630 DVDD.n15750 DVDD.n3516 4.5005
R9631 DVDD.n15711 DVDD.n4888 4.5005
R9632 DVDD.n4900 DVDD.n4888 4.5005
R9633 DVDD.n15712 DVDD.n4888 4.5005
R9634 DVDD.n4899 DVDD.n4888 4.5005
R9635 DVDD.n15714 DVDD.n4888 4.5005
R9636 DVDD.n4896 DVDD.n4888 4.5005
R9637 DVDD.n15750 DVDD.n4888 4.5005
R9638 DVDD.n4901 DVDD.n4888 4.5005
R9639 DVDD.n15710 DVDD.n4888 4.5005
R9640 DVDD.n4902 DVDD.n4888 4.5005
R9641 DVDD.n15709 DVDD.n4888 4.5005
R9642 DVDD.n4903 DVDD.n4888 4.5005
R9643 DVDD.n15707 DVDD.n4888 4.5005
R9644 DVDD.n4904 DVDD.n4888 4.5005
R9645 DVDD.n15752 DVDD.n4888 4.5005
R9646 DVDD.n15711 DVDD.n3515 4.5005
R9647 DVDD.n4900 DVDD.n3515 4.5005
R9648 DVDD.n15712 DVDD.n3515 4.5005
R9649 DVDD.n4899 DVDD.n3515 4.5005
R9650 DVDD.n15714 DVDD.n3515 4.5005
R9651 DVDD.n4896 DVDD.n3515 4.5005
R9652 DVDD.n15750 DVDD.n3515 4.5005
R9653 DVDD.n4901 DVDD.n3515 4.5005
R9654 DVDD.n15710 DVDD.n3515 4.5005
R9655 DVDD.n4902 DVDD.n3515 4.5005
R9656 DVDD.n15709 DVDD.n3515 4.5005
R9657 DVDD.n4903 DVDD.n3515 4.5005
R9658 DVDD.n15707 DVDD.n3515 4.5005
R9659 DVDD.n4904 DVDD.n3515 4.5005
R9660 DVDD.n15752 DVDD.n3515 4.5005
R9661 DVDD.n15711 DVDD.n4889 4.5005
R9662 DVDD.n4900 DVDD.n4889 4.5005
R9663 DVDD.n15712 DVDD.n4889 4.5005
R9664 DVDD.n4899 DVDD.n4889 4.5005
R9665 DVDD.n15714 DVDD.n4889 4.5005
R9666 DVDD.n4896 DVDD.n4889 4.5005
R9667 DVDD.n15750 DVDD.n4889 4.5005
R9668 DVDD.n4901 DVDD.n4889 4.5005
R9669 DVDD.n15710 DVDD.n4889 4.5005
R9670 DVDD.n4902 DVDD.n4889 4.5005
R9671 DVDD.n15709 DVDD.n4889 4.5005
R9672 DVDD.n4903 DVDD.n4889 4.5005
R9673 DVDD.n15707 DVDD.n4889 4.5005
R9674 DVDD.n4904 DVDD.n4889 4.5005
R9675 DVDD.n15752 DVDD.n4889 4.5005
R9676 DVDD.n15752 DVDD.n3514 4.5005
R9677 DVDD.n4904 DVDD.n3514 4.5005
R9678 DVDD.n15707 DVDD.n3514 4.5005
R9679 DVDD.n4903 DVDD.n3514 4.5005
R9680 DVDD.n15709 DVDD.n3514 4.5005
R9681 DVDD.n4902 DVDD.n3514 4.5005
R9682 DVDD.n15710 DVDD.n3514 4.5005
R9683 DVDD.n4901 DVDD.n3514 4.5005
R9684 DVDD.n15711 DVDD.n3514 4.5005
R9685 DVDD.n4900 DVDD.n3514 4.5005
R9686 DVDD.n15712 DVDD.n3514 4.5005
R9687 DVDD.n4899 DVDD.n3514 4.5005
R9688 DVDD.n15714 DVDD.n3514 4.5005
R9689 DVDD.n4896 DVDD.n3514 4.5005
R9690 DVDD.n15750 DVDD.n3514 4.5005
R9691 DVDD.n15752 DVDD.n4890 4.5005
R9692 DVDD.n4904 DVDD.n4890 4.5005
R9693 DVDD.n15707 DVDD.n4890 4.5005
R9694 DVDD.n4903 DVDD.n4890 4.5005
R9695 DVDD.n15709 DVDD.n4890 4.5005
R9696 DVDD.n4902 DVDD.n4890 4.5005
R9697 DVDD.n15710 DVDD.n4890 4.5005
R9698 DVDD.n4901 DVDD.n4890 4.5005
R9699 DVDD.n15711 DVDD.n4890 4.5005
R9700 DVDD.n4900 DVDD.n4890 4.5005
R9701 DVDD.n15712 DVDD.n4890 4.5005
R9702 DVDD.n4899 DVDD.n4890 4.5005
R9703 DVDD.n15714 DVDD.n4890 4.5005
R9704 DVDD.n4896 DVDD.n4890 4.5005
R9705 DVDD.n15750 DVDD.n4890 4.5005
R9706 DVDD.n15752 DVDD.n3513 4.5005
R9707 DVDD.n4904 DVDD.n3513 4.5005
R9708 DVDD.n15707 DVDD.n3513 4.5005
R9709 DVDD.n4903 DVDD.n3513 4.5005
R9710 DVDD.n15709 DVDD.n3513 4.5005
R9711 DVDD.n4902 DVDD.n3513 4.5005
R9712 DVDD.n15710 DVDD.n3513 4.5005
R9713 DVDD.n4901 DVDD.n3513 4.5005
R9714 DVDD.n15711 DVDD.n3513 4.5005
R9715 DVDD.n4900 DVDD.n3513 4.5005
R9716 DVDD.n15712 DVDD.n3513 4.5005
R9717 DVDD.n4899 DVDD.n3513 4.5005
R9718 DVDD.n15714 DVDD.n3513 4.5005
R9719 DVDD.n4896 DVDD.n3513 4.5005
R9720 DVDD.n15750 DVDD.n3513 4.5005
R9721 DVDD.n15752 DVDD.n4891 4.5005
R9722 DVDD.n4904 DVDD.n4891 4.5005
R9723 DVDD.n15707 DVDD.n4891 4.5005
R9724 DVDD.n4903 DVDD.n4891 4.5005
R9725 DVDD.n15709 DVDD.n4891 4.5005
R9726 DVDD.n4902 DVDD.n4891 4.5005
R9727 DVDD.n15710 DVDD.n4891 4.5005
R9728 DVDD.n4901 DVDD.n4891 4.5005
R9729 DVDD.n15711 DVDD.n4891 4.5005
R9730 DVDD.n4900 DVDD.n4891 4.5005
R9731 DVDD.n15712 DVDD.n4891 4.5005
R9732 DVDD.n4899 DVDD.n4891 4.5005
R9733 DVDD.n15714 DVDD.n4891 4.5005
R9734 DVDD.n4896 DVDD.n4891 4.5005
R9735 DVDD.n15750 DVDD.n4891 4.5005
R9736 DVDD.n15711 DVDD.n3512 4.5005
R9737 DVDD.n4900 DVDD.n3512 4.5005
R9738 DVDD.n15712 DVDD.n3512 4.5005
R9739 DVDD.n4899 DVDD.n3512 4.5005
R9740 DVDD.n15714 DVDD.n3512 4.5005
R9741 DVDD.n4896 DVDD.n3512 4.5005
R9742 DVDD.n15750 DVDD.n3512 4.5005
R9743 DVDD.n4901 DVDD.n3512 4.5005
R9744 DVDD.n15710 DVDD.n3512 4.5005
R9745 DVDD.n4902 DVDD.n3512 4.5005
R9746 DVDD.n15709 DVDD.n3512 4.5005
R9747 DVDD.n4903 DVDD.n3512 4.5005
R9748 DVDD.n15707 DVDD.n3512 4.5005
R9749 DVDD.n4904 DVDD.n3512 4.5005
R9750 DVDD.n15752 DVDD.n3512 4.5005
R9751 DVDD.n15711 DVDD.n4892 4.5005
R9752 DVDD.n4900 DVDD.n4892 4.5005
R9753 DVDD.n15712 DVDD.n4892 4.5005
R9754 DVDD.n4899 DVDD.n4892 4.5005
R9755 DVDD.n15714 DVDD.n4892 4.5005
R9756 DVDD.n4896 DVDD.n4892 4.5005
R9757 DVDD.n15750 DVDD.n4892 4.5005
R9758 DVDD.n4901 DVDD.n4892 4.5005
R9759 DVDD.n15710 DVDD.n4892 4.5005
R9760 DVDD.n4902 DVDD.n4892 4.5005
R9761 DVDD.n15709 DVDD.n4892 4.5005
R9762 DVDD.n4903 DVDD.n4892 4.5005
R9763 DVDD.n15707 DVDD.n4892 4.5005
R9764 DVDD.n4904 DVDD.n4892 4.5005
R9765 DVDD.n15752 DVDD.n4892 4.5005
R9766 DVDD.n15711 DVDD.n3511 4.5005
R9767 DVDD.n4900 DVDD.n3511 4.5005
R9768 DVDD.n15712 DVDD.n3511 4.5005
R9769 DVDD.n4899 DVDD.n3511 4.5005
R9770 DVDD.n15714 DVDD.n3511 4.5005
R9771 DVDD.n4896 DVDD.n3511 4.5005
R9772 DVDD.n15750 DVDD.n3511 4.5005
R9773 DVDD.n4901 DVDD.n3511 4.5005
R9774 DVDD.n15710 DVDD.n3511 4.5005
R9775 DVDD.n4902 DVDD.n3511 4.5005
R9776 DVDD.n15709 DVDD.n3511 4.5005
R9777 DVDD.n4903 DVDD.n3511 4.5005
R9778 DVDD.n15707 DVDD.n3511 4.5005
R9779 DVDD.n4904 DVDD.n3511 4.5005
R9780 DVDD.n15752 DVDD.n3511 4.5005
R9781 DVDD.n15752 DVDD.n15751 4.5005
R9782 DVDD.n15751 DVDD.n4904 4.5005
R9783 DVDD.n15751 DVDD.n15707 4.5005
R9784 DVDD.n15751 DVDD.n4903 4.5005
R9785 DVDD.n15751 DVDD.n15709 4.5005
R9786 DVDD.n15751 DVDD.n4902 4.5005
R9787 DVDD.n15751 DVDD.n15710 4.5005
R9788 DVDD.n15751 DVDD.n4901 4.5005
R9789 DVDD.n15751 DVDD.n15711 4.5005
R9790 DVDD.n15751 DVDD.n4900 4.5005
R9791 DVDD.n15751 DVDD.n15712 4.5005
R9792 DVDD.n15751 DVDD.n4899 4.5005
R9793 DVDD.n15751 DVDD.n15714 4.5005
R9794 DVDD.n15751 DVDD.n4896 4.5005
R9795 DVDD.n15751 DVDD.n15750 4.5005
R9796 DVDD.n15701 DVDD.n5048 4.5005
R9797 DVDD.n15701 DVDD.n5046 4.5005
R9798 DVDD.n15701 DVDD.n5049 4.5005
R9799 DVDD.n15701 DVDD.n5045 4.5005
R9800 DVDD.n15701 DVDD.n5050 4.5005
R9801 DVDD.n15701 DVDD.n5043 4.5005
R9802 DVDD.n15701 DVDD.n5051 4.5005
R9803 DVDD.n15701 DVDD.n5042 4.5005
R9804 DVDD.n15701 DVDD.n5052 4.5005
R9805 DVDD.n15701 DVDD.n5041 4.5005
R9806 DVDD.n15701 DVDD.n15700 4.5005
R9807 DVDD.n5066 DVDD.n5048 4.5005
R9808 DVDD.n5066 DVDD.n5046 4.5005
R9809 DVDD.n5066 DVDD.n5049 4.5005
R9810 DVDD.n5066 DVDD.n5045 4.5005
R9811 DVDD.n15698 DVDD.n5066 4.5005
R9812 DVDD.n5078 DVDD.n5066 4.5005
R9813 DVDD.n5066 DVDD.n5050 4.5005
R9814 DVDD.n5066 DVDD.n5043 4.5005
R9815 DVDD.n5066 DVDD.n5051 4.5005
R9816 DVDD.n5066 DVDD.n5042 4.5005
R9817 DVDD.n5066 DVDD.n5052 4.5005
R9818 DVDD.n5066 DVDD.n5041 4.5005
R9819 DVDD.n5081 DVDD.n5066 4.5005
R9820 DVDD.n5079 DVDD.n5066 4.5005
R9821 DVDD.n15700 DVDD.n5066 4.5005
R9822 DVDD.n5064 DVDD.n5051 4.5005
R9823 DVDD.n5064 DVDD.n5042 4.5005
R9824 DVDD.n5064 DVDD.n5052 4.5005
R9825 DVDD.n5064 DVDD.n5041 4.5005
R9826 DVDD.n5081 DVDD.n5064 4.5005
R9827 DVDD.n5079 DVDD.n5064 4.5005
R9828 DVDD.n15700 DVDD.n5064 4.5005
R9829 DVDD.n5064 DVDD.n5043 4.5005
R9830 DVDD.n5064 DVDD.n5050 4.5005
R9831 DVDD.n5078 DVDD.n5064 4.5005
R9832 DVDD.n15698 DVDD.n5064 4.5005
R9833 DVDD.n5064 DVDD.n5045 4.5005
R9834 DVDD.n5064 DVDD.n5049 4.5005
R9835 DVDD.n5064 DVDD.n5046 4.5005
R9836 DVDD.n5064 DVDD.n5048 4.5005
R9837 DVDD.n5067 DVDD.n5051 4.5005
R9838 DVDD.n5067 DVDD.n5042 4.5005
R9839 DVDD.n5067 DVDD.n5052 4.5005
R9840 DVDD.n5067 DVDD.n5041 4.5005
R9841 DVDD.n5081 DVDD.n5067 4.5005
R9842 DVDD.n5079 DVDD.n5067 4.5005
R9843 DVDD.n15700 DVDD.n5067 4.5005
R9844 DVDD.n5067 DVDD.n5043 4.5005
R9845 DVDD.n5067 DVDD.n5050 4.5005
R9846 DVDD.n5078 DVDD.n5067 4.5005
R9847 DVDD.n15698 DVDD.n5067 4.5005
R9848 DVDD.n5067 DVDD.n5045 4.5005
R9849 DVDD.n5067 DVDD.n5049 4.5005
R9850 DVDD.n5067 DVDD.n5046 4.5005
R9851 DVDD.n5067 DVDD.n5048 4.5005
R9852 DVDD.n5063 DVDD.n5051 4.5005
R9853 DVDD.n5063 DVDD.n5042 4.5005
R9854 DVDD.n5063 DVDD.n5052 4.5005
R9855 DVDD.n5063 DVDD.n5041 4.5005
R9856 DVDD.n5081 DVDD.n5063 4.5005
R9857 DVDD.n5079 DVDD.n5063 4.5005
R9858 DVDD.n15700 DVDD.n5063 4.5005
R9859 DVDD.n5063 DVDD.n5043 4.5005
R9860 DVDD.n5063 DVDD.n5050 4.5005
R9861 DVDD.n5078 DVDD.n5063 4.5005
R9862 DVDD.n15698 DVDD.n5063 4.5005
R9863 DVDD.n5063 DVDD.n5045 4.5005
R9864 DVDD.n5063 DVDD.n5049 4.5005
R9865 DVDD.n5063 DVDD.n5046 4.5005
R9866 DVDD.n5063 DVDD.n5048 4.5005
R9867 DVDD.n5068 DVDD.n5048 4.5005
R9868 DVDD.n5068 DVDD.n5046 4.5005
R9869 DVDD.n5068 DVDD.n5049 4.5005
R9870 DVDD.n5068 DVDD.n5045 4.5005
R9871 DVDD.n15698 DVDD.n5068 4.5005
R9872 DVDD.n5078 DVDD.n5068 4.5005
R9873 DVDD.n5068 DVDD.n5050 4.5005
R9874 DVDD.n5068 DVDD.n5043 4.5005
R9875 DVDD.n5068 DVDD.n5051 4.5005
R9876 DVDD.n5068 DVDD.n5042 4.5005
R9877 DVDD.n5068 DVDD.n5052 4.5005
R9878 DVDD.n5068 DVDD.n5041 4.5005
R9879 DVDD.n5081 DVDD.n5068 4.5005
R9880 DVDD.n5079 DVDD.n5068 4.5005
R9881 DVDD.n15700 DVDD.n5068 4.5005
R9882 DVDD.n5062 DVDD.n5048 4.5005
R9883 DVDD.n5062 DVDD.n5046 4.5005
R9884 DVDD.n5062 DVDD.n5049 4.5005
R9885 DVDD.n5062 DVDD.n5045 4.5005
R9886 DVDD.n15698 DVDD.n5062 4.5005
R9887 DVDD.n5078 DVDD.n5062 4.5005
R9888 DVDD.n5062 DVDD.n5050 4.5005
R9889 DVDD.n5062 DVDD.n5043 4.5005
R9890 DVDD.n5062 DVDD.n5051 4.5005
R9891 DVDD.n5062 DVDD.n5042 4.5005
R9892 DVDD.n5062 DVDD.n5052 4.5005
R9893 DVDD.n5062 DVDD.n5041 4.5005
R9894 DVDD.n5081 DVDD.n5062 4.5005
R9895 DVDD.n5079 DVDD.n5062 4.5005
R9896 DVDD.n15700 DVDD.n5062 4.5005
R9897 DVDD.n5069 DVDD.n5048 4.5005
R9898 DVDD.n5069 DVDD.n5046 4.5005
R9899 DVDD.n5069 DVDD.n5049 4.5005
R9900 DVDD.n5069 DVDD.n5045 4.5005
R9901 DVDD.n15698 DVDD.n5069 4.5005
R9902 DVDD.n5078 DVDD.n5069 4.5005
R9903 DVDD.n5069 DVDD.n5050 4.5005
R9904 DVDD.n5069 DVDD.n5043 4.5005
R9905 DVDD.n5069 DVDD.n5051 4.5005
R9906 DVDD.n5069 DVDD.n5042 4.5005
R9907 DVDD.n5069 DVDD.n5052 4.5005
R9908 DVDD.n5069 DVDD.n5041 4.5005
R9909 DVDD.n5081 DVDD.n5069 4.5005
R9910 DVDD.n5079 DVDD.n5069 4.5005
R9911 DVDD.n15700 DVDD.n5069 4.5005
R9912 DVDD.n5061 DVDD.n5048 4.5005
R9913 DVDD.n5061 DVDD.n5046 4.5005
R9914 DVDD.n5061 DVDD.n5049 4.5005
R9915 DVDD.n5061 DVDD.n5045 4.5005
R9916 DVDD.n15698 DVDD.n5061 4.5005
R9917 DVDD.n5078 DVDD.n5061 4.5005
R9918 DVDD.n5061 DVDD.n5050 4.5005
R9919 DVDD.n5061 DVDD.n5043 4.5005
R9920 DVDD.n5061 DVDD.n5051 4.5005
R9921 DVDD.n5061 DVDD.n5042 4.5005
R9922 DVDD.n5061 DVDD.n5052 4.5005
R9923 DVDD.n5061 DVDD.n5041 4.5005
R9924 DVDD.n5081 DVDD.n5061 4.5005
R9925 DVDD.n5079 DVDD.n5061 4.5005
R9926 DVDD.n15700 DVDD.n5061 4.5005
R9927 DVDD.n5070 DVDD.n5051 4.5005
R9928 DVDD.n5070 DVDD.n5042 4.5005
R9929 DVDD.n5070 DVDD.n5052 4.5005
R9930 DVDD.n5070 DVDD.n5041 4.5005
R9931 DVDD.n5081 DVDD.n5070 4.5005
R9932 DVDD.n5079 DVDD.n5070 4.5005
R9933 DVDD.n15700 DVDD.n5070 4.5005
R9934 DVDD.n5070 DVDD.n5043 4.5005
R9935 DVDD.n5070 DVDD.n5050 4.5005
R9936 DVDD.n5078 DVDD.n5070 4.5005
R9937 DVDD.n15698 DVDD.n5070 4.5005
R9938 DVDD.n5070 DVDD.n5045 4.5005
R9939 DVDD.n5070 DVDD.n5049 4.5005
R9940 DVDD.n5070 DVDD.n5046 4.5005
R9941 DVDD.n5070 DVDD.n5048 4.5005
R9942 DVDD.n5060 DVDD.n5051 4.5005
R9943 DVDD.n5060 DVDD.n5042 4.5005
R9944 DVDD.n5060 DVDD.n5052 4.5005
R9945 DVDD.n5060 DVDD.n5041 4.5005
R9946 DVDD.n5081 DVDD.n5060 4.5005
R9947 DVDD.n5079 DVDD.n5060 4.5005
R9948 DVDD.n15700 DVDD.n5060 4.5005
R9949 DVDD.n5060 DVDD.n5043 4.5005
R9950 DVDD.n5060 DVDD.n5050 4.5005
R9951 DVDD.n5078 DVDD.n5060 4.5005
R9952 DVDD.n15698 DVDD.n5060 4.5005
R9953 DVDD.n5060 DVDD.n5045 4.5005
R9954 DVDD.n5060 DVDD.n5049 4.5005
R9955 DVDD.n5060 DVDD.n5046 4.5005
R9956 DVDD.n5060 DVDD.n5048 4.5005
R9957 DVDD.n5071 DVDD.n5051 4.5005
R9958 DVDD.n5071 DVDD.n5042 4.5005
R9959 DVDD.n5071 DVDD.n5052 4.5005
R9960 DVDD.n5071 DVDD.n5041 4.5005
R9961 DVDD.n5081 DVDD.n5071 4.5005
R9962 DVDD.n5079 DVDD.n5071 4.5005
R9963 DVDD.n15700 DVDD.n5071 4.5005
R9964 DVDD.n5071 DVDD.n5043 4.5005
R9965 DVDD.n5071 DVDD.n5050 4.5005
R9966 DVDD.n5078 DVDD.n5071 4.5005
R9967 DVDD.n15698 DVDD.n5071 4.5005
R9968 DVDD.n5071 DVDD.n5045 4.5005
R9969 DVDD.n5071 DVDD.n5049 4.5005
R9970 DVDD.n5071 DVDD.n5046 4.5005
R9971 DVDD.n5071 DVDD.n5048 4.5005
R9972 DVDD.n5059 DVDD.n5048 4.5005
R9973 DVDD.n5059 DVDD.n5046 4.5005
R9974 DVDD.n5059 DVDD.n5049 4.5005
R9975 DVDD.n5059 DVDD.n5045 4.5005
R9976 DVDD.n15698 DVDD.n5059 4.5005
R9977 DVDD.n5078 DVDD.n5059 4.5005
R9978 DVDD.n5059 DVDD.n5050 4.5005
R9979 DVDD.n5059 DVDD.n5043 4.5005
R9980 DVDD.n5059 DVDD.n5051 4.5005
R9981 DVDD.n5059 DVDD.n5042 4.5005
R9982 DVDD.n5059 DVDD.n5052 4.5005
R9983 DVDD.n5059 DVDD.n5041 4.5005
R9984 DVDD.n5081 DVDD.n5059 4.5005
R9985 DVDD.n5079 DVDD.n5059 4.5005
R9986 DVDD.n15700 DVDD.n5059 4.5005
R9987 DVDD.n5072 DVDD.n5048 4.5005
R9988 DVDD.n5072 DVDD.n5046 4.5005
R9989 DVDD.n5072 DVDD.n5049 4.5005
R9990 DVDD.n5072 DVDD.n5045 4.5005
R9991 DVDD.n15698 DVDD.n5072 4.5005
R9992 DVDD.n5078 DVDD.n5072 4.5005
R9993 DVDD.n5072 DVDD.n5050 4.5005
R9994 DVDD.n5072 DVDD.n5043 4.5005
R9995 DVDD.n5072 DVDD.n5051 4.5005
R9996 DVDD.n5072 DVDD.n5042 4.5005
R9997 DVDD.n5072 DVDD.n5052 4.5005
R9998 DVDD.n5072 DVDD.n5041 4.5005
R9999 DVDD.n5081 DVDD.n5072 4.5005
R10000 DVDD.n5079 DVDD.n5072 4.5005
R10001 DVDD.n15700 DVDD.n5072 4.5005
R10002 DVDD.n5058 DVDD.n5048 4.5005
R10003 DVDD.n5058 DVDD.n5046 4.5005
R10004 DVDD.n5058 DVDD.n5049 4.5005
R10005 DVDD.n5058 DVDD.n5045 4.5005
R10006 DVDD.n15698 DVDD.n5058 4.5005
R10007 DVDD.n5078 DVDD.n5058 4.5005
R10008 DVDD.n5058 DVDD.n5050 4.5005
R10009 DVDD.n5058 DVDD.n5043 4.5005
R10010 DVDD.n5058 DVDD.n5051 4.5005
R10011 DVDD.n5058 DVDD.n5042 4.5005
R10012 DVDD.n5058 DVDD.n5052 4.5005
R10013 DVDD.n5058 DVDD.n5041 4.5005
R10014 DVDD.n5081 DVDD.n5058 4.5005
R10015 DVDD.n5079 DVDD.n5058 4.5005
R10016 DVDD.n15700 DVDD.n5058 4.5005
R10017 DVDD.n5073 DVDD.n5051 4.5005
R10018 DVDD.n5073 DVDD.n5042 4.5005
R10019 DVDD.n5073 DVDD.n5052 4.5005
R10020 DVDD.n5073 DVDD.n5041 4.5005
R10021 DVDD.n5081 DVDD.n5073 4.5005
R10022 DVDD.n5079 DVDD.n5073 4.5005
R10023 DVDD.n15700 DVDD.n5073 4.5005
R10024 DVDD.n5073 DVDD.n5043 4.5005
R10025 DVDD.n5073 DVDD.n5050 4.5005
R10026 DVDD.n5078 DVDD.n5073 4.5005
R10027 DVDD.n15698 DVDD.n5073 4.5005
R10028 DVDD.n5073 DVDD.n5045 4.5005
R10029 DVDD.n5073 DVDD.n5049 4.5005
R10030 DVDD.n5073 DVDD.n5046 4.5005
R10031 DVDD.n5073 DVDD.n5048 4.5005
R10032 DVDD.n5057 DVDD.n5051 4.5005
R10033 DVDD.n5057 DVDD.n5042 4.5005
R10034 DVDD.n5057 DVDD.n5052 4.5005
R10035 DVDD.n5057 DVDD.n5041 4.5005
R10036 DVDD.n5081 DVDD.n5057 4.5005
R10037 DVDD.n5079 DVDD.n5057 4.5005
R10038 DVDD.n15700 DVDD.n5057 4.5005
R10039 DVDD.n5057 DVDD.n5043 4.5005
R10040 DVDD.n5057 DVDD.n5050 4.5005
R10041 DVDD.n5078 DVDD.n5057 4.5005
R10042 DVDD.n15698 DVDD.n5057 4.5005
R10043 DVDD.n5057 DVDD.n5045 4.5005
R10044 DVDD.n5057 DVDD.n5049 4.5005
R10045 DVDD.n5057 DVDD.n5046 4.5005
R10046 DVDD.n5057 DVDD.n5048 4.5005
R10047 DVDD.n5074 DVDD.n5051 4.5005
R10048 DVDD.n5074 DVDD.n5042 4.5005
R10049 DVDD.n5074 DVDD.n5052 4.5005
R10050 DVDD.n5074 DVDD.n5041 4.5005
R10051 DVDD.n5081 DVDD.n5074 4.5005
R10052 DVDD.n5079 DVDD.n5074 4.5005
R10053 DVDD.n15700 DVDD.n5074 4.5005
R10054 DVDD.n5074 DVDD.n5043 4.5005
R10055 DVDD.n5074 DVDD.n5050 4.5005
R10056 DVDD.n5078 DVDD.n5074 4.5005
R10057 DVDD.n15698 DVDD.n5074 4.5005
R10058 DVDD.n5074 DVDD.n5045 4.5005
R10059 DVDD.n5074 DVDD.n5049 4.5005
R10060 DVDD.n5074 DVDD.n5046 4.5005
R10061 DVDD.n5074 DVDD.n5048 4.5005
R10062 DVDD.n5056 DVDD.n5051 4.5005
R10063 DVDD.n5056 DVDD.n5042 4.5005
R10064 DVDD.n5056 DVDD.n5052 4.5005
R10065 DVDD.n5056 DVDD.n5041 4.5005
R10066 DVDD.n5081 DVDD.n5056 4.5005
R10067 DVDD.n5079 DVDD.n5056 4.5005
R10068 DVDD.n15700 DVDD.n5056 4.5005
R10069 DVDD.n5056 DVDD.n5043 4.5005
R10070 DVDD.n5056 DVDD.n5050 4.5005
R10071 DVDD.n5078 DVDD.n5056 4.5005
R10072 DVDD.n15698 DVDD.n5056 4.5005
R10073 DVDD.n5056 DVDD.n5045 4.5005
R10074 DVDD.n5056 DVDD.n5049 4.5005
R10075 DVDD.n5056 DVDD.n5046 4.5005
R10076 DVDD.n5056 DVDD.n5048 4.5005
R10077 DVDD.n5075 DVDD.n5048 4.5005
R10078 DVDD.n5075 DVDD.n5046 4.5005
R10079 DVDD.n5075 DVDD.n5049 4.5005
R10080 DVDD.n5075 DVDD.n5045 4.5005
R10081 DVDD.n15698 DVDD.n5075 4.5005
R10082 DVDD.n5078 DVDD.n5075 4.5005
R10083 DVDD.n5075 DVDD.n5050 4.5005
R10084 DVDD.n5075 DVDD.n5043 4.5005
R10085 DVDD.n5075 DVDD.n5051 4.5005
R10086 DVDD.n5075 DVDD.n5042 4.5005
R10087 DVDD.n5075 DVDD.n5052 4.5005
R10088 DVDD.n5075 DVDD.n5041 4.5005
R10089 DVDD.n5081 DVDD.n5075 4.5005
R10090 DVDD.n5079 DVDD.n5075 4.5005
R10091 DVDD.n15700 DVDD.n5075 4.5005
R10092 DVDD.n5055 DVDD.n5048 4.5005
R10093 DVDD.n5055 DVDD.n5046 4.5005
R10094 DVDD.n5055 DVDD.n5049 4.5005
R10095 DVDD.n5055 DVDD.n5045 4.5005
R10096 DVDD.n15698 DVDD.n5055 4.5005
R10097 DVDD.n5078 DVDD.n5055 4.5005
R10098 DVDD.n5055 DVDD.n5050 4.5005
R10099 DVDD.n5055 DVDD.n5043 4.5005
R10100 DVDD.n5055 DVDD.n5051 4.5005
R10101 DVDD.n5055 DVDD.n5042 4.5005
R10102 DVDD.n5055 DVDD.n5052 4.5005
R10103 DVDD.n5055 DVDD.n5041 4.5005
R10104 DVDD.n5081 DVDD.n5055 4.5005
R10105 DVDD.n5079 DVDD.n5055 4.5005
R10106 DVDD.n15700 DVDD.n5055 4.5005
R10107 DVDD.n5076 DVDD.n5048 4.5005
R10108 DVDD.n5076 DVDD.n5046 4.5005
R10109 DVDD.n5076 DVDD.n5049 4.5005
R10110 DVDD.n5076 DVDD.n5045 4.5005
R10111 DVDD.n15698 DVDD.n5076 4.5005
R10112 DVDD.n5078 DVDD.n5076 4.5005
R10113 DVDD.n5076 DVDD.n5050 4.5005
R10114 DVDD.n5076 DVDD.n5043 4.5005
R10115 DVDD.n5076 DVDD.n5051 4.5005
R10116 DVDD.n5076 DVDD.n5042 4.5005
R10117 DVDD.n5076 DVDD.n5052 4.5005
R10118 DVDD.n5076 DVDD.n5041 4.5005
R10119 DVDD.n5081 DVDD.n5076 4.5005
R10120 DVDD.n5079 DVDD.n5076 4.5005
R10121 DVDD.n15700 DVDD.n5076 4.5005
R10122 DVDD.n5054 DVDD.n5051 4.5005
R10123 DVDD.n5054 DVDD.n5042 4.5005
R10124 DVDD.n5054 DVDD.n5052 4.5005
R10125 DVDD.n5054 DVDD.n5041 4.5005
R10126 DVDD.n5081 DVDD.n5054 4.5005
R10127 DVDD.n5079 DVDD.n5054 4.5005
R10128 DVDD.n15700 DVDD.n5054 4.5005
R10129 DVDD.n5054 DVDD.n5043 4.5005
R10130 DVDD.n5054 DVDD.n5050 4.5005
R10131 DVDD.n5078 DVDD.n5054 4.5005
R10132 DVDD.n15698 DVDD.n5054 4.5005
R10133 DVDD.n5054 DVDD.n5045 4.5005
R10134 DVDD.n5054 DVDD.n5049 4.5005
R10135 DVDD.n5054 DVDD.n5046 4.5005
R10136 DVDD.n5054 DVDD.n5048 4.5005
R10137 DVDD.n15699 DVDD.n5051 4.5005
R10138 DVDD.n15699 DVDD.n5042 4.5005
R10139 DVDD.n15699 DVDD.n5052 4.5005
R10140 DVDD.n15699 DVDD.n5041 4.5005
R10141 DVDD.n15699 DVDD.n5081 4.5005
R10142 DVDD.n15699 DVDD.n5079 4.5005
R10143 DVDD.n15700 DVDD.n15699 4.5005
R10144 DVDD.n15699 DVDD.n5043 4.5005
R10145 DVDD.n15699 DVDD.n5050 4.5005
R10146 DVDD.n15699 DVDD.n5078 4.5005
R10147 DVDD.n15699 DVDD.n15698 4.5005
R10148 DVDD.n15699 DVDD.n5045 4.5005
R10149 DVDD.n15699 DVDD.n5049 4.5005
R10150 DVDD.n15699 DVDD.n5046 4.5005
R10151 DVDD.n15699 DVDD.n5048 4.5005
R10152 DVDD.n15420 DVDD.n5241 4.5005
R10153 DVDD.n5256 DVDD.n5241 4.5005
R10154 DVDD.n15421 DVDD.n5241 4.5005
R10155 DVDD.n5255 DVDD.n5241 4.5005
R10156 DVDD.n15459 DVDD.n5241 4.5005
R10157 DVDD.n5257 DVDD.n5241 4.5005
R10158 DVDD.n15419 DVDD.n5241 4.5005
R10159 DVDD.n5259 DVDD.n5241 4.5005
R10160 DVDD.n15416 DVDD.n5241 4.5005
R10161 DVDD.n5260 DVDD.n5241 4.5005
R10162 DVDD.n15461 DVDD.n5241 4.5005
R10163 DVDD.n15461 DVDD.n5242 4.5005
R10164 DVDD.n5260 DVDD.n5242 4.5005
R10165 DVDD.n15416 DVDD.n5242 4.5005
R10166 DVDD.n5259 DVDD.n5242 4.5005
R10167 DVDD.n15418 DVDD.n5242 4.5005
R10168 DVDD.n5258 DVDD.n5242 4.5005
R10169 DVDD.n15419 DVDD.n5242 4.5005
R10170 DVDD.n5257 DVDD.n5242 4.5005
R10171 DVDD.n15420 DVDD.n5242 4.5005
R10172 DVDD.n5256 DVDD.n5242 4.5005
R10173 DVDD.n15421 DVDD.n5242 4.5005
R10174 DVDD.n5255 DVDD.n5242 4.5005
R10175 DVDD.n15423 DVDD.n5242 4.5005
R10176 DVDD.n5254 DVDD.n5242 4.5005
R10177 DVDD.n15459 DVDD.n5242 4.5005
R10178 DVDD.n15461 DVDD.n5240 4.5005
R10179 DVDD.n5260 DVDD.n5240 4.5005
R10180 DVDD.n15416 DVDD.n5240 4.5005
R10181 DVDD.n5259 DVDD.n5240 4.5005
R10182 DVDD.n15418 DVDD.n5240 4.5005
R10183 DVDD.n5258 DVDD.n5240 4.5005
R10184 DVDD.n15419 DVDD.n5240 4.5005
R10185 DVDD.n5257 DVDD.n5240 4.5005
R10186 DVDD.n15420 DVDD.n5240 4.5005
R10187 DVDD.n5256 DVDD.n5240 4.5005
R10188 DVDD.n15421 DVDD.n5240 4.5005
R10189 DVDD.n5255 DVDD.n5240 4.5005
R10190 DVDD.n15423 DVDD.n5240 4.5005
R10191 DVDD.n5254 DVDD.n5240 4.5005
R10192 DVDD.n15459 DVDD.n5240 4.5005
R10193 DVDD.n15461 DVDD.n5243 4.5005
R10194 DVDD.n5260 DVDD.n5243 4.5005
R10195 DVDD.n15416 DVDD.n5243 4.5005
R10196 DVDD.n5259 DVDD.n5243 4.5005
R10197 DVDD.n15418 DVDD.n5243 4.5005
R10198 DVDD.n5258 DVDD.n5243 4.5005
R10199 DVDD.n15419 DVDD.n5243 4.5005
R10200 DVDD.n5257 DVDD.n5243 4.5005
R10201 DVDD.n15420 DVDD.n5243 4.5005
R10202 DVDD.n5256 DVDD.n5243 4.5005
R10203 DVDD.n15421 DVDD.n5243 4.5005
R10204 DVDD.n5255 DVDD.n5243 4.5005
R10205 DVDD.n15423 DVDD.n5243 4.5005
R10206 DVDD.n5254 DVDD.n5243 4.5005
R10207 DVDD.n15459 DVDD.n5243 4.5005
R10208 DVDD.n15420 DVDD.n5239 4.5005
R10209 DVDD.n5256 DVDD.n5239 4.5005
R10210 DVDD.n15421 DVDD.n5239 4.5005
R10211 DVDD.n5255 DVDD.n5239 4.5005
R10212 DVDD.n15423 DVDD.n5239 4.5005
R10213 DVDD.n5254 DVDD.n5239 4.5005
R10214 DVDD.n15459 DVDD.n5239 4.5005
R10215 DVDD.n5257 DVDD.n5239 4.5005
R10216 DVDD.n15419 DVDD.n5239 4.5005
R10217 DVDD.n5258 DVDD.n5239 4.5005
R10218 DVDD.n15418 DVDD.n5239 4.5005
R10219 DVDD.n5259 DVDD.n5239 4.5005
R10220 DVDD.n15416 DVDD.n5239 4.5005
R10221 DVDD.n5260 DVDD.n5239 4.5005
R10222 DVDD.n15461 DVDD.n5239 4.5005
R10223 DVDD.n15420 DVDD.n5244 4.5005
R10224 DVDD.n5256 DVDD.n5244 4.5005
R10225 DVDD.n15421 DVDD.n5244 4.5005
R10226 DVDD.n5255 DVDD.n5244 4.5005
R10227 DVDD.n15423 DVDD.n5244 4.5005
R10228 DVDD.n5254 DVDD.n5244 4.5005
R10229 DVDD.n15459 DVDD.n5244 4.5005
R10230 DVDD.n5257 DVDD.n5244 4.5005
R10231 DVDD.n15419 DVDD.n5244 4.5005
R10232 DVDD.n5258 DVDD.n5244 4.5005
R10233 DVDD.n15418 DVDD.n5244 4.5005
R10234 DVDD.n5259 DVDD.n5244 4.5005
R10235 DVDD.n15416 DVDD.n5244 4.5005
R10236 DVDD.n5260 DVDD.n5244 4.5005
R10237 DVDD.n15461 DVDD.n5244 4.5005
R10238 DVDD.n15420 DVDD.n5238 4.5005
R10239 DVDD.n5256 DVDD.n5238 4.5005
R10240 DVDD.n15421 DVDD.n5238 4.5005
R10241 DVDD.n5255 DVDD.n5238 4.5005
R10242 DVDD.n15423 DVDD.n5238 4.5005
R10243 DVDD.n5254 DVDD.n5238 4.5005
R10244 DVDD.n15459 DVDD.n5238 4.5005
R10245 DVDD.n5257 DVDD.n5238 4.5005
R10246 DVDD.n15419 DVDD.n5238 4.5005
R10247 DVDD.n5258 DVDD.n5238 4.5005
R10248 DVDD.n15418 DVDD.n5238 4.5005
R10249 DVDD.n5259 DVDD.n5238 4.5005
R10250 DVDD.n15416 DVDD.n5238 4.5005
R10251 DVDD.n5260 DVDD.n5238 4.5005
R10252 DVDD.n15461 DVDD.n5238 4.5005
R10253 DVDD.n15420 DVDD.n5245 4.5005
R10254 DVDD.n5256 DVDD.n5245 4.5005
R10255 DVDD.n15421 DVDD.n5245 4.5005
R10256 DVDD.n5255 DVDD.n5245 4.5005
R10257 DVDD.n15423 DVDD.n5245 4.5005
R10258 DVDD.n5254 DVDD.n5245 4.5005
R10259 DVDD.n15459 DVDD.n5245 4.5005
R10260 DVDD.n5257 DVDD.n5245 4.5005
R10261 DVDD.n15419 DVDD.n5245 4.5005
R10262 DVDD.n5258 DVDD.n5245 4.5005
R10263 DVDD.n15418 DVDD.n5245 4.5005
R10264 DVDD.n5259 DVDD.n5245 4.5005
R10265 DVDD.n15416 DVDD.n5245 4.5005
R10266 DVDD.n5260 DVDD.n5245 4.5005
R10267 DVDD.n15461 DVDD.n5245 4.5005
R10268 DVDD.n15461 DVDD.n5237 4.5005
R10269 DVDD.n5260 DVDD.n5237 4.5005
R10270 DVDD.n15416 DVDD.n5237 4.5005
R10271 DVDD.n5259 DVDD.n5237 4.5005
R10272 DVDD.n15418 DVDD.n5237 4.5005
R10273 DVDD.n5258 DVDD.n5237 4.5005
R10274 DVDD.n15419 DVDD.n5237 4.5005
R10275 DVDD.n5257 DVDD.n5237 4.5005
R10276 DVDD.n15420 DVDD.n5237 4.5005
R10277 DVDD.n5256 DVDD.n5237 4.5005
R10278 DVDD.n15421 DVDD.n5237 4.5005
R10279 DVDD.n5255 DVDD.n5237 4.5005
R10280 DVDD.n15423 DVDD.n5237 4.5005
R10281 DVDD.n5254 DVDD.n5237 4.5005
R10282 DVDD.n15459 DVDD.n5237 4.5005
R10283 DVDD.n15461 DVDD.n5246 4.5005
R10284 DVDD.n5260 DVDD.n5246 4.5005
R10285 DVDD.n15416 DVDD.n5246 4.5005
R10286 DVDD.n5259 DVDD.n5246 4.5005
R10287 DVDD.n15418 DVDD.n5246 4.5005
R10288 DVDD.n5258 DVDD.n5246 4.5005
R10289 DVDD.n15419 DVDD.n5246 4.5005
R10290 DVDD.n5257 DVDD.n5246 4.5005
R10291 DVDD.n15420 DVDD.n5246 4.5005
R10292 DVDD.n5256 DVDD.n5246 4.5005
R10293 DVDD.n15421 DVDD.n5246 4.5005
R10294 DVDD.n5255 DVDD.n5246 4.5005
R10295 DVDD.n15423 DVDD.n5246 4.5005
R10296 DVDD.n5254 DVDD.n5246 4.5005
R10297 DVDD.n15459 DVDD.n5246 4.5005
R10298 DVDD.n15461 DVDD.n5236 4.5005
R10299 DVDD.n5260 DVDD.n5236 4.5005
R10300 DVDD.n15416 DVDD.n5236 4.5005
R10301 DVDD.n5259 DVDD.n5236 4.5005
R10302 DVDD.n15418 DVDD.n5236 4.5005
R10303 DVDD.n5258 DVDD.n5236 4.5005
R10304 DVDD.n15419 DVDD.n5236 4.5005
R10305 DVDD.n5257 DVDD.n5236 4.5005
R10306 DVDD.n15420 DVDD.n5236 4.5005
R10307 DVDD.n5256 DVDD.n5236 4.5005
R10308 DVDD.n15421 DVDD.n5236 4.5005
R10309 DVDD.n5255 DVDD.n5236 4.5005
R10310 DVDD.n15423 DVDD.n5236 4.5005
R10311 DVDD.n5254 DVDD.n5236 4.5005
R10312 DVDD.n15459 DVDD.n5236 4.5005
R10313 DVDD.n15420 DVDD.n5247 4.5005
R10314 DVDD.n5256 DVDD.n5247 4.5005
R10315 DVDD.n15421 DVDD.n5247 4.5005
R10316 DVDD.n5255 DVDD.n5247 4.5005
R10317 DVDD.n15423 DVDD.n5247 4.5005
R10318 DVDD.n5254 DVDD.n5247 4.5005
R10319 DVDD.n15459 DVDD.n5247 4.5005
R10320 DVDD.n5257 DVDD.n5247 4.5005
R10321 DVDD.n15419 DVDD.n5247 4.5005
R10322 DVDD.n5258 DVDD.n5247 4.5005
R10323 DVDD.n15418 DVDD.n5247 4.5005
R10324 DVDD.n5259 DVDD.n5247 4.5005
R10325 DVDD.n15416 DVDD.n5247 4.5005
R10326 DVDD.n5260 DVDD.n5247 4.5005
R10327 DVDD.n15461 DVDD.n5247 4.5005
R10328 DVDD.n15420 DVDD.n5235 4.5005
R10329 DVDD.n5256 DVDD.n5235 4.5005
R10330 DVDD.n15421 DVDD.n5235 4.5005
R10331 DVDD.n5255 DVDD.n5235 4.5005
R10332 DVDD.n15423 DVDD.n5235 4.5005
R10333 DVDD.n5254 DVDD.n5235 4.5005
R10334 DVDD.n15459 DVDD.n5235 4.5005
R10335 DVDD.n5257 DVDD.n5235 4.5005
R10336 DVDD.n15419 DVDD.n5235 4.5005
R10337 DVDD.n5258 DVDD.n5235 4.5005
R10338 DVDD.n15418 DVDD.n5235 4.5005
R10339 DVDD.n5259 DVDD.n5235 4.5005
R10340 DVDD.n15416 DVDD.n5235 4.5005
R10341 DVDD.n5260 DVDD.n5235 4.5005
R10342 DVDD.n15461 DVDD.n5235 4.5005
R10343 DVDD.n15420 DVDD.n5248 4.5005
R10344 DVDD.n5256 DVDD.n5248 4.5005
R10345 DVDD.n15421 DVDD.n5248 4.5005
R10346 DVDD.n5255 DVDD.n5248 4.5005
R10347 DVDD.n15423 DVDD.n5248 4.5005
R10348 DVDD.n5254 DVDD.n5248 4.5005
R10349 DVDD.n15459 DVDD.n5248 4.5005
R10350 DVDD.n5257 DVDD.n5248 4.5005
R10351 DVDD.n15419 DVDD.n5248 4.5005
R10352 DVDD.n5258 DVDD.n5248 4.5005
R10353 DVDD.n15418 DVDD.n5248 4.5005
R10354 DVDD.n5259 DVDD.n5248 4.5005
R10355 DVDD.n15416 DVDD.n5248 4.5005
R10356 DVDD.n5260 DVDD.n5248 4.5005
R10357 DVDD.n15461 DVDD.n5248 4.5005
R10358 DVDD.n15461 DVDD.n5234 4.5005
R10359 DVDD.n5260 DVDD.n5234 4.5005
R10360 DVDD.n15416 DVDD.n5234 4.5005
R10361 DVDD.n5259 DVDD.n5234 4.5005
R10362 DVDD.n15418 DVDD.n5234 4.5005
R10363 DVDD.n5258 DVDD.n5234 4.5005
R10364 DVDD.n15419 DVDD.n5234 4.5005
R10365 DVDD.n5257 DVDD.n5234 4.5005
R10366 DVDD.n15420 DVDD.n5234 4.5005
R10367 DVDD.n5256 DVDD.n5234 4.5005
R10368 DVDD.n15421 DVDD.n5234 4.5005
R10369 DVDD.n5255 DVDD.n5234 4.5005
R10370 DVDD.n15423 DVDD.n5234 4.5005
R10371 DVDD.n5254 DVDD.n5234 4.5005
R10372 DVDD.n15459 DVDD.n5234 4.5005
R10373 DVDD.n15461 DVDD.n5249 4.5005
R10374 DVDD.n5260 DVDD.n5249 4.5005
R10375 DVDD.n15416 DVDD.n5249 4.5005
R10376 DVDD.n5259 DVDD.n5249 4.5005
R10377 DVDD.n15418 DVDD.n5249 4.5005
R10378 DVDD.n5258 DVDD.n5249 4.5005
R10379 DVDD.n15419 DVDD.n5249 4.5005
R10380 DVDD.n5257 DVDD.n5249 4.5005
R10381 DVDD.n15420 DVDD.n5249 4.5005
R10382 DVDD.n5256 DVDD.n5249 4.5005
R10383 DVDD.n15421 DVDD.n5249 4.5005
R10384 DVDD.n5255 DVDD.n5249 4.5005
R10385 DVDD.n15423 DVDD.n5249 4.5005
R10386 DVDD.n5254 DVDD.n5249 4.5005
R10387 DVDD.n15459 DVDD.n5249 4.5005
R10388 DVDD.n15461 DVDD.n5233 4.5005
R10389 DVDD.n5260 DVDD.n5233 4.5005
R10390 DVDD.n15416 DVDD.n5233 4.5005
R10391 DVDD.n5259 DVDD.n5233 4.5005
R10392 DVDD.n15418 DVDD.n5233 4.5005
R10393 DVDD.n5258 DVDD.n5233 4.5005
R10394 DVDD.n15419 DVDD.n5233 4.5005
R10395 DVDD.n5257 DVDD.n5233 4.5005
R10396 DVDD.n15420 DVDD.n5233 4.5005
R10397 DVDD.n5256 DVDD.n5233 4.5005
R10398 DVDD.n15421 DVDD.n5233 4.5005
R10399 DVDD.n5255 DVDD.n5233 4.5005
R10400 DVDD.n15423 DVDD.n5233 4.5005
R10401 DVDD.n5254 DVDD.n5233 4.5005
R10402 DVDD.n15459 DVDD.n5233 4.5005
R10403 DVDD.n15461 DVDD.n5250 4.5005
R10404 DVDD.n5260 DVDD.n5250 4.5005
R10405 DVDD.n15416 DVDD.n5250 4.5005
R10406 DVDD.n5259 DVDD.n5250 4.5005
R10407 DVDD.n15418 DVDD.n5250 4.5005
R10408 DVDD.n5258 DVDD.n5250 4.5005
R10409 DVDD.n15419 DVDD.n5250 4.5005
R10410 DVDD.n5257 DVDD.n5250 4.5005
R10411 DVDD.n15420 DVDD.n5250 4.5005
R10412 DVDD.n5256 DVDD.n5250 4.5005
R10413 DVDD.n15421 DVDD.n5250 4.5005
R10414 DVDD.n5255 DVDD.n5250 4.5005
R10415 DVDD.n15423 DVDD.n5250 4.5005
R10416 DVDD.n5254 DVDD.n5250 4.5005
R10417 DVDD.n15459 DVDD.n5250 4.5005
R10418 DVDD.n15420 DVDD.n5232 4.5005
R10419 DVDD.n5256 DVDD.n5232 4.5005
R10420 DVDD.n15421 DVDD.n5232 4.5005
R10421 DVDD.n5255 DVDD.n5232 4.5005
R10422 DVDD.n15423 DVDD.n5232 4.5005
R10423 DVDD.n5254 DVDD.n5232 4.5005
R10424 DVDD.n15459 DVDD.n5232 4.5005
R10425 DVDD.n5257 DVDD.n5232 4.5005
R10426 DVDD.n15419 DVDD.n5232 4.5005
R10427 DVDD.n5258 DVDD.n5232 4.5005
R10428 DVDD.n15418 DVDD.n5232 4.5005
R10429 DVDD.n5259 DVDD.n5232 4.5005
R10430 DVDD.n15416 DVDD.n5232 4.5005
R10431 DVDD.n5260 DVDD.n5232 4.5005
R10432 DVDD.n15461 DVDD.n5232 4.5005
R10433 DVDD.n15420 DVDD.n5251 4.5005
R10434 DVDD.n5256 DVDD.n5251 4.5005
R10435 DVDD.n15421 DVDD.n5251 4.5005
R10436 DVDD.n5255 DVDD.n5251 4.5005
R10437 DVDD.n15423 DVDD.n5251 4.5005
R10438 DVDD.n5254 DVDD.n5251 4.5005
R10439 DVDD.n15459 DVDD.n5251 4.5005
R10440 DVDD.n5257 DVDD.n5251 4.5005
R10441 DVDD.n15419 DVDD.n5251 4.5005
R10442 DVDD.n5258 DVDD.n5251 4.5005
R10443 DVDD.n15418 DVDD.n5251 4.5005
R10444 DVDD.n5259 DVDD.n5251 4.5005
R10445 DVDD.n15416 DVDD.n5251 4.5005
R10446 DVDD.n5260 DVDD.n5251 4.5005
R10447 DVDD.n15461 DVDD.n5251 4.5005
R10448 DVDD.n15420 DVDD.n5231 4.5005
R10449 DVDD.n5256 DVDD.n5231 4.5005
R10450 DVDD.n15421 DVDD.n5231 4.5005
R10451 DVDD.n5255 DVDD.n5231 4.5005
R10452 DVDD.n15423 DVDD.n5231 4.5005
R10453 DVDD.n5254 DVDD.n5231 4.5005
R10454 DVDD.n15459 DVDD.n5231 4.5005
R10455 DVDD.n5257 DVDD.n5231 4.5005
R10456 DVDD.n15419 DVDD.n5231 4.5005
R10457 DVDD.n5258 DVDD.n5231 4.5005
R10458 DVDD.n15418 DVDD.n5231 4.5005
R10459 DVDD.n5259 DVDD.n5231 4.5005
R10460 DVDD.n15416 DVDD.n5231 4.5005
R10461 DVDD.n5260 DVDD.n5231 4.5005
R10462 DVDD.n15461 DVDD.n5231 4.5005
R10463 DVDD.n15461 DVDD.n5252 4.5005
R10464 DVDD.n5260 DVDD.n5252 4.5005
R10465 DVDD.n15416 DVDD.n5252 4.5005
R10466 DVDD.n5259 DVDD.n5252 4.5005
R10467 DVDD.n15418 DVDD.n5252 4.5005
R10468 DVDD.n5258 DVDD.n5252 4.5005
R10469 DVDD.n15419 DVDD.n5252 4.5005
R10470 DVDD.n5257 DVDD.n5252 4.5005
R10471 DVDD.n15420 DVDD.n5252 4.5005
R10472 DVDD.n5256 DVDD.n5252 4.5005
R10473 DVDD.n15421 DVDD.n5252 4.5005
R10474 DVDD.n5255 DVDD.n5252 4.5005
R10475 DVDD.n15423 DVDD.n5252 4.5005
R10476 DVDD.n5254 DVDD.n5252 4.5005
R10477 DVDD.n15459 DVDD.n5252 4.5005
R10478 DVDD.n15461 DVDD.n5230 4.5005
R10479 DVDD.n5260 DVDD.n5230 4.5005
R10480 DVDD.n15416 DVDD.n5230 4.5005
R10481 DVDD.n5259 DVDD.n5230 4.5005
R10482 DVDD.n15418 DVDD.n5230 4.5005
R10483 DVDD.n5258 DVDD.n5230 4.5005
R10484 DVDD.n15419 DVDD.n5230 4.5005
R10485 DVDD.n5257 DVDD.n5230 4.5005
R10486 DVDD.n15420 DVDD.n5230 4.5005
R10487 DVDD.n5256 DVDD.n5230 4.5005
R10488 DVDD.n15421 DVDD.n5230 4.5005
R10489 DVDD.n5255 DVDD.n5230 4.5005
R10490 DVDD.n15423 DVDD.n5230 4.5005
R10491 DVDD.n5254 DVDD.n5230 4.5005
R10492 DVDD.n15459 DVDD.n5230 4.5005
R10493 DVDD.n15461 DVDD.n15460 4.5005
R10494 DVDD.n15460 DVDD.n5260 4.5005
R10495 DVDD.n15460 DVDD.n15416 4.5005
R10496 DVDD.n15460 DVDD.n5259 4.5005
R10497 DVDD.n15460 DVDD.n15418 4.5005
R10498 DVDD.n15460 DVDD.n5258 4.5005
R10499 DVDD.n15460 DVDD.n15419 4.5005
R10500 DVDD.n15460 DVDD.n5257 4.5005
R10501 DVDD.n15460 DVDD.n15420 4.5005
R10502 DVDD.n15460 DVDD.n5256 4.5005
R10503 DVDD.n15460 DVDD.n15421 4.5005
R10504 DVDD.n15460 DVDD.n5255 4.5005
R10505 DVDD.n15460 DVDD.n15423 4.5005
R10506 DVDD.n15460 DVDD.n5254 4.5005
R10507 DVDD.n15460 DVDD.n15459 4.5005
R10508 DVDD.n15409 DVDD.n5377 4.5005
R10509 DVDD.n15409 DVDD.n5375 4.5005
R10510 DVDD.n15409 DVDD.n5378 4.5005
R10511 DVDD.n15409 DVDD.n5374 4.5005
R10512 DVDD.n15409 DVDD.n5379 4.5005
R10513 DVDD.n15409 DVDD.n5372 4.5005
R10514 DVDD.n15409 DVDD.n5380 4.5005
R10515 DVDD.n15409 DVDD.n5370 4.5005
R10516 DVDD.n15409 DVDD.n5381 4.5005
R10517 DVDD.n15409 DVDD.n5369 4.5005
R10518 DVDD.n15409 DVDD.n15408 4.5005
R10519 DVDD.n5395 DVDD.n5377 4.5005
R10520 DVDD.n5395 DVDD.n5375 4.5005
R10521 DVDD.n5395 DVDD.n5378 4.5005
R10522 DVDD.n5395 DVDD.n5374 4.5005
R10523 DVDD.n15317 DVDD.n5395 4.5005
R10524 DVDD.n5408 DVDD.n5395 4.5005
R10525 DVDD.n5395 DVDD.n5379 4.5005
R10526 DVDD.n5395 DVDD.n5372 4.5005
R10527 DVDD.n5395 DVDD.n5380 4.5005
R10528 DVDD.n5407 DVDD.n5395 4.5005
R10529 DVDD.n15406 DVDD.n5395 4.5005
R10530 DVDD.n5395 DVDD.n5370 4.5005
R10531 DVDD.n5395 DVDD.n5381 4.5005
R10532 DVDD.n5395 DVDD.n5369 4.5005
R10533 DVDD.n15408 DVDD.n5395 4.5005
R10534 DVDD.n5393 DVDD.n5377 4.5005
R10535 DVDD.n5393 DVDD.n5375 4.5005
R10536 DVDD.n5393 DVDD.n5378 4.5005
R10537 DVDD.n5393 DVDD.n5374 4.5005
R10538 DVDD.n15317 DVDD.n5393 4.5005
R10539 DVDD.n5408 DVDD.n5393 4.5005
R10540 DVDD.n5393 DVDD.n5379 4.5005
R10541 DVDD.n5393 DVDD.n5372 4.5005
R10542 DVDD.n5393 DVDD.n5380 4.5005
R10543 DVDD.n5407 DVDD.n5393 4.5005
R10544 DVDD.n15406 DVDD.n5393 4.5005
R10545 DVDD.n5393 DVDD.n5370 4.5005
R10546 DVDD.n5393 DVDD.n5381 4.5005
R10547 DVDD.n5393 DVDD.n5369 4.5005
R10548 DVDD.n15408 DVDD.n5393 4.5005
R10549 DVDD.n15408 DVDD.n5396 4.5005
R10550 DVDD.n5396 DVDD.n5369 4.5005
R10551 DVDD.n5396 DVDD.n5381 4.5005
R10552 DVDD.n5396 DVDD.n5370 4.5005
R10553 DVDD.n15406 DVDD.n5396 4.5005
R10554 DVDD.n5407 DVDD.n5396 4.5005
R10555 DVDD.n5396 DVDD.n5380 4.5005
R10556 DVDD.n5396 DVDD.n5372 4.5005
R10557 DVDD.n5396 DVDD.n5377 4.5005
R10558 DVDD.n5396 DVDD.n5375 4.5005
R10559 DVDD.n5396 DVDD.n5378 4.5005
R10560 DVDD.n5396 DVDD.n5374 4.5005
R10561 DVDD.n15317 DVDD.n5396 4.5005
R10562 DVDD.n5408 DVDD.n5396 4.5005
R10563 DVDD.n5396 DVDD.n5379 4.5005
R10564 DVDD.n15408 DVDD.n5392 4.5005
R10565 DVDD.n5392 DVDD.n5369 4.5005
R10566 DVDD.n5392 DVDD.n5381 4.5005
R10567 DVDD.n5392 DVDD.n5370 4.5005
R10568 DVDD.n15406 DVDD.n5392 4.5005
R10569 DVDD.n5407 DVDD.n5392 4.5005
R10570 DVDD.n5392 DVDD.n5380 4.5005
R10571 DVDD.n5392 DVDD.n5372 4.5005
R10572 DVDD.n5392 DVDD.n5377 4.5005
R10573 DVDD.n5392 DVDD.n5375 4.5005
R10574 DVDD.n5392 DVDD.n5378 4.5005
R10575 DVDD.n5392 DVDD.n5374 4.5005
R10576 DVDD.n15317 DVDD.n5392 4.5005
R10577 DVDD.n5408 DVDD.n5392 4.5005
R10578 DVDD.n5392 DVDD.n5379 4.5005
R10579 DVDD.n15408 DVDD.n5397 4.5005
R10580 DVDD.n5397 DVDD.n5369 4.5005
R10581 DVDD.n5397 DVDD.n5381 4.5005
R10582 DVDD.n5397 DVDD.n5370 4.5005
R10583 DVDD.n15406 DVDD.n5397 4.5005
R10584 DVDD.n5407 DVDD.n5397 4.5005
R10585 DVDD.n5397 DVDD.n5380 4.5005
R10586 DVDD.n5397 DVDD.n5372 4.5005
R10587 DVDD.n5397 DVDD.n5377 4.5005
R10588 DVDD.n5397 DVDD.n5375 4.5005
R10589 DVDD.n5397 DVDD.n5378 4.5005
R10590 DVDD.n5397 DVDD.n5374 4.5005
R10591 DVDD.n15317 DVDD.n5397 4.5005
R10592 DVDD.n5408 DVDD.n5397 4.5005
R10593 DVDD.n5397 DVDD.n5379 4.5005
R10594 DVDD.n15408 DVDD.n5391 4.5005
R10595 DVDD.n5391 DVDD.n5369 4.5005
R10596 DVDD.n5391 DVDD.n5381 4.5005
R10597 DVDD.n5391 DVDD.n5370 4.5005
R10598 DVDD.n15406 DVDD.n5391 4.5005
R10599 DVDD.n5407 DVDD.n5391 4.5005
R10600 DVDD.n5391 DVDD.n5380 4.5005
R10601 DVDD.n5391 DVDD.n5372 4.5005
R10602 DVDD.n5391 DVDD.n5377 4.5005
R10603 DVDD.n5391 DVDD.n5375 4.5005
R10604 DVDD.n5391 DVDD.n5378 4.5005
R10605 DVDD.n5391 DVDD.n5374 4.5005
R10606 DVDD.n15317 DVDD.n5391 4.5005
R10607 DVDD.n5408 DVDD.n5391 4.5005
R10608 DVDD.n5391 DVDD.n5379 4.5005
R10609 DVDD.n5398 DVDD.n5377 4.5005
R10610 DVDD.n5398 DVDD.n5375 4.5005
R10611 DVDD.n5398 DVDD.n5378 4.5005
R10612 DVDD.n5398 DVDD.n5374 4.5005
R10613 DVDD.n15317 DVDD.n5398 4.5005
R10614 DVDD.n5408 DVDD.n5398 4.5005
R10615 DVDD.n5398 DVDD.n5379 4.5005
R10616 DVDD.n5398 DVDD.n5372 4.5005
R10617 DVDD.n5398 DVDD.n5380 4.5005
R10618 DVDD.n5407 DVDD.n5398 4.5005
R10619 DVDD.n15406 DVDD.n5398 4.5005
R10620 DVDD.n5398 DVDD.n5370 4.5005
R10621 DVDD.n5398 DVDD.n5381 4.5005
R10622 DVDD.n5398 DVDD.n5369 4.5005
R10623 DVDD.n15408 DVDD.n5398 4.5005
R10624 DVDD.n5390 DVDD.n5377 4.5005
R10625 DVDD.n5390 DVDD.n5375 4.5005
R10626 DVDD.n5390 DVDD.n5378 4.5005
R10627 DVDD.n5390 DVDD.n5374 4.5005
R10628 DVDD.n15317 DVDD.n5390 4.5005
R10629 DVDD.n5408 DVDD.n5390 4.5005
R10630 DVDD.n5390 DVDD.n5379 4.5005
R10631 DVDD.n5390 DVDD.n5372 4.5005
R10632 DVDD.n5390 DVDD.n5380 4.5005
R10633 DVDD.n5407 DVDD.n5390 4.5005
R10634 DVDD.n15406 DVDD.n5390 4.5005
R10635 DVDD.n5390 DVDD.n5370 4.5005
R10636 DVDD.n5390 DVDD.n5381 4.5005
R10637 DVDD.n5390 DVDD.n5369 4.5005
R10638 DVDD.n15408 DVDD.n5390 4.5005
R10639 DVDD.n5399 DVDD.n5377 4.5005
R10640 DVDD.n5399 DVDD.n5375 4.5005
R10641 DVDD.n5399 DVDD.n5378 4.5005
R10642 DVDD.n5399 DVDD.n5374 4.5005
R10643 DVDD.n15317 DVDD.n5399 4.5005
R10644 DVDD.n5408 DVDD.n5399 4.5005
R10645 DVDD.n5399 DVDD.n5379 4.5005
R10646 DVDD.n5399 DVDD.n5372 4.5005
R10647 DVDD.n5399 DVDD.n5380 4.5005
R10648 DVDD.n5407 DVDD.n5399 4.5005
R10649 DVDD.n15406 DVDD.n5399 4.5005
R10650 DVDD.n5399 DVDD.n5370 4.5005
R10651 DVDD.n5399 DVDD.n5381 4.5005
R10652 DVDD.n5399 DVDD.n5369 4.5005
R10653 DVDD.n15408 DVDD.n5399 4.5005
R10654 DVDD.n15408 DVDD.n5389 4.5005
R10655 DVDD.n5389 DVDD.n5369 4.5005
R10656 DVDD.n5389 DVDD.n5381 4.5005
R10657 DVDD.n5389 DVDD.n5370 4.5005
R10658 DVDD.n15406 DVDD.n5389 4.5005
R10659 DVDD.n5407 DVDD.n5389 4.5005
R10660 DVDD.n5389 DVDD.n5380 4.5005
R10661 DVDD.n5389 DVDD.n5372 4.5005
R10662 DVDD.n5389 DVDD.n5377 4.5005
R10663 DVDD.n5389 DVDD.n5375 4.5005
R10664 DVDD.n5389 DVDD.n5378 4.5005
R10665 DVDD.n5389 DVDD.n5374 4.5005
R10666 DVDD.n15317 DVDD.n5389 4.5005
R10667 DVDD.n5408 DVDD.n5389 4.5005
R10668 DVDD.n5389 DVDD.n5379 4.5005
R10669 DVDD.n15408 DVDD.n5400 4.5005
R10670 DVDD.n5400 DVDD.n5369 4.5005
R10671 DVDD.n5400 DVDD.n5381 4.5005
R10672 DVDD.n5400 DVDD.n5370 4.5005
R10673 DVDD.n15406 DVDD.n5400 4.5005
R10674 DVDD.n5407 DVDD.n5400 4.5005
R10675 DVDD.n5400 DVDD.n5380 4.5005
R10676 DVDD.n5400 DVDD.n5372 4.5005
R10677 DVDD.n5400 DVDD.n5377 4.5005
R10678 DVDD.n5400 DVDD.n5375 4.5005
R10679 DVDD.n5400 DVDD.n5378 4.5005
R10680 DVDD.n5400 DVDD.n5374 4.5005
R10681 DVDD.n15317 DVDD.n5400 4.5005
R10682 DVDD.n5408 DVDD.n5400 4.5005
R10683 DVDD.n5400 DVDD.n5379 4.5005
R10684 DVDD.n15408 DVDD.n5388 4.5005
R10685 DVDD.n5388 DVDD.n5369 4.5005
R10686 DVDD.n5388 DVDD.n5381 4.5005
R10687 DVDD.n5388 DVDD.n5370 4.5005
R10688 DVDD.n15406 DVDD.n5388 4.5005
R10689 DVDD.n5407 DVDD.n5388 4.5005
R10690 DVDD.n5388 DVDD.n5380 4.5005
R10691 DVDD.n5388 DVDD.n5372 4.5005
R10692 DVDD.n5388 DVDD.n5377 4.5005
R10693 DVDD.n5388 DVDD.n5375 4.5005
R10694 DVDD.n5388 DVDD.n5378 4.5005
R10695 DVDD.n5388 DVDD.n5374 4.5005
R10696 DVDD.n15317 DVDD.n5388 4.5005
R10697 DVDD.n5408 DVDD.n5388 4.5005
R10698 DVDD.n5388 DVDD.n5379 4.5005
R10699 DVDD.n15408 DVDD.n5401 4.5005
R10700 DVDD.n5401 DVDD.n5369 4.5005
R10701 DVDD.n5401 DVDD.n5381 4.5005
R10702 DVDD.n5401 DVDD.n5370 4.5005
R10703 DVDD.n15406 DVDD.n5401 4.5005
R10704 DVDD.n5407 DVDD.n5401 4.5005
R10705 DVDD.n5401 DVDD.n5380 4.5005
R10706 DVDD.n5401 DVDD.n5372 4.5005
R10707 DVDD.n5401 DVDD.n5377 4.5005
R10708 DVDD.n5401 DVDD.n5375 4.5005
R10709 DVDD.n5401 DVDD.n5378 4.5005
R10710 DVDD.n5401 DVDD.n5374 4.5005
R10711 DVDD.n15317 DVDD.n5401 4.5005
R10712 DVDD.n5408 DVDD.n5401 4.5005
R10713 DVDD.n5401 DVDD.n5379 4.5005
R10714 DVDD.n5387 DVDD.n5377 4.5005
R10715 DVDD.n5387 DVDD.n5375 4.5005
R10716 DVDD.n5387 DVDD.n5378 4.5005
R10717 DVDD.n5387 DVDD.n5374 4.5005
R10718 DVDD.n15317 DVDD.n5387 4.5005
R10719 DVDD.n5408 DVDD.n5387 4.5005
R10720 DVDD.n5387 DVDD.n5379 4.5005
R10721 DVDD.n5387 DVDD.n5372 4.5005
R10722 DVDD.n5387 DVDD.n5380 4.5005
R10723 DVDD.n5407 DVDD.n5387 4.5005
R10724 DVDD.n15406 DVDD.n5387 4.5005
R10725 DVDD.n5387 DVDD.n5370 4.5005
R10726 DVDD.n5387 DVDD.n5381 4.5005
R10727 DVDD.n5387 DVDD.n5369 4.5005
R10728 DVDD.n15408 DVDD.n5387 4.5005
R10729 DVDD.n5402 DVDD.n5377 4.5005
R10730 DVDD.n5402 DVDD.n5375 4.5005
R10731 DVDD.n5402 DVDD.n5378 4.5005
R10732 DVDD.n5402 DVDD.n5374 4.5005
R10733 DVDD.n15317 DVDD.n5402 4.5005
R10734 DVDD.n5408 DVDD.n5402 4.5005
R10735 DVDD.n5402 DVDD.n5379 4.5005
R10736 DVDD.n5402 DVDD.n5372 4.5005
R10737 DVDD.n5402 DVDD.n5380 4.5005
R10738 DVDD.n5407 DVDD.n5402 4.5005
R10739 DVDD.n15406 DVDD.n5402 4.5005
R10740 DVDD.n5402 DVDD.n5370 4.5005
R10741 DVDD.n5402 DVDD.n5381 4.5005
R10742 DVDD.n5402 DVDD.n5369 4.5005
R10743 DVDD.n15408 DVDD.n5402 4.5005
R10744 DVDD.n5386 DVDD.n5377 4.5005
R10745 DVDD.n5386 DVDD.n5375 4.5005
R10746 DVDD.n5386 DVDD.n5378 4.5005
R10747 DVDD.n5386 DVDD.n5374 4.5005
R10748 DVDD.n15317 DVDD.n5386 4.5005
R10749 DVDD.n5408 DVDD.n5386 4.5005
R10750 DVDD.n5386 DVDD.n5379 4.5005
R10751 DVDD.n5386 DVDD.n5372 4.5005
R10752 DVDD.n5386 DVDD.n5380 4.5005
R10753 DVDD.n5407 DVDD.n5386 4.5005
R10754 DVDD.n15406 DVDD.n5386 4.5005
R10755 DVDD.n5386 DVDD.n5370 4.5005
R10756 DVDD.n5386 DVDD.n5381 4.5005
R10757 DVDD.n5386 DVDD.n5369 4.5005
R10758 DVDD.n15408 DVDD.n5386 4.5005
R10759 DVDD.n15408 DVDD.n5403 4.5005
R10760 DVDD.n5403 DVDD.n5369 4.5005
R10761 DVDD.n5403 DVDD.n5381 4.5005
R10762 DVDD.n5403 DVDD.n5370 4.5005
R10763 DVDD.n15406 DVDD.n5403 4.5005
R10764 DVDD.n5407 DVDD.n5403 4.5005
R10765 DVDD.n5403 DVDD.n5380 4.5005
R10766 DVDD.n5403 DVDD.n5372 4.5005
R10767 DVDD.n5403 DVDD.n5377 4.5005
R10768 DVDD.n5403 DVDD.n5375 4.5005
R10769 DVDD.n5403 DVDD.n5378 4.5005
R10770 DVDD.n5403 DVDD.n5374 4.5005
R10771 DVDD.n15317 DVDD.n5403 4.5005
R10772 DVDD.n5408 DVDD.n5403 4.5005
R10773 DVDD.n5403 DVDD.n5379 4.5005
R10774 DVDD.n15408 DVDD.n5385 4.5005
R10775 DVDD.n5385 DVDD.n5369 4.5005
R10776 DVDD.n5385 DVDD.n5381 4.5005
R10777 DVDD.n5385 DVDD.n5370 4.5005
R10778 DVDD.n15406 DVDD.n5385 4.5005
R10779 DVDD.n5407 DVDD.n5385 4.5005
R10780 DVDD.n5385 DVDD.n5380 4.5005
R10781 DVDD.n5385 DVDD.n5372 4.5005
R10782 DVDD.n5385 DVDD.n5377 4.5005
R10783 DVDD.n5385 DVDD.n5375 4.5005
R10784 DVDD.n5385 DVDD.n5378 4.5005
R10785 DVDD.n5385 DVDD.n5374 4.5005
R10786 DVDD.n15317 DVDD.n5385 4.5005
R10787 DVDD.n5408 DVDD.n5385 4.5005
R10788 DVDD.n5385 DVDD.n5379 4.5005
R10789 DVDD.n15408 DVDD.n5404 4.5005
R10790 DVDD.n5404 DVDD.n5369 4.5005
R10791 DVDD.n5404 DVDD.n5381 4.5005
R10792 DVDD.n5404 DVDD.n5370 4.5005
R10793 DVDD.n15406 DVDD.n5404 4.5005
R10794 DVDD.n5407 DVDD.n5404 4.5005
R10795 DVDD.n5404 DVDD.n5380 4.5005
R10796 DVDD.n5404 DVDD.n5372 4.5005
R10797 DVDD.n5404 DVDD.n5377 4.5005
R10798 DVDD.n5404 DVDD.n5375 4.5005
R10799 DVDD.n5404 DVDD.n5378 4.5005
R10800 DVDD.n5404 DVDD.n5374 4.5005
R10801 DVDD.n15317 DVDD.n5404 4.5005
R10802 DVDD.n5408 DVDD.n5404 4.5005
R10803 DVDD.n5404 DVDD.n5379 4.5005
R10804 DVDD.n5384 DVDD.n5377 4.5005
R10805 DVDD.n5384 DVDD.n5375 4.5005
R10806 DVDD.n5384 DVDD.n5378 4.5005
R10807 DVDD.n5384 DVDD.n5374 4.5005
R10808 DVDD.n15317 DVDD.n5384 4.5005
R10809 DVDD.n5408 DVDD.n5384 4.5005
R10810 DVDD.n5384 DVDD.n5379 4.5005
R10811 DVDD.n5384 DVDD.n5372 4.5005
R10812 DVDD.n5384 DVDD.n5380 4.5005
R10813 DVDD.n5407 DVDD.n5384 4.5005
R10814 DVDD.n15406 DVDD.n5384 4.5005
R10815 DVDD.n5384 DVDD.n5370 4.5005
R10816 DVDD.n5384 DVDD.n5381 4.5005
R10817 DVDD.n5384 DVDD.n5369 4.5005
R10818 DVDD.n15408 DVDD.n5384 4.5005
R10819 DVDD.n5405 DVDD.n5377 4.5005
R10820 DVDD.n5405 DVDD.n5375 4.5005
R10821 DVDD.n5405 DVDD.n5378 4.5005
R10822 DVDD.n5405 DVDD.n5374 4.5005
R10823 DVDD.n15317 DVDD.n5405 4.5005
R10824 DVDD.n5408 DVDD.n5405 4.5005
R10825 DVDD.n5405 DVDD.n5379 4.5005
R10826 DVDD.n5405 DVDD.n5372 4.5005
R10827 DVDD.n5405 DVDD.n5380 4.5005
R10828 DVDD.n5407 DVDD.n5405 4.5005
R10829 DVDD.n15406 DVDD.n5405 4.5005
R10830 DVDD.n5405 DVDD.n5370 4.5005
R10831 DVDD.n5405 DVDD.n5381 4.5005
R10832 DVDD.n5405 DVDD.n5369 4.5005
R10833 DVDD.n15408 DVDD.n5405 4.5005
R10834 DVDD.n5383 DVDD.n5377 4.5005
R10835 DVDD.n5383 DVDD.n5375 4.5005
R10836 DVDD.n5383 DVDD.n5378 4.5005
R10837 DVDD.n5383 DVDD.n5374 4.5005
R10838 DVDD.n15317 DVDD.n5383 4.5005
R10839 DVDD.n5408 DVDD.n5383 4.5005
R10840 DVDD.n5383 DVDD.n5379 4.5005
R10841 DVDD.n5383 DVDD.n5372 4.5005
R10842 DVDD.n5383 DVDD.n5380 4.5005
R10843 DVDD.n5407 DVDD.n5383 4.5005
R10844 DVDD.n15406 DVDD.n5383 4.5005
R10845 DVDD.n5383 DVDD.n5370 4.5005
R10846 DVDD.n5383 DVDD.n5381 4.5005
R10847 DVDD.n5383 DVDD.n5369 4.5005
R10848 DVDD.n15408 DVDD.n5383 4.5005
R10849 DVDD.n15407 DVDD.n5377 4.5005
R10850 DVDD.n15407 DVDD.n5375 4.5005
R10851 DVDD.n15407 DVDD.n5378 4.5005
R10852 DVDD.n15407 DVDD.n5374 4.5005
R10853 DVDD.n15407 DVDD.n15317 4.5005
R10854 DVDD.n15407 DVDD.n5408 4.5005
R10855 DVDD.n15407 DVDD.n5379 4.5005
R10856 DVDD.n15407 DVDD.n5372 4.5005
R10857 DVDD.n15407 DVDD.n5380 4.5005
R10858 DVDD.n15407 DVDD.n5407 4.5005
R10859 DVDD.n15407 DVDD.n15406 4.5005
R10860 DVDD.n15407 DVDD.n5370 4.5005
R10861 DVDD.n15407 DVDD.n5381 4.5005
R10862 DVDD.n15407 DVDD.n5369 4.5005
R10863 DVDD.n15408 DVDD.n15407 4.5005
R10864 DVDD.n5477 DVDD.n5468 4.5005
R10865 DVDD.n5475 DVDD.n5468 4.5005
R10866 DVDD.n5478 DVDD.n5468 4.5005
R10867 DVDD.n5474 DVDD.n5468 4.5005
R10868 DVDD.n5481 DVDD.n5468 4.5005
R10869 DVDD.n5472 DVDD.n5468 4.5005
R10870 DVDD.n5482 DVDD.n5468 4.5005
R10871 DVDD.n5471 DVDD.n5468 4.5005
R10872 DVDD.n5483 DVDD.n5468 4.5005
R10873 DVDD.n5470 DVDD.n5468 4.5005
R10874 DVDD.n15285 DVDD.n5468 4.5005
R10875 DVDD.n15286 DVDD.n5477 4.5005
R10876 DVDD.n15286 DVDD.n5475 4.5005
R10877 DVDD.n15286 DVDD.n5478 4.5005
R10878 DVDD.n15286 DVDD.n5474 4.5005
R10879 DVDD.n15286 DVDD.n5480 4.5005
R10880 DVDD.n15286 DVDD.n5473 4.5005
R10881 DVDD.n15286 DVDD.n5481 4.5005
R10882 DVDD.n15286 DVDD.n5472 4.5005
R10883 DVDD.n15286 DVDD.n5482 4.5005
R10884 DVDD.n15286 DVDD.n5471 4.5005
R10885 DVDD.n15286 DVDD.n5483 4.5005
R10886 DVDD.n15286 DVDD.n5470 4.5005
R10887 DVDD.n15286 DVDD.n5485 4.5005
R10888 DVDD.n15286 DVDD.n5469 4.5005
R10889 DVDD.n15286 DVDD.n15285 4.5005
R10890 DVDD.n5492 DVDD.n5477 4.5005
R10891 DVDD.n5492 DVDD.n5475 4.5005
R10892 DVDD.n5492 DVDD.n5478 4.5005
R10893 DVDD.n5492 DVDD.n5474 4.5005
R10894 DVDD.n5492 DVDD.n5480 4.5005
R10895 DVDD.n5492 DVDD.n5473 4.5005
R10896 DVDD.n5492 DVDD.n5481 4.5005
R10897 DVDD.n5492 DVDD.n5472 4.5005
R10898 DVDD.n5492 DVDD.n5482 4.5005
R10899 DVDD.n5492 DVDD.n5471 4.5005
R10900 DVDD.n5492 DVDD.n5483 4.5005
R10901 DVDD.n5492 DVDD.n5470 4.5005
R10902 DVDD.n5492 DVDD.n5485 4.5005
R10903 DVDD.n5492 DVDD.n5469 4.5005
R10904 DVDD.n15285 DVDD.n5492 4.5005
R10905 DVDD.n5490 DVDD.n5477 4.5005
R10906 DVDD.n5490 DVDD.n5475 4.5005
R10907 DVDD.n5490 DVDD.n5478 4.5005
R10908 DVDD.n5490 DVDD.n5474 4.5005
R10909 DVDD.n5490 DVDD.n5480 4.5005
R10910 DVDD.n5490 DVDD.n5473 4.5005
R10911 DVDD.n5490 DVDD.n5481 4.5005
R10912 DVDD.n5490 DVDD.n5472 4.5005
R10913 DVDD.n5490 DVDD.n5482 4.5005
R10914 DVDD.n5490 DVDD.n5471 4.5005
R10915 DVDD.n5490 DVDD.n5483 4.5005
R10916 DVDD.n5490 DVDD.n5470 4.5005
R10917 DVDD.n5490 DVDD.n5485 4.5005
R10918 DVDD.n5490 DVDD.n5469 4.5005
R10919 DVDD.n15285 DVDD.n5490 4.5005
R10920 DVDD.n5493 DVDD.n5482 4.5005
R10921 DVDD.n5493 DVDD.n5471 4.5005
R10922 DVDD.n5493 DVDD.n5483 4.5005
R10923 DVDD.n5493 DVDD.n5470 4.5005
R10924 DVDD.n5493 DVDD.n5485 4.5005
R10925 DVDD.n5493 DVDD.n5469 4.5005
R10926 DVDD.n15285 DVDD.n5493 4.5005
R10927 DVDD.n5493 DVDD.n5472 4.5005
R10928 DVDD.n5493 DVDD.n5481 4.5005
R10929 DVDD.n5493 DVDD.n5473 4.5005
R10930 DVDD.n5493 DVDD.n5480 4.5005
R10931 DVDD.n5493 DVDD.n5474 4.5005
R10932 DVDD.n5493 DVDD.n5478 4.5005
R10933 DVDD.n5493 DVDD.n5475 4.5005
R10934 DVDD.n5493 DVDD.n5477 4.5005
R10935 DVDD.n5489 DVDD.n5482 4.5005
R10936 DVDD.n5489 DVDD.n5471 4.5005
R10937 DVDD.n5489 DVDD.n5483 4.5005
R10938 DVDD.n5489 DVDD.n5470 4.5005
R10939 DVDD.n5489 DVDD.n5485 4.5005
R10940 DVDD.n5489 DVDD.n5469 4.5005
R10941 DVDD.n15285 DVDD.n5489 4.5005
R10942 DVDD.n5489 DVDD.n5472 4.5005
R10943 DVDD.n5489 DVDD.n5481 4.5005
R10944 DVDD.n5489 DVDD.n5473 4.5005
R10945 DVDD.n5489 DVDD.n5480 4.5005
R10946 DVDD.n5489 DVDD.n5474 4.5005
R10947 DVDD.n5489 DVDD.n5478 4.5005
R10948 DVDD.n5489 DVDD.n5475 4.5005
R10949 DVDD.n5489 DVDD.n5477 4.5005
R10950 DVDD.n5494 DVDD.n5482 4.5005
R10951 DVDD.n5494 DVDD.n5471 4.5005
R10952 DVDD.n5494 DVDD.n5483 4.5005
R10953 DVDD.n5494 DVDD.n5470 4.5005
R10954 DVDD.n5494 DVDD.n5485 4.5005
R10955 DVDD.n5494 DVDD.n5469 4.5005
R10956 DVDD.n15285 DVDD.n5494 4.5005
R10957 DVDD.n5494 DVDD.n5472 4.5005
R10958 DVDD.n5494 DVDD.n5481 4.5005
R10959 DVDD.n5494 DVDD.n5473 4.5005
R10960 DVDD.n5494 DVDD.n5480 4.5005
R10961 DVDD.n5494 DVDD.n5474 4.5005
R10962 DVDD.n5494 DVDD.n5478 4.5005
R10963 DVDD.n5494 DVDD.n5475 4.5005
R10964 DVDD.n5494 DVDD.n5477 4.5005
R10965 DVDD.n5488 DVDD.n5477 4.5005
R10966 DVDD.n5488 DVDD.n5475 4.5005
R10967 DVDD.n5488 DVDD.n5478 4.5005
R10968 DVDD.n5488 DVDD.n5474 4.5005
R10969 DVDD.n5488 DVDD.n5480 4.5005
R10970 DVDD.n5488 DVDD.n5473 4.5005
R10971 DVDD.n5488 DVDD.n5481 4.5005
R10972 DVDD.n5488 DVDD.n5472 4.5005
R10973 DVDD.n5488 DVDD.n5482 4.5005
R10974 DVDD.n5488 DVDD.n5471 4.5005
R10975 DVDD.n5488 DVDD.n5483 4.5005
R10976 DVDD.n5488 DVDD.n5470 4.5005
R10977 DVDD.n5488 DVDD.n5485 4.5005
R10978 DVDD.n5488 DVDD.n5469 4.5005
R10979 DVDD.n15285 DVDD.n5488 4.5005
R10980 DVDD.n5495 DVDD.n5477 4.5005
R10981 DVDD.n5495 DVDD.n5475 4.5005
R10982 DVDD.n5495 DVDD.n5478 4.5005
R10983 DVDD.n5495 DVDD.n5474 4.5005
R10984 DVDD.n5495 DVDD.n5480 4.5005
R10985 DVDD.n5495 DVDD.n5473 4.5005
R10986 DVDD.n5495 DVDD.n5481 4.5005
R10987 DVDD.n5495 DVDD.n5472 4.5005
R10988 DVDD.n5495 DVDD.n5482 4.5005
R10989 DVDD.n5495 DVDD.n5471 4.5005
R10990 DVDD.n5495 DVDD.n5483 4.5005
R10991 DVDD.n5495 DVDD.n5470 4.5005
R10992 DVDD.n5495 DVDD.n5485 4.5005
R10993 DVDD.n5495 DVDD.n5469 4.5005
R10994 DVDD.n15285 DVDD.n5495 4.5005
R10995 DVDD.n5487 DVDD.n5477 4.5005
R10996 DVDD.n5487 DVDD.n5475 4.5005
R10997 DVDD.n5487 DVDD.n5478 4.5005
R10998 DVDD.n5487 DVDD.n5474 4.5005
R10999 DVDD.n5487 DVDD.n5480 4.5005
R11000 DVDD.n5487 DVDD.n5473 4.5005
R11001 DVDD.n5487 DVDD.n5481 4.5005
R11002 DVDD.n5487 DVDD.n5472 4.5005
R11003 DVDD.n5487 DVDD.n5482 4.5005
R11004 DVDD.n5487 DVDD.n5471 4.5005
R11005 DVDD.n5487 DVDD.n5483 4.5005
R11006 DVDD.n5487 DVDD.n5470 4.5005
R11007 DVDD.n5487 DVDD.n5485 4.5005
R11008 DVDD.n5487 DVDD.n5469 4.5005
R11009 DVDD.n15285 DVDD.n5487 4.5005
R11010 DVDD.n15284 DVDD.n5482 4.5005
R11011 DVDD.n15284 DVDD.n5471 4.5005
R11012 DVDD.n15284 DVDD.n5483 4.5005
R11013 DVDD.n15284 DVDD.n5470 4.5005
R11014 DVDD.n15284 DVDD.n5485 4.5005
R11015 DVDD.n15284 DVDD.n5469 4.5005
R11016 DVDD.n15285 DVDD.n15284 4.5005
R11017 DVDD.n15284 DVDD.n5472 4.5005
R11018 DVDD.n15284 DVDD.n5481 4.5005
R11019 DVDD.n15284 DVDD.n5473 4.5005
R11020 DVDD.n15284 DVDD.n5480 4.5005
R11021 DVDD.n15284 DVDD.n5474 4.5005
R11022 DVDD.n15284 DVDD.n5478 4.5005
R11023 DVDD.n15284 DVDD.n5475 4.5005
R11024 DVDD.n15284 DVDD.n5477 4.5005
R11025 DVDD.n20609 DVDD.n19703 4.5005
R11026 DVDD.n20607 DVDD.n19703 4.5005
R11027 DVDD.n20612 DVDD.n19703 4.5005
R11028 DVDD.n20606 DVDD.n19703 4.5005
R11029 DVDD.n20613 DVDD.n19703 4.5005
R11030 DVDD.n20605 DVDD.n19703 4.5005
R11031 DVDD.n20614 DVDD.n19703 4.5005
R11032 DVDD.n20647 DVDD.n19703 4.5005
R11033 DVDD.n20655 DVDD.n19703 4.5005
R11034 DVDD.n20657 DVDD.n19703 4.5005
R11035 DVDD.n20609 DVDD.n19186 4.5005
R11036 DVDD.n20608 DVDD.n19186 4.5005
R11037 DVDD.n20611 DVDD.n19186 4.5005
R11038 DVDD.n20607 DVDD.n19186 4.5005
R11039 DVDD.n20612 DVDD.n19186 4.5005
R11040 DVDD.n20606 DVDD.n19186 4.5005
R11041 DVDD.n20613 DVDD.n19186 4.5005
R11042 DVDD.n20605 DVDD.n19186 4.5005
R11043 DVDD.n20614 DVDD.n19186 4.5005
R11044 DVDD.n20604 DVDD.n19186 4.5005
R11045 DVDD.n20616 DVDD.n19186 4.5005
R11046 DVDD.n20655 DVDD.n19186 4.5005
R11047 DVDD.n20657 DVDD.n19186 4.5005
R11048 DVDD.n20609 DVDD.n19704 4.5005
R11049 DVDD.n20608 DVDD.n19704 4.5005
R11050 DVDD.n20611 DVDD.n19704 4.5005
R11051 DVDD.n20607 DVDD.n19704 4.5005
R11052 DVDD.n20612 DVDD.n19704 4.5005
R11053 DVDD.n20606 DVDD.n19704 4.5005
R11054 DVDD.n20613 DVDD.n19704 4.5005
R11055 DVDD.n20605 DVDD.n19704 4.5005
R11056 DVDD.n20614 DVDD.n19704 4.5005
R11057 DVDD.n20604 DVDD.n19704 4.5005
R11058 DVDD.n20616 DVDD.n19704 4.5005
R11059 DVDD.n20655 DVDD.n19704 4.5005
R11060 DVDD.n20657 DVDD.n19704 4.5005
R11061 DVDD.n20609 DVDD.n19185 4.5005
R11062 DVDD.n20608 DVDD.n19185 4.5005
R11063 DVDD.n20611 DVDD.n19185 4.5005
R11064 DVDD.n20607 DVDD.n19185 4.5005
R11065 DVDD.n20612 DVDD.n19185 4.5005
R11066 DVDD.n20606 DVDD.n19185 4.5005
R11067 DVDD.n20613 DVDD.n19185 4.5005
R11068 DVDD.n20605 DVDD.n19185 4.5005
R11069 DVDD.n20614 DVDD.n19185 4.5005
R11070 DVDD.n20604 DVDD.n19185 4.5005
R11071 DVDD.n20616 DVDD.n19185 4.5005
R11072 DVDD.n20655 DVDD.n19185 4.5005
R11073 DVDD.n20657 DVDD.n19185 4.5005
R11074 DVDD.n20609 DVDD.n19705 4.5005
R11075 DVDD.n20608 DVDD.n19705 4.5005
R11076 DVDD.n20611 DVDD.n19705 4.5005
R11077 DVDD.n20607 DVDD.n19705 4.5005
R11078 DVDD.n20612 DVDD.n19705 4.5005
R11079 DVDD.n20606 DVDD.n19705 4.5005
R11080 DVDD.n20613 DVDD.n19705 4.5005
R11081 DVDD.n20605 DVDD.n19705 4.5005
R11082 DVDD.n20614 DVDD.n19705 4.5005
R11083 DVDD.n20604 DVDD.n19705 4.5005
R11084 DVDD.n20616 DVDD.n19705 4.5005
R11085 DVDD.n20655 DVDD.n19705 4.5005
R11086 DVDD.n20657 DVDD.n19705 4.5005
R11087 DVDD.n20609 DVDD.n19184 4.5005
R11088 DVDD.n20608 DVDD.n19184 4.5005
R11089 DVDD.n20611 DVDD.n19184 4.5005
R11090 DVDD.n20607 DVDD.n19184 4.5005
R11091 DVDD.n20612 DVDD.n19184 4.5005
R11092 DVDD.n20606 DVDD.n19184 4.5005
R11093 DVDD.n20613 DVDD.n19184 4.5005
R11094 DVDD.n20605 DVDD.n19184 4.5005
R11095 DVDD.n20614 DVDD.n19184 4.5005
R11096 DVDD.n20604 DVDD.n19184 4.5005
R11097 DVDD.n20616 DVDD.n19184 4.5005
R11098 DVDD.n20655 DVDD.n19184 4.5005
R11099 DVDD.n20657 DVDD.n19184 4.5005
R11100 DVDD.n20609 DVDD.n19706 4.5005
R11101 DVDD.n20608 DVDD.n19706 4.5005
R11102 DVDD.n20611 DVDD.n19706 4.5005
R11103 DVDD.n20607 DVDD.n19706 4.5005
R11104 DVDD.n20612 DVDD.n19706 4.5005
R11105 DVDD.n20606 DVDD.n19706 4.5005
R11106 DVDD.n20613 DVDD.n19706 4.5005
R11107 DVDD.n20605 DVDD.n19706 4.5005
R11108 DVDD.n20614 DVDD.n19706 4.5005
R11109 DVDD.n20604 DVDD.n19706 4.5005
R11110 DVDD.n20616 DVDD.n19706 4.5005
R11111 DVDD.n20655 DVDD.n19706 4.5005
R11112 DVDD.n20657 DVDD.n19706 4.5005
R11113 DVDD.n20609 DVDD.n19183 4.5005
R11114 DVDD.n20608 DVDD.n19183 4.5005
R11115 DVDD.n20611 DVDD.n19183 4.5005
R11116 DVDD.n20607 DVDD.n19183 4.5005
R11117 DVDD.n20612 DVDD.n19183 4.5005
R11118 DVDD.n20606 DVDD.n19183 4.5005
R11119 DVDD.n20613 DVDD.n19183 4.5005
R11120 DVDD.n20605 DVDD.n19183 4.5005
R11121 DVDD.n20614 DVDD.n19183 4.5005
R11122 DVDD.n20604 DVDD.n19183 4.5005
R11123 DVDD.n20616 DVDD.n19183 4.5005
R11124 DVDD.n20655 DVDD.n19183 4.5005
R11125 DVDD.n20657 DVDD.n19183 4.5005
R11126 DVDD.n20609 DVDD.n19707 4.5005
R11127 DVDD.n20608 DVDD.n19707 4.5005
R11128 DVDD.n20611 DVDD.n19707 4.5005
R11129 DVDD.n20607 DVDD.n19707 4.5005
R11130 DVDD.n20612 DVDD.n19707 4.5005
R11131 DVDD.n20606 DVDD.n19707 4.5005
R11132 DVDD.n20613 DVDD.n19707 4.5005
R11133 DVDD.n20605 DVDD.n19707 4.5005
R11134 DVDD.n20614 DVDD.n19707 4.5005
R11135 DVDD.n20604 DVDD.n19707 4.5005
R11136 DVDD.n20616 DVDD.n19707 4.5005
R11137 DVDD.n20655 DVDD.n19707 4.5005
R11138 DVDD.n20657 DVDD.n19707 4.5005
R11139 DVDD.n20609 DVDD.n19182 4.5005
R11140 DVDD.n20608 DVDD.n19182 4.5005
R11141 DVDD.n20611 DVDD.n19182 4.5005
R11142 DVDD.n20607 DVDD.n19182 4.5005
R11143 DVDD.n20612 DVDD.n19182 4.5005
R11144 DVDD.n20606 DVDD.n19182 4.5005
R11145 DVDD.n20613 DVDD.n19182 4.5005
R11146 DVDD.n20605 DVDD.n19182 4.5005
R11147 DVDD.n20614 DVDD.n19182 4.5005
R11148 DVDD.n20604 DVDD.n19182 4.5005
R11149 DVDD.n20616 DVDD.n19182 4.5005
R11150 DVDD.n20655 DVDD.n19182 4.5005
R11151 DVDD.n20657 DVDD.n19182 4.5005
R11152 DVDD.n20656 DVDD.n20609 4.5005
R11153 DVDD.n20656 DVDD.n20608 4.5005
R11154 DVDD.n20656 DVDD.n20611 4.5005
R11155 DVDD.n20656 DVDD.n20607 4.5005
R11156 DVDD.n20656 DVDD.n20612 4.5005
R11157 DVDD.n20656 DVDD.n20606 4.5005
R11158 DVDD.n20656 DVDD.n20613 4.5005
R11159 DVDD.n20656 DVDD.n20605 4.5005
R11160 DVDD.n20656 DVDD.n20614 4.5005
R11161 DVDD.n20656 DVDD.n20604 4.5005
R11162 DVDD.n20656 DVDD.n20616 4.5005
R11163 DVDD.n20656 DVDD.n20655 4.5005
R11164 DVDD.n20656 DVDD.n20602 4.5005
R11165 DVDD.n20657 DVDD.n20656 4.5005
R11166 DVDD.n20122 DVDD.n20065 4.5005
R11167 DVDD.n20076 DVDD.n20065 4.5005
R11168 DVDD.n20125 DVDD.n20065 4.5005
R11169 DVDD.n20075 DVDD.n20065 4.5005
R11170 DVDD.n20126 DVDD.n20065 4.5005
R11171 DVDD.n20074 DVDD.n20065 4.5005
R11172 DVDD.n20127 DVDD.n20065 4.5005
R11173 DVDD.n20072 DVDD.n20065 4.5005
R11174 DVDD.n20163 DVDD.n20065 4.5005
R11175 DVDD.n20071 DVDD.n20065 4.5005
R11176 DVDD.n20165 DVDD.n20065 4.5005
R11177 DVDD.n20122 DVDD.n20064 4.5005
R11178 DVDD.n20077 DVDD.n20064 4.5005
R11179 DVDD.n20124 DVDD.n20064 4.5005
R11180 DVDD.n20076 DVDD.n20064 4.5005
R11181 DVDD.n20125 DVDD.n20064 4.5005
R11182 DVDD.n20075 DVDD.n20064 4.5005
R11183 DVDD.n20126 DVDD.n20064 4.5005
R11184 DVDD.n20074 DVDD.n20064 4.5005
R11185 DVDD.n20127 DVDD.n20064 4.5005
R11186 DVDD.n20073 DVDD.n20064 4.5005
R11187 DVDD.n20129 DVDD.n20064 4.5005
R11188 DVDD.n20072 DVDD.n20064 4.5005
R11189 DVDD.n20163 DVDD.n20064 4.5005
R11190 DVDD.n20071 DVDD.n20064 4.5005
R11191 DVDD.n20165 DVDD.n20064 4.5005
R11192 DVDD.n20122 DVDD.n20066 4.5005
R11193 DVDD.n20077 DVDD.n20066 4.5005
R11194 DVDD.n20124 DVDD.n20066 4.5005
R11195 DVDD.n20076 DVDD.n20066 4.5005
R11196 DVDD.n20125 DVDD.n20066 4.5005
R11197 DVDD.n20075 DVDD.n20066 4.5005
R11198 DVDD.n20126 DVDD.n20066 4.5005
R11199 DVDD.n20074 DVDD.n20066 4.5005
R11200 DVDD.n20127 DVDD.n20066 4.5005
R11201 DVDD.n20073 DVDD.n20066 4.5005
R11202 DVDD.n20129 DVDD.n20066 4.5005
R11203 DVDD.n20072 DVDD.n20066 4.5005
R11204 DVDD.n20163 DVDD.n20066 4.5005
R11205 DVDD.n20071 DVDD.n20066 4.5005
R11206 DVDD.n20165 DVDD.n20066 4.5005
R11207 DVDD.n20122 DVDD.n20063 4.5005
R11208 DVDD.n20077 DVDD.n20063 4.5005
R11209 DVDD.n20124 DVDD.n20063 4.5005
R11210 DVDD.n20076 DVDD.n20063 4.5005
R11211 DVDD.n20125 DVDD.n20063 4.5005
R11212 DVDD.n20075 DVDD.n20063 4.5005
R11213 DVDD.n20126 DVDD.n20063 4.5005
R11214 DVDD.n20074 DVDD.n20063 4.5005
R11215 DVDD.n20127 DVDD.n20063 4.5005
R11216 DVDD.n20073 DVDD.n20063 4.5005
R11217 DVDD.n20129 DVDD.n20063 4.5005
R11218 DVDD.n20072 DVDD.n20063 4.5005
R11219 DVDD.n20163 DVDD.n20063 4.5005
R11220 DVDD.n20071 DVDD.n20063 4.5005
R11221 DVDD.n20165 DVDD.n20063 4.5005
R11222 DVDD.n20122 DVDD.n20067 4.5005
R11223 DVDD.n20077 DVDD.n20067 4.5005
R11224 DVDD.n20124 DVDD.n20067 4.5005
R11225 DVDD.n20076 DVDD.n20067 4.5005
R11226 DVDD.n20125 DVDD.n20067 4.5005
R11227 DVDD.n20075 DVDD.n20067 4.5005
R11228 DVDD.n20126 DVDD.n20067 4.5005
R11229 DVDD.n20074 DVDD.n20067 4.5005
R11230 DVDD.n20127 DVDD.n20067 4.5005
R11231 DVDD.n20073 DVDD.n20067 4.5005
R11232 DVDD.n20129 DVDD.n20067 4.5005
R11233 DVDD.n20072 DVDD.n20067 4.5005
R11234 DVDD.n20163 DVDD.n20067 4.5005
R11235 DVDD.n20071 DVDD.n20067 4.5005
R11236 DVDD.n20165 DVDD.n20067 4.5005
R11237 DVDD.n20122 DVDD.n20062 4.5005
R11238 DVDD.n20077 DVDD.n20062 4.5005
R11239 DVDD.n20124 DVDD.n20062 4.5005
R11240 DVDD.n20076 DVDD.n20062 4.5005
R11241 DVDD.n20125 DVDD.n20062 4.5005
R11242 DVDD.n20075 DVDD.n20062 4.5005
R11243 DVDD.n20126 DVDD.n20062 4.5005
R11244 DVDD.n20074 DVDD.n20062 4.5005
R11245 DVDD.n20127 DVDD.n20062 4.5005
R11246 DVDD.n20073 DVDD.n20062 4.5005
R11247 DVDD.n20129 DVDD.n20062 4.5005
R11248 DVDD.n20072 DVDD.n20062 4.5005
R11249 DVDD.n20163 DVDD.n20062 4.5005
R11250 DVDD.n20071 DVDD.n20062 4.5005
R11251 DVDD.n20165 DVDD.n20062 4.5005
R11252 DVDD.n20122 DVDD.n20068 4.5005
R11253 DVDD.n20077 DVDD.n20068 4.5005
R11254 DVDD.n20124 DVDD.n20068 4.5005
R11255 DVDD.n20076 DVDD.n20068 4.5005
R11256 DVDD.n20125 DVDD.n20068 4.5005
R11257 DVDD.n20075 DVDD.n20068 4.5005
R11258 DVDD.n20126 DVDD.n20068 4.5005
R11259 DVDD.n20074 DVDD.n20068 4.5005
R11260 DVDD.n20127 DVDD.n20068 4.5005
R11261 DVDD.n20073 DVDD.n20068 4.5005
R11262 DVDD.n20129 DVDD.n20068 4.5005
R11263 DVDD.n20072 DVDD.n20068 4.5005
R11264 DVDD.n20163 DVDD.n20068 4.5005
R11265 DVDD.n20071 DVDD.n20068 4.5005
R11266 DVDD.n20165 DVDD.n20068 4.5005
R11267 DVDD.n20122 DVDD.n20061 4.5005
R11268 DVDD.n20077 DVDD.n20061 4.5005
R11269 DVDD.n20124 DVDD.n20061 4.5005
R11270 DVDD.n20076 DVDD.n20061 4.5005
R11271 DVDD.n20125 DVDD.n20061 4.5005
R11272 DVDD.n20075 DVDD.n20061 4.5005
R11273 DVDD.n20126 DVDD.n20061 4.5005
R11274 DVDD.n20074 DVDD.n20061 4.5005
R11275 DVDD.n20127 DVDD.n20061 4.5005
R11276 DVDD.n20073 DVDD.n20061 4.5005
R11277 DVDD.n20129 DVDD.n20061 4.5005
R11278 DVDD.n20072 DVDD.n20061 4.5005
R11279 DVDD.n20163 DVDD.n20061 4.5005
R11280 DVDD.n20071 DVDD.n20061 4.5005
R11281 DVDD.n20165 DVDD.n20061 4.5005
R11282 DVDD.n20122 DVDD.n20069 4.5005
R11283 DVDD.n20077 DVDD.n20069 4.5005
R11284 DVDD.n20124 DVDD.n20069 4.5005
R11285 DVDD.n20076 DVDD.n20069 4.5005
R11286 DVDD.n20125 DVDD.n20069 4.5005
R11287 DVDD.n20075 DVDD.n20069 4.5005
R11288 DVDD.n20126 DVDD.n20069 4.5005
R11289 DVDD.n20074 DVDD.n20069 4.5005
R11290 DVDD.n20127 DVDD.n20069 4.5005
R11291 DVDD.n20073 DVDD.n20069 4.5005
R11292 DVDD.n20129 DVDD.n20069 4.5005
R11293 DVDD.n20072 DVDD.n20069 4.5005
R11294 DVDD.n20163 DVDD.n20069 4.5005
R11295 DVDD.n20071 DVDD.n20069 4.5005
R11296 DVDD.n20165 DVDD.n20069 4.5005
R11297 DVDD.n20122 DVDD.n20060 4.5005
R11298 DVDD.n20077 DVDD.n20060 4.5005
R11299 DVDD.n20124 DVDD.n20060 4.5005
R11300 DVDD.n20076 DVDD.n20060 4.5005
R11301 DVDD.n20125 DVDD.n20060 4.5005
R11302 DVDD.n20075 DVDD.n20060 4.5005
R11303 DVDD.n20126 DVDD.n20060 4.5005
R11304 DVDD.n20074 DVDD.n20060 4.5005
R11305 DVDD.n20127 DVDD.n20060 4.5005
R11306 DVDD.n20073 DVDD.n20060 4.5005
R11307 DVDD.n20129 DVDD.n20060 4.5005
R11308 DVDD.n20072 DVDD.n20060 4.5005
R11309 DVDD.n20163 DVDD.n20060 4.5005
R11310 DVDD.n20071 DVDD.n20060 4.5005
R11311 DVDD.n20165 DVDD.n20060 4.5005
R11312 DVDD.n20164 DVDD.n20122 4.5005
R11313 DVDD.n20164 DVDD.n20077 4.5005
R11314 DVDD.n20164 DVDD.n20124 4.5005
R11315 DVDD.n20164 DVDD.n20076 4.5005
R11316 DVDD.n20164 DVDD.n20125 4.5005
R11317 DVDD.n20164 DVDD.n20075 4.5005
R11318 DVDD.n20164 DVDD.n20126 4.5005
R11319 DVDD.n20164 DVDD.n20074 4.5005
R11320 DVDD.n20164 DVDD.n20127 4.5005
R11321 DVDD.n20164 DVDD.n20073 4.5005
R11322 DVDD.n20164 DVDD.n20129 4.5005
R11323 DVDD.n20164 DVDD.n20072 4.5005
R11324 DVDD.n20164 DVDD.n20163 4.5005
R11325 DVDD.n20164 DVDD.n20071 4.5005
R11326 DVDD.n20165 DVDD.n20164 4.5005
R11327 DVDD.n15143 DVDD.n5565 4.5005
R11328 DVDD.n15144 DVDD.n5568 4.5005
R11329 DVDD.n10222 DVDD.n10221 4.5005
R11330 DVDD.n10222 DVDD.n2291 4.5005
R11331 DVDD.n16429 DVDD.n2281 4.5005
R11332 DVDD.n16432 DVDD.n2281 4.5005
R11333 DVDD.n16451 DVDD.n2265 4.5005
R11334 DVDD.n16451 DVDD.n16450 4.5005
R11335 DVDD.n15146 DVDD.n5566 4.5005
R11336 DVDD.n10204 DVDD.n8960 4.5005
R11337 DVDD.n10221 DVDD.n8960 4.5005
R11338 DVDD.n8960 DVDD.n2291 4.5005
R11339 DVDD.n16406 DVDD.n2279 4.5005
R11340 DVDD.n16429 DVDD.n2279 4.5005
R11341 DVDD.n16432 DVDD.n2279 4.5005
R11342 DVDD.n16433 DVDD.n2267 4.5005
R11343 DVDD.n2267 DVDD.n2265 4.5005
R11344 DVDD.n16450 DVDD.n2267 4.5005
R11345 DVDD.n15147 DVDD.n5565 4.5005
R11346 DVDD.n15148 DVDD.n15147 4.5005
R11347 DVDD.n15147 DVDD.n15146 4.5005
R11348 DVDD.n5575 DVDD.n5563 4.5005
R11349 DVDD.n5574 DVDD.n5563 4.5005
R11350 DVDD.n5572 DVDD.n5563 4.5005
R11351 DVDD.n5570 DVDD.n5563 4.5005
R11352 DVDD.n5568 DVDD.n5563 4.5005
R11353 DVDD.n10219 DVDD.n10204 4.5005
R11354 DVDD.n10219 DVDD.n8970 4.5005
R11355 DVDD.n10219 DVDD.n10206 4.5005
R11356 DVDD.n10219 DVDD.n8969 4.5005
R11357 DVDD.n10219 DVDD.n10208 4.5005
R11358 DVDD.n10219 DVDD.n8968 4.5005
R11359 DVDD.n10219 DVDD.n10210 4.5005
R11360 DVDD.n10219 DVDD.n8967 4.5005
R11361 DVDD.n10219 DVDD.n10212 4.5005
R11362 DVDD.n10219 DVDD.n8966 4.5005
R11363 DVDD.n10219 DVDD.n10214 4.5005
R11364 DVDD.n10219 DVDD.n8965 4.5005
R11365 DVDD.n10219 DVDD.n10216 4.5005
R11366 DVDD.n10219 DVDD.n8964 4.5005
R11367 DVDD.n10219 DVDD.n10218 4.5005
R11368 DVDD.n10219 DVDD.n2291 4.5005
R11369 DVDD.n16431 DVDD.n16406 4.5005
R11370 DVDD.n16431 DVDD.n2290 4.5005
R11371 DVDD.n16431 DVDD.n16409 4.5005
R11372 DVDD.n16431 DVDD.n2289 4.5005
R11373 DVDD.n16431 DVDD.n16412 4.5005
R11374 DVDD.n16431 DVDD.n2288 4.5005
R11375 DVDD.n16431 DVDD.n16415 4.5005
R11376 DVDD.n16431 DVDD.n2287 4.5005
R11377 DVDD.n16431 DVDD.n16418 4.5005
R11378 DVDD.n16431 DVDD.n2286 4.5005
R11379 DVDD.n16431 DVDD.n16421 4.5005
R11380 DVDD.n16431 DVDD.n2285 4.5005
R11381 DVDD.n16431 DVDD.n16424 4.5005
R11382 DVDD.n16431 DVDD.n2284 4.5005
R11383 DVDD.n16431 DVDD.n16426 4.5005
R11384 DVDD.n16432 DVDD.n16431 4.5005
R11385 DVDD.n16449 DVDD.n16433 4.5005
R11386 DVDD.n16449 DVDD.n2277 4.5005
R11387 DVDD.n16449 DVDD.n16435 4.5005
R11388 DVDD.n16449 DVDD.n2276 4.5005
R11389 DVDD.n16449 DVDD.n16437 4.5005
R11390 DVDD.n16449 DVDD.n2275 4.5005
R11391 DVDD.n16449 DVDD.n16439 4.5005
R11392 DVDD.n16449 DVDD.n2274 4.5005
R11393 DVDD.n16449 DVDD.n16441 4.5005
R11394 DVDD.n16449 DVDD.n2273 4.5005
R11395 DVDD.n16449 DVDD.n16443 4.5005
R11396 DVDD.n16449 DVDD.n2272 4.5005
R11397 DVDD.n16449 DVDD.n16445 4.5005
R11398 DVDD.n16449 DVDD.n2271 4.5005
R11399 DVDD.n16449 DVDD.n16447 4.5005
R11400 DVDD.n16450 DVDD.n16449 4.5005
R11401 DVDD.n15145 DVDD.n5563 4.5005
R11402 DVDD.n15145 DVDD.n15144 4.5005
R11403 DVDD.n17734 DVDD.n888 4.5005
R11404 DVDD.n17734 DVDD.n17733 4.5005
R11405 DVDD.n17731 DVDD.n17730 4.5005
R11406 DVDD.n888 DVDD.n884 4.5005
R11407 DVDD.n886 DVDD.n885 4.5005
R11408 DVDD.n17737 DVDD.n879 4.5005
R11409 DVDD.n17737 DVDD.n882 4.5005
R11410 DVDD.n17737 DVDD.n878 4.5005
R11411 DVDD.n885 DVDD.n880 4.5005
R11412 DVDD.n17728 DVDD.n880 4.5005
R11413 DVDD.n17730 DVDD.n880 4.5005
R11414 DVDD.n18027 DVDD.n550 4.5005
R11415 DVDD.n18035 DVDD.n18034 4.5005
R11416 DVDD.n546 DVDD.n544 4.5005
R11417 DVDD.n550 DVDD.n543 4.5005
R11418 DVDD.n18025 DVDD.n543 4.5005
R11419 DVDD.n18024 DVDD.n543 4.5005
R11420 DVDD.n18028 DVDD.n543 4.5005
R11421 DVDD.n18030 DVDD.n543 4.5005
R11422 DVDD.n18036 DVDD.n544 4.5005
R11423 DVDD.n18036 DVDD.n542 4.5005
R11424 DVDD.n18036 DVDD.n18035 4.5005
R11425 DVDD.n17736 DVDD.n884 4.5005
R11426 DVDD.n17737 DVDD.n17736 4.5005
R11427 DVDD.n18027 DVDD.n549 4.5005
R11428 DVDD.n549 DVDD.n543 4.5005
R11429 DVDD.n17877 DVDD.n808 4.5005
R11430 DVDD.n808 DVDD.n785 4.5005
R11431 DVDD.n808 DVDD.n799 4.5005
R11432 DVDD.n808 DVDD.n786 4.5005
R11433 DVDD.n808 DVDD.n797 4.5005
R11434 DVDD.n808 DVDD.n788 4.5005
R11435 DVDD.n808 DVDD.n793 4.5005
R11436 DVDD.n808 DVDD.n791 4.5005
R11437 DVDD.n808 DVDD.n794 4.5005
R11438 DVDD.n808 DVDD.n790 4.5005
R11439 DVDD.n808 DVDD.n796 4.5005
R11440 DVDD.n17876 DVDD.n793 4.5005
R11441 DVDD.n17876 DVDD.n791 4.5005
R11442 DVDD.n17876 DVDD.n794 4.5005
R11443 DVDD.n17876 DVDD.n790 4.5005
R11444 DVDD.n17876 DVDD.n795 4.5005
R11445 DVDD.n17876 DVDD.n789 4.5005
R11446 DVDD.n17876 DVDD.n796 4.5005
R11447 DVDD.n801 DVDD.n793 4.5005
R11448 DVDD.n801 DVDD.n791 4.5005
R11449 DVDD.n801 DVDD.n794 4.5005
R11450 DVDD.n801 DVDD.n790 4.5005
R11451 DVDD.n801 DVDD.n795 4.5005
R11452 DVDD.n801 DVDD.n789 4.5005
R11453 DVDD.n801 DVDD.n796 4.5005
R11454 DVDD.n812 DVDD.n793 4.5005
R11455 DVDD.n812 DVDD.n791 4.5005
R11456 DVDD.n812 DVDD.n794 4.5005
R11457 DVDD.n812 DVDD.n790 4.5005
R11458 DVDD.n812 DVDD.n795 4.5005
R11459 DVDD.n812 DVDD.n789 4.5005
R11460 DVDD.n812 DVDD.n796 4.5005
R11461 DVDD.n17877 DVDD.n804 4.5005
R11462 DVDD.n804 DVDD.n785 4.5005
R11463 DVDD.n804 DVDD.n799 4.5005
R11464 DVDD.n804 DVDD.n786 4.5005
R11465 DVDD.n804 DVDD.n798 4.5005
R11466 DVDD.n804 DVDD.n787 4.5005
R11467 DVDD.n804 DVDD.n797 4.5005
R11468 DVDD.n804 DVDD.n788 4.5005
R11469 DVDD.n804 DVDD.n793 4.5005
R11470 DVDD.n804 DVDD.n791 4.5005
R11471 DVDD.n804 DVDD.n794 4.5005
R11472 DVDD.n804 DVDD.n790 4.5005
R11473 DVDD.n804 DVDD.n795 4.5005
R11474 DVDD.n804 DVDD.n789 4.5005
R11475 DVDD.n804 DVDD.n796 4.5005
R11476 DVDD.n17877 DVDD.n809 4.5005
R11477 DVDD.n809 DVDD.n785 4.5005
R11478 DVDD.n809 DVDD.n799 4.5005
R11479 DVDD.n809 DVDD.n786 4.5005
R11480 DVDD.n809 DVDD.n798 4.5005
R11481 DVDD.n809 DVDD.n787 4.5005
R11482 DVDD.n809 DVDD.n797 4.5005
R11483 DVDD.n809 DVDD.n788 4.5005
R11484 DVDD.n809 DVDD.n793 4.5005
R11485 DVDD.n809 DVDD.n791 4.5005
R11486 DVDD.n809 DVDD.n794 4.5005
R11487 DVDD.n809 DVDD.n790 4.5005
R11488 DVDD.n809 DVDD.n795 4.5005
R11489 DVDD.n809 DVDD.n789 4.5005
R11490 DVDD.n809 DVDD.n796 4.5005
R11491 DVDD.n17877 DVDD.n803 4.5005
R11492 DVDD.n803 DVDD.n785 4.5005
R11493 DVDD.n803 DVDD.n799 4.5005
R11494 DVDD.n803 DVDD.n786 4.5005
R11495 DVDD.n803 DVDD.n798 4.5005
R11496 DVDD.n803 DVDD.n787 4.5005
R11497 DVDD.n803 DVDD.n797 4.5005
R11498 DVDD.n803 DVDD.n788 4.5005
R11499 DVDD.n803 DVDD.n793 4.5005
R11500 DVDD.n803 DVDD.n791 4.5005
R11501 DVDD.n803 DVDD.n794 4.5005
R11502 DVDD.n803 DVDD.n790 4.5005
R11503 DVDD.n803 DVDD.n795 4.5005
R11504 DVDD.n803 DVDD.n789 4.5005
R11505 DVDD.n803 DVDD.n796 4.5005
R11506 DVDD.n17877 DVDD.n810 4.5005
R11507 DVDD.n810 DVDD.n785 4.5005
R11508 DVDD.n810 DVDD.n799 4.5005
R11509 DVDD.n810 DVDD.n786 4.5005
R11510 DVDD.n810 DVDD.n798 4.5005
R11511 DVDD.n810 DVDD.n787 4.5005
R11512 DVDD.n810 DVDD.n797 4.5005
R11513 DVDD.n810 DVDD.n788 4.5005
R11514 DVDD.n810 DVDD.n793 4.5005
R11515 DVDD.n810 DVDD.n791 4.5005
R11516 DVDD.n810 DVDD.n794 4.5005
R11517 DVDD.n810 DVDD.n790 4.5005
R11518 DVDD.n810 DVDD.n795 4.5005
R11519 DVDD.n810 DVDD.n789 4.5005
R11520 DVDD.n810 DVDD.n796 4.5005
R11521 DVDD.n802 DVDD.n793 4.5005
R11522 DVDD.n802 DVDD.n791 4.5005
R11523 DVDD.n802 DVDD.n794 4.5005
R11524 DVDD.n802 DVDD.n790 4.5005
R11525 DVDD.n802 DVDD.n795 4.5005
R11526 DVDD.n802 DVDD.n789 4.5005
R11527 DVDD.n802 DVDD.n796 4.5005
R11528 DVDD.n811 DVDD.n793 4.5005
R11529 DVDD.n811 DVDD.n791 4.5005
R11530 DVDD.n811 DVDD.n794 4.5005
R11531 DVDD.n811 DVDD.n790 4.5005
R11532 DVDD.n811 DVDD.n795 4.5005
R11533 DVDD.n811 DVDD.n789 4.5005
R11534 DVDD.n811 DVDD.n796 4.5005
R11535 DVDD.n17878 DVDD.n793 4.5005
R11536 DVDD.n17878 DVDD.n791 4.5005
R11537 DVDD.n17878 DVDD.n794 4.5005
R11538 DVDD.n17878 DVDD.n790 4.5005
R11539 DVDD.n17878 DVDD.n795 4.5005
R11540 DVDD.n17878 DVDD.n789 4.5005
R11541 DVDD.n17878 DVDD.n796 4.5005
R11542 DVDD.n760 DVDD.n739 4.5005
R11543 DVDD.n760 DVDD.n737 4.5005
R11544 DVDD.n760 DVDD.n740 4.5005
R11545 DVDD.n760 DVDD.n736 4.5005
R11546 DVDD.n760 DVDD.n742 4.5005
R11547 DVDD.n760 DVDD.n734 4.5005
R11548 DVDD.n760 DVDD.n743 4.5005
R11549 DVDD.n760 DVDD.n733 4.5005
R11550 DVDD.n760 DVDD.n744 4.5005
R11551 DVDD.n760 DVDD.n732 4.5005
R11552 DVDD.n17954 DVDD.n760 4.5005
R11553 DVDD.n762 DVDD.n739 4.5005
R11554 DVDD.n762 DVDD.n737 4.5005
R11555 DVDD.n762 DVDD.n740 4.5005
R11556 DVDD.n762 DVDD.n736 4.5005
R11557 DVDD.n762 DVDD.n741 4.5005
R11558 DVDD.n762 DVDD.n735 4.5005
R11559 DVDD.n762 DVDD.n742 4.5005
R11560 DVDD.n762 DVDD.n734 4.5005
R11561 DVDD.n762 DVDD.n743 4.5005
R11562 DVDD.n762 DVDD.n733 4.5005
R11563 DVDD.n762 DVDD.n744 4.5005
R11564 DVDD.n762 DVDD.n732 4.5005
R11565 DVDD.n762 DVDD.n745 4.5005
R11566 DVDD.n762 DVDD.n731 4.5005
R11567 DVDD.n17954 DVDD.n762 4.5005
R11568 DVDD.n757 DVDD.n739 4.5005
R11569 DVDD.n757 DVDD.n737 4.5005
R11570 DVDD.n757 DVDD.n740 4.5005
R11571 DVDD.n757 DVDD.n736 4.5005
R11572 DVDD.n757 DVDD.n741 4.5005
R11573 DVDD.n757 DVDD.n735 4.5005
R11574 DVDD.n757 DVDD.n742 4.5005
R11575 DVDD.n757 DVDD.n734 4.5005
R11576 DVDD.n757 DVDD.n743 4.5005
R11577 DVDD.n757 DVDD.n733 4.5005
R11578 DVDD.n757 DVDD.n744 4.5005
R11579 DVDD.n757 DVDD.n732 4.5005
R11580 DVDD.n757 DVDD.n745 4.5005
R11581 DVDD.n757 DVDD.n731 4.5005
R11582 DVDD.n17954 DVDD.n757 4.5005
R11583 DVDD.n763 DVDD.n739 4.5005
R11584 DVDD.n763 DVDD.n737 4.5005
R11585 DVDD.n763 DVDD.n740 4.5005
R11586 DVDD.n763 DVDD.n736 4.5005
R11587 DVDD.n763 DVDD.n741 4.5005
R11588 DVDD.n763 DVDD.n735 4.5005
R11589 DVDD.n763 DVDD.n742 4.5005
R11590 DVDD.n763 DVDD.n734 4.5005
R11591 DVDD.n763 DVDD.n743 4.5005
R11592 DVDD.n763 DVDD.n733 4.5005
R11593 DVDD.n763 DVDD.n744 4.5005
R11594 DVDD.n763 DVDD.n732 4.5005
R11595 DVDD.n763 DVDD.n745 4.5005
R11596 DVDD.n763 DVDD.n731 4.5005
R11597 DVDD.n17954 DVDD.n763 4.5005
R11598 DVDD.n756 DVDD.n743 4.5005
R11599 DVDD.n756 DVDD.n733 4.5005
R11600 DVDD.n756 DVDD.n744 4.5005
R11601 DVDD.n756 DVDD.n732 4.5005
R11602 DVDD.n756 DVDD.n745 4.5005
R11603 DVDD.n756 DVDD.n731 4.5005
R11604 DVDD.n17954 DVDD.n756 4.5005
R11605 DVDD.n764 DVDD.n743 4.5005
R11606 DVDD.n764 DVDD.n733 4.5005
R11607 DVDD.n764 DVDD.n744 4.5005
R11608 DVDD.n764 DVDD.n732 4.5005
R11609 DVDD.n764 DVDD.n745 4.5005
R11610 DVDD.n764 DVDD.n731 4.5005
R11611 DVDD.n17954 DVDD.n764 4.5005
R11612 DVDD.n755 DVDD.n743 4.5005
R11613 DVDD.n755 DVDD.n733 4.5005
R11614 DVDD.n755 DVDD.n744 4.5005
R11615 DVDD.n755 DVDD.n732 4.5005
R11616 DVDD.n755 DVDD.n745 4.5005
R11617 DVDD.n755 DVDD.n731 4.5005
R11618 DVDD.n17954 DVDD.n755 4.5005
R11619 DVDD.n765 DVDD.n739 4.5005
R11620 DVDD.n765 DVDD.n737 4.5005
R11621 DVDD.n765 DVDD.n740 4.5005
R11622 DVDD.n765 DVDD.n736 4.5005
R11623 DVDD.n765 DVDD.n741 4.5005
R11624 DVDD.n765 DVDD.n735 4.5005
R11625 DVDD.n765 DVDD.n742 4.5005
R11626 DVDD.n765 DVDD.n734 4.5005
R11627 DVDD.n765 DVDD.n743 4.5005
R11628 DVDD.n765 DVDD.n733 4.5005
R11629 DVDD.n765 DVDD.n744 4.5005
R11630 DVDD.n765 DVDD.n732 4.5005
R11631 DVDD.n765 DVDD.n745 4.5005
R11632 DVDD.n765 DVDD.n731 4.5005
R11633 DVDD.n17954 DVDD.n765 4.5005
R11634 DVDD.n754 DVDD.n739 4.5005
R11635 DVDD.n754 DVDD.n737 4.5005
R11636 DVDD.n754 DVDD.n740 4.5005
R11637 DVDD.n754 DVDD.n736 4.5005
R11638 DVDD.n754 DVDD.n741 4.5005
R11639 DVDD.n754 DVDD.n735 4.5005
R11640 DVDD.n754 DVDD.n742 4.5005
R11641 DVDD.n754 DVDD.n734 4.5005
R11642 DVDD.n754 DVDD.n743 4.5005
R11643 DVDD.n754 DVDD.n733 4.5005
R11644 DVDD.n754 DVDD.n744 4.5005
R11645 DVDD.n754 DVDD.n732 4.5005
R11646 DVDD.n754 DVDD.n745 4.5005
R11647 DVDD.n754 DVDD.n731 4.5005
R11648 DVDD.n17954 DVDD.n754 4.5005
R11649 DVDD.n766 DVDD.n739 4.5005
R11650 DVDD.n766 DVDD.n737 4.5005
R11651 DVDD.n766 DVDD.n740 4.5005
R11652 DVDD.n766 DVDD.n736 4.5005
R11653 DVDD.n766 DVDD.n741 4.5005
R11654 DVDD.n766 DVDD.n735 4.5005
R11655 DVDD.n766 DVDD.n742 4.5005
R11656 DVDD.n766 DVDD.n734 4.5005
R11657 DVDD.n766 DVDD.n743 4.5005
R11658 DVDD.n766 DVDD.n733 4.5005
R11659 DVDD.n766 DVDD.n744 4.5005
R11660 DVDD.n766 DVDD.n732 4.5005
R11661 DVDD.n766 DVDD.n745 4.5005
R11662 DVDD.n766 DVDD.n731 4.5005
R11663 DVDD.n17954 DVDD.n766 4.5005
R11664 DVDD.n753 DVDD.n739 4.5005
R11665 DVDD.n753 DVDD.n737 4.5005
R11666 DVDD.n753 DVDD.n740 4.5005
R11667 DVDD.n753 DVDD.n736 4.5005
R11668 DVDD.n753 DVDD.n741 4.5005
R11669 DVDD.n753 DVDD.n735 4.5005
R11670 DVDD.n753 DVDD.n742 4.5005
R11671 DVDD.n753 DVDD.n734 4.5005
R11672 DVDD.n753 DVDD.n743 4.5005
R11673 DVDD.n753 DVDD.n733 4.5005
R11674 DVDD.n753 DVDD.n744 4.5005
R11675 DVDD.n753 DVDD.n732 4.5005
R11676 DVDD.n753 DVDD.n745 4.5005
R11677 DVDD.n753 DVDD.n731 4.5005
R11678 DVDD.n17954 DVDD.n753 4.5005
R11679 DVDD.n767 DVDD.n743 4.5005
R11680 DVDD.n767 DVDD.n733 4.5005
R11681 DVDD.n767 DVDD.n744 4.5005
R11682 DVDD.n767 DVDD.n732 4.5005
R11683 DVDD.n767 DVDD.n745 4.5005
R11684 DVDD.n767 DVDD.n731 4.5005
R11685 DVDD.n17954 DVDD.n767 4.5005
R11686 DVDD.n752 DVDD.n743 4.5005
R11687 DVDD.n752 DVDD.n733 4.5005
R11688 DVDD.n752 DVDD.n744 4.5005
R11689 DVDD.n752 DVDD.n732 4.5005
R11690 DVDD.n752 DVDD.n745 4.5005
R11691 DVDD.n752 DVDD.n731 4.5005
R11692 DVDD.n17954 DVDD.n752 4.5005
R11693 DVDD.n768 DVDD.n743 4.5005
R11694 DVDD.n768 DVDD.n733 4.5005
R11695 DVDD.n768 DVDD.n744 4.5005
R11696 DVDD.n768 DVDD.n732 4.5005
R11697 DVDD.n768 DVDD.n745 4.5005
R11698 DVDD.n768 DVDD.n731 4.5005
R11699 DVDD.n17954 DVDD.n768 4.5005
R11700 DVDD.n751 DVDD.n739 4.5005
R11701 DVDD.n751 DVDD.n737 4.5005
R11702 DVDD.n751 DVDD.n740 4.5005
R11703 DVDD.n751 DVDD.n736 4.5005
R11704 DVDD.n751 DVDD.n741 4.5005
R11705 DVDD.n751 DVDD.n735 4.5005
R11706 DVDD.n751 DVDD.n742 4.5005
R11707 DVDD.n751 DVDD.n734 4.5005
R11708 DVDD.n751 DVDD.n743 4.5005
R11709 DVDD.n751 DVDD.n733 4.5005
R11710 DVDD.n751 DVDD.n744 4.5005
R11711 DVDD.n751 DVDD.n732 4.5005
R11712 DVDD.n751 DVDD.n745 4.5005
R11713 DVDD.n751 DVDD.n731 4.5005
R11714 DVDD.n17954 DVDD.n751 4.5005
R11715 DVDD.n769 DVDD.n739 4.5005
R11716 DVDD.n769 DVDD.n737 4.5005
R11717 DVDD.n769 DVDD.n740 4.5005
R11718 DVDD.n769 DVDD.n736 4.5005
R11719 DVDD.n769 DVDD.n741 4.5005
R11720 DVDD.n769 DVDD.n735 4.5005
R11721 DVDD.n769 DVDD.n742 4.5005
R11722 DVDD.n769 DVDD.n734 4.5005
R11723 DVDD.n769 DVDD.n743 4.5005
R11724 DVDD.n769 DVDD.n733 4.5005
R11725 DVDD.n769 DVDD.n744 4.5005
R11726 DVDD.n769 DVDD.n732 4.5005
R11727 DVDD.n769 DVDD.n745 4.5005
R11728 DVDD.n769 DVDD.n731 4.5005
R11729 DVDD.n17954 DVDD.n769 4.5005
R11730 DVDD.n750 DVDD.n739 4.5005
R11731 DVDD.n750 DVDD.n737 4.5005
R11732 DVDD.n750 DVDD.n740 4.5005
R11733 DVDD.n750 DVDD.n736 4.5005
R11734 DVDD.n750 DVDD.n741 4.5005
R11735 DVDD.n750 DVDD.n735 4.5005
R11736 DVDD.n750 DVDD.n742 4.5005
R11737 DVDD.n750 DVDD.n734 4.5005
R11738 DVDD.n750 DVDD.n743 4.5005
R11739 DVDD.n750 DVDD.n733 4.5005
R11740 DVDD.n750 DVDD.n744 4.5005
R11741 DVDD.n750 DVDD.n732 4.5005
R11742 DVDD.n750 DVDD.n745 4.5005
R11743 DVDD.n750 DVDD.n731 4.5005
R11744 DVDD.n17954 DVDD.n750 4.5005
R11745 DVDD.n770 DVDD.n743 4.5005
R11746 DVDD.n770 DVDD.n733 4.5005
R11747 DVDD.n770 DVDD.n744 4.5005
R11748 DVDD.n770 DVDD.n732 4.5005
R11749 DVDD.n770 DVDD.n745 4.5005
R11750 DVDD.n770 DVDD.n731 4.5005
R11751 DVDD.n17954 DVDD.n770 4.5005
R11752 DVDD.n749 DVDD.n743 4.5005
R11753 DVDD.n749 DVDD.n733 4.5005
R11754 DVDD.n749 DVDD.n744 4.5005
R11755 DVDD.n749 DVDD.n732 4.5005
R11756 DVDD.n749 DVDD.n745 4.5005
R11757 DVDD.n749 DVDD.n731 4.5005
R11758 DVDD.n17954 DVDD.n749 4.5005
R11759 DVDD.n771 DVDD.n743 4.5005
R11760 DVDD.n771 DVDD.n733 4.5005
R11761 DVDD.n771 DVDD.n744 4.5005
R11762 DVDD.n771 DVDD.n732 4.5005
R11763 DVDD.n771 DVDD.n745 4.5005
R11764 DVDD.n771 DVDD.n731 4.5005
R11765 DVDD.n17954 DVDD.n771 4.5005
R11766 DVDD.n748 DVDD.n743 4.5005
R11767 DVDD.n748 DVDD.n733 4.5005
R11768 DVDD.n748 DVDD.n744 4.5005
R11769 DVDD.n748 DVDD.n732 4.5005
R11770 DVDD.n748 DVDD.n745 4.5005
R11771 DVDD.n748 DVDD.n731 4.5005
R11772 DVDD.n17954 DVDD.n748 4.5005
R11773 DVDD.n17953 DVDD.n739 4.5005
R11774 DVDD.n17953 DVDD.n737 4.5005
R11775 DVDD.n17953 DVDD.n740 4.5005
R11776 DVDD.n17953 DVDD.n736 4.5005
R11777 DVDD.n17953 DVDD.n741 4.5005
R11778 DVDD.n17953 DVDD.n735 4.5005
R11779 DVDD.n17953 DVDD.n742 4.5005
R11780 DVDD.n17953 DVDD.n734 4.5005
R11781 DVDD.n17953 DVDD.n743 4.5005
R11782 DVDD.n17953 DVDD.n733 4.5005
R11783 DVDD.n17953 DVDD.n744 4.5005
R11784 DVDD.n17953 DVDD.n732 4.5005
R11785 DVDD.n17953 DVDD.n745 4.5005
R11786 DVDD.n17953 DVDD.n731 4.5005
R11787 DVDD.n17954 DVDD.n17953 4.5005
R11788 DVDD.n747 DVDD.n739 4.5005
R11789 DVDD.n747 DVDD.n737 4.5005
R11790 DVDD.n747 DVDD.n740 4.5005
R11791 DVDD.n747 DVDD.n736 4.5005
R11792 DVDD.n747 DVDD.n741 4.5005
R11793 DVDD.n747 DVDD.n735 4.5005
R11794 DVDD.n747 DVDD.n742 4.5005
R11795 DVDD.n747 DVDD.n734 4.5005
R11796 DVDD.n747 DVDD.n743 4.5005
R11797 DVDD.n747 DVDD.n733 4.5005
R11798 DVDD.n747 DVDD.n744 4.5005
R11799 DVDD.n747 DVDD.n732 4.5005
R11800 DVDD.n747 DVDD.n745 4.5005
R11801 DVDD.n747 DVDD.n731 4.5005
R11802 DVDD.n17954 DVDD.n747 4.5005
R11803 DVDD.n17955 DVDD.n739 4.5005
R11804 DVDD.n17955 DVDD.n737 4.5005
R11805 DVDD.n17955 DVDD.n740 4.5005
R11806 DVDD.n17955 DVDD.n736 4.5005
R11807 DVDD.n17955 DVDD.n741 4.5005
R11808 DVDD.n17955 DVDD.n735 4.5005
R11809 DVDD.n17955 DVDD.n742 4.5005
R11810 DVDD.n17955 DVDD.n734 4.5005
R11811 DVDD.n17955 DVDD.n743 4.5005
R11812 DVDD.n17955 DVDD.n733 4.5005
R11813 DVDD.n17955 DVDD.n744 4.5005
R11814 DVDD.n17955 DVDD.n732 4.5005
R11815 DVDD.n17955 DVDD.n745 4.5005
R11816 DVDD.n17955 DVDD.n731 4.5005
R11817 DVDD.n17955 DVDD.n17954 4.5005
R11818 DVDD.n17962 DVDD.n649 4.5005
R11819 DVDD.n17962 DVDD.n647 4.5005
R11820 DVDD.n17962 DVDD.n650 4.5005
R11821 DVDD.n17962 DVDD.n646 4.5005
R11822 DVDD.n17962 DVDD.n651 4.5005
R11823 DVDD.n17962 DVDD.n645 4.5005
R11824 DVDD.n17962 DVDD.n652 4.5005
R11825 DVDD.n657 DVDD.n649 4.5005
R11826 DVDD.n657 DVDD.n647 4.5005
R11827 DVDD.n657 DVDD.n650 4.5005
R11828 DVDD.n657 DVDD.n646 4.5005
R11829 DVDD.n657 DVDD.n651 4.5005
R11830 DVDD.n657 DVDD.n645 4.5005
R11831 DVDD.n657 DVDD.n652 4.5005
R11832 DVDD.n680 DVDD.n649 4.5005
R11833 DVDD.n680 DVDD.n647 4.5005
R11834 DVDD.n680 DVDD.n650 4.5005
R11835 DVDD.n680 DVDD.n646 4.5005
R11836 DVDD.n680 DVDD.n651 4.5005
R11837 DVDD.n680 DVDD.n645 4.5005
R11838 DVDD.n680 DVDD.n652 4.5005
R11839 DVDD.n17963 DVDD.n669 4.5005
R11840 DVDD.n669 DVDD.n641 4.5005
R11841 DVDD.n669 DVDD.n655 4.5005
R11842 DVDD.n669 DVDD.n642 4.5005
R11843 DVDD.n669 DVDD.n653 4.5005
R11844 DVDD.n669 DVDD.n644 4.5005
R11845 DVDD.n669 DVDD.n649 4.5005
R11846 DVDD.n669 DVDD.n647 4.5005
R11847 DVDD.n669 DVDD.n650 4.5005
R11848 DVDD.n669 DVDD.n646 4.5005
R11849 DVDD.n669 DVDD.n652 4.5005
R11850 DVDD.n17963 DVDD.n671 4.5005
R11851 DVDD.n671 DVDD.n641 4.5005
R11852 DVDD.n671 DVDD.n655 4.5005
R11853 DVDD.n671 DVDD.n642 4.5005
R11854 DVDD.n671 DVDD.n654 4.5005
R11855 DVDD.n671 DVDD.n643 4.5005
R11856 DVDD.n671 DVDD.n653 4.5005
R11857 DVDD.n671 DVDD.n644 4.5005
R11858 DVDD.n671 DVDD.n649 4.5005
R11859 DVDD.n671 DVDD.n647 4.5005
R11860 DVDD.n671 DVDD.n650 4.5005
R11861 DVDD.n671 DVDD.n646 4.5005
R11862 DVDD.n671 DVDD.n651 4.5005
R11863 DVDD.n671 DVDD.n645 4.5005
R11864 DVDD.n671 DVDD.n652 4.5005
R11865 DVDD.n17963 DVDD.n666 4.5005
R11866 DVDD.n666 DVDD.n641 4.5005
R11867 DVDD.n666 DVDD.n655 4.5005
R11868 DVDD.n666 DVDD.n642 4.5005
R11869 DVDD.n666 DVDD.n654 4.5005
R11870 DVDD.n666 DVDD.n643 4.5005
R11871 DVDD.n666 DVDD.n653 4.5005
R11872 DVDD.n666 DVDD.n644 4.5005
R11873 DVDD.n666 DVDD.n649 4.5005
R11874 DVDD.n666 DVDD.n647 4.5005
R11875 DVDD.n666 DVDD.n650 4.5005
R11876 DVDD.n666 DVDD.n646 4.5005
R11877 DVDD.n666 DVDD.n651 4.5005
R11878 DVDD.n666 DVDD.n645 4.5005
R11879 DVDD.n666 DVDD.n652 4.5005
R11880 DVDD.n658 DVDD.n649 4.5005
R11881 DVDD.n658 DVDD.n647 4.5005
R11882 DVDD.n658 DVDD.n650 4.5005
R11883 DVDD.n658 DVDD.n646 4.5005
R11884 DVDD.n658 DVDD.n651 4.5005
R11885 DVDD.n658 DVDD.n645 4.5005
R11886 DVDD.n658 DVDD.n652 4.5005
R11887 DVDD.n679 DVDD.n649 4.5005
R11888 DVDD.n679 DVDD.n647 4.5005
R11889 DVDD.n679 DVDD.n650 4.5005
R11890 DVDD.n679 DVDD.n646 4.5005
R11891 DVDD.n679 DVDD.n651 4.5005
R11892 DVDD.n679 DVDD.n645 4.5005
R11893 DVDD.n679 DVDD.n652 4.5005
R11894 DVDD.n659 DVDD.n649 4.5005
R11895 DVDD.n659 DVDD.n647 4.5005
R11896 DVDD.n659 DVDD.n650 4.5005
R11897 DVDD.n659 DVDD.n646 4.5005
R11898 DVDD.n659 DVDD.n651 4.5005
R11899 DVDD.n659 DVDD.n645 4.5005
R11900 DVDD.n659 DVDD.n652 4.5005
R11901 DVDD.n678 DVDD.n649 4.5005
R11902 DVDD.n678 DVDD.n647 4.5005
R11903 DVDD.n678 DVDD.n650 4.5005
R11904 DVDD.n678 DVDD.n646 4.5005
R11905 DVDD.n678 DVDD.n651 4.5005
R11906 DVDD.n678 DVDD.n645 4.5005
R11907 DVDD.n678 DVDD.n652 4.5005
R11908 DVDD.n17963 DVDD.n672 4.5005
R11909 DVDD.n672 DVDD.n641 4.5005
R11910 DVDD.n672 DVDD.n655 4.5005
R11911 DVDD.n672 DVDD.n642 4.5005
R11912 DVDD.n672 DVDD.n654 4.5005
R11913 DVDD.n672 DVDD.n643 4.5005
R11914 DVDD.n672 DVDD.n653 4.5005
R11915 DVDD.n672 DVDD.n644 4.5005
R11916 DVDD.n672 DVDD.n649 4.5005
R11917 DVDD.n672 DVDD.n647 4.5005
R11918 DVDD.n672 DVDD.n650 4.5005
R11919 DVDD.n672 DVDD.n646 4.5005
R11920 DVDD.n672 DVDD.n651 4.5005
R11921 DVDD.n672 DVDD.n645 4.5005
R11922 DVDD.n672 DVDD.n652 4.5005
R11923 DVDD.n17963 DVDD.n665 4.5005
R11924 DVDD.n665 DVDD.n641 4.5005
R11925 DVDD.n665 DVDD.n655 4.5005
R11926 DVDD.n665 DVDD.n642 4.5005
R11927 DVDD.n665 DVDD.n654 4.5005
R11928 DVDD.n665 DVDD.n643 4.5005
R11929 DVDD.n665 DVDD.n653 4.5005
R11930 DVDD.n665 DVDD.n644 4.5005
R11931 DVDD.n665 DVDD.n649 4.5005
R11932 DVDD.n665 DVDD.n647 4.5005
R11933 DVDD.n665 DVDD.n650 4.5005
R11934 DVDD.n665 DVDD.n646 4.5005
R11935 DVDD.n665 DVDD.n651 4.5005
R11936 DVDD.n665 DVDD.n645 4.5005
R11937 DVDD.n665 DVDD.n652 4.5005
R11938 DVDD.n17963 DVDD.n673 4.5005
R11939 DVDD.n673 DVDD.n641 4.5005
R11940 DVDD.n673 DVDD.n655 4.5005
R11941 DVDD.n673 DVDD.n642 4.5005
R11942 DVDD.n673 DVDD.n654 4.5005
R11943 DVDD.n673 DVDD.n643 4.5005
R11944 DVDD.n673 DVDD.n653 4.5005
R11945 DVDD.n673 DVDD.n644 4.5005
R11946 DVDD.n673 DVDD.n649 4.5005
R11947 DVDD.n673 DVDD.n647 4.5005
R11948 DVDD.n673 DVDD.n650 4.5005
R11949 DVDD.n673 DVDD.n646 4.5005
R11950 DVDD.n673 DVDD.n651 4.5005
R11951 DVDD.n673 DVDD.n645 4.5005
R11952 DVDD.n673 DVDD.n652 4.5005
R11953 DVDD.n660 DVDD.n649 4.5005
R11954 DVDD.n660 DVDD.n647 4.5005
R11955 DVDD.n660 DVDD.n650 4.5005
R11956 DVDD.n660 DVDD.n646 4.5005
R11957 DVDD.n660 DVDD.n651 4.5005
R11958 DVDD.n660 DVDD.n645 4.5005
R11959 DVDD.n660 DVDD.n652 4.5005
R11960 DVDD.n677 DVDD.n649 4.5005
R11961 DVDD.n677 DVDD.n647 4.5005
R11962 DVDD.n677 DVDD.n650 4.5005
R11963 DVDD.n677 DVDD.n646 4.5005
R11964 DVDD.n677 DVDD.n651 4.5005
R11965 DVDD.n677 DVDD.n645 4.5005
R11966 DVDD.n677 DVDD.n652 4.5005
R11967 DVDD.n661 DVDD.n649 4.5005
R11968 DVDD.n661 DVDD.n647 4.5005
R11969 DVDD.n661 DVDD.n650 4.5005
R11970 DVDD.n661 DVDD.n646 4.5005
R11971 DVDD.n661 DVDD.n651 4.5005
R11972 DVDD.n661 DVDD.n645 4.5005
R11973 DVDD.n661 DVDD.n652 4.5005
R11974 DVDD.n17963 DVDD.n664 4.5005
R11975 DVDD.n664 DVDD.n641 4.5005
R11976 DVDD.n664 DVDD.n655 4.5005
R11977 DVDD.n664 DVDD.n642 4.5005
R11978 DVDD.n664 DVDD.n654 4.5005
R11979 DVDD.n664 DVDD.n643 4.5005
R11980 DVDD.n664 DVDD.n653 4.5005
R11981 DVDD.n664 DVDD.n644 4.5005
R11982 DVDD.n664 DVDD.n649 4.5005
R11983 DVDD.n664 DVDD.n647 4.5005
R11984 DVDD.n664 DVDD.n650 4.5005
R11985 DVDD.n664 DVDD.n646 4.5005
R11986 DVDD.n664 DVDD.n651 4.5005
R11987 DVDD.n664 DVDD.n645 4.5005
R11988 DVDD.n664 DVDD.n652 4.5005
R11989 DVDD.n17963 DVDD.n674 4.5005
R11990 DVDD.n674 DVDD.n641 4.5005
R11991 DVDD.n674 DVDD.n655 4.5005
R11992 DVDD.n674 DVDD.n642 4.5005
R11993 DVDD.n674 DVDD.n654 4.5005
R11994 DVDD.n674 DVDD.n643 4.5005
R11995 DVDD.n674 DVDD.n653 4.5005
R11996 DVDD.n674 DVDD.n644 4.5005
R11997 DVDD.n674 DVDD.n649 4.5005
R11998 DVDD.n674 DVDD.n647 4.5005
R11999 DVDD.n674 DVDD.n650 4.5005
R12000 DVDD.n674 DVDD.n646 4.5005
R12001 DVDD.n674 DVDD.n651 4.5005
R12002 DVDD.n674 DVDD.n645 4.5005
R12003 DVDD.n674 DVDD.n652 4.5005
R12004 DVDD.n17963 DVDD.n663 4.5005
R12005 DVDD.n663 DVDD.n641 4.5005
R12006 DVDD.n663 DVDD.n655 4.5005
R12007 DVDD.n663 DVDD.n642 4.5005
R12008 DVDD.n663 DVDD.n654 4.5005
R12009 DVDD.n663 DVDD.n643 4.5005
R12010 DVDD.n663 DVDD.n653 4.5005
R12011 DVDD.n663 DVDD.n644 4.5005
R12012 DVDD.n663 DVDD.n649 4.5005
R12013 DVDD.n663 DVDD.n647 4.5005
R12014 DVDD.n663 DVDD.n650 4.5005
R12015 DVDD.n663 DVDD.n646 4.5005
R12016 DVDD.n663 DVDD.n651 4.5005
R12017 DVDD.n663 DVDD.n645 4.5005
R12018 DVDD.n663 DVDD.n652 4.5005
R12019 DVDD.n17963 DVDD.n675 4.5005
R12020 DVDD.n675 DVDD.n641 4.5005
R12021 DVDD.n675 DVDD.n655 4.5005
R12022 DVDD.n675 DVDD.n642 4.5005
R12023 DVDD.n675 DVDD.n654 4.5005
R12024 DVDD.n675 DVDD.n643 4.5005
R12025 DVDD.n675 DVDD.n653 4.5005
R12026 DVDD.n675 DVDD.n644 4.5005
R12027 DVDD.n675 DVDD.n649 4.5005
R12028 DVDD.n675 DVDD.n647 4.5005
R12029 DVDD.n675 DVDD.n650 4.5005
R12030 DVDD.n675 DVDD.n646 4.5005
R12031 DVDD.n675 DVDD.n651 4.5005
R12032 DVDD.n675 DVDD.n645 4.5005
R12033 DVDD.n675 DVDD.n652 4.5005
R12034 DVDD.n676 DVDD.n649 4.5005
R12035 DVDD.n676 DVDD.n647 4.5005
R12036 DVDD.n676 DVDD.n650 4.5005
R12037 DVDD.n676 DVDD.n646 4.5005
R12038 DVDD.n676 DVDD.n651 4.5005
R12039 DVDD.n676 DVDD.n645 4.5005
R12040 DVDD.n676 DVDD.n652 4.5005
R12041 DVDD.n662 DVDD.n649 4.5005
R12042 DVDD.n662 DVDD.n647 4.5005
R12043 DVDD.n662 DVDD.n650 4.5005
R12044 DVDD.n662 DVDD.n646 4.5005
R12045 DVDD.n662 DVDD.n651 4.5005
R12046 DVDD.n662 DVDD.n645 4.5005
R12047 DVDD.n662 DVDD.n652 4.5005
R12048 DVDD.n17964 DVDD.n649 4.5005
R12049 DVDD.n17964 DVDD.n647 4.5005
R12050 DVDD.n17964 DVDD.n650 4.5005
R12051 DVDD.n17964 DVDD.n646 4.5005
R12052 DVDD.n17964 DVDD.n651 4.5005
R12053 DVDD.n17964 DVDD.n645 4.5005
R12054 DVDD.n17964 DVDD.n652 4.5005
R12055 DVDD.n17963 DVDD.n639 4.5005
R12056 DVDD.n641 DVDD.n639 4.5005
R12057 DVDD.n655 DVDD.n639 4.5005
R12058 DVDD.n642 DVDD.n639 4.5005
R12059 DVDD.n654 DVDD.n639 4.5005
R12060 DVDD.n643 DVDD.n639 4.5005
R12061 DVDD.n653 DVDD.n639 4.5005
R12062 DVDD.n644 DVDD.n639 4.5005
R12063 DVDD.n649 DVDD.n639 4.5005
R12064 DVDD.n647 DVDD.n639 4.5005
R12065 DVDD.n650 DVDD.n639 4.5005
R12066 DVDD.n646 DVDD.n639 4.5005
R12067 DVDD.n651 DVDD.n639 4.5005
R12068 DVDD.n645 DVDD.n639 4.5005
R12069 DVDD.n652 DVDD.n639 4.5005
R12070 DVDD.n17978 DVDD.n582 4.5005
R12071 DVDD.n582 DVDD.n554 4.5005
R12072 DVDD.n582 DVDD.n568 4.5005
R12073 DVDD.n582 DVDD.n555 4.5005
R12074 DVDD.n582 DVDD.n566 4.5005
R12075 DVDD.n582 DVDD.n557 4.5005
R12076 DVDD.n582 DVDD.n562 4.5005
R12077 DVDD.n582 DVDD.n560 4.5005
R12078 DVDD.n582 DVDD.n563 4.5005
R12079 DVDD.n582 DVDD.n559 4.5005
R12080 DVDD.n582 DVDD.n565 4.5005
R12081 DVDD.n17978 DVDD.n584 4.5005
R12082 DVDD.n584 DVDD.n554 4.5005
R12083 DVDD.n584 DVDD.n568 4.5005
R12084 DVDD.n584 DVDD.n555 4.5005
R12085 DVDD.n584 DVDD.n567 4.5005
R12086 DVDD.n584 DVDD.n556 4.5005
R12087 DVDD.n584 DVDD.n566 4.5005
R12088 DVDD.n584 DVDD.n557 4.5005
R12089 DVDD.n584 DVDD.n562 4.5005
R12090 DVDD.n584 DVDD.n560 4.5005
R12091 DVDD.n584 DVDD.n563 4.5005
R12092 DVDD.n584 DVDD.n559 4.5005
R12093 DVDD.n584 DVDD.n564 4.5005
R12094 DVDD.n584 DVDD.n558 4.5005
R12095 DVDD.n584 DVDD.n565 4.5005
R12096 DVDD.n17977 DVDD.n562 4.5005
R12097 DVDD.n17977 DVDD.n560 4.5005
R12098 DVDD.n17977 DVDD.n563 4.5005
R12099 DVDD.n17977 DVDD.n559 4.5005
R12100 DVDD.n17977 DVDD.n564 4.5005
R12101 DVDD.n17977 DVDD.n558 4.5005
R12102 DVDD.n17977 DVDD.n565 4.5005
R12103 DVDD.n570 DVDD.n562 4.5005
R12104 DVDD.n570 DVDD.n560 4.5005
R12105 DVDD.n570 DVDD.n563 4.5005
R12106 DVDD.n570 DVDD.n559 4.5005
R12107 DVDD.n570 DVDD.n564 4.5005
R12108 DVDD.n570 DVDD.n558 4.5005
R12109 DVDD.n570 DVDD.n565 4.5005
R12110 DVDD.n593 DVDD.n562 4.5005
R12111 DVDD.n593 DVDD.n560 4.5005
R12112 DVDD.n593 DVDD.n563 4.5005
R12113 DVDD.n593 DVDD.n559 4.5005
R12114 DVDD.n593 DVDD.n564 4.5005
R12115 DVDD.n593 DVDD.n558 4.5005
R12116 DVDD.n593 DVDD.n565 4.5005
R12117 DVDD.n17978 DVDD.n579 4.5005
R12118 DVDD.n579 DVDD.n554 4.5005
R12119 DVDD.n579 DVDD.n568 4.5005
R12120 DVDD.n579 DVDD.n555 4.5005
R12121 DVDD.n579 DVDD.n567 4.5005
R12122 DVDD.n579 DVDD.n556 4.5005
R12123 DVDD.n579 DVDD.n566 4.5005
R12124 DVDD.n579 DVDD.n557 4.5005
R12125 DVDD.n579 DVDD.n562 4.5005
R12126 DVDD.n579 DVDD.n560 4.5005
R12127 DVDD.n579 DVDD.n563 4.5005
R12128 DVDD.n579 DVDD.n559 4.5005
R12129 DVDD.n579 DVDD.n564 4.5005
R12130 DVDD.n579 DVDD.n558 4.5005
R12131 DVDD.n579 DVDD.n565 4.5005
R12132 DVDD.n17978 DVDD.n585 4.5005
R12133 DVDD.n585 DVDD.n554 4.5005
R12134 DVDD.n585 DVDD.n568 4.5005
R12135 DVDD.n585 DVDD.n555 4.5005
R12136 DVDD.n585 DVDD.n567 4.5005
R12137 DVDD.n585 DVDD.n556 4.5005
R12138 DVDD.n585 DVDD.n566 4.5005
R12139 DVDD.n585 DVDD.n557 4.5005
R12140 DVDD.n585 DVDD.n562 4.5005
R12141 DVDD.n585 DVDD.n560 4.5005
R12142 DVDD.n585 DVDD.n563 4.5005
R12143 DVDD.n585 DVDD.n559 4.5005
R12144 DVDD.n585 DVDD.n564 4.5005
R12145 DVDD.n585 DVDD.n558 4.5005
R12146 DVDD.n585 DVDD.n565 4.5005
R12147 DVDD.n17978 DVDD.n578 4.5005
R12148 DVDD.n578 DVDD.n554 4.5005
R12149 DVDD.n578 DVDD.n568 4.5005
R12150 DVDD.n578 DVDD.n555 4.5005
R12151 DVDD.n578 DVDD.n567 4.5005
R12152 DVDD.n578 DVDD.n556 4.5005
R12153 DVDD.n578 DVDD.n566 4.5005
R12154 DVDD.n578 DVDD.n557 4.5005
R12155 DVDD.n578 DVDD.n562 4.5005
R12156 DVDD.n578 DVDD.n560 4.5005
R12157 DVDD.n578 DVDD.n563 4.5005
R12158 DVDD.n578 DVDD.n559 4.5005
R12159 DVDD.n578 DVDD.n564 4.5005
R12160 DVDD.n578 DVDD.n558 4.5005
R12161 DVDD.n578 DVDD.n565 4.5005
R12162 DVDD.n17978 DVDD.n586 4.5005
R12163 DVDD.n586 DVDD.n554 4.5005
R12164 DVDD.n586 DVDD.n568 4.5005
R12165 DVDD.n586 DVDD.n555 4.5005
R12166 DVDD.n586 DVDD.n567 4.5005
R12167 DVDD.n586 DVDD.n556 4.5005
R12168 DVDD.n586 DVDD.n566 4.5005
R12169 DVDD.n586 DVDD.n557 4.5005
R12170 DVDD.n586 DVDD.n562 4.5005
R12171 DVDD.n586 DVDD.n560 4.5005
R12172 DVDD.n586 DVDD.n563 4.5005
R12173 DVDD.n586 DVDD.n559 4.5005
R12174 DVDD.n586 DVDD.n564 4.5005
R12175 DVDD.n586 DVDD.n558 4.5005
R12176 DVDD.n586 DVDD.n565 4.5005
R12177 DVDD.n571 DVDD.n562 4.5005
R12178 DVDD.n571 DVDD.n560 4.5005
R12179 DVDD.n571 DVDD.n563 4.5005
R12180 DVDD.n571 DVDD.n559 4.5005
R12181 DVDD.n571 DVDD.n564 4.5005
R12182 DVDD.n571 DVDD.n558 4.5005
R12183 DVDD.n571 DVDD.n565 4.5005
R12184 DVDD.n592 DVDD.n562 4.5005
R12185 DVDD.n592 DVDD.n560 4.5005
R12186 DVDD.n592 DVDD.n563 4.5005
R12187 DVDD.n592 DVDD.n559 4.5005
R12188 DVDD.n592 DVDD.n564 4.5005
R12189 DVDD.n592 DVDD.n558 4.5005
R12190 DVDD.n592 DVDD.n565 4.5005
R12191 DVDD.n572 DVDD.n562 4.5005
R12192 DVDD.n572 DVDD.n560 4.5005
R12193 DVDD.n572 DVDD.n563 4.5005
R12194 DVDD.n572 DVDD.n559 4.5005
R12195 DVDD.n572 DVDD.n564 4.5005
R12196 DVDD.n572 DVDD.n558 4.5005
R12197 DVDD.n572 DVDD.n565 4.5005
R12198 DVDD.n17978 DVDD.n577 4.5005
R12199 DVDD.n577 DVDD.n554 4.5005
R12200 DVDD.n577 DVDD.n568 4.5005
R12201 DVDD.n577 DVDD.n555 4.5005
R12202 DVDD.n577 DVDD.n567 4.5005
R12203 DVDD.n577 DVDD.n556 4.5005
R12204 DVDD.n577 DVDD.n566 4.5005
R12205 DVDD.n577 DVDD.n557 4.5005
R12206 DVDD.n577 DVDD.n562 4.5005
R12207 DVDD.n577 DVDD.n560 4.5005
R12208 DVDD.n577 DVDD.n563 4.5005
R12209 DVDD.n577 DVDD.n559 4.5005
R12210 DVDD.n577 DVDD.n564 4.5005
R12211 DVDD.n577 DVDD.n558 4.5005
R12212 DVDD.n577 DVDD.n565 4.5005
R12213 DVDD.n17978 DVDD.n587 4.5005
R12214 DVDD.n587 DVDD.n554 4.5005
R12215 DVDD.n587 DVDD.n568 4.5005
R12216 DVDD.n587 DVDD.n555 4.5005
R12217 DVDD.n587 DVDD.n567 4.5005
R12218 DVDD.n587 DVDD.n556 4.5005
R12219 DVDD.n587 DVDD.n566 4.5005
R12220 DVDD.n587 DVDD.n557 4.5005
R12221 DVDD.n587 DVDD.n562 4.5005
R12222 DVDD.n587 DVDD.n560 4.5005
R12223 DVDD.n587 DVDD.n563 4.5005
R12224 DVDD.n587 DVDD.n559 4.5005
R12225 DVDD.n587 DVDD.n564 4.5005
R12226 DVDD.n587 DVDD.n558 4.5005
R12227 DVDD.n587 DVDD.n565 4.5005
R12228 DVDD.n17978 DVDD.n576 4.5005
R12229 DVDD.n576 DVDD.n554 4.5005
R12230 DVDD.n576 DVDD.n568 4.5005
R12231 DVDD.n576 DVDD.n555 4.5005
R12232 DVDD.n576 DVDD.n567 4.5005
R12233 DVDD.n576 DVDD.n556 4.5005
R12234 DVDD.n576 DVDD.n566 4.5005
R12235 DVDD.n576 DVDD.n557 4.5005
R12236 DVDD.n576 DVDD.n562 4.5005
R12237 DVDD.n576 DVDD.n560 4.5005
R12238 DVDD.n576 DVDD.n563 4.5005
R12239 DVDD.n576 DVDD.n559 4.5005
R12240 DVDD.n576 DVDD.n564 4.5005
R12241 DVDD.n576 DVDD.n558 4.5005
R12242 DVDD.n576 DVDD.n565 4.5005
R12243 DVDD.n17978 DVDD.n588 4.5005
R12244 DVDD.n588 DVDD.n554 4.5005
R12245 DVDD.n588 DVDD.n568 4.5005
R12246 DVDD.n588 DVDD.n555 4.5005
R12247 DVDD.n588 DVDD.n567 4.5005
R12248 DVDD.n588 DVDD.n556 4.5005
R12249 DVDD.n588 DVDD.n566 4.5005
R12250 DVDD.n588 DVDD.n557 4.5005
R12251 DVDD.n588 DVDD.n562 4.5005
R12252 DVDD.n588 DVDD.n560 4.5005
R12253 DVDD.n588 DVDD.n563 4.5005
R12254 DVDD.n588 DVDD.n559 4.5005
R12255 DVDD.n588 DVDD.n564 4.5005
R12256 DVDD.n588 DVDD.n558 4.5005
R12257 DVDD.n588 DVDD.n565 4.5005
R12258 DVDD.n591 DVDD.n562 4.5005
R12259 DVDD.n591 DVDD.n560 4.5005
R12260 DVDD.n591 DVDD.n563 4.5005
R12261 DVDD.n591 DVDD.n559 4.5005
R12262 DVDD.n591 DVDD.n564 4.5005
R12263 DVDD.n591 DVDD.n558 4.5005
R12264 DVDD.n591 DVDD.n565 4.5005
R12265 DVDD.n573 DVDD.n562 4.5005
R12266 DVDD.n573 DVDD.n560 4.5005
R12267 DVDD.n573 DVDD.n563 4.5005
R12268 DVDD.n573 DVDD.n559 4.5005
R12269 DVDD.n573 DVDD.n564 4.5005
R12270 DVDD.n573 DVDD.n558 4.5005
R12271 DVDD.n573 DVDD.n565 4.5005
R12272 DVDD.n590 DVDD.n562 4.5005
R12273 DVDD.n590 DVDD.n560 4.5005
R12274 DVDD.n590 DVDD.n563 4.5005
R12275 DVDD.n590 DVDD.n559 4.5005
R12276 DVDD.n590 DVDD.n564 4.5005
R12277 DVDD.n590 DVDD.n558 4.5005
R12278 DVDD.n590 DVDD.n565 4.5005
R12279 DVDD.n17978 DVDD.n575 4.5005
R12280 DVDD.n575 DVDD.n554 4.5005
R12281 DVDD.n575 DVDD.n568 4.5005
R12282 DVDD.n575 DVDD.n555 4.5005
R12283 DVDD.n575 DVDD.n567 4.5005
R12284 DVDD.n575 DVDD.n556 4.5005
R12285 DVDD.n575 DVDD.n566 4.5005
R12286 DVDD.n575 DVDD.n557 4.5005
R12287 DVDD.n575 DVDD.n562 4.5005
R12288 DVDD.n575 DVDD.n560 4.5005
R12289 DVDD.n575 DVDD.n563 4.5005
R12290 DVDD.n575 DVDD.n559 4.5005
R12291 DVDD.n575 DVDD.n564 4.5005
R12292 DVDD.n575 DVDD.n558 4.5005
R12293 DVDD.n575 DVDD.n565 4.5005
R12294 DVDD.n17978 DVDD.n589 4.5005
R12295 DVDD.n589 DVDD.n554 4.5005
R12296 DVDD.n589 DVDD.n568 4.5005
R12297 DVDD.n589 DVDD.n555 4.5005
R12298 DVDD.n589 DVDD.n567 4.5005
R12299 DVDD.n589 DVDD.n556 4.5005
R12300 DVDD.n589 DVDD.n566 4.5005
R12301 DVDD.n589 DVDD.n557 4.5005
R12302 DVDD.n589 DVDD.n562 4.5005
R12303 DVDD.n589 DVDD.n560 4.5005
R12304 DVDD.n589 DVDD.n563 4.5005
R12305 DVDD.n589 DVDD.n559 4.5005
R12306 DVDD.n589 DVDD.n564 4.5005
R12307 DVDD.n589 DVDD.n558 4.5005
R12308 DVDD.n589 DVDD.n565 4.5005
R12309 DVDD.n17978 DVDD.n574 4.5005
R12310 DVDD.n574 DVDD.n554 4.5005
R12311 DVDD.n574 DVDD.n568 4.5005
R12312 DVDD.n574 DVDD.n555 4.5005
R12313 DVDD.n574 DVDD.n567 4.5005
R12314 DVDD.n574 DVDD.n556 4.5005
R12315 DVDD.n574 DVDD.n566 4.5005
R12316 DVDD.n574 DVDD.n557 4.5005
R12317 DVDD.n574 DVDD.n562 4.5005
R12318 DVDD.n574 DVDD.n560 4.5005
R12319 DVDD.n574 DVDD.n563 4.5005
R12320 DVDD.n574 DVDD.n559 4.5005
R12321 DVDD.n574 DVDD.n564 4.5005
R12322 DVDD.n574 DVDD.n558 4.5005
R12323 DVDD.n574 DVDD.n565 4.5005
R12324 DVDD.n17979 DVDD.n562 4.5005
R12325 DVDD.n17979 DVDD.n560 4.5005
R12326 DVDD.n17979 DVDD.n563 4.5005
R12327 DVDD.n17979 DVDD.n559 4.5005
R12328 DVDD.n17979 DVDD.n564 4.5005
R12329 DVDD.n17979 DVDD.n558 4.5005
R12330 DVDD.n17979 DVDD.n565 4.5005
R12331 DVDD.n562 DVDD.n552 4.5005
R12332 DVDD.n560 DVDD.n552 4.5005
R12333 DVDD.n563 DVDD.n552 4.5005
R12334 DVDD.n559 DVDD.n552 4.5005
R12335 DVDD.n564 DVDD.n552 4.5005
R12336 DVDD.n558 DVDD.n552 4.5005
R12337 DVDD.n565 DVDD.n552 4.5005
R12338 DVDD.n529 DVDD.n514 4.5005
R12339 DVDD.n529 DVDD.n505 4.5005
R12340 DVDD.n529 DVDD.n515 4.5005
R12341 DVDD.n529 DVDD.n504 4.5005
R12342 DVDD.n529 DVDD.n516 4.5005
R12343 DVDD.n18040 DVDD.n529 4.5005
R12344 DVDD.n18043 DVDD.n529 4.5005
R12345 DVDD.n532 DVDD.n510 4.5005
R12346 DVDD.n532 DVDD.n509 4.5005
R12347 DVDD.n532 DVDD.n511 4.5005
R12348 DVDD.n532 DVDD.n508 4.5005
R12349 DVDD.n532 DVDD.n513 4.5005
R12350 DVDD.n532 DVDD.n506 4.5005
R12351 DVDD.n532 DVDD.n514 4.5005
R12352 DVDD.n532 DVDD.n505 4.5005
R12353 DVDD.n532 DVDD.n515 4.5005
R12354 DVDD.n532 DVDD.n504 4.5005
R12355 DVDD.n18043 DVDD.n532 4.5005
R12356 DVDD.n528 DVDD.n510 4.5005
R12357 DVDD.n528 DVDD.n509 4.5005
R12358 DVDD.n528 DVDD.n511 4.5005
R12359 DVDD.n528 DVDD.n508 4.5005
R12360 DVDD.n528 DVDD.n512 4.5005
R12361 DVDD.n528 DVDD.n507 4.5005
R12362 DVDD.n528 DVDD.n513 4.5005
R12363 DVDD.n528 DVDD.n506 4.5005
R12364 DVDD.n528 DVDD.n514 4.5005
R12365 DVDD.n528 DVDD.n505 4.5005
R12366 DVDD.n528 DVDD.n515 4.5005
R12367 DVDD.n528 DVDD.n504 4.5005
R12368 DVDD.n528 DVDD.n516 4.5005
R12369 DVDD.n18040 DVDD.n528 4.5005
R12370 DVDD.n18043 DVDD.n528 4.5005
R12371 DVDD.n533 DVDD.n510 4.5005
R12372 DVDD.n533 DVDD.n509 4.5005
R12373 DVDD.n533 DVDD.n511 4.5005
R12374 DVDD.n533 DVDD.n508 4.5005
R12375 DVDD.n533 DVDD.n512 4.5005
R12376 DVDD.n533 DVDD.n507 4.5005
R12377 DVDD.n533 DVDD.n513 4.5005
R12378 DVDD.n533 DVDD.n506 4.5005
R12379 DVDD.n533 DVDD.n514 4.5005
R12380 DVDD.n533 DVDD.n505 4.5005
R12381 DVDD.n533 DVDD.n515 4.5005
R12382 DVDD.n533 DVDD.n504 4.5005
R12383 DVDD.n533 DVDD.n516 4.5005
R12384 DVDD.n18040 DVDD.n533 4.5005
R12385 DVDD.n18043 DVDD.n533 4.5005
R12386 DVDD.n527 DVDD.n510 4.5005
R12387 DVDD.n527 DVDD.n509 4.5005
R12388 DVDD.n527 DVDD.n511 4.5005
R12389 DVDD.n527 DVDD.n508 4.5005
R12390 DVDD.n527 DVDD.n512 4.5005
R12391 DVDD.n527 DVDD.n507 4.5005
R12392 DVDD.n527 DVDD.n513 4.5005
R12393 DVDD.n527 DVDD.n506 4.5005
R12394 DVDD.n527 DVDD.n514 4.5005
R12395 DVDD.n527 DVDD.n505 4.5005
R12396 DVDD.n527 DVDD.n515 4.5005
R12397 DVDD.n527 DVDD.n504 4.5005
R12398 DVDD.n527 DVDD.n516 4.5005
R12399 DVDD.n18040 DVDD.n527 4.5005
R12400 DVDD.n18043 DVDD.n527 4.5005
R12401 DVDD.n534 DVDD.n514 4.5005
R12402 DVDD.n534 DVDD.n505 4.5005
R12403 DVDD.n534 DVDD.n515 4.5005
R12404 DVDD.n534 DVDD.n504 4.5005
R12405 DVDD.n534 DVDD.n516 4.5005
R12406 DVDD.n18040 DVDD.n534 4.5005
R12407 DVDD.n18043 DVDD.n534 4.5005
R12408 DVDD.n526 DVDD.n514 4.5005
R12409 DVDD.n526 DVDD.n505 4.5005
R12410 DVDD.n526 DVDD.n515 4.5005
R12411 DVDD.n526 DVDD.n504 4.5005
R12412 DVDD.n526 DVDD.n516 4.5005
R12413 DVDD.n18040 DVDD.n526 4.5005
R12414 DVDD.n18043 DVDD.n526 4.5005
R12415 DVDD.n535 DVDD.n514 4.5005
R12416 DVDD.n535 DVDD.n505 4.5005
R12417 DVDD.n535 DVDD.n515 4.5005
R12418 DVDD.n535 DVDD.n504 4.5005
R12419 DVDD.n535 DVDD.n516 4.5005
R12420 DVDD.n18040 DVDD.n535 4.5005
R12421 DVDD.n18043 DVDD.n535 4.5005
R12422 DVDD.n525 DVDD.n510 4.5005
R12423 DVDD.n525 DVDD.n509 4.5005
R12424 DVDD.n525 DVDD.n511 4.5005
R12425 DVDD.n525 DVDD.n508 4.5005
R12426 DVDD.n525 DVDD.n512 4.5005
R12427 DVDD.n525 DVDD.n507 4.5005
R12428 DVDD.n525 DVDD.n513 4.5005
R12429 DVDD.n525 DVDD.n506 4.5005
R12430 DVDD.n525 DVDD.n514 4.5005
R12431 DVDD.n525 DVDD.n505 4.5005
R12432 DVDD.n525 DVDD.n515 4.5005
R12433 DVDD.n525 DVDD.n504 4.5005
R12434 DVDD.n525 DVDD.n516 4.5005
R12435 DVDD.n18040 DVDD.n525 4.5005
R12436 DVDD.n18043 DVDD.n525 4.5005
R12437 DVDD.n536 DVDD.n510 4.5005
R12438 DVDD.n536 DVDD.n509 4.5005
R12439 DVDD.n536 DVDD.n511 4.5005
R12440 DVDD.n536 DVDD.n508 4.5005
R12441 DVDD.n536 DVDD.n512 4.5005
R12442 DVDD.n536 DVDD.n507 4.5005
R12443 DVDD.n536 DVDD.n513 4.5005
R12444 DVDD.n536 DVDD.n506 4.5005
R12445 DVDD.n536 DVDD.n514 4.5005
R12446 DVDD.n536 DVDD.n505 4.5005
R12447 DVDD.n536 DVDD.n515 4.5005
R12448 DVDD.n536 DVDD.n504 4.5005
R12449 DVDD.n536 DVDD.n516 4.5005
R12450 DVDD.n18040 DVDD.n536 4.5005
R12451 DVDD.n18043 DVDD.n536 4.5005
R12452 DVDD.n524 DVDD.n510 4.5005
R12453 DVDD.n524 DVDD.n509 4.5005
R12454 DVDD.n524 DVDD.n511 4.5005
R12455 DVDD.n524 DVDD.n508 4.5005
R12456 DVDD.n524 DVDD.n512 4.5005
R12457 DVDD.n524 DVDD.n507 4.5005
R12458 DVDD.n524 DVDD.n513 4.5005
R12459 DVDD.n524 DVDD.n506 4.5005
R12460 DVDD.n524 DVDD.n514 4.5005
R12461 DVDD.n524 DVDD.n505 4.5005
R12462 DVDD.n524 DVDD.n515 4.5005
R12463 DVDD.n524 DVDD.n504 4.5005
R12464 DVDD.n524 DVDD.n516 4.5005
R12465 DVDD.n18040 DVDD.n524 4.5005
R12466 DVDD.n18043 DVDD.n524 4.5005
R12467 DVDD.n537 DVDD.n514 4.5005
R12468 DVDD.n537 DVDD.n505 4.5005
R12469 DVDD.n537 DVDD.n515 4.5005
R12470 DVDD.n537 DVDD.n504 4.5005
R12471 DVDD.n537 DVDD.n516 4.5005
R12472 DVDD.n18040 DVDD.n537 4.5005
R12473 DVDD.n18043 DVDD.n537 4.5005
R12474 DVDD.n523 DVDD.n514 4.5005
R12475 DVDD.n523 DVDD.n505 4.5005
R12476 DVDD.n523 DVDD.n515 4.5005
R12477 DVDD.n523 DVDD.n504 4.5005
R12478 DVDD.n523 DVDD.n516 4.5005
R12479 DVDD.n18040 DVDD.n523 4.5005
R12480 DVDD.n18043 DVDD.n523 4.5005
R12481 DVDD.n538 DVDD.n514 4.5005
R12482 DVDD.n538 DVDD.n505 4.5005
R12483 DVDD.n538 DVDD.n515 4.5005
R12484 DVDD.n538 DVDD.n504 4.5005
R12485 DVDD.n538 DVDD.n516 4.5005
R12486 DVDD.n18040 DVDD.n538 4.5005
R12487 DVDD.n18043 DVDD.n538 4.5005
R12488 DVDD.n522 DVDD.n514 4.5005
R12489 DVDD.n522 DVDD.n505 4.5005
R12490 DVDD.n522 DVDD.n515 4.5005
R12491 DVDD.n522 DVDD.n504 4.5005
R12492 DVDD.n522 DVDD.n516 4.5005
R12493 DVDD.n18040 DVDD.n522 4.5005
R12494 DVDD.n18043 DVDD.n522 4.5005
R12495 DVDD.n539 DVDD.n510 4.5005
R12496 DVDD.n539 DVDD.n509 4.5005
R12497 DVDD.n539 DVDD.n511 4.5005
R12498 DVDD.n539 DVDD.n508 4.5005
R12499 DVDD.n539 DVDD.n512 4.5005
R12500 DVDD.n539 DVDD.n507 4.5005
R12501 DVDD.n539 DVDD.n513 4.5005
R12502 DVDD.n539 DVDD.n506 4.5005
R12503 DVDD.n539 DVDD.n514 4.5005
R12504 DVDD.n539 DVDD.n505 4.5005
R12505 DVDD.n539 DVDD.n515 4.5005
R12506 DVDD.n539 DVDD.n504 4.5005
R12507 DVDD.n539 DVDD.n516 4.5005
R12508 DVDD.n18040 DVDD.n539 4.5005
R12509 DVDD.n18043 DVDD.n539 4.5005
R12510 DVDD.n521 DVDD.n510 4.5005
R12511 DVDD.n521 DVDD.n509 4.5005
R12512 DVDD.n521 DVDD.n511 4.5005
R12513 DVDD.n521 DVDD.n508 4.5005
R12514 DVDD.n521 DVDD.n512 4.5005
R12515 DVDD.n521 DVDD.n507 4.5005
R12516 DVDD.n521 DVDD.n513 4.5005
R12517 DVDD.n521 DVDD.n506 4.5005
R12518 DVDD.n521 DVDD.n514 4.5005
R12519 DVDD.n521 DVDD.n505 4.5005
R12520 DVDD.n521 DVDD.n515 4.5005
R12521 DVDD.n521 DVDD.n504 4.5005
R12522 DVDD.n521 DVDD.n516 4.5005
R12523 DVDD.n18040 DVDD.n521 4.5005
R12524 DVDD.n18043 DVDD.n521 4.5005
R12525 DVDD.n540 DVDD.n507 4.5005
R12526 DVDD.n540 DVDD.n513 4.5005
R12527 DVDD.n540 DVDD.n506 4.5005
R12528 DVDD.n540 DVDD.n514 4.5005
R12529 DVDD.n540 DVDD.n505 4.5005
R12530 DVDD.n540 DVDD.n515 4.5005
R12531 DVDD.n540 DVDD.n504 4.5005
R12532 DVDD.n540 DVDD.n516 4.5005
R12533 DVDD.n18040 DVDD.n540 4.5005
R12534 DVDD.n18043 DVDD.n540 4.5005
R12535 DVDD.n520 DVDD.n514 4.5005
R12536 DVDD.n520 DVDD.n505 4.5005
R12537 DVDD.n520 DVDD.n515 4.5005
R12538 DVDD.n520 DVDD.n504 4.5005
R12539 DVDD.n520 DVDD.n516 4.5005
R12540 DVDD.n18040 DVDD.n520 4.5005
R12541 DVDD.n18043 DVDD.n520 4.5005
R12542 DVDD.n18037 DVDD.n514 4.5005
R12543 DVDD.n18037 DVDD.n505 4.5005
R12544 DVDD.n18037 DVDD.n515 4.5005
R12545 DVDD.n18037 DVDD.n516 4.5005
R12546 DVDD.n18040 DVDD.n18037 4.5005
R12547 DVDD.n18043 DVDD.n18037 4.5005
R12548 DVDD.n519 DVDD.n510 4.5005
R12549 DVDD.n519 DVDD.n509 4.5005
R12550 DVDD.n519 DVDD.n511 4.5005
R12551 DVDD.n519 DVDD.n508 4.5005
R12552 DVDD.n519 DVDD.n512 4.5005
R12553 DVDD.n519 DVDD.n507 4.5005
R12554 DVDD.n519 DVDD.n513 4.5005
R12555 DVDD.n519 DVDD.n506 4.5005
R12556 DVDD.n519 DVDD.n514 4.5005
R12557 DVDD.n519 DVDD.n505 4.5005
R12558 DVDD.n519 DVDD.n515 4.5005
R12559 DVDD.n519 DVDD.n516 4.5005
R12560 DVDD.n18043 DVDD.n519 4.5005
R12561 DVDD.n18042 DVDD.n510 4.5005
R12562 DVDD.n18042 DVDD.n509 4.5005
R12563 DVDD.n18042 DVDD.n511 4.5005
R12564 DVDD.n18042 DVDD.n508 4.5005
R12565 DVDD.n18042 DVDD.n512 4.5005
R12566 DVDD.n18042 DVDD.n507 4.5005
R12567 DVDD.n18042 DVDD.n513 4.5005
R12568 DVDD.n18042 DVDD.n506 4.5005
R12569 DVDD.n18042 DVDD.n514 4.5005
R12570 DVDD.n18042 DVDD.n505 4.5005
R12571 DVDD.n18042 DVDD.n515 4.5005
R12572 DVDD.n18042 DVDD.n516 4.5005
R12573 DVDD.n18043 DVDD.n18042 4.5005
R12574 DVDD.n518 DVDD.n510 4.5005
R12575 DVDD.n518 DVDD.n509 4.5005
R12576 DVDD.n518 DVDD.n511 4.5005
R12577 DVDD.n518 DVDD.n508 4.5005
R12578 DVDD.n518 DVDD.n512 4.5005
R12579 DVDD.n518 DVDD.n507 4.5005
R12580 DVDD.n518 DVDD.n513 4.5005
R12581 DVDD.n518 DVDD.n506 4.5005
R12582 DVDD.n518 DVDD.n514 4.5005
R12583 DVDD.n518 DVDD.n505 4.5005
R12584 DVDD.n518 DVDD.n515 4.5005
R12585 DVDD.n518 DVDD.n516 4.5005
R12586 DVDD.n18043 DVDD.n518 4.5005
R12587 DVDD.n18044 DVDD.n510 4.5005
R12588 DVDD.n18044 DVDD.n509 4.5005
R12589 DVDD.n18044 DVDD.n511 4.5005
R12590 DVDD.n18044 DVDD.n508 4.5005
R12591 DVDD.n18044 DVDD.n512 4.5005
R12592 DVDD.n18044 DVDD.n507 4.5005
R12593 DVDD.n18044 DVDD.n513 4.5005
R12594 DVDD.n18044 DVDD.n506 4.5005
R12595 DVDD.n18044 DVDD.n514 4.5005
R12596 DVDD.n18044 DVDD.n505 4.5005
R12597 DVDD.n18044 DVDD.n515 4.5005
R12598 DVDD.n18044 DVDD.n504 4.5005
R12599 DVDD.n18044 DVDD.n516 4.5005
R12600 DVDD.n18044 DVDD.n18043 4.5005
R12601 DVDD.n18045 DVDD.n496 4.5005
R12602 DVDD.n18126 DVDD.n18045 4.5005
R12603 DVDD.n18059 DVDD.n18045 4.5005
R12604 DVDD.n18058 DVDD.n18045 4.5005
R12605 DVDD.n18062 DVDD.n18045 4.5005
R12606 DVDD.n18085 DVDD.n18045 4.5005
R12607 DVDD.n18063 DVDD.n18045 4.5005
R12608 DVDD.n501 DVDD.n496 4.5005
R12609 DVDD.n18126 DVDD.n501 4.5005
R12610 DVDD.n18059 DVDD.n501 4.5005
R12611 DVDD.n18058 DVDD.n501 4.5005
R12612 DVDD.n18061 DVDD.n501 4.5005
R12613 DVDD.n18057 DVDD.n501 4.5005
R12614 DVDD.n18062 DVDD.n501 4.5005
R12615 DVDD.n18063 DVDD.n501 4.5005
R12616 DVDD.n18046 DVDD.n496 4.5005
R12617 DVDD.n18126 DVDD.n18046 4.5005
R12618 DVDD.n18059 DVDD.n18046 4.5005
R12619 DVDD.n18058 DVDD.n18046 4.5005
R12620 DVDD.n18061 DVDD.n18046 4.5005
R12621 DVDD.n18057 DVDD.n18046 4.5005
R12622 DVDD.n18062 DVDD.n18046 4.5005
R12623 DVDD.n18063 DVDD.n18046 4.5005
R12624 DVDD.n500 DVDD.n496 4.5005
R12625 DVDD.n18126 DVDD.n500 4.5005
R12626 DVDD.n18059 DVDD.n500 4.5005
R12627 DVDD.n18058 DVDD.n500 4.5005
R12628 DVDD.n18061 DVDD.n500 4.5005
R12629 DVDD.n18057 DVDD.n500 4.5005
R12630 DVDD.n18062 DVDD.n500 4.5005
R12631 DVDD.n18063 DVDD.n500 4.5005
R12632 DVDD.n18047 DVDD.n496 4.5005
R12633 DVDD.n18126 DVDD.n18047 4.5005
R12634 DVDD.n18059 DVDD.n18047 4.5005
R12635 DVDD.n18058 DVDD.n18047 4.5005
R12636 DVDD.n18061 DVDD.n18047 4.5005
R12637 DVDD.n18062 DVDD.n18047 4.5005
R12638 DVDD.n18063 DVDD.n18047 4.5005
R12639 DVDD.n18054 DVDD.n18047 4.5005
R12640 DVDD.n499 DVDD.n496 4.5005
R12641 DVDD.n18126 DVDD.n499 4.5005
R12642 DVDD.n18059 DVDD.n499 4.5005
R12643 DVDD.n18058 DVDD.n499 4.5005
R12644 DVDD.n18061 DVDD.n499 4.5005
R12645 DVDD.n18062 DVDD.n499 4.5005
R12646 DVDD.n18063 DVDD.n499 4.5005
R12647 DVDD.n18048 DVDD.n496 4.5005
R12648 DVDD.n18126 DVDD.n18048 4.5005
R12649 DVDD.n18059 DVDD.n18048 4.5005
R12650 DVDD.n18058 DVDD.n18048 4.5005
R12651 DVDD.n18061 DVDD.n18048 4.5005
R12652 DVDD.n18057 DVDD.n18048 4.5005
R12653 DVDD.n18062 DVDD.n18048 4.5005
R12654 DVDD.n18063 DVDD.n18048 4.5005
R12655 DVDD.n498 DVDD.n496 4.5005
R12656 DVDD.n18126 DVDD.n498 4.5005
R12657 DVDD.n18059 DVDD.n498 4.5005
R12658 DVDD.n18058 DVDD.n498 4.5005
R12659 DVDD.n18061 DVDD.n498 4.5005
R12660 DVDD.n18057 DVDD.n498 4.5005
R12661 DVDD.n18062 DVDD.n498 4.5005
R12662 DVDD.n18063 DVDD.n498 4.5005
R12663 DVDD.n18049 DVDD.n496 4.5005
R12664 DVDD.n18126 DVDD.n18049 4.5005
R12665 DVDD.n18059 DVDD.n18049 4.5005
R12666 DVDD.n18058 DVDD.n18049 4.5005
R12667 DVDD.n18061 DVDD.n18049 4.5005
R12668 DVDD.n18057 DVDD.n18049 4.5005
R12669 DVDD.n18062 DVDD.n18049 4.5005
R12670 DVDD.n18063 DVDD.n18049 4.5005
R12671 DVDD.n497 DVDD.n496 4.5005
R12672 DVDD.n18126 DVDD.n497 4.5005
R12673 DVDD.n18059 DVDD.n497 4.5005
R12674 DVDD.n18058 DVDD.n497 4.5005
R12675 DVDD.n18061 DVDD.n497 4.5005
R12676 DVDD.n18057 DVDD.n497 4.5005
R12677 DVDD.n18062 DVDD.n497 4.5005
R12678 DVDD.n18063 DVDD.n497 4.5005
R12679 DVDD.n18125 DVDD.n496 4.5005
R12680 DVDD.n18126 DVDD.n18125 4.5005
R12681 DVDD.n18125 DVDD.n18059 4.5005
R12682 DVDD.n18125 DVDD.n18058 4.5005
R12683 DVDD.n18125 DVDD.n18061 4.5005
R12684 DVDD.n18125 DVDD.n18057 4.5005
R12685 DVDD.n18125 DVDD.n18062 4.5005
R12686 DVDD.n18125 DVDD.n18063 4.5005
R12687 DVDD.n18125 DVDD.n18054 4.5005
R12688 DVDD.n474 DVDD.n454 4.5005
R12689 DVDD.n474 DVDD.n453 4.5005
R12690 DVDD.n474 DVDD.n455 4.5005
R12691 DVDD.n474 DVDD.n452 4.5005
R12692 DVDD.n474 DVDD.n457 4.5005
R12693 DVDD.n474 DVDD.n450 4.5005
R12694 DVDD.n474 DVDD.n458 4.5005
R12695 DVDD.n474 DVDD.n449 4.5005
R12696 DVDD.n474 DVDD.n459 4.5005
R12697 DVDD.n474 DVDD.n448 4.5005
R12698 DVDD.n474 DVDD.n460 4.5005
R12699 DVDD.n18197 DVDD.n474 4.5005
R12700 DVDD.n18164 DVDD.n454 4.5005
R12701 DVDD.n18164 DVDD.n453 4.5005
R12702 DVDD.n18164 DVDD.n455 4.5005
R12703 DVDD.n18164 DVDD.n452 4.5005
R12704 DVDD.n18164 DVDD.n456 4.5005
R12705 DVDD.n18164 DVDD.n451 4.5005
R12706 DVDD.n18164 DVDD.n457 4.5005
R12707 DVDD.n18164 DVDD.n450 4.5005
R12708 DVDD.n18164 DVDD.n458 4.5005
R12709 DVDD.n18164 DVDD.n449 4.5005
R12710 DVDD.n18164 DVDD.n459 4.5005
R12711 DVDD.n18164 DVDD.n460 4.5005
R12712 DVDD.n18197 DVDD.n18164 4.5005
R12713 DVDD.n472 DVDD.n454 4.5005
R12714 DVDD.n472 DVDD.n453 4.5005
R12715 DVDD.n472 DVDD.n455 4.5005
R12716 DVDD.n472 DVDD.n452 4.5005
R12717 DVDD.n472 DVDD.n456 4.5005
R12718 DVDD.n472 DVDD.n451 4.5005
R12719 DVDD.n472 DVDD.n457 4.5005
R12720 DVDD.n472 DVDD.n450 4.5005
R12721 DVDD.n472 DVDD.n458 4.5005
R12722 DVDD.n472 DVDD.n449 4.5005
R12723 DVDD.n472 DVDD.n459 4.5005
R12724 DVDD.n472 DVDD.n460 4.5005
R12725 DVDD.n18197 DVDD.n472 4.5005
R12726 DVDD.n18166 DVDD.n454 4.5005
R12727 DVDD.n18166 DVDD.n453 4.5005
R12728 DVDD.n18166 DVDD.n455 4.5005
R12729 DVDD.n18166 DVDD.n452 4.5005
R12730 DVDD.n18166 DVDD.n456 4.5005
R12731 DVDD.n18166 DVDD.n451 4.5005
R12732 DVDD.n18166 DVDD.n457 4.5005
R12733 DVDD.n18166 DVDD.n450 4.5005
R12734 DVDD.n18166 DVDD.n458 4.5005
R12735 DVDD.n18166 DVDD.n449 4.5005
R12736 DVDD.n18166 DVDD.n459 4.5005
R12737 DVDD.n18166 DVDD.n460 4.5005
R12738 DVDD.n18197 DVDD.n18166 4.5005
R12739 DVDD.n471 DVDD.n454 4.5005
R12740 DVDD.n471 DVDD.n453 4.5005
R12741 DVDD.n471 DVDD.n455 4.5005
R12742 DVDD.n471 DVDD.n452 4.5005
R12743 DVDD.n471 DVDD.n456 4.5005
R12744 DVDD.n471 DVDD.n451 4.5005
R12745 DVDD.n471 DVDD.n457 4.5005
R12746 DVDD.n471 DVDD.n450 4.5005
R12747 DVDD.n471 DVDD.n458 4.5005
R12748 DVDD.n471 DVDD.n449 4.5005
R12749 DVDD.n471 DVDD.n459 4.5005
R12750 DVDD.n471 DVDD.n460 4.5005
R12751 DVDD.n18197 DVDD.n471 4.5005
R12752 DVDD.n18168 DVDD.n454 4.5005
R12753 DVDD.n18168 DVDD.n453 4.5005
R12754 DVDD.n18168 DVDD.n455 4.5005
R12755 DVDD.n18168 DVDD.n452 4.5005
R12756 DVDD.n18168 DVDD.n456 4.5005
R12757 DVDD.n18168 DVDD.n451 4.5005
R12758 DVDD.n18168 DVDD.n457 4.5005
R12759 DVDD.n18168 DVDD.n450 4.5005
R12760 DVDD.n18168 DVDD.n458 4.5005
R12761 DVDD.n18168 DVDD.n449 4.5005
R12762 DVDD.n18168 DVDD.n459 4.5005
R12763 DVDD.n18168 DVDD.n460 4.5005
R12764 DVDD.n18197 DVDD.n18168 4.5005
R12765 DVDD.n470 DVDD.n454 4.5005
R12766 DVDD.n470 DVDD.n453 4.5005
R12767 DVDD.n470 DVDD.n455 4.5005
R12768 DVDD.n470 DVDD.n452 4.5005
R12769 DVDD.n470 DVDD.n456 4.5005
R12770 DVDD.n470 DVDD.n451 4.5005
R12771 DVDD.n470 DVDD.n457 4.5005
R12772 DVDD.n470 DVDD.n450 4.5005
R12773 DVDD.n470 DVDD.n458 4.5005
R12774 DVDD.n470 DVDD.n449 4.5005
R12775 DVDD.n470 DVDD.n459 4.5005
R12776 DVDD.n470 DVDD.n460 4.5005
R12777 DVDD.n18197 DVDD.n470 4.5005
R12778 DVDD.n18170 DVDD.n454 4.5005
R12779 DVDD.n18170 DVDD.n453 4.5005
R12780 DVDD.n18170 DVDD.n455 4.5005
R12781 DVDD.n18170 DVDD.n452 4.5005
R12782 DVDD.n18170 DVDD.n456 4.5005
R12783 DVDD.n18170 DVDD.n451 4.5005
R12784 DVDD.n18170 DVDD.n457 4.5005
R12785 DVDD.n18170 DVDD.n450 4.5005
R12786 DVDD.n18170 DVDD.n458 4.5005
R12787 DVDD.n18170 DVDD.n449 4.5005
R12788 DVDD.n18170 DVDD.n459 4.5005
R12789 DVDD.n18170 DVDD.n460 4.5005
R12790 DVDD.n18197 DVDD.n18170 4.5005
R12791 DVDD.n469 DVDD.n454 4.5005
R12792 DVDD.n469 DVDD.n453 4.5005
R12793 DVDD.n469 DVDD.n455 4.5005
R12794 DVDD.n469 DVDD.n452 4.5005
R12795 DVDD.n469 DVDD.n456 4.5005
R12796 DVDD.n469 DVDD.n451 4.5005
R12797 DVDD.n469 DVDD.n457 4.5005
R12798 DVDD.n469 DVDD.n450 4.5005
R12799 DVDD.n469 DVDD.n458 4.5005
R12800 DVDD.n469 DVDD.n449 4.5005
R12801 DVDD.n469 DVDD.n459 4.5005
R12802 DVDD.n469 DVDD.n460 4.5005
R12803 DVDD.n18197 DVDD.n469 4.5005
R12804 DVDD.n18172 DVDD.n454 4.5005
R12805 DVDD.n18172 DVDD.n453 4.5005
R12806 DVDD.n18172 DVDD.n455 4.5005
R12807 DVDD.n18172 DVDD.n452 4.5005
R12808 DVDD.n18172 DVDD.n456 4.5005
R12809 DVDD.n18172 DVDD.n451 4.5005
R12810 DVDD.n18172 DVDD.n457 4.5005
R12811 DVDD.n18172 DVDD.n450 4.5005
R12812 DVDD.n18172 DVDD.n458 4.5005
R12813 DVDD.n18172 DVDD.n449 4.5005
R12814 DVDD.n18172 DVDD.n459 4.5005
R12815 DVDD.n18172 DVDD.n460 4.5005
R12816 DVDD.n18197 DVDD.n18172 4.5005
R12817 DVDD.n468 DVDD.n454 4.5005
R12818 DVDD.n468 DVDD.n453 4.5005
R12819 DVDD.n468 DVDD.n455 4.5005
R12820 DVDD.n468 DVDD.n452 4.5005
R12821 DVDD.n468 DVDD.n456 4.5005
R12822 DVDD.n468 DVDD.n451 4.5005
R12823 DVDD.n468 DVDD.n457 4.5005
R12824 DVDD.n468 DVDD.n450 4.5005
R12825 DVDD.n468 DVDD.n458 4.5005
R12826 DVDD.n468 DVDD.n449 4.5005
R12827 DVDD.n468 DVDD.n459 4.5005
R12828 DVDD.n468 DVDD.n460 4.5005
R12829 DVDD.n18197 DVDD.n468 4.5005
R12830 DVDD.n18174 DVDD.n454 4.5005
R12831 DVDD.n18174 DVDD.n453 4.5005
R12832 DVDD.n18174 DVDD.n455 4.5005
R12833 DVDD.n18174 DVDD.n452 4.5005
R12834 DVDD.n18174 DVDD.n456 4.5005
R12835 DVDD.n18174 DVDD.n451 4.5005
R12836 DVDD.n18174 DVDD.n457 4.5005
R12837 DVDD.n18174 DVDD.n450 4.5005
R12838 DVDD.n18174 DVDD.n458 4.5005
R12839 DVDD.n18174 DVDD.n449 4.5005
R12840 DVDD.n18174 DVDD.n459 4.5005
R12841 DVDD.n18174 DVDD.n460 4.5005
R12842 DVDD.n18197 DVDD.n18174 4.5005
R12843 DVDD.n467 DVDD.n454 4.5005
R12844 DVDD.n467 DVDD.n453 4.5005
R12845 DVDD.n467 DVDD.n455 4.5005
R12846 DVDD.n467 DVDD.n452 4.5005
R12847 DVDD.n467 DVDD.n456 4.5005
R12848 DVDD.n467 DVDD.n451 4.5005
R12849 DVDD.n467 DVDD.n457 4.5005
R12850 DVDD.n467 DVDD.n450 4.5005
R12851 DVDD.n467 DVDD.n458 4.5005
R12852 DVDD.n467 DVDD.n449 4.5005
R12853 DVDD.n467 DVDD.n459 4.5005
R12854 DVDD.n467 DVDD.n460 4.5005
R12855 DVDD.n18197 DVDD.n467 4.5005
R12856 DVDD.n18176 DVDD.n454 4.5005
R12857 DVDD.n18176 DVDD.n453 4.5005
R12858 DVDD.n18176 DVDD.n455 4.5005
R12859 DVDD.n18176 DVDD.n452 4.5005
R12860 DVDD.n18176 DVDD.n456 4.5005
R12861 DVDD.n18176 DVDD.n451 4.5005
R12862 DVDD.n18176 DVDD.n457 4.5005
R12863 DVDD.n18176 DVDD.n450 4.5005
R12864 DVDD.n18176 DVDD.n458 4.5005
R12865 DVDD.n18176 DVDD.n449 4.5005
R12866 DVDD.n18176 DVDD.n459 4.5005
R12867 DVDD.n18176 DVDD.n460 4.5005
R12868 DVDD.n18197 DVDD.n18176 4.5005
R12869 DVDD.n466 DVDD.n454 4.5005
R12870 DVDD.n466 DVDD.n453 4.5005
R12871 DVDD.n466 DVDD.n455 4.5005
R12872 DVDD.n466 DVDD.n452 4.5005
R12873 DVDD.n466 DVDD.n456 4.5005
R12874 DVDD.n466 DVDD.n451 4.5005
R12875 DVDD.n466 DVDD.n457 4.5005
R12876 DVDD.n466 DVDD.n450 4.5005
R12877 DVDD.n466 DVDD.n458 4.5005
R12878 DVDD.n466 DVDD.n449 4.5005
R12879 DVDD.n466 DVDD.n459 4.5005
R12880 DVDD.n466 DVDD.n460 4.5005
R12881 DVDD.n18197 DVDD.n466 4.5005
R12882 DVDD.n18178 DVDD.n454 4.5005
R12883 DVDD.n18178 DVDD.n453 4.5005
R12884 DVDD.n18178 DVDD.n455 4.5005
R12885 DVDD.n18178 DVDD.n452 4.5005
R12886 DVDD.n18178 DVDD.n456 4.5005
R12887 DVDD.n18178 DVDD.n451 4.5005
R12888 DVDD.n18178 DVDD.n457 4.5005
R12889 DVDD.n18178 DVDD.n450 4.5005
R12890 DVDD.n18178 DVDD.n458 4.5005
R12891 DVDD.n18178 DVDD.n449 4.5005
R12892 DVDD.n18178 DVDD.n459 4.5005
R12893 DVDD.n18178 DVDD.n460 4.5005
R12894 DVDD.n18197 DVDD.n18178 4.5005
R12895 DVDD.n465 DVDD.n454 4.5005
R12896 DVDD.n465 DVDD.n453 4.5005
R12897 DVDD.n465 DVDD.n455 4.5005
R12898 DVDD.n465 DVDD.n452 4.5005
R12899 DVDD.n465 DVDD.n456 4.5005
R12900 DVDD.n465 DVDD.n451 4.5005
R12901 DVDD.n465 DVDD.n457 4.5005
R12902 DVDD.n465 DVDD.n450 4.5005
R12903 DVDD.n465 DVDD.n458 4.5005
R12904 DVDD.n465 DVDD.n449 4.5005
R12905 DVDD.n465 DVDD.n459 4.5005
R12906 DVDD.n465 DVDD.n460 4.5005
R12907 DVDD.n18197 DVDD.n465 4.5005
R12908 DVDD.n18180 DVDD.n454 4.5005
R12909 DVDD.n18180 DVDD.n453 4.5005
R12910 DVDD.n18180 DVDD.n455 4.5005
R12911 DVDD.n18180 DVDD.n452 4.5005
R12912 DVDD.n18180 DVDD.n456 4.5005
R12913 DVDD.n18180 DVDD.n451 4.5005
R12914 DVDD.n18180 DVDD.n457 4.5005
R12915 DVDD.n18180 DVDD.n450 4.5005
R12916 DVDD.n18180 DVDD.n458 4.5005
R12917 DVDD.n18180 DVDD.n449 4.5005
R12918 DVDD.n18180 DVDD.n459 4.5005
R12919 DVDD.n18180 DVDD.n460 4.5005
R12920 DVDD.n18197 DVDD.n18180 4.5005
R12921 DVDD.n464 DVDD.n454 4.5005
R12922 DVDD.n464 DVDD.n453 4.5005
R12923 DVDD.n464 DVDD.n455 4.5005
R12924 DVDD.n464 DVDD.n452 4.5005
R12925 DVDD.n464 DVDD.n456 4.5005
R12926 DVDD.n464 DVDD.n451 4.5005
R12927 DVDD.n464 DVDD.n457 4.5005
R12928 DVDD.n464 DVDD.n450 4.5005
R12929 DVDD.n464 DVDD.n458 4.5005
R12930 DVDD.n464 DVDD.n449 4.5005
R12931 DVDD.n464 DVDD.n459 4.5005
R12932 DVDD.n464 DVDD.n460 4.5005
R12933 DVDD.n18197 DVDD.n464 4.5005
R12934 DVDD.n18182 DVDD.n454 4.5005
R12935 DVDD.n18182 DVDD.n453 4.5005
R12936 DVDD.n18182 DVDD.n455 4.5005
R12937 DVDD.n18182 DVDD.n452 4.5005
R12938 DVDD.n18182 DVDD.n456 4.5005
R12939 DVDD.n18182 DVDD.n451 4.5005
R12940 DVDD.n18182 DVDD.n457 4.5005
R12941 DVDD.n18182 DVDD.n450 4.5005
R12942 DVDD.n18182 DVDD.n458 4.5005
R12943 DVDD.n18182 DVDD.n449 4.5005
R12944 DVDD.n18182 DVDD.n459 4.5005
R12945 DVDD.n18182 DVDD.n460 4.5005
R12946 DVDD.n18197 DVDD.n18182 4.5005
R12947 DVDD.n463 DVDD.n454 4.5005
R12948 DVDD.n463 DVDD.n453 4.5005
R12949 DVDD.n463 DVDD.n455 4.5005
R12950 DVDD.n463 DVDD.n452 4.5005
R12951 DVDD.n463 DVDD.n456 4.5005
R12952 DVDD.n463 DVDD.n451 4.5005
R12953 DVDD.n463 DVDD.n457 4.5005
R12954 DVDD.n463 DVDD.n450 4.5005
R12955 DVDD.n463 DVDD.n458 4.5005
R12956 DVDD.n463 DVDD.n449 4.5005
R12957 DVDD.n463 DVDD.n459 4.5005
R12958 DVDD.n463 DVDD.n460 4.5005
R12959 DVDD.n18197 DVDD.n463 4.5005
R12960 DVDD.n18196 DVDD.n454 4.5005
R12961 DVDD.n18196 DVDD.n453 4.5005
R12962 DVDD.n18196 DVDD.n455 4.5005
R12963 DVDD.n18196 DVDD.n452 4.5005
R12964 DVDD.n18196 DVDD.n456 4.5005
R12965 DVDD.n18196 DVDD.n451 4.5005
R12966 DVDD.n18196 DVDD.n457 4.5005
R12967 DVDD.n18196 DVDD.n450 4.5005
R12968 DVDD.n18196 DVDD.n458 4.5005
R12969 DVDD.n18196 DVDD.n449 4.5005
R12970 DVDD.n18196 DVDD.n459 4.5005
R12971 DVDD.n18196 DVDD.n460 4.5005
R12972 DVDD.n18197 DVDD.n18196 4.5005
R12973 DVDD.n462 DVDD.n454 4.5005
R12974 DVDD.n462 DVDD.n453 4.5005
R12975 DVDD.n462 DVDD.n455 4.5005
R12976 DVDD.n462 DVDD.n452 4.5005
R12977 DVDD.n462 DVDD.n456 4.5005
R12978 DVDD.n462 DVDD.n451 4.5005
R12979 DVDD.n462 DVDD.n457 4.5005
R12980 DVDD.n462 DVDD.n450 4.5005
R12981 DVDD.n462 DVDD.n458 4.5005
R12982 DVDD.n462 DVDD.n449 4.5005
R12983 DVDD.n462 DVDD.n459 4.5005
R12984 DVDD.n462 DVDD.n460 4.5005
R12985 DVDD.n18197 DVDD.n462 4.5005
R12986 DVDD.n18198 DVDD.n454 4.5005
R12987 DVDD.n18198 DVDD.n453 4.5005
R12988 DVDD.n18198 DVDD.n455 4.5005
R12989 DVDD.n18198 DVDD.n452 4.5005
R12990 DVDD.n18198 DVDD.n456 4.5005
R12991 DVDD.n18198 DVDD.n451 4.5005
R12992 DVDD.n18198 DVDD.n457 4.5005
R12993 DVDD.n18198 DVDD.n450 4.5005
R12994 DVDD.n18198 DVDD.n458 4.5005
R12995 DVDD.n18198 DVDD.n449 4.5005
R12996 DVDD.n18198 DVDD.n459 4.5005
R12997 DVDD.n18198 DVDD.n448 4.5005
R12998 DVDD.n18198 DVDD.n460 4.5005
R12999 DVDD.n18198 DVDD.n18197 4.5005
R13000 DVDD.n18199 DVDD.n435 4.5005
R13001 DVDD.n18199 DVDD.n440 4.5005
R13002 DVDD.n22122 DVDD.n18199 4.5005
R13003 DVDD.n22074 DVDD.n18199 4.5005
R13004 DVDD.n22077 DVDD.n18199 4.5005
R13005 DVDD.n22072 DVDD.n18199 4.5005
R13006 DVDD.n22078 DVDD.n18199 4.5005
R13007 DVDD.n22071 DVDD.n18199 4.5005
R13008 DVDD.n22079 DVDD.n18199 4.5005
R13009 DVDD.n22114 DVDD.n18199 4.5005
R13010 DVDD.n22115 DVDD.n18199 4.5005
R13011 DVDD.n22120 DVDD.n18199 4.5005
R13012 DVDD.n445 DVDD.n435 4.5005
R13013 DVDD.n445 DVDD.n440 4.5005
R13014 DVDD.n22122 DVDD.n445 4.5005
R13015 DVDD.n22074 DVDD.n445 4.5005
R13016 DVDD.n22076 DVDD.n445 4.5005
R13017 DVDD.n22073 DVDD.n445 4.5005
R13018 DVDD.n22077 DVDD.n445 4.5005
R13019 DVDD.n22072 DVDD.n445 4.5005
R13020 DVDD.n22078 DVDD.n445 4.5005
R13021 DVDD.n22071 DVDD.n445 4.5005
R13022 DVDD.n22079 DVDD.n445 4.5005
R13023 DVDD.n22115 DVDD.n445 4.5005
R13024 DVDD.n22120 DVDD.n445 4.5005
R13025 DVDD.n18200 DVDD.n435 4.5005
R13026 DVDD.n18200 DVDD.n440 4.5005
R13027 DVDD.n22122 DVDD.n18200 4.5005
R13028 DVDD.n22074 DVDD.n18200 4.5005
R13029 DVDD.n22076 DVDD.n18200 4.5005
R13030 DVDD.n22073 DVDD.n18200 4.5005
R13031 DVDD.n22077 DVDD.n18200 4.5005
R13032 DVDD.n22072 DVDD.n18200 4.5005
R13033 DVDD.n22078 DVDD.n18200 4.5005
R13034 DVDD.n22071 DVDD.n18200 4.5005
R13035 DVDD.n22079 DVDD.n18200 4.5005
R13036 DVDD.n22115 DVDD.n18200 4.5005
R13037 DVDD.n22120 DVDD.n18200 4.5005
R13038 DVDD.n444 DVDD.n435 4.5005
R13039 DVDD.n444 DVDD.n440 4.5005
R13040 DVDD.n22122 DVDD.n444 4.5005
R13041 DVDD.n22074 DVDD.n444 4.5005
R13042 DVDD.n22076 DVDD.n444 4.5005
R13043 DVDD.n22073 DVDD.n444 4.5005
R13044 DVDD.n22077 DVDD.n444 4.5005
R13045 DVDD.n22072 DVDD.n444 4.5005
R13046 DVDD.n22078 DVDD.n444 4.5005
R13047 DVDD.n22071 DVDD.n444 4.5005
R13048 DVDD.n22079 DVDD.n444 4.5005
R13049 DVDD.n22115 DVDD.n444 4.5005
R13050 DVDD.n22120 DVDD.n444 4.5005
R13051 DVDD.n18201 DVDD.n435 4.5005
R13052 DVDD.n18201 DVDD.n440 4.5005
R13053 DVDD.n22122 DVDD.n18201 4.5005
R13054 DVDD.n22074 DVDD.n18201 4.5005
R13055 DVDD.n22076 DVDD.n18201 4.5005
R13056 DVDD.n22073 DVDD.n18201 4.5005
R13057 DVDD.n22077 DVDD.n18201 4.5005
R13058 DVDD.n22072 DVDD.n18201 4.5005
R13059 DVDD.n22078 DVDD.n18201 4.5005
R13060 DVDD.n22071 DVDD.n18201 4.5005
R13061 DVDD.n22079 DVDD.n18201 4.5005
R13062 DVDD.n22115 DVDD.n18201 4.5005
R13063 DVDD.n22120 DVDD.n18201 4.5005
R13064 DVDD.n443 DVDD.n435 4.5005
R13065 DVDD.n443 DVDD.n440 4.5005
R13066 DVDD.n22122 DVDD.n443 4.5005
R13067 DVDD.n22074 DVDD.n443 4.5005
R13068 DVDD.n22076 DVDD.n443 4.5005
R13069 DVDD.n22073 DVDD.n443 4.5005
R13070 DVDD.n22077 DVDD.n443 4.5005
R13071 DVDD.n22072 DVDD.n443 4.5005
R13072 DVDD.n22078 DVDD.n443 4.5005
R13073 DVDD.n22071 DVDD.n443 4.5005
R13074 DVDD.n22079 DVDD.n443 4.5005
R13075 DVDD.n22115 DVDD.n443 4.5005
R13076 DVDD.n22120 DVDD.n443 4.5005
R13077 DVDD.n18202 DVDD.n435 4.5005
R13078 DVDD.n18202 DVDD.n440 4.5005
R13079 DVDD.n22122 DVDD.n18202 4.5005
R13080 DVDD.n22074 DVDD.n18202 4.5005
R13081 DVDD.n22076 DVDD.n18202 4.5005
R13082 DVDD.n22073 DVDD.n18202 4.5005
R13083 DVDD.n22077 DVDD.n18202 4.5005
R13084 DVDD.n22072 DVDD.n18202 4.5005
R13085 DVDD.n22078 DVDD.n18202 4.5005
R13086 DVDD.n22071 DVDD.n18202 4.5005
R13087 DVDD.n22079 DVDD.n18202 4.5005
R13088 DVDD.n22115 DVDD.n18202 4.5005
R13089 DVDD.n22120 DVDD.n18202 4.5005
R13090 DVDD.n442 DVDD.n435 4.5005
R13091 DVDD.n442 DVDD.n440 4.5005
R13092 DVDD.n22122 DVDD.n442 4.5005
R13093 DVDD.n22074 DVDD.n442 4.5005
R13094 DVDD.n22076 DVDD.n442 4.5005
R13095 DVDD.n22073 DVDD.n442 4.5005
R13096 DVDD.n22077 DVDD.n442 4.5005
R13097 DVDD.n22072 DVDD.n442 4.5005
R13098 DVDD.n22078 DVDD.n442 4.5005
R13099 DVDD.n22071 DVDD.n442 4.5005
R13100 DVDD.n22079 DVDD.n442 4.5005
R13101 DVDD.n22115 DVDD.n442 4.5005
R13102 DVDD.n22120 DVDD.n442 4.5005
R13103 DVDD.n18203 DVDD.n435 4.5005
R13104 DVDD.n18203 DVDD.n440 4.5005
R13105 DVDD.n22122 DVDD.n18203 4.5005
R13106 DVDD.n22074 DVDD.n18203 4.5005
R13107 DVDD.n22076 DVDD.n18203 4.5005
R13108 DVDD.n22073 DVDD.n18203 4.5005
R13109 DVDD.n22077 DVDD.n18203 4.5005
R13110 DVDD.n22072 DVDD.n18203 4.5005
R13111 DVDD.n22078 DVDD.n18203 4.5005
R13112 DVDD.n22071 DVDD.n18203 4.5005
R13113 DVDD.n22079 DVDD.n18203 4.5005
R13114 DVDD.n22115 DVDD.n18203 4.5005
R13115 DVDD.n22120 DVDD.n18203 4.5005
R13116 DVDD.n441 DVDD.n435 4.5005
R13117 DVDD.n441 DVDD.n440 4.5005
R13118 DVDD.n22122 DVDD.n441 4.5005
R13119 DVDD.n22074 DVDD.n441 4.5005
R13120 DVDD.n22076 DVDD.n441 4.5005
R13121 DVDD.n22073 DVDD.n441 4.5005
R13122 DVDD.n22077 DVDD.n441 4.5005
R13123 DVDD.n22072 DVDD.n441 4.5005
R13124 DVDD.n22078 DVDD.n441 4.5005
R13125 DVDD.n22071 DVDD.n441 4.5005
R13126 DVDD.n22079 DVDD.n441 4.5005
R13127 DVDD.n22115 DVDD.n441 4.5005
R13128 DVDD.n22120 DVDD.n441 4.5005
R13129 DVDD.n22121 DVDD.n435 4.5005
R13130 DVDD.n22121 DVDD.n440 4.5005
R13131 DVDD.n22122 DVDD.n22121 4.5005
R13132 DVDD.n22121 DVDD.n22074 4.5005
R13133 DVDD.n22121 DVDD.n22076 4.5005
R13134 DVDD.n22121 DVDD.n22073 4.5005
R13135 DVDD.n22121 DVDD.n22077 4.5005
R13136 DVDD.n22121 DVDD.n22072 4.5005
R13137 DVDD.n22121 DVDD.n22078 4.5005
R13138 DVDD.n22121 DVDD.n22071 4.5005
R13139 DVDD.n22121 DVDD.n22079 4.5005
R13140 DVDD.n22121 DVDD.n22120 4.5005
R13141 DVDD.n18981 DVDD.n18966 4.5005
R13142 DVDD.n18981 DVDD.n18965 4.5005
R13143 DVDD.n18981 DVDD.n18967 4.5005
R13144 DVDD.n18981 DVDD.n18964 4.5005
R13145 DVDD.n18981 DVDD.n18969 4.5005
R13146 DVDD.n18981 DVDD.n18962 4.5005
R13147 DVDD.n18981 DVDD.n18970 4.5005
R13148 DVDD.n18981 DVDD.n18961 4.5005
R13149 DVDD.n18981 DVDD.n18971 4.5005
R13150 DVDD.n18995 DVDD.n18981 4.5005
R13151 DVDD.n20852 DVDD.n18981 4.5005
R13152 DVDD.n20854 DVDD.n18981 4.5005
R13153 DVDD.n18978 DVDD.n18966 4.5005
R13154 DVDD.n18978 DVDD.n18965 4.5005
R13155 DVDD.n18978 DVDD.n18967 4.5005
R13156 DVDD.n18978 DVDD.n18964 4.5005
R13157 DVDD.n18978 DVDD.n18968 4.5005
R13158 DVDD.n18978 DVDD.n18963 4.5005
R13159 DVDD.n18978 DVDD.n18969 4.5005
R13160 DVDD.n18978 DVDD.n18962 4.5005
R13161 DVDD.n18978 DVDD.n18970 4.5005
R13162 DVDD.n18978 DVDD.n18961 4.5005
R13163 DVDD.n18978 DVDD.n18971 4.5005
R13164 DVDD.n20852 DVDD.n18978 4.5005
R13165 DVDD.n20854 DVDD.n18978 4.5005
R13166 DVDD.n18982 DVDD.n18966 4.5005
R13167 DVDD.n18982 DVDD.n18965 4.5005
R13168 DVDD.n18982 DVDD.n18967 4.5005
R13169 DVDD.n18982 DVDD.n18964 4.5005
R13170 DVDD.n18982 DVDD.n18968 4.5005
R13171 DVDD.n18982 DVDD.n18963 4.5005
R13172 DVDD.n18982 DVDD.n18969 4.5005
R13173 DVDD.n18982 DVDD.n18962 4.5005
R13174 DVDD.n18982 DVDD.n18970 4.5005
R13175 DVDD.n18982 DVDD.n18961 4.5005
R13176 DVDD.n18982 DVDD.n18971 4.5005
R13177 DVDD.n20852 DVDD.n18982 4.5005
R13178 DVDD.n20854 DVDD.n18982 4.5005
R13179 DVDD.n18977 DVDD.n18966 4.5005
R13180 DVDD.n18977 DVDD.n18965 4.5005
R13181 DVDD.n18977 DVDD.n18967 4.5005
R13182 DVDD.n18977 DVDD.n18964 4.5005
R13183 DVDD.n18977 DVDD.n18968 4.5005
R13184 DVDD.n18977 DVDD.n18963 4.5005
R13185 DVDD.n18977 DVDD.n18969 4.5005
R13186 DVDD.n18977 DVDD.n18962 4.5005
R13187 DVDD.n18977 DVDD.n18970 4.5005
R13188 DVDD.n18977 DVDD.n18961 4.5005
R13189 DVDD.n18977 DVDD.n18971 4.5005
R13190 DVDD.n20852 DVDD.n18977 4.5005
R13191 DVDD.n20854 DVDD.n18977 4.5005
R13192 DVDD.n18983 DVDD.n18966 4.5005
R13193 DVDD.n18983 DVDD.n18965 4.5005
R13194 DVDD.n18983 DVDD.n18967 4.5005
R13195 DVDD.n18983 DVDD.n18964 4.5005
R13196 DVDD.n18983 DVDD.n18968 4.5005
R13197 DVDD.n18983 DVDD.n18963 4.5005
R13198 DVDD.n18983 DVDD.n18969 4.5005
R13199 DVDD.n18983 DVDD.n18962 4.5005
R13200 DVDD.n18983 DVDD.n18970 4.5005
R13201 DVDD.n18983 DVDD.n18961 4.5005
R13202 DVDD.n18983 DVDD.n18971 4.5005
R13203 DVDD.n20852 DVDD.n18983 4.5005
R13204 DVDD.n20854 DVDD.n18983 4.5005
R13205 DVDD.n18976 DVDD.n18966 4.5005
R13206 DVDD.n18976 DVDD.n18965 4.5005
R13207 DVDD.n18976 DVDD.n18967 4.5005
R13208 DVDD.n18976 DVDD.n18964 4.5005
R13209 DVDD.n18976 DVDD.n18968 4.5005
R13210 DVDD.n18976 DVDD.n18963 4.5005
R13211 DVDD.n18976 DVDD.n18969 4.5005
R13212 DVDD.n18976 DVDD.n18962 4.5005
R13213 DVDD.n18976 DVDD.n18970 4.5005
R13214 DVDD.n18976 DVDD.n18961 4.5005
R13215 DVDD.n18976 DVDD.n18971 4.5005
R13216 DVDD.n20852 DVDD.n18976 4.5005
R13217 DVDD.n20854 DVDD.n18976 4.5005
R13218 DVDD.n18984 DVDD.n18966 4.5005
R13219 DVDD.n18984 DVDD.n18965 4.5005
R13220 DVDD.n18984 DVDD.n18967 4.5005
R13221 DVDD.n18984 DVDD.n18964 4.5005
R13222 DVDD.n18984 DVDD.n18968 4.5005
R13223 DVDD.n18984 DVDD.n18963 4.5005
R13224 DVDD.n18984 DVDD.n18969 4.5005
R13225 DVDD.n18984 DVDD.n18962 4.5005
R13226 DVDD.n18984 DVDD.n18970 4.5005
R13227 DVDD.n18984 DVDD.n18961 4.5005
R13228 DVDD.n18984 DVDD.n18971 4.5005
R13229 DVDD.n20852 DVDD.n18984 4.5005
R13230 DVDD.n20854 DVDD.n18984 4.5005
R13231 DVDD.n18975 DVDD.n18966 4.5005
R13232 DVDD.n18975 DVDD.n18965 4.5005
R13233 DVDD.n18975 DVDD.n18967 4.5005
R13234 DVDD.n18975 DVDD.n18964 4.5005
R13235 DVDD.n18975 DVDD.n18968 4.5005
R13236 DVDD.n18975 DVDD.n18963 4.5005
R13237 DVDD.n18975 DVDD.n18969 4.5005
R13238 DVDD.n18975 DVDD.n18962 4.5005
R13239 DVDD.n18975 DVDD.n18970 4.5005
R13240 DVDD.n18975 DVDD.n18961 4.5005
R13241 DVDD.n18975 DVDD.n18971 4.5005
R13242 DVDD.n20852 DVDD.n18975 4.5005
R13243 DVDD.n20854 DVDD.n18975 4.5005
R13244 DVDD.n20853 DVDD.n18966 4.5005
R13245 DVDD.n20853 DVDD.n18965 4.5005
R13246 DVDD.n20853 DVDD.n18967 4.5005
R13247 DVDD.n20853 DVDD.n18964 4.5005
R13248 DVDD.n20853 DVDD.n18968 4.5005
R13249 DVDD.n20853 DVDD.n18963 4.5005
R13250 DVDD.n20853 DVDD.n18969 4.5005
R13251 DVDD.n20853 DVDD.n18962 4.5005
R13252 DVDD.n20853 DVDD.n18970 4.5005
R13253 DVDD.n20853 DVDD.n18961 4.5005
R13254 DVDD.n20853 DVDD.n18971 4.5005
R13255 DVDD.n20853 DVDD.n20852 4.5005
R13256 DVDD.n20854 DVDD.n20853 4.5005
R13257 DVDD.n18974 DVDD.n18966 4.5005
R13258 DVDD.n18974 DVDD.n18965 4.5005
R13259 DVDD.n18974 DVDD.n18967 4.5005
R13260 DVDD.n18974 DVDD.n18964 4.5005
R13261 DVDD.n18974 DVDD.n18968 4.5005
R13262 DVDD.n18974 DVDD.n18963 4.5005
R13263 DVDD.n18974 DVDD.n18969 4.5005
R13264 DVDD.n18974 DVDD.n18962 4.5005
R13265 DVDD.n18974 DVDD.n18970 4.5005
R13266 DVDD.n18974 DVDD.n18961 4.5005
R13267 DVDD.n18974 DVDD.n18971 4.5005
R13268 DVDD.n20852 DVDD.n18974 4.5005
R13269 DVDD.n20854 DVDD.n18974 4.5005
R13270 DVDD.n20855 DVDD.n18966 4.5005
R13271 DVDD.n20855 DVDD.n18965 4.5005
R13272 DVDD.n20855 DVDD.n18967 4.5005
R13273 DVDD.n20855 DVDD.n18964 4.5005
R13274 DVDD.n20855 DVDD.n18968 4.5005
R13275 DVDD.n20855 DVDD.n18963 4.5005
R13276 DVDD.n20855 DVDD.n18969 4.5005
R13277 DVDD.n20855 DVDD.n18962 4.5005
R13278 DVDD.n20855 DVDD.n18970 4.5005
R13279 DVDD.n20855 DVDD.n18961 4.5005
R13280 DVDD.n20855 DVDD.n18971 4.5005
R13281 DVDD.n20855 DVDD.n20854 4.5005
R13282 DVDD.n18953 DVDD.n18938 4.5005
R13283 DVDD.n18953 DVDD.n18936 4.5005
R13284 DVDD.n18953 DVDD.n18939 4.5005
R13285 DVDD.n18953 DVDD.n18935 4.5005
R13286 DVDD.n18953 DVDD.n18941 4.5005
R13287 DVDD.n18953 DVDD.n18933 4.5005
R13288 DVDD.n18953 DVDD.n18942 4.5005
R13289 DVDD.n18953 DVDD.n18932 4.5005
R13290 DVDD.n18953 DVDD.n18943 4.5005
R13291 DVDD.n18953 DVDD.n18931 4.5005
R13292 DVDD.n20883 DVDD.n18953 4.5005
R13293 DVDD.n18949 DVDD.n18938 4.5005
R13294 DVDD.n18949 DVDD.n18936 4.5005
R13295 DVDD.n18949 DVDD.n18939 4.5005
R13296 DVDD.n18949 DVDD.n18935 4.5005
R13297 DVDD.n18949 DVDD.n18940 4.5005
R13298 DVDD.n18949 DVDD.n18934 4.5005
R13299 DVDD.n18949 DVDD.n18941 4.5005
R13300 DVDD.n18949 DVDD.n18933 4.5005
R13301 DVDD.n18949 DVDD.n18942 4.5005
R13302 DVDD.n18949 DVDD.n18932 4.5005
R13303 DVDD.n18949 DVDD.n18943 4.5005
R13304 DVDD.n18949 DVDD.n18931 4.5005
R13305 DVDD.n18949 DVDD.n18944 4.5005
R13306 DVDD.n18949 DVDD.n18930 4.5005
R13307 DVDD.n20883 DVDD.n18949 4.5005
R13308 DVDD.n18954 DVDD.n18938 4.5005
R13309 DVDD.n18954 DVDD.n18936 4.5005
R13310 DVDD.n18954 DVDD.n18939 4.5005
R13311 DVDD.n18954 DVDD.n18935 4.5005
R13312 DVDD.n18954 DVDD.n18940 4.5005
R13313 DVDD.n18954 DVDD.n18934 4.5005
R13314 DVDD.n18954 DVDD.n18941 4.5005
R13315 DVDD.n18954 DVDD.n18933 4.5005
R13316 DVDD.n18954 DVDD.n18942 4.5005
R13317 DVDD.n18954 DVDD.n18932 4.5005
R13318 DVDD.n18954 DVDD.n18943 4.5005
R13319 DVDD.n18954 DVDD.n18931 4.5005
R13320 DVDD.n18954 DVDD.n18944 4.5005
R13321 DVDD.n18954 DVDD.n18930 4.5005
R13322 DVDD.n20883 DVDD.n18954 4.5005
R13323 DVDD.n18948 DVDD.n18938 4.5005
R13324 DVDD.n18948 DVDD.n18936 4.5005
R13325 DVDD.n18948 DVDD.n18939 4.5005
R13326 DVDD.n18948 DVDD.n18935 4.5005
R13327 DVDD.n18948 DVDD.n18940 4.5005
R13328 DVDD.n18948 DVDD.n18934 4.5005
R13329 DVDD.n18948 DVDD.n18941 4.5005
R13330 DVDD.n18948 DVDD.n18933 4.5005
R13331 DVDD.n18948 DVDD.n18942 4.5005
R13332 DVDD.n18948 DVDD.n18932 4.5005
R13333 DVDD.n18948 DVDD.n18943 4.5005
R13334 DVDD.n18948 DVDD.n18931 4.5005
R13335 DVDD.n18948 DVDD.n18944 4.5005
R13336 DVDD.n18948 DVDD.n18930 4.5005
R13337 DVDD.n20883 DVDD.n18948 4.5005
R13338 DVDD.n18955 DVDD.n18938 4.5005
R13339 DVDD.n18955 DVDD.n18936 4.5005
R13340 DVDD.n18955 DVDD.n18939 4.5005
R13341 DVDD.n18955 DVDD.n18935 4.5005
R13342 DVDD.n18955 DVDD.n18940 4.5005
R13343 DVDD.n18955 DVDD.n18934 4.5005
R13344 DVDD.n18955 DVDD.n18941 4.5005
R13345 DVDD.n18955 DVDD.n18933 4.5005
R13346 DVDD.n18955 DVDD.n18942 4.5005
R13347 DVDD.n18955 DVDD.n18932 4.5005
R13348 DVDD.n18955 DVDD.n18943 4.5005
R13349 DVDD.n18955 DVDD.n18931 4.5005
R13350 DVDD.n18955 DVDD.n18944 4.5005
R13351 DVDD.n18955 DVDD.n18930 4.5005
R13352 DVDD.n20883 DVDD.n18955 4.5005
R13353 DVDD.n18947 DVDD.n18938 4.5005
R13354 DVDD.n18947 DVDD.n18936 4.5005
R13355 DVDD.n18947 DVDD.n18939 4.5005
R13356 DVDD.n18947 DVDD.n18935 4.5005
R13357 DVDD.n18947 DVDD.n18940 4.5005
R13358 DVDD.n18947 DVDD.n18934 4.5005
R13359 DVDD.n18947 DVDD.n18941 4.5005
R13360 DVDD.n18947 DVDD.n18933 4.5005
R13361 DVDD.n18947 DVDD.n18942 4.5005
R13362 DVDD.n18947 DVDD.n18932 4.5005
R13363 DVDD.n18947 DVDD.n18943 4.5005
R13364 DVDD.n18947 DVDD.n18931 4.5005
R13365 DVDD.n18947 DVDD.n18944 4.5005
R13366 DVDD.n18947 DVDD.n18930 4.5005
R13367 DVDD.n20883 DVDD.n18947 4.5005
R13368 DVDD.n18956 DVDD.n18938 4.5005
R13369 DVDD.n18956 DVDD.n18936 4.5005
R13370 DVDD.n18956 DVDD.n18939 4.5005
R13371 DVDD.n18956 DVDD.n18935 4.5005
R13372 DVDD.n18956 DVDD.n18940 4.5005
R13373 DVDD.n18956 DVDD.n18934 4.5005
R13374 DVDD.n18956 DVDD.n18941 4.5005
R13375 DVDD.n18956 DVDD.n18933 4.5005
R13376 DVDD.n18956 DVDD.n18942 4.5005
R13377 DVDD.n18956 DVDD.n18932 4.5005
R13378 DVDD.n18956 DVDD.n18943 4.5005
R13379 DVDD.n18956 DVDD.n18931 4.5005
R13380 DVDD.n18956 DVDD.n18944 4.5005
R13381 DVDD.n18956 DVDD.n18930 4.5005
R13382 DVDD.n20883 DVDD.n18956 4.5005
R13383 DVDD.n18946 DVDD.n18938 4.5005
R13384 DVDD.n18946 DVDD.n18936 4.5005
R13385 DVDD.n18946 DVDD.n18939 4.5005
R13386 DVDD.n18946 DVDD.n18935 4.5005
R13387 DVDD.n18946 DVDD.n18940 4.5005
R13388 DVDD.n18946 DVDD.n18934 4.5005
R13389 DVDD.n18946 DVDD.n18941 4.5005
R13390 DVDD.n18946 DVDD.n18933 4.5005
R13391 DVDD.n18946 DVDD.n18942 4.5005
R13392 DVDD.n18946 DVDD.n18932 4.5005
R13393 DVDD.n18946 DVDD.n18943 4.5005
R13394 DVDD.n18946 DVDD.n18931 4.5005
R13395 DVDD.n18946 DVDD.n18944 4.5005
R13396 DVDD.n18946 DVDD.n18930 4.5005
R13397 DVDD.n20883 DVDD.n18946 4.5005
R13398 DVDD.n20882 DVDD.n18938 4.5005
R13399 DVDD.n20882 DVDD.n18936 4.5005
R13400 DVDD.n20882 DVDD.n18939 4.5005
R13401 DVDD.n20882 DVDD.n18935 4.5005
R13402 DVDD.n20882 DVDD.n18940 4.5005
R13403 DVDD.n20882 DVDD.n18934 4.5005
R13404 DVDD.n20882 DVDD.n18941 4.5005
R13405 DVDD.n20882 DVDD.n18933 4.5005
R13406 DVDD.n20882 DVDD.n18942 4.5005
R13407 DVDD.n20882 DVDD.n18932 4.5005
R13408 DVDD.n20882 DVDD.n18943 4.5005
R13409 DVDD.n20882 DVDD.n18931 4.5005
R13410 DVDD.n20882 DVDD.n18944 4.5005
R13411 DVDD.n20882 DVDD.n18930 4.5005
R13412 DVDD.n20883 DVDD.n20882 4.5005
R13413 DVDD.n20884 DVDD.n18938 4.5005
R13414 DVDD.n20884 DVDD.n18936 4.5005
R13415 DVDD.n20884 DVDD.n18939 4.5005
R13416 DVDD.n20884 DVDD.n18935 4.5005
R13417 DVDD.n20884 DVDD.n18940 4.5005
R13418 DVDD.n20884 DVDD.n18934 4.5005
R13419 DVDD.n20884 DVDD.n18941 4.5005
R13420 DVDD.n20884 DVDD.n18933 4.5005
R13421 DVDD.n20884 DVDD.n18942 4.5005
R13422 DVDD.n20884 DVDD.n18932 4.5005
R13423 DVDD.n20884 DVDD.n18943 4.5005
R13424 DVDD.n20884 DVDD.n18931 4.5005
R13425 DVDD.n20884 DVDD.n18944 4.5005
R13426 DVDD.n20884 DVDD.n18930 4.5005
R13427 DVDD.n20884 DVDD.n20883 4.5005
R13428 DVDD.n18938 DVDD.n18929 4.5005
R13429 DVDD.n18936 DVDD.n18929 4.5005
R13430 DVDD.n18939 DVDD.n18929 4.5005
R13431 DVDD.n18935 DVDD.n18929 4.5005
R13432 DVDD.n18940 DVDD.n18929 4.5005
R13433 DVDD.n18934 DVDD.n18929 4.5005
R13434 DVDD.n18941 DVDD.n18929 4.5005
R13435 DVDD.n18933 DVDD.n18929 4.5005
R13436 DVDD.n18942 DVDD.n18929 4.5005
R13437 DVDD.n18932 DVDD.n18929 4.5005
R13438 DVDD.n18943 DVDD.n18929 4.5005
R13439 DVDD.n18931 DVDD.n18929 4.5005
R13440 DVDD.n18944 DVDD.n18929 4.5005
R13441 DVDD.n18930 DVDD.n18929 4.5005
R13442 DVDD.n20883 DVDD.n18929 4.5005
R13443 DVDD.n18037 DVDD.n506 4.5005
R13444 DVDD.n18037 DVDD.n513 4.5005
R13445 DVDD.n18037 DVDD.n507 4.5005
R13446 DVDD.n18037 DVDD.n512 4.5005
R13447 DVDD.n18037 DVDD.n508 4.5005
R13448 DVDD.n18037 DVDD.n511 4.5005
R13449 DVDD.n18037 DVDD.n509 4.5005
R13450 DVDD.n18037 DVDD.n510 4.5005
R13451 DVDD.n520 DVDD.n506 4.5005
R13452 DVDD.n520 DVDD.n513 4.5005
R13453 DVDD.n520 DVDD.n507 4.5005
R13454 DVDD.n520 DVDD.n512 4.5005
R13455 DVDD.n520 DVDD.n508 4.5005
R13456 DVDD.n520 DVDD.n511 4.5005
R13457 DVDD.n520 DVDD.n509 4.5005
R13458 DVDD.n520 DVDD.n510 4.5005
R13459 DVDD.n540 DVDD.n512 4.5005
R13460 DVDD.n540 DVDD.n508 4.5005
R13461 DVDD.n540 DVDD.n511 4.5005
R13462 DVDD.n540 DVDD.n509 4.5005
R13463 DVDD.n540 DVDD.n510 4.5005
R13464 DVDD.n522 DVDD.n506 4.5005
R13465 DVDD.n522 DVDD.n513 4.5005
R13466 DVDD.n522 DVDD.n507 4.5005
R13467 DVDD.n522 DVDD.n512 4.5005
R13468 DVDD.n522 DVDD.n508 4.5005
R13469 DVDD.n522 DVDD.n511 4.5005
R13470 DVDD.n522 DVDD.n509 4.5005
R13471 DVDD.n522 DVDD.n510 4.5005
R13472 DVDD.n538 DVDD.n506 4.5005
R13473 DVDD.n538 DVDD.n513 4.5005
R13474 DVDD.n538 DVDD.n507 4.5005
R13475 DVDD.n538 DVDD.n512 4.5005
R13476 DVDD.n538 DVDD.n508 4.5005
R13477 DVDD.n538 DVDD.n511 4.5005
R13478 DVDD.n538 DVDD.n509 4.5005
R13479 DVDD.n538 DVDD.n510 4.5005
R13480 DVDD.n523 DVDD.n506 4.5005
R13481 DVDD.n523 DVDD.n513 4.5005
R13482 DVDD.n523 DVDD.n507 4.5005
R13483 DVDD.n523 DVDD.n512 4.5005
R13484 DVDD.n523 DVDD.n508 4.5005
R13485 DVDD.n523 DVDD.n511 4.5005
R13486 DVDD.n523 DVDD.n509 4.5005
R13487 DVDD.n523 DVDD.n510 4.5005
R13488 DVDD.n537 DVDD.n506 4.5005
R13489 DVDD.n537 DVDD.n513 4.5005
R13490 DVDD.n537 DVDD.n507 4.5005
R13491 DVDD.n537 DVDD.n512 4.5005
R13492 DVDD.n537 DVDD.n508 4.5005
R13493 DVDD.n537 DVDD.n511 4.5005
R13494 DVDD.n537 DVDD.n509 4.5005
R13495 DVDD.n537 DVDD.n510 4.5005
R13496 DVDD.n535 DVDD.n506 4.5005
R13497 DVDD.n535 DVDD.n513 4.5005
R13498 DVDD.n535 DVDD.n507 4.5005
R13499 DVDD.n535 DVDD.n512 4.5005
R13500 DVDD.n535 DVDD.n508 4.5005
R13501 DVDD.n535 DVDD.n511 4.5005
R13502 DVDD.n535 DVDD.n509 4.5005
R13503 DVDD.n535 DVDD.n510 4.5005
R13504 DVDD.n526 DVDD.n506 4.5005
R13505 DVDD.n526 DVDD.n513 4.5005
R13506 DVDD.n526 DVDD.n507 4.5005
R13507 DVDD.n526 DVDD.n512 4.5005
R13508 DVDD.n526 DVDD.n508 4.5005
R13509 DVDD.n526 DVDD.n511 4.5005
R13510 DVDD.n526 DVDD.n509 4.5005
R13511 DVDD.n526 DVDD.n510 4.5005
R13512 DVDD.n534 DVDD.n506 4.5005
R13513 DVDD.n534 DVDD.n513 4.5005
R13514 DVDD.n534 DVDD.n507 4.5005
R13515 DVDD.n534 DVDD.n512 4.5005
R13516 DVDD.n534 DVDD.n508 4.5005
R13517 DVDD.n534 DVDD.n511 4.5005
R13518 DVDD.n534 DVDD.n509 4.5005
R13519 DVDD.n534 DVDD.n510 4.5005
R13520 DVDD.n529 DVDD.n506 4.5005
R13521 DVDD.n529 DVDD.n513 4.5005
R13522 DVDD.n529 DVDD.n507 4.5005
R13523 DVDD.n529 DVDD.n512 4.5005
R13524 DVDD.n529 DVDD.n508 4.5005
R13525 DVDD.n529 DVDD.n511 4.5005
R13526 DVDD.n529 DVDD.n509 4.5005
R13527 DVDD.n529 DVDD.n510 4.5005
R13528 DVDD.n557 DVDD.n552 4.5005
R13529 DVDD.n566 DVDD.n552 4.5005
R13530 DVDD.n556 DVDD.n552 4.5005
R13531 DVDD.n567 DVDD.n552 4.5005
R13532 DVDD.n555 DVDD.n552 4.5005
R13533 DVDD.n568 DVDD.n552 4.5005
R13534 DVDD.n554 DVDD.n552 4.5005
R13535 DVDD.n17978 DVDD.n552 4.5005
R13536 DVDD.n17979 DVDD.n557 4.5005
R13537 DVDD.n17979 DVDD.n566 4.5005
R13538 DVDD.n17979 DVDD.n556 4.5005
R13539 DVDD.n17979 DVDD.n567 4.5005
R13540 DVDD.n17979 DVDD.n555 4.5005
R13541 DVDD.n17979 DVDD.n568 4.5005
R13542 DVDD.n17979 DVDD.n554 4.5005
R13543 DVDD.n17979 DVDD.n17978 4.5005
R13544 DVDD.n590 DVDD.n557 4.5005
R13545 DVDD.n590 DVDD.n566 4.5005
R13546 DVDD.n590 DVDD.n556 4.5005
R13547 DVDD.n590 DVDD.n567 4.5005
R13548 DVDD.n590 DVDD.n555 4.5005
R13549 DVDD.n590 DVDD.n568 4.5005
R13550 DVDD.n590 DVDD.n554 4.5005
R13551 DVDD.n17978 DVDD.n590 4.5005
R13552 DVDD.n573 DVDD.n557 4.5005
R13553 DVDD.n573 DVDD.n566 4.5005
R13554 DVDD.n573 DVDD.n556 4.5005
R13555 DVDD.n573 DVDD.n567 4.5005
R13556 DVDD.n573 DVDD.n555 4.5005
R13557 DVDD.n573 DVDD.n568 4.5005
R13558 DVDD.n573 DVDD.n554 4.5005
R13559 DVDD.n17978 DVDD.n573 4.5005
R13560 DVDD.n591 DVDD.n557 4.5005
R13561 DVDD.n591 DVDD.n566 4.5005
R13562 DVDD.n591 DVDD.n556 4.5005
R13563 DVDD.n591 DVDD.n567 4.5005
R13564 DVDD.n591 DVDD.n555 4.5005
R13565 DVDD.n591 DVDD.n568 4.5005
R13566 DVDD.n591 DVDD.n554 4.5005
R13567 DVDD.n17978 DVDD.n591 4.5005
R13568 DVDD.n572 DVDD.n557 4.5005
R13569 DVDD.n572 DVDD.n566 4.5005
R13570 DVDD.n572 DVDD.n556 4.5005
R13571 DVDD.n572 DVDD.n567 4.5005
R13572 DVDD.n572 DVDD.n555 4.5005
R13573 DVDD.n572 DVDD.n568 4.5005
R13574 DVDD.n572 DVDD.n554 4.5005
R13575 DVDD.n17978 DVDD.n572 4.5005
R13576 DVDD.n592 DVDD.n557 4.5005
R13577 DVDD.n592 DVDD.n566 4.5005
R13578 DVDD.n592 DVDD.n556 4.5005
R13579 DVDD.n592 DVDD.n567 4.5005
R13580 DVDD.n592 DVDD.n555 4.5005
R13581 DVDD.n592 DVDD.n568 4.5005
R13582 DVDD.n592 DVDD.n554 4.5005
R13583 DVDD.n17978 DVDD.n592 4.5005
R13584 DVDD.n571 DVDD.n557 4.5005
R13585 DVDD.n571 DVDD.n566 4.5005
R13586 DVDD.n571 DVDD.n556 4.5005
R13587 DVDD.n571 DVDD.n567 4.5005
R13588 DVDD.n571 DVDD.n555 4.5005
R13589 DVDD.n571 DVDD.n568 4.5005
R13590 DVDD.n571 DVDD.n554 4.5005
R13591 DVDD.n17978 DVDD.n571 4.5005
R13592 DVDD.n593 DVDD.n557 4.5005
R13593 DVDD.n593 DVDD.n566 4.5005
R13594 DVDD.n593 DVDD.n556 4.5005
R13595 DVDD.n593 DVDD.n567 4.5005
R13596 DVDD.n593 DVDD.n555 4.5005
R13597 DVDD.n593 DVDD.n568 4.5005
R13598 DVDD.n593 DVDD.n554 4.5005
R13599 DVDD.n17978 DVDD.n593 4.5005
R13600 DVDD.n570 DVDD.n557 4.5005
R13601 DVDD.n570 DVDD.n566 4.5005
R13602 DVDD.n570 DVDD.n556 4.5005
R13603 DVDD.n570 DVDD.n567 4.5005
R13604 DVDD.n570 DVDD.n555 4.5005
R13605 DVDD.n570 DVDD.n568 4.5005
R13606 DVDD.n570 DVDD.n554 4.5005
R13607 DVDD.n17978 DVDD.n570 4.5005
R13608 DVDD.n17977 DVDD.n557 4.5005
R13609 DVDD.n17977 DVDD.n566 4.5005
R13610 DVDD.n17977 DVDD.n556 4.5005
R13611 DVDD.n17977 DVDD.n567 4.5005
R13612 DVDD.n17977 DVDD.n555 4.5005
R13613 DVDD.n17977 DVDD.n568 4.5005
R13614 DVDD.n17977 DVDD.n554 4.5005
R13615 DVDD.n17978 DVDD.n17977 4.5005
R13616 DVDD.n17964 DVDD.n644 4.5005
R13617 DVDD.n17964 DVDD.n653 4.5005
R13618 DVDD.n17964 DVDD.n643 4.5005
R13619 DVDD.n17964 DVDD.n654 4.5005
R13620 DVDD.n17964 DVDD.n642 4.5005
R13621 DVDD.n17964 DVDD.n655 4.5005
R13622 DVDD.n17964 DVDD.n641 4.5005
R13623 DVDD.n17964 DVDD.n17963 4.5005
R13624 DVDD.n662 DVDD.n644 4.5005
R13625 DVDD.n662 DVDD.n653 4.5005
R13626 DVDD.n662 DVDD.n643 4.5005
R13627 DVDD.n662 DVDD.n654 4.5005
R13628 DVDD.n662 DVDD.n642 4.5005
R13629 DVDD.n662 DVDD.n655 4.5005
R13630 DVDD.n662 DVDD.n641 4.5005
R13631 DVDD.n17963 DVDD.n662 4.5005
R13632 DVDD.n676 DVDD.n644 4.5005
R13633 DVDD.n676 DVDD.n653 4.5005
R13634 DVDD.n676 DVDD.n643 4.5005
R13635 DVDD.n676 DVDD.n654 4.5005
R13636 DVDD.n676 DVDD.n642 4.5005
R13637 DVDD.n676 DVDD.n655 4.5005
R13638 DVDD.n676 DVDD.n641 4.5005
R13639 DVDD.n17963 DVDD.n676 4.5005
R13640 DVDD.n661 DVDD.n644 4.5005
R13641 DVDD.n661 DVDD.n653 4.5005
R13642 DVDD.n661 DVDD.n643 4.5005
R13643 DVDD.n661 DVDD.n654 4.5005
R13644 DVDD.n661 DVDD.n642 4.5005
R13645 DVDD.n661 DVDD.n655 4.5005
R13646 DVDD.n661 DVDD.n641 4.5005
R13647 DVDD.n17963 DVDD.n661 4.5005
R13648 DVDD.n677 DVDD.n644 4.5005
R13649 DVDD.n677 DVDD.n653 4.5005
R13650 DVDD.n677 DVDD.n643 4.5005
R13651 DVDD.n677 DVDD.n654 4.5005
R13652 DVDD.n677 DVDD.n642 4.5005
R13653 DVDD.n677 DVDD.n655 4.5005
R13654 DVDD.n677 DVDD.n641 4.5005
R13655 DVDD.n17963 DVDD.n677 4.5005
R13656 DVDD.n660 DVDD.n644 4.5005
R13657 DVDD.n660 DVDD.n653 4.5005
R13658 DVDD.n660 DVDD.n643 4.5005
R13659 DVDD.n660 DVDD.n654 4.5005
R13660 DVDD.n660 DVDD.n642 4.5005
R13661 DVDD.n660 DVDD.n655 4.5005
R13662 DVDD.n660 DVDD.n641 4.5005
R13663 DVDD.n17963 DVDD.n660 4.5005
R13664 DVDD.n678 DVDD.n644 4.5005
R13665 DVDD.n678 DVDD.n653 4.5005
R13666 DVDD.n678 DVDD.n643 4.5005
R13667 DVDD.n678 DVDD.n654 4.5005
R13668 DVDD.n678 DVDD.n642 4.5005
R13669 DVDD.n678 DVDD.n655 4.5005
R13670 DVDD.n678 DVDD.n641 4.5005
R13671 DVDD.n17963 DVDD.n678 4.5005
R13672 DVDD.n659 DVDD.n644 4.5005
R13673 DVDD.n659 DVDD.n653 4.5005
R13674 DVDD.n659 DVDD.n643 4.5005
R13675 DVDD.n659 DVDD.n654 4.5005
R13676 DVDD.n659 DVDD.n642 4.5005
R13677 DVDD.n659 DVDD.n655 4.5005
R13678 DVDD.n659 DVDD.n641 4.5005
R13679 DVDD.n17963 DVDD.n659 4.5005
R13680 DVDD.n679 DVDD.n644 4.5005
R13681 DVDD.n679 DVDD.n653 4.5005
R13682 DVDD.n679 DVDD.n643 4.5005
R13683 DVDD.n679 DVDD.n654 4.5005
R13684 DVDD.n679 DVDD.n642 4.5005
R13685 DVDD.n679 DVDD.n655 4.5005
R13686 DVDD.n679 DVDD.n641 4.5005
R13687 DVDD.n17963 DVDD.n679 4.5005
R13688 DVDD.n658 DVDD.n644 4.5005
R13689 DVDD.n658 DVDD.n653 4.5005
R13690 DVDD.n658 DVDD.n643 4.5005
R13691 DVDD.n658 DVDD.n654 4.5005
R13692 DVDD.n658 DVDD.n642 4.5005
R13693 DVDD.n658 DVDD.n655 4.5005
R13694 DVDD.n658 DVDD.n641 4.5005
R13695 DVDD.n17963 DVDD.n658 4.5005
R13696 DVDD.n680 DVDD.n644 4.5005
R13697 DVDD.n680 DVDD.n653 4.5005
R13698 DVDD.n680 DVDD.n643 4.5005
R13699 DVDD.n680 DVDD.n654 4.5005
R13700 DVDD.n680 DVDD.n642 4.5005
R13701 DVDD.n680 DVDD.n655 4.5005
R13702 DVDD.n680 DVDD.n641 4.5005
R13703 DVDD.n17963 DVDD.n680 4.5005
R13704 DVDD.n657 DVDD.n644 4.5005
R13705 DVDD.n657 DVDD.n653 4.5005
R13706 DVDD.n657 DVDD.n643 4.5005
R13707 DVDD.n657 DVDD.n654 4.5005
R13708 DVDD.n657 DVDD.n642 4.5005
R13709 DVDD.n657 DVDD.n655 4.5005
R13710 DVDD.n657 DVDD.n641 4.5005
R13711 DVDD.n17963 DVDD.n657 4.5005
R13712 DVDD.n17962 DVDD.n644 4.5005
R13713 DVDD.n17962 DVDD.n653 4.5005
R13714 DVDD.n17962 DVDD.n643 4.5005
R13715 DVDD.n17962 DVDD.n654 4.5005
R13716 DVDD.n17962 DVDD.n642 4.5005
R13717 DVDD.n17962 DVDD.n655 4.5005
R13718 DVDD.n17962 DVDD.n641 4.5005
R13719 DVDD.n17963 DVDD.n17962 4.5005
R13720 DVDD.n748 DVDD.n734 4.5005
R13721 DVDD.n748 DVDD.n742 4.5005
R13722 DVDD.n748 DVDD.n735 4.5005
R13723 DVDD.n748 DVDD.n741 4.5005
R13724 DVDD.n748 DVDD.n736 4.5005
R13725 DVDD.n748 DVDD.n740 4.5005
R13726 DVDD.n748 DVDD.n737 4.5005
R13727 DVDD.n748 DVDD.n739 4.5005
R13728 DVDD.n771 DVDD.n734 4.5005
R13729 DVDD.n771 DVDD.n742 4.5005
R13730 DVDD.n771 DVDD.n735 4.5005
R13731 DVDD.n771 DVDD.n741 4.5005
R13732 DVDD.n771 DVDD.n736 4.5005
R13733 DVDD.n771 DVDD.n740 4.5005
R13734 DVDD.n771 DVDD.n737 4.5005
R13735 DVDD.n771 DVDD.n739 4.5005
R13736 DVDD.n749 DVDD.n734 4.5005
R13737 DVDD.n749 DVDD.n742 4.5005
R13738 DVDD.n749 DVDD.n735 4.5005
R13739 DVDD.n749 DVDD.n741 4.5005
R13740 DVDD.n749 DVDD.n736 4.5005
R13741 DVDD.n749 DVDD.n740 4.5005
R13742 DVDD.n749 DVDD.n737 4.5005
R13743 DVDD.n749 DVDD.n739 4.5005
R13744 DVDD.n770 DVDD.n734 4.5005
R13745 DVDD.n770 DVDD.n742 4.5005
R13746 DVDD.n770 DVDD.n735 4.5005
R13747 DVDD.n770 DVDD.n741 4.5005
R13748 DVDD.n770 DVDD.n736 4.5005
R13749 DVDD.n770 DVDD.n740 4.5005
R13750 DVDD.n770 DVDD.n737 4.5005
R13751 DVDD.n770 DVDD.n739 4.5005
R13752 DVDD.n768 DVDD.n734 4.5005
R13753 DVDD.n768 DVDD.n742 4.5005
R13754 DVDD.n768 DVDD.n735 4.5005
R13755 DVDD.n768 DVDD.n741 4.5005
R13756 DVDD.n768 DVDD.n736 4.5005
R13757 DVDD.n768 DVDD.n740 4.5005
R13758 DVDD.n768 DVDD.n737 4.5005
R13759 DVDD.n768 DVDD.n739 4.5005
R13760 DVDD.n752 DVDD.n734 4.5005
R13761 DVDD.n752 DVDD.n742 4.5005
R13762 DVDD.n752 DVDD.n735 4.5005
R13763 DVDD.n752 DVDD.n741 4.5005
R13764 DVDD.n752 DVDD.n736 4.5005
R13765 DVDD.n752 DVDD.n740 4.5005
R13766 DVDD.n752 DVDD.n737 4.5005
R13767 DVDD.n752 DVDD.n739 4.5005
R13768 DVDD.n767 DVDD.n734 4.5005
R13769 DVDD.n767 DVDD.n742 4.5005
R13770 DVDD.n767 DVDD.n735 4.5005
R13771 DVDD.n767 DVDD.n741 4.5005
R13772 DVDD.n767 DVDD.n736 4.5005
R13773 DVDD.n767 DVDD.n740 4.5005
R13774 DVDD.n767 DVDD.n737 4.5005
R13775 DVDD.n767 DVDD.n739 4.5005
R13776 DVDD.n755 DVDD.n734 4.5005
R13777 DVDD.n755 DVDD.n742 4.5005
R13778 DVDD.n755 DVDD.n735 4.5005
R13779 DVDD.n755 DVDD.n741 4.5005
R13780 DVDD.n755 DVDD.n736 4.5005
R13781 DVDD.n755 DVDD.n740 4.5005
R13782 DVDD.n755 DVDD.n737 4.5005
R13783 DVDD.n755 DVDD.n739 4.5005
R13784 DVDD.n764 DVDD.n734 4.5005
R13785 DVDD.n764 DVDD.n742 4.5005
R13786 DVDD.n764 DVDD.n735 4.5005
R13787 DVDD.n764 DVDD.n741 4.5005
R13788 DVDD.n764 DVDD.n736 4.5005
R13789 DVDD.n764 DVDD.n740 4.5005
R13790 DVDD.n764 DVDD.n737 4.5005
R13791 DVDD.n764 DVDD.n739 4.5005
R13792 DVDD.n756 DVDD.n734 4.5005
R13793 DVDD.n756 DVDD.n742 4.5005
R13794 DVDD.n756 DVDD.n735 4.5005
R13795 DVDD.n756 DVDD.n741 4.5005
R13796 DVDD.n756 DVDD.n736 4.5005
R13797 DVDD.n756 DVDD.n740 4.5005
R13798 DVDD.n756 DVDD.n737 4.5005
R13799 DVDD.n756 DVDD.n739 4.5005
R13800 DVDD.n17878 DVDD.n788 4.5005
R13801 DVDD.n17878 DVDD.n797 4.5005
R13802 DVDD.n17878 DVDD.n787 4.5005
R13803 DVDD.n17878 DVDD.n798 4.5005
R13804 DVDD.n17878 DVDD.n786 4.5005
R13805 DVDD.n17878 DVDD.n799 4.5005
R13806 DVDD.n17878 DVDD.n785 4.5005
R13807 DVDD.n17878 DVDD.n17877 4.5005
R13808 DVDD.n811 DVDD.n788 4.5005
R13809 DVDD.n811 DVDD.n797 4.5005
R13810 DVDD.n811 DVDD.n787 4.5005
R13811 DVDD.n811 DVDD.n798 4.5005
R13812 DVDD.n811 DVDD.n786 4.5005
R13813 DVDD.n811 DVDD.n799 4.5005
R13814 DVDD.n811 DVDD.n785 4.5005
R13815 DVDD.n17877 DVDD.n811 4.5005
R13816 DVDD.n802 DVDD.n788 4.5005
R13817 DVDD.n802 DVDD.n797 4.5005
R13818 DVDD.n802 DVDD.n787 4.5005
R13819 DVDD.n802 DVDD.n798 4.5005
R13820 DVDD.n802 DVDD.n786 4.5005
R13821 DVDD.n802 DVDD.n799 4.5005
R13822 DVDD.n802 DVDD.n785 4.5005
R13823 DVDD.n17877 DVDD.n802 4.5005
R13824 DVDD.n812 DVDD.n788 4.5005
R13825 DVDD.n812 DVDD.n797 4.5005
R13826 DVDD.n812 DVDD.n787 4.5005
R13827 DVDD.n812 DVDD.n798 4.5005
R13828 DVDD.n812 DVDD.n786 4.5005
R13829 DVDD.n812 DVDD.n799 4.5005
R13830 DVDD.n812 DVDD.n785 4.5005
R13831 DVDD.n17877 DVDD.n812 4.5005
R13832 DVDD.n801 DVDD.n788 4.5005
R13833 DVDD.n801 DVDD.n797 4.5005
R13834 DVDD.n801 DVDD.n787 4.5005
R13835 DVDD.n801 DVDD.n798 4.5005
R13836 DVDD.n801 DVDD.n786 4.5005
R13837 DVDD.n801 DVDD.n799 4.5005
R13838 DVDD.n801 DVDD.n785 4.5005
R13839 DVDD.n17877 DVDD.n801 4.5005
R13840 DVDD.n17876 DVDD.n788 4.5005
R13841 DVDD.n17876 DVDD.n797 4.5005
R13842 DVDD.n17876 DVDD.n787 4.5005
R13843 DVDD.n17876 DVDD.n798 4.5005
R13844 DVDD.n17876 DVDD.n786 4.5005
R13845 DVDD.n17876 DVDD.n799 4.5005
R13846 DVDD.n17876 DVDD.n785 4.5005
R13847 DVDD.n17877 DVDD.n17876 4.5005
R13848 DVDD.n15131 DVDD.n5643 4.5005
R13849 DVDD.n5986 DVDD.n5643 4.5005
R13850 DVDD.n5643 DVDD.n5593 4.5005
R13851 DVDD.n5740 DVDD.n5643 4.5005
R13852 DVDD.n17710 DVDD.n17371 4.5005
R13853 DVDD.n17371 DVDD.n17306 4.5005
R13854 DVDD.n17371 DVDD.n17309 4.5005
R13855 DVDD.n17371 DVDD.n17307 4.5005
R13856 DVDD.n15131 DVDD.n5641 4.5005
R13857 DVDD.n5641 DVDD.n5593 4.5005
R13858 DVDD.n5641 DVDD.n5592 4.5005
R13859 DVDD.n17710 DVDD.n17360 4.5005
R13860 DVDD.n17360 DVDD.n17306 4.5005
R13861 DVDD.n17360 DVDD.n17309 4.5005
R13862 DVDD.n17710 DVDD.n17374 4.5005
R13863 DVDD.n17374 DVDD.n17309 4.5005
R13864 DVDD.n17374 DVDD.n17308 4.5005
R13865 DVDD.n17710 DVDD.n17359 4.5005
R13866 DVDD.n17359 DVDD.n17309 4.5005
R13867 DVDD.n17359 DVDD.n17308 4.5005
R13868 DVDD.n17710 DVDD.n17377 4.5005
R13869 DVDD.n17377 DVDD.n17309 4.5005
R13870 DVDD.n17377 DVDD.n17308 4.5005
R13871 DVDD.n17710 DVDD.n17358 4.5005
R13872 DVDD.n17358 DVDD.n17309 4.5005
R13873 DVDD.n17358 DVDD.n17308 4.5005
R13874 DVDD.n17710 DVDD.n17380 4.5005
R13875 DVDD.n17380 DVDD.n17309 4.5005
R13876 DVDD.n17380 DVDD.n17308 4.5005
R13877 DVDD.n17710 DVDD.n17357 4.5005
R13878 DVDD.n17357 DVDD.n17309 4.5005
R13879 DVDD.n17357 DVDD.n17308 4.5005
R13880 DVDD.n17710 DVDD.n17383 4.5005
R13881 DVDD.n17383 DVDD.n17309 4.5005
R13882 DVDD.n17383 DVDD.n17308 4.5005
R13883 DVDD.n17710 DVDD.n17356 4.5005
R13884 DVDD.n17356 DVDD.n17309 4.5005
R13885 DVDD.n17356 DVDD.n17308 4.5005
R13886 DVDD.n17710 DVDD.n17386 4.5005
R13887 DVDD.n17386 DVDD.n17309 4.5005
R13888 DVDD.n17386 DVDD.n17308 4.5005
R13889 DVDD.n17710 DVDD.n17355 4.5005
R13890 DVDD.n17355 DVDD.n17309 4.5005
R13891 DVDD.n17355 DVDD.n17308 4.5005
R13892 DVDD.n17710 DVDD.n17389 4.5005
R13893 DVDD.n17389 DVDD.n17309 4.5005
R13894 DVDD.n17389 DVDD.n17308 4.5005
R13895 DVDD.n17710 DVDD.n17354 4.5005
R13896 DVDD.n17354 DVDD.n17309 4.5005
R13897 DVDD.n17354 DVDD.n17308 4.5005
R13898 DVDD.n17710 DVDD.n17392 4.5005
R13899 DVDD.n17392 DVDD.n17309 4.5005
R13900 DVDD.n17392 DVDD.n17308 4.5005
R13901 DVDD.n17710 DVDD.n17353 4.5005
R13902 DVDD.n17353 DVDD.n17309 4.5005
R13903 DVDD.n17353 DVDD.n17308 4.5005
R13904 DVDD.n17710 DVDD.n17395 4.5005
R13905 DVDD.n17395 DVDD.n17309 4.5005
R13906 DVDD.n17395 DVDD.n17308 4.5005
R13907 DVDD.n17710 DVDD.n17352 4.5005
R13908 DVDD.n17352 DVDD.n17309 4.5005
R13909 DVDD.n17352 DVDD.n17308 4.5005
R13910 DVDD.n17710 DVDD.n17398 4.5005
R13911 DVDD.n17398 DVDD.n17309 4.5005
R13912 DVDD.n17398 DVDD.n17308 4.5005
R13913 DVDD.n17710 DVDD.n17351 4.5005
R13914 DVDD.n17351 DVDD.n17309 4.5005
R13915 DVDD.n17351 DVDD.n17308 4.5005
R13916 DVDD.n17710 DVDD.n17401 4.5005
R13917 DVDD.n17401 DVDD.n17309 4.5005
R13918 DVDD.n17401 DVDD.n17308 4.5005
R13919 DVDD.n17710 DVDD.n17350 4.5005
R13920 DVDD.n17350 DVDD.n17309 4.5005
R13921 DVDD.n17350 DVDD.n17308 4.5005
R13922 DVDD.n17710 DVDD.n17404 4.5005
R13923 DVDD.n17404 DVDD.n17309 4.5005
R13924 DVDD.n17404 DVDD.n17308 4.5005
R13925 DVDD.n17710 DVDD.n17349 4.5005
R13926 DVDD.n17349 DVDD.n17309 4.5005
R13927 DVDD.n17349 DVDD.n17308 4.5005
R13928 DVDD.n17710 DVDD.n17407 4.5005
R13929 DVDD.n17407 DVDD.n17309 4.5005
R13930 DVDD.n17407 DVDD.n17308 4.5005
R13931 DVDD.n17710 DVDD.n17348 4.5005
R13932 DVDD.n17348 DVDD.n17309 4.5005
R13933 DVDD.n17348 DVDD.n17308 4.5005
R13934 DVDD.n17710 DVDD.n17410 4.5005
R13935 DVDD.n17410 DVDD.n17309 4.5005
R13936 DVDD.n17410 DVDD.n17308 4.5005
R13937 DVDD.n17710 DVDD.n17347 4.5005
R13938 DVDD.n17347 DVDD.n17309 4.5005
R13939 DVDD.n17347 DVDD.n17308 4.5005
R13940 DVDD.n17710 DVDD.n17413 4.5005
R13941 DVDD.n17413 DVDD.n17309 4.5005
R13942 DVDD.n17413 DVDD.n17308 4.5005
R13943 DVDD.n17710 DVDD.n17346 4.5005
R13944 DVDD.n17346 DVDD.n17309 4.5005
R13945 DVDD.n17346 DVDD.n17308 4.5005
R13946 DVDD.n17710 DVDD.n17416 4.5005
R13947 DVDD.n17416 DVDD.n17309 4.5005
R13948 DVDD.n17416 DVDD.n17308 4.5005
R13949 DVDD.n17710 DVDD.n17345 4.5005
R13950 DVDD.n17345 DVDD.n17309 4.5005
R13951 DVDD.n17345 DVDD.n17308 4.5005
R13952 DVDD.n17710 DVDD.n17419 4.5005
R13953 DVDD.n17419 DVDD.n17309 4.5005
R13954 DVDD.n17419 DVDD.n17308 4.5005
R13955 DVDD.n17710 DVDD.n17344 4.5005
R13956 DVDD.n17344 DVDD.n17309 4.5005
R13957 DVDD.n17344 DVDD.n17308 4.5005
R13958 DVDD.n17710 DVDD.n17422 4.5005
R13959 DVDD.n17422 DVDD.n17309 4.5005
R13960 DVDD.n17422 DVDD.n17308 4.5005
R13961 DVDD.n17710 DVDD.n17343 4.5005
R13962 DVDD.n17343 DVDD.n17309 4.5005
R13963 DVDD.n17343 DVDD.n17308 4.5005
R13964 DVDD.n17710 DVDD.n17425 4.5005
R13965 DVDD.n17425 DVDD.n17309 4.5005
R13966 DVDD.n17425 DVDD.n17308 4.5005
R13967 DVDD.n17710 DVDD.n17342 4.5005
R13968 DVDD.n17342 DVDD.n17309 4.5005
R13969 DVDD.n17342 DVDD.n17308 4.5005
R13970 DVDD.n17710 DVDD.n17428 4.5005
R13971 DVDD.n17428 DVDD.n17309 4.5005
R13972 DVDD.n17428 DVDD.n17308 4.5005
R13973 DVDD.n17710 DVDD.n17341 4.5005
R13974 DVDD.n17341 DVDD.n17309 4.5005
R13975 DVDD.n17341 DVDD.n17308 4.5005
R13976 DVDD.n17710 DVDD.n17431 4.5005
R13977 DVDD.n17431 DVDD.n17309 4.5005
R13978 DVDD.n17431 DVDD.n17308 4.5005
R13979 DVDD.n17710 DVDD.n17340 4.5005
R13980 DVDD.n17340 DVDD.n17309 4.5005
R13981 DVDD.n17340 DVDD.n17308 4.5005
R13982 DVDD.n17710 DVDD.n17434 4.5005
R13983 DVDD.n17434 DVDD.n17309 4.5005
R13984 DVDD.n17434 DVDD.n17308 4.5005
R13985 DVDD.n17710 DVDD.n17339 4.5005
R13986 DVDD.n17339 DVDD.n17309 4.5005
R13987 DVDD.n17339 DVDD.n17308 4.5005
R13988 DVDD.n17710 DVDD.n17437 4.5005
R13989 DVDD.n17437 DVDD.n17309 4.5005
R13990 DVDD.n17437 DVDD.n17308 4.5005
R13991 DVDD.n17710 DVDD.n17338 4.5005
R13992 DVDD.n17338 DVDD.n17309 4.5005
R13993 DVDD.n17338 DVDD.n17308 4.5005
R13994 DVDD.n17710 DVDD.n17440 4.5005
R13995 DVDD.n17440 DVDD.n17309 4.5005
R13996 DVDD.n17440 DVDD.n17308 4.5005
R13997 DVDD.n17710 DVDD.n17337 4.5005
R13998 DVDD.n17337 DVDD.n17309 4.5005
R13999 DVDD.n17337 DVDD.n17308 4.5005
R14000 DVDD.n17710 DVDD.n17443 4.5005
R14001 DVDD.n17443 DVDD.n17309 4.5005
R14002 DVDD.n17443 DVDD.n17308 4.5005
R14003 DVDD.n17710 DVDD.n17336 4.5005
R14004 DVDD.n17336 DVDD.n17309 4.5005
R14005 DVDD.n17336 DVDD.n17308 4.5005
R14006 DVDD.n17710 DVDD.n17446 4.5005
R14007 DVDD.n17446 DVDD.n17309 4.5005
R14008 DVDD.n17446 DVDD.n17308 4.5005
R14009 DVDD.n17710 DVDD.n17335 4.5005
R14010 DVDD.n17335 DVDD.n17309 4.5005
R14011 DVDD.n17335 DVDD.n17308 4.5005
R14012 DVDD.n17710 DVDD.n17449 4.5005
R14013 DVDD.n17449 DVDD.n17309 4.5005
R14014 DVDD.n17449 DVDD.n17308 4.5005
R14015 DVDD.n17710 DVDD.n17334 4.5005
R14016 DVDD.n17334 DVDD.n17309 4.5005
R14017 DVDD.n17334 DVDD.n17308 4.5005
R14018 DVDD.n17710 DVDD.n17452 4.5005
R14019 DVDD.n17452 DVDD.n17309 4.5005
R14020 DVDD.n17452 DVDD.n17308 4.5005
R14021 DVDD.n17710 DVDD.n17333 4.5005
R14022 DVDD.n17333 DVDD.n17309 4.5005
R14023 DVDD.n17333 DVDD.n17308 4.5005
R14024 DVDD.n17710 DVDD.n17455 4.5005
R14025 DVDD.n17455 DVDD.n17309 4.5005
R14026 DVDD.n17455 DVDD.n17308 4.5005
R14027 DVDD.n17710 DVDD.n17332 4.5005
R14028 DVDD.n17332 DVDD.n17309 4.5005
R14029 DVDD.n17332 DVDD.n17308 4.5005
R14030 DVDD.n17710 DVDD.n17458 4.5005
R14031 DVDD.n17458 DVDD.n17309 4.5005
R14032 DVDD.n17458 DVDD.n17308 4.5005
R14033 DVDD.n17710 DVDD.n17331 4.5005
R14034 DVDD.n17331 DVDD.n17309 4.5005
R14035 DVDD.n17331 DVDD.n17308 4.5005
R14036 DVDD.n17710 DVDD.n17461 4.5005
R14037 DVDD.n17461 DVDD.n17309 4.5005
R14038 DVDD.n17461 DVDD.n17308 4.5005
R14039 DVDD.n17710 DVDD.n17330 4.5005
R14040 DVDD.n17330 DVDD.n17309 4.5005
R14041 DVDD.n17330 DVDD.n17308 4.5005
R14042 DVDD.n17710 DVDD.n17464 4.5005
R14043 DVDD.n17464 DVDD.n17309 4.5005
R14044 DVDD.n17464 DVDD.n17308 4.5005
R14045 DVDD.n17710 DVDD.n17329 4.5005
R14046 DVDD.n17329 DVDD.n17309 4.5005
R14047 DVDD.n17329 DVDD.n17308 4.5005
R14048 DVDD.n17710 DVDD.n17467 4.5005
R14049 DVDD.n17467 DVDD.n17309 4.5005
R14050 DVDD.n17467 DVDD.n17308 4.5005
R14051 DVDD.n17710 DVDD.n17328 4.5005
R14052 DVDD.n17328 DVDD.n17309 4.5005
R14053 DVDD.n17328 DVDD.n17308 4.5005
R14054 DVDD.n17710 DVDD.n17470 4.5005
R14055 DVDD.n17470 DVDD.n17309 4.5005
R14056 DVDD.n17470 DVDD.n17308 4.5005
R14057 DVDD.n17710 DVDD.n17327 4.5005
R14058 DVDD.n17327 DVDD.n17309 4.5005
R14059 DVDD.n17327 DVDD.n17308 4.5005
R14060 DVDD.n17710 DVDD.n17473 4.5005
R14061 DVDD.n17473 DVDD.n17309 4.5005
R14062 DVDD.n17473 DVDD.n17308 4.5005
R14063 DVDD.n17710 DVDD.n17326 4.5005
R14064 DVDD.n17326 DVDD.n17309 4.5005
R14065 DVDD.n17326 DVDD.n17308 4.5005
R14066 DVDD.n17710 DVDD.n17476 4.5005
R14067 DVDD.n17476 DVDD.n17309 4.5005
R14068 DVDD.n17476 DVDD.n17308 4.5005
R14069 DVDD.n17710 DVDD.n17325 4.5005
R14070 DVDD.n17325 DVDD.n17309 4.5005
R14071 DVDD.n17325 DVDD.n17308 4.5005
R14072 DVDD.n17710 DVDD.n17479 4.5005
R14073 DVDD.n17479 DVDD.n17309 4.5005
R14074 DVDD.n17479 DVDD.n17308 4.5005
R14075 DVDD.n17710 DVDD.n17324 4.5005
R14076 DVDD.n17324 DVDD.n17309 4.5005
R14077 DVDD.n17324 DVDD.n17308 4.5005
R14078 DVDD.n17710 DVDD.n17482 4.5005
R14079 DVDD.n17482 DVDD.n17309 4.5005
R14080 DVDD.n17482 DVDD.n17308 4.5005
R14081 DVDD.n17710 DVDD.n17323 4.5005
R14082 DVDD.n17323 DVDD.n17309 4.5005
R14083 DVDD.n17323 DVDD.n17308 4.5005
R14084 DVDD.n17710 DVDD.n17485 4.5005
R14085 DVDD.n17485 DVDD.n17309 4.5005
R14086 DVDD.n17485 DVDD.n17308 4.5005
R14087 DVDD.n17710 DVDD.n17322 4.5005
R14088 DVDD.n17322 DVDD.n17309 4.5005
R14089 DVDD.n17322 DVDD.n17308 4.5005
R14090 DVDD.n17710 DVDD.n17488 4.5005
R14091 DVDD.n17488 DVDD.n17309 4.5005
R14092 DVDD.n17488 DVDD.n17308 4.5005
R14093 DVDD.n17710 DVDD.n17321 4.5005
R14094 DVDD.n17321 DVDD.n17309 4.5005
R14095 DVDD.n17321 DVDD.n17308 4.5005
R14096 DVDD.n17710 DVDD.n17491 4.5005
R14097 DVDD.n17491 DVDD.n17309 4.5005
R14098 DVDD.n17491 DVDD.n17308 4.5005
R14099 DVDD.n17710 DVDD.n17320 4.5005
R14100 DVDD.n17320 DVDD.n17309 4.5005
R14101 DVDD.n17320 DVDD.n17308 4.5005
R14102 DVDD.n17710 DVDD.n17494 4.5005
R14103 DVDD.n17494 DVDD.n17309 4.5005
R14104 DVDD.n17494 DVDD.n17308 4.5005
R14105 DVDD.n17710 DVDD.n17319 4.5005
R14106 DVDD.n17319 DVDD.n17309 4.5005
R14107 DVDD.n17319 DVDD.n17308 4.5005
R14108 DVDD.n17710 DVDD.n17497 4.5005
R14109 DVDD.n17497 DVDD.n17309 4.5005
R14110 DVDD.n17497 DVDD.n17308 4.5005
R14111 DVDD.n17710 DVDD.n17318 4.5005
R14112 DVDD.n17318 DVDD.n17309 4.5005
R14113 DVDD.n17318 DVDD.n17308 4.5005
R14114 DVDD.n17710 DVDD.n17500 4.5005
R14115 DVDD.n17500 DVDD.n17309 4.5005
R14116 DVDD.n17500 DVDD.n17308 4.5005
R14117 DVDD.n17710 DVDD.n17317 4.5005
R14118 DVDD.n17317 DVDD.n17309 4.5005
R14119 DVDD.n17317 DVDD.n17308 4.5005
R14120 DVDD.n17710 DVDD.n17503 4.5005
R14121 DVDD.n17503 DVDD.n17309 4.5005
R14122 DVDD.n17503 DVDD.n17308 4.5005
R14123 DVDD.n17710 DVDD.n17316 4.5005
R14124 DVDD.n17316 DVDD.n17309 4.5005
R14125 DVDD.n17316 DVDD.n17308 4.5005
R14126 DVDD.n17710 DVDD.n17506 4.5005
R14127 DVDD.n17506 DVDD.n17309 4.5005
R14128 DVDD.n17506 DVDD.n17308 4.5005
R14129 DVDD.n17710 DVDD.n17315 4.5005
R14130 DVDD.n17315 DVDD.n17309 4.5005
R14131 DVDD.n17315 DVDD.n17308 4.5005
R14132 DVDD.n17710 DVDD.n17509 4.5005
R14133 DVDD.n17509 DVDD.n17309 4.5005
R14134 DVDD.n17509 DVDD.n17308 4.5005
R14135 DVDD.n17710 DVDD.n17314 4.5005
R14136 DVDD.n17314 DVDD.n17309 4.5005
R14137 DVDD.n17314 DVDD.n17308 4.5005
R14138 DVDD.n17710 DVDD.n17512 4.5005
R14139 DVDD.n17512 DVDD.n17309 4.5005
R14140 DVDD.n17512 DVDD.n17308 4.5005
R14141 DVDD.n17710 DVDD.n17313 4.5005
R14142 DVDD.n17313 DVDD.n17309 4.5005
R14143 DVDD.n17313 DVDD.n17308 4.5005
R14144 DVDD.n17710 DVDD.n17709 4.5005
R14145 DVDD.n17709 DVDD.n17309 4.5005
R14146 DVDD.n17709 DVDD.n17308 4.5005
R14147 DVDD.n17710 DVDD.n17312 4.5005
R14148 DVDD.n17312 DVDD.n17309 4.5005
R14149 DVDD.n17312 DVDD.n17307 4.5005
R14150 DVDD.n17312 DVDD.n17308 4.5005
R14151 DVDD.n5642 DVDD.n5584 4.5005
R14152 DVDD.n5987 DVDD.n5584 4.5005
R14153 DVDD.n5938 DVDD.n5584 4.5005
R14154 DVDD.n5991 DVDD.n5584 4.5005
R14155 DVDD.n5934 DVDD.n5584 4.5005
R14156 DVDD.n17369 DVDD.n898 4.5005
R14157 DVDD.n17366 DVDD.n898 4.5005
R14158 DVDD.n17367 DVDD.n898 4.5005
R14159 DVDD.n5992 DVDD.n5642 4.5005
R14160 DVDD.n5992 DVDD.n5987 4.5005
R14161 DVDD.n5992 DVDD.n5938 4.5005
R14162 DVDD.n5992 DVDD.n5991 4.5005
R14163 DVDD.n5992 DVDD.n5934 4.5005
R14164 DVDD.n17362 DVDD.n907 4.5005
R14165 DVDD.n17362 DVDD.n17311 4.5005
R14166 DVDD.n17369 DVDD.n17362 4.5005
R14167 DVDD.n17366 DVDD.n17362 4.5005
R14168 DVDD.n17367 DVDD.n17362 4.5005
R14169 DVDD.n5936 DVDD.n5642 4.5005
R14170 DVDD.n5987 DVDD.n5936 4.5005
R14171 DVDD.n5938 DVDD.n5936 4.5005
R14172 DVDD.n5991 DVDD.n5936 4.5005
R14173 DVDD.n5936 DVDD.n5934 4.5005
R14174 DVDD.n17361 DVDD.n907 4.5005
R14175 DVDD.n17361 DVDD.n17311 4.5005
R14176 DVDD.n17369 DVDD.n17361 4.5005
R14177 DVDD.n17366 DVDD.n17361 4.5005
R14178 DVDD.n17367 DVDD.n17361 4.5005
R14179 DVDD.n5990 DVDD.n5642 4.5005
R14180 DVDD.n5990 DVDD.n5987 4.5005
R14181 DVDD.n5990 DVDD.n5938 4.5005
R14182 DVDD.n5991 DVDD.n5990 4.5005
R14183 DVDD.n5990 DVDD.n5934 4.5005
R14184 DVDD.n17368 DVDD.n907 4.5005
R14185 DVDD.n17368 DVDD.n17311 4.5005
R14186 DVDD.n17369 DVDD.n17368 4.5005
R14187 DVDD.n17368 DVDD.n17366 4.5005
R14188 DVDD.n17368 DVDD.n17367 4.5005
R14189 DVDD.n1603 DVDD.n1262 4.5005
R14190 DVDD.n1356 DVDD.n1262 4.5005
R14191 DVDD.n17262 DVDD.n1653 4.5005
R14192 DVDD.n17262 DVDD.n17261 4.5005
R14193 DVDD.n16994 DVDD.n1754 4.5005
R14194 DVDD.n16994 DVDD.n16993 4.5005
R14195 DVDD.n2154 DVDD.n1813 4.5005
R14196 DVDD.n1907 DVDD.n1813 4.5005
R14197 DVDD.n16704 DVDD.n2207 4.5005
R14198 DVDD.n16704 DVDD.n16703 4.5005
R14199 DVDD.n13254 DVDD.n12912 4.5005
R14200 DVDD.n13007 DVDD.n12912 4.5005
R14201 DVDD.n13471 DVDD.n13470 4.5005
R14202 DVDD.n13470 DVDD.n13469 4.5005
R14203 DVDD.n13485 DVDD.n13484 4.5005
R14204 DVDD.n13484 DVDD.n13483 4.5005
R14205 DVDD.n13744 DVDD.n12329 4.5005
R14206 DVDD.n13744 DVDD.n13743 4.5005
R14207 DVDD.n12028 DVDD.n11938 4.5005
R14208 DVDD.n12275 DVDD.n11938 4.5005
R14209 DVDD.n13777 DVDD.n11630 4.5005
R14210 DVDD.n13777 DVDD.n13776 4.5005
R14211 DVDD.n13799 DVDD.n11275 4.5005
R14212 DVDD.n13799 DVDD.n13798 4.5005
R14213 DVDD.n14001 DVDD.n14000 4.5005
R14214 DVDD.n14000 DVDD.n13999 4.5005
R14215 DVDD.n10801 DVDD.n10711 4.5005
R14216 DVDD.n11048 DVDD.n10711 4.5005
R14217 DVDD.n14269 DVDD.n10639 4.5005
R14218 DVDD.n14269 DVDD.n14268 4.5005
R14219 DVDD.n14282 DVDD.n14281 4.5005
R14220 DVDD.n14281 DVDD.n14280 4.5005
R14221 DVDD.n8947 DVDD.n8610 4.5005
R14222 DVDD.n8738 DVDD.n8610 4.5005
R14223 DVDD.n8349 DVDD.n8259 4.5005
R14224 DVDD.n8596 DVDD.n8259 4.5005
R14225 DVDD.n14559 DVDD.n8204 4.5005
R14226 DVDD.n14559 DVDD.n14558 4.5005
R14227 DVDD.n14825 DVDD.n8086 4.5005
R14228 DVDD.n14825 DVDD.n14824 4.5005
R14229 DVDD.n14838 DVDD.n14837 4.5005
R14230 DVDD.n14837 DVDD.n14836 4.5005
R14231 DVDD.n9556 DVDD.n7679 4.5005
R14232 DVDD.n9309 DVDD.n7679 4.5005
R14233 DVDD.n14861 DVDD.n14860 4.5005
R14234 DVDD.n14860 DVDD.n14859 4.5005
R14235 DVDD.n15058 DVDD.n15057 4.5005
R14236 DVDD.n15057 DVDD.n15056 4.5005
R14237 DVDD.n7404 DVDD.n7111 4.5005
R14238 DVDD.n7404 DVDD.n7403 4.5005
R14239 DVDD.n15090 DVDD.n15089 4.5005
R14240 DVDD.n15089 DVDD.n15088 4.5005
R14241 DVDD.n5644 DVDD.n5592 4.5005
R14242 DVDD.n5740 DVDD.n5644 4.5005
R14243 DVDD.n5644 DVDD.n5593 4.5005
R14244 DVDD.n15131 DVDD.n5644 4.5005
R14245 DVDD.n15132 DVDD.n5592 4.5005
R14246 DVDD.n15132 DVDD.n5593 4.5005
R14247 DVDD.n15132 DVDD.n15131 4.5005
R14248 DVDD.n5645 DVDD.n5592 4.5005
R14249 DVDD.n5645 DVDD.n5593 4.5005
R14250 DVDD.n15131 DVDD.n5645 4.5005
R14251 DVDD.n5640 DVDD.n5592 4.5005
R14252 DVDD.n5640 DVDD.n5593 4.5005
R14253 DVDD.n15131 DVDD.n5640 4.5005
R14254 DVDD.n5646 DVDD.n5592 4.5005
R14255 DVDD.n5646 DVDD.n5593 4.5005
R14256 DVDD.n15131 DVDD.n5646 4.5005
R14257 DVDD.n5639 DVDD.n5592 4.5005
R14258 DVDD.n5639 DVDD.n5593 4.5005
R14259 DVDD.n15131 DVDD.n5639 4.5005
R14260 DVDD.n5647 DVDD.n5592 4.5005
R14261 DVDD.n5647 DVDD.n5593 4.5005
R14262 DVDD.n15131 DVDD.n5647 4.5005
R14263 DVDD.n5638 DVDD.n5592 4.5005
R14264 DVDD.n5638 DVDD.n5593 4.5005
R14265 DVDD.n15131 DVDD.n5638 4.5005
R14266 DVDD.n5648 DVDD.n5592 4.5005
R14267 DVDD.n5648 DVDD.n5593 4.5005
R14268 DVDD.n15131 DVDD.n5648 4.5005
R14269 DVDD.n5637 DVDD.n5592 4.5005
R14270 DVDD.n5637 DVDD.n5593 4.5005
R14271 DVDD.n15131 DVDD.n5637 4.5005
R14272 DVDD.n5649 DVDD.n5592 4.5005
R14273 DVDD.n5649 DVDD.n5593 4.5005
R14274 DVDD.n15131 DVDD.n5649 4.5005
R14275 DVDD.n5636 DVDD.n5592 4.5005
R14276 DVDD.n5636 DVDD.n5593 4.5005
R14277 DVDD.n15131 DVDD.n5636 4.5005
R14278 DVDD.n5650 DVDD.n5592 4.5005
R14279 DVDD.n5650 DVDD.n5593 4.5005
R14280 DVDD.n15131 DVDD.n5650 4.5005
R14281 DVDD.n5635 DVDD.n5592 4.5005
R14282 DVDD.n5635 DVDD.n5593 4.5005
R14283 DVDD.n15131 DVDD.n5635 4.5005
R14284 DVDD.n5651 DVDD.n5592 4.5005
R14285 DVDD.n5651 DVDD.n5593 4.5005
R14286 DVDD.n15131 DVDD.n5651 4.5005
R14287 DVDD.n5634 DVDD.n5592 4.5005
R14288 DVDD.n5634 DVDD.n5593 4.5005
R14289 DVDD.n15131 DVDD.n5634 4.5005
R14290 DVDD.n5652 DVDD.n5592 4.5005
R14291 DVDD.n5652 DVDD.n5593 4.5005
R14292 DVDD.n15131 DVDD.n5652 4.5005
R14293 DVDD.n5633 DVDD.n5592 4.5005
R14294 DVDD.n5633 DVDD.n5593 4.5005
R14295 DVDD.n15131 DVDD.n5633 4.5005
R14296 DVDD.n5653 DVDD.n5592 4.5005
R14297 DVDD.n5653 DVDD.n5593 4.5005
R14298 DVDD.n15131 DVDD.n5653 4.5005
R14299 DVDD.n5632 DVDD.n5592 4.5005
R14300 DVDD.n5632 DVDD.n5593 4.5005
R14301 DVDD.n15131 DVDD.n5632 4.5005
R14302 DVDD.n5654 DVDD.n5592 4.5005
R14303 DVDD.n5654 DVDD.n5593 4.5005
R14304 DVDD.n15131 DVDD.n5654 4.5005
R14305 DVDD.n5631 DVDD.n5592 4.5005
R14306 DVDD.n5631 DVDD.n5593 4.5005
R14307 DVDD.n15131 DVDD.n5631 4.5005
R14308 DVDD.n5655 DVDD.n5592 4.5005
R14309 DVDD.n5655 DVDD.n5593 4.5005
R14310 DVDD.n15131 DVDD.n5655 4.5005
R14311 DVDD.n5630 DVDD.n5592 4.5005
R14312 DVDD.n5630 DVDD.n5593 4.5005
R14313 DVDD.n15131 DVDD.n5630 4.5005
R14314 DVDD.n5656 DVDD.n5592 4.5005
R14315 DVDD.n5656 DVDD.n5593 4.5005
R14316 DVDD.n15131 DVDD.n5656 4.5005
R14317 DVDD.n5629 DVDD.n5592 4.5005
R14318 DVDD.n5629 DVDD.n5593 4.5005
R14319 DVDD.n15131 DVDD.n5629 4.5005
R14320 DVDD.n5657 DVDD.n5592 4.5005
R14321 DVDD.n5657 DVDD.n5593 4.5005
R14322 DVDD.n15131 DVDD.n5657 4.5005
R14323 DVDD.n5628 DVDD.n5592 4.5005
R14324 DVDD.n5628 DVDD.n5593 4.5005
R14325 DVDD.n15131 DVDD.n5628 4.5005
R14326 DVDD.n5658 DVDD.n5592 4.5005
R14327 DVDD.n5658 DVDD.n5593 4.5005
R14328 DVDD.n15131 DVDD.n5658 4.5005
R14329 DVDD.n5627 DVDD.n5592 4.5005
R14330 DVDD.n5627 DVDD.n5593 4.5005
R14331 DVDD.n15131 DVDD.n5627 4.5005
R14332 DVDD.n5659 DVDD.n5592 4.5005
R14333 DVDD.n5659 DVDD.n5593 4.5005
R14334 DVDD.n15131 DVDD.n5659 4.5005
R14335 DVDD.n5626 DVDD.n5592 4.5005
R14336 DVDD.n5626 DVDD.n5593 4.5005
R14337 DVDD.n15131 DVDD.n5626 4.5005
R14338 DVDD.n5660 DVDD.n5592 4.5005
R14339 DVDD.n5660 DVDD.n5593 4.5005
R14340 DVDD.n15131 DVDD.n5660 4.5005
R14341 DVDD.n5625 DVDD.n5592 4.5005
R14342 DVDD.n5625 DVDD.n5593 4.5005
R14343 DVDD.n15131 DVDD.n5625 4.5005
R14344 DVDD.n5661 DVDD.n5592 4.5005
R14345 DVDD.n5661 DVDD.n5593 4.5005
R14346 DVDD.n15131 DVDD.n5661 4.5005
R14347 DVDD.n5624 DVDD.n5592 4.5005
R14348 DVDD.n5624 DVDD.n5593 4.5005
R14349 DVDD.n15131 DVDD.n5624 4.5005
R14350 DVDD.n5662 DVDD.n5592 4.5005
R14351 DVDD.n5662 DVDD.n5593 4.5005
R14352 DVDD.n15131 DVDD.n5662 4.5005
R14353 DVDD.n5623 DVDD.n5592 4.5005
R14354 DVDD.n5623 DVDD.n5593 4.5005
R14355 DVDD.n15131 DVDD.n5623 4.5005
R14356 DVDD.n5663 DVDD.n5592 4.5005
R14357 DVDD.n5663 DVDD.n5593 4.5005
R14358 DVDD.n15131 DVDD.n5663 4.5005
R14359 DVDD.n5622 DVDD.n5592 4.5005
R14360 DVDD.n5622 DVDD.n5593 4.5005
R14361 DVDD.n15131 DVDD.n5622 4.5005
R14362 DVDD.n5664 DVDD.n5592 4.5005
R14363 DVDD.n5664 DVDD.n5593 4.5005
R14364 DVDD.n15131 DVDD.n5664 4.5005
R14365 DVDD.n5621 DVDD.n5592 4.5005
R14366 DVDD.n5621 DVDD.n5593 4.5005
R14367 DVDD.n15131 DVDD.n5621 4.5005
R14368 DVDD.n5665 DVDD.n5592 4.5005
R14369 DVDD.n5665 DVDD.n5593 4.5005
R14370 DVDD.n15131 DVDD.n5665 4.5005
R14371 DVDD.n5620 DVDD.n5592 4.5005
R14372 DVDD.n5620 DVDD.n5593 4.5005
R14373 DVDD.n15131 DVDD.n5620 4.5005
R14374 DVDD.n5666 DVDD.n5592 4.5005
R14375 DVDD.n5666 DVDD.n5593 4.5005
R14376 DVDD.n15131 DVDD.n5666 4.5005
R14377 DVDD.n5619 DVDD.n5592 4.5005
R14378 DVDD.n5619 DVDD.n5593 4.5005
R14379 DVDD.n15131 DVDD.n5619 4.5005
R14380 DVDD.n5667 DVDD.n5592 4.5005
R14381 DVDD.n5667 DVDD.n5593 4.5005
R14382 DVDD.n15131 DVDD.n5667 4.5005
R14383 DVDD.n5618 DVDD.n5592 4.5005
R14384 DVDD.n5618 DVDD.n5593 4.5005
R14385 DVDD.n15131 DVDD.n5618 4.5005
R14386 DVDD.n5668 DVDD.n5592 4.5005
R14387 DVDD.n5668 DVDD.n5593 4.5005
R14388 DVDD.n15131 DVDD.n5668 4.5005
R14389 DVDD.n5617 DVDD.n5592 4.5005
R14390 DVDD.n5617 DVDD.n5593 4.5005
R14391 DVDD.n15131 DVDD.n5617 4.5005
R14392 DVDD.n5669 DVDD.n5592 4.5005
R14393 DVDD.n5669 DVDD.n5593 4.5005
R14394 DVDD.n15131 DVDD.n5669 4.5005
R14395 DVDD.n5616 DVDD.n5592 4.5005
R14396 DVDD.n5616 DVDD.n5593 4.5005
R14397 DVDD.n15131 DVDD.n5616 4.5005
R14398 DVDD.n5670 DVDD.n5592 4.5005
R14399 DVDD.n5670 DVDD.n5593 4.5005
R14400 DVDD.n15131 DVDD.n5670 4.5005
R14401 DVDD.n5615 DVDD.n5592 4.5005
R14402 DVDD.n5615 DVDD.n5593 4.5005
R14403 DVDD.n15131 DVDD.n5615 4.5005
R14404 DVDD.n5671 DVDD.n5592 4.5005
R14405 DVDD.n5671 DVDD.n5593 4.5005
R14406 DVDD.n15131 DVDD.n5671 4.5005
R14407 DVDD.n5614 DVDD.n5592 4.5005
R14408 DVDD.n5614 DVDD.n5593 4.5005
R14409 DVDD.n15131 DVDD.n5614 4.5005
R14410 DVDD.n5672 DVDD.n5592 4.5005
R14411 DVDD.n5672 DVDD.n5593 4.5005
R14412 DVDD.n15131 DVDD.n5672 4.5005
R14413 DVDD.n5613 DVDD.n5592 4.5005
R14414 DVDD.n5613 DVDD.n5593 4.5005
R14415 DVDD.n15131 DVDD.n5613 4.5005
R14416 DVDD.n5673 DVDD.n5592 4.5005
R14417 DVDD.n5673 DVDD.n5593 4.5005
R14418 DVDD.n15131 DVDD.n5673 4.5005
R14419 DVDD.n5612 DVDD.n5592 4.5005
R14420 DVDD.n5612 DVDD.n5593 4.5005
R14421 DVDD.n15131 DVDD.n5612 4.5005
R14422 DVDD.n5674 DVDD.n5592 4.5005
R14423 DVDD.n5674 DVDD.n5593 4.5005
R14424 DVDD.n15131 DVDD.n5674 4.5005
R14425 DVDD.n5611 DVDD.n5592 4.5005
R14426 DVDD.n5611 DVDD.n5593 4.5005
R14427 DVDD.n15131 DVDD.n5611 4.5005
R14428 DVDD.n5675 DVDD.n5592 4.5005
R14429 DVDD.n5675 DVDD.n5593 4.5005
R14430 DVDD.n15131 DVDD.n5675 4.5005
R14431 DVDD.n5610 DVDD.n5592 4.5005
R14432 DVDD.n5610 DVDD.n5593 4.5005
R14433 DVDD.n15131 DVDD.n5610 4.5005
R14434 DVDD.n5676 DVDD.n5592 4.5005
R14435 DVDD.n5676 DVDD.n5593 4.5005
R14436 DVDD.n15131 DVDD.n5676 4.5005
R14437 DVDD.n5609 DVDD.n5592 4.5005
R14438 DVDD.n5609 DVDD.n5593 4.5005
R14439 DVDD.n15131 DVDD.n5609 4.5005
R14440 DVDD.n5677 DVDD.n5592 4.5005
R14441 DVDD.n5677 DVDD.n5593 4.5005
R14442 DVDD.n15131 DVDD.n5677 4.5005
R14443 DVDD.n5608 DVDD.n5592 4.5005
R14444 DVDD.n5608 DVDD.n5593 4.5005
R14445 DVDD.n15131 DVDD.n5608 4.5005
R14446 DVDD.n5678 DVDD.n5592 4.5005
R14447 DVDD.n5678 DVDD.n5593 4.5005
R14448 DVDD.n15131 DVDD.n5678 4.5005
R14449 DVDD.n5607 DVDD.n5592 4.5005
R14450 DVDD.n5607 DVDD.n5593 4.5005
R14451 DVDD.n15131 DVDD.n5607 4.5005
R14452 DVDD.n5679 DVDD.n5592 4.5005
R14453 DVDD.n5679 DVDD.n5593 4.5005
R14454 DVDD.n15131 DVDD.n5679 4.5005
R14455 DVDD.n5606 DVDD.n5592 4.5005
R14456 DVDD.n5606 DVDD.n5593 4.5005
R14457 DVDD.n15131 DVDD.n5606 4.5005
R14458 DVDD.n5680 DVDD.n5592 4.5005
R14459 DVDD.n5680 DVDD.n5593 4.5005
R14460 DVDD.n15131 DVDD.n5680 4.5005
R14461 DVDD.n5605 DVDD.n5592 4.5005
R14462 DVDD.n5605 DVDD.n5593 4.5005
R14463 DVDD.n15131 DVDD.n5605 4.5005
R14464 DVDD.n5681 DVDD.n5592 4.5005
R14465 DVDD.n5681 DVDD.n5593 4.5005
R14466 DVDD.n15131 DVDD.n5681 4.5005
R14467 DVDD.n5604 DVDD.n5592 4.5005
R14468 DVDD.n5604 DVDD.n5593 4.5005
R14469 DVDD.n15131 DVDD.n5604 4.5005
R14470 DVDD.n5682 DVDD.n5592 4.5005
R14471 DVDD.n5682 DVDD.n5593 4.5005
R14472 DVDD.n15131 DVDD.n5682 4.5005
R14473 DVDD.n5603 DVDD.n5592 4.5005
R14474 DVDD.n5603 DVDD.n5593 4.5005
R14475 DVDD.n15131 DVDD.n5603 4.5005
R14476 DVDD.n5683 DVDD.n5592 4.5005
R14477 DVDD.n5683 DVDD.n5593 4.5005
R14478 DVDD.n15131 DVDD.n5683 4.5005
R14479 DVDD.n5602 DVDD.n5592 4.5005
R14480 DVDD.n5602 DVDD.n5593 4.5005
R14481 DVDD.n15131 DVDD.n5602 4.5005
R14482 DVDD.n5684 DVDD.n5592 4.5005
R14483 DVDD.n5684 DVDD.n5593 4.5005
R14484 DVDD.n15131 DVDD.n5684 4.5005
R14485 DVDD.n5601 DVDD.n5592 4.5005
R14486 DVDD.n5601 DVDD.n5593 4.5005
R14487 DVDD.n15131 DVDD.n5601 4.5005
R14488 DVDD.n5685 DVDD.n5592 4.5005
R14489 DVDD.n5685 DVDD.n5593 4.5005
R14490 DVDD.n15131 DVDD.n5685 4.5005
R14491 DVDD.n5600 DVDD.n5592 4.5005
R14492 DVDD.n5600 DVDD.n5593 4.5005
R14493 DVDD.n15131 DVDD.n5600 4.5005
R14494 DVDD.n5686 DVDD.n5592 4.5005
R14495 DVDD.n5686 DVDD.n5593 4.5005
R14496 DVDD.n15131 DVDD.n5686 4.5005
R14497 DVDD.n5599 DVDD.n5592 4.5005
R14498 DVDD.n5599 DVDD.n5593 4.5005
R14499 DVDD.n15131 DVDD.n5599 4.5005
R14500 DVDD.n5687 DVDD.n5592 4.5005
R14501 DVDD.n5687 DVDD.n5593 4.5005
R14502 DVDD.n15131 DVDD.n5687 4.5005
R14503 DVDD.n5598 DVDD.n5592 4.5005
R14504 DVDD.n5598 DVDD.n5593 4.5005
R14505 DVDD.n15131 DVDD.n5598 4.5005
R14506 DVDD.n5688 DVDD.n5592 4.5005
R14507 DVDD.n5688 DVDD.n5593 4.5005
R14508 DVDD.n15131 DVDD.n5688 4.5005
R14509 DVDD.n5597 DVDD.n5592 4.5005
R14510 DVDD.n5597 DVDD.n5593 4.5005
R14511 DVDD.n15131 DVDD.n5597 4.5005
R14512 DVDD.n5689 DVDD.n5592 4.5005
R14513 DVDD.n5689 DVDD.n5593 4.5005
R14514 DVDD.n15131 DVDD.n5689 4.5005
R14515 DVDD.n5596 DVDD.n5592 4.5005
R14516 DVDD.n5596 DVDD.n5593 4.5005
R14517 DVDD.n15131 DVDD.n5596 4.5005
R14518 DVDD.n5690 DVDD.n5592 4.5005
R14519 DVDD.n5690 DVDD.n5593 4.5005
R14520 DVDD.n15131 DVDD.n5690 4.5005
R14521 DVDD.n5595 DVDD.n5592 4.5005
R14522 DVDD.n5595 DVDD.n5593 4.5005
R14523 DVDD.n15131 DVDD.n5595 4.5005
R14524 DVDD.n5691 DVDD.n5592 4.5005
R14525 DVDD.n5691 DVDD.n5593 4.5005
R14526 DVDD.n15131 DVDD.n5691 4.5005
R14527 DVDD.n5594 DVDD.n5592 4.5005
R14528 DVDD.n5594 DVDD.n5593 4.5005
R14529 DVDD.n15131 DVDD.n5594 4.5005
R14530 DVDD.n15130 DVDD.n5592 4.5005
R14531 DVDD.n15130 DVDD.n5740 4.5005
R14532 DVDD.n15130 DVDD.n5593 4.5005
R14533 DVDD.n15131 DVDD.n15130 4.5005
R14534 DVDD.n17711 DVDD.n17308 4.5005
R14535 DVDD.n17711 DVDD.n17307 4.5005
R14536 DVDD.n17711 DVDD.n17309 4.5005
R14537 DVDD.n17711 DVDD.n17306 4.5005
R14538 DVDD.n17711 DVDD.n17710 4.5005
R14539 DVDD.n5643 DVDD.n5592 4.5005
R14540 DVDD.n6696 DVDD.n6404 4.5005
R14541 DVDD.n6696 DVDD.n6695 4.5005
R14542 DVDD.n963 DVDD.n915 4.5005
R14543 DVDD.n1068 DVDD.n915 4.5005
R14544 DVDD.n15112 DVDD.n6042 4.5005
R14545 DVDD.n15112 DVDD.n15111 4.5005
R14546 DVDD.n17726 DVDD.n892 4.5005
R14547 DVDD.n892 DVDD.n890 4.5005
R14548 DVDD.n17724 DVDD.n892 4.5005
R14549 DVDD.n5587 DVDD.n5582 4.5005
R14550 DVDD.n5587 DVDD.n5577 4.5005
R14551 DVDD.n15139 DVDD.n5587 4.5005
R14552 DVDD.n896 DVDD.n894 4.5005
R14553 DVDD.n900 DVDD.n894 4.5005
R14554 DVDD.n17726 DVDD.n894 4.5005
R14555 DVDD.n894 DVDD.n890 4.5005
R14556 DVDD.n17724 DVDD.n894 4.5005
R14557 DVDD.n15141 DVDD.n5580 4.5005
R14558 DVDD.n5580 DVDD.n5577 4.5005
R14559 DVDD.n15139 DVDD.n5580 4.5005
R14560 DVDD.n896 DVDD.n891 4.5005
R14561 DVDD.n900 DVDD.n891 4.5005
R14562 DVDD.n17726 DVDD.n891 4.5005
R14563 DVDD.n891 DVDD.n890 4.5005
R14564 DVDD.n17724 DVDD.n891 4.5005
R14565 DVDD.n5582 DVDD.n5578 4.5005
R14566 DVDD.n5586 DVDD.n5578 4.5005
R14567 DVDD.n15141 DVDD.n5578 4.5005
R14568 DVDD.n5578 DVDD.n5577 4.5005
R14569 DVDD.n15139 DVDD.n5578 4.5005
R14570 DVDD.n17725 DVDD.n896 4.5005
R14571 DVDD.n17725 DVDD.n900 4.5005
R14572 DVDD.n17726 DVDD.n17725 4.5005
R14573 DVDD.n17725 DVDD.n890 4.5005
R14574 DVDD.n17725 DVDD.n17724 4.5005
R14575 DVDD.n15140 DVDD.n5582 4.5005
R14576 DVDD.n15140 DVDD.n5586 4.5005
R14577 DVDD.n15141 DVDD.n15140 4.5005
R14578 DVDD.n15140 DVDD.n5577 4.5005
R14579 DVDD.n15140 DVDD.n15139 4.5005
R14580 DVDD.n10200 DVDD.n9572 4.5005
R14581 DVDD.n10203 DVDD.n9572 4.5005
R14582 DVDD.n10177 DVDD.n8972 4.5005
R14583 DVDD.n10200 DVDD.n8972 4.5005
R14584 DVDD.n10203 DVDD.n8972 4.5005
R14585 DVDD.n10202 DVDD.n10177 4.5005
R14586 DVDD.n10202 DVDD.n10175 4.5005
R14587 DVDD.n10202 DVDD.n10180 4.5005
R14588 DVDD.n10202 DVDD.n10174 4.5005
R14589 DVDD.n10202 DVDD.n10183 4.5005
R14590 DVDD.n10202 DVDD.n10173 4.5005
R14591 DVDD.n10202 DVDD.n10186 4.5005
R14592 DVDD.n10202 DVDD.n10172 4.5005
R14593 DVDD.n10202 DVDD.n10189 4.5005
R14594 DVDD.n10202 DVDD.n10171 4.5005
R14595 DVDD.n10202 DVDD.n10192 4.5005
R14596 DVDD.n10202 DVDD.n10170 4.5005
R14597 DVDD.n10202 DVDD.n10195 4.5005
R14598 DVDD.n10202 DVDD.n10169 4.5005
R14599 DVDD.n10202 DVDD.n10197 4.5005
R14600 DVDD.n10203 DVDD.n10202 4.5005
R14601 DVDD.n4979 DVDD.n3488 4.5005
R14602 DVDD.n4981 DVDD.n3473 4.5005
R14603 DVDD.n4981 DVDD.n4980 4.5005
R14604 DVDD.n4980 DVDD.n4916 4.5005
R14605 DVDD.n4980 DVDD.n4919 4.5005
R14606 DVDD.n4980 DVDD.n4915 4.5005
R14607 DVDD.n4980 DVDD.n4922 4.5005
R14608 DVDD.n4980 DVDD.n4914 4.5005
R14609 DVDD.n4980 DVDD.n4925 4.5005
R14610 DVDD.n4980 DVDD.n4913 4.5005
R14611 DVDD.n4980 DVDD.n4928 4.5005
R14612 DVDD.n4980 DVDD.n4912 4.5005
R14613 DVDD.n4980 DVDD.n4931 4.5005
R14614 DVDD.n4980 DVDD.n4911 4.5005
R14615 DVDD.n4980 DVDD.n4934 4.5005
R14616 DVDD.n4980 DVDD.n4910 4.5005
R14617 DVDD.n4980 DVDD.n4937 4.5005
R14618 DVDD.n4980 DVDD.n4909 4.5005
R14619 DVDD.n4980 DVDD.n4940 4.5005
R14620 DVDD.n4980 DVDD.n4908 4.5005
R14621 DVDD.n4980 DVDD.n4979 4.5005
R14622 DVDD.n21013 DVDD.n18703 4.5005
R14623 DVDD.n20983 DVDD.n18703 4.5005
R14624 DVDD.n21013 DVDD.n21012 4.5005
R14625 DVDD.n21012 DVDD.n20991 4.5005
R14626 DVDD.n21012 DVDD.n20989 4.5005
R14627 DVDD.n21012 DVDD.n20994 4.5005
R14628 DVDD.n21012 DVDD.n20988 4.5005
R14629 DVDD.n21012 DVDD.n20997 4.5005
R14630 DVDD.n21012 DVDD.n20987 4.5005
R14631 DVDD.n21012 DVDD.n21000 4.5005
R14632 DVDD.n21012 DVDD.n20986 4.5005
R14633 DVDD.n21012 DVDD.n21003 4.5005
R14634 DVDD.n21012 DVDD.n20985 4.5005
R14635 DVDD.n21012 DVDD.n21006 4.5005
R14636 DVDD.n21012 DVDD.n20984 4.5005
R14637 DVDD.n21012 DVDD.n21009 4.5005
R14638 DVDD.n21012 DVDD.n20983 4.5005
R14639 DVDD.n20978 DVDD.n18762 4.5005
R14640 DVDD.n20979 DVDD.n20978 4.5005
R14641 DVDD.n20981 DVDD.n20978 4.5005
R14642 DVDD.n20982 DVDD.n20981 4.5005
R14643 DVDD.n20532 DVDD.n20531 4.5005
R14644 DVDD.n20531 DVDD.n20524 4.5005
R14645 DVDD.n20531 DVDD.n20530 4.5005
R14646 DVDD.n20530 DVDD.n20529 4.5005
R14647 DVDD.n20519 DVDD.n18822 4.5005
R14648 DVDD.n20519 DVDD.n20488 4.5005
R14649 DVDD.n20516 DVDD.n18822 4.5005
R14650 DVDD.n20517 DVDD.n20516 4.5005
R14651 DVDD.n20516 DVDD.n20503 4.5005
R14652 DVDD.n20516 DVDD.n20505 4.5005
R14653 DVDD.n20516 DVDD.n20502 4.5005
R14654 DVDD.n20516 DVDD.n20507 4.5005
R14655 DVDD.n20516 DVDD.n20501 4.5005
R14656 DVDD.n20516 DVDD.n20509 4.5005
R14657 DVDD.n20516 DVDD.n20500 4.5005
R14658 DVDD.n20516 DVDD.n20511 4.5005
R14659 DVDD.n20516 DVDD.n20499 4.5005
R14660 DVDD.n20516 DVDD.n20513 4.5005
R14661 DVDD.n20516 DVDD.n20498 4.5005
R14662 DVDD.n20516 DVDD.n20515 4.5005
R14663 DVDD.n20516 DVDD.n20488 4.5005
R14664 DVDD.n20516 DVDD.n20496 4.5005
R14665 DVDD.n21012 DVDD.n21011 4.5005
R14666 DVDD.n9763 DVDD.n9610 4.5005
R14667 DVDD.n9764 DVDD.n9610 4.5005
R14668 DVDD.n9762 DVDD.n9610 4.5005
R14669 DVDD.n9765 DVDD.n9610 4.5005
R14670 DVDD.n9761 DVDD.n9610 4.5005
R14671 DVDD.n9768 DVDD.n9610 4.5005
R14672 DVDD.n9759 DVDD.n9610 4.5005
R14673 DVDD.n9769 DVDD.n9610 4.5005
R14674 DVDD.n9758 DVDD.n9610 4.5005
R14675 DVDD.n9770 DVDD.n9610 4.5005
R14676 DVDD.n9939 DVDD.n9610 4.5005
R14677 DVDD.n9948 DVDD.n9610 4.5005
R14678 DVDD.n9806 DVDD.n9763 4.5005
R14679 DVDD.n9806 DVDD.n9764 4.5005
R14680 DVDD.n9806 DVDD.n9762 4.5005
R14681 DVDD.n9806 DVDD.n9765 4.5005
R14682 DVDD.n9806 DVDD.n9761 4.5005
R14683 DVDD.n9806 DVDD.n9767 4.5005
R14684 DVDD.n9806 DVDD.n9760 4.5005
R14685 DVDD.n9806 DVDD.n9768 4.5005
R14686 DVDD.n9806 DVDD.n9759 4.5005
R14687 DVDD.n9806 DVDD.n9769 4.5005
R14688 DVDD.n9806 DVDD.n9758 4.5005
R14689 DVDD.n9806 DVDD.n9770 4.5005
R14690 DVDD.n9806 DVDD.n9772 4.5005
R14691 DVDD.n9948 DVDD.n9806 4.5005
R14692 DVDD.n9809 DVDD.n9763 4.5005
R14693 DVDD.n9809 DVDD.n9764 4.5005
R14694 DVDD.n9809 DVDD.n9762 4.5005
R14695 DVDD.n9809 DVDD.n9765 4.5005
R14696 DVDD.n9809 DVDD.n9761 4.5005
R14697 DVDD.n9809 DVDD.n9767 4.5005
R14698 DVDD.n9809 DVDD.n9760 4.5005
R14699 DVDD.n9809 DVDD.n9768 4.5005
R14700 DVDD.n9809 DVDD.n9759 4.5005
R14701 DVDD.n9809 DVDD.n9769 4.5005
R14702 DVDD.n9809 DVDD.n9758 4.5005
R14703 DVDD.n9809 DVDD.n9770 4.5005
R14704 DVDD.n9809 DVDD.n9772 4.5005
R14705 DVDD.n9948 DVDD.n9809 4.5005
R14706 DVDD.n9805 DVDD.n9763 4.5005
R14707 DVDD.n9805 DVDD.n9764 4.5005
R14708 DVDD.n9805 DVDD.n9762 4.5005
R14709 DVDD.n9805 DVDD.n9765 4.5005
R14710 DVDD.n9805 DVDD.n9761 4.5005
R14711 DVDD.n9805 DVDD.n9767 4.5005
R14712 DVDD.n9805 DVDD.n9760 4.5005
R14713 DVDD.n9805 DVDD.n9768 4.5005
R14714 DVDD.n9805 DVDD.n9759 4.5005
R14715 DVDD.n9805 DVDD.n9769 4.5005
R14716 DVDD.n9805 DVDD.n9758 4.5005
R14717 DVDD.n9805 DVDD.n9770 4.5005
R14718 DVDD.n9805 DVDD.n9772 4.5005
R14719 DVDD.n9805 DVDD.n9757 4.5005
R14720 DVDD.n9948 DVDD.n9805 4.5005
R14721 DVDD.n9811 DVDD.n9763 4.5005
R14722 DVDD.n9811 DVDD.n9764 4.5005
R14723 DVDD.n9811 DVDD.n9762 4.5005
R14724 DVDD.n9811 DVDD.n9765 4.5005
R14725 DVDD.n9811 DVDD.n9761 4.5005
R14726 DVDD.n9811 DVDD.n9767 4.5005
R14727 DVDD.n9811 DVDD.n9760 4.5005
R14728 DVDD.n9811 DVDD.n9768 4.5005
R14729 DVDD.n9811 DVDD.n9759 4.5005
R14730 DVDD.n9811 DVDD.n9769 4.5005
R14731 DVDD.n9811 DVDD.n9758 4.5005
R14732 DVDD.n9811 DVDD.n9770 4.5005
R14733 DVDD.n9811 DVDD.n9772 4.5005
R14734 DVDD.n9948 DVDD.n9811 4.5005
R14735 DVDD.n9797 DVDD.n9763 4.5005
R14736 DVDD.n9797 DVDD.n9764 4.5005
R14737 DVDD.n9797 DVDD.n9762 4.5005
R14738 DVDD.n9797 DVDD.n9765 4.5005
R14739 DVDD.n9797 DVDD.n9761 4.5005
R14740 DVDD.n9797 DVDD.n9767 4.5005
R14741 DVDD.n9797 DVDD.n9760 4.5005
R14742 DVDD.n9797 DVDD.n9768 4.5005
R14743 DVDD.n9797 DVDD.n9759 4.5005
R14744 DVDD.n9797 DVDD.n9769 4.5005
R14745 DVDD.n9797 DVDD.n9758 4.5005
R14746 DVDD.n9797 DVDD.n9770 4.5005
R14747 DVDD.n9797 DVDD.n9772 4.5005
R14748 DVDD.n9948 DVDD.n9797 4.5005
R14749 DVDD.n9812 DVDD.n9763 4.5005
R14750 DVDD.n9812 DVDD.n9764 4.5005
R14751 DVDD.n9812 DVDD.n9762 4.5005
R14752 DVDD.n9812 DVDD.n9765 4.5005
R14753 DVDD.n9812 DVDD.n9761 4.5005
R14754 DVDD.n9812 DVDD.n9767 4.5005
R14755 DVDD.n9812 DVDD.n9760 4.5005
R14756 DVDD.n9812 DVDD.n9768 4.5005
R14757 DVDD.n9812 DVDD.n9759 4.5005
R14758 DVDD.n9812 DVDD.n9769 4.5005
R14759 DVDD.n9812 DVDD.n9758 4.5005
R14760 DVDD.n9812 DVDD.n9770 4.5005
R14761 DVDD.n9812 DVDD.n9772 4.5005
R14762 DVDD.n9812 DVDD.n9757 4.5005
R14763 DVDD.n9948 DVDD.n9812 4.5005
R14764 DVDD.n9796 DVDD.n9763 4.5005
R14765 DVDD.n9796 DVDD.n9764 4.5005
R14766 DVDD.n9796 DVDD.n9762 4.5005
R14767 DVDD.n9796 DVDD.n9765 4.5005
R14768 DVDD.n9796 DVDD.n9761 4.5005
R14769 DVDD.n9796 DVDD.n9767 4.5005
R14770 DVDD.n9796 DVDD.n9760 4.5005
R14771 DVDD.n9796 DVDD.n9768 4.5005
R14772 DVDD.n9796 DVDD.n9759 4.5005
R14773 DVDD.n9796 DVDD.n9769 4.5005
R14774 DVDD.n9796 DVDD.n9758 4.5005
R14775 DVDD.n9796 DVDD.n9770 4.5005
R14776 DVDD.n9939 DVDD.n9796 4.5005
R14777 DVDD.n9796 DVDD.n9772 4.5005
R14778 DVDD.n9948 DVDD.n9796 4.5005
R14779 DVDD.n3136 DVDD.n3115 4.5005
R14780 DVDD.n3136 DVDD.n3116 4.5005
R14781 DVDD.n3136 DVDD.n3114 4.5005
R14782 DVDD.n3136 DVDD.n3117 4.5005
R14783 DVDD.n3136 DVDD.n3113 4.5005
R14784 DVDD.n3136 DVDD.n3119 4.5005
R14785 DVDD.n3136 DVDD.n3111 4.5005
R14786 DVDD.n3136 DVDD.n3120 4.5005
R14787 DVDD.n3136 DVDD.n3110 4.5005
R14788 DVDD.n3136 DVDD.n3121 4.5005
R14789 DVDD.n3136 DVDD.n3109 4.5005
R14790 DVDD.n3136 DVDD.n3122 4.5005
R14791 DVDD.n16067 DVDD.n3136 4.5005
R14792 DVDD.n16008 DVDD.n3115 4.5005
R14793 DVDD.n16008 DVDD.n3116 4.5005
R14794 DVDD.n16008 DVDD.n3114 4.5005
R14795 DVDD.n16008 DVDD.n3117 4.5005
R14796 DVDD.n16008 DVDD.n3113 4.5005
R14797 DVDD.n16008 DVDD.n3118 4.5005
R14798 DVDD.n16008 DVDD.n3112 4.5005
R14799 DVDD.n16008 DVDD.n3119 4.5005
R14800 DVDD.n16008 DVDD.n3111 4.5005
R14801 DVDD.n16008 DVDD.n3120 4.5005
R14802 DVDD.n16008 DVDD.n3110 4.5005
R14803 DVDD.n16008 DVDD.n3121 4.5005
R14804 DVDD.n16008 DVDD.n3122 4.5005
R14805 DVDD.n16067 DVDD.n16008 4.5005
R14806 DVDD.n3134 DVDD.n3115 4.5005
R14807 DVDD.n3134 DVDD.n3116 4.5005
R14808 DVDD.n3134 DVDD.n3114 4.5005
R14809 DVDD.n3134 DVDD.n3117 4.5005
R14810 DVDD.n3134 DVDD.n3113 4.5005
R14811 DVDD.n3134 DVDD.n3118 4.5005
R14812 DVDD.n3134 DVDD.n3112 4.5005
R14813 DVDD.n3134 DVDD.n3119 4.5005
R14814 DVDD.n3134 DVDD.n3111 4.5005
R14815 DVDD.n3134 DVDD.n3120 4.5005
R14816 DVDD.n3134 DVDD.n3110 4.5005
R14817 DVDD.n3134 DVDD.n3121 4.5005
R14818 DVDD.n16067 DVDD.n3134 4.5005
R14819 DVDD.n16009 DVDD.n3115 4.5005
R14820 DVDD.n16009 DVDD.n3116 4.5005
R14821 DVDD.n16009 DVDD.n3114 4.5005
R14822 DVDD.n16009 DVDD.n3117 4.5005
R14823 DVDD.n16009 DVDD.n3113 4.5005
R14824 DVDD.n16009 DVDD.n3118 4.5005
R14825 DVDD.n16009 DVDD.n3112 4.5005
R14826 DVDD.n16009 DVDD.n3119 4.5005
R14827 DVDD.n16009 DVDD.n3111 4.5005
R14828 DVDD.n16009 DVDD.n3120 4.5005
R14829 DVDD.n16009 DVDD.n3110 4.5005
R14830 DVDD.n16009 DVDD.n3121 4.5005
R14831 DVDD.n16009 DVDD.n3122 4.5005
R14832 DVDD.n16067 DVDD.n16009 4.5005
R14833 DVDD.n3133 DVDD.n3115 4.5005
R14834 DVDD.n3133 DVDD.n3116 4.5005
R14835 DVDD.n3133 DVDD.n3114 4.5005
R14836 DVDD.n3133 DVDD.n3117 4.5005
R14837 DVDD.n3133 DVDD.n3113 4.5005
R14838 DVDD.n3133 DVDD.n3118 4.5005
R14839 DVDD.n3133 DVDD.n3112 4.5005
R14840 DVDD.n3133 DVDD.n3119 4.5005
R14841 DVDD.n3133 DVDD.n3111 4.5005
R14842 DVDD.n3133 DVDD.n3120 4.5005
R14843 DVDD.n3133 DVDD.n3110 4.5005
R14844 DVDD.n3133 DVDD.n3121 4.5005
R14845 DVDD.n3133 DVDD.n3122 4.5005
R14846 DVDD.n16067 DVDD.n3133 4.5005
R14847 DVDD.n16018 DVDD.n3115 4.5005
R14848 DVDD.n16018 DVDD.n3116 4.5005
R14849 DVDD.n16018 DVDD.n3114 4.5005
R14850 DVDD.n16018 DVDD.n3117 4.5005
R14851 DVDD.n16018 DVDD.n3113 4.5005
R14852 DVDD.n16018 DVDD.n3118 4.5005
R14853 DVDD.n16018 DVDD.n3112 4.5005
R14854 DVDD.n16018 DVDD.n3119 4.5005
R14855 DVDD.n16018 DVDD.n3111 4.5005
R14856 DVDD.n16018 DVDD.n3120 4.5005
R14857 DVDD.n16018 DVDD.n3110 4.5005
R14858 DVDD.n16018 DVDD.n3121 4.5005
R14859 DVDD.n16018 DVDD.n3122 4.5005
R14860 DVDD.n16061 DVDD.n16018 4.5005
R14861 DVDD.n16067 DVDD.n16018 4.5005
R14862 DVDD.n3132 DVDD.n3115 4.5005
R14863 DVDD.n3132 DVDD.n3116 4.5005
R14864 DVDD.n3132 DVDD.n3114 4.5005
R14865 DVDD.n3132 DVDD.n3117 4.5005
R14866 DVDD.n3132 DVDD.n3113 4.5005
R14867 DVDD.n3132 DVDD.n3118 4.5005
R14868 DVDD.n3132 DVDD.n3112 4.5005
R14869 DVDD.n3132 DVDD.n3119 4.5005
R14870 DVDD.n3132 DVDD.n3111 4.5005
R14871 DVDD.n3132 DVDD.n3120 4.5005
R14872 DVDD.n3132 DVDD.n3110 4.5005
R14873 DVDD.n3132 DVDD.n3121 4.5005
R14874 DVDD.n3132 DVDD.n3122 4.5005
R14875 DVDD.n16067 DVDD.n3132 4.5005
R14876 DVDD.n16020 DVDD.n3115 4.5005
R14877 DVDD.n16020 DVDD.n3116 4.5005
R14878 DVDD.n16020 DVDD.n3114 4.5005
R14879 DVDD.n16020 DVDD.n3117 4.5005
R14880 DVDD.n16020 DVDD.n3113 4.5005
R14881 DVDD.n16020 DVDD.n3118 4.5005
R14882 DVDD.n16020 DVDD.n3112 4.5005
R14883 DVDD.n16020 DVDD.n3119 4.5005
R14884 DVDD.n16020 DVDD.n3111 4.5005
R14885 DVDD.n16020 DVDD.n3120 4.5005
R14886 DVDD.n16020 DVDD.n3110 4.5005
R14887 DVDD.n16020 DVDD.n3121 4.5005
R14888 DVDD.n16020 DVDD.n3122 4.5005
R14889 DVDD.n16067 DVDD.n16020 4.5005
R14890 DVDD.n3130 DVDD.n3115 4.5005
R14891 DVDD.n3130 DVDD.n3116 4.5005
R14892 DVDD.n3130 DVDD.n3114 4.5005
R14893 DVDD.n3130 DVDD.n3117 4.5005
R14894 DVDD.n3130 DVDD.n3113 4.5005
R14895 DVDD.n3130 DVDD.n3118 4.5005
R14896 DVDD.n3130 DVDD.n3112 4.5005
R14897 DVDD.n3130 DVDD.n3119 4.5005
R14898 DVDD.n3130 DVDD.n3111 4.5005
R14899 DVDD.n3130 DVDD.n3120 4.5005
R14900 DVDD.n3130 DVDD.n3110 4.5005
R14901 DVDD.n3130 DVDD.n3121 4.5005
R14902 DVDD.n3130 DVDD.n3122 4.5005
R14903 DVDD.n16061 DVDD.n3130 4.5005
R14904 DVDD.n16067 DVDD.n3130 4.5005
R14905 DVDD.n16021 DVDD.n3115 4.5005
R14906 DVDD.n16021 DVDD.n3116 4.5005
R14907 DVDD.n16021 DVDD.n3114 4.5005
R14908 DVDD.n16021 DVDD.n3117 4.5005
R14909 DVDD.n16021 DVDD.n3113 4.5005
R14910 DVDD.n16021 DVDD.n3118 4.5005
R14911 DVDD.n16021 DVDD.n3112 4.5005
R14912 DVDD.n16021 DVDD.n3119 4.5005
R14913 DVDD.n16021 DVDD.n3111 4.5005
R14914 DVDD.n16021 DVDD.n3120 4.5005
R14915 DVDD.n16021 DVDD.n3110 4.5005
R14916 DVDD.n16021 DVDD.n3121 4.5005
R14917 DVDD.n16021 DVDD.n3122 4.5005
R14918 DVDD.n16067 DVDD.n16021 4.5005
R14919 DVDD.n3129 DVDD.n3115 4.5005
R14920 DVDD.n3129 DVDD.n3116 4.5005
R14921 DVDD.n3129 DVDD.n3114 4.5005
R14922 DVDD.n3129 DVDD.n3117 4.5005
R14923 DVDD.n3129 DVDD.n3113 4.5005
R14924 DVDD.n3129 DVDD.n3118 4.5005
R14925 DVDD.n3129 DVDD.n3112 4.5005
R14926 DVDD.n3129 DVDD.n3119 4.5005
R14927 DVDD.n3129 DVDD.n3111 4.5005
R14928 DVDD.n3129 DVDD.n3120 4.5005
R14929 DVDD.n3129 DVDD.n3110 4.5005
R14930 DVDD.n3129 DVDD.n3121 4.5005
R14931 DVDD.n3129 DVDD.n3122 4.5005
R14932 DVDD.n16067 DVDD.n3129 4.5005
R14933 DVDD.n16030 DVDD.n3115 4.5005
R14934 DVDD.n16030 DVDD.n3116 4.5005
R14935 DVDD.n16030 DVDD.n3114 4.5005
R14936 DVDD.n16030 DVDD.n3117 4.5005
R14937 DVDD.n16030 DVDD.n3113 4.5005
R14938 DVDD.n16030 DVDD.n3118 4.5005
R14939 DVDD.n16030 DVDD.n3112 4.5005
R14940 DVDD.n16030 DVDD.n3119 4.5005
R14941 DVDD.n16030 DVDD.n3111 4.5005
R14942 DVDD.n16030 DVDD.n3120 4.5005
R14943 DVDD.n16030 DVDD.n3110 4.5005
R14944 DVDD.n16030 DVDD.n3121 4.5005
R14945 DVDD.n16030 DVDD.n3122 4.5005
R14946 DVDD.n16061 DVDD.n16030 4.5005
R14947 DVDD.n16067 DVDD.n16030 4.5005
R14948 DVDD.n3128 DVDD.n3115 4.5005
R14949 DVDD.n3128 DVDD.n3116 4.5005
R14950 DVDD.n3128 DVDD.n3114 4.5005
R14951 DVDD.n3128 DVDD.n3117 4.5005
R14952 DVDD.n3128 DVDD.n3113 4.5005
R14953 DVDD.n3128 DVDD.n3118 4.5005
R14954 DVDD.n3128 DVDD.n3112 4.5005
R14955 DVDD.n3128 DVDD.n3119 4.5005
R14956 DVDD.n3128 DVDD.n3111 4.5005
R14957 DVDD.n3128 DVDD.n3120 4.5005
R14958 DVDD.n3128 DVDD.n3110 4.5005
R14959 DVDD.n3128 DVDD.n3121 4.5005
R14960 DVDD.n3128 DVDD.n3109 4.5005
R14961 DVDD.n3128 DVDD.n3122 4.5005
R14962 DVDD.n16067 DVDD.n3128 4.5005
R14963 DVDD.n16032 DVDD.n3115 4.5005
R14964 DVDD.n16032 DVDD.n3116 4.5005
R14965 DVDD.n16032 DVDD.n3114 4.5005
R14966 DVDD.n16032 DVDD.n3117 4.5005
R14967 DVDD.n16032 DVDD.n3113 4.5005
R14968 DVDD.n16032 DVDD.n3118 4.5005
R14969 DVDD.n16032 DVDD.n3112 4.5005
R14970 DVDD.n16032 DVDD.n3119 4.5005
R14971 DVDD.n16032 DVDD.n3111 4.5005
R14972 DVDD.n16032 DVDD.n3120 4.5005
R14973 DVDD.n16032 DVDD.n3110 4.5005
R14974 DVDD.n16032 DVDD.n3121 4.5005
R14975 DVDD.n16032 DVDD.n3122 4.5005
R14976 DVDD.n16067 DVDD.n16032 4.5005
R14977 DVDD.n3127 DVDD.n3115 4.5005
R14978 DVDD.n3127 DVDD.n3116 4.5005
R14979 DVDD.n3127 DVDD.n3114 4.5005
R14980 DVDD.n3127 DVDD.n3117 4.5005
R14981 DVDD.n3127 DVDD.n3113 4.5005
R14982 DVDD.n3127 DVDD.n3118 4.5005
R14983 DVDD.n3127 DVDD.n3112 4.5005
R14984 DVDD.n3127 DVDD.n3119 4.5005
R14985 DVDD.n3127 DVDD.n3111 4.5005
R14986 DVDD.n3127 DVDD.n3120 4.5005
R14987 DVDD.n3127 DVDD.n3110 4.5005
R14988 DVDD.n3127 DVDD.n3121 4.5005
R14989 DVDD.n3127 DVDD.n3122 4.5005
R14990 DVDD.n16067 DVDD.n3127 4.5005
R14991 DVDD.n16040 DVDD.n3115 4.5005
R14992 DVDD.n16040 DVDD.n3116 4.5005
R14993 DVDD.n16040 DVDD.n3114 4.5005
R14994 DVDD.n16040 DVDD.n3117 4.5005
R14995 DVDD.n16040 DVDD.n3113 4.5005
R14996 DVDD.n16040 DVDD.n3118 4.5005
R14997 DVDD.n16040 DVDD.n3112 4.5005
R14998 DVDD.n16040 DVDD.n3119 4.5005
R14999 DVDD.n16040 DVDD.n3111 4.5005
R15000 DVDD.n16040 DVDD.n3120 4.5005
R15001 DVDD.n16040 DVDD.n3110 4.5005
R15002 DVDD.n16040 DVDD.n3121 4.5005
R15003 DVDD.n16040 DVDD.n3109 4.5005
R15004 DVDD.n16040 DVDD.n3122 4.5005
R15005 DVDD.n16067 DVDD.n16040 4.5005
R15006 DVDD.n3126 DVDD.n3115 4.5005
R15007 DVDD.n3126 DVDD.n3116 4.5005
R15008 DVDD.n3126 DVDD.n3114 4.5005
R15009 DVDD.n3126 DVDD.n3117 4.5005
R15010 DVDD.n3126 DVDD.n3113 4.5005
R15011 DVDD.n3126 DVDD.n3118 4.5005
R15012 DVDD.n3126 DVDD.n3112 4.5005
R15013 DVDD.n3126 DVDD.n3119 4.5005
R15014 DVDD.n3126 DVDD.n3111 4.5005
R15015 DVDD.n3126 DVDD.n3120 4.5005
R15016 DVDD.n3126 DVDD.n3110 4.5005
R15017 DVDD.n3126 DVDD.n3121 4.5005
R15018 DVDD.n3126 DVDD.n3109 4.5005
R15019 DVDD.n3126 DVDD.n3122 4.5005
R15020 DVDD.n16067 DVDD.n3126 4.5005
R15021 DVDD.n16042 DVDD.n3115 4.5005
R15022 DVDD.n16042 DVDD.n3116 4.5005
R15023 DVDD.n16042 DVDD.n3114 4.5005
R15024 DVDD.n16042 DVDD.n3117 4.5005
R15025 DVDD.n16042 DVDD.n3113 4.5005
R15026 DVDD.n16042 DVDD.n3118 4.5005
R15027 DVDD.n16042 DVDD.n3112 4.5005
R15028 DVDD.n16042 DVDD.n3119 4.5005
R15029 DVDD.n16042 DVDD.n3111 4.5005
R15030 DVDD.n16042 DVDD.n3120 4.5005
R15031 DVDD.n16042 DVDD.n3110 4.5005
R15032 DVDD.n16042 DVDD.n3121 4.5005
R15033 DVDD.n16042 DVDD.n3122 4.5005
R15034 DVDD.n16067 DVDD.n16042 4.5005
R15035 DVDD.n3125 DVDD.n3115 4.5005
R15036 DVDD.n3125 DVDD.n3116 4.5005
R15037 DVDD.n3125 DVDD.n3114 4.5005
R15038 DVDD.n3125 DVDD.n3117 4.5005
R15039 DVDD.n3125 DVDD.n3113 4.5005
R15040 DVDD.n3125 DVDD.n3118 4.5005
R15041 DVDD.n3125 DVDD.n3112 4.5005
R15042 DVDD.n3125 DVDD.n3119 4.5005
R15043 DVDD.n3125 DVDD.n3111 4.5005
R15044 DVDD.n3125 DVDD.n3120 4.5005
R15045 DVDD.n3125 DVDD.n3110 4.5005
R15046 DVDD.n3125 DVDD.n3121 4.5005
R15047 DVDD.n3125 DVDD.n3122 4.5005
R15048 DVDD.n16067 DVDD.n3125 4.5005
R15049 DVDD.n16068 DVDD.n3115 4.5005
R15050 DVDD.n16068 DVDD.n3116 4.5005
R15051 DVDD.n16068 DVDD.n3114 4.5005
R15052 DVDD.n16068 DVDD.n3117 4.5005
R15053 DVDD.n16068 DVDD.n3113 4.5005
R15054 DVDD.n16068 DVDD.n3118 4.5005
R15055 DVDD.n16068 DVDD.n3112 4.5005
R15056 DVDD.n16068 DVDD.n3119 4.5005
R15057 DVDD.n16068 DVDD.n3111 4.5005
R15058 DVDD.n16068 DVDD.n3120 4.5005
R15059 DVDD.n16068 DVDD.n3110 4.5005
R15060 DVDD.n16068 DVDD.n3121 4.5005
R15061 DVDD.n16068 DVDD.n3109 4.5005
R15062 DVDD.n16068 DVDD.n3122 4.5005
R15063 DVDD.n16068 DVDD.n16067 4.5005
R15064 DVDD.n3115 DVDD.n3107 4.5005
R15065 DVDD.n3116 DVDD.n3107 4.5005
R15066 DVDD.n3114 DVDD.n3107 4.5005
R15067 DVDD.n3117 DVDD.n3107 4.5005
R15068 DVDD.n3113 DVDD.n3107 4.5005
R15069 DVDD.n3118 DVDD.n3107 4.5005
R15070 DVDD.n3112 DVDD.n3107 4.5005
R15071 DVDD.n3119 DVDD.n3107 4.5005
R15072 DVDD.n3111 DVDD.n3107 4.5005
R15073 DVDD.n3120 DVDD.n3107 4.5005
R15074 DVDD.n3110 DVDD.n3107 4.5005
R15075 DVDD.n3121 DVDD.n3107 4.5005
R15076 DVDD.n3109 DVDD.n3107 4.5005
R15077 DVDD.n3122 DVDD.n3107 4.5005
R15078 DVDD.n16061 DVDD.n3107 4.5005
R15079 DVDD.n16067 DVDD.n3107 4.5005
R15080 DVDD.n5158 DVDD.n5136 4.5005
R15081 DVDD.n5158 DVDD.n5137 4.5005
R15082 DVDD.n5158 DVDD.n5135 4.5005
R15083 DVDD.n5158 DVDD.n5138 4.5005
R15084 DVDD.n5158 DVDD.n5134 4.5005
R15085 DVDD.n5158 DVDD.n5140 4.5005
R15086 DVDD.n5158 DVDD.n5132 4.5005
R15087 DVDD.n5158 DVDD.n5141 4.5005
R15088 DVDD.n5158 DVDD.n5131 4.5005
R15089 DVDD.n5158 DVDD.n5142 4.5005
R15090 DVDD.n15520 DVDD.n5158 4.5005
R15091 DVDD.n15528 DVDD.n5158 4.5005
R15092 DVDD.n5168 DVDD.n5136 4.5005
R15093 DVDD.n5168 DVDD.n5137 4.5005
R15094 DVDD.n5168 DVDD.n5135 4.5005
R15095 DVDD.n5168 DVDD.n5138 4.5005
R15096 DVDD.n5168 DVDD.n5134 4.5005
R15097 DVDD.n5168 DVDD.n5139 4.5005
R15098 DVDD.n5168 DVDD.n5133 4.5005
R15099 DVDD.n5168 DVDD.n5140 4.5005
R15100 DVDD.n5168 DVDD.n5132 4.5005
R15101 DVDD.n5168 DVDD.n5141 4.5005
R15102 DVDD.n5168 DVDD.n5131 4.5005
R15103 DVDD.n5168 DVDD.n5142 4.5005
R15104 DVDD.n15520 DVDD.n5168 4.5005
R15105 DVDD.n5168 DVDD.n5143 4.5005
R15106 DVDD.n15528 DVDD.n5168 4.5005
R15107 DVDD.n5155 DVDD.n5136 4.5005
R15108 DVDD.n5155 DVDD.n5137 4.5005
R15109 DVDD.n5155 DVDD.n5135 4.5005
R15110 DVDD.n5155 DVDD.n5138 4.5005
R15111 DVDD.n5155 DVDD.n5134 4.5005
R15112 DVDD.n5155 DVDD.n5139 4.5005
R15113 DVDD.n5155 DVDD.n5133 4.5005
R15114 DVDD.n5155 DVDD.n5140 4.5005
R15115 DVDD.n5155 DVDD.n5132 4.5005
R15116 DVDD.n5155 DVDD.n5141 4.5005
R15117 DVDD.n5155 DVDD.n5131 4.5005
R15118 DVDD.n5155 DVDD.n5142 4.5005
R15119 DVDD.n5155 DVDD.n5143 4.5005
R15120 DVDD.n15528 DVDD.n5155 4.5005
R15121 DVDD.n5170 DVDD.n5136 4.5005
R15122 DVDD.n5170 DVDD.n5137 4.5005
R15123 DVDD.n5170 DVDD.n5135 4.5005
R15124 DVDD.n5170 DVDD.n5138 4.5005
R15125 DVDD.n5170 DVDD.n5134 4.5005
R15126 DVDD.n5170 DVDD.n5139 4.5005
R15127 DVDD.n5170 DVDD.n5133 4.5005
R15128 DVDD.n5170 DVDD.n5140 4.5005
R15129 DVDD.n5170 DVDD.n5132 4.5005
R15130 DVDD.n5170 DVDD.n5141 4.5005
R15131 DVDD.n5170 DVDD.n5131 4.5005
R15132 DVDD.n5170 DVDD.n5142 4.5005
R15133 DVDD.n5170 DVDD.n5143 4.5005
R15134 DVDD.n15528 DVDD.n5170 4.5005
R15135 DVDD.n5154 DVDD.n5136 4.5005
R15136 DVDD.n5154 DVDD.n5137 4.5005
R15137 DVDD.n5154 DVDD.n5135 4.5005
R15138 DVDD.n5154 DVDD.n5138 4.5005
R15139 DVDD.n5154 DVDD.n5134 4.5005
R15140 DVDD.n5154 DVDD.n5139 4.5005
R15141 DVDD.n5154 DVDD.n5133 4.5005
R15142 DVDD.n5154 DVDD.n5140 4.5005
R15143 DVDD.n5154 DVDD.n5132 4.5005
R15144 DVDD.n5154 DVDD.n5141 4.5005
R15145 DVDD.n5154 DVDD.n5131 4.5005
R15146 DVDD.n5154 DVDD.n5142 4.5005
R15147 DVDD.n15520 DVDD.n5154 4.5005
R15148 DVDD.n5154 DVDD.n5143 4.5005
R15149 DVDD.n15528 DVDD.n5154 4.5005
R15150 DVDD.n5179 DVDD.n5136 4.5005
R15151 DVDD.n5179 DVDD.n5137 4.5005
R15152 DVDD.n5179 DVDD.n5135 4.5005
R15153 DVDD.n5179 DVDD.n5138 4.5005
R15154 DVDD.n5179 DVDD.n5134 4.5005
R15155 DVDD.n5179 DVDD.n5139 4.5005
R15156 DVDD.n5179 DVDD.n5133 4.5005
R15157 DVDD.n5179 DVDD.n5140 4.5005
R15158 DVDD.n5179 DVDD.n5132 4.5005
R15159 DVDD.n5179 DVDD.n5141 4.5005
R15160 DVDD.n5179 DVDD.n5131 4.5005
R15161 DVDD.n5179 DVDD.n5142 4.5005
R15162 DVDD.n15520 DVDD.n5179 4.5005
R15163 DVDD.n5179 DVDD.n5143 4.5005
R15164 DVDD.n15528 DVDD.n5179 4.5005
R15165 DVDD.n5153 DVDD.n5136 4.5005
R15166 DVDD.n5153 DVDD.n5137 4.5005
R15167 DVDD.n5153 DVDD.n5135 4.5005
R15168 DVDD.n5153 DVDD.n5138 4.5005
R15169 DVDD.n5153 DVDD.n5134 4.5005
R15170 DVDD.n5153 DVDD.n5139 4.5005
R15171 DVDD.n5153 DVDD.n5133 4.5005
R15172 DVDD.n5153 DVDD.n5140 4.5005
R15173 DVDD.n5153 DVDD.n5132 4.5005
R15174 DVDD.n5153 DVDD.n5141 4.5005
R15175 DVDD.n5153 DVDD.n5131 4.5005
R15176 DVDD.n5153 DVDD.n5142 4.5005
R15177 DVDD.n5153 DVDD.n5143 4.5005
R15178 DVDD.n15528 DVDD.n5153 4.5005
R15179 DVDD.n5181 DVDD.n5136 4.5005
R15180 DVDD.n5181 DVDD.n5137 4.5005
R15181 DVDD.n5181 DVDD.n5135 4.5005
R15182 DVDD.n5181 DVDD.n5138 4.5005
R15183 DVDD.n5181 DVDD.n5134 4.5005
R15184 DVDD.n5181 DVDD.n5139 4.5005
R15185 DVDD.n5181 DVDD.n5133 4.5005
R15186 DVDD.n5181 DVDD.n5140 4.5005
R15187 DVDD.n5181 DVDD.n5132 4.5005
R15188 DVDD.n5181 DVDD.n5141 4.5005
R15189 DVDD.n5181 DVDD.n5131 4.5005
R15190 DVDD.n5181 DVDD.n5142 4.5005
R15191 DVDD.n5181 DVDD.n5143 4.5005
R15192 DVDD.n15528 DVDD.n5181 4.5005
R15193 DVDD.n5152 DVDD.n5136 4.5005
R15194 DVDD.n5152 DVDD.n5137 4.5005
R15195 DVDD.n5152 DVDD.n5135 4.5005
R15196 DVDD.n5152 DVDD.n5138 4.5005
R15197 DVDD.n5152 DVDD.n5134 4.5005
R15198 DVDD.n5152 DVDD.n5139 4.5005
R15199 DVDD.n5152 DVDD.n5133 4.5005
R15200 DVDD.n5152 DVDD.n5140 4.5005
R15201 DVDD.n5152 DVDD.n5132 4.5005
R15202 DVDD.n5152 DVDD.n5141 4.5005
R15203 DVDD.n5152 DVDD.n5131 4.5005
R15204 DVDD.n5152 DVDD.n5142 4.5005
R15205 DVDD.n15520 DVDD.n5152 4.5005
R15206 DVDD.n5152 DVDD.n5143 4.5005
R15207 DVDD.n15528 DVDD.n5152 4.5005
R15208 DVDD.n5190 DVDD.n5136 4.5005
R15209 DVDD.n5190 DVDD.n5137 4.5005
R15210 DVDD.n5190 DVDD.n5135 4.5005
R15211 DVDD.n5190 DVDD.n5138 4.5005
R15212 DVDD.n5190 DVDD.n5134 4.5005
R15213 DVDD.n5190 DVDD.n5139 4.5005
R15214 DVDD.n5190 DVDD.n5133 4.5005
R15215 DVDD.n5190 DVDD.n5140 4.5005
R15216 DVDD.n5190 DVDD.n5132 4.5005
R15217 DVDD.n5190 DVDD.n5141 4.5005
R15218 DVDD.n5190 DVDD.n5131 4.5005
R15219 DVDD.n5190 DVDD.n5142 4.5005
R15220 DVDD.n15520 DVDD.n5190 4.5005
R15221 DVDD.n5190 DVDD.n5143 4.5005
R15222 DVDD.n15528 DVDD.n5190 4.5005
R15223 DVDD.n5151 DVDD.n5136 4.5005
R15224 DVDD.n5151 DVDD.n5137 4.5005
R15225 DVDD.n5151 DVDD.n5135 4.5005
R15226 DVDD.n5151 DVDD.n5138 4.5005
R15227 DVDD.n5151 DVDD.n5134 4.5005
R15228 DVDD.n5151 DVDD.n5139 4.5005
R15229 DVDD.n5151 DVDD.n5133 4.5005
R15230 DVDD.n5151 DVDD.n5140 4.5005
R15231 DVDD.n5151 DVDD.n5132 4.5005
R15232 DVDD.n5151 DVDD.n5141 4.5005
R15233 DVDD.n5151 DVDD.n5131 4.5005
R15234 DVDD.n5151 DVDD.n5142 4.5005
R15235 DVDD.n5151 DVDD.n5143 4.5005
R15236 DVDD.n15528 DVDD.n5151 4.5005
R15237 DVDD.n5192 DVDD.n5136 4.5005
R15238 DVDD.n5192 DVDD.n5137 4.5005
R15239 DVDD.n5192 DVDD.n5135 4.5005
R15240 DVDD.n5192 DVDD.n5138 4.5005
R15241 DVDD.n5192 DVDD.n5134 4.5005
R15242 DVDD.n5192 DVDD.n5139 4.5005
R15243 DVDD.n5192 DVDD.n5133 4.5005
R15244 DVDD.n5192 DVDD.n5140 4.5005
R15245 DVDD.n5192 DVDD.n5132 4.5005
R15246 DVDD.n5192 DVDD.n5141 4.5005
R15247 DVDD.n5192 DVDD.n5131 4.5005
R15248 DVDD.n5192 DVDD.n5142 4.5005
R15249 DVDD.n5192 DVDD.n5143 4.5005
R15250 DVDD.n15528 DVDD.n5192 4.5005
R15251 DVDD.n5150 DVDD.n5136 4.5005
R15252 DVDD.n5150 DVDD.n5137 4.5005
R15253 DVDD.n5150 DVDD.n5135 4.5005
R15254 DVDD.n5150 DVDD.n5138 4.5005
R15255 DVDD.n5150 DVDD.n5134 4.5005
R15256 DVDD.n5150 DVDD.n5139 4.5005
R15257 DVDD.n5150 DVDD.n5133 4.5005
R15258 DVDD.n5150 DVDD.n5140 4.5005
R15259 DVDD.n5150 DVDD.n5132 4.5005
R15260 DVDD.n5150 DVDD.n5141 4.5005
R15261 DVDD.n5150 DVDD.n5131 4.5005
R15262 DVDD.n5150 DVDD.n5142 4.5005
R15263 DVDD.n15520 DVDD.n5150 4.5005
R15264 DVDD.n5150 DVDD.n5143 4.5005
R15265 DVDD.n15528 DVDD.n5150 4.5005
R15266 DVDD.n5200 DVDD.n5136 4.5005
R15267 DVDD.n5200 DVDD.n5137 4.5005
R15268 DVDD.n5200 DVDD.n5135 4.5005
R15269 DVDD.n5200 DVDD.n5138 4.5005
R15270 DVDD.n5200 DVDD.n5134 4.5005
R15271 DVDD.n5200 DVDD.n5139 4.5005
R15272 DVDD.n5200 DVDD.n5133 4.5005
R15273 DVDD.n5200 DVDD.n5140 4.5005
R15274 DVDD.n5200 DVDD.n5132 4.5005
R15275 DVDD.n5200 DVDD.n5141 4.5005
R15276 DVDD.n5200 DVDD.n5131 4.5005
R15277 DVDD.n5200 DVDD.n5142 4.5005
R15278 DVDD.n15520 DVDD.n5200 4.5005
R15279 DVDD.n5200 DVDD.n5143 4.5005
R15280 DVDD.n15528 DVDD.n5200 4.5005
R15281 DVDD.n5149 DVDD.n5136 4.5005
R15282 DVDD.n5149 DVDD.n5137 4.5005
R15283 DVDD.n5149 DVDD.n5135 4.5005
R15284 DVDD.n5149 DVDD.n5138 4.5005
R15285 DVDD.n5149 DVDD.n5134 4.5005
R15286 DVDD.n5149 DVDD.n5139 4.5005
R15287 DVDD.n5149 DVDD.n5133 4.5005
R15288 DVDD.n5149 DVDD.n5140 4.5005
R15289 DVDD.n5149 DVDD.n5132 4.5005
R15290 DVDD.n5149 DVDD.n5141 4.5005
R15291 DVDD.n5149 DVDD.n5131 4.5005
R15292 DVDD.n5149 DVDD.n5142 4.5005
R15293 DVDD.n5149 DVDD.n5143 4.5005
R15294 DVDD.n15528 DVDD.n5149 4.5005
R15295 DVDD.n5202 DVDD.n5136 4.5005
R15296 DVDD.n5202 DVDD.n5137 4.5005
R15297 DVDD.n5202 DVDD.n5135 4.5005
R15298 DVDD.n5202 DVDD.n5138 4.5005
R15299 DVDD.n5202 DVDD.n5134 4.5005
R15300 DVDD.n5202 DVDD.n5139 4.5005
R15301 DVDD.n5202 DVDD.n5133 4.5005
R15302 DVDD.n5202 DVDD.n5140 4.5005
R15303 DVDD.n5202 DVDD.n5132 4.5005
R15304 DVDD.n5202 DVDD.n5141 4.5005
R15305 DVDD.n5202 DVDD.n5131 4.5005
R15306 DVDD.n5202 DVDD.n5142 4.5005
R15307 DVDD.n5202 DVDD.n5143 4.5005
R15308 DVDD.n15528 DVDD.n5202 4.5005
R15309 DVDD.n5148 DVDD.n5136 4.5005
R15310 DVDD.n5148 DVDD.n5137 4.5005
R15311 DVDD.n5148 DVDD.n5135 4.5005
R15312 DVDD.n5148 DVDD.n5138 4.5005
R15313 DVDD.n5148 DVDD.n5134 4.5005
R15314 DVDD.n5148 DVDD.n5139 4.5005
R15315 DVDD.n5148 DVDD.n5133 4.5005
R15316 DVDD.n5148 DVDD.n5140 4.5005
R15317 DVDD.n5148 DVDD.n5132 4.5005
R15318 DVDD.n5148 DVDD.n5141 4.5005
R15319 DVDD.n5148 DVDD.n5131 4.5005
R15320 DVDD.n5148 DVDD.n5142 4.5005
R15321 DVDD.n5148 DVDD.n5143 4.5005
R15322 DVDD.n15528 DVDD.n5148 4.5005
R15323 DVDD.n5204 DVDD.n5136 4.5005
R15324 DVDD.n5204 DVDD.n5137 4.5005
R15325 DVDD.n5204 DVDD.n5135 4.5005
R15326 DVDD.n5204 DVDD.n5138 4.5005
R15327 DVDD.n5204 DVDD.n5134 4.5005
R15328 DVDD.n5204 DVDD.n5139 4.5005
R15329 DVDD.n5204 DVDD.n5133 4.5005
R15330 DVDD.n5204 DVDD.n5140 4.5005
R15331 DVDD.n5204 DVDD.n5132 4.5005
R15332 DVDD.n5204 DVDD.n5141 4.5005
R15333 DVDD.n5204 DVDD.n5131 4.5005
R15334 DVDD.n5204 DVDD.n5142 4.5005
R15335 DVDD.n5204 DVDD.n5143 4.5005
R15336 DVDD.n15528 DVDD.n5204 4.5005
R15337 DVDD.n5147 DVDD.n5136 4.5005
R15338 DVDD.n5147 DVDD.n5137 4.5005
R15339 DVDD.n5147 DVDD.n5135 4.5005
R15340 DVDD.n5147 DVDD.n5138 4.5005
R15341 DVDD.n5147 DVDD.n5134 4.5005
R15342 DVDD.n5147 DVDD.n5139 4.5005
R15343 DVDD.n5147 DVDD.n5133 4.5005
R15344 DVDD.n5147 DVDD.n5140 4.5005
R15345 DVDD.n5147 DVDD.n5132 4.5005
R15346 DVDD.n5147 DVDD.n5141 4.5005
R15347 DVDD.n5147 DVDD.n5131 4.5005
R15348 DVDD.n5147 DVDD.n5142 4.5005
R15349 DVDD.n5147 DVDD.n5143 4.5005
R15350 DVDD.n15528 DVDD.n5147 4.5005
R15351 DVDD.n5206 DVDD.n5136 4.5005
R15352 DVDD.n5206 DVDD.n5137 4.5005
R15353 DVDD.n5206 DVDD.n5135 4.5005
R15354 DVDD.n5206 DVDD.n5138 4.5005
R15355 DVDD.n5206 DVDD.n5134 4.5005
R15356 DVDD.n5206 DVDD.n5139 4.5005
R15357 DVDD.n5206 DVDD.n5133 4.5005
R15358 DVDD.n5206 DVDD.n5140 4.5005
R15359 DVDD.n5206 DVDD.n5132 4.5005
R15360 DVDD.n5206 DVDD.n5141 4.5005
R15361 DVDD.n5206 DVDD.n5131 4.5005
R15362 DVDD.n5206 DVDD.n5142 4.5005
R15363 DVDD.n5206 DVDD.n5143 4.5005
R15364 DVDD.n15528 DVDD.n5206 4.5005
R15365 DVDD.n5146 DVDD.n5136 4.5005
R15366 DVDD.n5146 DVDD.n5137 4.5005
R15367 DVDD.n5146 DVDD.n5135 4.5005
R15368 DVDD.n5146 DVDD.n5138 4.5005
R15369 DVDD.n5146 DVDD.n5134 4.5005
R15370 DVDD.n5146 DVDD.n5139 4.5005
R15371 DVDD.n5146 DVDD.n5133 4.5005
R15372 DVDD.n5146 DVDD.n5140 4.5005
R15373 DVDD.n5146 DVDD.n5132 4.5005
R15374 DVDD.n5146 DVDD.n5141 4.5005
R15375 DVDD.n5146 DVDD.n5131 4.5005
R15376 DVDD.n5146 DVDD.n5142 4.5005
R15377 DVDD.n15520 DVDD.n5146 4.5005
R15378 DVDD.n5146 DVDD.n5143 4.5005
R15379 DVDD.n15528 DVDD.n5146 4.5005
R15380 DVDD.n15527 DVDD.n5136 4.5005
R15381 DVDD.n15527 DVDD.n5137 4.5005
R15382 DVDD.n15527 DVDD.n5135 4.5005
R15383 DVDD.n15527 DVDD.n5138 4.5005
R15384 DVDD.n15527 DVDD.n5134 4.5005
R15385 DVDD.n15527 DVDD.n5139 4.5005
R15386 DVDD.n15527 DVDD.n5133 4.5005
R15387 DVDD.n15527 DVDD.n5140 4.5005
R15388 DVDD.n15527 DVDD.n5132 4.5005
R15389 DVDD.n15527 DVDD.n5141 4.5005
R15390 DVDD.n15527 DVDD.n5131 4.5005
R15391 DVDD.n15527 DVDD.n5142 4.5005
R15392 DVDD.n15527 DVDD.n15520 4.5005
R15393 DVDD.n15527 DVDD.n5143 4.5005
R15394 DVDD.n15528 DVDD.n15527 4.5005
R15395 DVDD.n5145 DVDD.n5136 4.5005
R15396 DVDD.n5145 DVDD.n5137 4.5005
R15397 DVDD.n5145 DVDD.n5135 4.5005
R15398 DVDD.n5145 DVDD.n5138 4.5005
R15399 DVDD.n5145 DVDD.n5134 4.5005
R15400 DVDD.n5145 DVDD.n5139 4.5005
R15401 DVDD.n5145 DVDD.n5133 4.5005
R15402 DVDD.n5145 DVDD.n5140 4.5005
R15403 DVDD.n5145 DVDD.n5132 4.5005
R15404 DVDD.n5145 DVDD.n5141 4.5005
R15405 DVDD.n5145 DVDD.n5131 4.5005
R15406 DVDD.n5145 DVDD.n5142 4.5005
R15407 DVDD.n5145 DVDD.n5143 4.5005
R15408 DVDD.n15528 DVDD.n5145 4.5005
R15409 DVDD.n15529 DVDD.n5136 4.5005
R15410 DVDD.n15529 DVDD.n5137 4.5005
R15411 DVDD.n15529 DVDD.n5135 4.5005
R15412 DVDD.n15529 DVDD.n5138 4.5005
R15413 DVDD.n15529 DVDD.n5134 4.5005
R15414 DVDD.n15529 DVDD.n5139 4.5005
R15415 DVDD.n15529 DVDD.n5133 4.5005
R15416 DVDD.n15529 DVDD.n5140 4.5005
R15417 DVDD.n15529 DVDD.n5132 4.5005
R15418 DVDD.n15529 DVDD.n5141 4.5005
R15419 DVDD.n15529 DVDD.n5131 4.5005
R15420 DVDD.n15529 DVDD.n5142 4.5005
R15421 DVDD.n15529 DVDD.n5143 4.5005
R15422 DVDD.n15529 DVDD.n5129 4.5005
R15423 DVDD.n15529 DVDD.n15528 4.5005
R15424 DVDD.n15680 DVDD.n15534 4.5005
R15425 DVDD.n15610 DVDD.n15534 4.5005
R15426 DVDD.n15605 DVDD.n15534 4.5005
R15427 DVDD.n15611 DVDD.n15534 4.5005
R15428 DVDD.n15604 DVDD.n15534 4.5005
R15429 DVDD.n15614 DVDD.n15534 4.5005
R15430 DVDD.n15602 DVDD.n15534 4.5005
R15431 DVDD.n15615 DVDD.n15534 4.5005
R15432 DVDD.n15601 DVDD.n15534 4.5005
R15433 DVDD.n15616 DVDD.n15534 4.5005
R15434 DVDD.n15600 DVDD.n15534 4.5005
R15435 DVDD.n15618 DVDD.n15534 4.5005
R15436 DVDD.n15678 DVDD.n15534 4.5005
R15437 DVDD.n15680 DVDD.n15536 4.5005
R15438 DVDD.n15610 DVDD.n15536 4.5005
R15439 DVDD.n15605 DVDD.n15536 4.5005
R15440 DVDD.n15611 DVDD.n15536 4.5005
R15441 DVDD.n15604 DVDD.n15536 4.5005
R15442 DVDD.n15613 DVDD.n15536 4.5005
R15443 DVDD.n15603 DVDD.n15536 4.5005
R15444 DVDD.n15614 DVDD.n15536 4.5005
R15445 DVDD.n15602 DVDD.n15536 4.5005
R15446 DVDD.n15615 DVDD.n15536 4.5005
R15447 DVDD.n15601 DVDD.n15536 4.5005
R15448 DVDD.n15616 DVDD.n15536 4.5005
R15449 DVDD.n15618 DVDD.n15536 4.5005
R15450 DVDD.n15678 DVDD.n15536 4.5005
R15451 DVDD.n15680 DVDD.n5128 4.5005
R15452 DVDD.n15610 DVDD.n5128 4.5005
R15453 DVDD.n15605 DVDD.n5128 4.5005
R15454 DVDD.n15611 DVDD.n5128 4.5005
R15455 DVDD.n15604 DVDD.n5128 4.5005
R15456 DVDD.n15613 DVDD.n5128 4.5005
R15457 DVDD.n15603 DVDD.n5128 4.5005
R15458 DVDD.n15614 DVDD.n5128 4.5005
R15459 DVDD.n15602 DVDD.n5128 4.5005
R15460 DVDD.n15615 DVDD.n5128 4.5005
R15461 DVDD.n15601 DVDD.n5128 4.5005
R15462 DVDD.n15616 DVDD.n5128 4.5005
R15463 DVDD.n15678 DVDD.n5128 4.5005
R15464 DVDD.n15680 DVDD.n15544 4.5005
R15465 DVDD.n15610 DVDD.n15544 4.5005
R15466 DVDD.n15605 DVDD.n15544 4.5005
R15467 DVDD.n15611 DVDD.n15544 4.5005
R15468 DVDD.n15604 DVDD.n15544 4.5005
R15469 DVDD.n15613 DVDD.n15544 4.5005
R15470 DVDD.n15603 DVDD.n15544 4.5005
R15471 DVDD.n15614 DVDD.n15544 4.5005
R15472 DVDD.n15602 DVDD.n15544 4.5005
R15473 DVDD.n15615 DVDD.n15544 4.5005
R15474 DVDD.n15601 DVDD.n15544 4.5005
R15475 DVDD.n15616 DVDD.n15544 4.5005
R15476 DVDD.n15600 DVDD.n15544 4.5005
R15477 DVDD.n15618 DVDD.n15544 4.5005
R15478 DVDD.n15678 DVDD.n15544 4.5005
R15479 DVDD.n15680 DVDD.n5127 4.5005
R15480 DVDD.n15610 DVDD.n5127 4.5005
R15481 DVDD.n15605 DVDD.n5127 4.5005
R15482 DVDD.n15611 DVDD.n5127 4.5005
R15483 DVDD.n15604 DVDD.n5127 4.5005
R15484 DVDD.n15613 DVDD.n5127 4.5005
R15485 DVDD.n15603 DVDD.n5127 4.5005
R15486 DVDD.n15614 DVDD.n5127 4.5005
R15487 DVDD.n15602 DVDD.n5127 4.5005
R15488 DVDD.n15615 DVDD.n5127 4.5005
R15489 DVDD.n15601 DVDD.n5127 4.5005
R15490 DVDD.n15616 DVDD.n5127 4.5005
R15491 DVDD.n15618 DVDD.n5127 4.5005
R15492 DVDD.n15678 DVDD.n5127 4.5005
R15493 DVDD.n15680 DVDD.n15545 4.5005
R15494 DVDD.n15610 DVDD.n15545 4.5005
R15495 DVDD.n15605 DVDD.n15545 4.5005
R15496 DVDD.n15611 DVDD.n15545 4.5005
R15497 DVDD.n15604 DVDD.n15545 4.5005
R15498 DVDD.n15613 DVDD.n15545 4.5005
R15499 DVDD.n15603 DVDD.n15545 4.5005
R15500 DVDD.n15614 DVDD.n15545 4.5005
R15501 DVDD.n15602 DVDD.n15545 4.5005
R15502 DVDD.n15615 DVDD.n15545 4.5005
R15503 DVDD.n15601 DVDD.n15545 4.5005
R15504 DVDD.n15616 DVDD.n15545 4.5005
R15505 DVDD.n15618 DVDD.n15545 4.5005
R15506 DVDD.n15678 DVDD.n15545 4.5005
R15507 DVDD.n15680 DVDD.n5126 4.5005
R15508 DVDD.n15610 DVDD.n5126 4.5005
R15509 DVDD.n15605 DVDD.n5126 4.5005
R15510 DVDD.n15611 DVDD.n5126 4.5005
R15511 DVDD.n15604 DVDD.n5126 4.5005
R15512 DVDD.n15613 DVDD.n5126 4.5005
R15513 DVDD.n15603 DVDD.n5126 4.5005
R15514 DVDD.n15614 DVDD.n5126 4.5005
R15515 DVDD.n15602 DVDD.n5126 4.5005
R15516 DVDD.n15615 DVDD.n5126 4.5005
R15517 DVDD.n15601 DVDD.n5126 4.5005
R15518 DVDD.n15616 DVDD.n5126 4.5005
R15519 DVDD.n15600 DVDD.n5126 4.5005
R15520 DVDD.n15618 DVDD.n5126 4.5005
R15521 DVDD.n15678 DVDD.n5126 4.5005
R15522 DVDD.n15680 DVDD.n15553 4.5005
R15523 DVDD.n15610 DVDD.n15553 4.5005
R15524 DVDD.n15605 DVDD.n15553 4.5005
R15525 DVDD.n15611 DVDD.n15553 4.5005
R15526 DVDD.n15604 DVDD.n15553 4.5005
R15527 DVDD.n15613 DVDD.n15553 4.5005
R15528 DVDD.n15603 DVDD.n15553 4.5005
R15529 DVDD.n15614 DVDD.n15553 4.5005
R15530 DVDD.n15602 DVDD.n15553 4.5005
R15531 DVDD.n15615 DVDD.n15553 4.5005
R15532 DVDD.n15601 DVDD.n15553 4.5005
R15533 DVDD.n15616 DVDD.n15553 4.5005
R15534 DVDD.n15600 DVDD.n15553 4.5005
R15535 DVDD.n15618 DVDD.n15553 4.5005
R15536 DVDD.n15678 DVDD.n15553 4.5005
R15537 DVDD.n15680 DVDD.n5125 4.5005
R15538 DVDD.n15610 DVDD.n5125 4.5005
R15539 DVDD.n15605 DVDD.n5125 4.5005
R15540 DVDD.n15611 DVDD.n5125 4.5005
R15541 DVDD.n15604 DVDD.n5125 4.5005
R15542 DVDD.n15613 DVDD.n5125 4.5005
R15543 DVDD.n15603 DVDD.n5125 4.5005
R15544 DVDD.n15614 DVDD.n5125 4.5005
R15545 DVDD.n15602 DVDD.n5125 4.5005
R15546 DVDD.n15615 DVDD.n5125 4.5005
R15547 DVDD.n15601 DVDD.n5125 4.5005
R15548 DVDD.n15616 DVDD.n5125 4.5005
R15549 DVDD.n15618 DVDD.n5125 4.5005
R15550 DVDD.n15678 DVDD.n5125 4.5005
R15551 DVDD.n15680 DVDD.n15554 4.5005
R15552 DVDD.n15610 DVDD.n15554 4.5005
R15553 DVDD.n15605 DVDD.n15554 4.5005
R15554 DVDD.n15611 DVDD.n15554 4.5005
R15555 DVDD.n15604 DVDD.n15554 4.5005
R15556 DVDD.n15613 DVDD.n15554 4.5005
R15557 DVDD.n15603 DVDD.n15554 4.5005
R15558 DVDD.n15614 DVDD.n15554 4.5005
R15559 DVDD.n15602 DVDD.n15554 4.5005
R15560 DVDD.n15615 DVDD.n15554 4.5005
R15561 DVDD.n15601 DVDD.n15554 4.5005
R15562 DVDD.n15616 DVDD.n15554 4.5005
R15563 DVDD.n15618 DVDD.n15554 4.5005
R15564 DVDD.n15678 DVDD.n15554 4.5005
R15565 DVDD.n15680 DVDD.n5124 4.5005
R15566 DVDD.n15610 DVDD.n5124 4.5005
R15567 DVDD.n15605 DVDD.n5124 4.5005
R15568 DVDD.n15611 DVDD.n5124 4.5005
R15569 DVDD.n15604 DVDD.n5124 4.5005
R15570 DVDD.n15613 DVDD.n5124 4.5005
R15571 DVDD.n15603 DVDD.n5124 4.5005
R15572 DVDD.n15614 DVDD.n5124 4.5005
R15573 DVDD.n15602 DVDD.n5124 4.5005
R15574 DVDD.n15615 DVDD.n5124 4.5005
R15575 DVDD.n15601 DVDD.n5124 4.5005
R15576 DVDD.n15616 DVDD.n5124 4.5005
R15577 DVDD.n15600 DVDD.n5124 4.5005
R15578 DVDD.n15618 DVDD.n5124 4.5005
R15579 DVDD.n15678 DVDD.n5124 4.5005
R15580 DVDD.n15680 DVDD.n15562 4.5005
R15581 DVDD.n15610 DVDD.n15562 4.5005
R15582 DVDD.n15605 DVDD.n15562 4.5005
R15583 DVDD.n15611 DVDD.n15562 4.5005
R15584 DVDD.n15604 DVDD.n15562 4.5005
R15585 DVDD.n15613 DVDD.n15562 4.5005
R15586 DVDD.n15603 DVDD.n15562 4.5005
R15587 DVDD.n15614 DVDD.n15562 4.5005
R15588 DVDD.n15602 DVDD.n15562 4.5005
R15589 DVDD.n15615 DVDD.n15562 4.5005
R15590 DVDD.n15601 DVDD.n15562 4.5005
R15591 DVDD.n15616 DVDD.n15562 4.5005
R15592 DVDD.n15600 DVDD.n15562 4.5005
R15593 DVDD.n15618 DVDD.n15562 4.5005
R15594 DVDD.n15678 DVDD.n15562 4.5005
R15595 DVDD.n15680 DVDD.n5123 4.5005
R15596 DVDD.n15610 DVDD.n5123 4.5005
R15597 DVDD.n15605 DVDD.n5123 4.5005
R15598 DVDD.n15611 DVDD.n5123 4.5005
R15599 DVDD.n15604 DVDD.n5123 4.5005
R15600 DVDD.n15613 DVDD.n5123 4.5005
R15601 DVDD.n15603 DVDD.n5123 4.5005
R15602 DVDD.n15614 DVDD.n5123 4.5005
R15603 DVDD.n15602 DVDD.n5123 4.5005
R15604 DVDD.n15615 DVDD.n5123 4.5005
R15605 DVDD.n15601 DVDD.n5123 4.5005
R15606 DVDD.n15616 DVDD.n5123 4.5005
R15607 DVDD.n15618 DVDD.n5123 4.5005
R15608 DVDD.n15678 DVDD.n5123 4.5005
R15609 DVDD.n15680 DVDD.n15563 4.5005
R15610 DVDD.n15610 DVDD.n15563 4.5005
R15611 DVDD.n15605 DVDD.n15563 4.5005
R15612 DVDD.n15611 DVDD.n15563 4.5005
R15613 DVDD.n15604 DVDD.n15563 4.5005
R15614 DVDD.n15613 DVDD.n15563 4.5005
R15615 DVDD.n15603 DVDD.n15563 4.5005
R15616 DVDD.n15614 DVDD.n15563 4.5005
R15617 DVDD.n15602 DVDD.n15563 4.5005
R15618 DVDD.n15615 DVDD.n15563 4.5005
R15619 DVDD.n15601 DVDD.n15563 4.5005
R15620 DVDD.n15616 DVDD.n15563 4.5005
R15621 DVDD.n15618 DVDD.n15563 4.5005
R15622 DVDD.n15678 DVDD.n15563 4.5005
R15623 DVDD.n15680 DVDD.n5122 4.5005
R15624 DVDD.n15610 DVDD.n5122 4.5005
R15625 DVDD.n15605 DVDD.n5122 4.5005
R15626 DVDD.n15611 DVDD.n5122 4.5005
R15627 DVDD.n15604 DVDD.n5122 4.5005
R15628 DVDD.n15613 DVDD.n5122 4.5005
R15629 DVDD.n15603 DVDD.n5122 4.5005
R15630 DVDD.n15614 DVDD.n5122 4.5005
R15631 DVDD.n15602 DVDD.n5122 4.5005
R15632 DVDD.n15615 DVDD.n5122 4.5005
R15633 DVDD.n15601 DVDD.n5122 4.5005
R15634 DVDD.n15616 DVDD.n5122 4.5005
R15635 DVDD.n15600 DVDD.n5122 4.5005
R15636 DVDD.n15618 DVDD.n5122 4.5005
R15637 DVDD.n15678 DVDD.n5122 4.5005
R15638 DVDD.n15680 DVDD.n15571 4.5005
R15639 DVDD.n15610 DVDD.n15571 4.5005
R15640 DVDD.n15605 DVDD.n15571 4.5005
R15641 DVDD.n15611 DVDD.n15571 4.5005
R15642 DVDD.n15604 DVDD.n15571 4.5005
R15643 DVDD.n15613 DVDD.n15571 4.5005
R15644 DVDD.n15603 DVDD.n15571 4.5005
R15645 DVDD.n15614 DVDD.n15571 4.5005
R15646 DVDD.n15602 DVDD.n15571 4.5005
R15647 DVDD.n15615 DVDD.n15571 4.5005
R15648 DVDD.n15601 DVDD.n15571 4.5005
R15649 DVDD.n15616 DVDD.n15571 4.5005
R15650 DVDD.n15600 DVDD.n15571 4.5005
R15651 DVDD.n15618 DVDD.n15571 4.5005
R15652 DVDD.n15678 DVDD.n15571 4.5005
R15653 DVDD.n15680 DVDD.n5121 4.5005
R15654 DVDD.n15610 DVDD.n5121 4.5005
R15655 DVDD.n15605 DVDD.n5121 4.5005
R15656 DVDD.n15611 DVDD.n5121 4.5005
R15657 DVDD.n15604 DVDD.n5121 4.5005
R15658 DVDD.n15613 DVDD.n5121 4.5005
R15659 DVDD.n15603 DVDD.n5121 4.5005
R15660 DVDD.n15614 DVDD.n5121 4.5005
R15661 DVDD.n15602 DVDD.n5121 4.5005
R15662 DVDD.n15615 DVDD.n5121 4.5005
R15663 DVDD.n15601 DVDD.n5121 4.5005
R15664 DVDD.n15616 DVDD.n5121 4.5005
R15665 DVDD.n15618 DVDD.n5121 4.5005
R15666 DVDD.n15678 DVDD.n5121 4.5005
R15667 DVDD.n15680 DVDD.n15572 4.5005
R15668 DVDD.n15610 DVDD.n15572 4.5005
R15669 DVDD.n15605 DVDD.n15572 4.5005
R15670 DVDD.n15611 DVDD.n15572 4.5005
R15671 DVDD.n15604 DVDD.n15572 4.5005
R15672 DVDD.n15613 DVDD.n15572 4.5005
R15673 DVDD.n15603 DVDD.n15572 4.5005
R15674 DVDD.n15614 DVDD.n15572 4.5005
R15675 DVDD.n15602 DVDD.n15572 4.5005
R15676 DVDD.n15615 DVDD.n15572 4.5005
R15677 DVDD.n15601 DVDD.n15572 4.5005
R15678 DVDD.n15616 DVDD.n15572 4.5005
R15679 DVDD.n15618 DVDD.n15572 4.5005
R15680 DVDD.n15678 DVDD.n15572 4.5005
R15681 DVDD.n15680 DVDD.n5120 4.5005
R15682 DVDD.n15610 DVDD.n5120 4.5005
R15683 DVDD.n15605 DVDD.n5120 4.5005
R15684 DVDD.n15611 DVDD.n5120 4.5005
R15685 DVDD.n15604 DVDD.n5120 4.5005
R15686 DVDD.n15613 DVDD.n5120 4.5005
R15687 DVDD.n15603 DVDD.n5120 4.5005
R15688 DVDD.n15614 DVDD.n5120 4.5005
R15689 DVDD.n15602 DVDD.n5120 4.5005
R15690 DVDD.n15615 DVDD.n5120 4.5005
R15691 DVDD.n15601 DVDD.n5120 4.5005
R15692 DVDD.n15616 DVDD.n5120 4.5005
R15693 DVDD.n15600 DVDD.n5120 4.5005
R15694 DVDD.n15618 DVDD.n5120 4.5005
R15695 DVDD.n15678 DVDD.n5120 4.5005
R15696 DVDD.n15680 DVDD.n15580 4.5005
R15697 DVDD.n15610 DVDD.n15580 4.5005
R15698 DVDD.n15605 DVDD.n15580 4.5005
R15699 DVDD.n15611 DVDD.n15580 4.5005
R15700 DVDD.n15604 DVDD.n15580 4.5005
R15701 DVDD.n15613 DVDD.n15580 4.5005
R15702 DVDD.n15603 DVDD.n15580 4.5005
R15703 DVDD.n15614 DVDD.n15580 4.5005
R15704 DVDD.n15602 DVDD.n15580 4.5005
R15705 DVDD.n15615 DVDD.n15580 4.5005
R15706 DVDD.n15601 DVDD.n15580 4.5005
R15707 DVDD.n15616 DVDD.n15580 4.5005
R15708 DVDD.n15600 DVDD.n15580 4.5005
R15709 DVDD.n15618 DVDD.n15580 4.5005
R15710 DVDD.n15678 DVDD.n15580 4.5005
R15711 DVDD.n15680 DVDD.n5119 4.5005
R15712 DVDD.n15610 DVDD.n5119 4.5005
R15713 DVDD.n15605 DVDD.n5119 4.5005
R15714 DVDD.n15611 DVDD.n5119 4.5005
R15715 DVDD.n15604 DVDD.n5119 4.5005
R15716 DVDD.n15613 DVDD.n5119 4.5005
R15717 DVDD.n15603 DVDD.n5119 4.5005
R15718 DVDD.n15614 DVDD.n5119 4.5005
R15719 DVDD.n15602 DVDD.n5119 4.5005
R15720 DVDD.n15615 DVDD.n5119 4.5005
R15721 DVDD.n15601 DVDD.n5119 4.5005
R15722 DVDD.n15616 DVDD.n5119 4.5005
R15723 DVDD.n15618 DVDD.n5119 4.5005
R15724 DVDD.n15678 DVDD.n5119 4.5005
R15725 DVDD.n15680 DVDD.n15581 4.5005
R15726 DVDD.n15610 DVDD.n15581 4.5005
R15727 DVDD.n15605 DVDD.n15581 4.5005
R15728 DVDD.n15611 DVDD.n15581 4.5005
R15729 DVDD.n15604 DVDD.n15581 4.5005
R15730 DVDD.n15613 DVDD.n15581 4.5005
R15731 DVDD.n15603 DVDD.n15581 4.5005
R15732 DVDD.n15614 DVDD.n15581 4.5005
R15733 DVDD.n15602 DVDD.n15581 4.5005
R15734 DVDD.n15615 DVDD.n15581 4.5005
R15735 DVDD.n15601 DVDD.n15581 4.5005
R15736 DVDD.n15616 DVDD.n15581 4.5005
R15737 DVDD.n15618 DVDD.n15581 4.5005
R15738 DVDD.n15678 DVDD.n15581 4.5005
R15739 DVDD.n15680 DVDD.n5118 4.5005
R15740 DVDD.n15610 DVDD.n5118 4.5005
R15741 DVDD.n15605 DVDD.n5118 4.5005
R15742 DVDD.n15611 DVDD.n5118 4.5005
R15743 DVDD.n15604 DVDD.n5118 4.5005
R15744 DVDD.n15613 DVDD.n5118 4.5005
R15745 DVDD.n15603 DVDD.n5118 4.5005
R15746 DVDD.n15614 DVDD.n5118 4.5005
R15747 DVDD.n15602 DVDD.n5118 4.5005
R15748 DVDD.n15615 DVDD.n5118 4.5005
R15749 DVDD.n15601 DVDD.n5118 4.5005
R15750 DVDD.n15616 DVDD.n5118 4.5005
R15751 DVDD.n15600 DVDD.n5118 4.5005
R15752 DVDD.n15618 DVDD.n5118 4.5005
R15753 DVDD.n15678 DVDD.n5118 4.5005
R15754 DVDD.n15680 DVDD.n15679 4.5005
R15755 DVDD.n15679 DVDD.n15610 4.5005
R15756 DVDD.n15679 DVDD.n15605 4.5005
R15757 DVDD.n15679 DVDD.n15611 4.5005
R15758 DVDD.n15679 DVDD.n15604 4.5005
R15759 DVDD.n15679 DVDD.n15613 4.5005
R15760 DVDD.n15679 DVDD.n15603 4.5005
R15761 DVDD.n15679 DVDD.n15614 4.5005
R15762 DVDD.n15679 DVDD.n15602 4.5005
R15763 DVDD.n15679 DVDD.n15615 4.5005
R15764 DVDD.n15679 DVDD.n15601 4.5005
R15765 DVDD.n15679 DVDD.n15616 4.5005
R15766 DVDD.n15679 DVDD.n15600 4.5005
R15767 DVDD.n15679 DVDD.n15618 4.5005
R15768 DVDD.n15679 DVDD.n15593 4.5005
R15769 DVDD.n15679 DVDD.n15678 4.5005
R15770 DVDD.n3487 DVDD.n3431 4.5005
R15771 DVDD.n3489 DVDD.n3431 4.5005
R15772 DVDD.n3486 DVDD.n3431 4.5005
R15773 DVDD.n3490 DVDD.n3431 4.5005
R15774 DVDD.n3485 DVDD.n3431 4.5005
R15775 DVDD.n3493 DVDD.n3431 4.5005
R15776 DVDD.n3483 DVDD.n3431 4.5005
R15777 DVDD.n3494 DVDD.n3431 4.5005
R15778 DVDD.n3482 DVDD.n3431 4.5005
R15779 DVDD.n15790 DVDD.n3431 4.5005
R15780 DVDD.n3481 DVDD.n3431 4.5005
R15781 DVDD.n15795 DVDD.n3431 4.5005
R15782 DVDD.n3487 DVDD.n3440 4.5005
R15783 DVDD.n3489 DVDD.n3440 4.5005
R15784 DVDD.n3486 DVDD.n3440 4.5005
R15785 DVDD.n3490 DVDD.n3440 4.5005
R15786 DVDD.n3485 DVDD.n3440 4.5005
R15787 DVDD.n3492 DVDD.n3440 4.5005
R15788 DVDD.n3484 DVDD.n3440 4.5005
R15789 DVDD.n3493 DVDD.n3440 4.5005
R15790 DVDD.n3483 DVDD.n3440 4.5005
R15791 DVDD.n3494 DVDD.n3440 4.5005
R15792 DVDD.n3482 DVDD.n3440 4.5005
R15793 DVDD.n15790 DVDD.n3440 4.5005
R15794 DVDD.n3481 DVDD.n3440 4.5005
R15795 DVDD.n15793 DVDD.n3440 4.5005
R15796 DVDD.n15795 DVDD.n3440 4.5005
R15797 DVDD.n3487 DVDD.n3430 4.5005
R15798 DVDD.n3489 DVDD.n3430 4.5005
R15799 DVDD.n3486 DVDD.n3430 4.5005
R15800 DVDD.n3490 DVDD.n3430 4.5005
R15801 DVDD.n3485 DVDD.n3430 4.5005
R15802 DVDD.n3492 DVDD.n3430 4.5005
R15803 DVDD.n3484 DVDD.n3430 4.5005
R15804 DVDD.n3493 DVDD.n3430 4.5005
R15805 DVDD.n3483 DVDD.n3430 4.5005
R15806 DVDD.n3494 DVDD.n3430 4.5005
R15807 DVDD.n3482 DVDD.n3430 4.5005
R15808 DVDD.n15790 DVDD.n3430 4.5005
R15809 DVDD.n15793 DVDD.n3430 4.5005
R15810 DVDD.n15795 DVDD.n3430 4.5005
R15811 DVDD.n3487 DVDD.n3442 4.5005
R15812 DVDD.n3489 DVDD.n3442 4.5005
R15813 DVDD.n3486 DVDD.n3442 4.5005
R15814 DVDD.n3490 DVDD.n3442 4.5005
R15815 DVDD.n3485 DVDD.n3442 4.5005
R15816 DVDD.n3492 DVDD.n3442 4.5005
R15817 DVDD.n3484 DVDD.n3442 4.5005
R15818 DVDD.n3493 DVDD.n3442 4.5005
R15819 DVDD.n3483 DVDD.n3442 4.5005
R15820 DVDD.n3494 DVDD.n3442 4.5005
R15821 DVDD.n3482 DVDD.n3442 4.5005
R15822 DVDD.n15790 DVDD.n3442 4.5005
R15823 DVDD.n15793 DVDD.n3442 4.5005
R15824 DVDD.n15795 DVDD.n3442 4.5005
R15825 DVDD.n3487 DVDD.n3429 4.5005
R15826 DVDD.n3489 DVDD.n3429 4.5005
R15827 DVDD.n3486 DVDD.n3429 4.5005
R15828 DVDD.n3490 DVDD.n3429 4.5005
R15829 DVDD.n3485 DVDD.n3429 4.5005
R15830 DVDD.n3492 DVDD.n3429 4.5005
R15831 DVDD.n3484 DVDD.n3429 4.5005
R15832 DVDD.n3493 DVDD.n3429 4.5005
R15833 DVDD.n3483 DVDD.n3429 4.5005
R15834 DVDD.n3494 DVDD.n3429 4.5005
R15835 DVDD.n3482 DVDD.n3429 4.5005
R15836 DVDD.n15790 DVDD.n3429 4.5005
R15837 DVDD.n3481 DVDD.n3429 4.5005
R15838 DVDD.n15793 DVDD.n3429 4.5005
R15839 DVDD.n15795 DVDD.n3429 4.5005
R15840 DVDD.n3487 DVDD.n3451 4.5005
R15841 DVDD.n3489 DVDD.n3451 4.5005
R15842 DVDD.n3486 DVDD.n3451 4.5005
R15843 DVDD.n3490 DVDD.n3451 4.5005
R15844 DVDD.n3485 DVDD.n3451 4.5005
R15845 DVDD.n3492 DVDD.n3451 4.5005
R15846 DVDD.n3484 DVDD.n3451 4.5005
R15847 DVDD.n3493 DVDD.n3451 4.5005
R15848 DVDD.n3483 DVDD.n3451 4.5005
R15849 DVDD.n3494 DVDD.n3451 4.5005
R15850 DVDD.n3482 DVDD.n3451 4.5005
R15851 DVDD.n15790 DVDD.n3451 4.5005
R15852 DVDD.n3481 DVDD.n3451 4.5005
R15853 DVDD.n15793 DVDD.n3451 4.5005
R15854 DVDD.n15795 DVDD.n3451 4.5005
R15855 DVDD.n3487 DVDD.n3428 4.5005
R15856 DVDD.n3489 DVDD.n3428 4.5005
R15857 DVDD.n3486 DVDD.n3428 4.5005
R15858 DVDD.n3490 DVDD.n3428 4.5005
R15859 DVDD.n3485 DVDD.n3428 4.5005
R15860 DVDD.n3492 DVDD.n3428 4.5005
R15861 DVDD.n3484 DVDD.n3428 4.5005
R15862 DVDD.n3493 DVDD.n3428 4.5005
R15863 DVDD.n3483 DVDD.n3428 4.5005
R15864 DVDD.n3494 DVDD.n3428 4.5005
R15865 DVDD.n3482 DVDD.n3428 4.5005
R15866 DVDD.n15790 DVDD.n3428 4.5005
R15867 DVDD.n15793 DVDD.n3428 4.5005
R15868 DVDD.n15795 DVDD.n3428 4.5005
R15869 DVDD.n3487 DVDD.n3453 4.5005
R15870 DVDD.n3489 DVDD.n3453 4.5005
R15871 DVDD.n3486 DVDD.n3453 4.5005
R15872 DVDD.n3490 DVDD.n3453 4.5005
R15873 DVDD.n3485 DVDD.n3453 4.5005
R15874 DVDD.n3492 DVDD.n3453 4.5005
R15875 DVDD.n3484 DVDD.n3453 4.5005
R15876 DVDD.n3493 DVDD.n3453 4.5005
R15877 DVDD.n3483 DVDD.n3453 4.5005
R15878 DVDD.n3494 DVDD.n3453 4.5005
R15879 DVDD.n3482 DVDD.n3453 4.5005
R15880 DVDD.n15790 DVDD.n3453 4.5005
R15881 DVDD.n15793 DVDD.n3453 4.5005
R15882 DVDD.n15795 DVDD.n3453 4.5005
R15883 DVDD.n3487 DVDD.n3427 4.5005
R15884 DVDD.n3489 DVDD.n3427 4.5005
R15885 DVDD.n3486 DVDD.n3427 4.5005
R15886 DVDD.n3490 DVDD.n3427 4.5005
R15887 DVDD.n3485 DVDD.n3427 4.5005
R15888 DVDD.n3492 DVDD.n3427 4.5005
R15889 DVDD.n3484 DVDD.n3427 4.5005
R15890 DVDD.n3493 DVDD.n3427 4.5005
R15891 DVDD.n3483 DVDD.n3427 4.5005
R15892 DVDD.n3494 DVDD.n3427 4.5005
R15893 DVDD.n3482 DVDD.n3427 4.5005
R15894 DVDD.n15790 DVDD.n3427 4.5005
R15895 DVDD.n3481 DVDD.n3427 4.5005
R15896 DVDD.n15793 DVDD.n3427 4.5005
R15897 DVDD.n15795 DVDD.n3427 4.5005
R15898 DVDD.n3487 DVDD.n3461 4.5005
R15899 DVDD.n3489 DVDD.n3461 4.5005
R15900 DVDD.n3486 DVDD.n3461 4.5005
R15901 DVDD.n3490 DVDD.n3461 4.5005
R15902 DVDD.n3485 DVDD.n3461 4.5005
R15903 DVDD.n3492 DVDD.n3461 4.5005
R15904 DVDD.n3484 DVDD.n3461 4.5005
R15905 DVDD.n3493 DVDD.n3461 4.5005
R15906 DVDD.n3483 DVDD.n3461 4.5005
R15907 DVDD.n3494 DVDD.n3461 4.5005
R15908 DVDD.n3482 DVDD.n3461 4.5005
R15909 DVDD.n15790 DVDD.n3461 4.5005
R15910 DVDD.n3481 DVDD.n3461 4.5005
R15911 DVDD.n15793 DVDD.n3461 4.5005
R15912 DVDD.n15795 DVDD.n3461 4.5005
R15913 DVDD.n3487 DVDD.n3426 4.5005
R15914 DVDD.n3489 DVDD.n3426 4.5005
R15915 DVDD.n3486 DVDD.n3426 4.5005
R15916 DVDD.n3490 DVDD.n3426 4.5005
R15917 DVDD.n3485 DVDD.n3426 4.5005
R15918 DVDD.n3492 DVDD.n3426 4.5005
R15919 DVDD.n3484 DVDD.n3426 4.5005
R15920 DVDD.n3493 DVDD.n3426 4.5005
R15921 DVDD.n3483 DVDD.n3426 4.5005
R15922 DVDD.n3494 DVDD.n3426 4.5005
R15923 DVDD.n3482 DVDD.n3426 4.5005
R15924 DVDD.n15790 DVDD.n3426 4.5005
R15925 DVDD.n15793 DVDD.n3426 4.5005
R15926 DVDD.n15795 DVDD.n3426 4.5005
R15927 DVDD.n3487 DVDD.n3463 4.5005
R15928 DVDD.n3489 DVDD.n3463 4.5005
R15929 DVDD.n3486 DVDD.n3463 4.5005
R15930 DVDD.n3490 DVDD.n3463 4.5005
R15931 DVDD.n3485 DVDD.n3463 4.5005
R15932 DVDD.n3492 DVDD.n3463 4.5005
R15933 DVDD.n3484 DVDD.n3463 4.5005
R15934 DVDD.n3493 DVDD.n3463 4.5005
R15935 DVDD.n3483 DVDD.n3463 4.5005
R15936 DVDD.n3494 DVDD.n3463 4.5005
R15937 DVDD.n3482 DVDD.n3463 4.5005
R15938 DVDD.n15790 DVDD.n3463 4.5005
R15939 DVDD.n15793 DVDD.n3463 4.5005
R15940 DVDD.n15795 DVDD.n3463 4.5005
R15941 DVDD.n3487 DVDD.n3425 4.5005
R15942 DVDD.n3489 DVDD.n3425 4.5005
R15943 DVDD.n3486 DVDD.n3425 4.5005
R15944 DVDD.n3490 DVDD.n3425 4.5005
R15945 DVDD.n3485 DVDD.n3425 4.5005
R15946 DVDD.n3492 DVDD.n3425 4.5005
R15947 DVDD.n3484 DVDD.n3425 4.5005
R15948 DVDD.n3493 DVDD.n3425 4.5005
R15949 DVDD.n3483 DVDD.n3425 4.5005
R15950 DVDD.n3494 DVDD.n3425 4.5005
R15951 DVDD.n3482 DVDD.n3425 4.5005
R15952 DVDD.n15790 DVDD.n3425 4.5005
R15953 DVDD.n15793 DVDD.n3425 4.5005
R15954 DVDD.n15795 DVDD.n3425 4.5005
R15955 DVDD.n3487 DVDD.n3465 4.5005
R15956 DVDD.n3489 DVDD.n3465 4.5005
R15957 DVDD.n3486 DVDD.n3465 4.5005
R15958 DVDD.n3490 DVDD.n3465 4.5005
R15959 DVDD.n3485 DVDD.n3465 4.5005
R15960 DVDD.n3492 DVDD.n3465 4.5005
R15961 DVDD.n3484 DVDD.n3465 4.5005
R15962 DVDD.n3493 DVDD.n3465 4.5005
R15963 DVDD.n3483 DVDD.n3465 4.5005
R15964 DVDD.n3494 DVDD.n3465 4.5005
R15965 DVDD.n3482 DVDD.n3465 4.5005
R15966 DVDD.n15790 DVDD.n3465 4.5005
R15967 DVDD.n15793 DVDD.n3465 4.5005
R15968 DVDD.n15795 DVDD.n3465 4.5005
R15969 DVDD.n3487 DVDD.n3424 4.5005
R15970 DVDD.n3489 DVDD.n3424 4.5005
R15971 DVDD.n3486 DVDD.n3424 4.5005
R15972 DVDD.n3490 DVDD.n3424 4.5005
R15973 DVDD.n3485 DVDD.n3424 4.5005
R15974 DVDD.n3492 DVDD.n3424 4.5005
R15975 DVDD.n3484 DVDD.n3424 4.5005
R15976 DVDD.n3493 DVDD.n3424 4.5005
R15977 DVDD.n3483 DVDD.n3424 4.5005
R15978 DVDD.n3494 DVDD.n3424 4.5005
R15979 DVDD.n3482 DVDD.n3424 4.5005
R15980 DVDD.n15790 DVDD.n3424 4.5005
R15981 DVDD.n15793 DVDD.n3424 4.5005
R15982 DVDD.n15795 DVDD.n3424 4.5005
R15983 DVDD.n3487 DVDD.n3467 4.5005
R15984 DVDD.n3489 DVDD.n3467 4.5005
R15985 DVDD.n3486 DVDD.n3467 4.5005
R15986 DVDD.n3490 DVDD.n3467 4.5005
R15987 DVDD.n3485 DVDD.n3467 4.5005
R15988 DVDD.n3492 DVDD.n3467 4.5005
R15989 DVDD.n3484 DVDD.n3467 4.5005
R15990 DVDD.n3493 DVDD.n3467 4.5005
R15991 DVDD.n3483 DVDD.n3467 4.5005
R15992 DVDD.n3494 DVDD.n3467 4.5005
R15993 DVDD.n3482 DVDD.n3467 4.5005
R15994 DVDD.n15790 DVDD.n3467 4.5005
R15995 DVDD.n15793 DVDD.n3467 4.5005
R15996 DVDD.n15795 DVDD.n3467 4.5005
R15997 DVDD.n3487 DVDD.n3423 4.5005
R15998 DVDD.n3489 DVDD.n3423 4.5005
R15999 DVDD.n3486 DVDD.n3423 4.5005
R16000 DVDD.n3490 DVDD.n3423 4.5005
R16001 DVDD.n3485 DVDD.n3423 4.5005
R16002 DVDD.n3492 DVDD.n3423 4.5005
R16003 DVDD.n3484 DVDD.n3423 4.5005
R16004 DVDD.n3493 DVDD.n3423 4.5005
R16005 DVDD.n3483 DVDD.n3423 4.5005
R16006 DVDD.n3494 DVDD.n3423 4.5005
R16007 DVDD.n3482 DVDD.n3423 4.5005
R16008 DVDD.n15790 DVDD.n3423 4.5005
R16009 DVDD.n3481 DVDD.n3423 4.5005
R16010 DVDD.n15793 DVDD.n3423 4.5005
R16011 DVDD.n15795 DVDD.n3423 4.5005
R16012 DVDD.n3487 DVDD.n3469 4.5005
R16013 DVDD.n3489 DVDD.n3469 4.5005
R16014 DVDD.n3486 DVDD.n3469 4.5005
R16015 DVDD.n3490 DVDD.n3469 4.5005
R16016 DVDD.n3485 DVDD.n3469 4.5005
R16017 DVDD.n3492 DVDD.n3469 4.5005
R16018 DVDD.n3484 DVDD.n3469 4.5005
R16019 DVDD.n3493 DVDD.n3469 4.5005
R16020 DVDD.n3483 DVDD.n3469 4.5005
R16021 DVDD.n3494 DVDD.n3469 4.5005
R16022 DVDD.n3482 DVDD.n3469 4.5005
R16023 DVDD.n15790 DVDD.n3469 4.5005
R16024 DVDD.n15793 DVDD.n3469 4.5005
R16025 DVDD.n15795 DVDD.n3469 4.5005
R16026 DVDD.n3487 DVDD.n3422 4.5005
R16027 DVDD.n3489 DVDD.n3422 4.5005
R16028 DVDD.n3486 DVDD.n3422 4.5005
R16029 DVDD.n3490 DVDD.n3422 4.5005
R16030 DVDD.n3485 DVDD.n3422 4.5005
R16031 DVDD.n3492 DVDD.n3422 4.5005
R16032 DVDD.n3484 DVDD.n3422 4.5005
R16033 DVDD.n3493 DVDD.n3422 4.5005
R16034 DVDD.n3483 DVDD.n3422 4.5005
R16035 DVDD.n3494 DVDD.n3422 4.5005
R16036 DVDD.n3482 DVDD.n3422 4.5005
R16037 DVDD.n15790 DVDD.n3422 4.5005
R16038 DVDD.n15793 DVDD.n3422 4.5005
R16039 DVDD.n15795 DVDD.n3422 4.5005
R16040 DVDD.n3487 DVDD.n3471 4.5005
R16041 DVDD.n3489 DVDD.n3471 4.5005
R16042 DVDD.n3486 DVDD.n3471 4.5005
R16043 DVDD.n3490 DVDD.n3471 4.5005
R16044 DVDD.n3485 DVDD.n3471 4.5005
R16045 DVDD.n3492 DVDD.n3471 4.5005
R16046 DVDD.n3484 DVDD.n3471 4.5005
R16047 DVDD.n3493 DVDD.n3471 4.5005
R16048 DVDD.n3483 DVDD.n3471 4.5005
R16049 DVDD.n3494 DVDD.n3471 4.5005
R16050 DVDD.n3482 DVDD.n3471 4.5005
R16051 DVDD.n15790 DVDD.n3471 4.5005
R16052 DVDD.n15793 DVDD.n3471 4.5005
R16053 DVDD.n15795 DVDD.n3471 4.5005
R16054 DVDD.n3487 DVDD.n3421 4.5005
R16055 DVDD.n3489 DVDD.n3421 4.5005
R16056 DVDD.n3486 DVDD.n3421 4.5005
R16057 DVDD.n3490 DVDD.n3421 4.5005
R16058 DVDD.n3485 DVDD.n3421 4.5005
R16059 DVDD.n3492 DVDD.n3421 4.5005
R16060 DVDD.n3484 DVDD.n3421 4.5005
R16061 DVDD.n3493 DVDD.n3421 4.5005
R16062 DVDD.n3483 DVDD.n3421 4.5005
R16063 DVDD.n3494 DVDD.n3421 4.5005
R16064 DVDD.n3482 DVDD.n3421 4.5005
R16065 DVDD.n15790 DVDD.n3421 4.5005
R16066 DVDD.n3481 DVDD.n3421 4.5005
R16067 DVDD.n15793 DVDD.n3421 4.5005
R16068 DVDD.n15795 DVDD.n3421 4.5005
R16069 DVDD.n3647 DVDD.n3635 4.5005
R16070 DVDD.n3647 DVDD.n3640 4.5005
R16071 DVDD.n4769 DVDD.n3647 4.5005
R16072 DVDD.n3652 DVDD.n3647 4.5005
R16073 DVDD.n4767 DVDD.n3647 4.5005
R16074 DVDD.n3654 DVDD.n3647 4.5005
R16075 DVDD.n3665 DVDD.n3647 4.5005
R16076 DVDD.n3712 DVDD.n3647 4.5005
R16077 DVDD.n3656 DVDD.n3647 4.5005
R16078 DVDD.n4752 DVDD.n3647 4.5005
R16079 DVDD.n3645 DVDD.n3635 4.5005
R16080 DVDD.n3645 DVDD.n3640 4.5005
R16081 DVDD.n4769 DVDD.n3645 4.5005
R16082 DVDD.n3652 DVDD.n3645 4.5005
R16083 DVDD.n4767 DVDD.n3645 4.5005
R16084 DVDD.n3653 DVDD.n3645 4.5005
R16085 DVDD.n3667 DVDD.n3645 4.5005
R16086 DVDD.n3654 DVDD.n3645 4.5005
R16087 DVDD.n3665 DVDD.n3645 4.5005
R16088 DVDD.n3656 DVDD.n3645 4.5005
R16089 DVDD.n4752 DVDD.n3645 4.5005
R16090 DVDD.n4752 DVDD.n3650 4.5005
R16091 DVDD.n4752 DVDD.n3643 4.5005
R16092 DVDD.n4752 DVDD.n3648 4.5005
R16093 DVDD.n4085 DVDD.n3839 4.5005
R16094 DVDD.n4086 DVDD.n3839 4.5005
R16095 DVDD.n4084 DVDD.n3839 4.5005
R16096 DVDD.n4087 DVDD.n3839 4.5005
R16097 DVDD.n4083 DVDD.n3839 4.5005
R16098 DVDD.n4090 DVDD.n3839 4.5005
R16099 DVDD.n4081 DVDD.n3839 4.5005
R16100 DVDD.n4091 DVDD.n3839 4.5005
R16101 DVDD.n4080 DVDD.n3839 4.5005
R16102 DVDD.n4133 DVDD.n3839 4.5005
R16103 DVDD.n4079 DVDD.n3839 4.5005
R16104 DVDD.n4135 DVDD.n3839 4.5005
R16105 DVDD.n4137 DVDD.n3839 4.5005
R16106 DVDD.n4085 DVDD.n3841 4.5005
R16107 DVDD.n4086 DVDD.n3841 4.5005
R16108 DVDD.n4084 DVDD.n3841 4.5005
R16109 DVDD.n4087 DVDD.n3841 4.5005
R16110 DVDD.n4083 DVDD.n3841 4.5005
R16111 DVDD.n4089 DVDD.n3841 4.5005
R16112 DVDD.n4082 DVDD.n3841 4.5005
R16113 DVDD.n4090 DVDD.n3841 4.5005
R16114 DVDD.n4081 DVDD.n3841 4.5005
R16115 DVDD.n4091 DVDD.n3841 4.5005
R16116 DVDD.n4080 DVDD.n3841 4.5005
R16117 DVDD.n4133 DVDD.n3841 4.5005
R16118 DVDD.n4135 DVDD.n3841 4.5005
R16119 DVDD.n4137 DVDD.n3841 4.5005
R16120 DVDD.n4085 DVDD.n3838 4.5005
R16121 DVDD.n4086 DVDD.n3838 4.5005
R16122 DVDD.n4084 DVDD.n3838 4.5005
R16123 DVDD.n4087 DVDD.n3838 4.5005
R16124 DVDD.n4083 DVDD.n3838 4.5005
R16125 DVDD.n4089 DVDD.n3838 4.5005
R16126 DVDD.n4082 DVDD.n3838 4.5005
R16127 DVDD.n4090 DVDD.n3838 4.5005
R16128 DVDD.n4081 DVDD.n3838 4.5005
R16129 DVDD.n4091 DVDD.n3838 4.5005
R16130 DVDD.n4080 DVDD.n3838 4.5005
R16131 DVDD.n4133 DVDD.n3838 4.5005
R16132 DVDD.n4135 DVDD.n3838 4.5005
R16133 DVDD.n4137 DVDD.n3838 4.5005
R16134 DVDD.n4085 DVDD.n3843 4.5005
R16135 DVDD.n4086 DVDD.n3843 4.5005
R16136 DVDD.n4084 DVDD.n3843 4.5005
R16137 DVDD.n4087 DVDD.n3843 4.5005
R16138 DVDD.n4083 DVDD.n3843 4.5005
R16139 DVDD.n4089 DVDD.n3843 4.5005
R16140 DVDD.n4082 DVDD.n3843 4.5005
R16141 DVDD.n4090 DVDD.n3843 4.5005
R16142 DVDD.n4081 DVDD.n3843 4.5005
R16143 DVDD.n4091 DVDD.n3843 4.5005
R16144 DVDD.n4080 DVDD.n3843 4.5005
R16145 DVDD.n4133 DVDD.n3843 4.5005
R16146 DVDD.n4135 DVDD.n3843 4.5005
R16147 DVDD.n4137 DVDD.n3843 4.5005
R16148 DVDD.n4085 DVDD.n3837 4.5005
R16149 DVDD.n4086 DVDD.n3837 4.5005
R16150 DVDD.n4084 DVDD.n3837 4.5005
R16151 DVDD.n4087 DVDD.n3837 4.5005
R16152 DVDD.n4083 DVDD.n3837 4.5005
R16153 DVDD.n4089 DVDD.n3837 4.5005
R16154 DVDD.n4082 DVDD.n3837 4.5005
R16155 DVDD.n4090 DVDD.n3837 4.5005
R16156 DVDD.n4081 DVDD.n3837 4.5005
R16157 DVDD.n4091 DVDD.n3837 4.5005
R16158 DVDD.n4080 DVDD.n3837 4.5005
R16159 DVDD.n4133 DVDD.n3837 4.5005
R16160 DVDD.n4135 DVDD.n3837 4.5005
R16161 DVDD.n4137 DVDD.n3837 4.5005
R16162 DVDD.n4085 DVDD.n3845 4.5005
R16163 DVDD.n4086 DVDD.n3845 4.5005
R16164 DVDD.n4084 DVDD.n3845 4.5005
R16165 DVDD.n4087 DVDD.n3845 4.5005
R16166 DVDD.n4083 DVDD.n3845 4.5005
R16167 DVDD.n4089 DVDD.n3845 4.5005
R16168 DVDD.n4082 DVDD.n3845 4.5005
R16169 DVDD.n4090 DVDD.n3845 4.5005
R16170 DVDD.n4081 DVDD.n3845 4.5005
R16171 DVDD.n4091 DVDD.n3845 4.5005
R16172 DVDD.n4080 DVDD.n3845 4.5005
R16173 DVDD.n4133 DVDD.n3845 4.5005
R16174 DVDD.n4135 DVDD.n3845 4.5005
R16175 DVDD.n4137 DVDD.n3845 4.5005
R16176 DVDD.n4085 DVDD.n3836 4.5005
R16177 DVDD.n4086 DVDD.n3836 4.5005
R16178 DVDD.n4084 DVDD.n3836 4.5005
R16179 DVDD.n4087 DVDD.n3836 4.5005
R16180 DVDD.n4083 DVDD.n3836 4.5005
R16181 DVDD.n4089 DVDD.n3836 4.5005
R16182 DVDD.n4082 DVDD.n3836 4.5005
R16183 DVDD.n4090 DVDD.n3836 4.5005
R16184 DVDD.n4081 DVDD.n3836 4.5005
R16185 DVDD.n4091 DVDD.n3836 4.5005
R16186 DVDD.n4080 DVDD.n3836 4.5005
R16187 DVDD.n4133 DVDD.n3836 4.5005
R16188 DVDD.n4135 DVDD.n3836 4.5005
R16189 DVDD.n4137 DVDD.n3836 4.5005
R16190 DVDD.n4085 DVDD.n3847 4.5005
R16191 DVDD.n4086 DVDD.n3847 4.5005
R16192 DVDD.n4084 DVDD.n3847 4.5005
R16193 DVDD.n4087 DVDD.n3847 4.5005
R16194 DVDD.n4083 DVDD.n3847 4.5005
R16195 DVDD.n4089 DVDD.n3847 4.5005
R16196 DVDD.n4082 DVDD.n3847 4.5005
R16197 DVDD.n4090 DVDD.n3847 4.5005
R16198 DVDD.n4081 DVDD.n3847 4.5005
R16199 DVDD.n4091 DVDD.n3847 4.5005
R16200 DVDD.n4080 DVDD.n3847 4.5005
R16201 DVDD.n4133 DVDD.n3847 4.5005
R16202 DVDD.n4135 DVDD.n3847 4.5005
R16203 DVDD.n4137 DVDD.n3847 4.5005
R16204 DVDD.n4085 DVDD.n3835 4.5005
R16205 DVDD.n4086 DVDD.n3835 4.5005
R16206 DVDD.n4084 DVDD.n3835 4.5005
R16207 DVDD.n4087 DVDD.n3835 4.5005
R16208 DVDD.n4083 DVDD.n3835 4.5005
R16209 DVDD.n4089 DVDD.n3835 4.5005
R16210 DVDD.n4082 DVDD.n3835 4.5005
R16211 DVDD.n4090 DVDD.n3835 4.5005
R16212 DVDD.n4081 DVDD.n3835 4.5005
R16213 DVDD.n4091 DVDD.n3835 4.5005
R16214 DVDD.n4080 DVDD.n3835 4.5005
R16215 DVDD.n4133 DVDD.n3835 4.5005
R16216 DVDD.n4135 DVDD.n3835 4.5005
R16217 DVDD.n4137 DVDD.n3835 4.5005
R16218 DVDD.n4085 DVDD.n3849 4.5005
R16219 DVDD.n4086 DVDD.n3849 4.5005
R16220 DVDD.n4084 DVDD.n3849 4.5005
R16221 DVDD.n4087 DVDD.n3849 4.5005
R16222 DVDD.n4083 DVDD.n3849 4.5005
R16223 DVDD.n4089 DVDD.n3849 4.5005
R16224 DVDD.n4082 DVDD.n3849 4.5005
R16225 DVDD.n4090 DVDD.n3849 4.5005
R16226 DVDD.n4081 DVDD.n3849 4.5005
R16227 DVDD.n4091 DVDD.n3849 4.5005
R16228 DVDD.n4080 DVDD.n3849 4.5005
R16229 DVDD.n4133 DVDD.n3849 4.5005
R16230 DVDD.n4135 DVDD.n3849 4.5005
R16231 DVDD.n4137 DVDD.n3849 4.5005
R16232 DVDD.n4085 DVDD.n3834 4.5005
R16233 DVDD.n4086 DVDD.n3834 4.5005
R16234 DVDD.n4084 DVDD.n3834 4.5005
R16235 DVDD.n4087 DVDD.n3834 4.5005
R16236 DVDD.n4083 DVDD.n3834 4.5005
R16237 DVDD.n4089 DVDD.n3834 4.5005
R16238 DVDD.n4082 DVDD.n3834 4.5005
R16239 DVDD.n4090 DVDD.n3834 4.5005
R16240 DVDD.n4081 DVDD.n3834 4.5005
R16241 DVDD.n4091 DVDD.n3834 4.5005
R16242 DVDD.n4080 DVDD.n3834 4.5005
R16243 DVDD.n4133 DVDD.n3834 4.5005
R16244 DVDD.n4135 DVDD.n3834 4.5005
R16245 DVDD.n4137 DVDD.n3834 4.5005
R16246 DVDD.n4085 DVDD.n3851 4.5005
R16247 DVDD.n4086 DVDD.n3851 4.5005
R16248 DVDD.n4084 DVDD.n3851 4.5005
R16249 DVDD.n4087 DVDD.n3851 4.5005
R16250 DVDD.n4083 DVDD.n3851 4.5005
R16251 DVDD.n4089 DVDD.n3851 4.5005
R16252 DVDD.n4082 DVDD.n3851 4.5005
R16253 DVDD.n4090 DVDD.n3851 4.5005
R16254 DVDD.n4081 DVDD.n3851 4.5005
R16255 DVDD.n4091 DVDD.n3851 4.5005
R16256 DVDD.n4080 DVDD.n3851 4.5005
R16257 DVDD.n4133 DVDD.n3851 4.5005
R16258 DVDD.n4135 DVDD.n3851 4.5005
R16259 DVDD.n4137 DVDD.n3851 4.5005
R16260 DVDD.n4085 DVDD.n3833 4.5005
R16261 DVDD.n4086 DVDD.n3833 4.5005
R16262 DVDD.n4084 DVDD.n3833 4.5005
R16263 DVDD.n4087 DVDD.n3833 4.5005
R16264 DVDD.n4083 DVDD.n3833 4.5005
R16265 DVDD.n4089 DVDD.n3833 4.5005
R16266 DVDD.n4082 DVDD.n3833 4.5005
R16267 DVDD.n4090 DVDD.n3833 4.5005
R16268 DVDD.n4081 DVDD.n3833 4.5005
R16269 DVDD.n4091 DVDD.n3833 4.5005
R16270 DVDD.n4080 DVDD.n3833 4.5005
R16271 DVDD.n4133 DVDD.n3833 4.5005
R16272 DVDD.n4135 DVDD.n3833 4.5005
R16273 DVDD.n4137 DVDD.n3833 4.5005
R16274 DVDD.n4085 DVDD.n3853 4.5005
R16275 DVDD.n4086 DVDD.n3853 4.5005
R16276 DVDD.n4084 DVDD.n3853 4.5005
R16277 DVDD.n4087 DVDD.n3853 4.5005
R16278 DVDD.n4083 DVDD.n3853 4.5005
R16279 DVDD.n4089 DVDD.n3853 4.5005
R16280 DVDD.n4082 DVDD.n3853 4.5005
R16281 DVDD.n4090 DVDD.n3853 4.5005
R16282 DVDD.n4081 DVDD.n3853 4.5005
R16283 DVDD.n4091 DVDD.n3853 4.5005
R16284 DVDD.n4080 DVDD.n3853 4.5005
R16285 DVDD.n4133 DVDD.n3853 4.5005
R16286 DVDD.n4135 DVDD.n3853 4.5005
R16287 DVDD.n4137 DVDD.n3853 4.5005
R16288 DVDD.n4085 DVDD.n3832 4.5005
R16289 DVDD.n4086 DVDD.n3832 4.5005
R16290 DVDD.n4084 DVDD.n3832 4.5005
R16291 DVDD.n4087 DVDD.n3832 4.5005
R16292 DVDD.n4083 DVDD.n3832 4.5005
R16293 DVDD.n4089 DVDD.n3832 4.5005
R16294 DVDD.n4082 DVDD.n3832 4.5005
R16295 DVDD.n4090 DVDD.n3832 4.5005
R16296 DVDD.n4081 DVDD.n3832 4.5005
R16297 DVDD.n4091 DVDD.n3832 4.5005
R16298 DVDD.n4080 DVDD.n3832 4.5005
R16299 DVDD.n4133 DVDD.n3832 4.5005
R16300 DVDD.n4135 DVDD.n3832 4.5005
R16301 DVDD.n4137 DVDD.n3832 4.5005
R16302 DVDD.n4085 DVDD.n3855 4.5005
R16303 DVDD.n4086 DVDD.n3855 4.5005
R16304 DVDD.n4084 DVDD.n3855 4.5005
R16305 DVDD.n4087 DVDD.n3855 4.5005
R16306 DVDD.n4083 DVDD.n3855 4.5005
R16307 DVDD.n4089 DVDD.n3855 4.5005
R16308 DVDD.n4082 DVDD.n3855 4.5005
R16309 DVDD.n4090 DVDD.n3855 4.5005
R16310 DVDD.n4081 DVDD.n3855 4.5005
R16311 DVDD.n4091 DVDD.n3855 4.5005
R16312 DVDD.n4080 DVDD.n3855 4.5005
R16313 DVDD.n4133 DVDD.n3855 4.5005
R16314 DVDD.n4135 DVDD.n3855 4.5005
R16315 DVDD.n4137 DVDD.n3855 4.5005
R16316 DVDD.n4085 DVDD.n3831 4.5005
R16317 DVDD.n4086 DVDD.n3831 4.5005
R16318 DVDD.n4084 DVDD.n3831 4.5005
R16319 DVDD.n4087 DVDD.n3831 4.5005
R16320 DVDD.n4083 DVDD.n3831 4.5005
R16321 DVDD.n4089 DVDD.n3831 4.5005
R16322 DVDD.n4082 DVDD.n3831 4.5005
R16323 DVDD.n4090 DVDD.n3831 4.5005
R16324 DVDD.n4081 DVDD.n3831 4.5005
R16325 DVDD.n4091 DVDD.n3831 4.5005
R16326 DVDD.n4080 DVDD.n3831 4.5005
R16327 DVDD.n4133 DVDD.n3831 4.5005
R16328 DVDD.n4135 DVDD.n3831 4.5005
R16329 DVDD.n4137 DVDD.n3831 4.5005
R16330 DVDD.n4085 DVDD.n3857 4.5005
R16331 DVDD.n4086 DVDD.n3857 4.5005
R16332 DVDD.n4084 DVDD.n3857 4.5005
R16333 DVDD.n4087 DVDD.n3857 4.5005
R16334 DVDD.n4083 DVDD.n3857 4.5005
R16335 DVDD.n4089 DVDD.n3857 4.5005
R16336 DVDD.n4082 DVDD.n3857 4.5005
R16337 DVDD.n4090 DVDD.n3857 4.5005
R16338 DVDD.n4081 DVDD.n3857 4.5005
R16339 DVDD.n4091 DVDD.n3857 4.5005
R16340 DVDD.n4080 DVDD.n3857 4.5005
R16341 DVDD.n4133 DVDD.n3857 4.5005
R16342 DVDD.n4135 DVDD.n3857 4.5005
R16343 DVDD.n4137 DVDD.n3857 4.5005
R16344 DVDD.n4085 DVDD.n3830 4.5005
R16345 DVDD.n4086 DVDD.n3830 4.5005
R16346 DVDD.n4084 DVDD.n3830 4.5005
R16347 DVDD.n4087 DVDD.n3830 4.5005
R16348 DVDD.n4083 DVDD.n3830 4.5005
R16349 DVDD.n4089 DVDD.n3830 4.5005
R16350 DVDD.n4082 DVDD.n3830 4.5005
R16351 DVDD.n4090 DVDD.n3830 4.5005
R16352 DVDD.n4081 DVDD.n3830 4.5005
R16353 DVDD.n4091 DVDD.n3830 4.5005
R16354 DVDD.n4080 DVDD.n3830 4.5005
R16355 DVDD.n4133 DVDD.n3830 4.5005
R16356 DVDD.n4135 DVDD.n3830 4.5005
R16357 DVDD.n4137 DVDD.n3830 4.5005
R16358 DVDD.n4085 DVDD.n3859 4.5005
R16359 DVDD.n4086 DVDD.n3859 4.5005
R16360 DVDD.n4084 DVDD.n3859 4.5005
R16361 DVDD.n4087 DVDD.n3859 4.5005
R16362 DVDD.n4083 DVDD.n3859 4.5005
R16363 DVDD.n4089 DVDD.n3859 4.5005
R16364 DVDD.n4082 DVDD.n3859 4.5005
R16365 DVDD.n4090 DVDD.n3859 4.5005
R16366 DVDD.n4081 DVDD.n3859 4.5005
R16367 DVDD.n4091 DVDD.n3859 4.5005
R16368 DVDD.n4080 DVDD.n3859 4.5005
R16369 DVDD.n4133 DVDD.n3859 4.5005
R16370 DVDD.n4135 DVDD.n3859 4.5005
R16371 DVDD.n4137 DVDD.n3859 4.5005
R16372 DVDD.n4085 DVDD.n3829 4.5005
R16373 DVDD.n4086 DVDD.n3829 4.5005
R16374 DVDD.n4084 DVDD.n3829 4.5005
R16375 DVDD.n4087 DVDD.n3829 4.5005
R16376 DVDD.n4083 DVDD.n3829 4.5005
R16377 DVDD.n4089 DVDD.n3829 4.5005
R16378 DVDD.n4082 DVDD.n3829 4.5005
R16379 DVDD.n4090 DVDD.n3829 4.5005
R16380 DVDD.n4081 DVDD.n3829 4.5005
R16381 DVDD.n4091 DVDD.n3829 4.5005
R16382 DVDD.n4080 DVDD.n3829 4.5005
R16383 DVDD.n4133 DVDD.n3829 4.5005
R16384 DVDD.n4135 DVDD.n3829 4.5005
R16385 DVDD.n4137 DVDD.n3829 4.5005
R16386 DVDD.n4085 DVDD.n3861 4.5005
R16387 DVDD.n4086 DVDD.n3861 4.5005
R16388 DVDD.n4084 DVDD.n3861 4.5005
R16389 DVDD.n4087 DVDD.n3861 4.5005
R16390 DVDD.n4083 DVDD.n3861 4.5005
R16391 DVDD.n4089 DVDD.n3861 4.5005
R16392 DVDD.n4082 DVDD.n3861 4.5005
R16393 DVDD.n4090 DVDD.n3861 4.5005
R16394 DVDD.n4081 DVDD.n3861 4.5005
R16395 DVDD.n4091 DVDD.n3861 4.5005
R16396 DVDD.n4080 DVDD.n3861 4.5005
R16397 DVDD.n4133 DVDD.n3861 4.5005
R16398 DVDD.n4135 DVDD.n3861 4.5005
R16399 DVDD.n4137 DVDD.n3861 4.5005
R16400 DVDD.n4085 DVDD.n3828 4.5005
R16401 DVDD.n4086 DVDD.n3828 4.5005
R16402 DVDD.n4084 DVDD.n3828 4.5005
R16403 DVDD.n4087 DVDD.n3828 4.5005
R16404 DVDD.n4083 DVDD.n3828 4.5005
R16405 DVDD.n4089 DVDD.n3828 4.5005
R16406 DVDD.n4082 DVDD.n3828 4.5005
R16407 DVDD.n4090 DVDD.n3828 4.5005
R16408 DVDD.n4081 DVDD.n3828 4.5005
R16409 DVDD.n4091 DVDD.n3828 4.5005
R16410 DVDD.n4080 DVDD.n3828 4.5005
R16411 DVDD.n4133 DVDD.n3828 4.5005
R16412 DVDD.n4135 DVDD.n3828 4.5005
R16413 DVDD.n4137 DVDD.n3828 4.5005
R16414 DVDD.n4136 DVDD.n4085 4.5005
R16415 DVDD.n4136 DVDD.n4086 4.5005
R16416 DVDD.n4136 DVDD.n4084 4.5005
R16417 DVDD.n4136 DVDD.n4087 4.5005
R16418 DVDD.n4136 DVDD.n4083 4.5005
R16419 DVDD.n4136 DVDD.n4089 4.5005
R16420 DVDD.n4136 DVDD.n4082 4.5005
R16421 DVDD.n4136 DVDD.n4090 4.5005
R16422 DVDD.n4136 DVDD.n4081 4.5005
R16423 DVDD.n4136 DVDD.n4091 4.5005
R16424 DVDD.n4136 DVDD.n4080 4.5005
R16425 DVDD.n4136 DVDD.n4133 4.5005
R16426 DVDD.n4136 DVDD.n4079 4.5005
R16427 DVDD.n4136 DVDD.n4135 4.5005
R16428 DVDD.n4137 DVDD.n4136 4.5005
R16429 DVDD.n4066 DVDD.n3869 4.5005
R16430 DVDD.n4066 DVDD.n3870 4.5005
R16431 DVDD.n4066 DVDD.n3868 4.5005
R16432 DVDD.n4066 DVDD.n3871 4.5005
R16433 DVDD.n4066 DVDD.n3867 4.5005
R16434 DVDD.n4066 DVDD.n3872 4.5005
R16435 DVDD.n4066 DVDD.n3865 4.5005
R16436 DVDD.n4066 DVDD.n3873 4.5005
R16437 DVDD.n4066 DVDD.n3864 4.5005
R16438 DVDD.n4066 DVDD.n3874 4.5005
R16439 DVDD.n4066 DVDD.n3863 4.5005
R16440 DVDD.n4066 DVDD.n3875 4.5005
R16441 DVDD.n4066 DVDD.n4065 4.5005
R16442 DVDD.n3882 DVDD.n3869 4.5005
R16443 DVDD.n3882 DVDD.n3870 4.5005
R16444 DVDD.n3882 DVDD.n3868 4.5005
R16445 DVDD.n3882 DVDD.n3871 4.5005
R16446 DVDD.n3882 DVDD.n3867 4.5005
R16447 DVDD.n4063 DVDD.n3882 4.5005
R16448 DVDD.n3897 DVDD.n3882 4.5005
R16449 DVDD.n3882 DVDD.n3872 4.5005
R16450 DVDD.n3882 DVDD.n3865 4.5005
R16451 DVDD.n3882 DVDD.n3873 4.5005
R16452 DVDD.n3882 DVDD.n3864 4.5005
R16453 DVDD.n3882 DVDD.n3874 4.5005
R16454 DVDD.n3882 DVDD.n3875 4.5005
R16455 DVDD.n4065 DVDD.n3882 4.5005
R16456 DVDD.n3885 DVDD.n3869 4.5005
R16457 DVDD.n3885 DVDD.n3870 4.5005
R16458 DVDD.n3885 DVDD.n3868 4.5005
R16459 DVDD.n3885 DVDD.n3871 4.5005
R16460 DVDD.n3885 DVDD.n3867 4.5005
R16461 DVDD.n4063 DVDD.n3885 4.5005
R16462 DVDD.n3897 DVDD.n3885 4.5005
R16463 DVDD.n3885 DVDD.n3872 4.5005
R16464 DVDD.n3885 DVDD.n3865 4.5005
R16465 DVDD.n3885 DVDD.n3873 4.5005
R16466 DVDD.n3885 DVDD.n3864 4.5005
R16467 DVDD.n3885 DVDD.n3874 4.5005
R16468 DVDD.n3885 DVDD.n3875 4.5005
R16469 DVDD.n4065 DVDD.n3885 4.5005
R16470 DVDD.n3881 DVDD.n3869 4.5005
R16471 DVDD.n3881 DVDD.n3870 4.5005
R16472 DVDD.n3881 DVDD.n3868 4.5005
R16473 DVDD.n3881 DVDD.n3871 4.5005
R16474 DVDD.n3881 DVDD.n3867 4.5005
R16475 DVDD.n4063 DVDD.n3881 4.5005
R16476 DVDD.n3897 DVDD.n3881 4.5005
R16477 DVDD.n3881 DVDD.n3872 4.5005
R16478 DVDD.n3881 DVDD.n3865 4.5005
R16479 DVDD.n3881 DVDD.n3873 4.5005
R16480 DVDD.n3881 DVDD.n3864 4.5005
R16481 DVDD.n3881 DVDD.n3874 4.5005
R16482 DVDD.n3881 DVDD.n3875 4.5005
R16483 DVDD.n4065 DVDD.n3881 4.5005
R16484 DVDD.n3887 DVDD.n3869 4.5005
R16485 DVDD.n3887 DVDD.n3870 4.5005
R16486 DVDD.n3887 DVDD.n3868 4.5005
R16487 DVDD.n3887 DVDD.n3871 4.5005
R16488 DVDD.n3887 DVDD.n3867 4.5005
R16489 DVDD.n4063 DVDD.n3887 4.5005
R16490 DVDD.n3897 DVDD.n3887 4.5005
R16491 DVDD.n3887 DVDD.n3872 4.5005
R16492 DVDD.n3887 DVDD.n3865 4.5005
R16493 DVDD.n3887 DVDD.n3873 4.5005
R16494 DVDD.n3887 DVDD.n3864 4.5005
R16495 DVDD.n3887 DVDD.n3874 4.5005
R16496 DVDD.n3887 DVDD.n3875 4.5005
R16497 DVDD.n4065 DVDD.n3887 4.5005
R16498 DVDD.n3880 DVDD.n3869 4.5005
R16499 DVDD.n3880 DVDD.n3870 4.5005
R16500 DVDD.n3880 DVDD.n3868 4.5005
R16501 DVDD.n3880 DVDD.n3871 4.5005
R16502 DVDD.n3880 DVDD.n3867 4.5005
R16503 DVDD.n4063 DVDD.n3880 4.5005
R16504 DVDD.n3897 DVDD.n3880 4.5005
R16505 DVDD.n3880 DVDD.n3872 4.5005
R16506 DVDD.n3880 DVDD.n3865 4.5005
R16507 DVDD.n3880 DVDD.n3873 4.5005
R16508 DVDD.n3880 DVDD.n3864 4.5005
R16509 DVDD.n3880 DVDD.n3874 4.5005
R16510 DVDD.n3880 DVDD.n3875 4.5005
R16511 DVDD.n4065 DVDD.n3880 4.5005
R16512 DVDD.n3889 DVDD.n3869 4.5005
R16513 DVDD.n3889 DVDD.n3870 4.5005
R16514 DVDD.n3889 DVDD.n3868 4.5005
R16515 DVDD.n3889 DVDD.n3871 4.5005
R16516 DVDD.n3889 DVDD.n3867 4.5005
R16517 DVDD.n4063 DVDD.n3889 4.5005
R16518 DVDD.n3897 DVDD.n3889 4.5005
R16519 DVDD.n3889 DVDD.n3872 4.5005
R16520 DVDD.n3889 DVDD.n3865 4.5005
R16521 DVDD.n3889 DVDD.n3873 4.5005
R16522 DVDD.n3889 DVDD.n3864 4.5005
R16523 DVDD.n3889 DVDD.n3874 4.5005
R16524 DVDD.n3889 DVDD.n3875 4.5005
R16525 DVDD.n4065 DVDD.n3889 4.5005
R16526 DVDD.n3879 DVDD.n3869 4.5005
R16527 DVDD.n3879 DVDD.n3870 4.5005
R16528 DVDD.n3879 DVDD.n3868 4.5005
R16529 DVDD.n3879 DVDD.n3871 4.5005
R16530 DVDD.n3879 DVDD.n3867 4.5005
R16531 DVDD.n4063 DVDD.n3879 4.5005
R16532 DVDD.n3897 DVDD.n3879 4.5005
R16533 DVDD.n3879 DVDD.n3872 4.5005
R16534 DVDD.n3879 DVDD.n3865 4.5005
R16535 DVDD.n3879 DVDD.n3873 4.5005
R16536 DVDD.n3879 DVDD.n3864 4.5005
R16537 DVDD.n3879 DVDD.n3874 4.5005
R16538 DVDD.n3879 DVDD.n3875 4.5005
R16539 DVDD.n4065 DVDD.n3879 4.5005
R16540 DVDD.n4064 DVDD.n3869 4.5005
R16541 DVDD.n4064 DVDD.n3870 4.5005
R16542 DVDD.n4064 DVDD.n3868 4.5005
R16543 DVDD.n4064 DVDD.n3871 4.5005
R16544 DVDD.n4064 DVDD.n3867 4.5005
R16545 DVDD.n4064 DVDD.n4063 4.5005
R16546 DVDD.n4064 DVDD.n3897 4.5005
R16547 DVDD.n4064 DVDD.n3872 4.5005
R16548 DVDD.n4064 DVDD.n3865 4.5005
R16549 DVDD.n4064 DVDD.n3873 4.5005
R16550 DVDD.n4064 DVDD.n3864 4.5005
R16551 DVDD.n4064 DVDD.n3874 4.5005
R16552 DVDD.n4064 DVDD.n3875 4.5005
R16553 DVDD.n4065 DVDD.n4064 4.5005
R16554 DVDD.n3878 DVDD.n3869 4.5005
R16555 DVDD.n3878 DVDD.n3870 4.5005
R16556 DVDD.n3878 DVDD.n3868 4.5005
R16557 DVDD.n3878 DVDD.n3871 4.5005
R16558 DVDD.n3878 DVDD.n3867 4.5005
R16559 DVDD.n4063 DVDD.n3878 4.5005
R16560 DVDD.n3897 DVDD.n3878 4.5005
R16561 DVDD.n3878 DVDD.n3872 4.5005
R16562 DVDD.n3878 DVDD.n3865 4.5005
R16563 DVDD.n3878 DVDD.n3873 4.5005
R16564 DVDD.n3878 DVDD.n3864 4.5005
R16565 DVDD.n3878 DVDD.n3874 4.5005
R16566 DVDD.n3878 DVDD.n3875 4.5005
R16567 DVDD.n4065 DVDD.n3878 4.5005
R16568 DVDD.n3869 DVDD.n231 4.5005
R16569 DVDD.n3870 DVDD.n231 4.5005
R16570 DVDD.n3868 DVDD.n231 4.5005
R16571 DVDD.n3871 DVDD.n231 4.5005
R16572 DVDD.n3867 DVDD.n231 4.5005
R16573 DVDD.n4063 DVDD.n231 4.5005
R16574 DVDD.n3897 DVDD.n231 4.5005
R16575 DVDD.n3872 DVDD.n231 4.5005
R16576 DVDD.n3865 DVDD.n231 4.5005
R16577 DVDD.n3873 DVDD.n231 4.5005
R16578 DVDD.n3864 DVDD.n231 4.5005
R16579 DVDD.n3874 DVDD.n231 4.5005
R16580 DVDD.n4065 DVDD.n231 4.5005
R16581 DVDD.n18838 DVDD.n18829 4.5005
R16582 DVDD.n18839 DVDD.n18829 4.5005
R16583 DVDD.n18837 DVDD.n18829 4.5005
R16584 DVDD.n18840 DVDD.n18829 4.5005
R16585 DVDD.n18836 DVDD.n18829 4.5005
R16586 DVDD.n18843 DVDD.n18829 4.5005
R16587 DVDD.n18834 DVDD.n18829 4.5005
R16588 DVDD.n18844 DVDD.n18829 4.5005
R16589 DVDD.n18833 DVDD.n18829 4.5005
R16590 DVDD.n18845 DVDD.n18829 4.5005
R16591 DVDD.n18832 DVDD.n18829 4.5005
R16592 DVDD.n20970 DVDD.n18829 4.5005
R16593 DVDD.n20971 DVDD.n18838 4.5005
R16594 DVDD.n20971 DVDD.n18839 4.5005
R16595 DVDD.n20971 DVDD.n18837 4.5005
R16596 DVDD.n20971 DVDD.n18840 4.5005
R16597 DVDD.n20971 DVDD.n18836 4.5005
R16598 DVDD.n20971 DVDD.n18842 4.5005
R16599 DVDD.n20971 DVDD.n18835 4.5005
R16600 DVDD.n20971 DVDD.n18843 4.5005
R16601 DVDD.n20971 DVDD.n18834 4.5005
R16602 DVDD.n20971 DVDD.n18844 4.5005
R16603 DVDD.n20971 DVDD.n18833 4.5005
R16604 DVDD.n20971 DVDD.n18845 4.5005
R16605 DVDD.n20971 DVDD.n18832 4.5005
R16606 DVDD.n20971 DVDD.n18846 4.5005
R16607 DVDD.n20971 DVDD.n20970 4.5005
R16608 DVDD.n18855 DVDD.n18838 4.5005
R16609 DVDD.n18855 DVDD.n18839 4.5005
R16610 DVDD.n18855 DVDD.n18837 4.5005
R16611 DVDD.n18855 DVDD.n18840 4.5005
R16612 DVDD.n18855 DVDD.n18836 4.5005
R16613 DVDD.n18855 DVDD.n18842 4.5005
R16614 DVDD.n18855 DVDD.n18835 4.5005
R16615 DVDD.n18855 DVDD.n18843 4.5005
R16616 DVDD.n18855 DVDD.n18834 4.5005
R16617 DVDD.n18855 DVDD.n18844 4.5005
R16618 DVDD.n18855 DVDD.n18833 4.5005
R16619 DVDD.n18855 DVDD.n18845 4.5005
R16620 DVDD.n18855 DVDD.n18846 4.5005
R16621 DVDD.n20970 DVDD.n18855 4.5005
R16622 DVDD.n18852 DVDD.n18838 4.5005
R16623 DVDD.n18852 DVDD.n18839 4.5005
R16624 DVDD.n18852 DVDD.n18837 4.5005
R16625 DVDD.n18852 DVDD.n18840 4.5005
R16626 DVDD.n18852 DVDD.n18836 4.5005
R16627 DVDD.n18852 DVDD.n18842 4.5005
R16628 DVDD.n18852 DVDD.n18835 4.5005
R16629 DVDD.n18852 DVDD.n18843 4.5005
R16630 DVDD.n18852 DVDD.n18834 4.5005
R16631 DVDD.n18852 DVDD.n18844 4.5005
R16632 DVDD.n18852 DVDD.n18833 4.5005
R16633 DVDD.n18852 DVDD.n18845 4.5005
R16634 DVDD.n18852 DVDD.n18846 4.5005
R16635 DVDD.n20970 DVDD.n18852 4.5005
R16636 DVDD.n18857 DVDD.n18838 4.5005
R16637 DVDD.n18857 DVDD.n18839 4.5005
R16638 DVDD.n18857 DVDD.n18837 4.5005
R16639 DVDD.n18857 DVDD.n18840 4.5005
R16640 DVDD.n18857 DVDD.n18836 4.5005
R16641 DVDD.n18857 DVDD.n18842 4.5005
R16642 DVDD.n18857 DVDD.n18835 4.5005
R16643 DVDD.n18857 DVDD.n18843 4.5005
R16644 DVDD.n18857 DVDD.n18834 4.5005
R16645 DVDD.n18857 DVDD.n18844 4.5005
R16646 DVDD.n18857 DVDD.n18833 4.5005
R16647 DVDD.n18857 DVDD.n18845 4.5005
R16648 DVDD.n18857 DVDD.n18846 4.5005
R16649 DVDD.n20970 DVDD.n18857 4.5005
R16650 DVDD.n18851 DVDD.n18838 4.5005
R16651 DVDD.n18851 DVDD.n18839 4.5005
R16652 DVDD.n18851 DVDD.n18837 4.5005
R16653 DVDD.n18851 DVDD.n18840 4.5005
R16654 DVDD.n18851 DVDD.n18836 4.5005
R16655 DVDD.n18851 DVDD.n18842 4.5005
R16656 DVDD.n18851 DVDD.n18835 4.5005
R16657 DVDD.n18851 DVDD.n18843 4.5005
R16658 DVDD.n18851 DVDD.n18834 4.5005
R16659 DVDD.n18851 DVDD.n18844 4.5005
R16660 DVDD.n18851 DVDD.n18833 4.5005
R16661 DVDD.n18851 DVDD.n18845 4.5005
R16662 DVDD.n18851 DVDD.n18846 4.5005
R16663 DVDD.n20970 DVDD.n18851 4.5005
R16664 DVDD.n18858 DVDD.n18838 4.5005
R16665 DVDD.n18858 DVDD.n18839 4.5005
R16666 DVDD.n18858 DVDD.n18837 4.5005
R16667 DVDD.n18858 DVDD.n18840 4.5005
R16668 DVDD.n18858 DVDD.n18836 4.5005
R16669 DVDD.n18858 DVDD.n18842 4.5005
R16670 DVDD.n18858 DVDD.n18835 4.5005
R16671 DVDD.n18858 DVDD.n18843 4.5005
R16672 DVDD.n18858 DVDD.n18834 4.5005
R16673 DVDD.n18858 DVDD.n18844 4.5005
R16674 DVDD.n18858 DVDD.n18833 4.5005
R16675 DVDD.n18858 DVDD.n18845 4.5005
R16676 DVDD.n18858 DVDD.n18832 4.5005
R16677 DVDD.n18858 DVDD.n18846 4.5005
R16678 DVDD.n20970 DVDD.n18858 4.5005
R16679 DVDD.n18850 DVDD.n18838 4.5005
R16680 DVDD.n18850 DVDD.n18839 4.5005
R16681 DVDD.n18850 DVDD.n18837 4.5005
R16682 DVDD.n18850 DVDD.n18840 4.5005
R16683 DVDD.n18850 DVDD.n18836 4.5005
R16684 DVDD.n18850 DVDD.n18842 4.5005
R16685 DVDD.n18850 DVDD.n18835 4.5005
R16686 DVDD.n18850 DVDD.n18843 4.5005
R16687 DVDD.n18850 DVDD.n18834 4.5005
R16688 DVDD.n18850 DVDD.n18844 4.5005
R16689 DVDD.n18850 DVDD.n18833 4.5005
R16690 DVDD.n18850 DVDD.n18845 4.5005
R16691 DVDD.n18850 DVDD.n18846 4.5005
R16692 DVDD.n20970 DVDD.n18850 4.5005
R16693 DVDD.n18859 DVDD.n18838 4.5005
R16694 DVDD.n18859 DVDD.n18839 4.5005
R16695 DVDD.n18859 DVDD.n18837 4.5005
R16696 DVDD.n18859 DVDD.n18840 4.5005
R16697 DVDD.n18859 DVDD.n18836 4.5005
R16698 DVDD.n18859 DVDD.n18842 4.5005
R16699 DVDD.n18859 DVDD.n18835 4.5005
R16700 DVDD.n18859 DVDD.n18843 4.5005
R16701 DVDD.n18859 DVDD.n18834 4.5005
R16702 DVDD.n18859 DVDD.n18844 4.5005
R16703 DVDD.n18859 DVDD.n18833 4.5005
R16704 DVDD.n18859 DVDD.n18845 4.5005
R16705 DVDD.n18859 DVDD.n18832 4.5005
R16706 DVDD.n18859 DVDD.n18846 4.5005
R16707 DVDD.n20970 DVDD.n18859 4.5005
R16708 DVDD.n19748 DVDD.n19731 4.5005
R16709 DVDD.n19748 DVDD.n19733 4.5005
R16710 DVDD.n19748 DVDD.n19730 4.5005
R16711 DVDD.n19748 DVDD.n19734 4.5005
R16712 DVDD.n19748 DVDD.n19729 4.5005
R16713 DVDD.n19748 DVDD.n19736 4.5005
R16714 DVDD.n19748 DVDD.n19727 4.5005
R16715 DVDD.n19748 DVDD.n19737 4.5005
R16716 DVDD.n19748 DVDD.n19726 4.5005
R16717 DVDD.n19748 DVDD.n19738 4.5005
R16718 DVDD.n19748 DVDD.n19725 4.5005
R16719 DVDD.n20572 DVDD.n19748 4.5005
R16720 DVDD.n19744 DVDD.n19731 4.5005
R16721 DVDD.n19744 DVDD.n19733 4.5005
R16722 DVDD.n19744 DVDD.n19730 4.5005
R16723 DVDD.n19744 DVDD.n19734 4.5005
R16724 DVDD.n19744 DVDD.n19729 4.5005
R16725 DVDD.n19744 DVDD.n19735 4.5005
R16726 DVDD.n19744 DVDD.n19728 4.5005
R16727 DVDD.n19744 DVDD.n19736 4.5005
R16728 DVDD.n19744 DVDD.n19727 4.5005
R16729 DVDD.n19744 DVDD.n19737 4.5005
R16730 DVDD.n19744 DVDD.n19726 4.5005
R16731 DVDD.n19744 DVDD.n19738 4.5005
R16732 DVDD.n19744 DVDD.n19725 4.5005
R16733 DVDD.n19744 DVDD.n19739 4.5005
R16734 DVDD.n19744 DVDD.n19724 4.5005
R16735 DVDD.n20572 DVDD.n19744 4.5005
R16736 DVDD.n19749 DVDD.n19731 4.5005
R16737 DVDD.n19749 DVDD.n19733 4.5005
R16738 DVDD.n19749 DVDD.n19730 4.5005
R16739 DVDD.n19749 DVDD.n19734 4.5005
R16740 DVDD.n19749 DVDD.n19729 4.5005
R16741 DVDD.n19749 DVDD.n19735 4.5005
R16742 DVDD.n19749 DVDD.n19728 4.5005
R16743 DVDD.n19749 DVDD.n19736 4.5005
R16744 DVDD.n19749 DVDD.n19727 4.5005
R16745 DVDD.n19749 DVDD.n19737 4.5005
R16746 DVDD.n19749 DVDD.n19726 4.5005
R16747 DVDD.n19749 DVDD.n19738 4.5005
R16748 DVDD.n19749 DVDD.n19725 4.5005
R16749 DVDD.n19749 DVDD.n19739 4.5005
R16750 DVDD.n19749 DVDD.n19724 4.5005
R16751 DVDD.n20572 DVDD.n19749 4.5005
R16752 DVDD.n19743 DVDD.n19731 4.5005
R16753 DVDD.n19743 DVDD.n19733 4.5005
R16754 DVDD.n19743 DVDD.n19730 4.5005
R16755 DVDD.n19743 DVDD.n19734 4.5005
R16756 DVDD.n19743 DVDD.n19729 4.5005
R16757 DVDD.n19743 DVDD.n19735 4.5005
R16758 DVDD.n19743 DVDD.n19728 4.5005
R16759 DVDD.n19743 DVDD.n19736 4.5005
R16760 DVDD.n19743 DVDD.n19727 4.5005
R16761 DVDD.n19743 DVDD.n19737 4.5005
R16762 DVDD.n19743 DVDD.n19726 4.5005
R16763 DVDD.n19743 DVDD.n19738 4.5005
R16764 DVDD.n19743 DVDD.n19725 4.5005
R16765 DVDD.n19743 DVDD.n19739 4.5005
R16766 DVDD.n19743 DVDD.n19724 4.5005
R16767 DVDD.n20572 DVDD.n19743 4.5005
R16768 DVDD.n19750 DVDD.n19731 4.5005
R16769 DVDD.n19750 DVDD.n19733 4.5005
R16770 DVDD.n19750 DVDD.n19730 4.5005
R16771 DVDD.n19750 DVDD.n19734 4.5005
R16772 DVDD.n19750 DVDD.n19729 4.5005
R16773 DVDD.n19750 DVDD.n19735 4.5005
R16774 DVDD.n19750 DVDD.n19728 4.5005
R16775 DVDD.n19750 DVDD.n19736 4.5005
R16776 DVDD.n19750 DVDD.n19727 4.5005
R16777 DVDD.n19750 DVDD.n19737 4.5005
R16778 DVDD.n19750 DVDD.n19726 4.5005
R16779 DVDD.n19750 DVDD.n19738 4.5005
R16780 DVDD.n19750 DVDD.n19725 4.5005
R16781 DVDD.n19750 DVDD.n19739 4.5005
R16782 DVDD.n19750 DVDD.n19724 4.5005
R16783 DVDD.n20572 DVDD.n19750 4.5005
R16784 DVDD.n19742 DVDD.n19731 4.5005
R16785 DVDD.n19742 DVDD.n19733 4.5005
R16786 DVDD.n19742 DVDD.n19730 4.5005
R16787 DVDD.n19742 DVDD.n19734 4.5005
R16788 DVDD.n19742 DVDD.n19729 4.5005
R16789 DVDD.n19742 DVDD.n19735 4.5005
R16790 DVDD.n19742 DVDD.n19728 4.5005
R16791 DVDD.n19742 DVDD.n19736 4.5005
R16792 DVDD.n19742 DVDD.n19727 4.5005
R16793 DVDD.n19742 DVDD.n19737 4.5005
R16794 DVDD.n19742 DVDD.n19726 4.5005
R16795 DVDD.n19742 DVDD.n19738 4.5005
R16796 DVDD.n19742 DVDD.n19725 4.5005
R16797 DVDD.n19742 DVDD.n19739 4.5005
R16798 DVDD.n19742 DVDD.n19724 4.5005
R16799 DVDD.n20572 DVDD.n19742 4.5005
R16800 DVDD.n20571 DVDD.n19731 4.5005
R16801 DVDD.n20571 DVDD.n19733 4.5005
R16802 DVDD.n20571 DVDD.n19730 4.5005
R16803 DVDD.n20571 DVDD.n19734 4.5005
R16804 DVDD.n20571 DVDD.n19729 4.5005
R16805 DVDD.n20571 DVDD.n19735 4.5005
R16806 DVDD.n20571 DVDD.n19728 4.5005
R16807 DVDD.n20571 DVDD.n19736 4.5005
R16808 DVDD.n20571 DVDD.n19727 4.5005
R16809 DVDD.n20571 DVDD.n19737 4.5005
R16810 DVDD.n20571 DVDD.n19726 4.5005
R16811 DVDD.n20571 DVDD.n19738 4.5005
R16812 DVDD.n20571 DVDD.n19725 4.5005
R16813 DVDD.n20571 DVDD.n19739 4.5005
R16814 DVDD.n20571 DVDD.n19724 4.5005
R16815 DVDD.n20572 DVDD.n20571 4.5005
R16816 DVDD.n19741 DVDD.n19731 4.5005
R16817 DVDD.n19741 DVDD.n19733 4.5005
R16818 DVDD.n19741 DVDD.n19730 4.5005
R16819 DVDD.n19741 DVDD.n19734 4.5005
R16820 DVDD.n19741 DVDD.n19729 4.5005
R16821 DVDD.n19741 DVDD.n19735 4.5005
R16822 DVDD.n19741 DVDD.n19728 4.5005
R16823 DVDD.n19741 DVDD.n19736 4.5005
R16824 DVDD.n19741 DVDD.n19727 4.5005
R16825 DVDD.n19741 DVDD.n19737 4.5005
R16826 DVDD.n19741 DVDD.n19726 4.5005
R16827 DVDD.n19741 DVDD.n19738 4.5005
R16828 DVDD.n19741 DVDD.n19725 4.5005
R16829 DVDD.n19741 DVDD.n19739 4.5005
R16830 DVDD.n19741 DVDD.n19724 4.5005
R16831 DVDD.n20572 DVDD.n19741 4.5005
R16832 DVDD.n20573 DVDD.n19731 4.5005
R16833 DVDD.n20573 DVDD.n19733 4.5005
R16834 DVDD.n20573 DVDD.n19730 4.5005
R16835 DVDD.n20573 DVDD.n19734 4.5005
R16836 DVDD.n20573 DVDD.n19729 4.5005
R16837 DVDD.n20573 DVDD.n19735 4.5005
R16838 DVDD.n20573 DVDD.n19728 4.5005
R16839 DVDD.n20573 DVDD.n19736 4.5005
R16840 DVDD.n20573 DVDD.n19727 4.5005
R16841 DVDD.n20573 DVDD.n19737 4.5005
R16842 DVDD.n20573 DVDD.n19726 4.5005
R16843 DVDD.n20573 DVDD.n19738 4.5005
R16844 DVDD.n20573 DVDD.n19725 4.5005
R16845 DVDD.n20573 DVDD.n19739 4.5005
R16846 DVDD.n20573 DVDD.n19724 4.5005
R16847 DVDD.n20573 DVDD.n20572 4.5005
R16848 DVDD.n19731 DVDD.n19722 4.5005
R16849 DVDD.n19733 DVDD.n19722 4.5005
R16850 DVDD.n19730 DVDD.n19722 4.5005
R16851 DVDD.n19734 DVDD.n19722 4.5005
R16852 DVDD.n19729 DVDD.n19722 4.5005
R16853 DVDD.n19735 DVDD.n19722 4.5005
R16854 DVDD.n19728 DVDD.n19722 4.5005
R16855 DVDD.n19736 DVDD.n19722 4.5005
R16856 DVDD.n19727 DVDD.n19722 4.5005
R16857 DVDD.n19737 DVDD.n19722 4.5005
R16858 DVDD.n19726 DVDD.n19722 4.5005
R16859 DVDD.n19738 DVDD.n19722 4.5005
R16860 DVDD.n19725 DVDD.n19722 4.5005
R16861 DVDD.n19739 DVDD.n19722 4.5005
R16862 DVDD.n19724 DVDD.n19722 4.5005
R16863 DVDD.n20572 DVDD.n19722 4.5005
R16864 DVDD.n19731 DVDD.n19721 4.5005
R16865 DVDD.n19733 DVDD.n19721 4.5005
R16866 DVDD.n19730 DVDD.n19721 4.5005
R16867 DVDD.n19734 DVDD.n19721 4.5005
R16868 DVDD.n19729 DVDD.n19721 4.5005
R16869 DVDD.n19735 DVDD.n19721 4.5005
R16870 DVDD.n19728 DVDD.n19721 4.5005
R16871 DVDD.n19736 DVDD.n19721 4.5005
R16872 DVDD.n19727 DVDD.n19721 4.5005
R16873 DVDD.n19737 DVDD.n19721 4.5005
R16874 DVDD.n19726 DVDD.n19721 4.5005
R16875 DVDD.n19738 DVDD.n19721 4.5005
R16876 DVDD.n19725 DVDD.n19721 4.5005
R16877 DVDD.n19739 DVDD.n19721 4.5005
R16878 DVDD.n19724 DVDD.n19721 4.5005
R16879 DVDD.n20572 DVDD.n19721 4.5005
R16880 DVDD.n18848 DVDD.n18838 4.5005
R16881 DVDD.n18848 DVDD.n18839 4.5005
R16882 DVDD.n18848 DVDD.n18837 4.5005
R16883 DVDD.n18848 DVDD.n18840 4.5005
R16884 DVDD.n18848 DVDD.n18836 4.5005
R16885 DVDD.n18848 DVDD.n18842 4.5005
R16886 DVDD.n18848 DVDD.n18835 4.5005
R16887 DVDD.n18848 DVDD.n18843 4.5005
R16888 DVDD.n18848 DVDD.n18834 4.5005
R16889 DVDD.n18848 DVDD.n18844 4.5005
R16890 DVDD.n18848 DVDD.n18833 4.5005
R16891 DVDD.n18848 DVDD.n18845 4.5005
R16892 DVDD.n18848 DVDD.n18846 4.5005
R16893 DVDD.n18865 DVDD.n18848 4.5005
R16894 DVDD.n20970 DVDD.n18848 4.5005
R16895 DVDD.n20969 DVDD.n18838 4.5005
R16896 DVDD.n20969 DVDD.n18839 4.5005
R16897 DVDD.n20969 DVDD.n18837 4.5005
R16898 DVDD.n20969 DVDD.n18840 4.5005
R16899 DVDD.n20969 DVDD.n18836 4.5005
R16900 DVDD.n20969 DVDD.n18842 4.5005
R16901 DVDD.n20969 DVDD.n18835 4.5005
R16902 DVDD.n20969 DVDD.n18843 4.5005
R16903 DVDD.n20969 DVDD.n18834 4.5005
R16904 DVDD.n20969 DVDD.n18844 4.5005
R16905 DVDD.n20969 DVDD.n18833 4.5005
R16906 DVDD.n20969 DVDD.n18845 4.5005
R16907 DVDD.n20969 DVDD.n18832 4.5005
R16908 DVDD.n20969 DVDD.n18846 4.5005
R16909 DVDD.n20969 DVDD.n18865 4.5005
R16910 DVDD.n20970 DVDD.n20969 4.5005
R16911 DVDD.n3656 DVDD.n3648 4.5005
R16912 DVDD.n3712 DVDD.n3648 4.5005
R16913 DVDD.n3656 DVDD.n3644 4.5005
R16914 DVDD.n3712 DVDD.n3644 4.5005
R16915 DVDD.n3656 DVDD.n3649 4.5005
R16916 DVDD.n3712 DVDD.n3649 4.5005
R16917 DVDD.n3656 DVDD.n3643 4.5005
R16918 DVDD.n3712 DVDD.n3643 4.5005
R16919 DVDD.n3656 DVDD.n3650 4.5005
R16920 DVDD.n3712 DVDD.n3650 4.5005
R16921 DVDD.n3656 DVDD.n3642 4.5005
R16922 DVDD.n3712 DVDD.n3642 4.5005
R16923 DVDD.n3663 DVDD.n3651 4.5005
R16924 DVDD.n3656 DVDD.n3651 4.5005
R16925 DVDD.n4768 DVDD.n3663 4.5005
R16926 DVDD.n4768 DVDD.n3656 4.5005
R16927 DVDD.n3665 DVDD.n3648 4.5005
R16928 DVDD.n3654 DVDD.n3648 4.5005
R16929 DVDD.n3665 DVDD.n3644 4.5005
R16930 DVDD.n3654 DVDD.n3644 4.5005
R16931 DVDD.n3665 DVDD.n3649 4.5005
R16932 DVDD.n3654 DVDD.n3649 4.5005
R16933 DVDD.n3665 DVDD.n3643 4.5005
R16934 DVDD.n3654 DVDD.n3643 4.5005
R16935 DVDD.n3665 DVDD.n3650 4.5005
R16936 DVDD.n3654 DVDD.n3650 4.5005
R16937 DVDD.n3654 DVDD.n3642 4.5005
R16938 DVDD.n3665 DVDD.n3651 4.5005
R16939 DVDD.n3654 DVDD.n3651 4.5005
R16940 DVDD.n3665 DVDD.n3641 4.5005
R16941 DVDD.n3654 DVDD.n3641 4.5005
R16942 DVDD.n4768 DVDD.n3665 4.5005
R16943 DVDD.n4768 DVDD.n3654 4.5005
R16944 DVDD.n3667 DVDD.n3648 4.5005
R16945 DVDD.n3653 DVDD.n3648 4.5005
R16946 DVDD.n3667 DVDD.n3644 4.5005
R16947 DVDD.n3653 DVDD.n3644 4.5005
R16948 DVDD.n3667 DVDD.n3649 4.5005
R16949 DVDD.n3653 DVDD.n3649 4.5005
R16950 DVDD.n3667 DVDD.n3643 4.5005
R16951 DVDD.n3653 DVDD.n3643 4.5005
R16952 DVDD.n3667 DVDD.n3650 4.5005
R16953 DVDD.n3653 DVDD.n3650 4.5005
R16954 DVDD.n3667 DVDD.n3642 4.5005
R16955 DVDD.n3653 DVDD.n3642 4.5005
R16956 DVDD.n3667 DVDD.n3651 4.5005
R16957 DVDD.n3653 DVDD.n3651 4.5005
R16958 DVDD.n3667 DVDD.n3641 4.5005
R16959 DVDD.n3653 DVDD.n3641 4.5005
R16960 DVDD.n4768 DVDD.n3667 4.5005
R16961 DVDD.n4768 DVDD.n3653 4.5005
R16962 DVDD.n4768 DVDD.n4767 4.5005
R16963 DVDD.n4767 DVDD.n3641 4.5005
R16964 DVDD.n4767 DVDD.n3651 4.5005
R16965 DVDD.n4767 DVDD.n3642 4.5005
R16966 DVDD.n4767 DVDD.n3650 4.5005
R16967 DVDD.n4767 DVDD.n3643 4.5005
R16968 DVDD.n4767 DVDD.n3649 4.5005
R16969 DVDD.n4767 DVDD.n3644 4.5005
R16970 DVDD.n4767 DVDD.n3648 4.5005
R16971 DVDD.n3652 DVDD.n3648 4.5005
R16972 DVDD.n4769 DVDD.n3648 4.5005
R16973 DVDD.n3648 DVDD.n3640 4.5005
R16974 DVDD.n3648 DVDD.n3635 4.5005
R16975 DVDD.n3652 DVDD.n3644 4.5005
R16976 DVDD.n4769 DVDD.n3644 4.5005
R16977 DVDD.n3644 DVDD.n3640 4.5005
R16978 DVDD.n3644 DVDD.n3635 4.5005
R16979 DVDD.n3652 DVDD.n3649 4.5005
R16980 DVDD.n4769 DVDD.n3649 4.5005
R16981 DVDD.n3649 DVDD.n3640 4.5005
R16982 DVDD.n3649 DVDD.n3635 4.5005
R16983 DVDD.n3652 DVDD.n3643 4.5005
R16984 DVDD.n4769 DVDD.n3643 4.5005
R16985 DVDD.n3643 DVDD.n3640 4.5005
R16986 DVDD.n3643 DVDD.n3635 4.5005
R16987 DVDD.n3652 DVDD.n3650 4.5005
R16988 DVDD.n4769 DVDD.n3650 4.5005
R16989 DVDD.n3650 DVDD.n3640 4.5005
R16990 DVDD.n3650 DVDD.n3635 4.5005
R16991 DVDD.n3652 DVDD.n3642 4.5005
R16992 DVDD.n4769 DVDD.n3642 4.5005
R16993 DVDD.n3642 DVDD.n3640 4.5005
R16994 DVDD.n3642 DVDD.n3635 4.5005
R16995 DVDD.n3652 DVDD.n3651 4.5005
R16996 DVDD.n4769 DVDD.n3651 4.5005
R16997 DVDD.n3651 DVDD.n3640 4.5005
R16998 DVDD.n3651 DVDD.n3635 4.5005
R16999 DVDD.n3652 DVDD.n3641 4.5005
R17000 DVDD.n4769 DVDD.n3641 4.5005
R17001 DVDD.n3641 DVDD.n3640 4.5005
R17002 DVDD.n3641 DVDD.n3635 4.5005
R17003 DVDD.n4768 DVDD.n3652 4.5005
R17004 DVDD.n4769 DVDD.n4768 4.5005
R17005 DVDD.n4768 DVDD.n3640 4.5005
R17006 DVDD.n4768 DVDD.n3635 4.5005
R17007 DVDD.n3487 DVDD.n3472 4.5005
R17008 DVDD.n3489 DVDD.n3472 4.5005
R17009 DVDD.n3486 DVDD.n3472 4.5005
R17010 DVDD.n3490 DVDD.n3472 4.5005
R17011 DVDD.n3485 DVDD.n3472 4.5005
R17012 DVDD.n3492 DVDD.n3472 4.5005
R17013 DVDD.n3484 DVDD.n3472 4.5005
R17014 DVDD.n3493 DVDD.n3472 4.5005
R17015 DVDD.n3483 DVDD.n3472 4.5005
R17016 DVDD.n3494 DVDD.n3472 4.5005
R17017 DVDD.n3482 DVDD.n3472 4.5005
R17018 DVDD.n15790 DVDD.n3472 4.5005
R17019 DVDD.n15793 DVDD.n3472 4.5005
R17020 DVDD.n3472 DVDD.n3419 4.5005
R17021 DVDD.n15795 DVDD.n3472 4.5005
R17022 DVDD.n3487 DVDD.n3420 4.5005
R17023 DVDD.n3489 DVDD.n3420 4.5005
R17024 DVDD.n3486 DVDD.n3420 4.5005
R17025 DVDD.n3490 DVDD.n3420 4.5005
R17026 DVDD.n3485 DVDD.n3420 4.5005
R17027 DVDD.n3492 DVDD.n3420 4.5005
R17028 DVDD.n3484 DVDD.n3420 4.5005
R17029 DVDD.n3493 DVDD.n3420 4.5005
R17030 DVDD.n3483 DVDD.n3420 4.5005
R17031 DVDD.n3494 DVDD.n3420 4.5005
R17032 DVDD.n3482 DVDD.n3420 4.5005
R17033 DVDD.n15790 DVDD.n3420 4.5005
R17034 DVDD.n3481 DVDD.n3420 4.5005
R17035 DVDD.n15793 DVDD.n3420 4.5005
R17036 DVDD.n3420 DVDD.n3419 4.5005
R17037 DVDD.n15795 DVDD.n3420 4.5005
R17038 DVDD.n15794 DVDD.n3487 4.5005
R17039 DVDD.n15794 DVDD.n3489 4.5005
R17040 DVDD.n15794 DVDD.n3486 4.5005
R17041 DVDD.n15794 DVDD.n3490 4.5005
R17042 DVDD.n15794 DVDD.n3485 4.5005
R17043 DVDD.n15794 DVDD.n3492 4.5005
R17044 DVDD.n15794 DVDD.n3484 4.5005
R17045 DVDD.n15794 DVDD.n3493 4.5005
R17046 DVDD.n15794 DVDD.n3483 4.5005
R17047 DVDD.n15794 DVDD.n3494 4.5005
R17048 DVDD.n15794 DVDD.n3482 4.5005
R17049 DVDD.n15794 DVDD.n15790 4.5005
R17050 DVDD.n15794 DVDD.n3481 4.5005
R17051 DVDD.n15794 DVDD.n15793 4.5005
R17052 DVDD.n15794 DVDD.n3419 4.5005
R17053 DVDD.n15795 DVDD.n15794 4.5005
R17054 DVDD.n16051 DVDD.n3115 4.5005
R17055 DVDD.n16051 DVDD.n3116 4.5005
R17056 DVDD.n16051 DVDD.n3114 4.5005
R17057 DVDD.n16051 DVDD.n3117 4.5005
R17058 DVDD.n16051 DVDD.n3113 4.5005
R17059 DVDD.n16051 DVDD.n3118 4.5005
R17060 DVDD.n16051 DVDD.n3112 4.5005
R17061 DVDD.n16051 DVDD.n3119 4.5005
R17062 DVDD.n16051 DVDD.n3111 4.5005
R17063 DVDD.n16051 DVDD.n3120 4.5005
R17064 DVDD.n16051 DVDD.n3110 4.5005
R17065 DVDD.n16051 DVDD.n3121 4.5005
R17066 DVDD.n16051 DVDD.n3122 4.5005
R17067 DVDD.n16061 DVDD.n16051 4.5005
R17068 DVDD.n16067 DVDD.n16051 4.5005
R17069 DVDD.n3124 DVDD.n3115 4.5005
R17070 DVDD.n3124 DVDD.n3116 4.5005
R17071 DVDD.n3124 DVDD.n3114 4.5005
R17072 DVDD.n3124 DVDD.n3117 4.5005
R17073 DVDD.n3124 DVDD.n3113 4.5005
R17074 DVDD.n3124 DVDD.n3118 4.5005
R17075 DVDD.n3124 DVDD.n3112 4.5005
R17076 DVDD.n3124 DVDD.n3119 4.5005
R17077 DVDD.n3124 DVDD.n3111 4.5005
R17078 DVDD.n3124 DVDD.n3120 4.5005
R17079 DVDD.n3124 DVDD.n3110 4.5005
R17080 DVDD.n3124 DVDD.n3121 4.5005
R17081 DVDD.n3124 DVDD.n3122 4.5005
R17082 DVDD.n16061 DVDD.n3124 4.5005
R17083 DVDD.n16067 DVDD.n3124 4.5005
R17084 DVDD.n16066 DVDD.n3115 4.5005
R17085 DVDD.n16066 DVDD.n3116 4.5005
R17086 DVDD.n16066 DVDD.n3114 4.5005
R17087 DVDD.n16066 DVDD.n3117 4.5005
R17088 DVDD.n16066 DVDD.n3113 4.5005
R17089 DVDD.n16066 DVDD.n3118 4.5005
R17090 DVDD.n16066 DVDD.n3112 4.5005
R17091 DVDD.n16066 DVDD.n3119 4.5005
R17092 DVDD.n16066 DVDD.n3111 4.5005
R17093 DVDD.n16066 DVDD.n3120 4.5005
R17094 DVDD.n16066 DVDD.n3110 4.5005
R17095 DVDD.n16066 DVDD.n3121 4.5005
R17096 DVDD.n16066 DVDD.n3122 4.5005
R17097 DVDD.n16066 DVDD.n16061 4.5005
R17098 DVDD.n16067 DVDD.n16066 4.5005
R17099 DVDD.n9947 DVDD.n9763 4.5005
R17100 DVDD.n9947 DVDD.n9764 4.5005
R17101 DVDD.n9947 DVDD.n9762 4.5005
R17102 DVDD.n9947 DVDD.n9765 4.5005
R17103 DVDD.n9947 DVDD.n9761 4.5005
R17104 DVDD.n9947 DVDD.n9767 4.5005
R17105 DVDD.n9947 DVDD.n9760 4.5005
R17106 DVDD.n9947 DVDD.n9768 4.5005
R17107 DVDD.n9947 DVDD.n9759 4.5005
R17108 DVDD.n9947 DVDD.n9769 4.5005
R17109 DVDD.n9947 DVDD.n9758 4.5005
R17110 DVDD.n9947 DVDD.n9770 4.5005
R17111 DVDD.n9947 DVDD.n9939 4.5005
R17112 DVDD.n9947 DVDD.n9772 4.5005
R17113 DVDD.n9948 DVDD.n9947 4.5005
R17114 DVDD.n9774 DVDD.n9763 4.5005
R17115 DVDD.n9774 DVDD.n9764 4.5005
R17116 DVDD.n9774 DVDD.n9762 4.5005
R17117 DVDD.n9774 DVDD.n9765 4.5005
R17118 DVDD.n9774 DVDD.n9761 4.5005
R17119 DVDD.n9774 DVDD.n9767 4.5005
R17120 DVDD.n9774 DVDD.n9760 4.5005
R17121 DVDD.n9774 DVDD.n9768 4.5005
R17122 DVDD.n9774 DVDD.n9759 4.5005
R17123 DVDD.n9774 DVDD.n9769 4.5005
R17124 DVDD.n9774 DVDD.n9758 4.5005
R17125 DVDD.n9774 DVDD.n9770 4.5005
R17126 DVDD.n9774 DVDD.n9772 4.5005
R17127 DVDD.n9774 DVDD.n9757 4.5005
R17128 DVDD.n9948 DVDD.n9774 4.5005
R17129 DVDD.n9949 DVDD.n9763 4.5005
R17130 DVDD.n9949 DVDD.n9764 4.5005
R17131 DVDD.n9949 DVDD.n9762 4.5005
R17132 DVDD.n9949 DVDD.n9765 4.5005
R17133 DVDD.n9949 DVDD.n9761 4.5005
R17134 DVDD.n9949 DVDD.n9767 4.5005
R17135 DVDD.n9949 DVDD.n9760 4.5005
R17136 DVDD.n9949 DVDD.n9768 4.5005
R17137 DVDD.n9949 DVDD.n9759 4.5005
R17138 DVDD.n9949 DVDD.n9769 4.5005
R17139 DVDD.n9949 DVDD.n9758 4.5005
R17140 DVDD.n9949 DVDD.n9770 4.5005
R17141 DVDD.n9949 DVDD.n9772 4.5005
R17142 DVDD.n9949 DVDD.n9757 4.5005
R17143 DVDD.n9949 DVDD.n9948 4.5005
R17144 DVDD.n21214 DVDD.n21213 4.5005
R17145 DVDD.n21214 DVDD.n18684 4.5005
R17146 DVDD.n21214 DVDD.n18683 4.5005
R17147 DVDD.n21214 DVDD.n18682 4.5005
R17148 DVDD.n21214 DVDD.n18681 4.5005
R17149 DVDD.n21214 DVDD.n18679 4.5005
R17150 DVDD.n21214 DVDD.n18678 4.5005
R17151 DVDD.n21214 DVDD.n18677 4.5005
R17152 DVDD.n21214 DVDD.n18676 4.5005
R17153 DVDD.n21214 DVDD.n18675 4.5005
R17154 DVDD.n21214 DVDD.n18674 4.5005
R17155 DVDD.n21213 DVDD.n18690 4.5005
R17156 DVDD.n18690 DVDD.n18684 4.5005
R17157 DVDD.n18690 DVDD.n18683 4.5005
R17158 DVDD.n18690 DVDD.n18682 4.5005
R17159 DVDD.n18690 DVDD.n18681 4.5005
R17160 DVDD.n18700 DVDD.n18690 4.5005
R17161 DVDD.n21211 DVDD.n18690 4.5005
R17162 DVDD.n18690 DVDD.n18679 4.5005
R17163 DVDD.n18690 DVDD.n18678 4.5005
R17164 DVDD.n18690 DVDD.n18677 4.5005
R17165 DVDD.n18690 DVDD.n18676 4.5005
R17166 DVDD.n18690 DVDD.n18675 4.5005
R17167 DVDD.n18690 DVDD.n18674 4.5005
R17168 DVDD.n18701 DVDD.n18690 4.5005
R17169 DVDD.n21213 DVDD.n18693 4.5005
R17170 DVDD.n18693 DVDD.n18684 4.5005
R17171 DVDD.n18693 DVDD.n18683 4.5005
R17172 DVDD.n18693 DVDD.n18682 4.5005
R17173 DVDD.n18693 DVDD.n18681 4.5005
R17174 DVDD.n18700 DVDD.n18693 4.5005
R17175 DVDD.n21211 DVDD.n18693 4.5005
R17176 DVDD.n18693 DVDD.n18679 4.5005
R17177 DVDD.n18693 DVDD.n18678 4.5005
R17178 DVDD.n18693 DVDD.n18677 4.5005
R17179 DVDD.n18693 DVDD.n18676 4.5005
R17180 DVDD.n18693 DVDD.n18675 4.5005
R17181 DVDD.n18701 DVDD.n18693 4.5005
R17182 DVDD.n18702 DVDD.n18693 4.5005
R17183 DVDD.n21213 DVDD.n18689 4.5005
R17184 DVDD.n18689 DVDD.n18684 4.5005
R17185 DVDD.n18689 DVDD.n18683 4.5005
R17186 DVDD.n18689 DVDD.n18682 4.5005
R17187 DVDD.n18689 DVDD.n18681 4.5005
R17188 DVDD.n18700 DVDD.n18689 4.5005
R17189 DVDD.n21211 DVDD.n18689 4.5005
R17190 DVDD.n18689 DVDD.n18679 4.5005
R17191 DVDD.n18689 DVDD.n18678 4.5005
R17192 DVDD.n18689 DVDD.n18677 4.5005
R17193 DVDD.n18689 DVDD.n18676 4.5005
R17194 DVDD.n18689 DVDD.n18675 4.5005
R17195 DVDD.n18701 DVDD.n18689 4.5005
R17196 DVDD.n18702 DVDD.n18689 4.5005
R17197 DVDD.n21213 DVDD.n18694 4.5005
R17198 DVDD.n18694 DVDD.n18684 4.5005
R17199 DVDD.n18694 DVDD.n18683 4.5005
R17200 DVDD.n18694 DVDD.n18682 4.5005
R17201 DVDD.n18694 DVDD.n18681 4.5005
R17202 DVDD.n18700 DVDD.n18694 4.5005
R17203 DVDD.n21211 DVDD.n18694 4.5005
R17204 DVDD.n18694 DVDD.n18679 4.5005
R17205 DVDD.n18694 DVDD.n18678 4.5005
R17206 DVDD.n18694 DVDD.n18677 4.5005
R17207 DVDD.n18694 DVDD.n18676 4.5005
R17208 DVDD.n18694 DVDD.n18675 4.5005
R17209 DVDD.n18694 DVDD.n18674 4.5005
R17210 DVDD.n18701 DVDD.n18694 4.5005
R17211 DVDD.n18702 DVDD.n18694 4.5005
R17212 DVDD.n21213 DVDD.n18688 4.5005
R17213 DVDD.n18688 DVDD.n18684 4.5005
R17214 DVDD.n18688 DVDD.n18683 4.5005
R17215 DVDD.n18688 DVDD.n18682 4.5005
R17216 DVDD.n18688 DVDD.n18681 4.5005
R17217 DVDD.n18700 DVDD.n18688 4.5005
R17218 DVDD.n21211 DVDD.n18688 4.5005
R17219 DVDD.n18688 DVDD.n18679 4.5005
R17220 DVDD.n18688 DVDD.n18678 4.5005
R17221 DVDD.n18688 DVDD.n18677 4.5005
R17222 DVDD.n18688 DVDD.n18676 4.5005
R17223 DVDD.n18688 DVDD.n18675 4.5005
R17224 DVDD.n18688 DVDD.n18674 4.5005
R17225 DVDD.n18701 DVDD.n18688 4.5005
R17226 DVDD.n18702 DVDD.n18688 4.5005
R17227 DVDD.n21213 DVDD.n18696 4.5005
R17228 DVDD.n18696 DVDD.n18684 4.5005
R17229 DVDD.n18696 DVDD.n18683 4.5005
R17230 DVDD.n18696 DVDD.n18682 4.5005
R17231 DVDD.n18696 DVDD.n18681 4.5005
R17232 DVDD.n18700 DVDD.n18696 4.5005
R17233 DVDD.n21211 DVDD.n18696 4.5005
R17234 DVDD.n18696 DVDD.n18679 4.5005
R17235 DVDD.n18696 DVDD.n18678 4.5005
R17236 DVDD.n18696 DVDD.n18677 4.5005
R17237 DVDD.n18696 DVDD.n18676 4.5005
R17238 DVDD.n18696 DVDD.n18675 4.5005
R17239 DVDD.n18701 DVDD.n18696 4.5005
R17240 DVDD.n18702 DVDD.n18696 4.5005
R17241 DVDD.n21213 DVDD.n18687 4.5005
R17242 DVDD.n18687 DVDD.n18684 4.5005
R17243 DVDD.n18687 DVDD.n18683 4.5005
R17244 DVDD.n18687 DVDD.n18682 4.5005
R17245 DVDD.n18687 DVDD.n18681 4.5005
R17246 DVDD.n18700 DVDD.n18687 4.5005
R17247 DVDD.n21211 DVDD.n18687 4.5005
R17248 DVDD.n18687 DVDD.n18679 4.5005
R17249 DVDD.n18687 DVDD.n18678 4.5005
R17250 DVDD.n18687 DVDD.n18677 4.5005
R17251 DVDD.n18687 DVDD.n18676 4.5005
R17252 DVDD.n18687 DVDD.n18675 4.5005
R17253 DVDD.n18701 DVDD.n18687 4.5005
R17254 DVDD.n18702 DVDD.n18687 4.5005
R17255 DVDD.n21213 DVDD.n18698 4.5005
R17256 DVDD.n18698 DVDD.n18684 4.5005
R17257 DVDD.n18698 DVDD.n18683 4.5005
R17258 DVDD.n18698 DVDD.n18682 4.5005
R17259 DVDD.n18698 DVDD.n18681 4.5005
R17260 DVDD.n18700 DVDD.n18698 4.5005
R17261 DVDD.n21211 DVDD.n18698 4.5005
R17262 DVDD.n18698 DVDD.n18679 4.5005
R17263 DVDD.n18698 DVDD.n18678 4.5005
R17264 DVDD.n18698 DVDD.n18677 4.5005
R17265 DVDD.n18698 DVDD.n18676 4.5005
R17266 DVDD.n18698 DVDD.n18675 4.5005
R17267 DVDD.n18701 DVDD.n18698 4.5005
R17268 DVDD.n18702 DVDD.n18698 4.5005
R17269 DVDD.n21213 DVDD.n18686 4.5005
R17270 DVDD.n18686 DVDD.n18684 4.5005
R17271 DVDD.n18686 DVDD.n18683 4.5005
R17272 DVDD.n18686 DVDD.n18682 4.5005
R17273 DVDD.n18686 DVDD.n18681 4.5005
R17274 DVDD.n18700 DVDD.n18686 4.5005
R17275 DVDD.n21211 DVDD.n18686 4.5005
R17276 DVDD.n18686 DVDD.n18679 4.5005
R17277 DVDD.n18686 DVDD.n18678 4.5005
R17278 DVDD.n18686 DVDD.n18677 4.5005
R17279 DVDD.n18686 DVDD.n18676 4.5005
R17280 DVDD.n18686 DVDD.n18675 4.5005
R17281 DVDD.n18701 DVDD.n18686 4.5005
R17282 DVDD.n18708 DVDD.n18686 4.5005
R17283 DVDD.n18702 DVDD.n18686 4.5005
R17284 DVDD.n21212 DVDD.n18702 4.5005
R17285 DVDD.n21212 DVDD.n18708 4.5005
R17286 DVDD.n21212 DVDD.n18701 4.5005
R17287 DVDD.n21212 DVDD.n18674 4.5005
R17288 DVDD.n21212 DVDD.n18675 4.5005
R17289 DVDD.n21212 DVDD.n18676 4.5005
R17290 DVDD.n21212 DVDD.n18677 4.5005
R17291 DVDD.n21212 DVDD.n18678 4.5005
R17292 DVDD.n21212 DVDD.n18679 4.5005
R17293 DVDD.n21212 DVDD.n21211 4.5005
R17294 DVDD.n21212 DVDD.n18700 4.5005
R17295 DVDD.n21212 DVDD.n18681 4.5005
R17296 DVDD.n21212 DVDD.n18682 4.5005
R17297 DVDD.n21212 DVDD.n18683 4.5005
R17298 DVDD.n21212 DVDD.n18684 4.5005
R17299 DVDD.n21213 DVDD.n21212 4.5005
R17300 DVDD.n21186 DVDD.n18730 4.5005
R17301 DVDD.n18736 DVDD.n18730 4.5005
R17302 DVDD.n21184 DVDD.n18730 4.5005
R17303 DVDD.n18738 DVDD.n18730 4.5005
R17304 DVDD.n21097 DVDD.n18730 4.5005
R17305 DVDD.n18739 DVDD.n18730 4.5005
R17306 DVDD.n21096 DVDD.n18730 4.5005
R17307 DVDD.n18740 DVDD.n18730 4.5005
R17308 DVDD.n21095 DVDD.n18730 4.5005
R17309 DVDD.n18742 DVDD.n18730 4.5005
R17310 DVDD.n18743 DVDD.n18730 4.5005
R17311 DVDD.n21186 DVDD.n18728 4.5005
R17312 DVDD.n18736 DVDD.n18728 4.5005
R17313 DVDD.n21184 DVDD.n18728 4.5005
R17314 DVDD.n18737 DVDD.n18728 4.5005
R17315 DVDD.n21099 DVDD.n18728 4.5005
R17316 DVDD.n18738 DVDD.n18728 4.5005
R17317 DVDD.n21097 DVDD.n18728 4.5005
R17318 DVDD.n18739 DVDD.n18728 4.5005
R17319 DVDD.n21096 DVDD.n18728 4.5005
R17320 DVDD.n18740 DVDD.n18728 4.5005
R17321 DVDD.n21095 DVDD.n18728 4.5005
R17322 DVDD.n18741 DVDD.n18728 4.5005
R17323 DVDD.n18742 DVDD.n18728 4.5005
R17324 DVDD.n18743 DVDD.n18728 4.5005
R17325 DVDD.n21186 DVDD.n18731 4.5005
R17326 DVDD.n18736 DVDD.n18731 4.5005
R17327 DVDD.n21184 DVDD.n18731 4.5005
R17328 DVDD.n18737 DVDD.n18731 4.5005
R17329 DVDD.n21099 DVDD.n18731 4.5005
R17330 DVDD.n18738 DVDD.n18731 4.5005
R17331 DVDD.n21097 DVDD.n18731 4.5005
R17332 DVDD.n18739 DVDD.n18731 4.5005
R17333 DVDD.n21096 DVDD.n18731 4.5005
R17334 DVDD.n18740 DVDD.n18731 4.5005
R17335 DVDD.n21095 DVDD.n18731 4.5005
R17336 DVDD.n18741 DVDD.n18731 4.5005
R17337 DVDD.n18742 DVDD.n18731 4.5005
R17338 DVDD.n18743 DVDD.n18731 4.5005
R17339 DVDD.n21186 DVDD.n18727 4.5005
R17340 DVDD.n18736 DVDD.n18727 4.5005
R17341 DVDD.n21184 DVDD.n18727 4.5005
R17342 DVDD.n18737 DVDD.n18727 4.5005
R17343 DVDD.n21099 DVDD.n18727 4.5005
R17344 DVDD.n18738 DVDD.n18727 4.5005
R17345 DVDD.n21097 DVDD.n18727 4.5005
R17346 DVDD.n18739 DVDD.n18727 4.5005
R17347 DVDD.n21096 DVDD.n18727 4.5005
R17348 DVDD.n18740 DVDD.n18727 4.5005
R17349 DVDD.n21095 DVDD.n18727 4.5005
R17350 DVDD.n18741 DVDD.n18727 4.5005
R17351 DVDD.n18742 DVDD.n18727 4.5005
R17352 DVDD.n18743 DVDD.n18727 4.5005
R17353 DVDD.n21186 DVDD.n18732 4.5005
R17354 DVDD.n18736 DVDD.n18732 4.5005
R17355 DVDD.n21184 DVDD.n18732 4.5005
R17356 DVDD.n18737 DVDD.n18732 4.5005
R17357 DVDD.n21099 DVDD.n18732 4.5005
R17358 DVDD.n18738 DVDD.n18732 4.5005
R17359 DVDD.n21097 DVDD.n18732 4.5005
R17360 DVDD.n18739 DVDD.n18732 4.5005
R17361 DVDD.n21096 DVDD.n18732 4.5005
R17362 DVDD.n18740 DVDD.n18732 4.5005
R17363 DVDD.n21095 DVDD.n18732 4.5005
R17364 DVDD.n18741 DVDD.n18732 4.5005
R17365 DVDD.n18742 DVDD.n18732 4.5005
R17366 DVDD.n21088 DVDD.n18732 4.5005
R17367 DVDD.n18743 DVDD.n18732 4.5005
R17368 DVDD.n21186 DVDD.n18726 4.5005
R17369 DVDD.n18736 DVDD.n18726 4.5005
R17370 DVDD.n21184 DVDD.n18726 4.5005
R17371 DVDD.n18737 DVDD.n18726 4.5005
R17372 DVDD.n21099 DVDD.n18726 4.5005
R17373 DVDD.n18738 DVDD.n18726 4.5005
R17374 DVDD.n21097 DVDD.n18726 4.5005
R17375 DVDD.n18739 DVDD.n18726 4.5005
R17376 DVDD.n21096 DVDD.n18726 4.5005
R17377 DVDD.n18740 DVDD.n18726 4.5005
R17378 DVDD.n21095 DVDD.n18726 4.5005
R17379 DVDD.n18741 DVDD.n18726 4.5005
R17380 DVDD.n21094 DVDD.n18726 4.5005
R17381 DVDD.n18742 DVDD.n18726 4.5005
R17382 DVDD.n18743 DVDD.n18726 4.5005
R17383 DVDD.n21186 DVDD.n18733 4.5005
R17384 DVDD.n18736 DVDD.n18733 4.5005
R17385 DVDD.n21184 DVDD.n18733 4.5005
R17386 DVDD.n18737 DVDD.n18733 4.5005
R17387 DVDD.n21099 DVDD.n18733 4.5005
R17388 DVDD.n18738 DVDD.n18733 4.5005
R17389 DVDD.n21097 DVDD.n18733 4.5005
R17390 DVDD.n18739 DVDD.n18733 4.5005
R17391 DVDD.n21096 DVDD.n18733 4.5005
R17392 DVDD.n18740 DVDD.n18733 4.5005
R17393 DVDD.n21095 DVDD.n18733 4.5005
R17394 DVDD.n18741 DVDD.n18733 4.5005
R17395 DVDD.n18742 DVDD.n18733 4.5005
R17396 DVDD.n18743 DVDD.n18733 4.5005
R17397 DVDD.n21186 DVDD.n18725 4.5005
R17398 DVDD.n18736 DVDD.n18725 4.5005
R17399 DVDD.n21184 DVDD.n18725 4.5005
R17400 DVDD.n18737 DVDD.n18725 4.5005
R17401 DVDD.n21099 DVDD.n18725 4.5005
R17402 DVDD.n18738 DVDD.n18725 4.5005
R17403 DVDD.n21097 DVDD.n18725 4.5005
R17404 DVDD.n18739 DVDD.n18725 4.5005
R17405 DVDD.n21096 DVDD.n18725 4.5005
R17406 DVDD.n18740 DVDD.n18725 4.5005
R17407 DVDD.n21095 DVDD.n18725 4.5005
R17408 DVDD.n18741 DVDD.n18725 4.5005
R17409 DVDD.n18742 DVDD.n18725 4.5005
R17410 DVDD.n18743 DVDD.n18725 4.5005
R17411 DVDD.n21186 DVDD.n18734 4.5005
R17412 DVDD.n18736 DVDD.n18734 4.5005
R17413 DVDD.n21184 DVDD.n18734 4.5005
R17414 DVDD.n18737 DVDD.n18734 4.5005
R17415 DVDD.n21099 DVDD.n18734 4.5005
R17416 DVDD.n18738 DVDD.n18734 4.5005
R17417 DVDD.n21097 DVDD.n18734 4.5005
R17418 DVDD.n18739 DVDD.n18734 4.5005
R17419 DVDD.n21096 DVDD.n18734 4.5005
R17420 DVDD.n18740 DVDD.n18734 4.5005
R17421 DVDD.n21095 DVDD.n18734 4.5005
R17422 DVDD.n18741 DVDD.n18734 4.5005
R17423 DVDD.n18742 DVDD.n18734 4.5005
R17424 DVDD.n18743 DVDD.n18734 4.5005
R17425 DVDD.n21186 DVDD.n18724 4.5005
R17426 DVDD.n18736 DVDD.n18724 4.5005
R17427 DVDD.n21184 DVDD.n18724 4.5005
R17428 DVDD.n18737 DVDD.n18724 4.5005
R17429 DVDD.n21099 DVDD.n18724 4.5005
R17430 DVDD.n18738 DVDD.n18724 4.5005
R17431 DVDD.n21097 DVDD.n18724 4.5005
R17432 DVDD.n18739 DVDD.n18724 4.5005
R17433 DVDD.n21096 DVDD.n18724 4.5005
R17434 DVDD.n18740 DVDD.n18724 4.5005
R17435 DVDD.n21095 DVDD.n18724 4.5005
R17436 DVDD.n18741 DVDD.n18724 4.5005
R17437 DVDD.n18742 DVDD.n18724 4.5005
R17438 DVDD.n21088 DVDD.n18724 4.5005
R17439 DVDD.n18743 DVDD.n18724 4.5005
R17440 DVDD.n21185 DVDD.n18743 4.5005
R17441 DVDD.n21185 DVDD.n21088 4.5005
R17442 DVDD.n21185 DVDD.n18742 4.5005
R17443 DVDD.n21185 DVDD.n21094 4.5005
R17444 DVDD.n21185 DVDD.n18741 4.5005
R17445 DVDD.n21185 DVDD.n21095 4.5005
R17446 DVDD.n21185 DVDD.n18740 4.5005
R17447 DVDD.n21185 DVDD.n21096 4.5005
R17448 DVDD.n21185 DVDD.n18739 4.5005
R17449 DVDD.n21185 DVDD.n21097 4.5005
R17450 DVDD.n21185 DVDD.n18738 4.5005
R17451 DVDD.n21185 DVDD.n21099 4.5005
R17452 DVDD.n21185 DVDD.n18737 4.5005
R17453 DVDD.n21185 DVDD.n21184 4.5005
R17454 DVDD.n21185 DVDD.n18736 4.5005
R17455 DVDD.n21186 DVDD.n21185 4.5005
R17456 DVDD.n22251 DVDD.n22244 4.5005
R17457 DVDD.n22244 DVDD.n98 4.5005
R17458 DVDD.n22244 DVDD.n111 4.5005
R17459 DVDD.n22244 DVDD.n100 4.5005
R17460 DVDD.n22244 DVDD.n109 4.5005
R17461 DVDD.n22244 DVDD.n101 4.5005
R17462 DVDD.n22244 DVDD.n108 4.5005
R17463 DVDD.n22244 DVDD.n102 4.5005
R17464 DVDD.n22244 DVDD.n107 4.5005
R17465 DVDD.n22244 DVDD.n89 4.5005
R17466 DVDD.n22244 DVDD.n85 4.5005
R17467 DVDD.n22251 DVDD.n117 4.5005
R17468 DVDD.n117 DVDD.n98 4.5005
R17469 DVDD.n117 DVDD.n111 4.5005
R17470 DVDD.n117 DVDD.n99 4.5005
R17471 DVDD.n117 DVDD.n110 4.5005
R17472 DVDD.n117 DVDD.n100 4.5005
R17473 DVDD.n117 DVDD.n109 4.5005
R17474 DVDD.n117 DVDD.n101 4.5005
R17475 DVDD.n117 DVDD.n108 4.5005
R17476 DVDD.n117 DVDD.n102 4.5005
R17477 DVDD.n117 DVDD.n107 4.5005
R17478 DVDD.n117 DVDD.n103 4.5005
R17479 DVDD.n117 DVDD.n89 4.5005
R17480 DVDD.n117 DVDD.n85 4.5005
R17481 DVDD.n22251 DVDD.n22246 4.5005
R17482 DVDD.n22246 DVDD.n98 4.5005
R17483 DVDD.n22246 DVDD.n111 4.5005
R17484 DVDD.n22246 DVDD.n99 4.5005
R17485 DVDD.n22246 DVDD.n110 4.5005
R17486 DVDD.n22246 DVDD.n100 4.5005
R17487 DVDD.n22246 DVDD.n109 4.5005
R17488 DVDD.n22246 DVDD.n101 4.5005
R17489 DVDD.n22246 DVDD.n108 4.5005
R17490 DVDD.n22246 DVDD.n102 4.5005
R17491 DVDD.n22246 DVDD.n107 4.5005
R17492 DVDD.n22246 DVDD.n103 4.5005
R17493 DVDD.n22246 DVDD.n89 4.5005
R17494 DVDD.n22246 DVDD.n85 4.5005
R17495 DVDD.n22251 DVDD.n116 4.5005
R17496 DVDD.n116 DVDD.n98 4.5005
R17497 DVDD.n116 DVDD.n111 4.5005
R17498 DVDD.n116 DVDD.n99 4.5005
R17499 DVDD.n116 DVDD.n110 4.5005
R17500 DVDD.n116 DVDD.n100 4.5005
R17501 DVDD.n116 DVDD.n109 4.5005
R17502 DVDD.n116 DVDD.n101 4.5005
R17503 DVDD.n116 DVDD.n108 4.5005
R17504 DVDD.n116 DVDD.n102 4.5005
R17505 DVDD.n116 DVDD.n107 4.5005
R17506 DVDD.n116 DVDD.n103 4.5005
R17507 DVDD.n116 DVDD.n89 4.5005
R17508 DVDD.n116 DVDD.n85 4.5005
R17509 DVDD.n22251 DVDD.n96 4.5005
R17510 DVDD.n98 DVDD.n96 4.5005
R17511 DVDD.n111 DVDD.n96 4.5005
R17512 DVDD.n99 DVDD.n96 4.5005
R17513 DVDD.n110 DVDD.n96 4.5005
R17514 DVDD.n100 DVDD.n96 4.5005
R17515 DVDD.n109 DVDD.n96 4.5005
R17516 DVDD.n101 DVDD.n96 4.5005
R17517 DVDD.n108 DVDD.n96 4.5005
R17518 DVDD.n102 DVDD.n96 4.5005
R17519 DVDD.n107 DVDD.n96 4.5005
R17520 DVDD.n103 DVDD.n96 4.5005
R17521 DVDD.n96 DVDD.n89 4.5005
R17522 DVDD.n22253 DVDD.n96 4.5005
R17523 DVDD.n96 DVDD.n85 4.5005
R17524 DVDD.n22251 DVDD.n114 4.5005
R17525 DVDD.n114 DVDD.n98 4.5005
R17526 DVDD.n114 DVDD.n111 4.5005
R17527 DVDD.n114 DVDD.n99 4.5005
R17528 DVDD.n114 DVDD.n110 4.5005
R17529 DVDD.n114 DVDD.n100 4.5005
R17530 DVDD.n114 DVDD.n109 4.5005
R17531 DVDD.n114 DVDD.n101 4.5005
R17532 DVDD.n114 DVDD.n108 4.5005
R17533 DVDD.n114 DVDD.n102 4.5005
R17534 DVDD.n114 DVDD.n107 4.5005
R17535 DVDD.n114 DVDD.n103 4.5005
R17536 DVDD.n114 DVDD.n106 4.5005
R17537 DVDD.n114 DVDD.n89 4.5005
R17538 DVDD.n114 DVDD.n85 4.5005
R17539 DVDD.n22251 DVDD.n22248 4.5005
R17540 DVDD.n22248 DVDD.n98 4.5005
R17541 DVDD.n22248 DVDD.n111 4.5005
R17542 DVDD.n22248 DVDD.n99 4.5005
R17543 DVDD.n22248 DVDD.n110 4.5005
R17544 DVDD.n22248 DVDD.n100 4.5005
R17545 DVDD.n22248 DVDD.n109 4.5005
R17546 DVDD.n22248 DVDD.n101 4.5005
R17547 DVDD.n22248 DVDD.n108 4.5005
R17548 DVDD.n22248 DVDD.n102 4.5005
R17549 DVDD.n22248 DVDD.n107 4.5005
R17550 DVDD.n22248 DVDD.n103 4.5005
R17551 DVDD.n22248 DVDD.n89 4.5005
R17552 DVDD.n22248 DVDD.n85 4.5005
R17553 DVDD.n22251 DVDD.n113 4.5005
R17554 DVDD.n113 DVDD.n98 4.5005
R17555 DVDD.n113 DVDD.n111 4.5005
R17556 DVDD.n113 DVDD.n99 4.5005
R17557 DVDD.n113 DVDD.n110 4.5005
R17558 DVDD.n113 DVDD.n100 4.5005
R17559 DVDD.n113 DVDD.n109 4.5005
R17560 DVDD.n113 DVDD.n101 4.5005
R17561 DVDD.n113 DVDD.n108 4.5005
R17562 DVDD.n113 DVDD.n102 4.5005
R17563 DVDD.n113 DVDD.n107 4.5005
R17564 DVDD.n113 DVDD.n103 4.5005
R17565 DVDD.n113 DVDD.n89 4.5005
R17566 DVDD.n113 DVDD.n85 4.5005
R17567 DVDD.n22251 DVDD.n22250 4.5005
R17568 DVDD.n22250 DVDD.n98 4.5005
R17569 DVDD.n22250 DVDD.n111 4.5005
R17570 DVDD.n22250 DVDD.n99 4.5005
R17571 DVDD.n22250 DVDD.n110 4.5005
R17572 DVDD.n22250 DVDD.n100 4.5005
R17573 DVDD.n22250 DVDD.n109 4.5005
R17574 DVDD.n22250 DVDD.n101 4.5005
R17575 DVDD.n22250 DVDD.n108 4.5005
R17576 DVDD.n22250 DVDD.n102 4.5005
R17577 DVDD.n22250 DVDD.n107 4.5005
R17578 DVDD.n22250 DVDD.n103 4.5005
R17579 DVDD.n22250 DVDD.n89 4.5005
R17580 DVDD.n22250 DVDD.n85 4.5005
R17581 DVDD.n22251 DVDD.n90 4.5005
R17582 DVDD.n98 DVDD.n90 4.5005
R17583 DVDD.n111 DVDD.n90 4.5005
R17584 DVDD.n99 DVDD.n90 4.5005
R17585 DVDD.n110 DVDD.n90 4.5005
R17586 DVDD.n100 DVDD.n90 4.5005
R17587 DVDD.n109 DVDD.n90 4.5005
R17588 DVDD.n101 DVDD.n90 4.5005
R17589 DVDD.n108 DVDD.n90 4.5005
R17590 DVDD.n102 DVDD.n90 4.5005
R17591 DVDD.n107 DVDD.n90 4.5005
R17592 DVDD.n103 DVDD.n90 4.5005
R17593 DVDD.n90 DVDD.n89 4.5005
R17594 DVDD.n22253 DVDD.n90 4.5005
R17595 DVDD.n90 DVDD.n85 4.5005
R17596 DVDD.n22252 DVDD.n85 4.5005
R17597 DVDD.n22253 DVDD.n22252 4.5005
R17598 DVDD.n22252 DVDD.n89 4.5005
R17599 DVDD.n22252 DVDD.n106 4.5005
R17600 DVDD.n22252 DVDD.n103 4.5005
R17601 DVDD.n22252 DVDD.n107 4.5005
R17602 DVDD.n22252 DVDD.n102 4.5005
R17603 DVDD.n22252 DVDD.n108 4.5005
R17604 DVDD.n22252 DVDD.n101 4.5005
R17605 DVDD.n22252 DVDD.n109 4.5005
R17606 DVDD.n22252 DVDD.n100 4.5005
R17607 DVDD.n22252 DVDD.n110 4.5005
R17608 DVDD.n22252 DVDD.n99 4.5005
R17609 DVDD.n22252 DVDD.n111 4.5005
R17610 DVDD.n22252 DVDD.n98 4.5005
R17611 DVDD.n22252 DVDD.n22251 4.5005
R17612 DVDD.n22297 DVDD.n49 4.5005
R17613 DVDD.n59 DVDD.n49 4.5005
R17614 DVDD.n76 DVDD.n49 4.5005
R17615 DVDD.n60 DVDD.n49 4.5005
R17616 DVDD.n75 DVDD.n49 4.5005
R17617 DVDD.n61 DVDD.n49 4.5005
R17618 DVDD.n74 DVDD.n49 4.5005
R17619 DVDD.n63 DVDD.n49 4.5005
R17620 DVDD.n71 DVDD.n49 4.5005
R17621 DVDD.n65 DVDD.n49 4.5005
R17622 DVDD.n22299 DVDD.n49 4.5005
R17623 DVDD.n22297 DVDD.n47 4.5005
R17624 DVDD.n58 DVDD.n47 4.5005
R17625 DVDD.n78 DVDD.n47 4.5005
R17626 DVDD.n59 DVDD.n47 4.5005
R17627 DVDD.n76 DVDD.n47 4.5005
R17628 DVDD.n60 DVDD.n47 4.5005
R17629 DVDD.n75 DVDD.n47 4.5005
R17630 DVDD.n61 DVDD.n47 4.5005
R17631 DVDD.n74 DVDD.n47 4.5005
R17632 DVDD.n62 DVDD.n47 4.5005
R17633 DVDD.n73 DVDD.n47 4.5005
R17634 DVDD.n63 DVDD.n47 4.5005
R17635 DVDD.n65 DVDD.n47 4.5005
R17636 DVDD.n22299 DVDD.n47 4.5005
R17637 DVDD.n22297 DVDD.n51 4.5005
R17638 DVDD.n58 DVDD.n51 4.5005
R17639 DVDD.n78 DVDD.n51 4.5005
R17640 DVDD.n59 DVDD.n51 4.5005
R17641 DVDD.n76 DVDD.n51 4.5005
R17642 DVDD.n60 DVDD.n51 4.5005
R17643 DVDD.n75 DVDD.n51 4.5005
R17644 DVDD.n61 DVDD.n51 4.5005
R17645 DVDD.n74 DVDD.n51 4.5005
R17646 DVDD.n62 DVDD.n51 4.5005
R17647 DVDD.n73 DVDD.n51 4.5005
R17648 DVDD.n63 DVDD.n51 4.5005
R17649 DVDD.n65 DVDD.n51 4.5005
R17650 DVDD.n22299 DVDD.n51 4.5005
R17651 DVDD.n22297 DVDD.n46 4.5005
R17652 DVDD.n58 DVDD.n46 4.5005
R17653 DVDD.n78 DVDD.n46 4.5005
R17654 DVDD.n59 DVDD.n46 4.5005
R17655 DVDD.n76 DVDD.n46 4.5005
R17656 DVDD.n60 DVDD.n46 4.5005
R17657 DVDD.n75 DVDD.n46 4.5005
R17658 DVDD.n61 DVDD.n46 4.5005
R17659 DVDD.n74 DVDD.n46 4.5005
R17660 DVDD.n62 DVDD.n46 4.5005
R17661 DVDD.n73 DVDD.n46 4.5005
R17662 DVDD.n63 DVDD.n46 4.5005
R17663 DVDD.n65 DVDD.n46 4.5005
R17664 DVDD.n22299 DVDD.n46 4.5005
R17665 DVDD.n22297 DVDD.n52 4.5005
R17666 DVDD.n58 DVDD.n52 4.5005
R17667 DVDD.n78 DVDD.n52 4.5005
R17668 DVDD.n59 DVDD.n52 4.5005
R17669 DVDD.n76 DVDD.n52 4.5005
R17670 DVDD.n60 DVDD.n52 4.5005
R17671 DVDD.n75 DVDD.n52 4.5005
R17672 DVDD.n61 DVDD.n52 4.5005
R17673 DVDD.n74 DVDD.n52 4.5005
R17674 DVDD.n62 DVDD.n52 4.5005
R17675 DVDD.n73 DVDD.n52 4.5005
R17676 DVDD.n63 DVDD.n52 4.5005
R17677 DVDD.n65 DVDD.n52 4.5005
R17678 DVDD.n52 DVDD.n42 4.5005
R17679 DVDD.n22299 DVDD.n52 4.5005
R17680 DVDD.n22297 DVDD.n45 4.5005
R17681 DVDD.n58 DVDD.n45 4.5005
R17682 DVDD.n78 DVDD.n45 4.5005
R17683 DVDD.n59 DVDD.n45 4.5005
R17684 DVDD.n76 DVDD.n45 4.5005
R17685 DVDD.n60 DVDD.n45 4.5005
R17686 DVDD.n75 DVDD.n45 4.5005
R17687 DVDD.n61 DVDD.n45 4.5005
R17688 DVDD.n74 DVDD.n45 4.5005
R17689 DVDD.n62 DVDD.n45 4.5005
R17690 DVDD.n73 DVDD.n45 4.5005
R17691 DVDD.n63 DVDD.n45 4.5005
R17692 DVDD.n71 DVDD.n45 4.5005
R17693 DVDD.n65 DVDD.n45 4.5005
R17694 DVDD.n22299 DVDD.n45 4.5005
R17695 DVDD.n22297 DVDD.n54 4.5005
R17696 DVDD.n58 DVDD.n54 4.5005
R17697 DVDD.n78 DVDD.n54 4.5005
R17698 DVDD.n59 DVDD.n54 4.5005
R17699 DVDD.n76 DVDD.n54 4.5005
R17700 DVDD.n60 DVDD.n54 4.5005
R17701 DVDD.n75 DVDD.n54 4.5005
R17702 DVDD.n61 DVDD.n54 4.5005
R17703 DVDD.n74 DVDD.n54 4.5005
R17704 DVDD.n62 DVDD.n54 4.5005
R17705 DVDD.n73 DVDD.n54 4.5005
R17706 DVDD.n63 DVDD.n54 4.5005
R17707 DVDD.n65 DVDD.n54 4.5005
R17708 DVDD.n22299 DVDD.n54 4.5005
R17709 DVDD.n22297 DVDD.n44 4.5005
R17710 DVDD.n58 DVDD.n44 4.5005
R17711 DVDD.n78 DVDD.n44 4.5005
R17712 DVDD.n59 DVDD.n44 4.5005
R17713 DVDD.n76 DVDD.n44 4.5005
R17714 DVDD.n60 DVDD.n44 4.5005
R17715 DVDD.n75 DVDD.n44 4.5005
R17716 DVDD.n61 DVDD.n44 4.5005
R17717 DVDD.n74 DVDD.n44 4.5005
R17718 DVDD.n62 DVDD.n44 4.5005
R17719 DVDD.n73 DVDD.n44 4.5005
R17720 DVDD.n63 DVDD.n44 4.5005
R17721 DVDD.n65 DVDD.n44 4.5005
R17722 DVDD.n22299 DVDD.n44 4.5005
R17723 DVDD.n22297 DVDD.n56 4.5005
R17724 DVDD.n58 DVDD.n56 4.5005
R17725 DVDD.n78 DVDD.n56 4.5005
R17726 DVDD.n59 DVDD.n56 4.5005
R17727 DVDD.n76 DVDD.n56 4.5005
R17728 DVDD.n60 DVDD.n56 4.5005
R17729 DVDD.n75 DVDD.n56 4.5005
R17730 DVDD.n61 DVDD.n56 4.5005
R17731 DVDD.n74 DVDD.n56 4.5005
R17732 DVDD.n62 DVDD.n56 4.5005
R17733 DVDD.n73 DVDD.n56 4.5005
R17734 DVDD.n63 DVDD.n56 4.5005
R17735 DVDD.n65 DVDD.n56 4.5005
R17736 DVDD.n22299 DVDD.n56 4.5005
R17737 DVDD.n22297 DVDD.n43 4.5005
R17738 DVDD.n58 DVDD.n43 4.5005
R17739 DVDD.n78 DVDD.n43 4.5005
R17740 DVDD.n59 DVDD.n43 4.5005
R17741 DVDD.n76 DVDD.n43 4.5005
R17742 DVDD.n60 DVDD.n43 4.5005
R17743 DVDD.n75 DVDD.n43 4.5005
R17744 DVDD.n61 DVDD.n43 4.5005
R17745 DVDD.n74 DVDD.n43 4.5005
R17746 DVDD.n62 DVDD.n43 4.5005
R17747 DVDD.n73 DVDD.n43 4.5005
R17748 DVDD.n63 DVDD.n43 4.5005
R17749 DVDD.n65 DVDD.n43 4.5005
R17750 DVDD.n43 DVDD.n42 4.5005
R17751 DVDD.n22299 DVDD.n43 4.5005
R17752 DVDD.n22299 DVDD.n22298 4.5005
R17753 DVDD.n22298 DVDD.n42 4.5005
R17754 DVDD.n22298 DVDD.n65 4.5005
R17755 DVDD.n22298 DVDD.n71 4.5005
R17756 DVDD.n22298 DVDD.n63 4.5005
R17757 DVDD.n22298 DVDD.n73 4.5005
R17758 DVDD.n22298 DVDD.n62 4.5005
R17759 DVDD.n22298 DVDD.n74 4.5005
R17760 DVDD.n22298 DVDD.n61 4.5005
R17761 DVDD.n22298 DVDD.n75 4.5005
R17762 DVDD.n22298 DVDD.n60 4.5005
R17763 DVDD.n22298 DVDD.n76 4.5005
R17764 DVDD.n22298 DVDD.n59 4.5005
R17765 DVDD.n22298 DVDD.n78 4.5005
R17766 DVDD.n22298 DVDD.n58 4.5005
R17767 DVDD.n22298 DVDD.n22297 4.5005
R17768 DVDD.n22 DVDD.n11 4.5005
R17769 DVDD.n22344 DVDD.n11 4.5005
R17770 DVDD.n11 DVDD.n4 4.5005
R17771 DVDD.n22344 DVDD.n9 4.5005
R17772 DVDD.n9 DVDD.n4 4.5005
R17773 DVDD.n22344 DVDD.n12 4.5005
R17774 DVDD.n12 DVDD.n4 4.5005
R17775 DVDD.n22343 DVDD.n1 4.5005
R17776 DVDD.n22343 DVDD.n22 4.5005
R17777 DVDD.n22344 DVDD.n22343 4.5005
R17778 DVDD.n22342 DVDD.n22337 4.5005
R17779 DVDD.n22337 DVDD.n14 4.5005
R17780 DVDD.n22337 DVDD.n26 4.5005
R17781 DVDD.n22337 DVDD.n15 4.5005
R17782 DVDD.n22337 DVDD.n24 4.5005
R17783 DVDD.n22337 DVDD.n17 4.5005
R17784 DVDD.n22337 DVDD.n23 4.5005
R17785 DVDD.n22337 DVDD.n18 4.5005
R17786 DVDD.n22337 DVDD.n0 4.5005
R17787 DVDD.n22337 DVDD.n1 4.5005
R17788 DVDD.n22337 DVDD.n22 4.5005
R17789 DVDD.n22337 DVDD.n4 4.5005
R17790 DVDD.n22342 DVDD.n32 4.5005
R17791 DVDD.n32 DVDD.n14 4.5005
R17792 DVDD.n32 DVDD.n26 4.5005
R17793 DVDD.n32 DVDD.n15 4.5005
R17794 DVDD.n32 DVDD.n25 4.5005
R17795 DVDD.n32 DVDD.n16 4.5005
R17796 DVDD.n32 DVDD.n24 4.5005
R17797 DVDD.n32 DVDD.n17 4.5005
R17798 DVDD.n32 DVDD.n23 4.5005
R17799 DVDD.n32 DVDD.n18 4.5005
R17800 DVDD.n32 DVDD.n0 4.5005
R17801 DVDD.n32 DVDD.n22 4.5005
R17802 DVDD.n32 DVDD.n4 4.5005
R17803 DVDD.n22342 DVDD.n22339 4.5005
R17804 DVDD.n22339 DVDD.n14 4.5005
R17805 DVDD.n22339 DVDD.n26 4.5005
R17806 DVDD.n22339 DVDD.n15 4.5005
R17807 DVDD.n22339 DVDD.n25 4.5005
R17808 DVDD.n22339 DVDD.n16 4.5005
R17809 DVDD.n22339 DVDD.n24 4.5005
R17810 DVDD.n22339 DVDD.n17 4.5005
R17811 DVDD.n22339 DVDD.n23 4.5005
R17812 DVDD.n22339 DVDD.n18 4.5005
R17813 DVDD.n22339 DVDD.n0 4.5005
R17814 DVDD.n22339 DVDD.n22 4.5005
R17815 DVDD.n22339 DVDD.n4 4.5005
R17816 DVDD.n22342 DVDD.n31 4.5005
R17817 DVDD.n31 DVDD.n14 4.5005
R17818 DVDD.n31 DVDD.n26 4.5005
R17819 DVDD.n31 DVDD.n15 4.5005
R17820 DVDD.n31 DVDD.n25 4.5005
R17821 DVDD.n31 DVDD.n16 4.5005
R17822 DVDD.n31 DVDD.n24 4.5005
R17823 DVDD.n31 DVDD.n17 4.5005
R17824 DVDD.n31 DVDD.n23 4.5005
R17825 DVDD.n31 DVDD.n18 4.5005
R17826 DVDD.n31 DVDD.n0 4.5005
R17827 DVDD.n31 DVDD.n22 4.5005
R17828 DVDD.n31 DVDD.n4 4.5005
R17829 DVDD.n22342 DVDD.n22341 4.5005
R17830 DVDD.n22341 DVDD.n14 4.5005
R17831 DVDD.n22341 DVDD.n26 4.5005
R17832 DVDD.n22341 DVDD.n15 4.5005
R17833 DVDD.n22341 DVDD.n25 4.5005
R17834 DVDD.n22341 DVDD.n16 4.5005
R17835 DVDD.n22341 DVDD.n24 4.5005
R17836 DVDD.n22341 DVDD.n17 4.5005
R17837 DVDD.n22341 DVDD.n23 4.5005
R17838 DVDD.n22341 DVDD.n18 4.5005
R17839 DVDD.n22341 DVDD.n0 4.5005
R17840 DVDD.n22341 DVDD.n22 4.5005
R17841 DVDD.n22341 DVDD.n4 4.5005
R17842 DVDD.n22342 DVDD.n30 4.5005
R17843 DVDD.n30 DVDD.n14 4.5005
R17844 DVDD.n30 DVDD.n26 4.5005
R17845 DVDD.n30 DVDD.n15 4.5005
R17846 DVDD.n30 DVDD.n25 4.5005
R17847 DVDD.n30 DVDD.n16 4.5005
R17848 DVDD.n30 DVDD.n24 4.5005
R17849 DVDD.n30 DVDD.n17 4.5005
R17850 DVDD.n30 DVDD.n23 4.5005
R17851 DVDD.n30 DVDD.n18 4.5005
R17852 DVDD.n30 DVDD.n0 4.5005
R17853 DVDD.n30 DVDD.n1 4.5005
R17854 DVDD.n30 DVDD.n22 4.5005
R17855 DVDD.n30 DVDD.n4 4.5005
R17856 DVDD.n22343 DVDD.n0 4.5005
R17857 DVDD.n22343 DVDD.n18 4.5005
R17858 DVDD.n22343 DVDD.n23 4.5005
R17859 DVDD.n22343 DVDD.n17 4.5005
R17860 DVDD.n22343 DVDD.n24 4.5005
R17861 DVDD.n22343 DVDD.n16 4.5005
R17862 DVDD.n22343 DVDD.n25 4.5005
R17863 DVDD.n22343 DVDD.n15 4.5005
R17864 DVDD.n22343 DVDD.n26 4.5005
R17865 DVDD.n22343 DVDD.n14 4.5005
R17866 DVDD.n22343 DVDD.n22342 4.5005
R17867 DVDD.n29 DVDD.n0 4.5005
R17868 DVDD.n29 DVDD.n18 4.5005
R17869 DVDD.n29 DVDD.n23 4.5005
R17870 DVDD.n29 DVDD.n17 4.5005
R17871 DVDD.n29 DVDD.n24 4.5005
R17872 DVDD.n29 DVDD.n16 4.5005
R17873 DVDD.n29 DVDD.n25 4.5005
R17874 DVDD.n29 DVDD.n15 4.5005
R17875 DVDD.n29 DVDD.n26 4.5005
R17876 DVDD.n29 DVDD.n14 4.5005
R17877 DVDD.n22342 DVDD.n29 4.5005
R17878 DVDD.n12 DVDD.n0 4.5005
R17879 DVDD.n18 DVDD.n12 4.5005
R17880 DVDD.n23 DVDD.n12 4.5005
R17881 DVDD.n17 DVDD.n12 4.5005
R17882 DVDD.n24 DVDD.n12 4.5005
R17883 DVDD.n16 DVDD.n12 4.5005
R17884 DVDD.n25 DVDD.n12 4.5005
R17885 DVDD.n15 DVDD.n12 4.5005
R17886 DVDD.n26 DVDD.n12 4.5005
R17887 DVDD.n14 DVDD.n12 4.5005
R17888 DVDD.n22342 DVDD.n12 4.5005
R17889 DVDD.n9 DVDD.n0 4.5005
R17890 DVDD.n18 DVDD.n9 4.5005
R17891 DVDD.n23 DVDD.n9 4.5005
R17892 DVDD.n17 DVDD.n9 4.5005
R17893 DVDD.n24 DVDD.n9 4.5005
R17894 DVDD.n16 DVDD.n9 4.5005
R17895 DVDD.n25 DVDD.n9 4.5005
R17896 DVDD.n15 DVDD.n9 4.5005
R17897 DVDD.n26 DVDD.n9 4.5005
R17898 DVDD.n14 DVDD.n9 4.5005
R17899 DVDD.n22342 DVDD.n9 4.5005
R17900 DVDD.n11 DVDD.n0 4.5005
R17901 DVDD.n18 DVDD.n11 4.5005
R17902 DVDD.n23 DVDD.n11 4.5005
R17903 DVDD.n17 DVDD.n11 4.5005
R17904 DVDD.n24 DVDD.n11 4.5005
R17905 DVDD.n16 DVDD.n11 4.5005
R17906 DVDD.n25 DVDD.n11 4.5005
R17907 DVDD.n15 DVDD.n11 4.5005
R17908 DVDD.n26 DVDD.n11 4.5005
R17909 DVDD.n14 DVDD.n11 4.5005
R17910 DVDD.n22342 DVDD.n11 4.5005
R17911 DVDD.n19193 DVDD.n18653 4.5005
R17912 DVDD.n19195 DVDD.n18653 4.5005
R17913 DVDD.n19203 DVDD.n19195 4.5005
R17914 DVDD.n19700 DVDD.n19195 4.5005
R17915 DVDD.n19204 DVDD.n19195 4.5005
R17916 DVDD.n19635 DVDD.n19194 4.5005
R17917 DVDD.n19635 DVDD.n19195 4.5005
R17918 DVDD.n19210 DVDD.n19194 4.5005
R17919 DVDD.n19210 DVDD.n19192 4.5005
R17920 DVDD.n19210 DVDD.n19196 4.5005
R17921 DVDD.n19210 DVDD.n19191 4.5005
R17922 DVDD.n19210 DVDD.n19197 4.5005
R17923 DVDD.n19210 DVDD.n19190 4.5005
R17924 DVDD.n19210 DVDD.n19198 4.5005
R17925 DVDD.n19210 DVDD.n19188 4.5005
R17926 DVDD.n19210 DVDD.n19200 4.5005
R17927 DVDD.n19701 DVDD.n19210 4.5005
R17928 DVDD.n19206 DVDD.n19194 4.5005
R17929 DVDD.n19206 DVDD.n19193 4.5005
R17930 DVDD.n19206 DVDD.n19195 4.5005
R17931 DVDD.n19206 DVDD.n19192 4.5005
R17932 DVDD.n19206 DVDD.n19196 4.5005
R17933 DVDD.n19206 DVDD.n19191 4.5005
R17934 DVDD.n19206 DVDD.n19197 4.5005
R17935 DVDD.n19206 DVDD.n19190 4.5005
R17936 DVDD.n19206 DVDD.n19198 4.5005
R17937 DVDD.n19206 DVDD.n19189 4.5005
R17938 DVDD.n19206 DVDD.n19199 4.5005
R17939 DVDD.n19206 DVDD.n19200 4.5005
R17940 DVDD.n19701 DVDD.n19206 4.5005
R17941 DVDD.n19212 DVDD.n19194 4.5005
R17942 DVDD.n19212 DVDD.n19193 4.5005
R17943 DVDD.n19212 DVDD.n19195 4.5005
R17944 DVDD.n19212 DVDD.n19192 4.5005
R17945 DVDD.n19212 DVDD.n19196 4.5005
R17946 DVDD.n19212 DVDD.n19191 4.5005
R17947 DVDD.n19212 DVDD.n19197 4.5005
R17948 DVDD.n19212 DVDD.n19190 4.5005
R17949 DVDD.n19212 DVDD.n19198 4.5005
R17950 DVDD.n19212 DVDD.n19189 4.5005
R17951 DVDD.n19212 DVDD.n19199 4.5005
R17952 DVDD.n19212 DVDD.n19200 4.5005
R17953 DVDD.n19701 DVDD.n19212 4.5005
R17954 DVDD.n19205 DVDD.n19194 4.5005
R17955 DVDD.n19205 DVDD.n19193 4.5005
R17956 DVDD.n19205 DVDD.n19195 4.5005
R17957 DVDD.n19205 DVDD.n19192 4.5005
R17958 DVDD.n19205 DVDD.n19196 4.5005
R17959 DVDD.n19205 DVDD.n19191 4.5005
R17960 DVDD.n19205 DVDD.n19197 4.5005
R17961 DVDD.n19205 DVDD.n19190 4.5005
R17962 DVDD.n19205 DVDD.n19198 4.5005
R17963 DVDD.n19205 DVDD.n19189 4.5005
R17964 DVDD.n19205 DVDD.n19199 4.5005
R17965 DVDD.n19205 DVDD.n19200 4.5005
R17966 DVDD.n19701 DVDD.n19205 4.5005
R17967 DVDD.n19214 DVDD.n19194 4.5005
R17968 DVDD.n19214 DVDD.n19193 4.5005
R17969 DVDD.n19214 DVDD.n19195 4.5005
R17970 DVDD.n19214 DVDD.n19192 4.5005
R17971 DVDD.n19214 DVDD.n19196 4.5005
R17972 DVDD.n19214 DVDD.n19191 4.5005
R17973 DVDD.n19214 DVDD.n19197 4.5005
R17974 DVDD.n19214 DVDD.n19190 4.5005
R17975 DVDD.n19214 DVDD.n19198 4.5005
R17976 DVDD.n19214 DVDD.n19189 4.5005
R17977 DVDD.n19214 DVDD.n19199 4.5005
R17978 DVDD.n19214 DVDD.n19200 4.5005
R17979 DVDD.n19701 DVDD.n19214 4.5005
R17980 DVDD.n19702 DVDD.n19194 4.5005
R17981 DVDD.n19702 DVDD.n19193 4.5005
R17982 DVDD.n19702 DVDD.n19195 4.5005
R17983 DVDD.n19702 DVDD.n19192 4.5005
R17984 DVDD.n19702 DVDD.n19196 4.5005
R17985 DVDD.n19702 DVDD.n19191 4.5005
R17986 DVDD.n19702 DVDD.n19197 4.5005
R17987 DVDD.n19702 DVDD.n19190 4.5005
R17988 DVDD.n19702 DVDD.n19198 4.5005
R17989 DVDD.n19702 DVDD.n19189 4.5005
R17990 DVDD.n19702 DVDD.n19199 4.5005
R17991 DVDD.n19702 DVDD.n19188 4.5005
R17992 DVDD.n19702 DVDD.n19200 4.5005
R17993 DVDD.n19702 DVDD.n19701 4.5005
R17994 DVDD.n19701 DVDD.n19635 4.5005
R17995 DVDD.n19699 DVDD.n19635 4.5005
R17996 DVDD.n19635 DVDD.n19200 4.5005
R17997 DVDD.n19635 DVDD.n19188 4.5005
R17998 DVDD.n19635 DVDD.n19199 4.5005
R17999 DVDD.n19635 DVDD.n19189 4.5005
R18000 DVDD.n19635 DVDD.n19198 4.5005
R18001 DVDD.n19635 DVDD.n19190 4.5005
R18002 DVDD.n19635 DVDD.n19197 4.5005
R18003 DVDD.n19635 DVDD.n19191 4.5005
R18004 DVDD.n19635 DVDD.n19196 4.5005
R18005 DVDD.n19701 DVDD.n19204 4.5005
R18006 DVDD.n19699 DVDD.n19204 4.5005
R18007 DVDD.n19204 DVDD.n19200 4.5005
R18008 DVDD.n19204 DVDD.n19188 4.5005
R18009 DVDD.n19204 DVDD.n19199 4.5005
R18010 DVDD.n19204 DVDD.n19189 4.5005
R18011 DVDD.n19204 DVDD.n19198 4.5005
R18012 DVDD.n19204 DVDD.n19190 4.5005
R18013 DVDD.n19204 DVDD.n19197 4.5005
R18014 DVDD.n19204 DVDD.n19191 4.5005
R18015 DVDD.n19204 DVDD.n19196 4.5005
R18016 DVDD.n19701 DVDD.n19700 4.5005
R18017 DVDD.n19700 DVDD.n19699 4.5005
R18018 DVDD.n19700 DVDD.n19200 4.5005
R18019 DVDD.n19700 DVDD.n19188 4.5005
R18020 DVDD.n19700 DVDD.n19199 4.5005
R18021 DVDD.n19700 DVDD.n19189 4.5005
R18022 DVDD.n19700 DVDD.n19198 4.5005
R18023 DVDD.n19700 DVDD.n19190 4.5005
R18024 DVDD.n19700 DVDD.n19197 4.5005
R18025 DVDD.n19700 DVDD.n19191 4.5005
R18026 DVDD.n19700 DVDD.n19196 4.5005
R18027 DVDD.n19701 DVDD.n19203 4.5005
R18028 DVDD.n19699 DVDD.n19203 4.5005
R18029 DVDD.n19203 DVDD.n19200 4.5005
R18030 DVDD.n19203 DVDD.n19188 4.5005
R18031 DVDD.n19203 DVDD.n19199 4.5005
R18032 DVDD.n19203 DVDD.n19189 4.5005
R18033 DVDD.n19203 DVDD.n19198 4.5005
R18034 DVDD.n19203 DVDD.n19190 4.5005
R18035 DVDD.n19203 DVDD.n19197 4.5005
R18036 DVDD.n19203 DVDD.n19191 4.5005
R18037 DVDD.n19203 DVDD.n19196 4.5005
R18038 DVDD.n19701 DVDD.n18653 4.5005
R18039 DVDD.n19699 DVDD.n18653 4.5005
R18040 DVDD.n19200 DVDD.n18653 4.5005
R18041 DVDD.n19188 DVDD.n18653 4.5005
R18042 DVDD.n19199 DVDD.n18653 4.5005
R18043 DVDD.n19189 DVDD.n18653 4.5005
R18044 DVDD.n19198 DVDD.n18653 4.5005
R18045 DVDD.n19190 DVDD.n18653 4.5005
R18046 DVDD.n19197 DVDD.n18653 4.5005
R18047 DVDD.n19191 DVDD.n18653 4.5005
R18048 DVDD.n19196 DVDD.n18653 4.5005
R18049 DVDD.n19635 DVDD.n19192 4.5005
R18050 DVDD.n19204 DVDD.n19192 4.5005
R18051 DVDD.n19700 DVDD.n19192 4.5005
R18052 DVDD.n19203 DVDD.n19192 4.5005
R18053 DVDD.n19192 DVDD.n18653 4.5005
R18054 DVDD.t67 DVDD.n19384 4.06554
R18055 DVDD.n21282 DVDD.t66 4.06554
R18056 DVDD.t155 DVDD 4.04483
R18057 DVDD DVDD.t155 4.04483
R18058 DVDD DVDD.t157 4.04483
R18059 DVDD.t157 DVDD 4.04483
R18060 DVDD.t158 DVDD 4.04483
R18061 DVDD DVDD.t158 4.04483
R18062 DVDD.t161 DVDD 4.04483
R18063 DVDD DVDD.t161 4.04483
R18064 DVDD.n19385 DVDD.t67 3.48482
R18065 DVDD.n21289 DVDD.t66 3.48482
R18066 DVDD.n19401 DVDD.t62 2.9041
R18067 DVDD.n21314 DVDD.t69 2.9041
R18068 DVDD.n21503 DVDD.n21502 2.33866
R18069 DVDD.n19338 DVDD.t63 2.32338
R18070 DVDD.n21321 DVDD.t65 2.32338
R18071 DVDD.n19331 DVDD.n19330 2.30804
R18072 DVDD.n19326 DVDD.n19320 2.30804
R18073 DVDD.n19324 DVDD.n19323 2.30804
R18074 DVDD.n19630 DVDD.n19217 2.30804
R18075 DVDD.n19628 DVDD.n19627 2.30804
R18076 DVDD.n19623 DVDD.n19221 2.30804
R18077 DVDD.n19621 DVDD.n19620 2.30804
R18078 DVDD.n19616 DVDD.n19224 2.30804
R18079 DVDD.n19614 DVDD.n19613 2.30804
R18080 DVDD.n19609 DVDD.n19227 2.30804
R18081 DVDD.n19607 DVDD.n19606 2.30804
R18082 DVDD.n19602 DVDD.n19230 2.30804
R18083 DVDD.n19600 DVDD.n19599 2.30804
R18084 DVDD.n19595 DVDD.n19233 2.30804
R18085 DVDD.n19593 DVDD.n19592 2.30804
R18086 DVDD.n19588 DVDD.n19238 2.30804
R18087 DVDD.n19586 DVDD.n19585 2.30804
R18088 DVDD.n19581 DVDD.n19241 2.30804
R18089 DVDD.n19579 DVDD.n19578 2.30804
R18090 DVDD.n19574 DVDD.n19244 2.30804
R18091 DVDD.n19572 DVDD.n19571 2.30804
R18092 DVDD.n19567 DVDD.n19247 2.30804
R18093 DVDD.n19565 DVDD.n19564 2.30804
R18094 DVDD.n19560 DVDD.n19250 2.30804
R18095 DVDD.n19558 DVDD.n19557 2.30804
R18096 DVDD.n19551 DVDD.n19253 2.30804
R18097 DVDD.n19549 DVDD.n19548 2.30804
R18098 DVDD.n19544 DVDD.n19256 2.30804
R18099 DVDD.n19542 DVDD.n19541 2.30804
R18100 DVDD.n19537 DVDD.n19259 2.30804
R18101 DVDD.n19535 DVDD.n19534 2.30804
R18102 DVDD.n19530 DVDD.n19262 2.30804
R18103 DVDD.n19528 DVDD.n19527 2.30804
R18104 DVDD.n19523 DVDD.n19265 2.30804
R18105 DVDD.n19521 DVDD.n19520 2.30804
R18106 DVDD.n19516 DVDD.n19268 2.30804
R18107 DVDD.n19514 DVDD.n19513 2.30804
R18108 DVDD.n19509 DVDD.n19271 2.30804
R18109 DVDD.n19507 DVDD.n19506 2.30804
R18110 DVDD.n19500 DVDD.n19274 2.30804
R18111 DVDD.n19498 DVDD.n19497 2.30804
R18112 DVDD.n19493 DVDD.n19277 2.30804
R18113 DVDD.n19491 DVDD.n19490 2.30804
R18114 DVDD.n19486 DVDD.n19280 2.30804
R18115 DVDD.n19484 DVDD.n19483 2.30804
R18116 DVDD.n19479 DVDD.n19283 2.30804
R18117 DVDD.n19477 DVDD.n19476 2.30804
R18118 DVDD.n19472 DVDD.n19286 2.30804
R18119 DVDD.n19470 DVDD.n19469 2.30804
R18120 DVDD.n19465 DVDD.n19290 2.30804
R18121 DVDD.n19463 DVDD.n19462 2.30804
R18122 DVDD.n19458 DVDD.n19294 2.30804
R18123 DVDD.n19456 DVDD.n19455 2.30804
R18124 DVDD.n19451 DVDD.n19297 2.30804
R18125 DVDD.n19449 DVDD.n19448 2.30804
R18126 DVDD.n19444 DVDD.n19300 2.30804
R18127 DVDD.n19442 DVDD.n19441 2.30804
R18128 DVDD.n19437 DVDD.n19303 2.30804
R18129 DVDD.n19435 DVDD.n19434 2.30804
R18130 DVDD.n19430 DVDD.n19306 2.30804
R18131 DVDD.n19428 DVDD.n19427 2.30804
R18132 DVDD.n19422 DVDD.n19309 2.30804
R18133 DVDD.n19420 DVDD.n19419 2.30804
R18134 DVDD.n19415 DVDD.n19312 2.30804
R18135 DVDD.n21491 DVDD.n21490 2.30804
R18136 DVDD.n21488 DVDD.n21487 2.30804
R18137 DVDD.n21483 DVDD.n21329 2.30804
R18138 DVDD.n21481 DVDD.n21480 2.30804
R18139 DVDD.n21476 DVDD.n21373 2.30804
R18140 DVDD.n21474 DVDD.n21473 2.30804
R18141 DVDD.n21469 DVDD.n21376 2.30804
R18142 DVDD.n21467 DVDD.n21466 2.30804
R18143 DVDD.n21462 DVDD.n21379 2.30804
R18144 DVDD.n21460 DVDD.n21459 2.30804
R18145 DVDD.n21455 DVDD.n21382 2.30804
R18146 DVDD.n21453 DVDD.n21452 2.30804
R18147 DVDD.n21448 DVDD.n21385 2.30804
R18148 DVDD.n21446 DVDD.n21445 2.30804
R18149 DVDD.n21439 DVDD.n21388 2.30804
R18150 DVDD.n21437 DVDD.n21436 2.30804
R18151 DVDD.n21432 DVDD.n21391 2.30804
R18152 DVDD.n21430 DVDD.n21429 2.30804
R18153 DVDD.n21425 DVDD.n21394 2.30804
R18154 DVDD.n21423 DVDD.n21422 2.30804
R18155 DVDD.n21418 DVDD.n21397 2.30804
R18156 DVDD.n21416 DVDD.n21415 2.30804
R18157 DVDD.n21411 DVDD.n21400 2.30804
R18158 DVDD.n21409 DVDD.n21408 2.30804
R18159 DVDD.n21404 DVDD.n21402 2.30804
R18160 DVDD.n21643 DVDD.n18559 2.30804
R18161 DVDD.n21641 DVDD.n21640 2.30804
R18162 DVDD.n21636 DVDD.n18563 2.30804
R18163 DVDD.n21634 DVDD.n21633 2.30804
R18164 DVDD.n21629 DVDD.n18566 2.30804
R18165 DVDD.n21627 DVDD.n21626 2.30804
R18166 DVDD.n21622 DVDD.n18569 2.30804
R18167 DVDD.n21620 DVDD.n21619 2.30804
R18168 DVDD.n21615 DVDD.n18572 2.30804
R18169 DVDD.n21613 DVDD.n21612 2.30804
R18170 DVDD.n21608 DVDD.n18575 2.30804
R18171 DVDD.n21606 DVDD.n21605 2.30804
R18172 DVDD.n21601 DVDD.n18578 2.30804
R18173 DVDD.n21599 DVDD.n21598 2.30804
R18174 DVDD.n21579 DVDD.n18581 2.30804
R18175 DVDD.n21577 DVDD.n21576 2.30804
R18176 DVDD.n21572 DVDD.n18584 2.30804
R18177 DVDD.n21570 DVDD.n21569 2.30804
R18178 DVDD.n21565 DVDD.n18587 2.30804
R18179 DVDD.n21563 DVDD.n21562 2.30804
R18180 DVDD.n21558 DVDD.n18590 2.30804
R18181 DVDD.n21556 DVDD.n21555 2.30804
R18182 DVDD.n21551 DVDD.n18593 2.30804
R18183 DVDD.n21549 DVDD.n21548 2.30804
R18184 DVDD.n21544 DVDD.n18596 2.30804
R18185 DVDD.n21542 DVDD.n21541 2.30804
R18186 DVDD.n21537 DVDD.n18600 2.30804
R18187 DVDD.n21535 DVDD.n21534 2.30804
R18188 DVDD.n21530 DVDD.n18603 2.30804
R18189 DVDD.n21528 DVDD.n21527 2.30804
R18190 DVDD.n21523 DVDD.n18606 2.30804
R18191 DVDD.n21521 DVDD.n21520 2.30804
R18192 DVDD.n21516 DVDD.n18609 2.30804
R18193 DVDD.n21514 DVDD.n21513 2.30804
R18194 DVDD.n21509 DVDD.n18612 2.30804
R18195 DVDD.n21507 DVDD.n21506 2.30804
R18196 DVDD.n21500 DVDD.n21499 2.30804
R18197 DVDD.n21501 DVDD.n21500 2.30804
R18198 DVDD.n18615 DVDD.n18613 2.30804
R18199 DVDD.n21508 DVDD.n21507 2.30804
R18200 DVDD.n18612 DVDD.n18610 2.30804
R18201 DVDD.n21515 DVDD.n21514 2.30804
R18202 DVDD.n18609 DVDD.n18607 2.30804
R18203 DVDD.n21522 DVDD.n21521 2.30804
R18204 DVDD.n18606 DVDD.n18604 2.30804
R18205 DVDD.n21529 DVDD.n21528 2.30804
R18206 DVDD.n18603 DVDD.n18601 2.30804
R18207 DVDD.n21536 DVDD.n21535 2.30804
R18208 DVDD.n18600 DVDD.n18598 2.30804
R18209 DVDD.n21543 DVDD.n21542 2.30804
R18210 DVDD.n18596 DVDD.n18594 2.30804
R18211 DVDD.n21550 DVDD.n21549 2.30804
R18212 DVDD.n18593 DVDD.n18591 2.30804
R18213 DVDD.n21557 DVDD.n21556 2.30804
R18214 DVDD.n18590 DVDD.n18588 2.30804
R18215 DVDD.n21564 DVDD.n21563 2.30804
R18216 DVDD.n18587 DVDD.n18585 2.30804
R18217 DVDD.n21571 DVDD.n21570 2.30804
R18218 DVDD.n18584 DVDD.n18582 2.30804
R18219 DVDD.n21578 DVDD.n21577 2.30804
R18220 DVDD.n18581 DVDD.n18579 2.30804
R18221 DVDD.n21600 DVDD.n21599 2.30804
R18222 DVDD.n18578 DVDD.n18576 2.30804
R18223 DVDD.n21607 DVDD.n21606 2.30804
R18224 DVDD.n18575 DVDD.n18573 2.30804
R18225 DVDD.n21614 DVDD.n21613 2.30804
R18226 DVDD.n18572 DVDD.n18570 2.30804
R18227 DVDD.n21621 DVDD.n21620 2.30804
R18228 DVDD.n18569 DVDD.n18567 2.30804
R18229 DVDD.n21628 DVDD.n21627 2.30804
R18230 DVDD.n18566 DVDD.n18564 2.30804
R18231 DVDD.n21635 DVDD.n21634 2.30804
R18232 DVDD.n18563 DVDD.n18561 2.30804
R18233 DVDD.n21642 DVDD.n21641 2.30804
R18234 DVDD.n21403 DVDD.n18559 2.30804
R18235 DVDD.n21402 DVDD.n21401 2.30804
R18236 DVDD.n21410 DVDD.n21409 2.30804
R18237 DVDD.n21400 DVDD.n21398 2.30804
R18238 DVDD.n21417 DVDD.n21416 2.30804
R18239 DVDD.n21397 DVDD.n21395 2.30804
R18240 DVDD.n21424 DVDD.n21423 2.30804
R18241 DVDD.n21394 DVDD.n21392 2.30804
R18242 DVDD.n21431 DVDD.n21430 2.30804
R18243 DVDD.n21391 DVDD.n21389 2.30804
R18244 DVDD.n21438 DVDD.n21437 2.30804
R18245 DVDD.n21388 DVDD.n21386 2.30804
R18246 DVDD.n21447 DVDD.n21446 2.30804
R18247 DVDD.n21385 DVDD.n21383 2.30804
R18248 DVDD.n21454 DVDD.n21453 2.30804
R18249 DVDD.n21382 DVDD.n21380 2.30804
R18250 DVDD.n21461 DVDD.n21460 2.30804
R18251 DVDD.n21379 DVDD.n21377 2.30804
R18252 DVDD.n21468 DVDD.n21467 2.30804
R18253 DVDD.n21376 DVDD.n21374 2.30804
R18254 DVDD.n21475 DVDD.n21474 2.30804
R18255 DVDD.n21373 DVDD.n21330 2.30804
R18256 DVDD.n21482 DVDD.n21481 2.30804
R18257 DVDD.n21329 DVDD.n21327 2.30804
R18258 DVDD.n21489 DVDD.n21488 2.30804
R18259 DVDD.n21492 DVDD.n21491 2.30804
R18260 DVDD.n19414 DVDD.n19413 2.30804
R18261 DVDD.n19312 DVDD.n19310 2.30804
R18262 DVDD.n19421 DVDD.n19420 2.30804
R18263 DVDD.n19309 DVDD.n19307 2.30804
R18264 DVDD.n19429 DVDD.n19428 2.30804
R18265 DVDD.n19306 DVDD.n19304 2.30804
R18266 DVDD.n19436 DVDD.n19435 2.30804
R18267 DVDD.n19303 DVDD.n19301 2.30804
R18268 DVDD.n19443 DVDD.n19442 2.30804
R18269 DVDD.n19300 DVDD.n19298 2.30804
R18270 DVDD.n19450 DVDD.n19449 2.30804
R18271 DVDD.n19297 DVDD.n19295 2.30804
R18272 DVDD.n19457 DVDD.n19456 2.30804
R18273 DVDD.n19294 DVDD.n19292 2.30804
R18274 DVDD.n19464 DVDD.n19463 2.30804
R18275 DVDD.n19290 DVDD.n19287 2.30804
R18276 DVDD.n19471 DVDD.n19470 2.30804
R18277 DVDD.n19286 DVDD.n19284 2.30804
R18278 DVDD.n19478 DVDD.n19477 2.30804
R18279 DVDD.n19283 DVDD.n19281 2.30804
R18280 DVDD.n19485 DVDD.n19484 2.30804
R18281 DVDD.n19280 DVDD.n19278 2.30804
R18282 DVDD.n19492 DVDD.n19491 2.30804
R18283 DVDD.n19277 DVDD.n19275 2.30804
R18284 DVDD.n19499 DVDD.n19498 2.30804
R18285 DVDD.n19274 DVDD.n19272 2.30804
R18286 DVDD.n19508 DVDD.n19507 2.30804
R18287 DVDD.n19271 DVDD.n19269 2.30804
R18288 DVDD.n19515 DVDD.n19514 2.30804
R18289 DVDD.n19268 DVDD.n19266 2.30804
R18290 DVDD.n19522 DVDD.n19521 2.30804
R18291 DVDD.n19265 DVDD.n19263 2.30804
R18292 DVDD.n19529 DVDD.n19528 2.30804
R18293 DVDD.n19262 DVDD.n19260 2.30804
R18294 DVDD.n19536 DVDD.n19535 2.30804
R18295 DVDD.n19259 DVDD.n19257 2.30804
R18296 DVDD.n19543 DVDD.n19542 2.30804
R18297 DVDD.n19256 DVDD.n19254 2.30804
R18298 DVDD.n19550 DVDD.n19549 2.30804
R18299 DVDD.n19253 DVDD.n19251 2.30804
R18300 DVDD.n19559 DVDD.n19558 2.30804
R18301 DVDD.n19250 DVDD.n19248 2.30804
R18302 DVDD.n19566 DVDD.n19565 2.30804
R18303 DVDD.n19247 DVDD.n19245 2.30804
R18304 DVDD.n19573 DVDD.n19572 2.30804
R18305 DVDD.n19244 DVDD.n19242 2.30804
R18306 DVDD.n19580 DVDD.n19579 2.30804
R18307 DVDD.n19241 DVDD.n19239 2.30804
R18308 DVDD.n19587 DVDD.n19586 2.30804
R18309 DVDD.n19238 DVDD.n19234 2.30804
R18310 DVDD.n19594 DVDD.n19593 2.30804
R18311 DVDD.n19233 DVDD.n19231 2.30804
R18312 DVDD.n19601 DVDD.n19600 2.30804
R18313 DVDD.n19230 DVDD.n19228 2.30804
R18314 DVDD.n19608 DVDD.n19607 2.30804
R18315 DVDD.n19227 DVDD.n19225 2.30804
R18316 DVDD.n19615 DVDD.n19614 2.30804
R18317 DVDD.n19224 DVDD.n19222 2.30804
R18318 DVDD.n19622 DVDD.n19621 2.30804
R18319 DVDD.n19221 DVDD.n19219 2.30804
R18320 DVDD.n19629 DVDD.n19628 2.30804
R18321 DVDD.n19321 DVDD.n19217 2.30804
R18322 DVDD.n19325 DVDD.n19324 2.30804
R18323 DVDD.n19320 DVDD.n19318 2.30804
R18324 DVDD.n19332 DVDD.n19331 2.30804
R18325 DVDD.n17310 DVDD.n898 2.25086
R18326 DVDD.n15087 DVDD.n7042 2.2505
R18327 DVDD.n7041 DVDD.n6797 2.2505
R18328 DVDD.n7040 DVDD.n7039 2.2505
R18329 DVDD.n7037 DVDD.n6798 2.2505
R18330 DVDD.n7035 DVDD.n7033 2.2505
R18331 DVDD.n7032 DVDD.n6800 2.2505
R18332 DVDD.n7031 DVDD.n7030 2.2505
R18333 DVDD.n7028 DVDD.n6801 2.2505
R18334 DVDD.n7026 DVDD.n7024 2.2505
R18335 DVDD.n7023 DVDD.n6803 2.2505
R18336 DVDD.n7022 DVDD.n7021 2.2505
R18337 DVDD.n7019 DVDD.n6804 2.2505
R18338 DVDD.n7017 DVDD.n7015 2.2505
R18339 DVDD.n7014 DVDD.n6806 2.2505
R18340 DVDD.n7013 DVDD.n7012 2.2505
R18341 DVDD.n7010 DVDD.n6807 2.2505
R18342 DVDD.n7008 DVDD.n7006 2.2505
R18343 DVDD.n7005 DVDD.n6809 2.2505
R18344 DVDD.n7004 DVDD.n7003 2.2505
R18345 DVDD.n7001 DVDD.n6810 2.2505
R18346 DVDD.n6999 DVDD.n6997 2.2505
R18347 DVDD.n6996 DVDD.n6812 2.2505
R18348 DVDD.n6995 DVDD.n6994 2.2505
R18349 DVDD.n6992 DVDD.n6813 2.2505
R18350 DVDD.n6990 DVDD.n6988 2.2505
R18351 DVDD.n6987 DVDD.n6815 2.2505
R18352 DVDD.n6986 DVDD.n6985 2.2505
R18353 DVDD.n6983 DVDD.n6816 2.2505
R18354 DVDD.n6981 DVDD.n6979 2.2505
R18355 DVDD.n6978 DVDD.n6818 2.2505
R18356 DVDD.n6977 DVDD.n6976 2.2505
R18357 DVDD.n6974 DVDD.n6819 2.2505
R18358 DVDD.n6972 DVDD.n6970 2.2505
R18359 DVDD.n6969 DVDD.n6821 2.2505
R18360 DVDD.n6968 DVDD.n6967 2.2505
R18361 DVDD.n6965 DVDD.n6822 2.2505
R18362 DVDD.n6963 DVDD.n6961 2.2505
R18363 DVDD.n6960 DVDD.n6824 2.2505
R18364 DVDD.n6959 DVDD.n6958 2.2505
R18365 DVDD.n6956 DVDD.n6825 2.2505
R18366 DVDD.n6954 DVDD.n6952 2.2505
R18367 DVDD.n6951 DVDD.n6827 2.2505
R18368 DVDD.n6950 DVDD.n6949 2.2505
R18369 DVDD.n6947 DVDD.n6828 2.2505
R18370 DVDD.n6945 DVDD.n6943 2.2505
R18371 DVDD.n6942 DVDD.n6830 2.2505
R18372 DVDD.n6941 DVDD.n6940 2.2505
R18373 DVDD.n6938 DVDD.n6831 2.2505
R18374 DVDD.n6936 DVDD.n6934 2.2505
R18375 DVDD.n6933 DVDD.n6833 2.2505
R18376 DVDD.n6932 DVDD.n6931 2.2505
R18377 DVDD.n6929 DVDD.n6834 2.2505
R18378 DVDD.n6927 DVDD.n6925 2.2505
R18379 DVDD.n6924 DVDD.n6836 2.2505
R18380 DVDD.n6923 DVDD.n6922 2.2505
R18381 DVDD.n6920 DVDD.n6837 2.2505
R18382 DVDD.n6918 DVDD.n6916 2.2505
R18383 DVDD.n6915 DVDD.n6839 2.2505
R18384 DVDD.n6914 DVDD.n6913 2.2505
R18385 DVDD.n6911 DVDD.n6840 2.2505
R18386 DVDD.n6909 DVDD.n6907 2.2505
R18387 DVDD.n6906 DVDD.n6842 2.2505
R18388 DVDD.n6905 DVDD.n6904 2.2505
R18389 DVDD.n6902 DVDD.n6843 2.2505
R18390 DVDD.n6900 DVDD.n6898 2.2505
R18391 DVDD.n6897 DVDD.n6845 2.2505
R18392 DVDD.n6896 DVDD.n6895 2.2505
R18393 DVDD.n6893 DVDD.n6846 2.2505
R18394 DVDD.n6891 DVDD.n6889 2.2505
R18395 DVDD.n6888 DVDD.n6848 2.2505
R18396 DVDD.n6887 DVDD.n6886 2.2505
R18397 DVDD.n6884 DVDD.n6849 2.2505
R18398 DVDD.n6882 DVDD.n6880 2.2505
R18399 DVDD.n6879 DVDD.n6851 2.2505
R18400 DVDD.n6878 DVDD.n6877 2.2505
R18401 DVDD.n6875 DVDD.n6852 2.2505
R18402 DVDD.n6873 DVDD.n6871 2.2505
R18403 DVDD.n6870 DVDD.n6854 2.2505
R18404 DVDD.n6869 DVDD.n6868 2.2505
R18405 DVDD.n6866 DVDD.n6855 2.2505
R18406 DVDD.n6864 DVDD.n6862 2.2505
R18407 DVDD.n6861 DVDD.n6857 2.2505
R18408 DVDD.n6860 DVDD.n6859 2.2505
R18409 DVDD.n6858 DVDD.n6751 2.2505
R18410 DVDD.n15090 DVDD.n6751 2.2505
R18411 DVDD.n6859 DVDD.n6750 2.2505
R18412 DVDD.n6857 DVDD.n6856 2.2505
R18413 DVDD.n6864 DVDD.n6863 2.2505
R18414 DVDD.n6866 DVDD.n6865 2.2505
R18415 DVDD.n6868 DVDD.n6867 2.2505
R18416 DVDD.n6854 DVDD.n6853 2.2505
R18417 DVDD.n6873 DVDD.n6872 2.2505
R18418 DVDD.n6875 DVDD.n6874 2.2505
R18419 DVDD.n6877 DVDD.n6876 2.2505
R18420 DVDD.n6851 DVDD.n6850 2.2505
R18421 DVDD.n6882 DVDD.n6881 2.2505
R18422 DVDD.n6884 DVDD.n6883 2.2505
R18423 DVDD.n6886 DVDD.n6885 2.2505
R18424 DVDD.n6848 DVDD.n6847 2.2505
R18425 DVDD.n6891 DVDD.n6890 2.2505
R18426 DVDD.n6893 DVDD.n6892 2.2505
R18427 DVDD.n6895 DVDD.n6894 2.2505
R18428 DVDD.n6845 DVDD.n6844 2.2505
R18429 DVDD.n6900 DVDD.n6899 2.2505
R18430 DVDD.n6902 DVDD.n6901 2.2505
R18431 DVDD.n6904 DVDD.n6903 2.2505
R18432 DVDD.n6842 DVDD.n6841 2.2505
R18433 DVDD.n6909 DVDD.n6908 2.2505
R18434 DVDD.n6911 DVDD.n6910 2.2505
R18435 DVDD.n6913 DVDD.n6912 2.2505
R18436 DVDD.n6839 DVDD.n6838 2.2505
R18437 DVDD.n6918 DVDD.n6917 2.2505
R18438 DVDD.n6920 DVDD.n6919 2.2505
R18439 DVDD.n6922 DVDD.n6921 2.2505
R18440 DVDD.n6836 DVDD.n6835 2.2505
R18441 DVDD.n6927 DVDD.n6926 2.2505
R18442 DVDD.n6929 DVDD.n6928 2.2505
R18443 DVDD.n6931 DVDD.n6930 2.2505
R18444 DVDD.n6833 DVDD.n6832 2.2505
R18445 DVDD.n6936 DVDD.n6935 2.2505
R18446 DVDD.n6938 DVDD.n6937 2.2505
R18447 DVDD.n6940 DVDD.n6939 2.2505
R18448 DVDD.n6830 DVDD.n6829 2.2505
R18449 DVDD.n6945 DVDD.n6944 2.2505
R18450 DVDD.n6947 DVDD.n6946 2.2505
R18451 DVDD.n6949 DVDD.n6948 2.2505
R18452 DVDD.n6827 DVDD.n6826 2.2505
R18453 DVDD.n6954 DVDD.n6953 2.2505
R18454 DVDD.n6956 DVDD.n6955 2.2505
R18455 DVDD.n6958 DVDD.n6957 2.2505
R18456 DVDD.n6824 DVDD.n6823 2.2505
R18457 DVDD.n6963 DVDD.n6962 2.2505
R18458 DVDD.n6965 DVDD.n6964 2.2505
R18459 DVDD.n6967 DVDD.n6966 2.2505
R18460 DVDD.n6821 DVDD.n6820 2.2505
R18461 DVDD.n6972 DVDD.n6971 2.2505
R18462 DVDD.n6974 DVDD.n6973 2.2505
R18463 DVDD.n6976 DVDD.n6975 2.2505
R18464 DVDD.n6818 DVDD.n6817 2.2505
R18465 DVDD.n6981 DVDD.n6980 2.2505
R18466 DVDD.n6983 DVDD.n6982 2.2505
R18467 DVDD.n6985 DVDD.n6984 2.2505
R18468 DVDD.n6815 DVDD.n6814 2.2505
R18469 DVDD.n6990 DVDD.n6989 2.2505
R18470 DVDD.n6992 DVDD.n6991 2.2505
R18471 DVDD.n6994 DVDD.n6993 2.2505
R18472 DVDD.n6812 DVDD.n6811 2.2505
R18473 DVDD.n6999 DVDD.n6998 2.2505
R18474 DVDD.n7001 DVDD.n7000 2.2505
R18475 DVDD.n7003 DVDD.n7002 2.2505
R18476 DVDD.n6809 DVDD.n6808 2.2505
R18477 DVDD.n7008 DVDD.n7007 2.2505
R18478 DVDD.n7010 DVDD.n7009 2.2505
R18479 DVDD.n7012 DVDD.n7011 2.2505
R18480 DVDD.n6806 DVDD.n6805 2.2505
R18481 DVDD.n7017 DVDD.n7016 2.2505
R18482 DVDD.n7019 DVDD.n7018 2.2505
R18483 DVDD.n7021 DVDD.n7020 2.2505
R18484 DVDD.n6803 DVDD.n6802 2.2505
R18485 DVDD.n7026 DVDD.n7025 2.2505
R18486 DVDD.n7028 DVDD.n7027 2.2505
R18487 DVDD.n7030 DVDD.n7029 2.2505
R18488 DVDD.n6800 DVDD.n6799 2.2505
R18489 DVDD.n7035 DVDD.n7034 2.2505
R18490 DVDD.n7037 DVDD.n7036 2.2505
R18491 DVDD.n7039 DVDD.n7038 2.2505
R18492 DVDD.n6797 DVDD.n6796 2.2505
R18493 DVDD.n15088 DVDD.n15087 2.2505
R18494 DVDD.n7398 DVDD.n7112 2.2505
R18495 DVDD.n7400 DVDD.n7399 2.2505
R18496 DVDD.n7397 DVDD.n7113 2.2505
R18497 DVDD.n7396 DVDD.n7395 2.2505
R18498 DVDD.n7391 DVDD.n7114 2.2505
R18499 DVDD.n7387 DVDD.n7386 2.2505
R18500 DVDD.n7385 DVDD.n7115 2.2505
R18501 DVDD.n7384 DVDD.n7383 2.2505
R18502 DVDD.n7379 DVDD.n7116 2.2505
R18503 DVDD.n7375 DVDD.n7374 2.2505
R18504 DVDD.n7373 DVDD.n7117 2.2505
R18505 DVDD.n7372 DVDD.n7371 2.2505
R18506 DVDD.n7367 DVDD.n7118 2.2505
R18507 DVDD.n7363 DVDD.n7362 2.2505
R18508 DVDD.n7361 DVDD.n7119 2.2505
R18509 DVDD.n7360 DVDD.n7359 2.2505
R18510 DVDD.n7355 DVDD.n7120 2.2505
R18511 DVDD.n7351 DVDD.n7350 2.2505
R18512 DVDD.n7349 DVDD.n7121 2.2505
R18513 DVDD.n7348 DVDD.n7347 2.2505
R18514 DVDD.n7343 DVDD.n7122 2.2505
R18515 DVDD.n7339 DVDD.n7338 2.2505
R18516 DVDD.n7337 DVDD.n7123 2.2505
R18517 DVDD.n7336 DVDD.n7335 2.2505
R18518 DVDD.n7331 DVDD.n7124 2.2505
R18519 DVDD.n7327 DVDD.n7326 2.2505
R18520 DVDD.n7325 DVDD.n7125 2.2505
R18521 DVDD.n7324 DVDD.n7323 2.2505
R18522 DVDD.n7319 DVDD.n7126 2.2505
R18523 DVDD.n7315 DVDD.n7314 2.2505
R18524 DVDD.n7313 DVDD.n7127 2.2505
R18525 DVDD.n7312 DVDD.n7311 2.2505
R18526 DVDD.n7307 DVDD.n7128 2.2505
R18527 DVDD.n7303 DVDD.n7302 2.2505
R18528 DVDD.n7301 DVDD.n7129 2.2505
R18529 DVDD.n7300 DVDD.n7299 2.2505
R18530 DVDD.n7295 DVDD.n7130 2.2505
R18531 DVDD.n7291 DVDD.n7290 2.2505
R18532 DVDD.n7289 DVDD.n7131 2.2505
R18533 DVDD.n7288 DVDD.n7287 2.2505
R18534 DVDD.n7283 DVDD.n7132 2.2505
R18535 DVDD.n7279 DVDD.n7278 2.2505
R18536 DVDD.n7277 DVDD.n7133 2.2505
R18537 DVDD.n7276 DVDD.n7275 2.2505
R18538 DVDD.n7271 DVDD.n7134 2.2505
R18539 DVDD.n7267 DVDD.n7266 2.2505
R18540 DVDD.n7265 DVDD.n7135 2.2505
R18541 DVDD.n7264 DVDD.n7263 2.2505
R18542 DVDD.n7259 DVDD.n7136 2.2505
R18543 DVDD.n7255 DVDD.n7254 2.2505
R18544 DVDD.n7253 DVDD.n7137 2.2505
R18545 DVDD.n7252 DVDD.n7251 2.2505
R18546 DVDD.n7247 DVDD.n7138 2.2505
R18547 DVDD.n7243 DVDD.n7242 2.2505
R18548 DVDD.n7241 DVDD.n7139 2.2505
R18549 DVDD.n7240 DVDD.n7239 2.2505
R18550 DVDD.n7235 DVDD.n7140 2.2505
R18551 DVDD.n7231 DVDD.n7230 2.2505
R18552 DVDD.n7229 DVDD.n7141 2.2505
R18553 DVDD.n7228 DVDD.n7227 2.2505
R18554 DVDD.n7223 DVDD.n7142 2.2505
R18555 DVDD.n7219 DVDD.n7218 2.2505
R18556 DVDD.n7217 DVDD.n7143 2.2505
R18557 DVDD.n7216 DVDD.n7215 2.2505
R18558 DVDD.n7211 DVDD.n7144 2.2505
R18559 DVDD.n7207 DVDD.n7206 2.2505
R18560 DVDD.n7205 DVDD.n7145 2.2505
R18561 DVDD.n7204 DVDD.n7203 2.2505
R18562 DVDD.n7199 DVDD.n7146 2.2505
R18563 DVDD.n7195 DVDD.n7194 2.2505
R18564 DVDD.n7193 DVDD.n7147 2.2505
R18565 DVDD.n7192 DVDD.n7191 2.2505
R18566 DVDD.n7187 DVDD.n7148 2.2505
R18567 DVDD.n7183 DVDD.n7182 2.2505
R18568 DVDD.n7181 DVDD.n7149 2.2505
R18569 DVDD.n7180 DVDD.n7179 2.2505
R18570 DVDD.n7175 DVDD.n7150 2.2505
R18571 DVDD.n7171 DVDD.n7170 2.2505
R18572 DVDD.n7169 DVDD.n7151 2.2505
R18573 DVDD.n7168 DVDD.n7167 2.2505
R18574 DVDD.n7163 DVDD.n7152 2.2505
R18575 DVDD.n7159 DVDD.n7158 2.2505
R18576 DVDD.n7157 DVDD.n7156 2.2505
R18577 DVDD.n7153 DVDD.n7066 2.2505
R18578 DVDD.n7153 DVDD.n7111 2.2505
R18579 DVDD.n7156 DVDD.n7155 2.2505
R18580 DVDD.n7160 DVDD.n7159 2.2505
R18581 DVDD.n7163 DVDD.n7162 2.2505
R18582 DVDD.n7167 DVDD.n7166 2.2505
R18583 DVDD.n7164 DVDD.n7151 2.2505
R18584 DVDD.n7172 DVDD.n7171 2.2505
R18585 DVDD.n7175 DVDD.n7174 2.2505
R18586 DVDD.n7179 DVDD.n7178 2.2505
R18587 DVDD.n7176 DVDD.n7149 2.2505
R18588 DVDD.n7184 DVDD.n7183 2.2505
R18589 DVDD.n7187 DVDD.n7186 2.2505
R18590 DVDD.n7191 DVDD.n7190 2.2505
R18591 DVDD.n7188 DVDD.n7147 2.2505
R18592 DVDD.n7196 DVDD.n7195 2.2505
R18593 DVDD.n7199 DVDD.n7198 2.2505
R18594 DVDD.n7203 DVDD.n7202 2.2505
R18595 DVDD.n7200 DVDD.n7145 2.2505
R18596 DVDD.n7208 DVDD.n7207 2.2505
R18597 DVDD.n7211 DVDD.n7210 2.2505
R18598 DVDD.n7215 DVDD.n7214 2.2505
R18599 DVDD.n7212 DVDD.n7143 2.2505
R18600 DVDD.n7220 DVDD.n7219 2.2505
R18601 DVDD.n7223 DVDD.n7222 2.2505
R18602 DVDD.n7227 DVDD.n7226 2.2505
R18603 DVDD.n7224 DVDD.n7141 2.2505
R18604 DVDD.n7232 DVDD.n7231 2.2505
R18605 DVDD.n7235 DVDD.n7234 2.2505
R18606 DVDD.n7239 DVDD.n7238 2.2505
R18607 DVDD.n7236 DVDD.n7139 2.2505
R18608 DVDD.n7244 DVDD.n7243 2.2505
R18609 DVDD.n7247 DVDD.n7246 2.2505
R18610 DVDD.n7251 DVDD.n7250 2.2505
R18611 DVDD.n7248 DVDD.n7137 2.2505
R18612 DVDD.n7256 DVDD.n7255 2.2505
R18613 DVDD.n7259 DVDD.n7258 2.2505
R18614 DVDD.n7263 DVDD.n7262 2.2505
R18615 DVDD.n7260 DVDD.n7135 2.2505
R18616 DVDD.n7268 DVDD.n7267 2.2505
R18617 DVDD.n7271 DVDD.n7270 2.2505
R18618 DVDD.n7275 DVDD.n7274 2.2505
R18619 DVDD.n7272 DVDD.n7133 2.2505
R18620 DVDD.n7280 DVDD.n7279 2.2505
R18621 DVDD.n7283 DVDD.n7282 2.2505
R18622 DVDD.n7287 DVDD.n7286 2.2505
R18623 DVDD.n7284 DVDD.n7131 2.2505
R18624 DVDD.n7292 DVDD.n7291 2.2505
R18625 DVDD.n7295 DVDD.n7294 2.2505
R18626 DVDD.n7299 DVDD.n7298 2.2505
R18627 DVDD.n7296 DVDD.n7129 2.2505
R18628 DVDD.n7304 DVDD.n7303 2.2505
R18629 DVDD.n7307 DVDD.n7306 2.2505
R18630 DVDD.n7311 DVDD.n7310 2.2505
R18631 DVDD.n7308 DVDD.n7127 2.2505
R18632 DVDD.n7316 DVDD.n7315 2.2505
R18633 DVDD.n7319 DVDD.n7318 2.2505
R18634 DVDD.n7323 DVDD.n7322 2.2505
R18635 DVDD.n7320 DVDD.n7125 2.2505
R18636 DVDD.n7328 DVDD.n7327 2.2505
R18637 DVDD.n7331 DVDD.n7330 2.2505
R18638 DVDD.n7335 DVDD.n7334 2.2505
R18639 DVDD.n7332 DVDD.n7123 2.2505
R18640 DVDD.n7340 DVDD.n7339 2.2505
R18641 DVDD.n7343 DVDD.n7342 2.2505
R18642 DVDD.n7347 DVDD.n7346 2.2505
R18643 DVDD.n7344 DVDD.n7121 2.2505
R18644 DVDD.n7352 DVDD.n7351 2.2505
R18645 DVDD.n7355 DVDD.n7354 2.2505
R18646 DVDD.n7359 DVDD.n7358 2.2505
R18647 DVDD.n7356 DVDD.n7119 2.2505
R18648 DVDD.n7364 DVDD.n7363 2.2505
R18649 DVDD.n7367 DVDD.n7366 2.2505
R18650 DVDD.n7371 DVDD.n7370 2.2505
R18651 DVDD.n7368 DVDD.n7117 2.2505
R18652 DVDD.n7376 DVDD.n7375 2.2505
R18653 DVDD.n7379 DVDD.n7378 2.2505
R18654 DVDD.n7383 DVDD.n7382 2.2505
R18655 DVDD.n7380 DVDD.n7115 2.2505
R18656 DVDD.n7388 DVDD.n7387 2.2505
R18657 DVDD.n7391 DVDD.n7390 2.2505
R18658 DVDD.n7395 DVDD.n7394 2.2505
R18659 DVDD.n7392 DVDD.n7113 2.2505
R18660 DVDD.n7401 DVDD.n7400 2.2505
R18661 DVDD.n7403 DVDD.n7112 2.2505
R18662 DVDD.n15055 DVDD.n15054 2.2505
R18663 DVDD.n15053 DVDD.n7502 2.2505
R18664 DVDD.n15052 DVDD.n15051 2.2505
R18665 DVDD.n15049 DVDD.n7503 2.2505
R18666 DVDD.n15047 DVDD.n15045 2.2505
R18667 DVDD.n15044 DVDD.n7505 2.2505
R18668 DVDD.n15043 DVDD.n15042 2.2505
R18669 DVDD.n15040 DVDD.n7506 2.2505
R18670 DVDD.n15038 DVDD.n15036 2.2505
R18671 DVDD.n15035 DVDD.n7508 2.2505
R18672 DVDD.n15034 DVDD.n15033 2.2505
R18673 DVDD.n15031 DVDD.n7509 2.2505
R18674 DVDD.n15029 DVDD.n15027 2.2505
R18675 DVDD.n15026 DVDD.n7511 2.2505
R18676 DVDD.n15025 DVDD.n15024 2.2505
R18677 DVDD.n15022 DVDD.n7512 2.2505
R18678 DVDD.n15020 DVDD.n15018 2.2505
R18679 DVDD.n15017 DVDD.n7514 2.2505
R18680 DVDD.n15016 DVDD.n15015 2.2505
R18681 DVDD.n15013 DVDD.n7515 2.2505
R18682 DVDD.n15011 DVDD.n15009 2.2505
R18683 DVDD.n15008 DVDD.n7517 2.2505
R18684 DVDD.n15007 DVDD.n15006 2.2505
R18685 DVDD.n15004 DVDD.n7518 2.2505
R18686 DVDD.n15002 DVDD.n15000 2.2505
R18687 DVDD.n14999 DVDD.n7520 2.2505
R18688 DVDD.n14998 DVDD.n14997 2.2505
R18689 DVDD.n14995 DVDD.n7521 2.2505
R18690 DVDD.n14993 DVDD.n14991 2.2505
R18691 DVDD.n14990 DVDD.n7523 2.2505
R18692 DVDD.n14989 DVDD.n14988 2.2505
R18693 DVDD.n14986 DVDD.n7524 2.2505
R18694 DVDD.n14984 DVDD.n14982 2.2505
R18695 DVDD.n14981 DVDD.n7526 2.2505
R18696 DVDD.n14980 DVDD.n14979 2.2505
R18697 DVDD.n14977 DVDD.n7527 2.2505
R18698 DVDD.n14975 DVDD.n14973 2.2505
R18699 DVDD.n14972 DVDD.n7529 2.2505
R18700 DVDD.n14971 DVDD.n14970 2.2505
R18701 DVDD.n14968 DVDD.n7530 2.2505
R18702 DVDD.n14966 DVDD.n14964 2.2505
R18703 DVDD.n14963 DVDD.n7532 2.2505
R18704 DVDD.n14962 DVDD.n14961 2.2505
R18705 DVDD.n14959 DVDD.n7533 2.2505
R18706 DVDD.n14957 DVDD.n14955 2.2505
R18707 DVDD.n14954 DVDD.n7535 2.2505
R18708 DVDD.n14953 DVDD.n14952 2.2505
R18709 DVDD.n14950 DVDD.n7536 2.2505
R18710 DVDD.n14948 DVDD.n14946 2.2505
R18711 DVDD.n14945 DVDD.n7538 2.2505
R18712 DVDD.n14944 DVDD.n14943 2.2505
R18713 DVDD.n14941 DVDD.n7539 2.2505
R18714 DVDD.n14939 DVDD.n14937 2.2505
R18715 DVDD.n14936 DVDD.n7541 2.2505
R18716 DVDD.n14935 DVDD.n14934 2.2505
R18717 DVDD.n14932 DVDD.n7542 2.2505
R18718 DVDD.n14930 DVDD.n14928 2.2505
R18719 DVDD.n14927 DVDD.n7544 2.2505
R18720 DVDD.n14926 DVDD.n14925 2.2505
R18721 DVDD.n14923 DVDD.n7545 2.2505
R18722 DVDD.n14921 DVDD.n14919 2.2505
R18723 DVDD.n14918 DVDD.n7547 2.2505
R18724 DVDD.n14917 DVDD.n14916 2.2505
R18725 DVDD.n14914 DVDD.n7548 2.2505
R18726 DVDD.n14912 DVDD.n14910 2.2505
R18727 DVDD.n14909 DVDD.n7550 2.2505
R18728 DVDD.n14908 DVDD.n14907 2.2505
R18729 DVDD.n14905 DVDD.n7551 2.2505
R18730 DVDD.n14903 DVDD.n14901 2.2505
R18731 DVDD.n14900 DVDD.n7553 2.2505
R18732 DVDD.n14899 DVDD.n14898 2.2505
R18733 DVDD.n14896 DVDD.n7554 2.2505
R18734 DVDD.n14894 DVDD.n14892 2.2505
R18735 DVDD.n14891 DVDD.n7556 2.2505
R18736 DVDD.n14890 DVDD.n14889 2.2505
R18737 DVDD.n14887 DVDD.n7557 2.2505
R18738 DVDD.n14885 DVDD.n14883 2.2505
R18739 DVDD.n14882 DVDD.n7559 2.2505
R18740 DVDD.n14881 DVDD.n14880 2.2505
R18741 DVDD.n14878 DVDD.n7560 2.2505
R18742 DVDD.n14876 DVDD.n14874 2.2505
R18743 DVDD.n14873 DVDD.n7562 2.2505
R18744 DVDD.n14872 DVDD.n14871 2.2505
R18745 DVDD.n14870 DVDD.n7457 2.2505
R18746 DVDD.n15058 DVDD.n7457 2.2505
R18747 DVDD.n14871 DVDD.n7455 2.2505
R18748 DVDD.n7562 DVDD.n7561 2.2505
R18749 DVDD.n14876 DVDD.n14875 2.2505
R18750 DVDD.n14878 DVDD.n14877 2.2505
R18751 DVDD.n14880 DVDD.n14879 2.2505
R18752 DVDD.n7559 DVDD.n7558 2.2505
R18753 DVDD.n14885 DVDD.n14884 2.2505
R18754 DVDD.n14887 DVDD.n14886 2.2505
R18755 DVDD.n14889 DVDD.n14888 2.2505
R18756 DVDD.n7556 DVDD.n7555 2.2505
R18757 DVDD.n14894 DVDD.n14893 2.2505
R18758 DVDD.n14896 DVDD.n14895 2.2505
R18759 DVDD.n14898 DVDD.n14897 2.2505
R18760 DVDD.n7553 DVDD.n7552 2.2505
R18761 DVDD.n14903 DVDD.n14902 2.2505
R18762 DVDD.n14905 DVDD.n14904 2.2505
R18763 DVDD.n14907 DVDD.n14906 2.2505
R18764 DVDD.n7550 DVDD.n7549 2.2505
R18765 DVDD.n14912 DVDD.n14911 2.2505
R18766 DVDD.n14914 DVDD.n14913 2.2505
R18767 DVDD.n14916 DVDD.n14915 2.2505
R18768 DVDD.n7547 DVDD.n7546 2.2505
R18769 DVDD.n14921 DVDD.n14920 2.2505
R18770 DVDD.n14923 DVDD.n14922 2.2505
R18771 DVDD.n14925 DVDD.n14924 2.2505
R18772 DVDD.n7544 DVDD.n7543 2.2505
R18773 DVDD.n14930 DVDD.n14929 2.2505
R18774 DVDD.n14932 DVDD.n14931 2.2505
R18775 DVDD.n14934 DVDD.n14933 2.2505
R18776 DVDD.n7541 DVDD.n7540 2.2505
R18777 DVDD.n14939 DVDD.n14938 2.2505
R18778 DVDD.n14941 DVDD.n14940 2.2505
R18779 DVDD.n14943 DVDD.n14942 2.2505
R18780 DVDD.n7538 DVDD.n7537 2.2505
R18781 DVDD.n14948 DVDD.n14947 2.2505
R18782 DVDD.n14950 DVDD.n14949 2.2505
R18783 DVDD.n14952 DVDD.n14951 2.2505
R18784 DVDD.n7535 DVDD.n7534 2.2505
R18785 DVDD.n14957 DVDD.n14956 2.2505
R18786 DVDD.n14959 DVDD.n14958 2.2505
R18787 DVDD.n14961 DVDD.n14960 2.2505
R18788 DVDD.n7532 DVDD.n7531 2.2505
R18789 DVDD.n14966 DVDD.n14965 2.2505
R18790 DVDD.n14968 DVDD.n14967 2.2505
R18791 DVDD.n14970 DVDD.n14969 2.2505
R18792 DVDD.n7529 DVDD.n7528 2.2505
R18793 DVDD.n14975 DVDD.n14974 2.2505
R18794 DVDD.n14977 DVDD.n14976 2.2505
R18795 DVDD.n14979 DVDD.n14978 2.2505
R18796 DVDD.n7526 DVDD.n7525 2.2505
R18797 DVDD.n14984 DVDD.n14983 2.2505
R18798 DVDD.n14986 DVDD.n14985 2.2505
R18799 DVDD.n14988 DVDD.n14987 2.2505
R18800 DVDD.n7523 DVDD.n7522 2.2505
R18801 DVDD.n14993 DVDD.n14992 2.2505
R18802 DVDD.n14995 DVDD.n14994 2.2505
R18803 DVDD.n14997 DVDD.n14996 2.2505
R18804 DVDD.n7520 DVDD.n7519 2.2505
R18805 DVDD.n15002 DVDD.n15001 2.2505
R18806 DVDD.n15004 DVDD.n15003 2.2505
R18807 DVDD.n15006 DVDD.n15005 2.2505
R18808 DVDD.n7517 DVDD.n7516 2.2505
R18809 DVDD.n15011 DVDD.n15010 2.2505
R18810 DVDD.n15013 DVDD.n15012 2.2505
R18811 DVDD.n15015 DVDD.n15014 2.2505
R18812 DVDD.n7514 DVDD.n7513 2.2505
R18813 DVDD.n15020 DVDD.n15019 2.2505
R18814 DVDD.n15022 DVDD.n15021 2.2505
R18815 DVDD.n15024 DVDD.n15023 2.2505
R18816 DVDD.n7511 DVDD.n7510 2.2505
R18817 DVDD.n15029 DVDD.n15028 2.2505
R18818 DVDD.n15031 DVDD.n15030 2.2505
R18819 DVDD.n15033 DVDD.n15032 2.2505
R18820 DVDD.n7508 DVDD.n7507 2.2505
R18821 DVDD.n15038 DVDD.n15037 2.2505
R18822 DVDD.n15040 DVDD.n15039 2.2505
R18823 DVDD.n15042 DVDD.n15041 2.2505
R18824 DVDD.n7505 DVDD.n7504 2.2505
R18825 DVDD.n15047 DVDD.n15046 2.2505
R18826 DVDD.n15049 DVDD.n15048 2.2505
R18827 DVDD.n15051 DVDD.n15050 2.2505
R18828 DVDD.n7502 DVDD.n7501 2.2505
R18829 DVDD.n15056 DVDD.n15055 2.2505
R18830 DVDD.n14858 DVDD.n7661 2.2505
R18831 DVDD.n9035 DVDD.n7660 2.2505
R18832 DVDD.n9038 DVDD.n9037 2.2505
R18833 DVDD.n9039 DVDD.n9034 2.2505
R18834 DVDD.n9042 DVDD.n9040 2.2505
R18835 DVDD.n9044 DVDD.n9032 2.2505
R18836 DVDD.n9047 DVDD.n9046 2.2505
R18837 DVDD.n9048 DVDD.n9031 2.2505
R18838 DVDD.n9051 DVDD.n9049 2.2505
R18839 DVDD.n9053 DVDD.n9029 2.2505
R18840 DVDD.n9056 DVDD.n9055 2.2505
R18841 DVDD.n9057 DVDD.n9028 2.2505
R18842 DVDD.n9060 DVDD.n9058 2.2505
R18843 DVDD.n9062 DVDD.n9026 2.2505
R18844 DVDD.n9065 DVDD.n9064 2.2505
R18845 DVDD.n9066 DVDD.n9025 2.2505
R18846 DVDD.n9069 DVDD.n9067 2.2505
R18847 DVDD.n9071 DVDD.n9023 2.2505
R18848 DVDD.n9074 DVDD.n9073 2.2505
R18849 DVDD.n9075 DVDD.n9022 2.2505
R18850 DVDD.n9078 DVDD.n9076 2.2505
R18851 DVDD.n9080 DVDD.n9020 2.2505
R18852 DVDD.n9083 DVDD.n9082 2.2505
R18853 DVDD.n9084 DVDD.n9019 2.2505
R18854 DVDD.n9087 DVDD.n9085 2.2505
R18855 DVDD.n9089 DVDD.n9017 2.2505
R18856 DVDD.n9092 DVDD.n9091 2.2505
R18857 DVDD.n9093 DVDD.n9016 2.2505
R18858 DVDD.n9096 DVDD.n9094 2.2505
R18859 DVDD.n9098 DVDD.n9014 2.2505
R18860 DVDD.n9101 DVDD.n9100 2.2505
R18861 DVDD.n9102 DVDD.n9013 2.2505
R18862 DVDD.n9105 DVDD.n9103 2.2505
R18863 DVDD.n9107 DVDD.n9011 2.2505
R18864 DVDD.n9110 DVDD.n9109 2.2505
R18865 DVDD.n9111 DVDD.n9010 2.2505
R18866 DVDD.n9114 DVDD.n9112 2.2505
R18867 DVDD.n9116 DVDD.n9008 2.2505
R18868 DVDD.n9119 DVDD.n9118 2.2505
R18869 DVDD.n9120 DVDD.n9007 2.2505
R18870 DVDD.n9123 DVDD.n9121 2.2505
R18871 DVDD.n9125 DVDD.n9005 2.2505
R18872 DVDD.n9128 DVDD.n9127 2.2505
R18873 DVDD.n9129 DVDD.n9004 2.2505
R18874 DVDD.n9132 DVDD.n9130 2.2505
R18875 DVDD.n9134 DVDD.n9002 2.2505
R18876 DVDD.n9137 DVDD.n9136 2.2505
R18877 DVDD.n9138 DVDD.n9001 2.2505
R18878 DVDD.n9141 DVDD.n9139 2.2505
R18879 DVDD.n9143 DVDD.n8999 2.2505
R18880 DVDD.n9146 DVDD.n9145 2.2505
R18881 DVDD.n9147 DVDD.n8998 2.2505
R18882 DVDD.n9150 DVDD.n9148 2.2505
R18883 DVDD.n9152 DVDD.n8996 2.2505
R18884 DVDD.n9155 DVDD.n9154 2.2505
R18885 DVDD.n9156 DVDD.n8995 2.2505
R18886 DVDD.n9159 DVDD.n9157 2.2505
R18887 DVDD.n9161 DVDD.n8993 2.2505
R18888 DVDD.n9164 DVDD.n9163 2.2505
R18889 DVDD.n9165 DVDD.n8992 2.2505
R18890 DVDD.n9168 DVDD.n9166 2.2505
R18891 DVDD.n9170 DVDD.n8990 2.2505
R18892 DVDD.n9173 DVDD.n9172 2.2505
R18893 DVDD.n9174 DVDD.n8989 2.2505
R18894 DVDD.n9177 DVDD.n9175 2.2505
R18895 DVDD.n9179 DVDD.n8987 2.2505
R18896 DVDD.n9182 DVDD.n9181 2.2505
R18897 DVDD.n9183 DVDD.n8986 2.2505
R18898 DVDD.n9186 DVDD.n9184 2.2505
R18899 DVDD.n9188 DVDD.n8984 2.2505
R18900 DVDD.n9191 DVDD.n9190 2.2505
R18901 DVDD.n9192 DVDD.n8983 2.2505
R18902 DVDD.n9195 DVDD.n9193 2.2505
R18903 DVDD.n9197 DVDD.n8981 2.2505
R18904 DVDD.n9200 DVDD.n9199 2.2505
R18905 DVDD.n9201 DVDD.n8980 2.2505
R18906 DVDD.n9204 DVDD.n9202 2.2505
R18907 DVDD.n9206 DVDD.n8978 2.2505
R18908 DVDD.n9209 DVDD.n9208 2.2505
R18909 DVDD.n9210 DVDD.n8977 2.2505
R18910 DVDD.n9213 DVDD.n9211 2.2505
R18911 DVDD.n9215 DVDD.n8975 2.2505
R18912 DVDD.n9217 DVDD.n9216 2.2505
R18913 DVDD.n9218 DVDD.n7614 2.2505
R18914 DVDD.n14861 DVDD.n7614 2.2505
R18915 DVDD.n9216 DVDD.n7612 2.2505
R18916 DVDD.n9215 DVDD.n9214 2.2505
R18917 DVDD.n9213 DVDD.n9212 2.2505
R18918 DVDD.n8977 DVDD.n8976 2.2505
R18919 DVDD.n9208 DVDD.n9207 2.2505
R18920 DVDD.n9206 DVDD.n9205 2.2505
R18921 DVDD.n9204 DVDD.n9203 2.2505
R18922 DVDD.n8980 DVDD.n8979 2.2505
R18923 DVDD.n9199 DVDD.n9198 2.2505
R18924 DVDD.n9197 DVDD.n9196 2.2505
R18925 DVDD.n9195 DVDD.n9194 2.2505
R18926 DVDD.n8983 DVDD.n8982 2.2505
R18927 DVDD.n9190 DVDD.n9189 2.2505
R18928 DVDD.n9188 DVDD.n9187 2.2505
R18929 DVDD.n9186 DVDD.n9185 2.2505
R18930 DVDD.n8986 DVDD.n8985 2.2505
R18931 DVDD.n9181 DVDD.n9180 2.2505
R18932 DVDD.n9179 DVDD.n9178 2.2505
R18933 DVDD.n9177 DVDD.n9176 2.2505
R18934 DVDD.n8989 DVDD.n8988 2.2505
R18935 DVDD.n9172 DVDD.n9171 2.2505
R18936 DVDD.n9170 DVDD.n9169 2.2505
R18937 DVDD.n9168 DVDD.n9167 2.2505
R18938 DVDD.n8992 DVDD.n8991 2.2505
R18939 DVDD.n9163 DVDD.n9162 2.2505
R18940 DVDD.n9161 DVDD.n9160 2.2505
R18941 DVDD.n9159 DVDD.n9158 2.2505
R18942 DVDD.n8995 DVDD.n8994 2.2505
R18943 DVDD.n9154 DVDD.n9153 2.2505
R18944 DVDD.n9152 DVDD.n9151 2.2505
R18945 DVDD.n9150 DVDD.n9149 2.2505
R18946 DVDD.n8998 DVDD.n8997 2.2505
R18947 DVDD.n9145 DVDD.n9144 2.2505
R18948 DVDD.n9143 DVDD.n9142 2.2505
R18949 DVDD.n9141 DVDD.n9140 2.2505
R18950 DVDD.n9001 DVDD.n9000 2.2505
R18951 DVDD.n9136 DVDD.n9135 2.2505
R18952 DVDD.n9134 DVDD.n9133 2.2505
R18953 DVDD.n9132 DVDD.n9131 2.2505
R18954 DVDD.n9004 DVDD.n9003 2.2505
R18955 DVDD.n9127 DVDD.n9126 2.2505
R18956 DVDD.n9125 DVDD.n9124 2.2505
R18957 DVDD.n9123 DVDD.n9122 2.2505
R18958 DVDD.n9007 DVDD.n9006 2.2505
R18959 DVDD.n9118 DVDD.n9117 2.2505
R18960 DVDD.n9116 DVDD.n9115 2.2505
R18961 DVDD.n9114 DVDD.n9113 2.2505
R18962 DVDD.n9010 DVDD.n9009 2.2505
R18963 DVDD.n9109 DVDD.n9108 2.2505
R18964 DVDD.n9107 DVDD.n9106 2.2505
R18965 DVDD.n9105 DVDD.n9104 2.2505
R18966 DVDD.n9013 DVDD.n9012 2.2505
R18967 DVDD.n9100 DVDD.n9099 2.2505
R18968 DVDD.n9098 DVDD.n9097 2.2505
R18969 DVDD.n9096 DVDD.n9095 2.2505
R18970 DVDD.n9016 DVDD.n9015 2.2505
R18971 DVDD.n9091 DVDD.n9090 2.2505
R18972 DVDD.n9089 DVDD.n9088 2.2505
R18973 DVDD.n9087 DVDD.n9086 2.2505
R18974 DVDD.n9019 DVDD.n9018 2.2505
R18975 DVDD.n9082 DVDD.n9081 2.2505
R18976 DVDD.n9080 DVDD.n9079 2.2505
R18977 DVDD.n9078 DVDD.n9077 2.2505
R18978 DVDD.n9022 DVDD.n9021 2.2505
R18979 DVDD.n9073 DVDD.n9072 2.2505
R18980 DVDD.n9071 DVDD.n9070 2.2505
R18981 DVDD.n9069 DVDD.n9068 2.2505
R18982 DVDD.n9025 DVDD.n9024 2.2505
R18983 DVDD.n9064 DVDD.n9063 2.2505
R18984 DVDD.n9062 DVDD.n9061 2.2505
R18985 DVDD.n9060 DVDD.n9059 2.2505
R18986 DVDD.n9028 DVDD.n9027 2.2505
R18987 DVDD.n9055 DVDD.n9054 2.2505
R18988 DVDD.n9053 DVDD.n9052 2.2505
R18989 DVDD.n9051 DVDD.n9050 2.2505
R18990 DVDD.n9031 DVDD.n9030 2.2505
R18991 DVDD.n9046 DVDD.n9045 2.2505
R18992 DVDD.n9044 DVDD.n9043 2.2505
R18993 DVDD.n9042 DVDD.n9041 2.2505
R18994 DVDD.n9034 DVDD.n9033 2.2505
R18995 DVDD.n9037 DVDD.n9036 2.2505
R18996 DVDD.n7660 DVDD.n7659 2.2505
R18997 DVDD.n14859 DVDD.n14858 2.2505
R18998 DVDD.n9311 DVDD.n9310 2.2505
R18999 DVDD.n9312 DVDD.n9308 2.2505
R19000 DVDD.n9317 DVDD.n9313 2.2505
R19001 DVDD.n9318 DVDD.n9307 2.2505
R19002 DVDD.n9323 DVDD.n9322 2.2505
R19003 DVDD.n9324 DVDD.n9306 2.2505
R19004 DVDD.n9329 DVDD.n9325 2.2505
R19005 DVDD.n9330 DVDD.n9305 2.2505
R19006 DVDD.n9335 DVDD.n9334 2.2505
R19007 DVDD.n9336 DVDD.n9304 2.2505
R19008 DVDD.n9341 DVDD.n9337 2.2505
R19009 DVDD.n9342 DVDD.n9303 2.2505
R19010 DVDD.n9347 DVDD.n9346 2.2505
R19011 DVDD.n9348 DVDD.n9302 2.2505
R19012 DVDD.n9353 DVDD.n9349 2.2505
R19013 DVDD.n9354 DVDD.n9301 2.2505
R19014 DVDD.n9359 DVDD.n9358 2.2505
R19015 DVDD.n9360 DVDD.n9300 2.2505
R19016 DVDD.n9365 DVDD.n9361 2.2505
R19017 DVDD.n9366 DVDD.n9299 2.2505
R19018 DVDD.n9371 DVDD.n9370 2.2505
R19019 DVDD.n9372 DVDD.n9298 2.2505
R19020 DVDD.n9377 DVDD.n9373 2.2505
R19021 DVDD.n9378 DVDD.n9297 2.2505
R19022 DVDD.n9383 DVDD.n9382 2.2505
R19023 DVDD.n9384 DVDD.n9296 2.2505
R19024 DVDD.n9389 DVDD.n9385 2.2505
R19025 DVDD.n9390 DVDD.n9295 2.2505
R19026 DVDD.n9395 DVDD.n9394 2.2505
R19027 DVDD.n9396 DVDD.n9294 2.2505
R19028 DVDD.n9401 DVDD.n9397 2.2505
R19029 DVDD.n9402 DVDD.n9293 2.2505
R19030 DVDD.n9407 DVDD.n9406 2.2505
R19031 DVDD.n9408 DVDD.n9292 2.2505
R19032 DVDD.n9413 DVDD.n9409 2.2505
R19033 DVDD.n9414 DVDD.n9291 2.2505
R19034 DVDD.n9419 DVDD.n9418 2.2505
R19035 DVDD.n9420 DVDD.n9290 2.2505
R19036 DVDD.n9425 DVDD.n9421 2.2505
R19037 DVDD.n9426 DVDD.n9289 2.2505
R19038 DVDD.n9431 DVDD.n9430 2.2505
R19039 DVDD.n9432 DVDD.n9288 2.2505
R19040 DVDD.n9437 DVDD.n9433 2.2505
R19041 DVDD.n9438 DVDD.n9287 2.2505
R19042 DVDD.n9443 DVDD.n9442 2.2505
R19043 DVDD.n9444 DVDD.n9286 2.2505
R19044 DVDD.n9449 DVDD.n9445 2.2505
R19045 DVDD.n9450 DVDD.n9285 2.2505
R19046 DVDD.n9455 DVDD.n9454 2.2505
R19047 DVDD.n9456 DVDD.n9284 2.2505
R19048 DVDD.n9461 DVDD.n9457 2.2505
R19049 DVDD.n9462 DVDD.n9283 2.2505
R19050 DVDD.n9467 DVDD.n9466 2.2505
R19051 DVDD.n9468 DVDD.n9282 2.2505
R19052 DVDD.n9473 DVDD.n9469 2.2505
R19053 DVDD.n9474 DVDD.n9281 2.2505
R19054 DVDD.n9479 DVDD.n9478 2.2505
R19055 DVDD.n9480 DVDD.n9280 2.2505
R19056 DVDD.n9485 DVDD.n9481 2.2505
R19057 DVDD.n9486 DVDD.n9279 2.2505
R19058 DVDD.n9491 DVDD.n9490 2.2505
R19059 DVDD.n9492 DVDD.n9278 2.2505
R19060 DVDD.n9497 DVDD.n9493 2.2505
R19061 DVDD.n9498 DVDD.n9277 2.2505
R19062 DVDD.n9503 DVDD.n9502 2.2505
R19063 DVDD.n9504 DVDD.n9276 2.2505
R19064 DVDD.n9509 DVDD.n9505 2.2505
R19065 DVDD.n9510 DVDD.n9275 2.2505
R19066 DVDD.n9515 DVDD.n9514 2.2505
R19067 DVDD.n9516 DVDD.n9274 2.2505
R19068 DVDD.n9521 DVDD.n9517 2.2505
R19069 DVDD.n9522 DVDD.n9273 2.2505
R19070 DVDD.n9527 DVDD.n9526 2.2505
R19071 DVDD.n9528 DVDD.n9272 2.2505
R19072 DVDD.n9533 DVDD.n9529 2.2505
R19073 DVDD.n9534 DVDD.n9271 2.2505
R19074 DVDD.n9539 DVDD.n9538 2.2505
R19075 DVDD.n9540 DVDD.n9270 2.2505
R19076 DVDD.n9545 DVDD.n9541 2.2505
R19077 DVDD.n9546 DVDD.n9269 2.2505
R19078 DVDD.n9551 DVDD.n9550 2.2505
R19079 DVDD.n9552 DVDD.n9268 2.2505
R19080 DVDD.n9554 DVDD.n9553 2.2505
R19081 DVDD.n9555 DVDD.n9265 2.2505
R19082 DVDD.n9556 DVDD.n9555 2.2505
R19083 DVDD.n9554 DVDD.n9264 2.2505
R19084 DVDD.n9268 DVDD.n9267 2.2505
R19085 DVDD.n9550 DVDD.n9549 2.2505
R19086 DVDD.n9547 DVDD.n9546 2.2505
R19087 DVDD.n9545 DVDD.n9544 2.2505
R19088 DVDD.n9542 DVDD.n9270 2.2505
R19089 DVDD.n9538 DVDD.n9537 2.2505
R19090 DVDD.n9535 DVDD.n9534 2.2505
R19091 DVDD.n9533 DVDD.n9532 2.2505
R19092 DVDD.n9530 DVDD.n9272 2.2505
R19093 DVDD.n9526 DVDD.n9525 2.2505
R19094 DVDD.n9523 DVDD.n9522 2.2505
R19095 DVDD.n9521 DVDD.n9520 2.2505
R19096 DVDD.n9518 DVDD.n9274 2.2505
R19097 DVDD.n9514 DVDD.n9513 2.2505
R19098 DVDD.n9511 DVDD.n9510 2.2505
R19099 DVDD.n9509 DVDD.n9508 2.2505
R19100 DVDD.n9506 DVDD.n9276 2.2505
R19101 DVDD.n9502 DVDD.n9501 2.2505
R19102 DVDD.n9499 DVDD.n9498 2.2505
R19103 DVDD.n9497 DVDD.n9496 2.2505
R19104 DVDD.n9494 DVDD.n9278 2.2505
R19105 DVDD.n9490 DVDD.n9489 2.2505
R19106 DVDD.n9487 DVDD.n9486 2.2505
R19107 DVDD.n9485 DVDD.n9484 2.2505
R19108 DVDD.n9482 DVDD.n9280 2.2505
R19109 DVDD.n9478 DVDD.n9477 2.2505
R19110 DVDD.n9475 DVDD.n9474 2.2505
R19111 DVDD.n9473 DVDD.n9472 2.2505
R19112 DVDD.n9470 DVDD.n9282 2.2505
R19113 DVDD.n9466 DVDD.n9465 2.2505
R19114 DVDD.n9463 DVDD.n9462 2.2505
R19115 DVDD.n9461 DVDD.n9460 2.2505
R19116 DVDD.n9458 DVDD.n9284 2.2505
R19117 DVDD.n9454 DVDD.n9453 2.2505
R19118 DVDD.n9451 DVDD.n9450 2.2505
R19119 DVDD.n9449 DVDD.n9448 2.2505
R19120 DVDD.n9446 DVDD.n9286 2.2505
R19121 DVDD.n9442 DVDD.n9441 2.2505
R19122 DVDD.n9439 DVDD.n9438 2.2505
R19123 DVDD.n9437 DVDD.n9436 2.2505
R19124 DVDD.n9434 DVDD.n9288 2.2505
R19125 DVDD.n9430 DVDD.n9429 2.2505
R19126 DVDD.n9427 DVDD.n9426 2.2505
R19127 DVDD.n9425 DVDD.n9424 2.2505
R19128 DVDD.n9422 DVDD.n9290 2.2505
R19129 DVDD.n9418 DVDD.n9417 2.2505
R19130 DVDD.n9415 DVDD.n9414 2.2505
R19131 DVDD.n9413 DVDD.n9412 2.2505
R19132 DVDD.n9410 DVDD.n9292 2.2505
R19133 DVDD.n9406 DVDD.n9405 2.2505
R19134 DVDD.n9403 DVDD.n9402 2.2505
R19135 DVDD.n9401 DVDD.n9400 2.2505
R19136 DVDD.n9398 DVDD.n9294 2.2505
R19137 DVDD.n9394 DVDD.n9393 2.2505
R19138 DVDD.n9391 DVDD.n9390 2.2505
R19139 DVDD.n9389 DVDD.n9388 2.2505
R19140 DVDD.n9386 DVDD.n9296 2.2505
R19141 DVDD.n9382 DVDD.n9381 2.2505
R19142 DVDD.n9379 DVDD.n9378 2.2505
R19143 DVDD.n9377 DVDD.n9376 2.2505
R19144 DVDD.n9374 DVDD.n9298 2.2505
R19145 DVDD.n9370 DVDD.n9369 2.2505
R19146 DVDD.n9367 DVDD.n9366 2.2505
R19147 DVDD.n9365 DVDD.n9364 2.2505
R19148 DVDD.n9362 DVDD.n9300 2.2505
R19149 DVDD.n9358 DVDD.n9357 2.2505
R19150 DVDD.n9355 DVDD.n9354 2.2505
R19151 DVDD.n9353 DVDD.n9352 2.2505
R19152 DVDD.n9350 DVDD.n9302 2.2505
R19153 DVDD.n9346 DVDD.n9345 2.2505
R19154 DVDD.n9343 DVDD.n9342 2.2505
R19155 DVDD.n9341 DVDD.n9340 2.2505
R19156 DVDD.n9338 DVDD.n9304 2.2505
R19157 DVDD.n9334 DVDD.n9333 2.2505
R19158 DVDD.n9331 DVDD.n9330 2.2505
R19159 DVDD.n9329 DVDD.n9328 2.2505
R19160 DVDD.n9326 DVDD.n9306 2.2505
R19161 DVDD.n9322 DVDD.n9321 2.2505
R19162 DVDD.n9319 DVDD.n9318 2.2505
R19163 DVDD.n9317 DVDD.n9316 2.2505
R19164 DVDD.n9314 DVDD.n9308 2.2505
R19165 DVDD.n9310 DVDD.n9309 2.2505
R19166 DVDD.n14835 DVDD.n8023 2.2505
R19167 DVDD.n8022 DVDD.n7778 2.2505
R19168 DVDD.n8021 DVDD.n8020 2.2505
R19169 DVDD.n8018 DVDD.n7779 2.2505
R19170 DVDD.n8016 DVDD.n8014 2.2505
R19171 DVDD.n8013 DVDD.n7781 2.2505
R19172 DVDD.n8012 DVDD.n8011 2.2505
R19173 DVDD.n8009 DVDD.n7782 2.2505
R19174 DVDD.n8007 DVDD.n8005 2.2505
R19175 DVDD.n8004 DVDD.n7784 2.2505
R19176 DVDD.n8003 DVDD.n8002 2.2505
R19177 DVDD.n8000 DVDD.n7785 2.2505
R19178 DVDD.n7998 DVDD.n7996 2.2505
R19179 DVDD.n7995 DVDD.n7787 2.2505
R19180 DVDD.n7994 DVDD.n7993 2.2505
R19181 DVDD.n7991 DVDD.n7788 2.2505
R19182 DVDD.n7989 DVDD.n7987 2.2505
R19183 DVDD.n7986 DVDD.n7790 2.2505
R19184 DVDD.n7985 DVDD.n7984 2.2505
R19185 DVDD.n7982 DVDD.n7791 2.2505
R19186 DVDD.n7980 DVDD.n7978 2.2505
R19187 DVDD.n7977 DVDD.n7793 2.2505
R19188 DVDD.n7976 DVDD.n7975 2.2505
R19189 DVDD.n7973 DVDD.n7794 2.2505
R19190 DVDD.n7971 DVDD.n7969 2.2505
R19191 DVDD.n7968 DVDD.n7796 2.2505
R19192 DVDD.n7967 DVDD.n7966 2.2505
R19193 DVDD.n7964 DVDD.n7797 2.2505
R19194 DVDD.n7962 DVDD.n7960 2.2505
R19195 DVDD.n7959 DVDD.n7799 2.2505
R19196 DVDD.n7958 DVDD.n7957 2.2505
R19197 DVDD.n7955 DVDD.n7800 2.2505
R19198 DVDD.n7953 DVDD.n7951 2.2505
R19199 DVDD.n7950 DVDD.n7802 2.2505
R19200 DVDD.n7949 DVDD.n7948 2.2505
R19201 DVDD.n7946 DVDD.n7803 2.2505
R19202 DVDD.n7944 DVDD.n7942 2.2505
R19203 DVDD.n7941 DVDD.n7805 2.2505
R19204 DVDD.n7940 DVDD.n7939 2.2505
R19205 DVDD.n7937 DVDD.n7806 2.2505
R19206 DVDD.n7935 DVDD.n7933 2.2505
R19207 DVDD.n7932 DVDD.n7808 2.2505
R19208 DVDD.n7931 DVDD.n7930 2.2505
R19209 DVDD.n7928 DVDD.n7809 2.2505
R19210 DVDD.n7926 DVDD.n7924 2.2505
R19211 DVDD.n7923 DVDD.n7811 2.2505
R19212 DVDD.n7922 DVDD.n7921 2.2505
R19213 DVDD.n7919 DVDD.n7812 2.2505
R19214 DVDD.n7917 DVDD.n7915 2.2505
R19215 DVDD.n7914 DVDD.n7814 2.2505
R19216 DVDD.n7913 DVDD.n7912 2.2505
R19217 DVDD.n7910 DVDD.n7815 2.2505
R19218 DVDD.n7908 DVDD.n7906 2.2505
R19219 DVDD.n7905 DVDD.n7817 2.2505
R19220 DVDD.n7904 DVDD.n7903 2.2505
R19221 DVDD.n7901 DVDD.n7818 2.2505
R19222 DVDD.n7899 DVDD.n7897 2.2505
R19223 DVDD.n7896 DVDD.n7820 2.2505
R19224 DVDD.n7895 DVDD.n7894 2.2505
R19225 DVDD.n7892 DVDD.n7821 2.2505
R19226 DVDD.n7890 DVDD.n7888 2.2505
R19227 DVDD.n7887 DVDD.n7823 2.2505
R19228 DVDD.n7886 DVDD.n7885 2.2505
R19229 DVDD.n7883 DVDD.n7824 2.2505
R19230 DVDD.n7881 DVDD.n7879 2.2505
R19231 DVDD.n7878 DVDD.n7826 2.2505
R19232 DVDD.n7877 DVDD.n7876 2.2505
R19233 DVDD.n7874 DVDD.n7827 2.2505
R19234 DVDD.n7872 DVDD.n7870 2.2505
R19235 DVDD.n7869 DVDD.n7829 2.2505
R19236 DVDD.n7868 DVDD.n7867 2.2505
R19237 DVDD.n7865 DVDD.n7830 2.2505
R19238 DVDD.n7863 DVDD.n7861 2.2505
R19239 DVDD.n7860 DVDD.n7832 2.2505
R19240 DVDD.n7859 DVDD.n7858 2.2505
R19241 DVDD.n7856 DVDD.n7833 2.2505
R19242 DVDD.n7854 DVDD.n7852 2.2505
R19243 DVDD.n7851 DVDD.n7835 2.2505
R19244 DVDD.n7850 DVDD.n7849 2.2505
R19245 DVDD.n7847 DVDD.n7836 2.2505
R19246 DVDD.n7845 DVDD.n7843 2.2505
R19247 DVDD.n7842 DVDD.n7838 2.2505
R19248 DVDD.n7841 DVDD.n7840 2.2505
R19249 DVDD.n7839 DVDD.n7732 2.2505
R19250 DVDD.n14838 DVDD.n7732 2.2505
R19251 DVDD.n7840 DVDD.n7731 2.2505
R19252 DVDD.n7838 DVDD.n7837 2.2505
R19253 DVDD.n7845 DVDD.n7844 2.2505
R19254 DVDD.n7847 DVDD.n7846 2.2505
R19255 DVDD.n7849 DVDD.n7848 2.2505
R19256 DVDD.n7835 DVDD.n7834 2.2505
R19257 DVDD.n7854 DVDD.n7853 2.2505
R19258 DVDD.n7856 DVDD.n7855 2.2505
R19259 DVDD.n7858 DVDD.n7857 2.2505
R19260 DVDD.n7832 DVDD.n7831 2.2505
R19261 DVDD.n7863 DVDD.n7862 2.2505
R19262 DVDD.n7865 DVDD.n7864 2.2505
R19263 DVDD.n7867 DVDD.n7866 2.2505
R19264 DVDD.n7829 DVDD.n7828 2.2505
R19265 DVDD.n7872 DVDD.n7871 2.2505
R19266 DVDD.n7874 DVDD.n7873 2.2505
R19267 DVDD.n7876 DVDD.n7875 2.2505
R19268 DVDD.n7826 DVDD.n7825 2.2505
R19269 DVDD.n7881 DVDD.n7880 2.2505
R19270 DVDD.n7883 DVDD.n7882 2.2505
R19271 DVDD.n7885 DVDD.n7884 2.2505
R19272 DVDD.n7823 DVDD.n7822 2.2505
R19273 DVDD.n7890 DVDD.n7889 2.2505
R19274 DVDD.n7892 DVDD.n7891 2.2505
R19275 DVDD.n7894 DVDD.n7893 2.2505
R19276 DVDD.n7820 DVDD.n7819 2.2505
R19277 DVDD.n7899 DVDD.n7898 2.2505
R19278 DVDD.n7901 DVDD.n7900 2.2505
R19279 DVDD.n7903 DVDD.n7902 2.2505
R19280 DVDD.n7817 DVDD.n7816 2.2505
R19281 DVDD.n7908 DVDD.n7907 2.2505
R19282 DVDD.n7910 DVDD.n7909 2.2505
R19283 DVDD.n7912 DVDD.n7911 2.2505
R19284 DVDD.n7814 DVDD.n7813 2.2505
R19285 DVDD.n7917 DVDD.n7916 2.2505
R19286 DVDD.n7919 DVDD.n7918 2.2505
R19287 DVDD.n7921 DVDD.n7920 2.2505
R19288 DVDD.n7811 DVDD.n7810 2.2505
R19289 DVDD.n7926 DVDD.n7925 2.2505
R19290 DVDD.n7928 DVDD.n7927 2.2505
R19291 DVDD.n7930 DVDD.n7929 2.2505
R19292 DVDD.n7808 DVDD.n7807 2.2505
R19293 DVDD.n7935 DVDD.n7934 2.2505
R19294 DVDD.n7937 DVDD.n7936 2.2505
R19295 DVDD.n7939 DVDD.n7938 2.2505
R19296 DVDD.n7805 DVDD.n7804 2.2505
R19297 DVDD.n7944 DVDD.n7943 2.2505
R19298 DVDD.n7946 DVDD.n7945 2.2505
R19299 DVDD.n7948 DVDD.n7947 2.2505
R19300 DVDD.n7802 DVDD.n7801 2.2505
R19301 DVDD.n7953 DVDD.n7952 2.2505
R19302 DVDD.n7955 DVDD.n7954 2.2505
R19303 DVDD.n7957 DVDD.n7956 2.2505
R19304 DVDD.n7799 DVDD.n7798 2.2505
R19305 DVDD.n7962 DVDD.n7961 2.2505
R19306 DVDD.n7964 DVDD.n7963 2.2505
R19307 DVDD.n7966 DVDD.n7965 2.2505
R19308 DVDD.n7796 DVDD.n7795 2.2505
R19309 DVDD.n7971 DVDD.n7970 2.2505
R19310 DVDD.n7973 DVDD.n7972 2.2505
R19311 DVDD.n7975 DVDD.n7974 2.2505
R19312 DVDD.n7793 DVDD.n7792 2.2505
R19313 DVDD.n7980 DVDD.n7979 2.2505
R19314 DVDD.n7982 DVDD.n7981 2.2505
R19315 DVDD.n7984 DVDD.n7983 2.2505
R19316 DVDD.n7790 DVDD.n7789 2.2505
R19317 DVDD.n7989 DVDD.n7988 2.2505
R19318 DVDD.n7991 DVDD.n7990 2.2505
R19319 DVDD.n7993 DVDD.n7992 2.2505
R19320 DVDD.n7787 DVDD.n7786 2.2505
R19321 DVDD.n7998 DVDD.n7997 2.2505
R19322 DVDD.n8000 DVDD.n7999 2.2505
R19323 DVDD.n8002 DVDD.n8001 2.2505
R19324 DVDD.n7784 DVDD.n7783 2.2505
R19325 DVDD.n8007 DVDD.n8006 2.2505
R19326 DVDD.n8009 DVDD.n8008 2.2505
R19327 DVDD.n8011 DVDD.n8010 2.2505
R19328 DVDD.n7781 DVDD.n7780 2.2505
R19329 DVDD.n8016 DVDD.n8015 2.2505
R19330 DVDD.n8018 DVDD.n8017 2.2505
R19331 DVDD.n8020 DVDD.n8019 2.2505
R19332 DVDD.n7778 DVDD.n7777 2.2505
R19333 DVDD.n14836 DVDD.n14835 2.2505
R19334 DVDD.n8088 DVDD.n8038 2.2505
R19335 DVDD.n14821 DVDD.n14820 2.2505
R19336 DVDD.n14819 DVDD.n8090 2.2505
R19337 DVDD.n14818 DVDD.n14817 2.2505
R19338 DVDD.n14813 DVDD.n8091 2.2505
R19339 DVDD.n14809 DVDD.n14808 2.2505
R19340 DVDD.n14807 DVDD.n8092 2.2505
R19341 DVDD.n14806 DVDD.n14805 2.2505
R19342 DVDD.n14801 DVDD.n8093 2.2505
R19343 DVDD.n14797 DVDD.n14796 2.2505
R19344 DVDD.n14795 DVDD.n8094 2.2505
R19345 DVDD.n14794 DVDD.n14793 2.2505
R19346 DVDD.n14789 DVDD.n8095 2.2505
R19347 DVDD.n14785 DVDD.n14784 2.2505
R19348 DVDD.n14783 DVDD.n8096 2.2505
R19349 DVDD.n14782 DVDD.n14781 2.2505
R19350 DVDD.n14777 DVDD.n8097 2.2505
R19351 DVDD.n14773 DVDD.n14772 2.2505
R19352 DVDD.n14771 DVDD.n8098 2.2505
R19353 DVDD.n14770 DVDD.n14769 2.2505
R19354 DVDD.n14765 DVDD.n8099 2.2505
R19355 DVDD.n14761 DVDD.n14760 2.2505
R19356 DVDD.n14759 DVDD.n8100 2.2505
R19357 DVDD.n14758 DVDD.n14757 2.2505
R19358 DVDD.n14753 DVDD.n8101 2.2505
R19359 DVDD.n14749 DVDD.n14748 2.2505
R19360 DVDD.n14747 DVDD.n8102 2.2505
R19361 DVDD.n14746 DVDD.n14745 2.2505
R19362 DVDD.n14741 DVDD.n8103 2.2505
R19363 DVDD.n14737 DVDD.n14736 2.2505
R19364 DVDD.n14735 DVDD.n8104 2.2505
R19365 DVDD.n14734 DVDD.n14733 2.2505
R19366 DVDD.n14729 DVDD.n8105 2.2505
R19367 DVDD.n14725 DVDD.n14724 2.2505
R19368 DVDD.n14723 DVDD.n8106 2.2505
R19369 DVDD.n14722 DVDD.n14721 2.2505
R19370 DVDD.n14717 DVDD.n8107 2.2505
R19371 DVDD.n14713 DVDD.n14712 2.2505
R19372 DVDD.n14711 DVDD.n8108 2.2505
R19373 DVDD.n14710 DVDD.n14709 2.2505
R19374 DVDD.n14705 DVDD.n8109 2.2505
R19375 DVDD.n14701 DVDD.n14700 2.2505
R19376 DVDD.n14699 DVDD.n8110 2.2505
R19377 DVDD.n14698 DVDD.n14697 2.2505
R19378 DVDD.n14693 DVDD.n8111 2.2505
R19379 DVDD.n14689 DVDD.n14688 2.2505
R19380 DVDD.n14687 DVDD.n8112 2.2505
R19381 DVDD.n14686 DVDD.n14685 2.2505
R19382 DVDD.n14681 DVDD.n8113 2.2505
R19383 DVDD.n14677 DVDD.n14676 2.2505
R19384 DVDD.n14675 DVDD.n8114 2.2505
R19385 DVDD.n14674 DVDD.n14673 2.2505
R19386 DVDD.n14669 DVDD.n8115 2.2505
R19387 DVDD.n14665 DVDD.n14664 2.2505
R19388 DVDD.n14663 DVDD.n8116 2.2505
R19389 DVDD.n14662 DVDD.n14661 2.2505
R19390 DVDD.n14657 DVDD.n8117 2.2505
R19391 DVDD.n14653 DVDD.n14652 2.2505
R19392 DVDD.n14651 DVDD.n8118 2.2505
R19393 DVDD.n14650 DVDD.n14649 2.2505
R19394 DVDD.n14645 DVDD.n8119 2.2505
R19395 DVDD.n14641 DVDD.n14640 2.2505
R19396 DVDD.n14639 DVDD.n8120 2.2505
R19397 DVDD.n14638 DVDD.n14637 2.2505
R19398 DVDD.n14633 DVDD.n8121 2.2505
R19399 DVDD.n14629 DVDD.n14628 2.2505
R19400 DVDD.n14627 DVDD.n8122 2.2505
R19401 DVDD.n14626 DVDD.n14625 2.2505
R19402 DVDD.n14621 DVDD.n8123 2.2505
R19403 DVDD.n14617 DVDD.n14616 2.2505
R19404 DVDD.n14615 DVDD.n8124 2.2505
R19405 DVDD.n14614 DVDD.n14613 2.2505
R19406 DVDD.n14609 DVDD.n8125 2.2505
R19407 DVDD.n14605 DVDD.n14604 2.2505
R19408 DVDD.n14603 DVDD.n8126 2.2505
R19409 DVDD.n14602 DVDD.n14601 2.2505
R19410 DVDD.n14597 DVDD.n8127 2.2505
R19411 DVDD.n14593 DVDD.n14592 2.2505
R19412 DVDD.n14591 DVDD.n8128 2.2505
R19413 DVDD.n14590 DVDD.n14589 2.2505
R19414 DVDD.n14585 DVDD.n8129 2.2505
R19415 DVDD.n14581 DVDD.n14580 2.2505
R19416 DVDD.n14579 DVDD.n8132 2.2505
R19417 DVDD.n14578 DVDD.n14577 2.2505
R19418 DVDD.n14577 DVDD.n8086 2.2505
R19419 DVDD.n8132 DVDD.n8131 2.2505
R19420 DVDD.n14582 DVDD.n14581 2.2505
R19421 DVDD.n14585 DVDD.n14584 2.2505
R19422 DVDD.n14589 DVDD.n14588 2.2505
R19423 DVDD.n14586 DVDD.n8128 2.2505
R19424 DVDD.n14594 DVDD.n14593 2.2505
R19425 DVDD.n14597 DVDD.n14596 2.2505
R19426 DVDD.n14601 DVDD.n14600 2.2505
R19427 DVDD.n14598 DVDD.n8126 2.2505
R19428 DVDD.n14606 DVDD.n14605 2.2505
R19429 DVDD.n14609 DVDD.n14608 2.2505
R19430 DVDD.n14613 DVDD.n14612 2.2505
R19431 DVDD.n14610 DVDD.n8124 2.2505
R19432 DVDD.n14618 DVDD.n14617 2.2505
R19433 DVDD.n14621 DVDD.n14620 2.2505
R19434 DVDD.n14625 DVDD.n14624 2.2505
R19435 DVDD.n14622 DVDD.n8122 2.2505
R19436 DVDD.n14630 DVDD.n14629 2.2505
R19437 DVDD.n14633 DVDD.n14632 2.2505
R19438 DVDD.n14637 DVDD.n14636 2.2505
R19439 DVDD.n14634 DVDD.n8120 2.2505
R19440 DVDD.n14642 DVDD.n14641 2.2505
R19441 DVDD.n14645 DVDD.n14644 2.2505
R19442 DVDD.n14649 DVDD.n14648 2.2505
R19443 DVDD.n14646 DVDD.n8118 2.2505
R19444 DVDD.n14654 DVDD.n14653 2.2505
R19445 DVDD.n14657 DVDD.n14656 2.2505
R19446 DVDD.n14661 DVDD.n14660 2.2505
R19447 DVDD.n14658 DVDD.n8116 2.2505
R19448 DVDD.n14666 DVDD.n14665 2.2505
R19449 DVDD.n14669 DVDD.n14668 2.2505
R19450 DVDD.n14673 DVDD.n14672 2.2505
R19451 DVDD.n14670 DVDD.n8114 2.2505
R19452 DVDD.n14678 DVDD.n14677 2.2505
R19453 DVDD.n14681 DVDD.n14680 2.2505
R19454 DVDD.n14685 DVDD.n14684 2.2505
R19455 DVDD.n14682 DVDD.n8112 2.2505
R19456 DVDD.n14690 DVDD.n14689 2.2505
R19457 DVDD.n14693 DVDD.n14692 2.2505
R19458 DVDD.n14697 DVDD.n14696 2.2505
R19459 DVDD.n14694 DVDD.n8110 2.2505
R19460 DVDD.n14702 DVDD.n14701 2.2505
R19461 DVDD.n14705 DVDD.n14704 2.2505
R19462 DVDD.n14709 DVDD.n14708 2.2505
R19463 DVDD.n14706 DVDD.n8108 2.2505
R19464 DVDD.n14714 DVDD.n14713 2.2505
R19465 DVDD.n14717 DVDD.n14716 2.2505
R19466 DVDD.n14721 DVDD.n14720 2.2505
R19467 DVDD.n14718 DVDD.n8106 2.2505
R19468 DVDD.n14726 DVDD.n14725 2.2505
R19469 DVDD.n14729 DVDD.n14728 2.2505
R19470 DVDD.n14733 DVDD.n14732 2.2505
R19471 DVDD.n14730 DVDD.n8104 2.2505
R19472 DVDD.n14738 DVDD.n14737 2.2505
R19473 DVDD.n14741 DVDD.n14740 2.2505
R19474 DVDD.n14745 DVDD.n14744 2.2505
R19475 DVDD.n14742 DVDD.n8102 2.2505
R19476 DVDD.n14750 DVDD.n14749 2.2505
R19477 DVDD.n14753 DVDD.n14752 2.2505
R19478 DVDD.n14757 DVDD.n14756 2.2505
R19479 DVDD.n14754 DVDD.n8100 2.2505
R19480 DVDD.n14762 DVDD.n14761 2.2505
R19481 DVDD.n14765 DVDD.n14764 2.2505
R19482 DVDD.n14769 DVDD.n14768 2.2505
R19483 DVDD.n14766 DVDD.n8098 2.2505
R19484 DVDD.n14774 DVDD.n14773 2.2505
R19485 DVDD.n14777 DVDD.n14776 2.2505
R19486 DVDD.n14781 DVDD.n14780 2.2505
R19487 DVDD.n14778 DVDD.n8096 2.2505
R19488 DVDD.n14786 DVDD.n14785 2.2505
R19489 DVDD.n14789 DVDD.n14788 2.2505
R19490 DVDD.n14793 DVDD.n14792 2.2505
R19491 DVDD.n14790 DVDD.n8094 2.2505
R19492 DVDD.n14798 DVDD.n14797 2.2505
R19493 DVDD.n14801 DVDD.n14800 2.2505
R19494 DVDD.n14805 DVDD.n14804 2.2505
R19495 DVDD.n14802 DVDD.n8092 2.2505
R19496 DVDD.n14810 DVDD.n14809 2.2505
R19497 DVDD.n14813 DVDD.n14812 2.2505
R19498 DVDD.n14817 DVDD.n14816 2.2505
R19499 DVDD.n14814 DVDD.n8090 2.2505
R19500 DVDD.n14822 DVDD.n14821 2.2505
R19501 DVDD.n14824 DVDD.n8088 2.2505
R19502 DVDD.n8206 DVDD.n8158 2.2505
R19503 DVDD.n14555 DVDD.n14554 2.2505
R19504 DVDD.n14553 DVDD.n8207 2.2505
R19505 DVDD.n14552 DVDD.n14551 2.2505
R19506 DVDD.n14547 DVDD.n8208 2.2505
R19507 DVDD.n14543 DVDD.n14542 2.2505
R19508 DVDD.n14541 DVDD.n8209 2.2505
R19509 DVDD.n14540 DVDD.n14539 2.2505
R19510 DVDD.n14535 DVDD.n8210 2.2505
R19511 DVDD.n14531 DVDD.n14530 2.2505
R19512 DVDD.n14529 DVDD.n8211 2.2505
R19513 DVDD.n14528 DVDD.n14527 2.2505
R19514 DVDD.n14523 DVDD.n8212 2.2505
R19515 DVDD.n14519 DVDD.n14518 2.2505
R19516 DVDD.n14517 DVDD.n8213 2.2505
R19517 DVDD.n14516 DVDD.n14515 2.2505
R19518 DVDD.n14511 DVDD.n8214 2.2505
R19519 DVDD.n14507 DVDD.n14506 2.2505
R19520 DVDD.n14505 DVDD.n8215 2.2505
R19521 DVDD.n14504 DVDD.n14503 2.2505
R19522 DVDD.n14499 DVDD.n8216 2.2505
R19523 DVDD.n14495 DVDD.n14494 2.2505
R19524 DVDD.n14493 DVDD.n8217 2.2505
R19525 DVDD.n14492 DVDD.n14491 2.2505
R19526 DVDD.n14487 DVDD.n8218 2.2505
R19527 DVDD.n14483 DVDD.n14482 2.2505
R19528 DVDD.n14481 DVDD.n8219 2.2505
R19529 DVDD.n14480 DVDD.n14479 2.2505
R19530 DVDD.n14475 DVDD.n8220 2.2505
R19531 DVDD.n14471 DVDD.n14470 2.2505
R19532 DVDD.n14469 DVDD.n8221 2.2505
R19533 DVDD.n14468 DVDD.n14467 2.2505
R19534 DVDD.n14463 DVDD.n8222 2.2505
R19535 DVDD.n14459 DVDD.n14458 2.2505
R19536 DVDD.n14457 DVDD.n8223 2.2505
R19537 DVDD.n14456 DVDD.n14455 2.2505
R19538 DVDD.n14451 DVDD.n8224 2.2505
R19539 DVDD.n14447 DVDD.n14446 2.2505
R19540 DVDD.n14445 DVDD.n8225 2.2505
R19541 DVDD.n14444 DVDD.n14443 2.2505
R19542 DVDD.n14439 DVDD.n8226 2.2505
R19543 DVDD.n14435 DVDD.n14434 2.2505
R19544 DVDD.n14433 DVDD.n8227 2.2505
R19545 DVDD.n14432 DVDD.n14431 2.2505
R19546 DVDD.n14427 DVDD.n8228 2.2505
R19547 DVDD.n14423 DVDD.n14422 2.2505
R19548 DVDD.n14421 DVDD.n8229 2.2505
R19549 DVDD.n14420 DVDD.n14419 2.2505
R19550 DVDD.n14415 DVDD.n8230 2.2505
R19551 DVDD.n14411 DVDD.n14410 2.2505
R19552 DVDD.n14409 DVDD.n8231 2.2505
R19553 DVDD.n14408 DVDD.n14407 2.2505
R19554 DVDD.n14403 DVDD.n8232 2.2505
R19555 DVDD.n14399 DVDD.n14398 2.2505
R19556 DVDD.n14397 DVDD.n8233 2.2505
R19557 DVDD.n14396 DVDD.n14395 2.2505
R19558 DVDD.n14391 DVDD.n8234 2.2505
R19559 DVDD.n14387 DVDD.n14386 2.2505
R19560 DVDD.n14385 DVDD.n8235 2.2505
R19561 DVDD.n14384 DVDD.n14383 2.2505
R19562 DVDD.n14379 DVDD.n8236 2.2505
R19563 DVDD.n14375 DVDD.n14374 2.2505
R19564 DVDD.n14373 DVDD.n8237 2.2505
R19565 DVDD.n14372 DVDD.n14371 2.2505
R19566 DVDD.n14367 DVDD.n8238 2.2505
R19567 DVDD.n14363 DVDD.n14362 2.2505
R19568 DVDD.n14361 DVDD.n8239 2.2505
R19569 DVDD.n14360 DVDD.n14359 2.2505
R19570 DVDD.n14355 DVDD.n8240 2.2505
R19571 DVDD.n14351 DVDD.n14350 2.2505
R19572 DVDD.n14349 DVDD.n8241 2.2505
R19573 DVDD.n14348 DVDD.n14347 2.2505
R19574 DVDD.n14343 DVDD.n8242 2.2505
R19575 DVDD.n14339 DVDD.n14338 2.2505
R19576 DVDD.n14337 DVDD.n8243 2.2505
R19577 DVDD.n14336 DVDD.n14335 2.2505
R19578 DVDD.n14331 DVDD.n8244 2.2505
R19579 DVDD.n14327 DVDD.n14326 2.2505
R19580 DVDD.n14325 DVDD.n8245 2.2505
R19581 DVDD.n14324 DVDD.n14323 2.2505
R19582 DVDD.n14319 DVDD.n8246 2.2505
R19583 DVDD.n14315 DVDD.n14314 2.2505
R19584 DVDD.n14313 DVDD.n8249 2.2505
R19585 DVDD.n14312 DVDD.n14311 2.2505
R19586 DVDD.n14311 DVDD.n8204 2.2505
R19587 DVDD.n8249 DVDD.n8248 2.2505
R19588 DVDD.n14316 DVDD.n14315 2.2505
R19589 DVDD.n14319 DVDD.n14318 2.2505
R19590 DVDD.n14323 DVDD.n14322 2.2505
R19591 DVDD.n14320 DVDD.n8245 2.2505
R19592 DVDD.n14328 DVDD.n14327 2.2505
R19593 DVDD.n14331 DVDD.n14330 2.2505
R19594 DVDD.n14335 DVDD.n14334 2.2505
R19595 DVDD.n14332 DVDD.n8243 2.2505
R19596 DVDD.n14340 DVDD.n14339 2.2505
R19597 DVDD.n14343 DVDD.n14342 2.2505
R19598 DVDD.n14347 DVDD.n14346 2.2505
R19599 DVDD.n14344 DVDD.n8241 2.2505
R19600 DVDD.n14352 DVDD.n14351 2.2505
R19601 DVDD.n14355 DVDD.n14354 2.2505
R19602 DVDD.n14359 DVDD.n14358 2.2505
R19603 DVDD.n14356 DVDD.n8239 2.2505
R19604 DVDD.n14364 DVDD.n14363 2.2505
R19605 DVDD.n14367 DVDD.n14366 2.2505
R19606 DVDD.n14371 DVDD.n14370 2.2505
R19607 DVDD.n14368 DVDD.n8237 2.2505
R19608 DVDD.n14376 DVDD.n14375 2.2505
R19609 DVDD.n14379 DVDD.n14378 2.2505
R19610 DVDD.n14383 DVDD.n14382 2.2505
R19611 DVDD.n14380 DVDD.n8235 2.2505
R19612 DVDD.n14388 DVDD.n14387 2.2505
R19613 DVDD.n14391 DVDD.n14390 2.2505
R19614 DVDD.n14395 DVDD.n14394 2.2505
R19615 DVDD.n14392 DVDD.n8233 2.2505
R19616 DVDD.n14400 DVDD.n14399 2.2505
R19617 DVDD.n14403 DVDD.n14402 2.2505
R19618 DVDD.n14407 DVDD.n14406 2.2505
R19619 DVDD.n14404 DVDD.n8231 2.2505
R19620 DVDD.n14412 DVDD.n14411 2.2505
R19621 DVDD.n14415 DVDD.n14414 2.2505
R19622 DVDD.n14419 DVDD.n14418 2.2505
R19623 DVDD.n14416 DVDD.n8229 2.2505
R19624 DVDD.n14424 DVDD.n14423 2.2505
R19625 DVDD.n14427 DVDD.n14426 2.2505
R19626 DVDD.n14431 DVDD.n14430 2.2505
R19627 DVDD.n14428 DVDD.n8227 2.2505
R19628 DVDD.n14436 DVDD.n14435 2.2505
R19629 DVDD.n14439 DVDD.n14438 2.2505
R19630 DVDD.n14443 DVDD.n14442 2.2505
R19631 DVDD.n14440 DVDD.n8225 2.2505
R19632 DVDD.n14448 DVDD.n14447 2.2505
R19633 DVDD.n14451 DVDD.n14450 2.2505
R19634 DVDD.n14455 DVDD.n14454 2.2505
R19635 DVDD.n14452 DVDD.n8223 2.2505
R19636 DVDD.n14460 DVDD.n14459 2.2505
R19637 DVDD.n14463 DVDD.n14462 2.2505
R19638 DVDD.n14467 DVDD.n14466 2.2505
R19639 DVDD.n14464 DVDD.n8221 2.2505
R19640 DVDD.n14472 DVDD.n14471 2.2505
R19641 DVDD.n14475 DVDD.n14474 2.2505
R19642 DVDD.n14479 DVDD.n14478 2.2505
R19643 DVDD.n14476 DVDD.n8219 2.2505
R19644 DVDD.n14484 DVDD.n14483 2.2505
R19645 DVDD.n14487 DVDD.n14486 2.2505
R19646 DVDD.n14491 DVDD.n14490 2.2505
R19647 DVDD.n14488 DVDD.n8217 2.2505
R19648 DVDD.n14496 DVDD.n14495 2.2505
R19649 DVDD.n14499 DVDD.n14498 2.2505
R19650 DVDD.n14503 DVDD.n14502 2.2505
R19651 DVDD.n14500 DVDD.n8215 2.2505
R19652 DVDD.n14508 DVDD.n14507 2.2505
R19653 DVDD.n14511 DVDD.n14510 2.2505
R19654 DVDD.n14515 DVDD.n14514 2.2505
R19655 DVDD.n14512 DVDD.n8213 2.2505
R19656 DVDD.n14520 DVDD.n14519 2.2505
R19657 DVDD.n14523 DVDD.n14522 2.2505
R19658 DVDD.n14527 DVDD.n14526 2.2505
R19659 DVDD.n14524 DVDD.n8211 2.2505
R19660 DVDD.n14532 DVDD.n14531 2.2505
R19661 DVDD.n14535 DVDD.n14534 2.2505
R19662 DVDD.n14539 DVDD.n14538 2.2505
R19663 DVDD.n14536 DVDD.n8209 2.2505
R19664 DVDD.n14544 DVDD.n14543 2.2505
R19665 DVDD.n14547 DVDD.n14546 2.2505
R19666 DVDD.n14551 DVDD.n14550 2.2505
R19667 DVDD.n14548 DVDD.n8207 2.2505
R19668 DVDD.n14556 DVDD.n14555 2.2505
R19669 DVDD.n14558 DVDD.n8206 2.2505
R19670 DVDD.n8598 DVDD.n8597 2.2505
R19671 DVDD.n8265 DVDD.n8264 2.2505
R19672 DVDD.n8587 DVDD.n8266 2.2505
R19673 DVDD.n8589 DVDD.n8588 2.2505
R19674 DVDD.n8586 DVDD.n8268 2.2505
R19675 DVDD.n8585 DVDD.n8584 2.2505
R19676 DVDD.n8270 DVDD.n8269 2.2505
R19677 DVDD.n8576 DVDD.n8575 2.2505
R19678 DVDD.n8574 DVDD.n8272 2.2505
R19679 DVDD.n8573 DVDD.n8572 2.2505
R19680 DVDD.n8274 DVDD.n8273 2.2505
R19681 DVDD.n8564 DVDD.n8563 2.2505
R19682 DVDD.n8562 DVDD.n8276 2.2505
R19683 DVDD.n8561 DVDD.n8560 2.2505
R19684 DVDD.n8278 DVDD.n8277 2.2505
R19685 DVDD.n8552 DVDD.n8551 2.2505
R19686 DVDD.n8550 DVDD.n8280 2.2505
R19687 DVDD.n8549 DVDD.n8548 2.2505
R19688 DVDD.n8282 DVDD.n8281 2.2505
R19689 DVDD.n8540 DVDD.n8539 2.2505
R19690 DVDD.n8538 DVDD.n8284 2.2505
R19691 DVDD.n8537 DVDD.n8536 2.2505
R19692 DVDD.n8286 DVDD.n8285 2.2505
R19693 DVDD.n8528 DVDD.n8527 2.2505
R19694 DVDD.n8526 DVDD.n8288 2.2505
R19695 DVDD.n8525 DVDD.n8524 2.2505
R19696 DVDD.n8290 DVDD.n8289 2.2505
R19697 DVDD.n8516 DVDD.n8515 2.2505
R19698 DVDD.n8514 DVDD.n8292 2.2505
R19699 DVDD.n8513 DVDD.n8512 2.2505
R19700 DVDD.n8294 DVDD.n8293 2.2505
R19701 DVDD.n8504 DVDD.n8503 2.2505
R19702 DVDD.n8502 DVDD.n8296 2.2505
R19703 DVDD.n8501 DVDD.n8500 2.2505
R19704 DVDD.n8298 DVDD.n8297 2.2505
R19705 DVDD.n8492 DVDD.n8491 2.2505
R19706 DVDD.n8490 DVDD.n8300 2.2505
R19707 DVDD.n8489 DVDD.n8488 2.2505
R19708 DVDD.n8302 DVDD.n8301 2.2505
R19709 DVDD.n8480 DVDD.n8479 2.2505
R19710 DVDD.n8478 DVDD.n8304 2.2505
R19711 DVDD.n8477 DVDD.n8476 2.2505
R19712 DVDD.n8306 DVDD.n8305 2.2505
R19713 DVDD.n8468 DVDD.n8467 2.2505
R19714 DVDD.n8466 DVDD.n8308 2.2505
R19715 DVDD.n8465 DVDD.n8464 2.2505
R19716 DVDD.n8310 DVDD.n8309 2.2505
R19717 DVDD.n8456 DVDD.n8455 2.2505
R19718 DVDD.n8454 DVDD.n8312 2.2505
R19719 DVDD.n8453 DVDD.n8452 2.2505
R19720 DVDD.n8314 DVDD.n8313 2.2505
R19721 DVDD.n8444 DVDD.n8443 2.2505
R19722 DVDD.n8442 DVDD.n8316 2.2505
R19723 DVDD.n8441 DVDD.n8440 2.2505
R19724 DVDD.n8318 DVDD.n8317 2.2505
R19725 DVDD.n8432 DVDD.n8431 2.2505
R19726 DVDD.n8430 DVDD.n8320 2.2505
R19727 DVDD.n8429 DVDD.n8428 2.2505
R19728 DVDD.n8322 DVDD.n8321 2.2505
R19729 DVDD.n8420 DVDD.n8419 2.2505
R19730 DVDD.n8418 DVDD.n8324 2.2505
R19731 DVDD.n8417 DVDD.n8416 2.2505
R19732 DVDD.n8326 DVDD.n8325 2.2505
R19733 DVDD.n8408 DVDD.n8407 2.2505
R19734 DVDD.n8406 DVDD.n8328 2.2505
R19735 DVDD.n8405 DVDD.n8404 2.2505
R19736 DVDD.n8330 DVDD.n8329 2.2505
R19737 DVDD.n8396 DVDD.n8395 2.2505
R19738 DVDD.n8394 DVDD.n8332 2.2505
R19739 DVDD.n8393 DVDD.n8392 2.2505
R19740 DVDD.n8334 DVDD.n8333 2.2505
R19741 DVDD.n8384 DVDD.n8383 2.2505
R19742 DVDD.n8382 DVDD.n8336 2.2505
R19743 DVDD.n8381 DVDD.n8380 2.2505
R19744 DVDD.n8338 DVDD.n8337 2.2505
R19745 DVDD.n8372 DVDD.n8371 2.2505
R19746 DVDD.n8370 DVDD.n8340 2.2505
R19747 DVDD.n8369 DVDD.n8368 2.2505
R19748 DVDD.n8342 DVDD.n8341 2.2505
R19749 DVDD.n8360 DVDD.n8359 2.2505
R19750 DVDD.n8358 DVDD.n8344 2.2505
R19751 DVDD.n8357 DVDD.n8356 2.2505
R19752 DVDD.n8346 DVDD.n8345 2.2505
R19753 DVDD.n8348 DVDD.n8347 2.2505
R19754 DVDD.n8349 DVDD.n8348 2.2505
R19755 DVDD.n8351 DVDD.n8346 2.2505
R19756 DVDD.n8356 DVDD.n8355 2.2505
R19757 DVDD.n8353 DVDD.n8344 2.2505
R19758 DVDD.n8361 DVDD.n8360 2.2505
R19759 DVDD.n8363 DVDD.n8342 2.2505
R19760 DVDD.n8368 DVDD.n8367 2.2505
R19761 DVDD.n8365 DVDD.n8340 2.2505
R19762 DVDD.n8373 DVDD.n8372 2.2505
R19763 DVDD.n8375 DVDD.n8338 2.2505
R19764 DVDD.n8380 DVDD.n8379 2.2505
R19765 DVDD.n8377 DVDD.n8336 2.2505
R19766 DVDD.n8385 DVDD.n8384 2.2505
R19767 DVDD.n8387 DVDD.n8334 2.2505
R19768 DVDD.n8392 DVDD.n8391 2.2505
R19769 DVDD.n8389 DVDD.n8332 2.2505
R19770 DVDD.n8397 DVDD.n8396 2.2505
R19771 DVDD.n8399 DVDD.n8330 2.2505
R19772 DVDD.n8404 DVDD.n8403 2.2505
R19773 DVDD.n8401 DVDD.n8328 2.2505
R19774 DVDD.n8409 DVDD.n8408 2.2505
R19775 DVDD.n8411 DVDD.n8326 2.2505
R19776 DVDD.n8416 DVDD.n8415 2.2505
R19777 DVDD.n8413 DVDD.n8324 2.2505
R19778 DVDD.n8421 DVDD.n8420 2.2505
R19779 DVDD.n8423 DVDD.n8322 2.2505
R19780 DVDD.n8428 DVDD.n8427 2.2505
R19781 DVDD.n8425 DVDD.n8320 2.2505
R19782 DVDD.n8433 DVDD.n8432 2.2505
R19783 DVDD.n8435 DVDD.n8318 2.2505
R19784 DVDD.n8440 DVDD.n8439 2.2505
R19785 DVDD.n8437 DVDD.n8316 2.2505
R19786 DVDD.n8445 DVDD.n8444 2.2505
R19787 DVDD.n8447 DVDD.n8314 2.2505
R19788 DVDD.n8452 DVDD.n8451 2.2505
R19789 DVDD.n8449 DVDD.n8312 2.2505
R19790 DVDD.n8457 DVDD.n8456 2.2505
R19791 DVDD.n8459 DVDD.n8310 2.2505
R19792 DVDD.n8464 DVDD.n8463 2.2505
R19793 DVDD.n8461 DVDD.n8308 2.2505
R19794 DVDD.n8469 DVDD.n8468 2.2505
R19795 DVDD.n8471 DVDD.n8306 2.2505
R19796 DVDD.n8476 DVDD.n8475 2.2505
R19797 DVDD.n8473 DVDD.n8304 2.2505
R19798 DVDD.n8481 DVDD.n8480 2.2505
R19799 DVDD.n8483 DVDD.n8302 2.2505
R19800 DVDD.n8488 DVDD.n8487 2.2505
R19801 DVDD.n8485 DVDD.n8300 2.2505
R19802 DVDD.n8493 DVDD.n8492 2.2505
R19803 DVDD.n8495 DVDD.n8298 2.2505
R19804 DVDD.n8500 DVDD.n8499 2.2505
R19805 DVDD.n8497 DVDD.n8296 2.2505
R19806 DVDD.n8505 DVDD.n8504 2.2505
R19807 DVDD.n8507 DVDD.n8294 2.2505
R19808 DVDD.n8512 DVDD.n8511 2.2505
R19809 DVDD.n8509 DVDD.n8292 2.2505
R19810 DVDD.n8517 DVDD.n8516 2.2505
R19811 DVDD.n8519 DVDD.n8290 2.2505
R19812 DVDD.n8524 DVDD.n8523 2.2505
R19813 DVDD.n8521 DVDD.n8288 2.2505
R19814 DVDD.n8529 DVDD.n8528 2.2505
R19815 DVDD.n8531 DVDD.n8286 2.2505
R19816 DVDD.n8536 DVDD.n8535 2.2505
R19817 DVDD.n8533 DVDD.n8284 2.2505
R19818 DVDD.n8541 DVDD.n8540 2.2505
R19819 DVDD.n8543 DVDD.n8282 2.2505
R19820 DVDD.n8548 DVDD.n8547 2.2505
R19821 DVDD.n8545 DVDD.n8280 2.2505
R19822 DVDD.n8553 DVDD.n8552 2.2505
R19823 DVDD.n8555 DVDD.n8278 2.2505
R19824 DVDD.n8560 DVDD.n8559 2.2505
R19825 DVDD.n8557 DVDD.n8276 2.2505
R19826 DVDD.n8565 DVDD.n8564 2.2505
R19827 DVDD.n8567 DVDD.n8274 2.2505
R19828 DVDD.n8572 DVDD.n8571 2.2505
R19829 DVDD.n8569 DVDD.n8272 2.2505
R19830 DVDD.n8577 DVDD.n8576 2.2505
R19831 DVDD.n8579 DVDD.n8270 2.2505
R19832 DVDD.n8584 DVDD.n8583 2.2505
R19833 DVDD.n8581 DVDD.n8268 2.2505
R19834 DVDD.n8590 DVDD.n8589 2.2505
R19835 DVDD.n8592 DVDD.n8266 2.2505
R19836 DVDD.n8594 DVDD.n8265 2.2505
R19837 DVDD.n8597 DVDD.n8596 2.2505
R19838 DVDD.n8740 DVDD.n8739 2.2505
R19839 DVDD.n8742 DVDD.n8741 2.2505
R19840 DVDD.n8734 DVDD.n8733 2.2505
R19841 DVDD.n8749 DVDD.n8748 2.2505
R19842 DVDD.n8750 DVDD.n8732 2.2505
R19843 DVDD.n8752 DVDD.n8751 2.2505
R19844 DVDD.n8728 DVDD.n8727 2.2505
R19845 DVDD.n8759 DVDD.n8758 2.2505
R19846 DVDD.n8760 DVDD.n8726 2.2505
R19847 DVDD.n8762 DVDD.n8761 2.2505
R19848 DVDD.n8722 DVDD.n8721 2.2505
R19849 DVDD.n8769 DVDD.n8768 2.2505
R19850 DVDD.n8770 DVDD.n8720 2.2505
R19851 DVDD.n8772 DVDD.n8771 2.2505
R19852 DVDD.n8716 DVDD.n8715 2.2505
R19853 DVDD.n8779 DVDD.n8778 2.2505
R19854 DVDD.n8780 DVDD.n8714 2.2505
R19855 DVDD.n8782 DVDD.n8781 2.2505
R19856 DVDD.n8710 DVDD.n8709 2.2505
R19857 DVDD.n8789 DVDD.n8788 2.2505
R19858 DVDD.n8790 DVDD.n8708 2.2505
R19859 DVDD.n8792 DVDD.n8791 2.2505
R19860 DVDD.n8704 DVDD.n8703 2.2505
R19861 DVDD.n8799 DVDD.n8798 2.2505
R19862 DVDD.n8800 DVDD.n8702 2.2505
R19863 DVDD.n8802 DVDD.n8801 2.2505
R19864 DVDD.n8698 DVDD.n8697 2.2505
R19865 DVDD.n8809 DVDD.n8808 2.2505
R19866 DVDD.n8810 DVDD.n8696 2.2505
R19867 DVDD.n8812 DVDD.n8811 2.2505
R19868 DVDD.n8692 DVDD.n8691 2.2505
R19869 DVDD.n8819 DVDD.n8818 2.2505
R19870 DVDD.n8820 DVDD.n8690 2.2505
R19871 DVDD.n8822 DVDD.n8821 2.2505
R19872 DVDD.n8686 DVDD.n8685 2.2505
R19873 DVDD.n8829 DVDD.n8828 2.2505
R19874 DVDD.n8830 DVDD.n8684 2.2505
R19875 DVDD.n8832 DVDD.n8831 2.2505
R19876 DVDD.n8680 DVDD.n8679 2.2505
R19877 DVDD.n8839 DVDD.n8838 2.2505
R19878 DVDD.n8840 DVDD.n8678 2.2505
R19879 DVDD.n8842 DVDD.n8841 2.2505
R19880 DVDD.n8674 DVDD.n8673 2.2505
R19881 DVDD.n8849 DVDD.n8848 2.2505
R19882 DVDD.n8850 DVDD.n8672 2.2505
R19883 DVDD.n8852 DVDD.n8851 2.2505
R19884 DVDD.n8668 DVDD.n8667 2.2505
R19885 DVDD.n8859 DVDD.n8858 2.2505
R19886 DVDD.n8860 DVDD.n8666 2.2505
R19887 DVDD.n8862 DVDD.n8861 2.2505
R19888 DVDD.n8662 DVDD.n8661 2.2505
R19889 DVDD.n8869 DVDD.n8868 2.2505
R19890 DVDD.n8870 DVDD.n8660 2.2505
R19891 DVDD.n8872 DVDD.n8871 2.2505
R19892 DVDD.n8656 DVDD.n8655 2.2505
R19893 DVDD.n8879 DVDD.n8878 2.2505
R19894 DVDD.n8880 DVDD.n8654 2.2505
R19895 DVDD.n8882 DVDD.n8881 2.2505
R19896 DVDD.n8650 DVDD.n8649 2.2505
R19897 DVDD.n8889 DVDD.n8888 2.2505
R19898 DVDD.n8890 DVDD.n8648 2.2505
R19899 DVDD.n8892 DVDD.n8891 2.2505
R19900 DVDD.n8644 DVDD.n8643 2.2505
R19901 DVDD.n8899 DVDD.n8898 2.2505
R19902 DVDD.n8900 DVDD.n8642 2.2505
R19903 DVDD.n8902 DVDD.n8901 2.2505
R19904 DVDD.n8638 DVDD.n8637 2.2505
R19905 DVDD.n8909 DVDD.n8908 2.2505
R19906 DVDD.n8910 DVDD.n8636 2.2505
R19907 DVDD.n8912 DVDD.n8911 2.2505
R19908 DVDD.n8632 DVDD.n8631 2.2505
R19909 DVDD.n8919 DVDD.n8918 2.2505
R19910 DVDD.n8920 DVDD.n8630 2.2505
R19911 DVDD.n8922 DVDD.n8921 2.2505
R19912 DVDD.n8626 DVDD.n8625 2.2505
R19913 DVDD.n8929 DVDD.n8928 2.2505
R19914 DVDD.n8930 DVDD.n8624 2.2505
R19915 DVDD.n8932 DVDD.n8931 2.2505
R19916 DVDD.n8620 DVDD.n8619 2.2505
R19917 DVDD.n8939 DVDD.n8938 2.2505
R19918 DVDD.n8940 DVDD.n8618 2.2505
R19919 DVDD.n8942 DVDD.n8941 2.2505
R19920 DVDD.n8616 DVDD.n8615 2.2505
R19921 DVDD.n8949 DVDD.n8948 2.2505
R19922 DVDD.n8948 DVDD.n8947 2.2505
R19923 DVDD.n8945 DVDD.n8616 2.2505
R19924 DVDD.n8943 DVDD.n8942 2.2505
R19925 DVDD.n8621 DVDD.n8618 2.2505
R19926 DVDD.n8938 DVDD.n8937 2.2505
R19927 DVDD.n8935 DVDD.n8620 2.2505
R19928 DVDD.n8933 DVDD.n8932 2.2505
R19929 DVDD.n8627 DVDD.n8624 2.2505
R19930 DVDD.n8928 DVDD.n8927 2.2505
R19931 DVDD.n8925 DVDD.n8626 2.2505
R19932 DVDD.n8923 DVDD.n8922 2.2505
R19933 DVDD.n8633 DVDD.n8630 2.2505
R19934 DVDD.n8918 DVDD.n8917 2.2505
R19935 DVDD.n8915 DVDD.n8632 2.2505
R19936 DVDD.n8913 DVDD.n8912 2.2505
R19937 DVDD.n8639 DVDD.n8636 2.2505
R19938 DVDD.n8908 DVDD.n8907 2.2505
R19939 DVDD.n8905 DVDD.n8638 2.2505
R19940 DVDD.n8903 DVDD.n8902 2.2505
R19941 DVDD.n8645 DVDD.n8642 2.2505
R19942 DVDD.n8898 DVDD.n8897 2.2505
R19943 DVDD.n8895 DVDD.n8644 2.2505
R19944 DVDD.n8893 DVDD.n8892 2.2505
R19945 DVDD.n8651 DVDD.n8648 2.2505
R19946 DVDD.n8888 DVDD.n8887 2.2505
R19947 DVDD.n8885 DVDD.n8650 2.2505
R19948 DVDD.n8883 DVDD.n8882 2.2505
R19949 DVDD.n8657 DVDD.n8654 2.2505
R19950 DVDD.n8878 DVDD.n8877 2.2505
R19951 DVDD.n8875 DVDD.n8656 2.2505
R19952 DVDD.n8873 DVDD.n8872 2.2505
R19953 DVDD.n8663 DVDD.n8660 2.2505
R19954 DVDD.n8868 DVDD.n8867 2.2505
R19955 DVDD.n8865 DVDD.n8662 2.2505
R19956 DVDD.n8863 DVDD.n8862 2.2505
R19957 DVDD.n8669 DVDD.n8666 2.2505
R19958 DVDD.n8858 DVDD.n8857 2.2505
R19959 DVDD.n8855 DVDD.n8668 2.2505
R19960 DVDD.n8853 DVDD.n8852 2.2505
R19961 DVDD.n8675 DVDD.n8672 2.2505
R19962 DVDD.n8848 DVDD.n8847 2.2505
R19963 DVDD.n8845 DVDD.n8674 2.2505
R19964 DVDD.n8843 DVDD.n8842 2.2505
R19965 DVDD.n8681 DVDD.n8678 2.2505
R19966 DVDD.n8838 DVDD.n8837 2.2505
R19967 DVDD.n8835 DVDD.n8680 2.2505
R19968 DVDD.n8833 DVDD.n8832 2.2505
R19969 DVDD.n8687 DVDD.n8684 2.2505
R19970 DVDD.n8828 DVDD.n8827 2.2505
R19971 DVDD.n8825 DVDD.n8686 2.2505
R19972 DVDD.n8823 DVDD.n8822 2.2505
R19973 DVDD.n8693 DVDD.n8690 2.2505
R19974 DVDD.n8818 DVDD.n8817 2.2505
R19975 DVDD.n8815 DVDD.n8692 2.2505
R19976 DVDD.n8813 DVDD.n8812 2.2505
R19977 DVDD.n8699 DVDD.n8696 2.2505
R19978 DVDD.n8808 DVDD.n8807 2.2505
R19979 DVDD.n8805 DVDD.n8698 2.2505
R19980 DVDD.n8803 DVDD.n8802 2.2505
R19981 DVDD.n8705 DVDD.n8702 2.2505
R19982 DVDD.n8798 DVDD.n8797 2.2505
R19983 DVDD.n8795 DVDD.n8704 2.2505
R19984 DVDD.n8793 DVDD.n8792 2.2505
R19985 DVDD.n8711 DVDD.n8708 2.2505
R19986 DVDD.n8788 DVDD.n8787 2.2505
R19987 DVDD.n8785 DVDD.n8710 2.2505
R19988 DVDD.n8783 DVDD.n8782 2.2505
R19989 DVDD.n8717 DVDD.n8714 2.2505
R19990 DVDD.n8778 DVDD.n8777 2.2505
R19991 DVDD.n8775 DVDD.n8716 2.2505
R19992 DVDD.n8773 DVDD.n8772 2.2505
R19993 DVDD.n8723 DVDD.n8720 2.2505
R19994 DVDD.n8768 DVDD.n8767 2.2505
R19995 DVDD.n8765 DVDD.n8722 2.2505
R19996 DVDD.n8763 DVDD.n8762 2.2505
R19997 DVDD.n8729 DVDD.n8726 2.2505
R19998 DVDD.n8758 DVDD.n8757 2.2505
R19999 DVDD.n8755 DVDD.n8728 2.2505
R20000 DVDD.n8753 DVDD.n8752 2.2505
R20001 DVDD.n8735 DVDD.n8732 2.2505
R20002 DVDD.n8748 DVDD.n8747 2.2505
R20003 DVDD.n8745 DVDD.n8734 2.2505
R20004 DVDD.n8743 DVDD.n8742 2.2505
R20005 DVDD.n8739 DVDD.n8738 2.2505
R20006 DVDD.n14279 DVDD.n10576 2.2505
R20007 DVDD.n10575 DVDD.n10331 2.2505
R20008 DVDD.n10574 DVDD.n10573 2.2505
R20009 DVDD.n10571 DVDD.n10332 2.2505
R20010 DVDD.n10569 DVDD.n10567 2.2505
R20011 DVDD.n10566 DVDD.n10334 2.2505
R20012 DVDD.n10565 DVDD.n10564 2.2505
R20013 DVDD.n10562 DVDD.n10335 2.2505
R20014 DVDD.n10560 DVDD.n10558 2.2505
R20015 DVDD.n10557 DVDD.n10337 2.2505
R20016 DVDD.n10556 DVDD.n10555 2.2505
R20017 DVDD.n10553 DVDD.n10338 2.2505
R20018 DVDD.n10551 DVDD.n10549 2.2505
R20019 DVDD.n10548 DVDD.n10340 2.2505
R20020 DVDD.n10547 DVDD.n10546 2.2505
R20021 DVDD.n10544 DVDD.n10341 2.2505
R20022 DVDD.n10542 DVDD.n10540 2.2505
R20023 DVDD.n10539 DVDD.n10343 2.2505
R20024 DVDD.n10538 DVDD.n10537 2.2505
R20025 DVDD.n10535 DVDD.n10344 2.2505
R20026 DVDD.n10533 DVDD.n10531 2.2505
R20027 DVDD.n10530 DVDD.n10346 2.2505
R20028 DVDD.n10529 DVDD.n10528 2.2505
R20029 DVDD.n10526 DVDD.n10347 2.2505
R20030 DVDD.n10524 DVDD.n10522 2.2505
R20031 DVDD.n10521 DVDD.n10349 2.2505
R20032 DVDD.n10520 DVDD.n10519 2.2505
R20033 DVDD.n10517 DVDD.n10350 2.2505
R20034 DVDD.n10515 DVDD.n10513 2.2505
R20035 DVDD.n10512 DVDD.n10352 2.2505
R20036 DVDD.n10511 DVDD.n10510 2.2505
R20037 DVDD.n10508 DVDD.n10353 2.2505
R20038 DVDD.n10506 DVDD.n10504 2.2505
R20039 DVDD.n10503 DVDD.n10355 2.2505
R20040 DVDD.n10502 DVDD.n10501 2.2505
R20041 DVDD.n10499 DVDD.n10356 2.2505
R20042 DVDD.n10497 DVDD.n10495 2.2505
R20043 DVDD.n10494 DVDD.n10358 2.2505
R20044 DVDD.n10493 DVDD.n10492 2.2505
R20045 DVDD.n10490 DVDD.n10359 2.2505
R20046 DVDD.n10488 DVDD.n10486 2.2505
R20047 DVDD.n10485 DVDD.n10361 2.2505
R20048 DVDD.n10484 DVDD.n10483 2.2505
R20049 DVDD.n10481 DVDD.n10362 2.2505
R20050 DVDD.n10479 DVDD.n10477 2.2505
R20051 DVDD.n10476 DVDD.n10364 2.2505
R20052 DVDD.n10475 DVDD.n10474 2.2505
R20053 DVDD.n10472 DVDD.n10365 2.2505
R20054 DVDD.n10470 DVDD.n10468 2.2505
R20055 DVDD.n10467 DVDD.n10367 2.2505
R20056 DVDD.n10466 DVDD.n10465 2.2505
R20057 DVDD.n10463 DVDD.n10368 2.2505
R20058 DVDD.n10461 DVDD.n10459 2.2505
R20059 DVDD.n10458 DVDD.n10370 2.2505
R20060 DVDD.n10457 DVDD.n10456 2.2505
R20061 DVDD.n10454 DVDD.n10371 2.2505
R20062 DVDD.n10452 DVDD.n10450 2.2505
R20063 DVDD.n10449 DVDD.n10373 2.2505
R20064 DVDD.n10448 DVDD.n10447 2.2505
R20065 DVDD.n10445 DVDD.n10374 2.2505
R20066 DVDD.n10443 DVDD.n10441 2.2505
R20067 DVDD.n10440 DVDD.n10376 2.2505
R20068 DVDD.n10439 DVDD.n10438 2.2505
R20069 DVDD.n10436 DVDD.n10377 2.2505
R20070 DVDD.n10434 DVDD.n10432 2.2505
R20071 DVDD.n10431 DVDD.n10379 2.2505
R20072 DVDD.n10430 DVDD.n10429 2.2505
R20073 DVDD.n10427 DVDD.n10380 2.2505
R20074 DVDD.n10425 DVDD.n10423 2.2505
R20075 DVDD.n10422 DVDD.n10382 2.2505
R20076 DVDD.n10421 DVDD.n10420 2.2505
R20077 DVDD.n10418 DVDD.n10383 2.2505
R20078 DVDD.n10416 DVDD.n10414 2.2505
R20079 DVDD.n10413 DVDD.n10385 2.2505
R20080 DVDD.n10412 DVDD.n10411 2.2505
R20081 DVDD.n10409 DVDD.n10386 2.2505
R20082 DVDD.n10407 DVDD.n10405 2.2505
R20083 DVDD.n10404 DVDD.n10388 2.2505
R20084 DVDD.n10403 DVDD.n10402 2.2505
R20085 DVDD.n10400 DVDD.n10389 2.2505
R20086 DVDD.n10398 DVDD.n10396 2.2505
R20087 DVDD.n10395 DVDD.n10391 2.2505
R20088 DVDD.n10394 DVDD.n10393 2.2505
R20089 DVDD.n10392 DVDD.n10285 2.2505
R20090 DVDD.n14282 DVDD.n10285 2.2505
R20091 DVDD.n10393 DVDD.n10284 2.2505
R20092 DVDD.n10391 DVDD.n10390 2.2505
R20093 DVDD.n10398 DVDD.n10397 2.2505
R20094 DVDD.n10400 DVDD.n10399 2.2505
R20095 DVDD.n10402 DVDD.n10401 2.2505
R20096 DVDD.n10388 DVDD.n10387 2.2505
R20097 DVDD.n10407 DVDD.n10406 2.2505
R20098 DVDD.n10409 DVDD.n10408 2.2505
R20099 DVDD.n10411 DVDD.n10410 2.2505
R20100 DVDD.n10385 DVDD.n10384 2.2505
R20101 DVDD.n10416 DVDD.n10415 2.2505
R20102 DVDD.n10418 DVDD.n10417 2.2505
R20103 DVDD.n10420 DVDD.n10419 2.2505
R20104 DVDD.n10382 DVDD.n10381 2.2505
R20105 DVDD.n10425 DVDD.n10424 2.2505
R20106 DVDD.n10427 DVDD.n10426 2.2505
R20107 DVDD.n10429 DVDD.n10428 2.2505
R20108 DVDD.n10379 DVDD.n10378 2.2505
R20109 DVDD.n10434 DVDD.n10433 2.2505
R20110 DVDD.n10436 DVDD.n10435 2.2505
R20111 DVDD.n10438 DVDD.n10437 2.2505
R20112 DVDD.n10376 DVDD.n10375 2.2505
R20113 DVDD.n10443 DVDD.n10442 2.2505
R20114 DVDD.n10445 DVDD.n10444 2.2505
R20115 DVDD.n10447 DVDD.n10446 2.2505
R20116 DVDD.n10373 DVDD.n10372 2.2505
R20117 DVDD.n10452 DVDD.n10451 2.2505
R20118 DVDD.n10454 DVDD.n10453 2.2505
R20119 DVDD.n10456 DVDD.n10455 2.2505
R20120 DVDD.n10370 DVDD.n10369 2.2505
R20121 DVDD.n10461 DVDD.n10460 2.2505
R20122 DVDD.n10463 DVDD.n10462 2.2505
R20123 DVDD.n10465 DVDD.n10464 2.2505
R20124 DVDD.n10367 DVDD.n10366 2.2505
R20125 DVDD.n10470 DVDD.n10469 2.2505
R20126 DVDD.n10472 DVDD.n10471 2.2505
R20127 DVDD.n10474 DVDD.n10473 2.2505
R20128 DVDD.n10364 DVDD.n10363 2.2505
R20129 DVDD.n10479 DVDD.n10478 2.2505
R20130 DVDD.n10481 DVDD.n10480 2.2505
R20131 DVDD.n10483 DVDD.n10482 2.2505
R20132 DVDD.n10361 DVDD.n10360 2.2505
R20133 DVDD.n10488 DVDD.n10487 2.2505
R20134 DVDD.n10490 DVDD.n10489 2.2505
R20135 DVDD.n10492 DVDD.n10491 2.2505
R20136 DVDD.n10358 DVDD.n10357 2.2505
R20137 DVDD.n10497 DVDD.n10496 2.2505
R20138 DVDD.n10499 DVDD.n10498 2.2505
R20139 DVDD.n10501 DVDD.n10500 2.2505
R20140 DVDD.n10355 DVDD.n10354 2.2505
R20141 DVDD.n10506 DVDD.n10505 2.2505
R20142 DVDD.n10508 DVDD.n10507 2.2505
R20143 DVDD.n10510 DVDD.n10509 2.2505
R20144 DVDD.n10352 DVDD.n10351 2.2505
R20145 DVDD.n10515 DVDD.n10514 2.2505
R20146 DVDD.n10517 DVDD.n10516 2.2505
R20147 DVDD.n10519 DVDD.n10518 2.2505
R20148 DVDD.n10349 DVDD.n10348 2.2505
R20149 DVDD.n10524 DVDD.n10523 2.2505
R20150 DVDD.n10526 DVDD.n10525 2.2505
R20151 DVDD.n10528 DVDD.n10527 2.2505
R20152 DVDD.n10346 DVDD.n10345 2.2505
R20153 DVDD.n10533 DVDD.n10532 2.2505
R20154 DVDD.n10535 DVDD.n10534 2.2505
R20155 DVDD.n10537 DVDD.n10536 2.2505
R20156 DVDD.n10343 DVDD.n10342 2.2505
R20157 DVDD.n10542 DVDD.n10541 2.2505
R20158 DVDD.n10544 DVDD.n10543 2.2505
R20159 DVDD.n10546 DVDD.n10545 2.2505
R20160 DVDD.n10340 DVDD.n10339 2.2505
R20161 DVDD.n10551 DVDD.n10550 2.2505
R20162 DVDD.n10553 DVDD.n10552 2.2505
R20163 DVDD.n10555 DVDD.n10554 2.2505
R20164 DVDD.n10337 DVDD.n10336 2.2505
R20165 DVDD.n10560 DVDD.n10559 2.2505
R20166 DVDD.n10562 DVDD.n10561 2.2505
R20167 DVDD.n10564 DVDD.n10563 2.2505
R20168 DVDD.n10334 DVDD.n10333 2.2505
R20169 DVDD.n10569 DVDD.n10568 2.2505
R20170 DVDD.n10571 DVDD.n10570 2.2505
R20171 DVDD.n10573 DVDD.n10572 2.2505
R20172 DVDD.n10331 DVDD.n10330 2.2505
R20173 DVDD.n14280 DVDD.n14279 2.2505
R20174 DVDD.n10641 DVDD.n10591 2.2505
R20175 DVDD.n14265 DVDD.n14264 2.2505
R20176 DVDD.n14263 DVDD.n10643 2.2505
R20177 DVDD.n14262 DVDD.n14261 2.2505
R20178 DVDD.n14257 DVDD.n10644 2.2505
R20179 DVDD.n14253 DVDD.n14252 2.2505
R20180 DVDD.n14251 DVDD.n10645 2.2505
R20181 DVDD.n14250 DVDD.n14249 2.2505
R20182 DVDD.n14245 DVDD.n10646 2.2505
R20183 DVDD.n14241 DVDD.n14240 2.2505
R20184 DVDD.n14239 DVDD.n10647 2.2505
R20185 DVDD.n14238 DVDD.n14237 2.2505
R20186 DVDD.n14233 DVDD.n10648 2.2505
R20187 DVDD.n14229 DVDD.n14228 2.2505
R20188 DVDD.n14227 DVDD.n10649 2.2505
R20189 DVDD.n14226 DVDD.n14225 2.2505
R20190 DVDD.n14221 DVDD.n10650 2.2505
R20191 DVDD.n14217 DVDD.n14216 2.2505
R20192 DVDD.n14215 DVDD.n10651 2.2505
R20193 DVDD.n14214 DVDD.n14213 2.2505
R20194 DVDD.n14209 DVDD.n10652 2.2505
R20195 DVDD.n14205 DVDD.n14204 2.2505
R20196 DVDD.n14203 DVDD.n10653 2.2505
R20197 DVDD.n14202 DVDD.n14201 2.2505
R20198 DVDD.n14197 DVDD.n10654 2.2505
R20199 DVDD.n14193 DVDD.n14192 2.2505
R20200 DVDD.n14191 DVDD.n10655 2.2505
R20201 DVDD.n14190 DVDD.n14189 2.2505
R20202 DVDD.n14185 DVDD.n10656 2.2505
R20203 DVDD.n14181 DVDD.n14180 2.2505
R20204 DVDD.n14179 DVDD.n10657 2.2505
R20205 DVDD.n14178 DVDD.n14177 2.2505
R20206 DVDD.n14173 DVDD.n10658 2.2505
R20207 DVDD.n14169 DVDD.n14168 2.2505
R20208 DVDD.n14167 DVDD.n10659 2.2505
R20209 DVDD.n14166 DVDD.n14165 2.2505
R20210 DVDD.n14161 DVDD.n10660 2.2505
R20211 DVDD.n14157 DVDD.n14156 2.2505
R20212 DVDD.n14155 DVDD.n10661 2.2505
R20213 DVDD.n14154 DVDD.n14153 2.2505
R20214 DVDD.n14149 DVDD.n10662 2.2505
R20215 DVDD.n14145 DVDD.n14144 2.2505
R20216 DVDD.n14143 DVDD.n10663 2.2505
R20217 DVDD.n14142 DVDD.n14141 2.2505
R20218 DVDD.n14137 DVDD.n10664 2.2505
R20219 DVDD.n14133 DVDD.n14132 2.2505
R20220 DVDD.n14131 DVDD.n10665 2.2505
R20221 DVDD.n14130 DVDD.n14129 2.2505
R20222 DVDD.n14125 DVDD.n10666 2.2505
R20223 DVDD.n14121 DVDD.n14120 2.2505
R20224 DVDD.n14119 DVDD.n10667 2.2505
R20225 DVDD.n14118 DVDD.n14117 2.2505
R20226 DVDD.n14113 DVDD.n10668 2.2505
R20227 DVDD.n14109 DVDD.n14108 2.2505
R20228 DVDD.n14107 DVDD.n10669 2.2505
R20229 DVDD.n14106 DVDD.n14105 2.2505
R20230 DVDD.n14101 DVDD.n10670 2.2505
R20231 DVDD.n14097 DVDD.n14096 2.2505
R20232 DVDD.n14095 DVDD.n10671 2.2505
R20233 DVDD.n14094 DVDD.n14093 2.2505
R20234 DVDD.n14089 DVDD.n10672 2.2505
R20235 DVDD.n14085 DVDD.n14084 2.2505
R20236 DVDD.n14083 DVDD.n10673 2.2505
R20237 DVDD.n14082 DVDD.n14081 2.2505
R20238 DVDD.n14077 DVDD.n10674 2.2505
R20239 DVDD.n14073 DVDD.n14072 2.2505
R20240 DVDD.n14071 DVDD.n10675 2.2505
R20241 DVDD.n14070 DVDD.n14069 2.2505
R20242 DVDD.n14065 DVDD.n10676 2.2505
R20243 DVDD.n14061 DVDD.n14060 2.2505
R20244 DVDD.n14059 DVDD.n10677 2.2505
R20245 DVDD.n14058 DVDD.n14057 2.2505
R20246 DVDD.n14053 DVDD.n10678 2.2505
R20247 DVDD.n14049 DVDD.n14048 2.2505
R20248 DVDD.n14047 DVDD.n10679 2.2505
R20249 DVDD.n14046 DVDD.n14045 2.2505
R20250 DVDD.n14041 DVDD.n10680 2.2505
R20251 DVDD.n14037 DVDD.n14036 2.2505
R20252 DVDD.n14035 DVDD.n10681 2.2505
R20253 DVDD.n14034 DVDD.n14033 2.2505
R20254 DVDD.n14029 DVDD.n10682 2.2505
R20255 DVDD.n14025 DVDD.n14024 2.2505
R20256 DVDD.n14023 DVDD.n10685 2.2505
R20257 DVDD.n14022 DVDD.n14021 2.2505
R20258 DVDD.n14021 DVDD.n10639 2.2505
R20259 DVDD.n10685 DVDD.n10684 2.2505
R20260 DVDD.n14026 DVDD.n14025 2.2505
R20261 DVDD.n14029 DVDD.n14028 2.2505
R20262 DVDD.n14033 DVDD.n14032 2.2505
R20263 DVDD.n14030 DVDD.n10681 2.2505
R20264 DVDD.n14038 DVDD.n14037 2.2505
R20265 DVDD.n14041 DVDD.n14040 2.2505
R20266 DVDD.n14045 DVDD.n14044 2.2505
R20267 DVDD.n14042 DVDD.n10679 2.2505
R20268 DVDD.n14050 DVDD.n14049 2.2505
R20269 DVDD.n14053 DVDD.n14052 2.2505
R20270 DVDD.n14057 DVDD.n14056 2.2505
R20271 DVDD.n14054 DVDD.n10677 2.2505
R20272 DVDD.n14062 DVDD.n14061 2.2505
R20273 DVDD.n14065 DVDD.n14064 2.2505
R20274 DVDD.n14069 DVDD.n14068 2.2505
R20275 DVDD.n14066 DVDD.n10675 2.2505
R20276 DVDD.n14074 DVDD.n14073 2.2505
R20277 DVDD.n14077 DVDD.n14076 2.2505
R20278 DVDD.n14081 DVDD.n14080 2.2505
R20279 DVDD.n14078 DVDD.n10673 2.2505
R20280 DVDD.n14086 DVDD.n14085 2.2505
R20281 DVDD.n14089 DVDD.n14088 2.2505
R20282 DVDD.n14093 DVDD.n14092 2.2505
R20283 DVDD.n14090 DVDD.n10671 2.2505
R20284 DVDD.n14098 DVDD.n14097 2.2505
R20285 DVDD.n14101 DVDD.n14100 2.2505
R20286 DVDD.n14105 DVDD.n14104 2.2505
R20287 DVDD.n14102 DVDD.n10669 2.2505
R20288 DVDD.n14110 DVDD.n14109 2.2505
R20289 DVDD.n14113 DVDD.n14112 2.2505
R20290 DVDD.n14117 DVDD.n14116 2.2505
R20291 DVDD.n14114 DVDD.n10667 2.2505
R20292 DVDD.n14122 DVDD.n14121 2.2505
R20293 DVDD.n14125 DVDD.n14124 2.2505
R20294 DVDD.n14129 DVDD.n14128 2.2505
R20295 DVDD.n14126 DVDD.n10665 2.2505
R20296 DVDD.n14134 DVDD.n14133 2.2505
R20297 DVDD.n14137 DVDD.n14136 2.2505
R20298 DVDD.n14141 DVDD.n14140 2.2505
R20299 DVDD.n14138 DVDD.n10663 2.2505
R20300 DVDD.n14146 DVDD.n14145 2.2505
R20301 DVDD.n14149 DVDD.n14148 2.2505
R20302 DVDD.n14153 DVDD.n14152 2.2505
R20303 DVDD.n14150 DVDD.n10661 2.2505
R20304 DVDD.n14158 DVDD.n14157 2.2505
R20305 DVDD.n14161 DVDD.n14160 2.2505
R20306 DVDD.n14165 DVDD.n14164 2.2505
R20307 DVDD.n14162 DVDD.n10659 2.2505
R20308 DVDD.n14170 DVDD.n14169 2.2505
R20309 DVDD.n14173 DVDD.n14172 2.2505
R20310 DVDD.n14177 DVDD.n14176 2.2505
R20311 DVDD.n14174 DVDD.n10657 2.2505
R20312 DVDD.n14182 DVDD.n14181 2.2505
R20313 DVDD.n14185 DVDD.n14184 2.2505
R20314 DVDD.n14189 DVDD.n14188 2.2505
R20315 DVDD.n14186 DVDD.n10655 2.2505
R20316 DVDD.n14194 DVDD.n14193 2.2505
R20317 DVDD.n14197 DVDD.n14196 2.2505
R20318 DVDD.n14201 DVDD.n14200 2.2505
R20319 DVDD.n14198 DVDD.n10653 2.2505
R20320 DVDD.n14206 DVDD.n14205 2.2505
R20321 DVDD.n14209 DVDD.n14208 2.2505
R20322 DVDD.n14213 DVDD.n14212 2.2505
R20323 DVDD.n14210 DVDD.n10651 2.2505
R20324 DVDD.n14218 DVDD.n14217 2.2505
R20325 DVDD.n14221 DVDD.n14220 2.2505
R20326 DVDD.n14225 DVDD.n14224 2.2505
R20327 DVDD.n14222 DVDD.n10649 2.2505
R20328 DVDD.n14230 DVDD.n14229 2.2505
R20329 DVDD.n14233 DVDD.n14232 2.2505
R20330 DVDD.n14237 DVDD.n14236 2.2505
R20331 DVDD.n14234 DVDD.n10647 2.2505
R20332 DVDD.n14242 DVDD.n14241 2.2505
R20333 DVDD.n14245 DVDD.n14244 2.2505
R20334 DVDD.n14249 DVDD.n14248 2.2505
R20335 DVDD.n14246 DVDD.n10645 2.2505
R20336 DVDD.n14254 DVDD.n14253 2.2505
R20337 DVDD.n14257 DVDD.n14256 2.2505
R20338 DVDD.n14261 DVDD.n14260 2.2505
R20339 DVDD.n14258 DVDD.n10643 2.2505
R20340 DVDD.n14266 DVDD.n14265 2.2505
R20341 DVDD.n14268 DVDD.n10641 2.2505
R20342 DVDD.n11050 DVDD.n11049 2.2505
R20343 DVDD.n10717 DVDD.n10716 2.2505
R20344 DVDD.n11039 DVDD.n10718 2.2505
R20345 DVDD.n11041 DVDD.n11040 2.2505
R20346 DVDD.n11038 DVDD.n10720 2.2505
R20347 DVDD.n11037 DVDD.n11036 2.2505
R20348 DVDD.n10722 DVDD.n10721 2.2505
R20349 DVDD.n11028 DVDD.n11027 2.2505
R20350 DVDD.n11026 DVDD.n10724 2.2505
R20351 DVDD.n11025 DVDD.n11024 2.2505
R20352 DVDD.n10726 DVDD.n10725 2.2505
R20353 DVDD.n11016 DVDD.n11015 2.2505
R20354 DVDD.n11014 DVDD.n10728 2.2505
R20355 DVDD.n11013 DVDD.n11012 2.2505
R20356 DVDD.n10730 DVDD.n10729 2.2505
R20357 DVDD.n11004 DVDD.n11003 2.2505
R20358 DVDD.n11002 DVDD.n10732 2.2505
R20359 DVDD.n11001 DVDD.n11000 2.2505
R20360 DVDD.n10734 DVDD.n10733 2.2505
R20361 DVDD.n10992 DVDD.n10991 2.2505
R20362 DVDD.n10990 DVDD.n10736 2.2505
R20363 DVDD.n10989 DVDD.n10988 2.2505
R20364 DVDD.n10738 DVDD.n10737 2.2505
R20365 DVDD.n10980 DVDD.n10979 2.2505
R20366 DVDD.n10978 DVDD.n10740 2.2505
R20367 DVDD.n10977 DVDD.n10976 2.2505
R20368 DVDD.n10742 DVDD.n10741 2.2505
R20369 DVDD.n10968 DVDD.n10967 2.2505
R20370 DVDD.n10966 DVDD.n10744 2.2505
R20371 DVDD.n10965 DVDD.n10964 2.2505
R20372 DVDD.n10746 DVDD.n10745 2.2505
R20373 DVDD.n10956 DVDD.n10955 2.2505
R20374 DVDD.n10954 DVDD.n10748 2.2505
R20375 DVDD.n10953 DVDD.n10952 2.2505
R20376 DVDD.n10750 DVDD.n10749 2.2505
R20377 DVDD.n10944 DVDD.n10943 2.2505
R20378 DVDD.n10942 DVDD.n10752 2.2505
R20379 DVDD.n10941 DVDD.n10940 2.2505
R20380 DVDD.n10754 DVDD.n10753 2.2505
R20381 DVDD.n10932 DVDD.n10931 2.2505
R20382 DVDD.n10930 DVDD.n10756 2.2505
R20383 DVDD.n10929 DVDD.n10928 2.2505
R20384 DVDD.n10758 DVDD.n10757 2.2505
R20385 DVDD.n10920 DVDD.n10919 2.2505
R20386 DVDD.n10918 DVDD.n10760 2.2505
R20387 DVDD.n10917 DVDD.n10916 2.2505
R20388 DVDD.n10762 DVDD.n10761 2.2505
R20389 DVDD.n10908 DVDD.n10907 2.2505
R20390 DVDD.n10906 DVDD.n10764 2.2505
R20391 DVDD.n10905 DVDD.n10904 2.2505
R20392 DVDD.n10766 DVDD.n10765 2.2505
R20393 DVDD.n10896 DVDD.n10895 2.2505
R20394 DVDD.n10894 DVDD.n10768 2.2505
R20395 DVDD.n10893 DVDD.n10892 2.2505
R20396 DVDD.n10770 DVDD.n10769 2.2505
R20397 DVDD.n10884 DVDD.n10883 2.2505
R20398 DVDD.n10882 DVDD.n10772 2.2505
R20399 DVDD.n10881 DVDD.n10880 2.2505
R20400 DVDD.n10774 DVDD.n10773 2.2505
R20401 DVDD.n10872 DVDD.n10871 2.2505
R20402 DVDD.n10870 DVDD.n10776 2.2505
R20403 DVDD.n10869 DVDD.n10868 2.2505
R20404 DVDD.n10778 DVDD.n10777 2.2505
R20405 DVDD.n10860 DVDD.n10859 2.2505
R20406 DVDD.n10858 DVDD.n10780 2.2505
R20407 DVDD.n10857 DVDD.n10856 2.2505
R20408 DVDD.n10782 DVDD.n10781 2.2505
R20409 DVDD.n10848 DVDD.n10847 2.2505
R20410 DVDD.n10846 DVDD.n10784 2.2505
R20411 DVDD.n10845 DVDD.n10844 2.2505
R20412 DVDD.n10786 DVDD.n10785 2.2505
R20413 DVDD.n10836 DVDD.n10835 2.2505
R20414 DVDD.n10834 DVDD.n10788 2.2505
R20415 DVDD.n10833 DVDD.n10832 2.2505
R20416 DVDD.n10790 DVDD.n10789 2.2505
R20417 DVDD.n10824 DVDD.n10823 2.2505
R20418 DVDD.n10822 DVDD.n10792 2.2505
R20419 DVDD.n10821 DVDD.n10820 2.2505
R20420 DVDD.n10794 DVDD.n10793 2.2505
R20421 DVDD.n10812 DVDD.n10811 2.2505
R20422 DVDD.n10810 DVDD.n10796 2.2505
R20423 DVDD.n10809 DVDD.n10808 2.2505
R20424 DVDD.n10798 DVDD.n10797 2.2505
R20425 DVDD.n10800 DVDD.n10799 2.2505
R20426 DVDD.n10801 DVDD.n10800 2.2505
R20427 DVDD.n10803 DVDD.n10798 2.2505
R20428 DVDD.n10808 DVDD.n10807 2.2505
R20429 DVDD.n10805 DVDD.n10796 2.2505
R20430 DVDD.n10813 DVDD.n10812 2.2505
R20431 DVDD.n10815 DVDD.n10794 2.2505
R20432 DVDD.n10820 DVDD.n10819 2.2505
R20433 DVDD.n10817 DVDD.n10792 2.2505
R20434 DVDD.n10825 DVDD.n10824 2.2505
R20435 DVDD.n10827 DVDD.n10790 2.2505
R20436 DVDD.n10832 DVDD.n10831 2.2505
R20437 DVDD.n10829 DVDD.n10788 2.2505
R20438 DVDD.n10837 DVDD.n10836 2.2505
R20439 DVDD.n10839 DVDD.n10786 2.2505
R20440 DVDD.n10844 DVDD.n10843 2.2505
R20441 DVDD.n10841 DVDD.n10784 2.2505
R20442 DVDD.n10849 DVDD.n10848 2.2505
R20443 DVDD.n10851 DVDD.n10782 2.2505
R20444 DVDD.n10856 DVDD.n10855 2.2505
R20445 DVDD.n10853 DVDD.n10780 2.2505
R20446 DVDD.n10861 DVDD.n10860 2.2505
R20447 DVDD.n10863 DVDD.n10778 2.2505
R20448 DVDD.n10868 DVDD.n10867 2.2505
R20449 DVDD.n10865 DVDD.n10776 2.2505
R20450 DVDD.n10873 DVDD.n10872 2.2505
R20451 DVDD.n10875 DVDD.n10774 2.2505
R20452 DVDD.n10880 DVDD.n10879 2.2505
R20453 DVDD.n10877 DVDD.n10772 2.2505
R20454 DVDD.n10885 DVDD.n10884 2.2505
R20455 DVDD.n10887 DVDD.n10770 2.2505
R20456 DVDD.n10892 DVDD.n10891 2.2505
R20457 DVDD.n10889 DVDD.n10768 2.2505
R20458 DVDD.n10897 DVDD.n10896 2.2505
R20459 DVDD.n10899 DVDD.n10766 2.2505
R20460 DVDD.n10904 DVDD.n10903 2.2505
R20461 DVDD.n10901 DVDD.n10764 2.2505
R20462 DVDD.n10909 DVDD.n10908 2.2505
R20463 DVDD.n10911 DVDD.n10762 2.2505
R20464 DVDD.n10916 DVDD.n10915 2.2505
R20465 DVDD.n10913 DVDD.n10760 2.2505
R20466 DVDD.n10921 DVDD.n10920 2.2505
R20467 DVDD.n10923 DVDD.n10758 2.2505
R20468 DVDD.n10928 DVDD.n10927 2.2505
R20469 DVDD.n10925 DVDD.n10756 2.2505
R20470 DVDD.n10933 DVDD.n10932 2.2505
R20471 DVDD.n10935 DVDD.n10754 2.2505
R20472 DVDD.n10940 DVDD.n10939 2.2505
R20473 DVDD.n10937 DVDD.n10752 2.2505
R20474 DVDD.n10945 DVDD.n10944 2.2505
R20475 DVDD.n10947 DVDD.n10750 2.2505
R20476 DVDD.n10952 DVDD.n10951 2.2505
R20477 DVDD.n10949 DVDD.n10748 2.2505
R20478 DVDD.n10957 DVDD.n10956 2.2505
R20479 DVDD.n10959 DVDD.n10746 2.2505
R20480 DVDD.n10964 DVDD.n10963 2.2505
R20481 DVDD.n10961 DVDD.n10744 2.2505
R20482 DVDD.n10969 DVDD.n10968 2.2505
R20483 DVDD.n10971 DVDD.n10742 2.2505
R20484 DVDD.n10976 DVDD.n10975 2.2505
R20485 DVDD.n10973 DVDD.n10740 2.2505
R20486 DVDD.n10981 DVDD.n10980 2.2505
R20487 DVDD.n10983 DVDD.n10738 2.2505
R20488 DVDD.n10988 DVDD.n10987 2.2505
R20489 DVDD.n10985 DVDD.n10736 2.2505
R20490 DVDD.n10993 DVDD.n10992 2.2505
R20491 DVDD.n10995 DVDD.n10734 2.2505
R20492 DVDD.n11000 DVDD.n10999 2.2505
R20493 DVDD.n10997 DVDD.n10732 2.2505
R20494 DVDD.n11005 DVDD.n11004 2.2505
R20495 DVDD.n11007 DVDD.n10730 2.2505
R20496 DVDD.n11012 DVDD.n11011 2.2505
R20497 DVDD.n11009 DVDD.n10728 2.2505
R20498 DVDD.n11017 DVDD.n11016 2.2505
R20499 DVDD.n11019 DVDD.n10726 2.2505
R20500 DVDD.n11024 DVDD.n11023 2.2505
R20501 DVDD.n11021 DVDD.n10724 2.2505
R20502 DVDD.n11029 DVDD.n11028 2.2505
R20503 DVDD.n11031 DVDD.n10722 2.2505
R20504 DVDD.n11036 DVDD.n11035 2.2505
R20505 DVDD.n11033 DVDD.n10720 2.2505
R20506 DVDD.n11042 DVDD.n11041 2.2505
R20507 DVDD.n11044 DVDD.n10718 2.2505
R20508 DVDD.n11046 DVDD.n10717 2.2505
R20509 DVDD.n11049 DVDD.n11048 2.2505
R20510 DVDD.n13998 DVDD.n13997 2.2505
R20511 DVDD.n13996 DVDD.n11151 2.2505
R20512 DVDD.n13995 DVDD.n13994 2.2505
R20513 DVDD.n13992 DVDD.n11152 2.2505
R20514 DVDD.n13990 DVDD.n13988 2.2505
R20515 DVDD.n13987 DVDD.n11154 2.2505
R20516 DVDD.n13986 DVDD.n13985 2.2505
R20517 DVDD.n13983 DVDD.n11155 2.2505
R20518 DVDD.n13981 DVDD.n13979 2.2505
R20519 DVDD.n13978 DVDD.n11157 2.2505
R20520 DVDD.n13977 DVDD.n13976 2.2505
R20521 DVDD.n13974 DVDD.n11158 2.2505
R20522 DVDD.n13972 DVDD.n13970 2.2505
R20523 DVDD.n13969 DVDD.n11160 2.2505
R20524 DVDD.n13968 DVDD.n13967 2.2505
R20525 DVDD.n13965 DVDD.n11161 2.2505
R20526 DVDD.n13963 DVDD.n13961 2.2505
R20527 DVDD.n13960 DVDD.n11163 2.2505
R20528 DVDD.n13959 DVDD.n13958 2.2505
R20529 DVDD.n13956 DVDD.n11164 2.2505
R20530 DVDD.n13954 DVDD.n13952 2.2505
R20531 DVDD.n13951 DVDD.n11166 2.2505
R20532 DVDD.n13950 DVDD.n13949 2.2505
R20533 DVDD.n13947 DVDD.n11167 2.2505
R20534 DVDD.n13945 DVDD.n13943 2.2505
R20535 DVDD.n13942 DVDD.n11169 2.2505
R20536 DVDD.n13941 DVDD.n13940 2.2505
R20537 DVDD.n13938 DVDD.n11170 2.2505
R20538 DVDD.n13936 DVDD.n13934 2.2505
R20539 DVDD.n13933 DVDD.n11172 2.2505
R20540 DVDD.n13932 DVDD.n13931 2.2505
R20541 DVDD.n13929 DVDD.n11173 2.2505
R20542 DVDD.n13927 DVDD.n13925 2.2505
R20543 DVDD.n13924 DVDD.n11175 2.2505
R20544 DVDD.n13923 DVDD.n13922 2.2505
R20545 DVDD.n13920 DVDD.n11176 2.2505
R20546 DVDD.n13918 DVDD.n13916 2.2505
R20547 DVDD.n13915 DVDD.n11178 2.2505
R20548 DVDD.n13914 DVDD.n13913 2.2505
R20549 DVDD.n13911 DVDD.n11179 2.2505
R20550 DVDD.n13909 DVDD.n13907 2.2505
R20551 DVDD.n13906 DVDD.n11181 2.2505
R20552 DVDD.n13905 DVDD.n13904 2.2505
R20553 DVDD.n13902 DVDD.n11182 2.2505
R20554 DVDD.n13900 DVDD.n13898 2.2505
R20555 DVDD.n13897 DVDD.n11184 2.2505
R20556 DVDD.n13896 DVDD.n13895 2.2505
R20557 DVDD.n13893 DVDD.n11185 2.2505
R20558 DVDD.n13891 DVDD.n13889 2.2505
R20559 DVDD.n13888 DVDD.n11187 2.2505
R20560 DVDD.n13887 DVDD.n13886 2.2505
R20561 DVDD.n13884 DVDD.n11188 2.2505
R20562 DVDD.n13882 DVDD.n13880 2.2505
R20563 DVDD.n13879 DVDD.n11190 2.2505
R20564 DVDD.n13878 DVDD.n13877 2.2505
R20565 DVDD.n13875 DVDD.n11191 2.2505
R20566 DVDD.n13873 DVDD.n13871 2.2505
R20567 DVDD.n13870 DVDD.n11193 2.2505
R20568 DVDD.n13869 DVDD.n13868 2.2505
R20569 DVDD.n13866 DVDD.n11194 2.2505
R20570 DVDD.n13864 DVDD.n13862 2.2505
R20571 DVDD.n13861 DVDD.n11196 2.2505
R20572 DVDD.n13860 DVDD.n13859 2.2505
R20573 DVDD.n13857 DVDD.n11197 2.2505
R20574 DVDD.n13855 DVDD.n13853 2.2505
R20575 DVDD.n13852 DVDD.n11199 2.2505
R20576 DVDD.n13851 DVDD.n13850 2.2505
R20577 DVDD.n13848 DVDD.n11200 2.2505
R20578 DVDD.n13846 DVDD.n13844 2.2505
R20579 DVDD.n13843 DVDD.n11202 2.2505
R20580 DVDD.n13842 DVDD.n13841 2.2505
R20581 DVDD.n13839 DVDD.n11203 2.2505
R20582 DVDD.n13837 DVDD.n13835 2.2505
R20583 DVDD.n13834 DVDD.n11205 2.2505
R20584 DVDD.n13833 DVDD.n13832 2.2505
R20585 DVDD.n13830 DVDD.n11206 2.2505
R20586 DVDD.n13828 DVDD.n13826 2.2505
R20587 DVDD.n13825 DVDD.n11208 2.2505
R20588 DVDD.n13824 DVDD.n13823 2.2505
R20589 DVDD.n13821 DVDD.n11209 2.2505
R20590 DVDD.n13819 DVDD.n13817 2.2505
R20591 DVDD.n13816 DVDD.n11211 2.2505
R20592 DVDD.n13815 DVDD.n13814 2.2505
R20593 DVDD.n13813 DVDD.n11106 2.2505
R20594 DVDD.n14001 DVDD.n11106 2.2505
R20595 DVDD.n13814 DVDD.n11104 2.2505
R20596 DVDD.n11211 DVDD.n11210 2.2505
R20597 DVDD.n13819 DVDD.n13818 2.2505
R20598 DVDD.n13821 DVDD.n13820 2.2505
R20599 DVDD.n13823 DVDD.n13822 2.2505
R20600 DVDD.n11208 DVDD.n11207 2.2505
R20601 DVDD.n13828 DVDD.n13827 2.2505
R20602 DVDD.n13830 DVDD.n13829 2.2505
R20603 DVDD.n13832 DVDD.n13831 2.2505
R20604 DVDD.n11205 DVDD.n11204 2.2505
R20605 DVDD.n13837 DVDD.n13836 2.2505
R20606 DVDD.n13839 DVDD.n13838 2.2505
R20607 DVDD.n13841 DVDD.n13840 2.2505
R20608 DVDD.n11202 DVDD.n11201 2.2505
R20609 DVDD.n13846 DVDD.n13845 2.2505
R20610 DVDD.n13848 DVDD.n13847 2.2505
R20611 DVDD.n13850 DVDD.n13849 2.2505
R20612 DVDD.n11199 DVDD.n11198 2.2505
R20613 DVDD.n13855 DVDD.n13854 2.2505
R20614 DVDD.n13857 DVDD.n13856 2.2505
R20615 DVDD.n13859 DVDD.n13858 2.2505
R20616 DVDD.n11196 DVDD.n11195 2.2505
R20617 DVDD.n13864 DVDD.n13863 2.2505
R20618 DVDD.n13866 DVDD.n13865 2.2505
R20619 DVDD.n13868 DVDD.n13867 2.2505
R20620 DVDD.n11193 DVDD.n11192 2.2505
R20621 DVDD.n13873 DVDD.n13872 2.2505
R20622 DVDD.n13875 DVDD.n13874 2.2505
R20623 DVDD.n13877 DVDD.n13876 2.2505
R20624 DVDD.n11190 DVDD.n11189 2.2505
R20625 DVDD.n13882 DVDD.n13881 2.2505
R20626 DVDD.n13884 DVDD.n13883 2.2505
R20627 DVDD.n13886 DVDD.n13885 2.2505
R20628 DVDD.n11187 DVDD.n11186 2.2505
R20629 DVDD.n13891 DVDD.n13890 2.2505
R20630 DVDD.n13893 DVDD.n13892 2.2505
R20631 DVDD.n13895 DVDD.n13894 2.2505
R20632 DVDD.n11184 DVDD.n11183 2.2505
R20633 DVDD.n13900 DVDD.n13899 2.2505
R20634 DVDD.n13902 DVDD.n13901 2.2505
R20635 DVDD.n13904 DVDD.n13903 2.2505
R20636 DVDD.n11181 DVDD.n11180 2.2505
R20637 DVDD.n13909 DVDD.n13908 2.2505
R20638 DVDD.n13911 DVDD.n13910 2.2505
R20639 DVDD.n13913 DVDD.n13912 2.2505
R20640 DVDD.n11178 DVDD.n11177 2.2505
R20641 DVDD.n13918 DVDD.n13917 2.2505
R20642 DVDD.n13920 DVDD.n13919 2.2505
R20643 DVDD.n13922 DVDD.n13921 2.2505
R20644 DVDD.n11175 DVDD.n11174 2.2505
R20645 DVDD.n13927 DVDD.n13926 2.2505
R20646 DVDD.n13929 DVDD.n13928 2.2505
R20647 DVDD.n13931 DVDD.n13930 2.2505
R20648 DVDD.n11172 DVDD.n11171 2.2505
R20649 DVDD.n13936 DVDD.n13935 2.2505
R20650 DVDD.n13938 DVDD.n13937 2.2505
R20651 DVDD.n13940 DVDD.n13939 2.2505
R20652 DVDD.n11169 DVDD.n11168 2.2505
R20653 DVDD.n13945 DVDD.n13944 2.2505
R20654 DVDD.n13947 DVDD.n13946 2.2505
R20655 DVDD.n13949 DVDD.n13948 2.2505
R20656 DVDD.n11166 DVDD.n11165 2.2505
R20657 DVDD.n13954 DVDD.n13953 2.2505
R20658 DVDD.n13956 DVDD.n13955 2.2505
R20659 DVDD.n13958 DVDD.n13957 2.2505
R20660 DVDD.n11163 DVDD.n11162 2.2505
R20661 DVDD.n13963 DVDD.n13962 2.2505
R20662 DVDD.n13965 DVDD.n13964 2.2505
R20663 DVDD.n13967 DVDD.n13966 2.2505
R20664 DVDD.n11160 DVDD.n11159 2.2505
R20665 DVDD.n13972 DVDD.n13971 2.2505
R20666 DVDD.n13974 DVDD.n13973 2.2505
R20667 DVDD.n13976 DVDD.n13975 2.2505
R20668 DVDD.n11157 DVDD.n11156 2.2505
R20669 DVDD.n13981 DVDD.n13980 2.2505
R20670 DVDD.n13983 DVDD.n13982 2.2505
R20671 DVDD.n13985 DVDD.n13984 2.2505
R20672 DVDD.n11154 DVDD.n11153 2.2505
R20673 DVDD.n13990 DVDD.n13989 2.2505
R20674 DVDD.n13992 DVDD.n13991 2.2505
R20675 DVDD.n13994 DVDD.n13993 2.2505
R20676 DVDD.n11151 DVDD.n11150 2.2505
R20677 DVDD.n13999 DVDD.n13998 2.2505
R20678 DVDD.n13793 DVDD.n11278 2.2505
R20679 DVDD.n13795 DVDD.n13794 2.2505
R20680 DVDD.n11564 DVDD.n11280 2.2505
R20681 DVDD.n11563 DVDD.n11562 2.2505
R20682 DVDD.n11558 DVDD.n11281 2.2505
R20683 DVDD.n11554 DVDD.n11553 2.2505
R20684 DVDD.n11552 DVDD.n11282 2.2505
R20685 DVDD.n11551 DVDD.n11550 2.2505
R20686 DVDD.n11546 DVDD.n11283 2.2505
R20687 DVDD.n11542 DVDD.n11541 2.2505
R20688 DVDD.n11540 DVDD.n11284 2.2505
R20689 DVDD.n11539 DVDD.n11538 2.2505
R20690 DVDD.n11534 DVDD.n11285 2.2505
R20691 DVDD.n11530 DVDD.n11529 2.2505
R20692 DVDD.n11528 DVDD.n11286 2.2505
R20693 DVDD.n11527 DVDD.n11526 2.2505
R20694 DVDD.n11522 DVDD.n11287 2.2505
R20695 DVDD.n11518 DVDD.n11517 2.2505
R20696 DVDD.n11516 DVDD.n11288 2.2505
R20697 DVDD.n11515 DVDD.n11514 2.2505
R20698 DVDD.n11510 DVDD.n11289 2.2505
R20699 DVDD.n11506 DVDD.n11505 2.2505
R20700 DVDD.n11504 DVDD.n11290 2.2505
R20701 DVDD.n11503 DVDD.n11502 2.2505
R20702 DVDD.n11498 DVDD.n11291 2.2505
R20703 DVDD.n11494 DVDD.n11493 2.2505
R20704 DVDD.n11492 DVDD.n11292 2.2505
R20705 DVDD.n11491 DVDD.n11490 2.2505
R20706 DVDD.n11486 DVDD.n11293 2.2505
R20707 DVDD.n11482 DVDD.n11481 2.2505
R20708 DVDD.n11480 DVDD.n11294 2.2505
R20709 DVDD.n11479 DVDD.n11478 2.2505
R20710 DVDD.n11474 DVDD.n11295 2.2505
R20711 DVDD.n11470 DVDD.n11469 2.2505
R20712 DVDD.n11468 DVDD.n11296 2.2505
R20713 DVDD.n11467 DVDD.n11466 2.2505
R20714 DVDD.n11462 DVDD.n11297 2.2505
R20715 DVDD.n11458 DVDD.n11457 2.2505
R20716 DVDD.n11456 DVDD.n11298 2.2505
R20717 DVDD.n11455 DVDD.n11454 2.2505
R20718 DVDD.n11450 DVDD.n11299 2.2505
R20719 DVDD.n11446 DVDD.n11445 2.2505
R20720 DVDD.n11444 DVDD.n11300 2.2505
R20721 DVDD.n11443 DVDD.n11442 2.2505
R20722 DVDD.n11438 DVDD.n11301 2.2505
R20723 DVDD.n11434 DVDD.n11433 2.2505
R20724 DVDD.n11432 DVDD.n11302 2.2505
R20725 DVDD.n11431 DVDD.n11430 2.2505
R20726 DVDD.n11426 DVDD.n11303 2.2505
R20727 DVDD.n11422 DVDD.n11421 2.2505
R20728 DVDD.n11420 DVDD.n11304 2.2505
R20729 DVDD.n11419 DVDD.n11418 2.2505
R20730 DVDD.n11414 DVDD.n11305 2.2505
R20731 DVDD.n11410 DVDD.n11409 2.2505
R20732 DVDD.n11408 DVDD.n11306 2.2505
R20733 DVDD.n11407 DVDD.n11406 2.2505
R20734 DVDD.n11402 DVDD.n11307 2.2505
R20735 DVDD.n11398 DVDD.n11397 2.2505
R20736 DVDD.n11396 DVDD.n11308 2.2505
R20737 DVDD.n11395 DVDD.n11394 2.2505
R20738 DVDD.n11390 DVDD.n11309 2.2505
R20739 DVDD.n11386 DVDD.n11385 2.2505
R20740 DVDD.n11384 DVDD.n11310 2.2505
R20741 DVDD.n11383 DVDD.n11382 2.2505
R20742 DVDD.n11378 DVDD.n11311 2.2505
R20743 DVDD.n11374 DVDD.n11373 2.2505
R20744 DVDD.n11372 DVDD.n11312 2.2505
R20745 DVDD.n11371 DVDD.n11370 2.2505
R20746 DVDD.n11366 DVDD.n11313 2.2505
R20747 DVDD.n11362 DVDD.n11361 2.2505
R20748 DVDD.n11360 DVDD.n11314 2.2505
R20749 DVDD.n11359 DVDD.n11358 2.2505
R20750 DVDD.n11354 DVDD.n11315 2.2505
R20751 DVDD.n11350 DVDD.n11349 2.2505
R20752 DVDD.n11348 DVDD.n11316 2.2505
R20753 DVDD.n11347 DVDD.n11346 2.2505
R20754 DVDD.n11342 DVDD.n11317 2.2505
R20755 DVDD.n11338 DVDD.n11337 2.2505
R20756 DVDD.n11336 DVDD.n11318 2.2505
R20757 DVDD.n11335 DVDD.n11334 2.2505
R20758 DVDD.n11330 DVDD.n11319 2.2505
R20759 DVDD.n11326 DVDD.n11325 2.2505
R20760 DVDD.n11324 DVDD.n11323 2.2505
R20761 DVDD.n11320 DVDD.n11229 2.2505
R20762 DVDD.n11320 DVDD.n11275 2.2505
R20763 DVDD.n11323 DVDD.n11322 2.2505
R20764 DVDD.n11327 DVDD.n11326 2.2505
R20765 DVDD.n11330 DVDD.n11329 2.2505
R20766 DVDD.n11334 DVDD.n11333 2.2505
R20767 DVDD.n11331 DVDD.n11318 2.2505
R20768 DVDD.n11339 DVDD.n11338 2.2505
R20769 DVDD.n11342 DVDD.n11341 2.2505
R20770 DVDD.n11346 DVDD.n11345 2.2505
R20771 DVDD.n11343 DVDD.n11316 2.2505
R20772 DVDD.n11351 DVDD.n11350 2.2505
R20773 DVDD.n11354 DVDD.n11353 2.2505
R20774 DVDD.n11358 DVDD.n11357 2.2505
R20775 DVDD.n11355 DVDD.n11314 2.2505
R20776 DVDD.n11363 DVDD.n11362 2.2505
R20777 DVDD.n11366 DVDD.n11365 2.2505
R20778 DVDD.n11370 DVDD.n11369 2.2505
R20779 DVDD.n11367 DVDD.n11312 2.2505
R20780 DVDD.n11375 DVDD.n11374 2.2505
R20781 DVDD.n11378 DVDD.n11377 2.2505
R20782 DVDD.n11382 DVDD.n11381 2.2505
R20783 DVDD.n11379 DVDD.n11310 2.2505
R20784 DVDD.n11387 DVDD.n11386 2.2505
R20785 DVDD.n11390 DVDD.n11389 2.2505
R20786 DVDD.n11394 DVDD.n11393 2.2505
R20787 DVDD.n11391 DVDD.n11308 2.2505
R20788 DVDD.n11399 DVDD.n11398 2.2505
R20789 DVDD.n11402 DVDD.n11401 2.2505
R20790 DVDD.n11406 DVDD.n11405 2.2505
R20791 DVDD.n11403 DVDD.n11306 2.2505
R20792 DVDD.n11411 DVDD.n11410 2.2505
R20793 DVDD.n11414 DVDD.n11413 2.2505
R20794 DVDD.n11418 DVDD.n11417 2.2505
R20795 DVDD.n11415 DVDD.n11304 2.2505
R20796 DVDD.n11423 DVDD.n11422 2.2505
R20797 DVDD.n11426 DVDD.n11425 2.2505
R20798 DVDD.n11430 DVDD.n11429 2.2505
R20799 DVDD.n11427 DVDD.n11302 2.2505
R20800 DVDD.n11435 DVDD.n11434 2.2505
R20801 DVDD.n11438 DVDD.n11437 2.2505
R20802 DVDD.n11442 DVDD.n11441 2.2505
R20803 DVDD.n11439 DVDD.n11300 2.2505
R20804 DVDD.n11447 DVDD.n11446 2.2505
R20805 DVDD.n11450 DVDD.n11449 2.2505
R20806 DVDD.n11454 DVDD.n11453 2.2505
R20807 DVDD.n11451 DVDD.n11298 2.2505
R20808 DVDD.n11459 DVDD.n11458 2.2505
R20809 DVDD.n11462 DVDD.n11461 2.2505
R20810 DVDD.n11466 DVDD.n11465 2.2505
R20811 DVDD.n11463 DVDD.n11296 2.2505
R20812 DVDD.n11471 DVDD.n11470 2.2505
R20813 DVDD.n11474 DVDD.n11473 2.2505
R20814 DVDD.n11478 DVDD.n11477 2.2505
R20815 DVDD.n11475 DVDD.n11294 2.2505
R20816 DVDD.n11483 DVDD.n11482 2.2505
R20817 DVDD.n11486 DVDD.n11485 2.2505
R20818 DVDD.n11490 DVDD.n11489 2.2505
R20819 DVDD.n11487 DVDD.n11292 2.2505
R20820 DVDD.n11495 DVDD.n11494 2.2505
R20821 DVDD.n11498 DVDD.n11497 2.2505
R20822 DVDD.n11502 DVDD.n11501 2.2505
R20823 DVDD.n11499 DVDD.n11290 2.2505
R20824 DVDD.n11507 DVDD.n11506 2.2505
R20825 DVDD.n11510 DVDD.n11509 2.2505
R20826 DVDD.n11514 DVDD.n11513 2.2505
R20827 DVDD.n11511 DVDD.n11288 2.2505
R20828 DVDD.n11519 DVDD.n11518 2.2505
R20829 DVDD.n11522 DVDD.n11521 2.2505
R20830 DVDD.n11526 DVDD.n11525 2.2505
R20831 DVDD.n11523 DVDD.n11286 2.2505
R20832 DVDD.n11531 DVDD.n11530 2.2505
R20833 DVDD.n11534 DVDD.n11533 2.2505
R20834 DVDD.n11538 DVDD.n11537 2.2505
R20835 DVDD.n11535 DVDD.n11284 2.2505
R20836 DVDD.n11543 DVDD.n11542 2.2505
R20837 DVDD.n11546 DVDD.n11545 2.2505
R20838 DVDD.n11550 DVDD.n11549 2.2505
R20839 DVDD.n11547 DVDD.n11282 2.2505
R20840 DVDD.n11555 DVDD.n11554 2.2505
R20841 DVDD.n11558 DVDD.n11557 2.2505
R20842 DVDD.n11562 DVDD.n11561 2.2505
R20843 DVDD.n11559 DVDD.n11280 2.2505
R20844 DVDD.n13796 DVDD.n13795 2.2505
R20845 DVDD.n13798 DVDD.n11278 2.2505
R20846 DVDD.n13771 DVDD.n11633 2.2505
R20847 DVDD.n13773 DVDD.n13772 2.2505
R20848 DVDD.n11918 DVDD.n11634 2.2505
R20849 DVDD.n11917 DVDD.n11916 2.2505
R20850 DVDD.n11912 DVDD.n11635 2.2505
R20851 DVDD.n11908 DVDD.n11907 2.2505
R20852 DVDD.n11906 DVDD.n11636 2.2505
R20853 DVDD.n11905 DVDD.n11904 2.2505
R20854 DVDD.n11900 DVDD.n11637 2.2505
R20855 DVDD.n11896 DVDD.n11895 2.2505
R20856 DVDD.n11894 DVDD.n11638 2.2505
R20857 DVDD.n11893 DVDD.n11892 2.2505
R20858 DVDD.n11888 DVDD.n11639 2.2505
R20859 DVDD.n11884 DVDD.n11883 2.2505
R20860 DVDD.n11882 DVDD.n11640 2.2505
R20861 DVDD.n11881 DVDD.n11880 2.2505
R20862 DVDD.n11876 DVDD.n11641 2.2505
R20863 DVDD.n11872 DVDD.n11871 2.2505
R20864 DVDD.n11870 DVDD.n11642 2.2505
R20865 DVDD.n11869 DVDD.n11868 2.2505
R20866 DVDD.n11864 DVDD.n11643 2.2505
R20867 DVDD.n11860 DVDD.n11859 2.2505
R20868 DVDD.n11858 DVDD.n11644 2.2505
R20869 DVDD.n11857 DVDD.n11856 2.2505
R20870 DVDD.n11852 DVDD.n11645 2.2505
R20871 DVDD.n11848 DVDD.n11847 2.2505
R20872 DVDD.n11846 DVDD.n11646 2.2505
R20873 DVDD.n11845 DVDD.n11844 2.2505
R20874 DVDD.n11840 DVDD.n11647 2.2505
R20875 DVDD.n11836 DVDD.n11835 2.2505
R20876 DVDD.n11834 DVDD.n11648 2.2505
R20877 DVDD.n11833 DVDD.n11832 2.2505
R20878 DVDD.n11828 DVDD.n11649 2.2505
R20879 DVDD.n11824 DVDD.n11823 2.2505
R20880 DVDD.n11822 DVDD.n11650 2.2505
R20881 DVDD.n11821 DVDD.n11820 2.2505
R20882 DVDD.n11816 DVDD.n11651 2.2505
R20883 DVDD.n11812 DVDD.n11811 2.2505
R20884 DVDD.n11810 DVDD.n11652 2.2505
R20885 DVDD.n11809 DVDD.n11808 2.2505
R20886 DVDD.n11804 DVDD.n11653 2.2505
R20887 DVDD.n11800 DVDD.n11799 2.2505
R20888 DVDD.n11798 DVDD.n11654 2.2505
R20889 DVDD.n11797 DVDD.n11796 2.2505
R20890 DVDD.n11792 DVDD.n11655 2.2505
R20891 DVDD.n11788 DVDD.n11787 2.2505
R20892 DVDD.n11786 DVDD.n11656 2.2505
R20893 DVDD.n11785 DVDD.n11784 2.2505
R20894 DVDD.n11780 DVDD.n11657 2.2505
R20895 DVDD.n11776 DVDD.n11775 2.2505
R20896 DVDD.n11774 DVDD.n11658 2.2505
R20897 DVDD.n11773 DVDD.n11772 2.2505
R20898 DVDD.n11768 DVDD.n11659 2.2505
R20899 DVDD.n11764 DVDD.n11763 2.2505
R20900 DVDD.n11762 DVDD.n11660 2.2505
R20901 DVDD.n11761 DVDD.n11760 2.2505
R20902 DVDD.n11756 DVDD.n11661 2.2505
R20903 DVDD.n11752 DVDD.n11751 2.2505
R20904 DVDD.n11750 DVDD.n11662 2.2505
R20905 DVDD.n11749 DVDD.n11748 2.2505
R20906 DVDD.n11744 DVDD.n11663 2.2505
R20907 DVDD.n11740 DVDD.n11739 2.2505
R20908 DVDD.n11738 DVDD.n11664 2.2505
R20909 DVDD.n11737 DVDD.n11736 2.2505
R20910 DVDD.n11732 DVDD.n11665 2.2505
R20911 DVDD.n11728 DVDD.n11727 2.2505
R20912 DVDD.n11726 DVDD.n11666 2.2505
R20913 DVDD.n11725 DVDD.n11724 2.2505
R20914 DVDD.n11720 DVDD.n11667 2.2505
R20915 DVDD.n11716 DVDD.n11715 2.2505
R20916 DVDD.n11714 DVDD.n11668 2.2505
R20917 DVDD.n11713 DVDD.n11712 2.2505
R20918 DVDD.n11708 DVDD.n11669 2.2505
R20919 DVDD.n11704 DVDD.n11703 2.2505
R20920 DVDD.n11702 DVDD.n11670 2.2505
R20921 DVDD.n11701 DVDD.n11700 2.2505
R20922 DVDD.n11696 DVDD.n11671 2.2505
R20923 DVDD.n11692 DVDD.n11691 2.2505
R20924 DVDD.n11690 DVDD.n11672 2.2505
R20925 DVDD.n11689 DVDD.n11688 2.2505
R20926 DVDD.n11684 DVDD.n11673 2.2505
R20927 DVDD.n11680 DVDD.n11679 2.2505
R20928 DVDD.n11678 DVDD.n11677 2.2505
R20929 DVDD.n11674 DVDD.n11584 2.2505
R20930 DVDD.n11674 DVDD.n11630 2.2505
R20931 DVDD.n11677 DVDD.n11676 2.2505
R20932 DVDD.n11681 DVDD.n11680 2.2505
R20933 DVDD.n11684 DVDD.n11683 2.2505
R20934 DVDD.n11688 DVDD.n11687 2.2505
R20935 DVDD.n11685 DVDD.n11672 2.2505
R20936 DVDD.n11693 DVDD.n11692 2.2505
R20937 DVDD.n11696 DVDD.n11695 2.2505
R20938 DVDD.n11700 DVDD.n11699 2.2505
R20939 DVDD.n11697 DVDD.n11670 2.2505
R20940 DVDD.n11705 DVDD.n11704 2.2505
R20941 DVDD.n11708 DVDD.n11707 2.2505
R20942 DVDD.n11712 DVDD.n11711 2.2505
R20943 DVDD.n11709 DVDD.n11668 2.2505
R20944 DVDD.n11717 DVDD.n11716 2.2505
R20945 DVDD.n11720 DVDD.n11719 2.2505
R20946 DVDD.n11724 DVDD.n11723 2.2505
R20947 DVDD.n11721 DVDD.n11666 2.2505
R20948 DVDD.n11729 DVDD.n11728 2.2505
R20949 DVDD.n11732 DVDD.n11731 2.2505
R20950 DVDD.n11736 DVDD.n11735 2.2505
R20951 DVDD.n11733 DVDD.n11664 2.2505
R20952 DVDD.n11741 DVDD.n11740 2.2505
R20953 DVDD.n11744 DVDD.n11743 2.2505
R20954 DVDD.n11748 DVDD.n11747 2.2505
R20955 DVDD.n11745 DVDD.n11662 2.2505
R20956 DVDD.n11753 DVDD.n11752 2.2505
R20957 DVDD.n11756 DVDD.n11755 2.2505
R20958 DVDD.n11760 DVDD.n11759 2.2505
R20959 DVDD.n11757 DVDD.n11660 2.2505
R20960 DVDD.n11765 DVDD.n11764 2.2505
R20961 DVDD.n11768 DVDD.n11767 2.2505
R20962 DVDD.n11772 DVDD.n11771 2.2505
R20963 DVDD.n11769 DVDD.n11658 2.2505
R20964 DVDD.n11777 DVDD.n11776 2.2505
R20965 DVDD.n11780 DVDD.n11779 2.2505
R20966 DVDD.n11784 DVDD.n11783 2.2505
R20967 DVDD.n11781 DVDD.n11656 2.2505
R20968 DVDD.n11789 DVDD.n11788 2.2505
R20969 DVDD.n11792 DVDD.n11791 2.2505
R20970 DVDD.n11796 DVDD.n11795 2.2505
R20971 DVDD.n11793 DVDD.n11654 2.2505
R20972 DVDD.n11801 DVDD.n11800 2.2505
R20973 DVDD.n11804 DVDD.n11803 2.2505
R20974 DVDD.n11808 DVDD.n11807 2.2505
R20975 DVDD.n11805 DVDD.n11652 2.2505
R20976 DVDD.n11813 DVDD.n11812 2.2505
R20977 DVDD.n11816 DVDD.n11815 2.2505
R20978 DVDD.n11820 DVDD.n11819 2.2505
R20979 DVDD.n11817 DVDD.n11650 2.2505
R20980 DVDD.n11825 DVDD.n11824 2.2505
R20981 DVDD.n11828 DVDD.n11827 2.2505
R20982 DVDD.n11832 DVDD.n11831 2.2505
R20983 DVDD.n11829 DVDD.n11648 2.2505
R20984 DVDD.n11837 DVDD.n11836 2.2505
R20985 DVDD.n11840 DVDD.n11839 2.2505
R20986 DVDD.n11844 DVDD.n11843 2.2505
R20987 DVDD.n11841 DVDD.n11646 2.2505
R20988 DVDD.n11849 DVDD.n11848 2.2505
R20989 DVDD.n11852 DVDD.n11851 2.2505
R20990 DVDD.n11856 DVDD.n11855 2.2505
R20991 DVDD.n11853 DVDD.n11644 2.2505
R20992 DVDD.n11861 DVDD.n11860 2.2505
R20993 DVDD.n11864 DVDD.n11863 2.2505
R20994 DVDD.n11868 DVDD.n11867 2.2505
R20995 DVDD.n11865 DVDD.n11642 2.2505
R20996 DVDD.n11873 DVDD.n11872 2.2505
R20997 DVDD.n11876 DVDD.n11875 2.2505
R20998 DVDD.n11880 DVDD.n11879 2.2505
R20999 DVDD.n11877 DVDD.n11640 2.2505
R21000 DVDD.n11885 DVDD.n11884 2.2505
R21001 DVDD.n11888 DVDD.n11887 2.2505
R21002 DVDD.n11892 DVDD.n11891 2.2505
R21003 DVDD.n11889 DVDD.n11638 2.2505
R21004 DVDD.n11897 DVDD.n11896 2.2505
R21005 DVDD.n11900 DVDD.n11899 2.2505
R21006 DVDD.n11904 DVDD.n11903 2.2505
R21007 DVDD.n11901 DVDD.n11636 2.2505
R21008 DVDD.n11909 DVDD.n11908 2.2505
R21009 DVDD.n11912 DVDD.n11911 2.2505
R21010 DVDD.n11916 DVDD.n11915 2.2505
R21011 DVDD.n11913 DVDD.n11634 2.2505
R21012 DVDD.n13774 DVDD.n13773 2.2505
R21013 DVDD.n13776 DVDD.n11633 2.2505
R21014 DVDD.n12277 DVDD.n12276 2.2505
R21015 DVDD.n11945 DVDD.n11944 2.2505
R21016 DVDD.n12266 DVDD.n11946 2.2505
R21017 DVDD.n12268 DVDD.n12267 2.2505
R21018 DVDD.n12265 DVDD.n11948 2.2505
R21019 DVDD.n12264 DVDD.n12263 2.2505
R21020 DVDD.n11950 DVDD.n11949 2.2505
R21021 DVDD.n12255 DVDD.n12254 2.2505
R21022 DVDD.n12253 DVDD.n11952 2.2505
R21023 DVDD.n12252 DVDD.n12251 2.2505
R21024 DVDD.n11954 DVDD.n11953 2.2505
R21025 DVDD.n12243 DVDD.n12242 2.2505
R21026 DVDD.n12241 DVDD.n11956 2.2505
R21027 DVDD.n12240 DVDD.n12239 2.2505
R21028 DVDD.n11958 DVDD.n11957 2.2505
R21029 DVDD.n12231 DVDD.n12230 2.2505
R21030 DVDD.n12229 DVDD.n11960 2.2505
R21031 DVDD.n12228 DVDD.n12227 2.2505
R21032 DVDD.n11962 DVDD.n11961 2.2505
R21033 DVDD.n12219 DVDD.n12218 2.2505
R21034 DVDD.n12217 DVDD.n11964 2.2505
R21035 DVDD.n12216 DVDD.n12215 2.2505
R21036 DVDD.n11966 DVDD.n11965 2.2505
R21037 DVDD.n12207 DVDD.n12206 2.2505
R21038 DVDD.n12205 DVDD.n11968 2.2505
R21039 DVDD.n12204 DVDD.n12203 2.2505
R21040 DVDD.n11970 DVDD.n11969 2.2505
R21041 DVDD.n12195 DVDD.n12194 2.2505
R21042 DVDD.n12193 DVDD.n11972 2.2505
R21043 DVDD.n12192 DVDD.n12191 2.2505
R21044 DVDD.n11974 DVDD.n11973 2.2505
R21045 DVDD.n12183 DVDD.n12182 2.2505
R21046 DVDD.n12181 DVDD.n11976 2.2505
R21047 DVDD.n12180 DVDD.n12179 2.2505
R21048 DVDD.n11978 DVDD.n11977 2.2505
R21049 DVDD.n12171 DVDD.n12170 2.2505
R21050 DVDD.n12169 DVDD.n11980 2.2505
R21051 DVDD.n12168 DVDD.n12167 2.2505
R21052 DVDD.n11982 DVDD.n11981 2.2505
R21053 DVDD.n12159 DVDD.n12158 2.2505
R21054 DVDD.n12157 DVDD.n11984 2.2505
R21055 DVDD.n12156 DVDD.n12155 2.2505
R21056 DVDD.n11986 DVDD.n11985 2.2505
R21057 DVDD.n12147 DVDD.n12146 2.2505
R21058 DVDD.n12145 DVDD.n11988 2.2505
R21059 DVDD.n12144 DVDD.n12143 2.2505
R21060 DVDD.n11990 DVDD.n11989 2.2505
R21061 DVDD.n12135 DVDD.n12134 2.2505
R21062 DVDD.n12133 DVDD.n11992 2.2505
R21063 DVDD.n12132 DVDD.n12131 2.2505
R21064 DVDD.n11994 DVDD.n11993 2.2505
R21065 DVDD.n12123 DVDD.n12122 2.2505
R21066 DVDD.n12121 DVDD.n11996 2.2505
R21067 DVDD.n12120 DVDD.n12119 2.2505
R21068 DVDD.n11998 DVDD.n11997 2.2505
R21069 DVDD.n12111 DVDD.n12110 2.2505
R21070 DVDD.n12109 DVDD.n12000 2.2505
R21071 DVDD.n12108 DVDD.n12107 2.2505
R21072 DVDD.n12002 DVDD.n12001 2.2505
R21073 DVDD.n12099 DVDD.n12098 2.2505
R21074 DVDD.n12097 DVDD.n12004 2.2505
R21075 DVDD.n12096 DVDD.n12095 2.2505
R21076 DVDD.n12006 DVDD.n12005 2.2505
R21077 DVDD.n12087 DVDD.n12086 2.2505
R21078 DVDD.n12085 DVDD.n12008 2.2505
R21079 DVDD.n12084 DVDD.n12083 2.2505
R21080 DVDD.n12010 DVDD.n12009 2.2505
R21081 DVDD.n12075 DVDD.n12074 2.2505
R21082 DVDD.n12073 DVDD.n12012 2.2505
R21083 DVDD.n12072 DVDD.n12071 2.2505
R21084 DVDD.n12014 DVDD.n12013 2.2505
R21085 DVDD.n12063 DVDD.n12062 2.2505
R21086 DVDD.n12061 DVDD.n12016 2.2505
R21087 DVDD.n12060 DVDD.n12059 2.2505
R21088 DVDD.n12018 DVDD.n12017 2.2505
R21089 DVDD.n12051 DVDD.n12050 2.2505
R21090 DVDD.n12049 DVDD.n12020 2.2505
R21091 DVDD.n12048 DVDD.n12047 2.2505
R21092 DVDD.n12022 DVDD.n12021 2.2505
R21093 DVDD.n12039 DVDD.n12038 2.2505
R21094 DVDD.n12037 DVDD.n12024 2.2505
R21095 DVDD.n12036 DVDD.n12035 2.2505
R21096 DVDD.n12026 DVDD.n12025 2.2505
R21097 DVDD.n12027 DVDD.n11930 2.2505
R21098 DVDD.n12028 DVDD.n12027 2.2505
R21099 DVDD.n12030 DVDD.n12026 2.2505
R21100 DVDD.n12035 DVDD.n12034 2.2505
R21101 DVDD.n12032 DVDD.n12024 2.2505
R21102 DVDD.n12040 DVDD.n12039 2.2505
R21103 DVDD.n12042 DVDD.n12022 2.2505
R21104 DVDD.n12047 DVDD.n12046 2.2505
R21105 DVDD.n12044 DVDD.n12020 2.2505
R21106 DVDD.n12052 DVDD.n12051 2.2505
R21107 DVDD.n12054 DVDD.n12018 2.2505
R21108 DVDD.n12059 DVDD.n12058 2.2505
R21109 DVDD.n12056 DVDD.n12016 2.2505
R21110 DVDD.n12064 DVDD.n12063 2.2505
R21111 DVDD.n12066 DVDD.n12014 2.2505
R21112 DVDD.n12071 DVDD.n12070 2.2505
R21113 DVDD.n12068 DVDD.n12012 2.2505
R21114 DVDD.n12076 DVDD.n12075 2.2505
R21115 DVDD.n12078 DVDD.n12010 2.2505
R21116 DVDD.n12083 DVDD.n12082 2.2505
R21117 DVDD.n12080 DVDD.n12008 2.2505
R21118 DVDD.n12088 DVDD.n12087 2.2505
R21119 DVDD.n12090 DVDD.n12006 2.2505
R21120 DVDD.n12095 DVDD.n12094 2.2505
R21121 DVDD.n12092 DVDD.n12004 2.2505
R21122 DVDD.n12100 DVDD.n12099 2.2505
R21123 DVDD.n12102 DVDD.n12002 2.2505
R21124 DVDD.n12107 DVDD.n12106 2.2505
R21125 DVDD.n12104 DVDD.n12000 2.2505
R21126 DVDD.n12112 DVDD.n12111 2.2505
R21127 DVDD.n12114 DVDD.n11998 2.2505
R21128 DVDD.n12119 DVDD.n12118 2.2505
R21129 DVDD.n12116 DVDD.n11996 2.2505
R21130 DVDD.n12124 DVDD.n12123 2.2505
R21131 DVDD.n12126 DVDD.n11994 2.2505
R21132 DVDD.n12131 DVDD.n12130 2.2505
R21133 DVDD.n12128 DVDD.n11992 2.2505
R21134 DVDD.n12136 DVDD.n12135 2.2505
R21135 DVDD.n12138 DVDD.n11990 2.2505
R21136 DVDD.n12143 DVDD.n12142 2.2505
R21137 DVDD.n12140 DVDD.n11988 2.2505
R21138 DVDD.n12148 DVDD.n12147 2.2505
R21139 DVDD.n12150 DVDD.n11986 2.2505
R21140 DVDD.n12155 DVDD.n12154 2.2505
R21141 DVDD.n12152 DVDD.n11984 2.2505
R21142 DVDD.n12160 DVDD.n12159 2.2505
R21143 DVDD.n12162 DVDD.n11982 2.2505
R21144 DVDD.n12167 DVDD.n12166 2.2505
R21145 DVDD.n12164 DVDD.n11980 2.2505
R21146 DVDD.n12172 DVDD.n12171 2.2505
R21147 DVDD.n12174 DVDD.n11978 2.2505
R21148 DVDD.n12179 DVDD.n12178 2.2505
R21149 DVDD.n12176 DVDD.n11976 2.2505
R21150 DVDD.n12184 DVDD.n12183 2.2505
R21151 DVDD.n12186 DVDD.n11974 2.2505
R21152 DVDD.n12191 DVDD.n12190 2.2505
R21153 DVDD.n12188 DVDD.n11972 2.2505
R21154 DVDD.n12196 DVDD.n12195 2.2505
R21155 DVDD.n12198 DVDD.n11970 2.2505
R21156 DVDD.n12203 DVDD.n12202 2.2505
R21157 DVDD.n12200 DVDD.n11968 2.2505
R21158 DVDD.n12208 DVDD.n12207 2.2505
R21159 DVDD.n12210 DVDD.n11966 2.2505
R21160 DVDD.n12215 DVDD.n12214 2.2505
R21161 DVDD.n12212 DVDD.n11964 2.2505
R21162 DVDD.n12220 DVDD.n12219 2.2505
R21163 DVDD.n12222 DVDD.n11962 2.2505
R21164 DVDD.n12227 DVDD.n12226 2.2505
R21165 DVDD.n12224 DVDD.n11960 2.2505
R21166 DVDD.n12232 DVDD.n12231 2.2505
R21167 DVDD.n12234 DVDD.n11958 2.2505
R21168 DVDD.n12239 DVDD.n12238 2.2505
R21169 DVDD.n12236 DVDD.n11956 2.2505
R21170 DVDD.n12244 DVDD.n12243 2.2505
R21171 DVDD.n12246 DVDD.n11954 2.2505
R21172 DVDD.n12251 DVDD.n12250 2.2505
R21173 DVDD.n12248 DVDD.n11952 2.2505
R21174 DVDD.n12256 DVDD.n12255 2.2505
R21175 DVDD.n12258 DVDD.n11950 2.2505
R21176 DVDD.n12263 DVDD.n12262 2.2505
R21177 DVDD.n12260 DVDD.n11948 2.2505
R21178 DVDD.n12269 DVDD.n12268 2.2505
R21179 DVDD.n12271 DVDD.n11946 2.2505
R21180 DVDD.n12273 DVDD.n11945 2.2505
R21181 DVDD.n12276 DVDD.n12275 2.2505
R21182 DVDD.n12331 DVDD.n12281 2.2505
R21183 DVDD.n13740 DVDD.n13739 2.2505
R21184 DVDD.n13738 DVDD.n12334 2.2505
R21185 DVDD.n13737 DVDD.n13736 2.2505
R21186 DVDD.n13732 DVDD.n12335 2.2505
R21187 DVDD.n13728 DVDD.n13727 2.2505
R21188 DVDD.n13726 DVDD.n12336 2.2505
R21189 DVDD.n13725 DVDD.n13724 2.2505
R21190 DVDD.n13720 DVDD.n12337 2.2505
R21191 DVDD.n13716 DVDD.n13715 2.2505
R21192 DVDD.n13714 DVDD.n12338 2.2505
R21193 DVDD.n13713 DVDD.n13712 2.2505
R21194 DVDD.n13708 DVDD.n12339 2.2505
R21195 DVDD.n13704 DVDD.n13703 2.2505
R21196 DVDD.n13702 DVDD.n12340 2.2505
R21197 DVDD.n13701 DVDD.n13700 2.2505
R21198 DVDD.n13696 DVDD.n12341 2.2505
R21199 DVDD.n13692 DVDD.n13691 2.2505
R21200 DVDD.n13690 DVDD.n12342 2.2505
R21201 DVDD.n13689 DVDD.n13688 2.2505
R21202 DVDD.n13684 DVDD.n12343 2.2505
R21203 DVDD.n13680 DVDD.n13679 2.2505
R21204 DVDD.n13678 DVDD.n12344 2.2505
R21205 DVDD.n13677 DVDD.n13676 2.2505
R21206 DVDD.n13672 DVDD.n12345 2.2505
R21207 DVDD.n13668 DVDD.n13667 2.2505
R21208 DVDD.n13666 DVDD.n12346 2.2505
R21209 DVDD.n13665 DVDD.n13664 2.2505
R21210 DVDD.n13660 DVDD.n12347 2.2505
R21211 DVDD.n13656 DVDD.n13655 2.2505
R21212 DVDD.n13654 DVDD.n12348 2.2505
R21213 DVDD.n13653 DVDD.n13652 2.2505
R21214 DVDD.n13648 DVDD.n12349 2.2505
R21215 DVDD.n13644 DVDD.n13643 2.2505
R21216 DVDD.n13642 DVDD.n12350 2.2505
R21217 DVDD.n13641 DVDD.n13640 2.2505
R21218 DVDD.n13636 DVDD.n12351 2.2505
R21219 DVDD.n13632 DVDD.n13631 2.2505
R21220 DVDD.n13630 DVDD.n12352 2.2505
R21221 DVDD.n13629 DVDD.n13628 2.2505
R21222 DVDD.n13624 DVDD.n12353 2.2505
R21223 DVDD.n13620 DVDD.n13619 2.2505
R21224 DVDD.n13618 DVDD.n12354 2.2505
R21225 DVDD.n13617 DVDD.n13616 2.2505
R21226 DVDD.n13612 DVDD.n12355 2.2505
R21227 DVDD.n13608 DVDD.n13607 2.2505
R21228 DVDD.n13606 DVDD.n12356 2.2505
R21229 DVDD.n13605 DVDD.n13604 2.2505
R21230 DVDD.n13600 DVDD.n12357 2.2505
R21231 DVDD.n13596 DVDD.n13595 2.2505
R21232 DVDD.n13594 DVDD.n12358 2.2505
R21233 DVDD.n13593 DVDD.n13592 2.2505
R21234 DVDD.n13588 DVDD.n12359 2.2505
R21235 DVDD.n13584 DVDD.n13583 2.2505
R21236 DVDD.n13582 DVDD.n12360 2.2505
R21237 DVDD.n13581 DVDD.n13580 2.2505
R21238 DVDD.n13576 DVDD.n12361 2.2505
R21239 DVDD.n13572 DVDD.n13571 2.2505
R21240 DVDD.n13570 DVDD.n12362 2.2505
R21241 DVDD.n13569 DVDD.n13568 2.2505
R21242 DVDD.n13564 DVDD.n12363 2.2505
R21243 DVDD.n13560 DVDD.n13559 2.2505
R21244 DVDD.n13558 DVDD.n12364 2.2505
R21245 DVDD.n13557 DVDD.n13556 2.2505
R21246 DVDD.n13552 DVDD.n12365 2.2505
R21247 DVDD.n13548 DVDD.n13547 2.2505
R21248 DVDD.n13546 DVDD.n12366 2.2505
R21249 DVDD.n13545 DVDD.n13544 2.2505
R21250 DVDD.n13540 DVDD.n12367 2.2505
R21251 DVDD.n13536 DVDD.n13535 2.2505
R21252 DVDD.n13534 DVDD.n12368 2.2505
R21253 DVDD.n13533 DVDD.n13532 2.2505
R21254 DVDD.n13528 DVDD.n12369 2.2505
R21255 DVDD.n13524 DVDD.n13523 2.2505
R21256 DVDD.n13522 DVDD.n12370 2.2505
R21257 DVDD.n13521 DVDD.n13520 2.2505
R21258 DVDD.n13516 DVDD.n12371 2.2505
R21259 DVDD.n13512 DVDD.n13511 2.2505
R21260 DVDD.n13510 DVDD.n12372 2.2505
R21261 DVDD.n13509 DVDD.n13508 2.2505
R21262 DVDD.n13504 DVDD.n12373 2.2505
R21263 DVDD.n13500 DVDD.n13499 2.2505
R21264 DVDD.n13498 DVDD.n12376 2.2505
R21265 DVDD.n13497 DVDD.n13496 2.2505
R21266 DVDD.n13496 DVDD.n12329 2.2505
R21267 DVDD.n12376 DVDD.n12375 2.2505
R21268 DVDD.n13501 DVDD.n13500 2.2505
R21269 DVDD.n13504 DVDD.n13503 2.2505
R21270 DVDD.n13508 DVDD.n13507 2.2505
R21271 DVDD.n13505 DVDD.n12372 2.2505
R21272 DVDD.n13513 DVDD.n13512 2.2505
R21273 DVDD.n13516 DVDD.n13515 2.2505
R21274 DVDD.n13520 DVDD.n13519 2.2505
R21275 DVDD.n13517 DVDD.n12370 2.2505
R21276 DVDD.n13525 DVDD.n13524 2.2505
R21277 DVDD.n13528 DVDD.n13527 2.2505
R21278 DVDD.n13532 DVDD.n13531 2.2505
R21279 DVDD.n13529 DVDD.n12368 2.2505
R21280 DVDD.n13537 DVDD.n13536 2.2505
R21281 DVDD.n13540 DVDD.n13539 2.2505
R21282 DVDD.n13544 DVDD.n13543 2.2505
R21283 DVDD.n13541 DVDD.n12366 2.2505
R21284 DVDD.n13549 DVDD.n13548 2.2505
R21285 DVDD.n13552 DVDD.n13551 2.2505
R21286 DVDD.n13556 DVDD.n13555 2.2505
R21287 DVDD.n13553 DVDD.n12364 2.2505
R21288 DVDD.n13561 DVDD.n13560 2.2505
R21289 DVDD.n13564 DVDD.n13563 2.2505
R21290 DVDD.n13568 DVDD.n13567 2.2505
R21291 DVDD.n13565 DVDD.n12362 2.2505
R21292 DVDD.n13573 DVDD.n13572 2.2505
R21293 DVDD.n13576 DVDD.n13575 2.2505
R21294 DVDD.n13580 DVDD.n13579 2.2505
R21295 DVDD.n13577 DVDD.n12360 2.2505
R21296 DVDD.n13585 DVDD.n13584 2.2505
R21297 DVDD.n13588 DVDD.n13587 2.2505
R21298 DVDD.n13592 DVDD.n13591 2.2505
R21299 DVDD.n13589 DVDD.n12358 2.2505
R21300 DVDD.n13597 DVDD.n13596 2.2505
R21301 DVDD.n13600 DVDD.n13599 2.2505
R21302 DVDD.n13604 DVDD.n13603 2.2505
R21303 DVDD.n13601 DVDD.n12356 2.2505
R21304 DVDD.n13609 DVDD.n13608 2.2505
R21305 DVDD.n13612 DVDD.n13611 2.2505
R21306 DVDD.n13616 DVDD.n13615 2.2505
R21307 DVDD.n13613 DVDD.n12354 2.2505
R21308 DVDD.n13621 DVDD.n13620 2.2505
R21309 DVDD.n13624 DVDD.n13623 2.2505
R21310 DVDD.n13628 DVDD.n13627 2.2505
R21311 DVDD.n13625 DVDD.n12352 2.2505
R21312 DVDD.n13633 DVDD.n13632 2.2505
R21313 DVDD.n13636 DVDD.n13635 2.2505
R21314 DVDD.n13640 DVDD.n13639 2.2505
R21315 DVDD.n13637 DVDD.n12350 2.2505
R21316 DVDD.n13645 DVDD.n13644 2.2505
R21317 DVDD.n13648 DVDD.n13647 2.2505
R21318 DVDD.n13652 DVDD.n13651 2.2505
R21319 DVDD.n13649 DVDD.n12348 2.2505
R21320 DVDD.n13657 DVDD.n13656 2.2505
R21321 DVDD.n13660 DVDD.n13659 2.2505
R21322 DVDD.n13664 DVDD.n13663 2.2505
R21323 DVDD.n13661 DVDD.n12346 2.2505
R21324 DVDD.n13669 DVDD.n13668 2.2505
R21325 DVDD.n13672 DVDD.n13671 2.2505
R21326 DVDD.n13676 DVDD.n13675 2.2505
R21327 DVDD.n13673 DVDD.n12344 2.2505
R21328 DVDD.n13681 DVDD.n13680 2.2505
R21329 DVDD.n13684 DVDD.n13683 2.2505
R21330 DVDD.n13688 DVDD.n13687 2.2505
R21331 DVDD.n13685 DVDD.n12342 2.2505
R21332 DVDD.n13693 DVDD.n13692 2.2505
R21333 DVDD.n13696 DVDD.n13695 2.2505
R21334 DVDD.n13700 DVDD.n13699 2.2505
R21335 DVDD.n13697 DVDD.n12340 2.2505
R21336 DVDD.n13705 DVDD.n13704 2.2505
R21337 DVDD.n13708 DVDD.n13707 2.2505
R21338 DVDD.n13712 DVDD.n13711 2.2505
R21339 DVDD.n13709 DVDD.n12338 2.2505
R21340 DVDD.n13717 DVDD.n13716 2.2505
R21341 DVDD.n13720 DVDD.n13719 2.2505
R21342 DVDD.n13724 DVDD.n13723 2.2505
R21343 DVDD.n13721 DVDD.n12336 2.2505
R21344 DVDD.n13729 DVDD.n13728 2.2505
R21345 DVDD.n13732 DVDD.n13731 2.2505
R21346 DVDD.n13736 DVDD.n13735 2.2505
R21347 DVDD.n13733 DVDD.n12334 2.2505
R21348 DVDD.n13741 DVDD.n13740 2.2505
R21349 DVDD.n13743 DVDD.n12331 2.2505
R21350 DVDD.n13482 DVDD.n12725 2.2505
R21351 DVDD.n12724 DVDD.n12480 2.2505
R21352 DVDD.n12723 DVDD.n12722 2.2505
R21353 DVDD.n12720 DVDD.n12481 2.2505
R21354 DVDD.n12718 DVDD.n12716 2.2505
R21355 DVDD.n12715 DVDD.n12483 2.2505
R21356 DVDD.n12714 DVDD.n12713 2.2505
R21357 DVDD.n12711 DVDD.n12484 2.2505
R21358 DVDD.n12709 DVDD.n12707 2.2505
R21359 DVDD.n12706 DVDD.n12486 2.2505
R21360 DVDD.n12705 DVDD.n12704 2.2505
R21361 DVDD.n12702 DVDD.n12487 2.2505
R21362 DVDD.n12700 DVDD.n12698 2.2505
R21363 DVDD.n12697 DVDD.n12489 2.2505
R21364 DVDD.n12696 DVDD.n12695 2.2505
R21365 DVDD.n12693 DVDD.n12490 2.2505
R21366 DVDD.n12691 DVDD.n12689 2.2505
R21367 DVDD.n12688 DVDD.n12492 2.2505
R21368 DVDD.n12687 DVDD.n12686 2.2505
R21369 DVDD.n12684 DVDD.n12493 2.2505
R21370 DVDD.n12682 DVDD.n12680 2.2505
R21371 DVDD.n12679 DVDD.n12495 2.2505
R21372 DVDD.n12678 DVDD.n12677 2.2505
R21373 DVDD.n12675 DVDD.n12496 2.2505
R21374 DVDD.n12673 DVDD.n12671 2.2505
R21375 DVDD.n12670 DVDD.n12498 2.2505
R21376 DVDD.n12669 DVDD.n12668 2.2505
R21377 DVDD.n12666 DVDD.n12499 2.2505
R21378 DVDD.n12664 DVDD.n12662 2.2505
R21379 DVDD.n12661 DVDD.n12501 2.2505
R21380 DVDD.n12660 DVDD.n12659 2.2505
R21381 DVDD.n12657 DVDD.n12502 2.2505
R21382 DVDD.n12655 DVDD.n12653 2.2505
R21383 DVDD.n12652 DVDD.n12504 2.2505
R21384 DVDD.n12651 DVDD.n12650 2.2505
R21385 DVDD.n12648 DVDD.n12505 2.2505
R21386 DVDD.n12646 DVDD.n12644 2.2505
R21387 DVDD.n12643 DVDD.n12507 2.2505
R21388 DVDD.n12642 DVDD.n12641 2.2505
R21389 DVDD.n12639 DVDD.n12508 2.2505
R21390 DVDD.n12637 DVDD.n12635 2.2505
R21391 DVDD.n12634 DVDD.n12510 2.2505
R21392 DVDD.n12633 DVDD.n12632 2.2505
R21393 DVDD.n12630 DVDD.n12511 2.2505
R21394 DVDD.n12628 DVDD.n12626 2.2505
R21395 DVDD.n12625 DVDD.n12513 2.2505
R21396 DVDD.n12624 DVDD.n12623 2.2505
R21397 DVDD.n12621 DVDD.n12514 2.2505
R21398 DVDD.n12619 DVDD.n12617 2.2505
R21399 DVDD.n12616 DVDD.n12516 2.2505
R21400 DVDD.n12615 DVDD.n12614 2.2505
R21401 DVDD.n12612 DVDD.n12517 2.2505
R21402 DVDD.n12610 DVDD.n12608 2.2505
R21403 DVDD.n12607 DVDD.n12519 2.2505
R21404 DVDD.n12606 DVDD.n12605 2.2505
R21405 DVDD.n12603 DVDD.n12520 2.2505
R21406 DVDD.n12601 DVDD.n12599 2.2505
R21407 DVDD.n12598 DVDD.n12522 2.2505
R21408 DVDD.n12597 DVDD.n12596 2.2505
R21409 DVDD.n12594 DVDD.n12523 2.2505
R21410 DVDD.n12592 DVDD.n12590 2.2505
R21411 DVDD.n12589 DVDD.n12525 2.2505
R21412 DVDD.n12588 DVDD.n12587 2.2505
R21413 DVDD.n12585 DVDD.n12526 2.2505
R21414 DVDD.n12583 DVDD.n12581 2.2505
R21415 DVDD.n12580 DVDD.n12528 2.2505
R21416 DVDD.n12579 DVDD.n12578 2.2505
R21417 DVDD.n12576 DVDD.n12529 2.2505
R21418 DVDD.n12574 DVDD.n12572 2.2505
R21419 DVDD.n12571 DVDD.n12531 2.2505
R21420 DVDD.n12570 DVDD.n12569 2.2505
R21421 DVDD.n12567 DVDD.n12532 2.2505
R21422 DVDD.n12565 DVDD.n12563 2.2505
R21423 DVDD.n12562 DVDD.n12534 2.2505
R21424 DVDD.n12561 DVDD.n12560 2.2505
R21425 DVDD.n12558 DVDD.n12535 2.2505
R21426 DVDD.n12556 DVDD.n12554 2.2505
R21427 DVDD.n12553 DVDD.n12537 2.2505
R21428 DVDD.n12552 DVDD.n12551 2.2505
R21429 DVDD.n12549 DVDD.n12538 2.2505
R21430 DVDD.n12547 DVDD.n12545 2.2505
R21431 DVDD.n12544 DVDD.n12540 2.2505
R21432 DVDD.n12543 DVDD.n12542 2.2505
R21433 DVDD.n12541 DVDD.n12434 2.2505
R21434 DVDD.n13485 DVDD.n12434 2.2505
R21435 DVDD.n12542 DVDD.n12433 2.2505
R21436 DVDD.n12540 DVDD.n12539 2.2505
R21437 DVDD.n12547 DVDD.n12546 2.2505
R21438 DVDD.n12549 DVDD.n12548 2.2505
R21439 DVDD.n12551 DVDD.n12550 2.2505
R21440 DVDD.n12537 DVDD.n12536 2.2505
R21441 DVDD.n12556 DVDD.n12555 2.2505
R21442 DVDD.n12558 DVDD.n12557 2.2505
R21443 DVDD.n12560 DVDD.n12559 2.2505
R21444 DVDD.n12534 DVDD.n12533 2.2505
R21445 DVDD.n12565 DVDD.n12564 2.2505
R21446 DVDD.n12567 DVDD.n12566 2.2505
R21447 DVDD.n12569 DVDD.n12568 2.2505
R21448 DVDD.n12531 DVDD.n12530 2.2505
R21449 DVDD.n12574 DVDD.n12573 2.2505
R21450 DVDD.n12576 DVDD.n12575 2.2505
R21451 DVDD.n12578 DVDD.n12577 2.2505
R21452 DVDD.n12528 DVDD.n12527 2.2505
R21453 DVDD.n12583 DVDD.n12582 2.2505
R21454 DVDD.n12585 DVDD.n12584 2.2505
R21455 DVDD.n12587 DVDD.n12586 2.2505
R21456 DVDD.n12525 DVDD.n12524 2.2505
R21457 DVDD.n12592 DVDD.n12591 2.2505
R21458 DVDD.n12594 DVDD.n12593 2.2505
R21459 DVDD.n12596 DVDD.n12595 2.2505
R21460 DVDD.n12522 DVDD.n12521 2.2505
R21461 DVDD.n12601 DVDD.n12600 2.2505
R21462 DVDD.n12603 DVDD.n12602 2.2505
R21463 DVDD.n12605 DVDD.n12604 2.2505
R21464 DVDD.n12519 DVDD.n12518 2.2505
R21465 DVDD.n12610 DVDD.n12609 2.2505
R21466 DVDD.n12612 DVDD.n12611 2.2505
R21467 DVDD.n12614 DVDD.n12613 2.2505
R21468 DVDD.n12516 DVDD.n12515 2.2505
R21469 DVDD.n12619 DVDD.n12618 2.2505
R21470 DVDD.n12621 DVDD.n12620 2.2505
R21471 DVDD.n12623 DVDD.n12622 2.2505
R21472 DVDD.n12513 DVDD.n12512 2.2505
R21473 DVDD.n12628 DVDD.n12627 2.2505
R21474 DVDD.n12630 DVDD.n12629 2.2505
R21475 DVDD.n12632 DVDD.n12631 2.2505
R21476 DVDD.n12510 DVDD.n12509 2.2505
R21477 DVDD.n12637 DVDD.n12636 2.2505
R21478 DVDD.n12639 DVDD.n12638 2.2505
R21479 DVDD.n12641 DVDD.n12640 2.2505
R21480 DVDD.n12507 DVDD.n12506 2.2505
R21481 DVDD.n12646 DVDD.n12645 2.2505
R21482 DVDD.n12648 DVDD.n12647 2.2505
R21483 DVDD.n12650 DVDD.n12649 2.2505
R21484 DVDD.n12504 DVDD.n12503 2.2505
R21485 DVDD.n12655 DVDD.n12654 2.2505
R21486 DVDD.n12657 DVDD.n12656 2.2505
R21487 DVDD.n12659 DVDD.n12658 2.2505
R21488 DVDD.n12501 DVDD.n12500 2.2505
R21489 DVDD.n12664 DVDD.n12663 2.2505
R21490 DVDD.n12666 DVDD.n12665 2.2505
R21491 DVDD.n12668 DVDD.n12667 2.2505
R21492 DVDD.n12498 DVDD.n12497 2.2505
R21493 DVDD.n12673 DVDD.n12672 2.2505
R21494 DVDD.n12675 DVDD.n12674 2.2505
R21495 DVDD.n12677 DVDD.n12676 2.2505
R21496 DVDD.n12495 DVDD.n12494 2.2505
R21497 DVDD.n12682 DVDD.n12681 2.2505
R21498 DVDD.n12684 DVDD.n12683 2.2505
R21499 DVDD.n12686 DVDD.n12685 2.2505
R21500 DVDD.n12492 DVDD.n12491 2.2505
R21501 DVDD.n12691 DVDD.n12690 2.2505
R21502 DVDD.n12693 DVDD.n12692 2.2505
R21503 DVDD.n12695 DVDD.n12694 2.2505
R21504 DVDD.n12489 DVDD.n12488 2.2505
R21505 DVDD.n12700 DVDD.n12699 2.2505
R21506 DVDD.n12702 DVDD.n12701 2.2505
R21507 DVDD.n12704 DVDD.n12703 2.2505
R21508 DVDD.n12486 DVDD.n12485 2.2505
R21509 DVDD.n12709 DVDD.n12708 2.2505
R21510 DVDD.n12711 DVDD.n12710 2.2505
R21511 DVDD.n12713 DVDD.n12712 2.2505
R21512 DVDD.n12483 DVDD.n12482 2.2505
R21513 DVDD.n12718 DVDD.n12717 2.2505
R21514 DVDD.n12720 DVDD.n12719 2.2505
R21515 DVDD.n12722 DVDD.n12721 2.2505
R21516 DVDD.n12480 DVDD.n12479 2.2505
R21517 DVDD.n13483 DVDD.n13482 2.2505
R21518 DVDD.n13468 DVDD.n13467 2.2505
R21519 DVDD.n13466 DVDD.n12827 2.2505
R21520 DVDD.n13465 DVDD.n13464 2.2505
R21521 DVDD.n13462 DVDD.n12828 2.2505
R21522 DVDD.n13460 DVDD.n13458 2.2505
R21523 DVDD.n13457 DVDD.n12830 2.2505
R21524 DVDD.n13456 DVDD.n13455 2.2505
R21525 DVDD.n13453 DVDD.n12831 2.2505
R21526 DVDD.n13451 DVDD.n13449 2.2505
R21527 DVDD.n13448 DVDD.n12833 2.2505
R21528 DVDD.n13447 DVDD.n13446 2.2505
R21529 DVDD.n13444 DVDD.n12834 2.2505
R21530 DVDD.n13442 DVDD.n13440 2.2505
R21531 DVDD.n13439 DVDD.n12836 2.2505
R21532 DVDD.n13438 DVDD.n13437 2.2505
R21533 DVDD.n13435 DVDD.n12837 2.2505
R21534 DVDD.n13433 DVDD.n13431 2.2505
R21535 DVDD.n13430 DVDD.n12839 2.2505
R21536 DVDD.n13429 DVDD.n13428 2.2505
R21537 DVDD.n13426 DVDD.n12840 2.2505
R21538 DVDD.n13424 DVDD.n13422 2.2505
R21539 DVDD.n13421 DVDD.n12842 2.2505
R21540 DVDD.n13420 DVDD.n13419 2.2505
R21541 DVDD.n13417 DVDD.n12843 2.2505
R21542 DVDD.n13415 DVDD.n13413 2.2505
R21543 DVDD.n13412 DVDD.n12845 2.2505
R21544 DVDD.n13411 DVDD.n13410 2.2505
R21545 DVDD.n13408 DVDD.n12846 2.2505
R21546 DVDD.n13406 DVDD.n13404 2.2505
R21547 DVDD.n13403 DVDD.n12848 2.2505
R21548 DVDD.n13402 DVDD.n13401 2.2505
R21549 DVDD.n13399 DVDD.n12849 2.2505
R21550 DVDD.n13397 DVDD.n13395 2.2505
R21551 DVDD.n13394 DVDD.n12851 2.2505
R21552 DVDD.n13393 DVDD.n13392 2.2505
R21553 DVDD.n13390 DVDD.n12852 2.2505
R21554 DVDD.n13388 DVDD.n13386 2.2505
R21555 DVDD.n13385 DVDD.n12854 2.2505
R21556 DVDD.n13384 DVDD.n13383 2.2505
R21557 DVDD.n13381 DVDD.n12855 2.2505
R21558 DVDD.n13379 DVDD.n13377 2.2505
R21559 DVDD.n13376 DVDD.n12857 2.2505
R21560 DVDD.n13375 DVDD.n13374 2.2505
R21561 DVDD.n13372 DVDD.n12858 2.2505
R21562 DVDD.n13370 DVDD.n13368 2.2505
R21563 DVDD.n13367 DVDD.n12860 2.2505
R21564 DVDD.n13366 DVDD.n13365 2.2505
R21565 DVDD.n13363 DVDD.n12861 2.2505
R21566 DVDD.n13361 DVDD.n13359 2.2505
R21567 DVDD.n13358 DVDD.n12863 2.2505
R21568 DVDD.n13357 DVDD.n13356 2.2505
R21569 DVDD.n13354 DVDD.n12864 2.2505
R21570 DVDD.n13352 DVDD.n13350 2.2505
R21571 DVDD.n13349 DVDD.n12866 2.2505
R21572 DVDD.n13348 DVDD.n13347 2.2505
R21573 DVDD.n13345 DVDD.n12867 2.2505
R21574 DVDD.n13343 DVDD.n13341 2.2505
R21575 DVDD.n13340 DVDD.n12869 2.2505
R21576 DVDD.n13339 DVDD.n13338 2.2505
R21577 DVDD.n13336 DVDD.n12870 2.2505
R21578 DVDD.n13334 DVDD.n13332 2.2505
R21579 DVDD.n13331 DVDD.n12872 2.2505
R21580 DVDD.n13330 DVDD.n13329 2.2505
R21581 DVDD.n13327 DVDD.n12873 2.2505
R21582 DVDD.n13325 DVDD.n13323 2.2505
R21583 DVDD.n13322 DVDD.n12875 2.2505
R21584 DVDD.n13321 DVDD.n13320 2.2505
R21585 DVDD.n13318 DVDD.n12876 2.2505
R21586 DVDD.n13316 DVDD.n13314 2.2505
R21587 DVDD.n13313 DVDD.n12878 2.2505
R21588 DVDD.n13312 DVDD.n13311 2.2505
R21589 DVDD.n13309 DVDD.n12879 2.2505
R21590 DVDD.n13307 DVDD.n13305 2.2505
R21591 DVDD.n13304 DVDD.n12881 2.2505
R21592 DVDD.n13303 DVDD.n13302 2.2505
R21593 DVDD.n13300 DVDD.n12882 2.2505
R21594 DVDD.n13298 DVDD.n13296 2.2505
R21595 DVDD.n13295 DVDD.n12884 2.2505
R21596 DVDD.n13294 DVDD.n13293 2.2505
R21597 DVDD.n13291 DVDD.n12885 2.2505
R21598 DVDD.n13289 DVDD.n13287 2.2505
R21599 DVDD.n13286 DVDD.n12887 2.2505
R21600 DVDD.n13285 DVDD.n13284 2.2505
R21601 DVDD.n13283 DVDD.n12782 2.2505
R21602 DVDD.n13471 DVDD.n12782 2.2505
R21603 DVDD.n13284 DVDD.n12780 2.2505
R21604 DVDD.n12887 DVDD.n12886 2.2505
R21605 DVDD.n13289 DVDD.n13288 2.2505
R21606 DVDD.n13291 DVDD.n13290 2.2505
R21607 DVDD.n13293 DVDD.n13292 2.2505
R21608 DVDD.n12884 DVDD.n12883 2.2505
R21609 DVDD.n13298 DVDD.n13297 2.2505
R21610 DVDD.n13300 DVDD.n13299 2.2505
R21611 DVDD.n13302 DVDD.n13301 2.2505
R21612 DVDD.n12881 DVDD.n12880 2.2505
R21613 DVDD.n13307 DVDD.n13306 2.2505
R21614 DVDD.n13309 DVDD.n13308 2.2505
R21615 DVDD.n13311 DVDD.n13310 2.2505
R21616 DVDD.n12878 DVDD.n12877 2.2505
R21617 DVDD.n13316 DVDD.n13315 2.2505
R21618 DVDD.n13318 DVDD.n13317 2.2505
R21619 DVDD.n13320 DVDD.n13319 2.2505
R21620 DVDD.n12875 DVDD.n12874 2.2505
R21621 DVDD.n13325 DVDD.n13324 2.2505
R21622 DVDD.n13327 DVDD.n13326 2.2505
R21623 DVDD.n13329 DVDD.n13328 2.2505
R21624 DVDD.n12872 DVDD.n12871 2.2505
R21625 DVDD.n13334 DVDD.n13333 2.2505
R21626 DVDD.n13336 DVDD.n13335 2.2505
R21627 DVDD.n13338 DVDD.n13337 2.2505
R21628 DVDD.n12869 DVDD.n12868 2.2505
R21629 DVDD.n13343 DVDD.n13342 2.2505
R21630 DVDD.n13345 DVDD.n13344 2.2505
R21631 DVDD.n13347 DVDD.n13346 2.2505
R21632 DVDD.n12866 DVDD.n12865 2.2505
R21633 DVDD.n13352 DVDD.n13351 2.2505
R21634 DVDD.n13354 DVDD.n13353 2.2505
R21635 DVDD.n13356 DVDD.n13355 2.2505
R21636 DVDD.n12863 DVDD.n12862 2.2505
R21637 DVDD.n13361 DVDD.n13360 2.2505
R21638 DVDD.n13363 DVDD.n13362 2.2505
R21639 DVDD.n13365 DVDD.n13364 2.2505
R21640 DVDD.n12860 DVDD.n12859 2.2505
R21641 DVDD.n13370 DVDD.n13369 2.2505
R21642 DVDD.n13372 DVDD.n13371 2.2505
R21643 DVDD.n13374 DVDD.n13373 2.2505
R21644 DVDD.n12857 DVDD.n12856 2.2505
R21645 DVDD.n13379 DVDD.n13378 2.2505
R21646 DVDD.n13381 DVDD.n13380 2.2505
R21647 DVDD.n13383 DVDD.n13382 2.2505
R21648 DVDD.n12854 DVDD.n12853 2.2505
R21649 DVDD.n13388 DVDD.n13387 2.2505
R21650 DVDD.n13390 DVDD.n13389 2.2505
R21651 DVDD.n13392 DVDD.n13391 2.2505
R21652 DVDD.n12851 DVDD.n12850 2.2505
R21653 DVDD.n13397 DVDD.n13396 2.2505
R21654 DVDD.n13399 DVDD.n13398 2.2505
R21655 DVDD.n13401 DVDD.n13400 2.2505
R21656 DVDD.n12848 DVDD.n12847 2.2505
R21657 DVDD.n13406 DVDD.n13405 2.2505
R21658 DVDD.n13408 DVDD.n13407 2.2505
R21659 DVDD.n13410 DVDD.n13409 2.2505
R21660 DVDD.n12845 DVDD.n12844 2.2505
R21661 DVDD.n13415 DVDD.n13414 2.2505
R21662 DVDD.n13417 DVDD.n13416 2.2505
R21663 DVDD.n13419 DVDD.n13418 2.2505
R21664 DVDD.n12842 DVDD.n12841 2.2505
R21665 DVDD.n13424 DVDD.n13423 2.2505
R21666 DVDD.n13426 DVDD.n13425 2.2505
R21667 DVDD.n13428 DVDD.n13427 2.2505
R21668 DVDD.n12839 DVDD.n12838 2.2505
R21669 DVDD.n13433 DVDD.n13432 2.2505
R21670 DVDD.n13435 DVDD.n13434 2.2505
R21671 DVDD.n13437 DVDD.n13436 2.2505
R21672 DVDD.n12836 DVDD.n12835 2.2505
R21673 DVDD.n13442 DVDD.n13441 2.2505
R21674 DVDD.n13444 DVDD.n13443 2.2505
R21675 DVDD.n13446 DVDD.n13445 2.2505
R21676 DVDD.n12833 DVDD.n12832 2.2505
R21677 DVDD.n13451 DVDD.n13450 2.2505
R21678 DVDD.n13453 DVDD.n13452 2.2505
R21679 DVDD.n13455 DVDD.n13454 2.2505
R21680 DVDD.n12830 DVDD.n12829 2.2505
R21681 DVDD.n13460 DVDD.n13459 2.2505
R21682 DVDD.n13462 DVDD.n13461 2.2505
R21683 DVDD.n13464 DVDD.n13463 2.2505
R21684 DVDD.n12827 DVDD.n12826 2.2505
R21685 DVDD.n13469 DVDD.n13468 2.2505
R21686 DVDD.n13008 DVDD.n12915 2.2505
R21687 DVDD.n13010 DVDD.n13009 2.2505
R21688 DVDD.n13015 DVDD.n13011 2.2505
R21689 DVDD.n13016 DVDD.n13006 2.2505
R21690 DVDD.n13021 DVDD.n13020 2.2505
R21691 DVDD.n13022 DVDD.n13005 2.2505
R21692 DVDD.n13027 DVDD.n13023 2.2505
R21693 DVDD.n13028 DVDD.n13004 2.2505
R21694 DVDD.n13033 DVDD.n13032 2.2505
R21695 DVDD.n13034 DVDD.n13003 2.2505
R21696 DVDD.n13039 DVDD.n13035 2.2505
R21697 DVDD.n13040 DVDD.n13002 2.2505
R21698 DVDD.n13045 DVDD.n13044 2.2505
R21699 DVDD.n13046 DVDD.n13001 2.2505
R21700 DVDD.n13051 DVDD.n13047 2.2505
R21701 DVDD.n13052 DVDD.n13000 2.2505
R21702 DVDD.n13057 DVDD.n13056 2.2505
R21703 DVDD.n13058 DVDD.n12999 2.2505
R21704 DVDD.n13063 DVDD.n13059 2.2505
R21705 DVDD.n13064 DVDD.n12998 2.2505
R21706 DVDD.n13069 DVDD.n13068 2.2505
R21707 DVDD.n13070 DVDD.n12997 2.2505
R21708 DVDD.n13075 DVDD.n13071 2.2505
R21709 DVDD.n13076 DVDD.n12996 2.2505
R21710 DVDD.n13081 DVDD.n13080 2.2505
R21711 DVDD.n13082 DVDD.n12995 2.2505
R21712 DVDD.n13087 DVDD.n13083 2.2505
R21713 DVDD.n13088 DVDD.n12994 2.2505
R21714 DVDD.n13093 DVDD.n13092 2.2505
R21715 DVDD.n13094 DVDD.n12993 2.2505
R21716 DVDD.n13099 DVDD.n13095 2.2505
R21717 DVDD.n13100 DVDD.n12992 2.2505
R21718 DVDD.n13105 DVDD.n13104 2.2505
R21719 DVDD.n13106 DVDD.n12991 2.2505
R21720 DVDD.n13111 DVDD.n13107 2.2505
R21721 DVDD.n13112 DVDD.n12990 2.2505
R21722 DVDD.n13117 DVDD.n13116 2.2505
R21723 DVDD.n13118 DVDD.n12989 2.2505
R21724 DVDD.n13123 DVDD.n13119 2.2505
R21725 DVDD.n13124 DVDD.n12988 2.2505
R21726 DVDD.n13129 DVDD.n13128 2.2505
R21727 DVDD.n13130 DVDD.n12987 2.2505
R21728 DVDD.n13135 DVDD.n13131 2.2505
R21729 DVDD.n13136 DVDD.n12986 2.2505
R21730 DVDD.n13141 DVDD.n13140 2.2505
R21731 DVDD.n13142 DVDD.n12985 2.2505
R21732 DVDD.n13147 DVDD.n13143 2.2505
R21733 DVDD.n13148 DVDD.n12984 2.2505
R21734 DVDD.n13153 DVDD.n13152 2.2505
R21735 DVDD.n13154 DVDD.n12983 2.2505
R21736 DVDD.n13159 DVDD.n13155 2.2505
R21737 DVDD.n13160 DVDD.n12982 2.2505
R21738 DVDD.n13165 DVDD.n13164 2.2505
R21739 DVDD.n13166 DVDD.n12981 2.2505
R21740 DVDD.n13171 DVDD.n13167 2.2505
R21741 DVDD.n13172 DVDD.n12980 2.2505
R21742 DVDD.n13177 DVDD.n13176 2.2505
R21743 DVDD.n13178 DVDD.n12979 2.2505
R21744 DVDD.n13183 DVDD.n13179 2.2505
R21745 DVDD.n13184 DVDD.n12978 2.2505
R21746 DVDD.n13189 DVDD.n13188 2.2505
R21747 DVDD.n13190 DVDD.n12977 2.2505
R21748 DVDD.n13195 DVDD.n13191 2.2505
R21749 DVDD.n13196 DVDD.n12976 2.2505
R21750 DVDD.n13201 DVDD.n13200 2.2505
R21751 DVDD.n13202 DVDD.n12975 2.2505
R21752 DVDD.n13207 DVDD.n13203 2.2505
R21753 DVDD.n13208 DVDD.n12974 2.2505
R21754 DVDD.n13213 DVDD.n13212 2.2505
R21755 DVDD.n13214 DVDD.n12973 2.2505
R21756 DVDD.n13219 DVDD.n13215 2.2505
R21757 DVDD.n13220 DVDD.n12972 2.2505
R21758 DVDD.n13225 DVDD.n13224 2.2505
R21759 DVDD.n13226 DVDD.n12971 2.2505
R21760 DVDD.n13231 DVDD.n13227 2.2505
R21761 DVDD.n13232 DVDD.n12970 2.2505
R21762 DVDD.n13237 DVDD.n13236 2.2505
R21763 DVDD.n13238 DVDD.n12969 2.2505
R21764 DVDD.n13243 DVDD.n13239 2.2505
R21765 DVDD.n13244 DVDD.n12968 2.2505
R21766 DVDD.n13249 DVDD.n13248 2.2505
R21767 DVDD.n13250 DVDD.n12967 2.2505
R21768 DVDD.n13252 DVDD.n13251 2.2505
R21769 DVDD.n13253 DVDD.n12903 2.2505
R21770 DVDD.n13254 DVDD.n13253 2.2505
R21771 DVDD.n13252 DVDD.n12964 2.2505
R21772 DVDD.n12967 DVDD.n12966 2.2505
R21773 DVDD.n13248 DVDD.n13247 2.2505
R21774 DVDD.n13245 DVDD.n13244 2.2505
R21775 DVDD.n13243 DVDD.n13242 2.2505
R21776 DVDD.n13240 DVDD.n12969 2.2505
R21777 DVDD.n13236 DVDD.n13235 2.2505
R21778 DVDD.n13233 DVDD.n13232 2.2505
R21779 DVDD.n13231 DVDD.n13230 2.2505
R21780 DVDD.n13228 DVDD.n12971 2.2505
R21781 DVDD.n13224 DVDD.n13223 2.2505
R21782 DVDD.n13221 DVDD.n13220 2.2505
R21783 DVDD.n13219 DVDD.n13218 2.2505
R21784 DVDD.n13216 DVDD.n12973 2.2505
R21785 DVDD.n13212 DVDD.n13211 2.2505
R21786 DVDD.n13209 DVDD.n13208 2.2505
R21787 DVDD.n13207 DVDD.n13206 2.2505
R21788 DVDD.n13204 DVDD.n12975 2.2505
R21789 DVDD.n13200 DVDD.n13199 2.2505
R21790 DVDD.n13197 DVDD.n13196 2.2505
R21791 DVDD.n13195 DVDD.n13194 2.2505
R21792 DVDD.n13192 DVDD.n12977 2.2505
R21793 DVDD.n13188 DVDD.n13187 2.2505
R21794 DVDD.n13185 DVDD.n13184 2.2505
R21795 DVDD.n13183 DVDD.n13182 2.2505
R21796 DVDD.n13180 DVDD.n12979 2.2505
R21797 DVDD.n13176 DVDD.n13175 2.2505
R21798 DVDD.n13173 DVDD.n13172 2.2505
R21799 DVDD.n13171 DVDD.n13170 2.2505
R21800 DVDD.n13168 DVDD.n12981 2.2505
R21801 DVDD.n13164 DVDD.n13163 2.2505
R21802 DVDD.n13161 DVDD.n13160 2.2505
R21803 DVDD.n13159 DVDD.n13158 2.2505
R21804 DVDD.n13156 DVDD.n12983 2.2505
R21805 DVDD.n13152 DVDD.n13151 2.2505
R21806 DVDD.n13149 DVDD.n13148 2.2505
R21807 DVDD.n13147 DVDD.n13146 2.2505
R21808 DVDD.n13144 DVDD.n12985 2.2505
R21809 DVDD.n13140 DVDD.n13139 2.2505
R21810 DVDD.n13137 DVDD.n13136 2.2505
R21811 DVDD.n13135 DVDD.n13134 2.2505
R21812 DVDD.n13132 DVDD.n12987 2.2505
R21813 DVDD.n13128 DVDD.n13127 2.2505
R21814 DVDD.n13125 DVDD.n13124 2.2505
R21815 DVDD.n13123 DVDD.n13122 2.2505
R21816 DVDD.n13120 DVDD.n12989 2.2505
R21817 DVDD.n13116 DVDD.n13115 2.2505
R21818 DVDD.n13113 DVDD.n13112 2.2505
R21819 DVDD.n13111 DVDD.n13110 2.2505
R21820 DVDD.n13108 DVDD.n12991 2.2505
R21821 DVDD.n13104 DVDD.n13103 2.2505
R21822 DVDD.n13101 DVDD.n13100 2.2505
R21823 DVDD.n13099 DVDD.n13098 2.2505
R21824 DVDD.n13096 DVDD.n12993 2.2505
R21825 DVDD.n13092 DVDD.n13091 2.2505
R21826 DVDD.n13089 DVDD.n13088 2.2505
R21827 DVDD.n13087 DVDD.n13086 2.2505
R21828 DVDD.n13084 DVDD.n12995 2.2505
R21829 DVDD.n13080 DVDD.n13079 2.2505
R21830 DVDD.n13077 DVDD.n13076 2.2505
R21831 DVDD.n13075 DVDD.n13074 2.2505
R21832 DVDD.n13072 DVDD.n12997 2.2505
R21833 DVDD.n13068 DVDD.n13067 2.2505
R21834 DVDD.n13065 DVDD.n13064 2.2505
R21835 DVDD.n13063 DVDD.n13062 2.2505
R21836 DVDD.n13060 DVDD.n12999 2.2505
R21837 DVDD.n13056 DVDD.n13055 2.2505
R21838 DVDD.n13053 DVDD.n13052 2.2505
R21839 DVDD.n13051 DVDD.n13050 2.2505
R21840 DVDD.n13048 DVDD.n13001 2.2505
R21841 DVDD.n13044 DVDD.n13043 2.2505
R21842 DVDD.n13041 DVDD.n13040 2.2505
R21843 DVDD.n13039 DVDD.n13038 2.2505
R21844 DVDD.n13036 DVDD.n13003 2.2505
R21845 DVDD.n13032 DVDD.n13031 2.2505
R21846 DVDD.n13029 DVDD.n13028 2.2505
R21847 DVDD.n13027 DVDD.n13026 2.2505
R21848 DVDD.n13024 DVDD.n13005 2.2505
R21849 DVDD.n13020 DVDD.n13019 2.2505
R21850 DVDD.n13017 DVDD.n13016 2.2505
R21851 DVDD.n13015 DVDD.n13014 2.2505
R21852 DVDD.n13012 DVDD.n13009 2.2505
R21853 DVDD.n13008 DVDD.n13007 2.2505
R21854 DVDD.n2209 DVDD.n2159 2.2505
R21855 DVDD.n16700 DVDD.n16699 2.2505
R21856 DVDD.n16698 DVDD.n2211 2.2505
R21857 DVDD.n16697 DVDD.n16696 2.2505
R21858 DVDD.n16692 DVDD.n2212 2.2505
R21859 DVDD.n16688 DVDD.n16687 2.2505
R21860 DVDD.n16686 DVDD.n2213 2.2505
R21861 DVDD.n16685 DVDD.n16684 2.2505
R21862 DVDD.n16680 DVDD.n2214 2.2505
R21863 DVDD.n16676 DVDD.n16675 2.2505
R21864 DVDD.n16674 DVDD.n2215 2.2505
R21865 DVDD.n16673 DVDD.n16672 2.2505
R21866 DVDD.n16668 DVDD.n2216 2.2505
R21867 DVDD.n16664 DVDD.n16663 2.2505
R21868 DVDD.n16662 DVDD.n2217 2.2505
R21869 DVDD.n16661 DVDD.n16660 2.2505
R21870 DVDD.n16656 DVDD.n2218 2.2505
R21871 DVDD.n16652 DVDD.n16651 2.2505
R21872 DVDD.n16650 DVDD.n2219 2.2505
R21873 DVDD.n16649 DVDD.n16648 2.2505
R21874 DVDD.n16644 DVDD.n2220 2.2505
R21875 DVDD.n16640 DVDD.n16639 2.2505
R21876 DVDD.n16638 DVDD.n2221 2.2505
R21877 DVDD.n16637 DVDD.n16636 2.2505
R21878 DVDD.n16632 DVDD.n2222 2.2505
R21879 DVDD.n16628 DVDD.n16627 2.2505
R21880 DVDD.n16626 DVDD.n2223 2.2505
R21881 DVDD.n16625 DVDD.n16624 2.2505
R21882 DVDD.n16620 DVDD.n2224 2.2505
R21883 DVDD.n16616 DVDD.n16615 2.2505
R21884 DVDD.n16614 DVDD.n2225 2.2505
R21885 DVDD.n16613 DVDD.n16612 2.2505
R21886 DVDD.n16608 DVDD.n2226 2.2505
R21887 DVDD.n16604 DVDD.n16603 2.2505
R21888 DVDD.n16602 DVDD.n2227 2.2505
R21889 DVDD.n16601 DVDD.n16600 2.2505
R21890 DVDD.n16596 DVDD.n2228 2.2505
R21891 DVDD.n16592 DVDD.n16591 2.2505
R21892 DVDD.n16590 DVDD.n2229 2.2505
R21893 DVDD.n16589 DVDD.n16588 2.2505
R21894 DVDD.n16584 DVDD.n2230 2.2505
R21895 DVDD.n16580 DVDD.n16579 2.2505
R21896 DVDD.n16578 DVDD.n2231 2.2505
R21897 DVDD.n16577 DVDD.n16576 2.2505
R21898 DVDD.n16572 DVDD.n2232 2.2505
R21899 DVDD.n16568 DVDD.n16567 2.2505
R21900 DVDD.n16566 DVDD.n2233 2.2505
R21901 DVDD.n16565 DVDD.n16564 2.2505
R21902 DVDD.n16560 DVDD.n2234 2.2505
R21903 DVDD.n16556 DVDD.n16555 2.2505
R21904 DVDD.n16554 DVDD.n2235 2.2505
R21905 DVDD.n16553 DVDD.n16552 2.2505
R21906 DVDD.n16548 DVDD.n2236 2.2505
R21907 DVDD.n16544 DVDD.n16543 2.2505
R21908 DVDD.n16542 DVDD.n2237 2.2505
R21909 DVDD.n16541 DVDD.n16540 2.2505
R21910 DVDD.n16536 DVDD.n2238 2.2505
R21911 DVDD.n16532 DVDD.n16531 2.2505
R21912 DVDD.n16530 DVDD.n2239 2.2505
R21913 DVDD.n16529 DVDD.n16528 2.2505
R21914 DVDD.n16524 DVDD.n2240 2.2505
R21915 DVDD.n16520 DVDD.n16519 2.2505
R21916 DVDD.n16518 DVDD.n2241 2.2505
R21917 DVDD.n16517 DVDD.n16516 2.2505
R21918 DVDD.n16512 DVDD.n2242 2.2505
R21919 DVDD.n16508 DVDD.n16507 2.2505
R21920 DVDD.n16506 DVDD.n2243 2.2505
R21921 DVDD.n16505 DVDD.n16504 2.2505
R21922 DVDD.n16500 DVDD.n2244 2.2505
R21923 DVDD.n16496 DVDD.n16495 2.2505
R21924 DVDD.n16494 DVDD.n2245 2.2505
R21925 DVDD.n16493 DVDD.n16492 2.2505
R21926 DVDD.n16488 DVDD.n2246 2.2505
R21927 DVDD.n16484 DVDD.n16483 2.2505
R21928 DVDD.n16482 DVDD.n2247 2.2505
R21929 DVDD.n16481 DVDD.n16480 2.2505
R21930 DVDD.n16476 DVDD.n2248 2.2505
R21931 DVDD.n16472 DVDD.n16471 2.2505
R21932 DVDD.n16470 DVDD.n2249 2.2505
R21933 DVDD.n16469 DVDD.n16468 2.2505
R21934 DVDD.n16464 DVDD.n2250 2.2505
R21935 DVDD.n16460 DVDD.n16459 2.2505
R21936 DVDD.n16458 DVDD.n2253 2.2505
R21937 DVDD.n16457 DVDD.n16456 2.2505
R21938 DVDD.n16456 DVDD.n2207 2.2505
R21939 DVDD.n2253 DVDD.n2252 2.2505
R21940 DVDD.n16461 DVDD.n16460 2.2505
R21941 DVDD.n16464 DVDD.n16463 2.2505
R21942 DVDD.n16468 DVDD.n16467 2.2505
R21943 DVDD.n16465 DVDD.n2249 2.2505
R21944 DVDD.n16473 DVDD.n16472 2.2505
R21945 DVDD.n16476 DVDD.n16475 2.2505
R21946 DVDD.n16480 DVDD.n16479 2.2505
R21947 DVDD.n16477 DVDD.n2247 2.2505
R21948 DVDD.n16485 DVDD.n16484 2.2505
R21949 DVDD.n16488 DVDD.n16487 2.2505
R21950 DVDD.n16492 DVDD.n16491 2.2505
R21951 DVDD.n16489 DVDD.n2245 2.2505
R21952 DVDD.n16497 DVDD.n16496 2.2505
R21953 DVDD.n16500 DVDD.n16499 2.2505
R21954 DVDD.n16504 DVDD.n16503 2.2505
R21955 DVDD.n16501 DVDD.n2243 2.2505
R21956 DVDD.n16509 DVDD.n16508 2.2505
R21957 DVDD.n16512 DVDD.n16511 2.2505
R21958 DVDD.n16516 DVDD.n16515 2.2505
R21959 DVDD.n16513 DVDD.n2241 2.2505
R21960 DVDD.n16521 DVDD.n16520 2.2505
R21961 DVDD.n16524 DVDD.n16523 2.2505
R21962 DVDD.n16528 DVDD.n16527 2.2505
R21963 DVDD.n16525 DVDD.n2239 2.2505
R21964 DVDD.n16533 DVDD.n16532 2.2505
R21965 DVDD.n16536 DVDD.n16535 2.2505
R21966 DVDD.n16540 DVDD.n16539 2.2505
R21967 DVDD.n16537 DVDD.n2237 2.2505
R21968 DVDD.n16545 DVDD.n16544 2.2505
R21969 DVDD.n16548 DVDD.n16547 2.2505
R21970 DVDD.n16552 DVDD.n16551 2.2505
R21971 DVDD.n16549 DVDD.n2235 2.2505
R21972 DVDD.n16557 DVDD.n16556 2.2505
R21973 DVDD.n16560 DVDD.n16559 2.2505
R21974 DVDD.n16564 DVDD.n16563 2.2505
R21975 DVDD.n16561 DVDD.n2233 2.2505
R21976 DVDD.n16569 DVDD.n16568 2.2505
R21977 DVDD.n16572 DVDD.n16571 2.2505
R21978 DVDD.n16576 DVDD.n16575 2.2505
R21979 DVDD.n16573 DVDD.n2231 2.2505
R21980 DVDD.n16581 DVDD.n16580 2.2505
R21981 DVDD.n16584 DVDD.n16583 2.2505
R21982 DVDD.n16588 DVDD.n16587 2.2505
R21983 DVDD.n16585 DVDD.n2229 2.2505
R21984 DVDD.n16593 DVDD.n16592 2.2505
R21985 DVDD.n16596 DVDD.n16595 2.2505
R21986 DVDD.n16600 DVDD.n16599 2.2505
R21987 DVDD.n16597 DVDD.n2227 2.2505
R21988 DVDD.n16605 DVDD.n16604 2.2505
R21989 DVDD.n16608 DVDD.n16607 2.2505
R21990 DVDD.n16612 DVDD.n16611 2.2505
R21991 DVDD.n16609 DVDD.n2225 2.2505
R21992 DVDD.n16617 DVDD.n16616 2.2505
R21993 DVDD.n16620 DVDD.n16619 2.2505
R21994 DVDD.n16624 DVDD.n16623 2.2505
R21995 DVDD.n16621 DVDD.n2223 2.2505
R21996 DVDD.n16629 DVDD.n16628 2.2505
R21997 DVDD.n16632 DVDD.n16631 2.2505
R21998 DVDD.n16636 DVDD.n16635 2.2505
R21999 DVDD.n16633 DVDD.n2221 2.2505
R22000 DVDD.n16641 DVDD.n16640 2.2505
R22001 DVDD.n16644 DVDD.n16643 2.2505
R22002 DVDD.n16648 DVDD.n16647 2.2505
R22003 DVDD.n16645 DVDD.n2219 2.2505
R22004 DVDD.n16653 DVDD.n16652 2.2505
R22005 DVDD.n16656 DVDD.n16655 2.2505
R22006 DVDD.n16660 DVDD.n16659 2.2505
R22007 DVDD.n16657 DVDD.n2217 2.2505
R22008 DVDD.n16665 DVDD.n16664 2.2505
R22009 DVDD.n16668 DVDD.n16667 2.2505
R22010 DVDD.n16672 DVDD.n16671 2.2505
R22011 DVDD.n16669 DVDD.n2215 2.2505
R22012 DVDD.n16677 DVDD.n16676 2.2505
R22013 DVDD.n16680 DVDD.n16679 2.2505
R22014 DVDD.n16684 DVDD.n16683 2.2505
R22015 DVDD.n16681 DVDD.n2213 2.2505
R22016 DVDD.n16689 DVDD.n16688 2.2505
R22017 DVDD.n16692 DVDD.n16691 2.2505
R22018 DVDD.n16696 DVDD.n16695 2.2505
R22019 DVDD.n16693 DVDD.n2211 2.2505
R22020 DVDD.n16701 DVDD.n16700 2.2505
R22021 DVDD.n16703 DVDD.n2209 2.2505
R22022 DVDD.n1909 DVDD.n1908 2.2505
R22023 DVDD.n1910 DVDD.n1906 2.2505
R22024 DVDD.n1915 DVDD.n1911 2.2505
R22025 DVDD.n1916 DVDD.n1905 2.2505
R22026 DVDD.n1921 DVDD.n1920 2.2505
R22027 DVDD.n1922 DVDD.n1904 2.2505
R22028 DVDD.n1927 DVDD.n1923 2.2505
R22029 DVDD.n1928 DVDD.n1903 2.2505
R22030 DVDD.n1933 DVDD.n1932 2.2505
R22031 DVDD.n1934 DVDD.n1902 2.2505
R22032 DVDD.n1939 DVDD.n1935 2.2505
R22033 DVDD.n1940 DVDD.n1901 2.2505
R22034 DVDD.n1945 DVDD.n1944 2.2505
R22035 DVDD.n1946 DVDD.n1900 2.2505
R22036 DVDD.n1951 DVDD.n1947 2.2505
R22037 DVDD.n1952 DVDD.n1899 2.2505
R22038 DVDD.n1957 DVDD.n1956 2.2505
R22039 DVDD.n1958 DVDD.n1898 2.2505
R22040 DVDD.n1963 DVDD.n1959 2.2505
R22041 DVDD.n1964 DVDD.n1897 2.2505
R22042 DVDD.n1969 DVDD.n1968 2.2505
R22043 DVDD.n1970 DVDD.n1896 2.2505
R22044 DVDD.n1975 DVDD.n1971 2.2505
R22045 DVDD.n1976 DVDD.n1895 2.2505
R22046 DVDD.n1981 DVDD.n1980 2.2505
R22047 DVDD.n1982 DVDD.n1894 2.2505
R22048 DVDD.n1987 DVDD.n1983 2.2505
R22049 DVDD.n1988 DVDD.n1893 2.2505
R22050 DVDD.n1993 DVDD.n1992 2.2505
R22051 DVDD.n1994 DVDD.n1892 2.2505
R22052 DVDD.n1999 DVDD.n1995 2.2505
R22053 DVDD.n2000 DVDD.n1891 2.2505
R22054 DVDD.n2005 DVDD.n2004 2.2505
R22055 DVDD.n2006 DVDD.n1890 2.2505
R22056 DVDD.n2011 DVDD.n2007 2.2505
R22057 DVDD.n2012 DVDD.n1889 2.2505
R22058 DVDD.n2017 DVDD.n2016 2.2505
R22059 DVDD.n2018 DVDD.n1888 2.2505
R22060 DVDD.n2023 DVDD.n2019 2.2505
R22061 DVDD.n2024 DVDD.n1887 2.2505
R22062 DVDD.n2029 DVDD.n2028 2.2505
R22063 DVDD.n2030 DVDD.n1886 2.2505
R22064 DVDD.n2035 DVDD.n2031 2.2505
R22065 DVDD.n2036 DVDD.n1885 2.2505
R22066 DVDD.n2041 DVDD.n2040 2.2505
R22067 DVDD.n2042 DVDD.n1884 2.2505
R22068 DVDD.n2047 DVDD.n2043 2.2505
R22069 DVDD.n2048 DVDD.n1883 2.2505
R22070 DVDD.n2053 DVDD.n2052 2.2505
R22071 DVDD.n2054 DVDD.n1882 2.2505
R22072 DVDD.n2059 DVDD.n2055 2.2505
R22073 DVDD.n2060 DVDD.n1881 2.2505
R22074 DVDD.n2065 DVDD.n2064 2.2505
R22075 DVDD.n2066 DVDD.n1880 2.2505
R22076 DVDD.n2071 DVDD.n2067 2.2505
R22077 DVDD.n2072 DVDD.n1879 2.2505
R22078 DVDD.n2077 DVDD.n2076 2.2505
R22079 DVDD.n2078 DVDD.n1878 2.2505
R22080 DVDD.n2083 DVDD.n2079 2.2505
R22081 DVDD.n2084 DVDD.n1877 2.2505
R22082 DVDD.n2089 DVDD.n2088 2.2505
R22083 DVDD.n2090 DVDD.n1876 2.2505
R22084 DVDD.n2095 DVDD.n2091 2.2505
R22085 DVDD.n2096 DVDD.n1875 2.2505
R22086 DVDD.n2101 DVDD.n2100 2.2505
R22087 DVDD.n2102 DVDD.n1874 2.2505
R22088 DVDD.n2107 DVDD.n2103 2.2505
R22089 DVDD.n2108 DVDD.n1873 2.2505
R22090 DVDD.n2113 DVDD.n2112 2.2505
R22091 DVDD.n2114 DVDD.n1872 2.2505
R22092 DVDD.n2119 DVDD.n2115 2.2505
R22093 DVDD.n2120 DVDD.n1871 2.2505
R22094 DVDD.n2125 DVDD.n2124 2.2505
R22095 DVDD.n2126 DVDD.n1870 2.2505
R22096 DVDD.n2131 DVDD.n2127 2.2505
R22097 DVDD.n2132 DVDD.n1869 2.2505
R22098 DVDD.n2137 DVDD.n2136 2.2505
R22099 DVDD.n2138 DVDD.n1868 2.2505
R22100 DVDD.n2143 DVDD.n2139 2.2505
R22101 DVDD.n2144 DVDD.n1867 2.2505
R22102 DVDD.n2149 DVDD.n2148 2.2505
R22103 DVDD.n2150 DVDD.n1866 2.2505
R22104 DVDD.n2152 DVDD.n2151 2.2505
R22105 DVDD.n2153 DVDD.n1817 2.2505
R22106 DVDD.n2154 DVDD.n2153 2.2505
R22107 DVDD.n2152 DVDD.n1863 2.2505
R22108 DVDD.n1866 DVDD.n1865 2.2505
R22109 DVDD.n2148 DVDD.n2147 2.2505
R22110 DVDD.n2145 DVDD.n2144 2.2505
R22111 DVDD.n2143 DVDD.n2142 2.2505
R22112 DVDD.n2140 DVDD.n1868 2.2505
R22113 DVDD.n2136 DVDD.n2135 2.2505
R22114 DVDD.n2133 DVDD.n2132 2.2505
R22115 DVDD.n2131 DVDD.n2130 2.2505
R22116 DVDD.n2128 DVDD.n1870 2.2505
R22117 DVDD.n2124 DVDD.n2123 2.2505
R22118 DVDD.n2121 DVDD.n2120 2.2505
R22119 DVDD.n2119 DVDD.n2118 2.2505
R22120 DVDD.n2116 DVDD.n1872 2.2505
R22121 DVDD.n2112 DVDD.n2111 2.2505
R22122 DVDD.n2109 DVDD.n2108 2.2505
R22123 DVDD.n2107 DVDD.n2106 2.2505
R22124 DVDD.n2104 DVDD.n1874 2.2505
R22125 DVDD.n2100 DVDD.n2099 2.2505
R22126 DVDD.n2097 DVDD.n2096 2.2505
R22127 DVDD.n2095 DVDD.n2094 2.2505
R22128 DVDD.n2092 DVDD.n1876 2.2505
R22129 DVDD.n2088 DVDD.n2087 2.2505
R22130 DVDD.n2085 DVDD.n2084 2.2505
R22131 DVDD.n2083 DVDD.n2082 2.2505
R22132 DVDD.n2080 DVDD.n1878 2.2505
R22133 DVDD.n2076 DVDD.n2075 2.2505
R22134 DVDD.n2073 DVDD.n2072 2.2505
R22135 DVDD.n2071 DVDD.n2070 2.2505
R22136 DVDD.n2068 DVDD.n1880 2.2505
R22137 DVDD.n2064 DVDD.n2063 2.2505
R22138 DVDD.n2061 DVDD.n2060 2.2505
R22139 DVDD.n2059 DVDD.n2058 2.2505
R22140 DVDD.n2056 DVDD.n1882 2.2505
R22141 DVDD.n2052 DVDD.n2051 2.2505
R22142 DVDD.n2049 DVDD.n2048 2.2505
R22143 DVDD.n2047 DVDD.n2046 2.2505
R22144 DVDD.n2044 DVDD.n1884 2.2505
R22145 DVDD.n2040 DVDD.n2039 2.2505
R22146 DVDD.n2037 DVDD.n2036 2.2505
R22147 DVDD.n2035 DVDD.n2034 2.2505
R22148 DVDD.n2032 DVDD.n1886 2.2505
R22149 DVDD.n2028 DVDD.n2027 2.2505
R22150 DVDD.n2025 DVDD.n2024 2.2505
R22151 DVDD.n2023 DVDD.n2022 2.2505
R22152 DVDD.n2020 DVDD.n1888 2.2505
R22153 DVDD.n2016 DVDD.n2015 2.2505
R22154 DVDD.n2013 DVDD.n2012 2.2505
R22155 DVDD.n2011 DVDD.n2010 2.2505
R22156 DVDD.n2008 DVDD.n1890 2.2505
R22157 DVDD.n2004 DVDD.n2003 2.2505
R22158 DVDD.n2001 DVDD.n2000 2.2505
R22159 DVDD.n1999 DVDD.n1998 2.2505
R22160 DVDD.n1996 DVDD.n1892 2.2505
R22161 DVDD.n1992 DVDD.n1991 2.2505
R22162 DVDD.n1989 DVDD.n1988 2.2505
R22163 DVDD.n1987 DVDD.n1986 2.2505
R22164 DVDD.n1984 DVDD.n1894 2.2505
R22165 DVDD.n1980 DVDD.n1979 2.2505
R22166 DVDD.n1977 DVDD.n1976 2.2505
R22167 DVDD.n1975 DVDD.n1974 2.2505
R22168 DVDD.n1972 DVDD.n1896 2.2505
R22169 DVDD.n1968 DVDD.n1967 2.2505
R22170 DVDD.n1965 DVDD.n1964 2.2505
R22171 DVDD.n1963 DVDD.n1962 2.2505
R22172 DVDD.n1960 DVDD.n1898 2.2505
R22173 DVDD.n1956 DVDD.n1955 2.2505
R22174 DVDD.n1953 DVDD.n1952 2.2505
R22175 DVDD.n1951 DVDD.n1950 2.2505
R22176 DVDD.n1948 DVDD.n1900 2.2505
R22177 DVDD.n1944 DVDD.n1943 2.2505
R22178 DVDD.n1941 DVDD.n1940 2.2505
R22179 DVDD.n1939 DVDD.n1938 2.2505
R22180 DVDD.n1936 DVDD.n1902 2.2505
R22181 DVDD.n1932 DVDD.n1931 2.2505
R22182 DVDD.n1929 DVDD.n1928 2.2505
R22183 DVDD.n1927 DVDD.n1926 2.2505
R22184 DVDD.n1924 DVDD.n1904 2.2505
R22185 DVDD.n1920 DVDD.n1919 2.2505
R22186 DVDD.n1917 DVDD.n1916 2.2505
R22187 DVDD.n1915 DVDD.n1914 2.2505
R22188 DVDD.n1912 DVDD.n1906 2.2505
R22189 DVDD.n1908 DVDD.n1907 2.2505
R22190 DVDD.n16988 DVDD.n1756 2.2505
R22191 DVDD.n16990 DVDD.n16989 2.2505
R22192 DVDD.n16987 DVDD.n1758 2.2505
R22193 DVDD.n16986 DVDD.n16985 2.2505
R22194 DVDD.n16981 DVDD.n1759 2.2505
R22195 DVDD.n16977 DVDD.n16976 2.2505
R22196 DVDD.n16975 DVDD.n1760 2.2505
R22197 DVDD.n16974 DVDD.n16973 2.2505
R22198 DVDD.n16969 DVDD.n1761 2.2505
R22199 DVDD.n16965 DVDD.n16964 2.2505
R22200 DVDD.n16963 DVDD.n1762 2.2505
R22201 DVDD.n16962 DVDD.n16961 2.2505
R22202 DVDD.n16957 DVDD.n1763 2.2505
R22203 DVDD.n16953 DVDD.n16952 2.2505
R22204 DVDD.n16951 DVDD.n1764 2.2505
R22205 DVDD.n16950 DVDD.n16949 2.2505
R22206 DVDD.n16945 DVDD.n1765 2.2505
R22207 DVDD.n16941 DVDD.n16940 2.2505
R22208 DVDD.n16939 DVDD.n1766 2.2505
R22209 DVDD.n16938 DVDD.n16937 2.2505
R22210 DVDD.n16933 DVDD.n1767 2.2505
R22211 DVDD.n16929 DVDD.n16928 2.2505
R22212 DVDD.n16927 DVDD.n1768 2.2505
R22213 DVDD.n16926 DVDD.n16925 2.2505
R22214 DVDD.n16921 DVDD.n1769 2.2505
R22215 DVDD.n16917 DVDD.n16916 2.2505
R22216 DVDD.n16915 DVDD.n1770 2.2505
R22217 DVDD.n16914 DVDD.n16913 2.2505
R22218 DVDD.n16909 DVDD.n1771 2.2505
R22219 DVDD.n16905 DVDD.n16904 2.2505
R22220 DVDD.n16903 DVDD.n1772 2.2505
R22221 DVDD.n16902 DVDD.n16901 2.2505
R22222 DVDD.n16897 DVDD.n1773 2.2505
R22223 DVDD.n16893 DVDD.n16892 2.2505
R22224 DVDD.n16891 DVDD.n1774 2.2505
R22225 DVDD.n16890 DVDD.n16889 2.2505
R22226 DVDD.n16885 DVDD.n1775 2.2505
R22227 DVDD.n16881 DVDD.n16880 2.2505
R22228 DVDD.n16879 DVDD.n1776 2.2505
R22229 DVDD.n16878 DVDD.n16877 2.2505
R22230 DVDD.n16873 DVDD.n1777 2.2505
R22231 DVDD.n16869 DVDD.n16868 2.2505
R22232 DVDD.n16867 DVDD.n1778 2.2505
R22233 DVDD.n16866 DVDD.n16865 2.2505
R22234 DVDD.n16861 DVDD.n1779 2.2505
R22235 DVDD.n16857 DVDD.n16856 2.2505
R22236 DVDD.n16855 DVDD.n1780 2.2505
R22237 DVDD.n16854 DVDD.n16853 2.2505
R22238 DVDD.n16849 DVDD.n1781 2.2505
R22239 DVDD.n16845 DVDD.n16844 2.2505
R22240 DVDD.n16843 DVDD.n1782 2.2505
R22241 DVDD.n16842 DVDD.n16841 2.2505
R22242 DVDD.n16837 DVDD.n1783 2.2505
R22243 DVDD.n16833 DVDD.n16832 2.2505
R22244 DVDD.n16831 DVDD.n1784 2.2505
R22245 DVDD.n16830 DVDD.n16829 2.2505
R22246 DVDD.n16825 DVDD.n1785 2.2505
R22247 DVDD.n16821 DVDD.n16820 2.2505
R22248 DVDD.n16819 DVDD.n1786 2.2505
R22249 DVDD.n16818 DVDD.n16817 2.2505
R22250 DVDD.n16813 DVDD.n1787 2.2505
R22251 DVDD.n16809 DVDD.n16808 2.2505
R22252 DVDD.n16807 DVDD.n1788 2.2505
R22253 DVDD.n16806 DVDD.n16805 2.2505
R22254 DVDD.n16801 DVDD.n1789 2.2505
R22255 DVDD.n16797 DVDD.n16796 2.2505
R22256 DVDD.n16795 DVDD.n1790 2.2505
R22257 DVDD.n16794 DVDD.n16793 2.2505
R22258 DVDD.n16789 DVDD.n1791 2.2505
R22259 DVDD.n16785 DVDD.n16784 2.2505
R22260 DVDD.n16783 DVDD.n1792 2.2505
R22261 DVDD.n16782 DVDD.n16781 2.2505
R22262 DVDD.n16777 DVDD.n1793 2.2505
R22263 DVDD.n16773 DVDD.n16772 2.2505
R22264 DVDD.n16771 DVDD.n1794 2.2505
R22265 DVDD.n16770 DVDD.n16769 2.2505
R22266 DVDD.n16765 DVDD.n1795 2.2505
R22267 DVDD.n16761 DVDD.n16760 2.2505
R22268 DVDD.n16759 DVDD.n1796 2.2505
R22269 DVDD.n16758 DVDD.n16757 2.2505
R22270 DVDD.n16753 DVDD.n1797 2.2505
R22271 DVDD.n16749 DVDD.n16748 2.2505
R22272 DVDD.n16747 DVDD.n1800 2.2505
R22273 DVDD.n16746 DVDD.n16745 2.2505
R22274 DVDD.n16745 DVDD.n1754 2.2505
R22275 DVDD.n1800 DVDD.n1799 2.2505
R22276 DVDD.n16750 DVDD.n16749 2.2505
R22277 DVDD.n16753 DVDD.n16752 2.2505
R22278 DVDD.n16757 DVDD.n16756 2.2505
R22279 DVDD.n16754 DVDD.n1796 2.2505
R22280 DVDD.n16762 DVDD.n16761 2.2505
R22281 DVDD.n16765 DVDD.n16764 2.2505
R22282 DVDD.n16769 DVDD.n16768 2.2505
R22283 DVDD.n16766 DVDD.n1794 2.2505
R22284 DVDD.n16774 DVDD.n16773 2.2505
R22285 DVDD.n16777 DVDD.n16776 2.2505
R22286 DVDD.n16781 DVDD.n16780 2.2505
R22287 DVDD.n16778 DVDD.n1792 2.2505
R22288 DVDD.n16786 DVDD.n16785 2.2505
R22289 DVDD.n16789 DVDD.n16788 2.2505
R22290 DVDD.n16793 DVDD.n16792 2.2505
R22291 DVDD.n16790 DVDD.n1790 2.2505
R22292 DVDD.n16798 DVDD.n16797 2.2505
R22293 DVDD.n16801 DVDD.n16800 2.2505
R22294 DVDD.n16805 DVDD.n16804 2.2505
R22295 DVDD.n16802 DVDD.n1788 2.2505
R22296 DVDD.n16810 DVDD.n16809 2.2505
R22297 DVDD.n16813 DVDD.n16812 2.2505
R22298 DVDD.n16817 DVDD.n16816 2.2505
R22299 DVDD.n16814 DVDD.n1786 2.2505
R22300 DVDD.n16822 DVDD.n16821 2.2505
R22301 DVDD.n16825 DVDD.n16824 2.2505
R22302 DVDD.n16829 DVDD.n16828 2.2505
R22303 DVDD.n16826 DVDD.n1784 2.2505
R22304 DVDD.n16834 DVDD.n16833 2.2505
R22305 DVDD.n16837 DVDD.n16836 2.2505
R22306 DVDD.n16841 DVDD.n16840 2.2505
R22307 DVDD.n16838 DVDD.n1782 2.2505
R22308 DVDD.n16846 DVDD.n16845 2.2505
R22309 DVDD.n16849 DVDD.n16848 2.2505
R22310 DVDD.n16853 DVDD.n16852 2.2505
R22311 DVDD.n16850 DVDD.n1780 2.2505
R22312 DVDD.n16858 DVDD.n16857 2.2505
R22313 DVDD.n16861 DVDD.n16860 2.2505
R22314 DVDD.n16865 DVDD.n16864 2.2505
R22315 DVDD.n16862 DVDD.n1778 2.2505
R22316 DVDD.n16870 DVDD.n16869 2.2505
R22317 DVDD.n16873 DVDD.n16872 2.2505
R22318 DVDD.n16877 DVDD.n16876 2.2505
R22319 DVDD.n16874 DVDD.n1776 2.2505
R22320 DVDD.n16882 DVDD.n16881 2.2505
R22321 DVDD.n16885 DVDD.n16884 2.2505
R22322 DVDD.n16889 DVDD.n16888 2.2505
R22323 DVDD.n16886 DVDD.n1774 2.2505
R22324 DVDD.n16894 DVDD.n16893 2.2505
R22325 DVDD.n16897 DVDD.n16896 2.2505
R22326 DVDD.n16901 DVDD.n16900 2.2505
R22327 DVDD.n16898 DVDD.n1772 2.2505
R22328 DVDD.n16906 DVDD.n16905 2.2505
R22329 DVDD.n16909 DVDD.n16908 2.2505
R22330 DVDD.n16913 DVDD.n16912 2.2505
R22331 DVDD.n16910 DVDD.n1770 2.2505
R22332 DVDD.n16918 DVDD.n16917 2.2505
R22333 DVDD.n16921 DVDD.n16920 2.2505
R22334 DVDD.n16925 DVDD.n16924 2.2505
R22335 DVDD.n16922 DVDD.n1768 2.2505
R22336 DVDD.n16930 DVDD.n16929 2.2505
R22337 DVDD.n16933 DVDD.n16932 2.2505
R22338 DVDD.n16937 DVDD.n16936 2.2505
R22339 DVDD.n16934 DVDD.n1766 2.2505
R22340 DVDD.n16942 DVDD.n16941 2.2505
R22341 DVDD.n16945 DVDD.n16944 2.2505
R22342 DVDD.n16949 DVDD.n16948 2.2505
R22343 DVDD.n16946 DVDD.n1764 2.2505
R22344 DVDD.n16954 DVDD.n16953 2.2505
R22345 DVDD.n16957 DVDD.n16956 2.2505
R22346 DVDD.n16961 DVDD.n16960 2.2505
R22347 DVDD.n16958 DVDD.n1762 2.2505
R22348 DVDD.n16966 DVDD.n16965 2.2505
R22349 DVDD.n16969 DVDD.n16968 2.2505
R22350 DVDD.n16973 DVDD.n16972 2.2505
R22351 DVDD.n16970 DVDD.n1760 2.2505
R22352 DVDD.n16978 DVDD.n16977 2.2505
R22353 DVDD.n16981 DVDD.n16980 2.2505
R22354 DVDD.n16985 DVDD.n16984 2.2505
R22355 DVDD.n16982 DVDD.n1758 2.2505
R22356 DVDD.n16991 DVDD.n16990 2.2505
R22357 DVDD.n16993 DVDD.n1756 2.2505
R22358 DVDD.n17256 DVDD.n1657 2.2505
R22359 DVDD.n17258 DVDD.n17257 2.2505
R22360 DVDD.n17255 DVDD.n1659 2.2505
R22361 DVDD.n17254 DVDD.n17253 2.2505
R22362 DVDD.n17249 DVDD.n1660 2.2505
R22363 DVDD.n17245 DVDD.n17244 2.2505
R22364 DVDD.n17243 DVDD.n1661 2.2505
R22365 DVDD.n17242 DVDD.n17241 2.2505
R22366 DVDD.n17237 DVDD.n1662 2.2505
R22367 DVDD.n17233 DVDD.n17232 2.2505
R22368 DVDD.n17231 DVDD.n1663 2.2505
R22369 DVDD.n17230 DVDD.n17229 2.2505
R22370 DVDD.n17225 DVDD.n1664 2.2505
R22371 DVDD.n17221 DVDD.n17220 2.2505
R22372 DVDD.n17219 DVDD.n1665 2.2505
R22373 DVDD.n17218 DVDD.n17217 2.2505
R22374 DVDD.n17213 DVDD.n1666 2.2505
R22375 DVDD.n17209 DVDD.n17208 2.2505
R22376 DVDD.n17207 DVDD.n1667 2.2505
R22377 DVDD.n17206 DVDD.n17205 2.2505
R22378 DVDD.n17201 DVDD.n1668 2.2505
R22379 DVDD.n17197 DVDD.n17196 2.2505
R22380 DVDD.n17195 DVDD.n1669 2.2505
R22381 DVDD.n17194 DVDD.n17193 2.2505
R22382 DVDD.n17189 DVDD.n1670 2.2505
R22383 DVDD.n17185 DVDD.n17184 2.2505
R22384 DVDD.n17183 DVDD.n1671 2.2505
R22385 DVDD.n17182 DVDD.n17181 2.2505
R22386 DVDD.n17177 DVDD.n1672 2.2505
R22387 DVDD.n17173 DVDD.n17172 2.2505
R22388 DVDD.n17171 DVDD.n1673 2.2505
R22389 DVDD.n17170 DVDD.n17169 2.2505
R22390 DVDD.n17165 DVDD.n1674 2.2505
R22391 DVDD.n17161 DVDD.n17160 2.2505
R22392 DVDD.n17159 DVDD.n1675 2.2505
R22393 DVDD.n17158 DVDD.n17157 2.2505
R22394 DVDD.n17153 DVDD.n1676 2.2505
R22395 DVDD.n17149 DVDD.n17148 2.2505
R22396 DVDD.n17147 DVDD.n1677 2.2505
R22397 DVDD.n17146 DVDD.n17145 2.2505
R22398 DVDD.n17141 DVDD.n1678 2.2505
R22399 DVDD.n17137 DVDD.n17136 2.2505
R22400 DVDD.n17135 DVDD.n1679 2.2505
R22401 DVDD.n17134 DVDD.n17133 2.2505
R22402 DVDD.n17129 DVDD.n1680 2.2505
R22403 DVDD.n17125 DVDD.n17124 2.2505
R22404 DVDD.n17123 DVDD.n1681 2.2505
R22405 DVDD.n17122 DVDD.n17121 2.2505
R22406 DVDD.n17117 DVDD.n1682 2.2505
R22407 DVDD.n17113 DVDD.n17112 2.2505
R22408 DVDD.n17111 DVDD.n1683 2.2505
R22409 DVDD.n17110 DVDD.n17109 2.2505
R22410 DVDD.n17105 DVDD.n1684 2.2505
R22411 DVDD.n17101 DVDD.n17100 2.2505
R22412 DVDD.n17099 DVDD.n1685 2.2505
R22413 DVDD.n17098 DVDD.n17097 2.2505
R22414 DVDD.n17093 DVDD.n1686 2.2505
R22415 DVDD.n17089 DVDD.n17088 2.2505
R22416 DVDD.n17087 DVDD.n1687 2.2505
R22417 DVDD.n17086 DVDD.n17085 2.2505
R22418 DVDD.n17081 DVDD.n1688 2.2505
R22419 DVDD.n17077 DVDD.n17076 2.2505
R22420 DVDD.n17075 DVDD.n1689 2.2505
R22421 DVDD.n17074 DVDD.n17073 2.2505
R22422 DVDD.n17069 DVDD.n1690 2.2505
R22423 DVDD.n17065 DVDD.n17064 2.2505
R22424 DVDD.n17063 DVDD.n1691 2.2505
R22425 DVDD.n17062 DVDD.n17061 2.2505
R22426 DVDD.n17057 DVDD.n1692 2.2505
R22427 DVDD.n17053 DVDD.n17052 2.2505
R22428 DVDD.n17051 DVDD.n1693 2.2505
R22429 DVDD.n17050 DVDD.n17049 2.2505
R22430 DVDD.n17045 DVDD.n1694 2.2505
R22431 DVDD.n17041 DVDD.n17040 2.2505
R22432 DVDD.n17039 DVDD.n1695 2.2505
R22433 DVDD.n17038 DVDD.n17037 2.2505
R22434 DVDD.n17033 DVDD.n1696 2.2505
R22435 DVDD.n17029 DVDD.n17028 2.2505
R22436 DVDD.n17027 DVDD.n1697 2.2505
R22437 DVDD.n17026 DVDD.n17025 2.2505
R22438 DVDD.n17021 DVDD.n1698 2.2505
R22439 DVDD.n17017 DVDD.n17016 2.2505
R22440 DVDD.n17015 DVDD.n1701 2.2505
R22441 DVDD.n17014 DVDD.n17013 2.2505
R22442 DVDD.n17013 DVDD.n1653 2.2505
R22443 DVDD.n1701 DVDD.n1700 2.2505
R22444 DVDD.n17018 DVDD.n17017 2.2505
R22445 DVDD.n17021 DVDD.n17020 2.2505
R22446 DVDD.n17025 DVDD.n17024 2.2505
R22447 DVDD.n17022 DVDD.n1697 2.2505
R22448 DVDD.n17030 DVDD.n17029 2.2505
R22449 DVDD.n17033 DVDD.n17032 2.2505
R22450 DVDD.n17037 DVDD.n17036 2.2505
R22451 DVDD.n17034 DVDD.n1695 2.2505
R22452 DVDD.n17042 DVDD.n17041 2.2505
R22453 DVDD.n17045 DVDD.n17044 2.2505
R22454 DVDD.n17049 DVDD.n17048 2.2505
R22455 DVDD.n17046 DVDD.n1693 2.2505
R22456 DVDD.n17054 DVDD.n17053 2.2505
R22457 DVDD.n17057 DVDD.n17056 2.2505
R22458 DVDD.n17061 DVDD.n17060 2.2505
R22459 DVDD.n17058 DVDD.n1691 2.2505
R22460 DVDD.n17066 DVDD.n17065 2.2505
R22461 DVDD.n17069 DVDD.n17068 2.2505
R22462 DVDD.n17073 DVDD.n17072 2.2505
R22463 DVDD.n17070 DVDD.n1689 2.2505
R22464 DVDD.n17078 DVDD.n17077 2.2505
R22465 DVDD.n17081 DVDD.n17080 2.2505
R22466 DVDD.n17085 DVDD.n17084 2.2505
R22467 DVDD.n17082 DVDD.n1687 2.2505
R22468 DVDD.n17090 DVDD.n17089 2.2505
R22469 DVDD.n17093 DVDD.n17092 2.2505
R22470 DVDD.n17097 DVDD.n17096 2.2505
R22471 DVDD.n17094 DVDD.n1685 2.2505
R22472 DVDD.n17102 DVDD.n17101 2.2505
R22473 DVDD.n17105 DVDD.n17104 2.2505
R22474 DVDD.n17109 DVDD.n17108 2.2505
R22475 DVDD.n17106 DVDD.n1683 2.2505
R22476 DVDD.n17114 DVDD.n17113 2.2505
R22477 DVDD.n17117 DVDD.n17116 2.2505
R22478 DVDD.n17121 DVDD.n17120 2.2505
R22479 DVDD.n17118 DVDD.n1681 2.2505
R22480 DVDD.n17126 DVDD.n17125 2.2505
R22481 DVDD.n17129 DVDD.n17128 2.2505
R22482 DVDD.n17133 DVDD.n17132 2.2505
R22483 DVDD.n17130 DVDD.n1679 2.2505
R22484 DVDD.n17138 DVDD.n17137 2.2505
R22485 DVDD.n17141 DVDD.n17140 2.2505
R22486 DVDD.n17145 DVDD.n17144 2.2505
R22487 DVDD.n17142 DVDD.n1677 2.2505
R22488 DVDD.n17150 DVDD.n17149 2.2505
R22489 DVDD.n17153 DVDD.n17152 2.2505
R22490 DVDD.n17157 DVDD.n17156 2.2505
R22491 DVDD.n17154 DVDD.n1675 2.2505
R22492 DVDD.n17162 DVDD.n17161 2.2505
R22493 DVDD.n17165 DVDD.n17164 2.2505
R22494 DVDD.n17169 DVDD.n17168 2.2505
R22495 DVDD.n17166 DVDD.n1673 2.2505
R22496 DVDD.n17174 DVDD.n17173 2.2505
R22497 DVDD.n17177 DVDD.n17176 2.2505
R22498 DVDD.n17181 DVDD.n17180 2.2505
R22499 DVDD.n17178 DVDD.n1671 2.2505
R22500 DVDD.n17186 DVDD.n17185 2.2505
R22501 DVDD.n17189 DVDD.n17188 2.2505
R22502 DVDD.n17193 DVDD.n17192 2.2505
R22503 DVDD.n17190 DVDD.n1669 2.2505
R22504 DVDD.n17198 DVDD.n17197 2.2505
R22505 DVDD.n17201 DVDD.n17200 2.2505
R22506 DVDD.n17205 DVDD.n17204 2.2505
R22507 DVDD.n17202 DVDD.n1667 2.2505
R22508 DVDD.n17210 DVDD.n17209 2.2505
R22509 DVDD.n17213 DVDD.n17212 2.2505
R22510 DVDD.n17217 DVDD.n17216 2.2505
R22511 DVDD.n17214 DVDD.n1665 2.2505
R22512 DVDD.n17222 DVDD.n17221 2.2505
R22513 DVDD.n17225 DVDD.n17224 2.2505
R22514 DVDD.n17229 DVDD.n17228 2.2505
R22515 DVDD.n17226 DVDD.n1663 2.2505
R22516 DVDD.n17234 DVDD.n17233 2.2505
R22517 DVDD.n17237 DVDD.n17236 2.2505
R22518 DVDD.n17241 DVDD.n17240 2.2505
R22519 DVDD.n17238 DVDD.n1661 2.2505
R22520 DVDD.n17246 DVDD.n17245 2.2505
R22521 DVDD.n17249 DVDD.n17248 2.2505
R22522 DVDD.n17253 DVDD.n17252 2.2505
R22523 DVDD.n17250 DVDD.n1659 2.2505
R22524 DVDD.n17259 DVDD.n17258 2.2505
R22525 DVDD.n17261 DVDD.n1657 2.2505
R22526 DVDD.n6694 DVDD.n6693 2.2505
R22527 DVDD.n6692 DVDD.n6447 2.2505
R22528 DVDD.n6691 DVDD.n6690 2.2505
R22529 DVDD.n6688 DVDD.n6448 2.2505
R22530 DVDD.n6686 DVDD.n6684 2.2505
R22531 DVDD.n6683 DVDD.n6450 2.2505
R22532 DVDD.n6682 DVDD.n6681 2.2505
R22533 DVDD.n6679 DVDD.n6451 2.2505
R22534 DVDD.n6677 DVDD.n6675 2.2505
R22535 DVDD.n6674 DVDD.n6453 2.2505
R22536 DVDD.n6673 DVDD.n6672 2.2505
R22537 DVDD.n6670 DVDD.n6454 2.2505
R22538 DVDD.n6668 DVDD.n6666 2.2505
R22539 DVDD.n6665 DVDD.n6456 2.2505
R22540 DVDD.n6664 DVDD.n6663 2.2505
R22541 DVDD.n6661 DVDD.n6457 2.2505
R22542 DVDD.n6659 DVDD.n6657 2.2505
R22543 DVDD.n6656 DVDD.n6459 2.2505
R22544 DVDD.n6655 DVDD.n6654 2.2505
R22545 DVDD.n6652 DVDD.n6460 2.2505
R22546 DVDD.n6650 DVDD.n6648 2.2505
R22547 DVDD.n6647 DVDD.n6462 2.2505
R22548 DVDD.n6646 DVDD.n6645 2.2505
R22549 DVDD.n6643 DVDD.n6463 2.2505
R22550 DVDD.n6641 DVDD.n6639 2.2505
R22551 DVDD.n6638 DVDD.n6465 2.2505
R22552 DVDD.n6637 DVDD.n6636 2.2505
R22553 DVDD.n6634 DVDD.n6466 2.2505
R22554 DVDD.n6632 DVDD.n6630 2.2505
R22555 DVDD.n6629 DVDD.n6468 2.2505
R22556 DVDD.n6628 DVDD.n6627 2.2505
R22557 DVDD.n6625 DVDD.n6469 2.2505
R22558 DVDD.n6623 DVDD.n6621 2.2505
R22559 DVDD.n6620 DVDD.n6471 2.2505
R22560 DVDD.n6619 DVDD.n6618 2.2505
R22561 DVDD.n6616 DVDD.n6472 2.2505
R22562 DVDD.n6614 DVDD.n6612 2.2505
R22563 DVDD.n6611 DVDD.n6474 2.2505
R22564 DVDD.n6610 DVDD.n6609 2.2505
R22565 DVDD.n6607 DVDD.n6475 2.2505
R22566 DVDD.n6605 DVDD.n6603 2.2505
R22567 DVDD.n6602 DVDD.n6477 2.2505
R22568 DVDD.n6601 DVDD.n6600 2.2505
R22569 DVDD.n6598 DVDD.n6478 2.2505
R22570 DVDD.n6596 DVDD.n6594 2.2505
R22571 DVDD.n6593 DVDD.n6480 2.2505
R22572 DVDD.n6592 DVDD.n6591 2.2505
R22573 DVDD.n6589 DVDD.n6481 2.2505
R22574 DVDD.n6587 DVDD.n6585 2.2505
R22575 DVDD.n6584 DVDD.n6483 2.2505
R22576 DVDD.n6583 DVDD.n6582 2.2505
R22577 DVDD.n6580 DVDD.n6484 2.2505
R22578 DVDD.n6578 DVDD.n6576 2.2505
R22579 DVDD.n6575 DVDD.n6486 2.2505
R22580 DVDD.n6574 DVDD.n6573 2.2505
R22581 DVDD.n6571 DVDD.n6487 2.2505
R22582 DVDD.n6569 DVDD.n6567 2.2505
R22583 DVDD.n6566 DVDD.n6489 2.2505
R22584 DVDD.n6565 DVDD.n6564 2.2505
R22585 DVDD.n6562 DVDD.n6490 2.2505
R22586 DVDD.n6560 DVDD.n6558 2.2505
R22587 DVDD.n6557 DVDD.n6492 2.2505
R22588 DVDD.n6556 DVDD.n6555 2.2505
R22589 DVDD.n6553 DVDD.n6493 2.2505
R22590 DVDD.n6551 DVDD.n6549 2.2505
R22591 DVDD.n6548 DVDD.n6495 2.2505
R22592 DVDD.n6547 DVDD.n6546 2.2505
R22593 DVDD.n6544 DVDD.n6496 2.2505
R22594 DVDD.n6542 DVDD.n6540 2.2505
R22595 DVDD.n6539 DVDD.n6498 2.2505
R22596 DVDD.n6538 DVDD.n6537 2.2505
R22597 DVDD.n6535 DVDD.n6499 2.2505
R22598 DVDD.n6533 DVDD.n6531 2.2505
R22599 DVDD.n6530 DVDD.n6501 2.2505
R22600 DVDD.n6529 DVDD.n6528 2.2505
R22601 DVDD.n6526 DVDD.n6502 2.2505
R22602 DVDD.n6524 DVDD.n6522 2.2505
R22603 DVDD.n6521 DVDD.n6504 2.2505
R22604 DVDD.n6520 DVDD.n6519 2.2505
R22605 DVDD.n6517 DVDD.n6505 2.2505
R22606 DVDD.n6515 DVDD.n6513 2.2505
R22607 DVDD.n6512 DVDD.n6507 2.2505
R22608 DVDD.n6511 DVDD.n6510 2.2505
R22609 DVDD.n6508 DVDD.n6396 2.2505
R22610 DVDD.n6508 DVDD.n6404 2.2505
R22611 DVDD.n6510 DVDD.n6509 2.2505
R22612 DVDD.n6507 DVDD.n6506 2.2505
R22613 DVDD.n6515 DVDD.n6514 2.2505
R22614 DVDD.n6517 DVDD.n6516 2.2505
R22615 DVDD.n6519 DVDD.n6518 2.2505
R22616 DVDD.n6504 DVDD.n6503 2.2505
R22617 DVDD.n6524 DVDD.n6523 2.2505
R22618 DVDD.n6526 DVDD.n6525 2.2505
R22619 DVDD.n6528 DVDD.n6527 2.2505
R22620 DVDD.n6501 DVDD.n6500 2.2505
R22621 DVDD.n6533 DVDD.n6532 2.2505
R22622 DVDD.n6535 DVDD.n6534 2.2505
R22623 DVDD.n6537 DVDD.n6536 2.2505
R22624 DVDD.n6498 DVDD.n6497 2.2505
R22625 DVDD.n6542 DVDD.n6541 2.2505
R22626 DVDD.n6544 DVDD.n6543 2.2505
R22627 DVDD.n6546 DVDD.n6545 2.2505
R22628 DVDD.n6495 DVDD.n6494 2.2505
R22629 DVDD.n6551 DVDD.n6550 2.2505
R22630 DVDD.n6553 DVDD.n6552 2.2505
R22631 DVDD.n6555 DVDD.n6554 2.2505
R22632 DVDD.n6492 DVDD.n6491 2.2505
R22633 DVDD.n6560 DVDD.n6559 2.2505
R22634 DVDD.n6562 DVDD.n6561 2.2505
R22635 DVDD.n6564 DVDD.n6563 2.2505
R22636 DVDD.n6489 DVDD.n6488 2.2505
R22637 DVDD.n6569 DVDD.n6568 2.2505
R22638 DVDD.n6571 DVDD.n6570 2.2505
R22639 DVDD.n6573 DVDD.n6572 2.2505
R22640 DVDD.n6486 DVDD.n6485 2.2505
R22641 DVDD.n6578 DVDD.n6577 2.2505
R22642 DVDD.n6580 DVDD.n6579 2.2505
R22643 DVDD.n6582 DVDD.n6581 2.2505
R22644 DVDD.n6483 DVDD.n6482 2.2505
R22645 DVDD.n6587 DVDD.n6586 2.2505
R22646 DVDD.n6589 DVDD.n6588 2.2505
R22647 DVDD.n6591 DVDD.n6590 2.2505
R22648 DVDD.n6480 DVDD.n6479 2.2505
R22649 DVDD.n6596 DVDD.n6595 2.2505
R22650 DVDD.n6598 DVDD.n6597 2.2505
R22651 DVDD.n6600 DVDD.n6599 2.2505
R22652 DVDD.n6477 DVDD.n6476 2.2505
R22653 DVDD.n6605 DVDD.n6604 2.2505
R22654 DVDD.n6607 DVDD.n6606 2.2505
R22655 DVDD.n6609 DVDD.n6608 2.2505
R22656 DVDD.n6474 DVDD.n6473 2.2505
R22657 DVDD.n6614 DVDD.n6613 2.2505
R22658 DVDD.n6616 DVDD.n6615 2.2505
R22659 DVDD.n6618 DVDD.n6617 2.2505
R22660 DVDD.n6471 DVDD.n6470 2.2505
R22661 DVDD.n6623 DVDD.n6622 2.2505
R22662 DVDD.n6625 DVDD.n6624 2.2505
R22663 DVDD.n6627 DVDD.n6626 2.2505
R22664 DVDD.n6468 DVDD.n6467 2.2505
R22665 DVDD.n6632 DVDD.n6631 2.2505
R22666 DVDD.n6634 DVDD.n6633 2.2505
R22667 DVDD.n6636 DVDD.n6635 2.2505
R22668 DVDD.n6465 DVDD.n6464 2.2505
R22669 DVDD.n6641 DVDD.n6640 2.2505
R22670 DVDD.n6643 DVDD.n6642 2.2505
R22671 DVDD.n6645 DVDD.n6644 2.2505
R22672 DVDD.n6462 DVDD.n6461 2.2505
R22673 DVDD.n6650 DVDD.n6649 2.2505
R22674 DVDD.n6652 DVDD.n6651 2.2505
R22675 DVDD.n6654 DVDD.n6653 2.2505
R22676 DVDD.n6459 DVDD.n6458 2.2505
R22677 DVDD.n6659 DVDD.n6658 2.2505
R22678 DVDD.n6661 DVDD.n6660 2.2505
R22679 DVDD.n6663 DVDD.n6662 2.2505
R22680 DVDD.n6456 DVDD.n6455 2.2505
R22681 DVDD.n6668 DVDD.n6667 2.2505
R22682 DVDD.n6670 DVDD.n6669 2.2505
R22683 DVDD.n6672 DVDD.n6671 2.2505
R22684 DVDD.n6453 DVDD.n6452 2.2505
R22685 DVDD.n6677 DVDD.n6676 2.2505
R22686 DVDD.n6679 DVDD.n6678 2.2505
R22687 DVDD.n6681 DVDD.n6680 2.2505
R22688 DVDD.n6450 DVDD.n6449 2.2505
R22689 DVDD.n6686 DVDD.n6685 2.2505
R22690 DVDD.n6688 DVDD.n6687 2.2505
R22691 DVDD.n6690 DVDD.n6689 2.2505
R22692 DVDD.n6447 DVDD.n6446 2.2505
R22693 DVDD.n6695 DVDD.n6694 2.2505
R22694 DVDD.n15123 DVDD.n15122 2.2505
R22695 DVDD.n5935 DVDD.n5933 2.2505
R22696 DVDD.n6338 DVDD.n6000 2.2505
R22697 DVDD.n6341 DVDD.n6043 2.2505
R22698 DVDD.n6403 DVDD.n6346 2.2505
R22699 DVDD.n15103 DVDD.n15102 2.2505
R22700 DVDD.n7047 DVDD.n6391 2.2505
R22701 DVDD.n7046 DVDD.n6707 2.2505
R22702 DVDD.n7045 DVDD.n6749 2.2505
R22703 DVDD.n7054 DVDD.n6794 2.2505
R22704 DVDD.n15080 DVDD.n15079 2.2505
R22705 DVDD.n15069 DVDD.n15068 2.2505
R22706 DVDD.n7411 DVDD.n7405 2.2505
R22707 DVDD.n15062 DVDD.n15061 2.2505
R22708 DVDD.n7667 DVDD.n7458 2.2505
R22709 DVDD.n7669 DVDD.n7569 2.2505
R22710 DVDD.n7668 DVDD.n7611 2.2505
R22711 DVDD.n7664 DVDD.n7657 2.2505
R22712 DVDD.n9559 DVDD.n7676 2.2505
R22713 DVDD.n14851 DVDD.n14850 2.2505
R22714 DVDD.n8031 DVDD.n8030 2.2505
R22715 DVDD.n8033 DVDD.n7688 2.2505
R22716 DVDD.n8032 DVDD.n7730 2.2505
R22717 DVDD.n8026 DVDD.n7775 2.2505
R22718 DVDD.n8145 DVDD.n8144 2.2505
R22719 DVDD.n14827 DVDD.n14826 2.2505
R22720 DVDD.n8154 DVDD.n8043 2.2505
R22721 DVDD.n14568 DVDD.n14567 2.2505
R22722 DVDD.n14561 DVDD.n14560 2.2505
R22723 DVDD.n8599 DVDD.n8161 2.2505
R22724 DVDD.n8602 DVDD.n8601 2.2505
R22725 DVDD.n14302 DVDD.n14301 2.2505
R22726 DVDD.n10232 DVDD.n8261 2.2505
R22727 DVDD.n14295 DVDD.n14294 2.2505
R22728 DVDD.n10584 DVDD.n10583 2.2505
R22729 DVDD.n10586 DVDD.n10241 2.2505
R22730 DVDD.n10585 DVDD.n10283 2.2505
R22731 DVDD.n10579 DVDD.n10328 2.2505
R22732 DVDD.n10692 DVDD.n10691 2.2505
R22733 DVDD.n14271 DVDD.n14270 2.2505
R22734 DVDD.n11051 DVDD.n10596 2.2505
R22735 DVDD.n11054 DVDD.n11053 2.2505
R22736 DVDD.n14012 DVDD.n14011 2.2505
R22737 DVDD.n11215 DVDD.n10713 2.2505
R22738 DVDD.n14005 DVDD.n14004 2.2505
R22739 DVDD.n11572 DVDD.n11568 2.2505
R22740 DVDD.n11574 DVDD.n11573 2.2505
R22741 DVDD.n11575 DVDD.n11233 2.2505
R22742 DVDD.n13789 DVDD.n11276 2.2505
R22743 DVDD.n13788 DVDD.n13787 2.2505
R22744 DVDD.n11588 DVDD.n11579 2.2505
R22745 DVDD.n13767 DVDD.n11631 2.2505
R22746 DVDD.n13766 DVDD.n13765 2.2505
R22747 DVDD.n11937 DVDD.n11924 2.2505
R22748 DVDD.n13754 DVDD.n13753 2.2505
R22749 DVDD.n12332 DVDD.n11941 2.2505
R22750 DVDD.n13746 DVDD.n13745 2.2505
R22751 DVDD.n12388 DVDD.n12286 2.2505
R22752 DVDD.n12726 DVDD.n12390 2.2505
R22753 DVDD.n12729 DVDD.n12432 2.2505
R22754 DVDD.n12736 DVDD.n12734 2.2505
R22755 DVDD.n13475 DVDD.n13474 2.2505
R22756 DVDD.n12920 DVDD.n12783 2.2505
R22757 DVDD.n12922 DVDD.n12921 2.2505
R22758 DVDD.n13259 DVDD.n13258 2.2505
R22759 DVDD.n13266 DVDD.n13265 2.2505
R22760 DVDD.n13268 DVDD.n2163 2.2505
R22761 DVDD.n16706 DVDD.n16705 2.2505
R22762 DVDD.n2157 DVDD.n1821 2.2505
R22763 DVDD.n16714 DVDD.n16713 2.2505
R22764 DVDD.n16728 DVDD.n16727 2.2505
R22765 DVDD.n1812 DVDD.n1806 2.2505
R22766 DVDD.n16735 DVDD.n16734 2.2505
R22767 DVDD.n16996 DVDD.n16995 2.2505
R22768 DVDD.n1707 DVDD.n1706 2.2505
R22769 DVDD.n17003 DVDD.n17002 2.2505
R22770 DVDD.n17264 DVDD.n17263 2.2505
R22771 DVDD.n1655 DVDD.n1606 2.2505
R22772 DVDD.n17271 DVDD.n17270 2.2505
R22773 DVDD.n17282 DVDD.n17281 2.2505
R22774 DVDD.n1263 DVDD.n1257 2.2505
R22775 DVDD.n17289 DVDD.n17288 2.2505
R22776 DVDD.n17301 DVDD.n17300 2.2505
R22777 DVDD.n908 DVDD.n906 2.2505
R22778 DVDD.n17717 DVDD.n17716 2.2505
R22779 DVDD.n15110 DVDD.n6337 2.2505
R22780 DVDD.n6336 DVDD.n6047 2.2505
R22781 DVDD.n6335 DVDD.n6334 2.2505
R22782 DVDD.n6049 DVDD.n6048 2.2505
R22783 DVDD.n6154 DVDD.n6153 2.2505
R22784 DVDD.n6155 DVDD.n6151 2.2505
R22785 DVDD.n6158 DVDD.n6156 2.2505
R22786 DVDD.n6160 DVDD.n6149 2.2505
R22787 DVDD.n6163 DVDD.n6162 2.2505
R22788 DVDD.n6164 DVDD.n6148 2.2505
R22789 DVDD.n6167 DVDD.n6165 2.2505
R22790 DVDD.n6169 DVDD.n6146 2.2505
R22791 DVDD.n6172 DVDD.n6171 2.2505
R22792 DVDD.n6173 DVDD.n6145 2.2505
R22793 DVDD.n6176 DVDD.n6174 2.2505
R22794 DVDD.n6178 DVDD.n6143 2.2505
R22795 DVDD.n6181 DVDD.n6180 2.2505
R22796 DVDD.n6182 DVDD.n6142 2.2505
R22797 DVDD.n6185 DVDD.n6183 2.2505
R22798 DVDD.n6187 DVDD.n6140 2.2505
R22799 DVDD.n6190 DVDD.n6189 2.2505
R22800 DVDD.n6191 DVDD.n6139 2.2505
R22801 DVDD.n6194 DVDD.n6192 2.2505
R22802 DVDD.n6196 DVDD.n6137 2.2505
R22803 DVDD.n6199 DVDD.n6198 2.2505
R22804 DVDD.n6200 DVDD.n6136 2.2505
R22805 DVDD.n6203 DVDD.n6201 2.2505
R22806 DVDD.n6205 DVDD.n6134 2.2505
R22807 DVDD.n6208 DVDD.n6207 2.2505
R22808 DVDD.n6209 DVDD.n6133 2.2505
R22809 DVDD.n6212 DVDD.n6210 2.2505
R22810 DVDD.n6214 DVDD.n6131 2.2505
R22811 DVDD.n6217 DVDD.n6216 2.2505
R22812 DVDD.n6218 DVDD.n6130 2.2505
R22813 DVDD.n6221 DVDD.n6219 2.2505
R22814 DVDD.n6223 DVDD.n6128 2.2505
R22815 DVDD.n6226 DVDD.n6225 2.2505
R22816 DVDD.n6227 DVDD.n6127 2.2505
R22817 DVDD.n6230 DVDD.n6228 2.2505
R22818 DVDD.n6232 DVDD.n6125 2.2505
R22819 DVDD.n6235 DVDD.n6234 2.2505
R22820 DVDD.n6236 DVDD.n6124 2.2505
R22821 DVDD.n6239 DVDD.n6237 2.2505
R22822 DVDD.n6241 DVDD.n6122 2.2505
R22823 DVDD.n6244 DVDD.n6243 2.2505
R22824 DVDD.n6245 DVDD.n6121 2.2505
R22825 DVDD.n6248 DVDD.n6246 2.2505
R22826 DVDD.n6250 DVDD.n6119 2.2505
R22827 DVDD.n6253 DVDD.n6252 2.2505
R22828 DVDD.n6254 DVDD.n6118 2.2505
R22829 DVDD.n6257 DVDD.n6255 2.2505
R22830 DVDD.n6259 DVDD.n6116 2.2505
R22831 DVDD.n6262 DVDD.n6261 2.2505
R22832 DVDD.n6263 DVDD.n6115 2.2505
R22833 DVDD.n6266 DVDD.n6264 2.2505
R22834 DVDD.n6268 DVDD.n6113 2.2505
R22835 DVDD.n6271 DVDD.n6270 2.2505
R22836 DVDD.n6272 DVDD.n6112 2.2505
R22837 DVDD.n6275 DVDD.n6273 2.2505
R22838 DVDD.n6277 DVDD.n6110 2.2505
R22839 DVDD.n6280 DVDD.n6279 2.2505
R22840 DVDD.n6281 DVDD.n6109 2.2505
R22841 DVDD.n6284 DVDD.n6282 2.2505
R22842 DVDD.n6286 DVDD.n6107 2.2505
R22843 DVDD.n6289 DVDD.n6288 2.2505
R22844 DVDD.n6290 DVDD.n6106 2.2505
R22845 DVDD.n6293 DVDD.n6291 2.2505
R22846 DVDD.n6295 DVDD.n6104 2.2505
R22847 DVDD.n6298 DVDD.n6297 2.2505
R22848 DVDD.n6299 DVDD.n6103 2.2505
R22849 DVDD.n6302 DVDD.n6300 2.2505
R22850 DVDD.n6304 DVDD.n6101 2.2505
R22851 DVDD.n6307 DVDD.n6306 2.2505
R22852 DVDD.n6308 DVDD.n6100 2.2505
R22853 DVDD.n6311 DVDD.n6309 2.2505
R22854 DVDD.n6313 DVDD.n6098 2.2505
R22855 DVDD.n6316 DVDD.n6315 2.2505
R22856 DVDD.n6317 DVDD.n6097 2.2505
R22857 DVDD.n6320 DVDD.n6318 2.2505
R22858 DVDD.n6322 DVDD.n6095 2.2505
R22859 DVDD.n6325 DVDD.n6324 2.2505
R22860 DVDD.n6326 DVDD.n6093 2.2505
R22861 DVDD.n6328 DVDD.n6327 2.2505
R22862 DVDD.n6094 DVDD.n6091 2.2505
R22863 DVDD.n6091 DVDD.n6042 2.2505
R22864 DVDD.n6329 DVDD.n6328 2.2505
R22865 DVDD.n6093 DVDD.n6092 2.2505
R22866 DVDD.n6324 DVDD.n6323 2.2505
R22867 DVDD.n6322 DVDD.n6321 2.2505
R22868 DVDD.n6320 DVDD.n6319 2.2505
R22869 DVDD.n6097 DVDD.n6096 2.2505
R22870 DVDD.n6315 DVDD.n6314 2.2505
R22871 DVDD.n6313 DVDD.n6312 2.2505
R22872 DVDD.n6311 DVDD.n6310 2.2505
R22873 DVDD.n6100 DVDD.n6099 2.2505
R22874 DVDD.n6306 DVDD.n6305 2.2505
R22875 DVDD.n6304 DVDD.n6303 2.2505
R22876 DVDD.n6302 DVDD.n6301 2.2505
R22877 DVDD.n6103 DVDD.n6102 2.2505
R22878 DVDD.n6297 DVDD.n6296 2.2505
R22879 DVDD.n6295 DVDD.n6294 2.2505
R22880 DVDD.n6293 DVDD.n6292 2.2505
R22881 DVDD.n6106 DVDD.n6105 2.2505
R22882 DVDD.n6288 DVDD.n6287 2.2505
R22883 DVDD.n6286 DVDD.n6285 2.2505
R22884 DVDD.n6284 DVDD.n6283 2.2505
R22885 DVDD.n6109 DVDD.n6108 2.2505
R22886 DVDD.n6279 DVDD.n6278 2.2505
R22887 DVDD.n6277 DVDD.n6276 2.2505
R22888 DVDD.n6275 DVDD.n6274 2.2505
R22889 DVDD.n6112 DVDD.n6111 2.2505
R22890 DVDD.n6270 DVDD.n6269 2.2505
R22891 DVDD.n6268 DVDD.n6267 2.2505
R22892 DVDD.n6266 DVDD.n6265 2.2505
R22893 DVDD.n6115 DVDD.n6114 2.2505
R22894 DVDD.n6261 DVDD.n6260 2.2505
R22895 DVDD.n6259 DVDD.n6258 2.2505
R22896 DVDD.n6257 DVDD.n6256 2.2505
R22897 DVDD.n6118 DVDD.n6117 2.2505
R22898 DVDD.n6252 DVDD.n6251 2.2505
R22899 DVDD.n6250 DVDD.n6249 2.2505
R22900 DVDD.n6248 DVDD.n6247 2.2505
R22901 DVDD.n6121 DVDD.n6120 2.2505
R22902 DVDD.n6243 DVDD.n6242 2.2505
R22903 DVDD.n6241 DVDD.n6240 2.2505
R22904 DVDD.n6239 DVDD.n6238 2.2505
R22905 DVDD.n6124 DVDD.n6123 2.2505
R22906 DVDD.n6234 DVDD.n6233 2.2505
R22907 DVDD.n6232 DVDD.n6231 2.2505
R22908 DVDD.n6230 DVDD.n6229 2.2505
R22909 DVDD.n6127 DVDD.n6126 2.2505
R22910 DVDD.n6225 DVDD.n6224 2.2505
R22911 DVDD.n6223 DVDD.n6222 2.2505
R22912 DVDD.n6221 DVDD.n6220 2.2505
R22913 DVDD.n6130 DVDD.n6129 2.2505
R22914 DVDD.n6216 DVDD.n6215 2.2505
R22915 DVDD.n6214 DVDD.n6213 2.2505
R22916 DVDD.n6212 DVDD.n6211 2.2505
R22917 DVDD.n6133 DVDD.n6132 2.2505
R22918 DVDD.n6207 DVDD.n6206 2.2505
R22919 DVDD.n6205 DVDD.n6204 2.2505
R22920 DVDD.n6203 DVDD.n6202 2.2505
R22921 DVDD.n6136 DVDD.n6135 2.2505
R22922 DVDD.n6198 DVDD.n6197 2.2505
R22923 DVDD.n6196 DVDD.n6195 2.2505
R22924 DVDD.n6194 DVDD.n6193 2.2505
R22925 DVDD.n6139 DVDD.n6138 2.2505
R22926 DVDD.n6189 DVDD.n6188 2.2505
R22927 DVDD.n6187 DVDD.n6186 2.2505
R22928 DVDD.n6185 DVDD.n6184 2.2505
R22929 DVDD.n6142 DVDD.n6141 2.2505
R22930 DVDD.n6180 DVDD.n6179 2.2505
R22931 DVDD.n6178 DVDD.n6177 2.2505
R22932 DVDD.n6176 DVDD.n6175 2.2505
R22933 DVDD.n6145 DVDD.n6144 2.2505
R22934 DVDD.n6171 DVDD.n6170 2.2505
R22935 DVDD.n6169 DVDD.n6168 2.2505
R22936 DVDD.n6167 DVDD.n6166 2.2505
R22937 DVDD.n6148 DVDD.n6147 2.2505
R22938 DVDD.n6162 DVDD.n6161 2.2505
R22939 DVDD.n6160 DVDD.n6159 2.2505
R22940 DVDD.n6158 DVDD.n6157 2.2505
R22941 DVDD.n6151 DVDD.n6150 2.2505
R22942 DVDD.n6153 DVDD.n6152 2.2505
R22943 DVDD.n6050 DVDD.n6049 2.2505
R22944 DVDD.n6334 DVDD.n6333 2.2505
R22945 DVDD.n6047 DVDD.n6046 2.2505
R22946 DVDD.n15111 DVDD.n15110 2.2505
R22947 DVDD.n1358 DVDD.n1357 2.2505
R22948 DVDD.n1359 DVDD.n1355 2.2505
R22949 DVDD.n1364 DVDD.n1360 2.2505
R22950 DVDD.n1365 DVDD.n1354 2.2505
R22951 DVDD.n1370 DVDD.n1369 2.2505
R22952 DVDD.n1371 DVDD.n1353 2.2505
R22953 DVDD.n1376 DVDD.n1372 2.2505
R22954 DVDD.n1377 DVDD.n1352 2.2505
R22955 DVDD.n1382 DVDD.n1381 2.2505
R22956 DVDD.n1383 DVDD.n1351 2.2505
R22957 DVDD.n1388 DVDD.n1384 2.2505
R22958 DVDD.n1389 DVDD.n1350 2.2505
R22959 DVDD.n1394 DVDD.n1393 2.2505
R22960 DVDD.n1395 DVDD.n1349 2.2505
R22961 DVDD.n1400 DVDD.n1396 2.2505
R22962 DVDD.n1401 DVDD.n1348 2.2505
R22963 DVDD.n1406 DVDD.n1405 2.2505
R22964 DVDD.n1407 DVDD.n1347 2.2505
R22965 DVDD.n1412 DVDD.n1408 2.2505
R22966 DVDD.n1413 DVDD.n1346 2.2505
R22967 DVDD.n1418 DVDD.n1417 2.2505
R22968 DVDD.n1419 DVDD.n1345 2.2505
R22969 DVDD.n1424 DVDD.n1420 2.2505
R22970 DVDD.n1425 DVDD.n1344 2.2505
R22971 DVDD.n1430 DVDD.n1429 2.2505
R22972 DVDD.n1431 DVDD.n1343 2.2505
R22973 DVDD.n1436 DVDD.n1432 2.2505
R22974 DVDD.n1437 DVDD.n1342 2.2505
R22975 DVDD.n1442 DVDD.n1441 2.2505
R22976 DVDD.n1443 DVDD.n1341 2.2505
R22977 DVDD.n1448 DVDD.n1444 2.2505
R22978 DVDD.n1449 DVDD.n1340 2.2505
R22979 DVDD.n1454 DVDD.n1453 2.2505
R22980 DVDD.n1455 DVDD.n1339 2.2505
R22981 DVDD.n1460 DVDD.n1456 2.2505
R22982 DVDD.n1461 DVDD.n1338 2.2505
R22983 DVDD.n1466 DVDD.n1465 2.2505
R22984 DVDD.n1467 DVDD.n1337 2.2505
R22985 DVDD.n1472 DVDD.n1468 2.2505
R22986 DVDD.n1473 DVDD.n1336 2.2505
R22987 DVDD.n1478 DVDD.n1477 2.2505
R22988 DVDD.n1479 DVDD.n1335 2.2505
R22989 DVDD.n1484 DVDD.n1480 2.2505
R22990 DVDD.n1485 DVDD.n1334 2.2505
R22991 DVDD.n1490 DVDD.n1489 2.2505
R22992 DVDD.n1491 DVDD.n1333 2.2505
R22993 DVDD.n1496 DVDD.n1492 2.2505
R22994 DVDD.n1497 DVDD.n1332 2.2505
R22995 DVDD.n1502 DVDD.n1501 2.2505
R22996 DVDD.n1503 DVDD.n1331 2.2505
R22997 DVDD.n1508 DVDD.n1504 2.2505
R22998 DVDD.n1509 DVDD.n1330 2.2505
R22999 DVDD.n1514 DVDD.n1513 2.2505
R23000 DVDD.n1515 DVDD.n1329 2.2505
R23001 DVDD.n1520 DVDD.n1516 2.2505
R23002 DVDD.n1521 DVDD.n1328 2.2505
R23003 DVDD.n1526 DVDD.n1525 2.2505
R23004 DVDD.n1527 DVDD.n1327 2.2505
R23005 DVDD.n1532 DVDD.n1528 2.2505
R23006 DVDD.n1533 DVDD.n1326 2.2505
R23007 DVDD.n1538 DVDD.n1537 2.2505
R23008 DVDD.n1539 DVDD.n1325 2.2505
R23009 DVDD.n1544 DVDD.n1540 2.2505
R23010 DVDD.n1545 DVDD.n1324 2.2505
R23011 DVDD.n1550 DVDD.n1549 2.2505
R23012 DVDD.n1551 DVDD.n1323 2.2505
R23013 DVDD.n1556 DVDD.n1552 2.2505
R23014 DVDD.n1557 DVDD.n1322 2.2505
R23015 DVDD.n1562 DVDD.n1561 2.2505
R23016 DVDD.n1563 DVDD.n1321 2.2505
R23017 DVDD.n1568 DVDD.n1564 2.2505
R23018 DVDD.n1569 DVDD.n1320 2.2505
R23019 DVDD.n1574 DVDD.n1573 2.2505
R23020 DVDD.n1575 DVDD.n1319 2.2505
R23021 DVDD.n1580 DVDD.n1576 2.2505
R23022 DVDD.n1581 DVDD.n1318 2.2505
R23023 DVDD.n1586 DVDD.n1585 2.2505
R23024 DVDD.n1587 DVDD.n1317 2.2505
R23025 DVDD.n1592 DVDD.n1588 2.2505
R23026 DVDD.n1593 DVDD.n1316 2.2505
R23027 DVDD.n1598 DVDD.n1597 2.2505
R23028 DVDD.n1599 DVDD.n1315 2.2505
R23029 DVDD.n1601 DVDD.n1600 2.2505
R23030 DVDD.n1602 DVDD.n1267 2.2505
R23031 DVDD.n1603 DVDD.n1602 2.2505
R23032 DVDD.n1601 DVDD.n1312 2.2505
R23033 DVDD.n1315 DVDD.n1314 2.2505
R23034 DVDD.n1597 DVDD.n1596 2.2505
R23035 DVDD.n1594 DVDD.n1593 2.2505
R23036 DVDD.n1592 DVDD.n1591 2.2505
R23037 DVDD.n1589 DVDD.n1317 2.2505
R23038 DVDD.n1585 DVDD.n1584 2.2505
R23039 DVDD.n1582 DVDD.n1581 2.2505
R23040 DVDD.n1580 DVDD.n1579 2.2505
R23041 DVDD.n1577 DVDD.n1319 2.2505
R23042 DVDD.n1573 DVDD.n1572 2.2505
R23043 DVDD.n1570 DVDD.n1569 2.2505
R23044 DVDD.n1568 DVDD.n1567 2.2505
R23045 DVDD.n1565 DVDD.n1321 2.2505
R23046 DVDD.n1561 DVDD.n1560 2.2505
R23047 DVDD.n1558 DVDD.n1557 2.2505
R23048 DVDD.n1556 DVDD.n1555 2.2505
R23049 DVDD.n1553 DVDD.n1323 2.2505
R23050 DVDD.n1549 DVDD.n1548 2.2505
R23051 DVDD.n1546 DVDD.n1545 2.2505
R23052 DVDD.n1544 DVDD.n1543 2.2505
R23053 DVDD.n1541 DVDD.n1325 2.2505
R23054 DVDD.n1537 DVDD.n1536 2.2505
R23055 DVDD.n1534 DVDD.n1533 2.2505
R23056 DVDD.n1532 DVDD.n1531 2.2505
R23057 DVDD.n1529 DVDD.n1327 2.2505
R23058 DVDD.n1525 DVDD.n1524 2.2505
R23059 DVDD.n1522 DVDD.n1521 2.2505
R23060 DVDD.n1520 DVDD.n1519 2.2505
R23061 DVDD.n1517 DVDD.n1329 2.2505
R23062 DVDD.n1513 DVDD.n1512 2.2505
R23063 DVDD.n1510 DVDD.n1509 2.2505
R23064 DVDD.n1508 DVDD.n1507 2.2505
R23065 DVDD.n1505 DVDD.n1331 2.2505
R23066 DVDD.n1501 DVDD.n1500 2.2505
R23067 DVDD.n1498 DVDD.n1497 2.2505
R23068 DVDD.n1496 DVDD.n1495 2.2505
R23069 DVDD.n1493 DVDD.n1333 2.2505
R23070 DVDD.n1489 DVDD.n1488 2.2505
R23071 DVDD.n1486 DVDD.n1485 2.2505
R23072 DVDD.n1484 DVDD.n1483 2.2505
R23073 DVDD.n1481 DVDD.n1335 2.2505
R23074 DVDD.n1477 DVDD.n1476 2.2505
R23075 DVDD.n1474 DVDD.n1473 2.2505
R23076 DVDD.n1472 DVDD.n1471 2.2505
R23077 DVDD.n1469 DVDD.n1337 2.2505
R23078 DVDD.n1465 DVDD.n1464 2.2505
R23079 DVDD.n1462 DVDD.n1461 2.2505
R23080 DVDD.n1460 DVDD.n1459 2.2505
R23081 DVDD.n1457 DVDD.n1339 2.2505
R23082 DVDD.n1453 DVDD.n1452 2.2505
R23083 DVDD.n1450 DVDD.n1449 2.2505
R23084 DVDD.n1448 DVDD.n1447 2.2505
R23085 DVDD.n1445 DVDD.n1341 2.2505
R23086 DVDD.n1441 DVDD.n1440 2.2505
R23087 DVDD.n1438 DVDD.n1437 2.2505
R23088 DVDD.n1436 DVDD.n1435 2.2505
R23089 DVDD.n1433 DVDD.n1343 2.2505
R23090 DVDD.n1429 DVDD.n1428 2.2505
R23091 DVDD.n1426 DVDD.n1425 2.2505
R23092 DVDD.n1424 DVDD.n1423 2.2505
R23093 DVDD.n1421 DVDD.n1345 2.2505
R23094 DVDD.n1417 DVDD.n1416 2.2505
R23095 DVDD.n1414 DVDD.n1413 2.2505
R23096 DVDD.n1412 DVDD.n1411 2.2505
R23097 DVDD.n1409 DVDD.n1347 2.2505
R23098 DVDD.n1405 DVDD.n1404 2.2505
R23099 DVDD.n1402 DVDD.n1401 2.2505
R23100 DVDD.n1400 DVDD.n1399 2.2505
R23101 DVDD.n1397 DVDD.n1349 2.2505
R23102 DVDD.n1393 DVDD.n1392 2.2505
R23103 DVDD.n1390 DVDD.n1389 2.2505
R23104 DVDD.n1388 DVDD.n1387 2.2505
R23105 DVDD.n1385 DVDD.n1351 2.2505
R23106 DVDD.n1381 DVDD.n1380 2.2505
R23107 DVDD.n1378 DVDD.n1377 2.2505
R23108 DVDD.n1376 DVDD.n1375 2.2505
R23109 DVDD.n1373 DVDD.n1353 2.2505
R23110 DVDD.n1369 DVDD.n1368 2.2505
R23111 DVDD.n1366 DVDD.n1365 2.2505
R23112 DVDD.n1364 DVDD.n1363 2.2505
R23113 DVDD.n1361 DVDD.n1355 2.2505
R23114 DVDD.n1357 DVDD.n1356 2.2505
R23115 DVDD.n15124 DVDD.n15123 2.2505
R23116 DVDD.n5933 DVDD.n5932 2.2505
R23117 DVDD.n6339 DVDD.n6338 2.2505
R23118 DVDD.n15108 DVDD.n6341 2.2505
R23119 DVDD.n6346 DVDD.n6340 2.2505
R23120 DVDD.n15104 DVDD.n15103 2.2505
R23121 DVDD.n7048 DVDD.n7047 2.2505
R23122 DVDD.n7046 DVDD.n7043 2.2505
R23123 DVDD.n15085 DVDD.n7045 2.2505
R23124 DVDD.n7054 DVDD.n7044 2.2505
R23125 DVDD.n15081 DVDD.n15080 2.2505
R23126 DVDD.n15068 DVDD.n15067 2.2505
R23127 DVDD.n7406 DVDD.n7405 2.2505
R23128 DVDD.n15063 DVDD.n15062 2.2505
R23129 DVDD.n7667 DVDD.n7666 2.2505
R23130 DVDD.n7670 DVDD.n7669 2.2505
R23131 DVDD.n7668 DVDD.n7662 2.2505
R23132 DVDD.n14856 DVDD.n7664 2.2505
R23133 DVDD.n7676 DVDD.n7663 2.2505
R23134 DVDD.n14852 DVDD.n14851 2.2505
R23135 DVDD.n8031 DVDD.n8028 2.2505
R23136 DVDD.n8034 DVDD.n8033 2.2505
R23137 DVDD.n8032 DVDD.n8024 2.2505
R23138 DVDD.n14833 DVDD.n8026 2.2505
R23139 DVDD.n8144 DVDD.n8025 2.2505
R23140 DVDD.n14828 DVDD.n14827 2.2505
R23141 DVDD.n8043 DVDD.n8041 2.2505
R23142 DVDD.n14567 DVDD.n14566 2.2505
R23143 DVDD.n14562 DVDD.n14561 2.2505
R23144 DVDD.n8161 DVDD.n8160 2.2505
R23145 DVDD.n8603 DVDD.n8602 2.2505
R23146 DVDD.n14301 DVDD.n14300 2.2505
R23147 DVDD.n8263 DVDD.n8261 2.2505
R23148 DVDD.n14296 DVDD.n14295 2.2505
R23149 DVDD.n10584 DVDD.n10581 2.2505
R23150 DVDD.n10587 DVDD.n10586 2.2505
R23151 DVDD.n10585 DVDD.n10577 2.2505
R23152 DVDD.n14277 DVDD.n10579 2.2505
R23153 DVDD.n10691 DVDD.n10578 2.2505
R23154 DVDD.n14272 DVDD.n14271 2.2505
R23155 DVDD.n10596 DVDD.n10594 2.2505
R23156 DVDD.n11055 DVDD.n11054 2.2505
R23157 DVDD.n14011 DVDD.n14010 2.2505
R23158 DVDD.n10715 DVDD.n10713 2.2505
R23159 DVDD.n14006 DVDD.n14005 2.2505
R23160 DVDD.n11572 DVDD.n11571 2.2505
R23161 DVDD.n11574 DVDD.n11567 2.2505
R23162 DVDD.n11576 DVDD.n11575 2.2505
R23163 DVDD.n13790 DVDD.n13789 2.2505
R23164 DVDD.n13788 DVDD.n11578 2.2505
R23165 DVDD.n11921 DVDD.n11579 2.2505
R23166 DVDD.n13768 DVDD.n13767 2.2505
R23167 DVDD.n13766 DVDD.n11923 2.2505
R23168 DVDD.n12278 DVDD.n11924 2.2505
R23169 DVDD.n13753 DVDD.n13752 2.2505
R23170 DVDD.n11943 DVDD.n11941 2.2505
R23171 DVDD.n13747 DVDD.n13746 2.2505
R23172 DVDD.n12286 DVDD.n12284 2.2505
R23173 DVDD.n12727 DVDD.n12726 2.2505
R23174 DVDD.n13480 DVDD.n12729 2.2505
R23175 DVDD.n12734 DVDD.n12728 2.2505
R23176 DVDD.n13476 DVDD.n13475 2.2505
R23177 DVDD.n12920 DVDD.n12919 2.2505
R23178 DVDD.n12922 DVDD.n12917 2.2505
R23179 DVDD.n13260 DVDD.n13259 2.2505
R23180 DVDD.n13265 DVDD.n13264 2.2505
R23181 DVDD.n2163 DVDD.n2161 2.2505
R23182 DVDD.n16707 DVDD.n16706 2.2505
R23183 DVDD.n2158 DVDD.n2157 2.2505
R23184 DVDD.n16713 DVDD.n16712 2.2505
R23185 DVDD.n16729 DVDD.n16728 2.2505
R23186 DVDD.n1807 DVDD.n1806 2.2505
R23187 DVDD.n16734 DVDD.n16733 2.2505
R23188 DVDD.n16997 DVDD.n16996 2.2505
R23189 DVDD.n1708 DVDD.n1707 2.2505
R23190 DVDD.n17002 DVDD.n17001 2.2505
R23191 DVDD.n17265 DVDD.n17264 2.2505
R23192 DVDD.n1607 DVDD.n1606 2.2505
R23193 DVDD.n17270 DVDD.n17269 2.2505
R23194 DVDD.n17283 DVDD.n17282 2.2505
R23195 DVDD.n1258 DVDD.n1257 2.2505
R23196 DVDD.n17288 DVDD.n17287 2.2505
R23197 DVDD.n17302 DVDD.n17301 2.2505
R23198 DVDD.n910 DVDD.n908 2.2505
R23199 DVDD.n17716 DVDD.n17715 2.2505
R23200 DVDD.n965 DVDD.n963 2.2505
R23201 DVDD.n1254 DVDD.n1253 2.2505
R23202 DVDD.n967 DVDD.n966 2.2505
R23203 DVDD.n1249 DVDD.n1248 2.2505
R23204 DVDD.n1246 DVDD.n1245 2.2505
R23205 DVDD.n1244 DVDD.n972 2.2505
R23206 DVDD.n970 DVDD.n969 2.2505
R23207 DVDD.n1240 DVDD.n1239 2.2505
R23208 DVDD.n1237 DVDD.n1236 2.2505
R23209 DVDD.n1235 DVDD.n977 2.2505
R23210 DVDD.n975 DVDD.n974 2.2505
R23211 DVDD.n1231 DVDD.n1230 2.2505
R23212 DVDD.n1228 DVDD.n1227 2.2505
R23213 DVDD.n1226 DVDD.n982 2.2505
R23214 DVDD.n980 DVDD.n979 2.2505
R23215 DVDD.n1222 DVDD.n1221 2.2505
R23216 DVDD.n1219 DVDD.n1218 2.2505
R23217 DVDD.n1217 DVDD.n987 2.2505
R23218 DVDD.n985 DVDD.n984 2.2505
R23219 DVDD.n1213 DVDD.n1212 2.2505
R23220 DVDD.n1210 DVDD.n1209 2.2505
R23221 DVDD.n1208 DVDD.n992 2.2505
R23222 DVDD.n990 DVDD.n989 2.2505
R23223 DVDD.n1204 DVDD.n1203 2.2505
R23224 DVDD.n1201 DVDD.n1200 2.2505
R23225 DVDD.n1199 DVDD.n997 2.2505
R23226 DVDD.n995 DVDD.n994 2.2505
R23227 DVDD.n1195 DVDD.n1194 2.2505
R23228 DVDD.n1192 DVDD.n1191 2.2505
R23229 DVDD.n1190 DVDD.n1002 2.2505
R23230 DVDD.n1000 DVDD.n999 2.2505
R23231 DVDD.n1186 DVDD.n1185 2.2505
R23232 DVDD.n1183 DVDD.n1182 2.2505
R23233 DVDD.n1181 DVDD.n1007 2.2505
R23234 DVDD.n1005 DVDD.n1004 2.2505
R23235 DVDD.n1177 DVDD.n1176 2.2505
R23236 DVDD.n1174 DVDD.n1173 2.2505
R23237 DVDD.n1172 DVDD.n1012 2.2505
R23238 DVDD.n1010 DVDD.n1009 2.2505
R23239 DVDD.n1168 DVDD.n1167 2.2505
R23240 DVDD.n1165 DVDD.n1164 2.2505
R23241 DVDD.n1163 DVDD.n1017 2.2505
R23242 DVDD.n1015 DVDD.n1014 2.2505
R23243 DVDD.n1159 DVDD.n1158 2.2505
R23244 DVDD.n1156 DVDD.n1155 2.2505
R23245 DVDD.n1154 DVDD.n1022 2.2505
R23246 DVDD.n1020 DVDD.n1019 2.2505
R23247 DVDD.n1150 DVDD.n1149 2.2505
R23248 DVDD.n1147 DVDD.n1146 2.2505
R23249 DVDD.n1145 DVDD.n1027 2.2505
R23250 DVDD.n1025 DVDD.n1024 2.2505
R23251 DVDD.n1141 DVDD.n1140 2.2505
R23252 DVDD.n1138 DVDD.n1137 2.2505
R23253 DVDD.n1136 DVDD.n1032 2.2505
R23254 DVDD.n1030 DVDD.n1029 2.2505
R23255 DVDD.n1132 DVDD.n1131 2.2505
R23256 DVDD.n1129 DVDD.n1128 2.2505
R23257 DVDD.n1127 DVDD.n1037 2.2505
R23258 DVDD.n1035 DVDD.n1034 2.2505
R23259 DVDD.n1123 DVDD.n1122 2.2505
R23260 DVDD.n1120 DVDD.n1119 2.2505
R23261 DVDD.n1118 DVDD.n1042 2.2505
R23262 DVDD.n1040 DVDD.n1039 2.2505
R23263 DVDD.n1114 DVDD.n1113 2.2505
R23264 DVDD.n1111 DVDD.n1110 2.2505
R23265 DVDD.n1109 DVDD.n1047 2.2505
R23266 DVDD.n1045 DVDD.n1044 2.2505
R23267 DVDD.n1105 DVDD.n1104 2.2505
R23268 DVDD.n1102 DVDD.n1101 2.2505
R23269 DVDD.n1100 DVDD.n1052 2.2505
R23270 DVDD.n1050 DVDD.n1049 2.2505
R23271 DVDD.n1096 DVDD.n1095 2.2505
R23272 DVDD.n1093 DVDD.n1092 2.2505
R23273 DVDD.n1091 DVDD.n1057 2.2505
R23274 DVDD.n1055 DVDD.n1054 2.2505
R23275 DVDD.n1087 DVDD.n1086 2.2505
R23276 DVDD.n1084 DVDD.n1083 2.2505
R23277 DVDD.n1082 DVDD.n1062 2.2505
R23278 DVDD.n1060 DVDD.n1059 2.2505
R23279 DVDD.n1078 DVDD.n1077 2.2505
R23280 DVDD.n1075 DVDD.n1074 2.2505
R23281 DVDD.n1073 DVDD.n1067 2.2505
R23282 DVDD.n1065 DVDD.n1064 2.2505
R23283 DVDD.n1069 DVDD.n1068 2.2505
R23284 DVDD.n1070 DVDD.n1069 2.2505
R23285 DVDD.n1071 DVDD.n1064 2.2505
R23286 DVDD.n1073 DVDD.n1072 2.2505
R23287 DVDD.n1074 DVDD.n1063 2.2505
R23288 DVDD.n1079 DVDD.n1078 2.2505
R23289 DVDD.n1080 DVDD.n1059 2.2505
R23290 DVDD.n1082 DVDD.n1081 2.2505
R23291 DVDD.n1083 DVDD.n1058 2.2505
R23292 DVDD.n1088 DVDD.n1087 2.2505
R23293 DVDD.n1089 DVDD.n1054 2.2505
R23294 DVDD.n1091 DVDD.n1090 2.2505
R23295 DVDD.n1092 DVDD.n1053 2.2505
R23296 DVDD.n1097 DVDD.n1096 2.2505
R23297 DVDD.n1098 DVDD.n1049 2.2505
R23298 DVDD.n1100 DVDD.n1099 2.2505
R23299 DVDD.n1101 DVDD.n1048 2.2505
R23300 DVDD.n1106 DVDD.n1105 2.2505
R23301 DVDD.n1107 DVDD.n1044 2.2505
R23302 DVDD.n1109 DVDD.n1108 2.2505
R23303 DVDD.n1110 DVDD.n1043 2.2505
R23304 DVDD.n1115 DVDD.n1114 2.2505
R23305 DVDD.n1116 DVDD.n1039 2.2505
R23306 DVDD.n1118 DVDD.n1117 2.2505
R23307 DVDD.n1119 DVDD.n1038 2.2505
R23308 DVDD.n1124 DVDD.n1123 2.2505
R23309 DVDD.n1125 DVDD.n1034 2.2505
R23310 DVDD.n1127 DVDD.n1126 2.2505
R23311 DVDD.n1128 DVDD.n1033 2.2505
R23312 DVDD.n1133 DVDD.n1132 2.2505
R23313 DVDD.n1134 DVDD.n1029 2.2505
R23314 DVDD.n1136 DVDD.n1135 2.2505
R23315 DVDD.n1137 DVDD.n1028 2.2505
R23316 DVDD.n1142 DVDD.n1141 2.2505
R23317 DVDD.n1143 DVDD.n1024 2.2505
R23318 DVDD.n1145 DVDD.n1144 2.2505
R23319 DVDD.n1146 DVDD.n1023 2.2505
R23320 DVDD.n1151 DVDD.n1150 2.2505
R23321 DVDD.n1152 DVDD.n1019 2.2505
R23322 DVDD.n1154 DVDD.n1153 2.2505
R23323 DVDD.n1155 DVDD.n1018 2.2505
R23324 DVDD.n1160 DVDD.n1159 2.2505
R23325 DVDD.n1161 DVDD.n1014 2.2505
R23326 DVDD.n1163 DVDD.n1162 2.2505
R23327 DVDD.n1164 DVDD.n1013 2.2505
R23328 DVDD.n1169 DVDD.n1168 2.2505
R23329 DVDD.n1170 DVDD.n1009 2.2505
R23330 DVDD.n1172 DVDD.n1171 2.2505
R23331 DVDD.n1173 DVDD.n1008 2.2505
R23332 DVDD.n1178 DVDD.n1177 2.2505
R23333 DVDD.n1179 DVDD.n1004 2.2505
R23334 DVDD.n1181 DVDD.n1180 2.2505
R23335 DVDD.n1182 DVDD.n1003 2.2505
R23336 DVDD.n1187 DVDD.n1186 2.2505
R23337 DVDD.n1188 DVDD.n999 2.2505
R23338 DVDD.n1190 DVDD.n1189 2.2505
R23339 DVDD.n1191 DVDD.n998 2.2505
R23340 DVDD.n1196 DVDD.n1195 2.2505
R23341 DVDD.n1197 DVDD.n994 2.2505
R23342 DVDD.n1199 DVDD.n1198 2.2505
R23343 DVDD.n1200 DVDD.n993 2.2505
R23344 DVDD.n1205 DVDD.n1204 2.2505
R23345 DVDD.n1206 DVDD.n989 2.2505
R23346 DVDD.n1208 DVDD.n1207 2.2505
R23347 DVDD.n1209 DVDD.n988 2.2505
R23348 DVDD.n1214 DVDD.n1213 2.2505
R23349 DVDD.n1215 DVDD.n984 2.2505
R23350 DVDD.n1217 DVDD.n1216 2.2505
R23351 DVDD.n1218 DVDD.n983 2.2505
R23352 DVDD.n1223 DVDD.n1222 2.2505
R23353 DVDD.n1224 DVDD.n979 2.2505
R23354 DVDD.n1226 DVDD.n1225 2.2505
R23355 DVDD.n1227 DVDD.n978 2.2505
R23356 DVDD.n1232 DVDD.n1231 2.2505
R23357 DVDD.n1233 DVDD.n974 2.2505
R23358 DVDD.n1235 DVDD.n1234 2.2505
R23359 DVDD.n1236 DVDD.n973 2.2505
R23360 DVDD.n1241 DVDD.n1240 2.2505
R23361 DVDD.n1242 DVDD.n969 2.2505
R23362 DVDD.n1244 DVDD.n1243 2.2505
R23363 DVDD.n1245 DVDD.n968 2.2505
R23364 DVDD.n1250 DVDD.n1249 2.2505
R23365 DVDD.n1251 DVDD.n967 2.2505
R23366 DVDD.n1253 DVDD.n1252 2.2505
R23367 DVDD.n965 DVDD.n918 2.2505
R23368 DVDD.n15125 DVDD.n15124 2.2505
R23369 DVDD.n5932 DVDD.n5931 2.2505
R23370 DVDD.n6342 DVDD.n6339 2.2505
R23371 DVDD.n15108 DVDD.n15107 2.2505
R23372 DVDD.n15106 DVDD.n6340 2.2505
R23373 DVDD.n15105 DVDD.n15104 2.2505
R23374 DVDD.n7049 DVDD.n7048 2.2505
R23375 DVDD.n7050 DVDD.n7043 2.2505
R23376 DVDD.n15085 DVDD.n15084 2.2505
R23377 DVDD.n15083 DVDD.n7044 2.2505
R23378 DVDD.n15082 DVDD.n15081 2.2505
R23379 DVDD.n15067 DVDD.n15066 2.2505
R23380 DVDD.n15065 DVDD.n7406 2.2505
R23381 DVDD.n15064 DVDD.n15063 2.2505
R23382 DVDD.n7666 DVDD.n7665 2.2505
R23383 DVDD.n7671 DVDD.n7670 2.2505
R23384 DVDD.n7672 DVDD.n7662 2.2505
R23385 DVDD.n14856 DVDD.n14855 2.2505
R23386 DVDD.n14854 DVDD.n7663 2.2505
R23387 DVDD.n14853 DVDD.n14852 2.2505
R23388 DVDD.n8028 DVDD.n8027 2.2505
R23389 DVDD.n8035 DVDD.n8034 2.2505
R23390 DVDD.n8036 DVDD.n8024 2.2505
R23391 DVDD.n14833 DVDD.n14832 2.2505
R23392 DVDD.n14831 DVDD.n8025 2.2505
R23393 DVDD.n14829 DVDD.n14828 2.2505
R23394 DVDD.n8041 DVDD.n8039 2.2505
R23395 DVDD.n14566 DVDD.n14565 2.2505
R23396 DVDD.n14563 DVDD.n14562 2.2505
R23397 DVDD.n8160 DVDD.n8159 2.2505
R23398 DVDD.n8604 DVDD.n8603 2.2505
R23399 DVDD.n14300 DVDD.n14299 2.2505
R23400 DVDD.n14298 DVDD.n8263 2.2505
R23401 DVDD.n14297 DVDD.n14296 2.2505
R23402 DVDD.n10581 DVDD.n10580 2.2505
R23403 DVDD.n10588 DVDD.n10587 2.2505
R23404 DVDD.n10589 DVDD.n10577 2.2505
R23405 DVDD.n14277 DVDD.n14276 2.2505
R23406 DVDD.n14275 DVDD.n10578 2.2505
R23407 DVDD.n14273 DVDD.n14272 2.2505
R23408 DVDD.n10594 DVDD.n10592 2.2505
R23409 DVDD.n11056 DVDD.n11055 2.2505
R23410 DVDD.n14010 DVDD.n14009 2.2505
R23411 DVDD.n14008 DVDD.n10715 2.2505
R23412 DVDD.n14007 DVDD.n14006 2.2505
R23413 DVDD.n11571 DVDD.n11570 2.2505
R23414 DVDD.n11569 DVDD.n11567 2.2505
R23415 DVDD.n11576 DVDD.n11565 2.2505
R23416 DVDD.n13791 DVDD.n13790 2.2505
R23417 DVDD.n11578 DVDD.n11566 2.2505
R23418 DVDD.n11921 DVDD.n11919 2.2505
R23419 DVDD.n13769 DVDD.n13768 2.2505
R23420 DVDD.n11923 DVDD.n11920 2.2505
R23421 DVDD.n12279 DVDD.n12278 2.2505
R23422 DVDD.n13752 DVDD.n13751 2.2505
R23423 DVDD.n13750 DVDD.n11943 2.2505
R23424 DVDD.n13748 DVDD.n13747 2.2505
R23425 DVDD.n12284 DVDD.n12282 2.2505
R23426 DVDD.n12730 DVDD.n12727 2.2505
R23427 DVDD.n13480 DVDD.n13479 2.2505
R23428 DVDD.n13478 DVDD.n12728 2.2505
R23429 DVDD.n13477 DVDD.n13476 2.2505
R23430 DVDD.n12919 DVDD.n12918 2.2505
R23431 DVDD.n12917 DVDD.n12916 2.2505
R23432 DVDD.n13261 DVDD.n13260 2.2505
R23433 DVDD.n13264 DVDD.n13263 2.2505
R23434 DVDD.n2161 DVDD.n2160 2.2505
R23435 DVDD.n16708 DVDD.n16707 2.2505
R23436 DVDD.n16710 DVDD.n2158 2.2505
R23437 DVDD.n16712 DVDD.n16711 2.2505
R23438 DVDD.n16730 DVDD.n16729 2.2505
R23439 DVDD.n16731 DVDD.n1807 2.2505
R23440 DVDD.n16733 DVDD.n16732 2.2505
R23441 DVDD.n16998 DVDD.n16997 2.2505
R23442 DVDD.n16999 DVDD.n1708 2.2505
R23443 DVDD.n17001 DVDD.n17000 2.2505
R23444 DVDD.n17266 DVDD.n17265 2.2505
R23445 DVDD.n17267 DVDD.n1607 2.2505
R23446 DVDD.n17269 DVDD.n17268 2.2505
R23447 DVDD.n17284 DVDD.n17283 2.2505
R23448 DVDD.n17285 DVDD.n1258 2.2505
R23449 DVDD.n17287 DVDD.n17286 2.2505
R23450 DVDD.n17303 DVDD.n17302 2.2505
R23451 DVDD.n17304 DVDD.n910 2.2505
R23452 DVDD.n17715 DVDD.n17714 2.2505
R23453 DVDD.n3034 DVDD.n3007 2.25007
R23454 DVDD.n3039 DVDD.n3007 2.25007
R23455 DVDD.n2769 DVDD.n2768 2.25007
R23456 DVDD.n2769 DVDD.n2722 2.25007
R23457 DVDD.n2694 DVDD.n2656 2.25007
R23458 DVDD.n2699 DVDD.n2656 2.25007
R23459 DVDD.n2361 DVDD.n2360 2.25007
R23460 DVDD.n2361 DVDD.n2359 2.25007
R23461 DVDD.n4531 DVDD.n4530 2.25007
R23462 DVDD.n4531 DVDD.n4529 2.25007
R23463 DVDD.n2964 DVDD.n2936 2.25007
R23464 DVDD.n2969 DVDD.n2936 2.25007
R23465 DVDD.n2823 DVDD.n2791 2.25007
R23466 DVDD.n2828 DVDD.n2791 2.25007
R23467 DVDD.n2621 DVDD.n2583 2.25007
R23468 DVDD.n2626 DVDD.n2583 2.25007
R23469 DVDD.n2485 DVDD.n2401 2.25007
R23470 DVDD.n2485 DVDD.n2484 2.25007
R23471 DVDD.n4634 DVDD.n4602 2.25007
R23472 DVDD.n4641 DVDD.n4602 2.25007
R23473 DVDD.n9778 DVDD.n9777 2.25007
R23474 DVDD.n9778 DVDD.n3095 2.25007
R23475 DVDD.n3195 DVDD.n3161 2.25007
R23476 DVDD.n15930 DVDD.n3161 2.25007
R23477 DVDD.n3288 DVDD.n3247 2.25007
R23478 DVDD.n3292 DVDD.n3247 2.25007
R23479 DVDD.n3398 DVDD.n3260 2.25007
R23480 DVDD.n3403 DVDD.n3260 2.25007
R23481 DVDD.n3815 DVDD.n3783 2.25007
R23482 DVDD.n4162 DVDD.n3783 2.25007
R23483 DVDD.n3578 DVDD.n3577 2.25007
R23484 DVDD.n15708 DVDD.n4881 2.25007
R23485 DVDD.n15713 DVDD.n3520 2.25007
R23486 DVDD.n15701 DVDD.n5044 2.25007
R23487 DVDD.n15701 DVDD.n5040 2.25007
R23488 DVDD.n15422 DVDD.n5241 2.25007
R23489 DVDD.n15417 DVDD.n5241 2.25007
R23490 DVDD.n15409 DVDD.n5373 2.25007
R23491 DVDD.n15409 DVDD.n5371 2.25007
R23492 DVDD.n760 DVDD.n759 2.25007
R23493 DVDD.n760 DVDD.n758 2.25007
R23494 DVDD.n669 DVDD.n668 2.25007
R23495 DVDD.n669 DVDD.n667 2.25007
R23496 DVDD.n582 DVDD.n581 2.25007
R23497 DVDD.n582 DVDD.n580 2.25007
R23498 DVDD.n532 DVDD.n531 2.25007
R23499 DVDD.n18039 DVDD.n532 2.25007
R23500 DVDD.n474 DVDD.n473 2.25007
R23501 DVDD.n3136 DVDD.n3135 2.25007
R23502 DVDD.n16053 DVDD.n3134 2.25007
R23503 DVDD.n5158 DVDD.n5157 2.25007
R23504 DVDD.n5158 DVDD.n5156 2.25007
R23505 DVDD.n15612 DVDD.n15534 2.25007
R23506 DVDD.n15617 DVDD.n5128 2.25007
R23507 DVDD.n3491 DVDD.n3431 2.25007
R23508 DVDD.n15792 DVDD.n3431 2.25007
R23509 DVDD.n4088 DVDD.n3839 2.25007
R23510 DVDD.n8961 DVDD.n8950 2.24982
R23511 DVDD.n2280 DVDD.n2278 2.24982
R23512 DVDD.n2266 DVDD.n2256 2.24982
R23513 DVDD.n8963 DVDD.n8959 2.24982
R23514 DVDD.n16428 DVDD.n2283 2.24982
R23515 DVDD.n2270 DVDD.n2269 2.24982
R23516 DVDD.n8973 DVDD.n8971 2.24982
R23517 DVDD.n10199 DVDD.n10168 2.24982
R23518 DVDD.n18799 DVDD.n18796 2.24964
R23519 DVDD.n18772 DVDD.n18771 2.24964
R23520 DVDD.n20481 DVDD.n20480 2.24964
R23521 DVDD.n19819 DVDD.n19810 2.24964
R23522 DVDD.n20443 DVDD.n20442 2.24964
R23523 DVDD.n9680 DVDD.n9678 2.24964
R23524 DVDD.n9669 DVDD.n9661 2.24964
R23525 DVDD.n9680 DVDD.n9679 2.24964
R23526 DVDD.n9673 DVDD.n9661 2.24964
R23527 DVDD.n3008 DVDD.n2995 2.24964
R23528 DVDD.n16113 DVDD.n16112 2.24964
R23529 DVDD.n3010 DVDD.n2995 2.24964
R23530 DVDD.n16113 DVDD.n16111 2.24964
R23531 DVDD.n3013 DVDD.n2995 2.24964
R23532 DVDD.n16113 DVDD.n16110 2.24964
R23533 DVDD.n3015 DVDD.n2995 2.24964
R23534 DVDD.n16113 DVDD.n16109 2.24964
R23535 DVDD.n16113 DVDD.n16108 2.24964
R23536 DVDD.n3018 DVDD.n2995 2.24964
R23537 DVDD.n16113 DVDD.n16107 2.24964
R23538 DVDD.n16113 DVDD.n16106 2.24964
R23539 DVDD.n3021 DVDD.n2995 2.24964
R23540 DVDD.n16113 DVDD.n16105 2.24964
R23541 DVDD.n2746 DVDD.n2735 2.24964
R23542 DVDD.n2764 DVDD.n2763 2.24964
R23543 DVDD.n2746 DVDD.n2736 2.24964
R23544 DVDD.n2746 DVDD.n2737 2.24964
R23545 DVDD.n2764 DVDD.n2762 2.24964
R23546 DVDD.n2746 DVDD.n2738 2.24964
R23547 DVDD.n2746 DVDD.n2739 2.24964
R23548 DVDD.n2764 DVDD.n2761 2.24964
R23549 DVDD.n2746 DVDD.n2740 2.24964
R23550 DVDD.n2746 DVDD.n2741 2.24964
R23551 DVDD.n2764 DVDD.n2760 2.24964
R23552 DVDD.n2746 DVDD.n2742 2.24964
R23553 DVDD.n2764 DVDD.n2759 2.24964
R23554 DVDD.n2746 DVDD.n2743 2.24964
R23555 DVDD.n2764 DVDD.n2758 2.24964
R23556 DVDD.n2746 DVDD.n2744 2.24964
R23557 DVDD.n2746 DVDD.n2745 2.24964
R23558 DVDD.n2764 DVDD.n2747 2.24964
R23559 DVDD.n2657 DVDD.n2644 2.24964
R23560 DVDD.n2685 DVDD.n2684 2.24964
R23561 DVDD.n2659 DVDD.n2644 2.24964
R23562 DVDD.n2685 DVDD.n2683 2.24964
R23563 DVDD.n2661 DVDD.n2644 2.24964
R23564 DVDD.n2663 DVDD.n2644 2.24964
R23565 DVDD.n2685 DVDD.n2682 2.24964
R23566 DVDD.n2665 DVDD.n2644 2.24964
R23567 DVDD.n2667 DVDD.n2644 2.24964
R23568 DVDD.n2685 DVDD.n2681 2.24964
R23569 DVDD.n2669 DVDD.n2644 2.24964
R23570 DVDD.n2671 DVDD.n2644 2.24964
R23571 DVDD.n2685 DVDD.n2680 2.24964
R23572 DVDD.n2673 DVDD.n2644 2.24964
R23573 DVDD.n2675 DVDD.n2644 2.24964
R23574 DVDD.n2685 DVDD.n2679 2.24964
R23575 DVDD.n2677 DVDD.n2644 2.24964
R23576 DVDD.n16390 DVDD.n16382 2.24964
R23577 DVDD.n2364 DVDD.n2335 2.24964
R23578 DVDD.n16390 DVDD.n16383 2.24964
R23579 DVDD.n16390 DVDD.n16384 2.24964
R23580 DVDD.n2367 DVDD.n2335 2.24964
R23581 DVDD.n16390 DVDD.n16385 2.24964
R23582 DVDD.n16390 DVDD.n16386 2.24964
R23583 DVDD.n2370 DVDD.n2335 2.24964
R23584 DVDD.n16390 DVDD.n16387 2.24964
R23585 DVDD.n2372 DVDD.n2335 2.24964
R23586 DVDD.n16390 DVDD.n16388 2.24964
R23587 DVDD.n2374 DVDD.n2335 2.24964
R23588 DVDD.n16390 DVDD.n2334 2.24964
R23589 DVDD.n16390 DVDD.n16389 2.24964
R23590 DVDD.n16392 DVDD.n2335 2.24964
R23591 DVDD.n16391 DVDD.n16390 2.24964
R23592 DVDD.n4555 DVDD.n4411 2.24964
R23593 DVDD.n4330 DVDD.n4323 2.24964
R23594 DVDD.n4399 DVDD.n4397 2.24964
R23595 DVDD.n4399 DVDD.n4396 2.24964
R23596 DVDD.n4399 DVDD.n4395 2.24964
R23597 DVDD.n4517 DVDD.n4516 2.24964
R23598 DVDD.n4528 DVDD.n4518 2.24964
R23599 DVDD.n4516 DVDD.n4515 2.24964
R23600 DVDD.n4528 DVDD.n4519 2.24964
R23601 DVDD.n4516 DVDD.n4514 2.24964
R23602 DVDD.n4528 DVDD.n4520 2.24964
R23603 DVDD.n4516 DVDD.n4513 2.24964
R23604 DVDD.n4528 DVDD.n4521 2.24964
R23605 DVDD.n4516 DVDD.n4512 2.24964
R23606 DVDD.n4528 DVDD.n4522 2.24964
R23607 DVDD.n4516 DVDD.n4511 2.24964
R23608 DVDD.n4528 DVDD.n4523 2.24964
R23609 DVDD.n4516 DVDD.n4510 2.24964
R23610 DVDD.n4528 DVDD.n4524 2.24964
R23611 DVDD.n4516 DVDD.n4509 2.24964
R23612 DVDD.n4528 DVDD.n4525 2.24964
R23613 DVDD.n4516 DVDD.n4508 2.24964
R23614 DVDD.n4528 DVDD.n4526 2.24964
R23615 DVDD.n4516 DVDD.n4507 2.24964
R23616 DVDD.n4528 DVDD.n4527 2.24964
R23617 DVDD.n4516 DVDD.n4490 2.24964
R23618 DVDD.n4528 DVDD.n4489 2.24964
R23619 DVDD.n4516 DVDD.n4506 2.24964
R23620 DVDD.n320 DVDD.n291 2.24964
R23621 DVDD.n22160 DVDD.n289 2.24964
R23622 DVDD.n320 DVDD.n316 2.24964
R23623 DVDD.n22160 DVDD.n288 2.24964
R23624 DVDD.n320 DVDD.n317 2.24964
R23625 DVDD.n22160 DVDD.n287 2.24964
R23626 DVDD.n320 DVDD.n318 2.24964
R23627 DVDD.n22160 DVDD.n286 2.24964
R23628 DVDD.n320 DVDD.n319 2.24964
R23629 DVDD.n22160 DVDD.n285 2.24964
R23630 DVDD.n19045 DVDD.n19044 2.24964
R23631 DVDD.n19057 DVDD.n19055 2.24964
R23632 DVDD.n19045 DVDD.n19043 2.24964
R23633 DVDD.n19057 DVDD.n19056 2.24964
R23634 DVDD.n19045 DVDD.n19042 2.24964
R23635 DVDD.n19057 DVDD.n19034 2.24964
R23636 DVDD.n19045 DVDD.n19041 2.24964
R23637 DVDD.n4556 DVDD.n4555 2.24964
R23638 DVDD.n4555 DVDD.n4410 2.24964
R23639 DVDD.n4555 DVDD.n4409 2.24964
R23640 DVDD.n4555 DVDD.n4408 2.24964
R23641 DVDD.n2376 DVDD.n2335 2.24964
R23642 DVDD.n16113 DVDD.n16104 2.24964
R23643 DVDD.n16113 DVDD.n16103 2.24964
R23644 DVDD.n16113 DVDD.n3025 2.24964
R23645 DVDD.n9675 DVDD.n9661 2.24964
R23646 DVDD.n9671 DVDD.n9661 2.24964
R23647 DVDD.n9677 DVDD.n9661 2.24964
R23648 DVDD.n19099 DVDD.n19096 2.24964
R23649 DVDD.n20924 DVDD.n18905 2.24964
R23650 DVDD.n9750 DVDD.n9747 2.24964
R23651 DVDD.n10001 DVDD.n10000 2.24964
R23652 DVDD.n9750 DVDD.n9748 2.24964
R23653 DVDD.n10001 DVDD.n9999 2.24964
R23654 DVDD.n2937 DVDD.n2924 2.24964
R23655 DVDD.n2980 DVDD.n2975 2.24964
R23656 DVDD.n2939 DVDD.n2924 2.24964
R23657 DVDD.n2980 DVDD.n2974 2.24964
R23658 DVDD.n2942 DVDD.n2924 2.24964
R23659 DVDD.n2980 DVDD.n2976 2.24964
R23660 DVDD.n2944 DVDD.n2924 2.24964
R23661 DVDD.n2980 DVDD.n2973 2.24964
R23662 DVDD.n2947 DVDD.n2924 2.24964
R23663 DVDD.n2980 DVDD.n2977 2.24964
R23664 DVDD.n2949 DVDD.n2924 2.24964
R23665 DVDD.n2951 DVDD.n2924 2.24964
R23666 DVDD.n2980 DVDD.n2978 2.24964
R23667 DVDD.n2953 DVDD.n2924 2.24964
R23668 DVDD.n2816 DVDD.n2805 2.24964
R23669 DVDD.n2872 DVDD.n2871 2.24964
R23670 DVDD.n2816 DVDD.n2806 2.24964
R23671 DVDD.n2816 DVDD.n2807 2.24964
R23672 DVDD.n2872 DVDD.n2870 2.24964
R23673 DVDD.n2816 DVDD.n2808 2.24964
R23674 DVDD.n2816 DVDD.n2809 2.24964
R23675 DVDD.n2872 DVDD.n2869 2.24964
R23676 DVDD.n2816 DVDD.n2810 2.24964
R23677 DVDD.n2816 DVDD.n2811 2.24964
R23678 DVDD.n2872 DVDD.n2868 2.24964
R23679 DVDD.n2816 DVDD.n2812 2.24964
R23680 DVDD.n2872 DVDD.n2867 2.24964
R23681 DVDD.n2816 DVDD.n2813 2.24964
R23682 DVDD.n2872 DVDD.n2866 2.24964
R23683 DVDD.n2816 DVDD.n2814 2.24964
R23684 DVDD.n2816 DVDD.n2815 2.24964
R23685 DVDD.n2872 DVDD.n2817 2.24964
R23686 DVDD.n2606 DVDD.n2595 2.24964
R23687 DVDD.n2613 DVDD.n2612 2.24964
R23688 DVDD.n2606 DVDD.n2596 2.24964
R23689 DVDD.n2613 DVDD.n2611 2.24964
R23690 DVDD.n2606 DVDD.n2597 2.24964
R23691 DVDD.n2606 DVDD.n2598 2.24964
R23692 DVDD.n2613 DVDD.n2610 2.24964
R23693 DVDD.n2606 DVDD.n2599 2.24964
R23694 DVDD.n2606 DVDD.n2600 2.24964
R23695 DVDD.n2613 DVDD.n2609 2.24964
R23696 DVDD.n2606 DVDD.n2601 2.24964
R23697 DVDD.n2606 DVDD.n2602 2.24964
R23698 DVDD.n2613 DVDD.n2608 2.24964
R23699 DVDD.n2606 DVDD.n2603 2.24964
R23700 DVDD.n2606 DVDD.n2604 2.24964
R23701 DVDD.n2613 DVDD.n2607 2.24964
R23702 DVDD.n2606 DVDD.n2605 2.24964
R23703 DVDD.n2424 DVDD.n2414 2.24964
R23704 DVDD.n2432 DVDD.n2430 2.24964
R23705 DVDD.n2424 DVDD.n2415 2.24964
R23706 DVDD.n2424 DVDD.n2416 2.24964
R23707 DVDD.n2432 DVDD.n2429 2.24964
R23708 DVDD.n2424 DVDD.n2417 2.24964
R23709 DVDD.n2424 DVDD.n2418 2.24964
R23710 DVDD.n2432 DVDD.n2428 2.24964
R23711 DVDD.n2424 DVDD.n2419 2.24964
R23712 DVDD.n2432 DVDD.n2427 2.24964
R23713 DVDD.n2424 DVDD.n2420 2.24964
R23714 DVDD.n2432 DVDD.n2426 2.24964
R23715 DVDD.n2424 DVDD.n2421 2.24964
R23716 DVDD.n2424 DVDD.n2422 2.24964
R23717 DVDD.n2432 DVDD.n2425 2.24964
R23718 DVDD.n2424 DVDD.n2423 2.24964
R23719 DVDD.n4259 DVDD.n4245 2.24964
R23720 DVDD.n4270 DVDD.n4246 2.24964
R23721 DVDD.n4598 DVDD.n4597 2.24964
R23722 DVDD.n4266 DVDD.n4245 2.24964
R23723 DVDD.n4267 DVDD.n4246 2.24964
R23724 DVDD.n4597 DVDD.n4273 2.24964
R23725 DVDD.n4597 DVDD.n4272 2.24964
R23726 DVDD.n4263 DVDD.n4246 2.24964
R23727 DVDD.n4597 DVDD.n4247 2.24964
R23728 DVDD.n4655 DVDD.n4654 2.24964
R23729 DVDD.n4626 DVDD.n4615 2.24964
R23730 DVDD.n4655 DVDD.n4653 2.24964
R23731 DVDD.n4626 DVDD.n4616 2.24964
R23732 DVDD.n4655 DVDD.n4652 2.24964
R23733 DVDD.n4626 DVDD.n4617 2.24964
R23734 DVDD.n4655 DVDD.n4651 2.24964
R23735 DVDD.n4626 DVDD.n4618 2.24964
R23736 DVDD.n4655 DVDD.n4650 2.24964
R23737 DVDD.n4626 DVDD.n4619 2.24964
R23738 DVDD.n4655 DVDD.n4649 2.24964
R23739 DVDD.n4626 DVDD.n4620 2.24964
R23740 DVDD.n4655 DVDD.n4648 2.24964
R23741 DVDD.n4626 DVDD.n4621 2.24964
R23742 DVDD.n4655 DVDD.n4647 2.24964
R23743 DVDD.n4626 DVDD.n4622 2.24964
R23744 DVDD.n4655 DVDD.n4646 2.24964
R23745 DVDD.n4626 DVDD.n4623 2.24964
R23746 DVDD.n4655 DVDD.n4645 2.24964
R23747 DVDD.n4626 DVDD.n4624 2.24964
R23748 DVDD.n4655 DVDD.n4644 2.24964
R23749 DVDD.n4626 DVDD.n4625 2.24964
R23750 DVDD.n4655 DVDD.n4614 2.24964
R23751 DVDD.n372 DVDD.n367 2.24964
R23752 DVDD.n426 DVDD.n425 2.24964
R23753 DVDD.n372 DVDD.n368 2.24964
R23754 DVDD.n426 DVDD.n424 2.24964
R23755 DVDD.n372 DVDD.n369 2.24964
R23756 DVDD.n426 DVDD.n423 2.24964
R23757 DVDD.n372 DVDD.n370 2.24964
R23758 DVDD.n426 DVDD.n422 2.24964
R23759 DVDD.n372 DVDD.n371 2.24964
R23760 DVDD.n426 DVDD.n373 2.24964
R23761 DVDD.n18898 DVDD.n18882 2.24964
R23762 DVDD.n18897 DVDD.n18881 2.24964
R23763 DVDD.n18901 DVDD.n18882 2.24964
R23764 DVDD.n18900 DVDD.n18881 2.24964
R23765 DVDD.n18903 DVDD.n18882 2.24964
R23766 DVDD.n18888 DVDD.n18881 2.24964
R23767 DVDD.n20927 DVDD.n18882 2.24964
R23768 DVDD.n2432 DVDD.n2431 2.24964
R23769 DVDD.n2980 DVDD.n2979 2.24964
R23770 DVDD.n2980 DVDD.n2972 2.24964
R23771 DVDD.n2980 DVDD.n2956 2.24964
R23772 DVDD.n9750 DVDD.n9749 2.24964
R23773 DVDD.n10001 DVDD.n9998 2.24964
R23774 DVDD.n10001 DVDD.n9746 2.24964
R23775 DVDD.n21060 DVDD.n18752 2.24964
R23776 DVDD.n21057 DVDD.n18754 2.24964
R23777 DVDD.n20533 DVDD.n19797 2.24964
R23778 DVDD.n19790 DVDD.n19781 2.24964
R23779 DVDD.n20536 DVDD.n19767 2.24964
R23780 DVDD.n9633 DVDD.n9613 2.24964
R23781 DVDD.n9648 DVDD.n9647 2.24964
R23782 DVDD.n9635 DVDD.n9613 2.24964
R23783 DVDD.n9648 DVDD.n9646 2.24964
R23784 DVDD.n16085 DVDD.n3067 2.24964
R23785 DVDD.n16081 DVDD.n16076 2.24964
R23786 DVDD.n16085 DVDD.n3069 2.24964
R23787 DVDD.n16081 DVDD.n16074 2.24964
R23788 DVDD.n16085 DVDD.n3065 2.24964
R23789 DVDD.n16081 DVDD.n16077 2.24964
R23790 DVDD.n16085 DVDD.n3071 2.24964
R23791 DVDD.n16081 DVDD.n16073 2.24964
R23792 DVDD.n16085 DVDD.n3063 2.24964
R23793 DVDD.n16081 DVDD.n16078 2.24964
R23794 DVDD.n16085 DVDD.n3062 2.24964
R23795 DVDD.n16085 DVDD.n3061 2.24964
R23796 DVDD.n16081 DVDD.n16079 2.24964
R23797 DVDD.n16085 DVDD.n3060 2.24964
R23798 DVDD.n3186 DVDD.n3175 2.24964
R23799 DVDD.n15937 DVDD.n15936 2.24964
R23800 DVDD.n3186 DVDD.n3176 2.24964
R23801 DVDD.n3186 DVDD.n3177 2.24964
R23802 DVDD.n15937 DVDD.n15935 2.24964
R23803 DVDD.n3186 DVDD.n3178 2.24964
R23804 DVDD.n3186 DVDD.n3179 2.24964
R23805 DVDD.n15937 DVDD.n15934 2.24964
R23806 DVDD.n3186 DVDD.n3180 2.24964
R23807 DVDD.n3186 DVDD.n3181 2.24964
R23808 DVDD.n15937 DVDD.n15933 2.24964
R23809 DVDD.n3186 DVDD.n3182 2.24964
R23810 DVDD.n15937 DVDD.n15932 2.24964
R23811 DVDD.n3186 DVDD.n3183 2.24964
R23812 DVDD.n15937 DVDD.n15931 2.24964
R23813 DVDD.n3186 DVDD.n3184 2.24964
R23814 DVDD.n3186 DVDD.n3185 2.24964
R23815 DVDD.n15937 DVDD.n3187 2.24964
R23816 DVDD.n3272 DVDD.n3261 2.24964
R23817 DVDD.n3279 DVDD.n3278 2.24964
R23818 DVDD.n3272 DVDD.n3262 2.24964
R23819 DVDD.n3279 DVDD.n3277 2.24964
R23820 DVDD.n3272 DVDD.n3263 2.24964
R23821 DVDD.n3272 DVDD.n3264 2.24964
R23822 DVDD.n3279 DVDD.n3276 2.24964
R23823 DVDD.n3272 DVDD.n3265 2.24964
R23824 DVDD.n3272 DVDD.n3266 2.24964
R23825 DVDD.n3279 DVDD.n3275 2.24964
R23826 DVDD.n3272 DVDD.n3267 2.24964
R23827 DVDD.n3272 DVDD.n3268 2.24964
R23828 DVDD.n3279 DVDD.n3274 2.24964
R23829 DVDD.n3272 DVDD.n3269 2.24964
R23830 DVDD.n3272 DVDD.n3270 2.24964
R23831 DVDD.n3279 DVDD.n3273 2.24964
R23832 DVDD.n3272 DVDD.n3271 2.24964
R23833 DVDD.n3381 DVDD.n3371 2.24964
R23834 DVDD.n3389 DVDD.n3387 2.24964
R23835 DVDD.n3381 DVDD.n3372 2.24964
R23836 DVDD.n3381 DVDD.n3373 2.24964
R23837 DVDD.n3389 DVDD.n3386 2.24964
R23838 DVDD.n3381 DVDD.n3374 2.24964
R23839 DVDD.n3381 DVDD.n3375 2.24964
R23840 DVDD.n3389 DVDD.n3385 2.24964
R23841 DVDD.n3381 DVDD.n3376 2.24964
R23842 DVDD.n3389 DVDD.n3384 2.24964
R23843 DVDD.n3381 DVDD.n3377 2.24964
R23844 DVDD.n3389 DVDD.n3383 2.24964
R23845 DVDD.n3381 DVDD.n3378 2.24964
R23846 DVDD.n3381 DVDD.n3379 2.24964
R23847 DVDD.n3389 DVDD.n3382 2.24964
R23848 DVDD.n3381 DVDD.n3380 2.24964
R23849 DVDD.n3746 DVDD.n3745 2.24964
R23850 DVDD.n4441 DVDD.n3747 2.24964
R23851 DVDD.n4419 DVDD.n3740 2.24964
R23852 DVDD.n4419 DVDD.n4418 2.24964
R23853 DVDD.n4419 DVDD.n4417 2.24964
R23854 DVDD.n4175 DVDD.n4174 2.24964
R23855 DVDD.n3807 DVDD.n3796 2.24964
R23856 DVDD.n4175 DVDD.n4173 2.24964
R23857 DVDD.n3807 DVDD.n3797 2.24964
R23858 DVDD.n4175 DVDD.n4172 2.24964
R23859 DVDD.n3807 DVDD.n3798 2.24964
R23860 DVDD.n4175 DVDD.n4171 2.24964
R23861 DVDD.n3807 DVDD.n3799 2.24964
R23862 DVDD.n4175 DVDD.n4170 2.24964
R23863 DVDD.n3807 DVDD.n3800 2.24964
R23864 DVDD.n4175 DVDD.n4169 2.24964
R23865 DVDD.n3807 DVDD.n3801 2.24964
R23866 DVDD.n4175 DVDD.n4168 2.24964
R23867 DVDD.n3807 DVDD.n3802 2.24964
R23868 DVDD.n4175 DVDD.n4167 2.24964
R23869 DVDD.n3807 DVDD.n3803 2.24964
R23870 DVDD.n4175 DVDD.n4166 2.24964
R23871 DVDD.n3807 DVDD.n3804 2.24964
R23872 DVDD.n4175 DVDD.n4165 2.24964
R23873 DVDD.n3807 DVDD.n3805 2.24964
R23874 DVDD.n4175 DVDD.n4164 2.24964
R23875 DVDD.n3807 DVDD.n3806 2.24964
R23876 DVDD.n4175 DVDD.n3795 2.24964
R23877 DVDD.n258 DVDD.n236 2.24964
R23878 DVDD.n22178 DVDD.n271 2.24964
R23879 DVDD.n261 DVDD.n236 2.24964
R23880 DVDD.n22178 DVDD.n270 2.24964
R23881 DVDD.n263 DVDD.n236 2.24964
R23882 DVDD.n22178 DVDD.n269 2.24964
R23883 DVDD.n265 DVDD.n236 2.24964
R23884 DVDD.n22179 DVDD.n22178 2.24964
R23885 DVDD.n267 DVDD.n236 2.24964
R23886 DVDD.n22178 DVDD.n237 2.24964
R23887 DVDD.n19153 DVDD.n19152 2.24964
R23888 DVDD.n19134 DVDD.n19132 2.24964
R23889 DVDD.n19153 DVDD.n19151 2.24964
R23890 DVDD.n19134 DVDD.n19133 2.24964
R23891 DVDD.n19153 DVDD.n19150 2.24964
R23892 DVDD.n19153 DVDD.n19130 2.24964
R23893 DVDD.n19134 DVDD.n19131 2.24964
R23894 DVDD.n3746 DVDD.n3744 2.24964
R23895 DVDD.n3746 DVDD.n3743 2.24964
R23896 DVDD.n3746 DVDD.n3742 2.24964
R23897 DVDD.n3746 DVDD.n3741 2.24964
R23898 DVDD.n3389 DVDD.n3388 2.24964
R23899 DVDD.n16081 DVDD.n16080 2.24964
R23900 DVDD.n16081 DVDD.n16072 2.24964
R23901 DVDD.n16081 DVDD.n3074 2.24964
R23902 DVDD.n9638 DVDD.n9613 2.24964
R23903 DVDD.n9648 DVDD.n9645 2.24964
R23904 DVDD.n9648 DVDD.n9640 2.24964
R23905 DVDD.n20980 DVDD.n18824 2.24964
R23906 DVDD.n20525 DVDD.n20520 2.24964
R23907 DVDD.n9808 DVDD.n9757 2.24964
R23908 DVDD.n9939 DVDD.n9938 2.24964
R23909 DVDD.n9810 DVDD.n9757 2.24964
R23910 DVDD.n9939 DVDD.n9816 2.24964
R23911 DVDD.n16061 DVDD.n16058 2.24964
R23912 DVDD.n16007 DVDD.n3109 2.24964
R23913 DVDD.n16061 DVDD.n16059 2.24964
R23914 DVDD.n16017 DVDD.n3109 2.24964
R23915 DVDD.n16061 DVDD.n16057 2.24964
R23916 DVDD.n16019 DVDD.n3109 2.24964
R23917 DVDD.n16061 DVDD.n16060 2.24964
R23918 DVDD.n16029 DVDD.n3109 2.24964
R23919 DVDD.n16061 DVDD.n16056 2.24964
R23920 DVDD.n16031 DVDD.n3109 2.24964
R23921 DVDD.n16061 DVDD.n16055 2.24964
R23922 DVDD.n16061 DVDD.n16054 2.24964
R23923 DVDD.n16041 DVDD.n3109 2.24964
R23924 DVDD.n16061 DVDD.n3108 2.24964
R23925 DVDD.n5160 DVDD.n5129 2.24964
R23926 DVDD.n15520 DVDD.n5214 2.24964
R23927 DVDD.n5169 DVDD.n5129 2.24964
R23928 DVDD.n5171 DVDD.n5129 2.24964
R23929 DVDD.n15520 DVDD.n5213 2.24964
R23930 DVDD.n5180 DVDD.n5129 2.24964
R23931 DVDD.n5182 DVDD.n5129 2.24964
R23932 DVDD.n15520 DVDD.n5212 2.24964
R23933 DVDD.n5191 DVDD.n5129 2.24964
R23934 DVDD.n5193 DVDD.n5129 2.24964
R23935 DVDD.n15520 DVDD.n5211 2.24964
R23936 DVDD.n5201 DVDD.n5129 2.24964
R23937 DVDD.n15520 DVDD.n5210 2.24964
R23938 DVDD.n5203 DVDD.n5129 2.24964
R23939 DVDD.n15520 DVDD.n5209 2.24964
R23940 DVDD.n5205 DVDD.n5129 2.24964
R23941 DVDD.n5207 DVDD.n5129 2.24964
R23942 DVDD.n15520 DVDD.n5130 2.24964
R23943 DVDD.n15593 DVDD.n15582 2.24964
R23944 DVDD.n15600 DVDD.n15599 2.24964
R23945 DVDD.n15593 DVDD.n15583 2.24964
R23946 DVDD.n15600 DVDD.n15598 2.24964
R23947 DVDD.n15593 DVDD.n15584 2.24964
R23948 DVDD.n15593 DVDD.n15585 2.24964
R23949 DVDD.n15600 DVDD.n15597 2.24964
R23950 DVDD.n15593 DVDD.n15586 2.24964
R23951 DVDD.n15593 DVDD.n15587 2.24964
R23952 DVDD.n15600 DVDD.n15596 2.24964
R23953 DVDD.n15593 DVDD.n15588 2.24964
R23954 DVDD.n15593 DVDD.n15589 2.24964
R23955 DVDD.n15600 DVDD.n15595 2.24964
R23956 DVDD.n15593 DVDD.n15590 2.24964
R23957 DVDD.n15593 DVDD.n15591 2.24964
R23958 DVDD.n15600 DVDD.n15594 2.24964
R23959 DVDD.n15593 DVDD.n15592 2.24964
R23960 DVDD.n3432 DVDD.n3419 2.24964
R23961 DVDD.n3481 DVDD.n3479 2.24964
R23962 DVDD.n3441 DVDD.n3419 2.24964
R23963 DVDD.n3443 DVDD.n3419 2.24964
R23964 DVDD.n3481 DVDD.n3478 2.24964
R23965 DVDD.n3452 DVDD.n3419 2.24964
R23966 DVDD.n3454 DVDD.n3419 2.24964
R23967 DVDD.n3481 DVDD.n3477 2.24964
R23968 DVDD.n3462 DVDD.n3419 2.24964
R23969 DVDD.n3481 DVDD.n3476 2.24964
R23970 DVDD.n3464 DVDD.n3419 2.24964
R23971 DVDD.n3481 DVDD.n3475 2.24964
R23972 DVDD.n3466 DVDD.n3419 2.24964
R23973 DVDD.n3468 DVDD.n3419 2.24964
R23974 DVDD.n3481 DVDD.n3474 2.24964
R23975 DVDD.n3470 DVDD.n3419 2.24964
R23976 DVDD.n3663 DVDD.n3662 2.24964
R23977 DVDD.n3712 DVDD.n3664 2.24964
R23978 DVDD.n4752 DVDD.n3657 2.24964
R23979 DVDD.n4752 DVDD.n3717 2.24964
R23980 DVDD.n4752 DVDD.n3716 2.24964
R23981 DVDD.n3840 DVDD.n3827 2.24964
R23982 DVDD.n4079 DVDD.n4068 2.24964
R23983 DVDD.n3842 DVDD.n3827 2.24964
R23984 DVDD.n4079 DVDD.n4069 2.24964
R23985 DVDD.n3844 DVDD.n3827 2.24964
R23986 DVDD.n4079 DVDD.n4070 2.24964
R23987 DVDD.n3846 DVDD.n3827 2.24964
R23988 DVDD.n4079 DVDD.n4071 2.24964
R23989 DVDD.n3848 DVDD.n3827 2.24964
R23990 DVDD.n4079 DVDD.n4072 2.24964
R23991 DVDD.n3850 DVDD.n3827 2.24964
R23992 DVDD.n4079 DVDD.n4073 2.24964
R23993 DVDD.n3852 DVDD.n3827 2.24964
R23994 DVDD.n4079 DVDD.n4074 2.24964
R23995 DVDD.n3854 DVDD.n3827 2.24964
R23996 DVDD.n4079 DVDD.n4075 2.24964
R23997 DVDD.n3856 DVDD.n3827 2.24964
R23998 DVDD.n4079 DVDD.n4076 2.24964
R23999 DVDD.n3858 DVDD.n3827 2.24964
R24000 DVDD.n4079 DVDD.n4077 2.24964
R24001 DVDD.n3860 DVDD.n3827 2.24964
R24002 DVDD.n4079 DVDD.n4078 2.24964
R24003 DVDD.n4067 DVDD.n3827 2.24964
R24004 DVDD.n3894 DVDD.n3862 2.24964
R24005 DVDD.n3884 DVDD.n3863 2.24964
R24006 DVDD.n3894 DVDD.n3890 2.24964
R24007 DVDD.n3886 DVDD.n3863 2.24964
R24008 DVDD.n3894 DVDD.n3891 2.24964
R24009 DVDD.n3888 DVDD.n3863 2.24964
R24010 DVDD.n3894 DVDD.n3892 2.24964
R24011 DVDD.n3896 DVDD.n3863 2.24964
R24012 DVDD.n3895 DVDD.n3894 2.24964
R24013 DVDD.n3877 DVDD.n3863 2.24964
R24014 DVDD.n18865 DVDD.n18831 2.24964
R24015 DVDD.n18854 DVDD.n18832 2.24964
R24016 DVDD.n18865 DVDD.n18864 2.24964
R24017 DVDD.n18856 DVDD.n18832 2.24964
R24018 DVDD.n18865 DVDD.n18863 2.24964
R24019 DVDD.n18865 DVDD.n18862 2.24964
R24020 DVDD.n18849 DVDD.n18832 2.24964
R24021 DVDD.n3663 DVDD.n3661 2.24964
R24022 DVDD.n3663 DVDD.n3660 2.24964
R24023 DVDD.n3663 DVDD.n3659 2.24964
R24024 DVDD.n3712 DVDD.n3710 2.24964
R24025 DVDD.n3481 DVDD.n3480 2.24964
R24026 DVDD.n16043 DVDD.n3109 2.24964
R24027 DVDD.n3131 DVDD.n3109 2.24964
R24028 DVDD.n16052 DVDD.n3109 2.24964
R24029 DVDD.n9813 DVDD.n9757 2.24964
R24030 DVDD.n9939 DVDD.n9815 2.24964
R24031 DVDD.n9939 DVDD.n9756 2.24964
R24032 DVDD.n18702 DVDD.n18672 2.24964
R24033 DVDD.n18708 DVDD.n18707 2.24964
R24034 DVDD.n18692 DVDD.n18674 2.24964
R24035 DVDD.n18708 DVDD.n18706 2.24964
R24036 DVDD.n18708 DVDD.n18705 2.24964
R24037 DVDD.n18695 DVDD.n18674 2.24964
R24038 DVDD.n18708 DVDD.n18704 2.24964
R24039 DVDD.n18697 DVDD.n18674 2.24964
R24040 DVDD.n21088 DVDD.n21086 2.24964
R24041 DVDD.n21094 DVDD.n21091 2.24964
R24042 DVDD.n21088 DVDD.n21087 2.24964
R24043 DVDD.n21094 DVDD.n21090 2.24964
R24044 DVDD.n21088 DVDD.n21085 2.24964
R24045 DVDD.n21094 DVDD.n21092 2.24964
R24046 DVDD.n21088 DVDD.n21084 2.24964
R24047 DVDD.n21094 DVDD.n21093 2.24964
R24048 DVDD.n22253 DVDD.n94 2.24964
R24049 DVDD.n22245 DVDD.n106 2.24964
R24050 DVDD.n22253 DVDD.n95 2.24964
R24051 DVDD.n115 DVDD.n106 2.24964
R24052 DVDD.n22253 DVDD.n92 2.24964
R24053 DVDD.n22247 DVDD.n106 2.24964
R24054 DVDD.n22253 DVDD.n91 2.24964
R24055 DVDD.n22249 DVDD.n106 2.24964
R24056 DVDD.n48 DVDD.n42 2.24964
R24057 DVDD.n71 DVDD.n68 2.24964
R24058 DVDD.n50 DVDD.n42 2.24964
R24059 DVDD.n71 DVDD.n67 2.24964
R24060 DVDD.n53 DVDD.n42 2.24964
R24061 DVDD.n71 DVDD.n69 2.24964
R24062 DVDD.n55 DVDD.n42 2.24964
R24063 DVDD.n71 DVDD.n70 2.24964
R24064 DVDD.n3940 DVDD.n3939 2.24953
R24065 DVDD.n3971 DVDD.n3967 2.24953
R24066 DVDD.n3940 DVDD.n3938 2.24953
R24067 DVDD.n3971 DVDD.n3968 2.24953
R24068 DVDD.n3940 DVDD.n3937 2.24953
R24069 DVDD.n3971 DVDD.n3969 2.24953
R24070 DVDD.n3940 DVDD.n3936 2.24953
R24071 DVDD.n3971 DVDD.n3970 2.24953
R24072 DVDD.n3940 DVDD.n3935 2.24953
R24073 DVDD.n3971 DVDD.n3921 2.24953
R24074 DVDD.n4834 DVDD.n4824 2.24953
R24075 DVDD.n4804 DVDD.n3552 2.24953
R24076 DVDD.n4834 DVDD.n4825 2.24953
R24077 DVDD.n4806 DVDD.n3552 2.24953
R24078 DVDD.n4834 DVDD.n4826 2.24953
R24079 DVDD.n4808 DVDD.n3552 2.24953
R24080 DVDD.n4834 DVDD.n4827 2.24953
R24081 DVDD.n4810 DVDD.n3552 2.24953
R24082 DVDD.n4834 DVDD.n4828 2.24953
R24083 DVDD.n4812 DVDD.n3552 2.24953
R24084 DVDD.n4834 DVDD.n4829 2.24953
R24085 DVDD.n4814 DVDD.n3552 2.24953
R24086 DVDD.n4834 DVDD.n4830 2.24953
R24087 DVDD.n4816 DVDD.n3552 2.24953
R24088 DVDD.n4834 DVDD.n4831 2.24953
R24089 DVDD.n4818 DVDD.n3552 2.24953
R24090 DVDD.n4834 DVDD.n4832 2.24953
R24091 DVDD.n4820 DVDD.n3552 2.24953
R24092 DVDD.n4834 DVDD.n4833 2.24953
R24093 DVDD.n4822 DVDD.n3552 2.24953
R24094 DVDD.n4835 DVDD.n4834 2.24953
R24095 DVDD.n4836 DVDD.n3552 2.24953
R24096 DVDD.n4834 DVDD.n3551 2.24953
R24097 DVDD.n4843 DVDD.n3523 2.24953
R24098 DVDD.n4841 DVDD.n3538 2.24953
R24099 DVDD.n3546 DVDD.n3523 2.24953
R24100 DVDD.n4853 DVDD.n3538 2.24953
R24101 DVDD.n4855 DVDD.n3523 2.24953
R24102 DVDD.n3539 DVDD.n3538 2.24953
R24103 DVDD.n4868 DVDD.n3523 2.24953
R24104 DVDD.n4870 DVDD.n3538 2.24953
R24105 DVDD.n4872 DVDD.n3523 2.24953
R24106 DVDD.n3538 DVDD.n3522 2.24953
R24107 DVDD.n4896 DVDD.n4894 2.24953
R24108 DVDD.n4899 DVDD.n4898 2.24953
R24109 DVDD.n4896 DVDD.n4895 2.24953
R24110 DVDD.n4899 DVDD.n4897 2.24953
R24111 DVDD.n20602 DVDD.n20597 2.24953
R24112 DVDD.n20647 DVDD.n20646 2.24953
R24113 DVDD.n20602 DVDD.n20598 2.24953
R24114 DVDD.n20647 DVDD.n20645 2.24953
R24115 DVDD.n20602 DVDD.n20599 2.24953
R24116 DVDD.n20647 DVDD.n20644 2.24953
R24117 DVDD.n20602 DVDD.n20600 2.24953
R24118 DVDD.n20647 DVDD.n20643 2.24953
R24119 DVDD.n20602 DVDD.n20601 2.24953
R24120 DVDD.n20647 DVDD.n20603 2.24953
R24121 DVDD.n541 DVDD.n504 2.24953
R24122 DVDD.n18041 DVDD.n18040 2.24953
R24123 DVDD.n18038 DVDD.n504 2.24953
R24124 DVDD.n18040 DVDD.n503 2.24953
R24125 DVDD.n18054 DVDD.n18050 2.24953
R24126 DVDD.n18085 DVDD.n18083 2.24953
R24127 DVDD.n18054 DVDD.n18051 2.24953
R24128 DVDD.n18085 DVDD.n18082 2.24953
R24129 DVDD.n18057 DVDD.n18056 2.24953
R24130 DVDD.n18085 DVDD.n18081 2.24953
R24131 DVDD.n18054 DVDD.n18052 2.24953
R24132 DVDD.n18085 DVDD.n18080 2.24953
R24133 DVDD.n18054 DVDD.n18053 2.24953
R24134 DVDD.n18085 DVDD.n18055 2.24953
R24135 DVDD.n18194 DVDD.n18193 2.24953
R24136 DVDD.n18163 DVDD.n448 2.24953
R24137 DVDD.n18194 DVDD.n18192 2.24953
R24138 DVDD.n18165 DVDD.n448 2.24953
R24139 DVDD.n18194 DVDD.n18191 2.24953
R24140 DVDD.n18167 DVDD.n448 2.24953
R24141 DVDD.n18194 DVDD.n18190 2.24953
R24142 DVDD.n18169 DVDD.n448 2.24953
R24143 DVDD.n18194 DVDD.n18189 2.24953
R24144 DVDD.n18171 DVDD.n448 2.24953
R24145 DVDD.n18194 DVDD.n18188 2.24953
R24146 DVDD.n18173 DVDD.n448 2.24953
R24147 DVDD.n18194 DVDD.n18187 2.24953
R24148 DVDD.n18175 DVDD.n448 2.24953
R24149 DVDD.n18194 DVDD.n18186 2.24953
R24150 DVDD.n18177 DVDD.n448 2.24953
R24151 DVDD.n18194 DVDD.n18185 2.24953
R24152 DVDD.n18179 DVDD.n448 2.24953
R24153 DVDD.n18194 DVDD.n18184 2.24953
R24154 DVDD.n18181 DVDD.n448 2.24953
R24155 DVDD.n18195 DVDD.n18194 2.24953
R24156 DVDD.n18183 DVDD.n448 2.24953
R24157 DVDD.n18194 DVDD.n447 2.24953
R24158 DVDD.n22086 DVDD.n22081 2.24953
R24159 DVDD.n22114 DVDD.n22113 2.24953
R24160 DVDD.n22086 DVDD.n22082 2.24953
R24161 DVDD.n22114 DVDD.n22112 2.24953
R24162 DVDD.n22086 DVDD.n22083 2.24953
R24163 DVDD.n22114 DVDD.n22111 2.24953
R24164 DVDD.n22086 DVDD.n22084 2.24953
R24165 DVDD.n22114 DVDD.n22110 2.24953
R24166 DVDD.n22086 DVDD.n22085 2.24953
R24167 DVDD.n22114 DVDD.n22070 2.24953
R24168 DVDD.n18989 DVDD.n18985 2.24953
R24169 DVDD.n18995 DVDD.n18994 2.24953
R24170 DVDD.n18989 DVDD.n18986 2.24953
R24171 DVDD.n18995 DVDD.n18993 2.24953
R24172 DVDD.n18989 DVDD.n18987 2.24953
R24173 DVDD.n18995 DVDD.n18992 2.24953
R24174 DVDD.n18989 DVDD.n18988 2.24953
R24175 DVDD.n18995 DVDD.n18991 2.24953
R24176 DVDD.n18990 DVDD.n18989 2.24953
R24177 DVDD.n18995 DVDD.n18960 2.24953
R24178 DVDD.n22344 DVDD.n8 2.24953
R24179 DVDD.n22338 DVDD.n1 2.24953
R24180 DVDD.n22344 DVDD.n7 2.24953
R24181 DVDD.n22340 DVDD.n1 2.24953
R24182 DVDD.n22344 DVDD.n6 2.24953
R24183 DVDD.n19699 DVDD.n19697 2.24953
R24184 DVDD.n19211 DVDD.n19188 2.24953
R24185 DVDD.n19699 DVDD.n19698 2.24953
R24186 DVDD.n19213 DVDD.n19188 2.24953
R24187 DVDD.n19699 DVDD.n19187 2.24953
R24188 DVDD.n10 DVDD.n1 2.24953
R24189 DVDD.n22 DVDD.n21 2.24953
R24190 DVDD.n28 DVDD.n1 2.24953
R24191 DVDD.n19 DVDD.n4 2.24953
R24192 DVDD.n19202 DVDD.n19194 2.24953
R24193 DVDD.n19636 DVDD.n19193 2.24953
R24194 DVDD.n19637 DVDD.n19194 2.24953
R24195 DVDD.n19634 DVDD.n19193 2.24953
R24196 DVDD.n4404 DVDD.n4329 2.24926
R24197 DVDD.n4400 DVDD.n4329 2.24926
R24198 DVDD.n4262 DVDD.n4261 2.24926
R24199 DVDD.n4262 DVDD.n4260 2.24926
R24200 DVDD.n3751 DVDD.n3728 2.24926
R24201 DVDD.n4440 DVDD.n3728 2.24926
R24202 DVDD.n4845 DVDD.n4844 2.24926
R24203 DVDD.n18060 DVDD.n18045 2.24926
R24204 DVDD.n3666 DVDD.n3647 2.24926
R24205 DVDD.n3658 DVDD.n3641 2.24926
R24206 DVDD.n3977 DVDD.n3933 2.24901
R24207 DVDD.n22121 DVDD.n22080 2.24901
R24208 DVDD.n20855 DVDD.n18972 2.24901
R24209 DVDD.n3893 DVDD.n231 2.24901
R24210 DVDD.n29 DVDD.n5 2.24901
R24211 DVDD.n9688 DVDD.n9668 2.24901
R24212 DVDD.n9693 DVDD.n9668 2.24901
R24213 DVDD.n22159 DVDD.n296 2.24901
R24214 DVDD.n22159 DVDD.n292 2.24901
R24215 DVDD.n19047 DVDD.n19028 2.24901
R24216 DVDD.n19052 DVDD.n19028 2.24901
R24217 DVDD.n19937 DVDD.n19879 2.24901
R24218 DVDD.n19942 DVDD.n19879 2.24901
R24219 DVDD.n9955 DVDD.n9741 2.24901
R24220 DVDD.n9960 DVDD.n9741 2.24901
R24221 DVDD.n379 DVDD.n361 2.24901
R24222 DVDD.n384 DVDD.n361 2.24901
R24223 DVDD.n18896 DVDD.n18895 2.24901
R24224 DVDD.n18896 DVDD.n18894 2.24901
R24225 DVDD.n20374 DVDD.n20373 2.24901
R24226 DVDD.n20374 DVDD.n20372 2.24901
R24227 DVDD.n10094 DVDD.n9618 2.24901
R24228 DVDD.n10094 DVDD.n9614 2.24901
R24229 DVDD.n260 DVDD.n259 2.24901
R24230 DVDD.n268 DVDD.n260 2.24901
R24231 DVDD.n19142 DVDD.n19124 2.24901
R24232 DVDD.n19147 DVDD.n19124 2.24901
R24233 DVDD.n20024 DVDD.n19964 2.24901
R24234 DVDD.n20029 DVDD.n19964 2.24901
R24235 DVDD.n3928 DVDD.n3916 2.24901
R24236 DVDD.n5479 DVDD.n5468 2.24901
R24237 DVDD.n5484 DVDD.n5468 2.24901
R24238 DVDD.n20610 DVDD.n19703 2.24901
R24239 DVDD.n20615 DVDD.n19703 2.24901
R24240 DVDD.n20123 DVDD.n20065 2.24901
R24241 DVDD.n20128 DVDD.n20065 2.24901
R24242 DVDD.n808 DVDD.n807 2.24901
R24243 DVDD.n808 DVDD.n806 2.24901
R24244 DVDD.n22075 DVDD.n18199 2.24901
R24245 DVDD.n18981 DVDD.n18980 2.24901
R24246 DVDD.n18953 DVDD.n18952 2.24901
R24247 DVDD.n18953 DVDD.n18951 2.24901
R24248 DVDD.n9766 DVDD.n9610 2.24901
R24249 DVDD.n9771 DVDD.n9610 2.24901
R24250 DVDD.n4066 DVDD.n3866 2.24901
R24251 DVDD.n18841 DVDD.n18829 2.24901
R24252 DVDD.n18861 DVDD.n18829 2.24901
R24253 DVDD.n19748 DVDD.n19747 2.24901
R24254 DVDD.n19748 DVDD.n19746 2.24901
R24255 DVDD.n21214 DVDD.n18680 2.24901
R24256 DVDD.n21214 DVDD.n18673 2.24901
R24257 DVDD.n21098 DVDD.n18730 2.24901
R24258 DVDD.n21089 DVDD.n18730 2.24901
R24259 DVDD.n22244 DVDD.n120 2.24901
R24260 DVDD.n22244 DVDD.n119 2.24901
R24261 DVDD.n77 DVDD.n49 2.24901
R24262 DVDD.n72 DVDD.n49 2.24901
R24263 DVDD.n22337 DVDD.n22336 2.24901
R24264 DVDD.n19210 DVDD.n19209 2.24901
R24265 DVDD.n19210 DVDD.n19208 2.24901
R24266 DVDD.n17370 DVDD.n17308 2.24752
R24267 DVDD.n5740 DVDD.n5693 2.24752
R24268 DVDD.n17373 DVDD.n17307 2.24752
R24269 DVDD.n17372 DVDD.n17306 2.24752
R24270 DVDD.n17376 DVDD.n17307 2.24752
R24271 DVDD.n17375 DVDD.n17306 2.24752
R24272 DVDD.n17379 DVDD.n17307 2.24752
R24273 DVDD.n17378 DVDD.n17306 2.24752
R24274 DVDD.n17382 DVDD.n17307 2.24752
R24275 DVDD.n17381 DVDD.n17306 2.24752
R24276 DVDD.n17385 DVDD.n17307 2.24752
R24277 DVDD.n17384 DVDD.n17306 2.24752
R24278 DVDD.n17388 DVDD.n17307 2.24752
R24279 DVDD.n17387 DVDD.n17306 2.24752
R24280 DVDD.n17391 DVDD.n17307 2.24752
R24281 DVDD.n17390 DVDD.n17306 2.24752
R24282 DVDD.n17394 DVDD.n17307 2.24752
R24283 DVDD.n17393 DVDD.n17306 2.24752
R24284 DVDD.n17397 DVDD.n17307 2.24752
R24285 DVDD.n17396 DVDD.n17306 2.24752
R24286 DVDD.n17400 DVDD.n17307 2.24752
R24287 DVDD.n17399 DVDD.n17306 2.24752
R24288 DVDD.n17403 DVDD.n17307 2.24752
R24289 DVDD.n17402 DVDD.n17306 2.24752
R24290 DVDD.n17406 DVDD.n17307 2.24752
R24291 DVDD.n17405 DVDD.n17306 2.24752
R24292 DVDD.n17409 DVDD.n17307 2.24752
R24293 DVDD.n17408 DVDD.n17306 2.24752
R24294 DVDD.n17412 DVDD.n17307 2.24752
R24295 DVDD.n17411 DVDD.n17306 2.24752
R24296 DVDD.n17415 DVDD.n17307 2.24752
R24297 DVDD.n17414 DVDD.n17306 2.24752
R24298 DVDD.n17418 DVDD.n17307 2.24752
R24299 DVDD.n17417 DVDD.n17306 2.24752
R24300 DVDD.n17421 DVDD.n17307 2.24752
R24301 DVDD.n17420 DVDD.n17306 2.24752
R24302 DVDD.n17424 DVDD.n17307 2.24752
R24303 DVDD.n17423 DVDD.n17306 2.24752
R24304 DVDD.n17427 DVDD.n17307 2.24752
R24305 DVDD.n17426 DVDD.n17306 2.24752
R24306 DVDD.n17430 DVDD.n17307 2.24752
R24307 DVDD.n17429 DVDD.n17306 2.24752
R24308 DVDD.n17433 DVDD.n17307 2.24752
R24309 DVDD.n17432 DVDD.n17306 2.24752
R24310 DVDD.n17436 DVDD.n17307 2.24752
R24311 DVDD.n17435 DVDD.n17306 2.24752
R24312 DVDD.n17439 DVDD.n17307 2.24752
R24313 DVDD.n17438 DVDD.n17306 2.24752
R24314 DVDD.n17442 DVDD.n17307 2.24752
R24315 DVDD.n17441 DVDD.n17306 2.24752
R24316 DVDD.n17445 DVDD.n17307 2.24752
R24317 DVDD.n17444 DVDD.n17306 2.24752
R24318 DVDD.n17448 DVDD.n17307 2.24752
R24319 DVDD.n17447 DVDD.n17306 2.24752
R24320 DVDD.n17451 DVDD.n17307 2.24752
R24321 DVDD.n17450 DVDD.n17306 2.24752
R24322 DVDD.n17454 DVDD.n17307 2.24752
R24323 DVDD.n17453 DVDD.n17306 2.24752
R24324 DVDD.n17457 DVDD.n17307 2.24752
R24325 DVDD.n17456 DVDD.n17306 2.24752
R24326 DVDD.n17460 DVDD.n17307 2.24752
R24327 DVDD.n17459 DVDD.n17306 2.24752
R24328 DVDD.n17463 DVDD.n17307 2.24752
R24329 DVDD.n17462 DVDD.n17306 2.24752
R24330 DVDD.n17466 DVDD.n17307 2.24752
R24331 DVDD.n17465 DVDD.n17306 2.24752
R24332 DVDD.n17469 DVDD.n17307 2.24752
R24333 DVDD.n17468 DVDD.n17306 2.24752
R24334 DVDD.n17472 DVDD.n17307 2.24752
R24335 DVDD.n17471 DVDD.n17306 2.24752
R24336 DVDD.n17475 DVDD.n17307 2.24752
R24337 DVDD.n17474 DVDD.n17306 2.24752
R24338 DVDD.n17478 DVDD.n17307 2.24752
R24339 DVDD.n17477 DVDD.n17306 2.24752
R24340 DVDD.n17481 DVDD.n17307 2.24752
R24341 DVDD.n17480 DVDD.n17306 2.24752
R24342 DVDD.n17484 DVDD.n17307 2.24752
R24343 DVDD.n17483 DVDD.n17306 2.24752
R24344 DVDD.n17487 DVDD.n17307 2.24752
R24345 DVDD.n17486 DVDD.n17306 2.24752
R24346 DVDD.n17490 DVDD.n17307 2.24752
R24347 DVDD.n17489 DVDD.n17306 2.24752
R24348 DVDD.n17493 DVDD.n17307 2.24752
R24349 DVDD.n17492 DVDD.n17306 2.24752
R24350 DVDD.n17496 DVDD.n17307 2.24752
R24351 DVDD.n17495 DVDD.n17306 2.24752
R24352 DVDD.n17499 DVDD.n17307 2.24752
R24353 DVDD.n17498 DVDD.n17306 2.24752
R24354 DVDD.n17502 DVDD.n17307 2.24752
R24355 DVDD.n17501 DVDD.n17306 2.24752
R24356 DVDD.n17505 DVDD.n17307 2.24752
R24357 DVDD.n17504 DVDD.n17306 2.24752
R24358 DVDD.n17508 DVDD.n17307 2.24752
R24359 DVDD.n17507 DVDD.n17306 2.24752
R24360 DVDD.n17511 DVDD.n17307 2.24752
R24361 DVDD.n17510 DVDD.n17306 2.24752
R24362 DVDD.n17514 DVDD.n17307 2.24752
R24363 DVDD.n17513 DVDD.n17306 2.24752
R24364 DVDD.n5988 DVDD.n5937 2.24752
R24365 DVDD.n17364 DVDD.n17363 2.24752
R24366 DVDD.n5989 DVDD.n5988 2.24752
R24367 DVDD.n17365 DVDD.n17364 2.24752
R24368 DVDD.n5986 DVDD.n5590 2.24752
R24369 DVDD.n5740 DVDD.n5591 2.24752
R24370 DVDD.n5986 DVDD.n5985 2.24752
R24371 DVDD.n5740 DVDD.n5694 2.24752
R24372 DVDD.n5986 DVDD.n5984 2.24752
R24373 DVDD.n5740 DVDD.n5695 2.24752
R24374 DVDD.n5986 DVDD.n5983 2.24752
R24375 DVDD.n5740 DVDD.n5696 2.24752
R24376 DVDD.n5986 DVDD.n5982 2.24752
R24377 DVDD.n5740 DVDD.n5697 2.24752
R24378 DVDD.n5986 DVDD.n5981 2.24752
R24379 DVDD.n5740 DVDD.n5698 2.24752
R24380 DVDD.n5986 DVDD.n5980 2.24752
R24381 DVDD.n5740 DVDD.n5699 2.24752
R24382 DVDD.n5986 DVDD.n5979 2.24752
R24383 DVDD.n5740 DVDD.n5700 2.24752
R24384 DVDD.n5986 DVDD.n5978 2.24752
R24385 DVDD.n5740 DVDD.n5701 2.24752
R24386 DVDD.n5986 DVDD.n5977 2.24752
R24387 DVDD.n5740 DVDD.n5702 2.24752
R24388 DVDD.n5986 DVDD.n5976 2.24752
R24389 DVDD.n5740 DVDD.n5703 2.24752
R24390 DVDD.n5986 DVDD.n5975 2.24752
R24391 DVDD.n5740 DVDD.n5704 2.24752
R24392 DVDD.n5986 DVDD.n5974 2.24752
R24393 DVDD.n5740 DVDD.n5705 2.24752
R24394 DVDD.n5986 DVDD.n5973 2.24752
R24395 DVDD.n5740 DVDD.n5706 2.24752
R24396 DVDD.n5986 DVDD.n5972 2.24752
R24397 DVDD.n5740 DVDD.n5707 2.24752
R24398 DVDD.n5986 DVDD.n5971 2.24752
R24399 DVDD.n5740 DVDD.n5708 2.24752
R24400 DVDD.n5986 DVDD.n5970 2.24752
R24401 DVDD.n5740 DVDD.n5709 2.24752
R24402 DVDD.n5986 DVDD.n5969 2.24752
R24403 DVDD.n5740 DVDD.n5710 2.24752
R24404 DVDD.n5986 DVDD.n5968 2.24752
R24405 DVDD.n5740 DVDD.n5711 2.24752
R24406 DVDD.n5986 DVDD.n5967 2.24752
R24407 DVDD.n5740 DVDD.n5712 2.24752
R24408 DVDD.n5986 DVDD.n5966 2.24752
R24409 DVDD.n5740 DVDD.n5713 2.24752
R24410 DVDD.n5986 DVDD.n5965 2.24752
R24411 DVDD.n5740 DVDD.n5714 2.24752
R24412 DVDD.n5986 DVDD.n5964 2.24752
R24413 DVDD.n5740 DVDD.n5715 2.24752
R24414 DVDD.n5986 DVDD.n5963 2.24752
R24415 DVDD.n5740 DVDD.n5716 2.24752
R24416 DVDD.n5986 DVDD.n5962 2.24752
R24417 DVDD.n5740 DVDD.n5717 2.24752
R24418 DVDD.n5986 DVDD.n5961 2.24752
R24419 DVDD.n5740 DVDD.n5718 2.24752
R24420 DVDD.n5986 DVDD.n5960 2.24752
R24421 DVDD.n5740 DVDD.n5719 2.24752
R24422 DVDD.n5986 DVDD.n5959 2.24752
R24423 DVDD.n5740 DVDD.n5720 2.24752
R24424 DVDD.n5986 DVDD.n5958 2.24752
R24425 DVDD.n5740 DVDD.n5721 2.24752
R24426 DVDD.n5986 DVDD.n5957 2.24752
R24427 DVDD.n5740 DVDD.n5722 2.24752
R24428 DVDD.n5986 DVDD.n5956 2.24752
R24429 DVDD.n5740 DVDD.n5723 2.24752
R24430 DVDD.n5986 DVDD.n5955 2.24752
R24431 DVDD.n5740 DVDD.n5724 2.24752
R24432 DVDD.n5986 DVDD.n5954 2.24752
R24433 DVDD.n5740 DVDD.n5725 2.24752
R24434 DVDD.n5986 DVDD.n5953 2.24752
R24435 DVDD.n5740 DVDD.n5726 2.24752
R24436 DVDD.n5986 DVDD.n5952 2.24752
R24437 DVDD.n5740 DVDD.n5727 2.24752
R24438 DVDD.n5986 DVDD.n5951 2.24752
R24439 DVDD.n5740 DVDD.n5728 2.24752
R24440 DVDD.n5986 DVDD.n5950 2.24752
R24441 DVDD.n5740 DVDD.n5729 2.24752
R24442 DVDD.n5986 DVDD.n5949 2.24752
R24443 DVDD.n5740 DVDD.n5730 2.24752
R24444 DVDD.n5986 DVDD.n5948 2.24752
R24445 DVDD.n5740 DVDD.n5731 2.24752
R24446 DVDD.n5986 DVDD.n5947 2.24752
R24447 DVDD.n5740 DVDD.n5732 2.24752
R24448 DVDD.n5986 DVDD.n5946 2.24752
R24449 DVDD.n5740 DVDD.n5733 2.24752
R24450 DVDD.n5986 DVDD.n5945 2.24752
R24451 DVDD.n5740 DVDD.n5734 2.24752
R24452 DVDD.n5986 DVDD.n5944 2.24752
R24453 DVDD.n5740 DVDD.n5735 2.24752
R24454 DVDD.n5986 DVDD.n5943 2.24752
R24455 DVDD.n5740 DVDD.n5736 2.24752
R24456 DVDD.n5986 DVDD.n5942 2.24752
R24457 DVDD.n5740 DVDD.n5737 2.24752
R24458 DVDD.n5986 DVDD.n5941 2.24752
R24459 DVDD.n5740 DVDD.n5738 2.24752
R24460 DVDD.n5986 DVDD.n5940 2.24752
R24461 DVDD.n5740 DVDD.n5739 2.24752
R24462 DVDD.n5986 DVDD.n5939 2.24752
R24463 DVDD.n5986 DVDD.n5692 2.24752
R24464 DVDD.n17723 DVDD.n17722 2.24752
R24465 DVDD.n15138 DVDD.n15137 2.24752
R24466 DVDD.n17723 DVDD.n895 2.24752
R24467 DVDD.n15138 DVDD.n5581 2.24752
R24468 DVDD.n4534 DVDD.n4388 2.24712
R24469 DVDD.n899 DVDD.n892 2.24681
R24470 DVDD.n5587 DVDD.n5579 2.24681
R24471 DVDD.n5585 DVDD.n5580 2.24681
R24472 DVDD.n4953 DVDD.n3396 2.24442
R24473 DVDD.n4956 DVDD.n3396 2.24442
R24474 DVDD.n4959 DVDD.n3396 2.24442
R24475 DVDD.n4962 DVDD.n3396 2.24442
R24476 DVDD.n4965 DVDD.n3396 2.24442
R24477 DVDD.n4968 DVDD.n3396 2.24442
R24478 DVDD.n4971 DVDD.n3396 2.24442
R24479 DVDD.n4974 DVDD.n3396 2.24442
R24480 DVDD.n4943 DVDD.n3396 2.24442
R24481 DVDD.n16396 DVDD.n2295 2.24442
R24482 DVDD.n16396 DVDD.n2333 2.24442
R24483 DVDD.n16396 DVDD.n2332 2.24442
R24484 DVDD.n16396 DVDD.n2331 2.24442
R24485 DVDD.n16396 DVDD.n2330 2.24442
R24486 DVDD.n16396 DVDD.n2329 2.24442
R24487 DVDD.n16396 DVDD.n2328 2.24442
R24488 DVDD.n16396 DVDD.n2327 2.24442
R24489 DVDD.n16396 DVDD.n2326 2.24442
R24490 DVDD.n2475 DVDD.n2446 2.24442
R24491 DVDD.n2475 DVDD.n2445 2.24442
R24492 DVDD.n2475 DVDD.n2444 2.24442
R24493 DVDD.n2475 DVDD.n2443 2.24442
R24494 DVDD.n2475 DVDD.n2442 2.24442
R24495 DVDD.n2475 DVDD.n2441 2.24442
R24496 DVDD.n2475 DVDD.n2440 2.24442
R24497 DVDD.n2475 DVDD.n2439 2.24442
R24498 DVDD.n2475 DVDD.n2438 2.24442
R24499 DVDD.n4942 DVDD.n3370 2.24442
R24500 DVDD.n4954 DVDD.n3370 2.24442
R24501 DVDD.n4957 DVDD.n3370 2.24442
R24502 DVDD.n4960 DVDD.n3370 2.24442
R24503 DVDD.n4963 DVDD.n3370 2.24442
R24504 DVDD.n4966 DVDD.n3370 2.24442
R24505 DVDD.n4969 DVDD.n3370 2.24442
R24506 DVDD.n4972 DVDD.n3370 2.24442
R24507 DVDD.n4975 DVDD.n3370 2.24442
R24508 DVDD.n2307 DVDD.n2294 2.24442
R24509 DVDD.n2309 DVDD.n2294 2.24442
R24510 DVDD.n2311 DVDD.n2294 2.24442
R24511 DVDD.n2313 DVDD.n2294 2.24442
R24512 DVDD.n2315 DVDD.n2294 2.24442
R24513 DVDD.n2317 DVDD.n2294 2.24442
R24514 DVDD.n2319 DVDD.n2294 2.24442
R24515 DVDD.n2321 DVDD.n2294 2.24442
R24516 DVDD.n2323 DVDD.n2294 2.24442
R24517 DVDD.n2457 DVDD.n2413 2.24442
R24518 DVDD.n2459 DVDD.n2413 2.24442
R24519 DVDD.n2461 DVDD.n2413 2.24442
R24520 DVDD.n2463 DVDD.n2413 2.24442
R24521 DVDD.n2465 DVDD.n2413 2.24442
R24522 DVDD.n2467 DVDD.n2413 2.24442
R24523 DVDD.n2469 DVDD.n2413 2.24442
R24524 DVDD.n2471 DVDD.n2413 2.24442
R24525 DVDD.n2447 DVDD.n2413 2.24442
R24526 DVDD.n5002 DVDD.n4984 2.24442
R24527 DVDD.n5002 DVDD.n4983 2.24442
R24528 DVDD.n4992 DVDD.n4991 2.24442
R24529 DVDD.n4997 DVDD.n4986 2.24442
R24530 DVDD.n4997 DVDD.n4993 2.24442
R24531 DVDD.n4998 DVDD.n4997 2.24442
R24532 DVDD.n4994 DVDD.n4987 2.24442
R24533 DVDD.n15143 DVDD.n5562 2.24442
R24534 DVDD.n15144 DVDD.n5576 2.24442
R24535 DVDD.n15144 DVDD.n5571 2.24442
R24536 DVDD.n10222 DVDD.n8958 2.24442
R24537 DVDD.n10222 DVDD.n8957 2.24442
R24538 DVDD.n10222 DVDD.n8956 2.24442
R24539 DVDD.n10222 DVDD.n8955 2.24442
R24540 DVDD.n10222 DVDD.n8954 2.24442
R24541 DVDD.n10222 DVDD.n8953 2.24442
R24542 DVDD.n10222 DVDD.n8952 2.24442
R24543 DVDD.n10222 DVDD.n8951 2.24442
R24544 DVDD.n16405 DVDD.n2281 2.24442
R24545 DVDD.n16408 DVDD.n2281 2.24442
R24546 DVDD.n16411 DVDD.n2281 2.24442
R24547 DVDD.n16414 DVDD.n2281 2.24442
R24548 DVDD.n16417 DVDD.n2281 2.24442
R24549 DVDD.n16420 DVDD.n2281 2.24442
R24550 DVDD.n16423 DVDD.n2281 2.24442
R24551 DVDD.n16427 DVDD.n2281 2.24442
R24552 DVDD.n16451 DVDD.n2264 2.24442
R24553 DVDD.n16451 DVDD.n2263 2.24442
R24554 DVDD.n16451 DVDD.n2262 2.24442
R24555 DVDD.n16451 DVDD.n2261 2.24442
R24556 DVDD.n16451 DVDD.n2260 2.24442
R24557 DVDD.n16451 DVDD.n2259 2.24442
R24558 DVDD.n16451 DVDD.n2258 2.24442
R24559 DVDD.n16451 DVDD.n2257 2.24442
R24560 DVDD.n5566 DVDD.n5561 2.24442
R24561 DVDD.n5567 DVDD.n5564 2.24442
R24562 DVDD.n5573 DVDD.n5564 2.24442
R24563 DVDD.n5569 DVDD.n5564 2.24442
R24564 DVDD.n10205 DVDD.n8960 2.24442
R24565 DVDD.n10207 DVDD.n8960 2.24442
R24566 DVDD.n10209 DVDD.n8960 2.24442
R24567 DVDD.n10211 DVDD.n8960 2.24442
R24568 DVDD.n10213 DVDD.n8960 2.24442
R24569 DVDD.n10215 DVDD.n8960 2.24442
R24570 DVDD.n10217 DVDD.n8960 2.24442
R24571 DVDD.n16407 DVDD.n2279 2.24442
R24572 DVDD.n16410 DVDD.n2279 2.24442
R24573 DVDD.n16413 DVDD.n2279 2.24442
R24574 DVDD.n16416 DVDD.n2279 2.24442
R24575 DVDD.n16419 DVDD.n2279 2.24442
R24576 DVDD.n16422 DVDD.n2279 2.24442
R24577 DVDD.n16425 DVDD.n2279 2.24442
R24578 DVDD.n16434 DVDD.n2267 2.24442
R24579 DVDD.n16436 DVDD.n2267 2.24442
R24580 DVDD.n16438 DVDD.n2267 2.24442
R24581 DVDD.n16440 DVDD.n2267 2.24442
R24582 DVDD.n16442 DVDD.n2267 2.24442
R24583 DVDD.n16444 DVDD.n2267 2.24442
R24584 DVDD.n16446 DVDD.n2267 2.24442
R24585 DVDD.n10220 DVDD.n10219 2.24442
R24586 DVDD.n16431 DVDD.n16430 2.24442
R24587 DVDD.n16449 DVDD.n16448 2.24442
R24588 DVDD.n17734 DVDD.n887 2.24442
R24589 DVDD.n17735 DVDD.n17734 2.24442
R24590 DVDD.n17731 DVDD.n889 2.24442
R24591 DVDD.n17732 DVDD.n884 2.24442
R24592 DVDD.n884 DVDD.n883 2.24442
R24593 DVDD.n17729 DVDD.n886 2.24442
R24594 DVDD.n17737 DVDD.n881 2.24442
R24595 DVDD.n18027 DVDD.n18026 2.24442
R24596 DVDD.n18029 DVDD.n18027 2.24442
R24597 DVDD.n18034 DVDD.n18033 2.24442
R24598 DVDD.n18032 DVDD.n547 2.24442
R24599 DVDD.n18032 DVDD.n548 2.24442
R24600 DVDD.n546 DVDD.n545 2.24442
R24601 DVDD.n18032 DVDD.n18031 2.24442
R24602 DVDD.n10176 DVDD.n9572 2.24442
R24603 DVDD.n10179 DVDD.n9572 2.24442
R24604 DVDD.n10182 DVDD.n9572 2.24442
R24605 DVDD.n10185 DVDD.n9572 2.24442
R24606 DVDD.n10188 DVDD.n9572 2.24442
R24607 DVDD.n10191 DVDD.n9572 2.24442
R24608 DVDD.n10194 DVDD.n9572 2.24442
R24609 DVDD.n10198 DVDD.n9572 2.24442
R24610 DVDD.n10178 DVDD.n8972 2.24442
R24611 DVDD.n10181 DVDD.n8972 2.24442
R24612 DVDD.n10184 DVDD.n8972 2.24442
R24613 DVDD.n10187 DVDD.n8972 2.24442
R24614 DVDD.n10190 DVDD.n8972 2.24442
R24615 DVDD.n10193 DVDD.n8972 2.24442
R24616 DVDD.n10196 DVDD.n8972 2.24442
R24617 DVDD.n10202 DVDD.n10201 2.24442
R24618 DVDD.n4907 DVDD.n3488 2.24442
R24619 DVDD.n4918 DVDD.n3488 2.24442
R24620 DVDD.n4921 DVDD.n3488 2.24442
R24621 DVDD.n4924 DVDD.n3488 2.24442
R24622 DVDD.n4927 DVDD.n3488 2.24442
R24623 DVDD.n4930 DVDD.n3488 2.24442
R24624 DVDD.n4933 DVDD.n3488 2.24442
R24625 DVDD.n4936 DVDD.n3488 2.24442
R24626 DVDD.n4939 DVDD.n3488 2.24442
R24627 DVDD.n4917 DVDD.n3473 2.24442
R24628 DVDD.n4920 DVDD.n3473 2.24442
R24629 DVDD.n4923 DVDD.n3473 2.24442
R24630 DVDD.n4926 DVDD.n3473 2.24442
R24631 DVDD.n4929 DVDD.n3473 2.24442
R24632 DVDD.n4932 DVDD.n3473 2.24442
R24633 DVDD.n4935 DVDD.n3473 2.24442
R24634 DVDD.n4938 DVDD.n3473 2.24442
R24635 DVDD.n4941 DVDD.n3473 2.24442
R24636 DVDD.n18800 DVDD.n104 2.24344
R24637 DVDD.n18793 DVDD.n104 2.24344
R24638 DVDD.n18803 DVDD.n104 2.24344
R24639 DVDD.n18806 DVDD.n104 2.24344
R24640 DVDD.n18809 DVDD.n104 2.24344
R24641 DVDD.n18812 DVDD.n104 2.24344
R24642 DVDD.n18815 DVDD.n104 2.24344
R24643 DVDD.n18798 DVDD.n97 2.24344
R24644 DVDD.n18802 DVDD.n97 2.24344
R24645 DVDD.n18805 DVDD.n97 2.24344
R24646 DVDD.n18808 DVDD.n97 2.24344
R24647 DVDD.n18811 DVDD.n97 2.24344
R24648 DVDD.n18814 DVDD.n97 2.24344
R24649 DVDD.n18817 DVDD.n97 2.24344
R24650 DVDD.n21051 DVDD.n18795 2.24344
R24651 DVDD.n20464 DVDD.n19816 2.24344
R24652 DVDD.n20464 DVDD.n19815 2.24344
R24653 DVDD.n20464 DVDD.n19814 2.24344
R24654 DVDD.n20464 DVDD.n19813 2.24344
R24655 DVDD.n20464 DVDD.n19812 2.24344
R24656 DVDD.n20464 DVDD.n19811 2.24344
R24657 DVDD.n20449 DVDD.n19820 2.24344
R24658 DVDD.n20451 DVDD.n19820 2.24344
R24659 DVDD.n20453 DVDD.n19820 2.24344
R24660 DVDD.n20455 DVDD.n19820 2.24344
R24661 DVDD.n20457 DVDD.n19820 2.24344
R24662 DVDD.n20459 DVDD.n19820 2.24344
R24663 DVDD.n20462 DVDD.n20461 2.24344
R24664 DVDD.n21026 DVDD.n66 2.24344
R24665 DVDD.n21029 DVDD.n66 2.24344
R24666 DVDD.n21032 DVDD.n66 2.24344
R24667 DVDD.n21035 DVDD.n66 2.24344
R24668 DVDD.n21038 DVDD.n66 2.24344
R24669 DVDD.n21041 DVDD.n66 2.24344
R24670 DVDD.n21046 DVDD.n66 2.24344
R24671 DVDD.n18818 DVDD.n57 2.24344
R24672 DVDD.n21028 DVDD.n57 2.24344
R24673 DVDD.n21031 DVDD.n57 2.24344
R24674 DVDD.n21034 DVDD.n57 2.24344
R24675 DVDD.n21037 DVDD.n57 2.24344
R24676 DVDD.n21040 DVDD.n57 2.24344
R24677 DVDD.n21043 DVDD.n57 2.24344
R24678 DVDD.n21045 DVDD.n57 2.24344
R24679 DVDD.n20922 DVDD.n18910 2.24344
R24680 DVDD.n20922 DVDD.n18911 2.24344
R24681 DVDD.n20922 DVDD.n18912 2.24344
R24682 DVDD.n20922 DVDD.n18913 2.24344
R24683 DVDD.n20922 DVDD.n18914 2.24344
R24684 DVDD.n20922 DVDD.n18915 2.24344
R24685 DVDD.n20922 DVDD.n20921 2.24344
R24686 DVDD.n20907 DVDD.n18908 2.24344
R24687 DVDD.n20909 DVDD.n18908 2.24344
R24688 DVDD.n20911 DVDD.n18908 2.24344
R24689 DVDD.n20913 DVDD.n18908 2.24344
R24690 DVDD.n20915 DVDD.n18908 2.24344
R24691 DVDD.n20917 DVDD.n18908 2.24344
R24692 DVDD.n18918 DVDD.n18908 2.24344
R24693 DVDD.n18916 DVDD.n18908 2.24344
R24694 DVDD.n21083 DVDD.n18750 2.24344
R24695 DVDD.n21083 DVDD.n18749 2.24344
R24696 DVDD.n21083 DVDD.n18748 2.24344
R24697 DVDD.n21083 DVDD.n18747 2.24344
R24698 DVDD.n21083 DVDD.n18746 2.24344
R24699 DVDD.n21083 DVDD.n18745 2.24344
R24700 DVDD.n21083 DVDD.n18744 2.24344
R24701 DVDD.n21067 DVDD.n18735 2.24344
R24702 DVDD.n21069 DVDD.n18735 2.24344
R24703 DVDD.n21071 DVDD.n18735 2.24344
R24704 DVDD.n21073 DVDD.n18735 2.24344
R24705 DVDD.n21075 DVDD.n18735 2.24344
R24706 DVDD.n21077 DVDD.n18735 2.24344
R24707 DVDD.n21079 DVDD.n18735 2.24344
R24708 DVDD.n20538 DVDD.n19796 2.24344
R24709 DVDD.n20538 DVDD.n19795 2.24344
R24710 DVDD.n20538 DVDD.n19794 2.24344
R24711 DVDD.n20538 DVDD.n19793 2.24344
R24712 DVDD.n20538 DVDD.n19792 2.24344
R24713 DVDD.n20538 DVDD.n19791 2.24344
R24714 DVDD.n19788 DVDD.n19787 2.24344
R24715 DVDD.n19788 DVDD.n19786 2.24344
R24716 DVDD.n19788 DVDD.n19785 2.24344
R24717 DVDD.n19788 DVDD.n19784 2.24344
R24718 DVDD.n19788 DVDD.n19783 2.24344
R24719 DVDD.n19788 DVDD.n19782 2.24344
R24720 DVDD.n20540 DVDD.n19780 2.24344
R24721 DVDD.n21010 DVDD.n18703 2.24344
R24722 DVDD.n20993 DVDD.n18703 2.24344
R24723 DVDD.n20996 DVDD.n18703 2.24344
R24724 DVDD.n20999 DVDD.n18703 2.24344
R24725 DVDD.n21002 DVDD.n18703 2.24344
R24726 DVDD.n21005 DVDD.n18703 2.24344
R24727 DVDD.n21008 DVDD.n18703 2.24344
R24728 DVDD.n20990 DVDD.n18699 2.24344
R24729 DVDD.n20992 DVDD.n18699 2.24344
R24730 DVDD.n20995 DVDD.n18699 2.24344
R24731 DVDD.n20998 DVDD.n18699 2.24344
R24732 DVDD.n21001 DVDD.n18699 2.24344
R24733 DVDD.n21004 DVDD.n18699 2.24344
R24734 DVDD.n21007 DVDD.n18699 2.24344
R24735 DVDD.n20519 DVDD.n20518 2.24344
R24736 DVDD.n20519 DVDD.n20494 2.24344
R24737 DVDD.n20519 DVDD.n20493 2.24344
R24738 DVDD.n20519 DVDD.n20492 2.24344
R24739 DVDD.n20519 DVDD.n20491 2.24344
R24740 DVDD.n20519 DVDD.n20490 2.24344
R24741 DVDD.n20519 DVDD.n20489 2.24344
R24742 DVDD.n20497 DVDD.n20487 2.24344
R24743 DVDD.n20504 DVDD.n20487 2.24344
R24744 DVDD.n20506 DVDD.n20487 2.24344
R24745 DVDD.n20508 DVDD.n20487 2.24344
R24746 DVDD.n20510 DVDD.n20487 2.24344
R24747 DVDD.n20512 DVDD.n20487 2.24344
R24748 DVDD.n20514 DVDD.n20487 2.24344
R24749 DVDD.n20495 DVDD.n20487 2.24344
R24750 DVDD.n18823 DVDD.n18699 2.24344
R24751 DVDD.n1605 DVDD.n1604 2.24164
R24752 DVDD.n1313 DVDD.n1262 2.24164
R24753 DVDD.n1605 DVDD.n1311 2.24164
R24754 DVDD.n1595 DVDD.n1262 2.24164
R24755 DVDD.n1605 DVDD.n1310 2.24164
R24756 DVDD.n1590 DVDD.n1262 2.24164
R24757 DVDD.n1605 DVDD.n1309 2.24164
R24758 DVDD.n1583 DVDD.n1262 2.24164
R24759 DVDD.n1605 DVDD.n1308 2.24164
R24760 DVDD.n1578 DVDD.n1262 2.24164
R24761 DVDD.n1605 DVDD.n1307 2.24164
R24762 DVDD.n1571 DVDD.n1262 2.24164
R24763 DVDD.n1605 DVDD.n1306 2.24164
R24764 DVDD.n1566 DVDD.n1262 2.24164
R24765 DVDD.n1605 DVDD.n1305 2.24164
R24766 DVDD.n1559 DVDD.n1262 2.24164
R24767 DVDD.n1605 DVDD.n1304 2.24164
R24768 DVDD.n1554 DVDD.n1262 2.24164
R24769 DVDD.n1605 DVDD.n1303 2.24164
R24770 DVDD.n1547 DVDD.n1262 2.24164
R24771 DVDD.n1605 DVDD.n1302 2.24164
R24772 DVDD.n1542 DVDD.n1262 2.24164
R24773 DVDD.n1605 DVDD.n1301 2.24164
R24774 DVDD.n1535 DVDD.n1262 2.24164
R24775 DVDD.n1605 DVDD.n1300 2.24164
R24776 DVDD.n1530 DVDD.n1262 2.24164
R24777 DVDD.n1605 DVDD.n1299 2.24164
R24778 DVDD.n1523 DVDD.n1262 2.24164
R24779 DVDD.n1605 DVDD.n1298 2.24164
R24780 DVDD.n1518 DVDD.n1262 2.24164
R24781 DVDD.n1605 DVDD.n1297 2.24164
R24782 DVDD.n1511 DVDD.n1262 2.24164
R24783 DVDD.n1605 DVDD.n1296 2.24164
R24784 DVDD.n1506 DVDD.n1262 2.24164
R24785 DVDD.n1605 DVDD.n1295 2.24164
R24786 DVDD.n1499 DVDD.n1262 2.24164
R24787 DVDD.n1605 DVDD.n1294 2.24164
R24788 DVDD.n1494 DVDD.n1262 2.24164
R24789 DVDD.n1605 DVDD.n1293 2.24164
R24790 DVDD.n1487 DVDD.n1262 2.24164
R24791 DVDD.n1605 DVDD.n1292 2.24164
R24792 DVDD.n1482 DVDD.n1262 2.24164
R24793 DVDD.n1605 DVDD.n1291 2.24164
R24794 DVDD.n1475 DVDD.n1262 2.24164
R24795 DVDD.n1605 DVDD.n1290 2.24164
R24796 DVDD.n1470 DVDD.n1262 2.24164
R24797 DVDD.n1605 DVDD.n1289 2.24164
R24798 DVDD.n1463 DVDD.n1262 2.24164
R24799 DVDD.n1605 DVDD.n1288 2.24164
R24800 DVDD.n1458 DVDD.n1262 2.24164
R24801 DVDD.n1605 DVDD.n1287 2.24164
R24802 DVDD.n1451 DVDD.n1262 2.24164
R24803 DVDD.n1605 DVDD.n1286 2.24164
R24804 DVDD.n1446 DVDD.n1262 2.24164
R24805 DVDD.n1605 DVDD.n1285 2.24164
R24806 DVDD.n1439 DVDD.n1262 2.24164
R24807 DVDD.n1605 DVDD.n1284 2.24164
R24808 DVDD.n1434 DVDD.n1262 2.24164
R24809 DVDD.n1605 DVDD.n1283 2.24164
R24810 DVDD.n1427 DVDD.n1262 2.24164
R24811 DVDD.n1605 DVDD.n1282 2.24164
R24812 DVDD.n1422 DVDD.n1262 2.24164
R24813 DVDD.n1605 DVDD.n1281 2.24164
R24814 DVDD.n1415 DVDD.n1262 2.24164
R24815 DVDD.n1605 DVDD.n1280 2.24164
R24816 DVDD.n1410 DVDD.n1262 2.24164
R24817 DVDD.n1605 DVDD.n1279 2.24164
R24818 DVDD.n1403 DVDD.n1262 2.24164
R24819 DVDD.n1605 DVDD.n1278 2.24164
R24820 DVDD.n1398 DVDD.n1262 2.24164
R24821 DVDD.n1605 DVDD.n1277 2.24164
R24822 DVDD.n1391 DVDD.n1262 2.24164
R24823 DVDD.n1605 DVDD.n1276 2.24164
R24824 DVDD.n1386 DVDD.n1262 2.24164
R24825 DVDD.n1605 DVDD.n1275 2.24164
R24826 DVDD.n1379 DVDD.n1262 2.24164
R24827 DVDD.n1605 DVDD.n1274 2.24164
R24828 DVDD.n1374 DVDD.n1262 2.24164
R24829 DVDD.n1605 DVDD.n1273 2.24164
R24830 DVDD.n1367 DVDD.n1262 2.24164
R24831 DVDD.n1605 DVDD.n1272 2.24164
R24832 DVDD.n1362 DVDD.n1262 2.24164
R24833 DVDD.n1605 DVDD.n1271 2.24164
R24834 DVDD.n1699 DVDD.n1658 2.24164
R24835 DVDD.n17262 DVDD.n1652 2.24164
R24836 DVDD.n17019 DVDD.n1658 2.24164
R24837 DVDD.n17262 DVDD.n1651 2.24164
R24838 DVDD.n17023 DVDD.n1658 2.24164
R24839 DVDD.n17262 DVDD.n1650 2.24164
R24840 DVDD.n17031 DVDD.n1658 2.24164
R24841 DVDD.n17262 DVDD.n1649 2.24164
R24842 DVDD.n17035 DVDD.n1658 2.24164
R24843 DVDD.n17262 DVDD.n1648 2.24164
R24844 DVDD.n17043 DVDD.n1658 2.24164
R24845 DVDD.n17262 DVDD.n1647 2.24164
R24846 DVDD.n17047 DVDD.n1658 2.24164
R24847 DVDD.n17262 DVDD.n1646 2.24164
R24848 DVDD.n17055 DVDD.n1658 2.24164
R24849 DVDD.n17262 DVDD.n1645 2.24164
R24850 DVDD.n17059 DVDD.n1658 2.24164
R24851 DVDD.n17262 DVDD.n1644 2.24164
R24852 DVDD.n17067 DVDD.n1658 2.24164
R24853 DVDD.n17262 DVDD.n1643 2.24164
R24854 DVDD.n17071 DVDD.n1658 2.24164
R24855 DVDD.n17262 DVDD.n1642 2.24164
R24856 DVDD.n17079 DVDD.n1658 2.24164
R24857 DVDD.n17262 DVDD.n1641 2.24164
R24858 DVDD.n17083 DVDD.n1658 2.24164
R24859 DVDD.n17262 DVDD.n1640 2.24164
R24860 DVDD.n17091 DVDD.n1658 2.24164
R24861 DVDD.n17262 DVDD.n1639 2.24164
R24862 DVDD.n17095 DVDD.n1658 2.24164
R24863 DVDD.n17262 DVDD.n1638 2.24164
R24864 DVDD.n17103 DVDD.n1658 2.24164
R24865 DVDD.n17262 DVDD.n1637 2.24164
R24866 DVDD.n17107 DVDD.n1658 2.24164
R24867 DVDD.n17262 DVDD.n1636 2.24164
R24868 DVDD.n17115 DVDD.n1658 2.24164
R24869 DVDD.n17262 DVDD.n1635 2.24164
R24870 DVDD.n17119 DVDD.n1658 2.24164
R24871 DVDD.n17262 DVDD.n1634 2.24164
R24872 DVDD.n17127 DVDD.n1658 2.24164
R24873 DVDD.n17262 DVDD.n1633 2.24164
R24874 DVDD.n17131 DVDD.n1658 2.24164
R24875 DVDD.n17262 DVDD.n1632 2.24164
R24876 DVDD.n17139 DVDD.n1658 2.24164
R24877 DVDD.n17262 DVDD.n1631 2.24164
R24878 DVDD.n17143 DVDD.n1658 2.24164
R24879 DVDD.n17262 DVDD.n1630 2.24164
R24880 DVDD.n17151 DVDD.n1658 2.24164
R24881 DVDD.n17262 DVDD.n1629 2.24164
R24882 DVDD.n17155 DVDD.n1658 2.24164
R24883 DVDD.n17262 DVDD.n1628 2.24164
R24884 DVDD.n17163 DVDD.n1658 2.24164
R24885 DVDD.n17262 DVDD.n1627 2.24164
R24886 DVDD.n17167 DVDD.n1658 2.24164
R24887 DVDD.n17262 DVDD.n1626 2.24164
R24888 DVDD.n17175 DVDD.n1658 2.24164
R24889 DVDD.n17262 DVDD.n1625 2.24164
R24890 DVDD.n17179 DVDD.n1658 2.24164
R24891 DVDD.n17262 DVDD.n1624 2.24164
R24892 DVDD.n17187 DVDD.n1658 2.24164
R24893 DVDD.n17262 DVDD.n1623 2.24164
R24894 DVDD.n17191 DVDD.n1658 2.24164
R24895 DVDD.n17262 DVDD.n1622 2.24164
R24896 DVDD.n17199 DVDD.n1658 2.24164
R24897 DVDD.n17262 DVDD.n1621 2.24164
R24898 DVDD.n17203 DVDD.n1658 2.24164
R24899 DVDD.n17262 DVDD.n1620 2.24164
R24900 DVDD.n17211 DVDD.n1658 2.24164
R24901 DVDD.n17262 DVDD.n1619 2.24164
R24902 DVDD.n17215 DVDD.n1658 2.24164
R24903 DVDD.n17262 DVDD.n1618 2.24164
R24904 DVDD.n17223 DVDD.n1658 2.24164
R24905 DVDD.n17262 DVDD.n1617 2.24164
R24906 DVDD.n17227 DVDD.n1658 2.24164
R24907 DVDD.n17262 DVDD.n1616 2.24164
R24908 DVDD.n17235 DVDD.n1658 2.24164
R24909 DVDD.n17262 DVDD.n1615 2.24164
R24910 DVDD.n17239 DVDD.n1658 2.24164
R24911 DVDD.n17262 DVDD.n1614 2.24164
R24912 DVDD.n17247 DVDD.n1658 2.24164
R24913 DVDD.n17262 DVDD.n1613 2.24164
R24914 DVDD.n17251 DVDD.n1658 2.24164
R24915 DVDD.n17262 DVDD.n1612 2.24164
R24916 DVDD.n17260 DVDD.n1658 2.24164
R24917 DVDD.n1798 DVDD.n1757 2.24164
R24918 DVDD.n16994 DVDD.n1753 2.24164
R24919 DVDD.n16751 DVDD.n1757 2.24164
R24920 DVDD.n16994 DVDD.n1752 2.24164
R24921 DVDD.n16755 DVDD.n1757 2.24164
R24922 DVDD.n16994 DVDD.n1751 2.24164
R24923 DVDD.n16763 DVDD.n1757 2.24164
R24924 DVDD.n16994 DVDD.n1750 2.24164
R24925 DVDD.n16767 DVDD.n1757 2.24164
R24926 DVDD.n16994 DVDD.n1749 2.24164
R24927 DVDD.n16775 DVDD.n1757 2.24164
R24928 DVDD.n16994 DVDD.n1748 2.24164
R24929 DVDD.n16779 DVDD.n1757 2.24164
R24930 DVDD.n16994 DVDD.n1747 2.24164
R24931 DVDD.n16787 DVDD.n1757 2.24164
R24932 DVDD.n16994 DVDD.n1746 2.24164
R24933 DVDD.n16791 DVDD.n1757 2.24164
R24934 DVDD.n16994 DVDD.n1745 2.24164
R24935 DVDD.n16799 DVDD.n1757 2.24164
R24936 DVDD.n16994 DVDD.n1744 2.24164
R24937 DVDD.n16803 DVDD.n1757 2.24164
R24938 DVDD.n16994 DVDD.n1743 2.24164
R24939 DVDD.n16811 DVDD.n1757 2.24164
R24940 DVDD.n16994 DVDD.n1742 2.24164
R24941 DVDD.n16815 DVDD.n1757 2.24164
R24942 DVDD.n16994 DVDD.n1741 2.24164
R24943 DVDD.n16823 DVDD.n1757 2.24164
R24944 DVDD.n16994 DVDD.n1740 2.24164
R24945 DVDD.n16827 DVDD.n1757 2.24164
R24946 DVDD.n16994 DVDD.n1739 2.24164
R24947 DVDD.n16835 DVDD.n1757 2.24164
R24948 DVDD.n16994 DVDD.n1738 2.24164
R24949 DVDD.n16839 DVDD.n1757 2.24164
R24950 DVDD.n16994 DVDD.n1737 2.24164
R24951 DVDD.n16847 DVDD.n1757 2.24164
R24952 DVDD.n16994 DVDD.n1736 2.24164
R24953 DVDD.n16851 DVDD.n1757 2.24164
R24954 DVDD.n16994 DVDD.n1735 2.24164
R24955 DVDD.n16859 DVDD.n1757 2.24164
R24956 DVDD.n16994 DVDD.n1734 2.24164
R24957 DVDD.n16863 DVDD.n1757 2.24164
R24958 DVDD.n16994 DVDD.n1733 2.24164
R24959 DVDD.n16871 DVDD.n1757 2.24164
R24960 DVDD.n16994 DVDD.n1732 2.24164
R24961 DVDD.n16875 DVDD.n1757 2.24164
R24962 DVDD.n16994 DVDD.n1731 2.24164
R24963 DVDD.n16883 DVDD.n1757 2.24164
R24964 DVDD.n16994 DVDD.n1730 2.24164
R24965 DVDD.n16887 DVDD.n1757 2.24164
R24966 DVDD.n16994 DVDD.n1729 2.24164
R24967 DVDD.n16895 DVDD.n1757 2.24164
R24968 DVDD.n16994 DVDD.n1728 2.24164
R24969 DVDD.n16899 DVDD.n1757 2.24164
R24970 DVDD.n16994 DVDD.n1727 2.24164
R24971 DVDD.n16907 DVDD.n1757 2.24164
R24972 DVDD.n16994 DVDD.n1726 2.24164
R24973 DVDD.n16911 DVDD.n1757 2.24164
R24974 DVDD.n16994 DVDD.n1725 2.24164
R24975 DVDD.n16919 DVDD.n1757 2.24164
R24976 DVDD.n16994 DVDD.n1724 2.24164
R24977 DVDD.n16923 DVDD.n1757 2.24164
R24978 DVDD.n16994 DVDD.n1723 2.24164
R24979 DVDD.n16931 DVDD.n1757 2.24164
R24980 DVDD.n16994 DVDD.n1722 2.24164
R24981 DVDD.n16935 DVDD.n1757 2.24164
R24982 DVDD.n16994 DVDD.n1721 2.24164
R24983 DVDD.n16943 DVDD.n1757 2.24164
R24984 DVDD.n16994 DVDD.n1720 2.24164
R24985 DVDD.n16947 DVDD.n1757 2.24164
R24986 DVDD.n16994 DVDD.n1719 2.24164
R24987 DVDD.n16955 DVDD.n1757 2.24164
R24988 DVDD.n16994 DVDD.n1718 2.24164
R24989 DVDD.n16959 DVDD.n1757 2.24164
R24990 DVDD.n16994 DVDD.n1717 2.24164
R24991 DVDD.n16967 DVDD.n1757 2.24164
R24992 DVDD.n16994 DVDD.n1716 2.24164
R24993 DVDD.n16971 DVDD.n1757 2.24164
R24994 DVDD.n16994 DVDD.n1715 2.24164
R24995 DVDD.n16979 DVDD.n1757 2.24164
R24996 DVDD.n16994 DVDD.n1714 2.24164
R24997 DVDD.n16983 DVDD.n1757 2.24164
R24998 DVDD.n16994 DVDD.n1713 2.24164
R24999 DVDD.n16992 DVDD.n1757 2.24164
R25000 DVDD.n2156 DVDD.n2155 2.24164
R25001 DVDD.n1864 DVDD.n1813 2.24164
R25002 DVDD.n2156 DVDD.n1862 2.24164
R25003 DVDD.n2146 DVDD.n1813 2.24164
R25004 DVDD.n2156 DVDD.n1861 2.24164
R25005 DVDD.n2141 DVDD.n1813 2.24164
R25006 DVDD.n2156 DVDD.n1860 2.24164
R25007 DVDD.n2134 DVDD.n1813 2.24164
R25008 DVDD.n2156 DVDD.n1859 2.24164
R25009 DVDD.n2129 DVDD.n1813 2.24164
R25010 DVDD.n2156 DVDD.n1858 2.24164
R25011 DVDD.n2122 DVDD.n1813 2.24164
R25012 DVDD.n2156 DVDD.n1857 2.24164
R25013 DVDD.n2117 DVDD.n1813 2.24164
R25014 DVDD.n2156 DVDD.n1856 2.24164
R25015 DVDD.n2110 DVDD.n1813 2.24164
R25016 DVDD.n2156 DVDD.n1855 2.24164
R25017 DVDD.n2105 DVDD.n1813 2.24164
R25018 DVDD.n2156 DVDD.n1854 2.24164
R25019 DVDD.n2098 DVDD.n1813 2.24164
R25020 DVDD.n2156 DVDD.n1853 2.24164
R25021 DVDD.n2093 DVDD.n1813 2.24164
R25022 DVDD.n2156 DVDD.n1852 2.24164
R25023 DVDD.n2086 DVDD.n1813 2.24164
R25024 DVDD.n2156 DVDD.n1851 2.24164
R25025 DVDD.n2081 DVDD.n1813 2.24164
R25026 DVDD.n2156 DVDD.n1850 2.24164
R25027 DVDD.n2074 DVDD.n1813 2.24164
R25028 DVDD.n2156 DVDD.n1849 2.24164
R25029 DVDD.n2069 DVDD.n1813 2.24164
R25030 DVDD.n2156 DVDD.n1848 2.24164
R25031 DVDD.n2062 DVDD.n1813 2.24164
R25032 DVDD.n2156 DVDD.n1847 2.24164
R25033 DVDD.n2057 DVDD.n1813 2.24164
R25034 DVDD.n2156 DVDD.n1846 2.24164
R25035 DVDD.n2050 DVDD.n1813 2.24164
R25036 DVDD.n2156 DVDD.n1845 2.24164
R25037 DVDD.n2045 DVDD.n1813 2.24164
R25038 DVDD.n2156 DVDD.n1844 2.24164
R25039 DVDD.n2038 DVDD.n1813 2.24164
R25040 DVDD.n2156 DVDD.n1843 2.24164
R25041 DVDD.n2033 DVDD.n1813 2.24164
R25042 DVDD.n2156 DVDD.n1842 2.24164
R25043 DVDD.n2026 DVDD.n1813 2.24164
R25044 DVDD.n2156 DVDD.n1841 2.24164
R25045 DVDD.n2021 DVDD.n1813 2.24164
R25046 DVDD.n2156 DVDD.n1840 2.24164
R25047 DVDD.n2014 DVDD.n1813 2.24164
R25048 DVDD.n2156 DVDD.n1839 2.24164
R25049 DVDD.n2009 DVDD.n1813 2.24164
R25050 DVDD.n2156 DVDD.n1838 2.24164
R25051 DVDD.n2002 DVDD.n1813 2.24164
R25052 DVDD.n2156 DVDD.n1837 2.24164
R25053 DVDD.n1997 DVDD.n1813 2.24164
R25054 DVDD.n2156 DVDD.n1836 2.24164
R25055 DVDD.n1990 DVDD.n1813 2.24164
R25056 DVDD.n2156 DVDD.n1835 2.24164
R25057 DVDD.n1985 DVDD.n1813 2.24164
R25058 DVDD.n2156 DVDD.n1834 2.24164
R25059 DVDD.n1978 DVDD.n1813 2.24164
R25060 DVDD.n2156 DVDD.n1833 2.24164
R25061 DVDD.n1973 DVDD.n1813 2.24164
R25062 DVDD.n2156 DVDD.n1832 2.24164
R25063 DVDD.n1966 DVDD.n1813 2.24164
R25064 DVDD.n2156 DVDD.n1831 2.24164
R25065 DVDD.n1961 DVDD.n1813 2.24164
R25066 DVDD.n2156 DVDD.n1830 2.24164
R25067 DVDD.n1954 DVDD.n1813 2.24164
R25068 DVDD.n2156 DVDD.n1829 2.24164
R25069 DVDD.n1949 DVDD.n1813 2.24164
R25070 DVDD.n2156 DVDD.n1828 2.24164
R25071 DVDD.n1942 DVDD.n1813 2.24164
R25072 DVDD.n2156 DVDD.n1827 2.24164
R25073 DVDD.n1937 DVDD.n1813 2.24164
R25074 DVDD.n2156 DVDD.n1826 2.24164
R25075 DVDD.n1930 DVDD.n1813 2.24164
R25076 DVDD.n2156 DVDD.n1825 2.24164
R25077 DVDD.n1925 DVDD.n1813 2.24164
R25078 DVDD.n2156 DVDD.n1824 2.24164
R25079 DVDD.n1918 DVDD.n1813 2.24164
R25080 DVDD.n2156 DVDD.n1823 2.24164
R25081 DVDD.n1913 DVDD.n1813 2.24164
R25082 DVDD.n2156 DVDD.n1822 2.24164
R25083 DVDD.n2251 DVDD.n2210 2.24164
R25084 DVDD.n16704 DVDD.n2206 2.24164
R25085 DVDD.n16462 DVDD.n2210 2.24164
R25086 DVDD.n16704 DVDD.n2205 2.24164
R25087 DVDD.n16466 DVDD.n2210 2.24164
R25088 DVDD.n16704 DVDD.n2204 2.24164
R25089 DVDD.n16474 DVDD.n2210 2.24164
R25090 DVDD.n16704 DVDD.n2203 2.24164
R25091 DVDD.n16478 DVDD.n2210 2.24164
R25092 DVDD.n16704 DVDD.n2202 2.24164
R25093 DVDD.n16486 DVDD.n2210 2.24164
R25094 DVDD.n16704 DVDD.n2201 2.24164
R25095 DVDD.n16490 DVDD.n2210 2.24164
R25096 DVDD.n16704 DVDD.n2200 2.24164
R25097 DVDD.n16498 DVDD.n2210 2.24164
R25098 DVDD.n16704 DVDD.n2199 2.24164
R25099 DVDD.n16502 DVDD.n2210 2.24164
R25100 DVDD.n16704 DVDD.n2198 2.24164
R25101 DVDD.n16510 DVDD.n2210 2.24164
R25102 DVDD.n16704 DVDD.n2197 2.24164
R25103 DVDD.n16514 DVDD.n2210 2.24164
R25104 DVDD.n16704 DVDD.n2196 2.24164
R25105 DVDD.n16522 DVDD.n2210 2.24164
R25106 DVDD.n16704 DVDD.n2195 2.24164
R25107 DVDD.n16526 DVDD.n2210 2.24164
R25108 DVDD.n16704 DVDD.n2194 2.24164
R25109 DVDD.n16534 DVDD.n2210 2.24164
R25110 DVDD.n16704 DVDD.n2193 2.24164
R25111 DVDD.n16538 DVDD.n2210 2.24164
R25112 DVDD.n16704 DVDD.n2192 2.24164
R25113 DVDD.n16546 DVDD.n2210 2.24164
R25114 DVDD.n16704 DVDD.n2191 2.24164
R25115 DVDD.n16550 DVDD.n2210 2.24164
R25116 DVDD.n16704 DVDD.n2190 2.24164
R25117 DVDD.n16558 DVDD.n2210 2.24164
R25118 DVDD.n16704 DVDD.n2189 2.24164
R25119 DVDD.n16562 DVDD.n2210 2.24164
R25120 DVDD.n16704 DVDD.n2188 2.24164
R25121 DVDD.n16570 DVDD.n2210 2.24164
R25122 DVDD.n16704 DVDD.n2187 2.24164
R25123 DVDD.n16574 DVDD.n2210 2.24164
R25124 DVDD.n16704 DVDD.n2186 2.24164
R25125 DVDD.n16582 DVDD.n2210 2.24164
R25126 DVDD.n16704 DVDD.n2185 2.24164
R25127 DVDD.n16586 DVDD.n2210 2.24164
R25128 DVDD.n16704 DVDD.n2184 2.24164
R25129 DVDD.n16594 DVDD.n2210 2.24164
R25130 DVDD.n16704 DVDD.n2183 2.24164
R25131 DVDD.n16598 DVDD.n2210 2.24164
R25132 DVDD.n16704 DVDD.n2182 2.24164
R25133 DVDD.n16606 DVDD.n2210 2.24164
R25134 DVDD.n16704 DVDD.n2181 2.24164
R25135 DVDD.n16610 DVDD.n2210 2.24164
R25136 DVDD.n16704 DVDD.n2180 2.24164
R25137 DVDD.n16618 DVDD.n2210 2.24164
R25138 DVDD.n16704 DVDD.n2179 2.24164
R25139 DVDD.n16622 DVDD.n2210 2.24164
R25140 DVDD.n16704 DVDD.n2178 2.24164
R25141 DVDD.n16630 DVDD.n2210 2.24164
R25142 DVDD.n16704 DVDD.n2177 2.24164
R25143 DVDD.n16634 DVDD.n2210 2.24164
R25144 DVDD.n16704 DVDD.n2176 2.24164
R25145 DVDD.n16642 DVDD.n2210 2.24164
R25146 DVDD.n16704 DVDD.n2175 2.24164
R25147 DVDD.n16646 DVDD.n2210 2.24164
R25148 DVDD.n16704 DVDD.n2174 2.24164
R25149 DVDD.n16654 DVDD.n2210 2.24164
R25150 DVDD.n16704 DVDD.n2173 2.24164
R25151 DVDD.n16658 DVDD.n2210 2.24164
R25152 DVDD.n16704 DVDD.n2172 2.24164
R25153 DVDD.n16666 DVDD.n2210 2.24164
R25154 DVDD.n16704 DVDD.n2171 2.24164
R25155 DVDD.n16670 DVDD.n2210 2.24164
R25156 DVDD.n16704 DVDD.n2170 2.24164
R25157 DVDD.n16678 DVDD.n2210 2.24164
R25158 DVDD.n16704 DVDD.n2169 2.24164
R25159 DVDD.n16682 DVDD.n2210 2.24164
R25160 DVDD.n16704 DVDD.n2168 2.24164
R25161 DVDD.n16690 DVDD.n2210 2.24164
R25162 DVDD.n16704 DVDD.n2167 2.24164
R25163 DVDD.n16694 DVDD.n2210 2.24164
R25164 DVDD.n16704 DVDD.n2166 2.24164
R25165 DVDD.n16702 DVDD.n2210 2.24164
R25166 DVDD.n13256 DVDD.n13255 2.24164
R25167 DVDD.n12965 DVDD.n12912 2.24164
R25168 DVDD.n13256 DVDD.n12963 2.24164
R25169 DVDD.n13246 DVDD.n12912 2.24164
R25170 DVDD.n13256 DVDD.n12962 2.24164
R25171 DVDD.n13241 DVDD.n12912 2.24164
R25172 DVDD.n13256 DVDD.n12961 2.24164
R25173 DVDD.n13234 DVDD.n12912 2.24164
R25174 DVDD.n13256 DVDD.n12960 2.24164
R25175 DVDD.n13229 DVDD.n12912 2.24164
R25176 DVDD.n13256 DVDD.n12959 2.24164
R25177 DVDD.n13222 DVDD.n12912 2.24164
R25178 DVDD.n13256 DVDD.n12958 2.24164
R25179 DVDD.n13217 DVDD.n12912 2.24164
R25180 DVDD.n13256 DVDD.n12957 2.24164
R25181 DVDD.n13210 DVDD.n12912 2.24164
R25182 DVDD.n13256 DVDD.n12956 2.24164
R25183 DVDD.n13205 DVDD.n12912 2.24164
R25184 DVDD.n13256 DVDD.n12955 2.24164
R25185 DVDD.n13198 DVDD.n12912 2.24164
R25186 DVDD.n13256 DVDD.n12954 2.24164
R25187 DVDD.n13193 DVDD.n12912 2.24164
R25188 DVDD.n13256 DVDD.n12953 2.24164
R25189 DVDD.n13186 DVDD.n12912 2.24164
R25190 DVDD.n13256 DVDD.n12952 2.24164
R25191 DVDD.n13181 DVDD.n12912 2.24164
R25192 DVDD.n13256 DVDD.n12951 2.24164
R25193 DVDD.n13174 DVDD.n12912 2.24164
R25194 DVDD.n13256 DVDD.n12950 2.24164
R25195 DVDD.n13169 DVDD.n12912 2.24164
R25196 DVDD.n13256 DVDD.n12949 2.24164
R25197 DVDD.n13162 DVDD.n12912 2.24164
R25198 DVDD.n13256 DVDD.n12948 2.24164
R25199 DVDD.n13157 DVDD.n12912 2.24164
R25200 DVDD.n13256 DVDD.n12947 2.24164
R25201 DVDD.n13150 DVDD.n12912 2.24164
R25202 DVDD.n13256 DVDD.n12946 2.24164
R25203 DVDD.n13145 DVDD.n12912 2.24164
R25204 DVDD.n13256 DVDD.n12945 2.24164
R25205 DVDD.n13138 DVDD.n12912 2.24164
R25206 DVDD.n13256 DVDD.n12944 2.24164
R25207 DVDD.n13133 DVDD.n12912 2.24164
R25208 DVDD.n13256 DVDD.n12943 2.24164
R25209 DVDD.n13126 DVDD.n12912 2.24164
R25210 DVDD.n13256 DVDD.n12942 2.24164
R25211 DVDD.n13121 DVDD.n12912 2.24164
R25212 DVDD.n13256 DVDD.n12941 2.24164
R25213 DVDD.n13114 DVDD.n12912 2.24164
R25214 DVDD.n13256 DVDD.n12940 2.24164
R25215 DVDD.n13109 DVDD.n12912 2.24164
R25216 DVDD.n13256 DVDD.n12939 2.24164
R25217 DVDD.n13102 DVDD.n12912 2.24164
R25218 DVDD.n13256 DVDD.n12938 2.24164
R25219 DVDD.n13097 DVDD.n12912 2.24164
R25220 DVDD.n13256 DVDD.n12937 2.24164
R25221 DVDD.n13090 DVDD.n12912 2.24164
R25222 DVDD.n13256 DVDD.n12936 2.24164
R25223 DVDD.n13085 DVDD.n12912 2.24164
R25224 DVDD.n13256 DVDD.n12935 2.24164
R25225 DVDD.n13078 DVDD.n12912 2.24164
R25226 DVDD.n13256 DVDD.n12934 2.24164
R25227 DVDD.n13073 DVDD.n12912 2.24164
R25228 DVDD.n13256 DVDD.n12933 2.24164
R25229 DVDD.n13066 DVDD.n12912 2.24164
R25230 DVDD.n13256 DVDD.n12932 2.24164
R25231 DVDD.n13061 DVDD.n12912 2.24164
R25232 DVDD.n13256 DVDD.n12931 2.24164
R25233 DVDD.n13054 DVDD.n12912 2.24164
R25234 DVDD.n13256 DVDD.n12930 2.24164
R25235 DVDD.n13049 DVDD.n12912 2.24164
R25236 DVDD.n13256 DVDD.n12929 2.24164
R25237 DVDD.n13042 DVDD.n12912 2.24164
R25238 DVDD.n13256 DVDD.n12928 2.24164
R25239 DVDD.n13037 DVDD.n12912 2.24164
R25240 DVDD.n13256 DVDD.n12927 2.24164
R25241 DVDD.n13030 DVDD.n12912 2.24164
R25242 DVDD.n13256 DVDD.n12926 2.24164
R25243 DVDD.n13025 DVDD.n12912 2.24164
R25244 DVDD.n13256 DVDD.n12925 2.24164
R25245 DVDD.n13018 DVDD.n12912 2.24164
R25246 DVDD.n13256 DVDD.n12924 2.24164
R25247 DVDD.n13013 DVDD.n12912 2.24164
R25248 DVDD.n13256 DVDD.n12923 2.24164
R25249 DVDD.n13473 DVDD.n13472 2.24164
R25250 DVDD.n13470 DVDD.n12824 2.24164
R25251 DVDD.n13473 DVDD.n12778 2.24164
R25252 DVDD.n13470 DVDD.n12823 2.24164
R25253 DVDD.n13473 DVDD.n12777 2.24164
R25254 DVDD.n13470 DVDD.n12822 2.24164
R25255 DVDD.n13473 DVDD.n12776 2.24164
R25256 DVDD.n13470 DVDD.n12821 2.24164
R25257 DVDD.n13473 DVDD.n12775 2.24164
R25258 DVDD.n13470 DVDD.n12820 2.24164
R25259 DVDD.n13473 DVDD.n12774 2.24164
R25260 DVDD.n13470 DVDD.n12819 2.24164
R25261 DVDD.n13473 DVDD.n12773 2.24164
R25262 DVDD.n13470 DVDD.n12818 2.24164
R25263 DVDD.n13473 DVDD.n12772 2.24164
R25264 DVDD.n13470 DVDD.n12817 2.24164
R25265 DVDD.n13473 DVDD.n12771 2.24164
R25266 DVDD.n13470 DVDD.n12816 2.24164
R25267 DVDD.n13473 DVDD.n12770 2.24164
R25268 DVDD.n13470 DVDD.n12815 2.24164
R25269 DVDD.n13473 DVDD.n12769 2.24164
R25270 DVDD.n13470 DVDD.n12814 2.24164
R25271 DVDD.n13473 DVDD.n12768 2.24164
R25272 DVDD.n13470 DVDD.n12813 2.24164
R25273 DVDD.n13473 DVDD.n12767 2.24164
R25274 DVDD.n13470 DVDD.n12812 2.24164
R25275 DVDD.n13473 DVDD.n12766 2.24164
R25276 DVDD.n13470 DVDD.n12811 2.24164
R25277 DVDD.n13473 DVDD.n12765 2.24164
R25278 DVDD.n13470 DVDD.n12810 2.24164
R25279 DVDD.n13473 DVDD.n12764 2.24164
R25280 DVDD.n13470 DVDD.n12809 2.24164
R25281 DVDD.n13473 DVDD.n12763 2.24164
R25282 DVDD.n13470 DVDD.n12808 2.24164
R25283 DVDD.n13473 DVDD.n12762 2.24164
R25284 DVDD.n13470 DVDD.n12807 2.24164
R25285 DVDD.n13473 DVDD.n12761 2.24164
R25286 DVDD.n13470 DVDD.n12806 2.24164
R25287 DVDD.n13473 DVDD.n12760 2.24164
R25288 DVDD.n13470 DVDD.n12805 2.24164
R25289 DVDD.n13473 DVDD.n12759 2.24164
R25290 DVDD.n13470 DVDD.n12804 2.24164
R25291 DVDD.n13473 DVDD.n12758 2.24164
R25292 DVDD.n13470 DVDD.n12803 2.24164
R25293 DVDD.n13473 DVDD.n12757 2.24164
R25294 DVDD.n13470 DVDD.n12802 2.24164
R25295 DVDD.n13473 DVDD.n12756 2.24164
R25296 DVDD.n13470 DVDD.n12801 2.24164
R25297 DVDD.n13473 DVDD.n12755 2.24164
R25298 DVDD.n13470 DVDD.n12800 2.24164
R25299 DVDD.n13473 DVDD.n12754 2.24164
R25300 DVDD.n13470 DVDD.n12799 2.24164
R25301 DVDD.n13473 DVDD.n12753 2.24164
R25302 DVDD.n13470 DVDD.n12798 2.24164
R25303 DVDD.n13473 DVDD.n12752 2.24164
R25304 DVDD.n13470 DVDD.n12797 2.24164
R25305 DVDD.n13473 DVDD.n12751 2.24164
R25306 DVDD.n13470 DVDD.n12796 2.24164
R25307 DVDD.n13473 DVDD.n12750 2.24164
R25308 DVDD.n13470 DVDD.n12795 2.24164
R25309 DVDD.n13473 DVDD.n12749 2.24164
R25310 DVDD.n13470 DVDD.n12794 2.24164
R25311 DVDD.n13473 DVDD.n12748 2.24164
R25312 DVDD.n13470 DVDD.n12793 2.24164
R25313 DVDD.n13473 DVDD.n12747 2.24164
R25314 DVDD.n13470 DVDD.n12792 2.24164
R25315 DVDD.n13473 DVDD.n12746 2.24164
R25316 DVDD.n13470 DVDD.n12791 2.24164
R25317 DVDD.n13473 DVDD.n12745 2.24164
R25318 DVDD.n13470 DVDD.n12790 2.24164
R25319 DVDD.n13473 DVDD.n12744 2.24164
R25320 DVDD.n13470 DVDD.n12789 2.24164
R25321 DVDD.n13473 DVDD.n12743 2.24164
R25322 DVDD.n13470 DVDD.n12788 2.24164
R25323 DVDD.n13473 DVDD.n12742 2.24164
R25324 DVDD.n13470 DVDD.n12787 2.24164
R25325 DVDD.n13473 DVDD.n12741 2.24164
R25326 DVDD.n13470 DVDD.n12786 2.24164
R25327 DVDD.n13473 DVDD.n12740 2.24164
R25328 DVDD.n13470 DVDD.n12785 2.24164
R25329 DVDD.n13473 DVDD.n12739 2.24164
R25330 DVDD.n13470 DVDD.n12784 2.24164
R25331 DVDD.n13473 DVDD.n12738 2.24164
R25332 DVDD.n13487 DVDD.n13486 2.24164
R25333 DVDD.n13484 DVDD.n12476 2.24164
R25334 DVDD.n13487 DVDD.n12431 2.24164
R25335 DVDD.n13484 DVDD.n12475 2.24164
R25336 DVDD.n13487 DVDD.n12430 2.24164
R25337 DVDD.n13484 DVDD.n12474 2.24164
R25338 DVDD.n13487 DVDD.n12429 2.24164
R25339 DVDD.n13484 DVDD.n12473 2.24164
R25340 DVDD.n13487 DVDD.n12428 2.24164
R25341 DVDD.n13484 DVDD.n12472 2.24164
R25342 DVDD.n13487 DVDD.n12427 2.24164
R25343 DVDD.n13484 DVDD.n12471 2.24164
R25344 DVDD.n13487 DVDD.n12426 2.24164
R25345 DVDD.n13484 DVDD.n12470 2.24164
R25346 DVDD.n13487 DVDD.n12425 2.24164
R25347 DVDD.n13484 DVDD.n12469 2.24164
R25348 DVDD.n13487 DVDD.n12424 2.24164
R25349 DVDD.n13484 DVDD.n12468 2.24164
R25350 DVDD.n13487 DVDD.n12423 2.24164
R25351 DVDD.n13484 DVDD.n12467 2.24164
R25352 DVDD.n13487 DVDD.n12422 2.24164
R25353 DVDD.n13484 DVDD.n12466 2.24164
R25354 DVDD.n13487 DVDD.n12421 2.24164
R25355 DVDD.n13484 DVDD.n12465 2.24164
R25356 DVDD.n13487 DVDD.n12420 2.24164
R25357 DVDD.n13484 DVDD.n12464 2.24164
R25358 DVDD.n13487 DVDD.n12419 2.24164
R25359 DVDD.n13484 DVDD.n12463 2.24164
R25360 DVDD.n13487 DVDD.n12418 2.24164
R25361 DVDD.n13484 DVDD.n12462 2.24164
R25362 DVDD.n13487 DVDD.n12417 2.24164
R25363 DVDD.n13484 DVDD.n12461 2.24164
R25364 DVDD.n13487 DVDD.n12416 2.24164
R25365 DVDD.n13484 DVDD.n12460 2.24164
R25366 DVDD.n13487 DVDD.n12415 2.24164
R25367 DVDD.n13484 DVDD.n12459 2.24164
R25368 DVDD.n13487 DVDD.n12414 2.24164
R25369 DVDD.n13484 DVDD.n12458 2.24164
R25370 DVDD.n13487 DVDD.n12413 2.24164
R25371 DVDD.n13484 DVDD.n12457 2.24164
R25372 DVDD.n13487 DVDD.n12412 2.24164
R25373 DVDD.n13484 DVDD.n12456 2.24164
R25374 DVDD.n13487 DVDD.n12411 2.24164
R25375 DVDD.n13484 DVDD.n12455 2.24164
R25376 DVDD.n13487 DVDD.n12410 2.24164
R25377 DVDD.n13484 DVDD.n12454 2.24164
R25378 DVDD.n13487 DVDD.n12409 2.24164
R25379 DVDD.n13484 DVDD.n12453 2.24164
R25380 DVDD.n13487 DVDD.n12408 2.24164
R25381 DVDD.n13484 DVDD.n12452 2.24164
R25382 DVDD.n13487 DVDD.n12407 2.24164
R25383 DVDD.n13484 DVDD.n12451 2.24164
R25384 DVDD.n13487 DVDD.n12406 2.24164
R25385 DVDD.n13484 DVDD.n12450 2.24164
R25386 DVDD.n13487 DVDD.n12405 2.24164
R25387 DVDD.n13484 DVDD.n12449 2.24164
R25388 DVDD.n13487 DVDD.n12404 2.24164
R25389 DVDD.n13484 DVDD.n12448 2.24164
R25390 DVDD.n13487 DVDD.n12403 2.24164
R25391 DVDD.n13484 DVDD.n12447 2.24164
R25392 DVDD.n13487 DVDD.n12402 2.24164
R25393 DVDD.n13484 DVDD.n12446 2.24164
R25394 DVDD.n13487 DVDD.n12401 2.24164
R25395 DVDD.n13484 DVDD.n12445 2.24164
R25396 DVDD.n13487 DVDD.n12400 2.24164
R25397 DVDD.n13484 DVDD.n12444 2.24164
R25398 DVDD.n13487 DVDD.n12399 2.24164
R25399 DVDD.n13484 DVDD.n12443 2.24164
R25400 DVDD.n13487 DVDD.n12398 2.24164
R25401 DVDD.n13484 DVDD.n12442 2.24164
R25402 DVDD.n13487 DVDD.n12397 2.24164
R25403 DVDD.n13484 DVDD.n12441 2.24164
R25404 DVDD.n13487 DVDD.n12396 2.24164
R25405 DVDD.n13484 DVDD.n12440 2.24164
R25406 DVDD.n13487 DVDD.n12395 2.24164
R25407 DVDD.n13484 DVDD.n12439 2.24164
R25408 DVDD.n13487 DVDD.n12394 2.24164
R25409 DVDD.n13484 DVDD.n12438 2.24164
R25410 DVDD.n13487 DVDD.n12393 2.24164
R25411 DVDD.n13484 DVDD.n12437 2.24164
R25412 DVDD.n13487 DVDD.n12392 2.24164
R25413 DVDD.n13484 DVDD.n12436 2.24164
R25414 DVDD.n13487 DVDD.n12391 2.24164
R25415 DVDD.n12374 DVDD.n12333 2.24164
R25416 DVDD.n13744 DVDD.n12328 2.24164
R25417 DVDD.n13502 DVDD.n12333 2.24164
R25418 DVDD.n13744 DVDD.n12327 2.24164
R25419 DVDD.n13506 DVDD.n12333 2.24164
R25420 DVDD.n13744 DVDD.n12326 2.24164
R25421 DVDD.n13514 DVDD.n12333 2.24164
R25422 DVDD.n13744 DVDD.n12325 2.24164
R25423 DVDD.n13518 DVDD.n12333 2.24164
R25424 DVDD.n13744 DVDD.n12324 2.24164
R25425 DVDD.n13526 DVDD.n12333 2.24164
R25426 DVDD.n13744 DVDD.n12323 2.24164
R25427 DVDD.n13530 DVDD.n12333 2.24164
R25428 DVDD.n13744 DVDD.n12322 2.24164
R25429 DVDD.n13538 DVDD.n12333 2.24164
R25430 DVDD.n13744 DVDD.n12321 2.24164
R25431 DVDD.n13542 DVDD.n12333 2.24164
R25432 DVDD.n13744 DVDD.n12320 2.24164
R25433 DVDD.n13550 DVDD.n12333 2.24164
R25434 DVDD.n13744 DVDD.n12319 2.24164
R25435 DVDD.n13554 DVDD.n12333 2.24164
R25436 DVDD.n13744 DVDD.n12318 2.24164
R25437 DVDD.n13562 DVDD.n12333 2.24164
R25438 DVDD.n13744 DVDD.n12317 2.24164
R25439 DVDD.n13566 DVDD.n12333 2.24164
R25440 DVDD.n13744 DVDD.n12316 2.24164
R25441 DVDD.n13574 DVDD.n12333 2.24164
R25442 DVDD.n13744 DVDD.n12315 2.24164
R25443 DVDD.n13578 DVDD.n12333 2.24164
R25444 DVDD.n13744 DVDD.n12314 2.24164
R25445 DVDD.n13586 DVDD.n12333 2.24164
R25446 DVDD.n13744 DVDD.n12313 2.24164
R25447 DVDD.n13590 DVDD.n12333 2.24164
R25448 DVDD.n13744 DVDD.n12312 2.24164
R25449 DVDD.n13598 DVDD.n12333 2.24164
R25450 DVDD.n13744 DVDD.n12311 2.24164
R25451 DVDD.n13602 DVDD.n12333 2.24164
R25452 DVDD.n13744 DVDD.n12310 2.24164
R25453 DVDD.n13610 DVDD.n12333 2.24164
R25454 DVDD.n13744 DVDD.n12309 2.24164
R25455 DVDD.n13614 DVDD.n12333 2.24164
R25456 DVDD.n13744 DVDD.n12308 2.24164
R25457 DVDD.n13622 DVDD.n12333 2.24164
R25458 DVDD.n13744 DVDD.n12307 2.24164
R25459 DVDD.n13626 DVDD.n12333 2.24164
R25460 DVDD.n13744 DVDD.n12306 2.24164
R25461 DVDD.n13634 DVDD.n12333 2.24164
R25462 DVDD.n13744 DVDD.n12305 2.24164
R25463 DVDD.n13638 DVDD.n12333 2.24164
R25464 DVDD.n13744 DVDD.n12304 2.24164
R25465 DVDD.n13646 DVDD.n12333 2.24164
R25466 DVDD.n13744 DVDD.n12303 2.24164
R25467 DVDD.n13650 DVDD.n12333 2.24164
R25468 DVDD.n13744 DVDD.n12302 2.24164
R25469 DVDD.n13658 DVDD.n12333 2.24164
R25470 DVDD.n13744 DVDD.n12301 2.24164
R25471 DVDD.n13662 DVDD.n12333 2.24164
R25472 DVDD.n13744 DVDD.n12300 2.24164
R25473 DVDD.n13670 DVDD.n12333 2.24164
R25474 DVDD.n13744 DVDD.n12299 2.24164
R25475 DVDD.n13674 DVDD.n12333 2.24164
R25476 DVDD.n13744 DVDD.n12298 2.24164
R25477 DVDD.n13682 DVDD.n12333 2.24164
R25478 DVDD.n13744 DVDD.n12297 2.24164
R25479 DVDD.n13686 DVDD.n12333 2.24164
R25480 DVDD.n13744 DVDD.n12296 2.24164
R25481 DVDD.n13694 DVDD.n12333 2.24164
R25482 DVDD.n13744 DVDD.n12295 2.24164
R25483 DVDD.n13698 DVDD.n12333 2.24164
R25484 DVDD.n13744 DVDD.n12294 2.24164
R25485 DVDD.n13706 DVDD.n12333 2.24164
R25486 DVDD.n13744 DVDD.n12293 2.24164
R25487 DVDD.n13710 DVDD.n12333 2.24164
R25488 DVDD.n13744 DVDD.n12292 2.24164
R25489 DVDD.n13718 DVDD.n12333 2.24164
R25490 DVDD.n13744 DVDD.n12291 2.24164
R25491 DVDD.n13722 DVDD.n12333 2.24164
R25492 DVDD.n13744 DVDD.n12290 2.24164
R25493 DVDD.n13730 DVDD.n12333 2.24164
R25494 DVDD.n13744 DVDD.n12289 2.24164
R25495 DVDD.n13734 DVDD.n12333 2.24164
R25496 DVDD.n13744 DVDD.n12288 2.24164
R25497 DVDD.n13742 DVDD.n12333 2.24164
R25498 DVDD.n12029 DVDD.n11926 2.24164
R25499 DVDD.n12031 DVDD.n11938 2.24164
R25500 DVDD.n12033 DVDD.n11926 2.24164
R25501 DVDD.n12023 DVDD.n11938 2.24164
R25502 DVDD.n12041 DVDD.n11926 2.24164
R25503 DVDD.n12043 DVDD.n11938 2.24164
R25504 DVDD.n12045 DVDD.n11926 2.24164
R25505 DVDD.n12019 DVDD.n11938 2.24164
R25506 DVDD.n12053 DVDD.n11926 2.24164
R25507 DVDD.n12055 DVDD.n11938 2.24164
R25508 DVDD.n12057 DVDD.n11926 2.24164
R25509 DVDD.n12015 DVDD.n11938 2.24164
R25510 DVDD.n12065 DVDD.n11926 2.24164
R25511 DVDD.n12067 DVDD.n11938 2.24164
R25512 DVDD.n12069 DVDD.n11926 2.24164
R25513 DVDD.n12011 DVDD.n11938 2.24164
R25514 DVDD.n12077 DVDD.n11926 2.24164
R25515 DVDD.n12079 DVDD.n11938 2.24164
R25516 DVDD.n12081 DVDD.n11926 2.24164
R25517 DVDD.n12007 DVDD.n11938 2.24164
R25518 DVDD.n12089 DVDD.n11926 2.24164
R25519 DVDD.n12091 DVDD.n11938 2.24164
R25520 DVDD.n12093 DVDD.n11926 2.24164
R25521 DVDD.n12003 DVDD.n11938 2.24164
R25522 DVDD.n12101 DVDD.n11926 2.24164
R25523 DVDD.n12103 DVDD.n11938 2.24164
R25524 DVDD.n12105 DVDD.n11926 2.24164
R25525 DVDD.n11999 DVDD.n11938 2.24164
R25526 DVDD.n12113 DVDD.n11926 2.24164
R25527 DVDD.n12115 DVDD.n11938 2.24164
R25528 DVDD.n12117 DVDD.n11926 2.24164
R25529 DVDD.n11995 DVDD.n11938 2.24164
R25530 DVDD.n12125 DVDD.n11926 2.24164
R25531 DVDD.n12127 DVDD.n11938 2.24164
R25532 DVDD.n12129 DVDD.n11926 2.24164
R25533 DVDD.n11991 DVDD.n11938 2.24164
R25534 DVDD.n12137 DVDD.n11926 2.24164
R25535 DVDD.n12139 DVDD.n11938 2.24164
R25536 DVDD.n12141 DVDD.n11926 2.24164
R25537 DVDD.n11987 DVDD.n11938 2.24164
R25538 DVDD.n12149 DVDD.n11926 2.24164
R25539 DVDD.n12151 DVDD.n11938 2.24164
R25540 DVDD.n12153 DVDD.n11926 2.24164
R25541 DVDD.n11983 DVDD.n11938 2.24164
R25542 DVDD.n12161 DVDD.n11926 2.24164
R25543 DVDD.n12163 DVDD.n11938 2.24164
R25544 DVDD.n12165 DVDD.n11926 2.24164
R25545 DVDD.n11979 DVDD.n11938 2.24164
R25546 DVDD.n12173 DVDD.n11926 2.24164
R25547 DVDD.n12175 DVDD.n11938 2.24164
R25548 DVDD.n12177 DVDD.n11926 2.24164
R25549 DVDD.n11975 DVDD.n11938 2.24164
R25550 DVDD.n12185 DVDD.n11926 2.24164
R25551 DVDD.n12187 DVDD.n11938 2.24164
R25552 DVDD.n12189 DVDD.n11926 2.24164
R25553 DVDD.n11971 DVDD.n11938 2.24164
R25554 DVDD.n12197 DVDD.n11926 2.24164
R25555 DVDD.n12199 DVDD.n11938 2.24164
R25556 DVDD.n12201 DVDD.n11926 2.24164
R25557 DVDD.n11967 DVDD.n11938 2.24164
R25558 DVDD.n12209 DVDD.n11926 2.24164
R25559 DVDD.n12211 DVDD.n11938 2.24164
R25560 DVDD.n12213 DVDD.n11926 2.24164
R25561 DVDD.n11963 DVDD.n11938 2.24164
R25562 DVDD.n12221 DVDD.n11926 2.24164
R25563 DVDD.n12223 DVDD.n11938 2.24164
R25564 DVDD.n12225 DVDD.n11926 2.24164
R25565 DVDD.n11959 DVDD.n11938 2.24164
R25566 DVDD.n12233 DVDD.n11926 2.24164
R25567 DVDD.n12235 DVDD.n11938 2.24164
R25568 DVDD.n12237 DVDD.n11926 2.24164
R25569 DVDD.n11955 DVDD.n11938 2.24164
R25570 DVDD.n12245 DVDD.n11926 2.24164
R25571 DVDD.n12247 DVDD.n11938 2.24164
R25572 DVDD.n12249 DVDD.n11926 2.24164
R25573 DVDD.n11951 DVDD.n11938 2.24164
R25574 DVDD.n12257 DVDD.n11926 2.24164
R25575 DVDD.n12259 DVDD.n11938 2.24164
R25576 DVDD.n12261 DVDD.n11926 2.24164
R25577 DVDD.n11947 DVDD.n11938 2.24164
R25578 DVDD.n12270 DVDD.n11926 2.24164
R25579 DVDD.n12272 DVDD.n11938 2.24164
R25580 DVDD.n12274 DVDD.n11926 2.24164
R25581 DVDD.n11675 DVDD.n11581 2.24164
R25582 DVDD.n13777 DVDD.n11629 2.24164
R25583 DVDD.n11682 DVDD.n11581 2.24164
R25584 DVDD.n13777 DVDD.n11628 2.24164
R25585 DVDD.n11686 DVDD.n11581 2.24164
R25586 DVDD.n13777 DVDD.n11627 2.24164
R25587 DVDD.n11694 DVDD.n11581 2.24164
R25588 DVDD.n13777 DVDD.n11626 2.24164
R25589 DVDD.n11698 DVDD.n11581 2.24164
R25590 DVDD.n13777 DVDD.n11625 2.24164
R25591 DVDD.n11706 DVDD.n11581 2.24164
R25592 DVDD.n13777 DVDD.n11624 2.24164
R25593 DVDD.n11710 DVDD.n11581 2.24164
R25594 DVDD.n13777 DVDD.n11623 2.24164
R25595 DVDD.n11718 DVDD.n11581 2.24164
R25596 DVDD.n13777 DVDD.n11622 2.24164
R25597 DVDD.n11722 DVDD.n11581 2.24164
R25598 DVDD.n13777 DVDD.n11621 2.24164
R25599 DVDD.n11730 DVDD.n11581 2.24164
R25600 DVDD.n13777 DVDD.n11620 2.24164
R25601 DVDD.n11734 DVDD.n11581 2.24164
R25602 DVDD.n13777 DVDD.n11619 2.24164
R25603 DVDD.n11742 DVDD.n11581 2.24164
R25604 DVDD.n13777 DVDD.n11618 2.24164
R25605 DVDD.n11746 DVDD.n11581 2.24164
R25606 DVDD.n13777 DVDD.n11617 2.24164
R25607 DVDD.n11754 DVDD.n11581 2.24164
R25608 DVDD.n13777 DVDD.n11616 2.24164
R25609 DVDD.n11758 DVDD.n11581 2.24164
R25610 DVDD.n13777 DVDD.n11615 2.24164
R25611 DVDD.n11766 DVDD.n11581 2.24164
R25612 DVDD.n13777 DVDD.n11614 2.24164
R25613 DVDD.n11770 DVDD.n11581 2.24164
R25614 DVDD.n13777 DVDD.n11613 2.24164
R25615 DVDD.n11778 DVDD.n11581 2.24164
R25616 DVDD.n13777 DVDD.n11612 2.24164
R25617 DVDD.n11782 DVDD.n11581 2.24164
R25618 DVDD.n13777 DVDD.n11611 2.24164
R25619 DVDD.n11790 DVDD.n11581 2.24164
R25620 DVDD.n13777 DVDD.n11610 2.24164
R25621 DVDD.n11794 DVDD.n11581 2.24164
R25622 DVDD.n13777 DVDD.n11609 2.24164
R25623 DVDD.n11802 DVDD.n11581 2.24164
R25624 DVDD.n13777 DVDD.n11608 2.24164
R25625 DVDD.n11806 DVDD.n11581 2.24164
R25626 DVDD.n13777 DVDD.n11607 2.24164
R25627 DVDD.n11814 DVDD.n11581 2.24164
R25628 DVDD.n13777 DVDD.n11606 2.24164
R25629 DVDD.n11818 DVDD.n11581 2.24164
R25630 DVDD.n13777 DVDD.n11605 2.24164
R25631 DVDD.n11826 DVDD.n11581 2.24164
R25632 DVDD.n13777 DVDD.n11604 2.24164
R25633 DVDD.n11830 DVDD.n11581 2.24164
R25634 DVDD.n13777 DVDD.n11603 2.24164
R25635 DVDD.n11838 DVDD.n11581 2.24164
R25636 DVDD.n13777 DVDD.n11602 2.24164
R25637 DVDD.n11842 DVDD.n11581 2.24164
R25638 DVDD.n13777 DVDD.n11601 2.24164
R25639 DVDD.n11850 DVDD.n11581 2.24164
R25640 DVDD.n13777 DVDD.n11600 2.24164
R25641 DVDD.n11854 DVDD.n11581 2.24164
R25642 DVDD.n13777 DVDD.n11599 2.24164
R25643 DVDD.n11862 DVDD.n11581 2.24164
R25644 DVDD.n13777 DVDD.n11598 2.24164
R25645 DVDD.n11866 DVDD.n11581 2.24164
R25646 DVDD.n13777 DVDD.n11597 2.24164
R25647 DVDD.n11874 DVDD.n11581 2.24164
R25648 DVDD.n13777 DVDD.n11596 2.24164
R25649 DVDD.n11878 DVDD.n11581 2.24164
R25650 DVDD.n13777 DVDD.n11595 2.24164
R25651 DVDD.n11886 DVDD.n11581 2.24164
R25652 DVDD.n13777 DVDD.n11594 2.24164
R25653 DVDD.n11890 DVDD.n11581 2.24164
R25654 DVDD.n13777 DVDD.n11593 2.24164
R25655 DVDD.n11898 DVDD.n11581 2.24164
R25656 DVDD.n13777 DVDD.n11592 2.24164
R25657 DVDD.n11902 DVDD.n11581 2.24164
R25658 DVDD.n13777 DVDD.n11591 2.24164
R25659 DVDD.n11910 DVDD.n11581 2.24164
R25660 DVDD.n13777 DVDD.n11590 2.24164
R25661 DVDD.n11914 DVDD.n11581 2.24164
R25662 DVDD.n13777 DVDD.n11589 2.24164
R25663 DVDD.n13775 DVDD.n11581 2.24164
R25664 DVDD.n11321 DVDD.n11279 2.24164
R25665 DVDD.n13799 DVDD.n11274 2.24164
R25666 DVDD.n11328 DVDD.n11279 2.24164
R25667 DVDD.n13799 DVDD.n11273 2.24164
R25668 DVDD.n11332 DVDD.n11279 2.24164
R25669 DVDD.n13799 DVDD.n11272 2.24164
R25670 DVDD.n11340 DVDD.n11279 2.24164
R25671 DVDD.n13799 DVDD.n11271 2.24164
R25672 DVDD.n11344 DVDD.n11279 2.24164
R25673 DVDD.n13799 DVDD.n11270 2.24164
R25674 DVDD.n11352 DVDD.n11279 2.24164
R25675 DVDD.n13799 DVDD.n11269 2.24164
R25676 DVDD.n11356 DVDD.n11279 2.24164
R25677 DVDD.n13799 DVDD.n11268 2.24164
R25678 DVDD.n11364 DVDD.n11279 2.24164
R25679 DVDD.n13799 DVDD.n11267 2.24164
R25680 DVDD.n11368 DVDD.n11279 2.24164
R25681 DVDD.n13799 DVDD.n11266 2.24164
R25682 DVDD.n11376 DVDD.n11279 2.24164
R25683 DVDD.n13799 DVDD.n11265 2.24164
R25684 DVDD.n11380 DVDD.n11279 2.24164
R25685 DVDD.n13799 DVDD.n11264 2.24164
R25686 DVDD.n11388 DVDD.n11279 2.24164
R25687 DVDD.n13799 DVDD.n11263 2.24164
R25688 DVDD.n11392 DVDD.n11279 2.24164
R25689 DVDD.n13799 DVDD.n11262 2.24164
R25690 DVDD.n11400 DVDD.n11279 2.24164
R25691 DVDD.n13799 DVDD.n11261 2.24164
R25692 DVDD.n11404 DVDD.n11279 2.24164
R25693 DVDD.n13799 DVDD.n11260 2.24164
R25694 DVDD.n11412 DVDD.n11279 2.24164
R25695 DVDD.n13799 DVDD.n11259 2.24164
R25696 DVDD.n11416 DVDD.n11279 2.24164
R25697 DVDD.n13799 DVDD.n11258 2.24164
R25698 DVDD.n11424 DVDD.n11279 2.24164
R25699 DVDD.n13799 DVDD.n11257 2.24164
R25700 DVDD.n11428 DVDD.n11279 2.24164
R25701 DVDD.n13799 DVDD.n11256 2.24164
R25702 DVDD.n11436 DVDD.n11279 2.24164
R25703 DVDD.n13799 DVDD.n11255 2.24164
R25704 DVDD.n11440 DVDD.n11279 2.24164
R25705 DVDD.n13799 DVDD.n11254 2.24164
R25706 DVDD.n11448 DVDD.n11279 2.24164
R25707 DVDD.n13799 DVDD.n11253 2.24164
R25708 DVDD.n11452 DVDD.n11279 2.24164
R25709 DVDD.n13799 DVDD.n11252 2.24164
R25710 DVDD.n11460 DVDD.n11279 2.24164
R25711 DVDD.n13799 DVDD.n11251 2.24164
R25712 DVDD.n11464 DVDD.n11279 2.24164
R25713 DVDD.n13799 DVDD.n11250 2.24164
R25714 DVDD.n11472 DVDD.n11279 2.24164
R25715 DVDD.n13799 DVDD.n11249 2.24164
R25716 DVDD.n11476 DVDD.n11279 2.24164
R25717 DVDD.n13799 DVDD.n11248 2.24164
R25718 DVDD.n11484 DVDD.n11279 2.24164
R25719 DVDD.n13799 DVDD.n11247 2.24164
R25720 DVDD.n11488 DVDD.n11279 2.24164
R25721 DVDD.n13799 DVDD.n11246 2.24164
R25722 DVDD.n11496 DVDD.n11279 2.24164
R25723 DVDD.n13799 DVDD.n11245 2.24164
R25724 DVDD.n11500 DVDD.n11279 2.24164
R25725 DVDD.n13799 DVDD.n11244 2.24164
R25726 DVDD.n11508 DVDD.n11279 2.24164
R25727 DVDD.n13799 DVDD.n11243 2.24164
R25728 DVDD.n11512 DVDD.n11279 2.24164
R25729 DVDD.n13799 DVDD.n11242 2.24164
R25730 DVDD.n11520 DVDD.n11279 2.24164
R25731 DVDD.n13799 DVDD.n11241 2.24164
R25732 DVDD.n11524 DVDD.n11279 2.24164
R25733 DVDD.n13799 DVDD.n11240 2.24164
R25734 DVDD.n11532 DVDD.n11279 2.24164
R25735 DVDD.n13799 DVDD.n11239 2.24164
R25736 DVDD.n11536 DVDD.n11279 2.24164
R25737 DVDD.n13799 DVDD.n11238 2.24164
R25738 DVDD.n11544 DVDD.n11279 2.24164
R25739 DVDD.n13799 DVDD.n11237 2.24164
R25740 DVDD.n11548 DVDD.n11279 2.24164
R25741 DVDD.n13799 DVDD.n11236 2.24164
R25742 DVDD.n11556 DVDD.n11279 2.24164
R25743 DVDD.n13799 DVDD.n11235 2.24164
R25744 DVDD.n11560 DVDD.n11279 2.24164
R25745 DVDD.n13799 DVDD.n11234 2.24164
R25746 DVDD.n13797 DVDD.n11279 2.24164
R25747 DVDD.n14003 DVDD.n14002 2.24164
R25748 DVDD.n14000 DVDD.n11148 2.24164
R25749 DVDD.n14003 DVDD.n11102 2.24164
R25750 DVDD.n14000 DVDD.n11147 2.24164
R25751 DVDD.n14003 DVDD.n11101 2.24164
R25752 DVDD.n14000 DVDD.n11146 2.24164
R25753 DVDD.n14003 DVDD.n11100 2.24164
R25754 DVDD.n14000 DVDD.n11145 2.24164
R25755 DVDD.n14003 DVDD.n11099 2.24164
R25756 DVDD.n14000 DVDD.n11144 2.24164
R25757 DVDD.n14003 DVDD.n11098 2.24164
R25758 DVDD.n14000 DVDD.n11143 2.24164
R25759 DVDD.n14003 DVDD.n11097 2.24164
R25760 DVDD.n14000 DVDD.n11142 2.24164
R25761 DVDD.n14003 DVDD.n11096 2.24164
R25762 DVDD.n14000 DVDD.n11141 2.24164
R25763 DVDD.n14003 DVDD.n11095 2.24164
R25764 DVDD.n14000 DVDD.n11140 2.24164
R25765 DVDD.n14003 DVDD.n11094 2.24164
R25766 DVDD.n14000 DVDD.n11139 2.24164
R25767 DVDD.n14003 DVDD.n11093 2.24164
R25768 DVDD.n14000 DVDD.n11138 2.24164
R25769 DVDD.n14003 DVDD.n11092 2.24164
R25770 DVDD.n14000 DVDD.n11137 2.24164
R25771 DVDD.n14003 DVDD.n11091 2.24164
R25772 DVDD.n14000 DVDD.n11136 2.24164
R25773 DVDD.n14003 DVDD.n11090 2.24164
R25774 DVDD.n14000 DVDD.n11135 2.24164
R25775 DVDD.n14003 DVDD.n11089 2.24164
R25776 DVDD.n14000 DVDD.n11134 2.24164
R25777 DVDD.n14003 DVDD.n11088 2.24164
R25778 DVDD.n14000 DVDD.n11133 2.24164
R25779 DVDD.n14003 DVDD.n11087 2.24164
R25780 DVDD.n14000 DVDD.n11132 2.24164
R25781 DVDD.n14003 DVDD.n11086 2.24164
R25782 DVDD.n14000 DVDD.n11131 2.24164
R25783 DVDD.n14003 DVDD.n11085 2.24164
R25784 DVDD.n14000 DVDD.n11130 2.24164
R25785 DVDD.n14003 DVDD.n11084 2.24164
R25786 DVDD.n14000 DVDD.n11129 2.24164
R25787 DVDD.n14003 DVDD.n11083 2.24164
R25788 DVDD.n14000 DVDD.n11128 2.24164
R25789 DVDD.n14003 DVDD.n11082 2.24164
R25790 DVDD.n14000 DVDD.n11127 2.24164
R25791 DVDD.n14003 DVDD.n11081 2.24164
R25792 DVDD.n14000 DVDD.n11126 2.24164
R25793 DVDD.n14003 DVDD.n11080 2.24164
R25794 DVDD.n14000 DVDD.n11125 2.24164
R25795 DVDD.n14003 DVDD.n11079 2.24164
R25796 DVDD.n14000 DVDD.n11124 2.24164
R25797 DVDD.n14003 DVDD.n11078 2.24164
R25798 DVDD.n14000 DVDD.n11123 2.24164
R25799 DVDD.n14003 DVDD.n11077 2.24164
R25800 DVDD.n14000 DVDD.n11122 2.24164
R25801 DVDD.n14003 DVDD.n11076 2.24164
R25802 DVDD.n14000 DVDD.n11121 2.24164
R25803 DVDD.n14003 DVDD.n11075 2.24164
R25804 DVDD.n14000 DVDD.n11120 2.24164
R25805 DVDD.n14003 DVDD.n11074 2.24164
R25806 DVDD.n14000 DVDD.n11119 2.24164
R25807 DVDD.n14003 DVDD.n11073 2.24164
R25808 DVDD.n14000 DVDD.n11118 2.24164
R25809 DVDD.n14003 DVDD.n11072 2.24164
R25810 DVDD.n14000 DVDD.n11117 2.24164
R25811 DVDD.n14003 DVDD.n11071 2.24164
R25812 DVDD.n14000 DVDD.n11116 2.24164
R25813 DVDD.n14003 DVDD.n11070 2.24164
R25814 DVDD.n14000 DVDD.n11115 2.24164
R25815 DVDD.n14003 DVDD.n11069 2.24164
R25816 DVDD.n14000 DVDD.n11114 2.24164
R25817 DVDD.n14003 DVDD.n11068 2.24164
R25818 DVDD.n14000 DVDD.n11113 2.24164
R25819 DVDD.n14003 DVDD.n11067 2.24164
R25820 DVDD.n14000 DVDD.n11112 2.24164
R25821 DVDD.n14003 DVDD.n11066 2.24164
R25822 DVDD.n14000 DVDD.n11111 2.24164
R25823 DVDD.n14003 DVDD.n11065 2.24164
R25824 DVDD.n14000 DVDD.n11110 2.24164
R25825 DVDD.n14003 DVDD.n11064 2.24164
R25826 DVDD.n14000 DVDD.n11109 2.24164
R25827 DVDD.n14003 DVDD.n11063 2.24164
R25828 DVDD.n14000 DVDD.n11108 2.24164
R25829 DVDD.n14003 DVDD.n11062 2.24164
R25830 DVDD.n10802 DVDD.n10710 2.24164
R25831 DVDD.n10804 DVDD.n10711 2.24164
R25832 DVDD.n10806 DVDD.n10710 2.24164
R25833 DVDD.n10795 DVDD.n10711 2.24164
R25834 DVDD.n10814 DVDD.n10710 2.24164
R25835 DVDD.n10816 DVDD.n10711 2.24164
R25836 DVDD.n10818 DVDD.n10710 2.24164
R25837 DVDD.n10791 DVDD.n10711 2.24164
R25838 DVDD.n10826 DVDD.n10710 2.24164
R25839 DVDD.n10828 DVDD.n10711 2.24164
R25840 DVDD.n10830 DVDD.n10710 2.24164
R25841 DVDD.n10787 DVDD.n10711 2.24164
R25842 DVDD.n10838 DVDD.n10710 2.24164
R25843 DVDD.n10840 DVDD.n10711 2.24164
R25844 DVDD.n10842 DVDD.n10710 2.24164
R25845 DVDD.n10783 DVDD.n10711 2.24164
R25846 DVDD.n10850 DVDD.n10710 2.24164
R25847 DVDD.n10852 DVDD.n10711 2.24164
R25848 DVDD.n10854 DVDD.n10710 2.24164
R25849 DVDD.n10779 DVDD.n10711 2.24164
R25850 DVDD.n10862 DVDD.n10710 2.24164
R25851 DVDD.n10864 DVDD.n10711 2.24164
R25852 DVDD.n10866 DVDD.n10710 2.24164
R25853 DVDD.n10775 DVDD.n10711 2.24164
R25854 DVDD.n10874 DVDD.n10710 2.24164
R25855 DVDD.n10876 DVDD.n10711 2.24164
R25856 DVDD.n10878 DVDD.n10710 2.24164
R25857 DVDD.n10771 DVDD.n10711 2.24164
R25858 DVDD.n10886 DVDD.n10710 2.24164
R25859 DVDD.n10888 DVDD.n10711 2.24164
R25860 DVDD.n10890 DVDD.n10710 2.24164
R25861 DVDD.n10767 DVDD.n10711 2.24164
R25862 DVDD.n10898 DVDD.n10710 2.24164
R25863 DVDD.n10900 DVDD.n10711 2.24164
R25864 DVDD.n10902 DVDD.n10710 2.24164
R25865 DVDD.n10763 DVDD.n10711 2.24164
R25866 DVDD.n10910 DVDD.n10710 2.24164
R25867 DVDD.n10912 DVDD.n10711 2.24164
R25868 DVDD.n10914 DVDD.n10710 2.24164
R25869 DVDD.n10759 DVDD.n10711 2.24164
R25870 DVDD.n10922 DVDD.n10710 2.24164
R25871 DVDD.n10924 DVDD.n10711 2.24164
R25872 DVDD.n10926 DVDD.n10710 2.24164
R25873 DVDD.n10755 DVDD.n10711 2.24164
R25874 DVDD.n10934 DVDD.n10710 2.24164
R25875 DVDD.n10936 DVDD.n10711 2.24164
R25876 DVDD.n10938 DVDD.n10710 2.24164
R25877 DVDD.n10751 DVDD.n10711 2.24164
R25878 DVDD.n10946 DVDD.n10710 2.24164
R25879 DVDD.n10948 DVDD.n10711 2.24164
R25880 DVDD.n10950 DVDD.n10710 2.24164
R25881 DVDD.n10747 DVDD.n10711 2.24164
R25882 DVDD.n10958 DVDD.n10710 2.24164
R25883 DVDD.n10960 DVDD.n10711 2.24164
R25884 DVDD.n10962 DVDD.n10710 2.24164
R25885 DVDD.n10743 DVDD.n10711 2.24164
R25886 DVDD.n10970 DVDD.n10710 2.24164
R25887 DVDD.n10972 DVDD.n10711 2.24164
R25888 DVDD.n10974 DVDD.n10710 2.24164
R25889 DVDD.n10739 DVDD.n10711 2.24164
R25890 DVDD.n10982 DVDD.n10710 2.24164
R25891 DVDD.n10984 DVDD.n10711 2.24164
R25892 DVDD.n10986 DVDD.n10710 2.24164
R25893 DVDD.n10735 DVDD.n10711 2.24164
R25894 DVDD.n10994 DVDD.n10710 2.24164
R25895 DVDD.n10996 DVDD.n10711 2.24164
R25896 DVDD.n10998 DVDD.n10710 2.24164
R25897 DVDD.n10731 DVDD.n10711 2.24164
R25898 DVDD.n11006 DVDD.n10710 2.24164
R25899 DVDD.n11008 DVDD.n10711 2.24164
R25900 DVDD.n11010 DVDD.n10710 2.24164
R25901 DVDD.n10727 DVDD.n10711 2.24164
R25902 DVDD.n11018 DVDD.n10710 2.24164
R25903 DVDD.n11020 DVDD.n10711 2.24164
R25904 DVDD.n11022 DVDD.n10710 2.24164
R25905 DVDD.n10723 DVDD.n10711 2.24164
R25906 DVDD.n11030 DVDD.n10710 2.24164
R25907 DVDD.n11032 DVDD.n10711 2.24164
R25908 DVDD.n11034 DVDD.n10710 2.24164
R25909 DVDD.n10719 DVDD.n10711 2.24164
R25910 DVDD.n11043 DVDD.n10710 2.24164
R25911 DVDD.n11045 DVDD.n10711 2.24164
R25912 DVDD.n11047 DVDD.n10710 2.24164
R25913 DVDD.n10683 DVDD.n10642 2.24164
R25914 DVDD.n14269 DVDD.n10638 2.24164
R25915 DVDD.n14027 DVDD.n10642 2.24164
R25916 DVDD.n14269 DVDD.n10637 2.24164
R25917 DVDD.n14031 DVDD.n10642 2.24164
R25918 DVDD.n14269 DVDD.n10636 2.24164
R25919 DVDD.n14039 DVDD.n10642 2.24164
R25920 DVDD.n14269 DVDD.n10635 2.24164
R25921 DVDD.n14043 DVDD.n10642 2.24164
R25922 DVDD.n14269 DVDD.n10634 2.24164
R25923 DVDD.n14051 DVDD.n10642 2.24164
R25924 DVDD.n14269 DVDD.n10633 2.24164
R25925 DVDD.n14055 DVDD.n10642 2.24164
R25926 DVDD.n14269 DVDD.n10632 2.24164
R25927 DVDD.n14063 DVDD.n10642 2.24164
R25928 DVDD.n14269 DVDD.n10631 2.24164
R25929 DVDD.n14067 DVDD.n10642 2.24164
R25930 DVDD.n14269 DVDD.n10630 2.24164
R25931 DVDD.n14075 DVDD.n10642 2.24164
R25932 DVDD.n14269 DVDD.n10629 2.24164
R25933 DVDD.n14079 DVDD.n10642 2.24164
R25934 DVDD.n14269 DVDD.n10628 2.24164
R25935 DVDD.n14087 DVDD.n10642 2.24164
R25936 DVDD.n14269 DVDD.n10627 2.24164
R25937 DVDD.n14091 DVDD.n10642 2.24164
R25938 DVDD.n14269 DVDD.n10626 2.24164
R25939 DVDD.n14099 DVDD.n10642 2.24164
R25940 DVDD.n14269 DVDD.n10625 2.24164
R25941 DVDD.n14103 DVDD.n10642 2.24164
R25942 DVDD.n14269 DVDD.n10624 2.24164
R25943 DVDD.n14111 DVDD.n10642 2.24164
R25944 DVDD.n14269 DVDD.n10623 2.24164
R25945 DVDD.n14115 DVDD.n10642 2.24164
R25946 DVDD.n14269 DVDD.n10622 2.24164
R25947 DVDD.n14123 DVDD.n10642 2.24164
R25948 DVDD.n14269 DVDD.n10621 2.24164
R25949 DVDD.n14127 DVDD.n10642 2.24164
R25950 DVDD.n14269 DVDD.n10620 2.24164
R25951 DVDD.n14135 DVDD.n10642 2.24164
R25952 DVDD.n14269 DVDD.n10619 2.24164
R25953 DVDD.n14139 DVDD.n10642 2.24164
R25954 DVDD.n14269 DVDD.n10618 2.24164
R25955 DVDD.n14147 DVDD.n10642 2.24164
R25956 DVDD.n14269 DVDD.n10617 2.24164
R25957 DVDD.n14151 DVDD.n10642 2.24164
R25958 DVDD.n14269 DVDD.n10616 2.24164
R25959 DVDD.n14159 DVDD.n10642 2.24164
R25960 DVDD.n14269 DVDD.n10615 2.24164
R25961 DVDD.n14163 DVDD.n10642 2.24164
R25962 DVDD.n14269 DVDD.n10614 2.24164
R25963 DVDD.n14171 DVDD.n10642 2.24164
R25964 DVDD.n14269 DVDD.n10613 2.24164
R25965 DVDD.n14175 DVDD.n10642 2.24164
R25966 DVDD.n14269 DVDD.n10612 2.24164
R25967 DVDD.n14183 DVDD.n10642 2.24164
R25968 DVDD.n14269 DVDD.n10611 2.24164
R25969 DVDD.n14187 DVDD.n10642 2.24164
R25970 DVDD.n14269 DVDD.n10610 2.24164
R25971 DVDD.n14195 DVDD.n10642 2.24164
R25972 DVDD.n14269 DVDD.n10609 2.24164
R25973 DVDD.n14199 DVDD.n10642 2.24164
R25974 DVDD.n14269 DVDD.n10608 2.24164
R25975 DVDD.n14207 DVDD.n10642 2.24164
R25976 DVDD.n14269 DVDD.n10607 2.24164
R25977 DVDD.n14211 DVDD.n10642 2.24164
R25978 DVDD.n14269 DVDD.n10606 2.24164
R25979 DVDD.n14219 DVDD.n10642 2.24164
R25980 DVDD.n14269 DVDD.n10605 2.24164
R25981 DVDD.n14223 DVDD.n10642 2.24164
R25982 DVDD.n14269 DVDD.n10604 2.24164
R25983 DVDD.n14231 DVDD.n10642 2.24164
R25984 DVDD.n14269 DVDD.n10603 2.24164
R25985 DVDD.n14235 DVDD.n10642 2.24164
R25986 DVDD.n14269 DVDD.n10602 2.24164
R25987 DVDD.n14243 DVDD.n10642 2.24164
R25988 DVDD.n14269 DVDD.n10601 2.24164
R25989 DVDD.n14247 DVDD.n10642 2.24164
R25990 DVDD.n14269 DVDD.n10600 2.24164
R25991 DVDD.n14255 DVDD.n10642 2.24164
R25992 DVDD.n14269 DVDD.n10599 2.24164
R25993 DVDD.n14259 DVDD.n10642 2.24164
R25994 DVDD.n14269 DVDD.n10598 2.24164
R25995 DVDD.n14267 DVDD.n10642 2.24164
R25996 DVDD.n14284 DVDD.n14283 2.24164
R25997 DVDD.n14281 DVDD.n10327 2.24164
R25998 DVDD.n14284 DVDD.n10282 2.24164
R25999 DVDD.n14281 DVDD.n10326 2.24164
R26000 DVDD.n14284 DVDD.n10281 2.24164
R26001 DVDD.n14281 DVDD.n10325 2.24164
R26002 DVDD.n14284 DVDD.n10280 2.24164
R26003 DVDD.n14281 DVDD.n10324 2.24164
R26004 DVDD.n14284 DVDD.n10279 2.24164
R26005 DVDD.n14281 DVDD.n10323 2.24164
R26006 DVDD.n14284 DVDD.n10278 2.24164
R26007 DVDD.n14281 DVDD.n10322 2.24164
R26008 DVDD.n14284 DVDD.n10277 2.24164
R26009 DVDD.n14281 DVDD.n10321 2.24164
R26010 DVDD.n14284 DVDD.n10276 2.24164
R26011 DVDD.n14281 DVDD.n10320 2.24164
R26012 DVDD.n14284 DVDD.n10275 2.24164
R26013 DVDD.n14281 DVDD.n10319 2.24164
R26014 DVDD.n14284 DVDD.n10274 2.24164
R26015 DVDD.n14281 DVDD.n10318 2.24164
R26016 DVDD.n14284 DVDD.n10273 2.24164
R26017 DVDD.n14281 DVDD.n10317 2.24164
R26018 DVDD.n14284 DVDD.n10272 2.24164
R26019 DVDD.n14281 DVDD.n10316 2.24164
R26020 DVDD.n14284 DVDD.n10271 2.24164
R26021 DVDD.n14281 DVDD.n10315 2.24164
R26022 DVDD.n14284 DVDD.n10270 2.24164
R26023 DVDD.n14281 DVDD.n10314 2.24164
R26024 DVDD.n14284 DVDD.n10269 2.24164
R26025 DVDD.n14281 DVDD.n10313 2.24164
R26026 DVDD.n14284 DVDD.n10268 2.24164
R26027 DVDD.n14281 DVDD.n10312 2.24164
R26028 DVDD.n14284 DVDD.n10267 2.24164
R26029 DVDD.n14281 DVDD.n10311 2.24164
R26030 DVDD.n14284 DVDD.n10266 2.24164
R26031 DVDD.n14281 DVDD.n10310 2.24164
R26032 DVDD.n14284 DVDD.n10265 2.24164
R26033 DVDD.n14281 DVDD.n10309 2.24164
R26034 DVDD.n14284 DVDD.n10264 2.24164
R26035 DVDD.n14281 DVDD.n10308 2.24164
R26036 DVDD.n14284 DVDD.n10263 2.24164
R26037 DVDD.n14281 DVDD.n10307 2.24164
R26038 DVDD.n14284 DVDD.n10262 2.24164
R26039 DVDD.n14281 DVDD.n10306 2.24164
R26040 DVDD.n14284 DVDD.n10261 2.24164
R26041 DVDD.n14281 DVDD.n10305 2.24164
R26042 DVDD.n14284 DVDD.n10260 2.24164
R26043 DVDD.n14281 DVDD.n10304 2.24164
R26044 DVDD.n14284 DVDD.n10259 2.24164
R26045 DVDD.n14281 DVDD.n10303 2.24164
R26046 DVDD.n14284 DVDD.n10258 2.24164
R26047 DVDD.n14281 DVDD.n10302 2.24164
R26048 DVDD.n14284 DVDD.n10257 2.24164
R26049 DVDD.n14281 DVDD.n10301 2.24164
R26050 DVDD.n14284 DVDD.n10256 2.24164
R26051 DVDD.n14281 DVDD.n10300 2.24164
R26052 DVDD.n14284 DVDD.n10255 2.24164
R26053 DVDD.n14281 DVDD.n10299 2.24164
R26054 DVDD.n14284 DVDD.n10254 2.24164
R26055 DVDD.n14281 DVDD.n10298 2.24164
R26056 DVDD.n14284 DVDD.n10253 2.24164
R26057 DVDD.n14281 DVDD.n10297 2.24164
R26058 DVDD.n14284 DVDD.n10252 2.24164
R26059 DVDD.n14281 DVDD.n10296 2.24164
R26060 DVDD.n14284 DVDD.n10251 2.24164
R26061 DVDD.n14281 DVDD.n10295 2.24164
R26062 DVDD.n14284 DVDD.n10250 2.24164
R26063 DVDD.n14281 DVDD.n10294 2.24164
R26064 DVDD.n14284 DVDD.n10249 2.24164
R26065 DVDD.n14281 DVDD.n10293 2.24164
R26066 DVDD.n14284 DVDD.n10248 2.24164
R26067 DVDD.n14281 DVDD.n10292 2.24164
R26068 DVDD.n14284 DVDD.n10247 2.24164
R26069 DVDD.n14281 DVDD.n10291 2.24164
R26070 DVDD.n14284 DVDD.n10246 2.24164
R26071 DVDD.n14281 DVDD.n10290 2.24164
R26072 DVDD.n14284 DVDD.n10245 2.24164
R26073 DVDD.n14281 DVDD.n10289 2.24164
R26074 DVDD.n14284 DVDD.n10244 2.24164
R26075 DVDD.n14281 DVDD.n10288 2.24164
R26076 DVDD.n14284 DVDD.n10243 2.24164
R26077 DVDD.n14281 DVDD.n10287 2.24164
R26078 DVDD.n14284 DVDD.n10242 2.24164
R26079 DVDD.n8946 DVDD.n8609 2.24164
R26080 DVDD.n8944 DVDD.n8610 2.24164
R26081 DVDD.n8617 DVDD.n8609 2.24164
R26082 DVDD.n8622 DVDD.n8610 2.24164
R26083 DVDD.n8936 DVDD.n8609 2.24164
R26084 DVDD.n8934 DVDD.n8610 2.24164
R26085 DVDD.n8623 DVDD.n8609 2.24164
R26086 DVDD.n8628 DVDD.n8610 2.24164
R26087 DVDD.n8926 DVDD.n8609 2.24164
R26088 DVDD.n8924 DVDD.n8610 2.24164
R26089 DVDD.n8629 DVDD.n8609 2.24164
R26090 DVDD.n8634 DVDD.n8610 2.24164
R26091 DVDD.n8916 DVDD.n8609 2.24164
R26092 DVDD.n8914 DVDD.n8610 2.24164
R26093 DVDD.n8635 DVDD.n8609 2.24164
R26094 DVDD.n8640 DVDD.n8610 2.24164
R26095 DVDD.n8906 DVDD.n8609 2.24164
R26096 DVDD.n8904 DVDD.n8610 2.24164
R26097 DVDD.n8641 DVDD.n8609 2.24164
R26098 DVDD.n8646 DVDD.n8610 2.24164
R26099 DVDD.n8896 DVDD.n8609 2.24164
R26100 DVDD.n8894 DVDD.n8610 2.24164
R26101 DVDD.n8647 DVDD.n8609 2.24164
R26102 DVDD.n8652 DVDD.n8610 2.24164
R26103 DVDD.n8886 DVDD.n8609 2.24164
R26104 DVDD.n8884 DVDD.n8610 2.24164
R26105 DVDD.n8653 DVDD.n8609 2.24164
R26106 DVDD.n8658 DVDD.n8610 2.24164
R26107 DVDD.n8876 DVDD.n8609 2.24164
R26108 DVDD.n8874 DVDD.n8610 2.24164
R26109 DVDD.n8659 DVDD.n8609 2.24164
R26110 DVDD.n8664 DVDD.n8610 2.24164
R26111 DVDD.n8866 DVDD.n8609 2.24164
R26112 DVDD.n8864 DVDD.n8610 2.24164
R26113 DVDD.n8665 DVDD.n8609 2.24164
R26114 DVDD.n8670 DVDD.n8610 2.24164
R26115 DVDD.n8856 DVDD.n8609 2.24164
R26116 DVDD.n8854 DVDD.n8610 2.24164
R26117 DVDD.n8671 DVDD.n8609 2.24164
R26118 DVDD.n8676 DVDD.n8610 2.24164
R26119 DVDD.n8846 DVDD.n8609 2.24164
R26120 DVDD.n8844 DVDD.n8610 2.24164
R26121 DVDD.n8677 DVDD.n8609 2.24164
R26122 DVDD.n8682 DVDD.n8610 2.24164
R26123 DVDD.n8836 DVDD.n8609 2.24164
R26124 DVDD.n8834 DVDD.n8610 2.24164
R26125 DVDD.n8683 DVDD.n8609 2.24164
R26126 DVDD.n8688 DVDD.n8610 2.24164
R26127 DVDD.n8826 DVDD.n8609 2.24164
R26128 DVDD.n8824 DVDD.n8610 2.24164
R26129 DVDD.n8689 DVDD.n8609 2.24164
R26130 DVDD.n8694 DVDD.n8610 2.24164
R26131 DVDD.n8816 DVDD.n8609 2.24164
R26132 DVDD.n8814 DVDD.n8610 2.24164
R26133 DVDD.n8695 DVDD.n8609 2.24164
R26134 DVDD.n8700 DVDD.n8610 2.24164
R26135 DVDD.n8806 DVDD.n8609 2.24164
R26136 DVDD.n8804 DVDD.n8610 2.24164
R26137 DVDD.n8701 DVDD.n8609 2.24164
R26138 DVDD.n8706 DVDD.n8610 2.24164
R26139 DVDD.n8796 DVDD.n8609 2.24164
R26140 DVDD.n8794 DVDD.n8610 2.24164
R26141 DVDD.n8707 DVDD.n8609 2.24164
R26142 DVDD.n8712 DVDD.n8610 2.24164
R26143 DVDD.n8786 DVDD.n8609 2.24164
R26144 DVDD.n8784 DVDD.n8610 2.24164
R26145 DVDD.n8713 DVDD.n8609 2.24164
R26146 DVDD.n8718 DVDD.n8610 2.24164
R26147 DVDD.n8776 DVDD.n8609 2.24164
R26148 DVDD.n8774 DVDD.n8610 2.24164
R26149 DVDD.n8719 DVDD.n8609 2.24164
R26150 DVDD.n8724 DVDD.n8610 2.24164
R26151 DVDD.n8766 DVDD.n8609 2.24164
R26152 DVDD.n8764 DVDD.n8610 2.24164
R26153 DVDD.n8725 DVDD.n8609 2.24164
R26154 DVDD.n8730 DVDD.n8610 2.24164
R26155 DVDD.n8756 DVDD.n8609 2.24164
R26156 DVDD.n8754 DVDD.n8610 2.24164
R26157 DVDD.n8731 DVDD.n8609 2.24164
R26158 DVDD.n8736 DVDD.n8610 2.24164
R26159 DVDD.n8746 DVDD.n8609 2.24164
R26160 DVDD.n8744 DVDD.n8610 2.24164
R26161 DVDD.n8737 DVDD.n8609 2.24164
R26162 DVDD.n8350 DVDD.n8258 2.24164
R26163 DVDD.n8352 DVDD.n8259 2.24164
R26164 DVDD.n8354 DVDD.n8258 2.24164
R26165 DVDD.n8343 DVDD.n8259 2.24164
R26166 DVDD.n8362 DVDD.n8258 2.24164
R26167 DVDD.n8364 DVDD.n8259 2.24164
R26168 DVDD.n8366 DVDD.n8258 2.24164
R26169 DVDD.n8339 DVDD.n8259 2.24164
R26170 DVDD.n8374 DVDD.n8258 2.24164
R26171 DVDD.n8376 DVDD.n8259 2.24164
R26172 DVDD.n8378 DVDD.n8258 2.24164
R26173 DVDD.n8335 DVDD.n8259 2.24164
R26174 DVDD.n8386 DVDD.n8258 2.24164
R26175 DVDD.n8388 DVDD.n8259 2.24164
R26176 DVDD.n8390 DVDD.n8258 2.24164
R26177 DVDD.n8331 DVDD.n8259 2.24164
R26178 DVDD.n8398 DVDD.n8258 2.24164
R26179 DVDD.n8400 DVDD.n8259 2.24164
R26180 DVDD.n8402 DVDD.n8258 2.24164
R26181 DVDD.n8327 DVDD.n8259 2.24164
R26182 DVDD.n8410 DVDD.n8258 2.24164
R26183 DVDD.n8412 DVDD.n8259 2.24164
R26184 DVDD.n8414 DVDD.n8258 2.24164
R26185 DVDD.n8323 DVDD.n8259 2.24164
R26186 DVDD.n8422 DVDD.n8258 2.24164
R26187 DVDD.n8424 DVDD.n8259 2.24164
R26188 DVDD.n8426 DVDD.n8258 2.24164
R26189 DVDD.n8319 DVDD.n8259 2.24164
R26190 DVDD.n8434 DVDD.n8258 2.24164
R26191 DVDD.n8436 DVDD.n8259 2.24164
R26192 DVDD.n8438 DVDD.n8258 2.24164
R26193 DVDD.n8315 DVDD.n8259 2.24164
R26194 DVDD.n8446 DVDD.n8258 2.24164
R26195 DVDD.n8448 DVDD.n8259 2.24164
R26196 DVDD.n8450 DVDD.n8258 2.24164
R26197 DVDD.n8311 DVDD.n8259 2.24164
R26198 DVDD.n8458 DVDD.n8258 2.24164
R26199 DVDD.n8460 DVDD.n8259 2.24164
R26200 DVDD.n8462 DVDD.n8258 2.24164
R26201 DVDD.n8307 DVDD.n8259 2.24164
R26202 DVDD.n8470 DVDD.n8258 2.24164
R26203 DVDD.n8472 DVDD.n8259 2.24164
R26204 DVDD.n8474 DVDD.n8258 2.24164
R26205 DVDD.n8303 DVDD.n8259 2.24164
R26206 DVDD.n8482 DVDD.n8258 2.24164
R26207 DVDD.n8484 DVDD.n8259 2.24164
R26208 DVDD.n8486 DVDD.n8258 2.24164
R26209 DVDD.n8299 DVDD.n8259 2.24164
R26210 DVDD.n8494 DVDD.n8258 2.24164
R26211 DVDD.n8496 DVDD.n8259 2.24164
R26212 DVDD.n8498 DVDD.n8258 2.24164
R26213 DVDD.n8295 DVDD.n8259 2.24164
R26214 DVDD.n8506 DVDD.n8258 2.24164
R26215 DVDD.n8508 DVDD.n8259 2.24164
R26216 DVDD.n8510 DVDD.n8258 2.24164
R26217 DVDD.n8291 DVDD.n8259 2.24164
R26218 DVDD.n8518 DVDD.n8258 2.24164
R26219 DVDD.n8520 DVDD.n8259 2.24164
R26220 DVDD.n8522 DVDD.n8258 2.24164
R26221 DVDD.n8287 DVDD.n8259 2.24164
R26222 DVDD.n8530 DVDD.n8258 2.24164
R26223 DVDD.n8532 DVDD.n8259 2.24164
R26224 DVDD.n8534 DVDD.n8258 2.24164
R26225 DVDD.n8283 DVDD.n8259 2.24164
R26226 DVDD.n8542 DVDD.n8258 2.24164
R26227 DVDD.n8544 DVDD.n8259 2.24164
R26228 DVDD.n8546 DVDD.n8258 2.24164
R26229 DVDD.n8279 DVDD.n8259 2.24164
R26230 DVDD.n8554 DVDD.n8258 2.24164
R26231 DVDD.n8556 DVDD.n8259 2.24164
R26232 DVDD.n8558 DVDD.n8258 2.24164
R26233 DVDD.n8275 DVDD.n8259 2.24164
R26234 DVDD.n8566 DVDD.n8258 2.24164
R26235 DVDD.n8568 DVDD.n8259 2.24164
R26236 DVDD.n8570 DVDD.n8258 2.24164
R26237 DVDD.n8271 DVDD.n8259 2.24164
R26238 DVDD.n8578 DVDD.n8258 2.24164
R26239 DVDD.n8580 DVDD.n8259 2.24164
R26240 DVDD.n8582 DVDD.n8258 2.24164
R26241 DVDD.n8267 DVDD.n8259 2.24164
R26242 DVDD.n8591 DVDD.n8258 2.24164
R26243 DVDD.n8593 DVDD.n8259 2.24164
R26244 DVDD.n8595 DVDD.n8258 2.24164
R26245 DVDD.n8247 DVDD.n8155 2.24164
R26246 DVDD.n14559 DVDD.n8203 2.24164
R26247 DVDD.n14317 DVDD.n8155 2.24164
R26248 DVDD.n14559 DVDD.n8202 2.24164
R26249 DVDD.n14321 DVDD.n8155 2.24164
R26250 DVDD.n14559 DVDD.n8201 2.24164
R26251 DVDD.n14329 DVDD.n8155 2.24164
R26252 DVDD.n14559 DVDD.n8200 2.24164
R26253 DVDD.n14333 DVDD.n8155 2.24164
R26254 DVDD.n14559 DVDD.n8199 2.24164
R26255 DVDD.n14341 DVDD.n8155 2.24164
R26256 DVDD.n14559 DVDD.n8198 2.24164
R26257 DVDD.n14345 DVDD.n8155 2.24164
R26258 DVDD.n14559 DVDD.n8197 2.24164
R26259 DVDD.n14353 DVDD.n8155 2.24164
R26260 DVDD.n14559 DVDD.n8196 2.24164
R26261 DVDD.n14357 DVDD.n8155 2.24164
R26262 DVDD.n14559 DVDD.n8195 2.24164
R26263 DVDD.n14365 DVDD.n8155 2.24164
R26264 DVDD.n14559 DVDD.n8194 2.24164
R26265 DVDD.n14369 DVDD.n8155 2.24164
R26266 DVDD.n14559 DVDD.n8193 2.24164
R26267 DVDD.n14377 DVDD.n8155 2.24164
R26268 DVDD.n14559 DVDD.n8192 2.24164
R26269 DVDD.n14381 DVDD.n8155 2.24164
R26270 DVDD.n14559 DVDD.n8191 2.24164
R26271 DVDD.n14389 DVDD.n8155 2.24164
R26272 DVDD.n14559 DVDD.n8190 2.24164
R26273 DVDD.n14393 DVDD.n8155 2.24164
R26274 DVDD.n14559 DVDD.n8189 2.24164
R26275 DVDD.n14401 DVDD.n8155 2.24164
R26276 DVDD.n14559 DVDD.n8188 2.24164
R26277 DVDD.n14405 DVDD.n8155 2.24164
R26278 DVDD.n14559 DVDD.n8187 2.24164
R26279 DVDD.n14413 DVDD.n8155 2.24164
R26280 DVDD.n14559 DVDD.n8186 2.24164
R26281 DVDD.n14417 DVDD.n8155 2.24164
R26282 DVDD.n14559 DVDD.n8185 2.24164
R26283 DVDD.n14425 DVDD.n8155 2.24164
R26284 DVDD.n14559 DVDD.n8184 2.24164
R26285 DVDD.n14429 DVDD.n8155 2.24164
R26286 DVDD.n14559 DVDD.n8183 2.24164
R26287 DVDD.n14437 DVDD.n8155 2.24164
R26288 DVDD.n14559 DVDD.n8182 2.24164
R26289 DVDD.n14441 DVDD.n8155 2.24164
R26290 DVDD.n14559 DVDD.n8181 2.24164
R26291 DVDD.n14449 DVDD.n8155 2.24164
R26292 DVDD.n14559 DVDD.n8180 2.24164
R26293 DVDD.n14453 DVDD.n8155 2.24164
R26294 DVDD.n14559 DVDD.n8179 2.24164
R26295 DVDD.n14461 DVDD.n8155 2.24164
R26296 DVDD.n14559 DVDD.n8178 2.24164
R26297 DVDD.n14465 DVDD.n8155 2.24164
R26298 DVDD.n14559 DVDD.n8177 2.24164
R26299 DVDD.n14473 DVDD.n8155 2.24164
R26300 DVDD.n14559 DVDD.n8176 2.24164
R26301 DVDD.n14477 DVDD.n8155 2.24164
R26302 DVDD.n14559 DVDD.n8175 2.24164
R26303 DVDD.n14485 DVDD.n8155 2.24164
R26304 DVDD.n14559 DVDD.n8174 2.24164
R26305 DVDD.n14489 DVDD.n8155 2.24164
R26306 DVDD.n14559 DVDD.n8173 2.24164
R26307 DVDD.n14497 DVDD.n8155 2.24164
R26308 DVDD.n14559 DVDD.n8172 2.24164
R26309 DVDD.n14501 DVDD.n8155 2.24164
R26310 DVDD.n14559 DVDD.n8171 2.24164
R26311 DVDD.n14509 DVDD.n8155 2.24164
R26312 DVDD.n14559 DVDD.n8170 2.24164
R26313 DVDD.n14513 DVDD.n8155 2.24164
R26314 DVDD.n14559 DVDD.n8169 2.24164
R26315 DVDD.n14521 DVDD.n8155 2.24164
R26316 DVDD.n14559 DVDD.n8168 2.24164
R26317 DVDD.n14525 DVDD.n8155 2.24164
R26318 DVDD.n14559 DVDD.n8167 2.24164
R26319 DVDD.n14533 DVDD.n8155 2.24164
R26320 DVDD.n14559 DVDD.n8166 2.24164
R26321 DVDD.n14537 DVDD.n8155 2.24164
R26322 DVDD.n14559 DVDD.n8165 2.24164
R26323 DVDD.n14545 DVDD.n8155 2.24164
R26324 DVDD.n14559 DVDD.n8164 2.24164
R26325 DVDD.n14549 DVDD.n8155 2.24164
R26326 DVDD.n14559 DVDD.n8163 2.24164
R26327 DVDD.n14557 DVDD.n8155 2.24164
R26328 DVDD.n8130 DVDD.n8089 2.24164
R26329 DVDD.n14825 DVDD.n8085 2.24164
R26330 DVDD.n14583 DVDD.n8089 2.24164
R26331 DVDD.n14825 DVDD.n8084 2.24164
R26332 DVDD.n14587 DVDD.n8089 2.24164
R26333 DVDD.n14825 DVDD.n8083 2.24164
R26334 DVDD.n14595 DVDD.n8089 2.24164
R26335 DVDD.n14825 DVDD.n8082 2.24164
R26336 DVDD.n14599 DVDD.n8089 2.24164
R26337 DVDD.n14825 DVDD.n8081 2.24164
R26338 DVDD.n14607 DVDD.n8089 2.24164
R26339 DVDD.n14825 DVDD.n8080 2.24164
R26340 DVDD.n14611 DVDD.n8089 2.24164
R26341 DVDD.n14825 DVDD.n8079 2.24164
R26342 DVDD.n14619 DVDD.n8089 2.24164
R26343 DVDD.n14825 DVDD.n8078 2.24164
R26344 DVDD.n14623 DVDD.n8089 2.24164
R26345 DVDD.n14825 DVDD.n8077 2.24164
R26346 DVDD.n14631 DVDD.n8089 2.24164
R26347 DVDD.n14825 DVDD.n8076 2.24164
R26348 DVDD.n14635 DVDD.n8089 2.24164
R26349 DVDD.n14825 DVDD.n8075 2.24164
R26350 DVDD.n14643 DVDD.n8089 2.24164
R26351 DVDD.n14825 DVDD.n8074 2.24164
R26352 DVDD.n14647 DVDD.n8089 2.24164
R26353 DVDD.n14825 DVDD.n8073 2.24164
R26354 DVDD.n14655 DVDD.n8089 2.24164
R26355 DVDD.n14825 DVDD.n8072 2.24164
R26356 DVDD.n14659 DVDD.n8089 2.24164
R26357 DVDD.n14825 DVDD.n8071 2.24164
R26358 DVDD.n14667 DVDD.n8089 2.24164
R26359 DVDD.n14825 DVDD.n8070 2.24164
R26360 DVDD.n14671 DVDD.n8089 2.24164
R26361 DVDD.n14825 DVDD.n8069 2.24164
R26362 DVDD.n14679 DVDD.n8089 2.24164
R26363 DVDD.n14825 DVDD.n8068 2.24164
R26364 DVDD.n14683 DVDD.n8089 2.24164
R26365 DVDD.n14825 DVDD.n8067 2.24164
R26366 DVDD.n14691 DVDD.n8089 2.24164
R26367 DVDD.n14825 DVDD.n8066 2.24164
R26368 DVDD.n14695 DVDD.n8089 2.24164
R26369 DVDD.n14825 DVDD.n8065 2.24164
R26370 DVDD.n14703 DVDD.n8089 2.24164
R26371 DVDD.n14825 DVDD.n8064 2.24164
R26372 DVDD.n14707 DVDD.n8089 2.24164
R26373 DVDD.n14825 DVDD.n8063 2.24164
R26374 DVDD.n14715 DVDD.n8089 2.24164
R26375 DVDD.n14825 DVDD.n8062 2.24164
R26376 DVDD.n14719 DVDD.n8089 2.24164
R26377 DVDD.n14825 DVDD.n8061 2.24164
R26378 DVDD.n14727 DVDD.n8089 2.24164
R26379 DVDD.n14825 DVDD.n8060 2.24164
R26380 DVDD.n14731 DVDD.n8089 2.24164
R26381 DVDD.n14825 DVDD.n8059 2.24164
R26382 DVDD.n14739 DVDD.n8089 2.24164
R26383 DVDD.n14825 DVDD.n8058 2.24164
R26384 DVDD.n14743 DVDD.n8089 2.24164
R26385 DVDD.n14825 DVDD.n8057 2.24164
R26386 DVDD.n14751 DVDD.n8089 2.24164
R26387 DVDD.n14825 DVDD.n8056 2.24164
R26388 DVDD.n14755 DVDD.n8089 2.24164
R26389 DVDD.n14825 DVDD.n8055 2.24164
R26390 DVDD.n14763 DVDD.n8089 2.24164
R26391 DVDD.n14825 DVDD.n8054 2.24164
R26392 DVDD.n14767 DVDD.n8089 2.24164
R26393 DVDD.n14825 DVDD.n8053 2.24164
R26394 DVDD.n14775 DVDD.n8089 2.24164
R26395 DVDD.n14825 DVDD.n8052 2.24164
R26396 DVDD.n14779 DVDD.n8089 2.24164
R26397 DVDD.n14825 DVDD.n8051 2.24164
R26398 DVDD.n14787 DVDD.n8089 2.24164
R26399 DVDD.n14825 DVDD.n8050 2.24164
R26400 DVDD.n14791 DVDD.n8089 2.24164
R26401 DVDD.n14825 DVDD.n8049 2.24164
R26402 DVDD.n14799 DVDD.n8089 2.24164
R26403 DVDD.n14825 DVDD.n8048 2.24164
R26404 DVDD.n14803 DVDD.n8089 2.24164
R26405 DVDD.n14825 DVDD.n8047 2.24164
R26406 DVDD.n14811 DVDD.n8089 2.24164
R26407 DVDD.n14825 DVDD.n8046 2.24164
R26408 DVDD.n14815 DVDD.n8089 2.24164
R26409 DVDD.n14825 DVDD.n8045 2.24164
R26410 DVDD.n14823 DVDD.n8089 2.24164
R26411 DVDD.n14840 DVDD.n14839 2.24164
R26412 DVDD.n14837 DVDD.n7774 2.24164
R26413 DVDD.n14840 DVDD.n7729 2.24164
R26414 DVDD.n14837 DVDD.n7773 2.24164
R26415 DVDD.n14840 DVDD.n7728 2.24164
R26416 DVDD.n14837 DVDD.n7772 2.24164
R26417 DVDD.n14840 DVDD.n7727 2.24164
R26418 DVDD.n14837 DVDD.n7771 2.24164
R26419 DVDD.n14840 DVDD.n7726 2.24164
R26420 DVDD.n14837 DVDD.n7770 2.24164
R26421 DVDD.n14840 DVDD.n7725 2.24164
R26422 DVDD.n14837 DVDD.n7769 2.24164
R26423 DVDD.n14840 DVDD.n7724 2.24164
R26424 DVDD.n14837 DVDD.n7768 2.24164
R26425 DVDD.n14840 DVDD.n7723 2.24164
R26426 DVDD.n14837 DVDD.n7767 2.24164
R26427 DVDD.n14840 DVDD.n7722 2.24164
R26428 DVDD.n14837 DVDD.n7766 2.24164
R26429 DVDD.n14840 DVDD.n7721 2.24164
R26430 DVDD.n14837 DVDD.n7765 2.24164
R26431 DVDD.n14840 DVDD.n7720 2.24164
R26432 DVDD.n14837 DVDD.n7764 2.24164
R26433 DVDD.n14840 DVDD.n7719 2.24164
R26434 DVDD.n14837 DVDD.n7763 2.24164
R26435 DVDD.n14840 DVDD.n7718 2.24164
R26436 DVDD.n14837 DVDD.n7762 2.24164
R26437 DVDD.n14840 DVDD.n7717 2.24164
R26438 DVDD.n14837 DVDD.n7761 2.24164
R26439 DVDD.n14840 DVDD.n7716 2.24164
R26440 DVDD.n14837 DVDD.n7760 2.24164
R26441 DVDD.n14840 DVDD.n7715 2.24164
R26442 DVDD.n14837 DVDD.n7759 2.24164
R26443 DVDD.n14840 DVDD.n7714 2.24164
R26444 DVDD.n14837 DVDD.n7758 2.24164
R26445 DVDD.n14840 DVDD.n7713 2.24164
R26446 DVDD.n14837 DVDD.n7757 2.24164
R26447 DVDD.n14840 DVDD.n7712 2.24164
R26448 DVDD.n14837 DVDD.n7756 2.24164
R26449 DVDD.n14840 DVDD.n7711 2.24164
R26450 DVDD.n14837 DVDD.n7755 2.24164
R26451 DVDD.n14840 DVDD.n7710 2.24164
R26452 DVDD.n14837 DVDD.n7754 2.24164
R26453 DVDD.n14840 DVDD.n7709 2.24164
R26454 DVDD.n14837 DVDD.n7753 2.24164
R26455 DVDD.n14840 DVDD.n7708 2.24164
R26456 DVDD.n14837 DVDD.n7752 2.24164
R26457 DVDD.n14840 DVDD.n7707 2.24164
R26458 DVDD.n14837 DVDD.n7751 2.24164
R26459 DVDD.n14840 DVDD.n7706 2.24164
R26460 DVDD.n14837 DVDD.n7750 2.24164
R26461 DVDD.n14840 DVDD.n7705 2.24164
R26462 DVDD.n14837 DVDD.n7749 2.24164
R26463 DVDD.n14840 DVDD.n7704 2.24164
R26464 DVDD.n14837 DVDD.n7748 2.24164
R26465 DVDD.n14840 DVDD.n7703 2.24164
R26466 DVDD.n14837 DVDD.n7747 2.24164
R26467 DVDD.n14840 DVDD.n7702 2.24164
R26468 DVDD.n14837 DVDD.n7746 2.24164
R26469 DVDD.n14840 DVDD.n7701 2.24164
R26470 DVDD.n14837 DVDD.n7745 2.24164
R26471 DVDD.n14840 DVDD.n7700 2.24164
R26472 DVDD.n14837 DVDD.n7744 2.24164
R26473 DVDD.n14840 DVDD.n7699 2.24164
R26474 DVDD.n14837 DVDD.n7743 2.24164
R26475 DVDD.n14840 DVDD.n7698 2.24164
R26476 DVDD.n14837 DVDD.n7742 2.24164
R26477 DVDD.n14840 DVDD.n7697 2.24164
R26478 DVDD.n14837 DVDD.n7741 2.24164
R26479 DVDD.n14840 DVDD.n7696 2.24164
R26480 DVDD.n14837 DVDD.n7740 2.24164
R26481 DVDD.n14840 DVDD.n7695 2.24164
R26482 DVDD.n14837 DVDD.n7739 2.24164
R26483 DVDD.n14840 DVDD.n7694 2.24164
R26484 DVDD.n14837 DVDD.n7738 2.24164
R26485 DVDD.n14840 DVDD.n7693 2.24164
R26486 DVDD.n14837 DVDD.n7737 2.24164
R26487 DVDD.n14840 DVDD.n7692 2.24164
R26488 DVDD.n14837 DVDD.n7736 2.24164
R26489 DVDD.n14840 DVDD.n7691 2.24164
R26490 DVDD.n14837 DVDD.n7735 2.24164
R26491 DVDD.n14840 DVDD.n7690 2.24164
R26492 DVDD.n14837 DVDD.n7734 2.24164
R26493 DVDD.n14840 DVDD.n7689 2.24164
R26494 DVDD.n9558 DVDD.n9557 2.24164
R26495 DVDD.n9266 DVDD.n7679 2.24164
R26496 DVDD.n9558 DVDD.n9263 2.24164
R26497 DVDD.n9548 DVDD.n7679 2.24164
R26498 DVDD.n9558 DVDD.n9262 2.24164
R26499 DVDD.n9543 DVDD.n7679 2.24164
R26500 DVDD.n9558 DVDD.n9261 2.24164
R26501 DVDD.n9536 DVDD.n7679 2.24164
R26502 DVDD.n9558 DVDD.n9260 2.24164
R26503 DVDD.n9531 DVDD.n7679 2.24164
R26504 DVDD.n9558 DVDD.n9259 2.24164
R26505 DVDD.n9524 DVDD.n7679 2.24164
R26506 DVDD.n9558 DVDD.n9258 2.24164
R26507 DVDD.n9519 DVDD.n7679 2.24164
R26508 DVDD.n9558 DVDD.n9257 2.24164
R26509 DVDD.n9512 DVDD.n7679 2.24164
R26510 DVDD.n9558 DVDD.n9256 2.24164
R26511 DVDD.n9507 DVDD.n7679 2.24164
R26512 DVDD.n9558 DVDD.n9255 2.24164
R26513 DVDD.n9500 DVDD.n7679 2.24164
R26514 DVDD.n9558 DVDD.n9254 2.24164
R26515 DVDD.n9495 DVDD.n7679 2.24164
R26516 DVDD.n9558 DVDD.n9253 2.24164
R26517 DVDD.n9488 DVDD.n7679 2.24164
R26518 DVDD.n9558 DVDD.n9252 2.24164
R26519 DVDD.n9483 DVDD.n7679 2.24164
R26520 DVDD.n9558 DVDD.n9251 2.24164
R26521 DVDD.n9476 DVDD.n7679 2.24164
R26522 DVDD.n9558 DVDD.n9250 2.24164
R26523 DVDD.n9471 DVDD.n7679 2.24164
R26524 DVDD.n9558 DVDD.n9249 2.24164
R26525 DVDD.n9464 DVDD.n7679 2.24164
R26526 DVDD.n9558 DVDD.n9248 2.24164
R26527 DVDD.n9459 DVDD.n7679 2.24164
R26528 DVDD.n9558 DVDD.n9247 2.24164
R26529 DVDD.n9452 DVDD.n7679 2.24164
R26530 DVDD.n9558 DVDD.n9246 2.24164
R26531 DVDD.n9447 DVDD.n7679 2.24164
R26532 DVDD.n9558 DVDD.n9245 2.24164
R26533 DVDD.n9440 DVDD.n7679 2.24164
R26534 DVDD.n9558 DVDD.n9244 2.24164
R26535 DVDD.n9435 DVDD.n7679 2.24164
R26536 DVDD.n9558 DVDD.n9243 2.24164
R26537 DVDD.n9428 DVDD.n7679 2.24164
R26538 DVDD.n9558 DVDD.n9242 2.24164
R26539 DVDD.n9423 DVDD.n7679 2.24164
R26540 DVDD.n9558 DVDD.n9241 2.24164
R26541 DVDD.n9416 DVDD.n7679 2.24164
R26542 DVDD.n9558 DVDD.n9240 2.24164
R26543 DVDD.n9411 DVDD.n7679 2.24164
R26544 DVDD.n9558 DVDD.n9239 2.24164
R26545 DVDD.n9404 DVDD.n7679 2.24164
R26546 DVDD.n9558 DVDD.n9238 2.24164
R26547 DVDD.n9399 DVDD.n7679 2.24164
R26548 DVDD.n9558 DVDD.n9237 2.24164
R26549 DVDD.n9392 DVDD.n7679 2.24164
R26550 DVDD.n9558 DVDD.n9236 2.24164
R26551 DVDD.n9387 DVDD.n7679 2.24164
R26552 DVDD.n9558 DVDD.n9235 2.24164
R26553 DVDD.n9380 DVDD.n7679 2.24164
R26554 DVDD.n9558 DVDD.n9234 2.24164
R26555 DVDD.n9375 DVDD.n7679 2.24164
R26556 DVDD.n9558 DVDD.n9233 2.24164
R26557 DVDD.n9368 DVDD.n7679 2.24164
R26558 DVDD.n9558 DVDD.n9232 2.24164
R26559 DVDD.n9363 DVDD.n7679 2.24164
R26560 DVDD.n9558 DVDD.n9231 2.24164
R26561 DVDD.n9356 DVDD.n7679 2.24164
R26562 DVDD.n9558 DVDD.n9230 2.24164
R26563 DVDD.n9351 DVDD.n7679 2.24164
R26564 DVDD.n9558 DVDD.n9229 2.24164
R26565 DVDD.n9344 DVDD.n7679 2.24164
R26566 DVDD.n9558 DVDD.n9228 2.24164
R26567 DVDD.n9339 DVDD.n7679 2.24164
R26568 DVDD.n9558 DVDD.n9227 2.24164
R26569 DVDD.n9332 DVDD.n7679 2.24164
R26570 DVDD.n9558 DVDD.n9226 2.24164
R26571 DVDD.n9327 DVDD.n7679 2.24164
R26572 DVDD.n9558 DVDD.n9225 2.24164
R26573 DVDD.n9320 DVDD.n7679 2.24164
R26574 DVDD.n9558 DVDD.n9224 2.24164
R26575 DVDD.n9315 DVDD.n7679 2.24164
R26576 DVDD.n9558 DVDD.n9223 2.24164
R26577 DVDD.n14863 DVDD.n14862 2.24164
R26578 DVDD.n14860 DVDD.n7656 2.24164
R26579 DVDD.n14863 DVDD.n7610 2.24164
R26580 DVDD.n14860 DVDD.n7655 2.24164
R26581 DVDD.n14863 DVDD.n7609 2.24164
R26582 DVDD.n14860 DVDD.n7654 2.24164
R26583 DVDD.n14863 DVDD.n7608 2.24164
R26584 DVDD.n14860 DVDD.n7653 2.24164
R26585 DVDD.n14863 DVDD.n7607 2.24164
R26586 DVDD.n14860 DVDD.n7652 2.24164
R26587 DVDD.n14863 DVDD.n7606 2.24164
R26588 DVDD.n14860 DVDD.n7651 2.24164
R26589 DVDD.n14863 DVDD.n7605 2.24164
R26590 DVDD.n14860 DVDD.n7650 2.24164
R26591 DVDD.n14863 DVDD.n7604 2.24164
R26592 DVDD.n14860 DVDD.n7649 2.24164
R26593 DVDD.n14863 DVDD.n7603 2.24164
R26594 DVDD.n14860 DVDD.n7648 2.24164
R26595 DVDD.n14863 DVDD.n7602 2.24164
R26596 DVDD.n14860 DVDD.n7647 2.24164
R26597 DVDD.n14863 DVDD.n7601 2.24164
R26598 DVDD.n14860 DVDD.n7646 2.24164
R26599 DVDD.n14863 DVDD.n7600 2.24164
R26600 DVDD.n14860 DVDD.n7645 2.24164
R26601 DVDD.n14863 DVDD.n7599 2.24164
R26602 DVDD.n14860 DVDD.n7644 2.24164
R26603 DVDD.n14863 DVDD.n7598 2.24164
R26604 DVDD.n14860 DVDD.n7643 2.24164
R26605 DVDD.n14863 DVDD.n7597 2.24164
R26606 DVDD.n14860 DVDD.n7642 2.24164
R26607 DVDD.n14863 DVDD.n7596 2.24164
R26608 DVDD.n14860 DVDD.n7641 2.24164
R26609 DVDD.n14863 DVDD.n7595 2.24164
R26610 DVDD.n14860 DVDD.n7640 2.24164
R26611 DVDD.n14863 DVDD.n7594 2.24164
R26612 DVDD.n14860 DVDD.n7639 2.24164
R26613 DVDD.n14863 DVDD.n7593 2.24164
R26614 DVDD.n14860 DVDD.n7638 2.24164
R26615 DVDD.n14863 DVDD.n7592 2.24164
R26616 DVDD.n14860 DVDD.n7637 2.24164
R26617 DVDD.n14863 DVDD.n7591 2.24164
R26618 DVDD.n14860 DVDD.n7636 2.24164
R26619 DVDD.n14863 DVDD.n7590 2.24164
R26620 DVDD.n14860 DVDD.n7635 2.24164
R26621 DVDD.n14863 DVDD.n7589 2.24164
R26622 DVDD.n14860 DVDD.n7634 2.24164
R26623 DVDD.n14863 DVDD.n7588 2.24164
R26624 DVDD.n14860 DVDD.n7633 2.24164
R26625 DVDD.n14863 DVDD.n7587 2.24164
R26626 DVDD.n14860 DVDD.n7632 2.24164
R26627 DVDD.n14863 DVDD.n7586 2.24164
R26628 DVDD.n14860 DVDD.n7631 2.24164
R26629 DVDD.n14863 DVDD.n7585 2.24164
R26630 DVDD.n14860 DVDD.n7630 2.24164
R26631 DVDD.n14863 DVDD.n7584 2.24164
R26632 DVDD.n14860 DVDD.n7629 2.24164
R26633 DVDD.n14863 DVDD.n7583 2.24164
R26634 DVDD.n14860 DVDD.n7628 2.24164
R26635 DVDD.n14863 DVDD.n7582 2.24164
R26636 DVDD.n14860 DVDD.n7627 2.24164
R26637 DVDD.n14863 DVDD.n7581 2.24164
R26638 DVDD.n14860 DVDD.n7626 2.24164
R26639 DVDD.n14863 DVDD.n7580 2.24164
R26640 DVDD.n14860 DVDD.n7625 2.24164
R26641 DVDD.n14863 DVDD.n7579 2.24164
R26642 DVDD.n14860 DVDD.n7624 2.24164
R26643 DVDD.n14863 DVDD.n7578 2.24164
R26644 DVDD.n14860 DVDD.n7623 2.24164
R26645 DVDD.n14863 DVDD.n7577 2.24164
R26646 DVDD.n14860 DVDD.n7622 2.24164
R26647 DVDD.n14863 DVDD.n7576 2.24164
R26648 DVDD.n14860 DVDD.n7621 2.24164
R26649 DVDD.n14863 DVDD.n7575 2.24164
R26650 DVDD.n14860 DVDD.n7620 2.24164
R26651 DVDD.n14863 DVDD.n7574 2.24164
R26652 DVDD.n14860 DVDD.n7619 2.24164
R26653 DVDD.n14863 DVDD.n7573 2.24164
R26654 DVDD.n14860 DVDD.n7618 2.24164
R26655 DVDD.n14863 DVDD.n7572 2.24164
R26656 DVDD.n14860 DVDD.n7617 2.24164
R26657 DVDD.n14863 DVDD.n7571 2.24164
R26658 DVDD.n14860 DVDD.n7616 2.24164
R26659 DVDD.n14863 DVDD.n7570 2.24164
R26660 DVDD.n15060 DVDD.n15059 2.24164
R26661 DVDD.n15057 DVDD.n7499 2.24164
R26662 DVDD.n15060 DVDD.n7453 2.24164
R26663 DVDD.n15057 DVDD.n7498 2.24164
R26664 DVDD.n15060 DVDD.n7452 2.24164
R26665 DVDD.n15057 DVDD.n7497 2.24164
R26666 DVDD.n15060 DVDD.n7451 2.24164
R26667 DVDD.n15057 DVDD.n7496 2.24164
R26668 DVDD.n15060 DVDD.n7450 2.24164
R26669 DVDD.n15057 DVDD.n7495 2.24164
R26670 DVDD.n15060 DVDD.n7449 2.24164
R26671 DVDD.n15057 DVDD.n7494 2.24164
R26672 DVDD.n15060 DVDD.n7448 2.24164
R26673 DVDD.n15057 DVDD.n7493 2.24164
R26674 DVDD.n15060 DVDD.n7447 2.24164
R26675 DVDD.n15057 DVDD.n7492 2.24164
R26676 DVDD.n15060 DVDD.n7446 2.24164
R26677 DVDD.n15057 DVDD.n7491 2.24164
R26678 DVDD.n15060 DVDD.n7445 2.24164
R26679 DVDD.n15057 DVDD.n7490 2.24164
R26680 DVDD.n15060 DVDD.n7444 2.24164
R26681 DVDD.n15057 DVDD.n7489 2.24164
R26682 DVDD.n15060 DVDD.n7443 2.24164
R26683 DVDD.n15057 DVDD.n7488 2.24164
R26684 DVDD.n15060 DVDD.n7442 2.24164
R26685 DVDD.n15057 DVDD.n7487 2.24164
R26686 DVDD.n15060 DVDD.n7441 2.24164
R26687 DVDD.n15057 DVDD.n7486 2.24164
R26688 DVDD.n15060 DVDD.n7440 2.24164
R26689 DVDD.n15057 DVDD.n7485 2.24164
R26690 DVDD.n15060 DVDD.n7439 2.24164
R26691 DVDD.n15057 DVDD.n7484 2.24164
R26692 DVDD.n15060 DVDD.n7438 2.24164
R26693 DVDD.n15057 DVDD.n7483 2.24164
R26694 DVDD.n15060 DVDD.n7437 2.24164
R26695 DVDD.n15057 DVDD.n7482 2.24164
R26696 DVDD.n15060 DVDD.n7436 2.24164
R26697 DVDD.n15057 DVDD.n7481 2.24164
R26698 DVDD.n15060 DVDD.n7435 2.24164
R26699 DVDD.n15057 DVDD.n7480 2.24164
R26700 DVDD.n15060 DVDD.n7434 2.24164
R26701 DVDD.n15057 DVDD.n7479 2.24164
R26702 DVDD.n15060 DVDD.n7433 2.24164
R26703 DVDD.n15057 DVDD.n7478 2.24164
R26704 DVDD.n15060 DVDD.n7432 2.24164
R26705 DVDD.n15057 DVDD.n7477 2.24164
R26706 DVDD.n15060 DVDD.n7431 2.24164
R26707 DVDD.n15057 DVDD.n7476 2.24164
R26708 DVDD.n15060 DVDD.n7430 2.24164
R26709 DVDD.n15057 DVDD.n7475 2.24164
R26710 DVDD.n15060 DVDD.n7429 2.24164
R26711 DVDD.n15057 DVDD.n7474 2.24164
R26712 DVDD.n15060 DVDD.n7428 2.24164
R26713 DVDD.n15057 DVDD.n7473 2.24164
R26714 DVDD.n15060 DVDD.n7427 2.24164
R26715 DVDD.n15057 DVDD.n7472 2.24164
R26716 DVDD.n15060 DVDD.n7426 2.24164
R26717 DVDD.n15057 DVDD.n7471 2.24164
R26718 DVDD.n15060 DVDD.n7425 2.24164
R26719 DVDD.n15057 DVDD.n7470 2.24164
R26720 DVDD.n15060 DVDD.n7424 2.24164
R26721 DVDD.n15057 DVDD.n7469 2.24164
R26722 DVDD.n15060 DVDD.n7423 2.24164
R26723 DVDD.n15057 DVDD.n7468 2.24164
R26724 DVDD.n15060 DVDD.n7422 2.24164
R26725 DVDD.n15057 DVDD.n7467 2.24164
R26726 DVDD.n15060 DVDD.n7421 2.24164
R26727 DVDD.n15057 DVDD.n7466 2.24164
R26728 DVDD.n15060 DVDD.n7420 2.24164
R26729 DVDD.n15057 DVDD.n7465 2.24164
R26730 DVDD.n15060 DVDD.n7419 2.24164
R26731 DVDD.n15057 DVDD.n7464 2.24164
R26732 DVDD.n15060 DVDD.n7418 2.24164
R26733 DVDD.n15057 DVDD.n7463 2.24164
R26734 DVDD.n15060 DVDD.n7417 2.24164
R26735 DVDD.n15057 DVDD.n7462 2.24164
R26736 DVDD.n15060 DVDD.n7416 2.24164
R26737 DVDD.n15057 DVDD.n7461 2.24164
R26738 DVDD.n15060 DVDD.n7415 2.24164
R26739 DVDD.n15057 DVDD.n7460 2.24164
R26740 DVDD.n15060 DVDD.n7414 2.24164
R26741 DVDD.n15057 DVDD.n7459 2.24164
R26742 DVDD.n15060 DVDD.n7413 2.24164
R26743 DVDD.n7154 DVDD.n7057 2.24164
R26744 DVDD.n7404 DVDD.n7110 2.24164
R26745 DVDD.n7161 DVDD.n7057 2.24164
R26746 DVDD.n7404 DVDD.n7109 2.24164
R26747 DVDD.n7165 DVDD.n7057 2.24164
R26748 DVDD.n7404 DVDD.n7108 2.24164
R26749 DVDD.n7173 DVDD.n7057 2.24164
R26750 DVDD.n7404 DVDD.n7107 2.24164
R26751 DVDD.n7177 DVDD.n7057 2.24164
R26752 DVDD.n7404 DVDD.n7106 2.24164
R26753 DVDD.n7185 DVDD.n7057 2.24164
R26754 DVDD.n7404 DVDD.n7105 2.24164
R26755 DVDD.n7189 DVDD.n7057 2.24164
R26756 DVDD.n7404 DVDD.n7104 2.24164
R26757 DVDD.n7197 DVDD.n7057 2.24164
R26758 DVDD.n7404 DVDD.n7103 2.24164
R26759 DVDD.n7201 DVDD.n7057 2.24164
R26760 DVDD.n7404 DVDD.n7102 2.24164
R26761 DVDD.n7209 DVDD.n7057 2.24164
R26762 DVDD.n7404 DVDD.n7101 2.24164
R26763 DVDD.n7213 DVDD.n7057 2.24164
R26764 DVDD.n7404 DVDD.n7100 2.24164
R26765 DVDD.n7221 DVDD.n7057 2.24164
R26766 DVDD.n7404 DVDD.n7099 2.24164
R26767 DVDD.n7225 DVDD.n7057 2.24164
R26768 DVDD.n7404 DVDD.n7098 2.24164
R26769 DVDD.n7233 DVDD.n7057 2.24164
R26770 DVDD.n7404 DVDD.n7097 2.24164
R26771 DVDD.n7237 DVDD.n7057 2.24164
R26772 DVDD.n7404 DVDD.n7096 2.24164
R26773 DVDD.n7245 DVDD.n7057 2.24164
R26774 DVDD.n7404 DVDD.n7095 2.24164
R26775 DVDD.n7249 DVDD.n7057 2.24164
R26776 DVDD.n7404 DVDD.n7094 2.24164
R26777 DVDD.n7257 DVDD.n7057 2.24164
R26778 DVDD.n7404 DVDD.n7093 2.24164
R26779 DVDD.n7261 DVDD.n7057 2.24164
R26780 DVDD.n7404 DVDD.n7092 2.24164
R26781 DVDD.n7269 DVDD.n7057 2.24164
R26782 DVDD.n7404 DVDD.n7091 2.24164
R26783 DVDD.n7273 DVDD.n7057 2.24164
R26784 DVDD.n7404 DVDD.n7090 2.24164
R26785 DVDD.n7281 DVDD.n7057 2.24164
R26786 DVDD.n7404 DVDD.n7089 2.24164
R26787 DVDD.n7285 DVDD.n7057 2.24164
R26788 DVDD.n7404 DVDD.n7088 2.24164
R26789 DVDD.n7293 DVDD.n7057 2.24164
R26790 DVDD.n7404 DVDD.n7087 2.24164
R26791 DVDD.n7297 DVDD.n7057 2.24164
R26792 DVDD.n7404 DVDD.n7086 2.24164
R26793 DVDD.n7305 DVDD.n7057 2.24164
R26794 DVDD.n7404 DVDD.n7085 2.24164
R26795 DVDD.n7309 DVDD.n7057 2.24164
R26796 DVDD.n7404 DVDD.n7084 2.24164
R26797 DVDD.n7317 DVDD.n7057 2.24164
R26798 DVDD.n7404 DVDD.n7083 2.24164
R26799 DVDD.n7321 DVDD.n7057 2.24164
R26800 DVDD.n7404 DVDD.n7082 2.24164
R26801 DVDD.n7329 DVDD.n7057 2.24164
R26802 DVDD.n7404 DVDD.n7081 2.24164
R26803 DVDD.n7333 DVDD.n7057 2.24164
R26804 DVDD.n7404 DVDD.n7080 2.24164
R26805 DVDD.n7341 DVDD.n7057 2.24164
R26806 DVDD.n7404 DVDD.n7079 2.24164
R26807 DVDD.n7345 DVDD.n7057 2.24164
R26808 DVDD.n7404 DVDD.n7078 2.24164
R26809 DVDD.n7353 DVDD.n7057 2.24164
R26810 DVDD.n7404 DVDD.n7077 2.24164
R26811 DVDD.n7357 DVDD.n7057 2.24164
R26812 DVDD.n7404 DVDD.n7076 2.24164
R26813 DVDD.n7365 DVDD.n7057 2.24164
R26814 DVDD.n7404 DVDD.n7075 2.24164
R26815 DVDD.n7369 DVDD.n7057 2.24164
R26816 DVDD.n7404 DVDD.n7074 2.24164
R26817 DVDD.n7377 DVDD.n7057 2.24164
R26818 DVDD.n7404 DVDD.n7073 2.24164
R26819 DVDD.n7381 DVDD.n7057 2.24164
R26820 DVDD.n7404 DVDD.n7072 2.24164
R26821 DVDD.n7389 DVDD.n7057 2.24164
R26822 DVDD.n7404 DVDD.n7071 2.24164
R26823 DVDD.n7393 DVDD.n7057 2.24164
R26824 DVDD.n7404 DVDD.n7070 2.24164
R26825 DVDD.n7402 DVDD.n7057 2.24164
R26826 DVDD.n15092 DVDD.n15091 2.24164
R26827 DVDD.n15089 DVDD.n6793 2.24164
R26828 DVDD.n15092 DVDD.n6748 2.24164
R26829 DVDD.n15089 DVDD.n6792 2.24164
R26830 DVDD.n15092 DVDD.n6747 2.24164
R26831 DVDD.n15089 DVDD.n6791 2.24164
R26832 DVDD.n15092 DVDD.n6746 2.24164
R26833 DVDD.n15089 DVDD.n6790 2.24164
R26834 DVDD.n15092 DVDD.n6745 2.24164
R26835 DVDD.n15089 DVDD.n6789 2.24164
R26836 DVDD.n15092 DVDD.n6744 2.24164
R26837 DVDD.n15089 DVDD.n6788 2.24164
R26838 DVDD.n15092 DVDD.n6743 2.24164
R26839 DVDD.n15089 DVDD.n6787 2.24164
R26840 DVDD.n15092 DVDD.n6742 2.24164
R26841 DVDD.n15089 DVDD.n6786 2.24164
R26842 DVDD.n15092 DVDD.n6741 2.24164
R26843 DVDD.n15089 DVDD.n6785 2.24164
R26844 DVDD.n15092 DVDD.n6740 2.24164
R26845 DVDD.n15089 DVDD.n6784 2.24164
R26846 DVDD.n15092 DVDD.n6739 2.24164
R26847 DVDD.n15089 DVDD.n6783 2.24164
R26848 DVDD.n15092 DVDD.n6738 2.24164
R26849 DVDD.n15089 DVDD.n6782 2.24164
R26850 DVDD.n15092 DVDD.n6737 2.24164
R26851 DVDD.n15089 DVDD.n6781 2.24164
R26852 DVDD.n15092 DVDD.n6736 2.24164
R26853 DVDD.n15089 DVDD.n6780 2.24164
R26854 DVDD.n15092 DVDD.n6735 2.24164
R26855 DVDD.n15089 DVDD.n6779 2.24164
R26856 DVDD.n15092 DVDD.n6734 2.24164
R26857 DVDD.n15089 DVDD.n6778 2.24164
R26858 DVDD.n15092 DVDD.n6733 2.24164
R26859 DVDD.n15089 DVDD.n6777 2.24164
R26860 DVDD.n15092 DVDD.n6732 2.24164
R26861 DVDD.n15089 DVDD.n6776 2.24164
R26862 DVDD.n15092 DVDD.n6731 2.24164
R26863 DVDD.n15089 DVDD.n6775 2.24164
R26864 DVDD.n15092 DVDD.n6730 2.24164
R26865 DVDD.n15089 DVDD.n6774 2.24164
R26866 DVDD.n15092 DVDD.n6729 2.24164
R26867 DVDD.n15089 DVDD.n6773 2.24164
R26868 DVDD.n15092 DVDD.n6728 2.24164
R26869 DVDD.n15089 DVDD.n6772 2.24164
R26870 DVDD.n15092 DVDD.n6727 2.24164
R26871 DVDD.n15089 DVDD.n6771 2.24164
R26872 DVDD.n15092 DVDD.n6726 2.24164
R26873 DVDD.n15089 DVDD.n6770 2.24164
R26874 DVDD.n15092 DVDD.n6725 2.24164
R26875 DVDD.n15089 DVDD.n6769 2.24164
R26876 DVDD.n15092 DVDD.n6724 2.24164
R26877 DVDD.n15089 DVDD.n6768 2.24164
R26878 DVDD.n15092 DVDD.n6723 2.24164
R26879 DVDD.n15089 DVDD.n6767 2.24164
R26880 DVDD.n15092 DVDD.n6722 2.24164
R26881 DVDD.n15089 DVDD.n6766 2.24164
R26882 DVDD.n15092 DVDD.n6721 2.24164
R26883 DVDD.n15089 DVDD.n6765 2.24164
R26884 DVDD.n15092 DVDD.n6720 2.24164
R26885 DVDD.n15089 DVDD.n6764 2.24164
R26886 DVDD.n15092 DVDD.n6719 2.24164
R26887 DVDD.n15089 DVDD.n6763 2.24164
R26888 DVDD.n15092 DVDD.n6718 2.24164
R26889 DVDD.n15089 DVDD.n6762 2.24164
R26890 DVDD.n15092 DVDD.n6717 2.24164
R26891 DVDD.n15089 DVDD.n6761 2.24164
R26892 DVDD.n15092 DVDD.n6716 2.24164
R26893 DVDD.n15089 DVDD.n6760 2.24164
R26894 DVDD.n15092 DVDD.n6715 2.24164
R26895 DVDD.n15089 DVDD.n6759 2.24164
R26896 DVDD.n15092 DVDD.n6714 2.24164
R26897 DVDD.n15089 DVDD.n6758 2.24164
R26898 DVDD.n15092 DVDD.n6713 2.24164
R26899 DVDD.n15089 DVDD.n6757 2.24164
R26900 DVDD.n15092 DVDD.n6712 2.24164
R26901 DVDD.n15089 DVDD.n6756 2.24164
R26902 DVDD.n15092 DVDD.n6711 2.24164
R26903 DVDD.n15089 DVDD.n6755 2.24164
R26904 DVDD.n15092 DVDD.n6710 2.24164
R26905 DVDD.n15089 DVDD.n6754 2.24164
R26906 DVDD.n15092 DVDD.n6709 2.24164
R26907 DVDD.n15089 DVDD.n6753 2.24164
R26908 DVDD.n15092 DVDD.n6708 2.24164
R26909 DVDD.n15101 DVDD.n6390 2.24164
R26910 DVDD.n6696 DVDD.n6405 2.24164
R26911 DVDD.n15101 DVDD.n6389 2.24164
R26912 DVDD.n6696 DVDD.n6406 2.24164
R26913 DVDD.n15101 DVDD.n6388 2.24164
R26914 DVDD.n6696 DVDD.n6407 2.24164
R26915 DVDD.n15101 DVDD.n6387 2.24164
R26916 DVDD.n6696 DVDD.n6408 2.24164
R26917 DVDD.n15101 DVDD.n6386 2.24164
R26918 DVDD.n6696 DVDD.n6409 2.24164
R26919 DVDD.n15101 DVDD.n6385 2.24164
R26920 DVDD.n6696 DVDD.n6410 2.24164
R26921 DVDD.n15101 DVDD.n6384 2.24164
R26922 DVDD.n6696 DVDD.n6411 2.24164
R26923 DVDD.n15101 DVDD.n6383 2.24164
R26924 DVDD.n6696 DVDD.n6412 2.24164
R26925 DVDD.n15101 DVDD.n6382 2.24164
R26926 DVDD.n6696 DVDD.n6413 2.24164
R26927 DVDD.n15101 DVDD.n6381 2.24164
R26928 DVDD.n6696 DVDD.n6414 2.24164
R26929 DVDD.n15101 DVDD.n6380 2.24164
R26930 DVDD.n6696 DVDD.n6415 2.24164
R26931 DVDD.n15101 DVDD.n6379 2.24164
R26932 DVDD.n6696 DVDD.n6416 2.24164
R26933 DVDD.n15101 DVDD.n6378 2.24164
R26934 DVDD.n6696 DVDD.n6417 2.24164
R26935 DVDD.n15101 DVDD.n6377 2.24164
R26936 DVDD.n6696 DVDD.n6418 2.24164
R26937 DVDD.n15101 DVDD.n6376 2.24164
R26938 DVDD.n6696 DVDD.n6419 2.24164
R26939 DVDD.n15101 DVDD.n6375 2.24164
R26940 DVDD.n6696 DVDD.n6420 2.24164
R26941 DVDD.n15101 DVDD.n6374 2.24164
R26942 DVDD.n6696 DVDD.n6421 2.24164
R26943 DVDD.n15101 DVDD.n6373 2.24164
R26944 DVDD.n6696 DVDD.n6422 2.24164
R26945 DVDD.n15101 DVDD.n6372 2.24164
R26946 DVDD.n6696 DVDD.n6423 2.24164
R26947 DVDD.n15101 DVDD.n6371 2.24164
R26948 DVDD.n6696 DVDD.n6424 2.24164
R26949 DVDD.n15101 DVDD.n6370 2.24164
R26950 DVDD.n6696 DVDD.n6425 2.24164
R26951 DVDD.n15101 DVDD.n6369 2.24164
R26952 DVDD.n6696 DVDD.n6426 2.24164
R26953 DVDD.n15101 DVDD.n6368 2.24164
R26954 DVDD.n6696 DVDD.n6427 2.24164
R26955 DVDD.n15101 DVDD.n6367 2.24164
R26956 DVDD.n6696 DVDD.n6428 2.24164
R26957 DVDD.n15101 DVDD.n6366 2.24164
R26958 DVDD.n6696 DVDD.n6429 2.24164
R26959 DVDD.n15101 DVDD.n6365 2.24164
R26960 DVDD.n6696 DVDD.n6430 2.24164
R26961 DVDD.n15101 DVDD.n6364 2.24164
R26962 DVDD.n6696 DVDD.n6431 2.24164
R26963 DVDD.n15101 DVDD.n6363 2.24164
R26964 DVDD.n6696 DVDD.n6432 2.24164
R26965 DVDD.n15101 DVDD.n6362 2.24164
R26966 DVDD.n6696 DVDD.n6433 2.24164
R26967 DVDD.n15101 DVDD.n6361 2.24164
R26968 DVDD.n6696 DVDD.n6434 2.24164
R26969 DVDD.n15101 DVDD.n6360 2.24164
R26970 DVDD.n6696 DVDD.n6435 2.24164
R26971 DVDD.n15101 DVDD.n6359 2.24164
R26972 DVDD.n6696 DVDD.n6436 2.24164
R26973 DVDD.n15101 DVDD.n6358 2.24164
R26974 DVDD.n6696 DVDD.n6437 2.24164
R26975 DVDD.n15101 DVDD.n6357 2.24164
R26976 DVDD.n6696 DVDD.n6438 2.24164
R26977 DVDD.n15101 DVDD.n6356 2.24164
R26978 DVDD.n6696 DVDD.n6439 2.24164
R26979 DVDD.n15101 DVDD.n6355 2.24164
R26980 DVDD.n6696 DVDD.n6440 2.24164
R26981 DVDD.n15101 DVDD.n6354 2.24164
R26982 DVDD.n6696 DVDD.n6441 2.24164
R26983 DVDD.n15101 DVDD.n6353 2.24164
R26984 DVDD.n6696 DVDD.n6442 2.24164
R26985 DVDD.n15101 DVDD.n6352 2.24164
R26986 DVDD.n6696 DVDD.n6443 2.24164
R26987 DVDD.n15101 DVDD.n6351 2.24164
R26988 DVDD.n6696 DVDD.n6444 2.24164
R26989 DVDD.n15101 DVDD.n6350 2.24164
R26990 DVDD.n6696 DVDD.n6445 2.24164
R26991 DVDD.n15101 DVDD.n6349 2.24164
R26992 DVDD.n1256 DVDD.n1255 2.24164
R26993 DVDD.n964 DVDD.n915 2.24164
R26994 DVDD.n1256 DVDD.n962 2.24164
R26995 DVDD.n1247 DVDD.n915 2.24164
R26996 DVDD.n1256 DVDD.n961 2.24164
R26997 DVDD.n971 DVDD.n915 2.24164
R26998 DVDD.n1256 DVDD.n960 2.24164
R26999 DVDD.n1238 DVDD.n915 2.24164
R27000 DVDD.n1256 DVDD.n959 2.24164
R27001 DVDD.n976 DVDD.n915 2.24164
R27002 DVDD.n1256 DVDD.n958 2.24164
R27003 DVDD.n1229 DVDD.n915 2.24164
R27004 DVDD.n1256 DVDD.n957 2.24164
R27005 DVDD.n981 DVDD.n915 2.24164
R27006 DVDD.n1256 DVDD.n956 2.24164
R27007 DVDD.n1220 DVDD.n915 2.24164
R27008 DVDD.n1256 DVDD.n955 2.24164
R27009 DVDD.n986 DVDD.n915 2.24164
R27010 DVDD.n1256 DVDD.n954 2.24164
R27011 DVDD.n1211 DVDD.n915 2.24164
R27012 DVDD.n1256 DVDD.n953 2.24164
R27013 DVDD.n991 DVDD.n915 2.24164
R27014 DVDD.n1256 DVDD.n952 2.24164
R27015 DVDD.n1202 DVDD.n915 2.24164
R27016 DVDD.n1256 DVDD.n951 2.24164
R27017 DVDD.n996 DVDD.n915 2.24164
R27018 DVDD.n1256 DVDD.n950 2.24164
R27019 DVDD.n1193 DVDD.n915 2.24164
R27020 DVDD.n1256 DVDD.n949 2.24164
R27021 DVDD.n1001 DVDD.n915 2.24164
R27022 DVDD.n1256 DVDD.n948 2.24164
R27023 DVDD.n1184 DVDD.n915 2.24164
R27024 DVDD.n1256 DVDD.n947 2.24164
R27025 DVDD.n1006 DVDD.n915 2.24164
R27026 DVDD.n1256 DVDD.n946 2.24164
R27027 DVDD.n1175 DVDD.n915 2.24164
R27028 DVDD.n1256 DVDD.n945 2.24164
R27029 DVDD.n1011 DVDD.n915 2.24164
R27030 DVDD.n1256 DVDD.n944 2.24164
R27031 DVDD.n1166 DVDD.n915 2.24164
R27032 DVDD.n1256 DVDD.n943 2.24164
R27033 DVDD.n1016 DVDD.n915 2.24164
R27034 DVDD.n1256 DVDD.n942 2.24164
R27035 DVDD.n1157 DVDD.n915 2.24164
R27036 DVDD.n1256 DVDD.n941 2.24164
R27037 DVDD.n1021 DVDD.n915 2.24164
R27038 DVDD.n1256 DVDD.n940 2.24164
R27039 DVDD.n1148 DVDD.n915 2.24164
R27040 DVDD.n1256 DVDD.n939 2.24164
R27041 DVDD.n1026 DVDD.n915 2.24164
R27042 DVDD.n1256 DVDD.n938 2.24164
R27043 DVDD.n1139 DVDD.n915 2.24164
R27044 DVDD.n1256 DVDD.n937 2.24164
R27045 DVDD.n1031 DVDD.n915 2.24164
R27046 DVDD.n1256 DVDD.n936 2.24164
R27047 DVDD.n1130 DVDD.n915 2.24164
R27048 DVDD.n1256 DVDD.n935 2.24164
R27049 DVDD.n1036 DVDD.n915 2.24164
R27050 DVDD.n1256 DVDD.n934 2.24164
R27051 DVDD.n1121 DVDD.n915 2.24164
R27052 DVDD.n1256 DVDD.n933 2.24164
R27053 DVDD.n1041 DVDD.n915 2.24164
R27054 DVDD.n1256 DVDD.n932 2.24164
R27055 DVDD.n1112 DVDD.n915 2.24164
R27056 DVDD.n1256 DVDD.n931 2.24164
R27057 DVDD.n1046 DVDD.n915 2.24164
R27058 DVDD.n1256 DVDD.n930 2.24164
R27059 DVDD.n1103 DVDD.n915 2.24164
R27060 DVDD.n1256 DVDD.n929 2.24164
R27061 DVDD.n1051 DVDD.n915 2.24164
R27062 DVDD.n1256 DVDD.n928 2.24164
R27063 DVDD.n1094 DVDD.n915 2.24164
R27064 DVDD.n1256 DVDD.n927 2.24164
R27065 DVDD.n1056 DVDD.n915 2.24164
R27066 DVDD.n1256 DVDD.n926 2.24164
R27067 DVDD.n1085 DVDD.n915 2.24164
R27068 DVDD.n1256 DVDD.n925 2.24164
R27069 DVDD.n1061 DVDD.n915 2.24164
R27070 DVDD.n1256 DVDD.n924 2.24164
R27071 DVDD.n1076 DVDD.n915 2.24164
R27072 DVDD.n1256 DVDD.n923 2.24164
R27073 DVDD.n1066 DVDD.n915 2.24164
R27074 DVDD.n1256 DVDD.n922 2.24164
R27075 DVDD.n6331 DVDD.n6330 2.24164
R27076 DVDD.n15112 DVDD.n6041 2.24164
R27077 DVDD.n6331 DVDD.n6090 2.24164
R27078 DVDD.n15112 DVDD.n6040 2.24164
R27079 DVDD.n6331 DVDD.n6089 2.24164
R27080 DVDD.n15112 DVDD.n6039 2.24164
R27081 DVDD.n6331 DVDD.n6088 2.24164
R27082 DVDD.n15112 DVDD.n6038 2.24164
R27083 DVDD.n6331 DVDD.n6087 2.24164
R27084 DVDD.n15112 DVDD.n6037 2.24164
R27085 DVDD.n6331 DVDD.n6086 2.24164
R27086 DVDD.n15112 DVDD.n6036 2.24164
R27087 DVDD.n6331 DVDD.n6085 2.24164
R27088 DVDD.n15112 DVDD.n6035 2.24164
R27089 DVDD.n6331 DVDD.n6084 2.24164
R27090 DVDD.n15112 DVDD.n6034 2.24164
R27091 DVDD.n6331 DVDD.n6083 2.24164
R27092 DVDD.n15112 DVDD.n6033 2.24164
R27093 DVDD.n6331 DVDD.n6082 2.24164
R27094 DVDD.n15112 DVDD.n6032 2.24164
R27095 DVDD.n6331 DVDD.n6081 2.24164
R27096 DVDD.n15112 DVDD.n6031 2.24164
R27097 DVDD.n6331 DVDD.n6080 2.24164
R27098 DVDD.n15112 DVDD.n6030 2.24164
R27099 DVDD.n6331 DVDD.n6079 2.24164
R27100 DVDD.n15112 DVDD.n6029 2.24164
R27101 DVDD.n6331 DVDD.n6078 2.24164
R27102 DVDD.n15112 DVDD.n6028 2.24164
R27103 DVDD.n6331 DVDD.n6077 2.24164
R27104 DVDD.n15112 DVDD.n6027 2.24164
R27105 DVDD.n6331 DVDD.n6076 2.24164
R27106 DVDD.n15112 DVDD.n6026 2.24164
R27107 DVDD.n6331 DVDD.n6075 2.24164
R27108 DVDD.n15112 DVDD.n6025 2.24164
R27109 DVDD.n6331 DVDD.n6074 2.24164
R27110 DVDD.n15112 DVDD.n6024 2.24164
R27111 DVDD.n6331 DVDD.n6073 2.24164
R27112 DVDD.n15112 DVDD.n6023 2.24164
R27113 DVDD.n6331 DVDD.n6072 2.24164
R27114 DVDD.n15112 DVDD.n6022 2.24164
R27115 DVDD.n6331 DVDD.n6071 2.24164
R27116 DVDD.n15112 DVDD.n6021 2.24164
R27117 DVDD.n6331 DVDD.n6070 2.24164
R27118 DVDD.n15112 DVDD.n6020 2.24164
R27119 DVDD.n6331 DVDD.n6069 2.24164
R27120 DVDD.n15112 DVDD.n6019 2.24164
R27121 DVDD.n6331 DVDD.n6068 2.24164
R27122 DVDD.n15112 DVDD.n6018 2.24164
R27123 DVDD.n6331 DVDD.n6067 2.24164
R27124 DVDD.n15112 DVDD.n6017 2.24164
R27125 DVDD.n6331 DVDD.n6066 2.24164
R27126 DVDD.n15112 DVDD.n6016 2.24164
R27127 DVDD.n6331 DVDD.n6065 2.24164
R27128 DVDD.n15112 DVDD.n6015 2.24164
R27129 DVDD.n6331 DVDD.n6064 2.24164
R27130 DVDD.n15112 DVDD.n6014 2.24164
R27131 DVDD.n6331 DVDD.n6063 2.24164
R27132 DVDD.n15112 DVDD.n6013 2.24164
R27133 DVDD.n6331 DVDD.n6062 2.24164
R27134 DVDD.n15112 DVDD.n6012 2.24164
R27135 DVDD.n6331 DVDD.n6061 2.24164
R27136 DVDD.n15112 DVDD.n6011 2.24164
R27137 DVDD.n6331 DVDD.n6060 2.24164
R27138 DVDD.n15112 DVDD.n6010 2.24164
R27139 DVDD.n6331 DVDD.n6059 2.24164
R27140 DVDD.n15112 DVDD.n6009 2.24164
R27141 DVDD.n6331 DVDD.n6058 2.24164
R27142 DVDD.n15112 DVDD.n6008 2.24164
R27143 DVDD.n6331 DVDD.n6057 2.24164
R27144 DVDD.n15112 DVDD.n6007 2.24164
R27145 DVDD.n6331 DVDD.n6056 2.24164
R27146 DVDD.n15112 DVDD.n6006 2.24164
R27147 DVDD.n6331 DVDD.n6055 2.24164
R27148 DVDD.n15112 DVDD.n6005 2.24164
R27149 DVDD.n6331 DVDD.n6054 2.24164
R27150 DVDD.n15112 DVDD.n6004 2.24164
R27151 DVDD.n6331 DVDD.n6053 2.24164
R27152 DVDD.n15112 DVDD.n6003 2.24164
R27153 DVDD.n6331 DVDD.n6052 2.24164
R27154 DVDD.n15112 DVDD.n6002 2.24164
R27155 DVDD.n6332 DVDD.n6331 2.24164
R27156 DVDD.n15112 DVDD.n6001 2.24164
R27157 DVDD.n6331 DVDD.n6045 2.24164
R27158 DVDD.n18785 DVDD.n18770 2.23714
R27159 DVDD.n18783 DVDD.n18770 2.23714
R27160 DVDD.n18781 DVDD.n18770 2.23714
R27161 DVDD.n18779 DVDD.n18770 2.23714
R27162 DVDD.n18777 DVDD.n18770 2.23714
R27163 DVDD.n18775 DVDD.n18770 2.23714
R27164 DVDD.n21052 DVDD.n18786 2.23714
R27165 DVDD.n21052 DVDD.n18784 2.23714
R27166 DVDD.n21052 DVDD.n18782 2.23714
R27167 DVDD.n21052 DVDD.n18780 2.23714
R27168 DVDD.n21052 DVDD.n18778 2.23714
R27169 DVDD.n21052 DVDD.n18776 2.23714
R27170 DVDD.n21052 DVDD.n18774 2.23714
R27171 DVDD.n19107 DVDD.n19094 2.23714
R27172 DVDD.n19109 DVDD.n19094 2.23714
R27173 DVDD.n19111 DVDD.n19094 2.23714
R27174 DVDD.n19113 DVDD.n19094 2.23714
R27175 DVDD.n19115 DVDD.n19094 2.23714
R27176 DVDD.n19117 DVDD.n19094 2.23714
R27177 DVDD.n19119 DVDD.n19094 2.23714
R27178 DVDD.n19106 DVDD.n19095 2.23714
R27179 DVDD.n19108 DVDD.n19095 2.23714
R27180 DVDD.n19110 DVDD.n19095 2.23714
R27181 DVDD.n19112 DVDD.n19095 2.23714
R27182 DVDD.n19114 DVDD.n19095 2.23714
R27183 DVDD.n19116 DVDD.n19095 2.23714
R27184 DVDD.n19118 DVDD.n19095 2.23714
R27185 DVDD.n19120 DVDD.n19095 2.23714
R27186 DVDD.n20935 DVDD.n18868 2.23714
R27187 DVDD.n20937 DVDD.n18868 2.23714
R27188 DVDD.n20939 DVDD.n18868 2.23714
R27189 DVDD.n20941 DVDD.n18868 2.23714
R27190 DVDD.n20943 DVDD.n18868 2.23714
R27191 DVDD.n20945 DVDD.n18868 2.23714
R27192 DVDD.n20947 DVDD.n18868 2.23714
R27193 DVDD.n20934 DVDD.n18869 2.23714
R27194 DVDD.n20936 DVDD.n18869 2.23714
R27195 DVDD.n20938 DVDD.n18869 2.23714
R27196 DVDD.n20940 DVDD.n18869 2.23714
R27197 DVDD.n20942 DVDD.n18869 2.23714
R27198 DVDD.n20944 DVDD.n18869 2.23714
R27199 DVDD.n20946 DVDD.n18869 2.23714
R27200 DVDD.n20948 DVDD.n18869 2.23714
R27201 DVDD.n20467 DVDD.n20465 2.23714
R27202 DVDD.n20469 DVDD.n20465 2.23714
R27203 DVDD.n20471 DVDD.n20465 2.23714
R27204 DVDD.n20473 DVDD.n20465 2.23714
R27205 DVDD.n20475 DVDD.n20465 2.23714
R27206 DVDD.n20477 DVDD.n20465 2.23714
R27207 DVDD.n20466 DVDD.n19033 2.23714
R27208 DVDD.n20468 DVDD.n19033 2.23714
R27209 DVDD.n20470 DVDD.n19033 2.23714
R27210 DVDD.n20472 DVDD.n19033 2.23714
R27211 DVDD.n20474 DVDD.n19033 2.23714
R27212 DVDD.n20476 DVDD.n19033 2.23714
R27213 DVDD.n20478 DVDD.n19033 2.23714
R27214 DVDD.n21055 DVDD.n18769 2.23714
R27215 DVDD.n21055 DVDD.n18768 2.23714
R27216 DVDD.n21055 DVDD.n18767 2.23714
R27217 DVDD.n21055 DVDD.n18766 2.23714
R27218 DVDD.n21055 DVDD.n18765 2.23714
R27219 DVDD.n21055 DVDD.n18764 2.23714
R27220 DVDD.n21059 DVDD.n18761 2.23714
R27221 DVDD.n21059 DVDD.n18760 2.23714
R27222 DVDD.n21059 DVDD.n18759 2.23714
R27223 DVDD.n21059 DVDD.n18758 2.23714
R27224 DVDD.n21059 DVDD.n18757 2.23714
R27225 DVDD.n21059 DVDD.n18756 2.23714
R27226 DVDD.n21059 DVDD.n18755 2.23714
R27227 DVDD.n19123 DVDD.n19092 2.23714
R27228 DVDD.n19123 DVDD.n19090 2.23714
R27229 DVDD.n19123 DVDD.n19088 2.23714
R27230 DVDD.n19123 DVDD.n19086 2.23714
R27231 DVDD.n19123 DVDD.n19084 2.23714
R27232 DVDD.n19123 DVDD.n19082 2.23714
R27233 DVDD.n19123 DVDD.n19080 2.23714
R27234 DVDD.n19093 DVDD.n18763 2.23714
R27235 DVDD.n19091 DVDD.n18763 2.23714
R27236 DVDD.n19089 DVDD.n18763 2.23714
R27237 DVDD.n19087 DVDD.n18763 2.23714
R27238 DVDD.n19085 DVDD.n18763 2.23714
R27239 DVDD.n19083 DVDD.n18763 2.23714
R27240 DVDD.n19081 DVDD.n18763 2.23714
R27241 DVDD.n19079 DVDD.n18763 2.23714
R27242 DVDD.n20952 DVDD.n18866 2.23714
R27243 DVDD.n20954 DVDD.n18866 2.23714
R27244 DVDD.n20956 DVDD.n18866 2.23714
R27245 DVDD.n20958 DVDD.n18866 2.23714
R27246 DVDD.n20960 DVDD.n18866 2.23714
R27247 DVDD.n20962 DVDD.n18866 2.23714
R27248 DVDD.n20964 DVDD.n18866 2.23714
R27249 DVDD.n20951 DVDD.n18867 2.23714
R27250 DVDD.n20953 DVDD.n18867 2.23714
R27251 DVDD.n20955 DVDD.n18867 2.23714
R27252 DVDD.n20957 DVDD.n18867 2.23714
R27253 DVDD.n20959 DVDD.n18867 2.23714
R27254 DVDD.n20961 DVDD.n18867 2.23714
R27255 DVDD.n20963 DVDD.n18867 2.23714
R27256 DVDD.n20965 DVDD.n18867 2.23714
R27257 DVDD.n20535 DVDD.n19808 2.23714
R27258 DVDD.n20535 DVDD.n19806 2.23714
R27259 DVDD.n20535 DVDD.n19804 2.23714
R27260 DVDD.n20535 DVDD.n19802 2.23714
R27261 DVDD.n20535 DVDD.n19800 2.23714
R27262 DVDD.n20535 DVDD.n19798 2.23714
R27263 DVDD.n19809 DVDD.n19129 2.23714
R27264 DVDD.n19807 DVDD.n19129 2.23714
R27265 DVDD.n19805 DVDD.n19129 2.23714
R27266 DVDD.n19803 DVDD.n19129 2.23714
R27267 DVDD.n19801 DVDD.n19129 2.23714
R27268 DVDD.n19799 DVDD.n19129 2.23714
R27269 DVDD.n20484 DVDD.n19129 2.23714
R27270 DVDD.n20978 DVDD.n20977 2.23714
R27271 DVDD.n20978 DVDD.n20976 2.23714
R27272 DVDD.n20978 DVDD.n20975 2.23714
R27273 DVDD.n20982 DVDD.n18828 2.23714
R27274 DVDD.n20982 DVDD.n18827 2.23714
R27275 DVDD.n20982 DVDD.n18826 2.23714
R27276 DVDD.n20982 DVDD.n18825 2.23714
R27277 DVDD.n20531 DVDD.n20523 2.23714
R27278 DVDD.n20531 DVDD.n20522 2.23714
R27279 DVDD.n20531 DVDD.n20521 2.23714
R27280 DVDD.n20529 DVDD.n20486 2.23714
R27281 DVDD.n20529 DVDD.n20528 2.23714
R27282 DVDD.n20529 DVDD.n20527 2.23714
R27283 DVDD.n20529 DVDD.n20526 2.23714
R27284 DVDD.n21504 DVDD.n21503 2.14713
R27285 DVDD.n21500 DVDD.n18560 1.99748
R27286 DVDD.n18615 DVDD.n18560 1.99748
R27287 DVDD.n21507 DVDD.n18560 1.99748
R27288 DVDD.n18612 DVDD.n18560 1.99748
R27289 DVDD.n21514 DVDD.n18560 1.99748
R27290 DVDD.n18609 DVDD.n18560 1.99748
R27291 DVDD.n21521 DVDD.n18560 1.99748
R27292 DVDD.n18606 DVDD.n18560 1.99748
R27293 DVDD.n21528 DVDD.n18560 1.99748
R27294 DVDD.n18603 DVDD.n18560 1.99748
R27295 DVDD.n21535 DVDD.n18560 1.99748
R27296 DVDD.n18600 DVDD.n18560 1.99748
R27297 DVDD.n21542 DVDD.n18560 1.99748
R27298 DVDD.n18596 DVDD.n18560 1.99748
R27299 DVDD.n21549 DVDD.n18560 1.99748
R27300 DVDD.n18593 DVDD.n18560 1.99748
R27301 DVDD.n21556 DVDD.n18560 1.99748
R27302 DVDD.n18590 DVDD.n18560 1.99748
R27303 DVDD.n21563 DVDD.n18560 1.99748
R27304 DVDD.n18587 DVDD.n18560 1.99748
R27305 DVDD.n21570 DVDD.n18560 1.99748
R27306 DVDD.n18584 DVDD.n18560 1.99748
R27307 DVDD.n21577 DVDD.n18560 1.99748
R27308 DVDD.n18581 DVDD.n18560 1.99748
R27309 DVDD.n21599 DVDD.n18560 1.99748
R27310 DVDD.n18578 DVDD.n18560 1.99748
R27311 DVDD.n21606 DVDD.n18560 1.99748
R27312 DVDD.n18575 DVDD.n18560 1.99748
R27313 DVDD.n21613 DVDD.n18560 1.99748
R27314 DVDD.n18572 DVDD.n18560 1.99748
R27315 DVDD.n21620 DVDD.n18560 1.99748
R27316 DVDD.n18569 DVDD.n18560 1.99748
R27317 DVDD.n21627 DVDD.n18560 1.99748
R27318 DVDD.n18566 DVDD.n18560 1.99748
R27319 DVDD.n21634 DVDD.n18560 1.99748
R27320 DVDD.n18563 DVDD.n18560 1.99748
R27321 DVDD.n21641 DVDD.n18560 1.99748
R27322 DVDD.n18560 DVDD.n18559 1.99748
R27323 DVDD.n21402 DVDD.n18560 1.99748
R27324 DVDD.n21409 DVDD.n18560 1.99748
R27325 DVDD.n21400 DVDD.n18560 1.99748
R27326 DVDD.n21416 DVDD.n18560 1.99748
R27327 DVDD.n21397 DVDD.n18560 1.99748
R27328 DVDD.n21423 DVDD.n18560 1.99748
R27329 DVDD.n21394 DVDD.n18560 1.99748
R27330 DVDD.n21430 DVDD.n18560 1.99748
R27331 DVDD.n21391 DVDD.n18560 1.99748
R27332 DVDD.n21437 DVDD.n18560 1.99748
R27333 DVDD.n21388 DVDD.n18560 1.99748
R27334 DVDD.n21446 DVDD.n18560 1.99748
R27335 DVDD.n21385 DVDD.n18560 1.99748
R27336 DVDD.n21453 DVDD.n18560 1.99748
R27337 DVDD.n21382 DVDD.n18560 1.99748
R27338 DVDD.n21460 DVDD.n18560 1.99748
R27339 DVDD.n21379 DVDD.n18560 1.99748
R27340 DVDD.n21467 DVDD.n18560 1.99748
R27341 DVDD.n21376 DVDD.n18560 1.99748
R27342 DVDD.n21474 DVDD.n18560 1.99748
R27343 DVDD.n21373 DVDD.n18560 1.99748
R27344 DVDD.n21481 DVDD.n18560 1.99748
R27345 DVDD.n21329 DVDD.n18560 1.99748
R27346 DVDD.n21488 DVDD.n18560 1.99748
R27347 DVDD.n21491 DVDD.n18560 1.99748
R27348 DVDD.n19413 DVDD.n19218 1.99748
R27349 DVDD.n19312 DVDD.n19218 1.99748
R27350 DVDD.n19420 DVDD.n19218 1.99748
R27351 DVDD.n19309 DVDD.n19218 1.99748
R27352 DVDD.n19428 DVDD.n19218 1.99748
R27353 DVDD.n19306 DVDD.n19218 1.99748
R27354 DVDD.n19435 DVDD.n19218 1.99748
R27355 DVDD.n19303 DVDD.n19218 1.99748
R27356 DVDD.n19442 DVDD.n19218 1.99748
R27357 DVDD.n19300 DVDD.n19218 1.99748
R27358 DVDD.n19449 DVDD.n19218 1.99748
R27359 DVDD.n19297 DVDD.n19218 1.99748
R27360 DVDD.n19456 DVDD.n19218 1.99748
R27361 DVDD.n19294 DVDD.n19218 1.99748
R27362 DVDD.n19463 DVDD.n19218 1.99748
R27363 DVDD.n19290 DVDD.n19218 1.99748
R27364 DVDD.n19470 DVDD.n19218 1.99748
R27365 DVDD.n19286 DVDD.n19218 1.99748
R27366 DVDD.n19477 DVDD.n19218 1.99748
R27367 DVDD.n19283 DVDD.n19218 1.99748
R27368 DVDD.n19484 DVDD.n19218 1.99748
R27369 DVDD.n19280 DVDD.n19218 1.99748
R27370 DVDD.n19491 DVDD.n19218 1.99748
R27371 DVDD.n19277 DVDD.n19218 1.99748
R27372 DVDD.n19498 DVDD.n19218 1.99748
R27373 DVDD.n19274 DVDD.n19218 1.99748
R27374 DVDD.n19507 DVDD.n19218 1.99748
R27375 DVDD.n19271 DVDD.n19218 1.99748
R27376 DVDD.n19514 DVDD.n19218 1.99748
R27377 DVDD.n19268 DVDD.n19218 1.99748
R27378 DVDD.n19521 DVDD.n19218 1.99748
R27379 DVDD.n19265 DVDD.n19218 1.99748
R27380 DVDD.n19528 DVDD.n19218 1.99748
R27381 DVDD.n19262 DVDD.n19218 1.99748
R27382 DVDD.n19535 DVDD.n19218 1.99748
R27383 DVDD.n19259 DVDD.n19218 1.99748
R27384 DVDD.n19542 DVDD.n19218 1.99748
R27385 DVDD.n19256 DVDD.n19218 1.99748
R27386 DVDD.n19549 DVDD.n19218 1.99748
R27387 DVDD.n19253 DVDD.n19218 1.99748
R27388 DVDD.n19558 DVDD.n19218 1.99748
R27389 DVDD.n19250 DVDD.n19218 1.99748
R27390 DVDD.n19565 DVDD.n19218 1.99748
R27391 DVDD.n19247 DVDD.n19218 1.99748
R27392 DVDD.n19572 DVDD.n19218 1.99748
R27393 DVDD.n19244 DVDD.n19218 1.99748
R27394 DVDD.n19579 DVDD.n19218 1.99748
R27395 DVDD.n19241 DVDD.n19218 1.99748
R27396 DVDD.n19586 DVDD.n19218 1.99748
R27397 DVDD.n19238 DVDD.n19218 1.99748
R27398 DVDD.n19593 DVDD.n19218 1.99748
R27399 DVDD.n19233 DVDD.n19218 1.99748
R27400 DVDD.n19600 DVDD.n19218 1.99748
R27401 DVDD.n19230 DVDD.n19218 1.99748
R27402 DVDD.n19607 DVDD.n19218 1.99748
R27403 DVDD.n19227 DVDD.n19218 1.99748
R27404 DVDD.n19614 DVDD.n19218 1.99748
R27405 DVDD.n19224 DVDD.n19218 1.99748
R27406 DVDD.n19621 DVDD.n19218 1.99748
R27407 DVDD.n19221 DVDD.n19218 1.99748
R27408 DVDD.n19628 DVDD.n19218 1.99748
R27409 DVDD.n19218 DVDD.n19217 1.99748
R27410 DVDD.n19324 DVDD.n19218 1.99748
R27411 DVDD.n19320 DVDD.n19218 1.99748
R27412 DVDD.n19331 DVDD.n19218 1.99748
R27413 DVDD.n3460 DVDD.n3459 1.85434
R27414 DVDD.n3450 DVDD.n3449 1.85434
R27415 DVDD.n3439 DVDD.n3438 1.85434
R27416 DVDD.n15609 DVDD.n15608 1.85434
R27417 DVDD.n15579 DVDD.n15578 1.85434
R27418 DVDD.n15570 DVDD.n15569 1.85434
R27419 DVDD.n15561 DVDD.n15560 1.85434
R27420 DVDD.n15552 DVDD.n15551 1.85434
R27421 DVDD.n15543 DVDD.n15542 1.85434
R27422 DVDD.n15533 DVDD.n15532 1.85434
R27423 DVDD.n15526 DVDD.n15525 1.85434
R27424 DVDD.n5199 DVDD.n5198 1.85434
R27425 DVDD.n5189 DVDD.n5188 1.85434
R27426 DVDD.n5178 DVDD.n5177 1.85434
R27427 DVDD.n5167 DVDD.n5166 1.85434
R27428 DVDD.n16070 DVDD.n16069 1.85434
R27429 DVDD.n16039 DVDD.n16038 1.85434
R27430 DVDD.n16028 DVDD.n16027 1.85434
R27431 DVDD.n16050 DVDD.n16049 1.85434
R27432 DVDD.n16016 DVDD.n16015 1.85434
R27433 DVDD.n16065 DVDD.n16064 1.85434
R27434 DVDD.n9783 DVDD.n9782 1.85434
R27435 DVDD.n9791 DVDD.n9775 1.85434
R27436 DVDD.n9795 DVDD.n9794 1.85434
R27437 DVDD.n9946 DVDD.n9945 1.85434
R27438 DVDD.n9804 DVDD.n9803 1.85434
R27439 DVDD.n9951 DVDD.n9950 1.85434
R27440 DVDD.n10097 DVDD.n10096 1.85434
R27441 DVDD.n10099 DVDD.n10098 1.85434
R27442 DVDD.n10106 DVDD.n9602 1.85434
R27443 DVDD.n10110 DVDD.n10109 1.85434
R27444 DVDD.n10112 DVDD.n10111 1.85434
R27445 DVDD.n10118 DVDD.n9595 1.85434
R27446 DVDD.n10122 DVDD.n10121 1.85434
R27447 DVDD.n10124 DVDD.n10123 1.85434
R27448 DVDD.n10131 DVDD.n9587 1.85434
R27449 DVDD.n10135 DVDD.n10134 1.85434
R27450 DVDD.n10137 DVDD.n10136 1.85434
R27451 DVDD.n10144 DVDD.n9579 1.85434
R27452 DVDD.n10148 DVDD.n10147 1.85434
R27453 DVDD.n10150 DVDD.n10149 1.85434
R27454 DVDD.n10160 DVDD.n9573 1.85434
R27455 DVDD.n10164 DVDD.n10163 1.85434
R27456 DVDD.n10167 DVDD.n10166 1.85434
R27457 DVDD.n10165 DVDD.n2268 1.85238
R27458 DVDD.n3457 DVDD.n3455 1.85078
R27459 DVDD.n3446 DVDD.n3444 1.85078
R27460 DVDD.n3435 DVDD.n3433 1.85078
R27461 DVDD.n15606 DVDD.n2620 1.85078
R27462 DVDD.n15575 DVDD.n15573 1.85078
R27463 DVDD.n15566 DVDD.n15564 1.85078
R27464 DVDD.n15557 DVDD.n15555 1.85078
R27465 DVDD.n15548 DVDD.n15546 1.85078
R27466 DVDD.n15539 DVDD.n15537 1.85078
R27467 DVDD.n15530 DVDD.n2804 1.85078
R27468 DVDD.n15523 DVDD.n15521 1.85078
R27469 DVDD.n5196 DVDD.n5194 1.85078
R27470 DVDD.n5185 DVDD.n5183 1.85078
R27471 DVDD.n5174 DVDD.n5172 1.85078
R27472 DVDD.n5163 DVDD.n5161 1.85078
R27473 DVDD.n3105 DVDD.n3103 1.85078
R27474 DVDD.n16035 DVDD.n16033 1.85078
R27475 DVDD.n16024 DVDD.n16022 1.85078
R27476 DVDD.n16046 DVDD.n16044 1.85078
R27477 DVDD.n16012 DVDD.n16010 1.85078
R27478 DVDD.n16062 DVDD.n2963 1.85078
R27479 DVDD.n9784 DVDD.n9781 1.85078
R27480 DVDD.n9790 DVDD.n9780 1.85078
R27481 DVDD.n9787 DVDD.n9786 1.85078
R27482 DVDD.n9942 DVDD.n9940 1.85078
R27483 DVDD.n9800 DVDD.n9798 1.85078
R27484 DVDD.n9954 DVDD.n9953 1.85078
R27485 DVDD.n9740 DVDD.n9739 1.85078
R27486 DVDD.n10101 DVDD.n9609 1.85078
R27487 DVDD.n10104 DVDD.n9607 1.85078
R27488 DVDD.n9606 DVDD.n9605 1.85078
R27489 DVDD.n10114 DVDD.n9601 1.85078
R27490 DVDD.n10117 DVDD.n9599 1.85078
R27491 DVDD.n9598 DVDD.n9597 1.85078
R27492 DVDD.n10126 DVDD.n9594 1.85078
R27493 DVDD.n10129 DVDD.n9592 1.85078
R27494 DVDD.n9591 DVDD.n9590 1.85078
R27495 DVDD.n10139 DVDD.n9586 1.85078
R27496 DVDD.n10142 DVDD.n9584 1.85078
R27497 DVDD.n9583 DVDD.n9582 1.85078
R27498 DVDD.n10152 DVDD.n9578 1.85078
R27499 DVDD.n10158 DVDD.n9576 1.85078
R27500 DVDD.n10155 DVDD.n10154 1.85043
R27501 DVDD.n19352 DVDD.t70 1.74266
R27502 DVDD.n21295 DVDD.t71 1.74266
R27503 DVDD.n21969 DVDD.n21968 1.52276
R27504 DVDD.n21822 DVDD.n21812 1.52276
R27505 DVDD.n21853 DVDD.n21844 1.52209
R27506 DVDD.n21246 DVDD.n21218 1.52209
R27507 DVDD.n21956 DVDD.n18288 1.52209
R27508 DVDD.n18470 DVDD.n124 1.52209
R27509 DVDD.n4306 DVDD.n4301 1.52209
R27510 DVDD.n3702 DVDD.n3698 1.52209
R27511 DVDD.n21697 DVDD.n18523 1.52096
R27512 DVDD.n18423 DVDD.n18412 1.52096
R27513 DVDD.n22019 DVDD.n232 1.52029
R27514 DVDD.n21348 DVDD.n21344 1.52029
R27515 DVDD.n18258 DVDD.n18255 1.52029
R27516 DVDD.n18442 DVDD.n18411 1.52029
R27517 DVDD.n4285 DVDD.n4242 1.52029
R27518 DVDD.n3686 DVDD.n3680 1.52029
R27519 DVDD.n18421 DVDD.n18420 1.5005
R27520 DVDD.n18419 DVDD.n18413 1.5005
R27521 DVDD.n18415 DVDD.n18414 1.5005
R27522 DVDD.n18379 DVDD.n178 1.5005
R27523 DVDD.n18380 DVDD.n182 1.5005
R27524 DVDD.n21850 DVDD.n21849 1.5005
R27525 DVDD.n21846 DVDD.n21845 1.5005
R27526 DVDD.n21855 DVDD.n21854 1.5005
R27527 DVDD.n18279 DVDD.n18275 1.5005
R27528 DVDD.n21973 DVDD.n21972 1.5005
R27529 DVDD.n18278 DVDD.n18276 1.5005
R27530 DVDD.n18277 DVDD.n18246 1.5005
R27531 DVDD.n22013 DVDD.n18247 1.5005
R27532 DVDD.n22016 DVDD.n22015 1.5005
R27533 DVDD.n22012 DVDD.n22010 1.5005
R27534 DVDD.n22021 DVDD.n22020 1.5005
R27535 DVDD.n21972 DVDD.n21971 1.5005
R27536 DVDD.n21970 DVDD.n18278 1.5005
R27537 DVDD.n18277 DVDD.n209 1.5005
R27538 DVDD.n22013 DVDD.n220 1.5005
R27539 DVDD.n22017 DVDD.n22016 1.5005
R27540 DVDD.n22018 DVDD.n22012 1.5005
R27541 DVDD.n21341 DVDD.n140 1.5005
R27542 DVDD.n21239 DVDD.n141 1.5005
R27543 DVDD.n21240 DVDD.n21238 1.5005
R27544 DVDD.n21243 DVDD.n21236 1.5005
R27545 DVDD.n21245 DVDD.n21244 1.5005
R27546 DVDD.n21352 DVDD.n21351 1.5005
R27547 DVDD.n21343 DVDD.n21342 1.5005
R27548 DVDD.n21347 DVDD.n21346 1.5005
R27549 DVDD.n21349 DVDD.n21343 1.5005
R27550 DVDD.n21351 DVDD.n21350 1.5005
R27551 DVDD.n21341 DVDD.n18506 1.5005
R27552 DVDD.n21239 DVDD.n18503 1.5005
R27553 DVDD.n21241 DVDD.n21240 1.5005
R27554 DVDD.n21243 DVDD.n21242 1.5005
R27555 DVDD.n21696 DVDD.n21695 1.5005
R27556 DVDD.n18525 DVDD.n18522 1.5005
R27557 DVDD.n21702 DVDD.n21701 1.5005
R27558 DVDD.n18305 DVDD.n191 1.5005
R27559 DVDD.n18304 DVDD.n192 1.5005
R27560 DVDD.n21953 DVDD.n21952 1.5005
R27561 DVDD.n18292 DVDD.n18289 1.5005
R27562 DVDD.n21958 DVDD.n21957 1.5005
R27563 DVDD.n21698 DVDD.n18522 1.5005
R27564 DVDD.n21701 DVDD.n21700 1.5005
R27565 DVDD.n21699 DVDD.n191 1.5005
R27566 DVDD.n18290 DVDD.n192 1.5005
R27567 DVDD.n21954 DVDD.n21953 1.5005
R27568 DVDD.n21955 DVDD.n18289 1.5005
R27569 DVDD.n21818 DVDD.n21817 1.5005
R27570 DVDD.n21826 DVDD.n21825 1.5005
R27571 DVDD.n21821 DVDD.n21819 1.5005
R27572 DVDD.n21820 DVDD.n18250 1.5005
R27573 DVDD.n18263 DVDD.n18262 1.5005
R27574 DVDD.n18261 DVDD.n18251 1.5005
R27575 DVDD.n18254 DVDD.n18253 1.5005
R27576 DVDD.n18257 DVDD.n18256 1.5005
R27577 DVDD.n21825 DVDD.n21824 1.5005
R27578 DVDD.n21823 DVDD.n21821 1.5005
R27579 DVDD.n21820 DVDD.n216 1.5005
R27580 DVDD.n18262 DVDD.n212 1.5005
R27581 DVDD.n18261 DVDD.n18260 1.5005
R27582 DVDD.n18259 DVDD.n18254 1.5005
R27583 DVDD.n18419 DVDD.n18418 1.5005
R27584 DVDD.n18417 DVDD.n18415 1.5005
R27585 DVDD.n18416 DVDD.n178 1.5005
R27586 DVDD.n21847 DVDD.n182 1.5005
R27587 DVDD.n21851 DVDD.n21850 1.5005
R27588 DVDD.n21852 DVDD.n21846 1.5005
R27589 DVDD.n18446 DVDD.n152 1.5005
R27590 DVDD.n18468 DVDD.n153 1.5005
R27591 DVDD.n18469 DVDD.n18467 1.5005
R27592 DVDD.n18474 DVDD.n18473 1.5005
R27593 DVDD.n18466 DVDD.n18465 1.5005
R27594 DVDD.n18445 DVDD.n18436 1.5005
R27595 DVDD.n18444 DVDD.n18437 1.5005
R27596 DVDD.n18441 DVDD.n18440 1.5005
R27597 DVDD.n18444 DVDD.n18443 1.5005
R27598 DVDD.n18445 DVDD.n18435 1.5005
R27599 DVDD.n18447 DVDD.n18446 1.5005
R27600 DVDD.n18468 DVDD.n18448 1.5005
R27601 DVDD.n18471 DVDD.n18469 1.5005
R27602 DVDD.n18473 DVDD.n18472 1.5005
R27603 DVDD.n4288 DVDD.n4286 1.5005
R27604 DVDD.n4293 DVDD.n4292 1.5005
R27605 DVDD.n4290 DVDD.n4284 1.5005
R27606 DVDD.n4298 DVDD.n4297 1.5005
R27607 DVDD.n4314 DVDD.n4313 1.5005
R27608 DVDD.n4302 DVDD.n4300 1.5005
R27609 DVDD.n4309 DVDD.n4304 1.5005
R27610 DVDD.n4308 DVDD.n4307 1.5005
R27611 DVDD.n4294 DVDD.n4293 1.5005
R27612 DVDD.n4295 DVDD.n4284 1.5005
R27613 DVDD.n4297 DVDD.n4296 1.5005
R27614 DVDD.n4313 DVDD.n4312 1.5005
R27615 DVDD.n4311 DVDD.n4300 1.5005
R27616 DVDD.n4310 DVDD.n4309 1.5005
R27617 DVDD.n3685 DVDD.n3684 1.5005
R27618 DVDD.n3682 DVDD.n3679 1.5005
R27619 DVDD.n3691 DVDD.n3690 1.5005
R27620 DVDD.n3693 DVDD.n3674 1.5005
R27621 DVDD.n3708 DVDD.n3675 1.5005
R27622 DVDD.n3706 DVDD.n3705 1.5005
R27623 DVDD.n3696 DVDD.n3695 1.5005
R27624 DVDD.n3701 DVDD.n3700 1.5005
R27625 DVDD.n3687 DVDD.n3679 1.5005
R27626 DVDD.n3690 DVDD.n3689 1.5005
R27627 DVDD.n3688 DVDD.n3674 1.5005
R27628 DVDD.n3697 DVDD.n3675 1.5005
R27629 DVDD.n3705 DVDD.n3704 1.5005
R27630 DVDD.n3703 DVDD.n3696 1.5005
R27631 DVDD.n22056 DVDD.n366 1.5005
R27632 DVDD.n22059 DVDD.n22057 1.5005
R27633 DVDD.n22060 DVDD.n18217 1.5005
R27634 DVDD.n22051 DVDD.n18215 1.5005
R27635 DVDD.n22047 DVDD.n22046 1.5005
R27636 DVDD.n21917 DVDD.n21916 1.5005
R27637 DVDD.n21913 DVDD.n21800 1.5005
R27638 DVDD.n21828 DVDD.n21804 1.5005
R27639 DVDD.n21900 DVDD.n21815 1.5005
R27640 DVDD.n21902 DVDD.n21901 1.5005
R27641 DVDD.n21859 DVDD.n21811 1.5005
R27642 DVDD.n21875 DVDD.n21874 1.5005
R27643 DVDD.n21877 DVDD.n21843 1.5005
R27644 DVDD.n21878 DVDD.n21841 1.5005
R27645 DVDD.n21866 DVDD.n21839 1.5005
R27646 DVDD.n21759 DVDD.n21758 1.5005
R27647 DVDD.n21761 DVDD.n18400 1.5005
R27648 DVDD.n21762 DVDD.n18398 1.5005
R27649 DVDD.n21753 DVDD.n18396 1.5005
R27650 DVDD.n18424 DVDD.n18404 1.5005
R27651 DVDD.n21738 DVDD.n21737 1.5005
R27652 DVDD.n18426 DVDD.n18408 1.5005
R27653 DVDD.n21592 DVDD.n165 1.5005
R27654 DVDD.n22224 DVDD.n164 1.5005
R27655 DVDD.n22225 DVDD.n162 1.5005
R27656 DVDD.n18497 DVDD.n18496 1.5005
R27657 DVDD.n18493 DVDD.n18458 1.5005
R27658 DVDD.n18485 DVDD.n18484 1.5005
R27659 DVDD.n18462 DVDD.n125 1.5005
R27660 DVDD.n22242 DVDD.n22241 1.5005
R27661 DVDD.n15149 DVDD.n5560 1.5005
R27662 DVDD.n15151 DVDD.n15150 1.5005
R27663 DVDD.n15152 DVDD.n5559 1.5005
R27664 DVDD.n15154 DVDD.n15153 1.5005
R27665 DVDD.n15155 DVDD.n5558 1.5005
R27666 DVDD.n15157 DVDD.n15156 1.5005
R27667 DVDD.n15158 DVDD.n5557 1.5005
R27668 DVDD.n15160 DVDD.n15159 1.5005
R27669 DVDD.n15161 DVDD.n5556 1.5005
R27670 DVDD.n15163 DVDD.n15162 1.5005
R27671 DVDD.n15164 DVDD.n5555 1.5005
R27672 DVDD.n15166 DVDD.n15165 1.5005
R27673 DVDD.n15167 DVDD.n5554 1.5005
R27674 DVDD.n15169 DVDD.n15168 1.5005
R27675 DVDD.n15170 DVDD.n5553 1.5005
R27676 DVDD.n15172 DVDD.n15171 1.5005
R27677 DVDD.n15173 DVDD.n5552 1.5005
R27678 DVDD.n15175 DVDD.n15174 1.5005
R27679 DVDD.n15176 DVDD.n5551 1.5005
R27680 DVDD.n15178 DVDD.n15177 1.5005
R27681 DVDD.n15179 DVDD.n5550 1.5005
R27682 DVDD.n15181 DVDD.n15180 1.5005
R27683 DVDD.n15182 DVDD.n5549 1.5005
R27684 DVDD.n15184 DVDD.n15183 1.5005
R27685 DVDD.n15185 DVDD.n5548 1.5005
R27686 DVDD.n15187 DVDD.n15186 1.5005
R27687 DVDD.n15188 DVDD.n5547 1.5005
R27688 DVDD.n15190 DVDD.n15189 1.5005
R27689 DVDD.n15191 DVDD.n5546 1.5005
R27690 DVDD.n15193 DVDD.n15192 1.5005
R27691 DVDD.n15194 DVDD.n5545 1.5005
R27692 DVDD.n15196 DVDD.n15195 1.5005
R27693 DVDD.n15197 DVDD.n5544 1.5005
R27694 DVDD.n15199 DVDD.n15198 1.5005
R27695 DVDD.n15200 DVDD.n5543 1.5005
R27696 DVDD.n15202 DVDD.n15201 1.5005
R27697 DVDD.n15203 DVDD.n5542 1.5005
R27698 DVDD.n15205 DVDD.n15204 1.5005
R27699 DVDD.n15206 DVDD.n5541 1.5005
R27700 DVDD.n15208 DVDD.n15207 1.5005
R27701 DVDD.n15209 DVDD.n5540 1.5005
R27702 DVDD.n15211 DVDD.n15210 1.5005
R27703 DVDD.n15212 DVDD.n5539 1.5005
R27704 DVDD.n15214 DVDD.n15213 1.5005
R27705 DVDD.n15215 DVDD.n5538 1.5005
R27706 DVDD.n15217 DVDD.n15216 1.5005
R27707 DVDD.n15218 DVDD.n5537 1.5005
R27708 DVDD.n15220 DVDD.n15219 1.5005
R27709 DVDD.n15221 DVDD.n5536 1.5005
R27710 DVDD.n15223 DVDD.n15222 1.5005
R27711 DVDD.n15224 DVDD.n5535 1.5005
R27712 DVDD.n15226 DVDD.n15225 1.5005
R27713 DVDD.n15227 DVDD.n5534 1.5005
R27714 DVDD.n15229 DVDD.n15228 1.5005
R27715 DVDD.n15230 DVDD.n5533 1.5005
R27716 DVDD.n15232 DVDD.n15231 1.5005
R27717 DVDD.n15233 DVDD.n5532 1.5005
R27718 DVDD.n15235 DVDD.n15234 1.5005
R27719 DVDD.n15236 DVDD.n5531 1.5005
R27720 DVDD.n15238 DVDD.n15237 1.5005
R27721 DVDD.n15239 DVDD.n5530 1.5005
R27722 DVDD.n15241 DVDD.n15240 1.5005
R27723 DVDD.n15242 DVDD.n5529 1.5005
R27724 DVDD.n15244 DVDD.n15243 1.5005
R27725 DVDD.n15245 DVDD.n5528 1.5005
R27726 DVDD.n15247 DVDD.n15246 1.5005
R27727 DVDD.n15248 DVDD.n5527 1.5005
R27728 DVDD.n15250 DVDD.n15249 1.5005
R27729 DVDD.n15251 DVDD.n5526 1.5005
R27730 DVDD.n15253 DVDD.n15252 1.5005
R27731 DVDD.n15254 DVDD.n5525 1.5005
R27732 DVDD.n15256 DVDD.n15255 1.5005
R27733 DVDD.n15257 DVDD.n5524 1.5005
R27734 DVDD.n15259 DVDD.n15258 1.5005
R27735 DVDD.n15260 DVDD.n5523 1.5005
R27736 DVDD.n15262 DVDD.n15261 1.5005
R27737 DVDD.n15263 DVDD.n5522 1.5005
R27738 DVDD.n15265 DVDD.n15264 1.5005
R27739 DVDD.n15266 DVDD.n5521 1.5005
R27740 DVDD.n15268 DVDD.n15267 1.5005
R27741 DVDD.n15269 DVDD.n5520 1.5005
R27742 DVDD.n15271 DVDD.n15270 1.5005
R27743 DVDD.n15272 DVDD.n5519 1.5005
R27744 DVDD.n15274 DVDD.n15273 1.5005
R27745 DVDD.n15275 DVDD.n5518 1.5005
R27746 DVDD.n15277 DVDD.n15276 1.5005
R27747 DVDD.n15278 DVDD.n5517 1.5005
R27748 DVDD.n15280 DVDD.n15279 1.5005
R27749 DVDD.n15281 DVDD.n5497 1.5005
R27750 DVDD.n15283 DVDD.n15282 1.5005
R27751 DVDD.n5516 DVDD.n5496 1.5005
R27752 DVDD.n5515 DVDD.n5514 1.5005
R27753 DVDD.n5513 DVDD.n5512 1.5005
R27754 DVDD.n5511 DVDD.n5510 1.5005
R27755 DVDD.n5509 DVDD.n5508 1.5005
R27756 DVDD.n5507 DVDD.n5506 1.5005
R27757 DVDD.n5505 DVDD.n5504 1.5005
R27758 DVDD.n5503 DVDD.n5502 1.5005
R27759 DVDD.n5501 DVDD.n5500 1.5005
R27760 DVDD.n5499 DVDD.n5498 1.5005
R27761 DVDD.n5476 DVDD.n5467 1.5005
R27762 DVDD.n15288 DVDD.n15287 1.5005
R27763 DVDD.n15289 DVDD.n5466 1.5005
R27764 DVDD.n15291 DVDD.n15290 1.5005
R27765 DVDD.n15292 DVDD.n5465 1.5005
R27766 DVDD.n15294 DVDD.n15293 1.5005
R27767 DVDD.n15295 DVDD.n5464 1.5005
R27768 DVDD.n15297 DVDD.n15296 1.5005
R27769 DVDD.n15298 DVDD.n5463 1.5005
R27770 DVDD.n15300 DVDD.n15299 1.5005
R27771 DVDD.n15301 DVDD.n5462 1.5005
R27772 DVDD.n15303 DVDD.n15302 1.5005
R27773 DVDD.n15304 DVDD.n5461 1.5005
R27774 DVDD.n15306 DVDD.n15305 1.5005
R27775 DVDD.n15308 DVDD.n5460 1.5005
R27776 DVDD.n15310 DVDD.n15309 1.5005
R27777 DVDD.n15311 DVDD.n5459 1.5005
R27778 DVDD.n15313 DVDD.n15312 1.5005
R27779 DVDD.n15314 DVDD.n5409 1.5005
R27780 DVDD.n15316 DVDD.n15315 1.5005
R27781 DVDD.n5458 DVDD.n5406 1.5005
R27782 DVDD.n5457 DVDD.n5456 1.5005
R27783 DVDD.n5455 DVDD.n5454 1.5005
R27784 DVDD.n5453 DVDD.n5452 1.5005
R27785 DVDD.n5451 DVDD.n5450 1.5005
R27786 DVDD.n5449 DVDD.n5448 1.5005
R27787 DVDD.n5447 DVDD.n5446 1.5005
R27788 DVDD.n5445 DVDD.n5444 1.5005
R27789 DVDD.n5443 DVDD.n5442 1.5005
R27790 DVDD.n5441 DVDD.n5440 1.5005
R27791 DVDD.n5439 DVDD.n5438 1.5005
R27792 DVDD.n5437 DVDD.n5401 1.5005
R27793 DVDD.n5436 DVDD.n5435 1.5005
R27794 DVDD.n5434 DVDD.n5433 1.5005
R27795 DVDD.n5432 DVDD.n5431 1.5005
R27796 DVDD.n5430 DVDD.n5429 1.5005
R27797 DVDD.n5428 DVDD.n5427 1.5005
R27798 DVDD.n5426 DVDD.n5425 1.5005
R27799 DVDD.n5424 DVDD.n5423 1.5005
R27800 DVDD.n5422 DVDD.n5421 1.5005
R27801 DVDD.n5420 DVDD.n5419 1.5005
R27802 DVDD.n5418 DVDD.n5417 1.5005
R27803 DVDD.n5416 DVDD.n5415 1.5005
R27804 DVDD.n5414 DVDD.n5413 1.5005
R27805 DVDD.n5412 DVDD.n5411 1.5005
R27806 DVDD.n5410 DVDD.n5376 1.5005
R27807 DVDD.n15410 DVDD.n5368 1.5005
R27808 DVDD.n15412 DVDD.n15411 1.5005
R27809 DVDD.n15413 DVDD.n5261 1.5005
R27810 DVDD.n15415 DVDD.n15414 1.5005
R27811 DVDD.n5367 DVDD.n5253 1.5005
R27812 DVDD.n5366 DVDD.n5365 1.5005
R27813 DVDD.n5364 DVDD.n5363 1.5005
R27814 DVDD.n5362 DVDD.n5361 1.5005
R27815 DVDD.n5360 DVDD.n5359 1.5005
R27816 DVDD.n5358 DVDD.n5357 1.5005
R27817 DVDD.n5356 DVDD.n5355 1.5005
R27818 DVDD.n5354 DVDD.n5353 1.5005
R27819 DVDD.n5352 DVDD.n5351 1.5005
R27820 DVDD.n5350 DVDD.n5349 1.5005
R27821 DVDD.n5348 DVDD.n5347 1.5005
R27822 DVDD.n5346 DVDD.n5345 1.5005
R27823 DVDD.n5344 DVDD.n5343 1.5005
R27824 DVDD.n5342 DVDD.n5341 1.5005
R27825 DVDD.n5340 DVDD.n5339 1.5005
R27826 DVDD.n5338 DVDD.n5337 1.5005
R27827 DVDD.n5336 DVDD.n5335 1.5005
R27828 DVDD.n5334 DVDD.n5333 1.5005
R27829 DVDD.n5332 DVDD.n5331 1.5005
R27830 DVDD.n5330 DVDD.n5329 1.5005
R27831 DVDD.n5328 DVDD.n5327 1.5005
R27832 DVDD.n5326 DVDD.n5325 1.5005
R27833 DVDD.n5324 DVDD.n5323 1.5005
R27834 DVDD.n5322 DVDD.n5321 1.5005
R27835 DVDD.n5320 DVDD.n5319 1.5005
R27836 DVDD.n5318 DVDD.n5317 1.5005
R27837 DVDD.n5316 DVDD.n5315 1.5005
R27838 DVDD.n5314 DVDD.n5313 1.5005
R27839 DVDD.n5312 DVDD.n5080 1.5005
R27840 DVDD.n5311 DVDD.n5077 1.5005
R27841 DVDD.n5310 DVDD.n5309 1.5005
R27842 DVDD.n5308 DVDD.n5307 1.5005
R27843 DVDD.n5306 DVDD.n5305 1.5005
R27844 DVDD.n5304 DVDD.n5303 1.5005
R27845 DVDD.n5302 DVDD.n5301 1.5005
R27846 DVDD.n5300 DVDD.n5299 1.5005
R27847 DVDD.n5298 DVDD.n5297 1.5005
R27848 DVDD.n5296 DVDD.n5295 1.5005
R27849 DVDD.n5294 DVDD.n5293 1.5005
R27850 DVDD.n5292 DVDD.n5291 1.5005
R27851 DVDD.n5290 DVDD.n5289 1.5005
R27852 DVDD.n5288 DVDD.n5287 1.5005
R27853 DVDD.n5286 DVDD.n5285 1.5005
R27854 DVDD.n5284 DVDD.n5283 1.5005
R27855 DVDD.n5282 DVDD.n5281 1.5005
R27856 DVDD.n5280 DVDD.n5279 1.5005
R27857 DVDD.n5278 DVDD.n5061 1.5005
R27858 DVDD.n5277 DVDD.n5276 1.5005
R27859 DVDD.n5275 DVDD.n5274 1.5005
R27860 DVDD.n5273 DVDD.n5272 1.5005
R27861 DVDD.n5271 DVDD.n5270 1.5005
R27862 DVDD.n5269 DVDD.n5268 1.5005
R27863 DVDD.n5267 DVDD.n5266 1.5005
R27864 DVDD.n5265 DVDD.n5264 1.5005
R27865 DVDD.n5263 DVDD.n5262 1.5005
R27866 DVDD.n5047 DVDD.n5039 1.5005
R27867 DVDD.n15703 DVDD.n15702 1.5005
R27868 DVDD.n15704 DVDD.n4905 1.5005
R27869 DVDD.n15706 DVDD.n15705 1.5005
R27870 DVDD.n5038 DVDD.n4893 1.5005
R27871 DVDD.n5037 DVDD.n5036 1.5005
R27872 DVDD.n5035 DVDD.n5034 1.5005
R27873 DVDD.n5033 DVDD.n5032 1.5005
R27874 DVDD.n5031 DVDD.n4891 1.5005
R27875 DVDD.n5030 DVDD.n5029 1.5005
R27876 DVDD.n5028 DVDD.n5027 1.5005
R27877 DVDD.n5026 DVDD.n5025 1.5005
R27878 DVDD.n5024 DVDD.n5023 1.5005
R27879 DVDD.n5022 DVDD.n5021 1.5005
R27880 DVDD.n5020 DVDD.n5019 1.5005
R27881 DVDD.n5018 DVDD.n5017 1.5005
R27882 DVDD.n5016 DVDD.n5015 1.5005
R27883 DVDD.n5014 DVDD.n5013 1.5005
R27884 DVDD.n5012 DVDD.n5011 1.5005
R27885 DVDD.n5010 DVDD.n5009 1.5005
R27886 DVDD.n5008 DVDD.n5007 1.5005
R27887 DVDD.n5006 DVDD.n5005 1.5005
R27888 DVDD.n5004 DVDD.n5003 1.5005
R27889 DVDD.n17738 DVDD.n877 1.5005
R27890 DVDD.n17740 DVDD.n17739 1.5005
R27891 DVDD.n17741 DVDD.n876 1.5005
R27892 DVDD.n17743 DVDD.n17742 1.5005
R27893 DVDD.n17744 DVDD.n875 1.5005
R27894 DVDD.n17746 DVDD.n17745 1.5005
R27895 DVDD.n17747 DVDD.n874 1.5005
R27896 DVDD.n17749 DVDD.n17748 1.5005
R27897 DVDD.n17750 DVDD.n873 1.5005
R27898 DVDD.n17752 DVDD.n17751 1.5005
R27899 DVDD.n17753 DVDD.n872 1.5005
R27900 DVDD.n17755 DVDD.n17754 1.5005
R27901 DVDD.n17756 DVDD.n871 1.5005
R27902 DVDD.n17758 DVDD.n17757 1.5005
R27903 DVDD.n17759 DVDD.n870 1.5005
R27904 DVDD.n17761 DVDD.n17760 1.5005
R27905 DVDD.n17762 DVDD.n869 1.5005
R27906 DVDD.n17764 DVDD.n17763 1.5005
R27907 DVDD.n17765 DVDD.n868 1.5005
R27908 DVDD.n17767 DVDD.n17766 1.5005
R27909 DVDD.n17768 DVDD.n867 1.5005
R27910 DVDD.n17770 DVDD.n17769 1.5005
R27911 DVDD.n17771 DVDD.n866 1.5005
R27912 DVDD.n17773 DVDD.n17772 1.5005
R27913 DVDD.n17774 DVDD.n865 1.5005
R27914 DVDD.n17776 DVDD.n17775 1.5005
R27915 DVDD.n17777 DVDD.n864 1.5005
R27916 DVDD.n17779 DVDD.n17778 1.5005
R27917 DVDD.n17780 DVDD.n863 1.5005
R27918 DVDD.n17782 DVDD.n17781 1.5005
R27919 DVDD.n17783 DVDD.n862 1.5005
R27920 DVDD.n17785 DVDD.n17784 1.5005
R27921 DVDD.n17786 DVDD.n861 1.5005
R27922 DVDD.n17788 DVDD.n17787 1.5005
R27923 DVDD.n17789 DVDD.n860 1.5005
R27924 DVDD.n17791 DVDD.n17790 1.5005
R27925 DVDD.n17792 DVDD.n859 1.5005
R27926 DVDD.n17794 DVDD.n17793 1.5005
R27927 DVDD.n17795 DVDD.n858 1.5005
R27928 DVDD.n17797 DVDD.n17796 1.5005
R27929 DVDD.n17798 DVDD.n857 1.5005
R27930 DVDD.n17800 DVDD.n17799 1.5005
R27931 DVDD.n17801 DVDD.n856 1.5005
R27932 DVDD.n17803 DVDD.n17802 1.5005
R27933 DVDD.n17804 DVDD.n855 1.5005
R27934 DVDD.n17806 DVDD.n17805 1.5005
R27935 DVDD.n17807 DVDD.n854 1.5005
R27936 DVDD.n17809 DVDD.n17808 1.5005
R27937 DVDD.n17810 DVDD.n853 1.5005
R27938 DVDD.n17812 DVDD.n17811 1.5005
R27939 DVDD.n17813 DVDD.n852 1.5005
R27940 DVDD.n17815 DVDD.n17814 1.5005
R27941 DVDD.n17816 DVDD.n851 1.5005
R27942 DVDD.n17818 DVDD.n17817 1.5005
R27943 DVDD.n17819 DVDD.n850 1.5005
R27944 DVDD.n17821 DVDD.n17820 1.5005
R27945 DVDD.n17822 DVDD.n849 1.5005
R27946 DVDD.n17824 DVDD.n17823 1.5005
R27947 DVDD.n17825 DVDD.n848 1.5005
R27948 DVDD.n17827 DVDD.n17826 1.5005
R27949 DVDD.n17828 DVDD.n847 1.5005
R27950 DVDD.n17830 DVDD.n17829 1.5005
R27951 DVDD.n17831 DVDD.n846 1.5005
R27952 DVDD.n17833 DVDD.n17832 1.5005
R27953 DVDD.n17834 DVDD.n845 1.5005
R27954 DVDD.n17836 DVDD.n17835 1.5005
R27955 DVDD.n17837 DVDD.n844 1.5005
R27956 DVDD.n17839 DVDD.n17838 1.5005
R27957 DVDD.n17840 DVDD.n843 1.5005
R27958 DVDD.n17842 DVDD.n17841 1.5005
R27959 DVDD.n17843 DVDD.n842 1.5005
R27960 DVDD.n17845 DVDD.n17844 1.5005
R27961 DVDD.n17846 DVDD.n841 1.5005
R27962 DVDD.n17848 DVDD.n17847 1.5005
R27963 DVDD.n17849 DVDD.n840 1.5005
R27964 DVDD.n17851 DVDD.n17850 1.5005
R27965 DVDD.n17852 DVDD.n839 1.5005
R27966 DVDD.n17854 DVDD.n17853 1.5005
R27967 DVDD.n17855 DVDD.n838 1.5005
R27968 DVDD.n17857 DVDD.n17856 1.5005
R27969 DVDD.n17858 DVDD.n837 1.5005
R27970 DVDD.n17860 DVDD.n17859 1.5005
R27971 DVDD.n17861 DVDD.n836 1.5005
R27972 DVDD.n17863 DVDD.n17862 1.5005
R27973 DVDD.n17864 DVDD.n835 1.5005
R27974 DVDD.n17866 DVDD.n17865 1.5005
R27975 DVDD.n17867 DVDD.n834 1.5005
R27976 DVDD.n17869 DVDD.n17868 1.5005
R27977 DVDD.n17870 DVDD.n833 1.5005
R27978 DVDD.n17872 DVDD.n17871 1.5005
R27979 DVDD.n17873 DVDD.n814 1.5005
R27980 DVDD.n17875 DVDD.n17874 1.5005
R27981 DVDD.n832 DVDD.n813 1.5005
R27982 DVDD.n831 DVDD.n830 1.5005
R27983 DVDD.n829 DVDD.n828 1.5005
R27984 DVDD.n827 DVDD.n826 1.5005
R27985 DVDD.n825 DVDD.n824 1.5005
R27986 DVDD.n823 DVDD.n822 1.5005
R27987 DVDD.n821 DVDD.n820 1.5005
R27988 DVDD.n819 DVDD.n818 1.5005
R27989 DVDD.n817 DVDD.n816 1.5005
R27990 DVDD.n815 DVDD.n792 1.5005
R27991 DVDD.n17879 DVDD.n784 1.5005
R27992 DVDD.n17881 DVDD.n17880 1.5005
R27993 DVDD.n17882 DVDD.n783 1.5005
R27994 DVDD.n17884 DVDD.n17883 1.5005
R27995 DVDD.n17885 DVDD.n782 1.5005
R27996 DVDD.n17887 DVDD.n17886 1.5005
R27997 DVDD.n17888 DVDD.n781 1.5005
R27998 DVDD.n17890 DVDD.n17889 1.5005
R27999 DVDD.n17891 DVDD.n780 1.5005
R28000 DVDD.n17893 DVDD.n17892 1.5005
R28001 DVDD.n17894 DVDD.n778 1.5005
R28002 DVDD.n17896 DVDD.n17895 1.5005
R28003 DVDD.n17897 DVDD.n777 1.5005
R28004 DVDD.n17899 DVDD.n17898 1.5005
R28005 DVDD.n17900 DVDD.n776 1.5005
R28006 DVDD.n17902 DVDD.n17901 1.5005
R28007 DVDD.n17903 DVDD.n775 1.5005
R28008 DVDD.n17905 DVDD.n17904 1.5005
R28009 DVDD.n17907 DVDD.n17906 1.5005
R28010 DVDD.n17909 DVDD.n17908 1.5005
R28011 DVDD.n17911 DVDD.n17910 1.5005
R28012 DVDD.n17913 DVDD.n17912 1.5005
R28013 DVDD.n17915 DVDD.n17914 1.5005
R28014 DVDD.n17917 DVDD.n17916 1.5005
R28015 DVDD.n17919 DVDD.n17918 1.5005
R28016 DVDD.n17921 DVDD.n17920 1.5005
R28017 DVDD.n17923 DVDD.n17922 1.5005
R28018 DVDD.n17925 DVDD.n17924 1.5005
R28019 DVDD.n17927 DVDD.n17926 1.5005
R28020 DVDD.n17928 DVDD.n753 1.5005
R28021 DVDD.n17930 DVDD.n17929 1.5005
R28022 DVDD.n17932 DVDD.n17931 1.5005
R28023 DVDD.n17934 DVDD.n17933 1.5005
R28024 DVDD.n17936 DVDD.n17935 1.5005
R28025 DVDD.n17938 DVDD.n17937 1.5005
R28026 DVDD.n17940 DVDD.n17939 1.5005
R28027 DVDD.n17942 DVDD.n17941 1.5005
R28028 DVDD.n17944 DVDD.n17943 1.5005
R28029 DVDD.n17946 DVDD.n17945 1.5005
R28030 DVDD.n17948 DVDD.n17947 1.5005
R28031 DVDD.n17950 DVDD.n17949 1.5005
R28032 DVDD.n17952 DVDD.n17951 1.5005
R28033 DVDD.n774 DVDD.n772 1.5005
R28034 DVDD.n773 DVDD.n738 1.5005
R28035 DVDD.n17956 DVDD.n730 1.5005
R28036 DVDD.n17958 DVDD.n17957 1.5005
R28037 DVDD.n17959 DVDD.n682 1.5005
R28038 DVDD.n17961 DVDD.n17960 1.5005
R28039 DVDD.n729 DVDD.n681 1.5005
R28040 DVDD.n728 DVDD.n727 1.5005
R28041 DVDD.n726 DVDD.n725 1.5005
R28042 DVDD.n724 DVDD.n723 1.5005
R28043 DVDD.n722 DVDD.n721 1.5005
R28044 DVDD.n720 DVDD.n719 1.5005
R28045 DVDD.n718 DVDD.n717 1.5005
R28046 DVDD.n716 DVDD.n715 1.5005
R28047 DVDD.n714 DVDD.n713 1.5005
R28048 DVDD.n712 DVDD.n711 1.5005
R28049 DVDD.n710 DVDD.n709 1.5005
R28050 DVDD.n708 DVDD.n707 1.5005
R28051 DVDD.n706 DVDD.n705 1.5005
R28052 DVDD.n704 DVDD.n703 1.5005
R28053 DVDD.n702 DVDD.n701 1.5005
R28054 DVDD.n700 DVDD.n699 1.5005
R28055 DVDD.n698 DVDD.n697 1.5005
R28056 DVDD.n696 DVDD.n695 1.5005
R28057 DVDD.n694 DVDD.n693 1.5005
R28058 DVDD.n692 DVDD.n691 1.5005
R28059 DVDD.n690 DVDD.n689 1.5005
R28060 DVDD.n688 DVDD.n687 1.5005
R28061 DVDD.n686 DVDD.n685 1.5005
R28062 DVDD.n684 DVDD.n683 1.5005
R28063 DVDD.n648 DVDD.n640 1.5005
R28064 DVDD.n17966 DVDD.n17965 1.5005
R28065 DVDD.n17968 DVDD.n17967 1.5005
R28066 DVDD.n17969 DVDD.n638 1.5005
R28067 DVDD.n17971 DVDD.n17970 1.5005
R28068 DVDD.n17973 DVDD.n17972 1.5005
R28069 DVDD.n17974 DVDD.n595 1.5005
R28070 DVDD.n17976 DVDD.n17975 1.5005
R28071 DVDD.n637 DVDD.n594 1.5005
R28072 DVDD.n636 DVDD.n635 1.5005
R28073 DVDD.n634 DVDD.n633 1.5005
R28074 DVDD.n632 DVDD.n631 1.5005
R28075 DVDD.n630 DVDD.n629 1.5005
R28076 DVDD.n628 DVDD.n627 1.5005
R28077 DVDD.n626 DVDD.n625 1.5005
R28078 DVDD.n624 DVDD.n623 1.5005
R28079 DVDD.n622 DVDD.n621 1.5005
R28080 DVDD.n620 DVDD.n619 1.5005
R28081 DVDD.n618 DVDD.n617 1.5005
R28082 DVDD.n616 DVDD.n615 1.5005
R28083 DVDD.n614 DVDD.n613 1.5005
R28084 DVDD.n612 DVDD.n611 1.5005
R28085 DVDD.n610 DVDD.n588 1.5005
R28086 DVDD.n609 DVDD.n608 1.5005
R28087 DVDD.n607 DVDD.n606 1.5005
R28088 DVDD.n605 DVDD.n604 1.5005
R28089 DVDD.n603 DVDD.n602 1.5005
R28090 DVDD.n601 DVDD.n600 1.5005
R28091 DVDD.n599 DVDD.n598 1.5005
R28092 DVDD.n597 DVDD.n596 1.5005
R28093 DVDD.n561 DVDD.n553 1.5005
R28094 DVDD.n17981 DVDD.n17980 1.5005
R28095 DVDD.n17983 DVDD.n17982 1.5005
R28096 DVDD.n17984 DVDD.n551 1.5005
R28097 DVDD.n17986 DVDD.n17985 1.5005
R28098 DVDD.n17988 DVDD.n17987 1.5005
R28099 DVDD.n17990 DVDD.n17989 1.5005
R28100 DVDD.n17992 DVDD.n17991 1.5005
R28101 DVDD.n17994 DVDD.n17993 1.5005
R28102 DVDD.n17995 DVDD.n527 1.5005
R28103 DVDD.n17997 DVDD.n17996 1.5005
R28104 DVDD.n17999 DVDD.n17998 1.5005
R28105 DVDD.n18001 DVDD.n18000 1.5005
R28106 DVDD.n18003 DVDD.n18002 1.5005
R28107 DVDD.n18005 DVDD.n18004 1.5005
R28108 DVDD.n18007 DVDD.n18006 1.5005
R28109 DVDD.n18009 DVDD.n18008 1.5005
R28110 DVDD.n18011 DVDD.n18010 1.5005
R28111 DVDD.n18013 DVDD.n18012 1.5005
R28112 DVDD.n18015 DVDD.n18014 1.5005
R28113 DVDD.n18017 DVDD.n18016 1.5005
R28114 DVDD.n18019 DVDD.n18018 1.5005
R28115 DVDD.n18021 DVDD.n18020 1.5005
R28116 DVDD.n18023 DVDD.n18022 1.5005
R28117 DVDD.n3698 DVDD.n3647 1.5005
R28118 DVDD.n3699 DVDD.n3645 1.5005
R28119 DVDD.n22185 DVDD.n232 1.5005
R28120 DVDD.n22011 DVDD.n230 1.5005
R28121 DVDD.n22023 DVDD.n22022 1.5005
R28122 DVDD.n22014 DVDD.n21984 1.5005
R28123 DVDD.n22037 DVDD.n21985 1.5005
R28124 DVDD.n21982 DVDD.n18268 1.5005
R28125 DVDD.n18274 DVDD.n18266 1.5005
R28126 DVDD.n21975 DVDD.n21974 1.5005
R28127 DVDD.n18273 DVDD.n18271 1.5005
R28128 DVDD.n21968 DVDD.n21967 1.5005
R28129 DVDD.n18288 DVDD.n18280 1.5005
R28130 DVDD.n21960 DVDD.n21959 1.5005
R28131 DVDD.n18287 DVDD.n18285 1.5005
R28132 DVDD.n21951 DVDD.n21950 1.5005
R28133 DVDD.n18293 DVDD.n18291 1.5005
R28134 DVDD.n21704 DVDD.n21703 1.5005
R28135 DVDD.n18521 DVDD.n18519 1.5005
R28136 DVDD.n21694 DVDD.n21693 1.5005
R28137 DVDD.n18526 DVDD.n18524 1.5005
R28138 DVDD.n21686 DVDD.n18523 1.5005
R28139 DVDD.n21344 DVDD.n18530 1.5005
R28140 DVDD.n21345 DVDD.n18552 1.5005
R28141 DVDD.n21653 DVDD.n18553 1.5005
R28142 DVDD.n21340 DVDD.n18551 1.5005
R28143 DVDD.n21356 DVDD.n21353 1.5005
R28144 DVDD.n21258 DVDD.n18663 1.5005
R28145 DVDD.n21237 DVDD.n18662 1.5005
R28146 DVDD.n21235 DVDD.n21234 1.5005
R28147 DVDD.n21219 DVDD.n21217 1.5005
R28148 DVDD.n21247 DVDD.n21246 1.5005
R28149 DVDD.n3680 DVDD.n3648 1.5005
R28150 DVDD.n3681 DVDD.n3644 1.5005
R28151 DVDD.n3683 DVDD.n3649 1.5005
R28152 DVDD.n3678 DVDD.n3643 1.5005
R28153 DVDD.n3692 DVDD.n3650 1.5005
R28154 DVDD.n3707 DVDD.n3651 1.5005
R28155 DVDD.n3694 DVDD.n3641 1.5005
R28156 DVDD.n4768 DVDD.n3655 1.5005
R28157 DVDD.n19378 DVDD.t72 1.16194
R28158 DVDD.t13 DVDD.n18646 1.16194
R28159 DVDD.n4381 DVDD.n4355 1.15801
R28160 DVDD.n4376 DVDD.n4365 1.15801
R28161 DVDD.n4345 DVDD.n4342 1.15801
R28162 DVDD.n3677 DVDD.n3642 1.12575
R28163 DVDD.n20900 DVDD.n18920 1.1255
R28164 DVDD.n20386 DVDD.n18919 1.1255
R28165 DVDD.n20388 DVDD.n20387 1.1255
R28166 DVDD.n20393 DVDD.n20392 1.1255
R28167 DVDD.n20394 DVDD.n20385 1.1255
R28168 DVDD.n20396 DVDD.n20395 1.1255
R28169 DVDD.n20397 DVDD.n20383 1.1255
R28170 DVDD.n20401 DVDD.n20400 1.1255
R28171 DVDD.n20403 DVDD.n20402 1.1255
R28172 DVDD.n20405 DVDD.n20404 1.1255
R28173 DVDD.n20407 DVDD.n20381 1.1255
R28174 DVDD.n20411 DVDD.n20410 1.1255
R28175 DVDD.n20413 DVDD.n20412 1.1255
R28176 DVDD.n20415 DVDD.n20414 1.1255
R28177 DVDD.n20418 DVDD.n20378 1.1255
R28178 DVDD.n19842 DVDD.n19833 1.1255
R28179 DVDD.n20423 DVDD.n20422 1.1255
R28180 DVDD.n20425 DVDD.n20424 1.1255
R28181 DVDD.n19830 DVDD.n19829 1.1255
R28182 DVDD.n20430 DVDD.n20429 1.1255
R28183 DVDD.n20431 DVDD.n19827 1.1255
R28184 DVDD.n20433 DVDD.n20432 1.1255
R28185 DVDD.n19828 DVDD.n19825 1.1255
R28186 DVDD.n20437 DVDD.n19824 1.1255
R28187 DVDD.n20439 DVDD.n20438 1.1255
R28188 DVDD.n4306 DVDD.n4262 1.1255
R28189 DVDD.n4305 DVDD.n4257 1.1255
R28190 DVDD.n18255 DVDD.n366 1.1255
R28191 DVDD.n22059 DVDD.n18218 1.1255
R28192 DVDD.n22060 DVDD.n18216 1.1255
R28193 DVDD.n18252 DVDD.n18215 1.1255
R28194 DVDD.n22046 DVDD.n18229 1.1255
R28195 DVDD.n21917 DVDD.n21801 1.1255
R28196 DVDD.n21816 DVDD.n21800 1.1255
R28197 DVDD.n21828 DVDD.n21827 1.1255
R28198 DVDD.n21900 DVDD.n21813 1.1255
R28199 DVDD.n21901 DVDD.n21812 1.1255
R28200 DVDD.n21844 DVDD.n21811 1.1255
R28201 DVDD.n21875 DVDD.n21856 1.1255
R28202 DVDD.n21877 DVDD.n21842 1.1255
R28203 DVDD.n21878 DVDD.n21840 1.1255
R28204 DVDD.n21848 DVDD.n21839 1.1255
R28205 DVDD.n21759 DVDD.n18401 1.1255
R28206 DVDD.n21761 DVDD.n18399 1.1255
R28207 DVDD.n21762 DVDD.n18397 1.1255
R28208 DVDD.n18422 DVDD.n18396 1.1255
R28209 DVDD.n18424 DVDD.n18423 1.1255
R28210 DVDD.n21737 DVDD.n18411 1.1255
R28211 DVDD.n18439 DVDD.n18426 1.1255
R28212 DVDD.n18438 DVDD.n165 1.1255
R28213 DVDD.n22224 DVDD.n163 1.1255
R28214 DVDD.n22225 DVDD.n161 1.1255
R28215 DVDD.n18497 DVDD.n18459 1.1255
R28216 DVDD.n18464 DVDD.n18458 1.1255
R28217 DVDD.n18484 DVDD.n18475 1.1255
R28218 DVDD.n18463 DVDD.n125 1.1255
R28219 DVDD.n22241 DVDD.n124 1.1255
R28220 DVDD.n4599 DVDD.n4269 1.1255
R28221 DVDD.n4303 DVDD.n4253 1.1255
R28222 DVDD.n4299 DVDD.n4268 1.1255
R28223 DVDD.n4574 DVDD.n4254 1.1255
R28224 DVDD.n4283 DVDD.n4265 1.1255
R28225 DVDD.n4291 DVDD.n4255 1.1255
R28226 DVDD.n4289 DVDD.n4264 1.1255
R28227 DVDD.n4287 DVDD.n4256 1.1255
R28228 DVDD.n4601 DVDD.n4242 1.1255
R28229 DVDD.n15121 DVDD.n15120 1.1255
R28230 DVDD.n6051 DVDD.n5994 1.1255
R28231 DVDD.n15114 DVDD.n15113 1.1255
R28232 DVDD.n6402 DVDD.n6401 1.1255
R28233 DVDD.n6698 DVDD.n6697 1.1255
R28234 DVDD.n6699 DVDD.n6348 1.1255
R28235 DVDD.n15100 DVDD.n15099 1.1255
R28236 DVDD.n6706 DVDD.n6393 1.1255
R28237 DVDD.n15093 DVDD.n15092 1.1255
R28238 DVDD.n7062 DVDD.n6752 1.1255
R28239 DVDD.n7058 DVDD.n7056 1.1255
R28240 DVDD.n15078 DVDD.n15077 1.1255
R28241 DVDD.n15071 DVDD.n15070 1.1255
R28242 DVDD.n7410 DVDD.n7069 1.1255
R28243 DVDD.n7565 DVDD.n7412 1.1255
R28244 DVDD.n7456 DVDD.n7454 1.1255
R28245 DVDD.n14866 DVDD.n7500 1.1255
R28246 DVDD.n14865 DVDD.n14864 1.1255
R28247 DVDD.n7615 DVDD.n7568 1.1255
R28248 DVDD.n9222 DVDD.n9221 1.1255
R28249 DVDD.n9561 DVDD.n9560 1.1255
R28250 DVDD.n9562 DVDD.n7678 1.1255
R28251 DVDD.n14849 DVDD.n14848 1.1255
R28252 DVDD.n8029 DVDD.n7681 1.1255
R28253 DVDD.n14842 DVDD.n14841 1.1255
R28254 DVDD.n8136 DVDD.n7733 1.1255
R28255 DVDD.n8143 DVDD.n8142 1.1255
R28256 DVDD.n8147 DVDD.n8146 1.1255
R28257 DVDD.n8149 DVDD.n8044 1.1255
R28258 DVDD.n8152 DVDD.n8087 1.1255
R28259 DVDD.n14570 DVDD.n14569 1.1255
R28260 DVDD.n8162 DVDD.n8153 1.1255
R28261 DVDD.n8253 DVDD.n8205 1.1255
R28262 DVDD.n8600 DVDD.n8256 1.1255
R28263 DVDD.n14304 DVDD.n14303 1.1255
R28264 DVDD.n10230 DVDD.n10229 1.1255
R28265 DVDD.n10231 DVDD.n10225 1.1255
R28266 DVDD.n10234 DVDD.n10233 1.1255
R28267 DVDD.n14293 DVDD.n14292 1.1255
R28268 DVDD.n10582 DVDD.n8612 1.1255
R28269 DVDD.n14286 DVDD.n14285 1.1255
R28270 DVDD.n10695 DVDD.n10286 1.1255
R28271 DVDD.n10690 DVDD.n10689 1.1255
R28272 DVDD.n10702 DVDD.n10693 1.1255
R28273 DVDD.n10703 DVDD.n10597 1.1255
R28274 DVDD.n10705 DVDD.n10640 1.1255
R28275 DVDD.n11052 DVDD.n10708 1.1255
R28276 DVDD.n14014 DVDD.n14013 1.1255
R28277 DVDD.n11220 DVDD.n11216 1.1255
R28278 DVDD.n11221 DVDD.n11061 1.1255
R28279 DVDD.n11222 DVDD.n11103 1.1255
R28280 DVDD.n13809 DVDD.n11107 1.1255
R28281 DVDD.n13808 DVDD.n11149 1.1255
R28282 DVDD.n13807 DVDD.n11227 1.1255
R28283 DVDD.n13801 DVDD.n13800 1.1255
R28284 DVDD.n11580 DVDD.n11232 1.1255
R28285 DVDD.n13786 DVDD.n13785 1.1255
R28286 DVDD.n13779 DVDD.n13778 1.1255
R28287 DVDD.n11925 DVDD.n11587 1.1255
R28288 DVDD.n13764 DVDD.n13763 1.1255
R28289 DVDD.n11936 DVDD.n11927 1.1255
R28290 DVDD.n13756 DVDD.n13755 1.1255
R28291 DVDD.n11939 DVDD.n11935 1.1255
R28292 DVDD.n12381 DVDD.n12287 1.1255
R28293 DVDD.n12383 DVDD.n12330 1.1255
R28294 DVDD.n12389 DVDD.n12386 1.1255
R28295 DVDD.n13489 DVDD.n13488 1.1255
R28296 DVDD.n12894 DVDD.n12435 1.1255
R28297 DVDD.n12895 DVDD.n12477 1.1255
R28298 DVDD.n12896 DVDD.n12737 1.1255
R28299 DVDD.n13279 DVDD.n12779 1.1255
R28300 DVDD.n13278 DVDD.n12825 1.1255
R28301 DVDD.n13277 DVDD.n12901 1.1255
R28302 DVDD.n13257 DVDD.n12900 1.1255
R28303 DVDD.n13270 DVDD.n13269 1.1255
R28304 DVDD.n13267 DVDD.n12911 1.1255
R28305 DVDD.n12910 DVDD.n2165 1.1255
R28306 DVDD.n2208 DVDD.n1820 1.1255
R28307 DVDD.n16716 DVDD.n16715 1.1255
R28308 DVDD.n16717 DVDD.n1811 1.1255
R28309 DVDD.n16726 DVDD.n16725 1.1255
R28310 DVDD.n1805 DVDD.n1804 1.1255
R28311 DVDD.n16737 DVDD.n16736 1.1255
R28312 DVDD.n16739 DVDD.n1712 1.1255
R28313 DVDD.n1755 DVDD.n1705 1.1255
R28314 DVDD.n17005 DVDD.n17004 1.1255
R28315 DVDD.n17008 DVDD.n1611 1.1255
R28316 DVDD.n17007 DVDD.n1656 1.1255
R28317 DVDD.n1654 DVDD.n1270 1.1255
R28318 DVDD.n17273 DVDD.n17272 1.1255
R28319 DVDD.n17280 DVDD.n17279 1.1255
R28320 DVDD.n1264 DVDD.n921 1.1255
R28321 DVDD.n17291 DVDD.n17290 1.1255
R28322 DVDD.n17298 DVDD.n17297 1.1255
R28323 DVDD.n17299 DVDD.n904 1.1255
R28324 DVDD.n17719 DVDD.n17718 1.1255
R28325 DVDD.n15120 DVDD.n15119 1.1255
R28326 DVDD.n5996 DVDD.n5994 1.1255
R28327 DVDD.n15115 DVDD.n15114 1.1255
R28328 DVDD.n6401 DVDD.n6400 1.1255
R28329 DVDD.n6698 DVDD.n6398 1.1255
R28330 DVDD.n6700 DVDD.n6699 1.1255
R28331 DVDD.n15099 DVDD.n15098 1.1255
R28332 DVDD.n6395 DVDD.n6393 1.1255
R28333 DVDD.n15094 DVDD.n15093 1.1255
R28334 DVDD.n7063 DVDD.n7062 1.1255
R28335 DVDD.n7060 DVDD.n7058 1.1255
R28336 DVDD.n15077 DVDD.n15076 1.1255
R28337 DVDD.n15072 DVDD.n15071 1.1255
R28338 DVDD.n7069 DVDD.n7068 1.1255
R28339 DVDD.n7566 DVDD.n7565 1.1255
R28340 DVDD.n14868 DVDD.n7456 1.1255
R28341 DVDD.n14867 DVDD.n14866 1.1255
R28342 DVDD.n14865 DVDD.n7567 1.1255
R28343 DVDD.n9569 DVDD.n7568 1.1255
R28344 DVDD.n9567 DVDD.n9221 1.1255
R28345 DVDD.n9561 DVDD.n9220 1.1255
R28346 DVDD.n9563 DVDD.n9562 1.1255
R28347 DVDD.n14848 DVDD.n14847 1.1255
R28348 DVDD.n7683 DVDD.n7681 1.1255
R28349 DVDD.n14843 DVDD.n14842 1.1255
R28350 DVDD.n8137 DVDD.n8136 1.1255
R28351 DVDD.n8142 DVDD.n8141 1.1255
R28352 DVDD.n8147 DVDD.n8134 1.1255
R28353 DVDD.n14575 DVDD.n8149 1.1255
R28354 DVDD.n8152 DVDD.n8135 1.1255
R28355 DVDD.n14571 DVDD.n14570 1.1255
R28356 DVDD.n8153 DVDD.n8151 1.1255
R28357 DVDD.n14309 DVDD.n8253 1.1255
R28358 DVDD.n8256 DVDD.n8251 1.1255
R28359 DVDD.n14305 DVDD.n14304 1.1255
R28360 DVDD.n10229 DVDD.n10228 1.1255
R28361 DVDD.n10225 DVDD.n10224 1.1255
R28362 DVDD.n10235 DVDD.n10234 1.1255
R28363 DVDD.n14292 DVDD.n14291 1.1255
R28364 DVDD.n8614 DVDD.n8612 1.1255
R28365 DVDD.n14287 DVDD.n14286 1.1255
R28366 DVDD.n10696 DVDD.n10695 1.1255
R28367 DVDD.n10694 DVDD.n10689 1.1255
R28368 DVDD.n10702 DVDD.n10701 1.1255
R28369 DVDD.n10703 DVDD.n10687 1.1255
R28370 DVDD.n14019 DVDD.n10705 1.1255
R28371 DVDD.n10708 DVDD.n10688 1.1255
R28372 DVDD.n14015 DVDD.n14014 1.1255
R28373 DVDD.n11220 DVDD.n11219 1.1255
R28374 DVDD.n11221 DVDD.n11214 1.1255
R28375 DVDD.n11223 DVDD.n11222 1.1255
R28376 DVDD.n13810 DVDD.n13809 1.1255
R28377 DVDD.n13808 DVDD.n11225 1.1255
R28378 DVDD.n13807 DVDD.n13806 1.1255
R28379 DVDD.n13802 DVDD.n13801 1.1255
R28380 DVDD.n11232 DVDD.n11231 1.1255
R28381 DVDD.n13785 DVDD.n13784 1.1255
R28382 DVDD.n13780 DVDD.n13779 1.1255
R28383 DVDD.n11587 DVDD.n11586 1.1255
R28384 DVDD.n13763 DVDD.n13762 1.1255
R28385 DVDD.n11928 DVDD.n11927 1.1255
R28386 DVDD.n13757 DVDD.n13756 1.1255
R28387 DVDD.n11935 DVDD.n11933 1.1255
R28388 DVDD.n12381 DVDD.n12379 1.1255
R28389 DVDD.n13494 DVDD.n12383 1.1255
R28390 DVDD.n12386 DVDD.n12380 1.1255
R28391 DVDD.n13490 DVDD.n13489 1.1255
R28392 DVDD.n12894 DVDD.n12893 1.1255
R28393 DVDD.n12895 DVDD.n12890 1.1255
R28394 DVDD.n12897 DVDD.n12896 1.1255
R28395 DVDD.n13280 DVDD.n13279 1.1255
R28396 DVDD.n13278 DVDD.n12899 1.1255
R28397 DVDD.n13277 DVDD.n13276 1.1255
R28398 DVDD.n12902 DVDD.n12900 1.1255
R28399 DVDD.n13271 DVDD.n13270 1.1255
R28400 DVDD.n12911 DVDD.n12907 1.1255
R28401 DVDD.n12910 DVDD.n2255 1.1255
R28402 DVDD.n16454 DVDD.n1820 1.1255
R28403 DVDD.n16716 DVDD.n1819 1.1255
R28404 DVDD.n16718 DVDD.n16717 1.1255
R28405 DVDD.n16725 DVDD.n16724 1.1255
R28406 DVDD.n1816 DVDD.n1804 1.1255
R28407 DVDD.n16737 DVDD.n1802 1.1255
R28408 DVDD.n16743 DVDD.n16739 1.1255
R28409 DVDD.n1803 DVDD.n1705 1.1255
R28410 DVDD.n17005 DVDD.n1703 1.1255
R28411 DVDD.n17011 DVDD.n17008 1.1255
R28412 DVDD.n17007 DVDD.n1704 1.1255
R28413 DVDD.n1270 DVDD.n1269 1.1255
R28414 DVDD.n17274 DVDD.n17273 1.1255
R28415 DVDD.n17279 DVDD.n17278 1.1255
R28416 DVDD.n921 DVDD.n920 1.1255
R28417 DVDD.n17292 DVDD.n17291 1.1255
R28418 DVDD.n17297 DVDD.n17296 1.1255
R28419 DVDD.n904 DVDD.n902 1.1255
R28420 DVDD.n17720 DVDD.n17719 1.1255
R28421 DVDD.n17721 DVDD.n17720 1.1255
R28422 DVDD.n902 DVDD.n901 1.1255
R28423 DVDD.n17296 DVDD.n17295 1.1255
R28424 DVDD.n17293 DVDD.n17292 1.1255
R28425 DVDD.n920 DVDD.n919 1.1255
R28426 DVDD.n17278 DVDD.n17277 1.1255
R28427 DVDD.n17275 DVDD.n17274 1.1255
R28428 DVDD.n1269 DVDD.n1268 1.1255
R28429 DVDD.n17009 DVDD.n1704 1.1255
R28430 DVDD.n17011 DVDD.n17010 1.1255
R28431 DVDD.n16740 DVDD.n1703 1.1255
R28432 DVDD.n16741 DVDD.n1803 1.1255
R28433 DVDD.n16743 DVDD.n16742 1.1255
R28434 DVDD.n16721 DVDD.n1802 1.1255
R28435 DVDD.n16722 DVDD.n1816 1.1255
R28436 DVDD.n16724 DVDD.n16723 1.1255
R28437 DVDD.n16719 DVDD.n16718 1.1255
R28438 DVDD.n1819 DVDD.n1818 1.1255
R28439 DVDD.n16454 DVDD.n16453 1.1255
R28440 DVDD.n12904 DVDD.n2255 1.1255
R28441 DVDD.n12907 DVDD.n12905 1.1255
R28442 DVDD.n13272 DVDD.n13271 1.1255
R28443 DVDD.n13274 DVDD.n12902 1.1255
R28444 DVDD.n13276 DVDD.n13275 1.1255
R28445 DVDD.n12899 DVDD.n12889 1.1255
R28446 DVDD.n13281 DVDD.n13280 1.1255
R28447 DVDD.n12897 DVDD.n12888 1.1255
R28448 DVDD.n12891 DVDD.n12890 1.1255
R28449 DVDD.n12893 DVDD.n12892 1.1255
R28450 DVDD.n13491 DVDD.n13490 1.1255
R28451 DVDD.n13492 DVDD.n12380 1.1255
R28452 DVDD.n13494 DVDD.n13493 1.1255
R28453 DVDD.n12379 DVDD.n12378 1.1255
R28454 DVDD.n11933 DVDD.n11931 1.1255
R28455 DVDD.n13758 DVDD.n13757 1.1255
R28456 DVDD.n13760 DVDD.n11928 1.1255
R28457 DVDD.n13762 DVDD.n13761 1.1255
R28458 DVDD.n11586 DVDD.n11585 1.1255
R28459 DVDD.n13781 DVDD.n13780 1.1255
R28460 DVDD.n13784 DVDD.n13783 1.1255
R28461 DVDD.n11231 DVDD.n11230 1.1255
R28462 DVDD.n13803 DVDD.n13802 1.1255
R28463 DVDD.n13806 DVDD.n13805 1.1255
R28464 DVDD.n11225 DVDD.n11213 1.1255
R28465 DVDD.n13811 DVDD.n13810 1.1255
R28466 DVDD.n11223 DVDD.n11212 1.1255
R28467 DVDD.n11217 DVDD.n11214 1.1255
R28468 DVDD.n11219 DVDD.n11218 1.1255
R28469 DVDD.n14016 DVDD.n14015 1.1255
R28470 DVDD.n14017 DVDD.n10688 1.1255
R28471 DVDD.n14019 DVDD.n14018 1.1255
R28472 DVDD.n10699 DVDD.n10687 1.1255
R28473 DVDD.n10701 DVDD.n10700 1.1255
R28474 DVDD.n10698 DVDD.n10694 1.1255
R28475 DVDD.n10697 DVDD.n10696 1.1255
R28476 DVDD.n14288 DVDD.n14287 1.1255
R28477 DVDD.n14289 DVDD.n8614 1.1255
R28478 DVDD.n14291 DVDD.n14290 1.1255
R28479 DVDD.n10236 DVDD.n10235 1.1255
R28480 DVDD.n10226 DVDD.n10224 1.1255
R28481 DVDD.n10228 DVDD.n10227 1.1255
R28482 DVDD.n14306 DVDD.n14305 1.1255
R28483 DVDD.n14307 DVDD.n8251 1.1255
R28484 DVDD.n14309 DVDD.n14308 1.1255
R28485 DVDD.n8151 DVDD.n8150 1.1255
R28486 DVDD.n14572 DVDD.n14571 1.1255
R28487 DVDD.n14573 DVDD.n8135 1.1255
R28488 DVDD.n14575 DVDD.n14574 1.1255
R28489 DVDD.n8139 DVDD.n8134 1.1255
R28490 DVDD.n8141 DVDD.n8140 1.1255
R28491 DVDD.n8138 DVDD.n8137 1.1255
R28492 DVDD.n14844 DVDD.n14843 1.1255
R28493 DVDD.n14845 DVDD.n7683 1.1255
R28494 DVDD.n14847 DVDD.n14846 1.1255
R28495 DVDD.n9564 DVDD.n9563 1.1255
R28496 DVDD.n9565 DVDD.n9220 1.1255
R28497 DVDD.n9567 DVDD.n9566 1.1255
R28498 DVDD.n9570 DVDD.n9569 1.1255
R28499 DVDD.n8974 DVDD.n7567 1.1255
R28500 DVDD.n14867 DVDD.n7564 1.1255
R28501 DVDD.n14869 DVDD.n14868 1.1255
R28502 DVDD.n7566 DVDD.n7563 1.1255
R28503 DVDD.n7068 DVDD.n7067 1.1255
R28504 DVDD.n15073 DVDD.n15072 1.1255
R28505 DVDD.n15076 DVDD.n15075 1.1255
R28506 DVDD.n7065 DVDD.n7060 1.1255
R28507 DVDD.n7064 DVDD.n7063 1.1255
R28508 DVDD.n15095 DVDD.n15094 1.1255
R28509 DVDD.n15096 DVDD.n6395 1.1255
R28510 DVDD.n15098 DVDD.n15097 1.1255
R28511 DVDD.n6701 DVDD.n6700 1.1255
R28512 DVDD.n6398 DVDD.n6397 1.1255
R28513 DVDD.n6400 DVDD.n6399 1.1255
R28514 DVDD.n15116 DVDD.n15115 1.1255
R28515 DVDD.n15117 DVDD.n5996 1.1255
R28516 DVDD.n15119 DVDD.n15118 1.1255
R28517 DVDD.n20593 DVDD.n20592 1.1255
R28518 DVDD.n20591 DVDD.n19713 1.1255
R28519 DVDD.n20590 DVDD.n20589 1.1255
R28520 DVDD.n19715 DVDD.n19714 1.1255
R28521 DVDD.n20585 DVDD.n20584 1.1255
R28522 DVDD.n20583 DVDD.n19717 1.1255
R28523 DVDD.n20582 DVDD.n20581 1.1255
R28524 DVDD.n19719 DVDD.n19718 1.1255
R28525 DVDD.n20577 DVDD.n20576 1.1255
R28526 DVDD.n20575 DVDD.n20574 1.1255
R28527 DVDD.n19732 DVDD.n19723 1.1255
R28528 DVDD.n19755 DVDD.n19751 1.1255
R28529 DVDD.n20570 DVDD.n20569 1.1255
R28530 DVDD.n20568 DVDD.n20567 1.1255
R28531 DVDD.n20564 DVDD.n19756 1.1255
R28532 DVDD.n20562 DVDD.n20561 1.1255
R28533 DVDD.n20560 DVDD.n20559 1.1255
R28534 DVDD.n20558 DVDD.n20557 1.1255
R28535 DVDD.n20554 DVDD.n19758 1.1255
R28536 DVDD.n20553 DVDD.n20552 1.1255
R28537 DVDD.n20551 DVDD.n19760 1.1255
R28538 DVDD.n20550 DVDD.n20549 1.1255
R28539 DVDD.n19762 DVDD.n19761 1.1255
R28540 DVDD.n20545 DVDD.n20544 1.1255
R28541 DVDD.n20543 DVDD.n19764 1.1255
R28542 DVDD.n22185 DVDD.n22184 1.1255
R28543 DVDD.n233 DVDD.n230 1.1255
R28544 DVDD.n22024 DVDD.n22023 1.1255
R28545 DVDD.n22033 DVDD.n21984 1.1255
R28546 DVDD.n22037 DVDD.n22036 1.1255
R28547 DVDD.n21982 DVDD.n21981 1.1255
R28548 DVDD.n21978 DVDD.n18266 1.1255
R28549 DVDD.n21976 DVDD.n21975 1.1255
R28550 DVDD.n18271 DVDD.n18270 1.1255
R28551 DVDD.n21967 DVDD.n21966 1.1255
R28552 DVDD.n21963 DVDD.n18280 1.1255
R28553 DVDD.n21961 DVDD.n21960 1.1255
R28554 DVDD.n18285 DVDD.n18284 1.1255
R28555 DVDD.n21950 DVDD.n21949 1.1255
R28556 DVDD.n21946 DVDD.n18293 1.1255
R28557 DVDD.n21705 DVDD.n21704 1.1255
R28558 DVDD.n18519 DVDD.n18518 1.1255
R28559 DVDD.n21693 DVDD.n21692 1.1255
R28560 DVDD.n21688 DVDD.n18526 1.1255
R28561 DVDD.n21687 DVDD.n21686 1.1255
R28562 DVDD.n21648 DVDD.n18530 1.1255
R28563 DVDD.n21649 DVDD.n18552 1.1255
R28564 DVDD.n21653 DVDD.n21652 1.1255
R28565 DVDD.n18555 DVDD.n18551 1.1255
R28566 DVDD.n21356 DVDD.n21355 1.1255
R28567 DVDD.n21258 DVDD.n21257 1.1255
R28568 DVDD.n21254 DVDD.n18662 1.1255
R28569 DVDD.n21234 DVDD.n18666 1.1255
R28570 DVDD.n21217 DVDD.n21216 1.1255
R28571 DVDD.n21248 DVDD.n21247 1.1255
R28572 DVDD.n3459 DVDD 1.09758
R28573 DVDD.n3449 DVDD 1.09758
R28574 DVDD.n3438 DVDD 1.09758
R28575 DVDD.n15608 DVDD 1.09758
R28576 DVDD.n15578 DVDD 1.09758
R28577 DVDD.n15569 DVDD 1.09758
R28578 DVDD.n15560 DVDD 1.09758
R28579 DVDD.n15551 DVDD 1.09758
R28580 DVDD.n15542 DVDD 1.09758
R28581 DVDD.n15532 DVDD 1.09758
R28582 DVDD.n15525 DVDD 1.09758
R28583 DVDD.n5198 DVDD 1.09758
R28584 DVDD.n5188 DVDD 1.09758
R28585 DVDD.n5177 DVDD 1.09758
R28586 DVDD.n5166 DVDD 1.09758
R28587 DVDD.n16070 DVDD 1.09758
R28588 DVDD.n16038 DVDD 1.09758
R28589 DVDD.n16027 DVDD 1.09758
R28590 DVDD.n16049 DVDD 1.09758
R28591 DVDD.n16015 DVDD 1.09758
R28592 DVDD.n16064 DVDD 1.09758
R28593 DVDD DVDD.n9783 1.09758
R28594 DVDD.n9791 DVDD 1.09758
R28595 DVDD.n9794 DVDD 1.09758
R28596 DVDD.n9945 DVDD 1.09758
R28597 DVDD.n9803 DVDD 1.09758
R28598 DVDD DVDD.n9951 1.09758
R28599 DVDD.n10096 DVDD 1.09758
R28600 DVDD DVDD.n10099 1.09758
R28601 DVDD.n10106 DVDD 1.09758
R28602 DVDD.n10109 DVDD 1.09758
R28603 DVDD DVDD.n10112 1.09758
R28604 DVDD.n10118 DVDD 1.09758
R28605 DVDD.n10121 DVDD 1.09758
R28606 DVDD DVDD.n10124 1.09758
R28607 DVDD.n10131 DVDD 1.09758
R28608 DVDD.n10134 DVDD 1.09758
R28609 DVDD DVDD.n10137 1.09758
R28610 DVDD.n10144 DVDD 1.09758
R28611 DVDD.n10147 DVDD 1.09758
R28612 DVDD DVDD.n10150 1.09758
R28613 DVDD.n10160 DVDD 1.09758
R28614 DVDD.n10163 DVDD 1.09758
R28615 DVDD.n10166 DVDD 1.09758
R28616 DVDD.n10155 DVDD 1.09186
R28617 DVDD DVDD.n3457 1.09158
R28618 DVDD DVDD.n3446 1.09158
R28619 DVDD DVDD.n3435 1.09158
R28620 DVDD DVDD.n15606 1.09158
R28621 DVDD DVDD.n15575 1.09158
R28622 DVDD DVDD.n15566 1.09158
R28623 DVDD DVDD.n15557 1.09158
R28624 DVDD DVDD.n15548 1.09158
R28625 DVDD DVDD.n15539 1.09158
R28626 DVDD DVDD.n15530 1.09158
R28627 DVDD DVDD.n15523 1.09158
R28628 DVDD DVDD.n5196 1.09158
R28629 DVDD DVDD.n5185 1.09158
R28630 DVDD DVDD.n5174 1.09158
R28631 DVDD DVDD.n5163 1.09158
R28632 DVDD DVDD.n3105 1.09158
R28633 DVDD DVDD.n16035 1.09158
R28634 DVDD DVDD.n16024 1.09158
R28635 DVDD DVDD.n16046 1.09158
R28636 DVDD DVDD.n16012 1.09158
R28637 DVDD DVDD.n16062 1.09158
R28638 DVDD.n9784 DVDD 1.09158
R28639 DVDD DVDD.n9790 1.09158
R28640 DVDD.n9787 DVDD 1.09158
R28641 DVDD DVDD.n9942 1.09158
R28642 DVDD DVDD.n9800 1.09158
R28643 DVDD.n9953 DVDD 1.09158
R28644 DVDD.n9739 DVDD 1.09158
R28645 DVDD.n10101 DVDD 1.09158
R28646 DVDD DVDD.n10104 1.09158
R28647 DVDD.n9605 DVDD 1.09158
R28648 DVDD.n10114 DVDD 1.09158
R28649 DVDD DVDD.n10117 1.09158
R28650 DVDD.n9597 DVDD 1.09158
R28651 DVDD.n10126 DVDD 1.09158
R28652 DVDD DVDD.n10129 1.09158
R28653 DVDD.n9590 DVDD 1.09158
R28654 DVDD.n10139 DVDD 1.09158
R28655 DVDD DVDD.n10142 1.09158
R28656 DVDD.n9582 DVDD 1.09158
R28657 DVDD.n10152 DVDD 1.09158
R28658 DVDD DVDD.n10158 1.09158
R28659 DVDD DVDD.n10165 1.09158
R28660 DVDD.n4353 DVDD.n4339 1.086
R28661 DVDD.n4373 DVDD.n4372 1.06706
R28662 DVDD.n18344 DVDD.n18337 0.911483
R28663 DVDD.n18369 DVDD.n18311 0.910783
R28664 DVDD.n21270 DVDD.n18656 0.910783
R28665 DVDD.n4879 DVDD.n4878 0.910783
R28666 DVDD.n4847 DVDD.n4846 0.910649
R28667 DVDD.n21683 DVDD.n18535 0.909949
R28668 DVDD.n22004 DVDD.n21995 0.909949
R28669 DVDD.n21367 DVDD.n21366 0.909949
R28670 DVDD.n17713 DVDD.n17712 0.902975
R28671 DVDD.n15127 DVDD.n15126 0.902975
R28672 DVDD.n21681 DVDD.n21680 0.9005
R28673 DVDD.n21679 DVDD.n18537 0.9005
R28674 DVDD.n21675 DVDD.n21674 0.9005
R28675 DVDD.n18378 DVDD.n183 0.9005
R28676 DVDD.n18302 DVDD.n184 0.9005
R28677 DVDD.n18373 DVDD.n18372 0.9005
R28678 DVDD.n18312 DVDD.n18309 0.9005
R28679 DVDD.n18368 DVDD.n18367 0.9005
R28680 DVDD.n21679 DVDD.n21678 0.9005
R28681 DVDD.n21677 DVDD.n21675 0.9005
R28682 DVDD.n21676 DVDD.n183 0.9005
R28683 DVDD.n18310 DVDD.n184 0.9005
R28684 DVDD.n18372 DVDD.n18371 0.9005
R28685 DVDD.n18370 DVDD.n18309 0.9005
R28686 DVDD.n18343 DVDD.n18342 0.9005
R28687 DVDD.n18335 DVDD.n18333 0.9005
R28688 DVDD.n18348 DVDD.n18347 0.9005
R28689 DVDD.n18336 DVDD.n18245 0.9005
R28690 DVDD.n21996 DVDD.n18244 0.9005
R28691 DVDD.n22001 DVDD.n22000 0.9005
R28692 DVDD.n21994 DVDD.n21992 0.9005
R28693 DVDD.n22006 DVDD.n22005 0.9005
R28694 DVDD.n18345 DVDD.n18335 0.9005
R28695 DVDD.n18347 DVDD.n18346 0.9005
R28696 DVDD.n18336 DVDD.n207 0.9005
R28697 DVDD.n21996 DVDD.n208 0.9005
R28698 DVDD.n22002 DVDD.n22001 0.9005
R28699 DVDD.n22003 DVDD.n21994 0.9005
R28700 DVDD.n21336 DVDD.n138 0.9005
R28701 DVDD.n21263 DVDD.n143 0.9005
R28702 DVDD.n21264 DVDD.n21262 0.9005
R28703 DVDD.n21267 DVDD.n18658 0.9005
R28704 DVDD.n21269 DVDD.n21268 0.9005
R28705 DVDD.n21338 DVDD.n21337 0.9005
R28706 DVDD.n21364 DVDD.n21363 0.9005
R28707 DVDD.n21334 DVDD.n21333 0.9005
R28708 DVDD.n21365 DVDD.n21364 0.9005
R28709 DVDD.n21337 DVDD.n21335 0.9005
R28710 DVDD.n21336 DVDD.n18434 0.9005
R28711 DVDD.n21263 DVDD.n18433 0.9005
R28712 DVDD.n21265 DVDD.n21264 0.9005
R28713 DVDD.n21267 DVDD.n21266 0.9005
R28714 DVDD.n3549 DVDD.n3548 0.9005
R28715 DVDD.n4850 DVDD.n4849 0.9005
R28716 DVDD.n3545 DVDD.n3544 0.9005
R28717 DVDD.n4859 DVDD.n4858 0.9005
R28718 DVDD.n4864 DVDD.n4863 0.9005
R28719 DVDD.n4865 DVDD.n3535 0.9005
R28720 DVDD.n4876 DVDD.n4875 0.9005
R28721 DVDD.n3533 DVDD.n3532 0.9005
R28722 DVDD.n4849 DVDD.n4848 0.9005
R28723 DVDD.n3544 DVDD.n3543 0.9005
R28724 DVDD.n4860 DVDD.n4859 0.9005
R28725 DVDD.n4863 DVDD.n4862 0.9005
R28726 DVDD.n3535 DVDD.n3534 0.9005
R28727 DVDD.n4877 DVDD.n4876 0.9005
R28728 DVDD.n21684 DVDD.n21683 0.9005
R28729 DVDD.n21682 DVDD.n18534 0.9005
R28730 DVDD.n18539 DVDD.n18536 0.9005
R28731 DVDD.n21671 DVDD.n18538 0.9005
R28732 DVDD.n21673 DVDD.n21672 0.9005
R28733 DVDD.n18375 DVDD.n18374 0.9005
R28734 DVDD.n18308 DVDD.n18307 0.9005
R28735 DVDD.n18314 DVDD.n18313 0.9005
R28736 DVDD.n18366 DVDD.n18365 0.9005
R28737 DVDD.n18364 DVDD.n18311 0.9005
R28738 DVDD.n18337 DVDD.n18315 0.9005
R28739 DVDD.n18341 DVDD.n18340 0.9005
R28740 DVDD.n18338 DVDD.n18331 0.9005
R28741 DVDD.n18350 DVDD.n18349 0.9005
R28742 DVDD.n18334 DVDD.n18332 0.9005
R28743 DVDD.n21998 DVDD.n21997 0.9005
R28744 DVDD.n21999 DVDD.n21990 0.9005
R28745 DVDD.n22008 DVDD.n22007 0.9005
R28746 DVDD.n21993 DVDD.n21991 0.9005
R28747 DVDD.n21995 DVDD.n229 0.9005
R28748 DVDD.n4846 DVDD.n4845 0.9005
R28749 DVDD.n4842 DVDD.n3550 0.9005
R28750 DVDD.n4840 DVDD.n3547 0.9005
R28751 DVDD.n4852 DVDD.n4851 0.9005
R28752 DVDD.n4857 DVDD.n4856 0.9005
R28753 DVDD.n4854 DVDD.n3540 0.9005
R28754 DVDD.n4867 DVDD.n4866 0.9005
R28755 DVDD.n4869 DVDD.n3536 0.9005
R28756 DVDD.n4874 DVDD.n4873 0.9005
R28757 DVDD.n4871 DVDD.n3537 0.9005
R28758 DVDD.n4880 DVDD.n4879 0.9005
R28759 DVDD.n21271 DVDD.n21270 0.9005
R28760 DVDD.n18657 DVDD.n18654 0.9005
R28761 DVDD.n21222 DVDD.n21221 0.9005
R28762 DVDD.n18660 DVDD.n18659 0.9005
R28763 DVDD.n21261 DVDD.n21260 0.9005
R28764 DVDD.n21359 DVDD.n21358 0.9005
R28765 DVDD.n21361 DVDD.n21360 0.9005
R28766 DVDD.n21362 DVDD.n18549 0.9005
R28767 DVDD.n21369 DVDD.n21368 0.9005
R28768 DVDD.n21367 DVDD.n18533 0.9005
R28769 DVDD.n18103 DVDD.n18045 0.9005
R28770 DVDD.n18105 DVDD.n501 0.9005
R28771 DVDD.n18106 DVDD.n18046 0.9005
R28772 DVDD.n18102 DVDD.n500 0.9005
R28773 DVDD.n18097 DVDD.n18047 0.9005
R28774 DVDD.n18095 DVDD.n18048 0.9005
R28775 DVDD.n18093 DVDD.n498 0.9005
R28776 DVDD.n18065 DVDD.n18049 0.9005
R28777 DVDD.n18123 DVDD.n497 0.9005
R28778 DVDD.n18125 DVDD.n18124 0.9005
R28779 DVDD.n22069 DVDD.n22068 0.9005
R28780 DVDD.n18206 DVDD.n18204 0.9005
R28781 DVDD.n22063 DVDD.n22062 0.9005
R28782 DVDD.n18212 DVDD.n18210 0.9005
R28783 DVDD.n22044 DVDD.n22043 0.9005
R28784 DVDD.n21920 DVDD.n21919 0.9005
R28785 DVDD.n21798 DVDD.n21797 0.9005
R28786 DVDD.n21897 DVDD.n21896 0.9005
R28787 DVDD.n21793 DVDD.n21791 0.9005
R28788 DVDD.n21930 DVDD.n21929 0.9005
R28789 DVDD.n21931 DVDD.n21784 0.9005
R28790 DVDD.n21933 DVDD.n21932 0.9005
R28791 DVDD.n21787 DVDD.n21786 0.9005
R28792 DVDD.n21781 DVDD.n21780 0.9005
R28793 DVDD.n21942 DVDD.n21941 0.9005
R28794 DVDD.n21778 DVDD.n21777 0.9005
R28795 DVDD.n18388 DVDD.n18386 0.9005
R28796 DVDD.n21767 DVDD.n21766 0.9005
R28797 DVDD.n21768 DVDD.n18391 0.9005
R28798 DVDD.n21770 DVDD.n21769 0.9005
R28799 DVDD.n21732 DVDD.n18392 0.9005
R28800 DVDD.n22239 DVDD.n22238 0.9005
R28801 DVDD.n131 DVDD.n129 0.9005
R28802 DVDD.n18482 DVDD.n18481 0.9005
R28803 DVDD.n18480 DVDD.n18479 0.9005
R28804 DVDD.n157 DVDD.n134 0.9005
R28805 DVDD.n22227 DVDD.n159 0.9005
R28806 DVDD.n21726 DVDD.n158 0.9005
R28807 DVDD.n21727 DVDD.n18427 0.9005
R28808 DVDD.n21734 DVDD.n21733 0.9005
R28809 DVDD.n17613 DVDD.n17611 0.9005
R28810 DVDD.n17614 DVDD.n17610 0.9005
R28811 DVDD.n17615 DVDD.n17609 0.9005
R28812 DVDD.n17616 DVDD.n17608 0.9005
R28813 DVDD.n17617 DVDD.n17607 0.9005
R28814 DVDD.n17618 DVDD.n17606 0.9005
R28815 DVDD.n17619 DVDD.n17605 0.9005
R28816 DVDD.n17620 DVDD.n17604 0.9005
R28817 DVDD.n17621 DVDD.n17603 0.9005
R28818 DVDD.n17622 DVDD.n17602 0.9005
R28819 DVDD.n17623 DVDD.n17601 0.9005
R28820 DVDD.n17624 DVDD.n17600 0.9005
R28821 DVDD.n17625 DVDD.n17599 0.9005
R28822 DVDD.n17626 DVDD.n17598 0.9005
R28823 DVDD.n17627 DVDD.n17597 0.9005
R28824 DVDD.n17628 DVDD.n17596 0.9005
R28825 DVDD.n17629 DVDD.n17595 0.9005
R28826 DVDD.n17630 DVDD.n17594 0.9005
R28827 DVDD.n17631 DVDD.n17593 0.9005
R28828 DVDD.n17632 DVDD.n17592 0.9005
R28829 DVDD.n17633 DVDD.n17591 0.9005
R28830 DVDD.n17634 DVDD.n17590 0.9005
R28831 DVDD.n17635 DVDD.n17589 0.9005
R28832 DVDD.n17636 DVDD.n17588 0.9005
R28833 DVDD.n17637 DVDD.n17587 0.9005
R28834 DVDD.n17638 DVDD.n17586 0.9005
R28835 DVDD.n17639 DVDD.n17585 0.9005
R28836 DVDD.n17640 DVDD.n17584 0.9005
R28837 DVDD.n17641 DVDD.n17583 0.9005
R28838 DVDD.n17642 DVDD.n17582 0.9005
R28839 DVDD.n17643 DVDD.n17581 0.9005
R28840 DVDD.n17644 DVDD.n17580 0.9005
R28841 DVDD.n17645 DVDD.n17579 0.9005
R28842 DVDD.n17646 DVDD.n17578 0.9005
R28843 DVDD.n17647 DVDD.n17577 0.9005
R28844 DVDD.n17648 DVDD.n17576 0.9005
R28845 DVDD.n17649 DVDD.n17575 0.9005
R28846 DVDD.n17650 DVDD.n17574 0.9005
R28847 DVDD.n17651 DVDD.n17573 0.9005
R28848 DVDD.n17652 DVDD.n17572 0.9005
R28849 DVDD.n17653 DVDD.n17571 0.9005
R28850 DVDD.n17654 DVDD.n17570 0.9005
R28851 DVDD.n17655 DVDD.n17569 0.9005
R28852 DVDD.n17656 DVDD.n17568 0.9005
R28853 DVDD.n17657 DVDD.n17567 0.9005
R28854 DVDD.n17658 DVDD.n17566 0.9005
R28855 DVDD.n17659 DVDD.n17565 0.9005
R28856 DVDD.n17660 DVDD.n17564 0.9005
R28857 DVDD.n17661 DVDD.n17563 0.9005
R28858 DVDD.n17662 DVDD.n17562 0.9005
R28859 DVDD.n17663 DVDD.n17561 0.9005
R28860 DVDD.n17664 DVDD.n17560 0.9005
R28861 DVDD.n17665 DVDD.n17559 0.9005
R28862 DVDD.n17666 DVDD.n17558 0.9005
R28863 DVDD.n17667 DVDD.n17557 0.9005
R28864 DVDD.n17668 DVDD.n17556 0.9005
R28865 DVDD.n17669 DVDD.n17555 0.9005
R28866 DVDD.n17670 DVDD.n17554 0.9005
R28867 DVDD.n17671 DVDD.n17553 0.9005
R28868 DVDD.n17672 DVDD.n17552 0.9005
R28869 DVDD.n17673 DVDD.n17551 0.9005
R28870 DVDD.n17674 DVDD.n17550 0.9005
R28871 DVDD.n17675 DVDD.n17549 0.9005
R28872 DVDD.n17676 DVDD.n17548 0.9005
R28873 DVDD.n17677 DVDD.n17547 0.9005
R28874 DVDD.n17678 DVDD.n17546 0.9005
R28875 DVDD.n17679 DVDD.n17545 0.9005
R28876 DVDD.n17680 DVDD.n17544 0.9005
R28877 DVDD.n17681 DVDD.n17543 0.9005
R28878 DVDD.n17682 DVDD.n17542 0.9005
R28879 DVDD.n17683 DVDD.n17541 0.9005
R28880 DVDD.n17684 DVDD.n17540 0.9005
R28881 DVDD.n17685 DVDD.n17539 0.9005
R28882 DVDD.n17686 DVDD.n17538 0.9005
R28883 DVDD.n17687 DVDD.n17537 0.9005
R28884 DVDD.n17688 DVDD.n17536 0.9005
R28885 DVDD.n17689 DVDD.n17535 0.9005
R28886 DVDD.n17690 DVDD.n17534 0.9005
R28887 DVDD.n17691 DVDD.n17533 0.9005
R28888 DVDD.n17692 DVDD.n17532 0.9005
R28889 DVDD.n17693 DVDD.n17531 0.9005
R28890 DVDD.n17694 DVDD.n17530 0.9005
R28891 DVDD.n17695 DVDD.n17529 0.9005
R28892 DVDD.n17696 DVDD.n17528 0.9005
R28893 DVDD.n17697 DVDD.n17527 0.9005
R28894 DVDD.n17698 DVDD.n17526 0.9005
R28895 DVDD.n17699 DVDD.n17525 0.9005
R28896 DVDD.n17700 DVDD.n17524 0.9005
R28897 DVDD.n17701 DVDD.n17523 0.9005
R28898 DVDD.n17702 DVDD.n17522 0.9005
R28899 DVDD.n17703 DVDD.n17521 0.9005
R28900 DVDD.n17704 DVDD.n17520 0.9005
R28901 DVDD.n17705 DVDD.n17519 0.9005
R28902 DVDD.n17706 DVDD.n17518 0.9005
R28903 DVDD.n17707 DVDD.n17517 0.9005
R28904 DVDD.n17708 DVDD.n17516 0.9005
R28905 DVDD.n17515 DVDD.n897 0.9005
R28906 DVDD.n17612 DVDD.n17305 0.9005
R28907 DVDD.n17612 DVDD.n17371 0.9005
R28908 DVDD.n17613 DVDD.n17360 0.9005
R28909 DVDD.n17614 DVDD.n17374 0.9005
R28910 DVDD.n17615 DVDD.n17359 0.9005
R28911 DVDD.n17616 DVDD.n17377 0.9005
R28912 DVDD.n17617 DVDD.n17358 0.9005
R28913 DVDD.n17618 DVDD.n17380 0.9005
R28914 DVDD.n17619 DVDD.n17357 0.9005
R28915 DVDD.n17620 DVDD.n17383 0.9005
R28916 DVDD.n17621 DVDD.n17356 0.9005
R28917 DVDD.n17622 DVDD.n17386 0.9005
R28918 DVDD.n17623 DVDD.n17355 0.9005
R28919 DVDD.n17624 DVDD.n17389 0.9005
R28920 DVDD.n17625 DVDD.n17354 0.9005
R28921 DVDD.n17626 DVDD.n17392 0.9005
R28922 DVDD.n17627 DVDD.n17353 0.9005
R28923 DVDD.n17628 DVDD.n17395 0.9005
R28924 DVDD.n17629 DVDD.n17352 0.9005
R28925 DVDD.n17630 DVDD.n17398 0.9005
R28926 DVDD.n17631 DVDD.n17351 0.9005
R28927 DVDD.n17632 DVDD.n17401 0.9005
R28928 DVDD.n17633 DVDD.n17350 0.9005
R28929 DVDD.n17634 DVDD.n17404 0.9005
R28930 DVDD.n17635 DVDD.n17349 0.9005
R28931 DVDD.n17636 DVDD.n17407 0.9005
R28932 DVDD.n17637 DVDD.n17348 0.9005
R28933 DVDD.n17638 DVDD.n17410 0.9005
R28934 DVDD.n17639 DVDD.n17347 0.9005
R28935 DVDD.n17640 DVDD.n17413 0.9005
R28936 DVDD.n17641 DVDD.n17346 0.9005
R28937 DVDD.n17642 DVDD.n17416 0.9005
R28938 DVDD.n17643 DVDD.n17345 0.9005
R28939 DVDD.n17644 DVDD.n17419 0.9005
R28940 DVDD.n17645 DVDD.n17344 0.9005
R28941 DVDD.n17646 DVDD.n17422 0.9005
R28942 DVDD.n17647 DVDD.n17343 0.9005
R28943 DVDD.n17648 DVDD.n17425 0.9005
R28944 DVDD.n17649 DVDD.n17342 0.9005
R28945 DVDD.n17650 DVDD.n17428 0.9005
R28946 DVDD.n17651 DVDD.n17341 0.9005
R28947 DVDD.n17652 DVDD.n17431 0.9005
R28948 DVDD.n17653 DVDD.n17340 0.9005
R28949 DVDD.n17654 DVDD.n17434 0.9005
R28950 DVDD.n17655 DVDD.n17339 0.9005
R28951 DVDD.n17656 DVDD.n17437 0.9005
R28952 DVDD.n17657 DVDD.n17338 0.9005
R28953 DVDD.n17658 DVDD.n17440 0.9005
R28954 DVDD.n17659 DVDD.n17337 0.9005
R28955 DVDD.n17660 DVDD.n17443 0.9005
R28956 DVDD.n17661 DVDD.n17336 0.9005
R28957 DVDD.n17662 DVDD.n17446 0.9005
R28958 DVDD.n17663 DVDD.n17335 0.9005
R28959 DVDD.n17664 DVDD.n17449 0.9005
R28960 DVDD.n17665 DVDD.n17334 0.9005
R28961 DVDD.n17666 DVDD.n17452 0.9005
R28962 DVDD.n17667 DVDD.n17333 0.9005
R28963 DVDD.n17668 DVDD.n17455 0.9005
R28964 DVDD.n17669 DVDD.n17332 0.9005
R28965 DVDD.n17670 DVDD.n17458 0.9005
R28966 DVDD.n17671 DVDD.n17331 0.9005
R28967 DVDD.n17672 DVDD.n17461 0.9005
R28968 DVDD.n17673 DVDD.n17330 0.9005
R28969 DVDD.n17674 DVDD.n17464 0.9005
R28970 DVDD.n17675 DVDD.n17329 0.9005
R28971 DVDD.n17676 DVDD.n17467 0.9005
R28972 DVDD.n17677 DVDD.n17328 0.9005
R28973 DVDD.n17678 DVDD.n17470 0.9005
R28974 DVDD.n17679 DVDD.n17327 0.9005
R28975 DVDD.n17680 DVDD.n17473 0.9005
R28976 DVDD.n17681 DVDD.n17326 0.9005
R28977 DVDD.n17682 DVDD.n17476 0.9005
R28978 DVDD.n17683 DVDD.n17325 0.9005
R28979 DVDD.n17684 DVDD.n17479 0.9005
R28980 DVDD.n17685 DVDD.n17324 0.9005
R28981 DVDD.n17686 DVDD.n17482 0.9005
R28982 DVDD.n17687 DVDD.n17323 0.9005
R28983 DVDD.n17688 DVDD.n17485 0.9005
R28984 DVDD.n17689 DVDD.n17322 0.9005
R28985 DVDD.n17690 DVDD.n17488 0.9005
R28986 DVDD.n17691 DVDD.n17321 0.9005
R28987 DVDD.n17692 DVDD.n17491 0.9005
R28988 DVDD.n17693 DVDD.n17320 0.9005
R28989 DVDD.n17694 DVDD.n17494 0.9005
R28990 DVDD.n17695 DVDD.n17319 0.9005
R28991 DVDD.n17696 DVDD.n17497 0.9005
R28992 DVDD.n17697 DVDD.n17318 0.9005
R28993 DVDD.n17698 DVDD.n17500 0.9005
R28994 DVDD.n17699 DVDD.n17317 0.9005
R28995 DVDD.n17700 DVDD.n17503 0.9005
R28996 DVDD.n17701 DVDD.n17316 0.9005
R28997 DVDD.n17702 DVDD.n17506 0.9005
R28998 DVDD.n17703 DVDD.n17315 0.9005
R28999 DVDD.n17704 DVDD.n17509 0.9005
R29000 DVDD.n17705 DVDD.n17314 0.9005
R29001 DVDD.n17706 DVDD.n17512 0.9005
R29002 DVDD.n17707 DVDD.n17313 0.9005
R29003 DVDD.n17709 DVDD.n17708 0.9005
R29004 DVDD.n17312 DVDD.n897 0.9005
R29005 DVDD.n17712 DVDD.n17711 0.9005
R29006 DVDD.n15126 DVDD.n5643 0.9005
R29007 DVDD.n5742 DVDD.n5641 0.9005
R29008 DVDD.n5644 DVDD.n5583 0.9005
R29009 DVDD.n15133 DVDD.n15132 0.9005
R29010 DVDD.n5645 DVDD.n5589 0.9005
R29011 DVDD.n5790 DVDD.n5640 0.9005
R29012 DVDD.n5789 DVDD.n5646 0.9005
R29013 DVDD.n5794 DVDD.n5639 0.9005
R29014 DVDD.n5795 DVDD.n5647 0.9005
R29015 DVDD.n5796 DVDD.n5638 0.9005
R29016 DVDD.n5787 DVDD.n5648 0.9005
R29017 DVDD.n5800 DVDD.n5637 0.9005
R29018 DVDD.n5801 DVDD.n5649 0.9005
R29019 DVDD.n5802 DVDD.n5636 0.9005
R29020 DVDD.n5785 DVDD.n5650 0.9005
R29021 DVDD.n5806 DVDD.n5635 0.9005
R29022 DVDD.n5807 DVDD.n5651 0.9005
R29023 DVDD.n5808 DVDD.n5634 0.9005
R29024 DVDD.n5783 DVDD.n5652 0.9005
R29025 DVDD.n5812 DVDD.n5633 0.9005
R29026 DVDD.n5813 DVDD.n5653 0.9005
R29027 DVDD.n5814 DVDD.n5632 0.9005
R29028 DVDD.n5781 DVDD.n5654 0.9005
R29029 DVDD.n5818 DVDD.n5631 0.9005
R29030 DVDD.n5819 DVDD.n5655 0.9005
R29031 DVDD.n5820 DVDD.n5630 0.9005
R29032 DVDD.n5779 DVDD.n5656 0.9005
R29033 DVDD.n5824 DVDD.n5629 0.9005
R29034 DVDD.n5825 DVDD.n5657 0.9005
R29035 DVDD.n5826 DVDD.n5628 0.9005
R29036 DVDD.n5777 DVDD.n5658 0.9005
R29037 DVDD.n5830 DVDD.n5627 0.9005
R29038 DVDD.n5831 DVDD.n5659 0.9005
R29039 DVDD.n5832 DVDD.n5626 0.9005
R29040 DVDD.n5775 DVDD.n5660 0.9005
R29041 DVDD.n5836 DVDD.n5625 0.9005
R29042 DVDD.n5837 DVDD.n5661 0.9005
R29043 DVDD.n5838 DVDD.n5624 0.9005
R29044 DVDD.n5773 DVDD.n5662 0.9005
R29045 DVDD.n5842 DVDD.n5623 0.9005
R29046 DVDD.n5843 DVDD.n5663 0.9005
R29047 DVDD.n5844 DVDD.n5622 0.9005
R29048 DVDD.n5771 DVDD.n5664 0.9005
R29049 DVDD.n5848 DVDD.n5621 0.9005
R29050 DVDD.n5849 DVDD.n5665 0.9005
R29051 DVDD.n5850 DVDD.n5620 0.9005
R29052 DVDD.n5769 DVDD.n5666 0.9005
R29053 DVDD.n5854 DVDD.n5619 0.9005
R29054 DVDD.n5855 DVDD.n5667 0.9005
R29055 DVDD.n5856 DVDD.n5618 0.9005
R29056 DVDD.n5767 DVDD.n5668 0.9005
R29057 DVDD.n5860 DVDD.n5617 0.9005
R29058 DVDD.n5861 DVDD.n5669 0.9005
R29059 DVDD.n5862 DVDD.n5616 0.9005
R29060 DVDD.n5765 DVDD.n5670 0.9005
R29061 DVDD.n5866 DVDD.n5615 0.9005
R29062 DVDD.n5867 DVDD.n5671 0.9005
R29063 DVDD.n5868 DVDD.n5614 0.9005
R29064 DVDD.n5763 DVDD.n5672 0.9005
R29065 DVDD.n5872 DVDD.n5613 0.9005
R29066 DVDD.n5873 DVDD.n5673 0.9005
R29067 DVDD.n5874 DVDD.n5612 0.9005
R29068 DVDD.n5761 DVDD.n5674 0.9005
R29069 DVDD.n5878 DVDD.n5611 0.9005
R29070 DVDD.n5879 DVDD.n5675 0.9005
R29071 DVDD.n5880 DVDD.n5610 0.9005
R29072 DVDD.n5759 DVDD.n5676 0.9005
R29073 DVDD.n5884 DVDD.n5609 0.9005
R29074 DVDD.n5885 DVDD.n5677 0.9005
R29075 DVDD.n5886 DVDD.n5608 0.9005
R29076 DVDD.n5757 DVDD.n5678 0.9005
R29077 DVDD.n5890 DVDD.n5607 0.9005
R29078 DVDD.n5891 DVDD.n5679 0.9005
R29079 DVDD.n5892 DVDD.n5606 0.9005
R29080 DVDD.n5755 DVDD.n5680 0.9005
R29081 DVDD.n5896 DVDD.n5605 0.9005
R29082 DVDD.n5897 DVDD.n5681 0.9005
R29083 DVDD.n5898 DVDD.n5604 0.9005
R29084 DVDD.n5753 DVDD.n5682 0.9005
R29085 DVDD.n5902 DVDD.n5603 0.9005
R29086 DVDD.n5903 DVDD.n5683 0.9005
R29087 DVDD.n5904 DVDD.n5602 0.9005
R29088 DVDD.n5751 DVDD.n5684 0.9005
R29089 DVDD.n5908 DVDD.n5601 0.9005
R29090 DVDD.n5909 DVDD.n5685 0.9005
R29091 DVDD.n5910 DVDD.n5600 0.9005
R29092 DVDD.n5749 DVDD.n5686 0.9005
R29093 DVDD.n5914 DVDD.n5599 0.9005
R29094 DVDD.n5915 DVDD.n5687 0.9005
R29095 DVDD.n5916 DVDD.n5598 0.9005
R29096 DVDD.n5747 DVDD.n5688 0.9005
R29097 DVDD.n5920 DVDD.n5597 0.9005
R29098 DVDD.n5921 DVDD.n5689 0.9005
R29099 DVDD.n5922 DVDD.n5596 0.9005
R29100 DVDD.n5745 DVDD.n5690 0.9005
R29101 DVDD.n5926 DVDD.n5595 0.9005
R29102 DVDD.n5927 DVDD.n5691 0.9005
R29103 DVDD.n5928 DVDD.n5594 0.9005
R29104 DVDD.n15130 DVDD.n15129 0.9005
R29105 DVDD.n15135 DVDD.n5583 0.9005
R29106 DVDD.n15134 DVDD.n15133 0.9005
R29107 DVDD.n5589 DVDD.n5588 0.9005
R29108 DVDD.n5791 DVDD.n5790 0.9005
R29109 DVDD.n5792 DVDD.n5789 0.9005
R29110 DVDD.n5794 DVDD.n5793 0.9005
R29111 DVDD.n5795 DVDD.n5788 0.9005
R29112 DVDD.n5797 DVDD.n5796 0.9005
R29113 DVDD.n5798 DVDD.n5787 0.9005
R29114 DVDD.n5800 DVDD.n5799 0.9005
R29115 DVDD.n5801 DVDD.n5786 0.9005
R29116 DVDD.n5803 DVDD.n5802 0.9005
R29117 DVDD.n5804 DVDD.n5785 0.9005
R29118 DVDD.n5806 DVDD.n5805 0.9005
R29119 DVDD.n5807 DVDD.n5784 0.9005
R29120 DVDD.n5809 DVDD.n5808 0.9005
R29121 DVDD.n5810 DVDD.n5783 0.9005
R29122 DVDD.n5812 DVDD.n5811 0.9005
R29123 DVDD.n5813 DVDD.n5782 0.9005
R29124 DVDD.n5815 DVDD.n5814 0.9005
R29125 DVDD.n5816 DVDD.n5781 0.9005
R29126 DVDD.n5818 DVDD.n5817 0.9005
R29127 DVDD.n5819 DVDD.n5780 0.9005
R29128 DVDD.n5821 DVDD.n5820 0.9005
R29129 DVDD.n5822 DVDD.n5779 0.9005
R29130 DVDD.n5824 DVDD.n5823 0.9005
R29131 DVDD.n5825 DVDD.n5778 0.9005
R29132 DVDD.n5827 DVDD.n5826 0.9005
R29133 DVDD.n5828 DVDD.n5777 0.9005
R29134 DVDD.n5830 DVDD.n5829 0.9005
R29135 DVDD.n5831 DVDD.n5776 0.9005
R29136 DVDD.n5833 DVDD.n5832 0.9005
R29137 DVDD.n5834 DVDD.n5775 0.9005
R29138 DVDD.n5836 DVDD.n5835 0.9005
R29139 DVDD.n5837 DVDD.n5774 0.9005
R29140 DVDD.n5839 DVDD.n5838 0.9005
R29141 DVDD.n5840 DVDD.n5773 0.9005
R29142 DVDD.n5842 DVDD.n5841 0.9005
R29143 DVDD.n5843 DVDD.n5772 0.9005
R29144 DVDD.n5845 DVDD.n5844 0.9005
R29145 DVDD.n5846 DVDD.n5771 0.9005
R29146 DVDD.n5848 DVDD.n5847 0.9005
R29147 DVDD.n5849 DVDD.n5770 0.9005
R29148 DVDD.n5851 DVDD.n5850 0.9005
R29149 DVDD.n5852 DVDD.n5769 0.9005
R29150 DVDD.n5854 DVDD.n5853 0.9005
R29151 DVDD.n5855 DVDD.n5768 0.9005
R29152 DVDD.n5857 DVDD.n5856 0.9005
R29153 DVDD.n5858 DVDD.n5767 0.9005
R29154 DVDD.n5860 DVDD.n5859 0.9005
R29155 DVDD.n5861 DVDD.n5766 0.9005
R29156 DVDD.n5863 DVDD.n5862 0.9005
R29157 DVDD.n5864 DVDD.n5765 0.9005
R29158 DVDD.n5866 DVDD.n5865 0.9005
R29159 DVDD.n5867 DVDD.n5764 0.9005
R29160 DVDD.n5869 DVDD.n5868 0.9005
R29161 DVDD.n5870 DVDD.n5763 0.9005
R29162 DVDD.n5872 DVDD.n5871 0.9005
R29163 DVDD.n5873 DVDD.n5762 0.9005
R29164 DVDD.n5875 DVDD.n5874 0.9005
R29165 DVDD.n5876 DVDD.n5761 0.9005
R29166 DVDD.n5878 DVDD.n5877 0.9005
R29167 DVDD.n5879 DVDD.n5760 0.9005
R29168 DVDD.n5881 DVDD.n5880 0.9005
R29169 DVDD.n5882 DVDD.n5759 0.9005
R29170 DVDD.n5884 DVDD.n5883 0.9005
R29171 DVDD.n5885 DVDD.n5758 0.9005
R29172 DVDD.n5887 DVDD.n5886 0.9005
R29173 DVDD.n5888 DVDD.n5757 0.9005
R29174 DVDD.n5890 DVDD.n5889 0.9005
R29175 DVDD.n5891 DVDD.n5756 0.9005
R29176 DVDD.n5893 DVDD.n5892 0.9005
R29177 DVDD.n5894 DVDD.n5755 0.9005
R29178 DVDD.n5896 DVDD.n5895 0.9005
R29179 DVDD.n5897 DVDD.n5754 0.9005
R29180 DVDD.n5899 DVDD.n5898 0.9005
R29181 DVDD.n5900 DVDD.n5753 0.9005
R29182 DVDD.n5902 DVDD.n5901 0.9005
R29183 DVDD.n5903 DVDD.n5752 0.9005
R29184 DVDD.n5905 DVDD.n5904 0.9005
R29185 DVDD.n5906 DVDD.n5751 0.9005
R29186 DVDD.n5908 DVDD.n5907 0.9005
R29187 DVDD.n5909 DVDD.n5750 0.9005
R29188 DVDD.n5911 DVDD.n5910 0.9005
R29189 DVDD.n5912 DVDD.n5749 0.9005
R29190 DVDD.n5914 DVDD.n5913 0.9005
R29191 DVDD.n5915 DVDD.n5748 0.9005
R29192 DVDD.n5917 DVDD.n5916 0.9005
R29193 DVDD.n5918 DVDD.n5747 0.9005
R29194 DVDD.n5920 DVDD.n5919 0.9005
R29195 DVDD.n5921 DVDD.n5746 0.9005
R29196 DVDD.n5923 DVDD.n5922 0.9005
R29197 DVDD.n5924 DVDD.n5745 0.9005
R29198 DVDD.n5926 DVDD.n5925 0.9005
R29199 DVDD.n5927 DVDD.n5744 0.9005
R29200 DVDD.n5929 DVDD.n5928 0.9005
R29201 DVDD.n5930 DVDD.n5742 0.9005
R29202 DVDD.n15129 DVDD.n15128 0.9005
R29203 DVDD.n4335 DVDD.t35 0.896055
R29204 DVDD.n4370 DVDD.t55 0.896055
R29205 DVDD.n4350 DVDD.t1 0.896055
R29206 DVDD.n21971 DVDD.n21969 0.769795
R29207 DVDD.n21698 DVDD.n21697 0.769795
R29208 DVDD.n21824 DVDD.n21822 0.769795
R29209 DVDD.n18418 DVDD.n18412 0.769795
R29210 DVDD.n22019 DVDD.n22018 0.769684
R29211 DVDD.n21242 DVDD.n21218 0.769684
R29212 DVDD.n21349 DVDD.n21348 0.769684
R29213 DVDD.n21956 DVDD.n21955 0.769684
R29214 DVDD.n18259 DVDD.n18258 0.769684
R29215 DVDD.n21853 DVDD.n21852 0.769684
R29216 DVDD.n18472 DVDD.n18470 0.769684
R29217 DVDD.n18443 DVDD.n18442 0.769684
R29218 DVDD.n4294 DVDD.n4285 0.769684
R29219 DVDD.n4310 DVDD.n4301 0.769684
R29220 DVDD.n3687 DVDD.n3686 0.769684
R29221 DVDD.n3703 DVDD.n3702 0.769684
R29222 DVDD.n21929 DVDD.n21792 0.763137
R29223 DVDD.n21771 DVDD.n21770 0.762368
R29224 DVDD.n22238 DVDD.n130 0.760008
R29225 DVDD.n21936 DVDD.n21784 0.760008
R29226 DVDD.n18103 DVDD.n18099 0.760008
R29227 DVDD.n18124 DVDD.n18064 0.759948
R29228 DVDD.n21732 DVDD.n21731 0.75924
R29229 DVDD.n22068 DVDD.n22067 0.75924
R29230 DVDD.n18096 DVDD.n499 0.750711
R29231 DVDD.n18430 DVDD.n18429 0.7505
R29232 DVDD.n21723 DVDD.n155 0.7505
R29233 DVDD.n22231 DVDD.n22230 0.7505
R29234 DVDD.n18478 DVDD.n132 0.7505
R29235 DVDD.n22235 DVDD.n133 0.7505
R29236 DVDD.n22237 DVDD.n22236 0.7505
R29237 DVDD.n21725 DVDD.n21724 0.7505
R29238 DVDD.n21729 DVDD.n21728 0.7505
R29239 DVDD.n21730 DVDD.n21729 0.7505
R29240 DVDD.n21724 DVDD.n18431 0.7505
R29241 DVDD.n21723 DVDD.n21722 0.7505
R29242 DVDD.n22232 DVDD.n22231 0.7505
R29243 DVDD.n22233 DVDD.n132 0.7505
R29244 DVDD.n22235 DVDD.n22234 0.7505
R29245 DVDD.n21928 DVDD.n21927 0.7505
R29246 DVDD.n21926 DVDD.n21795 0.7505
R29247 DVDD.n21796 DVDD.n21794 0.7505
R29248 DVDD.n21922 DVDD.n21921 0.7505
R29249 DVDD.n22041 DVDD.n22040 0.7505
R29250 DVDD.n22042 DVDD.n18209 0.7505
R29251 DVDD.n22065 DVDD.n22064 0.7505
R29252 DVDD.n18211 DVDD.n18207 0.7505
R29253 DVDD.n21926 DVDD.n21925 0.7505
R29254 DVDD.n21924 DVDD.n21794 0.7505
R29255 DVDD.n21923 DVDD.n21922 0.7505
R29256 DVDD.n22040 DVDD.n213 0.7505
R29257 DVDD.n18209 DVDD.n18208 0.7505
R29258 DVDD.n22066 DVDD.n22065 0.7505
R29259 DVDD.n21764 DVDD.n18390 0.7505
R29260 DVDD.n21765 DVDD.n18389 0.7505
R29261 DVDD.n21776 DVDD.n21775 0.7505
R29262 DVDD.n18297 DVDD.n180 0.7505
R29263 DVDD.n18385 DVDD.n179 0.7505
R29264 DVDD.n21940 DVDD.n21939 0.7505
R29265 DVDD.n21785 DVDD.n21782 0.7505
R29266 DVDD.n21935 DVDD.n21934 0.7505
R29267 DVDD.n21772 DVDD.n18389 0.7505
R29268 DVDD.n21775 DVDD.n21774 0.7505
R29269 DVDD.n21773 DVDD.n180 0.7505
R29270 DVDD.n21783 DVDD.n179 0.7505
R29271 DVDD.n21939 DVDD.n21938 0.7505
R29272 DVDD.n21937 DVDD.n21782 0.7505
R29273 DVDD.n18122 DVDD.n18121 0.7505
R29274 DVDD.n18120 DVDD.n18067 0.7505
R29275 DVDD.n18094 DVDD.n18066 0.7505
R29276 DVDD.n18116 DVDD.n18115 0.7505
R29277 DVDD.n18113 DVDD.n18112 0.7505
R29278 DVDD.n18101 DVDD.n18098 0.7505
R29279 DVDD.n18108 DVDD.n18107 0.7505
R29280 DVDD.n18104 DVDD.n18100 0.7505
R29281 DVDD.n18120 DVDD.n18119 0.7505
R29282 DVDD.n18118 DVDD.n18066 0.7505
R29283 DVDD.n18117 DVDD.n18116 0.7505
R29284 DVDD.n18112 DVDD.n18111 0.7505
R29285 DVDD.n18110 DVDD.n18098 0.7505
R29286 DVDD.n18109 DVDD.n18108 0.7505
R29287 DVDD.n17725 DVDD.n898 0.7505
R29288 DVDD.n17362 DVDD.n891 0.7505
R29289 DVDD.n17361 DVDD.n894 0.7505
R29290 DVDD.n17368 DVDD.n892 0.7505
R29291 DVDD.n15140 DVDD.n5584 0.7505
R29292 DVDD.n5992 DVDD.n5578 0.7505
R29293 DVDD.n5936 DVDD.n5580 0.7505
R29294 DVDD.n5990 DVDD.n5587 0.7505
R29295 DVDD.n19895 DVDD.n19823 0.643357
R29296 DVDD.n19896 DVDD.n19894 0.643357
R29297 DVDD.n19898 DVDD.n19897 0.643357
R29298 DVDD.n19899 DVDD.n19893 0.643357
R29299 DVDD.n19901 DVDD.n19900 0.643357
R29300 DVDD.n19902 DVDD.n19892 0.643357
R29301 DVDD.n19904 DVDD.n19903 0.643357
R29302 DVDD.n19905 DVDD.n19884 0.643357
R29303 DVDD.n19935 DVDD.n19934 0.643357
R29304 DVDD.n19933 DVDD.n19932 0.643357
R29305 DVDD.n19931 DVDD.n19930 0.643357
R29306 DVDD.n19929 DVDD.n19928 0.643357
R29307 DVDD.n19927 DVDD.n19926 0.643357
R29308 DVDD.n19925 DVDD.n19924 0.643357
R29309 DVDD.n19923 DVDD.n19922 0.643357
R29310 DVDD.n19921 DVDD.n19920 0.643357
R29311 DVDD.n19919 DVDD.n19918 0.643357
R29312 DVDD.n19917 DVDD.n19916 0.643357
R29313 DVDD.n19915 DVDD.n19914 0.643357
R29314 DVDD.n19913 DVDD.n19906 0.643357
R29315 DVDD.n19912 DVDD.n19911 0.643357
R29316 DVDD.n19910 DVDD.n19907 0.643357
R29317 DVDD.n19909 DVDD.n19908 0.643357
R29318 DVDD.n19822 DVDD.n19821 0.643357
R29319 DVDD.n20441 DVDD.n20440 0.643357
R29320 DVDD.n20542 DVDD.n20541 0.643357
R29321 DVDD.n19766 DVDD.n19765 0.643357
R29322 DVDD.n19996 DVDD.n19995 0.643357
R29323 DVDD.n19997 DVDD.n19994 0.643357
R29324 DVDD.n19999 DVDD.n19998 0.643357
R29325 DVDD.n20000 DVDD.n19993 0.643357
R29326 DVDD.n20002 DVDD.n20001 0.643357
R29327 DVDD.n20004 DVDD.n20003 0.643357
R29328 DVDD.n20006 DVDD.n20005 0.643357
R29329 DVDD.n20008 DVDD.n20007 0.643357
R29330 DVDD.n20010 DVDD.n20009 0.643357
R29331 DVDD.n20012 DVDD.n20011 0.643357
R29332 DVDD.n20014 DVDD.n20013 0.643357
R29333 DVDD.n20016 DVDD.n20015 0.643357
R29334 DVDD.n20018 DVDD.n20017 0.643357
R29335 DVDD.n20020 DVDD.n20019 0.643357
R29336 DVDD.n20022 DVDD.n20021 0.643357
R29337 DVDD.n19992 DVDD.n19969 0.643357
R29338 DVDD.n19991 DVDD.n19990 0.643357
R29339 DVDD.n19989 DVDD.n19978 0.643357
R29340 DVDD.n19988 DVDD.n19987 0.643357
R29341 DVDD.n19986 DVDD.n19979 0.643357
R29342 DVDD.n19985 DVDD.n19984 0.643357
R29343 DVDD.n19983 DVDD.n19980 0.643357
R29344 DVDD.n19982 DVDD.n19981 0.643357
R29345 DVDD.n4373 DVDD.n4370 0.625181
R29346 DVDD.n4350 DVDD.n4339 0.625181
R29347 DVDD.n4344 DVDD.n4335 0.625181
R29348 DVDD.n4343 DVDD.n4337 0.625075
R29349 DVDD.n4338 DVDD.n4334 0.625075
R29350 DVDD.n4384 DVDD.n4382 0.625075
R29351 DVDD.n4380 DVDD.n4357 0.625075
R29352 DVDD.n4379 DVDD.n4359 0.625075
R29353 DVDD.n4378 DVDD.n4361 0.625075
R29354 DVDD.n4377 DVDD.n4364 0.625075
R29355 DVDD.n4375 DVDD.n4367 0.625075
R29356 DVDD.n4374 DVDD.n4369 0.625075
R29357 DVDD.n4349 DVDD.n4347 0.625075
R29358 DVDD.n4346 DVDD.n4341 0.625075
R29359 DVDD.n20595 DVDD 0.612796
R29360 DVDD DVDD.n19710 0.612796
R29361 DVDD DVDD.n20594 0.612796
R29362 DVDD DVDD.n19711 0.612796
R29363 DVDD.n20592 DVDD 0.612796
R29364 DVDD.n19981 DVDD 0.612796
R29365 DVDD.n20543 DVDD 0.612796
R29366 DVDD DVDD.n20542 0.612796
R29367 DVDD.n20899 DVDD 0.612796
R29368 DVDD DVDD.n18922 0.612796
R29369 DVDD DVDD.n20898 0.612796
R29370 DVDD DVDD.n18923 0.612796
R29371 DVDD.n20440 DVDD 0.612796
R29372 DVDD DVDD.n18920 0.612796
R29373 DVDD DVDD.n20439 0.612796
R29374 DVDD DVDD.n19823 0.612796
R29375 DVDD.n19394 DVDD.t68 0.58122
R29376 DVDD.t12 DVDD.n18631 0.58122
R29377 DVDD.n19097 DVDD.n18819 0.565091
R29378 DVDD.n20926 DVDD.n18906 0.565091
R29379 DVDD.n19101 DVDD.n19097 0.564924
R29380 DVDD.n20923 DVDD.n18906 0.564924
R29381 DVDD.n20438 DVDD.n18923 0.563
R29382 DVDD.n20437 DVDD.n20436 0.563
R29383 DVDD.n20435 DVDD.n19825 0.563
R29384 DVDD.n20434 DVDD.n20433 0.563
R29385 DVDD.n19827 DVDD.n19826 0.563
R29386 DVDD.n20429 DVDD.n20428 0.563
R29387 DVDD.n20427 DVDD.n19830 0.563
R29388 DVDD.n20426 DVDD.n20425 0.563
R29389 DVDD.n20422 DVDD.n19831 0.563
R29390 DVDD.n20379 DVDD.n19842 0.563
R29391 DVDD.n20418 DVDD.n20417 0.563
R29392 DVDD.n20416 DVDD.n20415 0.563
R29393 DVDD.n20412 DVDD.n20380 0.563
R29394 DVDD.n20410 DVDD.n20409 0.563
R29395 DVDD.n20408 DVDD.n20407 0.563
R29396 DVDD.n20406 DVDD.n20405 0.563
R29397 DVDD.n20402 DVDD.n20382 0.563
R29398 DVDD.n20400 DVDD.n20399 0.563
R29399 DVDD.n20398 DVDD.n20397 0.563
R29400 DVDD.n20396 DVDD.n20384 0.563
R29401 DVDD.n20389 DVDD.n20385 0.563
R29402 DVDD.n20392 DVDD.n20391 0.563
R29403 DVDD.n20390 DVDD.n20388 0.563
R29404 DVDD.n18921 DVDD.n18919 0.563
R29405 DVDD.n20900 DVDD.n20899 0.563
R29406 DVDD.n20081 DVDD.n19711 0.563
R29407 DVDD.n20082 DVDD.n20080 0.563
R29408 DVDD.n20084 DVDD.n20083 0.563
R29409 DVDD.n20085 DVDD.n20079 0.563
R29410 DVDD.n20087 DVDD.n20086 0.563
R29411 DVDD.n20088 DVDD.n20078 0.563
R29412 DVDD.n20090 DVDD.n20089 0.563
R29413 DVDD.n20091 DVDD.n20070 0.563
R29414 DVDD.n20121 DVDD.n20120 0.563
R29415 DVDD.n20119 DVDD.n20118 0.563
R29416 DVDD.n20117 DVDD.n20116 0.563
R29417 DVDD.n20115 DVDD.n20114 0.563
R29418 DVDD.n20113 DVDD.n20112 0.563
R29419 DVDD.n20111 DVDD.n20110 0.563
R29420 DVDD.n20109 DVDD.n20108 0.563
R29421 DVDD.n20107 DVDD.n20106 0.563
R29422 DVDD.n20105 DVDD.n20104 0.563
R29423 DVDD.n20103 DVDD.n20102 0.563
R29424 DVDD.n20101 DVDD.n20100 0.563
R29425 DVDD.n20099 DVDD.n20092 0.563
R29426 DVDD.n20098 DVDD.n20097 0.563
R29427 DVDD.n20096 DVDD.n20093 0.563
R29428 DVDD.n20095 DVDD.n20094 0.563
R29429 DVDD.n19709 DVDD.n19708 0.563
R29430 DVDD.n20596 DVDD.n20595 0.563
R29431 DVDD.n20856 DVDD.n18922 0.563
R29432 DVDD.n20857 DVDD.n18959 0.563
R29433 DVDD.n20859 DVDD.n20858 0.563
R29434 DVDD.n20860 DVDD.n18958 0.563
R29435 DVDD.n20862 DVDD.n20861 0.563
R29436 DVDD.n20863 DVDD.n18957 0.563
R29437 DVDD.n20865 DVDD.n20864 0.563
R29438 DVDD.n20867 DVDD.n20866 0.563
R29439 DVDD.n20869 DVDD.n20868 0.563
R29440 DVDD.n20871 DVDD.n20870 0.563
R29441 DVDD.n20873 DVDD.n20872 0.563
R29442 DVDD.n20875 DVDD.n20874 0.563
R29443 DVDD.n20877 DVDD.n20876 0.563
R29444 DVDD.n20879 DVDD.n20878 0.563
R29445 DVDD.n20881 DVDD.n20880 0.563
R29446 DVDD.n18937 DVDD.n18928 0.563
R29447 DVDD.n20886 DVDD.n20885 0.563
R29448 DVDD.n20887 DVDD.n18927 0.563
R29449 DVDD.n20889 DVDD.n20888 0.563
R29450 DVDD.n20890 DVDD.n18926 0.563
R29451 DVDD.n20892 DVDD.n20891 0.563
R29452 DVDD.n20893 DVDD.n18925 0.563
R29453 DVDD.n20895 DVDD.n20894 0.563
R29454 DVDD.n20896 DVDD.n18924 0.563
R29455 DVDD.n20898 DVDD.n20897 0.563
R29456 DVDD.n19764 DVDD.n19710 0.563
R29457 DVDD.n20546 DVDD.n20545 0.563
R29458 DVDD.n20547 DVDD.n19762 0.563
R29459 DVDD.n20549 DVDD.n20548 0.563
R29460 DVDD.n19763 DVDD.n19760 0.563
R29461 DVDD.n20553 DVDD.n19759 0.563
R29462 DVDD.n20555 DVDD.n20554 0.563
R29463 DVDD.n20557 DVDD.n20556 0.563
R29464 DVDD.n20559 DVDD.n19757 0.563
R29465 DVDD.n20563 DVDD.n20562 0.563
R29466 DVDD.n20565 DVDD.n20564 0.563
R29467 DVDD.n20567 DVDD.n20566 0.563
R29468 DVDD.n20570 DVDD.n19754 0.563
R29469 DVDD.n19753 DVDD.n19751 0.563
R29470 DVDD.n19752 DVDD.n19732 0.563
R29471 DVDD.n20574 DVDD.n19720 0.563
R29472 DVDD.n20578 DVDD.n20577 0.563
R29473 DVDD.n20579 DVDD.n19719 0.563
R29474 DVDD.n20581 DVDD.n20580 0.563
R29475 DVDD.n19717 DVDD.n19716 0.563
R29476 DVDD.n20586 DVDD.n20585 0.563
R29477 DVDD.n20587 DVDD.n19715 0.563
R29478 DVDD.n20589 DVDD.n20588 0.563
R29479 DVDD.n19713 DVDD.n19712 0.563
R29480 DVDD.n20594 DVDD.n20593 0.563
R29481 DVDD.n4343 DVDD.n4338 0.545794
R29482 DVDD.n4382 DVDD.n4338 0.545794
R29483 DVDD.n4382 DVDD.n4381 0.545794
R29484 DVDD.n4381 DVDD.n4380 0.545794
R29485 DVDD.n4380 DVDD.n4379 0.545794
R29486 DVDD.n4379 DVDD.n4378 0.545794
R29487 DVDD.n4378 DVDD.n4377 0.545794
R29488 DVDD.n4377 DVDD.n4376 0.545794
R29489 DVDD.n4376 DVDD.n4375 0.545794
R29490 DVDD.n4375 DVDD.n4374 0.545794
R29491 DVDD.n4374 DVDD.n4373 0.545794
R29492 DVDD.n4347 DVDD.n4339 0.545794
R29493 DVDD.n4347 DVDD.n4346 0.545794
R29494 DVDD.n4346 DVDD.n4345 0.545794
R29495 DVDD.n4344 DVDD.n4343 0.545794
R29496 DVDD.n21014 DVDD.n18822 0.542701
R29497 DVDD.n21014 DVDD.n21013 0.542701
R29498 DVDD.n21018 DVDD.n18820 0.542701
R29499 DVDD.n21019 DVDD.n21018 0.542701
R29500 DVDD.n4337 DVDD.n4336 0.532176
R29501 DVDD.n4334 DVDD.n4333 0.532176
R29502 DVDD.n4384 DVDD.n4383 0.532176
R29503 DVDD.n4357 DVDD.n4356 0.532176
R29504 DVDD.n4359 DVDD.n4358 0.532176
R29505 DVDD.n4361 DVDD.n4360 0.532176
R29506 DVDD.n4364 DVDD.n4363 0.532176
R29507 DVDD.n4367 DVDD.n4366 0.532176
R29508 DVDD.n4369 DVDD.n4368 0.532176
R29509 DVDD.n4349 DVDD.n4348 0.532176
R29510 DVDD.n4341 DVDD.n4340 0.532176
R29511 DVDD.n18205 DVDD.n366 0.5005
R29512 DVDD.n22059 DVDD.n22058 0.5005
R29513 DVDD.n22061 DVDD.n22060 0.5005
R29514 DVDD.n18231 DVDD.n18215 0.5005
R29515 DVDD.n22046 DVDD.n22045 0.5005
R29516 DVDD.n21918 DVDD.n21917 0.5005
R29517 DVDD.n21830 DVDD.n21800 0.5005
R29518 DVDD.n21898 DVDD.n21828 0.5005
R29519 DVDD.n21900 DVDD.n21899 0.5005
R29520 DVDD.n21901 DVDD.n21790 0.5005
R29521 DVDD.n21811 DVDD.n21789 0.5005
R29522 DVDD.n21875 DVDD.n21788 0.5005
R29523 DVDD.n21877 DVDD.n21876 0.5005
R29524 DVDD.n21879 DVDD.n21878 0.5005
R29525 DVDD.n21839 DVDD.n21779 0.5005
R29526 DVDD.n21759 DVDD.n18387 0.5005
R29527 DVDD.n21761 DVDD.n21760 0.5005
R29528 DVDD.n21763 DVDD.n21762 0.5005
R29529 DVDD.n18396 DVDD.n18394 0.5005
R29530 DVDD.n18424 DVDD.n18393 0.5005
R29531 DVDD.n21737 DVDD.n21736 0.5005
R29532 DVDD.n21735 DVDD.n18426 0.5005
R29533 DVDD.n166 DVDD.n165 0.5005
R29534 DVDD.n22224 DVDD.n22223 0.5005
R29535 DVDD.n22226 DVDD.n22225 0.5005
R29536 DVDD.n18498 DVDD.n18497 0.5005
R29537 DVDD.n18458 DVDD.n18457 0.5005
R29538 DVDD.n18484 DVDD.n18483 0.5005
R29539 DVDD.n18476 DVDD.n125 0.5005
R29540 DVDD.n22241 DVDD.n22240 0.5005
R29541 DVDD.n18614 DVDD.n18428 0.5005
R29542 DVDD.n22186 DVDD.n22185 0.5005
R29543 DVDD.n230 DVDD.n228 0.5005
R29544 DVDD.n22023 DVDD.n22009 0.5005
R29545 DVDD.n21989 DVDD.n21984 0.5005
R29546 DVDD.n22037 DVDD.n21983 0.5005
R29547 DVDD.n21982 DVDD.n18267 0.5005
R29548 DVDD.n18351 DVDD.n18266 0.5005
R29549 DVDD.n21975 DVDD.n18272 0.5005
R29550 DVDD.n18339 DVDD.n18271 0.5005
R29551 DVDD.n21967 DVDD.n18281 0.5005
R29552 DVDD.n18363 DVDD.n18280 0.5005
R29553 DVDD.n21960 DVDD.n18286 0.5005
R29554 DVDD.n18323 DVDD.n18285 0.5005
R29555 DVDD.n21950 DVDD.n18294 0.5005
R29556 DVDD.n18376 DVDD.n18293 0.5005
R29557 DVDD.n21704 DVDD.n18520 0.5005
R29558 DVDD.n21670 DVDD.n18519 0.5005
R29559 DVDD.n21693 DVDD.n18527 0.5005
R29560 DVDD.n18532 DVDD.n18526 0.5005
R29561 DVDD.n21686 DVDD.n21685 0.5005
R29562 DVDD.n21331 DVDD.n18530 0.5005
R29563 DVDD.n21332 DVDD.n18552 0.5005
R29564 DVDD.n21654 DVDD.n21653 0.5005
R29565 DVDD.n18551 DVDD.n18548 0.5005
R29566 DVDD.n21357 DVDD.n21356 0.5005
R29567 DVDD.n21259 DVDD.n21258 0.5005
R29568 DVDD.n21223 DVDD.n18662 0.5005
R29569 DVDD.n21234 DVDD.n21233 0.5005
R29570 DVDD.n21220 DVDD.n21217 0.5005
R29571 DVDD.n21247 DVDD.n18655 0.5005
R29572 DVDD.n4385 DVDD.n4337 0.475882
R29573 DVDD.n4385 DVDD.n4334 0.475882
R29574 DVDD.n4385 DVDD.n4384 0.475882
R29575 DVDD.n4362 DVDD.n4357 0.475882
R29576 DVDD.n4362 DVDD.n4359 0.475882
R29577 DVDD.n4362 DVDD.n4361 0.475882
R29578 DVDD.n4364 DVDD.n4362 0.475882
R29579 DVDD.n4371 DVDD.n4367 0.475882
R29580 DVDD.n4371 DVDD.n4369 0.475882
R29581 DVDD.n4351 DVDD.n4349 0.475882
R29582 DVDD.n4351 DVDD.n4341 0.475882
R29583 DVDD.n4371 DVDD.n4370 0.475785
R29584 DVDD.n4351 DVDD.n4350 0.475785
R29585 DVDD.n4385 DVDD.n4335 0.475785
R29586 DVDD.n18345 DVDD.n18344 0.459715
R29587 DVDD.n4848 DVDD.n4847 0.459715
R29588 DVDD.n21678 DVDD.n18535 0.459655
R29589 DVDD.n18370 DVDD.n18369 0.459655
R29590 DVDD.n22004 DVDD.n22003 0.459655
R29591 DVDD.n21266 DVDD.n18656 0.459655
R29592 DVDD.n21366 DVDD.n21365 0.459655
R29593 DVDD.n4878 DVDD.n4877 0.459655
R29594 DVDD.n19104 DVDD.n19102 0.452883
R29595 DVDD.n20932 DVDD.n18870 0.452883
R29596 DVDD.n20974 DVDD.n20973 0.452883
R29597 DVDD.n20968 DVDD.n20967 0.452883
R29598 DVDD.n19104 DVDD.n19103 0.452744
R29599 DVDD.n20932 DVDD.n20931 0.452744
R29600 DVDD.n20973 DVDD.n20972 0.452744
R29601 DVDD.n20967 DVDD.n18860 0.452744
R29602 DVDD.n20338 DVDD.n20336 0.4505
R29603 DVDD.n20341 DVDD.n20340 0.4505
R29604 DVDD.n20342 DVDD.n20334 0.4505
R29605 DVDD.n20345 DVDD.n20343 0.4505
R29606 DVDD.n20347 DVDD.n20332 0.4505
R29607 DVDD.n20350 DVDD.n20349 0.4505
R29608 DVDD.n20351 DVDD.n20331 0.4505
R29609 DVDD.n20354 DVDD.n20352 0.4505
R29610 DVDD.n20356 DVDD.n20329 0.4505
R29611 DVDD.n20359 DVDD.n20358 0.4505
R29612 DVDD.n20360 DVDD.n20328 0.4505
R29613 DVDD.n20362 DVDD.n20361 0.4505
R29614 DVDD.n20326 DVDD.n20325 0.4505
R29615 DVDD.n20367 DVDD.n20366 0.4505
R29616 DVDD.n20368 DVDD.n19857 0.4505
R29617 DVDD.n20370 DVDD.n20369 0.4505
R29618 DVDD.n20324 DVDD.n19856 0.4505
R29619 DVDD.n20323 DVDD.n20322 0.4505
R29620 DVDD.n20320 DVDD.n19858 0.4505
R29621 DVDD.n20318 DVDD.n20316 0.4505
R29622 DVDD.n20315 DVDD.n19860 0.4505
R29623 DVDD.n20314 DVDD.n20313 0.4505
R29624 DVDD.n20311 DVDD.n19861 0.4505
R29625 DVDD.n20309 DVDD.n20307 0.4505
R29626 DVDD.n20306 DVDD.n19863 0.4505
R29627 DVDD.n20305 DVDD.n20304 0.4505
R29628 DVDD.n20302 DVDD.n19864 0.4505
R29629 DVDD.n20300 DVDD.n20298 0.4505
R29630 DVDD.n20297 DVDD.n19866 0.4505
R29631 DVDD.n20296 DVDD.n20295 0.4505
R29632 DVDD.n19868 DVDD.n19867 0.4505
R29633 DVDD.n20291 DVDD.n20290 0.4505
R29634 DVDD.n20289 DVDD.n19870 0.4505
R29635 DVDD.n20288 DVDD.n20287 0.4505
R29636 DVDD.n19872 DVDD.n19871 0.4505
R29637 DVDD.n20280 DVDD.n20279 0.4505
R29638 DVDD.n20278 DVDD.n19945 0.4505
R29639 DVDD.n20277 DVDD.n20276 0.4505
R29640 DVDD.n20274 DVDD.n19946 0.4505
R29641 DVDD.n20272 DVDD.n20270 0.4505
R29642 DVDD.n20269 DVDD.n19948 0.4505
R29643 DVDD.n20268 DVDD.n20267 0.4505
R29644 DVDD.n20265 DVDD.n19949 0.4505
R29645 DVDD.n20263 DVDD.n20261 0.4505
R29646 DVDD.n20260 DVDD.n19951 0.4505
R29647 DVDD.n20259 DVDD.n20258 0.4505
R29648 DVDD.n20256 DVDD.n19952 0.4505
R29649 DVDD.n20250 DVDD.n19953 0.4505
R29650 DVDD.n20252 DVDD.n20251 0.4505
R29651 DVDD.n20249 DVDD.n19955 0.4505
R29652 DVDD.n20248 DVDD.n20247 0.4505
R29653 DVDD.n19957 DVDD.n19956 0.4505
R29654 DVDD.n20238 DVDD.n20033 0.4505
R29655 DVDD.n20240 DVDD.n20239 0.4505
R29656 DVDD.n20237 DVDD.n20032 0.4505
R29657 DVDD.n20236 DVDD.n20235 0.4505
R29658 DVDD.n20233 DVDD.n20034 0.4505
R29659 DVDD.n20231 DVDD.n20229 0.4505
R29660 DVDD.n20228 DVDD.n20036 0.4505
R29661 DVDD.n20227 DVDD.n20226 0.4505
R29662 DVDD.n20224 DVDD.n20037 0.4505
R29663 DVDD.n20222 DVDD.n20220 0.4505
R29664 DVDD.n20219 DVDD.n20039 0.4505
R29665 DVDD.n20218 DVDD.n20217 0.4505
R29666 DVDD.n20215 DVDD.n20040 0.4505
R29667 DVDD.n20213 DVDD.n20042 0.4505
R29668 DVDD.n20207 DVDD.n20041 0.4505
R29669 DVDD.n20209 DVDD.n20208 0.4505
R29670 DVDD.n20206 DVDD.n20043 0.4505
R29671 DVDD.n20205 DVDD.n20204 0.4505
R29672 DVDD.n20203 DVDD.n20044 0.4505
R29673 DVDD.n20201 DVDD.n20199 0.4505
R29674 DVDD.n20198 DVDD.n20046 0.4505
R29675 DVDD.n20197 DVDD.n20196 0.4505
R29676 DVDD.n20194 DVDD.n20047 0.4505
R29677 DVDD.n20192 DVDD.n20190 0.4505
R29678 DVDD.n20189 DVDD.n20049 0.4505
R29679 DVDD.n20188 DVDD.n20187 0.4505
R29680 DVDD.n20185 DVDD.n20050 0.4505
R29681 DVDD.n20183 DVDD.n20181 0.4505
R29682 DVDD.n20180 DVDD.n20052 0.4505
R29683 DVDD.n20179 DVDD.n20178 0.4505
R29684 DVDD.n20176 DVDD.n20053 0.4505
R29685 DVDD.n20170 DVDD.n20054 0.4505
R29686 DVDD.n20172 DVDD.n20171 0.4505
R29687 DVDD.n20169 DVDD.n20056 0.4505
R29688 DVDD.n20168 DVDD.n20167 0.4505
R29689 DVDD.n20058 DVDD.n20057 0.4505
R29690 DVDD.n20141 DVDD.n20137 0.4505
R29691 DVDD.n20144 DVDD.n20142 0.4505
R29692 DVDD.n20146 DVDD.n20135 0.4505
R29693 DVDD.n20149 DVDD.n20148 0.4505
R29694 DVDD.n20150 DVDD.n20134 0.4505
R29695 DVDD.n20153 DVDD.n20151 0.4505
R29696 DVDD.n20155 DVDD.n20132 0.4505
R29697 DVDD.n20158 DVDD.n20157 0.4505
R29698 DVDD.n20159 DVDD.n20131 0.4505
R29699 DVDD.n20161 DVDD.n20160 0.4505
R29700 DVDD.n20335 DVDD.n18945 0.4505
R29701 DVDD.n20338 DVDD.n20337 0.4505
R29702 DVDD.n20340 DVDD.n20339 0.4505
R29703 DVDD.n20334 DVDD.n20333 0.4505
R29704 DVDD.n20345 DVDD.n20344 0.4505
R29705 DVDD.n20347 DVDD.n20346 0.4505
R29706 DVDD.n20349 DVDD.n20348 0.4505
R29707 DVDD.n20331 DVDD.n20330 0.4505
R29708 DVDD.n20354 DVDD.n20353 0.4505
R29709 DVDD.n20356 DVDD.n20355 0.4505
R29710 DVDD.n20358 DVDD.n20357 0.4505
R29711 DVDD.n20328 DVDD.n20327 0.4505
R29712 DVDD.n20363 DVDD.n20362 0.4505
R29713 DVDD.n20364 DVDD.n20326 0.4505
R29714 DVDD.n20366 DVDD.n20365 0.4505
R29715 DVDD.n19857 DVDD.n19855 0.4505
R29716 DVDD.n20371 DVDD.n20370 0.4505
R29717 DVDD.n19856 DVDD.n19850 0.4505
R29718 DVDD.n20322 DVDD.n20321 0.4505
R29719 DVDD.n20320 DVDD.n20319 0.4505
R29720 DVDD.n20318 DVDD.n20317 0.4505
R29721 DVDD.n19860 DVDD.n19859 0.4505
R29722 DVDD.n20313 DVDD.n20312 0.4505
R29723 DVDD.n20311 DVDD.n20310 0.4505
R29724 DVDD.n20309 DVDD.n20308 0.4505
R29725 DVDD.n19863 DVDD.n19862 0.4505
R29726 DVDD.n20304 DVDD.n20303 0.4505
R29727 DVDD.n20302 DVDD.n20301 0.4505
R29728 DVDD.n20300 DVDD.n20299 0.4505
R29729 DVDD.n19866 DVDD.n19865 0.4505
R29730 DVDD.n20295 DVDD.n20294 0.4505
R29731 DVDD.n20293 DVDD.n19868 0.4505
R29732 DVDD.n20292 DVDD.n20291 0.4505
R29733 DVDD.n19870 DVDD.n19869 0.4505
R29734 DVDD.n20287 DVDD.n20286 0.4505
R29735 DVDD.n20282 DVDD.n19872 0.4505
R29736 DVDD.n20281 DVDD.n20280 0.4505
R29737 DVDD.n19945 DVDD.n19944 0.4505
R29738 DVDD.n20276 DVDD.n20275 0.4505
R29739 DVDD.n20274 DVDD.n20273 0.4505
R29740 DVDD.n20272 DVDD.n20271 0.4505
R29741 DVDD.n19948 DVDD.n19947 0.4505
R29742 DVDD.n20267 DVDD.n20266 0.4505
R29743 DVDD.n20265 DVDD.n20264 0.4505
R29744 DVDD.n20263 DVDD.n20262 0.4505
R29745 DVDD.n19951 DVDD.n19950 0.4505
R29746 DVDD.n20258 DVDD.n20257 0.4505
R29747 DVDD.n20256 DVDD.n20255 0.4505
R29748 DVDD.n20254 DVDD.n19953 0.4505
R29749 DVDD.n20253 DVDD.n20252 0.4505
R29750 DVDD.n19955 DVDD.n19954 0.4505
R29751 DVDD.n20247 DVDD.n20246 0.4505
R29752 DVDD.n20245 DVDD.n19957 0.4505
R29753 DVDD.n20033 DVDD.n19958 0.4505
R29754 DVDD.n20241 DVDD.n20240 0.4505
R29755 DVDD.n20032 DVDD.n20031 0.4505
R29756 DVDD.n20235 DVDD.n20234 0.4505
R29757 DVDD.n20233 DVDD.n20232 0.4505
R29758 DVDD.n20231 DVDD.n20230 0.4505
R29759 DVDD.n20036 DVDD.n20035 0.4505
R29760 DVDD.n20226 DVDD.n20225 0.4505
R29761 DVDD.n20224 DVDD.n20223 0.4505
R29762 DVDD.n20222 DVDD.n20221 0.4505
R29763 DVDD.n20039 DVDD.n20038 0.4505
R29764 DVDD.n20217 DVDD.n20216 0.4505
R29765 DVDD.n20215 DVDD.n20214 0.4505
R29766 DVDD.n20213 DVDD.n20212 0.4505
R29767 DVDD.n20211 DVDD.n20041 0.4505
R29768 DVDD.n20210 DVDD.n20209 0.4505
R29769 DVDD.n20043 DVDD.n19745 0.4505
R29770 DVDD.n20204 DVDD.n19740 0.4505
R29771 DVDD.n20203 DVDD.n20202 0.4505
R29772 DVDD.n20201 DVDD.n20200 0.4505
R29773 DVDD.n20046 DVDD.n20045 0.4505
R29774 DVDD.n20196 DVDD.n20195 0.4505
R29775 DVDD.n20194 DVDD.n20193 0.4505
R29776 DVDD.n20192 DVDD.n20191 0.4505
R29777 DVDD.n20049 DVDD.n20048 0.4505
R29778 DVDD.n20187 DVDD.n20186 0.4505
R29779 DVDD.n20185 DVDD.n20184 0.4505
R29780 DVDD.n20183 DVDD.n20182 0.4505
R29781 DVDD.n20052 DVDD.n20051 0.4505
R29782 DVDD.n20178 DVDD.n20177 0.4505
R29783 DVDD.n20176 DVDD.n20175 0.4505
R29784 DVDD.n20174 DVDD.n20054 0.4505
R29785 DVDD.n20173 DVDD.n20172 0.4505
R29786 DVDD.n20056 DVDD.n20055 0.4505
R29787 DVDD.n20167 DVDD.n20166 0.4505
R29788 DVDD.n20059 DVDD.n20058 0.4505
R29789 DVDD.n20139 DVDD.n20138 0.4505
R29790 DVDD.n20137 DVDD.n20136 0.4505
R29791 DVDD.n20144 DVDD.n20143 0.4505
R29792 DVDD.n20146 DVDD.n20145 0.4505
R29793 DVDD.n20148 DVDD.n20147 0.4505
R29794 DVDD.n20134 DVDD.n20133 0.4505
R29795 DVDD.n20153 DVDD.n20152 0.4505
R29796 DVDD.n20155 DVDD.n20154 0.4505
R29797 DVDD.n20157 DVDD.n20156 0.4505
R29798 DVDD.n20131 DVDD.n20130 0.4505
R29799 DVDD.n20162 DVDD.n20161 0.4505
R29800 DVDD.n20850 DVDD.n20849 0.4505
R29801 DVDD.n20848 DVDD.n18997 0.4505
R29802 DVDD.n20847 DVDD.n20846 0.4505
R29803 DVDD.n20844 DVDD.n18999 0.4505
R29804 DVDD.n20842 DVDD.n20840 0.4505
R29805 DVDD.n20839 DVDD.n19001 0.4505
R29806 DVDD.n20838 DVDD.n20837 0.4505
R29807 DVDD.n20835 DVDD.n19002 0.4505
R29808 DVDD.n20833 DVDD.n20831 0.4505
R29809 DVDD.n20830 DVDD.n19004 0.4505
R29810 DVDD.n20829 DVDD.n20828 0.4505
R29811 DVDD.n20826 DVDD.n19005 0.4505
R29812 DVDD.n20820 DVDD.n19006 0.4505
R29813 DVDD.n20822 DVDD.n20821 0.4505
R29814 DVDD.n20819 DVDD.n19008 0.4505
R29815 DVDD.n20818 DVDD.n20817 0.4505
R29816 DVDD.n20815 DVDD.n19009 0.4505
R29817 DVDD.n20813 DVDD.n20811 0.4505
R29818 DVDD.n20810 DVDD.n19011 0.4505
R29819 DVDD.n20809 DVDD.n20808 0.4505
R29820 DVDD.n20806 DVDD.n19012 0.4505
R29821 DVDD.n20804 DVDD.n20802 0.4505
R29822 DVDD.n20801 DVDD.n19014 0.4505
R29823 DVDD.n20800 DVDD.n20799 0.4505
R29824 DVDD.n20797 DVDD.n19015 0.4505
R29825 DVDD.n20795 DVDD.n20793 0.4505
R29826 DVDD.n20792 DVDD.n19017 0.4505
R29827 DVDD.n20791 DVDD.n20790 0.4505
R29828 DVDD.n20788 DVDD.n19018 0.4505
R29829 DVDD.n20787 DVDD.n20786 0.4505
R29830 DVDD.n20785 DVDD.n19019 0.4505
R29831 DVDD.n20784 DVDD.n20783 0.4505
R29832 DVDD.n19021 DVDD.n19020 0.4505
R29833 DVDD.n20773 DVDD.n19059 0.4505
R29834 DVDD.n20775 DVDD.n20774 0.4505
R29835 DVDD.n20772 DVDD.n19058 0.4505
R29836 DVDD.n20771 DVDD.n20770 0.4505
R29837 DVDD.n20768 DVDD.n19060 0.4505
R29838 DVDD.n20766 DVDD.n20764 0.4505
R29839 DVDD.n20763 DVDD.n19062 0.4505
R29840 DVDD.n20762 DVDD.n20761 0.4505
R29841 DVDD.n20759 DVDD.n19063 0.4505
R29842 DVDD.n20757 DVDD.n20755 0.4505
R29843 DVDD.n20754 DVDD.n19065 0.4505
R29844 DVDD.n20753 DVDD.n20752 0.4505
R29845 DVDD.n20750 DVDD.n19066 0.4505
R29846 DVDD.n20748 DVDD.n19068 0.4505
R29847 DVDD.n20742 DVDD.n19067 0.4505
R29848 DVDD.n20744 DVDD.n20743 0.4505
R29849 DVDD.n20741 DVDD.n19070 0.4505
R29850 DVDD.n20740 DVDD.n20739 0.4505
R29851 DVDD.n19072 DVDD.n19071 0.4505
R29852 DVDD.n20730 DVDD.n19155 0.4505
R29853 DVDD.n20732 DVDD.n20731 0.4505
R29854 DVDD.n20729 DVDD.n19154 0.4505
R29855 DVDD.n20728 DVDD.n20727 0.4505
R29856 DVDD.n20725 DVDD.n19156 0.4505
R29857 DVDD.n20723 DVDD.n20721 0.4505
R29858 DVDD.n20720 DVDD.n19158 0.4505
R29859 DVDD.n20719 DVDD.n20718 0.4505
R29860 DVDD.n20716 DVDD.n19159 0.4505
R29861 DVDD.n20714 DVDD.n20712 0.4505
R29862 DVDD.n20711 DVDD.n19161 0.4505
R29863 DVDD.n20710 DVDD.n20709 0.4505
R29864 DVDD.n20707 DVDD.n19162 0.4505
R29865 DVDD.n20705 DVDD.n19164 0.4505
R29866 DVDD.n20699 DVDD.n19163 0.4505
R29867 DVDD.n20701 DVDD.n20700 0.4505
R29868 DVDD.n20698 DVDD.n19165 0.4505
R29869 DVDD.n20697 DVDD.n20696 0.4505
R29870 DVDD.n20695 DVDD.n19166 0.4505
R29871 DVDD.n20693 DVDD.n20691 0.4505
R29872 DVDD.n20690 DVDD.n19168 0.4505
R29873 DVDD.n20689 DVDD.n20688 0.4505
R29874 DVDD.n20686 DVDD.n19169 0.4505
R29875 DVDD.n20684 DVDD.n20682 0.4505
R29876 DVDD.n20681 DVDD.n19171 0.4505
R29877 DVDD.n20680 DVDD.n20679 0.4505
R29878 DVDD.n20677 DVDD.n19172 0.4505
R29879 DVDD.n20675 DVDD.n20673 0.4505
R29880 DVDD.n20672 DVDD.n19174 0.4505
R29881 DVDD.n20671 DVDD.n20670 0.4505
R29882 DVDD.n20668 DVDD.n19175 0.4505
R29883 DVDD.n20662 DVDD.n19176 0.4505
R29884 DVDD.n20664 DVDD.n20663 0.4505
R29885 DVDD.n20661 DVDD.n19178 0.4505
R29886 DVDD.n20660 DVDD.n20659 0.4505
R29887 DVDD.n19180 DVDD.n19179 0.4505
R29888 DVDD.n20628 DVDD.n20624 0.4505
R29889 DVDD.n20631 DVDD.n20629 0.4505
R29890 DVDD.n20633 DVDD.n20622 0.4505
R29891 DVDD.n20636 DVDD.n20635 0.4505
R29892 DVDD.n20637 DVDD.n20621 0.4505
R29893 DVDD.n20640 DVDD.n20638 0.4505
R29894 DVDD.n20642 DVDD.n20619 0.4505
R29895 DVDD.n20650 DVDD.n20649 0.4505
R29896 DVDD.n20651 DVDD.n20618 0.4505
R29897 DVDD.n20653 DVDD.n20652 0.4505
R29898 DVDD.n18998 DVDD.n18973 0.4505
R29899 DVDD.n20851 DVDD.n20850 0.4505
R29900 DVDD.n18997 DVDD.n18996 0.4505
R29901 DVDD.n20846 DVDD.n20845 0.4505
R29902 DVDD.n20844 DVDD.n20843 0.4505
R29903 DVDD.n20842 DVDD.n20841 0.4505
R29904 DVDD.n19001 DVDD.n19000 0.4505
R29905 DVDD.n20837 DVDD.n20836 0.4505
R29906 DVDD.n20835 DVDD.n20834 0.4505
R29907 DVDD.n20833 DVDD.n20832 0.4505
R29908 DVDD.n19004 DVDD.n19003 0.4505
R29909 DVDD.n20828 DVDD.n20827 0.4505
R29910 DVDD.n20826 DVDD.n20825 0.4505
R29911 DVDD.n20824 DVDD.n19006 0.4505
R29912 DVDD.n20823 DVDD.n20822 0.4505
R29913 DVDD.n19008 DVDD.n19007 0.4505
R29914 DVDD.n20817 DVDD.n20816 0.4505
R29915 DVDD.n20815 DVDD.n20814 0.4505
R29916 DVDD.n20813 DVDD.n20812 0.4505
R29917 DVDD.n19011 DVDD.n19010 0.4505
R29918 DVDD.n20808 DVDD.n20807 0.4505
R29919 DVDD.n20806 DVDD.n20805 0.4505
R29920 DVDD.n20804 DVDD.n20803 0.4505
R29921 DVDD.n19014 DVDD.n19013 0.4505
R29922 DVDD.n20799 DVDD.n20798 0.4505
R29923 DVDD.n20797 DVDD.n20796 0.4505
R29924 DVDD.n20795 DVDD.n20794 0.4505
R29925 DVDD.n19017 DVDD.n19016 0.4505
R29926 DVDD.n20790 DVDD.n20789 0.4505
R29927 DVDD.n20788 DVDD.n18893 0.4505
R29928 DVDD.n20787 DVDD.n18887 0.4505
R29929 DVDD.n20781 DVDD.n19019 0.4505
R29930 DVDD.n20783 DVDD.n20782 0.4505
R29931 DVDD.n20780 DVDD.n19021 0.4505
R29932 DVDD.n19059 DVDD.n19022 0.4505
R29933 DVDD.n20776 DVDD.n20775 0.4505
R29934 DVDD.n19058 DVDD.n19054 0.4505
R29935 DVDD.n20770 DVDD.n20769 0.4505
R29936 DVDD.n20768 DVDD.n20767 0.4505
R29937 DVDD.n20766 DVDD.n20765 0.4505
R29938 DVDD.n19062 DVDD.n19061 0.4505
R29939 DVDD.n20761 DVDD.n20760 0.4505
R29940 DVDD.n20759 DVDD.n20758 0.4505
R29941 DVDD.n20757 DVDD.n20756 0.4505
R29942 DVDD.n19065 DVDD.n19064 0.4505
R29943 DVDD.n20752 DVDD.n20751 0.4505
R29944 DVDD.n20750 DVDD.n20749 0.4505
R29945 DVDD.n20748 DVDD.n20747 0.4505
R29946 DVDD.n20746 DVDD.n19067 0.4505
R29947 DVDD.n20745 DVDD.n20744 0.4505
R29948 DVDD.n19070 DVDD.n19069 0.4505
R29949 DVDD.n20739 DVDD.n20738 0.4505
R29950 DVDD.n20737 DVDD.n19072 0.4505
R29951 DVDD.n19155 DVDD.n19073 0.4505
R29952 DVDD.n20733 DVDD.n20732 0.4505
R29953 DVDD.n19154 DVDD.n19149 0.4505
R29954 DVDD.n20727 DVDD.n20726 0.4505
R29955 DVDD.n20725 DVDD.n20724 0.4505
R29956 DVDD.n20723 DVDD.n20722 0.4505
R29957 DVDD.n19158 DVDD.n19157 0.4505
R29958 DVDD.n20718 DVDD.n20717 0.4505
R29959 DVDD.n20716 DVDD.n20715 0.4505
R29960 DVDD.n20714 DVDD.n20713 0.4505
R29961 DVDD.n19161 DVDD.n19160 0.4505
R29962 DVDD.n20709 DVDD.n20708 0.4505
R29963 DVDD.n20707 DVDD.n20706 0.4505
R29964 DVDD.n20705 DVDD.n20704 0.4505
R29965 DVDD.n20703 DVDD.n19163 0.4505
R29966 DVDD.n20702 DVDD.n20701 0.4505
R29967 DVDD.n19165 DVDD.n18853 0.4505
R29968 DVDD.n20696 DVDD.n18847 0.4505
R29969 DVDD.n20695 DVDD.n20694 0.4505
R29970 DVDD.n20693 DVDD.n20692 0.4505
R29971 DVDD.n19168 DVDD.n19167 0.4505
R29972 DVDD.n20688 DVDD.n20687 0.4505
R29973 DVDD.n20686 DVDD.n20685 0.4505
R29974 DVDD.n20684 DVDD.n20683 0.4505
R29975 DVDD.n19171 DVDD.n19170 0.4505
R29976 DVDD.n20679 DVDD.n20678 0.4505
R29977 DVDD.n20677 DVDD.n20676 0.4505
R29978 DVDD.n20675 DVDD.n20674 0.4505
R29979 DVDD.n19174 DVDD.n19173 0.4505
R29980 DVDD.n20670 DVDD.n20669 0.4505
R29981 DVDD.n20668 DVDD.n20667 0.4505
R29982 DVDD.n20666 DVDD.n19176 0.4505
R29983 DVDD.n20665 DVDD.n20664 0.4505
R29984 DVDD.n19178 DVDD.n19177 0.4505
R29985 DVDD.n20659 DVDD.n20658 0.4505
R29986 DVDD.n19181 DVDD.n19180 0.4505
R29987 DVDD.n20626 DVDD.n20625 0.4505
R29988 DVDD.n20624 DVDD.n20623 0.4505
R29989 DVDD.n20631 DVDD.n20630 0.4505
R29990 DVDD.n20633 DVDD.n20632 0.4505
R29991 DVDD.n20635 DVDD.n20634 0.4505
R29992 DVDD.n20621 DVDD.n20620 0.4505
R29993 DVDD.n20640 DVDD.n20639 0.4505
R29994 DVDD.n20642 DVDD.n20641 0.4505
R29995 DVDD.n20649 DVDD.n20648 0.4505
R29996 DVDD.n20618 DVDD.n20617 0.4505
R29997 DVDD.n20654 DVDD.n20653 0.4505
R29998 DVDD.n3973 DVDD.n3964 0.4505
R29999 DVDD.n3963 DVDD.n3941 0.4505
R30000 DVDD.n3962 DVDD.n3961 0.4505
R30001 DVDD.n3959 DVDD.n3942 0.4505
R30002 DVDD.n3957 DVDD.n3955 0.4505
R30003 DVDD.n3954 DVDD.n3944 0.4505
R30004 DVDD.n3953 DVDD.n3952 0.4505
R30005 DVDD.n3950 DVDD.n3945 0.4505
R30006 DVDD.n3948 DVDD.n3946 0.4505
R30007 DVDD.n3909 DVDD.n3908 0.4505
R30008 DVDD.n3981 DVDD.n3980 0.4505
R30009 DVDD.n3982 DVDD.n3907 0.4505
R30010 DVDD.n3984 DVDD.n3983 0.4505
R30011 DVDD.n3905 DVDD.n3904 0.4505
R30012 DVDD.n3990 DVDD.n3989 0.4505
R30013 DVDD.n3991 DVDD.n3903 0.4505
R30014 DVDD.n3994 DVDD.n3992 0.4505
R30015 DVDD.n3996 DVDD.n3902 0.4505
R30016 DVDD.n3999 DVDD.n3998 0.4505
R30017 DVDD.n4000 DVDD.n3899 0.4505
R30018 DVDD.n4061 DVDD.n4060 0.4505
R30019 DVDD.n4059 DVDD.n3901 0.4505
R30020 DVDD.n4058 DVDD.n4057 0.4505
R30021 DVDD.n4055 DVDD.n4001 0.4505
R30022 DVDD.n4053 DVDD.n4051 0.4505
R30023 DVDD.n4050 DVDD.n4003 0.4505
R30024 DVDD.n4049 DVDD.n4048 0.4505
R30025 DVDD.n4046 DVDD.n4004 0.4505
R30026 DVDD.n4044 DVDD.n4043 0.4505
R30027 DVDD.n4042 DVDD.n4005 0.4505
R30028 DVDD.n4041 DVDD.n4040 0.4505
R30029 DVDD.n4007 DVDD.n4006 0.4505
R30030 DVDD.n4036 DVDD.n4035 0.4505
R30031 DVDD.n4034 DVDD.n4009 0.4505
R30032 DVDD.n4033 DVDD.n4032 0.4505
R30033 DVDD.n4030 DVDD.n4010 0.4505
R30034 DVDD.n4028 DVDD.n4026 0.4505
R30035 DVDD.n4025 DVDD.n4012 0.4505
R30036 DVDD.n4024 DVDD.n4023 0.4505
R30037 DVDD.n4021 DVDD.n4013 0.4505
R30038 DVDD.n4019 DVDD.n4017 0.4505
R30039 DVDD.n4016 DVDD.n4015 0.4505
R30040 DVDD.n276 DVDD.n273 0.4505
R30041 DVDD.n22176 DVDD.n22175 0.4505
R30042 DVDD.n22174 DVDD.n275 0.4505
R30043 DVDD.n22173 DVDD.n22172 0.4505
R30044 DVDD.n22171 DVDD.n277 0.4505
R30045 DVDD.n22170 DVDD.n279 0.4505
R30046 DVDD.n282 DVDD.n278 0.4505
R30047 DVDD.n22166 DVDD.n22165 0.4505
R30048 DVDD.n22164 DVDD.n281 0.4505
R30049 DVDD.n22163 DVDD.n22162 0.4505
R30050 DVDD.n284 DVDD.n283 0.4505
R30051 DVDD.n334 DVDD.n332 0.4505
R30052 DVDD.n336 DVDD.n331 0.4505
R30053 DVDD.n339 DVDD.n338 0.4505
R30054 DVDD.n340 DVDD.n330 0.4505
R30055 DVDD.n343 DVDD.n341 0.4505
R30056 DVDD.n345 DVDD.n328 0.4505
R30057 DVDD.n348 DVDD.n347 0.4505
R30058 DVDD.n349 DVDD.n325 0.4505
R30059 DVDD.n22154 DVDD.n22153 0.4505
R30060 DVDD.n22152 DVDD.n327 0.4505
R30061 DVDD.n22151 DVDD.n22150 0.4505
R30062 DVDD.n22148 DVDD.n350 0.4505
R30063 DVDD.n22147 DVDD.n22146 0.4505
R30064 DVDD.n22145 DVDD.n351 0.4505
R30065 DVDD.n22144 DVDD.n22143 0.4505
R30066 DVDD.n353 DVDD.n352 0.4505
R30067 DVDD.n400 DVDD.n399 0.4505
R30068 DVDD.n403 DVDD.n401 0.4505
R30069 DVDD.n405 DVDD.n398 0.4505
R30070 DVDD.n408 DVDD.n407 0.4505
R30071 DVDD.n409 DVDD.n397 0.4505
R30072 DVDD.n412 DVDD.n410 0.4505
R30073 DVDD.n414 DVDD.n395 0.4505
R30074 DVDD.n417 DVDD.n416 0.4505
R30075 DVDD.n418 DVDD.n394 0.4505
R30076 DVDD.n420 DVDD.n419 0.4505
R30077 DVDD.n428 DVDD.n392 0.4505
R30078 DVDD.n431 DVDD.n430 0.4505
R30079 DVDD.n432 DVDD.n390 0.4505
R30080 DVDD.n22136 DVDD.n22135 0.4505
R30081 DVDD.n22134 DVDD.n391 0.4505
R30082 DVDD.n22133 DVDD.n22132 0.4505
R30083 DVDD.n434 DVDD.n433 0.4505
R30084 DVDD.n22128 DVDD.n22127 0.4505
R30085 DVDD.n22126 DVDD.n436 0.4505
R30086 DVDD.n22125 DVDD.n22124 0.4505
R30087 DVDD.n438 DVDD.n437 0.4505
R30088 DVDD.n22094 DVDD.n22092 0.4505
R30089 DVDD.n22097 DVDD.n22096 0.4505
R30090 DVDD.n22098 DVDD.n22091 0.4505
R30091 DVDD.n22101 DVDD.n22099 0.4505
R30092 DVDD.n22103 DVDD.n22089 0.4505
R30093 DVDD.n22106 DVDD.n22105 0.4505
R30094 DVDD.n22108 DVDD.n22107 0.4505
R30095 DVDD.n22117 DVDD.n22088 0.4505
R30096 DVDD.n3975 DVDD.n3974 0.4505
R30097 DVDD.n3973 DVDD.n3972 0.4505
R30098 DVDD.n3966 DVDD.n3941 0.4505
R30099 DVDD.n3961 DVDD.n3960 0.4505
R30100 DVDD.n3959 DVDD.n3958 0.4505
R30101 DVDD.n3957 DVDD.n3956 0.4505
R30102 DVDD.n3944 DVDD.n3943 0.4505
R30103 DVDD.n3952 DVDD.n3951 0.4505
R30104 DVDD.n3950 DVDD.n3949 0.4505
R30105 DVDD.n3948 DVDD.n3947 0.4505
R30106 DVDD.n3926 DVDD.n3909 0.4505
R30107 DVDD.n3980 DVDD.n3979 0.4505
R30108 DVDD.n3907 DVDD.n3906 0.4505
R30109 DVDD.n3985 DVDD.n3984 0.4505
R30110 DVDD.n3986 DVDD.n3905 0.4505
R30111 DVDD.n3989 DVDD.n3988 0.4505
R30112 DVDD.n3987 DVDD.n3903 0.4505
R30113 DVDD.n3994 DVDD.n3993 0.4505
R30114 DVDD.n3996 DVDD.n3995 0.4505
R30115 DVDD.n3998 DVDD.n3997 0.4505
R30116 DVDD.n3899 DVDD.n3898 0.4505
R30117 DVDD.n4062 DVDD.n4061 0.4505
R30118 DVDD.n3901 DVDD.n3900 0.4505
R30119 DVDD.n4057 DVDD.n4056 0.4505
R30120 DVDD.n4055 DVDD.n4054 0.4505
R30121 DVDD.n4053 DVDD.n4052 0.4505
R30122 DVDD.n4003 DVDD.n4002 0.4505
R30123 DVDD.n4048 DVDD.n4047 0.4505
R30124 DVDD.n4046 DVDD.n4045 0.4505
R30125 DVDD.n4044 DVDD.n3876 0.4505
R30126 DVDD.n4005 DVDD.n3883 0.4505
R30127 DVDD.n4040 DVDD.n4039 0.4505
R30128 DVDD.n4038 DVDD.n4007 0.4505
R30129 DVDD.n4037 DVDD.n4036 0.4505
R30130 DVDD.n4009 DVDD.n4008 0.4505
R30131 DVDD.n4032 DVDD.n4031 0.4505
R30132 DVDD.n4030 DVDD.n4029 0.4505
R30133 DVDD.n4028 DVDD.n4027 0.4505
R30134 DVDD.n4012 DVDD.n4011 0.4505
R30135 DVDD.n4023 DVDD.n4022 0.4505
R30136 DVDD.n4021 DVDD.n4020 0.4505
R30137 DVDD.n4019 DVDD.n4018 0.4505
R30138 DVDD.n4015 DVDD.n4014 0.4505
R30139 DVDD.n273 DVDD.n272 0.4505
R30140 DVDD.n22177 DVDD.n22176 0.4505
R30141 DVDD.n275 DVDD.n274 0.4505
R30142 DVDD.n22172 DVDD.n251 0.4505
R30143 DVDD.n22171 DVDD.n257 0.4505
R30144 DVDD.n22170 DVDD.n22169 0.4505
R30145 DVDD.n22168 DVDD.n278 0.4505
R30146 DVDD.n22167 DVDD.n22166 0.4505
R30147 DVDD.n281 DVDD.n280 0.4505
R30148 DVDD.n22162 DVDD.n22161 0.4505
R30149 DVDD.n290 DVDD.n284 0.4505
R30150 DVDD.n334 DVDD.n333 0.4505
R30151 DVDD.n336 DVDD.n335 0.4505
R30152 DVDD.n338 DVDD.n337 0.4505
R30153 DVDD.n330 DVDD.n329 0.4505
R30154 DVDD.n343 DVDD.n342 0.4505
R30155 DVDD.n345 DVDD.n344 0.4505
R30156 DVDD.n347 DVDD.n346 0.4505
R30157 DVDD.n325 DVDD.n324 0.4505
R30158 DVDD.n22155 DVDD.n22154 0.4505
R30159 DVDD.n327 DVDD.n326 0.4505
R30160 DVDD.n22150 DVDD.n22149 0.4505
R30161 DVDD.n22148 DVDD.n304 0.4505
R30162 DVDD.n22147 DVDD.n310 0.4505
R30163 DVDD.n354 DVDD.n351 0.4505
R30164 DVDD.n22143 DVDD.n22142 0.4505
R30165 DVDD.n22141 DVDD.n353 0.4505
R30166 DVDD.n399 DVDD.n360 0.4505
R30167 DVDD.n403 DVDD.n402 0.4505
R30168 DVDD.n405 DVDD.n404 0.4505
R30169 DVDD.n407 DVDD.n406 0.4505
R30170 DVDD.n397 DVDD.n396 0.4505
R30171 DVDD.n412 DVDD.n411 0.4505
R30172 DVDD.n414 DVDD.n413 0.4505
R30173 DVDD.n416 DVDD.n415 0.4505
R30174 DVDD.n394 DVDD.n393 0.4505
R30175 DVDD.n421 DVDD.n420 0.4505
R30176 DVDD.n428 DVDD.n427 0.4505
R30177 DVDD.n430 DVDD.n429 0.4505
R30178 DVDD.n390 DVDD.n388 0.4505
R30179 DVDD.n22137 DVDD.n22136 0.4505
R30180 DVDD.n391 DVDD.n389 0.4505
R30181 DVDD.n22132 DVDD.n22131 0.4505
R30182 DVDD.n22130 DVDD.n434 0.4505
R30183 DVDD.n22129 DVDD.n22128 0.4505
R30184 DVDD.n439 DVDD.n436 0.4505
R30185 DVDD.n22124 DVDD.n22123 0.4505
R30186 DVDD.n446 DVDD.n438 0.4505
R30187 DVDD.n22094 DVDD.n22093 0.4505
R30188 DVDD.n22096 DVDD.n22095 0.4505
R30189 DVDD.n22091 DVDD.n22090 0.4505
R30190 DVDD.n22101 DVDD.n22100 0.4505
R30191 DVDD.n22103 DVDD.n22102 0.4505
R30192 DVDD.n22105 DVDD.n22104 0.4505
R30193 DVDD.n22109 DVDD.n22108 0.4505
R30194 DVDD.n22117 DVDD.n22116 0.4505
R30195 DVDD.n22118 DVDD.n22087 0.4505
R30196 DVDD.n18091 DVDD.n18070 0.4505
R30197 DVDD.n4576 DVDD.n4575 0.4505
R30198 DVDD.n4279 DVDD.n4278 0.4505
R30199 DVDD.n4580 DVDD.n4280 0.4505
R30200 DVDD.n4581 DVDD.n4252 0.4505
R30201 DVDD.n4582 DVDD.n4258 0.4505
R30202 DVDD.n4274 DVDD.n4271 0.4505
R30203 DVDD.n4596 DVDD.n4595 0.4505
R30204 DVDD.n4276 DVDD.n4275 0.4505
R30205 DVDD.n4591 DVDD.n4590 0.4505
R30206 DVDD.n4589 DVDD.n4588 0.4505
R30207 DVDD.n4587 DVDD.n488 0.4505
R30208 DVDD.n18133 DVDD.n18132 0.4505
R30209 DVDD.n491 DVDD.n489 0.4505
R30210 DVDD.n18128 DVDD.n18127 0.4505
R30211 DVDD.n502 DVDD.n495 0.4505
R30212 DVDD.n18073 DVDD.n18072 0.4505
R30213 DVDD.n18077 DVDD.n18074 0.4505
R30214 DVDD.n18079 DVDD.n18078 0.4505
R30215 DVDD.n18087 DVDD.n18086 0.4505
R30216 DVDD.n18084 DVDD.n18069 0.4505
R30217 DVDD.n18091 DVDD.n18090 0.4505
R30218 DVDD.n18089 DVDD.n18069 0.4505
R30219 DVDD.n18088 DVDD.n18087 0.4505
R30220 DVDD.n18079 DVDD.n18071 0.4505
R30221 DVDD.n18077 DVDD.n18076 0.4505
R30222 DVDD.n18075 DVDD.n18073 0.4505
R30223 DVDD.n495 DVDD.n494 0.4505
R30224 DVDD.n18129 DVDD.n18128 0.4505
R30225 DVDD.n18130 DVDD.n491 0.4505
R30226 DVDD.n18132 DVDD.n18131 0.4505
R30227 DVDD.n4587 DVDD.n4586 0.4505
R30228 DVDD.n4588 DVDD.n4585 0.4505
R30229 DVDD.n4592 DVDD.n4591 0.4505
R30230 DVDD.n4593 DVDD.n4276 0.4505
R30231 DVDD.n4595 DVDD.n4594 0.4505
R30232 DVDD.n4584 DVDD.n4274 0.4505
R30233 DVDD.n4583 DVDD.n4582 0.4505
R30234 DVDD.n4581 DVDD.n4277 0.4505
R30235 DVDD.n4580 DVDD.n4579 0.4505
R30236 DVDD.n4578 DVDD.n4279 0.4505
R30237 DVDD.n4577 DVDD.n4576 0.4505
R30238 DVDD.n3612 DVDD.n3611 0.4505
R30239 DVDD.n3615 DVDD.n3613 0.4505
R30240 DVDD.n3617 DVDD.n3616 0.4505
R30241 DVDD.n3619 DVDD.n3618 0.4505
R30242 DVDD.n3608 DVDD.n3607 0.4505
R30243 DVDD.n3623 DVDD.n3609 0.4505
R30244 DVDD.n3625 DVDD.n3624 0.4505
R30245 DVDD.n3627 DVDD.n3626 0.4505
R30246 DVDD.n3605 DVDD.n3604 0.4505
R30247 DVDD.n3631 DVDD.n3603 0.4505
R30248 DVDD.n3633 DVDD.n3632 0.4505
R30249 DVDD.n4779 DVDD.n4778 0.4505
R30250 DVDD.n4777 DVDD.n3602 0.4505
R30251 DVDD.n4776 DVDD.n4775 0.4505
R30252 DVDD.n3639 DVDD.n3636 0.4505
R30253 DVDD.n4771 DVDD.n4770 0.4505
R30254 DVDD.n3646 DVDD.n3638 0.4505
R30255 DVDD.n3669 DVDD.n3668 0.4505
R30256 DVDD.n4766 DVDD.n4765 0.4505
R30257 DVDD.n3671 DVDD.n3670 0.4505
R30258 DVDD.n4761 DVDD.n4760 0.4505
R30259 DVDD.n4762 DVDD.n4761 0.4505
R30260 DVDD.n4763 DVDD.n3671 0.4505
R30261 DVDD.n4765 DVDD.n4764 0.4505
R30262 DVDD.n3672 DVDD.n3669 0.4505
R30263 DVDD.n3638 DVDD.n3637 0.4505
R30264 DVDD.n4772 DVDD.n4771 0.4505
R30265 DVDD.n4773 DVDD.n3636 0.4505
R30266 DVDD.n4775 DVDD.n4774 0.4505
R30267 DVDD.n3602 DVDD.n3601 0.4505
R30268 DVDD.n4780 DVDD.n4779 0.4505
R30269 DVDD.n3632 DVDD.n3600 0.4505
R30270 DVDD.n3631 DVDD.n3630 0.4505
R30271 DVDD.n3629 DVDD.n3605 0.4505
R30272 DVDD.n3628 DVDD.n3627 0.4505
R30273 DVDD.n3625 DVDD.n3606 0.4505
R30274 DVDD.n3623 DVDD.n3622 0.4505
R30275 DVDD.n3621 DVDD.n3608 0.4505
R30276 DVDD.n3620 DVDD.n3619 0.4505
R30277 DVDD.n3617 DVDD.n3610 0.4505
R30278 DVDD.n3615 DVDD.n3614 0.4505
R30279 DVDD.n3612 DVDD.n3542 0.4505
R30280 DVDD.n4572 DVDD.n4571 0.4505
R30281 DVDD.n4570 DVDD.n4316 0.4505
R30282 DVDD.n4569 DVDD.n4568 0.4505
R30283 DVDD.n4318 DVDD.n4317 0.4505
R30284 DVDD.n4564 DVDD.n4563 0.4505
R30285 DVDD.n4562 DVDD.n4320 0.4505
R30286 DVDD.n4561 DVDD.n4560 0.4505
R30287 DVDD.n4322 DVDD.n4321 0.4505
R30288 DVDD.n4476 DVDD.n4474 0.4505
R30289 DVDD.n4477 DVDD.n4200 0.4505
R30290 DVDD.n4536 DVDD.n4199 0.4505
R30291 DVDD.n4538 DVDD.n4461 0.4505
R30292 DVDD.n4541 DVDD.n4540 0.4505
R30293 DVDD.n4542 DVDD.n4460 0.4505
R30294 DVDD.n4545 DVDD.n4543 0.4505
R30295 DVDD.n4547 DVDD.n4458 0.4505
R30296 DVDD.n4550 DVDD.n4549 0.4505
R30297 DVDD.n4551 DVDD.n4414 0.4505
R30298 DVDD.n4553 DVDD.n4552 0.4505
R30299 DVDD.n4457 DVDD.n4412 0.4505
R30300 DVDD.n4456 DVDD.n4455 0.4505
R30301 DVDD.n4758 DVDD.n3713 0.4505
R30302 DVDD.n3711 DVDD.n3676 0.4505
R30303 DVDD.n4754 DVDD.n4753 0.4505
R30304 DVDD.n4751 DVDD.n3715 0.4505
R30305 DVDD.n4750 DVDD.n4749 0.4505
R30306 DVDD.n3719 DVDD.n3718 0.4505
R30307 DVDD.n4745 DVDD.n4744 0.4505
R30308 DVDD.n3727 DVDD.n3721 0.4505
R30309 DVDD.n3754 DVDD.n3753 0.4505
R30310 DVDD.n4740 DVDD.n4739 0.4505
R30311 DVDD.n3817 DVDD.n3755 0.4505
R30312 DVDD.n4428 DVDD.n4427 0.4505
R30313 DVDD.n4431 DVDD.n4429 0.4505
R30314 DVDD.n4433 DVDD.n4432 0.4505
R30315 DVDD.n4435 DVDD.n4434 0.4505
R30316 DVDD.n4424 DVDD.n4423 0.4505
R30317 DVDD.n4439 DVDD.n4425 0.4505
R30318 DVDD.n4443 DVDD.n4442 0.4505
R30319 DVDD.n4445 DVDD.n4444 0.4505
R30320 DVDD.n4421 DVDD.n4420 0.4505
R30321 DVDD.n4450 DVDD.n4449 0.4505
R30322 DVDD.n4449 DVDD.n4448 0.4505
R30323 DVDD.n4447 DVDD.n4421 0.4505
R30324 DVDD.n4446 DVDD.n4445 0.4505
R30325 DVDD.n4443 DVDD.n4422 0.4505
R30326 DVDD.n4439 DVDD.n4438 0.4505
R30327 DVDD.n4437 DVDD.n4424 0.4505
R30328 DVDD.n4436 DVDD.n4435 0.4505
R30329 DVDD.n4433 DVDD.n4426 0.4505
R30330 DVDD.n4431 DVDD.n4430 0.4505
R30331 DVDD.n4428 DVDD.n3757 0.4505
R30332 DVDD.n4737 DVDD.n3755 0.4505
R30333 DVDD.n4739 DVDD.n4738 0.4505
R30334 DVDD.n3756 DVDD.n3754 0.4505
R30335 DVDD.n3721 DVDD.n3720 0.4505
R30336 DVDD.n4746 DVDD.n4745 0.4505
R30337 DVDD.n4747 DVDD.n3719 0.4505
R30338 DVDD.n4749 DVDD.n4748 0.4505
R30339 DVDD.n3715 DVDD.n3714 0.4505
R30340 DVDD.n4755 DVDD.n4754 0.4505
R30341 DVDD.n4756 DVDD.n3676 0.4505
R30342 DVDD.n4758 DVDD.n4757 0.4505
R30343 DVDD.n4455 DVDD.n4454 0.4505
R30344 DVDD.n4412 DVDD.n4407 0.4505
R30345 DVDD.n4554 DVDD.n4553 0.4505
R30346 DVDD.n4414 DVDD.n4413 0.4505
R30347 DVDD.n4549 DVDD.n4548 0.4505
R30348 DVDD.n4547 DVDD.n4546 0.4505
R30349 DVDD.n4545 DVDD.n4544 0.4505
R30350 DVDD.n4460 DVDD.n4459 0.4505
R30351 DVDD.n4540 DVDD.n4539 0.4505
R30352 DVDD.n4538 DVDD.n4537 0.4505
R30353 DVDD.n4536 DVDD.n4535 0.4505
R30354 DVDD.n4478 DVDD.n4477 0.4505
R30355 DVDD.n4476 DVDD.n4475 0.4505
R30356 DVDD.n4398 DVDD.n4322 0.4505
R30357 DVDD.n4560 DVDD.n4559 0.4505
R30358 DVDD.n4320 DVDD.n4319 0.4505
R30359 DVDD.n4565 DVDD.n4564 0.4505
R30360 DVDD.n4566 DVDD.n4318 0.4505
R30361 DVDD.n4568 DVDD.n4567 0.4505
R30362 DVDD.n4316 DVDD.n4315 0.4505
R30363 DVDD.n4573 DVDD.n4572 0.4505
R30364 DVDD.n10021 DVDD.n10019 0.4505
R30365 DVDD.n10024 DVDD.n10023 0.4505
R30366 DVDD.n10025 DVDD.n10015 0.4505
R30367 DVDD.n10028 DVDD.n10026 0.4505
R30368 DVDD.n10030 DVDD.n10013 0.4505
R30369 DVDD.n10033 DVDD.n10032 0.4505
R30370 DVDD.n10034 DVDD.n10012 0.4505
R30371 DVDD.n10037 DVDD.n10035 0.4505
R30372 DVDD.n10039 DVDD.n10010 0.4505
R30373 DVDD.n10042 DVDD.n10041 0.4505
R30374 DVDD.n9840 DVDD.n9839 0.4505
R30375 DVDD.n9843 DVDD.n9841 0.4505
R30376 DVDD.n9845 DVDD.n9836 0.4505
R30377 DVDD.n9848 DVDD.n9847 0.4505
R30378 DVDD.n9849 DVDD.n9835 0.4505
R30379 DVDD.n9852 DVDD.n9850 0.4505
R30380 DVDD.n9854 DVDD.n9833 0.4505
R30381 DVDD.n9857 DVDD.n9856 0.4505
R30382 DVDD.n9858 DVDD.n9832 0.4505
R30383 DVDD.n9861 DVDD.n9859 0.4505
R30384 DVDD.n9863 DVDD.n9830 0.4505
R30385 DVDD.n9866 DVDD.n9865 0.4505
R30386 DVDD.n9867 DVDD.n9829 0.4505
R30387 DVDD.n9870 DVDD.n9869 0.4505
R30388 DVDD.n9868 DVDD.n9826 0.4505
R30389 DVDD.n9874 DVDD.n9827 0.4505
R30390 DVDD.n9876 DVDD.n9825 0.4505
R30391 DVDD.n9879 DVDD.n9878 0.4505
R30392 DVDD.n9880 DVDD.n9824 0.4505
R30393 DVDD.n9883 DVDD.n9881 0.4505
R30394 DVDD.n9885 DVDD.n9822 0.4505
R30395 DVDD.n9888 DVDD.n9887 0.4505
R30396 DVDD.n9889 DVDD.n9821 0.4505
R30397 DVDD.n9892 DVDD.n9890 0.4505
R30398 DVDD.n9894 DVDD.n9819 0.4505
R30399 DVDD.n9897 DVDD.n9896 0.4505
R30400 DVDD.n9898 DVDD.n9817 0.4505
R30401 DVDD.n9936 DVDD.n9935 0.4505
R30402 DVDD.n9934 DVDD.n9818 0.4505
R30403 DVDD.n9933 DVDD.n9932 0.4505
R30404 DVDD.n9931 DVDD.n9899 0.4505
R30405 DVDD.n9903 DVDD.n9900 0.4505
R30406 DVDD.n9927 DVDD.n9926 0.4505
R30407 DVDD.n9925 DVDD.n9902 0.4505
R30408 DVDD.n9924 DVDD.n9923 0.4505
R30409 DVDD.n9921 DVDD.n9904 0.4505
R30410 DVDD.n9919 DVDD.n9917 0.4505
R30411 DVDD.n9916 DVDD.n9906 0.4505
R30412 DVDD.n9915 DVDD.n9914 0.4505
R30413 DVDD.n9912 DVDD.n9907 0.4505
R30414 DVDD.n9910 DVDD.n9908 0.4505
R30415 DVDD.n9651 DVDD.n9644 0.4505
R30416 DVDD.n10089 DVDD.n10088 0.4505
R30417 DVDD.n10087 DVDD.n9650 0.4505
R30418 DVDD.n10086 DVDD.n10085 0.4505
R30419 DVDD.n10083 DVDD.n9652 0.4505
R30420 DVDD.n10082 DVDD.n10081 0.4505
R30421 DVDD.n10080 DVDD.n9653 0.4505
R30422 DVDD.n10079 DVDD.n10078 0.4505
R30423 DVDD.n9655 DVDD.n9654 0.4505
R30424 DVDD.n10074 DVDD.n10073 0.4505
R30425 DVDD.n10072 DVDD.n9658 0.4505
R30426 DVDD.n10071 DVDD.n10070 0.4505
R30427 DVDD.n9660 DVDD.n9659 0.4505
R30428 DVDD.n9708 DVDD.n9706 0.4505
R30429 DVDD.n9711 DVDD.n9710 0.4505
R30430 DVDD.n9712 DVDD.n9705 0.4505
R30431 DVDD.n9715 DVDD.n9713 0.4505
R30432 DVDD.n9717 DVDD.n9703 0.4505
R30433 DVDD.n9720 DVDD.n9719 0.4505
R30434 DVDD.n9721 DVDD.n9702 0.4505
R30435 DVDD.n9724 DVDD.n9722 0.4505
R30436 DVDD.n9726 DVDD.n9700 0.4505
R30437 DVDD.n9729 DVDD.n9728 0.4505
R30438 DVDD.n9730 DVDD.n9698 0.4505
R30439 DVDD.n10064 DVDD.n10063 0.4505
R30440 DVDD.n10062 DVDD.n9699 0.4505
R30441 DVDD.n10061 DVDD.n10060 0.4505
R30442 DVDD.n9732 DVDD.n9731 0.4505
R30443 DVDD.n9976 DVDD.n9975 0.4505
R30444 DVDD.n9979 DVDD.n9977 0.4505
R30445 DVDD.n9981 DVDD.n9974 0.4505
R30446 DVDD.n9984 DVDD.n9983 0.4505
R30447 DVDD.n9985 DVDD.n9973 0.4505
R30448 DVDD.n9988 DVDD.n9986 0.4505
R30449 DVDD.n9990 DVDD.n9971 0.4505
R30450 DVDD.n9993 DVDD.n9992 0.4505
R30451 DVDD.n9994 DVDD.n9970 0.4505
R30452 DVDD.n9996 DVDD.n9995 0.4505
R30453 DVDD.n10003 DVDD.n9968 0.4505
R30454 DVDD.n10006 DVDD.n10005 0.4505
R30455 DVDD.n10007 DVDD.n9966 0.4505
R30456 DVDD.n10053 DVDD.n10052 0.4505
R30457 DVDD.n10051 DVDD.n9967 0.4505
R30458 DVDD.n10050 DVDD.n10049 0.4505
R30459 DVDD.n10046 DVDD.n10008 0.4505
R30460 DVDD.n10045 DVDD.n10044 0.4505
R30461 DVDD.n10043 DVDD.n10009 0.4505
R30462 DVDD.n10017 DVDD.n10016 0.4505
R30463 DVDD.n10021 DVDD.n10020 0.4505
R30464 DVDD.n10023 DVDD.n10022 0.4505
R30465 DVDD.n10015 DVDD.n10014 0.4505
R30466 DVDD.n10028 DVDD.n10027 0.4505
R30467 DVDD.n10030 DVDD.n10029 0.4505
R30468 DVDD.n10032 DVDD.n10031 0.4505
R30469 DVDD.n10012 DVDD.n10011 0.4505
R30470 DVDD.n10037 DVDD.n10036 0.4505
R30471 DVDD.n10039 DVDD.n10038 0.4505
R30472 DVDD.n10041 DVDD.n10040 0.4505
R30473 DVDD.n9837 DVDD.n5491 0.4505
R30474 DVDD.n9839 DVDD.n9838 0.4505
R30475 DVDD.n9843 DVDD.n9842 0.4505
R30476 DVDD.n9845 DVDD.n9844 0.4505
R30477 DVDD.n9847 DVDD.n9846 0.4505
R30478 DVDD.n9835 DVDD.n9834 0.4505
R30479 DVDD.n9852 DVDD.n9851 0.4505
R30480 DVDD.n9854 DVDD.n9853 0.4505
R30481 DVDD.n9856 DVDD.n9855 0.4505
R30482 DVDD.n9832 DVDD.n9831 0.4505
R30483 DVDD.n9861 DVDD.n9860 0.4505
R30484 DVDD.n9863 DVDD.n9862 0.4505
R30485 DVDD.n9865 DVDD.n9864 0.4505
R30486 DVDD.n9829 DVDD.n9828 0.4505
R30487 DVDD.n9871 DVDD.n9870 0.4505
R30488 DVDD.n9872 DVDD.n9826 0.4505
R30489 DVDD.n9874 DVDD.n9873 0.4505
R30490 DVDD.n9876 DVDD.n9875 0.4505
R30491 DVDD.n9878 DVDD.n9877 0.4505
R30492 DVDD.n9824 DVDD.n9823 0.4505
R30493 DVDD.n9883 DVDD.n9882 0.4505
R30494 DVDD.n9885 DVDD.n9884 0.4505
R30495 DVDD.n9887 DVDD.n9886 0.4505
R30496 DVDD.n9821 DVDD.n9820 0.4505
R30497 DVDD.n9892 DVDD.n9891 0.4505
R30498 DVDD.n9894 DVDD.n9893 0.4505
R30499 DVDD.n9896 DVDD.n9895 0.4505
R30500 DVDD.n9817 DVDD.n9814 0.4505
R30501 DVDD.n9937 DVDD.n9936 0.4505
R30502 DVDD.n9818 DVDD.n9773 0.4505
R30503 DVDD.n9932 DVDD.n9807 0.4505
R30504 DVDD.n9931 DVDD.n9930 0.4505
R30505 DVDD.n9929 DVDD.n9900 0.4505
R30506 DVDD.n9928 DVDD.n9927 0.4505
R30507 DVDD.n9902 DVDD.n9901 0.4505
R30508 DVDD.n9923 DVDD.n9922 0.4505
R30509 DVDD.n9921 DVDD.n9920 0.4505
R30510 DVDD.n9919 DVDD.n9918 0.4505
R30511 DVDD.n9906 DVDD.n9905 0.4505
R30512 DVDD.n9914 DVDD.n9913 0.4505
R30513 DVDD.n9912 DVDD.n9911 0.4505
R30514 DVDD.n9910 DVDD.n9909 0.4505
R30515 DVDD.n9644 DVDD.n9643 0.4505
R30516 DVDD.n10090 DVDD.n10089 0.4505
R30517 DVDD.n9650 DVDD.n9649 0.4505
R30518 DVDD.n10085 DVDD.n10084 0.4505
R30519 DVDD.n10083 DVDD.n9626 0.4505
R30520 DVDD.n10082 DVDD.n9632 0.4505
R30521 DVDD.n9656 DVDD.n9653 0.4505
R30522 DVDD.n10078 DVDD.n10077 0.4505
R30523 DVDD.n10076 DVDD.n9655 0.4505
R30524 DVDD.n10075 DVDD.n10074 0.4505
R30525 DVDD.n9658 DVDD.n9657 0.4505
R30526 DVDD.n10070 DVDD.n10069 0.4505
R30527 DVDD.n9667 DVDD.n9660 0.4505
R30528 DVDD.n9708 DVDD.n9707 0.4505
R30529 DVDD.n9710 DVDD.n9709 0.4505
R30530 DVDD.n9705 DVDD.n9704 0.4505
R30531 DVDD.n9715 DVDD.n9714 0.4505
R30532 DVDD.n9717 DVDD.n9716 0.4505
R30533 DVDD.n9719 DVDD.n9718 0.4505
R30534 DVDD.n9702 DVDD.n9701 0.4505
R30535 DVDD.n9724 DVDD.n9723 0.4505
R30536 DVDD.n9726 DVDD.n9725 0.4505
R30537 DVDD.n9728 DVDD.n9727 0.4505
R30538 DVDD.n9698 DVDD.n9696 0.4505
R30539 DVDD.n10065 DVDD.n10064 0.4505
R30540 DVDD.n9699 DVDD.n9697 0.4505
R30541 DVDD.n10060 DVDD.n10059 0.4505
R30542 DVDD.n10058 DVDD.n9732 0.4505
R30543 DVDD.n9975 DVDD.n9738 0.4505
R30544 DVDD.n9979 DVDD.n9978 0.4505
R30545 DVDD.n9981 DVDD.n9980 0.4505
R30546 DVDD.n9983 DVDD.n9982 0.4505
R30547 DVDD.n9973 DVDD.n9972 0.4505
R30548 DVDD.n9988 DVDD.n9987 0.4505
R30549 DVDD.n9990 DVDD.n9989 0.4505
R30550 DVDD.n9992 DVDD.n9991 0.4505
R30551 DVDD.n9970 DVDD.n9969 0.4505
R30552 DVDD.n9997 DVDD.n9996 0.4505
R30553 DVDD.n10003 DVDD.n10002 0.4505
R30554 DVDD.n10005 DVDD.n10004 0.4505
R30555 DVDD.n9966 DVDD.n9964 0.4505
R30556 DVDD.n10054 DVDD.n10053 0.4505
R30557 DVDD.n9967 DVDD.n9965 0.4505
R30558 DVDD.n10049 DVDD.n10048 0.4505
R30559 DVDD.n10047 DVDD.n10046 0.4505
R30560 DVDD.n10045 DVDD.n800 0.4505
R30561 DVDD.n10009 DVDD.n805 0.4505
R30562 DVDD.n4345 DVDD.n4344 0.4505
R30563 DVDD.n21685 DVDD.n21684 0.4505
R30564 DVDD.n18534 DVDD.n18532 0.4505
R30565 DVDD.n18539 DVDD.n18527 0.4505
R30566 DVDD.n21671 DVDD.n21670 0.4505
R30567 DVDD.n21672 DVDD.n18520 0.4505
R30568 DVDD.n18376 DVDD.n18375 0.4505
R30569 DVDD.n18307 DVDD.n18294 0.4505
R30570 DVDD.n18323 DVDD.n18314 0.4505
R30571 DVDD.n18365 DVDD.n18286 0.4505
R30572 DVDD.n18364 DVDD.n18363 0.4505
R30573 DVDD.n18315 DVDD.n18281 0.4505
R30574 DVDD.n18340 DVDD.n18339 0.4505
R30575 DVDD.n18331 DVDD.n18272 0.4505
R30576 DVDD.n18351 DVDD.n18350 0.4505
R30577 DVDD.n18332 DVDD.n18267 0.4505
R30578 DVDD.n21997 DVDD.n21983 0.4505
R30579 DVDD.n21990 DVDD.n21989 0.4505
R30580 DVDD.n22009 DVDD.n22008 0.4505
R30581 DVDD.n21991 DVDD.n228 0.4505
R30582 DVDD.n22186 DVDD.n229 0.4505
R30583 DVDD.n21271 DVDD.n18655 0.4505
R30584 DVDD.n21220 DVDD.n18654 0.4505
R30585 DVDD.n21233 DVDD.n21222 0.4505
R30586 DVDD.n21223 DVDD.n18660 0.4505
R30587 DVDD.n21260 DVDD.n21259 0.4505
R30588 DVDD.n21359 DVDD.n21357 0.4505
R30589 DVDD.n21360 DVDD.n18548 0.4505
R30590 DVDD.n21654 DVDD.n18549 0.4505
R30591 DVDD.n21369 DVDD.n21332 0.4505
R30592 DVDD.n21331 DVDD.n18533 0.4505
R30593 DVDD.n22069 DVDD.n18205 0.4505
R30594 DVDD.n22058 DVDD.n18204 0.4505
R30595 DVDD.n22062 DVDD.n22061 0.4505
R30596 DVDD.n18231 DVDD.n18212 0.4505
R30597 DVDD.n22045 DVDD.n22044 0.4505
R30598 DVDD.n21919 DVDD.n21918 0.4505
R30599 DVDD.n21830 DVDD.n21798 0.4505
R30600 DVDD.n21898 DVDD.n21897 0.4505
R30601 DVDD.n21899 DVDD.n21791 0.4505
R30602 DVDD.n21930 DVDD.n21790 0.4505
R30603 DVDD.n21931 DVDD.n21789 0.4505
R30604 DVDD.n21932 DVDD.n21788 0.4505
R30605 DVDD.n21876 DVDD.n21787 0.4505
R30606 DVDD.n21879 DVDD.n21780 0.4505
R30607 DVDD.n21942 DVDD.n21779 0.4505
R30608 DVDD.n21778 DVDD.n18387 0.4505
R30609 DVDD.n21760 DVDD.n18386 0.4505
R30610 DVDD.n21767 DVDD.n21763 0.4505
R30611 DVDD.n21768 DVDD.n18394 0.4505
R30612 DVDD.n21769 DVDD.n18393 0.4505
R30613 DVDD.n21736 DVDD.n18392 0.4505
R30614 DVDD.n22240 DVDD.n22239 0.4505
R30615 DVDD.n18476 DVDD.n129 0.4505
R30616 DVDD.n18483 DVDD.n18482 0.4505
R30617 DVDD.n18480 DVDD.n18457 0.4505
R30618 DVDD.n18498 DVDD.n157 0.4505
R30619 DVDD.n22227 DVDD.n22226 0.4505
R30620 DVDD.n22223 DVDD.n158 0.4505
R30621 DVDD.n18427 DVDD.n166 0.4505
R30622 DVDD.n21735 DVDD.n21734 0.4505
R30623 DVDD.n22346 DVDD.n22345 0.4505
R30624 DVDD.n20 DVDD.n2 0.4505
R30625 DVDD.n22351 DVDD.n22350 0.4505
R30626 DVDD.n22318 DVDD.n22317 0.4505
R30627 DVDD.n22320 DVDD.n22319 0.4505
R30628 DVDD.n22322 DVDD.n22321 0.4505
R30629 DVDD.n22314 DVDD.n22313 0.4505
R30630 DVDD.n22326 DVDD.n22315 0.4505
R30631 DVDD.n22328 DVDD.n22327 0.4505
R30632 DVDD.n22330 DVDD.n22329 0.4505
R30633 DVDD.n35 DVDD.n34 0.4505
R30634 DVDD.n22335 DVDD.n22334 0.4505
R30635 DVDD.n33 DVDD.n27 0.4505
R30636 DVDD.n22309 DVDD.n22308 0.4505
R30637 DVDD.n22307 DVDD.n37 0.4505
R30638 DVDD.n22306 DVDD.n22305 0.4505
R30639 DVDD.n39 DVDD.n38 0.4505
R30640 DVDD.n22301 DVDD.n22300 0.4505
R30641 DVDD.n64 DVDD.n41 0.4505
R30642 DVDD.n22275 DVDD.n22274 0.4505
R30643 DVDD.n22272 DVDD.n22271 0.4505
R30644 DVDD.n22279 DVDD.n22273 0.4505
R30645 DVDD.n22281 DVDD.n22280 0.4505
R30646 DVDD.n22283 DVDD.n22282 0.4505
R30647 DVDD.n22268 DVDD.n22267 0.4505
R30648 DVDD.n22287 DVDD.n22269 0.4505
R30649 DVDD.n22289 DVDD.n22288 0.4505
R30650 DVDD.n22291 DVDD.n22290 0.4505
R30651 DVDD.n82 DVDD.n81 0.4505
R30652 DVDD.n22296 DVDD.n22295 0.4505
R30653 DVDD.n80 DVDD.n79 0.4505
R30654 DVDD.n22263 DVDD.n22262 0.4505
R30655 DVDD.n22261 DVDD.n84 0.4505
R30656 DVDD.n22260 DVDD.n22259 0.4505
R30657 DVDD.n93 DVDD.n86 0.4505
R30658 DVDD.n22255 DVDD.n22254 0.4505
R30659 DVDD.n105 DVDD.n88 0.4505
R30660 DVDD.n21129 DVDD.n21128 0.4505
R30661 DVDD.n21133 DVDD.n21130 0.4505
R30662 DVDD.n21135 DVDD.n21134 0.4505
R30663 DVDD.n21137 DVDD.n21136 0.4505
R30664 DVDD.n21125 DVDD.n21124 0.4505
R30665 DVDD.n21141 DVDD.n21126 0.4505
R30666 DVDD.n21143 DVDD.n21142 0.4505
R30667 DVDD.n21145 DVDD.n21144 0.4505
R30668 DVDD.n21122 DVDD.n21121 0.4505
R30669 DVDD.n21149 DVDD.n118 0.4505
R30670 DVDD.n21150 DVDD.n112 0.4505
R30671 DVDD.n21152 DVDD.n21151 0.4505
R30672 DVDD.n21118 DVDD.n21117 0.4505
R30673 DVDD.n21157 DVDD.n21156 0.4505
R30674 DVDD.n21158 DVDD.n21116 0.4505
R30675 DVDD.n21160 DVDD.n21159 0.4505
R30676 DVDD.n21162 DVDD.n21161 0.4505
R30677 DVDD.n21113 DVDD.n21112 0.4505
R30678 DVDD.n21166 DVDD.n21114 0.4505
R30679 DVDD.n21168 DVDD.n21167 0.4505
R30680 DVDD.n21170 DVDD.n21169 0.4505
R30681 DVDD.n21109 DVDD.n21108 0.4505
R30682 DVDD.n21174 DVDD.n21110 0.4505
R30683 DVDD.n21176 DVDD.n21175 0.4505
R30684 DVDD.n21178 DVDD.n21177 0.4505
R30685 DVDD.n21103 DVDD.n21102 0.4505
R30686 DVDD.n21183 DVDD.n21182 0.4505
R30687 DVDD.n21101 DVDD.n21100 0.4505
R30688 DVDD.n21104 DVDD.n18729 0.4505
R30689 DVDD.n21187 DVDD.n18722 0.4505
R30690 DVDD.n21189 DVDD.n21188 0.4505
R30691 DVDD.n18723 DVDD.n18719 0.4505
R30692 DVDD.n21193 DVDD.n18720 0.4505
R30693 DVDD.n21195 DVDD.n21194 0.4505
R30694 DVDD.n21197 DVDD.n21196 0.4505
R30695 DVDD.n18716 DVDD.n18715 0.4505
R30696 DVDD.n21201 DVDD.n18717 0.4505
R30697 DVDD.n21203 DVDD.n21202 0.4505
R30698 DVDD.n21205 DVDD.n21204 0.4505
R30699 DVDD.n18712 DVDD.n18711 0.4505
R30700 DVDD.n21210 DVDD.n21209 0.4505
R30701 DVDD.n18710 DVDD.n18709 0.4505
R30702 DVDD.n19675 DVDD.n19674 0.4505
R30703 DVDD.n19679 DVDD.n19676 0.4505
R30704 DVDD.n19681 DVDD.n19680 0.4505
R30705 DVDD.n19682 DVDD.n18691 0.4505
R30706 DVDD.n19671 DVDD.n18685 0.4505
R30707 DVDD.n19687 DVDD.n19686 0.4505
R30708 DVDD.n19688 DVDD.n19670 0.4505
R30709 DVDD.n19690 DVDD.n19689 0.4505
R30710 DVDD.n19691 DVDD.n19207 0.4505
R30711 DVDD.n19640 DVDD.n19201 0.4505
R30712 DVDD.n19696 DVDD.n19695 0.4505
R30713 DVDD.n19639 DVDD.n19638 0.4505
R30714 DVDD.n19666 DVDD.n19665 0.4505
R30715 DVDD.n19664 DVDD.n19663 0.4505
R30716 DVDD.n19662 DVDD.n19644 0.4505
R30717 DVDD.n19643 DVDD.n19642 0.4505
R30718 DVDD.n19658 DVDD.n19657 0.4505
R30719 DVDD.n19656 DVDD.n19655 0.4505
R30720 DVDD.n19649 DVDD.n19648 0.4505
R30721 DVDD.n19647 DVDD.n19646 0.4505
R30722 DVDD.n19656 DVDD.n19645 0.4505
R30723 DVDD.n19659 DVDD.n19658 0.4505
R30724 DVDD.n19660 DVDD.n19643 0.4505
R30725 DVDD.n19662 DVDD.n19661 0.4505
R30726 DVDD.n19664 DVDD.n19641 0.4505
R30727 DVDD.n19667 DVDD.n19666 0.4505
R30728 DVDD.n19668 DVDD.n19639 0.4505
R30729 DVDD.n19695 DVDD.n19694 0.4505
R30730 DVDD.n19693 DVDD.n19640 0.4505
R30731 DVDD.n19692 DVDD.n19691 0.4505
R30732 DVDD.n19690 DVDD.n19669 0.4505
R30733 DVDD.n19672 DVDD.n19670 0.4505
R30734 DVDD.n19686 DVDD.n19685 0.4505
R30735 DVDD.n19684 DVDD.n19671 0.4505
R30736 DVDD.n19683 DVDD.n19682 0.4505
R30737 DVDD.n19681 DVDD.n19673 0.4505
R30738 DVDD.n19679 DVDD.n19678 0.4505
R30739 DVDD.n19677 DVDD.n19675 0.4505
R30740 DVDD.n18713 DVDD.n18710 0.4505
R30741 DVDD.n21209 DVDD.n21208 0.4505
R30742 DVDD.n21207 DVDD.n18712 0.4505
R30743 DVDD.n21206 DVDD.n21205 0.4505
R30744 DVDD.n21203 DVDD.n18714 0.4505
R30745 DVDD.n21201 DVDD.n21200 0.4505
R30746 DVDD.n21199 DVDD.n18716 0.4505
R30747 DVDD.n21198 DVDD.n21197 0.4505
R30748 DVDD.n21195 DVDD.n18718 0.4505
R30749 DVDD.n21193 DVDD.n21192 0.4505
R30750 DVDD.n21191 DVDD.n18719 0.4505
R30751 DVDD.n21190 DVDD.n21189 0.4505
R30752 DVDD.n18722 DVDD.n18721 0.4505
R30753 DVDD.n21105 DVDD.n21104 0.4505
R30754 DVDD.n21106 DVDD.n21101 0.4505
R30755 DVDD.n21182 DVDD.n21181 0.4505
R30756 DVDD.n21180 DVDD.n21103 0.4505
R30757 DVDD.n21179 DVDD.n21178 0.4505
R30758 DVDD.n21176 DVDD.n21107 0.4505
R30759 DVDD.n21174 DVDD.n21173 0.4505
R30760 DVDD.n21172 DVDD.n21109 0.4505
R30761 DVDD.n21171 DVDD.n21170 0.4505
R30762 DVDD.n21168 DVDD.n21111 0.4505
R30763 DVDD.n21166 DVDD.n21165 0.4505
R30764 DVDD.n21164 DVDD.n21113 0.4505
R30765 DVDD.n21163 DVDD.n21162 0.4505
R30766 DVDD.n21160 DVDD.n21115 0.4505
R30767 DVDD.n21119 DVDD.n21116 0.4505
R30768 DVDD.n21156 DVDD.n21155 0.4505
R30769 DVDD.n21154 DVDD.n21118 0.4505
R30770 DVDD.n21153 DVDD.n21152 0.4505
R30771 DVDD.n21150 DVDD.n21120 0.4505
R30772 DVDD.n21149 DVDD.n21148 0.4505
R30773 DVDD.n21147 DVDD.n21122 0.4505
R30774 DVDD.n21146 DVDD.n21145 0.4505
R30775 DVDD.n21143 DVDD.n21123 0.4505
R30776 DVDD.n21141 DVDD.n21140 0.4505
R30777 DVDD.n21139 DVDD.n21125 0.4505
R30778 DVDD.n21138 DVDD.n21137 0.4505
R30779 DVDD.n21135 DVDD.n21127 0.4505
R30780 DVDD.n21133 DVDD.n21132 0.4505
R30781 DVDD.n21131 DVDD.n21129 0.4505
R30782 DVDD.n88 DVDD.n87 0.4505
R30783 DVDD.n22256 DVDD.n22255 0.4505
R30784 DVDD.n22257 DVDD.n86 0.4505
R30785 DVDD.n22259 DVDD.n22258 0.4505
R30786 DVDD.n84 DVDD.n83 0.4505
R30787 DVDD.n22264 DVDD.n22263 0.4505
R30788 DVDD.n22265 DVDD.n80 0.4505
R30789 DVDD.n22295 DVDD.n22294 0.4505
R30790 DVDD.n22293 DVDD.n82 0.4505
R30791 DVDD.n22292 DVDD.n22291 0.4505
R30792 DVDD.n22289 DVDD.n22266 0.4505
R30793 DVDD.n22287 DVDD.n22286 0.4505
R30794 DVDD.n22285 DVDD.n22268 0.4505
R30795 DVDD.n22284 DVDD.n22283 0.4505
R30796 DVDD.n22281 DVDD.n22270 0.4505
R30797 DVDD.n22279 DVDD.n22278 0.4505
R30798 DVDD.n22277 DVDD.n22272 0.4505
R30799 DVDD.n22276 DVDD.n22275 0.4505
R30800 DVDD.n41 DVDD.n40 0.4505
R30801 DVDD.n22302 DVDD.n22301 0.4505
R30802 DVDD.n22303 DVDD.n39 0.4505
R30803 DVDD.n22305 DVDD.n22304 0.4505
R30804 DVDD.n37 DVDD.n36 0.4505
R30805 DVDD.n22310 DVDD.n22309 0.4505
R30806 DVDD.n22311 DVDD.n33 0.4505
R30807 DVDD.n22334 DVDD.n22333 0.4505
R30808 DVDD.n22332 DVDD.n35 0.4505
R30809 DVDD.n22331 DVDD.n22330 0.4505
R30810 DVDD.n22328 DVDD.n22312 0.4505
R30811 DVDD.n22326 DVDD.n22325 0.4505
R30812 DVDD.n22324 DVDD.n22314 0.4505
R30813 DVDD.n22323 DVDD.n22322 0.4505
R30814 DVDD.n22320 DVDD.n22316 0.4505
R30815 DVDD.n22318 DVDD.n3 0.4505
R30816 DVDD.n22350 DVDD.n22349 0.4505
R30817 DVDD.n22348 DVDD.n2 0.4505
R30818 DVDD.n19651 DVDD.n19647 0.4505
R30819 DVDD.n19654 DVDD.n19652 0.4505
R30820 DVDD.n19654 DVDD.n19653 0.4505
R30821 DVDD.n19417 DVDD 0.386971
R30822 DVDD.n21925 DVDD.n21792 0.384978
R30823 DVDD.n21772 DVDD.n21771 0.384978
R30824 DVDD.n18119 DVDD.n18064 0.384022
R30825 DVDD.n22234 DVDD.n130 0.383973
R30826 DVDD.n21731 DVDD.n21730 0.383973
R30827 DVDD.n22067 DVDD.n22066 0.383973
R30828 DVDD.n21937 DVDD.n21936 0.383973
R30829 DVDD.n18109 DVDD.n18099 0.383973
R30830 DVDD.n21371 DVDD.n21370 0.3755
R30831 DVDD.n19633 DVDD.n19632 0.3755
R30832 DVDD.n19425 DVDD.n13 0.3755
R30833 DVDD.n4372 DVDD.n4371 0.3755
R30834 DVDD.n20933 DVDD.n20932 0.365842
R30835 DVDD.n19105 DVDD.n19104 0.365842
R30836 DVDD.n20973 DVDD.n18830 0.365842
R30837 DVDD.n20967 DVDD.n20966 0.365842
R30838 DVDD.n4336 DVDD.t23 0.3645
R30839 DVDD.n4336 DVDD.t37 0.3645
R30840 DVDD.n4333 DVDD.t53 0.3645
R30841 DVDD.n4333 DVDD.t41 0.3645
R30842 DVDD.n4383 DVDD.t27 0.3645
R30843 DVDD.n4383 DVDD.t19 0.3645
R30844 DVDD.n4355 DVDD.t59 0.3645
R30845 DVDD.n4355 DVDD.t57 0.3645
R30846 DVDD.n4356 DVDD.t47 0.3645
R30847 DVDD.n4356 DVDD.t39 0.3645
R30848 DVDD.n4358 DVDD.t43 0.3645
R30849 DVDD.n4358 DVDD.t15 0.3645
R30850 DVDD.n4360 DVDD.t21 0.3645
R30851 DVDD.n4360 DVDD.t45 0.3645
R30852 DVDD.n4363 DVDD.t49 0.3645
R30853 DVDD.n4363 DVDD.t29 0.3645
R30854 DVDD.n4365 DVDD.t25 0.3645
R30855 DVDD.n4365 DVDD.t61 0.3645
R30856 DVDD.n4366 DVDD.t51 0.3645
R30857 DVDD.n4366 DVDD.t33 0.3645
R30858 DVDD.n4368 DVDD.t31 0.3645
R30859 DVDD.n4368 DVDD.t17 0.3645
R30860 DVDD.n4348 DVDD.t3 0.3645
R30861 DVDD.n4348 DVDD.t7 0.3645
R30862 DVDD.n4340 DVDD.t9 0.3645
R30863 DVDD.n4340 DVDD.t5 0.3645
R30864 DVDD.n4342 DVDD.t154 0.3645
R30865 DVDD.n4342 DVDD.t11 0.3645
R30866 DVDD.n22039 DVDD.n218 0.356216
R30867 DVDD.n21944 DVDD.n190 0.35585
R30868 DVDD.n22229 DVDD.n135 0.355277
R30869 DVDD.n4453 DVDD.n4452 0.35492
R30870 DVDD.n21944 DVDD.n187 0.354416
R30871 DVDD.n22229 DVDD.n147 0.35405
R30872 DVDD.n22039 DVDD.n217 0.35405
R30873 DVDD.n4453 DVDD.n4451 0.35312
R30874 DVDD.n4353 DVDD.n4352 0.346654
R30875 DVDD.n22193 DVDD.n218 0.33977
R30876 DVDD.n4452 DVDD.n4415 0.339393
R30877 DVDD.n21721 DVDD.n135 0.339029
R30878 DVDD.n196 DVDD.n187 0.33857
R30879 DVDD.n196 DVDD.n190 0.338454
R30880 DVDD.n4451 DVDD.n4415 0.338193
R30881 DVDD.n21721 DVDD.n147 0.337254
R30882 DVDD.n22193 DVDD.n217 0.337254
R30883 DVDD.n21944 DVDD.n18301 0.3005
R30884 DVDD.n22039 DVDD.n18243 0.3005
R30885 DVDD.n22229 DVDD.n137 0.3005
R30886 DVDD.n22039 DVDD.n18240 0.3005
R30887 DVDD.n21944 DVDD.n21943 0.3005
R30888 DVDD.n22229 DVDD.n22228 0.3005
R30889 DVDD.n22056 DVDD.n315 0.28175
R30890 DVDD.n22057 DVDD.n18220 0.28175
R30891 DVDD.n22049 DVDD.n18217 0.28175
R30892 DVDD.n22051 DVDD.n22050 0.28175
R30893 DVDD.n22048 DVDD.n22047 0.28175
R30894 DVDD.n22039 DVDD.n18225 0.28175
R30895 DVDD.n21916 DVDD.n21915 0.28175
R30896 DVDD.n21914 DVDD.n21913 0.28175
R30897 DVDD.n21804 DVDD.n21803 0.28175
R30898 DVDD.n21815 DVDD.n21814 0.28175
R30899 DVDD.n21902 DVDD.n21809 0.28175
R30900 DVDD.n21859 DVDD.n21858 0.28175
R30901 DVDD.n21874 DVDD.n21857 0.28175
R30902 DVDD.n21863 DVDD.n21843 0.28175
R30903 DVDD.n21864 DVDD.n21841 0.28175
R30904 DVDD.n21866 DVDD.n21865 0.28175
R30905 DVDD.n21944 DVDD.n18382 0.28175
R30906 DVDD.n21758 DVDD.n21757 0.28175
R30907 DVDD.n21756 DVDD.n18400 0.28175
R30908 DVDD.n21755 DVDD.n18398 0.28175
R30909 DVDD.n21754 DVDD.n21753 0.28175
R30910 DVDD.n18404 DVDD.n18403 0.28175
R30911 DVDD.n21738 DVDD.n18409 0.28175
R30912 DVDD.n21594 DVDD.n18408 0.28175
R30913 DVDD.n21593 DVDD.n21592 0.28175
R30914 DVDD.n21583 DVDD.n164 0.28175
R30915 DVDD.n21582 DVDD.n162 0.28175
R30916 DVDD.n22229 DVDD.n150 0.28175
R30917 DVDD.n18496 DVDD.n18495 0.28175
R30918 DVDD.n18494 DVDD.n18493 0.28175
R30919 DVDD.n18485 DVDD.n18461 0.28175
R30920 DVDD.n18462 DVDD.n121 0.28175
R30921 DVDD.n22243 DVDD.n22242 0.28175
R30922 DVDD.n22039 DVDD.n18228 0.28175
R30923 DVDD.n21944 DVDD.n18298 0.28175
R30924 DVDD.n22229 DVDD.n156 0.28175
R30925 DVDD.n22184 DVDD.n22183 0.28175
R30926 DVDD.n235 DVDD.n233 0.28175
R30927 DVDD.n22024 DVDD.n21987 0.28175
R30928 DVDD.n22034 DVDD.n22033 0.28175
R30929 DVDD.n22036 DVDD.n22035 0.28175
R30930 DVDD.n22039 DVDD.n18265 0.28175
R30931 DVDD.n21981 DVDD.n21980 0.28175
R30932 DVDD.n21979 DVDD.n21978 0.28175
R30933 DVDD.n21977 DVDD.n21976 0.28175
R30934 DVDD.n18270 DVDD.n18269 0.28175
R30935 DVDD.n21966 DVDD.n21965 0.28175
R30936 DVDD.n21964 DVDD.n21963 0.28175
R30937 DVDD.n21962 DVDD.n21961 0.28175
R30938 DVDD.n18284 DVDD.n18283 0.28175
R30939 DVDD.n21949 DVDD.n21948 0.28175
R30940 DVDD.n21947 DVDD.n21946 0.28175
R30941 DVDD.n21945 DVDD.n21944 0.28175
R30942 DVDD.n21705 DVDD.n18296 0.28175
R30943 DVDD.n21690 DVDD.n18518 0.28175
R30944 DVDD.n21692 DVDD.n21691 0.28175
R30945 DVDD.n21689 DVDD.n21688 0.28175
R30946 DVDD.n21687 DVDD.n18529 0.28175
R30947 DVDD.n21648 DVDD.n21647 0.28175
R30948 DVDD.n21650 DVDD.n21649 0.28175
R30949 DVDD.n21652 DVDD.n21651 0.28175
R30950 DVDD.n18556 DVDD.n18555 0.28175
R30951 DVDD.n21355 DVDD.n21354 0.28175
R30952 DVDD.n22229 DVDD.n136 0.28175
R30953 DVDD.n21257 DVDD.n21256 0.28175
R30954 DVDD.n21255 DVDD.n21254 0.28175
R30955 DVDD.n18666 DVDD.n18665 0.28175
R30956 DVDD.n21216 DVDD.n21215 0.28175
R30957 DVDD.n21248 DVDD.n18671 0.28175
R30958 DVDD.n22039 DVDD.n22038 0.28175
R30959 DVDD.n21944 DVDD.n18384 0.28175
R30960 DVDD.n22229 DVDD.n145 0.28175
R30961 DVDD.n3977 DVDD.n3578 0.244637
R30962 DVDD.n18199 DVDD.n18198 0.244637
R30963 DVDD.n19504 DVDD.n19503 0.237342
R30964 DVDD.n21596 DVDD.n21595 0.237342
R30965 DVDD.n19289 DVDD.n19288 0.237342
R30966 DVDD.n18595 DVDD.n18410 0.237342
R30967 DVDD.n19554 DVDD.n19553 0.237342
R30968 DVDD.n21646 DVDD.n21645 0.237342
R30969 DVDD.n19236 DVDD.n19235 0.237342
R30970 DVDD.n21442 DVDD.n21441 0.237342
R30971 DVDD.n19650 DVDD.n19194 0.235287
R30972 DVDD.n22347 DVDD.n4 0.23503
R30973 DVDD.n20140 DVDD.n20122 0.234541
R30974 DVDD.n20627 DVDD.n20609 0.234541
R30975 DVDD.n3976 DVDD.n3934 0.234541
R30976 DVDD.n15285 DVDD.n5486 0.234541
R30977 DVDD.n20883 DVDD.n18950 0.234284
R30978 DVDD.n20854 DVDD.n18979 0.234284
R30979 DVDD.n22120 DVDD.n22119 0.234284
R30980 DVDD.n10018 DVDD.n796 0.234284
R30981 DVDD.n20534 DVDD.n20532 0.22775
R30982 DVDD.n20925 DVDD.n18907 0.22775
R30983 DVDD.n21058 DVDD.n18762 0.22775
R30984 DVDD.n19100 DVDD.n19098 0.22775
R30985 DVDD.n22159 DVDD.n298 0.226773
R30986 DVDD.n4658 DVDD.n361 0.226773
R30987 DVDD.n4178 DVDD.n260 0.226773
R30988 DVDD.n4136 DVDD.n4066 0.226773
R30989 DVDD.n22240 DVDD.n126 0.218099
R30990 DVDD.n21249 DVDD.n21248 0.218099
R30991 DVDD.n21228 DVDD.n18655 0.218099
R30992 DVDD.n22242 DVDD.n122 0.218099
R30993 DVDD.n22187 DVDD.n22186 0.217859
R30994 DVDD.n22184 DVDD.n234 0.217859
R30995 DVDD.n18235 DVDD.n18205 0.217859
R30996 DVDD.n22056 DVDD.n22055 0.217859
R30997 DVDD.n21661 DVDD.n18531 0.214786
R30998 DVDD.n21663 DVDD.n21662 0.214786
R30999 DVDD.n18541 DVDD.n18540 0.214786
R31000 DVDD.n21669 DVDD.n21668 0.214786
R31001 DVDD.n18303 DVDD.n185 0.214786
R31002 DVDD.n18377 DVDD.n186 0.214786
R31003 DVDD.n18322 DVDD.n18306 0.214786
R31004 DVDD.n18325 DVDD.n18324 0.214786
R31005 DVDD.n18318 DVDD.n18316 0.214786
R31006 DVDD.n18362 DVDD.n18361 0.214786
R31007 DVDD.n18319 DVDD.n18317 0.214786
R31008 DVDD.n18357 DVDD.n18329 0.214786
R31009 DVDD.n18356 DVDD.n18330 0.214786
R31010 DVDD.n18355 DVDD.n18352 0.214786
R31011 DVDD.n18353 DVDD.n18248 0.214786
R31012 DVDD.n22191 DVDD.n224 0.214786
R31013 DVDD.n22190 DVDD.n225 0.214786
R31014 DVDD.n22189 DVDD.n226 0.214786
R31015 DVDD.n21988 DVDD.n227 0.214786
R31016 DVDD.n18546 DVDD.n142 0.214786
R31017 DVDD.n21226 DVDD.n139 0.214786
R31018 DVDD.n21227 DVDD.n18661 0.214786
R31019 DVDD.n21232 DVDD.n21231 0.214786
R31020 DVDD.n21225 DVDD.n21224 0.214786
R31021 DVDD.n21339 DVDD.n18547 0.214786
R31022 DVDD.n21656 DVDD.n21655 0.214786
R31023 DVDD.n18550 DVDD.n18543 0.214786
R31024 DVDD.n21660 DVDD.n18544 0.214786
R31025 DVDD.n21658 DVDD.n18543 0.214786
R31026 DVDD.n21657 DVDD.n21656 0.214786
R31027 DVDD.n18547 DVDD.n18545 0.214786
R31028 DVDD.n18546 DVDD.n18504 0.214786
R31029 DVDD.n21226 DVDD.n18505 0.214786
R31030 DVDD.n21229 DVDD.n21227 0.214786
R31031 DVDD.n21231 DVDD.n21230 0.214786
R31032 DVDD.n21661 DVDD.n18542 0.214786
R31033 DVDD.n21664 DVDD.n21663 0.214786
R31034 DVDD.n21665 DVDD.n18541 0.214786
R31035 DVDD.n21668 DVDD.n21667 0.214786
R31036 DVDD.n21666 DVDD.n185 0.214786
R31037 DVDD.n18320 DVDD.n186 0.214786
R31038 DVDD.n18322 DVDD.n18321 0.214786
R31039 DVDD.n18326 DVDD.n18325 0.214786
R31040 DVDD.n18327 DVDD.n18318 0.214786
R31041 DVDD.n18361 DVDD.n18360 0.214786
R31042 DVDD.n18359 DVDD.n18319 0.214786
R31043 DVDD.n18358 DVDD.n18357 0.214786
R31044 DVDD.n18356 DVDD.n18328 0.214786
R31045 DVDD.n18355 DVDD.n18354 0.214786
R31046 DVDD.n18353 DVDD.n221 0.214786
R31047 DVDD.n22192 DVDD.n22191 0.214786
R31048 DVDD.n22190 DVDD.n222 0.214786
R31049 DVDD.n22189 DVDD.n22188 0.214786
R31050 DVDD.n21660 DVDD.n21659 0.214786
R31051 DVDD.n21712 DVDD.n18514 0.214786
R31052 DVDD.n21711 DVDD.n18515 0.214786
R31053 DVDD.n18528 DVDD.n18516 0.214786
R31054 DVDD.n21707 DVDD.n21706 0.214786
R31055 DVDD.n18300 DVDD.n193 0.214786
R31056 DVDD.n22208 DVDD.n194 0.214786
R31057 DVDD.n18295 DVDD.n195 0.214786
R31058 DVDD.n22204 DVDD.n198 0.214786
R31059 DVDD.n22203 DVDD.n199 0.214786
R31060 DVDD.n22202 DVDD.n200 0.214786
R31061 DVDD.n18282 DVDD.n201 0.214786
R31062 DVDD.n22198 DVDD.n203 0.214786
R31063 DVDD.n22197 DVDD.n204 0.214786
R31064 DVDD.n22196 DVDD.n205 0.214786
R31065 DVDD.n18242 DVDD.n206 0.214786
R31066 DVDD.n22025 DVDD.n18249 0.214786
R31067 DVDD.n22026 DVDD.n21986 0.214786
R31068 DVDD.n22032 DVDD.n22031 0.214786
R31069 DVDD.n22028 DVDD.n22027 0.214786
R31070 DVDD.n21719 DVDD.n144 0.214786
R31071 DVDD.n18668 DVDD.n146 0.214786
R31072 DVDD.n18669 DVDD.n18664 0.214786
R31073 DVDD.n21253 DVDD.n21252 0.214786
R31074 DVDD.n18670 DVDD.n18667 0.214786
R31075 DVDD.n21718 DVDD.n18509 0.214786
R31076 DVDD.n21717 DVDD.n18510 0.214786
R31077 DVDD.n18554 DVDD.n18511 0.214786
R31078 DVDD.n21713 DVDD.n18513 0.214786
R31079 DVDD.n21715 DVDD.n18511 0.214786
R31080 DVDD.n21717 DVDD.n21716 0.214786
R31081 DVDD.n21718 DVDD.n18508 0.214786
R31082 DVDD.n21720 DVDD.n21719 0.214786
R31083 DVDD.n18668 DVDD.n18507 0.214786
R31084 DVDD.n21250 DVDD.n18669 0.214786
R31085 DVDD.n21252 DVDD.n21251 0.214786
R31086 DVDD.n21714 DVDD.n21713 0.214786
R31087 DVDD.n21712 DVDD.n18512 0.214786
R31088 DVDD.n21711 DVDD.n21710 0.214786
R31089 DVDD.n21709 DVDD.n18516 0.214786
R31090 DVDD.n21708 DVDD.n21707 0.214786
R31091 DVDD.n18517 DVDD.n193 0.214786
R31092 DVDD.n22208 DVDD.n22207 0.214786
R31093 DVDD.n22206 DVDD.n195 0.214786
R31094 DVDD.n22205 DVDD.n22204 0.214786
R31095 DVDD.n22203 DVDD.n197 0.214786
R31096 DVDD.n22202 DVDD.n22201 0.214786
R31097 DVDD.n22200 DVDD.n201 0.214786
R31098 DVDD.n22199 DVDD.n22198 0.214786
R31099 DVDD.n22197 DVDD.n202 0.214786
R31100 DVDD.n22196 DVDD.n22195 0.214786
R31101 DVDD.n22194 DVDD.n206 0.214786
R31102 DVDD.n22025 DVDD.n219 0.214786
R31103 DVDD.n22029 DVDD.n22026 0.214786
R31104 DVDD.n22031 DVDD.n22030 0.214786
R31105 DVDD.n22216 DVDD.n172 0.214786
R31106 DVDD.n22215 DVDD.n173 0.214786
R31107 DVDD.n18395 DVDD.n174 0.214786
R31108 DVDD.n22211 DVDD.n176 0.214786
R31109 DVDD.n22210 DVDD.n177 0.214786
R31110 DVDD.n18299 DVDD.n181 0.214786
R31111 DVDD.n21881 DVDD.n21880 0.214786
R31112 DVDD.n21838 DVDD.n21835 0.214786
R31113 DVDD.n21885 DVDD.n21836 0.214786
R31114 DVDD.n21887 DVDD.n21886 0.214786
R31115 DVDD.n21889 DVDD.n21888 0.214786
R31116 DVDD.n21831 DVDD.n21829 0.214786
R31117 DVDD.n21895 DVDD.n21894 0.214786
R31118 DVDD.n21833 DVDD.n21799 0.214786
R31119 DVDD.n21832 DVDD.n18241 0.214786
R31120 DVDD.n18232 DVDD.n18230 0.214786
R31121 DVDD.n18239 DVDD.n18238 0.214786
R31122 DVDD.n18233 DVDD.n18213 0.214786
R31123 DVDD.n18234 DVDD.n18214 0.214786
R31124 DVDD.n18451 DVDD.n154 0.214786
R31125 DVDD.n18501 DVDD.n148 0.214786
R31126 DVDD.n18500 DVDD.n18499 0.214786
R31127 DVDD.n18477 DVDD.n18456 0.214786
R31128 DVDD.n18454 DVDD.n127 0.214786
R31129 DVDD.n167 DVDD.n160 0.214786
R31130 DVDD.n22222 DVDD.n22221 0.214786
R31131 DVDD.n18425 DVDD.n168 0.214786
R31132 DVDD.n22217 DVDD.n171 0.214786
R31133 DVDD.n22219 DVDD.n168 0.214786
R31134 DVDD.n22221 DVDD.n22220 0.214786
R31135 DVDD.n169 DVDD.n167 0.214786
R31136 DVDD.n18452 DVDD.n18451 0.214786
R31137 DVDD.n18502 DVDD.n18501 0.214786
R31138 DVDD.n18500 DVDD.n18453 0.214786
R31139 DVDD.n18456 DVDD.n18455 0.214786
R31140 DVDD.n22218 DVDD.n22217 0.214786
R31141 DVDD.n22216 DVDD.n170 0.214786
R31142 DVDD.n22215 DVDD.n22214 0.214786
R31143 DVDD.n22213 DVDD.n174 0.214786
R31144 DVDD.n22212 DVDD.n22211 0.214786
R31145 DVDD.n22210 DVDD.n175 0.214786
R31146 DVDD.n21837 DVDD.n181 0.214786
R31147 DVDD.n21882 DVDD.n21881 0.214786
R31148 DVDD.n21883 DVDD.n21835 0.214786
R31149 DVDD.n21885 DVDD.n21884 0.214786
R31150 DVDD.n21886 DVDD.n21834 0.214786
R31151 DVDD.n21890 DVDD.n21889 0.214786
R31152 DVDD.n21891 DVDD.n21831 0.214786
R31153 DVDD.n21894 DVDD.n21893 0.214786
R31154 DVDD.n21892 DVDD.n21833 0.214786
R31155 DVDD.n21832 DVDD.n214 0.214786
R31156 DVDD.n18232 DVDD.n215 0.214786
R31157 DVDD.n18238 DVDD.n18237 0.214786
R31158 DVDD.n18236 DVDD.n18233 0.214786
R31159 DVDD.n18407 DVDD.n18406 0.214786
R31160 DVDD.n21589 DVDD.n21588 0.214786
R31161 DVDD.n21587 DVDD.n21586 0.214786
R31162 DVDD.n21584 DVDD.n18449 0.214786
R31163 DVDD.n18489 DVDD.n18450 0.214786
R31164 DVDD.n18490 DVDD.n18488 0.214786
R31165 DVDD.n18491 DVDD.n18487 0.214786
R31166 DVDD.n21742 DVDD.n21741 0.214786
R31167 DVDD.n21743 DVDD.n18405 0.214786
R31168 DVDD.n21751 DVDD.n21744 0.214786
R31169 DVDD.n21750 DVDD.n21745 0.214786
R31170 DVDD.n21748 DVDD.n21747 0.214786
R31171 DVDD.n21746 DVDD.n189 0.214786
R31172 DVDD.n21862 DVDD.n188 0.214786
R31173 DVDD.n21869 DVDD.n21868 0.214786
R31174 DVDD.n21870 DVDD.n21861 0.214786
R31175 DVDD.n21872 DVDD.n21871 0.214786
R31176 DVDD.n21807 DVDD.n21806 0.214786
R31177 DVDD.n21905 DVDD.n21904 0.214786
R31178 DVDD.n21906 DVDD.n21805 0.214786
R31179 DVDD.n21911 DVDD.n21907 0.214786
R31180 DVDD.n21910 DVDD.n21908 0.214786
R31181 DVDD.n21909 DVDD.n211 0.214786
R31182 DVDD.n18226 DVDD.n210 0.214786
R31183 DVDD.n18223 DVDD.n18222 0.214786
R31184 DVDD.n22054 DVDD.n22053 0.214786
R31185 DVDD.n21739 DVDD.n18405 0.214786
R31186 DVDD.n21752 DVDD.n21751 0.214786
R31187 DVDD.n21750 DVDD.n21749 0.214786
R31188 DVDD.n21748 DVDD.n18402 0.214786
R31189 DVDD.n18381 DVDD.n189 0.214786
R31190 DVDD.n18383 DVDD.n188 0.214786
R31191 DVDD.n21868 DVDD.n21867 0.214786
R31192 DVDD.n21861 DVDD.n21860 0.214786
R31193 DVDD.n21873 DVDD.n21872 0.214786
R31194 DVDD.n21808 DVDD.n21807 0.214786
R31195 DVDD.n21904 DVDD.n21903 0.214786
R31196 DVDD.n21810 DVDD.n21805 0.214786
R31197 DVDD.n21912 DVDD.n21911 0.214786
R31198 DVDD.n21910 DVDD.n21802 0.214786
R31199 DVDD.n21909 DVDD.n18264 0.214786
R31200 DVDD.n18227 DVDD.n18226 0.214786
R31201 DVDD.n18224 DVDD.n18223 0.214786
R31202 DVDD.n22053 DVDD.n22052 0.214786
R31203 DVDD.n18221 DVDD.n18219 0.214786
R31204 DVDD.n21584 DVDD.n149 0.214786
R31205 DVDD.n18489 DVDD.n151 0.214786
R31206 DVDD.n18490 DVDD.n18460 0.214786
R31207 DVDD.n18492 DVDD.n18491 0.214786
R31208 DVDD.n18486 DVDD.n123 0.214786
R31209 DVDD.n21586 DVDD.n21585 0.214786
R31210 DVDD.n21590 DVDD.n21589 0.214786
R31211 DVDD.n21591 DVDD.n18407 0.214786
R31212 DVDD.n21741 DVDD.n21740 0.214786
R31213 DVDD.n4803 DVDD.n4802 0.214786
R31214 DVDD.n4801 DVDD.n3579 0.214786
R31215 DVDD.n3581 DVDD.n3580 0.214786
R31216 DVDD.n4797 DVDD.n3583 0.214786
R31217 DVDD.n4796 DVDD.n3584 0.214786
R31218 DVDD.n4795 DVDD.n3585 0.214786
R31219 DVDD.n3587 DVDD.n3586 0.214786
R31220 DVDD.n4791 DVDD.n3589 0.214786
R31221 DVDD.n4790 DVDD.n3590 0.214786
R31222 DVDD.n4789 DVDD.n3591 0.214786
R31223 DVDD.n3593 DVDD.n3592 0.214786
R31224 DVDD.n4785 DVDD.n3595 0.214786
R31225 DVDD.n4784 DVDD.n3596 0.214786
R31226 DVDD.n4783 DVDD.n3597 0.214786
R31227 DVDD.n4106 DVDD.n4105 0.214786
R31228 DVDD.n4107 DVDD.n4104 0.214786
R31229 DVDD.n4109 DVDD.n4108 0.214786
R31230 DVDD.n4111 DVDD.n4110 0.214786
R31231 DVDD.n4100 DVDD.n4099 0.214786
R31232 DVDD.n4115 DVDD.n4101 0.214786
R31233 DVDD.n4117 DVDD.n4116 0.214786
R31234 DVDD.n4119 DVDD.n4118 0.214786
R31235 DVDD.n4096 DVDD.n4095 0.214786
R31236 DVDD.n4123 DVDD.n4097 0.214786
R31237 DVDD.n4125 DVDD.n4124 0.214786
R31238 DVDD.n4127 DVDD.n4126 0.214786
R31239 DVDD.n4093 DVDD.n4092 0.214786
R31240 DVDD.n4132 DVDD.n4131 0.214786
R31241 DVDD.n4134 DVDD.n3826 0.214786
R31242 DVDD.n4139 DVDD.n4138 0.214786
R31243 DVDD.n3824 DVDD.n3823 0.214786
R31244 DVDD.n4145 DVDD.n4144 0.214786
R31245 DVDD.n4146 DVDD.n3822 0.214786
R31246 DVDD.n4148 DVDD.n4147 0.214786
R31247 DVDD.n4150 DVDD.n4149 0.214786
R31248 DVDD.n3819 DVDD.n3818 0.214786
R31249 DVDD.n4154 DVDD.n3820 0.214786
R31250 DVDD.n4156 DVDD.n4155 0.214786
R31251 DVDD.n4734 DVDD.n3761 0.214786
R31252 DVDD.n4733 DVDD.n3762 0.214786
R31253 DVDD.n4732 DVDD.n3763 0.214786
R31254 DVDD.n4160 DVDD.n3764 0.214786
R31255 DVDD.n4728 DVDD.n3766 0.214786
R31256 DVDD.n4727 DVDD.n3767 0.214786
R31257 DVDD.n4726 DVDD.n3768 0.214786
R31258 DVDD.n4176 DVDD.n3769 0.214786
R31259 DVDD.n4722 DVDD.n3771 0.214786
R31260 DVDD.n4721 DVDD.n4180 0.214786
R31261 DVDD.n4720 DVDD.n4181 0.214786
R31262 DVDD.n4184 DVDD.n4182 0.214786
R31263 DVDD.n4716 DVDD.n4185 0.214786
R31264 DVDD.n4715 DVDD.n4186 0.214786
R31265 DVDD.n4714 DVDD.n4187 0.214786
R31266 DVDD.n4496 DVDD.n4188 0.214786
R31267 DVDD.n4710 DVDD.n4190 0.214786
R31268 DVDD.n4709 DVDD.n4191 0.214786
R31269 DVDD.n4708 DVDD.n4192 0.214786
R31270 DVDD.n4499 DVDD.n4193 0.214786
R31271 DVDD.n4704 DVDD.n4195 0.214786
R31272 DVDD.n4703 DVDD.n4196 0.214786
R31273 DVDD.n4702 DVDD.n4197 0.214786
R31274 DVDD.n4462 DVDD.n4198 0.214786
R31275 DVDD.n4697 DVDD.n4203 0.214786
R31276 DVDD.n4696 DVDD.n4204 0.214786
R31277 DVDD.n4695 DVDD.n4205 0.214786
R31278 DVDD.n4505 DVDD.n4206 0.214786
R31279 DVDD.n4691 DVDD.n4208 0.214786
R31280 DVDD.n4690 DVDD.n4209 0.214786
R31281 DVDD.n4689 DVDD.n4210 0.214786
R31282 DVDD.n4632 DVDD.n4211 0.214786
R31283 DVDD.n4685 DVDD.n4213 0.214786
R31284 DVDD.n4684 DVDD.n4214 0.214786
R31285 DVDD.n4683 DVDD.n4215 0.214786
R31286 DVDD.n4637 DVDD.n4216 0.214786
R31287 DVDD.n4679 DVDD.n4218 0.214786
R31288 DVDD.n4678 DVDD.n4219 0.214786
R31289 DVDD.n4677 DVDD.n4220 0.214786
R31290 DVDD.n4640 DVDD.n4221 0.214786
R31291 DVDD.n4673 DVDD.n4223 0.214786
R31292 DVDD.n4672 DVDD.n4224 0.214786
R31293 DVDD.n4671 DVDD.n4225 0.214786
R31294 DVDD.n4656 DVDD.n4226 0.214786
R31295 DVDD.n4667 DVDD.n4228 0.214786
R31296 DVDD.n4666 DVDD.n4660 0.214786
R31297 DVDD.n4665 DVDD.n4661 0.214786
R31298 DVDD.n4662 DVDD.n487 0.214786
R31299 DVDD.n18135 DVDD.n486 0.214786
R31300 DVDD.n18137 DVDD.n18136 0.214786
R31301 DVDD.n18139 DVDD.n18138 0.214786
R31302 DVDD.n483 DVDD.n482 0.214786
R31303 DVDD.n18143 DVDD.n484 0.214786
R31304 DVDD.n18145 DVDD.n18144 0.214786
R31305 DVDD.n18147 DVDD.n18146 0.214786
R31306 DVDD.n479 DVDD.n478 0.214786
R31307 DVDD.n18151 DVDD.n480 0.214786
R31308 DVDD.n18153 DVDD.n18152 0.214786
R31309 DVDD.n18155 DVDD.n18154 0.214786
R31310 DVDD.n18158 DVDD.n476 0.214786
R31311 DVDD.n18160 DVDD.n18159 0.214786
R31312 DVDD.n18161 DVDD.n461 0.214786
R31313 DVDD.n4801 DVDD.n4800 0.214786
R31314 DVDD.n4799 DVDD.n3581 0.214786
R31315 DVDD.n4798 DVDD.n4797 0.214786
R31316 DVDD.n4796 DVDD.n3582 0.214786
R31317 DVDD.n4795 DVDD.n4794 0.214786
R31318 DVDD.n4793 DVDD.n3587 0.214786
R31319 DVDD.n4792 DVDD.n4791 0.214786
R31320 DVDD.n4790 DVDD.n3588 0.214786
R31321 DVDD.n4789 DVDD.n4788 0.214786
R31322 DVDD.n4787 DVDD.n3593 0.214786
R31323 DVDD.n4786 DVDD.n4785 0.214786
R31324 DVDD.n4784 DVDD.n3594 0.214786
R31325 DVDD.n4783 DVDD.n4782 0.214786
R31326 DVDD.n4105 DVDD.n3599 0.214786
R31327 DVDD.n4104 DVDD.n4103 0.214786
R31328 DVDD.n4109 DVDD.n4102 0.214786
R31329 DVDD.n4112 DVDD.n4111 0.214786
R31330 DVDD.n4113 DVDD.n4100 0.214786
R31331 DVDD.n4115 DVDD.n4114 0.214786
R31332 DVDD.n4117 DVDD.n4098 0.214786
R31333 DVDD.n4120 DVDD.n4119 0.214786
R31334 DVDD.n4121 DVDD.n4096 0.214786
R31335 DVDD.n4123 DVDD.n4122 0.214786
R31336 DVDD.n4125 DVDD.n4094 0.214786
R31337 DVDD.n4128 DVDD.n4127 0.214786
R31338 DVDD.n4129 DVDD.n4093 0.214786
R31339 DVDD.n4131 DVDD.n4130 0.214786
R31340 DVDD.n3826 DVDD.n3825 0.214786
R31341 DVDD.n4140 DVDD.n4139 0.214786
R31342 DVDD.n4141 DVDD.n3824 0.214786
R31343 DVDD.n4144 DVDD.n4143 0.214786
R31344 DVDD.n4142 DVDD.n3822 0.214786
R31345 DVDD.n4148 DVDD.n3821 0.214786
R31346 DVDD.n4151 DVDD.n4150 0.214786
R31347 DVDD.n4152 DVDD.n3819 0.214786
R31348 DVDD.n4154 DVDD.n4153 0.214786
R31349 DVDD.n4155 DVDD.n3758 0.214786
R31350 DVDD.n4735 DVDD.n4734 0.214786
R31351 DVDD.n4733 DVDD.n3759 0.214786
R31352 DVDD.n4732 DVDD.n4731 0.214786
R31353 DVDD.n4730 DVDD.n3764 0.214786
R31354 DVDD.n4729 DVDD.n4728 0.214786
R31355 DVDD.n4727 DVDD.n3765 0.214786
R31356 DVDD.n4726 DVDD.n4725 0.214786
R31357 DVDD.n4724 DVDD.n3769 0.214786
R31358 DVDD.n4723 DVDD.n4722 0.214786
R31359 DVDD.n4721 DVDD.n3770 0.214786
R31360 DVDD.n4720 DVDD.n4719 0.214786
R31361 DVDD.n4718 DVDD.n4182 0.214786
R31362 DVDD.n4717 DVDD.n4716 0.214786
R31363 DVDD.n4715 DVDD.n4183 0.214786
R31364 DVDD.n4714 DVDD.n4713 0.214786
R31365 DVDD.n4712 DVDD.n4188 0.214786
R31366 DVDD.n4711 DVDD.n4710 0.214786
R31367 DVDD.n4709 DVDD.n4189 0.214786
R31368 DVDD.n4708 DVDD.n4707 0.214786
R31369 DVDD.n4706 DVDD.n4193 0.214786
R31370 DVDD.n4705 DVDD.n4704 0.214786
R31371 DVDD.n4703 DVDD.n4194 0.214786
R31372 DVDD.n4702 DVDD.n4701 0.214786
R31373 DVDD.n4700 DVDD.n4198 0.214786
R31374 DVDD.n4698 DVDD.n4697 0.214786
R31375 DVDD.n4696 DVDD.n4201 0.214786
R31376 DVDD.n4695 DVDD.n4694 0.214786
R31377 DVDD.n4693 DVDD.n4206 0.214786
R31378 DVDD.n4692 DVDD.n4691 0.214786
R31379 DVDD.n4690 DVDD.n4207 0.214786
R31380 DVDD.n4689 DVDD.n4688 0.214786
R31381 DVDD.n4687 DVDD.n4211 0.214786
R31382 DVDD.n4686 DVDD.n4685 0.214786
R31383 DVDD.n4684 DVDD.n4212 0.214786
R31384 DVDD.n4683 DVDD.n4682 0.214786
R31385 DVDD.n4681 DVDD.n4216 0.214786
R31386 DVDD.n4680 DVDD.n4679 0.214786
R31387 DVDD.n4678 DVDD.n4217 0.214786
R31388 DVDD.n4677 DVDD.n4676 0.214786
R31389 DVDD.n4675 DVDD.n4221 0.214786
R31390 DVDD.n4674 DVDD.n4673 0.214786
R31391 DVDD.n4672 DVDD.n4222 0.214786
R31392 DVDD.n4671 DVDD.n4670 0.214786
R31393 DVDD.n4669 DVDD.n4226 0.214786
R31394 DVDD.n4668 DVDD.n4667 0.214786
R31395 DVDD.n4666 DVDD.n4227 0.214786
R31396 DVDD.n4665 DVDD.n4664 0.214786
R31397 DVDD.n4663 DVDD.n4662 0.214786
R31398 DVDD.n492 DVDD.n486 0.214786
R31399 DVDD.n18137 DVDD.n485 0.214786
R31400 DVDD.n18140 DVDD.n18139 0.214786
R31401 DVDD.n18141 DVDD.n483 0.214786
R31402 DVDD.n18143 DVDD.n18142 0.214786
R31403 DVDD.n18145 DVDD.n481 0.214786
R31404 DVDD.n18148 DVDD.n18147 0.214786
R31405 DVDD.n18149 DVDD.n479 0.214786
R31406 DVDD.n18151 DVDD.n18150 0.214786
R31407 DVDD.n18153 DVDD.n477 0.214786
R31408 DVDD.n18156 DVDD.n18155 0.214786
R31409 DVDD.n18158 DVDD.n18157 0.214786
R31410 DVDD.n18160 DVDD.n475 0.214786
R31411 DVDD.n2898 DVDD.n2895 0.214786
R31412 DVDD.n2900 DVDD.n2894 0.214786
R31413 DVDD.n2902 DVDD.n2893 0.214786
R31414 DVDD.n2904 DVDD.n2892 0.214786
R31415 DVDD.n2906 DVDD.n2891 0.214786
R31416 DVDD.n2908 DVDD.n2890 0.214786
R31417 DVDD.n2910 DVDD.n2889 0.214786
R31418 DVDD.n2912 DVDD.n2888 0.214786
R31419 DVDD.n2914 DVDD.n2887 0.214786
R31420 DVDD.n2916 DVDD.n2886 0.214786
R31421 DVDD.n15328 DVDD.n15323 0.214786
R31422 DVDD.n15331 DVDD.n15330 0.214786
R31423 DVDD.n15332 DVDD.n15322 0.214786
R31424 DVDD.n15335 DVDD.n15333 0.214786
R31425 DVDD.n15337 DVDD.n15320 0.214786
R31426 DVDD.n15340 DVDD.n15339 0.214786
R31427 DVDD.n15341 DVDD.n15319 0.214786
R31428 DVDD.n15404 DVDD.n15342 0.214786
R31429 DVDD.n15403 DVDD.n15343 0.214786
R31430 DVDD.n15401 DVDD.n15344 0.214786
R31431 DVDD.n15399 DVDD.n15345 0.214786
R31432 DVDD.n15398 DVDD.n15346 0.214786
R31433 DVDD.n15397 DVDD.n15347 0.214786
R31434 DVDD.n15393 DVDD.n15350 0.214786
R31435 DVDD.n15392 DVDD.n15351 0.214786
R31436 DVDD.n15391 DVDD.n15352 0.214786
R31437 DVDD.n15389 DVDD.n15353 0.214786
R31438 DVDD.n15387 DVDD.n15354 0.214786
R31439 DVDD.n15385 DVDD.n15355 0.214786
R31440 DVDD.n15383 DVDD.n15356 0.214786
R31441 DVDD.n15381 DVDD.n15357 0.214786
R31442 DVDD.n15379 DVDD.n15358 0.214786
R31443 DVDD.n15377 DVDD.n15359 0.214786
R31444 DVDD.n15375 DVDD.n15360 0.214786
R31445 DVDD.n15373 DVDD.n15361 0.214786
R31446 DVDD.n15371 DVDD.n15362 0.214786
R31447 DVDD.n15369 DVDD.n15363 0.214786
R31448 DVDD.n15367 DVDD.n15365 0.214786
R31449 DVDD.n15364 DVDD.n3138 0.214786
R31450 DVDD.n16005 DVDD.n3139 0.214786
R31451 DVDD.n16004 DVDD.n3140 0.214786
R31452 DVDD.n16003 DVDD.n3141 0.214786
R31453 DVDD.n16000 DVDD.n3142 0.214786
R31454 DVDD.n15999 DVDD.n3143 0.214786
R31455 DVDD.n15997 DVDD.n3144 0.214786
R31456 DVDD.n15995 DVDD.n3145 0.214786
R31457 DVDD.n15993 DVDD.n3146 0.214786
R31458 DVDD.n3225 DVDD.n3224 0.214786
R31459 DVDD.n3222 DVDD.n3209 0.214786
R31460 DVDD.n3220 DVDD.n3210 0.214786
R31461 DVDD.n3218 DVDD.n3211 0.214786
R31462 DVDD.n3216 DVDD.n3212 0.214786
R31463 DVDD.n3214 DVDD.n3213 0.214786
R31464 DVDD.n3056 DVDD.n3055 0.214786
R31465 DVDD.n16088 DVDD.n16087 0.214786
R31466 DVDD.n16089 DVDD.n3054 0.214786
R31467 DVDD.n16091 DVDD.n16090 0.214786
R31468 DVDD.n3052 DVDD.n3051 0.214786
R31469 DVDD.n16096 DVDD.n16095 0.214786
R31470 DVDD.n16097 DVDD.n3050 0.214786
R31471 DVDD.n16100 DVDD.n16099 0.214786
R31472 DVDD.n16098 DVDD.n3047 0.214786
R31473 DVDD.n16115 DVDD.n3048 0.214786
R31474 DVDD.n16117 DVDD.n3046 0.214786
R31475 DVDD.n16120 DVDD.n16119 0.214786
R31476 DVDD.n16121 DVDD.n3045 0.214786
R31477 DVDD.n16124 DVDD.n16122 0.214786
R31478 DVDD.n16126 DVDD.n3043 0.214786
R31479 DVDD.n16129 DVDD.n16128 0.214786
R31480 DVDD.n16130 DVDD.n3042 0.214786
R31481 DVDD.n16133 DVDD.n16131 0.214786
R31482 DVDD.n16137 DVDD.n16136 0.214786
R31483 DVDD.n16139 DVDD.n16138 0.214786
R31484 DVDD.n2994 DVDD.n2993 0.214786
R31485 DVDD.n16147 DVDD.n16146 0.214786
R31486 DVDD.n16148 DVDD.n2992 0.214786
R31487 DVDD.n16151 DVDD.n16150 0.214786
R31488 DVDD.n16149 DVDD.n2990 0.214786
R31489 DVDD.n16155 DVDD.n2989 0.214786
R31490 DVDD.n16158 DVDD.n16157 0.214786
R31491 DVDD.n16159 DVDD.n2988 0.214786
R31492 DVDD.n16162 DVDD.n16160 0.214786
R31493 DVDD.n16164 DVDD.n2986 0.214786
R31494 DVDD.n16167 DVDD.n16166 0.214786
R31495 DVDD.n16168 DVDD.n2985 0.214786
R31496 DVDD.n16171 DVDD.n16169 0.214786
R31497 DVDD.n16173 DVDD.n2983 0.214786
R31498 DVDD.n16176 DVDD.n16175 0.214786
R31499 DVDD.n16177 DVDD.n2982 0.214786
R31500 DVDD.n16179 DVDD.n16178 0.214786
R31501 DVDD.n2923 DVDD.n2922 0.214786
R31502 DVDD.n16187 DVDD.n16186 0.214786
R31503 DVDD.n16188 DVDD.n2921 0.214786
R31504 DVDD.n16192 DVDD.n16191 0.214786
R31505 DVDD.n16190 DVDD.n2882 0.214786
R31506 DVDD.n16198 DVDD.n2883 0.214786
R31507 DVDD.n2919 DVDD.n2884 0.214786
R31508 DVDD.n2918 DVDD.n2885 0.214786
R31509 DVDD.n15456 DVDD.n15425 0.214786
R31510 DVDD.n15454 DVDD.n15426 0.214786
R31511 DVDD.n15452 DVDD.n15427 0.214786
R31512 DVDD.n15450 DVDD.n15428 0.214786
R31513 DVDD.n15448 DVDD.n15429 0.214786
R31514 DVDD.n15446 DVDD.n15430 0.214786
R31515 DVDD.n15444 DVDD.n15431 0.214786
R31516 DVDD.n15442 DVDD.n15432 0.214786
R31517 DVDD.n15440 DVDD.n15433 0.214786
R31518 DVDD.n15438 DVDD.n15434 0.214786
R31519 DVDD.n15436 DVDD.n15435 0.214786
R31520 DVDD.n5228 DVDD.n5227 0.214786
R31521 DVDD.n15465 DVDD.n15464 0.214786
R31522 DVDD.n15469 DVDD.n15468 0.214786
R31523 DVDD.n15467 DVDD.n5223 0.214786
R31524 DVDD.n15473 DVDD.n5224 0.214786
R31525 DVDD.n15475 DVDD.n5222 0.214786
R31526 DVDD.n15478 DVDD.n15477 0.214786
R31527 DVDD.n15479 DVDD.n5221 0.214786
R31528 DVDD.n15482 DVDD.n15480 0.214786
R31529 DVDD.n15484 DVDD.n5219 0.214786
R31530 DVDD.n15487 DVDD.n15486 0.214786
R31531 DVDD.n15488 DVDD.n5218 0.214786
R31532 DVDD.n15491 DVDD.n15489 0.214786
R31533 DVDD.n15493 DVDD.n5216 0.214786
R31534 DVDD.n15496 DVDD.n15495 0.214786
R31535 DVDD.n15497 DVDD.n5215 0.214786
R31536 DVDD.n15518 DVDD.n15498 0.214786
R31537 DVDD.n15517 DVDD.n15499 0.214786
R31538 DVDD.n15516 DVDD.n15500 0.214786
R31539 DVDD.n15515 DVDD.n15501 0.214786
R31540 DVDD.n15503 DVDD.n15502 0.214786
R31541 DVDD.n15511 DVDD.n15504 0.214786
R31542 DVDD.n15510 DVDD.n15505 0.214786
R31543 DVDD.n15508 DVDD.n15506 0.214786
R31544 DVDD.n3230 DVDD.n3228 0.214786
R31545 DVDD.n15915 DVDD.n15914 0.214786
R31546 DVDD.n15917 DVDD.n3208 0.214786
R31547 DVDD.n15920 DVDD.n15918 0.214786
R31548 DVDD.n15922 DVDD.n3207 0.214786
R31549 DVDD.n15925 DVDD.n15924 0.214786
R31550 DVDD.n15926 DVDD.n3206 0.214786
R31551 DVDD.n15929 DVDD.n15927 0.214786
R31552 DVDD.n15939 DVDD.n3204 0.214786
R31553 DVDD.n15942 DVDD.n15941 0.214786
R31554 DVDD.n15943 DVDD.n3203 0.214786
R31555 DVDD.n15985 DVDD.n15944 0.214786
R31556 DVDD.n15984 DVDD.n15945 0.214786
R31557 DVDD.n15983 DVDD.n15946 0.214786
R31558 DVDD.n15949 DVDD.n15947 0.214786
R31559 DVDD.n15979 DVDD.n15950 0.214786
R31560 DVDD.n15978 DVDD.n15951 0.214786
R31561 DVDD.n15977 DVDD.n15952 0.214786
R31562 DVDD.n15975 DVDD.n15953 0.214786
R31563 DVDD.n15973 DVDD.n15954 0.214786
R31564 DVDD.n15971 DVDD.n15955 0.214786
R31565 DVDD.n15969 DVDD.n15956 0.214786
R31566 DVDD.n15967 DVDD.n15957 0.214786
R31567 DVDD.n15965 DVDD.n15958 0.214786
R31568 DVDD.n15963 DVDD.n15959 0.214786
R31569 DVDD.n15961 DVDD.n2706 0.214786
R31570 DVDD.n16260 DVDD.n16259 0.214786
R31571 DVDD.n2709 DVDD.n2707 0.214786
R31572 DVDD.n2774 DVDD.n2773 0.214786
R31573 DVDD.n2775 DVDD.n2771 0.214786
R31574 DVDD.n16253 DVDD.n2776 0.214786
R31575 DVDD.n16252 DVDD.n2777 0.214786
R31576 DVDD.n16251 DVDD.n2778 0.214786
R31577 DVDD.n2843 DVDD.n2779 0.214786
R31578 DVDD.n2844 DVDD.n2842 0.214786
R31579 DVDD.n2847 DVDD.n2845 0.214786
R31580 DVDD.n2849 DVDD.n2841 0.214786
R31581 DVDD.n2852 DVDD.n2851 0.214786
R31582 DVDD.n2853 DVDD.n2840 0.214786
R31583 DVDD.n2856 DVDD.n2854 0.214786
R31584 DVDD.n2858 DVDD.n2838 0.214786
R31585 DVDD.n2861 DVDD.n2860 0.214786
R31586 DVDD.n2862 DVDD.n2837 0.214786
R31587 DVDD.n2864 DVDD.n2863 0.214786
R31588 DVDD.n2874 DVDD.n2835 0.214786
R31589 DVDD.n2877 DVDD.n2876 0.214786
R31590 DVDD.n2878 DVDD.n2834 0.214786
R31591 DVDD.n16244 DVDD.n2879 0.214786
R31592 DVDD.n16243 DVDD.n2880 0.214786
R31593 DVDD.n16242 DVDD.n2881 0.214786
R31594 DVDD.n16239 DVDD.n16200 0.214786
R31595 DVDD.n16237 DVDD.n16201 0.214786
R31596 DVDD.n16236 DVDD.n16202 0.214786
R31597 DVDD.n16235 DVDD.n16203 0.214786
R31598 DVDD.n16233 DVDD.n16204 0.214786
R31599 DVDD.n16231 DVDD.n16205 0.214786
R31600 DVDD.n16229 DVDD.n16206 0.214786
R31601 DVDD.n16227 DVDD.n16207 0.214786
R31602 DVDD.n16225 DVDD.n16208 0.214786
R31603 DVDD.n16223 DVDD.n16209 0.214786
R31604 DVDD.n16221 DVDD.n16210 0.214786
R31605 DVDD.n16219 DVDD.n16211 0.214786
R31606 DVDD.n16217 DVDD.n16212 0.214786
R31607 DVDD.n5090 DVDD.n5087 0.214786
R31608 DVDD.n5093 DVDD.n5092 0.214786
R31609 DVDD.n5094 DVDD.n5086 0.214786
R31610 DVDD.n5097 DVDD.n5095 0.214786
R31611 DVDD.n5099 DVDD.n5084 0.214786
R31612 DVDD.n5102 DVDD.n5101 0.214786
R31613 DVDD.n5103 DVDD.n5083 0.214786
R31614 DVDD.n15696 DVDD.n5104 0.214786
R31615 DVDD.n15695 DVDD.n5105 0.214786
R31616 DVDD.n15693 DVDD.n5106 0.214786
R31617 DVDD.n15691 DVDD.n5107 0.214786
R31618 DVDD.n15689 DVDD.n5108 0.214786
R31619 DVDD.n5110 DVDD.n5109 0.214786
R31620 DVDD.n15684 DVDD.n5114 0.214786
R31621 DVDD.n15683 DVDD.n5115 0.214786
R31622 DVDD.n15682 DVDD.n5116 0.214786
R31623 DVDD.n15629 DVDD.n5117 0.214786
R31624 DVDD.n15632 DVDD.n15630 0.214786
R31625 DVDD.n15634 DVDD.n15628 0.214786
R31626 DVDD.n15637 DVDD.n15636 0.214786
R31627 DVDD.n15638 DVDD.n15627 0.214786
R31628 DVDD.n15641 DVDD.n15639 0.214786
R31629 DVDD.n15643 DVDD.n15625 0.214786
R31630 DVDD.n15646 DVDD.n15645 0.214786
R31631 DVDD.n15647 DVDD.n15624 0.214786
R31632 DVDD.n15650 DVDD.n15648 0.214786
R31633 DVDD.n15652 DVDD.n15622 0.214786
R31634 DVDD.n15655 DVDD.n15654 0.214786
R31635 DVDD.n15656 DVDD.n15621 0.214786
R31636 DVDD.n15676 DVDD.n15657 0.214786
R31637 DVDD.n15675 DVDD.n15658 0.214786
R31638 DVDD.n15674 DVDD.n15659 0.214786
R31639 DVDD.n15671 DVDD.n15660 0.214786
R31640 DVDD.n15670 DVDD.n15661 0.214786
R31641 DVDD.n15668 DVDD.n15662 0.214786
R31642 DVDD.n15666 DVDD.n15664 0.214786
R31643 DVDD.n15663 DVDD.n3232 0.214786
R31644 DVDD.n15911 DVDD.n3233 0.214786
R31645 DVDD.n3301 DVDD.n3234 0.214786
R31646 DVDD.n3304 DVDD.n3302 0.214786
R31647 DVDD.n3307 DVDD.n3306 0.214786
R31648 DVDD.n3308 DVDD.n3300 0.214786
R31649 DVDD.n3311 DVDD.n3309 0.214786
R31650 DVDD.n3313 DVDD.n3298 0.214786
R31651 DVDD.n3316 DVDD.n3315 0.214786
R31652 DVDD.n3317 DVDD.n3297 0.214786
R31653 DVDD.n15905 DVDD.n3318 0.214786
R31654 DVDD.n15904 DVDD.n3319 0.214786
R31655 DVDD.n15903 DVDD.n3320 0.214786
R31656 DVDD.n3323 DVDD.n3321 0.214786
R31657 DVDD.n15899 DVDD.n3324 0.214786
R31658 DVDD.n15898 DVDD.n3325 0.214786
R31659 DVDD.n15897 DVDD.n3326 0.214786
R31660 DVDD.n15895 DVDD.n3327 0.214786
R31661 DVDD.n15893 DVDD.n3328 0.214786
R31662 DVDD.n15891 DVDD.n3329 0.214786
R31663 DVDD.n15889 DVDD.n3330 0.214786
R31664 DVDD.n15887 DVDD.n3331 0.214786
R31665 DVDD.n15885 DVDD.n3332 0.214786
R31666 DVDD.n15883 DVDD.n3333 0.214786
R31667 DVDD.n15881 DVDD.n2704 0.214786
R31668 DVDD.n16263 DVDD.n2702 0.214786
R31669 DVDD.n16265 DVDD.n16264 0.214786
R31670 DVDD.n2643 DVDD.n2642 0.214786
R31671 DVDD.n16273 DVDD.n16272 0.214786
R31672 DVDD.n16274 DVDD.n2641 0.214786
R31673 DVDD.n16277 DVDD.n16276 0.214786
R31674 DVDD.n16275 DVDD.n2638 0.214786
R31675 DVDD.n16281 DVDD.n2639 0.214786
R31676 DVDD.n16283 DVDD.n2637 0.214786
R31677 DVDD.n16286 DVDD.n16285 0.214786
R31678 DVDD.n16287 DVDD.n2636 0.214786
R31679 DVDD.n16290 DVDD.n16288 0.214786
R31680 DVDD.n16292 DVDD.n2634 0.214786
R31681 DVDD.n16295 DVDD.n16294 0.214786
R31682 DVDD.n16296 DVDD.n2633 0.214786
R31683 DVDD.n16299 DVDD.n16297 0.214786
R31684 DVDD.n16301 DVDD.n2631 0.214786
R31685 DVDD.n16304 DVDD.n16303 0.214786
R31686 DVDD.n16305 DVDD.n2630 0.214786
R31687 DVDD.n16310 DVDD.n16306 0.214786
R31688 DVDD.n16309 DVDD.n16308 0.214786
R31689 DVDD.n16307 DVDD.n2570 0.214786
R31690 DVDD.n16317 DVDD.n2569 0.214786
R31691 DVDD.n16319 DVDD.n16318 0.214786
R31692 DVDD.n16359 DVDD.n16321 0.214786
R31693 DVDD.n16358 DVDD.n16322 0.214786
R31694 DVDD.n16357 DVDD.n16323 0.214786
R31695 DVDD.n16356 DVDD.n16324 0.214786
R31696 DVDD.n16354 DVDD.n16325 0.214786
R31697 DVDD.n16352 DVDD.n16326 0.214786
R31698 DVDD.n16350 DVDD.n16327 0.214786
R31699 DVDD.n16348 DVDD.n16328 0.214786
R31700 DVDD.n16346 DVDD.n16329 0.214786
R31701 DVDD.n16344 DVDD.n16330 0.214786
R31702 DVDD.n16342 DVDD.n16331 0.214786
R31703 DVDD.n16340 DVDD.n16332 0.214786
R31704 DVDD.n16338 DVDD.n16333 0.214786
R31705 DVDD.n15747 DVDD.n15716 0.214786
R31706 DVDD.n15745 DVDD.n15717 0.214786
R31707 DVDD.n15743 DVDD.n15718 0.214786
R31708 DVDD.n15741 DVDD.n15719 0.214786
R31709 DVDD.n15739 DVDD.n15720 0.214786
R31710 DVDD.n15737 DVDD.n15721 0.214786
R31711 DVDD.n15735 DVDD.n15722 0.214786
R31712 DVDD.n15733 DVDD.n15723 0.214786
R31713 DVDD.n15731 DVDD.n15724 0.214786
R31714 DVDD.n15729 DVDD.n15725 0.214786
R31715 DVDD.n15727 DVDD.n15726 0.214786
R31716 DVDD.n3509 DVDD.n3508 0.214786
R31717 DVDD.n15756 DVDD.n15755 0.214786
R31718 DVDD.n15760 DVDD.n15759 0.214786
R31719 DVDD.n15758 DVDD.n3504 0.214786
R31720 DVDD.n15764 DVDD.n3503 0.214786
R31721 DVDD.n15767 DVDD.n15766 0.214786
R31722 DVDD.n15768 DVDD.n3502 0.214786
R31723 DVDD.n15771 DVDD.n15769 0.214786
R31724 DVDD.n15773 DVDD.n3500 0.214786
R31725 DVDD.n15776 DVDD.n15775 0.214786
R31726 DVDD.n15777 DVDD.n3499 0.214786
R31727 DVDD.n15780 DVDD.n15778 0.214786
R31728 DVDD.n15782 DVDD.n3497 0.214786
R31729 DVDD.n15785 DVDD.n15784 0.214786
R31730 DVDD.n15786 DVDD.n3496 0.214786
R31731 DVDD.n15788 DVDD.n15787 0.214786
R31732 DVDD.n3418 DVDD.n3417 0.214786
R31733 DVDD.n15798 DVDD.n15797 0.214786
R31734 DVDD.n15799 DVDD.n3416 0.214786
R31735 DVDD.n15801 DVDD.n15800 0.214786
R31736 DVDD.n3414 DVDD.n3413 0.214786
R31737 DVDD.n15806 DVDD.n15805 0.214786
R31738 DVDD.n15807 DVDD.n3412 0.214786
R31739 DVDD.n15810 DVDD.n15808 0.214786
R31740 DVDD.n15812 DVDD.n3410 0.214786
R31741 DVDD.n15816 DVDD.n15815 0.214786
R31742 DVDD.n15820 DVDD.n15818 0.214786
R31743 DVDD.n15823 DVDD.n15822 0.214786
R31744 DVDD.n15824 DVDD.n3409 0.214786
R31745 DVDD.n15827 DVDD.n15825 0.214786
R31746 DVDD.n15829 DVDD.n3407 0.214786
R31747 DVDD.n15832 DVDD.n15831 0.214786
R31748 DVDD.n15833 DVDD.n3406 0.214786
R31749 DVDD.n15835 DVDD.n15834 0.214786
R31750 DVDD.n3346 DVDD.n3345 0.214786
R31751 DVDD.n15842 DVDD.n15841 0.214786
R31752 DVDD.n15843 DVDD.n3344 0.214786
R31753 DVDD.n15845 DVDD.n15844 0.214786
R31754 DVDD.n3342 DVDD.n3341 0.214786
R31755 DVDD.n15851 DVDD.n15850 0.214786
R31756 DVDD.n15852 DVDD.n3340 0.214786
R31757 DVDD.n15855 DVDD.n15853 0.214786
R31758 DVDD.n15857 DVDD.n3339 0.214786
R31759 DVDD.n15860 DVDD.n15859 0.214786
R31760 DVDD.n15861 DVDD.n3338 0.214786
R31761 DVDD.n15864 DVDD.n15862 0.214786
R31762 DVDD.n15866 DVDD.n3336 0.214786
R31763 DVDD.n15869 DVDD.n15868 0.214786
R31764 DVDD.n15870 DVDD.n3335 0.214786
R31765 DVDD.n15873 DVDD.n15871 0.214786
R31766 DVDD.n15877 DVDD.n15875 0.214786
R31767 DVDD.n15874 DVDD.n2379 0.214786
R31768 DVDD.n16380 DVDD.n2380 0.214786
R31769 DVDD.n16379 DVDD.n2381 0.214786
R31770 DVDD.n16378 DVDD.n2382 0.214786
R31771 DVDD.n16377 DVDD.n2383 0.214786
R31772 DVDD.n2386 DVDD.n2384 0.214786
R31773 DVDD.n16373 DVDD.n2387 0.214786
R31774 DVDD.n16372 DVDD.n2388 0.214786
R31775 DVDD.n2494 DVDD.n2389 0.214786
R31776 DVDD.n2497 DVDD.n2495 0.214786
R31777 DVDD.n2500 DVDD.n2499 0.214786
R31778 DVDD.n2501 DVDD.n2493 0.214786
R31779 DVDD.n2504 DVDD.n2502 0.214786
R31780 DVDD.n2506 DVDD.n2491 0.214786
R31781 DVDD.n2509 DVDD.n2508 0.214786
R31782 DVDD.n2510 DVDD.n2490 0.214786
R31783 DVDD.n2513 DVDD.n2511 0.214786
R31784 DVDD.n2515 DVDD.n2488 0.214786
R31785 DVDD.n2518 DVDD.n2517 0.214786
R31786 DVDD.n2519 DVDD.n2487 0.214786
R31787 DVDD.n16366 DVDD.n2520 0.214786
R31788 DVDD.n16365 DVDD.n2521 0.214786
R31789 DVDD.n16364 DVDD.n2522 0.214786
R31790 DVDD.n2566 DVDD.n2565 0.214786
R31791 DVDD.n2564 DVDD.n2528 0.214786
R31792 DVDD.n2562 DVDD.n2529 0.214786
R31793 DVDD.n2560 DVDD.n2530 0.214786
R31794 DVDD.n2558 DVDD.n2531 0.214786
R31795 DVDD.n2556 DVDD.n2532 0.214786
R31796 DVDD.n2554 DVDD.n2533 0.214786
R31797 DVDD.n2552 DVDD.n2534 0.214786
R31798 DVDD.n2550 DVDD.n2535 0.214786
R31799 DVDD.n2548 DVDD.n2536 0.214786
R31800 DVDD.n2546 DVDD.n2537 0.214786
R31801 DVDD.n2544 DVDD.n2538 0.214786
R31802 DVDD.n2542 DVDD.n2539 0.214786
R31803 DVDD.n2540 DVDD.n517 0.214786
R31804 DVDD.n2542 DVDD.n2541 0.214786
R31805 DVDD.n2544 DVDD.n2543 0.214786
R31806 DVDD.n2546 DVDD.n2545 0.214786
R31807 DVDD.n2548 DVDD.n2547 0.214786
R31808 DVDD.n2550 DVDD.n2549 0.214786
R31809 DVDD.n2552 DVDD.n2551 0.214786
R31810 DVDD.n2554 DVDD.n2553 0.214786
R31811 DVDD.n2556 DVDD.n2555 0.214786
R31812 DVDD.n2558 DVDD.n2557 0.214786
R31813 DVDD.n2560 DVDD.n2559 0.214786
R31814 DVDD.n2562 DVDD.n2561 0.214786
R31815 DVDD.n2564 DVDD.n2563 0.214786
R31816 DVDD.n2565 DVDD.n2524 0.214786
R31817 DVDD.n16364 DVDD.n16363 0.214786
R31818 DVDD.n16365 DVDD.n2486 0.214786
R31819 DVDD.n16367 DVDD.n16366 0.214786
R31820 DVDD.n2487 DVDD.n2483 0.214786
R31821 DVDD.n2517 DVDD.n2516 0.214786
R31822 DVDD.n2515 DVDD.n2514 0.214786
R31823 DVDD.n2513 DVDD.n2512 0.214786
R31824 DVDD.n2490 DVDD.n2489 0.214786
R31825 DVDD.n2508 DVDD.n2507 0.214786
R31826 DVDD.n2506 DVDD.n2505 0.214786
R31827 DVDD.n2504 DVDD.n2503 0.214786
R31828 DVDD.n2493 DVDD.n2492 0.214786
R31829 DVDD.n2499 DVDD.n2498 0.214786
R31830 DVDD.n2497 DVDD.n2496 0.214786
R31831 DVDD.n2476 DVDD.n2389 0.214786
R31832 DVDD.n16372 DVDD.n16371 0.214786
R31833 DVDD.n16374 DVDD.n16373 0.214786
R31834 DVDD.n16375 DVDD.n2384 0.214786
R31835 DVDD.n16377 DVDD.n16376 0.214786
R31836 DVDD.n16378 DVDD.n2362 0.214786
R31837 DVDD.n16379 DVDD.n2349 0.214786
R31838 DVDD.n16381 DVDD.n16380 0.214786
R31839 DVDD.n2379 DVDD.n2378 0.214786
R31840 DVDD.n15877 DVDD.n15876 0.214786
R31841 DVDD.n15873 DVDD.n15872 0.214786
R31842 DVDD.n3335 DVDD.n3334 0.214786
R31843 DVDD.n15868 DVDD.n15867 0.214786
R31844 DVDD.n15866 DVDD.n15865 0.214786
R31845 DVDD.n15864 DVDD.n15863 0.214786
R31846 DVDD.n3338 DVDD.n3337 0.214786
R31847 DVDD.n15859 DVDD.n15858 0.214786
R31848 DVDD.n15857 DVDD.n15856 0.214786
R31849 DVDD.n15855 DVDD.n15854 0.214786
R31850 DVDD.n15848 DVDD.n3340 0.214786
R31851 DVDD.n15850 DVDD.n15849 0.214786
R31852 DVDD.n15847 DVDD.n3342 0.214786
R31853 DVDD.n15846 DVDD.n15845 0.214786
R31854 DVDD.n3344 DVDD.n3343 0.214786
R31855 DVDD.n15841 DVDD.n15840 0.214786
R31856 DVDD.n3347 DVDD.n3346 0.214786
R31857 DVDD.n15836 DVDD.n15835 0.214786
R31858 DVDD.n3406 DVDD.n3405 0.214786
R31859 DVDD.n15831 DVDD.n15830 0.214786
R31860 DVDD.n15829 DVDD.n15828 0.214786
R31861 DVDD.n15827 DVDD.n15826 0.214786
R31862 DVDD.n3409 DVDD.n3408 0.214786
R31863 DVDD.n15822 DVDD.n15821 0.214786
R31864 DVDD.n15820 DVDD.n15819 0.214786
R31865 DVDD.n15815 DVDD.n15814 0.214786
R31866 DVDD.n15812 DVDD.n15811 0.214786
R31867 DVDD.n15810 DVDD.n15809 0.214786
R31868 DVDD.n3412 DVDD.n3411 0.214786
R31869 DVDD.n15805 DVDD.n15804 0.214786
R31870 DVDD.n15803 DVDD.n3414 0.214786
R31871 DVDD.n15802 DVDD.n15801 0.214786
R31872 DVDD.n3416 DVDD.n3415 0.214786
R31873 DVDD.n15797 DVDD.n15796 0.214786
R31874 DVDD.n15791 DVDD.n3418 0.214786
R31875 DVDD.n15789 DVDD.n15788 0.214786
R31876 DVDD.n3496 DVDD.n3495 0.214786
R31877 DVDD.n15784 DVDD.n15783 0.214786
R31878 DVDD.n15782 DVDD.n15781 0.214786
R31879 DVDD.n15780 DVDD.n15779 0.214786
R31880 DVDD.n3499 DVDD.n3498 0.214786
R31881 DVDD.n15775 DVDD.n15774 0.214786
R31882 DVDD.n15773 DVDD.n15772 0.214786
R31883 DVDD.n15771 DVDD.n15770 0.214786
R31884 DVDD.n3502 DVDD.n3501 0.214786
R31885 DVDD.n15766 DVDD.n15765 0.214786
R31886 DVDD.n15764 DVDD.n15763 0.214786
R31887 DVDD.n15762 DVDD.n3504 0.214786
R31888 DVDD.n15761 DVDD.n15760 0.214786
R31889 DVDD.n15755 DVDD.n15754 0.214786
R31890 DVDD.n15753 DVDD.n3509 0.214786
R31891 DVDD.n15727 DVDD.n3510 0.214786
R31892 DVDD.n15729 DVDD.n15728 0.214786
R31893 DVDD.n15731 DVDD.n15730 0.214786
R31894 DVDD.n15733 DVDD.n15732 0.214786
R31895 DVDD.n15735 DVDD.n15734 0.214786
R31896 DVDD.n15737 DVDD.n15736 0.214786
R31897 DVDD.n15739 DVDD.n15738 0.214786
R31898 DVDD.n15741 DVDD.n15740 0.214786
R31899 DVDD.n15743 DVDD.n15742 0.214786
R31900 DVDD.n15745 DVDD.n15744 0.214786
R31901 DVDD.n15747 DVDD.n15746 0.214786
R31902 DVDD.n15749 DVDD.n15748 0.214786
R31903 DVDD.n16336 DVDD.n16335 0.214786
R31904 DVDD.n16338 DVDD.n16337 0.214786
R31905 DVDD.n16340 DVDD.n16339 0.214786
R31906 DVDD.n16342 DVDD.n16341 0.214786
R31907 DVDD.n16344 DVDD.n16343 0.214786
R31908 DVDD.n16346 DVDD.n16345 0.214786
R31909 DVDD.n16348 DVDD.n16347 0.214786
R31910 DVDD.n16350 DVDD.n16349 0.214786
R31911 DVDD.n16352 DVDD.n16351 0.214786
R31912 DVDD.n16354 DVDD.n16353 0.214786
R31913 DVDD.n16356 DVDD.n16355 0.214786
R31914 DVDD.n16357 DVDD.n583 0.214786
R31915 DVDD.n16358 DVDD.n569 0.214786
R31916 DVDD.n16360 DVDD.n16359 0.214786
R31917 DVDD.n16318 DVDD.n2526 0.214786
R31918 DVDD.n16317 DVDD.n16316 0.214786
R31919 DVDD.n16315 DVDD.n2570 0.214786
R31920 DVDD.n16309 DVDD.n2571 0.214786
R31921 DVDD.n16311 DVDD.n16310 0.214786
R31922 DVDD.n2630 DVDD.n2629 0.214786
R31923 DVDD.n16303 DVDD.n16302 0.214786
R31924 DVDD.n16301 DVDD.n16300 0.214786
R31925 DVDD.n16299 DVDD.n16298 0.214786
R31926 DVDD.n2633 DVDD.n2632 0.214786
R31927 DVDD.n16294 DVDD.n16293 0.214786
R31928 DVDD.n16292 DVDD.n16291 0.214786
R31929 DVDD.n16290 DVDD.n16289 0.214786
R31930 DVDD.n2636 DVDD.n2635 0.214786
R31931 DVDD.n16285 DVDD.n16284 0.214786
R31932 DVDD.n16283 DVDD.n16282 0.214786
R31933 DVDD.n16281 DVDD.n16280 0.214786
R31934 DVDD.n16279 DVDD.n2638 0.214786
R31935 DVDD.n16278 DVDD.n16277 0.214786
R31936 DVDD.n2641 DVDD.n2640 0.214786
R31937 DVDD.n16272 DVDD.n16271 0.214786
R31938 DVDD.n16267 DVDD.n2643 0.214786
R31939 DVDD.n16266 DVDD.n16265 0.214786
R31940 DVDD.n2702 DVDD.n2701 0.214786
R31941 DVDD.n15881 DVDD.n15880 0.214786
R31942 DVDD.n15883 DVDD.n15882 0.214786
R31943 DVDD.n15885 DVDD.n15884 0.214786
R31944 DVDD.n15887 DVDD.n15886 0.214786
R31945 DVDD.n15889 DVDD.n15888 0.214786
R31946 DVDD.n15891 DVDD.n15890 0.214786
R31947 DVDD.n15893 DVDD.n15892 0.214786
R31948 DVDD.n15895 DVDD.n15894 0.214786
R31949 DVDD.n15897 DVDD.n15896 0.214786
R31950 DVDD.n15898 DVDD.n3322 0.214786
R31951 DVDD.n15900 DVDD.n15899 0.214786
R31952 DVDD.n15901 DVDD.n3321 0.214786
R31953 DVDD.n15903 DVDD.n15902 0.214786
R31954 DVDD.n15904 DVDD.n3296 0.214786
R31955 DVDD.n15906 DVDD.n15905 0.214786
R31956 DVDD.n3297 DVDD.n3295 0.214786
R31957 DVDD.n3315 DVDD.n3314 0.214786
R31958 DVDD.n3313 DVDD.n3312 0.214786
R31959 DVDD.n3311 DVDD.n3310 0.214786
R31960 DVDD.n3300 DVDD.n3299 0.214786
R31961 DVDD.n3306 DVDD.n3305 0.214786
R31962 DVDD.n3304 DVDD.n3303 0.214786
R31963 DVDD.n3248 DVDD.n3234 0.214786
R31964 DVDD.n15911 DVDD.n15910 0.214786
R31965 DVDD.n3282 DVDD.n3232 0.214786
R31966 DVDD.n15666 DVDD.n15665 0.214786
R31967 DVDD.n15668 DVDD.n15667 0.214786
R31968 DVDD.n15670 DVDD.n15669 0.214786
R31969 DVDD.n15672 DVDD.n15671 0.214786
R31970 DVDD.n15674 DVDD.n15673 0.214786
R31971 DVDD.n15675 DVDD.n15620 0.214786
R31972 DVDD.n15677 DVDD.n15676 0.214786
R31973 DVDD.n15621 DVDD.n15619 0.214786
R31974 DVDD.n15654 DVDD.n15653 0.214786
R31975 DVDD.n15652 DVDD.n15651 0.214786
R31976 DVDD.n15650 DVDD.n15649 0.214786
R31977 DVDD.n15624 DVDD.n15623 0.214786
R31978 DVDD.n15645 DVDD.n15644 0.214786
R31979 DVDD.n15643 DVDD.n15642 0.214786
R31980 DVDD.n15641 DVDD.n15640 0.214786
R31981 DVDD.n15627 DVDD.n15626 0.214786
R31982 DVDD.n15636 DVDD.n15635 0.214786
R31983 DVDD.n15634 DVDD.n15633 0.214786
R31984 DVDD.n15632 DVDD.n15631 0.214786
R31985 DVDD.n15535 DVDD.n5117 0.214786
R31986 DVDD.n15682 DVDD.n15681 0.214786
R31987 DVDD.n15683 DVDD.n5112 0.214786
R31988 DVDD.n15685 DVDD.n15684 0.214786
R31989 DVDD.n15687 DVDD.n5110 0.214786
R31990 DVDD.n15689 DVDD.n15688 0.214786
R31991 DVDD.n15691 DVDD.n15690 0.214786
R31992 DVDD.n15693 DVDD.n15692 0.214786
R31993 DVDD.n15695 DVDD.n15694 0.214786
R31994 DVDD.n15697 DVDD.n15696 0.214786
R31995 DVDD.n5083 DVDD.n5082 0.214786
R31996 DVDD.n5101 DVDD.n5100 0.214786
R31997 DVDD.n5099 DVDD.n5098 0.214786
R31998 DVDD.n5097 DVDD.n5096 0.214786
R31999 DVDD.n5086 DVDD.n5085 0.214786
R32000 DVDD.n5092 DVDD.n5091 0.214786
R32001 DVDD.n5090 DVDD.n5089 0.214786
R32002 DVDD.n5088 DVDD.n5065 0.214786
R32003 DVDD.n16215 DVDD.n16214 0.214786
R32004 DVDD.n16217 DVDD.n16216 0.214786
R32005 DVDD.n16219 DVDD.n16218 0.214786
R32006 DVDD.n16221 DVDD.n16220 0.214786
R32007 DVDD.n16223 DVDD.n16222 0.214786
R32008 DVDD.n16225 DVDD.n16224 0.214786
R32009 DVDD.n16227 DVDD.n16226 0.214786
R32010 DVDD.n16229 DVDD.n16228 0.214786
R32011 DVDD.n16231 DVDD.n16230 0.214786
R32012 DVDD.n16233 DVDD.n16232 0.214786
R32013 DVDD.n16235 DVDD.n16234 0.214786
R32014 DVDD.n16236 DVDD.n670 0.214786
R32015 DVDD.n16237 DVDD.n656 0.214786
R32016 DVDD.n16239 DVDD.n16238 0.214786
R32017 DVDD.n16242 DVDD.n16241 0.214786
R32018 DVDD.n16243 DVDD.n2833 0.214786
R32019 DVDD.n16245 DVDD.n16244 0.214786
R32020 DVDD.n2834 DVDD.n2832 0.214786
R32021 DVDD.n2876 DVDD.n2875 0.214786
R32022 DVDD.n2874 DVDD.n2873 0.214786
R32023 DVDD.n2865 DVDD.n2864 0.214786
R32024 DVDD.n2837 DVDD.n2836 0.214786
R32025 DVDD.n2860 DVDD.n2859 0.214786
R32026 DVDD.n2858 DVDD.n2857 0.214786
R32027 DVDD.n2856 DVDD.n2855 0.214786
R32028 DVDD.n2840 DVDD.n2839 0.214786
R32029 DVDD.n2851 DVDD.n2850 0.214786
R32030 DVDD.n2849 DVDD.n2848 0.214786
R32031 DVDD.n2847 DVDD.n2846 0.214786
R32032 DVDD.n2842 DVDD.n2792 0.214786
R32033 DVDD.n16249 DVDD.n2779 0.214786
R32034 DVDD.n16251 DVDD.n16250 0.214786
R32035 DVDD.n16252 DVDD.n2770 0.214786
R32036 DVDD.n16254 DVDD.n16253 0.214786
R32037 DVDD.n2771 DVDD.n2767 0.214786
R32038 DVDD.n2773 DVDD.n2772 0.214786
R32039 DVDD.n2765 DVDD.n2709 0.214786
R32040 DVDD.n16259 DVDD.n16258 0.214786
R32041 DVDD.n15961 DVDD.n15960 0.214786
R32042 DVDD.n15963 DVDD.n15962 0.214786
R32043 DVDD.n15965 DVDD.n15964 0.214786
R32044 DVDD.n15967 DVDD.n15966 0.214786
R32045 DVDD.n15969 DVDD.n15968 0.214786
R32046 DVDD.n15971 DVDD.n15970 0.214786
R32047 DVDD.n15973 DVDD.n15972 0.214786
R32048 DVDD.n15975 DVDD.n15974 0.214786
R32049 DVDD.n15977 DVDD.n15976 0.214786
R32050 DVDD.n15978 DVDD.n15948 0.214786
R32051 DVDD.n15980 DVDD.n15979 0.214786
R32052 DVDD.n15981 DVDD.n15947 0.214786
R32053 DVDD.n15983 DVDD.n15982 0.214786
R32054 DVDD.n15984 DVDD.n3202 0.214786
R32055 DVDD.n15986 DVDD.n15985 0.214786
R32056 DVDD.n3203 DVDD.n3201 0.214786
R32057 DVDD.n15941 DVDD.n15940 0.214786
R32058 DVDD.n15939 DVDD.n15938 0.214786
R32059 DVDD.n15929 DVDD.n15928 0.214786
R32060 DVDD.n3206 DVDD.n3205 0.214786
R32061 DVDD.n15924 DVDD.n15923 0.214786
R32062 DVDD.n15922 DVDD.n15921 0.214786
R32063 DVDD.n15920 DVDD.n15919 0.214786
R32064 DVDD.n3208 DVDD.n3162 0.214786
R32065 DVDD.n15914 DVDD.n3149 0.214786
R32066 DVDD.n3230 DVDD.n3229 0.214786
R32067 DVDD.n15508 DVDD.n15507 0.214786
R32068 DVDD.n15510 DVDD.n15509 0.214786
R32069 DVDD.n15512 DVDD.n15511 0.214786
R32070 DVDD.n15513 DVDD.n15502 0.214786
R32071 DVDD.n15515 DVDD.n15514 0.214786
R32072 DVDD.n15516 DVDD.n5159 0.214786
R32073 DVDD.n15517 DVDD.n5144 0.214786
R32074 DVDD.n15519 DVDD.n15518 0.214786
R32075 DVDD.n5215 DVDD.n5208 0.214786
R32076 DVDD.n15495 DVDD.n15494 0.214786
R32077 DVDD.n15493 DVDD.n15492 0.214786
R32078 DVDD.n15491 DVDD.n15490 0.214786
R32079 DVDD.n5218 DVDD.n5217 0.214786
R32080 DVDD.n15486 DVDD.n15485 0.214786
R32081 DVDD.n15484 DVDD.n15483 0.214786
R32082 DVDD.n15482 DVDD.n15481 0.214786
R32083 DVDD.n5221 DVDD.n5220 0.214786
R32084 DVDD.n15477 DVDD.n15476 0.214786
R32085 DVDD.n15475 DVDD.n15474 0.214786
R32086 DVDD.n15473 DVDD.n15472 0.214786
R32087 DVDD.n15471 DVDD.n5223 0.214786
R32088 DVDD.n15470 DVDD.n15469 0.214786
R32089 DVDD.n15464 DVDD.n15463 0.214786
R32090 DVDD.n15462 DVDD.n5228 0.214786
R32091 DVDD.n15436 DVDD.n5229 0.214786
R32092 DVDD.n15438 DVDD.n15437 0.214786
R32093 DVDD.n15440 DVDD.n15439 0.214786
R32094 DVDD.n15442 DVDD.n15441 0.214786
R32095 DVDD.n15444 DVDD.n15443 0.214786
R32096 DVDD.n15446 DVDD.n15445 0.214786
R32097 DVDD.n15448 DVDD.n15447 0.214786
R32098 DVDD.n15450 DVDD.n15449 0.214786
R32099 DVDD.n15452 DVDD.n15451 0.214786
R32100 DVDD.n15454 DVDD.n15453 0.214786
R32101 DVDD.n15456 DVDD.n15455 0.214786
R32102 DVDD.n15458 DVDD.n15457 0.214786
R32103 DVDD.n2896 DVDD.n746 0.214786
R32104 DVDD.n2898 DVDD.n2897 0.214786
R32105 DVDD.n2900 DVDD.n2899 0.214786
R32106 DVDD.n2902 DVDD.n2901 0.214786
R32107 DVDD.n2904 DVDD.n2903 0.214786
R32108 DVDD.n2906 DVDD.n2905 0.214786
R32109 DVDD.n2908 DVDD.n2907 0.214786
R32110 DVDD.n2910 DVDD.n2909 0.214786
R32111 DVDD.n2912 DVDD.n2911 0.214786
R32112 DVDD.n2914 DVDD.n2913 0.214786
R32113 DVDD.n2916 DVDD.n2915 0.214786
R32114 DVDD.n15326 DVDD.n15325 0.214786
R32115 DVDD.n15328 DVDD.n15327 0.214786
R32116 DVDD.n15330 DVDD.n15329 0.214786
R32117 DVDD.n15322 DVDD.n15321 0.214786
R32118 DVDD.n15335 DVDD.n15334 0.214786
R32119 DVDD.n15337 DVDD.n15336 0.214786
R32120 DVDD.n15339 DVDD.n15338 0.214786
R32121 DVDD.n15319 DVDD.n15318 0.214786
R32122 DVDD.n15405 DVDD.n15404 0.214786
R32123 DVDD.n15403 DVDD.n15402 0.214786
R32124 DVDD.n15401 DVDD.n15400 0.214786
R32125 DVDD.n15399 DVDD.n5382 0.214786
R32126 DVDD.n15398 DVDD.n5394 0.214786
R32127 DVDD.n15397 DVDD.n15396 0.214786
R32128 DVDD.n15394 DVDD.n15393 0.214786
R32129 DVDD.n15392 DVDD.n15349 0.214786
R32130 DVDD.n15391 DVDD.n15390 0.214786
R32131 DVDD.n15389 DVDD.n15388 0.214786
R32132 DVDD.n15387 DVDD.n15386 0.214786
R32133 DVDD.n15385 DVDD.n15384 0.214786
R32134 DVDD.n15383 DVDD.n15382 0.214786
R32135 DVDD.n15381 DVDD.n15380 0.214786
R32136 DVDD.n15379 DVDD.n15378 0.214786
R32137 DVDD.n15377 DVDD.n15376 0.214786
R32138 DVDD.n15375 DVDD.n15374 0.214786
R32139 DVDD.n15373 DVDD.n15372 0.214786
R32140 DVDD.n15371 DVDD.n15370 0.214786
R32141 DVDD.n15369 DVDD.n15368 0.214786
R32142 DVDD.n15367 DVDD.n15366 0.214786
R32143 DVDD.n3138 DVDD.n3123 0.214786
R32144 DVDD.n16006 DVDD.n16005 0.214786
R32145 DVDD.n16004 DVDD.n3137 0.214786
R32146 DVDD.n16003 DVDD.n16002 0.214786
R32147 DVDD.n16001 DVDD.n16000 0.214786
R32148 DVDD.n15999 DVDD.n15998 0.214786
R32149 DVDD.n15997 DVDD.n15996 0.214786
R32150 DVDD.n15995 DVDD.n15994 0.214786
R32151 DVDD.n15993 DVDD.n15992 0.214786
R32152 DVDD.n3224 DVDD.n3223 0.214786
R32153 DVDD.n3222 DVDD.n3221 0.214786
R32154 DVDD.n3220 DVDD.n3219 0.214786
R32155 DVDD.n3218 DVDD.n3217 0.214786
R32156 DVDD.n3216 DVDD.n3215 0.214786
R32157 DVDD.n3214 DVDD.n3087 0.214786
R32158 DVDD.n16075 DVDD.n3056 0.214786
R32159 DVDD.n16087 DVDD.n16086 0.214786
R32160 DVDD.n3068 DVDD.n3054 0.214786
R32161 DVDD.n16092 DVDD.n16091 0.214786
R32162 DVDD.n16093 DVDD.n3052 0.214786
R32163 DVDD.n16095 DVDD.n16094 0.214786
R32164 DVDD.n3050 DVDD.n3049 0.214786
R32165 DVDD.n16101 DVDD.n16100 0.214786
R32166 DVDD.n16102 DVDD.n3047 0.214786
R32167 DVDD.n16115 DVDD.n16114 0.214786
R32168 DVDD.n16117 DVDD.n16116 0.214786
R32169 DVDD.n16119 DVDD.n16118 0.214786
R32170 DVDD.n3045 DVDD.n3044 0.214786
R32171 DVDD.n16124 DVDD.n16123 0.214786
R32172 DVDD.n16126 DVDD.n16125 0.214786
R32173 DVDD.n16128 DVDD.n16127 0.214786
R32174 DVDD.n3042 DVDD.n3041 0.214786
R32175 DVDD.n16133 DVDD.n16132 0.214786
R32176 DVDD.n16136 DVDD.n16135 0.214786
R32177 DVDD.n16140 DVDD.n16139 0.214786
R32178 DVDD.n16141 DVDD.n2994 0.214786
R32179 DVDD.n16146 DVDD.n16145 0.214786
R32180 DVDD.n2992 DVDD.n2991 0.214786
R32181 DVDD.n16152 DVDD.n16151 0.214786
R32182 DVDD.n16153 DVDD.n2990 0.214786
R32183 DVDD.n16155 DVDD.n16154 0.214786
R32184 DVDD.n16157 DVDD.n16156 0.214786
R32185 DVDD.n2988 DVDD.n2987 0.214786
R32186 DVDD.n16162 DVDD.n16161 0.214786
R32187 DVDD.n16164 DVDD.n16163 0.214786
R32188 DVDD.n16166 DVDD.n16165 0.214786
R32189 DVDD.n2985 DVDD.n2984 0.214786
R32190 DVDD.n16171 DVDD.n16170 0.214786
R32191 DVDD.n16173 DVDD.n16172 0.214786
R32192 DVDD.n16175 DVDD.n16174 0.214786
R32193 DVDD.n2982 DVDD.n2981 0.214786
R32194 DVDD.n16180 DVDD.n16179 0.214786
R32195 DVDD.n16181 DVDD.n2923 0.214786
R32196 DVDD.n16186 DVDD.n16185 0.214786
R32197 DVDD.n2921 DVDD.n2920 0.214786
R32198 DVDD.n16193 DVDD.n16192 0.214786
R32199 DVDD.n16194 DVDD.n2882 0.214786
R32200 DVDD.n16198 DVDD.n16197 0.214786
R32201 DVDD.n16196 DVDD.n2919 0.214786
R32202 DVDD.n2918 DVDD.n2917 0.214786
R32203 DVDD.n20483 DVDD 0.19085
R32204 DVDD DVDD.n20482 0.19085
R32205 DVDD.n20950 DVDD 0.19085
R32206 DVDD DVDD.n20949 0.19085
R32207 DVDD.n19122 DVDD 0.19085
R32208 DVDD DVDD.n19121 0.19085
R32209 DVDD.n21054 DVDD 0.19085
R32210 DVDD DVDD.n21053 0.19085
R32211 DVDD.n18618 DVDD.n18616 0.182868
R32212 DVDD.n4982 DVDD.n4981 0.177076
R32213 DVDD.n2474 DVDD.n550 0.177076
R32214 DVDD.n10177 DVDD.n5568 0.177076
R32215 DVDD.n16450 DVDD.n888 0.177076
R32216 DVDD.n20924 DVDD.n18906 0.168198
R32217 DVDD.n19099 DVDD.n19097 0.168198
R32218 DVDD.n20141 DVDD.n20140 0.158302
R32219 DVDD.n20336 DVDD.n18950 0.158302
R32220 DVDD.n20628 DVDD.n20627 0.158302
R32221 DVDD.n20849 DVDD.n18979 0.158302
R32222 DVDD.n3964 DVDD.n3934 0.158302
R32223 DVDD.n22119 DVDD.n22088 0.158302
R32224 DVDD.n9840 DVDD.n5486 0.158302
R32225 DVDD.n10019 DVDD.n10018 0.158302
R32226 DVDD.n22348 DVDD.n22347 0.157978
R32227 DVDD.n19651 DVDD.n19650 0.157978
R32228 DVDD.n19412 DVDD.n19411 0.142605
R32229 DVDD.n21495 DVDD.n21494 0.142605
R32230 DVDD.n19335 DVDD.n19334 0.142605
R32231 DVDD.n4381 DVDD.n4354 0.1405
R32232 DVDD.n4838 DVDD.n3565 0.140149
R32233 DVDD.n18197 DVDD.n18162 0.137029
R32234 DVDD.n20656 DVDD.n20596 0.130621
R32235 DVDD.n20856 DVDD.n20855 0.130621
R32236 DVDD.n20488 DVDD.n19773 0.125228
R32237 DVDD.n20463 DVDD.n18909 0.125228
R32238 DVDD.n20983 DVDD.n18751 0.125228
R32239 DVDD.n21050 DVDD.n21049 0.125228
R32240 DVDD.n19411 DVDD.n19313 0.123658
R32241 DVDD.n19360 DVDD.n19313 0.123658
R32242 DVDD.n19361 DVDD.n19360 0.123658
R32243 DVDD.n19362 DVDD.n19361 0.123658
R32244 DVDD.n19363 DVDD.n19362 0.123658
R32245 DVDD.n19365 DVDD.n19363 0.123658
R32246 DVDD.n19366 DVDD.n19365 0.123658
R32247 DVDD.n19367 DVDD.n19366 0.123658
R32248 DVDD.n19368 DVDD.n19367 0.123658
R32249 DVDD.n19370 DVDD.n19368 0.123658
R32250 DVDD.n19371 DVDD.n19370 0.123658
R32251 DVDD.n19372 DVDD.n19371 0.123658
R32252 DVDD.n19373 DVDD.n19372 0.123658
R32253 DVDD.n19374 DVDD.n19373 0.123658
R32254 DVDD.n19376 DVDD.n19374 0.123658
R32255 DVDD.n19376 DVDD.n19375 0.123658
R32256 DVDD.n21279 DVDD.n21278 0.123658
R32257 DVDD.n21280 DVDD.n21279 0.123658
R32258 DVDD.n21280 DVDD.n18641 0.123658
R32259 DVDD.n21291 DVDD.n18641 0.123658
R32260 DVDD.n21292 DVDD.n21291 0.123658
R32261 DVDD.n21293 DVDD.n21292 0.123658
R32262 DVDD.n21293 DVDD.n18633 0.123658
R32263 DVDD.n21303 DVDD.n18633 0.123658
R32264 DVDD.n21304 DVDD.n21303 0.123658
R32265 DVDD.n21305 DVDD.n21304 0.123658
R32266 DVDD.n21305 DVDD.n18626 0.123658
R32267 DVDD.n21316 DVDD.n18626 0.123658
R32268 DVDD.n21317 DVDD.n21316 0.123658
R32269 DVDD.n21319 DVDD.n21317 0.123658
R32270 DVDD.n21319 DVDD.n21318 0.123658
R32271 DVDD.n21318 DVDD.n18618 0.123658
R32272 DVDD.n21494 DVDD.n21493 0.123658
R32273 DVDD.n21493 DVDD.n21325 0.123658
R32274 DVDD.n21326 DVDD.n21325 0.123658
R32275 DVDD.n21486 DVDD.n21326 0.123658
R32276 DVDD.n21486 DVDD.n21485 0.123658
R32277 DVDD.n21485 DVDD.n21484 0.123658
R32278 DVDD.n21484 DVDD.n21328 0.123658
R32279 DVDD.n21479 DVDD.n21478 0.123658
R32280 DVDD.n21478 DVDD.n21477 0.123658
R32281 DVDD.n21477 DVDD.n21372 0.123658
R32282 DVDD.n21472 DVDD.n21372 0.123658
R32283 DVDD.n21472 DVDD.n21471 0.123658
R32284 DVDD.n21471 DVDD.n21470 0.123658
R32285 DVDD.n21470 DVDD.n21375 0.123658
R32286 DVDD.n21465 DVDD.n21375 0.123658
R32287 DVDD.n21465 DVDD.n21464 0.123658
R32288 DVDD.n21464 DVDD.n21463 0.123658
R32289 DVDD.n21463 DVDD.n21378 0.123658
R32290 DVDD.n21458 DVDD.n21378 0.123658
R32291 DVDD.n21458 DVDD.n21457 0.123658
R32292 DVDD.n21457 DVDD.n21456 0.123658
R32293 DVDD.n21456 DVDD.n21381 0.123658
R32294 DVDD.n21451 DVDD.n21381 0.123658
R32295 DVDD.n21451 DVDD.n21450 0.123658
R32296 DVDD.n21450 DVDD.n21449 0.123658
R32297 DVDD.n21449 DVDD.n21384 0.123658
R32298 DVDD.n21444 DVDD.n21384 0.123658
R32299 DVDD.n21444 DVDD.n21443 0.123658
R32300 DVDD.n21440 DVDD.n21387 0.123658
R32301 DVDD.n21435 DVDD.n21387 0.123658
R32302 DVDD.n21435 DVDD.n21434 0.123658
R32303 DVDD.n21434 DVDD.n21433 0.123658
R32304 DVDD.n21433 DVDD.n21390 0.123658
R32305 DVDD.n21428 DVDD.n21390 0.123658
R32306 DVDD.n21428 DVDD.n21427 0.123658
R32307 DVDD.n21427 DVDD.n21426 0.123658
R32308 DVDD.n21426 DVDD.n21393 0.123658
R32309 DVDD.n21421 DVDD.n21393 0.123658
R32310 DVDD.n21421 DVDD.n21420 0.123658
R32311 DVDD.n21420 DVDD.n21419 0.123658
R32312 DVDD.n21419 DVDD.n21396 0.123658
R32313 DVDD.n21414 DVDD.n21396 0.123658
R32314 DVDD.n21414 DVDD.n21413 0.123658
R32315 DVDD.n21413 DVDD.n21412 0.123658
R32316 DVDD.n21412 DVDD.n21399 0.123658
R32317 DVDD.n21407 DVDD.n21399 0.123658
R32318 DVDD.n21407 DVDD.n21406 0.123658
R32319 DVDD.n21406 DVDD.n21405 0.123658
R32320 DVDD.n21405 DVDD.n18557 0.123658
R32321 DVDD.n21644 DVDD.n18558 0.123658
R32322 DVDD.n21639 DVDD.n18558 0.123658
R32323 DVDD.n21639 DVDD.n21638 0.123658
R32324 DVDD.n21638 DVDD.n21637 0.123658
R32325 DVDD.n21637 DVDD.n18562 0.123658
R32326 DVDD.n21632 DVDD.n18562 0.123658
R32327 DVDD.n21632 DVDD.n21631 0.123658
R32328 DVDD.n21631 DVDD.n21630 0.123658
R32329 DVDD.n21630 DVDD.n18565 0.123658
R32330 DVDD.n21625 DVDD.n18565 0.123658
R32331 DVDD.n21625 DVDD.n21624 0.123658
R32332 DVDD.n21624 DVDD.n21623 0.123658
R32333 DVDD.n21623 DVDD.n18568 0.123658
R32334 DVDD.n21618 DVDD.n18568 0.123658
R32335 DVDD.n21618 DVDD.n21617 0.123658
R32336 DVDD.n21617 DVDD.n21616 0.123658
R32337 DVDD.n21616 DVDD.n18571 0.123658
R32338 DVDD.n21611 DVDD.n18571 0.123658
R32339 DVDD.n21611 DVDD.n21610 0.123658
R32340 DVDD.n21610 DVDD.n21609 0.123658
R32341 DVDD.n21609 DVDD.n18574 0.123658
R32342 DVDD.n21604 DVDD.n18574 0.123658
R32343 DVDD.n21604 DVDD.n21603 0.123658
R32344 DVDD.n21603 DVDD.n21602 0.123658
R32345 DVDD.n21602 DVDD.n18577 0.123658
R32346 DVDD.n21597 DVDD.n18577 0.123658
R32347 DVDD.n21581 DVDD.n21580 0.123658
R32348 DVDD.n21580 DVDD.n18580 0.123658
R32349 DVDD.n21575 DVDD.n18580 0.123658
R32350 DVDD.n21575 DVDD.n21574 0.123658
R32351 DVDD.n21574 DVDD.n21573 0.123658
R32352 DVDD.n21573 DVDD.n18583 0.123658
R32353 DVDD.n21568 DVDD.n18583 0.123658
R32354 DVDD.n21568 DVDD.n21567 0.123658
R32355 DVDD.n21567 DVDD.n21566 0.123658
R32356 DVDD.n21566 DVDD.n18586 0.123658
R32357 DVDD.n21561 DVDD.n18586 0.123658
R32358 DVDD.n21561 DVDD.n21560 0.123658
R32359 DVDD.n21560 DVDD.n21559 0.123658
R32360 DVDD.n21559 DVDD.n18589 0.123658
R32361 DVDD.n21554 DVDD.n18589 0.123658
R32362 DVDD.n21554 DVDD.n21553 0.123658
R32363 DVDD.n21553 DVDD.n21552 0.123658
R32364 DVDD.n21552 DVDD.n18592 0.123658
R32365 DVDD.n21547 DVDD.n18592 0.123658
R32366 DVDD.n21547 DVDD.n21546 0.123658
R32367 DVDD.n21546 DVDD.n21545 0.123658
R32368 DVDD.n21540 DVDD.n18597 0.123658
R32369 DVDD.n21540 DVDD.n21539 0.123658
R32370 DVDD.n21539 DVDD.n21538 0.123658
R32371 DVDD.n21538 DVDD.n18599 0.123658
R32372 DVDD.n21533 DVDD.n18599 0.123658
R32373 DVDD.n21533 DVDD.n21532 0.123658
R32374 DVDD.n21532 DVDD.n21531 0.123658
R32375 DVDD.n21531 DVDD.n18602 0.123658
R32376 DVDD.n21526 DVDD.n18602 0.123658
R32377 DVDD.n21526 DVDD.n21525 0.123658
R32378 DVDD.n21525 DVDD.n21524 0.123658
R32379 DVDD.n21524 DVDD.n18605 0.123658
R32380 DVDD.n21519 DVDD.n18605 0.123658
R32381 DVDD.n21519 DVDD.n21518 0.123658
R32382 DVDD.n21518 DVDD.n21517 0.123658
R32383 DVDD.n21517 DVDD.n18608 0.123658
R32384 DVDD.n21512 DVDD.n18608 0.123658
R32385 DVDD.n21512 DVDD.n21511 0.123658
R32386 DVDD.n21511 DVDD.n21510 0.123658
R32387 DVDD.n21510 DVDD.n18611 0.123658
R32388 DVDD.n21505 DVDD.n21504 0.123658
R32389 DVDD.n19406 DVDD.n19335 0.123658
R32390 DVDD.n19406 DVDD.n19405 0.123658
R32391 DVDD.n19405 DVDD.n19404 0.123658
R32392 DVDD.n19404 DVDD.n19336 0.123658
R32393 DVDD.n19398 DVDD.n19336 0.123658
R32394 DVDD.n19398 DVDD.n19397 0.123658
R32395 DVDD.n19397 DVDD.n19396 0.123658
R32396 DVDD.n19396 DVDD.n19344 0.123658
R32397 DVDD.n19390 DVDD.n19344 0.123658
R32398 DVDD.n19390 DVDD.n19389 0.123658
R32399 DVDD.n19389 DVDD.n19388 0.123658
R32400 DVDD.n19388 DVDD.n19350 0.123658
R32401 DVDD.n19382 DVDD.n19350 0.123658
R32402 DVDD.n19382 DVDD.n19381 0.123658
R32403 DVDD.n19381 DVDD.n19380 0.123658
R32404 DVDD.n19380 DVDD.n18652 0.123658
R32405 DVDD.n21274 DVDD.n18644 0.123658
R32406 DVDD.n21285 DVDD.n18644 0.123658
R32407 DVDD.n21286 DVDD.n21285 0.123658
R32408 DVDD.n21287 DVDD.n21286 0.123658
R32409 DVDD.n21287 DVDD.n18637 0.123658
R32410 DVDD.n21297 DVDD.n18637 0.123658
R32411 DVDD.n21298 DVDD.n21297 0.123658
R32412 DVDD.n21299 DVDD.n21298 0.123658
R32413 DVDD.n21299 DVDD.n18629 0.123658
R32414 DVDD.n21310 DVDD.n18629 0.123658
R32415 DVDD.n21311 DVDD.n21310 0.123658
R32416 DVDD.n21312 DVDD.n21311 0.123658
R32417 DVDD.n21312 DVDD.n18622 0.123658
R32418 DVDD.n21323 DVDD.n18622 0.123658
R32419 DVDD.n21324 DVDD.n21323 0.123658
R32420 DVDD.n21495 DVDD.n21324 0.123658
R32421 DVDD.n19334 DVDD.n19317 0.123658
R32422 DVDD.n19329 DVDD.n19317 0.123658
R32423 DVDD.n19329 DVDD.n19328 0.123658
R32424 DVDD.n19328 DVDD.n19327 0.123658
R32425 DVDD.n19327 DVDD.n19319 0.123658
R32426 DVDD.n19322 DVDD.n19319 0.123658
R32427 DVDD.n19322 DVDD.n19215 0.123658
R32428 DVDD.n19631 DVDD.n19216 0.123658
R32429 DVDD.n19626 DVDD.n19216 0.123658
R32430 DVDD.n19626 DVDD.n19625 0.123658
R32431 DVDD.n19625 DVDD.n19624 0.123658
R32432 DVDD.n19624 DVDD.n19220 0.123658
R32433 DVDD.n19619 DVDD.n19220 0.123658
R32434 DVDD.n19619 DVDD.n19618 0.123658
R32435 DVDD.n19618 DVDD.n19617 0.123658
R32436 DVDD.n19617 DVDD.n19223 0.123658
R32437 DVDD.n19612 DVDD.n19223 0.123658
R32438 DVDD.n19612 DVDD.n19611 0.123658
R32439 DVDD.n19611 DVDD.n19610 0.123658
R32440 DVDD.n19610 DVDD.n19226 0.123658
R32441 DVDD.n19605 DVDD.n19226 0.123658
R32442 DVDD.n19605 DVDD.n19604 0.123658
R32443 DVDD.n19604 DVDD.n19603 0.123658
R32444 DVDD.n19603 DVDD.n19229 0.123658
R32445 DVDD.n19598 DVDD.n19229 0.123658
R32446 DVDD.n19598 DVDD.n19597 0.123658
R32447 DVDD.n19597 DVDD.n19596 0.123658
R32448 DVDD.n19596 DVDD.n19232 0.123658
R32449 DVDD.n19591 DVDD.n19590 0.123658
R32450 DVDD.n19590 DVDD.n19589 0.123658
R32451 DVDD.n19589 DVDD.n19237 0.123658
R32452 DVDD.n19584 DVDD.n19237 0.123658
R32453 DVDD.n19584 DVDD.n19583 0.123658
R32454 DVDD.n19583 DVDD.n19582 0.123658
R32455 DVDD.n19582 DVDD.n19240 0.123658
R32456 DVDD.n19577 DVDD.n19240 0.123658
R32457 DVDD.n19577 DVDD.n19576 0.123658
R32458 DVDD.n19576 DVDD.n19575 0.123658
R32459 DVDD.n19575 DVDD.n19243 0.123658
R32460 DVDD.n19570 DVDD.n19243 0.123658
R32461 DVDD.n19570 DVDD.n19569 0.123658
R32462 DVDD.n19569 DVDD.n19568 0.123658
R32463 DVDD.n19568 DVDD.n19246 0.123658
R32464 DVDD.n19563 DVDD.n19246 0.123658
R32465 DVDD.n19563 DVDD.n19562 0.123658
R32466 DVDD.n19562 DVDD.n19561 0.123658
R32467 DVDD.n19561 DVDD.n19249 0.123658
R32468 DVDD.n19556 DVDD.n19249 0.123658
R32469 DVDD.n19556 DVDD.n19555 0.123658
R32470 DVDD.n19552 DVDD.n19252 0.123658
R32471 DVDD.n19547 DVDD.n19252 0.123658
R32472 DVDD.n19547 DVDD.n19546 0.123658
R32473 DVDD.n19546 DVDD.n19545 0.123658
R32474 DVDD.n19545 DVDD.n19255 0.123658
R32475 DVDD.n19540 DVDD.n19255 0.123658
R32476 DVDD.n19540 DVDD.n19539 0.123658
R32477 DVDD.n19539 DVDD.n19538 0.123658
R32478 DVDD.n19538 DVDD.n19258 0.123658
R32479 DVDD.n19533 DVDD.n19258 0.123658
R32480 DVDD.n19533 DVDD.n19532 0.123658
R32481 DVDD.n19532 DVDD.n19531 0.123658
R32482 DVDD.n19531 DVDD.n19261 0.123658
R32483 DVDD.n19526 DVDD.n19261 0.123658
R32484 DVDD.n19526 DVDD.n19525 0.123658
R32485 DVDD.n19525 DVDD.n19524 0.123658
R32486 DVDD.n19524 DVDD.n19264 0.123658
R32487 DVDD.n19519 DVDD.n19264 0.123658
R32488 DVDD.n19519 DVDD.n19518 0.123658
R32489 DVDD.n19518 DVDD.n19517 0.123658
R32490 DVDD.n19517 DVDD.n19267 0.123658
R32491 DVDD.n19512 DVDD.n19267 0.123658
R32492 DVDD.n19512 DVDD.n19511 0.123658
R32493 DVDD.n19511 DVDD.n19510 0.123658
R32494 DVDD.n19510 DVDD.n19270 0.123658
R32495 DVDD.n19505 DVDD.n19270 0.123658
R32496 DVDD.n19502 DVDD.n19501 0.123658
R32497 DVDD.n19501 DVDD.n19273 0.123658
R32498 DVDD.n19496 DVDD.n19273 0.123658
R32499 DVDD.n19496 DVDD.n19495 0.123658
R32500 DVDD.n19495 DVDD.n19494 0.123658
R32501 DVDD.n19494 DVDD.n19276 0.123658
R32502 DVDD.n19489 DVDD.n19276 0.123658
R32503 DVDD.n19489 DVDD.n19488 0.123658
R32504 DVDD.n19488 DVDD.n19487 0.123658
R32505 DVDD.n19487 DVDD.n19279 0.123658
R32506 DVDD.n19482 DVDD.n19279 0.123658
R32507 DVDD.n19482 DVDD.n19481 0.123658
R32508 DVDD.n19481 DVDD.n19480 0.123658
R32509 DVDD.n19480 DVDD.n19282 0.123658
R32510 DVDD.n19475 DVDD.n19282 0.123658
R32511 DVDD.n19475 DVDD.n19474 0.123658
R32512 DVDD.n19474 DVDD.n19473 0.123658
R32513 DVDD.n19473 DVDD.n19285 0.123658
R32514 DVDD.n19468 DVDD.n19285 0.123658
R32515 DVDD.n19468 DVDD.n19467 0.123658
R32516 DVDD.n19467 DVDD.n19466 0.123658
R32517 DVDD.n19461 DVDD.n19291 0.123658
R32518 DVDD.n19461 DVDD.n19460 0.123658
R32519 DVDD.n19460 DVDD.n19459 0.123658
R32520 DVDD.n19459 DVDD.n19293 0.123658
R32521 DVDD.n19454 DVDD.n19293 0.123658
R32522 DVDD.n19454 DVDD.n19453 0.123658
R32523 DVDD.n19453 DVDD.n19452 0.123658
R32524 DVDD.n19452 DVDD.n19296 0.123658
R32525 DVDD.n19447 DVDD.n19296 0.123658
R32526 DVDD.n19447 DVDD.n19446 0.123658
R32527 DVDD.n19446 DVDD.n19445 0.123658
R32528 DVDD.n19445 DVDD.n19299 0.123658
R32529 DVDD.n19440 DVDD.n19299 0.123658
R32530 DVDD.n19440 DVDD.n19439 0.123658
R32531 DVDD.n19439 DVDD.n19438 0.123658
R32532 DVDD.n19438 DVDD.n19302 0.123658
R32533 DVDD.n19433 DVDD.n19302 0.123658
R32534 DVDD.n19433 DVDD.n19432 0.123658
R32535 DVDD.n19432 DVDD.n19431 0.123658
R32536 DVDD.n19431 DVDD.n19305 0.123658
R32537 DVDD.n19426 DVDD.n19305 0.123658
R32538 DVDD.n19424 DVDD.n19423 0.123658
R32539 DVDD.n19423 DVDD.n19308 0.123658
R32540 DVDD.n19418 DVDD.n19308 0.123658
R32541 DVDD.n19417 DVDD.n19416 0.123658
R32542 DVDD.n19416 DVDD.n19311 0.123658
R32543 DVDD.n19412 DVDD.n19311 0.123658
R32544 DVDD.n21645 DVDD.n18557 0.122474
R32545 DVDD.n21596 DVDD.n21581 0.122474
R32546 DVDD.n19555 DVDD.n19554 0.122474
R32547 DVDD.n19504 DVDD.n19502 0.122474
R32548 DVDD.n21273 DVDD.n21272 0.122122
R32549 DVDD.n18648 DVDD.n128 0.122122
R32550 DVDD.n15459 DVDD.n15424 0.112533
R32551 DVDD.n15700 DVDD.n5053 0.112533
R32552 DVDD.n15750 DVDD.n15715 0.112533
R32553 DVDD.n15324 DVDD.n5379 0.112533
R32554 DVDD.n16213 DVDD.n652 0.112413
R32555 DVDD.n16334 DVDD.n565 0.112413
R32556 DVDD.n18043 DVDD.n530 0.112413
R32557 DVDD.n17954 DVDD.n761 0.112413
R32558 DVDD.n21251 DVDD.n21249 0.110634
R32559 DVDD.n22030 DVDD.n234 0.110634
R32560 DVDD.n21230 DVDD.n21228 0.110634
R32561 DVDD.n22188 DVDD.n22187 0.110634
R32562 DVDD.n18455 DVDD.n126 0.110634
R32563 DVDD.n18236 DVDD.n18235 0.110634
R32564 DVDD.n18487 DVDD.n122 0.110634
R32565 DVDD.n22055 DVDD.n22054 0.110634
R32566 DVDD.n21505 DVDD.n18614 0.109447
R32567 DVDD.n4979 DVDD.n4978 0.104685
R32568 DVDD.n16397 DVDD.n2324 0.104685
R32569 DVDD.n10204 DVDD.n10203 0.104685
R32570 DVDD.n16433 DVDD.n16432 0.104685
R32571 DVDD.n20539 DVDD.n19789 0.103951
R32572 DVDD.n19817 DVDD.n19789 0.103951
R32573 DVDD.n21082 DVDD.n18753 0.103951
R32574 DVDD.n18799 DVDD.n18753 0.103951
R32575 DVDD DVDD.n19417 0.102342
R32576 DVDD.n21442 DVDD.n21440 0.0987895
R32577 DVDD.n21545 DVDD.n18595 0.0987895
R32578 DVDD.n19591 DVDD.n19236 0.0987895
R32579 DVDD.n19466 DVDD.n19289 0.0987895
R32580 DVDD.n16400 DVDD.n2293 0.0936793
R32581 DVDD.n16400 DVDD.n16399 0.0936793
R32582 DVDD.n16404 DVDD.n2291 0.0936793
R32583 DVDD.n16406 DVDD.n16404 0.0936793
R32584 DVDD.n19703 DVDD.n19702 0.0933421
R32585 DVDD.n18981 DVDD.n30 0.0933421
R32586 DVDD.n4881 DVDD.n4880 0.0930579
R32587 DVDD.n18045 DVDD.n18044 0.0930579
R32588 DVDD DVDD.t132 0.092694
R32589 DVDD DVDD.t122 0.092694
R32590 DVDD DVDD.t79 0.092694
R32591 DVDD DVDD.t139 0.092694
R32592 DVDD DVDD.t100 0.092694
R32593 DVDD DVDD.t77 0.092694
R32594 DVDD DVDD.t94 0.092694
R32595 DVDD DVDD.t99 0.092694
R32596 DVDD.n22244 DVDD.n22243 0.0865488
R32597 DVDD.n22241 DVDD.n49 0.0865488
R32598 DVDD.n18730 DVDD.n18671 0.0865488
R32599 DVDD.n21247 DVDD.n21214 0.0865488
R32600 DVDD.n4329 DVDD.n2350 0.0862854
R32601 DVDD.n4262 DVDD.n2391 0.0862854
R32602 DVDD.n3728 DVDD.n3349 0.0862854
R32603 DVDD.n3647 DVDD.n3421 0.0862854
R32604 DVDD.n21479 DVDD.n21371 0.0857632
R32605 DVDD.n19632 DVDD.n19631 0.0857632
R32606 DVDD.n4800 DVDD.n3565 0.0813407
R32607 DVDD.n15716 DVDD.n15715 0.0760366
R32608 DVDD.n2539 DVDD.n530 0.0760366
R32609 DVDD.n5087 DVDD.n5053 0.0760366
R32610 DVDD.n16334 DVDD.n16333 0.0760366
R32611 DVDD.n15425 DVDD.n15424 0.0760366
R32612 DVDD.n16213 DVDD.n16212 0.0760366
R32613 DVDD.n15324 DVDD.n15323 0.0760366
R32614 DVDD.n2895 DVDD.n761 0.0760366
R32615 DVDD.n18162 DVDD.n475 0.0756776
R32616 DVDD.n19426 DVDD.n19425 0.0703684
R32617 DVDD.n19375 DVDD.n18648 0.0644474
R32618 DVDD.n21273 DVDD.n18652 0.0644474
R32619 DVDD.n10158 DVDD.n10157 0.0640746
R32620 DVDD.n10153 DVDD.n10152 0.0640746
R32621 DVDD.n9582 DVDD.n9577 0.0640746
R32622 DVDD.n10142 DVDD.n10141 0.0640746
R32623 DVDD.n10140 DVDD.n10139 0.0640746
R32624 DVDD.n9590 DVDD.n9585 0.0640746
R32625 DVDD.n10129 DVDD.n10128 0.0640746
R32626 DVDD.n10127 DVDD.n10126 0.0640746
R32627 DVDD.n9597 DVDD.n9593 0.0640746
R32628 DVDD.n10117 DVDD.n10116 0.0640746
R32629 DVDD.n10115 DVDD.n10114 0.0640746
R32630 DVDD.n9605 DVDD.n9600 0.0640746
R32631 DVDD.n10104 DVDD.n10103 0.0640746
R32632 DVDD.n10102 DVDD.n10101 0.0640746
R32633 DVDD.n9739 DVDD.n9608 0.0640746
R32634 DVDD.n9953 DVDD.n9687 0.0640746
R32635 DVDD.n9800 DVDD.n9799 0.0640746
R32636 DVDD.n9942 DVDD.n9941 0.0640746
R32637 DVDD.n9788 DVDD.n9787 0.0640746
R32638 DVDD.n9790 DVDD.n9789 0.0640746
R32639 DVDD.n9785 DVDD.n9784 0.0640746
R32640 DVDD.n16062 DVDD.n3032 0.0640746
R32641 DVDD.n16012 DVDD.n16011 0.0640746
R32642 DVDD.n16046 DVDD.n16045 0.0640746
R32643 DVDD.n16024 DVDD.n16023 0.0640746
R32644 DVDD.n16035 DVDD.n16034 0.0640746
R32645 DVDD.n3105 DVDD.n3104 0.0640746
R32646 DVDD.n5163 DVDD.n5162 0.0640746
R32647 DVDD.n5174 DVDD.n5173 0.0640746
R32648 DVDD.n5185 DVDD.n5184 0.0640746
R32649 DVDD.n5196 DVDD.n5195 0.0640746
R32650 DVDD.n15523 DVDD.n15522 0.0640746
R32651 DVDD.n15530 DVDD.n2734 0.0640746
R32652 DVDD.n15539 DVDD.n15538 0.0640746
R32653 DVDD.n15548 DVDD.n15547 0.0640746
R32654 DVDD.n15557 DVDD.n15556 0.0640746
R32655 DVDD.n15566 DVDD.n15565 0.0640746
R32656 DVDD.n15575 DVDD.n15574 0.0640746
R32657 DVDD.n15606 DVDD.n2692 0.0640746
R32658 DVDD.n3435 DVDD.n3434 0.0640746
R32659 DVDD.n3446 DVDD.n3445 0.0640746
R32660 DVDD.n3457 DVDD.n3456 0.0640746
R32661 DVDD.n10165 DVDD.n2282 0.0640746
R32662 DVDD.n10166 DVDD.n8962 0.0640746
R32663 DVDD.n10163 DVDD.n10162 0.0640746
R32664 DVDD.n10161 DVDD.n10160 0.0640746
R32665 DVDD.n10150 DVDD.n9575 0.0640746
R32666 DVDD.n10147 DVDD.n10146 0.0640746
R32667 DVDD.n10145 DVDD.n10144 0.0640746
R32668 DVDD.n10137 DVDD.n9581 0.0640746
R32669 DVDD.n10134 DVDD.n10133 0.0640746
R32670 DVDD.n10132 DVDD.n10131 0.0640746
R32671 DVDD.n10124 DVDD.n9589 0.0640746
R32672 DVDD.n10121 DVDD.n10120 0.0640746
R32673 DVDD.n10119 DVDD.n10118 0.0640746
R32674 DVDD.n10112 DVDD.n9596 0.0640746
R32675 DVDD.n10109 DVDD.n10108 0.0640746
R32676 DVDD.n10107 DVDD.n10106 0.0640746
R32677 DVDD.n10099 DVDD.n9604 0.0640746
R32678 DVDD.n10096 DVDD.n10095 0.0640746
R32679 DVDD.n9951 DVDD.n9612 0.0640746
R32680 DVDD.n9803 DVDD.n9802 0.0640746
R32681 DVDD.n9945 DVDD.n9944 0.0640746
R32682 DVDD.n9794 DVDD.n9793 0.0640746
R32683 DVDD.n9792 DVDD.n9791 0.0640746
R32684 DVDD.n9783 DVDD.n9779 0.0640746
R32685 DVDD.n16064 DVDD.n3081 0.0640746
R32686 DVDD.n16015 DVDD.n16014 0.0640746
R32687 DVDD.n16049 DVDD.n16048 0.0640746
R32688 DVDD.n16027 DVDD.n16026 0.0640746
R32689 DVDD.n16038 DVDD.n16037 0.0640746
R32690 DVDD.n16071 DVDD.n16070 0.0640746
R32691 DVDD.n5166 DVDD.n5165 0.0640746
R32692 DVDD.n5177 DVDD.n5176 0.0640746
R32693 DVDD.n5188 DVDD.n5187 0.0640746
R32694 DVDD.n5198 DVDD.n5197 0.0640746
R32695 DVDD.n15525 DVDD.n15524 0.0640746
R32696 DVDD.n15532 DVDD.n3174 0.0640746
R32697 DVDD.n15542 DVDD.n15541 0.0640746
R32698 DVDD.n15551 DVDD.n15550 0.0640746
R32699 DVDD.n15560 DVDD.n15559 0.0640746
R32700 DVDD.n15569 DVDD.n15568 0.0640746
R32701 DVDD.n15578 DVDD.n15577 0.0640746
R32702 DVDD.n15608 DVDD.n3286 0.0640746
R32703 DVDD.n3438 DVDD.n3437 0.0640746
R32704 DVDD.n3449 DVDD.n3448 0.0640746
R32705 DVDD.n3459 DVDD.n3458 0.0640746
R32706 DVDD.n10156 DVDD.n10155 0.0638464
R32707 DVDD.n21272 DVDD.n18653 0.0628842
R32708 DVDD.n128 DVDD.n11 0.0628842
R32709 DVDD.n21015 DVDD.n21014 0.059934
R32710 DVDD.n21018 DVDD.n21017 0.059934
R32711 DVDD DVDD.n3447 0.059934
R32712 DVDD DVDD.n3436 0.059934
R32713 DVDD DVDD.n15607 0.059934
R32714 DVDD DVDD.n15576 0.059934
R32715 DVDD DVDD.n15567 0.059934
R32716 DVDD DVDD.n15558 0.059934
R32717 DVDD DVDD.n15549 0.059934
R32718 DVDD DVDD.n15540 0.059934
R32719 DVDD DVDD.n15531 0.059934
R32720 DVDD DVDD.n5186 0.059934
R32721 DVDD DVDD.n5175 0.059934
R32722 DVDD DVDD.n5164 0.059934
R32723 DVDD DVDD.n3106 0.059934
R32724 DVDD DVDD.n16036 0.059934
R32725 DVDD DVDD.n16025 0.059934
R32726 DVDD DVDD.n16047 0.059934
R32727 DVDD DVDD.n16013 0.059934
R32728 DVDD DVDD.n16063 0.059934
R32729 DVDD DVDD.n9776 0.059934
R32730 DVDD DVDD.n9943 0.059934
R32731 DVDD DVDD.n9801 0.059934
R32732 DVDD DVDD.n9952 0.059934
R32733 DVDD DVDD.n9611 0.059934
R32734 DVDD DVDD.n10100 0.059934
R32735 DVDD DVDD.n10105 0.059934
R32736 DVDD DVDD.n9603 0.059934
R32737 DVDD DVDD.n10113 0.059934
R32738 DVDD DVDD.n10125 0.059934
R32739 DVDD DVDD.n10130 0.059934
R32740 DVDD DVDD.n9588 0.059934
R32741 DVDD DVDD.n10138 0.059934
R32742 DVDD DVDD.n10143 0.059934
R32743 DVDD DVDD.n9580 0.059934
R32744 DVDD DVDD.n10151 0.059934
R32745 DVDD DVDD.n10159 0.059934
R32746 DVDD DVDD.n9574 0.059934
R32747 DVDD.n21278 DVDD.n18648 0.0597105
R32748 DVDD.n21274 DVDD.n21273 0.0597105
R32749 DVDD.n20526 DVDD.n20521 0.0569562
R32750 DVDD.n20527 DVDD.n20522 0.0569562
R32751 DVDD.n20528 DVDD.n20523 0.0569562
R32752 DVDD.n20484 DVDD.n19798 0.0569562
R32753 DVDD.n19800 DVDD.n19799 0.0569562
R32754 DVDD.n19802 DVDD.n19801 0.0569562
R32755 DVDD.n19804 DVDD.n19803 0.0569562
R32756 DVDD.n19806 DVDD.n19805 0.0569562
R32757 DVDD.n19808 DVDD.n19807 0.0569562
R32758 DVDD.n20478 DVDD.n20477 0.0569562
R32759 DVDD.n20476 DVDD.n20475 0.0569562
R32760 DVDD.n20474 DVDD.n20473 0.0569562
R32761 DVDD.n20472 DVDD.n20471 0.0569562
R32762 DVDD.n20470 DVDD.n20469 0.0569562
R32763 DVDD.n20468 DVDD.n20467 0.0569562
R32764 DVDD.n20965 DVDD.n20964 0.0569562
R32765 DVDD.n20963 DVDD.n20962 0.0569562
R32766 DVDD.n20961 DVDD.n20960 0.0569562
R32767 DVDD.n20959 DVDD.n20958 0.0569562
R32768 DVDD.n20957 DVDD.n20956 0.0569562
R32769 DVDD.n20955 DVDD.n20954 0.0569562
R32770 DVDD.n20953 DVDD.n20952 0.0569562
R32771 DVDD.n20948 DVDD.n20947 0.0569562
R32772 DVDD.n20946 DVDD.n20945 0.0569562
R32773 DVDD.n20944 DVDD.n20943 0.0569562
R32774 DVDD.n20942 DVDD.n20941 0.0569562
R32775 DVDD.n20940 DVDD.n20939 0.0569562
R32776 DVDD.n20938 DVDD.n20937 0.0569562
R32777 DVDD.n20936 DVDD.n20935 0.0569562
R32778 DVDD.n19080 DVDD.n19079 0.0569562
R32779 DVDD.n19082 DVDD.n19081 0.0569562
R32780 DVDD.n19084 DVDD.n19083 0.0569562
R32781 DVDD.n19086 DVDD.n19085 0.0569562
R32782 DVDD.n19088 DVDD.n19087 0.0569562
R32783 DVDD.n19090 DVDD.n19089 0.0569562
R32784 DVDD.n19092 DVDD.n19091 0.0569562
R32785 DVDD.n19120 DVDD.n19119 0.0569562
R32786 DVDD.n19118 DVDD.n19117 0.0569562
R32787 DVDD.n19116 DVDD.n19115 0.0569562
R32788 DVDD.n19114 DVDD.n19113 0.0569562
R32789 DVDD.n19112 DVDD.n19111 0.0569562
R32790 DVDD.n19110 DVDD.n19109 0.0569562
R32791 DVDD.n19108 DVDD.n19107 0.0569562
R32792 DVDD.n20975 DVDD.n18825 0.0569562
R32793 DVDD.n20976 DVDD.n18826 0.0569562
R32794 DVDD.n20977 DVDD.n18827 0.0569562
R32795 DVDD.n18764 DVDD.n18755 0.0569562
R32796 DVDD.n18765 DVDD.n18756 0.0569562
R32797 DVDD.n18766 DVDD.n18757 0.0569562
R32798 DVDD.n18767 DVDD.n18758 0.0569562
R32799 DVDD.n18768 DVDD.n18759 0.0569562
R32800 DVDD.n18769 DVDD.n18760 0.0569562
R32801 DVDD.n18775 DVDD.n18774 0.0569562
R32802 DVDD.n18777 DVDD.n18776 0.0569562
R32803 DVDD.n18779 DVDD.n18778 0.0569562
R32804 DVDD.n18781 DVDD.n18780 0.0569562
R32805 DVDD.n18783 DVDD.n18782 0.0569562
R32806 DVDD.n18785 DVDD.n18784 0.0569562
R32807 DVDD.n18786 DVDD.n18785 0.0569562
R32808 DVDD.n18784 DVDD.n18783 0.0569562
R32809 DVDD.n18782 DVDD.n18781 0.0569562
R32810 DVDD.n18780 DVDD.n18779 0.0569562
R32811 DVDD.n18778 DVDD.n18777 0.0569562
R32812 DVDD.n18776 DVDD.n18775 0.0569562
R32813 DVDD.n19107 DVDD.n19106 0.0569562
R32814 DVDD.n19109 DVDD.n19108 0.0569562
R32815 DVDD.n19111 DVDD.n19110 0.0569562
R32816 DVDD.n19113 DVDD.n19112 0.0569562
R32817 DVDD.n19115 DVDD.n19114 0.0569562
R32818 DVDD.n19117 DVDD.n19116 0.0569562
R32819 DVDD.n19119 DVDD.n19118 0.0569562
R32820 DVDD.n20935 DVDD.n20934 0.0569562
R32821 DVDD.n20937 DVDD.n20936 0.0569562
R32822 DVDD.n20939 DVDD.n20938 0.0569562
R32823 DVDD.n20941 DVDD.n20940 0.0569562
R32824 DVDD.n20943 DVDD.n20942 0.0569562
R32825 DVDD.n20945 DVDD.n20944 0.0569562
R32826 DVDD.n20947 DVDD.n20946 0.0569562
R32827 DVDD.n20467 DVDD.n20466 0.0569562
R32828 DVDD.n20469 DVDD.n20468 0.0569562
R32829 DVDD.n20471 DVDD.n20470 0.0569562
R32830 DVDD.n20473 DVDD.n20472 0.0569562
R32831 DVDD.n20475 DVDD.n20474 0.0569562
R32832 DVDD.n20477 DVDD.n20476 0.0569562
R32833 DVDD.n18769 DVDD.n18761 0.0569562
R32834 DVDD.n18768 DVDD.n18760 0.0569562
R32835 DVDD.n18767 DVDD.n18759 0.0569562
R32836 DVDD.n18766 DVDD.n18758 0.0569562
R32837 DVDD.n18765 DVDD.n18757 0.0569562
R32838 DVDD.n18764 DVDD.n18756 0.0569562
R32839 DVDD.n19093 DVDD.n19092 0.0569562
R32840 DVDD.n19091 DVDD.n19090 0.0569562
R32841 DVDD.n19089 DVDD.n19088 0.0569562
R32842 DVDD.n19087 DVDD.n19086 0.0569562
R32843 DVDD.n19085 DVDD.n19084 0.0569562
R32844 DVDD.n19083 DVDD.n19082 0.0569562
R32845 DVDD.n19081 DVDD.n19080 0.0569562
R32846 DVDD.n20952 DVDD.n20951 0.0569562
R32847 DVDD.n20954 DVDD.n20953 0.0569562
R32848 DVDD.n20956 DVDD.n20955 0.0569562
R32849 DVDD.n20958 DVDD.n20957 0.0569562
R32850 DVDD.n20960 DVDD.n20959 0.0569562
R32851 DVDD.n20962 DVDD.n20961 0.0569562
R32852 DVDD.n20964 DVDD.n20963 0.0569562
R32853 DVDD.n19809 DVDD.n19808 0.0569562
R32854 DVDD.n19807 DVDD.n19806 0.0569562
R32855 DVDD.n19805 DVDD.n19804 0.0569562
R32856 DVDD.n19803 DVDD.n19802 0.0569562
R32857 DVDD.n19801 DVDD.n19800 0.0569562
R32858 DVDD.n19799 DVDD.n19798 0.0569562
R32859 DVDD.n20977 DVDD.n18828 0.0569562
R32860 DVDD.n20976 DVDD.n18827 0.0569562
R32861 DVDD.n20975 DVDD.n18826 0.0569562
R32862 DVDD.n20523 DVDD.n20486 0.0569562
R32863 DVDD.n20528 DVDD.n20522 0.0569562
R32864 DVDD.n20527 DVDD.n20521 0.0569562
R32865 DVDD.n20530 DVDD.n20525 0.0563
R32866 DVDD.n20525 DVDD.n20524 0.0563
R32867 DVDD.n20534 DVDD.n20533 0.0563
R32868 DVDD.n20533 DVDD.n20485 0.0563
R32869 DVDD.n20482 DVDD.n20481 0.0563
R32870 DVDD.n20481 DVDD.n20479 0.0563
R32871 DVDD.n20925 DVDD.n20924 0.0563
R32872 DVDD.n20981 DVDD.n20980 0.0563
R32873 DVDD.n20980 DVDD.n20979 0.0563
R32874 DVDD.n21058 DVDD.n21057 0.0563
R32875 DVDD.n21057 DVDD.n21056 0.0563
R32876 DVDD.n21053 DVDD.n18771 0.0563
R32877 DVDD.n18773 DVDD.n18771 0.0563
R32878 DVDD.n19100 DVDD.n19099 0.0563
R32879 DVDD.n19425 DVDD.n19424 0.0537895
R32880 DVDD.n223 DVDD.n218 0.0521876
R32881 DVDD.n22209 DVDD.n190 0.0515891
R32882 DVDD.n18432 DVDD.n135 0.0515849
R32883 DVDD.n4452 DVDD.n4416 0.0515834
R32884 DVDD.n22209 DVDD.n187 0.0503876
R32885 DVDD.n223 DVDD.n217 0.0497891
R32886 DVDD.n18432 DVDD.n147 0.0497891
R32887 DVDD.n4451 DVDD.n4416 0.0497834
R32888 DVDD.n20462 DVDD.n20441 0.0490122
R32889 DVDD.n20919 DVDD.n20900 0.0490122
R32890 DVDD.n20541 DVDD.n20540 0.0490122
R32891 DVDD.n20516 DVDD.n19764 0.0490122
R32892 DVDD.n16431 DVDD.n2282 0.0485293
R32893 DVDD.n16449 DVDD.n2268 0.0485293
R32894 DVDD.n10219 DVDD.n8962 0.0485293
R32895 DVDD.n10202 DVDD.n10167 0.0485293
R32896 DVDD.n5001 DVDD.n4985 0.0467228
R32897 DVDD.n549 DVDD.n544 0.0467228
R32898 DVDD.n15146 DVDD.n15145 0.0467228
R32899 DVDD.n17736 DVDD.n885 0.0467228
R32900 DVDD.n9789 DVDD.n9785 0.0440512
R32901 DVDD.n10116 DVDD.n9593 0.0440512
R32902 DVDD.n9781 DVDD.n9780 0.0440512
R32903 DVDD.n9599 DVDD.n9598 0.0440512
R32904 DVDD.n9792 DVDD.n9779 0.0440512
R32905 DVDD.n10120 DVDD.n10119 0.0440512
R32906 DVDD.n9782 DVDD.n9775 0.0440512
R32907 DVDD.n10122 DVDD.n9595 0.0440512
R32908 DVDD.n20081 DVDD 0.0410947
R32909 DVDD.n20897 DVDD 0.0410947
R32910 DVDD.n21371 DVDD.n21328 0.0383947
R32911 DVDD.n19632 DVDD.n19215 0.0383947
R32912 DVDD.n19895 DVDD 0.0381244
R32913 DVDD.n20438 DVDD 0.0381244
R32914 DVDD.n19982 DVDD 0.0381244
R32915 DVDD.n20593 DVDD 0.0381244
R32916 DVDD.n1600 DVDD.n1267 0.0380882
R32917 DVDD.n1600 DVDD.n1599 0.0380882
R32918 DVDD.n1599 DVDD.n1598 0.0380882
R32919 DVDD.n1598 DVDD.n1316 0.0380882
R32920 DVDD.n1588 DVDD.n1316 0.0380882
R32921 DVDD.n1588 DVDD.n1587 0.0380882
R32922 DVDD.n1587 DVDD.n1586 0.0380882
R32923 DVDD.n1586 DVDD.n1318 0.0380882
R32924 DVDD.n1576 DVDD.n1318 0.0380882
R32925 DVDD.n1576 DVDD.n1575 0.0380882
R32926 DVDD.n1575 DVDD.n1574 0.0380882
R32927 DVDD.n1574 DVDD.n1320 0.0380882
R32928 DVDD.n1564 DVDD.n1320 0.0380882
R32929 DVDD.n1564 DVDD.n1563 0.0380882
R32930 DVDD.n1563 DVDD.n1562 0.0380882
R32931 DVDD.n1562 DVDD.n1322 0.0380882
R32932 DVDD.n1552 DVDD.n1322 0.0380882
R32933 DVDD.n1552 DVDD.n1551 0.0380882
R32934 DVDD.n1551 DVDD.n1550 0.0380882
R32935 DVDD.n1550 DVDD.n1324 0.0380882
R32936 DVDD.n1540 DVDD.n1324 0.0380882
R32937 DVDD.n1540 DVDD.n1539 0.0380882
R32938 DVDD.n1539 DVDD.n1538 0.0380882
R32939 DVDD.n1538 DVDD.n1326 0.0380882
R32940 DVDD.n1528 DVDD.n1326 0.0380882
R32941 DVDD.n1528 DVDD.n1527 0.0380882
R32942 DVDD.n1527 DVDD.n1526 0.0380882
R32943 DVDD.n1526 DVDD.n1328 0.0380882
R32944 DVDD.n1516 DVDD.n1328 0.0380882
R32945 DVDD.n1516 DVDD.n1515 0.0380882
R32946 DVDD.n1515 DVDD.n1514 0.0380882
R32947 DVDD.n1514 DVDD.n1330 0.0380882
R32948 DVDD.n1504 DVDD.n1330 0.0380882
R32949 DVDD.n1504 DVDD.n1503 0.0380882
R32950 DVDD.n1503 DVDD.n1502 0.0380882
R32951 DVDD.n1502 DVDD.n1332 0.0380882
R32952 DVDD.n1492 DVDD.n1332 0.0380882
R32953 DVDD.n1492 DVDD.n1491 0.0380882
R32954 DVDD.n1491 DVDD.n1490 0.0380882
R32955 DVDD.n1490 DVDD.n1334 0.0380882
R32956 DVDD.n1480 DVDD.n1334 0.0380882
R32957 DVDD.n1480 DVDD.n1479 0.0380882
R32958 DVDD.n1479 DVDD.n1478 0.0380882
R32959 DVDD.n1478 DVDD.n1336 0.0380882
R32960 DVDD.n1468 DVDD.n1336 0.0380882
R32961 DVDD.n1468 DVDD.n1467 0.0380882
R32962 DVDD.n1467 DVDD.n1466 0.0380882
R32963 DVDD.n1466 DVDD.n1338 0.0380882
R32964 DVDD.n1456 DVDD.n1338 0.0380882
R32965 DVDD.n1456 DVDD.n1455 0.0380882
R32966 DVDD.n1455 DVDD.n1454 0.0380882
R32967 DVDD.n1454 DVDD.n1340 0.0380882
R32968 DVDD.n1444 DVDD.n1340 0.0380882
R32969 DVDD.n1444 DVDD.n1443 0.0380882
R32970 DVDD.n1443 DVDD.n1442 0.0380882
R32971 DVDD.n1442 DVDD.n1342 0.0380882
R32972 DVDD.n1432 DVDD.n1342 0.0380882
R32973 DVDD.n1432 DVDD.n1431 0.0380882
R32974 DVDD.n1431 DVDD.n1430 0.0380882
R32975 DVDD.n1430 DVDD.n1344 0.0380882
R32976 DVDD.n1420 DVDD.n1344 0.0380882
R32977 DVDD.n1420 DVDD.n1419 0.0380882
R32978 DVDD.n1419 DVDD.n1418 0.0380882
R32979 DVDD.n1418 DVDD.n1346 0.0380882
R32980 DVDD.n1408 DVDD.n1346 0.0380882
R32981 DVDD.n1408 DVDD.n1407 0.0380882
R32982 DVDD.n1407 DVDD.n1406 0.0380882
R32983 DVDD.n1406 DVDD.n1348 0.0380882
R32984 DVDD.n1396 DVDD.n1348 0.0380882
R32985 DVDD.n1396 DVDD.n1395 0.0380882
R32986 DVDD.n1395 DVDD.n1394 0.0380882
R32987 DVDD.n1394 DVDD.n1350 0.0380882
R32988 DVDD.n1384 DVDD.n1350 0.0380882
R32989 DVDD.n1384 DVDD.n1383 0.0380882
R32990 DVDD.n1383 DVDD.n1382 0.0380882
R32991 DVDD.n1382 DVDD.n1352 0.0380882
R32992 DVDD.n1372 DVDD.n1352 0.0380882
R32993 DVDD.n1372 DVDD.n1371 0.0380882
R32994 DVDD.n1371 DVDD.n1370 0.0380882
R32995 DVDD.n1370 DVDD.n1354 0.0380882
R32996 DVDD.n1360 DVDD.n1354 0.0380882
R32997 DVDD.n1360 DVDD.n1359 0.0380882
R32998 DVDD.n1359 DVDD.n1358 0.0380882
R32999 DVDD.n6860 DVDD.n6858 0.0380882
R33000 DVDD.n6861 DVDD.n6860 0.0380882
R33001 DVDD.n6862 DVDD.n6861 0.0380882
R33002 DVDD.n6862 DVDD.n6855 0.0380882
R33003 DVDD.n6869 DVDD.n6855 0.0380882
R33004 DVDD.n6870 DVDD.n6869 0.0380882
R33005 DVDD.n6871 DVDD.n6870 0.0380882
R33006 DVDD.n6871 DVDD.n6852 0.0380882
R33007 DVDD.n6878 DVDD.n6852 0.0380882
R33008 DVDD.n6879 DVDD.n6878 0.0380882
R33009 DVDD.n6880 DVDD.n6879 0.0380882
R33010 DVDD.n6880 DVDD.n6849 0.0380882
R33011 DVDD.n6887 DVDD.n6849 0.0380882
R33012 DVDD.n6888 DVDD.n6887 0.0380882
R33013 DVDD.n6889 DVDD.n6888 0.0380882
R33014 DVDD.n6889 DVDD.n6846 0.0380882
R33015 DVDD.n6896 DVDD.n6846 0.0380882
R33016 DVDD.n6897 DVDD.n6896 0.0380882
R33017 DVDD.n6898 DVDD.n6897 0.0380882
R33018 DVDD.n6898 DVDD.n6843 0.0380882
R33019 DVDD.n6905 DVDD.n6843 0.0380882
R33020 DVDD.n6906 DVDD.n6905 0.0380882
R33021 DVDD.n6907 DVDD.n6906 0.0380882
R33022 DVDD.n6907 DVDD.n6840 0.0380882
R33023 DVDD.n6914 DVDD.n6840 0.0380882
R33024 DVDD.n6915 DVDD.n6914 0.0380882
R33025 DVDD.n6916 DVDD.n6915 0.0380882
R33026 DVDD.n6916 DVDD.n6837 0.0380882
R33027 DVDD.n6923 DVDD.n6837 0.0380882
R33028 DVDD.n6924 DVDD.n6923 0.0380882
R33029 DVDD.n6925 DVDD.n6924 0.0380882
R33030 DVDD.n6925 DVDD.n6834 0.0380882
R33031 DVDD.n6932 DVDD.n6834 0.0380882
R33032 DVDD.n6933 DVDD.n6932 0.0380882
R33033 DVDD.n6934 DVDD.n6933 0.0380882
R33034 DVDD.n6934 DVDD.n6831 0.0380882
R33035 DVDD.n6941 DVDD.n6831 0.0380882
R33036 DVDD.n6942 DVDD.n6941 0.0380882
R33037 DVDD.n6943 DVDD.n6942 0.0380882
R33038 DVDD.n6943 DVDD.n6828 0.0380882
R33039 DVDD.n6950 DVDD.n6828 0.0380882
R33040 DVDD.n6951 DVDD.n6950 0.0380882
R33041 DVDD.n6952 DVDD.n6951 0.0380882
R33042 DVDD.n6952 DVDD.n6825 0.0380882
R33043 DVDD.n6959 DVDD.n6825 0.0380882
R33044 DVDD.n6960 DVDD.n6959 0.0380882
R33045 DVDD.n6961 DVDD.n6960 0.0380882
R33046 DVDD.n6961 DVDD.n6822 0.0380882
R33047 DVDD.n6968 DVDD.n6822 0.0380882
R33048 DVDD.n6969 DVDD.n6968 0.0380882
R33049 DVDD.n6970 DVDD.n6969 0.0380882
R33050 DVDD.n6970 DVDD.n6819 0.0380882
R33051 DVDD.n6977 DVDD.n6819 0.0380882
R33052 DVDD.n6978 DVDD.n6977 0.0380882
R33053 DVDD.n6979 DVDD.n6978 0.0380882
R33054 DVDD.n6979 DVDD.n6816 0.0380882
R33055 DVDD.n6986 DVDD.n6816 0.0380882
R33056 DVDD.n6987 DVDD.n6986 0.0380882
R33057 DVDD.n6988 DVDD.n6987 0.0380882
R33058 DVDD.n6988 DVDD.n6813 0.0380882
R33059 DVDD.n6995 DVDD.n6813 0.0380882
R33060 DVDD.n6996 DVDD.n6995 0.0380882
R33061 DVDD.n6997 DVDD.n6996 0.0380882
R33062 DVDD.n6997 DVDD.n6810 0.0380882
R33063 DVDD.n7004 DVDD.n6810 0.0380882
R33064 DVDD.n7005 DVDD.n7004 0.0380882
R33065 DVDD.n7006 DVDD.n7005 0.0380882
R33066 DVDD.n7006 DVDD.n6807 0.0380882
R33067 DVDD.n7013 DVDD.n6807 0.0380882
R33068 DVDD.n7014 DVDD.n7013 0.0380882
R33069 DVDD.n7015 DVDD.n7014 0.0380882
R33070 DVDD.n7015 DVDD.n6804 0.0380882
R33071 DVDD.n7022 DVDD.n6804 0.0380882
R33072 DVDD.n7023 DVDD.n7022 0.0380882
R33073 DVDD.n7024 DVDD.n7023 0.0380882
R33074 DVDD.n7024 DVDD.n6801 0.0380882
R33075 DVDD.n7031 DVDD.n6801 0.0380882
R33076 DVDD.n7032 DVDD.n7031 0.0380882
R33077 DVDD.n7033 DVDD.n7032 0.0380882
R33078 DVDD.n7033 DVDD.n6798 0.0380882
R33079 DVDD.n7040 DVDD.n6798 0.0380882
R33080 DVDD.n7041 DVDD.n7040 0.0380882
R33081 DVDD.n7042 DVDD.n7041 0.0380882
R33082 DVDD.n6859 DVDD.n6751 0.0380882
R33083 DVDD.n6859 DVDD.n6857 0.0380882
R33084 DVDD.n6864 DVDD.n6857 0.0380882
R33085 DVDD.n6866 DVDD.n6864 0.0380882
R33086 DVDD.n6868 DVDD.n6866 0.0380882
R33087 DVDD.n6868 DVDD.n6854 0.0380882
R33088 DVDD.n6873 DVDD.n6854 0.0380882
R33089 DVDD.n6875 DVDD.n6873 0.0380882
R33090 DVDD.n6877 DVDD.n6875 0.0380882
R33091 DVDD.n6877 DVDD.n6851 0.0380882
R33092 DVDD.n6882 DVDD.n6851 0.0380882
R33093 DVDD.n6884 DVDD.n6882 0.0380882
R33094 DVDD.n6886 DVDD.n6884 0.0380882
R33095 DVDD.n6886 DVDD.n6848 0.0380882
R33096 DVDD.n6891 DVDD.n6848 0.0380882
R33097 DVDD.n6893 DVDD.n6891 0.0380882
R33098 DVDD.n6895 DVDD.n6893 0.0380882
R33099 DVDD.n6895 DVDD.n6845 0.0380882
R33100 DVDD.n6900 DVDD.n6845 0.0380882
R33101 DVDD.n6902 DVDD.n6900 0.0380882
R33102 DVDD.n6904 DVDD.n6902 0.0380882
R33103 DVDD.n6904 DVDD.n6842 0.0380882
R33104 DVDD.n6909 DVDD.n6842 0.0380882
R33105 DVDD.n6911 DVDD.n6909 0.0380882
R33106 DVDD.n6913 DVDD.n6911 0.0380882
R33107 DVDD.n6913 DVDD.n6839 0.0380882
R33108 DVDD.n6918 DVDD.n6839 0.0380882
R33109 DVDD.n6920 DVDD.n6918 0.0380882
R33110 DVDD.n6922 DVDD.n6920 0.0380882
R33111 DVDD.n6922 DVDD.n6836 0.0380882
R33112 DVDD.n6927 DVDD.n6836 0.0380882
R33113 DVDD.n6929 DVDD.n6927 0.0380882
R33114 DVDD.n6931 DVDD.n6929 0.0380882
R33115 DVDD.n6931 DVDD.n6833 0.0380882
R33116 DVDD.n6936 DVDD.n6833 0.0380882
R33117 DVDD.n6938 DVDD.n6936 0.0380882
R33118 DVDD.n6940 DVDD.n6938 0.0380882
R33119 DVDD.n6940 DVDD.n6830 0.0380882
R33120 DVDD.n6945 DVDD.n6830 0.0380882
R33121 DVDD.n6947 DVDD.n6945 0.0380882
R33122 DVDD.n6949 DVDD.n6947 0.0380882
R33123 DVDD.n6949 DVDD.n6827 0.0380882
R33124 DVDD.n6954 DVDD.n6827 0.0380882
R33125 DVDD.n6956 DVDD.n6954 0.0380882
R33126 DVDD.n6958 DVDD.n6956 0.0380882
R33127 DVDD.n6958 DVDD.n6824 0.0380882
R33128 DVDD.n6963 DVDD.n6824 0.0380882
R33129 DVDD.n6965 DVDD.n6963 0.0380882
R33130 DVDD.n6967 DVDD.n6965 0.0380882
R33131 DVDD.n6967 DVDD.n6821 0.0380882
R33132 DVDD.n6972 DVDD.n6821 0.0380882
R33133 DVDD.n6974 DVDD.n6972 0.0380882
R33134 DVDD.n6976 DVDD.n6974 0.0380882
R33135 DVDD.n6976 DVDD.n6818 0.0380882
R33136 DVDD.n6981 DVDD.n6818 0.0380882
R33137 DVDD.n6983 DVDD.n6981 0.0380882
R33138 DVDD.n6985 DVDD.n6983 0.0380882
R33139 DVDD.n6985 DVDD.n6815 0.0380882
R33140 DVDD.n6990 DVDD.n6815 0.0380882
R33141 DVDD.n6992 DVDD.n6990 0.0380882
R33142 DVDD.n6994 DVDD.n6992 0.0380882
R33143 DVDD.n6994 DVDD.n6812 0.0380882
R33144 DVDD.n6999 DVDD.n6812 0.0380882
R33145 DVDD.n7001 DVDD.n6999 0.0380882
R33146 DVDD.n7003 DVDD.n7001 0.0380882
R33147 DVDD.n7003 DVDD.n6809 0.0380882
R33148 DVDD.n7008 DVDD.n6809 0.0380882
R33149 DVDD.n7010 DVDD.n7008 0.0380882
R33150 DVDD.n7012 DVDD.n7010 0.0380882
R33151 DVDD.n7012 DVDD.n6806 0.0380882
R33152 DVDD.n7017 DVDD.n6806 0.0380882
R33153 DVDD.n7019 DVDD.n7017 0.0380882
R33154 DVDD.n7021 DVDD.n7019 0.0380882
R33155 DVDD.n7021 DVDD.n6803 0.0380882
R33156 DVDD.n7026 DVDD.n6803 0.0380882
R33157 DVDD.n7028 DVDD.n7026 0.0380882
R33158 DVDD.n7030 DVDD.n7028 0.0380882
R33159 DVDD.n7030 DVDD.n6800 0.0380882
R33160 DVDD.n7035 DVDD.n6800 0.0380882
R33161 DVDD.n7037 DVDD.n7035 0.0380882
R33162 DVDD.n7039 DVDD.n7037 0.0380882
R33163 DVDD.n7039 DVDD.n6797 0.0380882
R33164 DVDD.n15087 DVDD.n6797 0.0380882
R33165 DVDD.n7157 DVDD.n7066 0.0380882
R33166 DVDD.n7158 DVDD.n7157 0.0380882
R33167 DVDD.n7158 DVDD.n7152 0.0380882
R33168 DVDD.n7168 DVDD.n7152 0.0380882
R33169 DVDD.n7169 DVDD.n7168 0.0380882
R33170 DVDD.n7170 DVDD.n7169 0.0380882
R33171 DVDD.n7170 DVDD.n7150 0.0380882
R33172 DVDD.n7180 DVDD.n7150 0.0380882
R33173 DVDD.n7181 DVDD.n7180 0.0380882
R33174 DVDD.n7182 DVDD.n7181 0.0380882
R33175 DVDD.n7182 DVDD.n7148 0.0380882
R33176 DVDD.n7192 DVDD.n7148 0.0380882
R33177 DVDD.n7193 DVDD.n7192 0.0380882
R33178 DVDD.n7194 DVDD.n7193 0.0380882
R33179 DVDD.n7194 DVDD.n7146 0.0380882
R33180 DVDD.n7204 DVDD.n7146 0.0380882
R33181 DVDD.n7205 DVDD.n7204 0.0380882
R33182 DVDD.n7206 DVDD.n7205 0.0380882
R33183 DVDD.n7206 DVDD.n7144 0.0380882
R33184 DVDD.n7216 DVDD.n7144 0.0380882
R33185 DVDD.n7217 DVDD.n7216 0.0380882
R33186 DVDD.n7218 DVDD.n7217 0.0380882
R33187 DVDD.n7218 DVDD.n7142 0.0380882
R33188 DVDD.n7228 DVDD.n7142 0.0380882
R33189 DVDD.n7229 DVDD.n7228 0.0380882
R33190 DVDD.n7230 DVDD.n7229 0.0380882
R33191 DVDD.n7230 DVDD.n7140 0.0380882
R33192 DVDD.n7240 DVDD.n7140 0.0380882
R33193 DVDD.n7241 DVDD.n7240 0.0380882
R33194 DVDD.n7242 DVDD.n7241 0.0380882
R33195 DVDD.n7242 DVDD.n7138 0.0380882
R33196 DVDD.n7252 DVDD.n7138 0.0380882
R33197 DVDD.n7253 DVDD.n7252 0.0380882
R33198 DVDD.n7254 DVDD.n7253 0.0380882
R33199 DVDD.n7254 DVDD.n7136 0.0380882
R33200 DVDD.n7264 DVDD.n7136 0.0380882
R33201 DVDD.n7265 DVDD.n7264 0.0380882
R33202 DVDD.n7266 DVDD.n7265 0.0380882
R33203 DVDD.n7266 DVDD.n7134 0.0380882
R33204 DVDD.n7276 DVDD.n7134 0.0380882
R33205 DVDD.n7277 DVDD.n7276 0.0380882
R33206 DVDD.n7278 DVDD.n7277 0.0380882
R33207 DVDD.n7278 DVDD.n7132 0.0380882
R33208 DVDD.n7288 DVDD.n7132 0.0380882
R33209 DVDD.n7289 DVDD.n7288 0.0380882
R33210 DVDD.n7290 DVDD.n7289 0.0380882
R33211 DVDD.n7290 DVDD.n7130 0.0380882
R33212 DVDD.n7300 DVDD.n7130 0.0380882
R33213 DVDD.n7301 DVDD.n7300 0.0380882
R33214 DVDD.n7302 DVDD.n7301 0.0380882
R33215 DVDD.n7302 DVDD.n7128 0.0380882
R33216 DVDD.n7312 DVDD.n7128 0.0380882
R33217 DVDD.n7313 DVDD.n7312 0.0380882
R33218 DVDD.n7314 DVDD.n7313 0.0380882
R33219 DVDD.n7314 DVDD.n7126 0.0380882
R33220 DVDD.n7324 DVDD.n7126 0.0380882
R33221 DVDD.n7325 DVDD.n7324 0.0380882
R33222 DVDD.n7326 DVDD.n7325 0.0380882
R33223 DVDD.n7326 DVDD.n7124 0.0380882
R33224 DVDD.n7336 DVDD.n7124 0.0380882
R33225 DVDD.n7337 DVDD.n7336 0.0380882
R33226 DVDD.n7338 DVDD.n7337 0.0380882
R33227 DVDD.n7338 DVDD.n7122 0.0380882
R33228 DVDD.n7348 DVDD.n7122 0.0380882
R33229 DVDD.n7349 DVDD.n7348 0.0380882
R33230 DVDD.n7350 DVDD.n7349 0.0380882
R33231 DVDD.n7350 DVDD.n7120 0.0380882
R33232 DVDD.n7360 DVDD.n7120 0.0380882
R33233 DVDD.n7361 DVDD.n7360 0.0380882
R33234 DVDD.n7362 DVDD.n7361 0.0380882
R33235 DVDD.n7362 DVDD.n7118 0.0380882
R33236 DVDD.n7372 DVDD.n7118 0.0380882
R33237 DVDD.n7373 DVDD.n7372 0.0380882
R33238 DVDD.n7374 DVDD.n7373 0.0380882
R33239 DVDD.n7374 DVDD.n7116 0.0380882
R33240 DVDD.n7384 DVDD.n7116 0.0380882
R33241 DVDD.n7385 DVDD.n7384 0.0380882
R33242 DVDD.n7386 DVDD.n7385 0.0380882
R33243 DVDD.n7386 DVDD.n7114 0.0380882
R33244 DVDD.n7396 DVDD.n7114 0.0380882
R33245 DVDD.n7397 DVDD.n7396 0.0380882
R33246 DVDD.n7399 DVDD.n7397 0.0380882
R33247 DVDD.n7399 DVDD.n7398 0.0380882
R33248 DVDD.n7156 DVDD.n7153 0.0380882
R33249 DVDD.n7159 DVDD.n7156 0.0380882
R33250 DVDD.n7163 DVDD.n7159 0.0380882
R33251 DVDD.n7167 DVDD.n7163 0.0380882
R33252 DVDD.n7167 DVDD.n7151 0.0380882
R33253 DVDD.n7171 DVDD.n7151 0.0380882
R33254 DVDD.n7175 DVDD.n7171 0.0380882
R33255 DVDD.n7179 DVDD.n7175 0.0380882
R33256 DVDD.n7179 DVDD.n7149 0.0380882
R33257 DVDD.n7183 DVDD.n7149 0.0380882
R33258 DVDD.n7187 DVDD.n7183 0.0380882
R33259 DVDD.n7191 DVDD.n7187 0.0380882
R33260 DVDD.n7191 DVDD.n7147 0.0380882
R33261 DVDD.n7195 DVDD.n7147 0.0380882
R33262 DVDD.n7199 DVDD.n7195 0.0380882
R33263 DVDD.n7203 DVDD.n7199 0.0380882
R33264 DVDD.n7203 DVDD.n7145 0.0380882
R33265 DVDD.n7207 DVDD.n7145 0.0380882
R33266 DVDD.n7211 DVDD.n7207 0.0380882
R33267 DVDD.n7215 DVDD.n7211 0.0380882
R33268 DVDD.n7215 DVDD.n7143 0.0380882
R33269 DVDD.n7219 DVDD.n7143 0.0380882
R33270 DVDD.n7223 DVDD.n7219 0.0380882
R33271 DVDD.n7227 DVDD.n7223 0.0380882
R33272 DVDD.n7227 DVDD.n7141 0.0380882
R33273 DVDD.n7231 DVDD.n7141 0.0380882
R33274 DVDD.n7235 DVDD.n7231 0.0380882
R33275 DVDD.n7239 DVDD.n7235 0.0380882
R33276 DVDD.n7239 DVDD.n7139 0.0380882
R33277 DVDD.n7243 DVDD.n7139 0.0380882
R33278 DVDD.n7247 DVDD.n7243 0.0380882
R33279 DVDD.n7251 DVDD.n7247 0.0380882
R33280 DVDD.n7251 DVDD.n7137 0.0380882
R33281 DVDD.n7255 DVDD.n7137 0.0380882
R33282 DVDD.n7259 DVDD.n7255 0.0380882
R33283 DVDD.n7263 DVDD.n7259 0.0380882
R33284 DVDD.n7263 DVDD.n7135 0.0380882
R33285 DVDD.n7267 DVDD.n7135 0.0380882
R33286 DVDD.n7271 DVDD.n7267 0.0380882
R33287 DVDD.n7275 DVDD.n7271 0.0380882
R33288 DVDD.n7275 DVDD.n7133 0.0380882
R33289 DVDD.n7279 DVDD.n7133 0.0380882
R33290 DVDD.n7283 DVDD.n7279 0.0380882
R33291 DVDD.n7287 DVDD.n7283 0.0380882
R33292 DVDD.n7287 DVDD.n7131 0.0380882
R33293 DVDD.n7291 DVDD.n7131 0.0380882
R33294 DVDD.n7295 DVDD.n7291 0.0380882
R33295 DVDD.n7299 DVDD.n7295 0.0380882
R33296 DVDD.n7299 DVDD.n7129 0.0380882
R33297 DVDD.n7303 DVDD.n7129 0.0380882
R33298 DVDD.n7307 DVDD.n7303 0.0380882
R33299 DVDD.n7311 DVDD.n7307 0.0380882
R33300 DVDD.n7311 DVDD.n7127 0.0380882
R33301 DVDD.n7315 DVDD.n7127 0.0380882
R33302 DVDD.n7319 DVDD.n7315 0.0380882
R33303 DVDD.n7323 DVDD.n7319 0.0380882
R33304 DVDD.n7323 DVDD.n7125 0.0380882
R33305 DVDD.n7327 DVDD.n7125 0.0380882
R33306 DVDD.n7331 DVDD.n7327 0.0380882
R33307 DVDD.n7335 DVDD.n7331 0.0380882
R33308 DVDD.n7335 DVDD.n7123 0.0380882
R33309 DVDD.n7339 DVDD.n7123 0.0380882
R33310 DVDD.n7343 DVDD.n7339 0.0380882
R33311 DVDD.n7347 DVDD.n7343 0.0380882
R33312 DVDD.n7347 DVDD.n7121 0.0380882
R33313 DVDD.n7351 DVDD.n7121 0.0380882
R33314 DVDD.n7355 DVDD.n7351 0.0380882
R33315 DVDD.n7359 DVDD.n7355 0.0380882
R33316 DVDD.n7359 DVDD.n7119 0.0380882
R33317 DVDD.n7363 DVDD.n7119 0.0380882
R33318 DVDD.n7367 DVDD.n7363 0.0380882
R33319 DVDD.n7371 DVDD.n7367 0.0380882
R33320 DVDD.n7371 DVDD.n7117 0.0380882
R33321 DVDD.n7375 DVDD.n7117 0.0380882
R33322 DVDD.n7379 DVDD.n7375 0.0380882
R33323 DVDD.n7383 DVDD.n7379 0.0380882
R33324 DVDD.n7383 DVDD.n7115 0.0380882
R33325 DVDD.n7387 DVDD.n7115 0.0380882
R33326 DVDD.n7391 DVDD.n7387 0.0380882
R33327 DVDD.n7395 DVDD.n7391 0.0380882
R33328 DVDD.n7395 DVDD.n7113 0.0380882
R33329 DVDD.n7400 DVDD.n7113 0.0380882
R33330 DVDD.n7400 DVDD.n7112 0.0380882
R33331 DVDD.n14872 DVDD.n14870 0.0380882
R33332 DVDD.n14873 DVDD.n14872 0.0380882
R33333 DVDD.n14874 DVDD.n14873 0.0380882
R33334 DVDD.n14874 DVDD.n7560 0.0380882
R33335 DVDD.n14881 DVDD.n7560 0.0380882
R33336 DVDD.n14882 DVDD.n14881 0.0380882
R33337 DVDD.n14883 DVDD.n14882 0.0380882
R33338 DVDD.n14883 DVDD.n7557 0.0380882
R33339 DVDD.n14890 DVDD.n7557 0.0380882
R33340 DVDD.n14891 DVDD.n14890 0.0380882
R33341 DVDD.n14892 DVDD.n14891 0.0380882
R33342 DVDD.n14892 DVDD.n7554 0.0380882
R33343 DVDD.n14899 DVDD.n7554 0.0380882
R33344 DVDD.n14900 DVDD.n14899 0.0380882
R33345 DVDD.n14901 DVDD.n14900 0.0380882
R33346 DVDD.n14901 DVDD.n7551 0.0380882
R33347 DVDD.n14908 DVDD.n7551 0.0380882
R33348 DVDD.n14909 DVDD.n14908 0.0380882
R33349 DVDD.n14910 DVDD.n14909 0.0380882
R33350 DVDD.n14910 DVDD.n7548 0.0380882
R33351 DVDD.n14917 DVDD.n7548 0.0380882
R33352 DVDD.n14918 DVDD.n14917 0.0380882
R33353 DVDD.n14919 DVDD.n14918 0.0380882
R33354 DVDD.n14919 DVDD.n7545 0.0380882
R33355 DVDD.n14926 DVDD.n7545 0.0380882
R33356 DVDD.n14927 DVDD.n14926 0.0380882
R33357 DVDD.n14928 DVDD.n14927 0.0380882
R33358 DVDD.n14928 DVDD.n7542 0.0380882
R33359 DVDD.n14935 DVDD.n7542 0.0380882
R33360 DVDD.n14936 DVDD.n14935 0.0380882
R33361 DVDD.n14937 DVDD.n14936 0.0380882
R33362 DVDD.n14937 DVDD.n7539 0.0380882
R33363 DVDD.n14944 DVDD.n7539 0.0380882
R33364 DVDD.n14945 DVDD.n14944 0.0380882
R33365 DVDD.n14946 DVDD.n14945 0.0380882
R33366 DVDD.n14946 DVDD.n7536 0.0380882
R33367 DVDD.n14953 DVDD.n7536 0.0380882
R33368 DVDD.n14954 DVDD.n14953 0.0380882
R33369 DVDD.n14955 DVDD.n14954 0.0380882
R33370 DVDD.n14955 DVDD.n7533 0.0380882
R33371 DVDD.n14962 DVDD.n7533 0.0380882
R33372 DVDD.n14963 DVDD.n14962 0.0380882
R33373 DVDD.n14964 DVDD.n14963 0.0380882
R33374 DVDD.n14964 DVDD.n7530 0.0380882
R33375 DVDD.n14971 DVDD.n7530 0.0380882
R33376 DVDD.n14972 DVDD.n14971 0.0380882
R33377 DVDD.n14973 DVDD.n14972 0.0380882
R33378 DVDD.n14973 DVDD.n7527 0.0380882
R33379 DVDD.n14980 DVDD.n7527 0.0380882
R33380 DVDD.n14981 DVDD.n14980 0.0380882
R33381 DVDD.n14982 DVDD.n14981 0.0380882
R33382 DVDD.n14982 DVDD.n7524 0.0380882
R33383 DVDD.n14989 DVDD.n7524 0.0380882
R33384 DVDD.n14990 DVDD.n14989 0.0380882
R33385 DVDD.n14991 DVDD.n14990 0.0380882
R33386 DVDD.n14991 DVDD.n7521 0.0380882
R33387 DVDD.n14998 DVDD.n7521 0.0380882
R33388 DVDD.n14999 DVDD.n14998 0.0380882
R33389 DVDD.n15000 DVDD.n14999 0.0380882
R33390 DVDD.n15000 DVDD.n7518 0.0380882
R33391 DVDD.n15007 DVDD.n7518 0.0380882
R33392 DVDD.n15008 DVDD.n15007 0.0380882
R33393 DVDD.n15009 DVDD.n15008 0.0380882
R33394 DVDD.n15009 DVDD.n7515 0.0380882
R33395 DVDD.n15016 DVDD.n7515 0.0380882
R33396 DVDD.n15017 DVDD.n15016 0.0380882
R33397 DVDD.n15018 DVDD.n15017 0.0380882
R33398 DVDD.n15018 DVDD.n7512 0.0380882
R33399 DVDD.n15025 DVDD.n7512 0.0380882
R33400 DVDD.n15026 DVDD.n15025 0.0380882
R33401 DVDD.n15027 DVDD.n15026 0.0380882
R33402 DVDD.n15027 DVDD.n7509 0.0380882
R33403 DVDD.n15034 DVDD.n7509 0.0380882
R33404 DVDD.n15035 DVDD.n15034 0.0380882
R33405 DVDD.n15036 DVDD.n15035 0.0380882
R33406 DVDD.n15036 DVDD.n7506 0.0380882
R33407 DVDD.n15043 DVDD.n7506 0.0380882
R33408 DVDD.n15044 DVDD.n15043 0.0380882
R33409 DVDD.n15045 DVDD.n15044 0.0380882
R33410 DVDD.n15045 DVDD.n7503 0.0380882
R33411 DVDD.n15052 DVDD.n7503 0.0380882
R33412 DVDD.n15053 DVDD.n15052 0.0380882
R33413 DVDD.n15054 DVDD.n15053 0.0380882
R33414 DVDD.n14871 DVDD.n7457 0.0380882
R33415 DVDD.n14871 DVDD.n7562 0.0380882
R33416 DVDD.n14876 DVDD.n7562 0.0380882
R33417 DVDD.n14878 DVDD.n14876 0.0380882
R33418 DVDD.n14880 DVDD.n14878 0.0380882
R33419 DVDD.n14880 DVDD.n7559 0.0380882
R33420 DVDD.n14885 DVDD.n7559 0.0380882
R33421 DVDD.n14887 DVDD.n14885 0.0380882
R33422 DVDD.n14889 DVDD.n14887 0.0380882
R33423 DVDD.n14889 DVDD.n7556 0.0380882
R33424 DVDD.n14894 DVDD.n7556 0.0380882
R33425 DVDD.n14896 DVDD.n14894 0.0380882
R33426 DVDD.n14898 DVDD.n14896 0.0380882
R33427 DVDD.n14898 DVDD.n7553 0.0380882
R33428 DVDD.n14903 DVDD.n7553 0.0380882
R33429 DVDD.n14905 DVDD.n14903 0.0380882
R33430 DVDD.n14907 DVDD.n14905 0.0380882
R33431 DVDD.n14907 DVDD.n7550 0.0380882
R33432 DVDD.n14912 DVDD.n7550 0.0380882
R33433 DVDD.n14914 DVDD.n14912 0.0380882
R33434 DVDD.n14916 DVDD.n14914 0.0380882
R33435 DVDD.n14916 DVDD.n7547 0.0380882
R33436 DVDD.n14921 DVDD.n7547 0.0380882
R33437 DVDD.n14923 DVDD.n14921 0.0380882
R33438 DVDD.n14925 DVDD.n14923 0.0380882
R33439 DVDD.n14925 DVDD.n7544 0.0380882
R33440 DVDD.n14930 DVDD.n7544 0.0380882
R33441 DVDD.n14932 DVDD.n14930 0.0380882
R33442 DVDD.n14934 DVDD.n14932 0.0380882
R33443 DVDD.n14934 DVDD.n7541 0.0380882
R33444 DVDD.n14939 DVDD.n7541 0.0380882
R33445 DVDD.n14941 DVDD.n14939 0.0380882
R33446 DVDD.n14943 DVDD.n14941 0.0380882
R33447 DVDD.n14943 DVDD.n7538 0.0380882
R33448 DVDD.n14948 DVDD.n7538 0.0380882
R33449 DVDD.n14950 DVDD.n14948 0.0380882
R33450 DVDD.n14952 DVDD.n14950 0.0380882
R33451 DVDD.n14952 DVDD.n7535 0.0380882
R33452 DVDD.n14957 DVDD.n7535 0.0380882
R33453 DVDD.n14959 DVDD.n14957 0.0380882
R33454 DVDD.n14961 DVDD.n14959 0.0380882
R33455 DVDD.n14961 DVDD.n7532 0.0380882
R33456 DVDD.n14966 DVDD.n7532 0.0380882
R33457 DVDD.n14968 DVDD.n14966 0.0380882
R33458 DVDD.n14970 DVDD.n14968 0.0380882
R33459 DVDD.n14970 DVDD.n7529 0.0380882
R33460 DVDD.n14975 DVDD.n7529 0.0380882
R33461 DVDD.n14977 DVDD.n14975 0.0380882
R33462 DVDD.n14979 DVDD.n14977 0.0380882
R33463 DVDD.n14979 DVDD.n7526 0.0380882
R33464 DVDD.n14984 DVDD.n7526 0.0380882
R33465 DVDD.n14986 DVDD.n14984 0.0380882
R33466 DVDD.n14988 DVDD.n14986 0.0380882
R33467 DVDD.n14988 DVDD.n7523 0.0380882
R33468 DVDD.n14993 DVDD.n7523 0.0380882
R33469 DVDD.n14995 DVDD.n14993 0.0380882
R33470 DVDD.n14997 DVDD.n14995 0.0380882
R33471 DVDD.n14997 DVDD.n7520 0.0380882
R33472 DVDD.n15002 DVDD.n7520 0.0380882
R33473 DVDD.n15004 DVDD.n15002 0.0380882
R33474 DVDD.n15006 DVDD.n15004 0.0380882
R33475 DVDD.n15006 DVDD.n7517 0.0380882
R33476 DVDD.n15011 DVDD.n7517 0.0380882
R33477 DVDD.n15013 DVDD.n15011 0.0380882
R33478 DVDD.n15015 DVDD.n15013 0.0380882
R33479 DVDD.n15015 DVDD.n7514 0.0380882
R33480 DVDD.n15020 DVDD.n7514 0.0380882
R33481 DVDD.n15022 DVDD.n15020 0.0380882
R33482 DVDD.n15024 DVDD.n15022 0.0380882
R33483 DVDD.n15024 DVDD.n7511 0.0380882
R33484 DVDD.n15029 DVDD.n7511 0.0380882
R33485 DVDD.n15031 DVDD.n15029 0.0380882
R33486 DVDD.n15033 DVDD.n15031 0.0380882
R33487 DVDD.n15033 DVDD.n7508 0.0380882
R33488 DVDD.n15038 DVDD.n7508 0.0380882
R33489 DVDD.n15040 DVDD.n15038 0.0380882
R33490 DVDD.n15042 DVDD.n15040 0.0380882
R33491 DVDD.n15042 DVDD.n7505 0.0380882
R33492 DVDD.n15047 DVDD.n7505 0.0380882
R33493 DVDD.n15049 DVDD.n15047 0.0380882
R33494 DVDD.n15051 DVDD.n15049 0.0380882
R33495 DVDD.n15051 DVDD.n7502 0.0380882
R33496 DVDD.n15055 DVDD.n7502 0.0380882
R33497 DVDD.n9218 DVDD.n9217 0.0380882
R33498 DVDD.n9217 DVDD.n8975 0.0380882
R33499 DVDD.n9211 DVDD.n8975 0.0380882
R33500 DVDD.n9211 DVDD.n9210 0.0380882
R33501 DVDD.n9210 DVDD.n9209 0.0380882
R33502 DVDD.n9209 DVDD.n8978 0.0380882
R33503 DVDD.n9202 DVDD.n8978 0.0380882
R33504 DVDD.n9202 DVDD.n9201 0.0380882
R33505 DVDD.n9201 DVDD.n9200 0.0380882
R33506 DVDD.n9200 DVDD.n8981 0.0380882
R33507 DVDD.n9193 DVDD.n8981 0.0380882
R33508 DVDD.n9193 DVDD.n9192 0.0380882
R33509 DVDD.n9192 DVDD.n9191 0.0380882
R33510 DVDD.n9191 DVDD.n8984 0.0380882
R33511 DVDD.n9184 DVDD.n8984 0.0380882
R33512 DVDD.n9184 DVDD.n9183 0.0380882
R33513 DVDD.n9183 DVDD.n9182 0.0380882
R33514 DVDD.n9182 DVDD.n8987 0.0380882
R33515 DVDD.n9175 DVDD.n8987 0.0380882
R33516 DVDD.n9175 DVDD.n9174 0.0380882
R33517 DVDD.n9174 DVDD.n9173 0.0380882
R33518 DVDD.n9173 DVDD.n8990 0.0380882
R33519 DVDD.n9166 DVDD.n8990 0.0380882
R33520 DVDD.n9166 DVDD.n9165 0.0380882
R33521 DVDD.n9165 DVDD.n9164 0.0380882
R33522 DVDD.n9164 DVDD.n8993 0.0380882
R33523 DVDD.n9157 DVDD.n8993 0.0380882
R33524 DVDD.n9157 DVDD.n9156 0.0380882
R33525 DVDD.n9156 DVDD.n9155 0.0380882
R33526 DVDD.n9155 DVDD.n8996 0.0380882
R33527 DVDD.n9148 DVDD.n8996 0.0380882
R33528 DVDD.n9148 DVDD.n9147 0.0380882
R33529 DVDD.n9147 DVDD.n9146 0.0380882
R33530 DVDD.n9146 DVDD.n8999 0.0380882
R33531 DVDD.n9139 DVDD.n8999 0.0380882
R33532 DVDD.n9139 DVDD.n9138 0.0380882
R33533 DVDD.n9138 DVDD.n9137 0.0380882
R33534 DVDD.n9137 DVDD.n9002 0.0380882
R33535 DVDD.n9130 DVDD.n9002 0.0380882
R33536 DVDD.n9130 DVDD.n9129 0.0380882
R33537 DVDD.n9129 DVDD.n9128 0.0380882
R33538 DVDD.n9128 DVDD.n9005 0.0380882
R33539 DVDD.n9121 DVDD.n9005 0.0380882
R33540 DVDD.n9121 DVDD.n9120 0.0380882
R33541 DVDD.n9120 DVDD.n9119 0.0380882
R33542 DVDD.n9119 DVDD.n9008 0.0380882
R33543 DVDD.n9112 DVDD.n9008 0.0380882
R33544 DVDD.n9112 DVDD.n9111 0.0380882
R33545 DVDD.n9111 DVDD.n9110 0.0380882
R33546 DVDD.n9110 DVDD.n9011 0.0380882
R33547 DVDD.n9103 DVDD.n9011 0.0380882
R33548 DVDD.n9103 DVDD.n9102 0.0380882
R33549 DVDD.n9102 DVDD.n9101 0.0380882
R33550 DVDD.n9101 DVDD.n9014 0.0380882
R33551 DVDD.n9094 DVDD.n9014 0.0380882
R33552 DVDD.n9094 DVDD.n9093 0.0380882
R33553 DVDD.n9093 DVDD.n9092 0.0380882
R33554 DVDD.n9092 DVDD.n9017 0.0380882
R33555 DVDD.n9085 DVDD.n9017 0.0380882
R33556 DVDD.n9085 DVDD.n9084 0.0380882
R33557 DVDD.n9084 DVDD.n9083 0.0380882
R33558 DVDD.n9083 DVDD.n9020 0.0380882
R33559 DVDD.n9076 DVDD.n9020 0.0380882
R33560 DVDD.n9076 DVDD.n9075 0.0380882
R33561 DVDD.n9075 DVDD.n9074 0.0380882
R33562 DVDD.n9074 DVDD.n9023 0.0380882
R33563 DVDD.n9067 DVDD.n9023 0.0380882
R33564 DVDD.n9067 DVDD.n9066 0.0380882
R33565 DVDD.n9066 DVDD.n9065 0.0380882
R33566 DVDD.n9065 DVDD.n9026 0.0380882
R33567 DVDD.n9058 DVDD.n9026 0.0380882
R33568 DVDD.n9058 DVDD.n9057 0.0380882
R33569 DVDD.n9057 DVDD.n9056 0.0380882
R33570 DVDD.n9056 DVDD.n9029 0.0380882
R33571 DVDD.n9049 DVDD.n9029 0.0380882
R33572 DVDD.n9049 DVDD.n9048 0.0380882
R33573 DVDD.n9048 DVDD.n9047 0.0380882
R33574 DVDD.n9047 DVDD.n9032 0.0380882
R33575 DVDD.n9040 DVDD.n9032 0.0380882
R33576 DVDD.n9040 DVDD.n9039 0.0380882
R33577 DVDD.n9039 DVDD.n9038 0.0380882
R33578 DVDD.n9038 DVDD.n9035 0.0380882
R33579 DVDD.n9035 DVDD.n7661 0.0380882
R33580 DVDD.n9216 DVDD.n7614 0.0380882
R33581 DVDD.n9216 DVDD.n9215 0.0380882
R33582 DVDD.n9215 DVDD.n9213 0.0380882
R33583 DVDD.n9213 DVDD.n8977 0.0380882
R33584 DVDD.n9208 DVDD.n8977 0.0380882
R33585 DVDD.n9208 DVDD.n9206 0.0380882
R33586 DVDD.n9206 DVDD.n9204 0.0380882
R33587 DVDD.n9204 DVDD.n8980 0.0380882
R33588 DVDD.n9199 DVDD.n8980 0.0380882
R33589 DVDD.n9199 DVDD.n9197 0.0380882
R33590 DVDD.n9197 DVDD.n9195 0.0380882
R33591 DVDD.n9195 DVDD.n8983 0.0380882
R33592 DVDD.n9190 DVDD.n8983 0.0380882
R33593 DVDD.n9190 DVDD.n9188 0.0380882
R33594 DVDD.n9188 DVDD.n9186 0.0380882
R33595 DVDD.n9186 DVDD.n8986 0.0380882
R33596 DVDD.n9181 DVDD.n8986 0.0380882
R33597 DVDD.n9181 DVDD.n9179 0.0380882
R33598 DVDD.n9179 DVDD.n9177 0.0380882
R33599 DVDD.n9177 DVDD.n8989 0.0380882
R33600 DVDD.n9172 DVDD.n8989 0.0380882
R33601 DVDD.n9172 DVDD.n9170 0.0380882
R33602 DVDD.n9170 DVDD.n9168 0.0380882
R33603 DVDD.n9168 DVDD.n8992 0.0380882
R33604 DVDD.n9163 DVDD.n8992 0.0380882
R33605 DVDD.n9163 DVDD.n9161 0.0380882
R33606 DVDD.n9161 DVDD.n9159 0.0380882
R33607 DVDD.n9159 DVDD.n8995 0.0380882
R33608 DVDD.n9154 DVDD.n8995 0.0380882
R33609 DVDD.n9154 DVDD.n9152 0.0380882
R33610 DVDD.n9152 DVDD.n9150 0.0380882
R33611 DVDD.n9150 DVDD.n8998 0.0380882
R33612 DVDD.n9145 DVDD.n8998 0.0380882
R33613 DVDD.n9145 DVDD.n9143 0.0380882
R33614 DVDD.n9143 DVDD.n9141 0.0380882
R33615 DVDD.n9141 DVDD.n9001 0.0380882
R33616 DVDD.n9136 DVDD.n9001 0.0380882
R33617 DVDD.n9136 DVDD.n9134 0.0380882
R33618 DVDD.n9134 DVDD.n9132 0.0380882
R33619 DVDD.n9132 DVDD.n9004 0.0380882
R33620 DVDD.n9127 DVDD.n9004 0.0380882
R33621 DVDD.n9127 DVDD.n9125 0.0380882
R33622 DVDD.n9125 DVDD.n9123 0.0380882
R33623 DVDD.n9123 DVDD.n9007 0.0380882
R33624 DVDD.n9118 DVDD.n9007 0.0380882
R33625 DVDD.n9118 DVDD.n9116 0.0380882
R33626 DVDD.n9116 DVDD.n9114 0.0380882
R33627 DVDD.n9114 DVDD.n9010 0.0380882
R33628 DVDD.n9109 DVDD.n9010 0.0380882
R33629 DVDD.n9109 DVDD.n9107 0.0380882
R33630 DVDD.n9107 DVDD.n9105 0.0380882
R33631 DVDD.n9105 DVDD.n9013 0.0380882
R33632 DVDD.n9100 DVDD.n9013 0.0380882
R33633 DVDD.n9100 DVDD.n9098 0.0380882
R33634 DVDD.n9098 DVDD.n9096 0.0380882
R33635 DVDD.n9096 DVDD.n9016 0.0380882
R33636 DVDD.n9091 DVDD.n9016 0.0380882
R33637 DVDD.n9091 DVDD.n9089 0.0380882
R33638 DVDD.n9089 DVDD.n9087 0.0380882
R33639 DVDD.n9087 DVDD.n9019 0.0380882
R33640 DVDD.n9082 DVDD.n9019 0.0380882
R33641 DVDD.n9082 DVDD.n9080 0.0380882
R33642 DVDD.n9080 DVDD.n9078 0.0380882
R33643 DVDD.n9078 DVDD.n9022 0.0380882
R33644 DVDD.n9073 DVDD.n9022 0.0380882
R33645 DVDD.n9073 DVDD.n9071 0.0380882
R33646 DVDD.n9071 DVDD.n9069 0.0380882
R33647 DVDD.n9069 DVDD.n9025 0.0380882
R33648 DVDD.n9064 DVDD.n9025 0.0380882
R33649 DVDD.n9064 DVDD.n9062 0.0380882
R33650 DVDD.n9062 DVDD.n9060 0.0380882
R33651 DVDD.n9060 DVDD.n9028 0.0380882
R33652 DVDD.n9055 DVDD.n9028 0.0380882
R33653 DVDD.n9055 DVDD.n9053 0.0380882
R33654 DVDD.n9053 DVDD.n9051 0.0380882
R33655 DVDD.n9051 DVDD.n9031 0.0380882
R33656 DVDD.n9046 DVDD.n9031 0.0380882
R33657 DVDD.n9046 DVDD.n9044 0.0380882
R33658 DVDD.n9044 DVDD.n9042 0.0380882
R33659 DVDD.n9042 DVDD.n9034 0.0380882
R33660 DVDD.n9037 DVDD.n9034 0.0380882
R33661 DVDD.n9037 DVDD.n7660 0.0380882
R33662 DVDD.n14858 DVDD.n7660 0.0380882
R33663 DVDD.n9553 DVDD.n9265 0.0380882
R33664 DVDD.n9553 DVDD.n9552 0.0380882
R33665 DVDD.n9552 DVDD.n9551 0.0380882
R33666 DVDD.n9551 DVDD.n9269 0.0380882
R33667 DVDD.n9541 DVDD.n9269 0.0380882
R33668 DVDD.n9541 DVDD.n9540 0.0380882
R33669 DVDD.n9540 DVDD.n9539 0.0380882
R33670 DVDD.n9539 DVDD.n9271 0.0380882
R33671 DVDD.n9529 DVDD.n9271 0.0380882
R33672 DVDD.n9529 DVDD.n9528 0.0380882
R33673 DVDD.n9528 DVDD.n9527 0.0380882
R33674 DVDD.n9527 DVDD.n9273 0.0380882
R33675 DVDD.n9517 DVDD.n9273 0.0380882
R33676 DVDD.n9517 DVDD.n9516 0.0380882
R33677 DVDD.n9516 DVDD.n9515 0.0380882
R33678 DVDD.n9515 DVDD.n9275 0.0380882
R33679 DVDD.n9505 DVDD.n9275 0.0380882
R33680 DVDD.n9505 DVDD.n9504 0.0380882
R33681 DVDD.n9504 DVDD.n9503 0.0380882
R33682 DVDD.n9503 DVDD.n9277 0.0380882
R33683 DVDD.n9493 DVDD.n9277 0.0380882
R33684 DVDD.n9493 DVDD.n9492 0.0380882
R33685 DVDD.n9492 DVDD.n9491 0.0380882
R33686 DVDD.n9491 DVDD.n9279 0.0380882
R33687 DVDD.n9481 DVDD.n9279 0.0380882
R33688 DVDD.n9481 DVDD.n9480 0.0380882
R33689 DVDD.n9480 DVDD.n9479 0.0380882
R33690 DVDD.n9479 DVDD.n9281 0.0380882
R33691 DVDD.n9469 DVDD.n9281 0.0380882
R33692 DVDD.n9469 DVDD.n9468 0.0380882
R33693 DVDD.n9468 DVDD.n9467 0.0380882
R33694 DVDD.n9467 DVDD.n9283 0.0380882
R33695 DVDD.n9457 DVDD.n9283 0.0380882
R33696 DVDD.n9457 DVDD.n9456 0.0380882
R33697 DVDD.n9456 DVDD.n9455 0.0380882
R33698 DVDD.n9455 DVDD.n9285 0.0380882
R33699 DVDD.n9445 DVDD.n9285 0.0380882
R33700 DVDD.n9445 DVDD.n9444 0.0380882
R33701 DVDD.n9444 DVDD.n9443 0.0380882
R33702 DVDD.n9443 DVDD.n9287 0.0380882
R33703 DVDD.n9433 DVDD.n9287 0.0380882
R33704 DVDD.n9433 DVDD.n9432 0.0380882
R33705 DVDD.n9432 DVDD.n9431 0.0380882
R33706 DVDD.n9431 DVDD.n9289 0.0380882
R33707 DVDD.n9421 DVDD.n9289 0.0380882
R33708 DVDD.n9421 DVDD.n9420 0.0380882
R33709 DVDD.n9420 DVDD.n9419 0.0380882
R33710 DVDD.n9419 DVDD.n9291 0.0380882
R33711 DVDD.n9409 DVDD.n9291 0.0380882
R33712 DVDD.n9409 DVDD.n9408 0.0380882
R33713 DVDD.n9408 DVDD.n9407 0.0380882
R33714 DVDD.n9407 DVDD.n9293 0.0380882
R33715 DVDD.n9397 DVDD.n9293 0.0380882
R33716 DVDD.n9397 DVDD.n9396 0.0380882
R33717 DVDD.n9396 DVDD.n9395 0.0380882
R33718 DVDD.n9395 DVDD.n9295 0.0380882
R33719 DVDD.n9385 DVDD.n9295 0.0380882
R33720 DVDD.n9385 DVDD.n9384 0.0380882
R33721 DVDD.n9384 DVDD.n9383 0.0380882
R33722 DVDD.n9383 DVDD.n9297 0.0380882
R33723 DVDD.n9373 DVDD.n9297 0.0380882
R33724 DVDD.n9373 DVDD.n9372 0.0380882
R33725 DVDD.n9372 DVDD.n9371 0.0380882
R33726 DVDD.n9371 DVDD.n9299 0.0380882
R33727 DVDD.n9361 DVDD.n9299 0.0380882
R33728 DVDD.n9361 DVDD.n9360 0.0380882
R33729 DVDD.n9360 DVDD.n9359 0.0380882
R33730 DVDD.n9359 DVDD.n9301 0.0380882
R33731 DVDD.n9349 DVDD.n9301 0.0380882
R33732 DVDD.n9349 DVDD.n9348 0.0380882
R33733 DVDD.n9348 DVDD.n9347 0.0380882
R33734 DVDD.n9347 DVDD.n9303 0.0380882
R33735 DVDD.n9337 DVDD.n9303 0.0380882
R33736 DVDD.n9337 DVDD.n9336 0.0380882
R33737 DVDD.n9336 DVDD.n9335 0.0380882
R33738 DVDD.n9335 DVDD.n9305 0.0380882
R33739 DVDD.n9325 DVDD.n9305 0.0380882
R33740 DVDD.n9325 DVDD.n9324 0.0380882
R33741 DVDD.n9324 DVDD.n9323 0.0380882
R33742 DVDD.n9323 DVDD.n9307 0.0380882
R33743 DVDD.n9313 DVDD.n9307 0.0380882
R33744 DVDD.n9313 DVDD.n9312 0.0380882
R33745 DVDD.n9312 DVDD.n9311 0.0380882
R33746 DVDD.n9555 DVDD.n9554 0.0380882
R33747 DVDD.n9554 DVDD.n9268 0.0380882
R33748 DVDD.n9550 DVDD.n9268 0.0380882
R33749 DVDD.n9550 DVDD.n9546 0.0380882
R33750 DVDD.n9546 DVDD.n9545 0.0380882
R33751 DVDD.n9545 DVDD.n9270 0.0380882
R33752 DVDD.n9538 DVDD.n9270 0.0380882
R33753 DVDD.n9538 DVDD.n9534 0.0380882
R33754 DVDD.n9534 DVDD.n9533 0.0380882
R33755 DVDD.n9533 DVDD.n9272 0.0380882
R33756 DVDD.n9526 DVDD.n9272 0.0380882
R33757 DVDD.n9526 DVDD.n9522 0.0380882
R33758 DVDD.n9522 DVDD.n9521 0.0380882
R33759 DVDD.n9521 DVDD.n9274 0.0380882
R33760 DVDD.n9514 DVDD.n9274 0.0380882
R33761 DVDD.n9514 DVDD.n9510 0.0380882
R33762 DVDD.n9510 DVDD.n9509 0.0380882
R33763 DVDD.n9509 DVDD.n9276 0.0380882
R33764 DVDD.n9502 DVDD.n9276 0.0380882
R33765 DVDD.n9502 DVDD.n9498 0.0380882
R33766 DVDD.n9498 DVDD.n9497 0.0380882
R33767 DVDD.n9497 DVDD.n9278 0.0380882
R33768 DVDD.n9490 DVDD.n9278 0.0380882
R33769 DVDD.n9490 DVDD.n9486 0.0380882
R33770 DVDD.n9486 DVDD.n9485 0.0380882
R33771 DVDD.n9485 DVDD.n9280 0.0380882
R33772 DVDD.n9478 DVDD.n9280 0.0380882
R33773 DVDD.n9478 DVDD.n9474 0.0380882
R33774 DVDD.n9474 DVDD.n9473 0.0380882
R33775 DVDD.n9473 DVDD.n9282 0.0380882
R33776 DVDD.n9466 DVDD.n9282 0.0380882
R33777 DVDD.n9466 DVDD.n9462 0.0380882
R33778 DVDD.n9462 DVDD.n9461 0.0380882
R33779 DVDD.n9461 DVDD.n9284 0.0380882
R33780 DVDD.n9454 DVDD.n9284 0.0380882
R33781 DVDD.n9454 DVDD.n9450 0.0380882
R33782 DVDD.n9450 DVDD.n9449 0.0380882
R33783 DVDD.n9449 DVDD.n9286 0.0380882
R33784 DVDD.n9442 DVDD.n9286 0.0380882
R33785 DVDD.n9442 DVDD.n9438 0.0380882
R33786 DVDD.n9438 DVDD.n9437 0.0380882
R33787 DVDD.n9437 DVDD.n9288 0.0380882
R33788 DVDD.n9430 DVDD.n9288 0.0380882
R33789 DVDD.n9430 DVDD.n9426 0.0380882
R33790 DVDD.n9426 DVDD.n9425 0.0380882
R33791 DVDD.n9425 DVDD.n9290 0.0380882
R33792 DVDD.n9418 DVDD.n9290 0.0380882
R33793 DVDD.n9418 DVDD.n9414 0.0380882
R33794 DVDD.n9414 DVDD.n9413 0.0380882
R33795 DVDD.n9413 DVDD.n9292 0.0380882
R33796 DVDD.n9406 DVDD.n9292 0.0380882
R33797 DVDD.n9406 DVDD.n9402 0.0380882
R33798 DVDD.n9402 DVDD.n9401 0.0380882
R33799 DVDD.n9401 DVDD.n9294 0.0380882
R33800 DVDD.n9394 DVDD.n9294 0.0380882
R33801 DVDD.n9394 DVDD.n9390 0.0380882
R33802 DVDD.n9390 DVDD.n9389 0.0380882
R33803 DVDD.n9389 DVDD.n9296 0.0380882
R33804 DVDD.n9382 DVDD.n9296 0.0380882
R33805 DVDD.n9382 DVDD.n9378 0.0380882
R33806 DVDD.n9378 DVDD.n9377 0.0380882
R33807 DVDD.n9377 DVDD.n9298 0.0380882
R33808 DVDD.n9370 DVDD.n9298 0.0380882
R33809 DVDD.n9370 DVDD.n9366 0.0380882
R33810 DVDD.n9366 DVDD.n9365 0.0380882
R33811 DVDD.n9365 DVDD.n9300 0.0380882
R33812 DVDD.n9358 DVDD.n9300 0.0380882
R33813 DVDD.n9358 DVDD.n9354 0.0380882
R33814 DVDD.n9354 DVDD.n9353 0.0380882
R33815 DVDD.n9353 DVDD.n9302 0.0380882
R33816 DVDD.n9346 DVDD.n9302 0.0380882
R33817 DVDD.n9346 DVDD.n9342 0.0380882
R33818 DVDD.n9342 DVDD.n9341 0.0380882
R33819 DVDD.n9341 DVDD.n9304 0.0380882
R33820 DVDD.n9334 DVDD.n9304 0.0380882
R33821 DVDD.n9334 DVDD.n9330 0.0380882
R33822 DVDD.n9330 DVDD.n9329 0.0380882
R33823 DVDD.n9329 DVDD.n9306 0.0380882
R33824 DVDD.n9322 DVDD.n9306 0.0380882
R33825 DVDD.n9322 DVDD.n9318 0.0380882
R33826 DVDD.n9318 DVDD.n9317 0.0380882
R33827 DVDD.n9317 DVDD.n9308 0.0380882
R33828 DVDD.n9310 DVDD.n9308 0.0380882
R33829 DVDD.n7841 DVDD.n7839 0.0380882
R33830 DVDD.n7842 DVDD.n7841 0.0380882
R33831 DVDD.n7843 DVDD.n7842 0.0380882
R33832 DVDD.n7843 DVDD.n7836 0.0380882
R33833 DVDD.n7850 DVDD.n7836 0.0380882
R33834 DVDD.n7851 DVDD.n7850 0.0380882
R33835 DVDD.n7852 DVDD.n7851 0.0380882
R33836 DVDD.n7852 DVDD.n7833 0.0380882
R33837 DVDD.n7859 DVDD.n7833 0.0380882
R33838 DVDD.n7860 DVDD.n7859 0.0380882
R33839 DVDD.n7861 DVDD.n7860 0.0380882
R33840 DVDD.n7861 DVDD.n7830 0.0380882
R33841 DVDD.n7868 DVDD.n7830 0.0380882
R33842 DVDD.n7869 DVDD.n7868 0.0380882
R33843 DVDD.n7870 DVDD.n7869 0.0380882
R33844 DVDD.n7870 DVDD.n7827 0.0380882
R33845 DVDD.n7877 DVDD.n7827 0.0380882
R33846 DVDD.n7878 DVDD.n7877 0.0380882
R33847 DVDD.n7879 DVDD.n7878 0.0380882
R33848 DVDD.n7879 DVDD.n7824 0.0380882
R33849 DVDD.n7886 DVDD.n7824 0.0380882
R33850 DVDD.n7887 DVDD.n7886 0.0380882
R33851 DVDD.n7888 DVDD.n7887 0.0380882
R33852 DVDD.n7888 DVDD.n7821 0.0380882
R33853 DVDD.n7895 DVDD.n7821 0.0380882
R33854 DVDD.n7896 DVDD.n7895 0.0380882
R33855 DVDD.n7897 DVDD.n7896 0.0380882
R33856 DVDD.n7897 DVDD.n7818 0.0380882
R33857 DVDD.n7904 DVDD.n7818 0.0380882
R33858 DVDD.n7905 DVDD.n7904 0.0380882
R33859 DVDD.n7906 DVDD.n7905 0.0380882
R33860 DVDD.n7906 DVDD.n7815 0.0380882
R33861 DVDD.n7913 DVDD.n7815 0.0380882
R33862 DVDD.n7914 DVDD.n7913 0.0380882
R33863 DVDD.n7915 DVDD.n7914 0.0380882
R33864 DVDD.n7915 DVDD.n7812 0.0380882
R33865 DVDD.n7922 DVDD.n7812 0.0380882
R33866 DVDD.n7923 DVDD.n7922 0.0380882
R33867 DVDD.n7924 DVDD.n7923 0.0380882
R33868 DVDD.n7924 DVDD.n7809 0.0380882
R33869 DVDD.n7931 DVDD.n7809 0.0380882
R33870 DVDD.n7932 DVDD.n7931 0.0380882
R33871 DVDD.n7933 DVDD.n7932 0.0380882
R33872 DVDD.n7933 DVDD.n7806 0.0380882
R33873 DVDD.n7940 DVDD.n7806 0.0380882
R33874 DVDD.n7941 DVDD.n7940 0.0380882
R33875 DVDD.n7942 DVDD.n7941 0.0380882
R33876 DVDD.n7942 DVDD.n7803 0.0380882
R33877 DVDD.n7949 DVDD.n7803 0.0380882
R33878 DVDD.n7950 DVDD.n7949 0.0380882
R33879 DVDD.n7951 DVDD.n7950 0.0380882
R33880 DVDD.n7951 DVDD.n7800 0.0380882
R33881 DVDD.n7958 DVDD.n7800 0.0380882
R33882 DVDD.n7959 DVDD.n7958 0.0380882
R33883 DVDD.n7960 DVDD.n7959 0.0380882
R33884 DVDD.n7960 DVDD.n7797 0.0380882
R33885 DVDD.n7967 DVDD.n7797 0.0380882
R33886 DVDD.n7968 DVDD.n7967 0.0380882
R33887 DVDD.n7969 DVDD.n7968 0.0380882
R33888 DVDD.n7969 DVDD.n7794 0.0380882
R33889 DVDD.n7976 DVDD.n7794 0.0380882
R33890 DVDD.n7977 DVDD.n7976 0.0380882
R33891 DVDD.n7978 DVDD.n7977 0.0380882
R33892 DVDD.n7978 DVDD.n7791 0.0380882
R33893 DVDD.n7985 DVDD.n7791 0.0380882
R33894 DVDD.n7986 DVDD.n7985 0.0380882
R33895 DVDD.n7987 DVDD.n7986 0.0380882
R33896 DVDD.n7987 DVDD.n7788 0.0380882
R33897 DVDD.n7994 DVDD.n7788 0.0380882
R33898 DVDD.n7995 DVDD.n7994 0.0380882
R33899 DVDD.n7996 DVDD.n7995 0.0380882
R33900 DVDD.n7996 DVDD.n7785 0.0380882
R33901 DVDD.n8003 DVDD.n7785 0.0380882
R33902 DVDD.n8004 DVDD.n8003 0.0380882
R33903 DVDD.n8005 DVDD.n8004 0.0380882
R33904 DVDD.n8005 DVDD.n7782 0.0380882
R33905 DVDD.n8012 DVDD.n7782 0.0380882
R33906 DVDD.n8013 DVDD.n8012 0.0380882
R33907 DVDD.n8014 DVDD.n8013 0.0380882
R33908 DVDD.n8014 DVDD.n7779 0.0380882
R33909 DVDD.n8021 DVDD.n7779 0.0380882
R33910 DVDD.n8022 DVDD.n8021 0.0380882
R33911 DVDD.n8023 DVDD.n8022 0.0380882
R33912 DVDD.n7840 DVDD.n7732 0.0380882
R33913 DVDD.n7840 DVDD.n7838 0.0380882
R33914 DVDD.n7845 DVDD.n7838 0.0380882
R33915 DVDD.n7847 DVDD.n7845 0.0380882
R33916 DVDD.n7849 DVDD.n7847 0.0380882
R33917 DVDD.n7849 DVDD.n7835 0.0380882
R33918 DVDD.n7854 DVDD.n7835 0.0380882
R33919 DVDD.n7856 DVDD.n7854 0.0380882
R33920 DVDD.n7858 DVDD.n7856 0.0380882
R33921 DVDD.n7858 DVDD.n7832 0.0380882
R33922 DVDD.n7863 DVDD.n7832 0.0380882
R33923 DVDD.n7865 DVDD.n7863 0.0380882
R33924 DVDD.n7867 DVDD.n7865 0.0380882
R33925 DVDD.n7867 DVDD.n7829 0.0380882
R33926 DVDD.n7872 DVDD.n7829 0.0380882
R33927 DVDD.n7874 DVDD.n7872 0.0380882
R33928 DVDD.n7876 DVDD.n7874 0.0380882
R33929 DVDD.n7876 DVDD.n7826 0.0380882
R33930 DVDD.n7881 DVDD.n7826 0.0380882
R33931 DVDD.n7883 DVDD.n7881 0.0380882
R33932 DVDD.n7885 DVDD.n7883 0.0380882
R33933 DVDD.n7885 DVDD.n7823 0.0380882
R33934 DVDD.n7890 DVDD.n7823 0.0380882
R33935 DVDD.n7892 DVDD.n7890 0.0380882
R33936 DVDD.n7894 DVDD.n7892 0.0380882
R33937 DVDD.n7894 DVDD.n7820 0.0380882
R33938 DVDD.n7899 DVDD.n7820 0.0380882
R33939 DVDD.n7901 DVDD.n7899 0.0380882
R33940 DVDD.n7903 DVDD.n7901 0.0380882
R33941 DVDD.n7903 DVDD.n7817 0.0380882
R33942 DVDD.n7908 DVDD.n7817 0.0380882
R33943 DVDD.n7910 DVDD.n7908 0.0380882
R33944 DVDD.n7912 DVDD.n7910 0.0380882
R33945 DVDD.n7912 DVDD.n7814 0.0380882
R33946 DVDD.n7917 DVDD.n7814 0.0380882
R33947 DVDD.n7919 DVDD.n7917 0.0380882
R33948 DVDD.n7921 DVDD.n7919 0.0380882
R33949 DVDD.n7921 DVDD.n7811 0.0380882
R33950 DVDD.n7926 DVDD.n7811 0.0380882
R33951 DVDD.n7928 DVDD.n7926 0.0380882
R33952 DVDD.n7930 DVDD.n7928 0.0380882
R33953 DVDD.n7930 DVDD.n7808 0.0380882
R33954 DVDD.n7935 DVDD.n7808 0.0380882
R33955 DVDD.n7937 DVDD.n7935 0.0380882
R33956 DVDD.n7939 DVDD.n7937 0.0380882
R33957 DVDD.n7939 DVDD.n7805 0.0380882
R33958 DVDD.n7944 DVDD.n7805 0.0380882
R33959 DVDD.n7946 DVDD.n7944 0.0380882
R33960 DVDD.n7948 DVDD.n7946 0.0380882
R33961 DVDD.n7948 DVDD.n7802 0.0380882
R33962 DVDD.n7953 DVDD.n7802 0.0380882
R33963 DVDD.n7955 DVDD.n7953 0.0380882
R33964 DVDD.n7957 DVDD.n7955 0.0380882
R33965 DVDD.n7957 DVDD.n7799 0.0380882
R33966 DVDD.n7962 DVDD.n7799 0.0380882
R33967 DVDD.n7964 DVDD.n7962 0.0380882
R33968 DVDD.n7966 DVDD.n7964 0.0380882
R33969 DVDD.n7966 DVDD.n7796 0.0380882
R33970 DVDD.n7971 DVDD.n7796 0.0380882
R33971 DVDD.n7973 DVDD.n7971 0.0380882
R33972 DVDD.n7975 DVDD.n7973 0.0380882
R33973 DVDD.n7975 DVDD.n7793 0.0380882
R33974 DVDD.n7980 DVDD.n7793 0.0380882
R33975 DVDD.n7982 DVDD.n7980 0.0380882
R33976 DVDD.n7984 DVDD.n7982 0.0380882
R33977 DVDD.n7984 DVDD.n7790 0.0380882
R33978 DVDD.n7989 DVDD.n7790 0.0380882
R33979 DVDD.n7991 DVDD.n7989 0.0380882
R33980 DVDD.n7993 DVDD.n7991 0.0380882
R33981 DVDD.n7993 DVDD.n7787 0.0380882
R33982 DVDD.n7998 DVDD.n7787 0.0380882
R33983 DVDD.n8000 DVDD.n7998 0.0380882
R33984 DVDD.n8002 DVDD.n8000 0.0380882
R33985 DVDD.n8002 DVDD.n7784 0.0380882
R33986 DVDD.n8007 DVDD.n7784 0.0380882
R33987 DVDD.n8009 DVDD.n8007 0.0380882
R33988 DVDD.n8011 DVDD.n8009 0.0380882
R33989 DVDD.n8011 DVDD.n7781 0.0380882
R33990 DVDD.n8016 DVDD.n7781 0.0380882
R33991 DVDD.n8018 DVDD.n8016 0.0380882
R33992 DVDD.n8020 DVDD.n8018 0.0380882
R33993 DVDD.n8020 DVDD.n7778 0.0380882
R33994 DVDD.n14835 DVDD.n7778 0.0380882
R33995 DVDD.n14579 DVDD.n14578 0.0380882
R33996 DVDD.n14580 DVDD.n14579 0.0380882
R33997 DVDD.n14580 DVDD.n8129 0.0380882
R33998 DVDD.n14590 DVDD.n8129 0.0380882
R33999 DVDD.n14591 DVDD.n14590 0.0380882
R34000 DVDD.n14592 DVDD.n14591 0.0380882
R34001 DVDD.n14592 DVDD.n8127 0.0380882
R34002 DVDD.n14602 DVDD.n8127 0.0380882
R34003 DVDD.n14603 DVDD.n14602 0.0380882
R34004 DVDD.n14604 DVDD.n14603 0.0380882
R34005 DVDD.n14604 DVDD.n8125 0.0380882
R34006 DVDD.n14614 DVDD.n8125 0.0380882
R34007 DVDD.n14615 DVDD.n14614 0.0380882
R34008 DVDD.n14616 DVDD.n14615 0.0380882
R34009 DVDD.n14616 DVDD.n8123 0.0380882
R34010 DVDD.n14626 DVDD.n8123 0.0380882
R34011 DVDD.n14627 DVDD.n14626 0.0380882
R34012 DVDD.n14628 DVDD.n14627 0.0380882
R34013 DVDD.n14628 DVDD.n8121 0.0380882
R34014 DVDD.n14638 DVDD.n8121 0.0380882
R34015 DVDD.n14639 DVDD.n14638 0.0380882
R34016 DVDD.n14640 DVDD.n14639 0.0380882
R34017 DVDD.n14640 DVDD.n8119 0.0380882
R34018 DVDD.n14650 DVDD.n8119 0.0380882
R34019 DVDD.n14651 DVDD.n14650 0.0380882
R34020 DVDD.n14652 DVDD.n14651 0.0380882
R34021 DVDD.n14652 DVDD.n8117 0.0380882
R34022 DVDD.n14662 DVDD.n8117 0.0380882
R34023 DVDD.n14663 DVDD.n14662 0.0380882
R34024 DVDD.n14664 DVDD.n14663 0.0380882
R34025 DVDD.n14664 DVDD.n8115 0.0380882
R34026 DVDD.n14674 DVDD.n8115 0.0380882
R34027 DVDD.n14675 DVDD.n14674 0.0380882
R34028 DVDD.n14676 DVDD.n14675 0.0380882
R34029 DVDD.n14676 DVDD.n8113 0.0380882
R34030 DVDD.n14686 DVDD.n8113 0.0380882
R34031 DVDD.n14687 DVDD.n14686 0.0380882
R34032 DVDD.n14688 DVDD.n14687 0.0380882
R34033 DVDD.n14688 DVDD.n8111 0.0380882
R34034 DVDD.n14698 DVDD.n8111 0.0380882
R34035 DVDD.n14699 DVDD.n14698 0.0380882
R34036 DVDD.n14700 DVDD.n14699 0.0380882
R34037 DVDD.n14700 DVDD.n8109 0.0380882
R34038 DVDD.n14710 DVDD.n8109 0.0380882
R34039 DVDD.n14711 DVDD.n14710 0.0380882
R34040 DVDD.n14712 DVDD.n14711 0.0380882
R34041 DVDD.n14712 DVDD.n8107 0.0380882
R34042 DVDD.n14722 DVDD.n8107 0.0380882
R34043 DVDD.n14723 DVDD.n14722 0.0380882
R34044 DVDD.n14724 DVDD.n14723 0.0380882
R34045 DVDD.n14724 DVDD.n8105 0.0380882
R34046 DVDD.n14734 DVDD.n8105 0.0380882
R34047 DVDD.n14735 DVDD.n14734 0.0380882
R34048 DVDD.n14736 DVDD.n14735 0.0380882
R34049 DVDD.n14736 DVDD.n8103 0.0380882
R34050 DVDD.n14746 DVDD.n8103 0.0380882
R34051 DVDD.n14747 DVDD.n14746 0.0380882
R34052 DVDD.n14748 DVDD.n14747 0.0380882
R34053 DVDD.n14748 DVDD.n8101 0.0380882
R34054 DVDD.n14758 DVDD.n8101 0.0380882
R34055 DVDD.n14759 DVDD.n14758 0.0380882
R34056 DVDD.n14760 DVDD.n14759 0.0380882
R34057 DVDD.n14760 DVDD.n8099 0.0380882
R34058 DVDD.n14770 DVDD.n8099 0.0380882
R34059 DVDD.n14771 DVDD.n14770 0.0380882
R34060 DVDD.n14772 DVDD.n14771 0.0380882
R34061 DVDD.n14772 DVDD.n8097 0.0380882
R34062 DVDD.n14782 DVDD.n8097 0.0380882
R34063 DVDD.n14783 DVDD.n14782 0.0380882
R34064 DVDD.n14784 DVDD.n14783 0.0380882
R34065 DVDD.n14784 DVDD.n8095 0.0380882
R34066 DVDD.n14794 DVDD.n8095 0.0380882
R34067 DVDD.n14795 DVDD.n14794 0.0380882
R34068 DVDD.n14796 DVDD.n14795 0.0380882
R34069 DVDD.n14796 DVDD.n8093 0.0380882
R34070 DVDD.n14806 DVDD.n8093 0.0380882
R34071 DVDD.n14807 DVDD.n14806 0.0380882
R34072 DVDD.n14808 DVDD.n14807 0.0380882
R34073 DVDD.n14808 DVDD.n8091 0.0380882
R34074 DVDD.n14818 DVDD.n8091 0.0380882
R34075 DVDD.n14819 DVDD.n14818 0.0380882
R34076 DVDD.n14820 DVDD.n14819 0.0380882
R34077 DVDD.n14820 DVDD.n8038 0.0380882
R34078 DVDD.n14577 DVDD.n8132 0.0380882
R34079 DVDD.n14581 DVDD.n8132 0.0380882
R34080 DVDD.n14585 DVDD.n14581 0.0380882
R34081 DVDD.n14589 DVDD.n14585 0.0380882
R34082 DVDD.n14589 DVDD.n8128 0.0380882
R34083 DVDD.n14593 DVDD.n8128 0.0380882
R34084 DVDD.n14597 DVDD.n14593 0.0380882
R34085 DVDD.n14601 DVDD.n14597 0.0380882
R34086 DVDD.n14601 DVDD.n8126 0.0380882
R34087 DVDD.n14605 DVDD.n8126 0.0380882
R34088 DVDD.n14609 DVDD.n14605 0.0380882
R34089 DVDD.n14613 DVDD.n14609 0.0380882
R34090 DVDD.n14613 DVDD.n8124 0.0380882
R34091 DVDD.n14617 DVDD.n8124 0.0380882
R34092 DVDD.n14621 DVDD.n14617 0.0380882
R34093 DVDD.n14625 DVDD.n14621 0.0380882
R34094 DVDD.n14625 DVDD.n8122 0.0380882
R34095 DVDD.n14629 DVDD.n8122 0.0380882
R34096 DVDD.n14633 DVDD.n14629 0.0380882
R34097 DVDD.n14637 DVDD.n14633 0.0380882
R34098 DVDD.n14637 DVDD.n8120 0.0380882
R34099 DVDD.n14641 DVDD.n8120 0.0380882
R34100 DVDD.n14645 DVDD.n14641 0.0380882
R34101 DVDD.n14649 DVDD.n14645 0.0380882
R34102 DVDD.n14649 DVDD.n8118 0.0380882
R34103 DVDD.n14653 DVDD.n8118 0.0380882
R34104 DVDD.n14657 DVDD.n14653 0.0380882
R34105 DVDD.n14661 DVDD.n14657 0.0380882
R34106 DVDD.n14661 DVDD.n8116 0.0380882
R34107 DVDD.n14665 DVDD.n8116 0.0380882
R34108 DVDD.n14669 DVDD.n14665 0.0380882
R34109 DVDD.n14673 DVDD.n14669 0.0380882
R34110 DVDD.n14673 DVDD.n8114 0.0380882
R34111 DVDD.n14677 DVDD.n8114 0.0380882
R34112 DVDD.n14681 DVDD.n14677 0.0380882
R34113 DVDD.n14685 DVDD.n14681 0.0380882
R34114 DVDD.n14685 DVDD.n8112 0.0380882
R34115 DVDD.n14689 DVDD.n8112 0.0380882
R34116 DVDD.n14693 DVDD.n14689 0.0380882
R34117 DVDD.n14697 DVDD.n14693 0.0380882
R34118 DVDD.n14697 DVDD.n8110 0.0380882
R34119 DVDD.n14701 DVDD.n8110 0.0380882
R34120 DVDD.n14705 DVDD.n14701 0.0380882
R34121 DVDD.n14709 DVDD.n14705 0.0380882
R34122 DVDD.n14709 DVDD.n8108 0.0380882
R34123 DVDD.n14713 DVDD.n8108 0.0380882
R34124 DVDD.n14717 DVDD.n14713 0.0380882
R34125 DVDD.n14721 DVDD.n14717 0.0380882
R34126 DVDD.n14721 DVDD.n8106 0.0380882
R34127 DVDD.n14725 DVDD.n8106 0.0380882
R34128 DVDD.n14729 DVDD.n14725 0.0380882
R34129 DVDD.n14733 DVDD.n14729 0.0380882
R34130 DVDD.n14733 DVDD.n8104 0.0380882
R34131 DVDD.n14737 DVDD.n8104 0.0380882
R34132 DVDD.n14741 DVDD.n14737 0.0380882
R34133 DVDD.n14745 DVDD.n14741 0.0380882
R34134 DVDD.n14745 DVDD.n8102 0.0380882
R34135 DVDD.n14749 DVDD.n8102 0.0380882
R34136 DVDD.n14753 DVDD.n14749 0.0380882
R34137 DVDD.n14757 DVDD.n14753 0.0380882
R34138 DVDD.n14757 DVDD.n8100 0.0380882
R34139 DVDD.n14761 DVDD.n8100 0.0380882
R34140 DVDD.n14765 DVDD.n14761 0.0380882
R34141 DVDD.n14769 DVDD.n14765 0.0380882
R34142 DVDD.n14769 DVDD.n8098 0.0380882
R34143 DVDD.n14773 DVDD.n8098 0.0380882
R34144 DVDD.n14777 DVDD.n14773 0.0380882
R34145 DVDD.n14781 DVDD.n14777 0.0380882
R34146 DVDD.n14781 DVDD.n8096 0.0380882
R34147 DVDD.n14785 DVDD.n8096 0.0380882
R34148 DVDD.n14789 DVDD.n14785 0.0380882
R34149 DVDD.n14793 DVDD.n14789 0.0380882
R34150 DVDD.n14793 DVDD.n8094 0.0380882
R34151 DVDD.n14797 DVDD.n8094 0.0380882
R34152 DVDD.n14801 DVDD.n14797 0.0380882
R34153 DVDD.n14805 DVDD.n14801 0.0380882
R34154 DVDD.n14805 DVDD.n8092 0.0380882
R34155 DVDD.n14809 DVDD.n8092 0.0380882
R34156 DVDD.n14813 DVDD.n14809 0.0380882
R34157 DVDD.n14817 DVDD.n14813 0.0380882
R34158 DVDD.n14817 DVDD.n8090 0.0380882
R34159 DVDD.n14821 DVDD.n8090 0.0380882
R34160 DVDD.n14821 DVDD.n8088 0.0380882
R34161 DVDD.n14313 DVDD.n14312 0.0380882
R34162 DVDD.n14314 DVDD.n14313 0.0380882
R34163 DVDD.n14314 DVDD.n8246 0.0380882
R34164 DVDD.n14324 DVDD.n8246 0.0380882
R34165 DVDD.n14325 DVDD.n14324 0.0380882
R34166 DVDD.n14326 DVDD.n14325 0.0380882
R34167 DVDD.n14326 DVDD.n8244 0.0380882
R34168 DVDD.n14336 DVDD.n8244 0.0380882
R34169 DVDD.n14337 DVDD.n14336 0.0380882
R34170 DVDD.n14338 DVDD.n14337 0.0380882
R34171 DVDD.n14338 DVDD.n8242 0.0380882
R34172 DVDD.n14348 DVDD.n8242 0.0380882
R34173 DVDD.n14349 DVDD.n14348 0.0380882
R34174 DVDD.n14350 DVDD.n14349 0.0380882
R34175 DVDD.n14350 DVDD.n8240 0.0380882
R34176 DVDD.n14360 DVDD.n8240 0.0380882
R34177 DVDD.n14361 DVDD.n14360 0.0380882
R34178 DVDD.n14362 DVDD.n14361 0.0380882
R34179 DVDD.n14362 DVDD.n8238 0.0380882
R34180 DVDD.n14372 DVDD.n8238 0.0380882
R34181 DVDD.n14373 DVDD.n14372 0.0380882
R34182 DVDD.n14374 DVDD.n14373 0.0380882
R34183 DVDD.n14374 DVDD.n8236 0.0380882
R34184 DVDD.n14384 DVDD.n8236 0.0380882
R34185 DVDD.n14385 DVDD.n14384 0.0380882
R34186 DVDD.n14386 DVDD.n14385 0.0380882
R34187 DVDD.n14386 DVDD.n8234 0.0380882
R34188 DVDD.n14396 DVDD.n8234 0.0380882
R34189 DVDD.n14397 DVDD.n14396 0.0380882
R34190 DVDD.n14398 DVDD.n14397 0.0380882
R34191 DVDD.n14398 DVDD.n8232 0.0380882
R34192 DVDD.n14408 DVDD.n8232 0.0380882
R34193 DVDD.n14409 DVDD.n14408 0.0380882
R34194 DVDD.n14410 DVDD.n14409 0.0380882
R34195 DVDD.n14410 DVDD.n8230 0.0380882
R34196 DVDD.n14420 DVDD.n8230 0.0380882
R34197 DVDD.n14421 DVDD.n14420 0.0380882
R34198 DVDD.n14422 DVDD.n14421 0.0380882
R34199 DVDD.n14422 DVDD.n8228 0.0380882
R34200 DVDD.n14432 DVDD.n8228 0.0380882
R34201 DVDD.n14433 DVDD.n14432 0.0380882
R34202 DVDD.n14434 DVDD.n14433 0.0380882
R34203 DVDD.n14434 DVDD.n8226 0.0380882
R34204 DVDD.n14444 DVDD.n8226 0.0380882
R34205 DVDD.n14445 DVDD.n14444 0.0380882
R34206 DVDD.n14446 DVDD.n14445 0.0380882
R34207 DVDD.n14446 DVDD.n8224 0.0380882
R34208 DVDD.n14456 DVDD.n8224 0.0380882
R34209 DVDD.n14457 DVDD.n14456 0.0380882
R34210 DVDD.n14458 DVDD.n14457 0.0380882
R34211 DVDD.n14458 DVDD.n8222 0.0380882
R34212 DVDD.n14468 DVDD.n8222 0.0380882
R34213 DVDD.n14469 DVDD.n14468 0.0380882
R34214 DVDD.n14470 DVDD.n14469 0.0380882
R34215 DVDD.n14470 DVDD.n8220 0.0380882
R34216 DVDD.n14480 DVDD.n8220 0.0380882
R34217 DVDD.n14481 DVDD.n14480 0.0380882
R34218 DVDD.n14482 DVDD.n14481 0.0380882
R34219 DVDD.n14482 DVDD.n8218 0.0380882
R34220 DVDD.n14492 DVDD.n8218 0.0380882
R34221 DVDD.n14493 DVDD.n14492 0.0380882
R34222 DVDD.n14494 DVDD.n14493 0.0380882
R34223 DVDD.n14494 DVDD.n8216 0.0380882
R34224 DVDD.n14504 DVDD.n8216 0.0380882
R34225 DVDD.n14505 DVDD.n14504 0.0380882
R34226 DVDD.n14506 DVDD.n14505 0.0380882
R34227 DVDD.n14506 DVDD.n8214 0.0380882
R34228 DVDD.n14516 DVDD.n8214 0.0380882
R34229 DVDD.n14517 DVDD.n14516 0.0380882
R34230 DVDD.n14518 DVDD.n14517 0.0380882
R34231 DVDD.n14518 DVDD.n8212 0.0380882
R34232 DVDD.n14528 DVDD.n8212 0.0380882
R34233 DVDD.n14529 DVDD.n14528 0.0380882
R34234 DVDD.n14530 DVDD.n14529 0.0380882
R34235 DVDD.n14530 DVDD.n8210 0.0380882
R34236 DVDD.n14540 DVDD.n8210 0.0380882
R34237 DVDD.n14541 DVDD.n14540 0.0380882
R34238 DVDD.n14542 DVDD.n14541 0.0380882
R34239 DVDD.n14542 DVDD.n8208 0.0380882
R34240 DVDD.n14552 DVDD.n8208 0.0380882
R34241 DVDD.n14553 DVDD.n14552 0.0380882
R34242 DVDD.n14554 DVDD.n14553 0.0380882
R34243 DVDD.n14554 DVDD.n8158 0.0380882
R34244 DVDD.n14311 DVDD.n8249 0.0380882
R34245 DVDD.n14315 DVDD.n8249 0.0380882
R34246 DVDD.n14319 DVDD.n14315 0.0380882
R34247 DVDD.n14323 DVDD.n14319 0.0380882
R34248 DVDD.n14323 DVDD.n8245 0.0380882
R34249 DVDD.n14327 DVDD.n8245 0.0380882
R34250 DVDD.n14331 DVDD.n14327 0.0380882
R34251 DVDD.n14335 DVDD.n14331 0.0380882
R34252 DVDD.n14335 DVDD.n8243 0.0380882
R34253 DVDD.n14339 DVDD.n8243 0.0380882
R34254 DVDD.n14343 DVDD.n14339 0.0380882
R34255 DVDD.n14347 DVDD.n14343 0.0380882
R34256 DVDD.n14347 DVDD.n8241 0.0380882
R34257 DVDD.n14351 DVDD.n8241 0.0380882
R34258 DVDD.n14355 DVDD.n14351 0.0380882
R34259 DVDD.n14359 DVDD.n14355 0.0380882
R34260 DVDD.n14359 DVDD.n8239 0.0380882
R34261 DVDD.n14363 DVDD.n8239 0.0380882
R34262 DVDD.n14367 DVDD.n14363 0.0380882
R34263 DVDD.n14371 DVDD.n14367 0.0380882
R34264 DVDD.n14371 DVDD.n8237 0.0380882
R34265 DVDD.n14375 DVDD.n8237 0.0380882
R34266 DVDD.n14379 DVDD.n14375 0.0380882
R34267 DVDD.n14383 DVDD.n14379 0.0380882
R34268 DVDD.n14383 DVDD.n8235 0.0380882
R34269 DVDD.n14387 DVDD.n8235 0.0380882
R34270 DVDD.n14391 DVDD.n14387 0.0380882
R34271 DVDD.n14395 DVDD.n14391 0.0380882
R34272 DVDD.n14395 DVDD.n8233 0.0380882
R34273 DVDD.n14399 DVDD.n8233 0.0380882
R34274 DVDD.n14403 DVDD.n14399 0.0380882
R34275 DVDD.n14407 DVDD.n14403 0.0380882
R34276 DVDD.n14407 DVDD.n8231 0.0380882
R34277 DVDD.n14411 DVDD.n8231 0.0380882
R34278 DVDD.n14415 DVDD.n14411 0.0380882
R34279 DVDD.n14419 DVDD.n14415 0.0380882
R34280 DVDD.n14419 DVDD.n8229 0.0380882
R34281 DVDD.n14423 DVDD.n8229 0.0380882
R34282 DVDD.n14427 DVDD.n14423 0.0380882
R34283 DVDD.n14431 DVDD.n14427 0.0380882
R34284 DVDD.n14431 DVDD.n8227 0.0380882
R34285 DVDD.n14435 DVDD.n8227 0.0380882
R34286 DVDD.n14439 DVDD.n14435 0.0380882
R34287 DVDD.n14443 DVDD.n14439 0.0380882
R34288 DVDD.n14443 DVDD.n8225 0.0380882
R34289 DVDD.n14447 DVDD.n8225 0.0380882
R34290 DVDD.n14451 DVDD.n14447 0.0380882
R34291 DVDD.n14455 DVDD.n14451 0.0380882
R34292 DVDD.n14455 DVDD.n8223 0.0380882
R34293 DVDD.n14459 DVDD.n8223 0.0380882
R34294 DVDD.n14463 DVDD.n14459 0.0380882
R34295 DVDD.n14467 DVDD.n14463 0.0380882
R34296 DVDD.n14467 DVDD.n8221 0.0380882
R34297 DVDD.n14471 DVDD.n8221 0.0380882
R34298 DVDD.n14475 DVDD.n14471 0.0380882
R34299 DVDD.n14479 DVDD.n14475 0.0380882
R34300 DVDD.n14479 DVDD.n8219 0.0380882
R34301 DVDD.n14483 DVDD.n8219 0.0380882
R34302 DVDD.n14487 DVDD.n14483 0.0380882
R34303 DVDD.n14491 DVDD.n14487 0.0380882
R34304 DVDD.n14491 DVDD.n8217 0.0380882
R34305 DVDD.n14495 DVDD.n8217 0.0380882
R34306 DVDD.n14499 DVDD.n14495 0.0380882
R34307 DVDD.n14503 DVDD.n14499 0.0380882
R34308 DVDD.n14503 DVDD.n8215 0.0380882
R34309 DVDD.n14507 DVDD.n8215 0.0380882
R34310 DVDD.n14511 DVDD.n14507 0.0380882
R34311 DVDD.n14515 DVDD.n14511 0.0380882
R34312 DVDD.n14515 DVDD.n8213 0.0380882
R34313 DVDD.n14519 DVDD.n8213 0.0380882
R34314 DVDD.n14523 DVDD.n14519 0.0380882
R34315 DVDD.n14527 DVDD.n14523 0.0380882
R34316 DVDD.n14527 DVDD.n8211 0.0380882
R34317 DVDD.n14531 DVDD.n8211 0.0380882
R34318 DVDD.n14535 DVDD.n14531 0.0380882
R34319 DVDD.n14539 DVDD.n14535 0.0380882
R34320 DVDD.n14539 DVDD.n8209 0.0380882
R34321 DVDD.n14543 DVDD.n8209 0.0380882
R34322 DVDD.n14547 DVDD.n14543 0.0380882
R34323 DVDD.n14551 DVDD.n14547 0.0380882
R34324 DVDD.n14551 DVDD.n8207 0.0380882
R34325 DVDD.n14555 DVDD.n8207 0.0380882
R34326 DVDD.n14555 DVDD.n8206 0.0380882
R34327 DVDD.n8347 DVDD.n8345 0.0380882
R34328 DVDD.n8357 DVDD.n8345 0.0380882
R34329 DVDD.n8358 DVDD.n8357 0.0380882
R34330 DVDD.n8359 DVDD.n8358 0.0380882
R34331 DVDD.n8359 DVDD.n8341 0.0380882
R34332 DVDD.n8369 DVDD.n8341 0.0380882
R34333 DVDD.n8370 DVDD.n8369 0.0380882
R34334 DVDD.n8371 DVDD.n8370 0.0380882
R34335 DVDD.n8371 DVDD.n8337 0.0380882
R34336 DVDD.n8381 DVDD.n8337 0.0380882
R34337 DVDD.n8382 DVDD.n8381 0.0380882
R34338 DVDD.n8383 DVDD.n8382 0.0380882
R34339 DVDD.n8383 DVDD.n8333 0.0380882
R34340 DVDD.n8393 DVDD.n8333 0.0380882
R34341 DVDD.n8394 DVDD.n8393 0.0380882
R34342 DVDD.n8395 DVDD.n8394 0.0380882
R34343 DVDD.n8395 DVDD.n8329 0.0380882
R34344 DVDD.n8405 DVDD.n8329 0.0380882
R34345 DVDD.n8406 DVDD.n8405 0.0380882
R34346 DVDD.n8407 DVDD.n8406 0.0380882
R34347 DVDD.n8407 DVDD.n8325 0.0380882
R34348 DVDD.n8417 DVDD.n8325 0.0380882
R34349 DVDD.n8418 DVDD.n8417 0.0380882
R34350 DVDD.n8419 DVDD.n8418 0.0380882
R34351 DVDD.n8419 DVDD.n8321 0.0380882
R34352 DVDD.n8429 DVDD.n8321 0.0380882
R34353 DVDD.n8430 DVDD.n8429 0.0380882
R34354 DVDD.n8431 DVDD.n8430 0.0380882
R34355 DVDD.n8431 DVDD.n8317 0.0380882
R34356 DVDD.n8441 DVDD.n8317 0.0380882
R34357 DVDD.n8442 DVDD.n8441 0.0380882
R34358 DVDD.n8443 DVDD.n8442 0.0380882
R34359 DVDD.n8443 DVDD.n8313 0.0380882
R34360 DVDD.n8453 DVDD.n8313 0.0380882
R34361 DVDD.n8454 DVDD.n8453 0.0380882
R34362 DVDD.n8455 DVDD.n8454 0.0380882
R34363 DVDD.n8455 DVDD.n8309 0.0380882
R34364 DVDD.n8465 DVDD.n8309 0.0380882
R34365 DVDD.n8466 DVDD.n8465 0.0380882
R34366 DVDD.n8467 DVDD.n8466 0.0380882
R34367 DVDD.n8467 DVDD.n8305 0.0380882
R34368 DVDD.n8477 DVDD.n8305 0.0380882
R34369 DVDD.n8478 DVDD.n8477 0.0380882
R34370 DVDD.n8479 DVDD.n8478 0.0380882
R34371 DVDD.n8479 DVDD.n8301 0.0380882
R34372 DVDD.n8489 DVDD.n8301 0.0380882
R34373 DVDD.n8490 DVDD.n8489 0.0380882
R34374 DVDD.n8491 DVDD.n8490 0.0380882
R34375 DVDD.n8491 DVDD.n8297 0.0380882
R34376 DVDD.n8501 DVDD.n8297 0.0380882
R34377 DVDD.n8502 DVDD.n8501 0.0380882
R34378 DVDD.n8503 DVDD.n8502 0.0380882
R34379 DVDD.n8503 DVDD.n8293 0.0380882
R34380 DVDD.n8513 DVDD.n8293 0.0380882
R34381 DVDD.n8514 DVDD.n8513 0.0380882
R34382 DVDD.n8515 DVDD.n8514 0.0380882
R34383 DVDD.n8515 DVDD.n8289 0.0380882
R34384 DVDD.n8525 DVDD.n8289 0.0380882
R34385 DVDD.n8526 DVDD.n8525 0.0380882
R34386 DVDD.n8527 DVDD.n8526 0.0380882
R34387 DVDD.n8527 DVDD.n8285 0.0380882
R34388 DVDD.n8537 DVDD.n8285 0.0380882
R34389 DVDD.n8538 DVDD.n8537 0.0380882
R34390 DVDD.n8539 DVDD.n8538 0.0380882
R34391 DVDD.n8539 DVDD.n8281 0.0380882
R34392 DVDD.n8549 DVDD.n8281 0.0380882
R34393 DVDD.n8550 DVDD.n8549 0.0380882
R34394 DVDD.n8551 DVDD.n8550 0.0380882
R34395 DVDD.n8551 DVDD.n8277 0.0380882
R34396 DVDD.n8561 DVDD.n8277 0.0380882
R34397 DVDD.n8562 DVDD.n8561 0.0380882
R34398 DVDD.n8563 DVDD.n8562 0.0380882
R34399 DVDD.n8563 DVDD.n8273 0.0380882
R34400 DVDD.n8573 DVDD.n8273 0.0380882
R34401 DVDD.n8574 DVDD.n8573 0.0380882
R34402 DVDD.n8575 DVDD.n8574 0.0380882
R34403 DVDD.n8575 DVDD.n8269 0.0380882
R34404 DVDD.n8585 DVDD.n8269 0.0380882
R34405 DVDD.n8586 DVDD.n8585 0.0380882
R34406 DVDD.n8588 DVDD.n8586 0.0380882
R34407 DVDD.n8588 DVDD.n8587 0.0380882
R34408 DVDD.n8587 DVDD.n8264 0.0380882
R34409 DVDD.n8598 DVDD.n8264 0.0380882
R34410 DVDD.n8348 DVDD.n8346 0.0380882
R34411 DVDD.n8356 DVDD.n8346 0.0380882
R34412 DVDD.n8356 DVDD.n8344 0.0380882
R34413 DVDD.n8360 DVDD.n8344 0.0380882
R34414 DVDD.n8360 DVDD.n8342 0.0380882
R34415 DVDD.n8368 DVDD.n8342 0.0380882
R34416 DVDD.n8368 DVDD.n8340 0.0380882
R34417 DVDD.n8372 DVDD.n8340 0.0380882
R34418 DVDD.n8372 DVDD.n8338 0.0380882
R34419 DVDD.n8380 DVDD.n8338 0.0380882
R34420 DVDD.n8380 DVDD.n8336 0.0380882
R34421 DVDD.n8384 DVDD.n8336 0.0380882
R34422 DVDD.n8384 DVDD.n8334 0.0380882
R34423 DVDD.n8392 DVDD.n8334 0.0380882
R34424 DVDD.n8392 DVDD.n8332 0.0380882
R34425 DVDD.n8396 DVDD.n8332 0.0380882
R34426 DVDD.n8396 DVDD.n8330 0.0380882
R34427 DVDD.n8404 DVDD.n8330 0.0380882
R34428 DVDD.n8404 DVDD.n8328 0.0380882
R34429 DVDD.n8408 DVDD.n8328 0.0380882
R34430 DVDD.n8408 DVDD.n8326 0.0380882
R34431 DVDD.n8416 DVDD.n8326 0.0380882
R34432 DVDD.n8416 DVDD.n8324 0.0380882
R34433 DVDD.n8420 DVDD.n8324 0.0380882
R34434 DVDD.n8420 DVDD.n8322 0.0380882
R34435 DVDD.n8428 DVDD.n8322 0.0380882
R34436 DVDD.n8428 DVDD.n8320 0.0380882
R34437 DVDD.n8432 DVDD.n8320 0.0380882
R34438 DVDD.n8432 DVDD.n8318 0.0380882
R34439 DVDD.n8440 DVDD.n8318 0.0380882
R34440 DVDD.n8440 DVDD.n8316 0.0380882
R34441 DVDD.n8444 DVDD.n8316 0.0380882
R34442 DVDD.n8444 DVDD.n8314 0.0380882
R34443 DVDD.n8452 DVDD.n8314 0.0380882
R34444 DVDD.n8452 DVDD.n8312 0.0380882
R34445 DVDD.n8456 DVDD.n8312 0.0380882
R34446 DVDD.n8456 DVDD.n8310 0.0380882
R34447 DVDD.n8464 DVDD.n8310 0.0380882
R34448 DVDD.n8464 DVDD.n8308 0.0380882
R34449 DVDD.n8468 DVDD.n8308 0.0380882
R34450 DVDD.n8468 DVDD.n8306 0.0380882
R34451 DVDD.n8476 DVDD.n8306 0.0380882
R34452 DVDD.n8476 DVDD.n8304 0.0380882
R34453 DVDD.n8480 DVDD.n8304 0.0380882
R34454 DVDD.n8480 DVDD.n8302 0.0380882
R34455 DVDD.n8488 DVDD.n8302 0.0380882
R34456 DVDD.n8488 DVDD.n8300 0.0380882
R34457 DVDD.n8492 DVDD.n8300 0.0380882
R34458 DVDD.n8492 DVDD.n8298 0.0380882
R34459 DVDD.n8500 DVDD.n8298 0.0380882
R34460 DVDD.n8500 DVDD.n8296 0.0380882
R34461 DVDD.n8504 DVDD.n8296 0.0380882
R34462 DVDD.n8504 DVDD.n8294 0.0380882
R34463 DVDD.n8512 DVDD.n8294 0.0380882
R34464 DVDD.n8512 DVDD.n8292 0.0380882
R34465 DVDD.n8516 DVDD.n8292 0.0380882
R34466 DVDD.n8516 DVDD.n8290 0.0380882
R34467 DVDD.n8524 DVDD.n8290 0.0380882
R34468 DVDD.n8524 DVDD.n8288 0.0380882
R34469 DVDD.n8528 DVDD.n8288 0.0380882
R34470 DVDD.n8528 DVDD.n8286 0.0380882
R34471 DVDD.n8536 DVDD.n8286 0.0380882
R34472 DVDD.n8536 DVDD.n8284 0.0380882
R34473 DVDD.n8540 DVDD.n8284 0.0380882
R34474 DVDD.n8540 DVDD.n8282 0.0380882
R34475 DVDD.n8548 DVDD.n8282 0.0380882
R34476 DVDD.n8548 DVDD.n8280 0.0380882
R34477 DVDD.n8552 DVDD.n8280 0.0380882
R34478 DVDD.n8552 DVDD.n8278 0.0380882
R34479 DVDD.n8560 DVDD.n8278 0.0380882
R34480 DVDD.n8560 DVDD.n8276 0.0380882
R34481 DVDD.n8564 DVDD.n8276 0.0380882
R34482 DVDD.n8564 DVDD.n8274 0.0380882
R34483 DVDD.n8572 DVDD.n8274 0.0380882
R34484 DVDD.n8572 DVDD.n8272 0.0380882
R34485 DVDD.n8576 DVDD.n8272 0.0380882
R34486 DVDD.n8576 DVDD.n8270 0.0380882
R34487 DVDD.n8584 DVDD.n8270 0.0380882
R34488 DVDD.n8584 DVDD.n8268 0.0380882
R34489 DVDD.n8589 DVDD.n8268 0.0380882
R34490 DVDD.n8589 DVDD.n8266 0.0380882
R34491 DVDD.n8266 DVDD.n8265 0.0380882
R34492 DVDD.n8597 DVDD.n8265 0.0380882
R34493 DVDD.n8949 DVDD.n8615 0.0380882
R34494 DVDD.n8941 DVDD.n8615 0.0380882
R34495 DVDD.n8941 DVDD.n8940 0.0380882
R34496 DVDD.n8940 DVDD.n8939 0.0380882
R34497 DVDD.n8939 DVDD.n8619 0.0380882
R34498 DVDD.n8931 DVDD.n8619 0.0380882
R34499 DVDD.n8931 DVDD.n8930 0.0380882
R34500 DVDD.n8930 DVDD.n8929 0.0380882
R34501 DVDD.n8929 DVDD.n8625 0.0380882
R34502 DVDD.n8921 DVDD.n8625 0.0380882
R34503 DVDD.n8921 DVDD.n8920 0.0380882
R34504 DVDD.n8920 DVDD.n8919 0.0380882
R34505 DVDD.n8919 DVDD.n8631 0.0380882
R34506 DVDD.n8911 DVDD.n8631 0.0380882
R34507 DVDD.n8911 DVDD.n8910 0.0380882
R34508 DVDD.n8910 DVDD.n8909 0.0380882
R34509 DVDD.n8909 DVDD.n8637 0.0380882
R34510 DVDD.n8901 DVDD.n8637 0.0380882
R34511 DVDD.n8901 DVDD.n8900 0.0380882
R34512 DVDD.n8900 DVDD.n8899 0.0380882
R34513 DVDD.n8899 DVDD.n8643 0.0380882
R34514 DVDD.n8891 DVDD.n8643 0.0380882
R34515 DVDD.n8891 DVDD.n8890 0.0380882
R34516 DVDD.n8890 DVDD.n8889 0.0380882
R34517 DVDD.n8889 DVDD.n8649 0.0380882
R34518 DVDD.n8881 DVDD.n8649 0.0380882
R34519 DVDD.n8881 DVDD.n8880 0.0380882
R34520 DVDD.n8880 DVDD.n8879 0.0380882
R34521 DVDD.n8879 DVDD.n8655 0.0380882
R34522 DVDD.n8871 DVDD.n8655 0.0380882
R34523 DVDD.n8871 DVDD.n8870 0.0380882
R34524 DVDD.n8870 DVDD.n8869 0.0380882
R34525 DVDD.n8869 DVDD.n8661 0.0380882
R34526 DVDD.n8861 DVDD.n8661 0.0380882
R34527 DVDD.n8861 DVDD.n8860 0.0380882
R34528 DVDD.n8860 DVDD.n8859 0.0380882
R34529 DVDD.n8859 DVDD.n8667 0.0380882
R34530 DVDD.n8851 DVDD.n8667 0.0380882
R34531 DVDD.n8851 DVDD.n8850 0.0380882
R34532 DVDD.n8850 DVDD.n8849 0.0380882
R34533 DVDD.n8849 DVDD.n8673 0.0380882
R34534 DVDD.n8841 DVDD.n8673 0.0380882
R34535 DVDD.n8841 DVDD.n8840 0.0380882
R34536 DVDD.n8840 DVDD.n8839 0.0380882
R34537 DVDD.n8839 DVDD.n8679 0.0380882
R34538 DVDD.n8831 DVDD.n8679 0.0380882
R34539 DVDD.n8831 DVDD.n8830 0.0380882
R34540 DVDD.n8830 DVDD.n8829 0.0380882
R34541 DVDD.n8829 DVDD.n8685 0.0380882
R34542 DVDD.n8821 DVDD.n8685 0.0380882
R34543 DVDD.n8821 DVDD.n8820 0.0380882
R34544 DVDD.n8820 DVDD.n8819 0.0380882
R34545 DVDD.n8819 DVDD.n8691 0.0380882
R34546 DVDD.n8811 DVDD.n8691 0.0380882
R34547 DVDD.n8811 DVDD.n8810 0.0380882
R34548 DVDD.n8810 DVDD.n8809 0.0380882
R34549 DVDD.n8809 DVDD.n8697 0.0380882
R34550 DVDD.n8801 DVDD.n8697 0.0380882
R34551 DVDD.n8801 DVDD.n8800 0.0380882
R34552 DVDD.n8800 DVDD.n8799 0.0380882
R34553 DVDD.n8799 DVDD.n8703 0.0380882
R34554 DVDD.n8791 DVDD.n8703 0.0380882
R34555 DVDD.n8791 DVDD.n8790 0.0380882
R34556 DVDD.n8790 DVDD.n8789 0.0380882
R34557 DVDD.n8789 DVDD.n8709 0.0380882
R34558 DVDD.n8781 DVDD.n8709 0.0380882
R34559 DVDD.n8781 DVDD.n8780 0.0380882
R34560 DVDD.n8780 DVDD.n8779 0.0380882
R34561 DVDD.n8779 DVDD.n8715 0.0380882
R34562 DVDD.n8771 DVDD.n8715 0.0380882
R34563 DVDD.n8771 DVDD.n8770 0.0380882
R34564 DVDD.n8770 DVDD.n8769 0.0380882
R34565 DVDD.n8769 DVDD.n8721 0.0380882
R34566 DVDD.n8761 DVDD.n8721 0.0380882
R34567 DVDD.n8761 DVDD.n8760 0.0380882
R34568 DVDD.n8760 DVDD.n8759 0.0380882
R34569 DVDD.n8759 DVDD.n8727 0.0380882
R34570 DVDD.n8751 DVDD.n8727 0.0380882
R34571 DVDD.n8751 DVDD.n8750 0.0380882
R34572 DVDD.n8750 DVDD.n8749 0.0380882
R34573 DVDD.n8749 DVDD.n8733 0.0380882
R34574 DVDD.n8741 DVDD.n8733 0.0380882
R34575 DVDD.n8741 DVDD.n8740 0.0380882
R34576 DVDD.n8948 DVDD.n8616 0.0380882
R34577 DVDD.n8942 DVDD.n8616 0.0380882
R34578 DVDD.n8942 DVDD.n8618 0.0380882
R34579 DVDD.n8938 DVDD.n8618 0.0380882
R34580 DVDD.n8938 DVDD.n8620 0.0380882
R34581 DVDD.n8932 DVDD.n8620 0.0380882
R34582 DVDD.n8932 DVDD.n8624 0.0380882
R34583 DVDD.n8928 DVDD.n8624 0.0380882
R34584 DVDD.n8928 DVDD.n8626 0.0380882
R34585 DVDD.n8922 DVDD.n8626 0.0380882
R34586 DVDD.n8922 DVDD.n8630 0.0380882
R34587 DVDD.n8918 DVDD.n8630 0.0380882
R34588 DVDD.n8918 DVDD.n8632 0.0380882
R34589 DVDD.n8912 DVDD.n8632 0.0380882
R34590 DVDD.n8912 DVDD.n8636 0.0380882
R34591 DVDD.n8908 DVDD.n8636 0.0380882
R34592 DVDD.n8908 DVDD.n8638 0.0380882
R34593 DVDD.n8902 DVDD.n8638 0.0380882
R34594 DVDD.n8902 DVDD.n8642 0.0380882
R34595 DVDD.n8898 DVDD.n8642 0.0380882
R34596 DVDD.n8898 DVDD.n8644 0.0380882
R34597 DVDD.n8892 DVDD.n8644 0.0380882
R34598 DVDD.n8892 DVDD.n8648 0.0380882
R34599 DVDD.n8888 DVDD.n8648 0.0380882
R34600 DVDD.n8888 DVDD.n8650 0.0380882
R34601 DVDD.n8882 DVDD.n8650 0.0380882
R34602 DVDD.n8882 DVDD.n8654 0.0380882
R34603 DVDD.n8878 DVDD.n8654 0.0380882
R34604 DVDD.n8878 DVDD.n8656 0.0380882
R34605 DVDD.n8872 DVDD.n8656 0.0380882
R34606 DVDD.n8872 DVDD.n8660 0.0380882
R34607 DVDD.n8868 DVDD.n8660 0.0380882
R34608 DVDD.n8868 DVDD.n8662 0.0380882
R34609 DVDD.n8862 DVDD.n8662 0.0380882
R34610 DVDD.n8862 DVDD.n8666 0.0380882
R34611 DVDD.n8858 DVDD.n8666 0.0380882
R34612 DVDD.n8858 DVDD.n8668 0.0380882
R34613 DVDD.n8852 DVDD.n8668 0.0380882
R34614 DVDD.n8852 DVDD.n8672 0.0380882
R34615 DVDD.n8848 DVDD.n8672 0.0380882
R34616 DVDD.n8848 DVDD.n8674 0.0380882
R34617 DVDD.n8842 DVDD.n8674 0.0380882
R34618 DVDD.n8842 DVDD.n8678 0.0380882
R34619 DVDD.n8838 DVDD.n8678 0.0380882
R34620 DVDD.n8838 DVDD.n8680 0.0380882
R34621 DVDD.n8832 DVDD.n8680 0.0380882
R34622 DVDD.n8832 DVDD.n8684 0.0380882
R34623 DVDD.n8828 DVDD.n8684 0.0380882
R34624 DVDD.n8828 DVDD.n8686 0.0380882
R34625 DVDD.n8822 DVDD.n8686 0.0380882
R34626 DVDD.n8822 DVDD.n8690 0.0380882
R34627 DVDD.n8818 DVDD.n8690 0.0380882
R34628 DVDD.n8818 DVDD.n8692 0.0380882
R34629 DVDD.n8812 DVDD.n8692 0.0380882
R34630 DVDD.n8812 DVDD.n8696 0.0380882
R34631 DVDD.n8808 DVDD.n8696 0.0380882
R34632 DVDD.n8808 DVDD.n8698 0.0380882
R34633 DVDD.n8802 DVDD.n8698 0.0380882
R34634 DVDD.n8802 DVDD.n8702 0.0380882
R34635 DVDD.n8798 DVDD.n8702 0.0380882
R34636 DVDD.n8798 DVDD.n8704 0.0380882
R34637 DVDD.n8792 DVDD.n8704 0.0380882
R34638 DVDD.n8792 DVDD.n8708 0.0380882
R34639 DVDD.n8788 DVDD.n8708 0.0380882
R34640 DVDD.n8788 DVDD.n8710 0.0380882
R34641 DVDD.n8782 DVDD.n8710 0.0380882
R34642 DVDD.n8782 DVDD.n8714 0.0380882
R34643 DVDD.n8778 DVDD.n8714 0.0380882
R34644 DVDD.n8778 DVDD.n8716 0.0380882
R34645 DVDD.n8772 DVDD.n8716 0.0380882
R34646 DVDD.n8772 DVDD.n8720 0.0380882
R34647 DVDD.n8768 DVDD.n8720 0.0380882
R34648 DVDD.n8768 DVDD.n8722 0.0380882
R34649 DVDD.n8762 DVDD.n8722 0.0380882
R34650 DVDD.n8762 DVDD.n8726 0.0380882
R34651 DVDD.n8758 DVDD.n8726 0.0380882
R34652 DVDD.n8758 DVDD.n8728 0.0380882
R34653 DVDD.n8752 DVDD.n8728 0.0380882
R34654 DVDD.n8752 DVDD.n8732 0.0380882
R34655 DVDD.n8748 DVDD.n8732 0.0380882
R34656 DVDD.n8748 DVDD.n8734 0.0380882
R34657 DVDD.n8742 DVDD.n8734 0.0380882
R34658 DVDD.n8742 DVDD.n8739 0.0380882
R34659 DVDD.n10394 DVDD.n10392 0.0380882
R34660 DVDD.n10395 DVDD.n10394 0.0380882
R34661 DVDD.n10396 DVDD.n10395 0.0380882
R34662 DVDD.n10396 DVDD.n10389 0.0380882
R34663 DVDD.n10403 DVDD.n10389 0.0380882
R34664 DVDD.n10404 DVDD.n10403 0.0380882
R34665 DVDD.n10405 DVDD.n10404 0.0380882
R34666 DVDD.n10405 DVDD.n10386 0.0380882
R34667 DVDD.n10412 DVDD.n10386 0.0380882
R34668 DVDD.n10413 DVDD.n10412 0.0380882
R34669 DVDD.n10414 DVDD.n10413 0.0380882
R34670 DVDD.n10414 DVDD.n10383 0.0380882
R34671 DVDD.n10421 DVDD.n10383 0.0380882
R34672 DVDD.n10422 DVDD.n10421 0.0380882
R34673 DVDD.n10423 DVDD.n10422 0.0380882
R34674 DVDD.n10423 DVDD.n10380 0.0380882
R34675 DVDD.n10430 DVDD.n10380 0.0380882
R34676 DVDD.n10431 DVDD.n10430 0.0380882
R34677 DVDD.n10432 DVDD.n10431 0.0380882
R34678 DVDD.n10432 DVDD.n10377 0.0380882
R34679 DVDD.n10439 DVDD.n10377 0.0380882
R34680 DVDD.n10440 DVDD.n10439 0.0380882
R34681 DVDD.n10441 DVDD.n10440 0.0380882
R34682 DVDD.n10441 DVDD.n10374 0.0380882
R34683 DVDD.n10448 DVDD.n10374 0.0380882
R34684 DVDD.n10449 DVDD.n10448 0.0380882
R34685 DVDD.n10450 DVDD.n10449 0.0380882
R34686 DVDD.n10450 DVDD.n10371 0.0380882
R34687 DVDD.n10457 DVDD.n10371 0.0380882
R34688 DVDD.n10458 DVDD.n10457 0.0380882
R34689 DVDD.n10459 DVDD.n10458 0.0380882
R34690 DVDD.n10459 DVDD.n10368 0.0380882
R34691 DVDD.n10466 DVDD.n10368 0.0380882
R34692 DVDD.n10467 DVDD.n10466 0.0380882
R34693 DVDD.n10468 DVDD.n10467 0.0380882
R34694 DVDD.n10468 DVDD.n10365 0.0380882
R34695 DVDD.n10475 DVDD.n10365 0.0380882
R34696 DVDD.n10476 DVDD.n10475 0.0380882
R34697 DVDD.n10477 DVDD.n10476 0.0380882
R34698 DVDD.n10477 DVDD.n10362 0.0380882
R34699 DVDD.n10484 DVDD.n10362 0.0380882
R34700 DVDD.n10485 DVDD.n10484 0.0380882
R34701 DVDD.n10486 DVDD.n10485 0.0380882
R34702 DVDD.n10486 DVDD.n10359 0.0380882
R34703 DVDD.n10493 DVDD.n10359 0.0380882
R34704 DVDD.n10494 DVDD.n10493 0.0380882
R34705 DVDD.n10495 DVDD.n10494 0.0380882
R34706 DVDD.n10495 DVDD.n10356 0.0380882
R34707 DVDD.n10502 DVDD.n10356 0.0380882
R34708 DVDD.n10503 DVDD.n10502 0.0380882
R34709 DVDD.n10504 DVDD.n10503 0.0380882
R34710 DVDD.n10504 DVDD.n10353 0.0380882
R34711 DVDD.n10511 DVDD.n10353 0.0380882
R34712 DVDD.n10512 DVDD.n10511 0.0380882
R34713 DVDD.n10513 DVDD.n10512 0.0380882
R34714 DVDD.n10513 DVDD.n10350 0.0380882
R34715 DVDD.n10520 DVDD.n10350 0.0380882
R34716 DVDD.n10521 DVDD.n10520 0.0380882
R34717 DVDD.n10522 DVDD.n10521 0.0380882
R34718 DVDD.n10522 DVDD.n10347 0.0380882
R34719 DVDD.n10529 DVDD.n10347 0.0380882
R34720 DVDD.n10530 DVDD.n10529 0.0380882
R34721 DVDD.n10531 DVDD.n10530 0.0380882
R34722 DVDD.n10531 DVDD.n10344 0.0380882
R34723 DVDD.n10538 DVDD.n10344 0.0380882
R34724 DVDD.n10539 DVDD.n10538 0.0380882
R34725 DVDD.n10540 DVDD.n10539 0.0380882
R34726 DVDD.n10540 DVDD.n10341 0.0380882
R34727 DVDD.n10547 DVDD.n10341 0.0380882
R34728 DVDD.n10548 DVDD.n10547 0.0380882
R34729 DVDD.n10549 DVDD.n10548 0.0380882
R34730 DVDD.n10549 DVDD.n10338 0.0380882
R34731 DVDD.n10556 DVDD.n10338 0.0380882
R34732 DVDD.n10557 DVDD.n10556 0.0380882
R34733 DVDD.n10558 DVDD.n10557 0.0380882
R34734 DVDD.n10558 DVDD.n10335 0.0380882
R34735 DVDD.n10565 DVDD.n10335 0.0380882
R34736 DVDD.n10566 DVDD.n10565 0.0380882
R34737 DVDD.n10567 DVDD.n10566 0.0380882
R34738 DVDD.n10567 DVDD.n10332 0.0380882
R34739 DVDD.n10574 DVDD.n10332 0.0380882
R34740 DVDD.n10575 DVDD.n10574 0.0380882
R34741 DVDD.n10576 DVDD.n10575 0.0380882
R34742 DVDD.n10393 DVDD.n10285 0.0380882
R34743 DVDD.n10393 DVDD.n10391 0.0380882
R34744 DVDD.n10398 DVDD.n10391 0.0380882
R34745 DVDD.n10400 DVDD.n10398 0.0380882
R34746 DVDD.n10402 DVDD.n10400 0.0380882
R34747 DVDD.n10402 DVDD.n10388 0.0380882
R34748 DVDD.n10407 DVDD.n10388 0.0380882
R34749 DVDD.n10409 DVDD.n10407 0.0380882
R34750 DVDD.n10411 DVDD.n10409 0.0380882
R34751 DVDD.n10411 DVDD.n10385 0.0380882
R34752 DVDD.n10416 DVDD.n10385 0.0380882
R34753 DVDD.n10418 DVDD.n10416 0.0380882
R34754 DVDD.n10420 DVDD.n10418 0.0380882
R34755 DVDD.n10420 DVDD.n10382 0.0380882
R34756 DVDD.n10425 DVDD.n10382 0.0380882
R34757 DVDD.n10427 DVDD.n10425 0.0380882
R34758 DVDD.n10429 DVDD.n10427 0.0380882
R34759 DVDD.n10429 DVDD.n10379 0.0380882
R34760 DVDD.n10434 DVDD.n10379 0.0380882
R34761 DVDD.n10436 DVDD.n10434 0.0380882
R34762 DVDD.n10438 DVDD.n10436 0.0380882
R34763 DVDD.n10438 DVDD.n10376 0.0380882
R34764 DVDD.n10443 DVDD.n10376 0.0380882
R34765 DVDD.n10445 DVDD.n10443 0.0380882
R34766 DVDD.n10447 DVDD.n10445 0.0380882
R34767 DVDD.n10447 DVDD.n10373 0.0380882
R34768 DVDD.n10452 DVDD.n10373 0.0380882
R34769 DVDD.n10454 DVDD.n10452 0.0380882
R34770 DVDD.n10456 DVDD.n10454 0.0380882
R34771 DVDD.n10456 DVDD.n10370 0.0380882
R34772 DVDD.n10461 DVDD.n10370 0.0380882
R34773 DVDD.n10463 DVDD.n10461 0.0380882
R34774 DVDD.n10465 DVDD.n10463 0.0380882
R34775 DVDD.n10465 DVDD.n10367 0.0380882
R34776 DVDD.n10470 DVDD.n10367 0.0380882
R34777 DVDD.n10472 DVDD.n10470 0.0380882
R34778 DVDD.n10474 DVDD.n10472 0.0380882
R34779 DVDD.n10474 DVDD.n10364 0.0380882
R34780 DVDD.n10479 DVDD.n10364 0.0380882
R34781 DVDD.n10481 DVDD.n10479 0.0380882
R34782 DVDD.n10483 DVDD.n10481 0.0380882
R34783 DVDD.n10483 DVDD.n10361 0.0380882
R34784 DVDD.n10488 DVDD.n10361 0.0380882
R34785 DVDD.n10490 DVDD.n10488 0.0380882
R34786 DVDD.n10492 DVDD.n10490 0.0380882
R34787 DVDD.n10492 DVDD.n10358 0.0380882
R34788 DVDD.n10497 DVDD.n10358 0.0380882
R34789 DVDD.n10499 DVDD.n10497 0.0380882
R34790 DVDD.n10501 DVDD.n10499 0.0380882
R34791 DVDD.n10501 DVDD.n10355 0.0380882
R34792 DVDD.n10506 DVDD.n10355 0.0380882
R34793 DVDD.n10508 DVDD.n10506 0.0380882
R34794 DVDD.n10510 DVDD.n10508 0.0380882
R34795 DVDD.n10510 DVDD.n10352 0.0380882
R34796 DVDD.n10515 DVDD.n10352 0.0380882
R34797 DVDD.n10517 DVDD.n10515 0.0380882
R34798 DVDD.n10519 DVDD.n10517 0.0380882
R34799 DVDD.n10519 DVDD.n10349 0.0380882
R34800 DVDD.n10524 DVDD.n10349 0.0380882
R34801 DVDD.n10526 DVDD.n10524 0.0380882
R34802 DVDD.n10528 DVDD.n10526 0.0380882
R34803 DVDD.n10528 DVDD.n10346 0.0380882
R34804 DVDD.n10533 DVDD.n10346 0.0380882
R34805 DVDD.n10535 DVDD.n10533 0.0380882
R34806 DVDD.n10537 DVDD.n10535 0.0380882
R34807 DVDD.n10537 DVDD.n10343 0.0380882
R34808 DVDD.n10542 DVDD.n10343 0.0380882
R34809 DVDD.n10544 DVDD.n10542 0.0380882
R34810 DVDD.n10546 DVDD.n10544 0.0380882
R34811 DVDD.n10546 DVDD.n10340 0.0380882
R34812 DVDD.n10551 DVDD.n10340 0.0380882
R34813 DVDD.n10553 DVDD.n10551 0.0380882
R34814 DVDD.n10555 DVDD.n10553 0.0380882
R34815 DVDD.n10555 DVDD.n10337 0.0380882
R34816 DVDD.n10560 DVDD.n10337 0.0380882
R34817 DVDD.n10562 DVDD.n10560 0.0380882
R34818 DVDD.n10564 DVDD.n10562 0.0380882
R34819 DVDD.n10564 DVDD.n10334 0.0380882
R34820 DVDD.n10569 DVDD.n10334 0.0380882
R34821 DVDD.n10571 DVDD.n10569 0.0380882
R34822 DVDD.n10573 DVDD.n10571 0.0380882
R34823 DVDD.n10573 DVDD.n10331 0.0380882
R34824 DVDD.n14279 DVDD.n10331 0.0380882
R34825 DVDD.n14023 DVDD.n14022 0.0380882
R34826 DVDD.n14024 DVDD.n14023 0.0380882
R34827 DVDD.n14024 DVDD.n10682 0.0380882
R34828 DVDD.n14034 DVDD.n10682 0.0380882
R34829 DVDD.n14035 DVDD.n14034 0.0380882
R34830 DVDD.n14036 DVDD.n14035 0.0380882
R34831 DVDD.n14036 DVDD.n10680 0.0380882
R34832 DVDD.n14046 DVDD.n10680 0.0380882
R34833 DVDD.n14047 DVDD.n14046 0.0380882
R34834 DVDD.n14048 DVDD.n14047 0.0380882
R34835 DVDD.n14048 DVDD.n10678 0.0380882
R34836 DVDD.n14058 DVDD.n10678 0.0380882
R34837 DVDD.n14059 DVDD.n14058 0.0380882
R34838 DVDD.n14060 DVDD.n14059 0.0380882
R34839 DVDD.n14060 DVDD.n10676 0.0380882
R34840 DVDD.n14070 DVDD.n10676 0.0380882
R34841 DVDD.n14071 DVDD.n14070 0.0380882
R34842 DVDD.n14072 DVDD.n14071 0.0380882
R34843 DVDD.n14072 DVDD.n10674 0.0380882
R34844 DVDD.n14082 DVDD.n10674 0.0380882
R34845 DVDD.n14083 DVDD.n14082 0.0380882
R34846 DVDD.n14084 DVDD.n14083 0.0380882
R34847 DVDD.n14084 DVDD.n10672 0.0380882
R34848 DVDD.n14094 DVDD.n10672 0.0380882
R34849 DVDD.n14095 DVDD.n14094 0.0380882
R34850 DVDD.n14096 DVDD.n14095 0.0380882
R34851 DVDD.n14096 DVDD.n10670 0.0380882
R34852 DVDD.n14106 DVDD.n10670 0.0380882
R34853 DVDD.n14107 DVDD.n14106 0.0380882
R34854 DVDD.n14108 DVDD.n14107 0.0380882
R34855 DVDD.n14108 DVDD.n10668 0.0380882
R34856 DVDD.n14118 DVDD.n10668 0.0380882
R34857 DVDD.n14119 DVDD.n14118 0.0380882
R34858 DVDD.n14120 DVDD.n14119 0.0380882
R34859 DVDD.n14120 DVDD.n10666 0.0380882
R34860 DVDD.n14130 DVDD.n10666 0.0380882
R34861 DVDD.n14131 DVDD.n14130 0.0380882
R34862 DVDD.n14132 DVDD.n14131 0.0380882
R34863 DVDD.n14132 DVDD.n10664 0.0380882
R34864 DVDD.n14142 DVDD.n10664 0.0380882
R34865 DVDD.n14143 DVDD.n14142 0.0380882
R34866 DVDD.n14144 DVDD.n14143 0.0380882
R34867 DVDD.n14144 DVDD.n10662 0.0380882
R34868 DVDD.n14154 DVDD.n10662 0.0380882
R34869 DVDD.n14155 DVDD.n14154 0.0380882
R34870 DVDD.n14156 DVDD.n14155 0.0380882
R34871 DVDD.n14156 DVDD.n10660 0.0380882
R34872 DVDD.n14166 DVDD.n10660 0.0380882
R34873 DVDD.n14167 DVDD.n14166 0.0380882
R34874 DVDD.n14168 DVDD.n14167 0.0380882
R34875 DVDD.n14168 DVDD.n10658 0.0380882
R34876 DVDD.n14178 DVDD.n10658 0.0380882
R34877 DVDD.n14179 DVDD.n14178 0.0380882
R34878 DVDD.n14180 DVDD.n14179 0.0380882
R34879 DVDD.n14180 DVDD.n10656 0.0380882
R34880 DVDD.n14190 DVDD.n10656 0.0380882
R34881 DVDD.n14191 DVDD.n14190 0.0380882
R34882 DVDD.n14192 DVDD.n14191 0.0380882
R34883 DVDD.n14192 DVDD.n10654 0.0380882
R34884 DVDD.n14202 DVDD.n10654 0.0380882
R34885 DVDD.n14203 DVDD.n14202 0.0380882
R34886 DVDD.n14204 DVDD.n14203 0.0380882
R34887 DVDD.n14204 DVDD.n10652 0.0380882
R34888 DVDD.n14214 DVDD.n10652 0.0380882
R34889 DVDD.n14215 DVDD.n14214 0.0380882
R34890 DVDD.n14216 DVDD.n14215 0.0380882
R34891 DVDD.n14216 DVDD.n10650 0.0380882
R34892 DVDD.n14226 DVDD.n10650 0.0380882
R34893 DVDD.n14227 DVDD.n14226 0.0380882
R34894 DVDD.n14228 DVDD.n14227 0.0380882
R34895 DVDD.n14228 DVDD.n10648 0.0380882
R34896 DVDD.n14238 DVDD.n10648 0.0380882
R34897 DVDD.n14239 DVDD.n14238 0.0380882
R34898 DVDD.n14240 DVDD.n14239 0.0380882
R34899 DVDD.n14240 DVDD.n10646 0.0380882
R34900 DVDD.n14250 DVDD.n10646 0.0380882
R34901 DVDD.n14251 DVDD.n14250 0.0380882
R34902 DVDD.n14252 DVDD.n14251 0.0380882
R34903 DVDD.n14252 DVDD.n10644 0.0380882
R34904 DVDD.n14262 DVDD.n10644 0.0380882
R34905 DVDD.n14263 DVDD.n14262 0.0380882
R34906 DVDD.n14264 DVDD.n14263 0.0380882
R34907 DVDD.n14264 DVDD.n10591 0.0380882
R34908 DVDD.n14021 DVDD.n10685 0.0380882
R34909 DVDD.n14025 DVDD.n10685 0.0380882
R34910 DVDD.n14029 DVDD.n14025 0.0380882
R34911 DVDD.n14033 DVDD.n14029 0.0380882
R34912 DVDD.n14033 DVDD.n10681 0.0380882
R34913 DVDD.n14037 DVDD.n10681 0.0380882
R34914 DVDD.n14041 DVDD.n14037 0.0380882
R34915 DVDD.n14045 DVDD.n14041 0.0380882
R34916 DVDD.n14045 DVDD.n10679 0.0380882
R34917 DVDD.n14049 DVDD.n10679 0.0380882
R34918 DVDD.n14053 DVDD.n14049 0.0380882
R34919 DVDD.n14057 DVDD.n14053 0.0380882
R34920 DVDD.n14057 DVDD.n10677 0.0380882
R34921 DVDD.n14061 DVDD.n10677 0.0380882
R34922 DVDD.n14065 DVDD.n14061 0.0380882
R34923 DVDD.n14069 DVDD.n14065 0.0380882
R34924 DVDD.n14069 DVDD.n10675 0.0380882
R34925 DVDD.n14073 DVDD.n10675 0.0380882
R34926 DVDD.n14077 DVDD.n14073 0.0380882
R34927 DVDD.n14081 DVDD.n14077 0.0380882
R34928 DVDD.n14081 DVDD.n10673 0.0380882
R34929 DVDD.n14085 DVDD.n10673 0.0380882
R34930 DVDD.n14089 DVDD.n14085 0.0380882
R34931 DVDD.n14093 DVDD.n14089 0.0380882
R34932 DVDD.n14093 DVDD.n10671 0.0380882
R34933 DVDD.n14097 DVDD.n10671 0.0380882
R34934 DVDD.n14101 DVDD.n14097 0.0380882
R34935 DVDD.n14105 DVDD.n14101 0.0380882
R34936 DVDD.n14105 DVDD.n10669 0.0380882
R34937 DVDD.n14109 DVDD.n10669 0.0380882
R34938 DVDD.n14113 DVDD.n14109 0.0380882
R34939 DVDD.n14117 DVDD.n14113 0.0380882
R34940 DVDD.n14117 DVDD.n10667 0.0380882
R34941 DVDD.n14121 DVDD.n10667 0.0380882
R34942 DVDD.n14125 DVDD.n14121 0.0380882
R34943 DVDD.n14129 DVDD.n14125 0.0380882
R34944 DVDD.n14129 DVDD.n10665 0.0380882
R34945 DVDD.n14133 DVDD.n10665 0.0380882
R34946 DVDD.n14137 DVDD.n14133 0.0380882
R34947 DVDD.n14141 DVDD.n14137 0.0380882
R34948 DVDD.n14141 DVDD.n10663 0.0380882
R34949 DVDD.n14145 DVDD.n10663 0.0380882
R34950 DVDD.n14149 DVDD.n14145 0.0380882
R34951 DVDD.n14153 DVDD.n14149 0.0380882
R34952 DVDD.n14153 DVDD.n10661 0.0380882
R34953 DVDD.n14157 DVDD.n10661 0.0380882
R34954 DVDD.n14161 DVDD.n14157 0.0380882
R34955 DVDD.n14165 DVDD.n14161 0.0380882
R34956 DVDD.n14165 DVDD.n10659 0.0380882
R34957 DVDD.n14169 DVDD.n10659 0.0380882
R34958 DVDD.n14173 DVDD.n14169 0.0380882
R34959 DVDD.n14177 DVDD.n14173 0.0380882
R34960 DVDD.n14177 DVDD.n10657 0.0380882
R34961 DVDD.n14181 DVDD.n10657 0.0380882
R34962 DVDD.n14185 DVDD.n14181 0.0380882
R34963 DVDD.n14189 DVDD.n14185 0.0380882
R34964 DVDD.n14189 DVDD.n10655 0.0380882
R34965 DVDD.n14193 DVDD.n10655 0.0380882
R34966 DVDD.n14197 DVDD.n14193 0.0380882
R34967 DVDD.n14201 DVDD.n14197 0.0380882
R34968 DVDD.n14201 DVDD.n10653 0.0380882
R34969 DVDD.n14205 DVDD.n10653 0.0380882
R34970 DVDD.n14209 DVDD.n14205 0.0380882
R34971 DVDD.n14213 DVDD.n14209 0.0380882
R34972 DVDD.n14213 DVDD.n10651 0.0380882
R34973 DVDD.n14217 DVDD.n10651 0.0380882
R34974 DVDD.n14221 DVDD.n14217 0.0380882
R34975 DVDD.n14225 DVDD.n14221 0.0380882
R34976 DVDD.n14225 DVDD.n10649 0.0380882
R34977 DVDD.n14229 DVDD.n10649 0.0380882
R34978 DVDD.n14233 DVDD.n14229 0.0380882
R34979 DVDD.n14237 DVDD.n14233 0.0380882
R34980 DVDD.n14237 DVDD.n10647 0.0380882
R34981 DVDD.n14241 DVDD.n10647 0.0380882
R34982 DVDD.n14245 DVDD.n14241 0.0380882
R34983 DVDD.n14249 DVDD.n14245 0.0380882
R34984 DVDD.n14249 DVDD.n10645 0.0380882
R34985 DVDD.n14253 DVDD.n10645 0.0380882
R34986 DVDD.n14257 DVDD.n14253 0.0380882
R34987 DVDD.n14261 DVDD.n14257 0.0380882
R34988 DVDD.n14261 DVDD.n10643 0.0380882
R34989 DVDD.n14265 DVDD.n10643 0.0380882
R34990 DVDD.n14265 DVDD.n10641 0.0380882
R34991 DVDD.n10799 DVDD.n10797 0.0380882
R34992 DVDD.n10809 DVDD.n10797 0.0380882
R34993 DVDD.n10810 DVDD.n10809 0.0380882
R34994 DVDD.n10811 DVDD.n10810 0.0380882
R34995 DVDD.n10811 DVDD.n10793 0.0380882
R34996 DVDD.n10821 DVDD.n10793 0.0380882
R34997 DVDD.n10822 DVDD.n10821 0.0380882
R34998 DVDD.n10823 DVDD.n10822 0.0380882
R34999 DVDD.n10823 DVDD.n10789 0.0380882
R35000 DVDD.n10833 DVDD.n10789 0.0380882
R35001 DVDD.n10834 DVDD.n10833 0.0380882
R35002 DVDD.n10835 DVDD.n10834 0.0380882
R35003 DVDD.n10835 DVDD.n10785 0.0380882
R35004 DVDD.n10845 DVDD.n10785 0.0380882
R35005 DVDD.n10846 DVDD.n10845 0.0380882
R35006 DVDD.n10847 DVDD.n10846 0.0380882
R35007 DVDD.n10847 DVDD.n10781 0.0380882
R35008 DVDD.n10857 DVDD.n10781 0.0380882
R35009 DVDD.n10858 DVDD.n10857 0.0380882
R35010 DVDD.n10859 DVDD.n10858 0.0380882
R35011 DVDD.n10859 DVDD.n10777 0.0380882
R35012 DVDD.n10869 DVDD.n10777 0.0380882
R35013 DVDD.n10870 DVDD.n10869 0.0380882
R35014 DVDD.n10871 DVDD.n10870 0.0380882
R35015 DVDD.n10871 DVDD.n10773 0.0380882
R35016 DVDD.n10881 DVDD.n10773 0.0380882
R35017 DVDD.n10882 DVDD.n10881 0.0380882
R35018 DVDD.n10883 DVDD.n10882 0.0380882
R35019 DVDD.n10883 DVDD.n10769 0.0380882
R35020 DVDD.n10893 DVDD.n10769 0.0380882
R35021 DVDD.n10894 DVDD.n10893 0.0380882
R35022 DVDD.n10895 DVDD.n10894 0.0380882
R35023 DVDD.n10895 DVDD.n10765 0.0380882
R35024 DVDD.n10905 DVDD.n10765 0.0380882
R35025 DVDD.n10906 DVDD.n10905 0.0380882
R35026 DVDD.n10907 DVDD.n10906 0.0380882
R35027 DVDD.n10907 DVDD.n10761 0.0380882
R35028 DVDD.n10917 DVDD.n10761 0.0380882
R35029 DVDD.n10918 DVDD.n10917 0.0380882
R35030 DVDD.n10919 DVDD.n10918 0.0380882
R35031 DVDD.n10919 DVDD.n10757 0.0380882
R35032 DVDD.n10929 DVDD.n10757 0.0380882
R35033 DVDD.n10930 DVDD.n10929 0.0380882
R35034 DVDD.n10931 DVDD.n10930 0.0380882
R35035 DVDD.n10931 DVDD.n10753 0.0380882
R35036 DVDD.n10941 DVDD.n10753 0.0380882
R35037 DVDD.n10942 DVDD.n10941 0.0380882
R35038 DVDD.n10943 DVDD.n10942 0.0380882
R35039 DVDD.n10943 DVDD.n10749 0.0380882
R35040 DVDD.n10953 DVDD.n10749 0.0380882
R35041 DVDD.n10954 DVDD.n10953 0.0380882
R35042 DVDD.n10955 DVDD.n10954 0.0380882
R35043 DVDD.n10955 DVDD.n10745 0.0380882
R35044 DVDD.n10965 DVDD.n10745 0.0380882
R35045 DVDD.n10966 DVDD.n10965 0.0380882
R35046 DVDD.n10967 DVDD.n10966 0.0380882
R35047 DVDD.n10967 DVDD.n10741 0.0380882
R35048 DVDD.n10977 DVDD.n10741 0.0380882
R35049 DVDD.n10978 DVDD.n10977 0.0380882
R35050 DVDD.n10979 DVDD.n10978 0.0380882
R35051 DVDD.n10979 DVDD.n10737 0.0380882
R35052 DVDD.n10989 DVDD.n10737 0.0380882
R35053 DVDD.n10990 DVDD.n10989 0.0380882
R35054 DVDD.n10991 DVDD.n10990 0.0380882
R35055 DVDD.n10991 DVDD.n10733 0.0380882
R35056 DVDD.n11001 DVDD.n10733 0.0380882
R35057 DVDD.n11002 DVDD.n11001 0.0380882
R35058 DVDD.n11003 DVDD.n11002 0.0380882
R35059 DVDD.n11003 DVDD.n10729 0.0380882
R35060 DVDD.n11013 DVDD.n10729 0.0380882
R35061 DVDD.n11014 DVDD.n11013 0.0380882
R35062 DVDD.n11015 DVDD.n11014 0.0380882
R35063 DVDD.n11015 DVDD.n10725 0.0380882
R35064 DVDD.n11025 DVDD.n10725 0.0380882
R35065 DVDD.n11026 DVDD.n11025 0.0380882
R35066 DVDD.n11027 DVDD.n11026 0.0380882
R35067 DVDD.n11027 DVDD.n10721 0.0380882
R35068 DVDD.n11037 DVDD.n10721 0.0380882
R35069 DVDD.n11038 DVDD.n11037 0.0380882
R35070 DVDD.n11040 DVDD.n11038 0.0380882
R35071 DVDD.n11040 DVDD.n11039 0.0380882
R35072 DVDD.n11039 DVDD.n10716 0.0380882
R35073 DVDD.n11050 DVDD.n10716 0.0380882
R35074 DVDD.n10800 DVDD.n10798 0.0380882
R35075 DVDD.n10808 DVDD.n10798 0.0380882
R35076 DVDD.n10808 DVDD.n10796 0.0380882
R35077 DVDD.n10812 DVDD.n10796 0.0380882
R35078 DVDD.n10812 DVDD.n10794 0.0380882
R35079 DVDD.n10820 DVDD.n10794 0.0380882
R35080 DVDD.n10820 DVDD.n10792 0.0380882
R35081 DVDD.n10824 DVDD.n10792 0.0380882
R35082 DVDD.n10824 DVDD.n10790 0.0380882
R35083 DVDD.n10832 DVDD.n10790 0.0380882
R35084 DVDD.n10832 DVDD.n10788 0.0380882
R35085 DVDD.n10836 DVDD.n10788 0.0380882
R35086 DVDD.n10836 DVDD.n10786 0.0380882
R35087 DVDD.n10844 DVDD.n10786 0.0380882
R35088 DVDD.n10844 DVDD.n10784 0.0380882
R35089 DVDD.n10848 DVDD.n10784 0.0380882
R35090 DVDD.n10848 DVDD.n10782 0.0380882
R35091 DVDD.n10856 DVDD.n10782 0.0380882
R35092 DVDD.n10856 DVDD.n10780 0.0380882
R35093 DVDD.n10860 DVDD.n10780 0.0380882
R35094 DVDD.n10860 DVDD.n10778 0.0380882
R35095 DVDD.n10868 DVDD.n10778 0.0380882
R35096 DVDD.n10868 DVDD.n10776 0.0380882
R35097 DVDD.n10872 DVDD.n10776 0.0380882
R35098 DVDD.n10872 DVDD.n10774 0.0380882
R35099 DVDD.n10880 DVDD.n10774 0.0380882
R35100 DVDD.n10880 DVDD.n10772 0.0380882
R35101 DVDD.n10884 DVDD.n10772 0.0380882
R35102 DVDD.n10884 DVDD.n10770 0.0380882
R35103 DVDD.n10892 DVDD.n10770 0.0380882
R35104 DVDD.n10892 DVDD.n10768 0.0380882
R35105 DVDD.n10896 DVDD.n10768 0.0380882
R35106 DVDD.n10896 DVDD.n10766 0.0380882
R35107 DVDD.n10904 DVDD.n10766 0.0380882
R35108 DVDD.n10904 DVDD.n10764 0.0380882
R35109 DVDD.n10908 DVDD.n10764 0.0380882
R35110 DVDD.n10908 DVDD.n10762 0.0380882
R35111 DVDD.n10916 DVDD.n10762 0.0380882
R35112 DVDD.n10916 DVDD.n10760 0.0380882
R35113 DVDD.n10920 DVDD.n10760 0.0380882
R35114 DVDD.n10920 DVDD.n10758 0.0380882
R35115 DVDD.n10928 DVDD.n10758 0.0380882
R35116 DVDD.n10928 DVDD.n10756 0.0380882
R35117 DVDD.n10932 DVDD.n10756 0.0380882
R35118 DVDD.n10932 DVDD.n10754 0.0380882
R35119 DVDD.n10940 DVDD.n10754 0.0380882
R35120 DVDD.n10940 DVDD.n10752 0.0380882
R35121 DVDD.n10944 DVDD.n10752 0.0380882
R35122 DVDD.n10944 DVDD.n10750 0.0380882
R35123 DVDD.n10952 DVDD.n10750 0.0380882
R35124 DVDD.n10952 DVDD.n10748 0.0380882
R35125 DVDD.n10956 DVDD.n10748 0.0380882
R35126 DVDD.n10956 DVDD.n10746 0.0380882
R35127 DVDD.n10964 DVDD.n10746 0.0380882
R35128 DVDD.n10964 DVDD.n10744 0.0380882
R35129 DVDD.n10968 DVDD.n10744 0.0380882
R35130 DVDD.n10968 DVDD.n10742 0.0380882
R35131 DVDD.n10976 DVDD.n10742 0.0380882
R35132 DVDD.n10976 DVDD.n10740 0.0380882
R35133 DVDD.n10980 DVDD.n10740 0.0380882
R35134 DVDD.n10980 DVDD.n10738 0.0380882
R35135 DVDD.n10988 DVDD.n10738 0.0380882
R35136 DVDD.n10988 DVDD.n10736 0.0380882
R35137 DVDD.n10992 DVDD.n10736 0.0380882
R35138 DVDD.n10992 DVDD.n10734 0.0380882
R35139 DVDD.n11000 DVDD.n10734 0.0380882
R35140 DVDD.n11000 DVDD.n10732 0.0380882
R35141 DVDD.n11004 DVDD.n10732 0.0380882
R35142 DVDD.n11004 DVDD.n10730 0.0380882
R35143 DVDD.n11012 DVDD.n10730 0.0380882
R35144 DVDD.n11012 DVDD.n10728 0.0380882
R35145 DVDD.n11016 DVDD.n10728 0.0380882
R35146 DVDD.n11016 DVDD.n10726 0.0380882
R35147 DVDD.n11024 DVDD.n10726 0.0380882
R35148 DVDD.n11024 DVDD.n10724 0.0380882
R35149 DVDD.n11028 DVDD.n10724 0.0380882
R35150 DVDD.n11028 DVDD.n10722 0.0380882
R35151 DVDD.n11036 DVDD.n10722 0.0380882
R35152 DVDD.n11036 DVDD.n10720 0.0380882
R35153 DVDD.n11041 DVDD.n10720 0.0380882
R35154 DVDD.n11041 DVDD.n10718 0.0380882
R35155 DVDD.n10718 DVDD.n10717 0.0380882
R35156 DVDD.n11049 DVDD.n10717 0.0380882
R35157 DVDD.n13815 DVDD.n13813 0.0380882
R35158 DVDD.n13816 DVDD.n13815 0.0380882
R35159 DVDD.n13817 DVDD.n13816 0.0380882
R35160 DVDD.n13817 DVDD.n11209 0.0380882
R35161 DVDD.n13824 DVDD.n11209 0.0380882
R35162 DVDD.n13825 DVDD.n13824 0.0380882
R35163 DVDD.n13826 DVDD.n13825 0.0380882
R35164 DVDD.n13826 DVDD.n11206 0.0380882
R35165 DVDD.n13833 DVDD.n11206 0.0380882
R35166 DVDD.n13834 DVDD.n13833 0.0380882
R35167 DVDD.n13835 DVDD.n13834 0.0380882
R35168 DVDD.n13835 DVDD.n11203 0.0380882
R35169 DVDD.n13842 DVDD.n11203 0.0380882
R35170 DVDD.n13843 DVDD.n13842 0.0380882
R35171 DVDD.n13844 DVDD.n13843 0.0380882
R35172 DVDD.n13844 DVDD.n11200 0.0380882
R35173 DVDD.n13851 DVDD.n11200 0.0380882
R35174 DVDD.n13852 DVDD.n13851 0.0380882
R35175 DVDD.n13853 DVDD.n13852 0.0380882
R35176 DVDD.n13853 DVDD.n11197 0.0380882
R35177 DVDD.n13860 DVDD.n11197 0.0380882
R35178 DVDD.n13861 DVDD.n13860 0.0380882
R35179 DVDD.n13862 DVDD.n13861 0.0380882
R35180 DVDD.n13862 DVDD.n11194 0.0380882
R35181 DVDD.n13869 DVDD.n11194 0.0380882
R35182 DVDD.n13870 DVDD.n13869 0.0380882
R35183 DVDD.n13871 DVDD.n13870 0.0380882
R35184 DVDD.n13871 DVDD.n11191 0.0380882
R35185 DVDD.n13878 DVDD.n11191 0.0380882
R35186 DVDD.n13879 DVDD.n13878 0.0380882
R35187 DVDD.n13880 DVDD.n13879 0.0380882
R35188 DVDD.n13880 DVDD.n11188 0.0380882
R35189 DVDD.n13887 DVDD.n11188 0.0380882
R35190 DVDD.n13888 DVDD.n13887 0.0380882
R35191 DVDD.n13889 DVDD.n13888 0.0380882
R35192 DVDD.n13889 DVDD.n11185 0.0380882
R35193 DVDD.n13896 DVDD.n11185 0.0380882
R35194 DVDD.n13897 DVDD.n13896 0.0380882
R35195 DVDD.n13898 DVDD.n13897 0.0380882
R35196 DVDD.n13898 DVDD.n11182 0.0380882
R35197 DVDD.n13905 DVDD.n11182 0.0380882
R35198 DVDD.n13906 DVDD.n13905 0.0380882
R35199 DVDD.n13907 DVDD.n13906 0.0380882
R35200 DVDD.n13907 DVDD.n11179 0.0380882
R35201 DVDD.n13914 DVDD.n11179 0.0380882
R35202 DVDD.n13915 DVDD.n13914 0.0380882
R35203 DVDD.n13916 DVDD.n13915 0.0380882
R35204 DVDD.n13916 DVDD.n11176 0.0380882
R35205 DVDD.n13923 DVDD.n11176 0.0380882
R35206 DVDD.n13924 DVDD.n13923 0.0380882
R35207 DVDD.n13925 DVDD.n13924 0.0380882
R35208 DVDD.n13925 DVDD.n11173 0.0380882
R35209 DVDD.n13932 DVDD.n11173 0.0380882
R35210 DVDD.n13933 DVDD.n13932 0.0380882
R35211 DVDD.n13934 DVDD.n13933 0.0380882
R35212 DVDD.n13934 DVDD.n11170 0.0380882
R35213 DVDD.n13941 DVDD.n11170 0.0380882
R35214 DVDD.n13942 DVDD.n13941 0.0380882
R35215 DVDD.n13943 DVDD.n13942 0.0380882
R35216 DVDD.n13943 DVDD.n11167 0.0380882
R35217 DVDD.n13950 DVDD.n11167 0.0380882
R35218 DVDD.n13951 DVDD.n13950 0.0380882
R35219 DVDD.n13952 DVDD.n13951 0.0380882
R35220 DVDD.n13952 DVDD.n11164 0.0380882
R35221 DVDD.n13959 DVDD.n11164 0.0380882
R35222 DVDD.n13960 DVDD.n13959 0.0380882
R35223 DVDD.n13961 DVDD.n13960 0.0380882
R35224 DVDD.n13961 DVDD.n11161 0.0380882
R35225 DVDD.n13968 DVDD.n11161 0.0380882
R35226 DVDD.n13969 DVDD.n13968 0.0380882
R35227 DVDD.n13970 DVDD.n13969 0.0380882
R35228 DVDD.n13970 DVDD.n11158 0.0380882
R35229 DVDD.n13977 DVDD.n11158 0.0380882
R35230 DVDD.n13978 DVDD.n13977 0.0380882
R35231 DVDD.n13979 DVDD.n13978 0.0380882
R35232 DVDD.n13979 DVDD.n11155 0.0380882
R35233 DVDD.n13986 DVDD.n11155 0.0380882
R35234 DVDD.n13987 DVDD.n13986 0.0380882
R35235 DVDD.n13988 DVDD.n13987 0.0380882
R35236 DVDD.n13988 DVDD.n11152 0.0380882
R35237 DVDD.n13995 DVDD.n11152 0.0380882
R35238 DVDD.n13996 DVDD.n13995 0.0380882
R35239 DVDD.n13997 DVDD.n13996 0.0380882
R35240 DVDD.n13814 DVDD.n11106 0.0380882
R35241 DVDD.n13814 DVDD.n11211 0.0380882
R35242 DVDD.n13819 DVDD.n11211 0.0380882
R35243 DVDD.n13821 DVDD.n13819 0.0380882
R35244 DVDD.n13823 DVDD.n13821 0.0380882
R35245 DVDD.n13823 DVDD.n11208 0.0380882
R35246 DVDD.n13828 DVDD.n11208 0.0380882
R35247 DVDD.n13830 DVDD.n13828 0.0380882
R35248 DVDD.n13832 DVDD.n13830 0.0380882
R35249 DVDD.n13832 DVDD.n11205 0.0380882
R35250 DVDD.n13837 DVDD.n11205 0.0380882
R35251 DVDD.n13839 DVDD.n13837 0.0380882
R35252 DVDD.n13841 DVDD.n13839 0.0380882
R35253 DVDD.n13841 DVDD.n11202 0.0380882
R35254 DVDD.n13846 DVDD.n11202 0.0380882
R35255 DVDD.n13848 DVDD.n13846 0.0380882
R35256 DVDD.n13850 DVDD.n13848 0.0380882
R35257 DVDD.n13850 DVDD.n11199 0.0380882
R35258 DVDD.n13855 DVDD.n11199 0.0380882
R35259 DVDD.n13857 DVDD.n13855 0.0380882
R35260 DVDD.n13859 DVDD.n13857 0.0380882
R35261 DVDD.n13859 DVDD.n11196 0.0380882
R35262 DVDD.n13864 DVDD.n11196 0.0380882
R35263 DVDD.n13866 DVDD.n13864 0.0380882
R35264 DVDD.n13868 DVDD.n13866 0.0380882
R35265 DVDD.n13868 DVDD.n11193 0.0380882
R35266 DVDD.n13873 DVDD.n11193 0.0380882
R35267 DVDD.n13875 DVDD.n13873 0.0380882
R35268 DVDD.n13877 DVDD.n13875 0.0380882
R35269 DVDD.n13877 DVDD.n11190 0.0380882
R35270 DVDD.n13882 DVDD.n11190 0.0380882
R35271 DVDD.n13884 DVDD.n13882 0.0380882
R35272 DVDD.n13886 DVDD.n13884 0.0380882
R35273 DVDD.n13886 DVDD.n11187 0.0380882
R35274 DVDD.n13891 DVDD.n11187 0.0380882
R35275 DVDD.n13893 DVDD.n13891 0.0380882
R35276 DVDD.n13895 DVDD.n13893 0.0380882
R35277 DVDD.n13895 DVDD.n11184 0.0380882
R35278 DVDD.n13900 DVDD.n11184 0.0380882
R35279 DVDD.n13902 DVDD.n13900 0.0380882
R35280 DVDD.n13904 DVDD.n13902 0.0380882
R35281 DVDD.n13904 DVDD.n11181 0.0380882
R35282 DVDD.n13909 DVDD.n11181 0.0380882
R35283 DVDD.n13911 DVDD.n13909 0.0380882
R35284 DVDD.n13913 DVDD.n13911 0.0380882
R35285 DVDD.n13913 DVDD.n11178 0.0380882
R35286 DVDD.n13918 DVDD.n11178 0.0380882
R35287 DVDD.n13920 DVDD.n13918 0.0380882
R35288 DVDD.n13922 DVDD.n13920 0.0380882
R35289 DVDD.n13922 DVDD.n11175 0.0380882
R35290 DVDD.n13927 DVDD.n11175 0.0380882
R35291 DVDD.n13929 DVDD.n13927 0.0380882
R35292 DVDD.n13931 DVDD.n13929 0.0380882
R35293 DVDD.n13931 DVDD.n11172 0.0380882
R35294 DVDD.n13936 DVDD.n11172 0.0380882
R35295 DVDD.n13938 DVDD.n13936 0.0380882
R35296 DVDD.n13940 DVDD.n13938 0.0380882
R35297 DVDD.n13940 DVDD.n11169 0.0380882
R35298 DVDD.n13945 DVDD.n11169 0.0380882
R35299 DVDD.n13947 DVDD.n13945 0.0380882
R35300 DVDD.n13949 DVDD.n13947 0.0380882
R35301 DVDD.n13949 DVDD.n11166 0.0380882
R35302 DVDD.n13954 DVDD.n11166 0.0380882
R35303 DVDD.n13956 DVDD.n13954 0.0380882
R35304 DVDD.n13958 DVDD.n13956 0.0380882
R35305 DVDD.n13958 DVDD.n11163 0.0380882
R35306 DVDD.n13963 DVDD.n11163 0.0380882
R35307 DVDD.n13965 DVDD.n13963 0.0380882
R35308 DVDD.n13967 DVDD.n13965 0.0380882
R35309 DVDD.n13967 DVDD.n11160 0.0380882
R35310 DVDD.n13972 DVDD.n11160 0.0380882
R35311 DVDD.n13974 DVDD.n13972 0.0380882
R35312 DVDD.n13976 DVDD.n13974 0.0380882
R35313 DVDD.n13976 DVDD.n11157 0.0380882
R35314 DVDD.n13981 DVDD.n11157 0.0380882
R35315 DVDD.n13983 DVDD.n13981 0.0380882
R35316 DVDD.n13985 DVDD.n13983 0.0380882
R35317 DVDD.n13985 DVDD.n11154 0.0380882
R35318 DVDD.n13990 DVDD.n11154 0.0380882
R35319 DVDD.n13992 DVDD.n13990 0.0380882
R35320 DVDD.n13994 DVDD.n13992 0.0380882
R35321 DVDD.n13994 DVDD.n11151 0.0380882
R35322 DVDD.n13998 DVDD.n11151 0.0380882
R35323 DVDD.n11324 DVDD.n11229 0.0380882
R35324 DVDD.n11325 DVDD.n11324 0.0380882
R35325 DVDD.n11325 DVDD.n11319 0.0380882
R35326 DVDD.n11335 DVDD.n11319 0.0380882
R35327 DVDD.n11336 DVDD.n11335 0.0380882
R35328 DVDD.n11337 DVDD.n11336 0.0380882
R35329 DVDD.n11337 DVDD.n11317 0.0380882
R35330 DVDD.n11347 DVDD.n11317 0.0380882
R35331 DVDD.n11348 DVDD.n11347 0.0380882
R35332 DVDD.n11349 DVDD.n11348 0.0380882
R35333 DVDD.n11349 DVDD.n11315 0.0380882
R35334 DVDD.n11359 DVDD.n11315 0.0380882
R35335 DVDD.n11360 DVDD.n11359 0.0380882
R35336 DVDD.n11361 DVDD.n11360 0.0380882
R35337 DVDD.n11361 DVDD.n11313 0.0380882
R35338 DVDD.n11371 DVDD.n11313 0.0380882
R35339 DVDD.n11372 DVDD.n11371 0.0380882
R35340 DVDD.n11373 DVDD.n11372 0.0380882
R35341 DVDD.n11373 DVDD.n11311 0.0380882
R35342 DVDD.n11383 DVDD.n11311 0.0380882
R35343 DVDD.n11384 DVDD.n11383 0.0380882
R35344 DVDD.n11385 DVDD.n11384 0.0380882
R35345 DVDD.n11385 DVDD.n11309 0.0380882
R35346 DVDD.n11395 DVDD.n11309 0.0380882
R35347 DVDD.n11396 DVDD.n11395 0.0380882
R35348 DVDD.n11397 DVDD.n11396 0.0380882
R35349 DVDD.n11397 DVDD.n11307 0.0380882
R35350 DVDD.n11407 DVDD.n11307 0.0380882
R35351 DVDD.n11408 DVDD.n11407 0.0380882
R35352 DVDD.n11409 DVDD.n11408 0.0380882
R35353 DVDD.n11409 DVDD.n11305 0.0380882
R35354 DVDD.n11419 DVDD.n11305 0.0380882
R35355 DVDD.n11420 DVDD.n11419 0.0380882
R35356 DVDD.n11421 DVDD.n11420 0.0380882
R35357 DVDD.n11421 DVDD.n11303 0.0380882
R35358 DVDD.n11431 DVDD.n11303 0.0380882
R35359 DVDD.n11432 DVDD.n11431 0.0380882
R35360 DVDD.n11433 DVDD.n11432 0.0380882
R35361 DVDD.n11433 DVDD.n11301 0.0380882
R35362 DVDD.n11443 DVDD.n11301 0.0380882
R35363 DVDD.n11444 DVDD.n11443 0.0380882
R35364 DVDD.n11445 DVDD.n11444 0.0380882
R35365 DVDD.n11445 DVDD.n11299 0.0380882
R35366 DVDD.n11455 DVDD.n11299 0.0380882
R35367 DVDD.n11456 DVDD.n11455 0.0380882
R35368 DVDD.n11457 DVDD.n11456 0.0380882
R35369 DVDD.n11457 DVDD.n11297 0.0380882
R35370 DVDD.n11467 DVDD.n11297 0.0380882
R35371 DVDD.n11468 DVDD.n11467 0.0380882
R35372 DVDD.n11469 DVDD.n11468 0.0380882
R35373 DVDD.n11469 DVDD.n11295 0.0380882
R35374 DVDD.n11479 DVDD.n11295 0.0380882
R35375 DVDD.n11480 DVDD.n11479 0.0380882
R35376 DVDD.n11481 DVDD.n11480 0.0380882
R35377 DVDD.n11481 DVDD.n11293 0.0380882
R35378 DVDD.n11491 DVDD.n11293 0.0380882
R35379 DVDD.n11492 DVDD.n11491 0.0380882
R35380 DVDD.n11493 DVDD.n11492 0.0380882
R35381 DVDD.n11493 DVDD.n11291 0.0380882
R35382 DVDD.n11503 DVDD.n11291 0.0380882
R35383 DVDD.n11504 DVDD.n11503 0.0380882
R35384 DVDD.n11505 DVDD.n11504 0.0380882
R35385 DVDD.n11505 DVDD.n11289 0.0380882
R35386 DVDD.n11515 DVDD.n11289 0.0380882
R35387 DVDD.n11516 DVDD.n11515 0.0380882
R35388 DVDD.n11517 DVDD.n11516 0.0380882
R35389 DVDD.n11517 DVDD.n11287 0.0380882
R35390 DVDD.n11527 DVDD.n11287 0.0380882
R35391 DVDD.n11528 DVDD.n11527 0.0380882
R35392 DVDD.n11529 DVDD.n11528 0.0380882
R35393 DVDD.n11529 DVDD.n11285 0.0380882
R35394 DVDD.n11539 DVDD.n11285 0.0380882
R35395 DVDD.n11540 DVDD.n11539 0.0380882
R35396 DVDD.n11541 DVDD.n11540 0.0380882
R35397 DVDD.n11541 DVDD.n11283 0.0380882
R35398 DVDD.n11551 DVDD.n11283 0.0380882
R35399 DVDD.n11552 DVDD.n11551 0.0380882
R35400 DVDD.n11553 DVDD.n11552 0.0380882
R35401 DVDD.n11553 DVDD.n11281 0.0380882
R35402 DVDD.n11563 DVDD.n11281 0.0380882
R35403 DVDD.n11564 DVDD.n11563 0.0380882
R35404 DVDD.n13794 DVDD.n11564 0.0380882
R35405 DVDD.n13794 DVDD.n13793 0.0380882
R35406 DVDD.n11323 DVDD.n11320 0.0380882
R35407 DVDD.n11326 DVDD.n11323 0.0380882
R35408 DVDD.n11330 DVDD.n11326 0.0380882
R35409 DVDD.n11334 DVDD.n11330 0.0380882
R35410 DVDD.n11334 DVDD.n11318 0.0380882
R35411 DVDD.n11338 DVDD.n11318 0.0380882
R35412 DVDD.n11342 DVDD.n11338 0.0380882
R35413 DVDD.n11346 DVDD.n11342 0.0380882
R35414 DVDD.n11346 DVDD.n11316 0.0380882
R35415 DVDD.n11350 DVDD.n11316 0.0380882
R35416 DVDD.n11354 DVDD.n11350 0.0380882
R35417 DVDD.n11358 DVDD.n11354 0.0380882
R35418 DVDD.n11358 DVDD.n11314 0.0380882
R35419 DVDD.n11362 DVDD.n11314 0.0380882
R35420 DVDD.n11366 DVDD.n11362 0.0380882
R35421 DVDD.n11370 DVDD.n11366 0.0380882
R35422 DVDD.n11370 DVDD.n11312 0.0380882
R35423 DVDD.n11374 DVDD.n11312 0.0380882
R35424 DVDD.n11378 DVDD.n11374 0.0380882
R35425 DVDD.n11382 DVDD.n11378 0.0380882
R35426 DVDD.n11382 DVDD.n11310 0.0380882
R35427 DVDD.n11386 DVDD.n11310 0.0380882
R35428 DVDD.n11390 DVDD.n11386 0.0380882
R35429 DVDD.n11394 DVDD.n11390 0.0380882
R35430 DVDD.n11394 DVDD.n11308 0.0380882
R35431 DVDD.n11398 DVDD.n11308 0.0380882
R35432 DVDD.n11402 DVDD.n11398 0.0380882
R35433 DVDD.n11406 DVDD.n11402 0.0380882
R35434 DVDD.n11406 DVDD.n11306 0.0380882
R35435 DVDD.n11410 DVDD.n11306 0.0380882
R35436 DVDD.n11414 DVDD.n11410 0.0380882
R35437 DVDD.n11418 DVDD.n11414 0.0380882
R35438 DVDD.n11418 DVDD.n11304 0.0380882
R35439 DVDD.n11422 DVDD.n11304 0.0380882
R35440 DVDD.n11426 DVDD.n11422 0.0380882
R35441 DVDD.n11430 DVDD.n11426 0.0380882
R35442 DVDD.n11430 DVDD.n11302 0.0380882
R35443 DVDD.n11434 DVDD.n11302 0.0380882
R35444 DVDD.n11438 DVDD.n11434 0.0380882
R35445 DVDD.n11442 DVDD.n11438 0.0380882
R35446 DVDD.n11442 DVDD.n11300 0.0380882
R35447 DVDD.n11446 DVDD.n11300 0.0380882
R35448 DVDD.n11450 DVDD.n11446 0.0380882
R35449 DVDD.n11454 DVDD.n11450 0.0380882
R35450 DVDD.n11454 DVDD.n11298 0.0380882
R35451 DVDD.n11458 DVDD.n11298 0.0380882
R35452 DVDD.n11462 DVDD.n11458 0.0380882
R35453 DVDD.n11466 DVDD.n11462 0.0380882
R35454 DVDD.n11466 DVDD.n11296 0.0380882
R35455 DVDD.n11470 DVDD.n11296 0.0380882
R35456 DVDD.n11474 DVDD.n11470 0.0380882
R35457 DVDD.n11478 DVDD.n11474 0.0380882
R35458 DVDD.n11478 DVDD.n11294 0.0380882
R35459 DVDD.n11482 DVDD.n11294 0.0380882
R35460 DVDD.n11486 DVDD.n11482 0.0380882
R35461 DVDD.n11490 DVDD.n11486 0.0380882
R35462 DVDD.n11490 DVDD.n11292 0.0380882
R35463 DVDD.n11494 DVDD.n11292 0.0380882
R35464 DVDD.n11498 DVDD.n11494 0.0380882
R35465 DVDD.n11502 DVDD.n11498 0.0380882
R35466 DVDD.n11502 DVDD.n11290 0.0380882
R35467 DVDD.n11506 DVDD.n11290 0.0380882
R35468 DVDD.n11510 DVDD.n11506 0.0380882
R35469 DVDD.n11514 DVDD.n11510 0.0380882
R35470 DVDD.n11514 DVDD.n11288 0.0380882
R35471 DVDD.n11518 DVDD.n11288 0.0380882
R35472 DVDD.n11522 DVDD.n11518 0.0380882
R35473 DVDD.n11526 DVDD.n11522 0.0380882
R35474 DVDD.n11526 DVDD.n11286 0.0380882
R35475 DVDD.n11530 DVDD.n11286 0.0380882
R35476 DVDD.n11534 DVDD.n11530 0.0380882
R35477 DVDD.n11538 DVDD.n11534 0.0380882
R35478 DVDD.n11538 DVDD.n11284 0.0380882
R35479 DVDD.n11542 DVDD.n11284 0.0380882
R35480 DVDD.n11546 DVDD.n11542 0.0380882
R35481 DVDD.n11550 DVDD.n11546 0.0380882
R35482 DVDD.n11550 DVDD.n11282 0.0380882
R35483 DVDD.n11554 DVDD.n11282 0.0380882
R35484 DVDD.n11558 DVDD.n11554 0.0380882
R35485 DVDD.n11562 DVDD.n11558 0.0380882
R35486 DVDD.n11562 DVDD.n11280 0.0380882
R35487 DVDD.n13795 DVDD.n11280 0.0380882
R35488 DVDD.n13795 DVDD.n11278 0.0380882
R35489 DVDD.n11678 DVDD.n11584 0.0380882
R35490 DVDD.n11679 DVDD.n11678 0.0380882
R35491 DVDD.n11679 DVDD.n11673 0.0380882
R35492 DVDD.n11689 DVDD.n11673 0.0380882
R35493 DVDD.n11690 DVDD.n11689 0.0380882
R35494 DVDD.n11691 DVDD.n11690 0.0380882
R35495 DVDD.n11691 DVDD.n11671 0.0380882
R35496 DVDD.n11701 DVDD.n11671 0.0380882
R35497 DVDD.n11702 DVDD.n11701 0.0380882
R35498 DVDD.n11703 DVDD.n11702 0.0380882
R35499 DVDD.n11703 DVDD.n11669 0.0380882
R35500 DVDD.n11713 DVDD.n11669 0.0380882
R35501 DVDD.n11714 DVDD.n11713 0.0380882
R35502 DVDD.n11715 DVDD.n11714 0.0380882
R35503 DVDD.n11715 DVDD.n11667 0.0380882
R35504 DVDD.n11725 DVDD.n11667 0.0380882
R35505 DVDD.n11726 DVDD.n11725 0.0380882
R35506 DVDD.n11727 DVDD.n11726 0.0380882
R35507 DVDD.n11727 DVDD.n11665 0.0380882
R35508 DVDD.n11737 DVDD.n11665 0.0380882
R35509 DVDD.n11738 DVDD.n11737 0.0380882
R35510 DVDD.n11739 DVDD.n11738 0.0380882
R35511 DVDD.n11739 DVDD.n11663 0.0380882
R35512 DVDD.n11749 DVDD.n11663 0.0380882
R35513 DVDD.n11750 DVDD.n11749 0.0380882
R35514 DVDD.n11751 DVDD.n11750 0.0380882
R35515 DVDD.n11751 DVDD.n11661 0.0380882
R35516 DVDD.n11761 DVDD.n11661 0.0380882
R35517 DVDD.n11762 DVDD.n11761 0.0380882
R35518 DVDD.n11763 DVDD.n11762 0.0380882
R35519 DVDD.n11763 DVDD.n11659 0.0380882
R35520 DVDD.n11773 DVDD.n11659 0.0380882
R35521 DVDD.n11774 DVDD.n11773 0.0380882
R35522 DVDD.n11775 DVDD.n11774 0.0380882
R35523 DVDD.n11775 DVDD.n11657 0.0380882
R35524 DVDD.n11785 DVDD.n11657 0.0380882
R35525 DVDD.n11786 DVDD.n11785 0.0380882
R35526 DVDD.n11787 DVDD.n11786 0.0380882
R35527 DVDD.n11787 DVDD.n11655 0.0380882
R35528 DVDD.n11797 DVDD.n11655 0.0380882
R35529 DVDD.n11798 DVDD.n11797 0.0380882
R35530 DVDD.n11799 DVDD.n11798 0.0380882
R35531 DVDD.n11799 DVDD.n11653 0.0380882
R35532 DVDD.n11809 DVDD.n11653 0.0380882
R35533 DVDD.n11810 DVDD.n11809 0.0380882
R35534 DVDD.n11811 DVDD.n11810 0.0380882
R35535 DVDD.n11811 DVDD.n11651 0.0380882
R35536 DVDD.n11821 DVDD.n11651 0.0380882
R35537 DVDD.n11822 DVDD.n11821 0.0380882
R35538 DVDD.n11823 DVDD.n11822 0.0380882
R35539 DVDD.n11823 DVDD.n11649 0.0380882
R35540 DVDD.n11833 DVDD.n11649 0.0380882
R35541 DVDD.n11834 DVDD.n11833 0.0380882
R35542 DVDD.n11835 DVDD.n11834 0.0380882
R35543 DVDD.n11835 DVDD.n11647 0.0380882
R35544 DVDD.n11845 DVDD.n11647 0.0380882
R35545 DVDD.n11846 DVDD.n11845 0.0380882
R35546 DVDD.n11847 DVDD.n11846 0.0380882
R35547 DVDD.n11847 DVDD.n11645 0.0380882
R35548 DVDD.n11857 DVDD.n11645 0.0380882
R35549 DVDD.n11858 DVDD.n11857 0.0380882
R35550 DVDD.n11859 DVDD.n11858 0.0380882
R35551 DVDD.n11859 DVDD.n11643 0.0380882
R35552 DVDD.n11869 DVDD.n11643 0.0380882
R35553 DVDD.n11870 DVDD.n11869 0.0380882
R35554 DVDD.n11871 DVDD.n11870 0.0380882
R35555 DVDD.n11871 DVDD.n11641 0.0380882
R35556 DVDD.n11881 DVDD.n11641 0.0380882
R35557 DVDD.n11882 DVDD.n11881 0.0380882
R35558 DVDD.n11883 DVDD.n11882 0.0380882
R35559 DVDD.n11883 DVDD.n11639 0.0380882
R35560 DVDD.n11893 DVDD.n11639 0.0380882
R35561 DVDD.n11894 DVDD.n11893 0.0380882
R35562 DVDD.n11895 DVDD.n11894 0.0380882
R35563 DVDD.n11895 DVDD.n11637 0.0380882
R35564 DVDD.n11905 DVDD.n11637 0.0380882
R35565 DVDD.n11906 DVDD.n11905 0.0380882
R35566 DVDD.n11907 DVDD.n11906 0.0380882
R35567 DVDD.n11907 DVDD.n11635 0.0380882
R35568 DVDD.n11917 DVDD.n11635 0.0380882
R35569 DVDD.n11918 DVDD.n11917 0.0380882
R35570 DVDD.n13772 DVDD.n11918 0.0380882
R35571 DVDD.n13772 DVDD.n13771 0.0380882
R35572 DVDD.n11677 DVDD.n11674 0.0380882
R35573 DVDD.n11680 DVDD.n11677 0.0380882
R35574 DVDD.n11684 DVDD.n11680 0.0380882
R35575 DVDD.n11688 DVDD.n11684 0.0380882
R35576 DVDD.n11688 DVDD.n11672 0.0380882
R35577 DVDD.n11692 DVDD.n11672 0.0380882
R35578 DVDD.n11696 DVDD.n11692 0.0380882
R35579 DVDD.n11700 DVDD.n11696 0.0380882
R35580 DVDD.n11700 DVDD.n11670 0.0380882
R35581 DVDD.n11704 DVDD.n11670 0.0380882
R35582 DVDD.n11708 DVDD.n11704 0.0380882
R35583 DVDD.n11712 DVDD.n11708 0.0380882
R35584 DVDD.n11712 DVDD.n11668 0.0380882
R35585 DVDD.n11716 DVDD.n11668 0.0380882
R35586 DVDD.n11720 DVDD.n11716 0.0380882
R35587 DVDD.n11724 DVDD.n11720 0.0380882
R35588 DVDD.n11724 DVDD.n11666 0.0380882
R35589 DVDD.n11728 DVDD.n11666 0.0380882
R35590 DVDD.n11732 DVDD.n11728 0.0380882
R35591 DVDD.n11736 DVDD.n11732 0.0380882
R35592 DVDD.n11736 DVDD.n11664 0.0380882
R35593 DVDD.n11740 DVDD.n11664 0.0380882
R35594 DVDD.n11744 DVDD.n11740 0.0380882
R35595 DVDD.n11748 DVDD.n11744 0.0380882
R35596 DVDD.n11748 DVDD.n11662 0.0380882
R35597 DVDD.n11752 DVDD.n11662 0.0380882
R35598 DVDD.n11756 DVDD.n11752 0.0380882
R35599 DVDD.n11760 DVDD.n11756 0.0380882
R35600 DVDD.n11760 DVDD.n11660 0.0380882
R35601 DVDD.n11764 DVDD.n11660 0.0380882
R35602 DVDD.n11768 DVDD.n11764 0.0380882
R35603 DVDD.n11772 DVDD.n11768 0.0380882
R35604 DVDD.n11772 DVDD.n11658 0.0380882
R35605 DVDD.n11776 DVDD.n11658 0.0380882
R35606 DVDD.n11780 DVDD.n11776 0.0380882
R35607 DVDD.n11784 DVDD.n11780 0.0380882
R35608 DVDD.n11784 DVDD.n11656 0.0380882
R35609 DVDD.n11788 DVDD.n11656 0.0380882
R35610 DVDD.n11792 DVDD.n11788 0.0380882
R35611 DVDD.n11796 DVDD.n11792 0.0380882
R35612 DVDD.n11796 DVDD.n11654 0.0380882
R35613 DVDD.n11800 DVDD.n11654 0.0380882
R35614 DVDD.n11804 DVDD.n11800 0.0380882
R35615 DVDD.n11808 DVDD.n11804 0.0380882
R35616 DVDD.n11808 DVDD.n11652 0.0380882
R35617 DVDD.n11812 DVDD.n11652 0.0380882
R35618 DVDD.n11816 DVDD.n11812 0.0380882
R35619 DVDD.n11820 DVDD.n11816 0.0380882
R35620 DVDD.n11820 DVDD.n11650 0.0380882
R35621 DVDD.n11824 DVDD.n11650 0.0380882
R35622 DVDD.n11828 DVDD.n11824 0.0380882
R35623 DVDD.n11832 DVDD.n11828 0.0380882
R35624 DVDD.n11832 DVDD.n11648 0.0380882
R35625 DVDD.n11836 DVDD.n11648 0.0380882
R35626 DVDD.n11840 DVDD.n11836 0.0380882
R35627 DVDD.n11844 DVDD.n11840 0.0380882
R35628 DVDD.n11844 DVDD.n11646 0.0380882
R35629 DVDD.n11848 DVDD.n11646 0.0380882
R35630 DVDD.n11852 DVDD.n11848 0.0380882
R35631 DVDD.n11856 DVDD.n11852 0.0380882
R35632 DVDD.n11856 DVDD.n11644 0.0380882
R35633 DVDD.n11860 DVDD.n11644 0.0380882
R35634 DVDD.n11864 DVDD.n11860 0.0380882
R35635 DVDD.n11868 DVDD.n11864 0.0380882
R35636 DVDD.n11868 DVDD.n11642 0.0380882
R35637 DVDD.n11872 DVDD.n11642 0.0380882
R35638 DVDD.n11876 DVDD.n11872 0.0380882
R35639 DVDD.n11880 DVDD.n11876 0.0380882
R35640 DVDD.n11880 DVDD.n11640 0.0380882
R35641 DVDD.n11884 DVDD.n11640 0.0380882
R35642 DVDD.n11888 DVDD.n11884 0.0380882
R35643 DVDD.n11892 DVDD.n11888 0.0380882
R35644 DVDD.n11892 DVDD.n11638 0.0380882
R35645 DVDD.n11896 DVDD.n11638 0.0380882
R35646 DVDD.n11900 DVDD.n11896 0.0380882
R35647 DVDD.n11904 DVDD.n11900 0.0380882
R35648 DVDD.n11904 DVDD.n11636 0.0380882
R35649 DVDD.n11908 DVDD.n11636 0.0380882
R35650 DVDD.n11912 DVDD.n11908 0.0380882
R35651 DVDD.n11916 DVDD.n11912 0.0380882
R35652 DVDD.n11916 DVDD.n11634 0.0380882
R35653 DVDD.n13773 DVDD.n11634 0.0380882
R35654 DVDD.n13773 DVDD.n11633 0.0380882
R35655 DVDD.n12025 DVDD.n11930 0.0380882
R35656 DVDD.n12036 DVDD.n12025 0.0380882
R35657 DVDD.n12037 DVDD.n12036 0.0380882
R35658 DVDD.n12038 DVDD.n12037 0.0380882
R35659 DVDD.n12038 DVDD.n12021 0.0380882
R35660 DVDD.n12048 DVDD.n12021 0.0380882
R35661 DVDD.n12049 DVDD.n12048 0.0380882
R35662 DVDD.n12050 DVDD.n12049 0.0380882
R35663 DVDD.n12050 DVDD.n12017 0.0380882
R35664 DVDD.n12060 DVDD.n12017 0.0380882
R35665 DVDD.n12061 DVDD.n12060 0.0380882
R35666 DVDD.n12062 DVDD.n12061 0.0380882
R35667 DVDD.n12062 DVDD.n12013 0.0380882
R35668 DVDD.n12072 DVDD.n12013 0.0380882
R35669 DVDD.n12073 DVDD.n12072 0.0380882
R35670 DVDD.n12074 DVDD.n12073 0.0380882
R35671 DVDD.n12074 DVDD.n12009 0.0380882
R35672 DVDD.n12084 DVDD.n12009 0.0380882
R35673 DVDD.n12085 DVDD.n12084 0.0380882
R35674 DVDD.n12086 DVDD.n12085 0.0380882
R35675 DVDD.n12086 DVDD.n12005 0.0380882
R35676 DVDD.n12096 DVDD.n12005 0.0380882
R35677 DVDD.n12097 DVDD.n12096 0.0380882
R35678 DVDD.n12098 DVDD.n12097 0.0380882
R35679 DVDD.n12098 DVDD.n12001 0.0380882
R35680 DVDD.n12108 DVDD.n12001 0.0380882
R35681 DVDD.n12109 DVDD.n12108 0.0380882
R35682 DVDD.n12110 DVDD.n12109 0.0380882
R35683 DVDD.n12110 DVDD.n11997 0.0380882
R35684 DVDD.n12120 DVDD.n11997 0.0380882
R35685 DVDD.n12121 DVDD.n12120 0.0380882
R35686 DVDD.n12122 DVDD.n12121 0.0380882
R35687 DVDD.n12122 DVDD.n11993 0.0380882
R35688 DVDD.n12132 DVDD.n11993 0.0380882
R35689 DVDD.n12133 DVDD.n12132 0.0380882
R35690 DVDD.n12134 DVDD.n12133 0.0380882
R35691 DVDD.n12134 DVDD.n11989 0.0380882
R35692 DVDD.n12144 DVDD.n11989 0.0380882
R35693 DVDD.n12145 DVDD.n12144 0.0380882
R35694 DVDD.n12146 DVDD.n12145 0.0380882
R35695 DVDD.n12146 DVDD.n11985 0.0380882
R35696 DVDD.n12156 DVDD.n11985 0.0380882
R35697 DVDD.n12157 DVDD.n12156 0.0380882
R35698 DVDD.n12158 DVDD.n12157 0.0380882
R35699 DVDD.n12158 DVDD.n11981 0.0380882
R35700 DVDD.n12168 DVDD.n11981 0.0380882
R35701 DVDD.n12169 DVDD.n12168 0.0380882
R35702 DVDD.n12170 DVDD.n12169 0.0380882
R35703 DVDD.n12170 DVDD.n11977 0.0380882
R35704 DVDD.n12180 DVDD.n11977 0.0380882
R35705 DVDD.n12181 DVDD.n12180 0.0380882
R35706 DVDD.n12182 DVDD.n12181 0.0380882
R35707 DVDD.n12182 DVDD.n11973 0.0380882
R35708 DVDD.n12192 DVDD.n11973 0.0380882
R35709 DVDD.n12193 DVDD.n12192 0.0380882
R35710 DVDD.n12194 DVDD.n12193 0.0380882
R35711 DVDD.n12194 DVDD.n11969 0.0380882
R35712 DVDD.n12204 DVDD.n11969 0.0380882
R35713 DVDD.n12205 DVDD.n12204 0.0380882
R35714 DVDD.n12206 DVDD.n12205 0.0380882
R35715 DVDD.n12206 DVDD.n11965 0.0380882
R35716 DVDD.n12216 DVDD.n11965 0.0380882
R35717 DVDD.n12217 DVDD.n12216 0.0380882
R35718 DVDD.n12218 DVDD.n12217 0.0380882
R35719 DVDD.n12218 DVDD.n11961 0.0380882
R35720 DVDD.n12228 DVDD.n11961 0.0380882
R35721 DVDD.n12229 DVDD.n12228 0.0380882
R35722 DVDD.n12230 DVDD.n12229 0.0380882
R35723 DVDD.n12230 DVDD.n11957 0.0380882
R35724 DVDD.n12240 DVDD.n11957 0.0380882
R35725 DVDD.n12241 DVDD.n12240 0.0380882
R35726 DVDD.n12242 DVDD.n12241 0.0380882
R35727 DVDD.n12242 DVDD.n11953 0.0380882
R35728 DVDD.n12252 DVDD.n11953 0.0380882
R35729 DVDD.n12253 DVDD.n12252 0.0380882
R35730 DVDD.n12254 DVDD.n12253 0.0380882
R35731 DVDD.n12254 DVDD.n11949 0.0380882
R35732 DVDD.n12264 DVDD.n11949 0.0380882
R35733 DVDD.n12265 DVDD.n12264 0.0380882
R35734 DVDD.n12267 DVDD.n12265 0.0380882
R35735 DVDD.n12267 DVDD.n12266 0.0380882
R35736 DVDD.n12266 DVDD.n11944 0.0380882
R35737 DVDD.n12277 DVDD.n11944 0.0380882
R35738 DVDD.n12027 DVDD.n12026 0.0380882
R35739 DVDD.n12035 DVDD.n12026 0.0380882
R35740 DVDD.n12035 DVDD.n12024 0.0380882
R35741 DVDD.n12039 DVDD.n12024 0.0380882
R35742 DVDD.n12039 DVDD.n12022 0.0380882
R35743 DVDD.n12047 DVDD.n12022 0.0380882
R35744 DVDD.n12047 DVDD.n12020 0.0380882
R35745 DVDD.n12051 DVDD.n12020 0.0380882
R35746 DVDD.n12051 DVDD.n12018 0.0380882
R35747 DVDD.n12059 DVDD.n12018 0.0380882
R35748 DVDD.n12059 DVDD.n12016 0.0380882
R35749 DVDD.n12063 DVDD.n12016 0.0380882
R35750 DVDD.n12063 DVDD.n12014 0.0380882
R35751 DVDD.n12071 DVDD.n12014 0.0380882
R35752 DVDD.n12071 DVDD.n12012 0.0380882
R35753 DVDD.n12075 DVDD.n12012 0.0380882
R35754 DVDD.n12075 DVDD.n12010 0.0380882
R35755 DVDD.n12083 DVDD.n12010 0.0380882
R35756 DVDD.n12083 DVDD.n12008 0.0380882
R35757 DVDD.n12087 DVDD.n12008 0.0380882
R35758 DVDD.n12087 DVDD.n12006 0.0380882
R35759 DVDD.n12095 DVDD.n12006 0.0380882
R35760 DVDD.n12095 DVDD.n12004 0.0380882
R35761 DVDD.n12099 DVDD.n12004 0.0380882
R35762 DVDD.n12099 DVDD.n12002 0.0380882
R35763 DVDD.n12107 DVDD.n12002 0.0380882
R35764 DVDD.n12107 DVDD.n12000 0.0380882
R35765 DVDD.n12111 DVDD.n12000 0.0380882
R35766 DVDD.n12111 DVDD.n11998 0.0380882
R35767 DVDD.n12119 DVDD.n11998 0.0380882
R35768 DVDD.n12119 DVDD.n11996 0.0380882
R35769 DVDD.n12123 DVDD.n11996 0.0380882
R35770 DVDD.n12123 DVDD.n11994 0.0380882
R35771 DVDD.n12131 DVDD.n11994 0.0380882
R35772 DVDD.n12131 DVDD.n11992 0.0380882
R35773 DVDD.n12135 DVDD.n11992 0.0380882
R35774 DVDD.n12135 DVDD.n11990 0.0380882
R35775 DVDD.n12143 DVDD.n11990 0.0380882
R35776 DVDD.n12143 DVDD.n11988 0.0380882
R35777 DVDD.n12147 DVDD.n11988 0.0380882
R35778 DVDD.n12147 DVDD.n11986 0.0380882
R35779 DVDD.n12155 DVDD.n11986 0.0380882
R35780 DVDD.n12155 DVDD.n11984 0.0380882
R35781 DVDD.n12159 DVDD.n11984 0.0380882
R35782 DVDD.n12159 DVDD.n11982 0.0380882
R35783 DVDD.n12167 DVDD.n11982 0.0380882
R35784 DVDD.n12167 DVDD.n11980 0.0380882
R35785 DVDD.n12171 DVDD.n11980 0.0380882
R35786 DVDD.n12171 DVDD.n11978 0.0380882
R35787 DVDD.n12179 DVDD.n11978 0.0380882
R35788 DVDD.n12179 DVDD.n11976 0.0380882
R35789 DVDD.n12183 DVDD.n11976 0.0380882
R35790 DVDD.n12183 DVDD.n11974 0.0380882
R35791 DVDD.n12191 DVDD.n11974 0.0380882
R35792 DVDD.n12191 DVDD.n11972 0.0380882
R35793 DVDD.n12195 DVDD.n11972 0.0380882
R35794 DVDD.n12195 DVDD.n11970 0.0380882
R35795 DVDD.n12203 DVDD.n11970 0.0380882
R35796 DVDD.n12203 DVDD.n11968 0.0380882
R35797 DVDD.n12207 DVDD.n11968 0.0380882
R35798 DVDD.n12207 DVDD.n11966 0.0380882
R35799 DVDD.n12215 DVDD.n11966 0.0380882
R35800 DVDD.n12215 DVDD.n11964 0.0380882
R35801 DVDD.n12219 DVDD.n11964 0.0380882
R35802 DVDD.n12219 DVDD.n11962 0.0380882
R35803 DVDD.n12227 DVDD.n11962 0.0380882
R35804 DVDD.n12227 DVDD.n11960 0.0380882
R35805 DVDD.n12231 DVDD.n11960 0.0380882
R35806 DVDD.n12231 DVDD.n11958 0.0380882
R35807 DVDD.n12239 DVDD.n11958 0.0380882
R35808 DVDD.n12239 DVDD.n11956 0.0380882
R35809 DVDD.n12243 DVDD.n11956 0.0380882
R35810 DVDD.n12243 DVDD.n11954 0.0380882
R35811 DVDD.n12251 DVDD.n11954 0.0380882
R35812 DVDD.n12251 DVDD.n11952 0.0380882
R35813 DVDD.n12255 DVDD.n11952 0.0380882
R35814 DVDD.n12255 DVDD.n11950 0.0380882
R35815 DVDD.n12263 DVDD.n11950 0.0380882
R35816 DVDD.n12263 DVDD.n11948 0.0380882
R35817 DVDD.n12268 DVDD.n11948 0.0380882
R35818 DVDD.n12268 DVDD.n11946 0.0380882
R35819 DVDD.n11946 DVDD.n11945 0.0380882
R35820 DVDD.n12276 DVDD.n11945 0.0380882
R35821 DVDD.n13498 DVDD.n13497 0.0380882
R35822 DVDD.n13499 DVDD.n13498 0.0380882
R35823 DVDD.n13499 DVDD.n12373 0.0380882
R35824 DVDD.n13509 DVDD.n12373 0.0380882
R35825 DVDD.n13510 DVDD.n13509 0.0380882
R35826 DVDD.n13511 DVDD.n13510 0.0380882
R35827 DVDD.n13511 DVDD.n12371 0.0380882
R35828 DVDD.n13521 DVDD.n12371 0.0380882
R35829 DVDD.n13522 DVDD.n13521 0.0380882
R35830 DVDD.n13523 DVDD.n13522 0.0380882
R35831 DVDD.n13523 DVDD.n12369 0.0380882
R35832 DVDD.n13533 DVDD.n12369 0.0380882
R35833 DVDD.n13534 DVDD.n13533 0.0380882
R35834 DVDD.n13535 DVDD.n13534 0.0380882
R35835 DVDD.n13535 DVDD.n12367 0.0380882
R35836 DVDD.n13545 DVDD.n12367 0.0380882
R35837 DVDD.n13546 DVDD.n13545 0.0380882
R35838 DVDD.n13547 DVDD.n13546 0.0380882
R35839 DVDD.n13547 DVDD.n12365 0.0380882
R35840 DVDD.n13557 DVDD.n12365 0.0380882
R35841 DVDD.n13558 DVDD.n13557 0.0380882
R35842 DVDD.n13559 DVDD.n13558 0.0380882
R35843 DVDD.n13559 DVDD.n12363 0.0380882
R35844 DVDD.n13569 DVDD.n12363 0.0380882
R35845 DVDD.n13570 DVDD.n13569 0.0380882
R35846 DVDD.n13571 DVDD.n13570 0.0380882
R35847 DVDD.n13571 DVDD.n12361 0.0380882
R35848 DVDD.n13581 DVDD.n12361 0.0380882
R35849 DVDD.n13582 DVDD.n13581 0.0380882
R35850 DVDD.n13583 DVDD.n13582 0.0380882
R35851 DVDD.n13583 DVDD.n12359 0.0380882
R35852 DVDD.n13593 DVDD.n12359 0.0380882
R35853 DVDD.n13594 DVDD.n13593 0.0380882
R35854 DVDD.n13595 DVDD.n13594 0.0380882
R35855 DVDD.n13595 DVDD.n12357 0.0380882
R35856 DVDD.n13605 DVDD.n12357 0.0380882
R35857 DVDD.n13606 DVDD.n13605 0.0380882
R35858 DVDD.n13607 DVDD.n13606 0.0380882
R35859 DVDD.n13607 DVDD.n12355 0.0380882
R35860 DVDD.n13617 DVDD.n12355 0.0380882
R35861 DVDD.n13618 DVDD.n13617 0.0380882
R35862 DVDD.n13619 DVDD.n13618 0.0380882
R35863 DVDD.n13619 DVDD.n12353 0.0380882
R35864 DVDD.n13629 DVDD.n12353 0.0380882
R35865 DVDD.n13630 DVDD.n13629 0.0380882
R35866 DVDD.n13631 DVDD.n13630 0.0380882
R35867 DVDD.n13631 DVDD.n12351 0.0380882
R35868 DVDD.n13641 DVDD.n12351 0.0380882
R35869 DVDD.n13642 DVDD.n13641 0.0380882
R35870 DVDD.n13643 DVDD.n13642 0.0380882
R35871 DVDD.n13643 DVDD.n12349 0.0380882
R35872 DVDD.n13653 DVDD.n12349 0.0380882
R35873 DVDD.n13654 DVDD.n13653 0.0380882
R35874 DVDD.n13655 DVDD.n13654 0.0380882
R35875 DVDD.n13655 DVDD.n12347 0.0380882
R35876 DVDD.n13665 DVDD.n12347 0.0380882
R35877 DVDD.n13666 DVDD.n13665 0.0380882
R35878 DVDD.n13667 DVDD.n13666 0.0380882
R35879 DVDD.n13667 DVDD.n12345 0.0380882
R35880 DVDD.n13677 DVDD.n12345 0.0380882
R35881 DVDD.n13678 DVDD.n13677 0.0380882
R35882 DVDD.n13679 DVDD.n13678 0.0380882
R35883 DVDD.n13679 DVDD.n12343 0.0380882
R35884 DVDD.n13689 DVDD.n12343 0.0380882
R35885 DVDD.n13690 DVDD.n13689 0.0380882
R35886 DVDD.n13691 DVDD.n13690 0.0380882
R35887 DVDD.n13691 DVDD.n12341 0.0380882
R35888 DVDD.n13701 DVDD.n12341 0.0380882
R35889 DVDD.n13702 DVDD.n13701 0.0380882
R35890 DVDD.n13703 DVDD.n13702 0.0380882
R35891 DVDD.n13703 DVDD.n12339 0.0380882
R35892 DVDD.n13713 DVDD.n12339 0.0380882
R35893 DVDD.n13714 DVDD.n13713 0.0380882
R35894 DVDD.n13715 DVDD.n13714 0.0380882
R35895 DVDD.n13715 DVDD.n12337 0.0380882
R35896 DVDD.n13725 DVDD.n12337 0.0380882
R35897 DVDD.n13726 DVDD.n13725 0.0380882
R35898 DVDD.n13727 DVDD.n13726 0.0380882
R35899 DVDD.n13727 DVDD.n12335 0.0380882
R35900 DVDD.n13737 DVDD.n12335 0.0380882
R35901 DVDD.n13738 DVDD.n13737 0.0380882
R35902 DVDD.n13739 DVDD.n13738 0.0380882
R35903 DVDD.n13739 DVDD.n12281 0.0380882
R35904 DVDD.n13496 DVDD.n12376 0.0380882
R35905 DVDD.n13500 DVDD.n12376 0.0380882
R35906 DVDD.n13504 DVDD.n13500 0.0380882
R35907 DVDD.n13508 DVDD.n13504 0.0380882
R35908 DVDD.n13508 DVDD.n12372 0.0380882
R35909 DVDD.n13512 DVDD.n12372 0.0380882
R35910 DVDD.n13516 DVDD.n13512 0.0380882
R35911 DVDD.n13520 DVDD.n13516 0.0380882
R35912 DVDD.n13520 DVDD.n12370 0.0380882
R35913 DVDD.n13524 DVDD.n12370 0.0380882
R35914 DVDD.n13528 DVDD.n13524 0.0380882
R35915 DVDD.n13532 DVDD.n13528 0.0380882
R35916 DVDD.n13532 DVDD.n12368 0.0380882
R35917 DVDD.n13536 DVDD.n12368 0.0380882
R35918 DVDD.n13540 DVDD.n13536 0.0380882
R35919 DVDD.n13544 DVDD.n13540 0.0380882
R35920 DVDD.n13544 DVDD.n12366 0.0380882
R35921 DVDD.n13548 DVDD.n12366 0.0380882
R35922 DVDD.n13552 DVDD.n13548 0.0380882
R35923 DVDD.n13556 DVDD.n13552 0.0380882
R35924 DVDD.n13556 DVDD.n12364 0.0380882
R35925 DVDD.n13560 DVDD.n12364 0.0380882
R35926 DVDD.n13564 DVDD.n13560 0.0380882
R35927 DVDD.n13568 DVDD.n13564 0.0380882
R35928 DVDD.n13568 DVDD.n12362 0.0380882
R35929 DVDD.n13572 DVDD.n12362 0.0380882
R35930 DVDD.n13576 DVDD.n13572 0.0380882
R35931 DVDD.n13580 DVDD.n13576 0.0380882
R35932 DVDD.n13580 DVDD.n12360 0.0380882
R35933 DVDD.n13584 DVDD.n12360 0.0380882
R35934 DVDD.n13588 DVDD.n13584 0.0380882
R35935 DVDD.n13592 DVDD.n13588 0.0380882
R35936 DVDD.n13592 DVDD.n12358 0.0380882
R35937 DVDD.n13596 DVDD.n12358 0.0380882
R35938 DVDD.n13600 DVDD.n13596 0.0380882
R35939 DVDD.n13604 DVDD.n13600 0.0380882
R35940 DVDD.n13604 DVDD.n12356 0.0380882
R35941 DVDD.n13608 DVDD.n12356 0.0380882
R35942 DVDD.n13612 DVDD.n13608 0.0380882
R35943 DVDD.n13616 DVDD.n13612 0.0380882
R35944 DVDD.n13616 DVDD.n12354 0.0380882
R35945 DVDD.n13620 DVDD.n12354 0.0380882
R35946 DVDD.n13624 DVDD.n13620 0.0380882
R35947 DVDD.n13628 DVDD.n13624 0.0380882
R35948 DVDD.n13628 DVDD.n12352 0.0380882
R35949 DVDD.n13632 DVDD.n12352 0.0380882
R35950 DVDD.n13636 DVDD.n13632 0.0380882
R35951 DVDD.n13640 DVDD.n13636 0.0380882
R35952 DVDD.n13640 DVDD.n12350 0.0380882
R35953 DVDD.n13644 DVDD.n12350 0.0380882
R35954 DVDD.n13648 DVDD.n13644 0.0380882
R35955 DVDD.n13652 DVDD.n13648 0.0380882
R35956 DVDD.n13652 DVDD.n12348 0.0380882
R35957 DVDD.n13656 DVDD.n12348 0.0380882
R35958 DVDD.n13660 DVDD.n13656 0.0380882
R35959 DVDD.n13664 DVDD.n13660 0.0380882
R35960 DVDD.n13664 DVDD.n12346 0.0380882
R35961 DVDD.n13668 DVDD.n12346 0.0380882
R35962 DVDD.n13672 DVDD.n13668 0.0380882
R35963 DVDD.n13676 DVDD.n13672 0.0380882
R35964 DVDD.n13676 DVDD.n12344 0.0380882
R35965 DVDD.n13680 DVDD.n12344 0.0380882
R35966 DVDD.n13684 DVDD.n13680 0.0380882
R35967 DVDD.n13688 DVDD.n13684 0.0380882
R35968 DVDD.n13688 DVDD.n12342 0.0380882
R35969 DVDD.n13692 DVDD.n12342 0.0380882
R35970 DVDD.n13696 DVDD.n13692 0.0380882
R35971 DVDD.n13700 DVDD.n13696 0.0380882
R35972 DVDD.n13700 DVDD.n12340 0.0380882
R35973 DVDD.n13704 DVDD.n12340 0.0380882
R35974 DVDD.n13708 DVDD.n13704 0.0380882
R35975 DVDD.n13712 DVDD.n13708 0.0380882
R35976 DVDD.n13712 DVDD.n12338 0.0380882
R35977 DVDD.n13716 DVDD.n12338 0.0380882
R35978 DVDD.n13720 DVDD.n13716 0.0380882
R35979 DVDD.n13724 DVDD.n13720 0.0380882
R35980 DVDD.n13724 DVDD.n12336 0.0380882
R35981 DVDD.n13728 DVDD.n12336 0.0380882
R35982 DVDD.n13732 DVDD.n13728 0.0380882
R35983 DVDD.n13736 DVDD.n13732 0.0380882
R35984 DVDD.n13736 DVDD.n12334 0.0380882
R35985 DVDD.n13740 DVDD.n12334 0.0380882
R35986 DVDD.n13740 DVDD.n12331 0.0380882
R35987 DVDD.n12543 DVDD.n12541 0.0380882
R35988 DVDD.n12544 DVDD.n12543 0.0380882
R35989 DVDD.n12545 DVDD.n12544 0.0380882
R35990 DVDD.n12545 DVDD.n12538 0.0380882
R35991 DVDD.n12552 DVDD.n12538 0.0380882
R35992 DVDD.n12553 DVDD.n12552 0.0380882
R35993 DVDD.n12554 DVDD.n12553 0.0380882
R35994 DVDD.n12554 DVDD.n12535 0.0380882
R35995 DVDD.n12561 DVDD.n12535 0.0380882
R35996 DVDD.n12562 DVDD.n12561 0.0380882
R35997 DVDD.n12563 DVDD.n12562 0.0380882
R35998 DVDD.n12563 DVDD.n12532 0.0380882
R35999 DVDD.n12570 DVDD.n12532 0.0380882
R36000 DVDD.n12571 DVDD.n12570 0.0380882
R36001 DVDD.n12572 DVDD.n12571 0.0380882
R36002 DVDD.n12572 DVDD.n12529 0.0380882
R36003 DVDD.n12579 DVDD.n12529 0.0380882
R36004 DVDD.n12580 DVDD.n12579 0.0380882
R36005 DVDD.n12581 DVDD.n12580 0.0380882
R36006 DVDD.n12581 DVDD.n12526 0.0380882
R36007 DVDD.n12588 DVDD.n12526 0.0380882
R36008 DVDD.n12589 DVDD.n12588 0.0380882
R36009 DVDD.n12590 DVDD.n12589 0.0380882
R36010 DVDD.n12590 DVDD.n12523 0.0380882
R36011 DVDD.n12597 DVDD.n12523 0.0380882
R36012 DVDD.n12598 DVDD.n12597 0.0380882
R36013 DVDD.n12599 DVDD.n12598 0.0380882
R36014 DVDD.n12599 DVDD.n12520 0.0380882
R36015 DVDD.n12606 DVDD.n12520 0.0380882
R36016 DVDD.n12607 DVDD.n12606 0.0380882
R36017 DVDD.n12608 DVDD.n12607 0.0380882
R36018 DVDD.n12608 DVDD.n12517 0.0380882
R36019 DVDD.n12615 DVDD.n12517 0.0380882
R36020 DVDD.n12616 DVDD.n12615 0.0380882
R36021 DVDD.n12617 DVDD.n12616 0.0380882
R36022 DVDD.n12617 DVDD.n12514 0.0380882
R36023 DVDD.n12624 DVDD.n12514 0.0380882
R36024 DVDD.n12625 DVDD.n12624 0.0380882
R36025 DVDD.n12626 DVDD.n12625 0.0380882
R36026 DVDD.n12626 DVDD.n12511 0.0380882
R36027 DVDD.n12633 DVDD.n12511 0.0380882
R36028 DVDD.n12634 DVDD.n12633 0.0380882
R36029 DVDD.n12635 DVDD.n12634 0.0380882
R36030 DVDD.n12635 DVDD.n12508 0.0380882
R36031 DVDD.n12642 DVDD.n12508 0.0380882
R36032 DVDD.n12643 DVDD.n12642 0.0380882
R36033 DVDD.n12644 DVDD.n12643 0.0380882
R36034 DVDD.n12644 DVDD.n12505 0.0380882
R36035 DVDD.n12651 DVDD.n12505 0.0380882
R36036 DVDD.n12652 DVDD.n12651 0.0380882
R36037 DVDD.n12653 DVDD.n12652 0.0380882
R36038 DVDD.n12653 DVDD.n12502 0.0380882
R36039 DVDD.n12660 DVDD.n12502 0.0380882
R36040 DVDD.n12661 DVDD.n12660 0.0380882
R36041 DVDD.n12662 DVDD.n12661 0.0380882
R36042 DVDD.n12662 DVDD.n12499 0.0380882
R36043 DVDD.n12669 DVDD.n12499 0.0380882
R36044 DVDD.n12670 DVDD.n12669 0.0380882
R36045 DVDD.n12671 DVDD.n12670 0.0380882
R36046 DVDD.n12671 DVDD.n12496 0.0380882
R36047 DVDD.n12678 DVDD.n12496 0.0380882
R36048 DVDD.n12679 DVDD.n12678 0.0380882
R36049 DVDD.n12680 DVDD.n12679 0.0380882
R36050 DVDD.n12680 DVDD.n12493 0.0380882
R36051 DVDD.n12687 DVDD.n12493 0.0380882
R36052 DVDD.n12688 DVDD.n12687 0.0380882
R36053 DVDD.n12689 DVDD.n12688 0.0380882
R36054 DVDD.n12689 DVDD.n12490 0.0380882
R36055 DVDD.n12696 DVDD.n12490 0.0380882
R36056 DVDD.n12697 DVDD.n12696 0.0380882
R36057 DVDD.n12698 DVDD.n12697 0.0380882
R36058 DVDD.n12698 DVDD.n12487 0.0380882
R36059 DVDD.n12705 DVDD.n12487 0.0380882
R36060 DVDD.n12706 DVDD.n12705 0.0380882
R36061 DVDD.n12707 DVDD.n12706 0.0380882
R36062 DVDD.n12707 DVDD.n12484 0.0380882
R36063 DVDD.n12714 DVDD.n12484 0.0380882
R36064 DVDD.n12715 DVDD.n12714 0.0380882
R36065 DVDD.n12716 DVDD.n12715 0.0380882
R36066 DVDD.n12716 DVDD.n12481 0.0380882
R36067 DVDD.n12723 DVDD.n12481 0.0380882
R36068 DVDD.n12724 DVDD.n12723 0.0380882
R36069 DVDD.n12725 DVDD.n12724 0.0380882
R36070 DVDD.n12542 DVDD.n12434 0.0380882
R36071 DVDD.n12542 DVDD.n12540 0.0380882
R36072 DVDD.n12547 DVDD.n12540 0.0380882
R36073 DVDD.n12549 DVDD.n12547 0.0380882
R36074 DVDD.n12551 DVDD.n12549 0.0380882
R36075 DVDD.n12551 DVDD.n12537 0.0380882
R36076 DVDD.n12556 DVDD.n12537 0.0380882
R36077 DVDD.n12558 DVDD.n12556 0.0380882
R36078 DVDD.n12560 DVDD.n12558 0.0380882
R36079 DVDD.n12560 DVDD.n12534 0.0380882
R36080 DVDD.n12565 DVDD.n12534 0.0380882
R36081 DVDD.n12567 DVDD.n12565 0.0380882
R36082 DVDD.n12569 DVDD.n12567 0.0380882
R36083 DVDD.n12569 DVDD.n12531 0.0380882
R36084 DVDD.n12574 DVDD.n12531 0.0380882
R36085 DVDD.n12576 DVDD.n12574 0.0380882
R36086 DVDD.n12578 DVDD.n12576 0.0380882
R36087 DVDD.n12578 DVDD.n12528 0.0380882
R36088 DVDD.n12583 DVDD.n12528 0.0380882
R36089 DVDD.n12585 DVDD.n12583 0.0380882
R36090 DVDD.n12587 DVDD.n12585 0.0380882
R36091 DVDD.n12587 DVDD.n12525 0.0380882
R36092 DVDD.n12592 DVDD.n12525 0.0380882
R36093 DVDD.n12594 DVDD.n12592 0.0380882
R36094 DVDD.n12596 DVDD.n12594 0.0380882
R36095 DVDD.n12596 DVDD.n12522 0.0380882
R36096 DVDD.n12601 DVDD.n12522 0.0380882
R36097 DVDD.n12603 DVDD.n12601 0.0380882
R36098 DVDD.n12605 DVDD.n12603 0.0380882
R36099 DVDD.n12605 DVDD.n12519 0.0380882
R36100 DVDD.n12610 DVDD.n12519 0.0380882
R36101 DVDD.n12612 DVDD.n12610 0.0380882
R36102 DVDD.n12614 DVDD.n12612 0.0380882
R36103 DVDD.n12614 DVDD.n12516 0.0380882
R36104 DVDD.n12619 DVDD.n12516 0.0380882
R36105 DVDD.n12621 DVDD.n12619 0.0380882
R36106 DVDD.n12623 DVDD.n12621 0.0380882
R36107 DVDD.n12623 DVDD.n12513 0.0380882
R36108 DVDD.n12628 DVDD.n12513 0.0380882
R36109 DVDD.n12630 DVDD.n12628 0.0380882
R36110 DVDD.n12632 DVDD.n12630 0.0380882
R36111 DVDD.n12632 DVDD.n12510 0.0380882
R36112 DVDD.n12637 DVDD.n12510 0.0380882
R36113 DVDD.n12639 DVDD.n12637 0.0380882
R36114 DVDD.n12641 DVDD.n12639 0.0380882
R36115 DVDD.n12641 DVDD.n12507 0.0380882
R36116 DVDD.n12646 DVDD.n12507 0.0380882
R36117 DVDD.n12648 DVDD.n12646 0.0380882
R36118 DVDD.n12650 DVDD.n12648 0.0380882
R36119 DVDD.n12650 DVDD.n12504 0.0380882
R36120 DVDD.n12655 DVDD.n12504 0.0380882
R36121 DVDD.n12657 DVDD.n12655 0.0380882
R36122 DVDD.n12659 DVDD.n12657 0.0380882
R36123 DVDD.n12659 DVDD.n12501 0.0380882
R36124 DVDD.n12664 DVDD.n12501 0.0380882
R36125 DVDD.n12666 DVDD.n12664 0.0380882
R36126 DVDD.n12668 DVDD.n12666 0.0380882
R36127 DVDD.n12668 DVDD.n12498 0.0380882
R36128 DVDD.n12673 DVDD.n12498 0.0380882
R36129 DVDD.n12675 DVDD.n12673 0.0380882
R36130 DVDD.n12677 DVDD.n12675 0.0380882
R36131 DVDD.n12677 DVDD.n12495 0.0380882
R36132 DVDD.n12682 DVDD.n12495 0.0380882
R36133 DVDD.n12684 DVDD.n12682 0.0380882
R36134 DVDD.n12686 DVDD.n12684 0.0380882
R36135 DVDD.n12686 DVDD.n12492 0.0380882
R36136 DVDD.n12691 DVDD.n12492 0.0380882
R36137 DVDD.n12693 DVDD.n12691 0.0380882
R36138 DVDD.n12695 DVDD.n12693 0.0380882
R36139 DVDD.n12695 DVDD.n12489 0.0380882
R36140 DVDD.n12700 DVDD.n12489 0.0380882
R36141 DVDD.n12702 DVDD.n12700 0.0380882
R36142 DVDD.n12704 DVDD.n12702 0.0380882
R36143 DVDD.n12704 DVDD.n12486 0.0380882
R36144 DVDD.n12709 DVDD.n12486 0.0380882
R36145 DVDD.n12711 DVDD.n12709 0.0380882
R36146 DVDD.n12713 DVDD.n12711 0.0380882
R36147 DVDD.n12713 DVDD.n12483 0.0380882
R36148 DVDD.n12718 DVDD.n12483 0.0380882
R36149 DVDD.n12720 DVDD.n12718 0.0380882
R36150 DVDD.n12722 DVDD.n12720 0.0380882
R36151 DVDD.n12722 DVDD.n12480 0.0380882
R36152 DVDD.n13482 DVDD.n12480 0.0380882
R36153 DVDD.n13285 DVDD.n13283 0.0380882
R36154 DVDD.n13286 DVDD.n13285 0.0380882
R36155 DVDD.n13287 DVDD.n13286 0.0380882
R36156 DVDD.n13287 DVDD.n12885 0.0380882
R36157 DVDD.n13294 DVDD.n12885 0.0380882
R36158 DVDD.n13295 DVDD.n13294 0.0380882
R36159 DVDD.n13296 DVDD.n13295 0.0380882
R36160 DVDD.n13296 DVDD.n12882 0.0380882
R36161 DVDD.n13303 DVDD.n12882 0.0380882
R36162 DVDD.n13304 DVDD.n13303 0.0380882
R36163 DVDD.n13305 DVDD.n13304 0.0380882
R36164 DVDD.n13305 DVDD.n12879 0.0380882
R36165 DVDD.n13312 DVDD.n12879 0.0380882
R36166 DVDD.n13313 DVDD.n13312 0.0380882
R36167 DVDD.n13314 DVDD.n13313 0.0380882
R36168 DVDD.n13314 DVDD.n12876 0.0380882
R36169 DVDD.n13321 DVDD.n12876 0.0380882
R36170 DVDD.n13322 DVDD.n13321 0.0380882
R36171 DVDD.n13323 DVDD.n13322 0.0380882
R36172 DVDD.n13323 DVDD.n12873 0.0380882
R36173 DVDD.n13330 DVDD.n12873 0.0380882
R36174 DVDD.n13331 DVDD.n13330 0.0380882
R36175 DVDD.n13332 DVDD.n13331 0.0380882
R36176 DVDD.n13332 DVDD.n12870 0.0380882
R36177 DVDD.n13339 DVDD.n12870 0.0380882
R36178 DVDD.n13340 DVDD.n13339 0.0380882
R36179 DVDD.n13341 DVDD.n13340 0.0380882
R36180 DVDD.n13341 DVDD.n12867 0.0380882
R36181 DVDD.n13348 DVDD.n12867 0.0380882
R36182 DVDD.n13349 DVDD.n13348 0.0380882
R36183 DVDD.n13350 DVDD.n13349 0.0380882
R36184 DVDD.n13350 DVDD.n12864 0.0380882
R36185 DVDD.n13357 DVDD.n12864 0.0380882
R36186 DVDD.n13358 DVDD.n13357 0.0380882
R36187 DVDD.n13359 DVDD.n13358 0.0380882
R36188 DVDD.n13359 DVDD.n12861 0.0380882
R36189 DVDD.n13366 DVDD.n12861 0.0380882
R36190 DVDD.n13367 DVDD.n13366 0.0380882
R36191 DVDD.n13368 DVDD.n13367 0.0380882
R36192 DVDD.n13368 DVDD.n12858 0.0380882
R36193 DVDD.n13375 DVDD.n12858 0.0380882
R36194 DVDD.n13376 DVDD.n13375 0.0380882
R36195 DVDD.n13377 DVDD.n13376 0.0380882
R36196 DVDD.n13377 DVDD.n12855 0.0380882
R36197 DVDD.n13384 DVDD.n12855 0.0380882
R36198 DVDD.n13385 DVDD.n13384 0.0380882
R36199 DVDD.n13386 DVDD.n13385 0.0380882
R36200 DVDD.n13386 DVDD.n12852 0.0380882
R36201 DVDD.n13393 DVDD.n12852 0.0380882
R36202 DVDD.n13394 DVDD.n13393 0.0380882
R36203 DVDD.n13395 DVDD.n13394 0.0380882
R36204 DVDD.n13395 DVDD.n12849 0.0380882
R36205 DVDD.n13402 DVDD.n12849 0.0380882
R36206 DVDD.n13403 DVDD.n13402 0.0380882
R36207 DVDD.n13404 DVDD.n13403 0.0380882
R36208 DVDD.n13404 DVDD.n12846 0.0380882
R36209 DVDD.n13411 DVDD.n12846 0.0380882
R36210 DVDD.n13412 DVDD.n13411 0.0380882
R36211 DVDD.n13413 DVDD.n13412 0.0380882
R36212 DVDD.n13413 DVDD.n12843 0.0380882
R36213 DVDD.n13420 DVDD.n12843 0.0380882
R36214 DVDD.n13421 DVDD.n13420 0.0380882
R36215 DVDD.n13422 DVDD.n13421 0.0380882
R36216 DVDD.n13422 DVDD.n12840 0.0380882
R36217 DVDD.n13429 DVDD.n12840 0.0380882
R36218 DVDD.n13430 DVDD.n13429 0.0380882
R36219 DVDD.n13431 DVDD.n13430 0.0380882
R36220 DVDD.n13431 DVDD.n12837 0.0380882
R36221 DVDD.n13438 DVDD.n12837 0.0380882
R36222 DVDD.n13439 DVDD.n13438 0.0380882
R36223 DVDD.n13440 DVDD.n13439 0.0380882
R36224 DVDD.n13440 DVDD.n12834 0.0380882
R36225 DVDD.n13447 DVDD.n12834 0.0380882
R36226 DVDD.n13448 DVDD.n13447 0.0380882
R36227 DVDD.n13449 DVDD.n13448 0.0380882
R36228 DVDD.n13449 DVDD.n12831 0.0380882
R36229 DVDD.n13456 DVDD.n12831 0.0380882
R36230 DVDD.n13457 DVDD.n13456 0.0380882
R36231 DVDD.n13458 DVDD.n13457 0.0380882
R36232 DVDD.n13458 DVDD.n12828 0.0380882
R36233 DVDD.n13465 DVDD.n12828 0.0380882
R36234 DVDD.n13466 DVDD.n13465 0.0380882
R36235 DVDD.n13467 DVDD.n13466 0.0380882
R36236 DVDD.n13284 DVDD.n12782 0.0380882
R36237 DVDD.n13284 DVDD.n12887 0.0380882
R36238 DVDD.n13289 DVDD.n12887 0.0380882
R36239 DVDD.n13291 DVDD.n13289 0.0380882
R36240 DVDD.n13293 DVDD.n13291 0.0380882
R36241 DVDD.n13293 DVDD.n12884 0.0380882
R36242 DVDD.n13298 DVDD.n12884 0.0380882
R36243 DVDD.n13300 DVDD.n13298 0.0380882
R36244 DVDD.n13302 DVDD.n13300 0.0380882
R36245 DVDD.n13302 DVDD.n12881 0.0380882
R36246 DVDD.n13307 DVDD.n12881 0.0380882
R36247 DVDD.n13309 DVDD.n13307 0.0380882
R36248 DVDD.n13311 DVDD.n13309 0.0380882
R36249 DVDD.n13311 DVDD.n12878 0.0380882
R36250 DVDD.n13316 DVDD.n12878 0.0380882
R36251 DVDD.n13318 DVDD.n13316 0.0380882
R36252 DVDD.n13320 DVDD.n13318 0.0380882
R36253 DVDD.n13320 DVDD.n12875 0.0380882
R36254 DVDD.n13325 DVDD.n12875 0.0380882
R36255 DVDD.n13327 DVDD.n13325 0.0380882
R36256 DVDD.n13329 DVDD.n13327 0.0380882
R36257 DVDD.n13329 DVDD.n12872 0.0380882
R36258 DVDD.n13334 DVDD.n12872 0.0380882
R36259 DVDD.n13336 DVDD.n13334 0.0380882
R36260 DVDD.n13338 DVDD.n13336 0.0380882
R36261 DVDD.n13338 DVDD.n12869 0.0380882
R36262 DVDD.n13343 DVDD.n12869 0.0380882
R36263 DVDD.n13345 DVDD.n13343 0.0380882
R36264 DVDD.n13347 DVDD.n13345 0.0380882
R36265 DVDD.n13347 DVDD.n12866 0.0380882
R36266 DVDD.n13352 DVDD.n12866 0.0380882
R36267 DVDD.n13354 DVDD.n13352 0.0380882
R36268 DVDD.n13356 DVDD.n13354 0.0380882
R36269 DVDD.n13356 DVDD.n12863 0.0380882
R36270 DVDD.n13361 DVDD.n12863 0.0380882
R36271 DVDD.n13363 DVDD.n13361 0.0380882
R36272 DVDD.n13365 DVDD.n13363 0.0380882
R36273 DVDD.n13365 DVDD.n12860 0.0380882
R36274 DVDD.n13370 DVDD.n12860 0.0380882
R36275 DVDD.n13372 DVDD.n13370 0.0380882
R36276 DVDD.n13374 DVDD.n13372 0.0380882
R36277 DVDD.n13374 DVDD.n12857 0.0380882
R36278 DVDD.n13379 DVDD.n12857 0.0380882
R36279 DVDD.n13381 DVDD.n13379 0.0380882
R36280 DVDD.n13383 DVDD.n13381 0.0380882
R36281 DVDD.n13383 DVDD.n12854 0.0380882
R36282 DVDD.n13388 DVDD.n12854 0.0380882
R36283 DVDD.n13390 DVDD.n13388 0.0380882
R36284 DVDD.n13392 DVDD.n13390 0.0380882
R36285 DVDD.n13392 DVDD.n12851 0.0380882
R36286 DVDD.n13397 DVDD.n12851 0.0380882
R36287 DVDD.n13399 DVDD.n13397 0.0380882
R36288 DVDD.n13401 DVDD.n13399 0.0380882
R36289 DVDD.n13401 DVDD.n12848 0.0380882
R36290 DVDD.n13406 DVDD.n12848 0.0380882
R36291 DVDD.n13408 DVDD.n13406 0.0380882
R36292 DVDD.n13410 DVDD.n13408 0.0380882
R36293 DVDD.n13410 DVDD.n12845 0.0380882
R36294 DVDD.n13415 DVDD.n12845 0.0380882
R36295 DVDD.n13417 DVDD.n13415 0.0380882
R36296 DVDD.n13419 DVDD.n13417 0.0380882
R36297 DVDD.n13419 DVDD.n12842 0.0380882
R36298 DVDD.n13424 DVDD.n12842 0.0380882
R36299 DVDD.n13426 DVDD.n13424 0.0380882
R36300 DVDD.n13428 DVDD.n13426 0.0380882
R36301 DVDD.n13428 DVDD.n12839 0.0380882
R36302 DVDD.n13433 DVDD.n12839 0.0380882
R36303 DVDD.n13435 DVDD.n13433 0.0380882
R36304 DVDD.n13437 DVDD.n13435 0.0380882
R36305 DVDD.n13437 DVDD.n12836 0.0380882
R36306 DVDD.n13442 DVDD.n12836 0.0380882
R36307 DVDD.n13444 DVDD.n13442 0.0380882
R36308 DVDD.n13446 DVDD.n13444 0.0380882
R36309 DVDD.n13446 DVDD.n12833 0.0380882
R36310 DVDD.n13451 DVDD.n12833 0.0380882
R36311 DVDD.n13453 DVDD.n13451 0.0380882
R36312 DVDD.n13455 DVDD.n13453 0.0380882
R36313 DVDD.n13455 DVDD.n12830 0.0380882
R36314 DVDD.n13460 DVDD.n12830 0.0380882
R36315 DVDD.n13462 DVDD.n13460 0.0380882
R36316 DVDD.n13464 DVDD.n13462 0.0380882
R36317 DVDD.n13464 DVDD.n12827 0.0380882
R36318 DVDD.n13468 DVDD.n12827 0.0380882
R36319 DVDD.n13251 DVDD.n12903 0.0380882
R36320 DVDD.n13251 DVDD.n13250 0.0380882
R36321 DVDD.n13250 DVDD.n13249 0.0380882
R36322 DVDD.n13249 DVDD.n12968 0.0380882
R36323 DVDD.n13239 DVDD.n12968 0.0380882
R36324 DVDD.n13239 DVDD.n13238 0.0380882
R36325 DVDD.n13238 DVDD.n13237 0.0380882
R36326 DVDD.n13237 DVDD.n12970 0.0380882
R36327 DVDD.n13227 DVDD.n12970 0.0380882
R36328 DVDD.n13227 DVDD.n13226 0.0380882
R36329 DVDD.n13226 DVDD.n13225 0.0380882
R36330 DVDD.n13225 DVDD.n12972 0.0380882
R36331 DVDD.n13215 DVDD.n12972 0.0380882
R36332 DVDD.n13215 DVDD.n13214 0.0380882
R36333 DVDD.n13214 DVDD.n13213 0.0380882
R36334 DVDD.n13213 DVDD.n12974 0.0380882
R36335 DVDD.n13203 DVDD.n12974 0.0380882
R36336 DVDD.n13203 DVDD.n13202 0.0380882
R36337 DVDD.n13202 DVDD.n13201 0.0380882
R36338 DVDD.n13201 DVDD.n12976 0.0380882
R36339 DVDD.n13191 DVDD.n12976 0.0380882
R36340 DVDD.n13191 DVDD.n13190 0.0380882
R36341 DVDD.n13190 DVDD.n13189 0.0380882
R36342 DVDD.n13189 DVDD.n12978 0.0380882
R36343 DVDD.n13179 DVDD.n12978 0.0380882
R36344 DVDD.n13179 DVDD.n13178 0.0380882
R36345 DVDD.n13178 DVDD.n13177 0.0380882
R36346 DVDD.n13177 DVDD.n12980 0.0380882
R36347 DVDD.n13167 DVDD.n12980 0.0380882
R36348 DVDD.n13167 DVDD.n13166 0.0380882
R36349 DVDD.n13166 DVDD.n13165 0.0380882
R36350 DVDD.n13165 DVDD.n12982 0.0380882
R36351 DVDD.n13155 DVDD.n12982 0.0380882
R36352 DVDD.n13155 DVDD.n13154 0.0380882
R36353 DVDD.n13154 DVDD.n13153 0.0380882
R36354 DVDD.n13153 DVDD.n12984 0.0380882
R36355 DVDD.n13143 DVDD.n12984 0.0380882
R36356 DVDD.n13143 DVDD.n13142 0.0380882
R36357 DVDD.n13142 DVDD.n13141 0.0380882
R36358 DVDD.n13141 DVDD.n12986 0.0380882
R36359 DVDD.n13131 DVDD.n12986 0.0380882
R36360 DVDD.n13131 DVDD.n13130 0.0380882
R36361 DVDD.n13130 DVDD.n13129 0.0380882
R36362 DVDD.n13129 DVDD.n12988 0.0380882
R36363 DVDD.n13119 DVDD.n12988 0.0380882
R36364 DVDD.n13119 DVDD.n13118 0.0380882
R36365 DVDD.n13118 DVDD.n13117 0.0380882
R36366 DVDD.n13117 DVDD.n12990 0.0380882
R36367 DVDD.n13107 DVDD.n12990 0.0380882
R36368 DVDD.n13107 DVDD.n13106 0.0380882
R36369 DVDD.n13106 DVDD.n13105 0.0380882
R36370 DVDD.n13105 DVDD.n12992 0.0380882
R36371 DVDD.n13095 DVDD.n12992 0.0380882
R36372 DVDD.n13095 DVDD.n13094 0.0380882
R36373 DVDD.n13094 DVDD.n13093 0.0380882
R36374 DVDD.n13093 DVDD.n12994 0.0380882
R36375 DVDD.n13083 DVDD.n12994 0.0380882
R36376 DVDD.n13083 DVDD.n13082 0.0380882
R36377 DVDD.n13082 DVDD.n13081 0.0380882
R36378 DVDD.n13081 DVDD.n12996 0.0380882
R36379 DVDD.n13071 DVDD.n12996 0.0380882
R36380 DVDD.n13071 DVDD.n13070 0.0380882
R36381 DVDD.n13070 DVDD.n13069 0.0380882
R36382 DVDD.n13069 DVDD.n12998 0.0380882
R36383 DVDD.n13059 DVDD.n12998 0.0380882
R36384 DVDD.n13059 DVDD.n13058 0.0380882
R36385 DVDD.n13058 DVDD.n13057 0.0380882
R36386 DVDD.n13057 DVDD.n13000 0.0380882
R36387 DVDD.n13047 DVDD.n13000 0.0380882
R36388 DVDD.n13047 DVDD.n13046 0.0380882
R36389 DVDD.n13046 DVDD.n13045 0.0380882
R36390 DVDD.n13045 DVDD.n13002 0.0380882
R36391 DVDD.n13035 DVDD.n13002 0.0380882
R36392 DVDD.n13035 DVDD.n13034 0.0380882
R36393 DVDD.n13034 DVDD.n13033 0.0380882
R36394 DVDD.n13033 DVDD.n13004 0.0380882
R36395 DVDD.n13023 DVDD.n13004 0.0380882
R36396 DVDD.n13023 DVDD.n13022 0.0380882
R36397 DVDD.n13022 DVDD.n13021 0.0380882
R36398 DVDD.n13021 DVDD.n13006 0.0380882
R36399 DVDD.n13011 DVDD.n13006 0.0380882
R36400 DVDD.n13011 DVDD.n13010 0.0380882
R36401 DVDD.n13010 DVDD.n12915 0.0380882
R36402 DVDD.n13253 DVDD.n13252 0.0380882
R36403 DVDD.n13252 DVDD.n12967 0.0380882
R36404 DVDD.n13248 DVDD.n12967 0.0380882
R36405 DVDD.n13248 DVDD.n13244 0.0380882
R36406 DVDD.n13244 DVDD.n13243 0.0380882
R36407 DVDD.n13243 DVDD.n12969 0.0380882
R36408 DVDD.n13236 DVDD.n12969 0.0380882
R36409 DVDD.n13236 DVDD.n13232 0.0380882
R36410 DVDD.n13232 DVDD.n13231 0.0380882
R36411 DVDD.n13231 DVDD.n12971 0.0380882
R36412 DVDD.n13224 DVDD.n12971 0.0380882
R36413 DVDD.n13224 DVDD.n13220 0.0380882
R36414 DVDD.n13220 DVDD.n13219 0.0380882
R36415 DVDD.n13219 DVDD.n12973 0.0380882
R36416 DVDD.n13212 DVDD.n12973 0.0380882
R36417 DVDD.n13212 DVDD.n13208 0.0380882
R36418 DVDD.n13208 DVDD.n13207 0.0380882
R36419 DVDD.n13207 DVDD.n12975 0.0380882
R36420 DVDD.n13200 DVDD.n12975 0.0380882
R36421 DVDD.n13200 DVDD.n13196 0.0380882
R36422 DVDD.n13196 DVDD.n13195 0.0380882
R36423 DVDD.n13195 DVDD.n12977 0.0380882
R36424 DVDD.n13188 DVDD.n12977 0.0380882
R36425 DVDD.n13188 DVDD.n13184 0.0380882
R36426 DVDD.n13184 DVDD.n13183 0.0380882
R36427 DVDD.n13183 DVDD.n12979 0.0380882
R36428 DVDD.n13176 DVDD.n12979 0.0380882
R36429 DVDD.n13176 DVDD.n13172 0.0380882
R36430 DVDD.n13172 DVDD.n13171 0.0380882
R36431 DVDD.n13171 DVDD.n12981 0.0380882
R36432 DVDD.n13164 DVDD.n12981 0.0380882
R36433 DVDD.n13164 DVDD.n13160 0.0380882
R36434 DVDD.n13160 DVDD.n13159 0.0380882
R36435 DVDD.n13159 DVDD.n12983 0.0380882
R36436 DVDD.n13152 DVDD.n12983 0.0380882
R36437 DVDD.n13152 DVDD.n13148 0.0380882
R36438 DVDD.n13148 DVDD.n13147 0.0380882
R36439 DVDD.n13147 DVDD.n12985 0.0380882
R36440 DVDD.n13140 DVDD.n12985 0.0380882
R36441 DVDD.n13140 DVDD.n13136 0.0380882
R36442 DVDD.n13136 DVDD.n13135 0.0380882
R36443 DVDD.n13135 DVDD.n12987 0.0380882
R36444 DVDD.n13128 DVDD.n12987 0.0380882
R36445 DVDD.n13128 DVDD.n13124 0.0380882
R36446 DVDD.n13124 DVDD.n13123 0.0380882
R36447 DVDD.n13123 DVDD.n12989 0.0380882
R36448 DVDD.n13116 DVDD.n12989 0.0380882
R36449 DVDD.n13116 DVDD.n13112 0.0380882
R36450 DVDD.n13112 DVDD.n13111 0.0380882
R36451 DVDD.n13111 DVDD.n12991 0.0380882
R36452 DVDD.n13104 DVDD.n12991 0.0380882
R36453 DVDD.n13104 DVDD.n13100 0.0380882
R36454 DVDD.n13100 DVDD.n13099 0.0380882
R36455 DVDD.n13099 DVDD.n12993 0.0380882
R36456 DVDD.n13092 DVDD.n12993 0.0380882
R36457 DVDD.n13092 DVDD.n13088 0.0380882
R36458 DVDD.n13088 DVDD.n13087 0.0380882
R36459 DVDD.n13087 DVDD.n12995 0.0380882
R36460 DVDD.n13080 DVDD.n12995 0.0380882
R36461 DVDD.n13080 DVDD.n13076 0.0380882
R36462 DVDD.n13076 DVDD.n13075 0.0380882
R36463 DVDD.n13075 DVDD.n12997 0.0380882
R36464 DVDD.n13068 DVDD.n12997 0.0380882
R36465 DVDD.n13068 DVDD.n13064 0.0380882
R36466 DVDD.n13064 DVDD.n13063 0.0380882
R36467 DVDD.n13063 DVDD.n12999 0.0380882
R36468 DVDD.n13056 DVDD.n12999 0.0380882
R36469 DVDD.n13056 DVDD.n13052 0.0380882
R36470 DVDD.n13052 DVDD.n13051 0.0380882
R36471 DVDD.n13051 DVDD.n13001 0.0380882
R36472 DVDD.n13044 DVDD.n13001 0.0380882
R36473 DVDD.n13044 DVDD.n13040 0.0380882
R36474 DVDD.n13040 DVDD.n13039 0.0380882
R36475 DVDD.n13039 DVDD.n13003 0.0380882
R36476 DVDD.n13032 DVDD.n13003 0.0380882
R36477 DVDD.n13032 DVDD.n13028 0.0380882
R36478 DVDD.n13028 DVDD.n13027 0.0380882
R36479 DVDD.n13027 DVDD.n13005 0.0380882
R36480 DVDD.n13020 DVDD.n13005 0.0380882
R36481 DVDD.n13020 DVDD.n13016 0.0380882
R36482 DVDD.n13016 DVDD.n13015 0.0380882
R36483 DVDD.n13015 DVDD.n13009 0.0380882
R36484 DVDD.n13009 DVDD.n13008 0.0380882
R36485 DVDD.n16458 DVDD.n16457 0.0380882
R36486 DVDD.n16459 DVDD.n16458 0.0380882
R36487 DVDD.n16459 DVDD.n2250 0.0380882
R36488 DVDD.n16469 DVDD.n2250 0.0380882
R36489 DVDD.n16470 DVDD.n16469 0.0380882
R36490 DVDD.n16471 DVDD.n16470 0.0380882
R36491 DVDD.n16471 DVDD.n2248 0.0380882
R36492 DVDD.n16481 DVDD.n2248 0.0380882
R36493 DVDD.n16482 DVDD.n16481 0.0380882
R36494 DVDD.n16483 DVDD.n16482 0.0380882
R36495 DVDD.n16483 DVDD.n2246 0.0380882
R36496 DVDD.n16493 DVDD.n2246 0.0380882
R36497 DVDD.n16494 DVDD.n16493 0.0380882
R36498 DVDD.n16495 DVDD.n16494 0.0380882
R36499 DVDD.n16495 DVDD.n2244 0.0380882
R36500 DVDD.n16505 DVDD.n2244 0.0380882
R36501 DVDD.n16506 DVDD.n16505 0.0380882
R36502 DVDD.n16507 DVDD.n16506 0.0380882
R36503 DVDD.n16507 DVDD.n2242 0.0380882
R36504 DVDD.n16517 DVDD.n2242 0.0380882
R36505 DVDD.n16518 DVDD.n16517 0.0380882
R36506 DVDD.n16519 DVDD.n16518 0.0380882
R36507 DVDD.n16519 DVDD.n2240 0.0380882
R36508 DVDD.n16529 DVDD.n2240 0.0380882
R36509 DVDD.n16530 DVDD.n16529 0.0380882
R36510 DVDD.n16531 DVDD.n16530 0.0380882
R36511 DVDD.n16531 DVDD.n2238 0.0380882
R36512 DVDD.n16541 DVDD.n2238 0.0380882
R36513 DVDD.n16542 DVDD.n16541 0.0380882
R36514 DVDD.n16543 DVDD.n16542 0.0380882
R36515 DVDD.n16543 DVDD.n2236 0.0380882
R36516 DVDD.n16553 DVDD.n2236 0.0380882
R36517 DVDD.n16554 DVDD.n16553 0.0380882
R36518 DVDD.n16555 DVDD.n16554 0.0380882
R36519 DVDD.n16555 DVDD.n2234 0.0380882
R36520 DVDD.n16565 DVDD.n2234 0.0380882
R36521 DVDD.n16566 DVDD.n16565 0.0380882
R36522 DVDD.n16567 DVDD.n16566 0.0380882
R36523 DVDD.n16567 DVDD.n2232 0.0380882
R36524 DVDD.n16577 DVDD.n2232 0.0380882
R36525 DVDD.n16578 DVDD.n16577 0.0380882
R36526 DVDD.n16579 DVDD.n16578 0.0380882
R36527 DVDD.n16579 DVDD.n2230 0.0380882
R36528 DVDD.n16589 DVDD.n2230 0.0380882
R36529 DVDD.n16590 DVDD.n16589 0.0380882
R36530 DVDD.n16591 DVDD.n16590 0.0380882
R36531 DVDD.n16591 DVDD.n2228 0.0380882
R36532 DVDD.n16601 DVDD.n2228 0.0380882
R36533 DVDD.n16602 DVDD.n16601 0.0380882
R36534 DVDD.n16603 DVDD.n16602 0.0380882
R36535 DVDD.n16603 DVDD.n2226 0.0380882
R36536 DVDD.n16613 DVDD.n2226 0.0380882
R36537 DVDD.n16614 DVDD.n16613 0.0380882
R36538 DVDD.n16615 DVDD.n16614 0.0380882
R36539 DVDD.n16615 DVDD.n2224 0.0380882
R36540 DVDD.n16625 DVDD.n2224 0.0380882
R36541 DVDD.n16626 DVDD.n16625 0.0380882
R36542 DVDD.n16627 DVDD.n16626 0.0380882
R36543 DVDD.n16627 DVDD.n2222 0.0380882
R36544 DVDD.n16637 DVDD.n2222 0.0380882
R36545 DVDD.n16638 DVDD.n16637 0.0380882
R36546 DVDD.n16639 DVDD.n16638 0.0380882
R36547 DVDD.n16639 DVDD.n2220 0.0380882
R36548 DVDD.n16649 DVDD.n2220 0.0380882
R36549 DVDD.n16650 DVDD.n16649 0.0380882
R36550 DVDD.n16651 DVDD.n16650 0.0380882
R36551 DVDD.n16651 DVDD.n2218 0.0380882
R36552 DVDD.n16661 DVDD.n2218 0.0380882
R36553 DVDD.n16662 DVDD.n16661 0.0380882
R36554 DVDD.n16663 DVDD.n16662 0.0380882
R36555 DVDD.n16663 DVDD.n2216 0.0380882
R36556 DVDD.n16673 DVDD.n2216 0.0380882
R36557 DVDD.n16674 DVDD.n16673 0.0380882
R36558 DVDD.n16675 DVDD.n16674 0.0380882
R36559 DVDD.n16675 DVDD.n2214 0.0380882
R36560 DVDD.n16685 DVDD.n2214 0.0380882
R36561 DVDD.n16686 DVDD.n16685 0.0380882
R36562 DVDD.n16687 DVDD.n16686 0.0380882
R36563 DVDD.n16687 DVDD.n2212 0.0380882
R36564 DVDD.n16697 DVDD.n2212 0.0380882
R36565 DVDD.n16698 DVDD.n16697 0.0380882
R36566 DVDD.n16699 DVDD.n16698 0.0380882
R36567 DVDD.n16699 DVDD.n2159 0.0380882
R36568 DVDD.n16456 DVDD.n2253 0.0380882
R36569 DVDD.n16460 DVDD.n2253 0.0380882
R36570 DVDD.n16464 DVDD.n16460 0.0380882
R36571 DVDD.n16468 DVDD.n16464 0.0380882
R36572 DVDD.n16468 DVDD.n2249 0.0380882
R36573 DVDD.n16472 DVDD.n2249 0.0380882
R36574 DVDD.n16476 DVDD.n16472 0.0380882
R36575 DVDD.n16480 DVDD.n16476 0.0380882
R36576 DVDD.n16480 DVDD.n2247 0.0380882
R36577 DVDD.n16484 DVDD.n2247 0.0380882
R36578 DVDD.n16488 DVDD.n16484 0.0380882
R36579 DVDD.n16492 DVDD.n16488 0.0380882
R36580 DVDD.n16492 DVDD.n2245 0.0380882
R36581 DVDD.n16496 DVDD.n2245 0.0380882
R36582 DVDD.n16500 DVDD.n16496 0.0380882
R36583 DVDD.n16504 DVDD.n16500 0.0380882
R36584 DVDD.n16504 DVDD.n2243 0.0380882
R36585 DVDD.n16508 DVDD.n2243 0.0380882
R36586 DVDD.n16512 DVDD.n16508 0.0380882
R36587 DVDD.n16516 DVDD.n16512 0.0380882
R36588 DVDD.n16516 DVDD.n2241 0.0380882
R36589 DVDD.n16520 DVDD.n2241 0.0380882
R36590 DVDD.n16524 DVDD.n16520 0.0380882
R36591 DVDD.n16528 DVDD.n16524 0.0380882
R36592 DVDD.n16528 DVDD.n2239 0.0380882
R36593 DVDD.n16532 DVDD.n2239 0.0380882
R36594 DVDD.n16536 DVDD.n16532 0.0380882
R36595 DVDD.n16540 DVDD.n16536 0.0380882
R36596 DVDD.n16540 DVDD.n2237 0.0380882
R36597 DVDD.n16544 DVDD.n2237 0.0380882
R36598 DVDD.n16548 DVDD.n16544 0.0380882
R36599 DVDD.n16552 DVDD.n16548 0.0380882
R36600 DVDD.n16552 DVDD.n2235 0.0380882
R36601 DVDD.n16556 DVDD.n2235 0.0380882
R36602 DVDD.n16560 DVDD.n16556 0.0380882
R36603 DVDD.n16564 DVDD.n16560 0.0380882
R36604 DVDD.n16564 DVDD.n2233 0.0380882
R36605 DVDD.n16568 DVDD.n2233 0.0380882
R36606 DVDD.n16572 DVDD.n16568 0.0380882
R36607 DVDD.n16576 DVDD.n16572 0.0380882
R36608 DVDD.n16576 DVDD.n2231 0.0380882
R36609 DVDD.n16580 DVDD.n2231 0.0380882
R36610 DVDD.n16584 DVDD.n16580 0.0380882
R36611 DVDD.n16588 DVDD.n16584 0.0380882
R36612 DVDD.n16588 DVDD.n2229 0.0380882
R36613 DVDD.n16592 DVDD.n2229 0.0380882
R36614 DVDD.n16596 DVDD.n16592 0.0380882
R36615 DVDD.n16600 DVDD.n16596 0.0380882
R36616 DVDD.n16600 DVDD.n2227 0.0380882
R36617 DVDD.n16604 DVDD.n2227 0.0380882
R36618 DVDD.n16608 DVDD.n16604 0.0380882
R36619 DVDD.n16612 DVDD.n16608 0.0380882
R36620 DVDD.n16612 DVDD.n2225 0.0380882
R36621 DVDD.n16616 DVDD.n2225 0.0380882
R36622 DVDD.n16620 DVDD.n16616 0.0380882
R36623 DVDD.n16624 DVDD.n16620 0.0380882
R36624 DVDD.n16624 DVDD.n2223 0.0380882
R36625 DVDD.n16628 DVDD.n2223 0.0380882
R36626 DVDD.n16632 DVDD.n16628 0.0380882
R36627 DVDD.n16636 DVDD.n16632 0.0380882
R36628 DVDD.n16636 DVDD.n2221 0.0380882
R36629 DVDD.n16640 DVDD.n2221 0.0380882
R36630 DVDD.n16644 DVDD.n16640 0.0380882
R36631 DVDD.n16648 DVDD.n16644 0.0380882
R36632 DVDD.n16648 DVDD.n2219 0.0380882
R36633 DVDD.n16652 DVDD.n2219 0.0380882
R36634 DVDD.n16656 DVDD.n16652 0.0380882
R36635 DVDD.n16660 DVDD.n16656 0.0380882
R36636 DVDD.n16660 DVDD.n2217 0.0380882
R36637 DVDD.n16664 DVDD.n2217 0.0380882
R36638 DVDD.n16668 DVDD.n16664 0.0380882
R36639 DVDD.n16672 DVDD.n16668 0.0380882
R36640 DVDD.n16672 DVDD.n2215 0.0380882
R36641 DVDD.n16676 DVDD.n2215 0.0380882
R36642 DVDD.n16680 DVDD.n16676 0.0380882
R36643 DVDD.n16684 DVDD.n16680 0.0380882
R36644 DVDD.n16684 DVDD.n2213 0.0380882
R36645 DVDD.n16688 DVDD.n2213 0.0380882
R36646 DVDD.n16692 DVDD.n16688 0.0380882
R36647 DVDD.n16696 DVDD.n16692 0.0380882
R36648 DVDD.n16696 DVDD.n2211 0.0380882
R36649 DVDD.n16700 DVDD.n2211 0.0380882
R36650 DVDD.n16700 DVDD.n2209 0.0380882
R36651 DVDD.n2151 DVDD.n1817 0.0380882
R36652 DVDD.n2151 DVDD.n2150 0.0380882
R36653 DVDD.n2150 DVDD.n2149 0.0380882
R36654 DVDD.n2149 DVDD.n1867 0.0380882
R36655 DVDD.n2139 DVDD.n1867 0.0380882
R36656 DVDD.n2139 DVDD.n2138 0.0380882
R36657 DVDD.n2138 DVDD.n2137 0.0380882
R36658 DVDD.n2137 DVDD.n1869 0.0380882
R36659 DVDD.n2127 DVDD.n1869 0.0380882
R36660 DVDD.n2127 DVDD.n2126 0.0380882
R36661 DVDD.n2126 DVDD.n2125 0.0380882
R36662 DVDD.n2125 DVDD.n1871 0.0380882
R36663 DVDD.n2115 DVDD.n1871 0.0380882
R36664 DVDD.n2115 DVDD.n2114 0.0380882
R36665 DVDD.n2114 DVDD.n2113 0.0380882
R36666 DVDD.n2113 DVDD.n1873 0.0380882
R36667 DVDD.n2103 DVDD.n1873 0.0380882
R36668 DVDD.n2103 DVDD.n2102 0.0380882
R36669 DVDD.n2102 DVDD.n2101 0.0380882
R36670 DVDD.n2101 DVDD.n1875 0.0380882
R36671 DVDD.n2091 DVDD.n1875 0.0380882
R36672 DVDD.n2091 DVDD.n2090 0.0380882
R36673 DVDD.n2090 DVDD.n2089 0.0380882
R36674 DVDD.n2089 DVDD.n1877 0.0380882
R36675 DVDD.n2079 DVDD.n1877 0.0380882
R36676 DVDD.n2079 DVDD.n2078 0.0380882
R36677 DVDD.n2078 DVDD.n2077 0.0380882
R36678 DVDD.n2077 DVDD.n1879 0.0380882
R36679 DVDD.n2067 DVDD.n1879 0.0380882
R36680 DVDD.n2067 DVDD.n2066 0.0380882
R36681 DVDD.n2066 DVDD.n2065 0.0380882
R36682 DVDD.n2065 DVDD.n1881 0.0380882
R36683 DVDD.n2055 DVDD.n1881 0.0380882
R36684 DVDD.n2055 DVDD.n2054 0.0380882
R36685 DVDD.n2054 DVDD.n2053 0.0380882
R36686 DVDD.n2053 DVDD.n1883 0.0380882
R36687 DVDD.n2043 DVDD.n1883 0.0380882
R36688 DVDD.n2043 DVDD.n2042 0.0380882
R36689 DVDD.n2042 DVDD.n2041 0.0380882
R36690 DVDD.n2041 DVDD.n1885 0.0380882
R36691 DVDD.n2031 DVDD.n1885 0.0380882
R36692 DVDD.n2031 DVDD.n2030 0.0380882
R36693 DVDD.n2030 DVDD.n2029 0.0380882
R36694 DVDD.n2029 DVDD.n1887 0.0380882
R36695 DVDD.n2019 DVDD.n1887 0.0380882
R36696 DVDD.n2019 DVDD.n2018 0.0380882
R36697 DVDD.n2018 DVDD.n2017 0.0380882
R36698 DVDD.n2017 DVDD.n1889 0.0380882
R36699 DVDD.n2007 DVDD.n1889 0.0380882
R36700 DVDD.n2007 DVDD.n2006 0.0380882
R36701 DVDD.n2006 DVDD.n2005 0.0380882
R36702 DVDD.n2005 DVDD.n1891 0.0380882
R36703 DVDD.n1995 DVDD.n1891 0.0380882
R36704 DVDD.n1995 DVDD.n1994 0.0380882
R36705 DVDD.n1994 DVDD.n1993 0.0380882
R36706 DVDD.n1993 DVDD.n1893 0.0380882
R36707 DVDD.n1983 DVDD.n1893 0.0380882
R36708 DVDD.n1983 DVDD.n1982 0.0380882
R36709 DVDD.n1982 DVDD.n1981 0.0380882
R36710 DVDD.n1981 DVDD.n1895 0.0380882
R36711 DVDD.n1971 DVDD.n1895 0.0380882
R36712 DVDD.n1971 DVDD.n1970 0.0380882
R36713 DVDD.n1970 DVDD.n1969 0.0380882
R36714 DVDD.n1969 DVDD.n1897 0.0380882
R36715 DVDD.n1959 DVDD.n1897 0.0380882
R36716 DVDD.n1959 DVDD.n1958 0.0380882
R36717 DVDD.n1958 DVDD.n1957 0.0380882
R36718 DVDD.n1957 DVDD.n1899 0.0380882
R36719 DVDD.n1947 DVDD.n1899 0.0380882
R36720 DVDD.n1947 DVDD.n1946 0.0380882
R36721 DVDD.n1946 DVDD.n1945 0.0380882
R36722 DVDD.n1945 DVDD.n1901 0.0380882
R36723 DVDD.n1935 DVDD.n1901 0.0380882
R36724 DVDD.n1935 DVDD.n1934 0.0380882
R36725 DVDD.n1934 DVDD.n1933 0.0380882
R36726 DVDD.n1933 DVDD.n1903 0.0380882
R36727 DVDD.n1923 DVDD.n1903 0.0380882
R36728 DVDD.n1923 DVDD.n1922 0.0380882
R36729 DVDD.n1922 DVDD.n1921 0.0380882
R36730 DVDD.n1921 DVDD.n1905 0.0380882
R36731 DVDD.n1911 DVDD.n1905 0.0380882
R36732 DVDD.n1911 DVDD.n1910 0.0380882
R36733 DVDD.n1910 DVDD.n1909 0.0380882
R36734 DVDD.n2153 DVDD.n2152 0.0380882
R36735 DVDD.n2152 DVDD.n1866 0.0380882
R36736 DVDD.n2148 DVDD.n1866 0.0380882
R36737 DVDD.n2148 DVDD.n2144 0.0380882
R36738 DVDD.n2144 DVDD.n2143 0.0380882
R36739 DVDD.n2143 DVDD.n1868 0.0380882
R36740 DVDD.n2136 DVDD.n1868 0.0380882
R36741 DVDD.n2136 DVDD.n2132 0.0380882
R36742 DVDD.n2132 DVDD.n2131 0.0380882
R36743 DVDD.n2131 DVDD.n1870 0.0380882
R36744 DVDD.n2124 DVDD.n1870 0.0380882
R36745 DVDD.n2124 DVDD.n2120 0.0380882
R36746 DVDD.n2120 DVDD.n2119 0.0380882
R36747 DVDD.n2119 DVDD.n1872 0.0380882
R36748 DVDD.n2112 DVDD.n1872 0.0380882
R36749 DVDD.n2112 DVDD.n2108 0.0380882
R36750 DVDD.n2108 DVDD.n2107 0.0380882
R36751 DVDD.n2107 DVDD.n1874 0.0380882
R36752 DVDD.n2100 DVDD.n1874 0.0380882
R36753 DVDD.n2100 DVDD.n2096 0.0380882
R36754 DVDD.n2096 DVDD.n2095 0.0380882
R36755 DVDD.n2095 DVDD.n1876 0.0380882
R36756 DVDD.n2088 DVDD.n1876 0.0380882
R36757 DVDD.n2088 DVDD.n2084 0.0380882
R36758 DVDD.n2084 DVDD.n2083 0.0380882
R36759 DVDD.n2083 DVDD.n1878 0.0380882
R36760 DVDD.n2076 DVDD.n1878 0.0380882
R36761 DVDD.n2076 DVDD.n2072 0.0380882
R36762 DVDD.n2072 DVDD.n2071 0.0380882
R36763 DVDD.n2071 DVDD.n1880 0.0380882
R36764 DVDD.n2064 DVDD.n1880 0.0380882
R36765 DVDD.n2064 DVDD.n2060 0.0380882
R36766 DVDD.n2060 DVDD.n2059 0.0380882
R36767 DVDD.n2059 DVDD.n1882 0.0380882
R36768 DVDD.n2052 DVDD.n1882 0.0380882
R36769 DVDD.n2052 DVDD.n2048 0.0380882
R36770 DVDD.n2048 DVDD.n2047 0.0380882
R36771 DVDD.n2047 DVDD.n1884 0.0380882
R36772 DVDD.n2040 DVDD.n1884 0.0380882
R36773 DVDD.n2040 DVDD.n2036 0.0380882
R36774 DVDD.n2036 DVDD.n2035 0.0380882
R36775 DVDD.n2035 DVDD.n1886 0.0380882
R36776 DVDD.n2028 DVDD.n1886 0.0380882
R36777 DVDD.n2028 DVDD.n2024 0.0380882
R36778 DVDD.n2024 DVDD.n2023 0.0380882
R36779 DVDD.n2023 DVDD.n1888 0.0380882
R36780 DVDD.n2016 DVDD.n1888 0.0380882
R36781 DVDD.n2016 DVDD.n2012 0.0380882
R36782 DVDD.n2012 DVDD.n2011 0.0380882
R36783 DVDD.n2011 DVDD.n1890 0.0380882
R36784 DVDD.n2004 DVDD.n1890 0.0380882
R36785 DVDD.n2004 DVDD.n2000 0.0380882
R36786 DVDD.n2000 DVDD.n1999 0.0380882
R36787 DVDD.n1999 DVDD.n1892 0.0380882
R36788 DVDD.n1992 DVDD.n1892 0.0380882
R36789 DVDD.n1992 DVDD.n1988 0.0380882
R36790 DVDD.n1988 DVDD.n1987 0.0380882
R36791 DVDD.n1987 DVDD.n1894 0.0380882
R36792 DVDD.n1980 DVDD.n1894 0.0380882
R36793 DVDD.n1980 DVDD.n1976 0.0380882
R36794 DVDD.n1976 DVDD.n1975 0.0380882
R36795 DVDD.n1975 DVDD.n1896 0.0380882
R36796 DVDD.n1968 DVDD.n1896 0.0380882
R36797 DVDD.n1968 DVDD.n1964 0.0380882
R36798 DVDD.n1964 DVDD.n1963 0.0380882
R36799 DVDD.n1963 DVDD.n1898 0.0380882
R36800 DVDD.n1956 DVDD.n1898 0.0380882
R36801 DVDD.n1956 DVDD.n1952 0.0380882
R36802 DVDD.n1952 DVDD.n1951 0.0380882
R36803 DVDD.n1951 DVDD.n1900 0.0380882
R36804 DVDD.n1944 DVDD.n1900 0.0380882
R36805 DVDD.n1944 DVDD.n1940 0.0380882
R36806 DVDD.n1940 DVDD.n1939 0.0380882
R36807 DVDD.n1939 DVDD.n1902 0.0380882
R36808 DVDD.n1932 DVDD.n1902 0.0380882
R36809 DVDD.n1932 DVDD.n1928 0.0380882
R36810 DVDD.n1928 DVDD.n1927 0.0380882
R36811 DVDD.n1927 DVDD.n1904 0.0380882
R36812 DVDD.n1920 DVDD.n1904 0.0380882
R36813 DVDD.n1920 DVDD.n1916 0.0380882
R36814 DVDD.n1916 DVDD.n1915 0.0380882
R36815 DVDD.n1915 DVDD.n1906 0.0380882
R36816 DVDD.n1908 DVDD.n1906 0.0380882
R36817 DVDD.n16747 DVDD.n16746 0.0380882
R36818 DVDD.n16748 DVDD.n16747 0.0380882
R36819 DVDD.n16748 DVDD.n1797 0.0380882
R36820 DVDD.n16758 DVDD.n1797 0.0380882
R36821 DVDD.n16759 DVDD.n16758 0.0380882
R36822 DVDD.n16760 DVDD.n16759 0.0380882
R36823 DVDD.n16760 DVDD.n1795 0.0380882
R36824 DVDD.n16770 DVDD.n1795 0.0380882
R36825 DVDD.n16771 DVDD.n16770 0.0380882
R36826 DVDD.n16772 DVDD.n16771 0.0380882
R36827 DVDD.n16772 DVDD.n1793 0.0380882
R36828 DVDD.n16782 DVDD.n1793 0.0380882
R36829 DVDD.n16783 DVDD.n16782 0.0380882
R36830 DVDD.n16784 DVDD.n16783 0.0380882
R36831 DVDD.n16784 DVDD.n1791 0.0380882
R36832 DVDD.n16794 DVDD.n1791 0.0380882
R36833 DVDD.n16795 DVDD.n16794 0.0380882
R36834 DVDD.n16796 DVDD.n16795 0.0380882
R36835 DVDD.n16796 DVDD.n1789 0.0380882
R36836 DVDD.n16806 DVDD.n1789 0.0380882
R36837 DVDD.n16807 DVDD.n16806 0.0380882
R36838 DVDD.n16808 DVDD.n16807 0.0380882
R36839 DVDD.n16808 DVDD.n1787 0.0380882
R36840 DVDD.n16818 DVDD.n1787 0.0380882
R36841 DVDD.n16819 DVDD.n16818 0.0380882
R36842 DVDD.n16820 DVDD.n16819 0.0380882
R36843 DVDD.n16820 DVDD.n1785 0.0380882
R36844 DVDD.n16830 DVDD.n1785 0.0380882
R36845 DVDD.n16831 DVDD.n16830 0.0380882
R36846 DVDD.n16832 DVDD.n16831 0.0380882
R36847 DVDD.n16832 DVDD.n1783 0.0380882
R36848 DVDD.n16842 DVDD.n1783 0.0380882
R36849 DVDD.n16843 DVDD.n16842 0.0380882
R36850 DVDD.n16844 DVDD.n16843 0.0380882
R36851 DVDD.n16844 DVDD.n1781 0.0380882
R36852 DVDD.n16854 DVDD.n1781 0.0380882
R36853 DVDD.n16855 DVDD.n16854 0.0380882
R36854 DVDD.n16856 DVDD.n16855 0.0380882
R36855 DVDD.n16856 DVDD.n1779 0.0380882
R36856 DVDD.n16866 DVDD.n1779 0.0380882
R36857 DVDD.n16867 DVDD.n16866 0.0380882
R36858 DVDD.n16868 DVDD.n16867 0.0380882
R36859 DVDD.n16868 DVDD.n1777 0.0380882
R36860 DVDD.n16878 DVDD.n1777 0.0380882
R36861 DVDD.n16879 DVDD.n16878 0.0380882
R36862 DVDD.n16880 DVDD.n16879 0.0380882
R36863 DVDD.n16880 DVDD.n1775 0.0380882
R36864 DVDD.n16890 DVDD.n1775 0.0380882
R36865 DVDD.n16891 DVDD.n16890 0.0380882
R36866 DVDD.n16892 DVDD.n16891 0.0380882
R36867 DVDD.n16892 DVDD.n1773 0.0380882
R36868 DVDD.n16902 DVDD.n1773 0.0380882
R36869 DVDD.n16903 DVDD.n16902 0.0380882
R36870 DVDD.n16904 DVDD.n16903 0.0380882
R36871 DVDD.n16904 DVDD.n1771 0.0380882
R36872 DVDD.n16914 DVDD.n1771 0.0380882
R36873 DVDD.n16915 DVDD.n16914 0.0380882
R36874 DVDD.n16916 DVDD.n16915 0.0380882
R36875 DVDD.n16916 DVDD.n1769 0.0380882
R36876 DVDD.n16926 DVDD.n1769 0.0380882
R36877 DVDD.n16927 DVDD.n16926 0.0380882
R36878 DVDD.n16928 DVDD.n16927 0.0380882
R36879 DVDD.n16928 DVDD.n1767 0.0380882
R36880 DVDD.n16938 DVDD.n1767 0.0380882
R36881 DVDD.n16939 DVDD.n16938 0.0380882
R36882 DVDD.n16940 DVDD.n16939 0.0380882
R36883 DVDD.n16940 DVDD.n1765 0.0380882
R36884 DVDD.n16950 DVDD.n1765 0.0380882
R36885 DVDD.n16951 DVDD.n16950 0.0380882
R36886 DVDD.n16952 DVDD.n16951 0.0380882
R36887 DVDD.n16952 DVDD.n1763 0.0380882
R36888 DVDD.n16962 DVDD.n1763 0.0380882
R36889 DVDD.n16963 DVDD.n16962 0.0380882
R36890 DVDD.n16964 DVDD.n16963 0.0380882
R36891 DVDD.n16964 DVDD.n1761 0.0380882
R36892 DVDD.n16974 DVDD.n1761 0.0380882
R36893 DVDD.n16975 DVDD.n16974 0.0380882
R36894 DVDD.n16976 DVDD.n16975 0.0380882
R36895 DVDD.n16976 DVDD.n1759 0.0380882
R36896 DVDD.n16986 DVDD.n1759 0.0380882
R36897 DVDD.n16987 DVDD.n16986 0.0380882
R36898 DVDD.n16989 DVDD.n16987 0.0380882
R36899 DVDD.n16989 DVDD.n16988 0.0380882
R36900 DVDD.n16745 DVDD.n1800 0.0380882
R36901 DVDD.n16749 DVDD.n1800 0.0380882
R36902 DVDD.n16753 DVDD.n16749 0.0380882
R36903 DVDD.n16757 DVDD.n16753 0.0380882
R36904 DVDD.n16757 DVDD.n1796 0.0380882
R36905 DVDD.n16761 DVDD.n1796 0.0380882
R36906 DVDD.n16765 DVDD.n16761 0.0380882
R36907 DVDD.n16769 DVDD.n16765 0.0380882
R36908 DVDD.n16769 DVDD.n1794 0.0380882
R36909 DVDD.n16773 DVDD.n1794 0.0380882
R36910 DVDD.n16777 DVDD.n16773 0.0380882
R36911 DVDD.n16781 DVDD.n16777 0.0380882
R36912 DVDD.n16781 DVDD.n1792 0.0380882
R36913 DVDD.n16785 DVDD.n1792 0.0380882
R36914 DVDD.n16789 DVDD.n16785 0.0380882
R36915 DVDD.n16793 DVDD.n16789 0.0380882
R36916 DVDD.n16793 DVDD.n1790 0.0380882
R36917 DVDD.n16797 DVDD.n1790 0.0380882
R36918 DVDD.n16801 DVDD.n16797 0.0380882
R36919 DVDD.n16805 DVDD.n16801 0.0380882
R36920 DVDD.n16805 DVDD.n1788 0.0380882
R36921 DVDD.n16809 DVDD.n1788 0.0380882
R36922 DVDD.n16813 DVDD.n16809 0.0380882
R36923 DVDD.n16817 DVDD.n16813 0.0380882
R36924 DVDD.n16817 DVDD.n1786 0.0380882
R36925 DVDD.n16821 DVDD.n1786 0.0380882
R36926 DVDD.n16825 DVDD.n16821 0.0380882
R36927 DVDD.n16829 DVDD.n16825 0.0380882
R36928 DVDD.n16829 DVDD.n1784 0.0380882
R36929 DVDD.n16833 DVDD.n1784 0.0380882
R36930 DVDD.n16837 DVDD.n16833 0.0380882
R36931 DVDD.n16841 DVDD.n16837 0.0380882
R36932 DVDD.n16841 DVDD.n1782 0.0380882
R36933 DVDD.n16845 DVDD.n1782 0.0380882
R36934 DVDD.n16849 DVDD.n16845 0.0380882
R36935 DVDD.n16853 DVDD.n16849 0.0380882
R36936 DVDD.n16853 DVDD.n1780 0.0380882
R36937 DVDD.n16857 DVDD.n1780 0.0380882
R36938 DVDD.n16861 DVDD.n16857 0.0380882
R36939 DVDD.n16865 DVDD.n16861 0.0380882
R36940 DVDD.n16865 DVDD.n1778 0.0380882
R36941 DVDD.n16869 DVDD.n1778 0.0380882
R36942 DVDD.n16873 DVDD.n16869 0.0380882
R36943 DVDD.n16877 DVDD.n16873 0.0380882
R36944 DVDD.n16877 DVDD.n1776 0.0380882
R36945 DVDD.n16881 DVDD.n1776 0.0380882
R36946 DVDD.n16885 DVDD.n16881 0.0380882
R36947 DVDD.n16889 DVDD.n16885 0.0380882
R36948 DVDD.n16889 DVDD.n1774 0.0380882
R36949 DVDD.n16893 DVDD.n1774 0.0380882
R36950 DVDD.n16897 DVDD.n16893 0.0380882
R36951 DVDD.n16901 DVDD.n16897 0.0380882
R36952 DVDD.n16901 DVDD.n1772 0.0380882
R36953 DVDD.n16905 DVDD.n1772 0.0380882
R36954 DVDD.n16909 DVDD.n16905 0.0380882
R36955 DVDD.n16913 DVDD.n16909 0.0380882
R36956 DVDD.n16913 DVDD.n1770 0.0380882
R36957 DVDD.n16917 DVDD.n1770 0.0380882
R36958 DVDD.n16921 DVDD.n16917 0.0380882
R36959 DVDD.n16925 DVDD.n16921 0.0380882
R36960 DVDD.n16925 DVDD.n1768 0.0380882
R36961 DVDD.n16929 DVDD.n1768 0.0380882
R36962 DVDD.n16933 DVDD.n16929 0.0380882
R36963 DVDD.n16937 DVDD.n16933 0.0380882
R36964 DVDD.n16937 DVDD.n1766 0.0380882
R36965 DVDD.n16941 DVDD.n1766 0.0380882
R36966 DVDD.n16945 DVDD.n16941 0.0380882
R36967 DVDD.n16949 DVDD.n16945 0.0380882
R36968 DVDD.n16949 DVDD.n1764 0.0380882
R36969 DVDD.n16953 DVDD.n1764 0.0380882
R36970 DVDD.n16957 DVDD.n16953 0.0380882
R36971 DVDD.n16961 DVDD.n16957 0.0380882
R36972 DVDD.n16961 DVDD.n1762 0.0380882
R36973 DVDD.n16965 DVDD.n1762 0.0380882
R36974 DVDD.n16969 DVDD.n16965 0.0380882
R36975 DVDD.n16973 DVDD.n16969 0.0380882
R36976 DVDD.n16973 DVDD.n1760 0.0380882
R36977 DVDD.n16977 DVDD.n1760 0.0380882
R36978 DVDD.n16981 DVDD.n16977 0.0380882
R36979 DVDD.n16985 DVDD.n16981 0.0380882
R36980 DVDD.n16985 DVDD.n1758 0.0380882
R36981 DVDD.n16990 DVDD.n1758 0.0380882
R36982 DVDD.n16990 DVDD.n1756 0.0380882
R36983 DVDD.n17015 DVDD.n17014 0.0380882
R36984 DVDD.n17016 DVDD.n17015 0.0380882
R36985 DVDD.n17016 DVDD.n1698 0.0380882
R36986 DVDD.n17026 DVDD.n1698 0.0380882
R36987 DVDD.n17027 DVDD.n17026 0.0380882
R36988 DVDD.n17028 DVDD.n17027 0.0380882
R36989 DVDD.n17028 DVDD.n1696 0.0380882
R36990 DVDD.n17038 DVDD.n1696 0.0380882
R36991 DVDD.n17039 DVDD.n17038 0.0380882
R36992 DVDD.n17040 DVDD.n17039 0.0380882
R36993 DVDD.n17040 DVDD.n1694 0.0380882
R36994 DVDD.n17050 DVDD.n1694 0.0380882
R36995 DVDD.n17051 DVDD.n17050 0.0380882
R36996 DVDD.n17052 DVDD.n17051 0.0380882
R36997 DVDD.n17052 DVDD.n1692 0.0380882
R36998 DVDD.n17062 DVDD.n1692 0.0380882
R36999 DVDD.n17063 DVDD.n17062 0.0380882
R37000 DVDD.n17064 DVDD.n17063 0.0380882
R37001 DVDD.n17064 DVDD.n1690 0.0380882
R37002 DVDD.n17074 DVDD.n1690 0.0380882
R37003 DVDD.n17075 DVDD.n17074 0.0380882
R37004 DVDD.n17076 DVDD.n17075 0.0380882
R37005 DVDD.n17076 DVDD.n1688 0.0380882
R37006 DVDD.n17086 DVDD.n1688 0.0380882
R37007 DVDD.n17087 DVDD.n17086 0.0380882
R37008 DVDD.n17088 DVDD.n17087 0.0380882
R37009 DVDD.n17088 DVDD.n1686 0.0380882
R37010 DVDD.n17098 DVDD.n1686 0.0380882
R37011 DVDD.n17099 DVDD.n17098 0.0380882
R37012 DVDD.n17100 DVDD.n17099 0.0380882
R37013 DVDD.n17100 DVDD.n1684 0.0380882
R37014 DVDD.n17110 DVDD.n1684 0.0380882
R37015 DVDD.n17111 DVDD.n17110 0.0380882
R37016 DVDD.n17112 DVDD.n17111 0.0380882
R37017 DVDD.n17112 DVDD.n1682 0.0380882
R37018 DVDD.n17122 DVDD.n1682 0.0380882
R37019 DVDD.n17123 DVDD.n17122 0.0380882
R37020 DVDD.n17124 DVDD.n17123 0.0380882
R37021 DVDD.n17124 DVDD.n1680 0.0380882
R37022 DVDD.n17134 DVDD.n1680 0.0380882
R37023 DVDD.n17135 DVDD.n17134 0.0380882
R37024 DVDD.n17136 DVDD.n17135 0.0380882
R37025 DVDD.n17136 DVDD.n1678 0.0380882
R37026 DVDD.n17146 DVDD.n1678 0.0380882
R37027 DVDD.n17147 DVDD.n17146 0.0380882
R37028 DVDD.n17148 DVDD.n17147 0.0380882
R37029 DVDD.n17148 DVDD.n1676 0.0380882
R37030 DVDD.n17158 DVDD.n1676 0.0380882
R37031 DVDD.n17159 DVDD.n17158 0.0380882
R37032 DVDD.n17160 DVDD.n17159 0.0380882
R37033 DVDD.n17160 DVDD.n1674 0.0380882
R37034 DVDD.n17170 DVDD.n1674 0.0380882
R37035 DVDD.n17171 DVDD.n17170 0.0380882
R37036 DVDD.n17172 DVDD.n17171 0.0380882
R37037 DVDD.n17172 DVDD.n1672 0.0380882
R37038 DVDD.n17182 DVDD.n1672 0.0380882
R37039 DVDD.n17183 DVDD.n17182 0.0380882
R37040 DVDD.n17184 DVDD.n17183 0.0380882
R37041 DVDD.n17184 DVDD.n1670 0.0380882
R37042 DVDD.n17194 DVDD.n1670 0.0380882
R37043 DVDD.n17195 DVDD.n17194 0.0380882
R37044 DVDD.n17196 DVDD.n17195 0.0380882
R37045 DVDD.n17196 DVDD.n1668 0.0380882
R37046 DVDD.n17206 DVDD.n1668 0.0380882
R37047 DVDD.n17207 DVDD.n17206 0.0380882
R37048 DVDD.n17208 DVDD.n17207 0.0380882
R37049 DVDD.n17208 DVDD.n1666 0.0380882
R37050 DVDD.n17218 DVDD.n1666 0.0380882
R37051 DVDD.n17219 DVDD.n17218 0.0380882
R37052 DVDD.n17220 DVDD.n17219 0.0380882
R37053 DVDD.n17220 DVDD.n1664 0.0380882
R37054 DVDD.n17230 DVDD.n1664 0.0380882
R37055 DVDD.n17231 DVDD.n17230 0.0380882
R37056 DVDD.n17232 DVDD.n17231 0.0380882
R37057 DVDD.n17232 DVDD.n1662 0.0380882
R37058 DVDD.n17242 DVDD.n1662 0.0380882
R37059 DVDD.n17243 DVDD.n17242 0.0380882
R37060 DVDD.n17244 DVDD.n17243 0.0380882
R37061 DVDD.n17244 DVDD.n1660 0.0380882
R37062 DVDD.n17254 DVDD.n1660 0.0380882
R37063 DVDD.n17255 DVDD.n17254 0.0380882
R37064 DVDD.n17257 DVDD.n17255 0.0380882
R37065 DVDD.n17257 DVDD.n17256 0.0380882
R37066 DVDD.n17013 DVDD.n1701 0.0380882
R37067 DVDD.n17017 DVDD.n1701 0.0380882
R37068 DVDD.n17021 DVDD.n17017 0.0380882
R37069 DVDD.n17025 DVDD.n17021 0.0380882
R37070 DVDD.n17025 DVDD.n1697 0.0380882
R37071 DVDD.n17029 DVDD.n1697 0.0380882
R37072 DVDD.n17033 DVDD.n17029 0.0380882
R37073 DVDD.n17037 DVDD.n17033 0.0380882
R37074 DVDD.n17037 DVDD.n1695 0.0380882
R37075 DVDD.n17041 DVDD.n1695 0.0380882
R37076 DVDD.n17045 DVDD.n17041 0.0380882
R37077 DVDD.n17049 DVDD.n17045 0.0380882
R37078 DVDD.n17049 DVDD.n1693 0.0380882
R37079 DVDD.n17053 DVDD.n1693 0.0380882
R37080 DVDD.n17057 DVDD.n17053 0.0380882
R37081 DVDD.n17061 DVDD.n17057 0.0380882
R37082 DVDD.n17061 DVDD.n1691 0.0380882
R37083 DVDD.n17065 DVDD.n1691 0.0380882
R37084 DVDD.n17069 DVDD.n17065 0.0380882
R37085 DVDD.n17073 DVDD.n17069 0.0380882
R37086 DVDD.n17073 DVDD.n1689 0.0380882
R37087 DVDD.n17077 DVDD.n1689 0.0380882
R37088 DVDD.n17081 DVDD.n17077 0.0380882
R37089 DVDD.n17085 DVDD.n17081 0.0380882
R37090 DVDD.n17085 DVDD.n1687 0.0380882
R37091 DVDD.n17089 DVDD.n1687 0.0380882
R37092 DVDD.n17093 DVDD.n17089 0.0380882
R37093 DVDD.n17097 DVDD.n17093 0.0380882
R37094 DVDD.n17097 DVDD.n1685 0.0380882
R37095 DVDD.n17101 DVDD.n1685 0.0380882
R37096 DVDD.n17105 DVDD.n17101 0.0380882
R37097 DVDD.n17109 DVDD.n17105 0.0380882
R37098 DVDD.n17109 DVDD.n1683 0.0380882
R37099 DVDD.n17113 DVDD.n1683 0.0380882
R37100 DVDD.n17117 DVDD.n17113 0.0380882
R37101 DVDD.n17121 DVDD.n17117 0.0380882
R37102 DVDD.n17121 DVDD.n1681 0.0380882
R37103 DVDD.n17125 DVDD.n1681 0.0380882
R37104 DVDD.n17129 DVDD.n17125 0.0380882
R37105 DVDD.n17133 DVDD.n17129 0.0380882
R37106 DVDD.n17133 DVDD.n1679 0.0380882
R37107 DVDD.n17137 DVDD.n1679 0.0380882
R37108 DVDD.n17141 DVDD.n17137 0.0380882
R37109 DVDD.n17145 DVDD.n17141 0.0380882
R37110 DVDD.n17145 DVDD.n1677 0.0380882
R37111 DVDD.n17149 DVDD.n1677 0.0380882
R37112 DVDD.n17153 DVDD.n17149 0.0380882
R37113 DVDD.n17157 DVDD.n17153 0.0380882
R37114 DVDD.n17157 DVDD.n1675 0.0380882
R37115 DVDD.n17161 DVDD.n1675 0.0380882
R37116 DVDD.n17165 DVDD.n17161 0.0380882
R37117 DVDD.n17169 DVDD.n17165 0.0380882
R37118 DVDD.n17169 DVDD.n1673 0.0380882
R37119 DVDD.n17173 DVDD.n1673 0.0380882
R37120 DVDD.n17177 DVDD.n17173 0.0380882
R37121 DVDD.n17181 DVDD.n17177 0.0380882
R37122 DVDD.n17181 DVDD.n1671 0.0380882
R37123 DVDD.n17185 DVDD.n1671 0.0380882
R37124 DVDD.n17189 DVDD.n17185 0.0380882
R37125 DVDD.n17193 DVDD.n17189 0.0380882
R37126 DVDD.n17193 DVDD.n1669 0.0380882
R37127 DVDD.n17197 DVDD.n1669 0.0380882
R37128 DVDD.n17201 DVDD.n17197 0.0380882
R37129 DVDD.n17205 DVDD.n17201 0.0380882
R37130 DVDD.n17205 DVDD.n1667 0.0380882
R37131 DVDD.n17209 DVDD.n1667 0.0380882
R37132 DVDD.n17213 DVDD.n17209 0.0380882
R37133 DVDD.n17217 DVDD.n17213 0.0380882
R37134 DVDD.n17217 DVDD.n1665 0.0380882
R37135 DVDD.n17221 DVDD.n1665 0.0380882
R37136 DVDD.n17225 DVDD.n17221 0.0380882
R37137 DVDD.n17229 DVDD.n17225 0.0380882
R37138 DVDD.n17229 DVDD.n1663 0.0380882
R37139 DVDD.n17233 DVDD.n1663 0.0380882
R37140 DVDD.n17237 DVDD.n17233 0.0380882
R37141 DVDD.n17241 DVDD.n17237 0.0380882
R37142 DVDD.n17241 DVDD.n1661 0.0380882
R37143 DVDD.n17245 DVDD.n1661 0.0380882
R37144 DVDD.n17249 DVDD.n17245 0.0380882
R37145 DVDD.n17253 DVDD.n17249 0.0380882
R37146 DVDD.n17253 DVDD.n1659 0.0380882
R37147 DVDD.n17258 DVDD.n1659 0.0380882
R37148 DVDD.n17258 DVDD.n1657 0.0380882
R37149 DVDD.n6511 DVDD.n6396 0.0380882
R37150 DVDD.n6512 DVDD.n6511 0.0380882
R37151 DVDD.n6513 DVDD.n6512 0.0380882
R37152 DVDD.n6513 DVDD.n6505 0.0380882
R37153 DVDD.n6520 DVDD.n6505 0.0380882
R37154 DVDD.n6521 DVDD.n6520 0.0380882
R37155 DVDD.n6522 DVDD.n6521 0.0380882
R37156 DVDD.n6522 DVDD.n6502 0.0380882
R37157 DVDD.n6529 DVDD.n6502 0.0380882
R37158 DVDD.n6530 DVDD.n6529 0.0380882
R37159 DVDD.n6531 DVDD.n6530 0.0380882
R37160 DVDD.n6531 DVDD.n6499 0.0380882
R37161 DVDD.n6538 DVDD.n6499 0.0380882
R37162 DVDD.n6539 DVDD.n6538 0.0380882
R37163 DVDD.n6540 DVDD.n6539 0.0380882
R37164 DVDD.n6540 DVDD.n6496 0.0380882
R37165 DVDD.n6547 DVDD.n6496 0.0380882
R37166 DVDD.n6548 DVDD.n6547 0.0380882
R37167 DVDD.n6549 DVDD.n6548 0.0380882
R37168 DVDD.n6549 DVDD.n6493 0.0380882
R37169 DVDD.n6556 DVDD.n6493 0.0380882
R37170 DVDD.n6557 DVDD.n6556 0.0380882
R37171 DVDD.n6558 DVDD.n6557 0.0380882
R37172 DVDD.n6558 DVDD.n6490 0.0380882
R37173 DVDD.n6565 DVDD.n6490 0.0380882
R37174 DVDD.n6566 DVDD.n6565 0.0380882
R37175 DVDD.n6567 DVDD.n6566 0.0380882
R37176 DVDD.n6567 DVDD.n6487 0.0380882
R37177 DVDD.n6574 DVDD.n6487 0.0380882
R37178 DVDD.n6575 DVDD.n6574 0.0380882
R37179 DVDD.n6576 DVDD.n6575 0.0380882
R37180 DVDD.n6576 DVDD.n6484 0.0380882
R37181 DVDD.n6583 DVDD.n6484 0.0380882
R37182 DVDD.n6584 DVDD.n6583 0.0380882
R37183 DVDD.n6585 DVDD.n6584 0.0380882
R37184 DVDD.n6585 DVDD.n6481 0.0380882
R37185 DVDD.n6592 DVDD.n6481 0.0380882
R37186 DVDD.n6593 DVDD.n6592 0.0380882
R37187 DVDD.n6594 DVDD.n6593 0.0380882
R37188 DVDD.n6594 DVDD.n6478 0.0380882
R37189 DVDD.n6601 DVDD.n6478 0.0380882
R37190 DVDD.n6602 DVDD.n6601 0.0380882
R37191 DVDD.n6603 DVDD.n6602 0.0380882
R37192 DVDD.n6603 DVDD.n6475 0.0380882
R37193 DVDD.n6610 DVDD.n6475 0.0380882
R37194 DVDD.n6611 DVDD.n6610 0.0380882
R37195 DVDD.n6612 DVDD.n6611 0.0380882
R37196 DVDD.n6612 DVDD.n6472 0.0380882
R37197 DVDD.n6619 DVDD.n6472 0.0380882
R37198 DVDD.n6620 DVDD.n6619 0.0380882
R37199 DVDD.n6621 DVDD.n6620 0.0380882
R37200 DVDD.n6621 DVDD.n6469 0.0380882
R37201 DVDD.n6628 DVDD.n6469 0.0380882
R37202 DVDD.n6629 DVDD.n6628 0.0380882
R37203 DVDD.n6630 DVDD.n6629 0.0380882
R37204 DVDD.n6630 DVDD.n6466 0.0380882
R37205 DVDD.n6637 DVDD.n6466 0.0380882
R37206 DVDD.n6638 DVDD.n6637 0.0380882
R37207 DVDD.n6639 DVDD.n6638 0.0380882
R37208 DVDD.n6639 DVDD.n6463 0.0380882
R37209 DVDD.n6646 DVDD.n6463 0.0380882
R37210 DVDD.n6647 DVDD.n6646 0.0380882
R37211 DVDD.n6648 DVDD.n6647 0.0380882
R37212 DVDD.n6648 DVDD.n6460 0.0380882
R37213 DVDD.n6655 DVDD.n6460 0.0380882
R37214 DVDD.n6656 DVDD.n6655 0.0380882
R37215 DVDD.n6657 DVDD.n6656 0.0380882
R37216 DVDD.n6657 DVDD.n6457 0.0380882
R37217 DVDD.n6664 DVDD.n6457 0.0380882
R37218 DVDD.n6665 DVDD.n6664 0.0380882
R37219 DVDD.n6666 DVDD.n6665 0.0380882
R37220 DVDD.n6666 DVDD.n6454 0.0380882
R37221 DVDD.n6673 DVDD.n6454 0.0380882
R37222 DVDD.n6674 DVDD.n6673 0.0380882
R37223 DVDD.n6675 DVDD.n6674 0.0380882
R37224 DVDD.n6675 DVDD.n6451 0.0380882
R37225 DVDD.n6682 DVDD.n6451 0.0380882
R37226 DVDD.n6683 DVDD.n6682 0.0380882
R37227 DVDD.n6684 DVDD.n6683 0.0380882
R37228 DVDD.n6684 DVDD.n6448 0.0380882
R37229 DVDD.n6691 DVDD.n6448 0.0380882
R37230 DVDD.n6692 DVDD.n6691 0.0380882
R37231 DVDD.n6693 DVDD.n6692 0.0380882
R37232 DVDD.n6510 DVDD.n6508 0.0380882
R37233 DVDD.n6510 DVDD.n6507 0.0380882
R37234 DVDD.n6515 DVDD.n6507 0.0380882
R37235 DVDD.n6517 DVDD.n6515 0.0380882
R37236 DVDD.n6519 DVDD.n6517 0.0380882
R37237 DVDD.n6519 DVDD.n6504 0.0380882
R37238 DVDD.n6524 DVDD.n6504 0.0380882
R37239 DVDD.n6526 DVDD.n6524 0.0380882
R37240 DVDD.n6528 DVDD.n6526 0.0380882
R37241 DVDD.n6528 DVDD.n6501 0.0380882
R37242 DVDD.n6533 DVDD.n6501 0.0380882
R37243 DVDD.n6535 DVDD.n6533 0.0380882
R37244 DVDD.n6537 DVDD.n6535 0.0380882
R37245 DVDD.n6537 DVDD.n6498 0.0380882
R37246 DVDD.n6542 DVDD.n6498 0.0380882
R37247 DVDD.n6544 DVDD.n6542 0.0380882
R37248 DVDD.n6546 DVDD.n6544 0.0380882
R37249 DVDD.n6546 DVDD.n6495 0.0380882
R37250 DVDD.n6551 DVDD.n6495 0.0380882
R37251 DVDD.n6553 DVDD.n6551 0.0380882
R37252 DVDD.n6555 DVDD.n6553 0.0380882
R37253 DVDD.n6555 DVDD.n6492 0.0380882
R37254 DVDD.n6560 DVDD.n6492 0.0380882
R37255 DVDD.n6562 DVDD.n6560 0.0380882
R37256 DVDD.n6564 DVDD.n6562 0.0380882
R37257 DVDD.n6564 DVDD.n6489 0.0380882
R37258 DVDD.n6569 DVDD.n6489 0.0380882
R37259 DVDD.n6571 DVDD.n6569 0.0380882
R37260 DVDD.n6573 DVDD.n6571 0.0380882
R37261 DVDD.n6573 DVDD.n6486 0.0380882
R37262 DVDD.n6578 DVDD.n6486 0.0380882
R37263 DVDD.n6580 DVDD.n6578 0.0380882
R37264 DVDD.n6582 DVDD.n6580 0.0380882
R37265 DVDD.n6582 DVDD.n6483 0.0380882
R37266 DVDD.n6587 DVDD.n6483 0.0380882
R37267 DVDD.n6589 DVDD.n6587 0.0380882
R37268 DVDD.n6591 DVDD.n6589 0.0380882
R37269 DVDD.n6591 DVDD.n6480 0.0380882
R37270 DVDD.n6596 DVDD.n6480 0.0380882
R37271 DVDD.n6598 DVDD.n6596 0.0380882
R37272 DVDD.n6600 DVDD.n6598 0.0380882
R37273 DVDD.n6600 DVDD.n6477 0.0380882
R37274 DVDD.n6605 DVDD.n6477 0.0380882
R37275 DVDD.n6607 DVDD.n6605 0.0380882
R37276 DVDD.n6609 DVDD.n6607 0.0380882
R37277 DVDD.n6609 DVDD.n6474 0.0380882
R37278 DVDD.n6614 DVDD.n6474 0.0380882
R37279 DVDD.n6616 DVDD.n6614 0.0380882
R37280 DVDD.n6618 DVDD.n6616 0.0380882
R37281 DVDD.n6618 DVDD.n6471 0.0380882
R37282 DVDD.n6623 DVDD.n6471 0.0380882
R37283 DVDD.n6625 DVDD.n6623 0.0380882
R37284 DVDD.n6627 DVDD.n6625 0.0380882
R37285 DVDD.n6627 DVDD.n6468 0.0380882
R37286 DVDD.n6632 DVDD.n6468 0.0380882
R37287 DVDD.n6634 DVDD.n6632 0.0380882
R37288 DVDD.n6636 DVDD.n6634 0.0380882
R37289 DVDD.n6636 DVDD.n6465 0.0380882
R37290 DVDD.n6641 DVDD.n6465 0.0380882
R37291 DVDD.n6643 DVDD.n6641 0.0380882
R37292 DVDD.n6645 DVDD.n6643 0.0380882
R37293 DVDD.n6645 DVDD.n6462 0.0380882
R37294 DVDD.n6650 DVDD.n6462 0.0380882
R37295 DVDD.n6652 DVDD.n6650 0.0380882
R37296 DVDD.n6654 DVDD.n6652 0.0380882
R37297 DVDD.n6654 DVDD.n6459 0.0380882
R37298 DVDD.n6659 DVDD.n6459 0.0380882
R37299 DVDD.n6661 DVDD.n6659 0.0380882
R37300 DVDD.n6663 DVDD.n6661 0.0380882
R37301 DVDD.n6663 DVDD.n6456 0.0380882
R37302 DVDD.n6668 DVDD.n6456 0.0380882
R37303 DVDD.n6670 DVDD.n6668 0.0380882
R37304 DVDD.n6672 DVDD.n6670 0.0380882
R37305 DVDD.n6672 DVDD.n6453 0.0380882
R37306 DVDD.n6677 DVDD.n6453 0.0380882
R37307 DVDD.n6679 DVDD.n6677 0.0380882
R37308 DVDD.n6681 DVDD.n6679 0.0380882
R37309 DVDD.n6681 DVDD.n6450 0.0380882
R37310 DVDD.n6686 DVDD.n6450 0.0380882
R37311 DVDD.n6688 DVDD.n6686 0.0380882
R37312 DVDD.n6690 DVDD.n6688 0.0380882
R37313 DVDD.n6690 DVDD.n6447 0.0380882
R37314 DVDD.n6694 DVDD.n6447 0.0380882
R37315 DVDD.n6327 DVDD.n6094 0.0380882
R37316 DVDD.n6327 DVDD.n6326 0.0380882
R37317 DVDD.n6326 DVDD.n6325 0.0380882
R37318 DVDD.n6325 DVDD.n6095 0.0380882
R37319 DVDD.n6318 DVDD.n6095 0.0380882
R37320 DVDD.n6318 DVDD.n6317 0.0380882
R37321 DVDD.n6317 DVDD.n6316 0.0380882
R37322 DVDD.n6316 DVDD.n6098 0.0380882
R37323 DVDD.n6309 DVDD.n6098 0.0380882
R37324 DVDD.n6309 DVDD.n6308 0.0380882
R37325 DVDD.n6308 DVDD.n6307 0.0380882
R37326 DVDD.n6307 DVDD.n6101 0.0380882
R37327 DVDD.n6300 DVDD.n6101 0.0380882
R37328 DVDD.n6300 DVDD.n6299 0.0380882
R37329 DVDD.n6299 DVDD.n6298 0.0380882
R37330 DVDD.n6298 DVDD.n6104 0.0380882
R37331 DVDD.n6291 DVDD.n6104 0.0380882
R37332 DVDD.n6291 DVDD.n6290 0.0380882
R37333 DVDD.n6290 DVDD.n6289 0.0380882
R37334 DVDD.n6289 DVDD.n6107 0.0380882
R37335 DVDD.n6282 DVDD.n6107 0.0380882
R37336 DVDD.n6282 DVDD.n6281 0.0380882
R37337 DVDD.n6281 DVDD.n6280 0.0380882
R37338 DVDD.n6280 DVDD.n6110 0.0380882
R37339 DVDD.n6273 DVDD.n6110 0.0380882
R37340 DVDD.n6273 DVDD.n6272 0.0380882
R37341 DVDD.n6272 DVDD.n6271 0.0380882
R37342 DVDD.n6271 DVDD.n6113 0.0380882
R37343 DVDD.n6264 DVDD.n6113 0.0380882
R37344 DVDD.n6264 DVDD.n6263 0.0380882
R37345 DVDD.n6263 DVDD.n6262 0.0380882
R37346 DVDD.n6262 DVDD.n6116 0.0380882
R37347 DVDD.n6255 DVDD.n6116 0.0380882
R37348 DVDD.n6255 DVDD.n6254 0.0380882
R37349 DVDD.n6254 DVDD.n6253 0.0380882
R37350 DVDD.n6253 DVDD.n6119 0.0380882
R37351 DVDD.n6246 DVDD.n6119 0.0380882
R37352 DVDD.n6246 DVDD.n6245 0.0380882
R37353 DVDD.n6245 DVDD.n6244 0.0380882
R37354 DVDD.n6244 DVDD.n6122 0.0380882
R37355 DVDD.n6237 DVDD.n6122 0.0380882
R37356 DVDD.n6237 DVDD.n6236 0.0380882
R37357 DVDD.n6236 DVDD.n6235 0.0380882
R37358 DVDD.n6235 DVDD.n6125 0.0380882
R37359 DVDD.n6228 DVDD.n6125 0.0380882
R37360 DVDD.n6228 DVDD.n6227 0.0380882
R37361 DVDD.n6227 DVDD.n6226 0.0380882
R37362 DVDD.n6226 DVDD.n6128 0.0380882
R37363 DVDD.n6219 DVDD.n6128 0.0380882
R37364 DVDD.n6219 DVDD.n6218 0.0380882
R37365 DVDD.n6218 DVDD.n6217 0.0380882
R37366 DVDD.n6217 DVDD.n6131 0.0380882
R37367 DVDD.n6210 DVDD.n6131 0.0380882
R37368 DVDD.n6210 DVDD.n6209 0.0380882
R37369 DVDD.n6209 DVDD.n6208 0.0380882
R37370 DVDD.n6208 DVDD.n6134 0.0380882
R37371 DVDD.n6201 DVDD.n6134 0.0380882
R37372 DVDD.n6201 DVDD.n6200 0.0380882
R37373 DVDD.n6200 DVDD.n6199 0.0380882
R37374 DVDD.n6199 DVDD.n6137 0.0380882
R37375 DVDD.n6192 DVDD.n6137 0.0380882
R37376 DVDD.n6192 DVDD.n6191 0.0380882
R37377 DVDD.n6191 DVDD.n6190 0.0380882
R37378 DVDD.n6190 DVDD.n6140 0.0380882
R37379 DVDD.n6183 DVDD.n6140 0.0380882
R37380 DVDD.n6183 DVDD.n6182 0.0380882
R37381 DVDD.n6182 DVDD.n6181 0.0380882
R37382 DVDD.n6181 DVDD.n6143 0.0380882
R37383 DVDD.n6174 DVDD.n6143 0.0380882
R37384 DVDD.n6174 DVDD.n6173 0.0380882
R37385 DVDD.n6173 DVDD.n6172 0.0380882
R37386 DVDD.n6172 DVDD.n6146 0.0380882
R37387 DVDD.n6165 DVDD.n6146 0.0380882
R37388 DVDD.n6165 DVDD.n6164 0.0380882
R37389 DVDD.n6164 DVDD.n6163 0.0380882
R37390 DVDD.n6163 DVDD.n6149 0.0380882
R37391 DVDD.n6156 DVDD.n6149 0.0380882
R37392 DVDD.n6156 DVDD.n6155 0.0380882
R37393 DVDD.n6155 DVDD.n6154 0.0380882
R37394 DVDD.n6154 DVDD.n6048 0.0380882
R37395 DVDD.n6335 DVDD.n6048 0.0380882
R37396 DVDD.n6336 DVDD.n6335 0.0380882
R37397 DVDD.n6337 DVDD.n6336 0.0380882
R37398 DVDD.n6328 DVDD.n6091 0.0380882
R37399 DVDD.n6328 DVDD.n6093 0.0380882
R37400 DVDD.n6324 DVDD.n6093 0.0380882
R37401 DVDD.n6324 DVDD.n6322 0.0380882
R37402 DVDD.n6322 DVDD.n6320 0.0380882
R37403 DVDD.n6320 DVDD.n6097 0.0380882
R37404 DVDD.n6315 DVDD.n6097 0.0380882
R37405 DVDD.n6315 DVDD.n6313 0.0380882
R37406 DVDD.n6313 DVDD.n6311 0.0380882
R37407 DVDD.n6311 DVDD.n6100 0.0380882
R37408 DVDD.n6306 DVDD.n6100 0.0380882
R37409 DVDD.n6306 DVDD.n6304 0.0380882
R37410 DVDD.n6304 DVDD.n6302 0.0380882
R37411 DVDD.n6302 DVDD.n6103 0.0380882
R37412 DVDD.n6297 DVDD.n6103 0.0380882
R37413 DVDD.n6297 DVDD.n6295 0.0380882
R37414 DVDD.n6295 DVDD.n6293 0.0380882
R37415 DVDD.n6293 DVDD.n6106 0.0380882
R37416 DVDD.n6288 DVDD.n6106 0.0380882
R37417 DVDD.n6288 DVDD.n6286 0.0380882
R37418 DVDD.n6286 DVDD.n6284 0.0380882
R37419 DVDD.n6284 DVDD.n6109 0.0380882
R37420 DVDD.n6279 DVDD.n6109 0.0380882
R37421 DVDD.n6279 DVDD.n6277 0.0380882
R37422 DVDD.n6277 DVDD.n6275 0.0380882
R37423 DVDD.n6275 DVDD.n6112 0.0380882
R37424 DVDD.n6270 DVDD.n6112 0.0380882
R37425 DVDD.n6270 DVDD.n6268 0.0380882
R37426 DVDD.n6268 DVDD.n6266 0.0380882
R37427 DVDD.n6266 DVDD.n6115 0.0380882
R37428 DVDD.n6261 DVDD.n6115 0.0380882
R37429 DVDD.n6261 DVDD.n6259 0.0380882
R37430 DVDD.n6259 DVDD.n6257 0.0380882
R37431 DVDD.n6257 DVDD.n6118 0.0380882
R37432 DVDD.n6252 DVDD.n6118 0.0380882
R37433 DVDD.n6252 DVDD.n6250 0.0380882
R37434 DVDD.n6250 DVDD.n6248 0.0380882
R37435 DVDD.n6248 DVDD.n6121 0.0380882
R37436 DVDD.n6243 DVDD.n6121 0.0380882
R37437 DVDD.n6243 DVDD.n6241 0.0380882
R37438 DVDD.n6241 DVDD.n6239 0.0380882
R37439 DVDD.n6239 DVDD.n6124 0.0380882
R37440 DVDD.n6234 DVDD.n6124 0.0380882
R37441 DVDD.n6234 DVDD.n6232 0.0380882
R37442 DVDD.n6232 DVDD.n6230 0.0380882
R37443 DVDD.n6230 DVDD.n6127 0.0380882
R37444 DVDD.n6225 DVDD.n6127 0.0380882
R37445 DVDD.n6225 DVDD.n6223 0.0380882
R37446 DVDD.n6223 DVDD.n6221 0.0380882
R37447 DVDD.n6221 DVDD.n6130 0.0380882
R37448 DVDD.n6216 DVDD.n6130 0.0380882
R37449 DVDD.n6216 DVDD.n6214 0.0380882
R37450 DVDD.n6214 DVDD.n6212 0.0380882
R37451 DVDD.n6212 DVDD.n6133 0.0380882
R37452 DVDD.n6207 DVDD.n6133 0.0380882
R37453 DVDD.n6207 DVDD.n6205 0.0380882
R37454 DVDD.n6205 DVDD.n6203 0.0380882
R37455 DVDD.n6203 DVDD.n6136 0.0380882
R37456 DVDD.n6198 DVDD.n6136 0.0380882
R37457 DVDD.n6198 DVDD.n6196 0.0380882
R37458 DVDD.n6196 DVDD.n6194 0.0380882
R37459 DVDD.n6194 DVDD.n6139 0.0380882
R37460 DVDD.n6189 DVDD.n6139 0.0380882
R37461 DVDD.n6189 DVDD.n6187 0.0380882
R37462 DVDD.n6187 DVDD.n6185 0.0380882
R37463 DVDD.n6185 DVDD.n6142 0.0380882
R37464 DVDD.n6180 DVDD.n6142 0.0380882
R37465 DVDD.n6180 DVDD.n6178 0.0380882
R37466 DVDD.n6178 DVDD.n6176 0.0380882
R37467 DVDD.n6176 DVDD.n6145 0.0380882
R37468 DVDD.n6171 DVDD.n6145 0.0380882
R37469 DVDD.n6171 DVDD.n6169 0.0380882
R37470 DVDD.n6169 DVDD.n6167 0.0380882
R37471 DVDD.n6167 DVDD.n6148 0.0380882
R37472 DVDD.n6162 DVDD.n6148 0.0380882
R37473 DVDD.n6162 DVDD.n6160 0.0380882
R37474 DVDD.n6160 DVDD.n6158 0.0380882
R37475 DVDD.n6158 DVDD.n6151 0.0380882
R37476 DVDD.n6153 DVDD.n6151 0.0380882
R37477 DVDD.n6153 DVDD.n6049 0.0380882
R37478 DVDD.n6334 DVDD.n6049 0.0380882
R37479 DVDD.n6334 DVDD.n6047 0.0380882
R37480 DVDD.n15110 DVDD.n6047 0.0380882
R37481 DVDD.n1602 DVDD.n1601 0.0380882
R37482 DVDD.n1601 DVDD.n1315 0.0380882
R37483 DVDD.n1597 DVDD.n1315 0.0380882
R37484 DVDD.n1597 DVDD.n1593 0.0380882
R37485 DVDD.n1593 DVDD.n1592 0.0380882
R37486 DVDD.n1592 DVDD.n1317 0.0380882
R37487 DVDD.n1585 DVDD.n1317 0.0380882
R37488 DVDD.n1585 DVDD.n1581 0.0380882
R37489 DVDD.n1581 DVDD.n1580 0.0380882
R37490 DVDD.n1580 DVDD.n1319 0.0380882
R37491 DVDD.n1573 DVDD.n1319 0.0380882
R37492 DVDD.n1573 DVDD.n1569 0.0380882
R37493 DVDD.n1569 DVDD.n1568 0.0380882
R37494 DVDD.n1568 DVDD.n1321 0.0380882
R37495 DVDD.n1561 DVDD.n1321 0.0380882
R37496 DVDD.n1561 DVDD.n1557 0.0380882
R37497 DVDD.n1557 DVDD.n1556 0.0380882
R37498 DVDD.n1556 DVDD.n1323 0.0380882
R37499 DVDD.n1549 DVDD.n1323 0.0380882
R37500 DVDD.n1549 DVDD.n1545 0.0380882
R37501 DVDD.n1545 DVDD.n1544 0.0380882
R37502 DVDD.n1544 DVDD.n1325 0.0380882
R37503 DVDD.n1537 DVDD.n1325 0.0380882
R37504 DVDD.n1537 DVDD.n1533 0.0380882
R37505 DVDD.n1533 DVDD.n1532 0.0380882
R37506 DVDD.n1532 DVDD.n1327 0.0380882
R37507 DVDD.n1525 DVDD.n1327 0.0380882
R37508 DVDD.n1525 DVDD.n1521 0.0380882
R37509 DVDD.n1521 DVDD.n1520 0.0380882
R37510 DVDD.n1520 DVDD.n1329 0.0380882
R37511 DVDD.n1513 DVDD.n1329 0.0380882
R37512 DVDD.n1513 DVDD.n1509 0.0380882
R37513 DVDD.n1509 DVDD.n1508 0.0380882
R37514 DVDD.n1508 DVDD.n1331 0.0380882
R37515 DVDD.n1501 DVDD.n1331 0.0380882
R37516 DVDD.n1501 DVDD.n1497 0.0380882
R37517 DVDD.n1497 DVDD.n1496 0.0380882
R37518 DVDD.n1496 DVDD.n1333 0.0380882
R37519 DVDD.n1489 DVDD.n1333 0.0380882
R37520 DVDD.n1489 DVDD.n1485 0.0380882
R37521 DVDD.n1485 DVDD.n1484 0.0380882
R37522 DVDD.n1484 DVDD.n1335 0.0380882
R37523 DVDD.n1477 DVDD.n1335 0.0380882
R37524 DVDD.n1477 DVDD.n1473 0.0380882
R37525 DVDD.n1473 DVDD.n1472 0.0380882
R37526 DVDD.n1472 DVDD.n1337 0.0380882
R37527 DVDD.n1465 DVDD.n1337 0.0380882
R37528 DVDD.n1465 DVDD.n1461 0.0380882
R37529 DVDD.n1461 DVDD.n1460 0.0380882
R37530 DVDD.n1460 DVDD.n1339 0.0380882
R37531 DVDD.n1453 DVDD.n1339 0.0380882
R37532 DVDD.n1453 DVDD.n1449 0.0380882
R37533 DVDD.n1449 DVDD.n1448 0.0380882
R37534 DVDD.n1448 DVDD.n1341 0.0380882
R37535 DVDD.n1441 DVDD.n1341 0.0380882
R37536 DVDD.n1441 DVDD.n1437 0.0380882
R37537 DVDD.n1437 DVDD.n1436 0.0380882
R37538 DVDD.n1436 DVDD.n1343 0.0380882
R37539 DVDD.n1429 DVDD.n1343 0.0380882
R37540 DVDD.n1429 DVDD.n1425 0.0380882
R37541 DVDD.n1425 DVDD.n1424 0.0380882
R37542 DVDD.n1424 DVDD.n1345 0.0380882
R37543 DVDD.n1417 DVDD.n1345 0.0380882
R37544 DVDD.n1417 DVDD.n1413 0.0380882
R37545 DVDD.n1413 DVDD.n1412 0.0380882
R37546 DVDD.n1412 DVDD.n1347 0.0380882
R37547 DVDD.n1405 DVDD.n1347 0.0380882
R37548 DVDD.n1405 DVDD.n1401 0.0380882
R37549 DVDD.n1401 DVDD.n1400 0.0380882
R37550 DVDD.n1400 DVDD.n1349 0.0380882
R37551 DVDD.n1393 DVDD.n1349 0.0380882
R37552 DVDD.n1393 DVDD.n1389 0.0380882
R37553 DVDD.n1389 DVDD.n1388 0.0380882
R37554 DVDD.n1388 DVDD.n1351 0.0380882
R37555 DVDD.n1381 DVDD.n1351 0.0380882
R37556 DVDD.n1381 DVDD.n1377 0.0380882
R37557 DVDD.n1377 DVDD.n1376 0.0380882
R37558 DVDD.n1376 DVDD.n1353 0.0380882
R37559 DVDD.n1369 DVDD.n1353 0.0380882
R37560 DVDD.n1369 DVDD.n1365 0.0380882
R37561 DVDD.n1365 DVDD.n1364 0.0380882
R37562 DVDD.n1364 DVDD.n1355 0.0380882
R37563 DVDD.n1357 DVDD.n1355 0.0380882
R37564 DVDD.n1253 DVDD.n965 0.0380882
R37565 DVDD.n1253 DVDD.n967 0.0380882
R37566 DVDD.n1249 DVDD.n967 0.0380882
R37567 DVDD.n1249 DVDD.n1245 0.0380882
R37568 DVDD.n1245 DVDD.n1244 0.0380882
R37569 DVDD.n1244 DVDD.n969 0.0380882
R37570 DVDD.n1240 DVDD.n969 0.0380882
R37571 DVDD.n1240 DVDD.n1236 0.0380882
R37572 DVDD.n1236 DVDD.n1235 0.0380882
R37573 DVDD.n1235 DVDD.n974 0.0380882
R37574 DVDD.n1231 DVDD.n974 0.0380882
R37575 DVDD.n1231 DVDD.n1227 0.0380882
R37576 DVDD.n1227 DVDD.n1226 0.0380882
R37577 DVDD.n1226 DVDD.n979 0.0380882
R37578 DVDD.n1222 DVDD.n979 0.0380882
R37579 DVDD.n1222 DVDD.n1218 0.0380882
R37580 DVDD.n1218 DVDD.n1217 0.0380882
R37581 DVDD.n1217 DVDD.n984 0.0380882
R37582 DVDD.n1213 DVDD.n984 0.0380882
R37583 DVDD.n1213 DVDD.n1209 0.0380882
R37584 DVDD.n1209 DVDD.n1208 0.0380882
R37585 DVDD.n1208 DVDD.n989 0.0380882
R37586 DVDD.n1204 DVDD.n989 0.0380882
R37587 DVDD.n1204 DVDD.n1200 0.0380882
R37588 DVDD.n1200 DVDD.n1199 0.0380882
R37589 DVDD.n1199 DVDD.n994 0.0380882
R37590 DVDD.n1195 DVDD.n994 0.0380882
R37591 DVDD.n1195 DVDD.n1191 0.0380882
R37592 DVDD.n1191 DVDD.n1190 0.0380882
R37593 DVDD.n1190 DVDD.n999 0.0380882
R37594 DVDD.n1186 DVDD.n999 0.0380882
R37595 DVDD.n1186 DVDD.n1182 0.0380882
R37596 DVDD.n1182 DVDD.n1181 0.0380882
R37597 DVDD.n1181 DVDD.n1004 0.0380882
R37598 DVDD.n1177 DVDD.n1004 0.0380882
R37599 DVDD.n1177 DVDD.n1173 0.0380882
R37600 DVDD.n1173 DVDD.n1172 0.0380882
R37601 DVDD.n1172 DVDD.n1009 0.0380882
R37602 DVDD.n1168 DVDD.n1009 0.0380882
R37603 DVDD.n1168 DVDD.n1164 0.0380882
R37604 DVDD.n1164 DVDD.n1163 0.0380882
R37605 DVDD.n1163 DVDD.n1014 0.0380882
R37606 DVDD.n1159 DVDD.n1014 0.0380882
R37607 DVDD.n1159 DVDD.n1155 0.0380882
R37608 DVDD.n1155 DVDD.n1154 0.0380882
R37609 DVDD.n1154 DVDD.n1019 0.0380882
R37610 DVDD.n1150 DVDD.n1019 0.0380882
R37611 DVDD.n1150 DVDD.n1146 0.0380882
R37612 DVDD.n1146 DVDD.n1145 0.0380882
R37613 DVDD.n1145 DVDD.n1024 0.0380882
R37614 DVDD.n1141 DVDD.n1024 0.0380882
R37615 DVDD.n1141 DVDD.n1137 0.0380882
R37616 DVDD.n1137 DVDD.n1136 0.0380882
R37617 DVDD.n1136 DVDD.n1029 0.0380882
R37618 DVDD.n1132 DVDD.n1029 0.0380882
R37619 DVDD.n1132 DVDD.n1128 0.0380882
R37620 DVDD.n1128 DVDD.n1127 0.0380882
R37621 DVDD.n1127 DVDD.n1034 0.0380882
R37622 DVDD.n1123 DVDD.n1034 0.0380882
R37623 DVDD.n1123 DVDD.n1119 0.0380882
R37624 DVDD.n1119 DVDD.n1118 0.0380882
R37625 DVDD.n1118 DVDD.n1039 0.0380882
R37626 DVDD.n1114 DVDD.n1039 0.0380882
R37627 DVDD.n1114 DVDD.n1110 0.0380882
R37628 DVDD.n1110 DVDD.n1109 0.0380882
R37629 DVDD.n1109 DVDD.n1044 0.0380882
R37630 DVDD.n1105 DVDD.n1044 0.0380882
R37631 DVDD.n1105 DVDD.n1101 0.0380882
R37632 DVDD.n1101 DVDD.n1100 0.0380882
R37633 DVDD.n1100 DVDD.n1049 0.0380882
R37634 DVDD.n1096 DVDD.n1049 0.0380882
R37635 DVDD.n1096 DVDD.n1092 0.0380882
R37636 DVDD.n1092 DVDD.n1091 0.0380882
R37637 DVDD.n1091 DVDD.n1054 0.0380882
R37638 DVDD.n1087 DVDD.n1054 0.0380882
R37639 DVDD.n1087 DVDD.n1083 0.0380882
R37640 DVDD.n1083 DVDD.n1082 0.0380882
R37641 DVDD.n1082 DVDD.n1059 0.0380882
R37642 DVDD.n1078 DVDD.n1059 0.0380882
R37643 DVDD.n1078 DVDD.n1074 0.0380882
R37644 DVDD.n1074 DVDD.n1073 0.0380882
R37645 DVDD.n1073 DVDD.n1064 0.0380882
R37646 DVDD.n1069 DVDD.n1064 0.0380882
R37647 DVDD.n1252 DVDD.n918 0.0380882
R37648 DVDD.n1252 DVDD.n1251 0.0380882
R37649 DVDD.n1251 DVDD.n1250 0.0380882
R37650 DVDD.n1250 DVDD.n968 0.0380882
R37651 DVDD.n1243 DVDD.n968 0.0380882
R37652 DVDD.n1243 DVDD.n1242 0.0380882
R37653 DVDD.n1242 DVDD.n1241 0.0380882
R37654 DVDD.n1241 DVDD.n973 0.0380882
R37655 DVDD.n1234 DVDD.n973 0.0380882
R37656 DVDD.n1234 DVDD.n1233 0.0380882
R37657 DVDD.n1233 DVDD.n1232 0.0380882
R37658 DVDD.n1232 DVDD.n978 0.0380882
R37659 DVDD.n1225 DVDD.n978 0.0380882
R37660 DVDD.n1225 DVDD.n1224 0.0380882
R37661 DVDD.n1224 DVDD.n1223 0.0380882
R37662 DVDD.n1223 DVDD.n983 0.0380882
R37663 DVDD.n1216 DVDD.n983 0.0380882
R37664 DVDD.n1216 DVDD.n1215 0.0380882
R37665 DVDD.n1215 DVDD.n1214 0.0380882
R37666 DVDD.n1214 DVDD.n988 0.0380882
R37667 DVDD.n1207 DVDD.n988 0.0380882
R37668 DVDD.n1207 DVDD.n1206 0.0380882
R37669 DVDD.n1206 DVDD.n1205 0.0380882
R37670 DVDD.n1205 DVDD.n993 0.0380882
R37671 DVDD.n1198 DVDD.n993 0.0380882
R37672 DVDD.n1198 DVDD.n1197 0.0380882
R37673 DVDD.n1197 DVDD.n1196 0.0380882
R37674 DVDD.n1196 DVDD.n998 0.0380882
R37675 DVDD.n1189 DVDD.n998 0.0380882
R37676 DVDD.n1189 DVDD.n1188 0.0380882
R37677 DVDD.n1188 DVDD.n1187 0.0380882
R37678 DVDD.n1187 DVDD.n1003 0.0380882
R37679 DVDD.n1180 DVDD.n1003 0.0380882
R37680 DVDD.n1180 DVDD.n1179 0.0380882
R37681 DVDD.n1179 DVDD.n1178 0.0380882
R37682 DVDD.n1178 DVDD.n1008 0.0380882
R37683 DVDD.n1171 DVDD.n1008 0.0380882
R37684 DVDD.n1171 DVDD.n1170 0.0380882
R37685 DVDD.n1170 DVDD.n1169 0.0380882
R37686 DVDD.n1169 DVDD.n1013 0.0380882
R37687 DVDD.n1162 DVDD.n1013 0.0380882
R37688 DVDD.n1162 DVDD.n1161 0.0380882
R37689 DVDD.n1161 DVDD.n1160 0.0380882
R37690 DVDD.n1160 DVDD.n1018 0.0380882
R37691 DVDD.n1153 DVDD.n1018 0.0380882
R37692 DVDD.n1153 DVDD.n1152 0.0380882
R37693 DVDD.n1152 DVDD.n1151 0.0380882
R37694 DVDD.n1151 DVDD.n1023 0.0380882
R37695 DVDD.n1144 DVDD.n1023 0.0380882
R37696 DVDD.n1144 DVDD.n1143 0.0380882
R37697 DVDD.n1143 DVDD.n1142 0.0380882
R37698 DVDD.n1142 DVDD.n1028 0.0380882
R37699 DVDD.n1135 DVDD.n1028 0.0380882
R37700 DVDD.n1135 DVDD.n1134 0.0380882
R37701 DVDD.n1134 DVDD.n1133 0.0380882
R37702 DVDD.n1133 DVDD.n1033 0.0380882
R37703 DVDD.n1126 DVDD.n1033 0.0380882
R37704 DVDD.n1126 DVDD.n1125 0.0380882
R37705 DVDD.n1125 DVDD.n1124 0.0380882
R37706 DVDD.n1124 DVDD.n1038 0.0380882
R37707 DVDD.n1117 DVDD.n1038 0.0380882
R37708 DVDD.n1117 DVDD.n1116 0.0380882
R37709 DVDD.n1116 DVDD.n1115 0.0380882
R37710 DVDD.n1115 DVDD.n1043 0.0380882
R37711 DVDD.n1108 DVDD.n1043 0.0380882
R37712 DVDD.n1108 DVDD.n1107 0.0380882
R37713 DVDD.n1107 DVDD.n1106 0.0380882
R37714 DVDD.n1106 DVDD.n1048 0.0380882
R37715 DVDD.n1099 DVDD.n1048 0.0380882
R37716 DVDD.n1099 DVDD.n1098 0.0380882
R37717 DVDD.n1098 DVDD.n1097 0.0380882
R37718 DVDD.n1097 DVDD.n1053 0.0380882
R37719 DVDD.n1090 DVDD.n1053 0.0380882
R37720 DVDD.n1090 DVDD.n1089 0.0380882
R37721 DVDD.n1089 DVDD.n1088 0.0380882
R37722 DVDD.n1088 DVDD.n1058 0.0380882
R37723 DVDD.n1081 DVDD.n1058 0.0380882
R37724 DVDD.n1081 DVDD.n1080 0.0380882
R37725 DVDD.n1080 DVDD.n1079 0.0380882
R37726 DVDD.n1079 DVDD.n1063 0.0380882
R37727 DVDD.n1072 DVDD.n1063 0.0380882
R37728 DVDD.n1072 DVDD.n1071 0.0380882
R37729 DVDD.n1071 DVDD.n1070 0.0380882
R37730 DVDD DVDD.t162 0.0375588
R37731 DVDD DVDD.t156 0.0375588
R37732 DVDD DVDD.t159 0.0375588
R37733 DVDD DVDD.t160 0.0375588
R37734 DVDD.n19095 DVDD.n18770 0.036061
R37735 DVDD.n19102 DVDD.n19101 0.036061
R37736 DVDD.n21055 DVDD.n18763 0.036061
R37737 DVDD.n20978 DVDD.n20974 0.036061
R37738 DVDD.n19789 DVDD.n18821 0.0336579
R37739 DVDD.n21016 DVDD.n18753 0.0336579
R37740 DVDD.n9574 DVDD.t123 0.03326
R37741 DVDD.n9574 DVDD.t144 0.03326
R37742 DVDD.n3447 DVDD.t107 0.03326
R37743 DVDD.n3447 DVDD.t133 0.03326
R37744 DVDD.n3436 DVDD.t117 0.03326
R37745 DVDD.n3436 DVDD.t76 0.03326
R37746 DVDD.n15607 DVDD.t102 0.03326
R37747 DVDD.n15607 DVDD.t90 0.03326
R37748 DVDD.n15576 DVDD.t112 0.03326
R37749 DVDD.n15576 DVDD.t97 0.03326
R37750 DVDD.n15567 DVDD.t118 0.03326
R37751 DVDD.n15567 DVDD.t83 0.03326
R37752 DVDD.n15558 DVDD.t129 0.03326
R37753 DVDD.n15558 DVDD.t91 0.03326
R37754 DVDD.n15549 DVDD.t73 0.03326
R37755 DVDD.n15549 DVDD.t104 0.03326
R37756 DVDD.n15540 DVDD.t140 0.03326
R37757 DVDD.n15540 DVDD.t108 0.03326
R37758 DVDD.n15531 DVDD.t145 0.03326
R37759 DVDD.n15531 DVDD.t119 0.03326
R37760 DVDD.n5186 DVDD.t82 0.03326
R37761 DVDD.n5186 DVDD.t125 0.03326
R37762 DVDD.n5175 DVDD.t93 0.03326
R37763 DVDD.n5175 DVDD.t134 0.03326
R37764 DVDD.n5164 DVDD.t101 0.03326
R37765 DVDD.n5164 DVDD.t109 0.03326
R37766 DVDD.n3106 DVDD.t147 0.03326
R37767 DVDD.n3106 DVDD.t114 0.03326
R37768 DVDD.n16036 DVDD.t74 0.03326
R37769 DVDD.n16036 DVDD.t124 0.03326
R37770 DVDD.n16025 DVDD.t85 0.03326
R37771 DVDD.n16025 DVDD.t110 0.03326
R37772 DVDD.n16047 DVDD.t95 0.03326
R37773 DVDD.n16047 DVDD.t120 0.03326
R37774 DVDD.n16013 DVDD.t105 0.03326
R37775 DVDD.n16013 DVDD.t142 0.03326
R37776 DVDD.n16063 DVDD.t88 0.03326
R37777 DVDD.n16063 DVDD.t150 0.03326
R37778 DVDD.n9776 DVDD.t103 0.03326
R37779 DVDD.n9776 DVDD.t84 0.03326
R37780 DVDD.n9943 DVDD.t130 0.03326
R37781 DVDD.n9943 DVDD.t152 0.03326
R37782 DVDD.n9801 DVDD.t136 0.03326
R37783 DVDD.n9801 DVDD.t78 0.03326
R37784 DVDD.n9952 DVDD.t146 0.03326
R37785 DVDD.n9952 DVDD.t92 0.03326
R37786 DVDD.n9611 DVDD.t131 0.03326
R37787 DVDD.n9611 DVDD.t98 0.03326
R37788 DVDD.n10100 DVDD.t141 0.03326
R37789 DVDD.n10100 DVDD.t126 0.03326
R37790 DVDD.n10105 DVDD.t148 0.03326
R37791 DVDD.n10105 DVDD.t111 0.03326
R37792 DVDD.n9603 DVDD.t80 0.03326
R37793 DVDD.n9603 DVDD.t121 0.03326
R37794 DVDD.n10113 DVDD.t86 0.03326
R37795 DVDD.n10113 DVDD.t127 0.03326
R37796 DVDD.n10125 DVDD.t137 0.03326
R37797 DVDD.n10125 DVDD.t106 0.03326
R37798 DVDD.n10130 DVDD.t149 0.03326
R37799 DVDD.n10130 DVDD.t115 0.03326
R37800 DVDD.n9588 DVDD.t75 0.03326
R37801 DVDD.n9588 DVDD.t116 0.03326
R37802 DVDD.n10138 DVDD.t87 0.03326
R37803 DVDD.n10138 DVDD.t128 0.03326
R37804 DVDD.n10143 DVDD.t96 0.03326
R37805 DVDD.n10143 DVDD.t135 0.03326
R37806 DVDD.n9580 DVDD.t81 0.03326
R37807 DVDD.n9580 DVDD.t143 0.03326
R37808 DVDD.n10151 DVDD.t89 0.03326
R37809 DVDD.n10151 DVDD.t151 0.03326
R37810 DVDD.n10159 DVDD.t113 0.03326
R37811 DVDD.n10159 DVDD.t138 0.03326
R37812 DVDD.n18420 DVDD.n18419 0.03245
R37813 DVDD.n18419 DVDD.n18415 0.03245
R37814 DVDD.n18415 DVDD.n178 0.03245
R37815 DVDD.n21850 DVDD.n182 0.03245
R37816 DVDD.n21850 DVDD.n21846 0.03245
R37817 DVDD.n21854 DVDD.n21846 0.03245
R37818 DVDD.n21972 DVDD.n18275 0.03245
R37819 DVDD.n21972 DVDD.n18278 0.03245
R37820 DVDD.n18278 DVDD.n18277 0.03245
R37821 DVDD.n22016 DVDD.n22013 0.03245
R37822 DVDD.n22016 DVDD.n22012 0.03245
R37823 DVDD.n22020 DVDD.n22012 0.03245
R37824 DVDD.n21244 DVDD.n21243 0.03245
R37825 DVDD.n21243 DVDD.n21240 0.03245
R37826 DVDD.n21240 DVDD.n21239 0.03245
R37827 DVDD.n21351 DVDD.n21341 0.03245
R37828 DVDD.n21351 DVDD.n21343 0.03245
R37829 DVDD.n21347 DVDD.n21343 0.03245
R37830 DVDD.n21696 DVDD.n18522 0.03245
R37831 DVDD.n21701 DVDD.n18522 0.03245
R37832 DVDD.n21701 DVDD.n191 0.03245
R37833 DVDD.n21953 DVDD.n192 0.03245
R37834 DVDD.n21953 DVDD.n18289 0.03245
R37835 DVDD.n21957 DVDD.n18289 0.03245
R37836 DVDD.n21825 DVDD.n21818 0.03245
R37837 DVDD.n21825 DVDD.n21821 0.03245
R37838 DVDD.n21821 DVDD.n21820 0.03245
R37839 DVDD.n18262 DVDD.n18261 0.03245
R37840 DVDD.n18261 DVDD.n18254 0.03245
R37841 DVDD.n18257 DVDD.n18254 0.03245
R37842 DVDD.n18473 DVDD.n18466 0.03245
R37843 DVDD.n18473 DVDD.n18469 0.03245
R37844 DVDD.n18469 DVDD.n18468 0.03245
R37845 DVDD.n18446 DVDD.n18445 0.03245
R37846 DVDD.n18445 DVDD.n18444 0.03245
R37847 DVDD.n18444 DVDD.n18441 0.03245
R37848 DVDD.n4293 DVDD.n4286 0.03245
R37849 DVDD.n4293 DVDD.n4284 0.03245
R37850 DVDD.n4297 DVDD.n4284 0.03245
R37851 DVDD.n4313 DVDD.n4300 0.03245
R37852 DVDD.n4309 DVDD.n4300 0.03245
R37853 DVDD.n4309 DVDD.n4308 0.03245
R37854 DVDD.n3685 DVDD.n3679 0.03245
R37855 DVDD.n3690 DVDD.n3679 0.03245
R37856 DVDD.n3690 DVDD.n3674 0.03245
R37857 DVDD.n3705 DVDD.n3675 0.03245
R37858 DVDD.n3705 DVDD.n3696 0.03245
R37859 DVDD.n3701 DVDD.n3696 0.03245
R37860 DVDD.n15125 DVDD.n5931 0.03245
R37861 DVDD.n6342 DVDD.n5931 0.03245
R37862 DVDD.n15107 DVDD.n15106 0.03245
R37863 DVDD.n15106 DVDD.n15105 0.03245
R37864 DVDD.n7050 DVDD.n7049 0.03245
R37865 DVDD.n15084 DVDD.n15083 0.03245
R37866 DVDD.n15083 DVDD.n15082 0.03245
R37867 DVDD.n15066 DVDD.n15065 0.03245
R37868 DVDD.n15065 DVDD.n15064 0.03245
R37869 DVDD.n7671 DVDD.n7665 0.03245
R37870 DVDD.n7672 DVDD.n7671 0.03245
R37871 DVDD.n14855 DVDD.n14854 0.03245
R37872 DVDD.n14854 DVDD.n14853 0.03245
R37873 DVDD.n8035 DVDD.n8027 0.03245
R37874 DVDD.n8036 DVDD.n8035 0.03245
R37875 DVDD.n14832 DVDD.n14831 0.03245
R37876 DVDD.n14829 DVDD.n8039 0.03245
R37877 DVDD.n14565 DVDD.n8039 0.03245
R37878 DVDD.n14563 DVDD.n8159 0.03245
R37879 DVDD.n8604 DVDD.n8159 0.03245
R37880 DVDD.n14299 DVDD.n14298 0.03245
R37881 DVDD.n14298 DVDD.n14297 0.03245
R37882 DVDD.n10588 DVDD.n10580 0.03245
R37883 DVDD.n10589 DVDD.n10588 0.03245
R37884 DVDD.n14276 DVDD.n14275 0.03245
R37885 DVDD.n14273 DVDD.n10592 0.03245
R37886 DVDD.n11056 DVDD.n10592 0.03245
R37887 DVDD.n14009 DVDD.n14008 0.03245
R37888 DVDD.n14008 DVDD.n14007 0.03245
R37889 DVDD.n11570 DVDD.n11569 0.03245
R37890 DVDD.n11569 DVDD.n11565 0.03245
R37891 DVDD.n13791 DVDD.n11566 0.03245
R37892 DVDD.n11919 DVDD.n11566 0.03245
R37893 DVDD.n13769 DVDD.n11920 0.03245
R37894 DVDD.n12279 DVDD.n11920 0.03245
R37895 DVDD.n13751 DVDD.n13750 0.03245
R37896 DVDD.n13748 DVDD.n12282 0.03245
R37897 DVDD.n12730 DVDD.n12282 0.03245
R37898 DVDD.n13479 DVDD.n13478 0.03245
R37899 DVDD.n13478 DVDD.n13477 0.03245
R37900 DVDD.n12918 DVDD.n12916 0.03245
R37901 DVDD.n13261 DVDD.n12916 0.03245
R37902 DVDD.n13263 DVDD.n2160 0.03245
R37903 DVDD.n16708 DVDD.n2160 0.03245
R37904 DVDD.n16711 DVDD.n16710 0.03245
R37905 DVDD.n16731 DVDD.n16730 0.03245
R37906 DVDD.n16732 DVDD.n16731 0.03245
R37907 DVDD.n16999 DVDD.n16998 0.03245
R37908 DVDD.n17000 DVDD.n16999 0.03245
R37909 DVDD.n17267 DVDD.n17266 0.03245
R37910 DVDD.n17268 DVDD.n17267 0.03245
R37911 DVDD.n17285 DVDD.n17284 0.03245
R37912 DVDD.n17286 DVDD.n17285 0.03245
R37913 DVDD.n17304 DVDD.n17303 0.03245
R37914 DVDD.n17714 DVDD.n17304 0.03245
R37915 DVDD.n20465 DVDD.n20464 0.0318024
R37916 DVDD.n21052 DVDD.n21051 0.0318024
R37917 DVDD.n20923 DVDD.n20922 0.0318024
R37918 DVDD.n21048 DVDD.n18819 0.0318024
R37919 DVDD.n20538 DVDD.n20535 0.0318024
R37920 DVDD.n21081 DVDD.n21059 0.0318024
R37921 DVDD.n20531 DVDD.n20519 0.0318024
R37922 DVDD.n21012 DVDD.n20982 0.0318024
R37923 DVDD.n7051 DVDD.n7050 0.031775
R37924 DVDD.n17276 DVDD.n1267 0.0317353
R37925 DVDD.n6858 DVDD.n6703 0.0317353
R37926 DVDD.n15074 DVDD.n7066 0.0317353
R37927 DVDD.n14870 DVDD.n14869 0.0317353
R37928 DVDD.n9219 DVDD.n9218 0.0317353
R37929 DVDD.n9265 DVDD.n7684 0.0317353
R37930 DVDD.n7839 DVDD.n7685 0.0317353
R37931 DVDD.n14578 DVDD.n8133 0.0317353
R37932 DVDD.n14312 DVDD.n8250 0.0317353
R37933 DVDD.n8347 DVDD.n8254 0.0317353
R37934 DVDD.n10237 DVDD.n8949 0.0317353
R37935 DVDD.n10392 DVDD.n10238 0.0317353
R37936 DVDD.n14022 DVDD.n10686 0.0317353
R37937 DVDD.n10799 DVDD.n10706 0.0317353
R37938 DVDD.n13813 DVDD.n13812 0.0317353
R37939 DVDD.n13804 DVDD.n11229 0.0317353
R37940 DVDD.n13782 DVDD.n11584 0.0317353
R37941 DVDD.n13759 DVDD.n11930 0.0317353
R37942 DVDD.n13497 DVDD.n12377 0.0317353
R37943 DVDD.n12541 DVDD.n12384 0.0317353
R37944 DVDD.n13283 DVDD.n13282 0.0317353
R37945 DVDD.n13273 DVDD.n12903 0.0317353
R37946 DVDD.n16457 DVDD.n2254 0.0317353
R37947 DVDD.n16720 DVDD.n1817 0.0317353
R37948 DVDD.n16746 DVDD.n1801 0.0317353
R37949 DVDD.n17014 DVDD.n1702 0.0317353
R37950 DVDD.n6702 DVDD.n6396 0.0317353
R37951 DVDD.n6094 DVDD.n5997 0.0317353
R37952 DVDD.n17294 DVDD.n918 0.0317353
R37953 DVDD.n14275 DVDD.n14274 0.031325
R37954 DVDD.n21272 DVDD.n21271 0.0309579
R37955 DVDD.n22239 DVDD.n128 0.0309579
R37956 DVDD.n13751 DVDD.n12280 0.030875
R37957 DVDD.n16711 DVDD.n1808 0.030875
R37958 DVDD.n20537 DVDD.n20536 0.0308261
R37959 DVDD.n20539 DVDD.n19781 0.0308261
R37960 DVDD.n20442 DVDD.n19818 0.0308261
R37961 DVDD.n20463 DVDD.n19819 0.0308261
R37962 DVDD.n21082 DVDD.n18752 0.0308261
R37963 DVDD.n14832 DVDD.n8037 0.030425
R37964 DVDD.n20532 DVDD.n20486 0.0287281
R37965 DVDD.n20483 DVDD.n19809 0.0287281
R37966 DVDD.n20466 DVDD.n18907 0.0287281
R37967 DVDD.n20951 DVDD.n20950 0.0287281
R37968 DVDD.n20934 DVDD.n20933 0.0287281
R37969 DVDD.n19122 DVDD.n19093 0.0287281
R37970 DVDD.n19106 DVDD.n19105 0.0287281
R37971 DVDD.n18828 DVDD.n18762 0.0287281
R37972 DVDD.n21054 DVDD.n18761 0.0287281
R37973 DVDD.n19098 DVDD.n18786 0.0287281
R37974 DVDD.n18774 DVDD.n18773 0.0287281
R37975 DVDD.n19121 DVDD.n19120 0.0287281
R37976 DVDD.n20949 DVDD.n20948 0.0287281
R37977 DVDD.n20479 DVDD.n20478 0.0287281
R37978 DVDD.n21056 DVDD.n18755 0.0287281
R37979 DVDD.n19079 DVDD.n18830 0.0287281
R37980 DVDD.n20966 DVDD.n20965 0.0287281
R37981 DVDD.n20485 DVDD.n20484 0.0287281
R37982 DVDD.n20979 DVDD.n18825 0.0287281
R37983 DVDD.n20526 DVDD.n20524 0.0287281
R37984 DVDD.n14831 DVDD.n14830 0.028625
R37985 DVDD.n15123 DVDD.n5933 0.0284039
R37986 DVDD.n6338 DVDD.n5933 0.0284039
R37987 DVDD.n6346 DVDD.n6341 0.0284039
R37988 DVDD.n15103 DVDD.n6346 0.0284039
R37989 DVDD.n7047 DVDD.n7046 0.0284039
R37990 DVDD.n7054 DVDD.n7045 0.0284039
R37991 DVDD.n15080 DVDD.n7054 0.0284039
R37992 DVDD.n15068 DVDD.n7405 0.0284039
R37993 DVDD.n15062 DVDD.n7405 0.0284039
R37994 DVDD.n7669 DVDD.n7667 0.0284039
R37995 DVDD.n7669 DVDD.n7668 0.0284039
R37996 DVDD.n7676 DVDD.n7664 0.0284039
R37997 DVDD.n14851 DVDD.n7676 0.0284039
R37998 DVDD.n8033 DVDD.n8031 0.0284039
R37999 DVDD.n8033 DVDD.n8032 0.0284039
R38000 DVDD.n8144 DVDD.n8026 0.0284039
R38001 DVDD.n14827 DVDD.n8043 0.0284039
R38002 DVDD.n14567 DVDD.n8043 0.0284039
R38003 DVDD.n14561 DVDD.n8161 0.0284039
R38004 DVDD.n8602 DVDD.n8161 0.0284039
R38005 DVDD.n14301 DVDD.n8261 0.0284039
R38006 DVDD.n14295 DVDD.n8261 0.0284039
R38007 DVDD.n10586 DVDD.n10584 0.0284039
R38008 DVDD.n10586 DVDD.n10585 0.0284039
R38009 DVDD.n10691 DVDD.n10579 0.0284039
R38010 DVDD.n14271 DVDD.n10596 0.0284039
R38011 DVDD.n11054 DVDD.n10596 0.0284039
R38012 DVDD.n14011 DVDD.n10713 0.0284039
R38013 DVDD.n14005 DVDD.n10713 0.0284039
R38014 DVDD.n11574 DVDD.n11572 0.0284039
R38015 DVDD.n11575 DVDD.n11574 0.0284039
R38016 DVDD.n13789 DVDD.n13788 0.0284039
R38017 DVDD.n13788 DVDD.n11579 0.0284039
R38018 DVDD.n13767 DVDD.n13766 0.0284039
R38019 DVDD.n13766 DVDD.n11924 0.0284039
R38020 DVDD.n13753 DVDD.n11941 0.0284039
R38021 DVDD.n13746 DVDD.n12286 0.0284039
R38022 DVDD.n12726 DVDD.n12286 0.0284039
R38023 DVDD.n12734 DVDD.n12729 0.0284039
R38024 DVDD.n13475 DVDD.n12734 0.0284039
R38025 DVDD.n12922 DVDD.n12920 0.0284039
R38026 DVDD.n13259 DVDD.n12922 0.0284039
R38027 DVDD.n13265 DVDD.n2163 0.0284039
R38028 DVDD.n16706 DVDD.n2163 0.0284039
R38029 DVDD.n16713 DVDD.n2157 0.0284039
R38030 DVDD.n16728 DVDD.n1806 0.0284039
R38031 DVDD.n16734 DVDD.n1806 0.0284039
R38032 DVDD.n16996 DVDD.n1707 0.0284039
R38033 DVDD.n17002 DVDD.n1707 0.0284039
R38034 DVDD.n17264 DVDD.n1606 0.0284039
R38035 DVDD.n17270 DVDD.n1606 0.0284039
R38036 DVDD.n17282 DVDD.n1257 0.0284039
R38037 DVDD.n17288 DVDD.n1257 0.0284039
R38038 DVDD.n17301 DVDD.n908 0.0284039
R38039 DVDD.n17716 DVDD.n908 0.0284039
R38040 DVDD.n15124 DVDD.n5932 0.0284039
R38041 DVDD.n6339 DVDD.n5932 0.0284039
R38042 DVDD.n15108 DVDD.n6340 0.0284039
R38043 DVDD.n15104 DVDD.n6340 0.0284039
R38044 DVDD.n7048 DVDD.n7043 0.0284039
R38045 DVDD.n15085 DVDD.n7044 0.0284039
R38046 DVDD.n15081 DVDD.n7044 0.0284039
R38047 DVDD.n15067 DVDD.n7406 0.0284039
R38048 DVDD.n15063 DVDD.n7406 0.0284039
R38049 DVDD.n7670 DVDD.n7666 0.0284039
R38050 DVDD.n7670 DVDD.n7662 0.0284039
R38051 DVDD.n14856 DVDD.n7663 0.0284039
R38052 DVDD.n14852 DVDD.n7663 0.0284039
R38053 DVDD.n8034 DVDD.n8028 0.0284039
R38054 DVDD.n8034 DVDD.n8024 0.0284039
R38055 DVDD.n14833 DVDD.n8025 0.0284039
R38056 DVDD.n14828 DVDD.n8041 0.0284039
R38057 DVDD.n14566 DVDD.n8041 0.0284039
R38058 DVDD.n14562 DVDD.n8160 0.0284039
R38059 DVDD.n8603 DVDD.n8160 0.0284039
R38060 DVDD.n14300 DVDD.n8263 0.0284039
R38061 DVDD.n14296 DVDD.n8263 0.0284039
R38062 DVDD.n10587 DVDD.n10581 0.0284039
R38063 DVDD.n10587 DVDD.n10577 0.0284039
R38064 DVDD.n14277 DVDD.n10578 0.0284039
R38065 DVDD.n14272 DVDD.n10594 0.0284039
R38066 DVDD.n11055 DVDD.n10594 0.0284039
R38067 DVDD.n14010 DVDD.n10715 0.0284039
R38068 DVDD.n14006 DVDD.n10715 0.0284039
R38069 DVDD.n11571 DVDD.n11567 0.0284039
R38070 DVDD.n11576 DVDD.n11567 0.0284039
R38071 DVDD.n13790 DVDD.n11578 0.0284039
R38072 DVDD.n11921 DVDD.n11578 0.0284039
R38073 DVDD.n13768 DVDD.n11923 0.0284039
R38074 DVDD.n12278 DVDD.n11923 0.0284039
R38075 DVDD.n13752 DVDD.n11943 0.0284039
R38076 DVDD.n13747 DVDD.n12284 0.0284039
R38077 DVDD.n12727 DVDD.n12284 0.0284039
R38078 DVDD.n13480 DVDD.n12728 0.0284039
R38079 DVDD.n13476 DVDD.n12728 0.0284039
R38080 DVDD.n12919 DVDD.n12917 0.0284039
R38081 DVDD.n13260 DVDD.n12917 0.0284039
R38082 DVDD.n13264 DVDD.n2161 0.0284039
R38083 DVDD.n16707 DVDD.n2161 0.0284039
R38084 DVDD.n16712 DVDD.n2158 0.0284039
R38085 DVDD.n16729 DVDD.n1807 0.0284039
R38086 DVDD.n16733 DVDD.n1807 0.0284039
R38087 DVDD.n16997 DVDD.n1708 0.0284039
R38088 DVDD.n17001 DVDD.n1708 0.0284039
R38089 DVDD.n17265 DVDD.n1607 0.0284039
R38090 DVDD.n17269 DVDD.n1607 0.0284039
R38091 DVDD.n17283 DVDD.n1258 0.0284039
R38092 DVDD.n17287 DVDD.n1258 0.0284039
R38093 DVDD.n17302 DVDD.n910 0.0284039
R38094 DVDD.n17715 DVDD.n910 0.0284039
R38095 DVDD.n18423 DVDD.n18422 0.0284
R38096 DVDD.n21856 DVDD.n21842 0.0284
R38097 DVDD.n21974 DVDD.n18273 0.0284
R38098 DVDD.n22011 DVDD.n232 0.0284
R38099 DVDD.n21235 DVDD.n21219 0.0284
R38100 DVDD.n21345 DVDD.n21344 0.0284
R38101 DVDD.n18524 DVDD.n18523 0.0284
R38102 DVDD.n21959 DVDD.n18287 0.0284
R38103 DVDD.n21827 DVDD.n21813 0.0284
R38104 DVDD.n18255 DVDD.n18218 0.0284
R38105 DVDD.n18475 DVDD.n18463 0.0284
R38106 DVDD.n18439 DVDD.n18411 0.0284
R38107 DVDD.n4287 DVDD.n4242 0.0284
R38108 DVDD.n4305 DVDD.n4269 0.0284
R38109 DVDD.n3681 DVDD.n3680 0.0284
R38110 DVDD.n3699 DVDD.n3655 0.0284
R38111 DVDD.n13750 DVDD.n13749 0.028175
R38112 DVDD.n16710 DVDD.n16709 0.028175
R38113 DVDD.n15143 DVDD.n15142 0.0278316
R38114 DVDD.n17731 DVDD.n17727 0.0278316
R38115 DVDD.n7046 DVDD.n6795 0.0278144
R38116 DVDD.n15086 DVDD.n7043 0.0278144
R38117 DVDD.n18421 DVDD.n18397 0.027725
R38118 DVDD.n22022 DVDD.n22021 0.027725
R38119 DVDD.n21346 DVDD.n18553 0.027725
R38120 DVDD.n21695 DVDD.n21694 0.027725
R38121 DVDD.n18256 DVDD.n18216 0.027725
R38122 DVDD.n18440 DVDD.n18438 0.027725
R38123 DVDD.n4289 DVDD.n4288 0.027725
R38124 DVDD.n3684 DVDD.n3683 0.027725
R38125 DVDD.n14276 DVDD.n10590 0.027725
R38126 DVDD.n10691 DVDD.n10595 0.0274214
R38127 DVDD.n10593 DVDD.n10578 0.0274214
R38128 DVDD.n21855 DVDD.n21844 0.027275
R38129 DVDD.n21968 DVDD.n18279 0.027275
R38130 DVDD.n21246 DVDD.n21245 0.027275
R38131 DVDD.n21958 DVDD.n18288 0.027275
R38132 DVDD.n21817 DVDD.n21812 0.027275
R38133 DVDD.n18465 DVDD.n124 0.027275
R38134 DVDD.n4307 DVDD.n4306 0.027275
R38135 DVDD.n3700 DVDD.n3698 0.027275
R38136 DVDD.n7049 DVDD.n6344 0.027275
R38137 DVDD.n13753 DVDD.n11940 0.0270284
R38138 DVDD.n16713 DVDD.n1810 0.0270284
R38139 DVDD.n13752 DVDD.n11942 0.0270284
R38140 DVDD.n16712 DVDD.n1809 0.0270284
R38141 DVDD.n18022 DVDD.n18021 0.026913
R38142 DVDD.n18021 DVDD.n18019 0.026913
R38143 DVDD.n18019 DVDD.n18017 0.026913
R38144 DVDD.n18017 DVDD.n18015 0.026913
R38145 DVDD.n18015 DVDD.n18013 0.026913
R38146 DVDD.n18013 DVDD.n18011 0.026913
R38147 DVDD.n18011 DVDD.n18008 0.026913
R38148 DVDD.n18008 DVDD.n18007 0.026913
R38149 DVDD.n18007 DVDD.n18005 0.026913
R38150 DVDD.n18005 DVDD.n18003 0.026913
R38151 DVDD.n18003 DVDD.n18001 0.026913
R38152 DVDD.n18001 DVDD.n17999 0.026913
R38153 DVDD.n17999 DVDD.n17997 0.026913
R38154 DVDD.n17997 DVDD.n17995 0.026913
R38155 DVDD.n17995 DVDD.n17994 0.026913
R38156 DVDD.n17994 DVDD.n17992 0.026913
R38157 DVDD.n17992 DVDD.n17990 0.026913
R38158 DVDD.n17990 DVDD.n17988 0.026913
R38159 DVDD.n17988 DVDD.n17986 0.026913
R38160 DVDD.n17986 DVDD.n551 0.026913
R38161 DVDD.n17982 DVDD.n551 0.026913
R38162 DVDD.n17982 DVDD.n17981 0.026913
R38163 DVDD.n17981 DVDD.n553 0.026913
R38164 DVDD.n597 DVDD.n553 0.026913
R38165 DVDD.n599 DVDD.n597 0.026913
R38166 DVDD.n601 DVDD.n599 0.026913
R38167 DVDD.n603 DVDD.n601 0.026913
R38168 DVDD.n605 DVDD.n603 0.026913
R38169 DVDD.n607 DVDD.n605 0.026913
R38170 DVDD.n609 DVDD.n607 0.026913
R38171 DVDD.n610 DVDD.n609 0.026913
R38172 DVDD.n612 DVDD.n610 0.026913
R38173 DVDD.n614 DVDD.n612 0.026913
R38174 DVDD.n616 DVDD.n614 0.026913
R38175 DVDD.n618 DVDD.n616 0.026913
R38176 DVDD.n620 DVDD.n618 0.026913
R38177 DVDD.n622 DVDD.n620 0.026913
R38178 DVDD.n623 DVDD.n622 0.026913
R38179 DVDD.n626 DVDD.n623 0.026913
R38180 DVDD.n628 DVDD.n626 0.026913
R38181 DVDD.n630 DVDD.n628 0.026913
R38182 DVDD.n632 DVDD.n630 0.026913
R38183 DVDD.n634 DVDD.n632 0.026913
R38184 DVDD.n636 DVDD.n634 0.026913
R38185 DVDD.n637 DVDD.n636 0.026913
R38186 DVDD.n17975 DVDD.n637 0.026913
R38187 DVDD.n17975 DVDD.n17974 0.026913
R38188 DVDD.n17974 DVDD.n17973 0.026913
R38189 DVDD.n17973 DVDD.n17971 0.026913
R38190 DVDD.n17971 DVDD.n638 0.026913
R38191 DVDD.n17967 DVDD.n638 0.026913
R38192 DVDD.n17967 DVDD.n17966 0.026913
R38193 DVDD.n17966 DVDD.n640 0.026913
R38194 DVDD.n684 DVDD.n640 0.026913
R38195 DVDD.n685 DVDD.n684 0.026913
R38196 DVDD.n688 DVDD.n685 0.026913
R38197 DVDD.n690 DVDD.n688 0.026913
R38198 DVDD.n692 DVDD.n690 0.026913
R38199 DVDD.n694 DVDD.n692 0.026913
R38200 DVDD.n696 DVDD.n694 0.026913
R38201 DVDD.n698 DVDD.n696 0.026913
R38202 DVDD.n700 DVDD.n698 0.026913
R38203 DVDD.n701 DVDD.n700 0.026913
R38204 DVDD.n704 DVDD.n701 0.026913
R38205 DVDD.n706 DVDD.n704 0.026913
R38206 DVDD.n708 DVDD.n706 0.026913
R38207 DVDD.n710 DVDD.n708 0.026913
R38208 DVDD.n712 DVDD.n710 0.026913
R38209 DVDD.n714 DVDD.n712 0.026913
R38210 DVDD.n716 DVDD.n714 0.026913
R38211 DVDD.n717 DVDD.n716 0.026913
R38212 DVDD.n720 DVDD.n717 0.026913
R38213 DVDD.n722 DVDD.n720 0.026913
R38214 DVDD.n724 DVDD.n722 0.026913
R38215 DVDD.n726 DVDD.n724 0.026913
R38216 DVDD.n728 DVDD.n726 0.026913
R38217 DVDD.n729 DVDD.n728 0.026913
R38218 DVDD.n17960 DVDD.n729 0.026913
R38219 DVDD.n17960 DVDD.n17959 0.026913
R38220 DVDD.n17959 DVDD.n17958 0.026913
R38221 DVDD.n17958 DVDD.n730 0.026913
R38222 DVDD.n773 DVDD.n730 0.026913
R38223 DVDD.n774 DVDD.n773 0.026913
R38224 DVDD.n17951 DVDD.n774 0.026913
R38225 DVDD.n17951 DVDD.n17950 0.026913
R38226 DVDD.n17950 DVDD.n17948 0.026913
R38227 DVDD.n17948 DVDD.n17946 0.026913
R38228 DVDD.n17946 DVDD.n17944 0.026913
R38229 DVDD.n17944 DVDD.n17941 0.026913
R38230 DVDD.n17941 DVDD.n17940 0.026913
R38231 DVDD.n17940 DVDD.n17938 0.026913
R38232 DVDD.n17938 DVDD.n17936 0.026913
R38233 DVDD.n17936 DVDD.n17934 0.026913
R38234 DVDD.n17934 DVDD.n17932 0.026913
R38235 DVDD.n17932 DVDD.n17930 0.026913
R38236 DVDD.n17930 DVDD.n17928 0.026913
R38237 DVDD.n17928 DVDD.n17927 0.026913
R38238 DVDD.n17927 DVDD.n17925 0.026913
R38239 DVDD.n17925 DVDD.n17923 0.026913
R38240 DVDD.n17923 DVDD.n17921 0.026913
R38241 DVDD.n17921 DVDD.n17919 0.026913
R38242 DVDD.n17919 DVDD.n17917 0.026913
R38243 DVDD.n17917 DVDD.n17915 0.026913
R38244 DVDD.n17915 DVDD.n17912 0.026913
R38245 DVDD.n17912 DVDD.n17911 0.026913
R38246 DVDD.n17911 DVDD.n17909 0.026913
R38247 DVDD.n17909 DVDD.n17907 0.026913
R38248 DVDD.n17907 DVDD.n17905 0.026913
R38249 DVDD.n17905 DVDD.n775 0.026913
R38250 DVDD.n17901 DVDD.n775 0.026913
R38251 DVDD.n17901 DVDD.n17900 0.026913
R38252 DVDD.n17900 DVDD.n17899 0.026913
R38253 DVDD.n17899 DVDD.n777 0.026913
R38254 DVDD.n17895 DVDD.n17894 0.026913
R38255 DVDD.n17894 DVDD.n17893 0.026913
R38256 DVDD.n17893 DVDD.n780 0.026913
R38257 DVDD.n17889 DVDD.n780 0.026913
R38258 DVDD.n17889 DVDD.n17888 0.026913
R38259 DVDD.n17888 DVDD.n17887 0.026913
R38260 DVDD.n17887 DVDD.n782 0.026913
R38261 DVDD.n17883 DVDD.n782 0.026913
R38262 DVDD.n17883 DVDD.n17882 0.026913
R38263 DVDD.n17882 DVDD.n17881 0.026913
R38264 DVDD.n17881 DVDD.n784 0.026913
R38265 DVDD.n815 DVDD.n784 0.026913
R38266 DVDD.n817 DVDD.n815 0.026913
R38267 DVDD.n818 DVDD.n817 0.026913
R38268 DVDD.n821 DVDD.n818 0.026913
R38269 DVDD.n823 DVDD.n821 0.026913
R38270 DVDD.n825 DVDD.n823 0.026913
R38271 DVDD.n827 DVDD.n825 0.026913
R38272 DVDD.n829 DVDD.n827 0.026913
R38273 DVDD.n831 DVDD.n829 0.026913
R38274 DVDD.n832 DVDD.n831 0.026913
R38275 DVDD.n17874 DVDD.n832 0.026913
R38276 DVDD.n17874 DVDD.n17873 0.026913
R38277 DVDD.n17873 DVDD.n17872 0.026913
R38278 DVDD.n17872 DVDD.n833 0.026913
R38279 DVDD.n17868 DVDD.n833 0.026913
R38280 DVDD.n17868 DVDD.n17867 0.026913
R38281 DVDD.n17867 DVDD.n17866 0.026913
R38282 DVDD.n17866 DVDD.n835 0.026913
R38283 DVDD.n17862 DVDD.n835 0.026913
R38284 DVDD.n17862 DVDD.n17861 0.026913
R38285 DVDD.n17861 DVDD.n17860 0.026913
R38286 DVDD.n17860 DVDD.n837 0.026913
R38287 DVDD.n17856 DVDD.n837 0.026913
R38288 DVDD.n17856 DVDD.n17855 0.026913
R38289 DVDD.n17855 DVDD.n17854 0.026913
R38290 DVDD.n17854 DVDD.n839 0.026913
R38291 DVDD.n17850 DVDD.n839 0.026913
R38292 DVDD.n17850 DVDD.n17849 0.026913
R38293 DVDD.n17849 DVDD.n17848 0.026913
R38294 DVDD.n17848 DVDD.n841 0.026913
R38295 DVDD.n17844 DVDD.n841 0.026913
R38296 DVDD.n17844 DVDD.n17843 0.026913
R38297 DVDD.n17843 DVDD.n17842 0.026913
R38298 DVDD.n17842 DVDD.n843 0.026913
R38299 DVDD.n17838 DVDD.n843 0.026913
R38300 DVDD.n17838 DVDD.n17837 0.026913
R38301 DVDD.n17837 DVDD.n17836 0.026913
R38302 DVDD.n17836 DVDD.n845 0.026913
R38303 DVDD.n17832 DVDD.n845 0.026913
R38304 DVDD.n17832 DVDD.n17831 0.026913
R38305 DVDD.n17831 DVDD.n17830 0.026913
R38306 DVDD.n17830 DVDD.n847 0.026913
R38307 DVDD.n17826 DVDD.n847 0.026913
R38308 DVDD.n17826 DVDD.n17825 0.026913
R38309 DVDD.n17825 DVDD.n17824 0.026913
R38310 DVDD.n17824 DVDD.n849 0.026913
R38311 DVDD.n17820 DVDD.n849 0.026913
R38312 DVDD.n17820 DVDD.n17819 0.026913
R38313 DVDD.n17819 DVDD.n17818 0.026913
R38314 DVDD.n17818 DVDD.n851 0.026913
R38315 DVDD.n17814 DVDD.n851 0.026913
R38316 DVDD.n17814 DVDD.n17813 0.026913
R38317 DVDD.n17813 DVDD.n17812 0.026913
R38318 DVDD.n17812 DVDD.n853 0.026913
R38319 DVDD.n17808 DVDD.n853 0.026913
R38320 DVDD.n17808 DVDD.n17807 0.026913
R38321 DVDD.n17807 DVDD.n17806 0.026913
R38322 DVDD.n17806 DVDD.n855 0.026913
R38323 DVDD.n17802 DVDD.n855 0.026913
R38324 DVDD.n17802 DVDD.n17801 0.026913
R38325 DVDD.n17801 DVDD.n17800 0.026913
R38326 DVDD.n17800 DVDD.n857 0.026913
R38327 DVDD.n17796 DVDD.n857 0.026913
R38328 DVDD.n17796 DVDD.n17795 0.026913
R38329 DVDD.n17795 DVDD.n17794 0.026913
R38330 DVDD.n17794 DVDD.n859 0.026913
R38331 DVDD.n17790 DVDD.n859 0.026913
R38332 DVDD.n17790 DVDD.n17789 0.026913
R38333 DVDD.n17789 DVDD.n17788 0.026913
R38334 DVDD.n17788 DVDD.n861 0.026913
R38335 DVDD.n17784 DVDD.n861 0.026913
R38336 DVDD.n17784 DVDD.n17783 0.026913
R38337 DVDD.n17783 DVDD.n17782 0.026913
R38338 DVDD.n17782 DVDD.n863 0.026913
R38339 DVDD.n17778 DVDD.n863 0.026913
R38340 DVDD.n17778 DVDD.n17777 0.026913
R38341 DVDD.n17777 DVDD.n17776 0.026913
R38342 DVDD.n17776 DVDD.n865 0.026913
R38343 DVDD.n17772 DVDD.n865 0.026913
R38344 DVDD.n17772 DVDD.n17771 0.026913
R38345 DVDD.n17771 DVDD.n17770 0.026913
R38346 DVDD.n17770 DVDD.n867 0.026913
R38347 DVDD.n17766 DVDD.n867 0.026913
R38348 DVDD.n17766 DVDD.n17765 0.026913
R38349 DVDD.n17765 DVDD.n17764 0.026913
R38350 DVDD.n17764 DVDD.n869 0.026913
R38351 DVDD.n17760 DVDD.n869 0.026913
R38352 DVDD.n17760 DVDD.n17759 0.026913
R38353 DVDD.n17759 DVDD.n17758 0.026913
R38354 DVDD.n17758 DVDD.n871 0.026913
R38355 DVDD.n17754 DVDD.n871 0.026913
R38356 DVDD.n17754 DVDD.n17753 0.026913
R38357 DVDD.n17753 DVDD.n17752 0.026913
R38358 DVDD.n17752 DVDD.n873 0.026913
R38359 DVDD.n17748 DVDD.n873 0.026913
R38360 DVDD.n17748 DVDD.n17747 0.026913
R38361 DVDD.n17747 DVDD.n17746 0.026913
R38362 DVDD.n17746 DVDD.n875 0.026913
R38363 DVDD.n17742 DVDD.n875 0.026913
R38364 DVDD.n17742 DVDD.n17741 0.026913
R38365 DVDD.n17741 DVDD.n17740 0.026913
R38366 DVDD.n17740 DVDD.n877 0.026913
R38367 DVDD.n5006 DVDD.n5004 0.026913
R38368 DVDD.n5008 DVDD.n5006 0.026913
R38369 DVDD.n5010 DVDD.n5008 0.026913
R38370 DVDD.n5012 DVDD.n5010 0.026913
R38371 DVDD.n5014 DVDD.n5012 0.026913
R38372 DVDD.n5015 DVDD.n5014 0.026913
R38373 DVDD.n5018 DVDD.n5015 0.026913
R38374 DVDD.n5020 DVDD.n5018 0.026913
R38375 DVDD.n5022 DVDD.n5020 0.026913
R38376 DVDD.n5024 DVDD.n5022 0.026913
R38377 DVDD.n5026 DVDD.n5024 0.026913
R38378 DVDD.n5028 DVDD.n5026 0.026913
R38379 DVDD.n5030 DVDD.n5028 0.026913
R38380 DVDD.n5031 DVDD.n5030 0.026913
R38381 DVDD.n5033 DVDD.n5031 0.026913
R38382 DVDD.n5035 DVDD.n5033 0.026913
R38383 DVDD.n5037 DVDD.n5035 0.026913
R38384 DVDD.n5038 DVDD.n5037 0.026913
R38385 DVDD.n15705 DVDD.n5038 0.026913
R38386 DVDD.n15705 DVDD.n15704 0.026913
R38387 DVDD.n15704 DVDD.n15703 0.026913
R38388 DVDD.n15703 DVDD.n5039 0.026913
R38389 DVDD.n5262 DVDD.n5039 0.026913
R38390 DVDD.n5265 DVDD.n5262 0.026913
R38391 DVDD.n5267 DVDD.n5265 0.026913
R38392 DVDD.n5269 DVDD.n5267 0.026913
R38393 DVDD.n5271 DVDD.n5269 0.026913
R38394 DVDD.n5273 DVDD.n5271 0.026913
R38395 DVDD.n5275 DVDD.n5273 0.026913
R38396 DVDD.n5277 DVDD.n5275 0.026913
R38397 DVDD.n5278 DVDD.n5277 0.026913
R38398 DVDD.n5280 DVDD.n5278 0.026913
R38399 DVDD.n5282 DVDD.n5280 0.026913
R38400 DVDD.n5284 DVDD.n5282 0.026913
R38401 DVDD.n5286 DVDD.n5284 0.026913
R38402 DVDD.n5288 DVDD.n5286 0.026913
R38403 DVDD.n5290 DVDD.n5288 0.026913
R38404 DVDD.n5291 DVDD.n5290 0.026913
R38405 DVDD.n5294 DVDD.n5291 0.026913
R38406 DVDD.n5296 DVDD.n5294 0.026913
R38407 DVDD.n5298 DVDD.n5296 0.026913
R38408 DVDD.n5300 DVDD.n5298 0.026913
R38409 DVDD.n5302 DVDD.n5300 0.026913
R38410 DVDD.n5304 DVDD.n5302 0.026913
R38411 DVDD.n5306 DVDD.n5304 0.026913
R38412 DVDD.n5307 DVDD.n5306 0.026913
R38413 DVDD.n5310 DVDD.n5307 0.026913
R38414 DVDD.n5311 DVDD.n5310 0.026913
R38415 DVDD.n5312 DVDD.n5311 0.026913
R38416 DVDD.n5313 DVDD.n5312 0.026913
R38417 DVDD.n5316 DVDD.n5313 0.026913
R38418 DVDD.n5318 DVDD.n5316 0.026913
R38419 DVDD.n5320 DVDD.n5318 0.026913
R38420 DVDD.n5322 DVDD.n5320 0.026913
R38421 DVDD.n5323 DVDD.n5322 0.026913
R38422 DVDD.n5326 DVDD.n5323 0.026913
R38423 DVDD.n5328 DVDD.n5326 0.026913
R38424 DVDD.n5330 DVDD.n5328 0.026913
R38425 DVDD.n5332 DVDD.n5330 0.026913
R38426 DVDD.n5334 DVDD.n5332 0.026913
R38427 DVDD.n5336 DVDD.n5334 0.026913
R38428 DVDD.n5338 DVDD.n5336 0.026913
R38429 DVDD.n5339 DVDD.n5338 0.026913
R38430 DVDD.n5342 DVDD.n5339 0.026913
R38431 DVDD.n5344 DVDD.n5342 0.026913
R38432 DVDD.n5346 DVDD.n5344 0.026913
R38433 DVDD.n5348 DVDD.n5346 0.026913
R38434 DVDD.n5350 DVDD.n5348 0.026913
R38435 DVDD.n5352 DVDD.n5350 0.026913
R38436 DVDD.n5354 DVDD.n5352 0.026913
R38437 DVDD.n5355 DVDD.n5354 0.026913
R38438 DVDD.n5358 DVDD.n5355 0.026913
R38439 DVDD.n5360 DVDD.n5358 0.026913
R38440 DVDD.n5362 DVDD.n5360 0.026913
R38441 DVDD.n5364 DVDD.n5362 0.026913
R38442 DVDD.n5366 DVDD.n5364 0.026913
R38443 DVDD.n5367 DVDD.n5366 0.026913
R38444 DVDD.n15414 DVDD.n5367 0.026913
R38445 DVDD.n15414 DVDD.n15413 0.026913
R38446 DVDD.n15413 DVDD.n15412 0.026913
R38447 DVDD.n15412 DVDD.n5368 0.026913
R38448 DVDD.n5410 DVDD.n5368 0.026913
R38449 DVDD.n5412 DVDD.n5410 0.026913
R38450 DVDD.n5414 DVDD.n5412 0.026913
R38451 DVDD.n5416 DVDD.n5414 0.026913
R38452 DVDD.n5418 DVDD.n5416 0.026913
R38453 DVDD.n5420 DVDD.n5418 0.026913
R38454 DVDD.n5421 DVDD.n5420 0.026913
R38455 DVDD.n5424 DVDD.n5421 0.026913
R38456 DVDD.n5426 DVDD.n5424 0.026913
R38457 DVDD.n5428 DVDD.n5426 0.026913
R38458 DVDD.n5430 DVDD.n5428 0.026913
R38459 DVDD.n5432 DVDD.n5430 0.026913
R38460 DVDD.n5434 DVDD.n5432 0.026913
R38461 DVDD.n5436 DVDD.n5434 0.026913
R38462 DVDD.n5437 DVDD.n5436 0.026913
R38463 DVDD.n5439 DVDD.n5437 0.026913
R38464 DVDD.n5441 DVDD.n5439 0.026913
R38465 DVDD.n5443 DVDD.n5441 0.026913
R38466 DVDD.n5445 DVDD.n5443 0.026913
R38467 DVDD.n5447 DVDD.n5445 0.026913
R38468 DVDD.n5449 DVDD.n5447 0.026913
R38469 DVDD.n5450 DVDD.n5449 0.026913
R38470 DVDD.n5453 DVDD.n5450 0.026913
R38471 DVDD.n5455 DVDD.n5453 0.026913
R38472 DVDD.n5457 DVDD.n5455 0.026913
R38473 DVDD.n5458 DVDD.n5457 0.026913
R38474 DVDD.n15315 DVDD.n5458 0.026913
R38475 DVDD.n15315 DVDD.n15314 0.026913
R38476 DVDD.n15314 DVDD.n15313 0.026913
R38477 DVDD.n15313 DVDD.n5459 0.026913
R38478 DVDD.n15309 DVDD.n5459 0.026913
R38479 DVDD.n15309 DVDD.n15308 0.026913
R38480 DVDD.n15306 DVDD.n5461 0.026913
R38481 DVDD.n15302 DVDD.n5461 0.026913
R38482 DVDD.n15302 DVDD.n15301 0.026913
R38483 DVDD.n15301 DVDD.n15300 0.026913
R38484 DVDD.n15300 DVDD.n5463 0.026913
R38485 DVDD.n15296 DVDD.n5463 0.026913
R38486 DVDD.n15296 DVDD.n15295 0.026913
R38487 DVDD.n15295 DVDD.n15294 0.026913
R38488 DVDD.n15294 DVDD.n5465 0.026913
R38489 DVDD.n15290 DVDD.n5465 0.026913
R38490 DVDD.n15290 DVDD.n15289 0.026913
R38491 DVDD.n15289 DVDD.n15288 0.026913
R38492 DVDD.n15288 DVDD.n5467 0.026913
R38493 DVDD.n5498 DVDD.n5467 0.026913
R38494 DVDD.n5501 DVDD.n5498 0.026913
R38495 DVDD.n5503 DVDD.n5501 0.026913
R38496 DVDD.n5505 DVDD.n5503 0.026913
R38497 DVDD.n5507 DVDD.n5505 0.026913
R38498 DVDD.n5509 DVDD.n5507 0.026913
R38499 DVDD.n5511 DVDD.n5509 0.026913
R38500 DVDD.n5513 DVDD.n5511 0.026913
R38501 DVDD.n5515 DVDD.n5513 0.026913
R38502 DVDD.n5516 DVDD.n5515 0.026913
R38503 DVDD.n15282 DVDD.n5516 0.026913
R38504 DVDD.n15282 DVDD.n15281 0.026913
R38505 DVDD.n15281 DVDD.n15280 0.026913
R38506 DVDD.n15280 DVDD.n5517 0.026913
R38507 DVDD.n15276 DVDD.n5517 0.026913
R38508 DVDD.n15276 DVDD.n15275 0.026913
R38509 DVDD.n15275 DVDD.n15274 0.026913
R38510 DVDD.n15274 DVDD.n5519 0.026913
R38511 DVDD.n15270 DVDD.n5519 0.026913
R38512 DVDD.n15270 DVDD.n15269 0.026913
R38513 DVDD.n15269 DVDD.n15268 0.026913
R38514 DVDD.n15268 DVDD.n5521 0.026913
R38515 DVDD.n15264 DVDD.n5521 0.026913
R38516 DVDD.n15264 DVDD.n15263 0.026913
R38517 DVDD.n15263 DVDD.n15262 0.026913
R38518 DVDD.n15262 DVDD.n5523 0.026913
R38519 DVDD.n15258 DVDD.n5523 0.026913
R38520 DVDD.n15258 DVDD.n15257 0.026913
R38521 DVDD.n15257 DVDD.n15256 0.026913
R38522 DVDD.n15256 DVDD.n5525 0.026913
R38523 DVDD.n15252 DVDD.n5525 0.026913
R38524 DVDD.n15252 DVDD.n15251 0.026913
R38525 DVDD.n15251 DVDD.n15250 0.026913
R38526 DVDD.n15250 DVDD.n5527 0.026913
R38527 DVDD.n15246 DVDD.n5527 0.026913
R38528 DVDD.n15246 DVDD.n15245 0.026913
R38529 DVDD.n15245 DVDD.n15244 0.026913
R38530 DVDD.n15244 DVDD.n5529 0.026913
R38531 DVDD.n15240 DVDD.n5529 0.026913
R38532 DVDD.n15240 DVDD.n15239 0.026913
R38533 DVDD.n15239 DVDD.n15238 0.026913
R38534 DVDD.n15238 DVDD.n5531 0.026913
R38535 DVDD.n15234 DVDD.n5531 0.026913
R38536 DVDD.n15234 DVDD.n15233 0.026913
R38537 DVDD.n15233 DVDD.n15232 0.026913
R38538 DVDD.n15232 DVDD.n5533 0.026913
R38539 DVDD.n15228 DVDD.n5533 0.026913
R38540 DVDD.n15228 DVDD.n15227 0.026913
R38541 DVDD.n15227 DVDD.n15226 0.026913
R38542 DVDD.n15226 DVDD.n5535 0.026913
R38543 DVDD.n15222 DVDD.n5535 0.026913
R38544 DVDD.n15222 DVDD.n15221 0.026913
R38545 DVDD.n15221 DVDD.n15220 0.026913
R38546 DVDD.n15220 DVDD.n5537 0.026913
R38547 DVDD.n15216 DVDD.n5537 0.026913
R38548 DVDD.n15216 DVDD.n15215 0.026913
R38549 DVDD.n15215 DVDD.n15214 0.026913
R38550 DVDD.n15214 DVDD.n5539 0.026913
R38551 DVDD.n15210 DVDD.n5539 0.026913
R38552 DVDD.n15210 DVDD.n15209 0.026913
R38553 DVDD.n15209 DVDD.n15208 0.026913
R38554 DVDD.n15208 DVDD.n5541 0.026913
R38555 DVDD.n15204 DVDD.n5541 0.026913
R38556 DVDD.n15204 DVDD.n15203 0.026913
R38557 DVDD.n15203 DVDD.n15202 0.026913
R38558 DVDD.n15202 DVDD.n5543 0.026913
R38559 DVDD.n15198 DVDD.n5543 0.026913
R38560 DVDD.n15198 DVDD.n15197 0.026913
R38561 DVDD.n15197 DVDD.n15196 0.026913
R38562 DVDD.n15196 DVDD.n5545 0.026913
R38563 DVDD.n15192 DVDD.n5545 0.026913
R38564 DVDD.n15192 DVDD.n15191 0.026913
R38565 DVDD.n15191 DVDD.n15190 0.026913
R38566 DVDD.n15190 DVDD.n5547 0.026913
R38567 DVDD.n15186 DVDD.n5547 0.026913
R38568 DVDD.n15186 DVDD.n15185 0.026913
R38569 DVDD.n15185 DVDD.n15184 0.026913
R38570 DVDD.n15184 DVDD.n5549 0.026913
R38571 DVDD.n15180 DVDD.n5549 0.026913
R38572 DVDD.n15180 DVDD.n15179 0.026913
R38573 DVDD.n15179 DVDD.n15178 0.026913
R38574 DVDD.n15178 DVDD.n5551 0.026913
R38575 DVDD.n15174 DVDD.n5551 0.026913
R38576 DVDD.n15174 DVDD.n15173 0.026913
R38577 DVDD.n15173 DVDD.n15172 0.026913
R38578 DVDD.n15172 DVDD.n5553 0.026913
R38579 DVDD.n15168 DVDD.n5553 0.026913
R38580 DVDD.n15168 DVDD.n15167 0.026913
R38581 DVDD.n15167 DVDD.n15166 0.026913
R38582 DVDD.n15166 DVDD.n5555 0.026913
R38583 DVDD.n15162 DVDD.n5555 0.026913
R38584 DVDD.n15162 DVDD.n15161 0.026913
R38585 DVDD.n15161 DVDD.n15160 0.026913
R38586 DVDD.n15160 DVDD.n5557 0.026913
R38587 DVDD.n15156 DVDD.n5557 0.026913
R38588 DVDD.n15156 DVDD.n15155 0.026913
R38589 DVDD.n15155 DVDD.n15154 0.026913
R38590 DVDD.n15154 DVDD.n5559 0.026913
R38591 DVDD.n15150 DVDD.n5559 0.026913
R38592 DVDD.n15150 DVDD.n15149 0.026913
R38593 DVDD.n10200 DVDD.n10199 0.026913
R38594 DVDD.n10203 DVDD.n8971 0.026913
R38595 DVDD.n10221 DVDD.n8959 0.026913
R38596 DVDD.n8961 DVDD.n2291 0.026913
R38597 DVDD.n16429 DVDD.n16428 0.026913
R38598 DVDD.n16432 DVDD.n2278 0.026913
R38599 DVDD.n2269 DVDD.n2265 0.026913
R38600 DVDD.n16450 DVDD.n2266 0.026913
R38601 DVDD.n11929 DVDD.n2281 0.0268854
R38602 DVDD.n16452 DVDD.n16451 0.0268854
R38603 DVDD.n10223 DVDD.n10222 0.0268854
R38604 DVDD.n9572 DVDD.n9571 0.0268854
R38605 DVDD.n8026 DVDD.n7776 0.0266354
R38606 DVDD.n14834 DVDD.n14833 0.0266354
R38607 DVDD.n15082 DVDD.n7052 0.025925
R38608 DVDD.n1358 DVDD.n1259 0.0259118
R38609 DVDD.n7051 DVDD.n7042 0.0259118
R38610 DVDD.n7398 DVDD.n7052 0.0259118
R38611 DVDD.n15054 DVDD.n7407 0.0259118
R38612 DVDD.n7673 DVDD.n7661 0.0259118
R38613 DVDD.n9311 DVDD.n7674 0.0259118
R38614 DVDD.n8037 DVDD.n8023 0.0259118
R38615 DVDD.n14830 DVDD.n8038 0.0259118
R38616 DVDD.n14564 DVDD.n8158 0.0259118
R38617 DVDD.n8605 DVDD.n8598 0.0259118
R38618 DVDD.n8740 DVDD.n8606 0.0259118
R38619 DVDD.n10590 DVDD.n10576 0.0259118
R38620 DVDD.n14274 DVDD.n10591 0.0259118
R38621 DVDD.n11057 DVDD.n11050 0.0259118
R38622 DVDD.n13997 DVDD.n11058 0.0259118
R38623 DVDD.n13793 DVDD.n13792 0.0259118
R38624 DVDD.n13771 DVDD.n13770 0.0259118
R38625 DVDD.n12280 DVDD.n12277 0.0259118
R38626 DVDD.n13749 DVDD.n12281 0.0259118
R38627 DVDD.n12731 DVDD.n12725 0.0259118
R38628 DVDD.n13467 DVDD.n12732 0.0259118
R38629 DVDD.n13262 DVDD.n12915 0.0259118
R38630 DVDD.n16709 DVDD.n2159 0.0259118
R38631 DVDD.n1909 DVDD.n1808 0.0259118
R38632 DVDD.n16988 DVDD.n1709 0.0259118
R38633 DVDD.n17256 DVDD.n1608 0.0259118
R38634 DVDD.n6693 DVDD.n6344 0.0259118
R38635 DVDD.n6343 DVDD.n6337 0.0259118
R38636 DVDD.n1070 DVDD.n912 0.0259118
R38637 DVDD.n21845 DVDD.n21840 0.025475
R38638 DVDD.n21973 DVDD.n18274 0.025475
R38639 DVDD.n21237 DVDD.n21236 0.025475
R38640 DVDD.n21951 DVDD.n18292 0.025475
R38641 DVDD.n21826 DVDD.n21816 0.025475
R38642 DVDD.n18474 DVDD.n18464 0.025475
R38643 DVDD.n4304 DVDD.n4303 0.025475
R38644 DVDD.n3695 DVDD.n3694 0.025475
R38645 DVDD.n11057 DVDD.n11056 0.025475
R38646 DVDD.n17303 DVDD.n912 0.025475
R38647 DVDD.n21443 DVDD.n21442 0.0253684
R38648 DVDD.n18597 DVDD.n18595 0.0253684
R38649 DVDD.n19236 DVDD.n19232 0.0253684
R38650 DVDD.n19291 DVDD.n19289 0.0253684
R38651 DVDD.n16401 DVDD.n16400 0.0253032
R38652 DVDD.n16404 DVDD.n16403 0.0253032
R38653 DVDD.n17725 DVDD.n897 0.0251375
R38654 DVDD.n17312 DVDD.n898 0.0251375
R38655 DVDD.n15140 DVDD.n5583 0.0251375
R38656 DVDD.n5644 DVDD.n5584 0.0251375
R38657 DVDD.n8144 DVDD.n8042 0.0250633
R38658 DVDD.n8040 DVDD.n8025 0.0250633
R38659 DVDD.n13770 DVDD.n13769 0.025025
R38660 DVDD.n16732 DVDD.n1709 0.025025
R38661 DVDD.n20778 DVDD.n19033 0.0249537
R38662 DVDD.n20928 DVDD.n20926 0.0249537
R38663 DVDD.n20735 DVDD.n19129 0.0249537
R38664 DVDD.n20529 DVDD.n18859 0.0249537
R38665 DVDD.n12285 DVDD.n11941 0.0246703
R38666 DVDD.n2164 DVDD.n2157 0.0246703
R38667 DVDD.n12283 DVDD.n11943 0.0246703
R38668 DVDD.n2162 DVDD.n2158 0.0246703
R38669 DVDD.n8027 DVDD.n7674 0.024575
R38670 DVDD.n10579 DVDD.n10329 0.0242773
R38671 DVDD.n14278 DVDD.n14277 0.0242773
R38672 DVDD.n7047 DVDD.n6347 0.0238843
R38673 DVDD.n7048 DVDD.n6345 0.0238843
R38674 DVDD.n18413 DVDD.n18399 0.023675
R38675 DVDD.n22014 DVDD.n22010 0.023675
R38676 DVDD.n21342 DVDD.n21340 0.023675
R38677 DVDD.n18525 DVDD.n18521 0.023675
R38678 DVDD.n18253 DVDD.n18252 0.023675
R38679 DVDD.n18437 DVDD.n163 0.023675
R38680 DVDD.n4292 DVDD.n4291 0.023675
R38681 DVDD.n3682 DVDD.n3678 0.023675
R38682 DVDD.n14565 DVDD.n14564 0.022775
R38683 DVDD.n15080 DVDD.n7055 0.0227052
R38684 DVDD.n15081 DVDD.n7053 0.0227052
R38685 DVDD.n12731 DVDD.n12730 0.022325
R38686 DVDD.n13263 DVDD.n13262 0.022325
R38687 DVDD.n11054 DVDD.n10712 0.0223122
R38688 DVDD.n17301 DVDD.n914 0.0223122
R38689 DVDD.n11055 DVDD.n10714 0.0223122
R38690 DVDD.n17302 DVDD.n913 0.0223122
R38691 DVDD.n9789 DVDD.n9788 0.0219244
R38692 DVDD.n10102 DVDD.n9608 0.0219244
R38693 DVDD.n10103 DVDD.n10102 0.0219244
R38694 DVDD.n10103 DVDD.n9600 0.0219244
R38695 DVDD.n10115 DVDD.n9600 0.0219244
R38696 DVDD.n10116 DVDD.n10115 0.0219244
R38697 DVDD.n10127 DVDD.n9593 0.0219244
R38698 DVDD.n10128 DVDD.n10127 0.0219244
R38699 DVDD.n10128 DVDD.n9585 0.0219244
R38700 DVDD.n10140 DVDD.n9585 0.0219244
R38701 DVDD.n10141 DVDD.n10140 0.0219244
R38702 DVDD.n10141 DVDD.n9577 0.0219244
R38703 DVDD.n10153 DVDD.n9577 0.0219244
R38704 DVDD.n10157 DVDD.n10153 0.0219244
R38705 DVDD.n10157 DVDD.n10156 0.0219244
R38706 DVDD.n10156 DVDD.n2282 0.0219244
R38707 DVDD.n9786 DVDD.n9780 0.0219244
R38708 DVDD.n9740 DVDD.n9609 0.0219244
R38709 DVDD.n9609 DVDD.n9607 0.0219244
R38710 DVDD.n9607 DVDD.n9606 0.0219244
R38711 DVDD.n9606 DVDD.n9601 0.0219244
R38712 DVDD.n9601 DVDD.n9599 0.0219244
R38713 DVDD.n9598 DVDD.n9594 0.0219244
R38714 DVDD.n9594 DVDD.n9592 0.0219244
R38715 DVDD.n9592 DVDD.n9591 0.0219244
R38716 DVDD.n9591 DVDD.n9586 0.0219244
R38717 DVDD.n9586 DVDD.n9584 0.0219244
R38718 DVDD.n9584 DVDD.n9583 0.0219244
R38719 DVDD.n9583 DVDD.n9578 0.0219244
R38720 DVDD.n9578 DVDD.n9576 0.0219244
R38721 DVDD.n10154 DVDD.n9576 0.0219244
R38722 DVDD.n10154 DVDD.n2268 0.0219244
R38723 DVDD.n9793 DVDD.n9792 0.0219244
R38724 DVDD.n10095 DVDD.n9604 0.0219244
R38725 DVDD.n10107 DVDD.n9604 0.0219244
R38726 DVDD.n10108 DVDD.n10107 0.0219244
R38727 DVDD.n10108 DVDD.n9596 0.0219244
R38728 DVDD.n10119 DVDD.n9596 0.0219244
R38729 DVDD.n10120 DVDD.n9589 0.0219244
R38730 DVDD.n10132 DVDD.n9589 0.0219244
R38731 DVDD.n10133 DVDD.n10132 0.0219244
R38732 DVDD.n10133 DVDD.n9581 0.0219244
R38733 DVDD.n10145 DVDD.n9581 0.0219244
R38734 DVDD.n10146 DVDD.n10145 0.0219244
R38735 DVDD.n10146 DVDD.n9575 0.0219244
R38736 DVDD.n10161 DVDD.n9575 0.0219244
R38737 DVDD.n10162 DVDD.n10161 0.0219244
R38738 DVDD.n10162 DVDD.n8962 0.0219244
R38739 DVDD.n9795 DVDD.n9775 0.0219244
R38740 DVDD.n10098 DVDD.n10097 0.0219244
R38741 DVDD.n10098 DVDD.n9602 0.0219244
R38742 DVDD.n10110 DVDD.n9602 0.0219244
R38743 DVDD.n10111 DVDD.n10110 0.0219244
R38744 DVDD.n10111 DVDD.n9595 0.0219244
R38745 DVDD.n10123 DVDD.n10122 0.0219244
R38746 DVDD.n10123 DVDD.n9587 0.0219244
R38747 DVDD.n10135 DVDD.n9587 0.0219244
R38748 DVDD.n10136 DVDD.n10135 0.0219244
R38749 DVDD.n10136 DVDD.n9579 0.0219244
R38750 DVDD.n10148 DVDD.n9579 0.0219244
R38751 DVDD.n10149 DVDD.n10148 0.0219244
R38752 DVDD.n10149 DVDD.n9573 0.0219244
R38753 DVDD.n10164 DVDD.n9573 0.0219244
R38754 DVDD.n10167 DVDD.n10164 0.0219244
R38755 DVDD.n13767 DVDD.n11632 0.0219192
R38756 DVDD.n16734 DVDD.n1711 0.0219192
R38757 DVDD.n13768 DVDD.n11922 0.0219192
R38758 DVDD.n16733 DVDD.n1710 0.0219192
R38759 DVDD.n10580 DVDD.n8606 0.021875
R38760 DVDD.n19418 DVDD 0.0218158
R38761 DVDD.n21971 DVDD.n21970 0.0218
R38762 DVDD.n21970 DVDD.n209 0.0218
R38763 DVDD.n22017 DVDD.n220 0.0218
R38764 DVDD.n22018 DVDD.n22017 0.0218
R38765 DVDD.n21242 DVDD.n21241 0.0218
R38766 DVDD.n21241 DVDD.n18503 0.0218
R38767 DVDD.n21350 DVDD.n18506 0.0218
R38768 DVDD.n21350 DVDD.n21349 0.0218
R38769 DVDD.n21700 DVDD.n21698 0.0218
R38770 DVDD.n21700 DVDD.n21699 0.0218
R38771 DVDD.n21954 DVDD.n18290 0.0218
R38772 DVDD.n21955 DVDD.n21954 0.0218
R38773 DVDD.n21824 DVDD.n21823 0.0218
R38774 DVDD.n21823 DVDD.n216 0.0218
R38775 DVDD.n18260 DVDD.n212 0.0218
R38776 DVDD.n18260 DVDD.n18259 0.0218
R38777 DVDD.n18418 DVDD.n18417 0.0218
R38778 DVDD.n18417 DVDD.n18416 0.0218
R38779 DVDD.n21851 DVDD.n21847 0.0218
R38780 DVDD.n21852 DVDD.n21851 0.0218
R38781 DVDD.n18472 DVDD.n18471 0.0218
R38782 DVDD.n18471 DVDD.n18448 0.0218
R38783 DVDD.n18447 DVDD.n18435 0.0218
R38784 DVDD.n18443 DVDD.n18435 0.0218
R38785 DVDD.n4295 DVDD.n4294 0.0218
R38786 DVDD.n4296 DVDD.n4295 0.0218
R38787 DVDD.n4312 DVDD.n4311 0.0218
R38788 DVDD.n4311 DVDD.n4310 0.0218
R38789 DVDD.n3689 DVDD.n3687 0.0218
R38790 DVDD.n3689 DVDD.n3688 0.0218
R38791 DVDD.n3704 DVDD.n3697 0.0218
R38792 DVDD.n3704 DVDD.n3703 0.0218
R38793 DVDD.n8031 DVDD.n7677 0.0215262
R38794 DVDD.n8028 DVDD.n7675 0.0215262
R38795 DVDD.n21849 DVDD.n21848 0.021425
R38796 DVDD.n18276 DVDD.n18268 0.021425
R38797 DVDD.n21238 DVDD.n18663 0.021425
R38798 DVDD.n21952 DVDD.n18291 0.021425
R38799 DVDD.n21819 DVDD.n21801 0.021425
R38800 DVDD.n18467 DVDD.n18459 0.021425
R38801 DVDD.n4302 DVDD.n4299 0.021425
R38802 DVDD.n3707 DVDD.n3706 0.021425
R38803 DVDD.n15107 DVDD.n6343 0.021425
R38804 DVDD.n15064 DVDD.n7407 0.020075
R38805 DVDD.n14567 DVDD.n8156 0.0199541
R38806 DVDD.n14566 DVDD.n8157 0.0199541
R38807 DVDD.n15091 DVDD.n6750 0.019716
R38808 DVDD.n6856 DVDD.n6793 0.019716
R38809 DVDD.n6856 DVDD.n6748 0.019716
R38810 DVDD.n6865 DVDD.n6792 0.019716
R38811 DVDD.n6865 DVDD.n6747 0.019716
R38812 DVDD.n6853 DVDD.n6791 0.019716
R38813 DVDD.n6853 DVDD.n6746 0.019716
R38814 DVDD.n6874 DVDD.n6790 0.019716
R38815 DVDD.n6874 DVDD.n6745 0.019716
R38816 DVDD.n6850 DVDD.n6789 0.019716
R38817 DVDD.n6850 DVDD.n6744 0.019716
R38818 DVDD.n6883 DVDD.n6788 0.019716
R38819 DVDD.n6883 DVDD.n6743 0.019716
R38820 DVDD.n6847 DVDD.n6787 0.019716
R38821 DVDD.n6847 DVDD.n6742 0.019716
R38822 DVDD.n6892 DVDD.n6786 0.019716
R38823 DVDD.n6892 DVDD.n6741 0.019716
R38824 DVDD.n6844 DVDD.n6785 0.019716
R38825 DVDD.n6844 DVDD.n6740 0.019716
R38826 DVDD.n6901 DVDD.n6784 0.019716
R38827 DVDD.n6901 DVDD.n6739 0.019716
R38828 DVDD.n6841 DVDD.n6783 0.019716
R38829 DVDD.n6841 DVDD.n6738 0.019716
R38830 DVDD.n6910 DVDD.n6782 0.019716
R38831 DVDD.n6910 DVDD.n6737 0.019716
R38832 DVDD.n6838 DVDD.n6781 0.019716
R38833 DVDD.n6838 DVDD.n6736 0.019716
R38834 DVDD.n6919 DVDD.n6780 0.019716
R38835 DVDD.n6919 DVDD.n6735 0.019716
R38836 DVDD.n6835 DVDD.n6779 0.019716
R38837 DVDD.n6835 DVDD.n6734 0.019716
R38838 DVDD.n6928 DVDD.n6778 0.019716
R38839 DVDD.n6928 DVDD.n6733 0.019716
R38840 DVDD.n6832 DVDD.n6777 0.019716
R38841 DVDD.n6832 DVDD.n6732 0.019716
R38842 DVDD.n6937 DVDD.n6776 0.019716
R38843 DVDD.n6937 DVDD.n6731 0.019716
R38844 DVDD.n6829 DVDD.n6775 0.019716
R38845 DVDD.n6829 DVDD.n6730 0.019716
R38846 DVDD.n6946 DVDD.n6774 0.019716
R38847 DVDD.n6946 DVDD.n6729 0.019716
R38848 DVDD.n6826 DVDD.n6773 0.019716
R38849 DVDD.n6826 DVDD.n6728 0.019716
R38850 DVDD.n6955 DVDD.n6772 0.019716
R38851 DVDD.n6955 DVDD.n6727 0.019716
R38852 DVDD.n6823 DVDD.n6771 0.019716
R38853 DVDD.n6823 DVDD.n6726 0.019716
R38854 DVDD.n6964 DVDD.n6770 0.019716
R38855 DVDD.n6964 DVDD.n6725 0.019716
R38856 DVDD.n6820 DVDD.n6769 0.019716
R38857 DVDD.n6820 DVDD.n6724 0.019716
R38858 DVDD.n6973 DVDD.n6768 0.019716
R38859 DVDD.n6973 DVDD.n6723 0.019716
R38860 DVDD.n6817 DVDD.n6767 0.019716
R38861 DVDD.n6817 DVDD.n6722 0.019716
R38862 DVDD.n6982 DVDD.n6766 0.019716
R38863 DVDD.n6982 DVDD.n6721 0.019716
R38864 DVDD.n6814 DVDD.n6765 0.019716
R38865 DVDD.n6814 DVDD.n6720 0.019716
R38866 DVDD.n6991 DVDD.n6764 0.019716
R38867 DVDD.n6991 DVDD.n6719 0.019716
R38868 DVDD.n6811 DVDD.n6763 0.019716
R38869 DVDD.n6811 DVDD.n6718 0.019716
R38870 DVDD.n7000 DVDD.n6762 0.019716
R38871 DVDD.n7000 DVDD.n6717 0.019716
R38872 DVDD.n6808 DVDD.n6761 0.019716
R38873 DVDD.n6808 DVDD.n6716 0.019716
R38874 DVDD.n7009 DVDD.n6760 0.019716
R38875 DVDD.n7009 DVDD.n6715 0.019716
R38876 DVDD.n6805 DVDD.n6759 0.019716
R38877 DVDD.n6805 DVDD.n6714 0.019716
R38878 DVDD.n7018 DVDD.n6758 0.019716
R38879 DVDD.n7018 DVDD.n6713 0.019716
R38880 DVDD.n6802 DVDD.n6757 0.019716
R38881 DVDD.n6802 DVDD.n6712 0.019716
R38882 DVDD.n7027 DVDD.n6756 0.019716
R38883 DVDD.n7027 DVDD.n6711 0.019716
R38884 DVDD.n6799 DVDD.n6755 0.019716
R38885 DVDD.n6799 DVDD.n6710 0.019716
R38886 DVDD.n7036 DVDD.n6754 0.019716
R38887 DVDD.n7036 DVDD.n6709 0.019716
R38888 DVDD.n6796 DVDD.n6753 0.019716
R38889 DVDD.n6796 DVDD.n6708 0.019716
R38890 DVDD.n7155 DVDD.n7154 0.019716
R38891 DVDD.n7160 DVDD.n7110 0.019716
R38892 DVDD.n7161 DVDD.n7160 0.019716
R38893 DVDD.n7166 DVDD.n7109 0.019716
R38894 DVDD.n7166 DVDD.n7165 0.019716
R38895 DVDD.n7172 DVDD.n7108 0.019716
R38896 DVDD.n7173 DVDD.n7172 0.019716
R38897 DVDD.n7178 DVDD.n7107 0.019716
R38898 DVDD.n7178 DVDD.n7177 0.019716
R38899 DVDD.n7184 DVDD.n7106 0.019716
R38900 DVDD.n7185 DVDD.n7184 0.019716
R38901 DVDD.n7190 DVDD.n7105 0.019716
R38902 DVDD.n7190 DVDD.n7189 0.019716
R38903 DVDD.n7196 DVDD.n7104 0.019716
R38904 DVDD.n7197 DVDD.n7196 0.019716
R38905 DVDD.n7202 DVDD.n7103 0.019716
R38906 DVDD.n7202 DVDD.n7201 0.019716
R38907 DVDD.n7208 DVDD.n7102 0.019716
R38908 DVDD.n7209 DVDD.n7208 0.019716
R38909 DVDD.n7214 DVDD.n7101 0.019716
R38910 DVDD.n7214 DVDD.n7213 0.019716
R38911 DVDD.n7220 DVDD.n7100 0.019716
R38912 DVDD.n7221 DVDD.n7220 0.019716
R38913 DVDD.n7226 DVDD.n7099 0.019716
R38914 DVDD.n7226 DVDD.n7225 0.019716
R38915 DVDD.n7232 DVDD.n7098 0.019716
R38916 DVDD.n7233 DVDD.n7232 0.019716
R38917 DVDD.n7238 DVDD.n7097 0.019716
R38918 DVDD.n7238 DVDD.n7237 0.019716
R38919 DVDD.n7244 DVDD.n7096 0.019716
R38920 DVDD.n7245 DVDD.n7244 0.019716
R38921 DVDD.n7250 DVDD.n7095 0.019716
R38922 DVDD.n7250 DVDD.n7249 0.019716
R38923 DVDD.n7256 DVDD.n7094 0.019716
R38924 DVDD.n7257 DVDD.n7256 0.019716
R38925 DVDD.n7262 DVDD.n7093 0.019716
R38926 DVDD.n7262 DVDD.n7261 0.019716
R38927 DVDD.n7268 DVDD.n7092 0.019716
R38928 DVDD.n7269 DVDD.n7268 0.019716
R38929 DVDD.n7274 DVDD.n7091 0.019716
R38930 DVDD.n7274 DVDD.n7273 0.019716
R38931 DVDD.n7280 DVDD.n7090 0.019716
R38932 DVDD.n7281 DVDD.n7280 0.019716
R38933 DVDD.n7286 DVDD.n7089 0.019716
R38934 DVDD.n7286 DVDD.n7285 0.019716
R38935 DVDD.n7292 DVDD.n7088 0.019716
R38936 DVDD.n7293 DVDD.n7292 0.019716
R38937 DVDD.n7298 DVDD.n7087 0.019716
R38938 DVDD.n7298 DVDD.n7297 0.019716
R38939 DVDD.n7304 DVDD.n7086 0.019716
R38940 DVDD.n7305 DVDD.n7304 0.019716
R38941 DVDD.n7310 DVDD.n7085 0.019716
R38942 DVDD.n7310 DVDD.n7309 0.019716
R38943 DVDD.n7316 DVDD.n7084 0.019716
R38944 DVDD.n7317 DVDD.n7316 0.019716
R38945 DVDD.n7322 DVDD.n7083 0.019716
R38946 DVDD.n7322 DVDD.n7321 0.019716
R38947 DVDD.n7328 DVDD.n7082 0.019716
R38948 DVDD.n7329 DVDD.n7328 0.019716
R38949 DVDD.n7334 DVDD.n7081 0.019716
R38950 DVDD.n7334 DVDD.n7333 0.019716
R38951 DVDD.n7340 DVDD.n7080 0.019716
R38952 DVDD.n7341 DVDD.n7340 0.019716
R38953 DVDD.n7346 DVDD.n7079 0.019716
R38954 DVDD.n7346 DVDD.n7345 0.019716
R38955 DVDD.n7352 DVDD.n7078 0.019716
R38956 DVDD.n7353 DVDD.n7352 0.019716
R38957 DVDD.n7358 DVDD.n7077 0.019716
R38958 DVDD.n7358 DVDD.n7357 0.019716
R38959 DVDD.n7364 DVDD.n7076 0.019716
R38960 DVDD.n7365 DVDD.n7364 0.019716
R38961 DVDD.n7370 DVDD.n7075 0.019716
R38962 DVDD.n7370 DVDD.n7369 0.019716
R38963 DVDD.n7376 DVDD.n7074 0.019716
R38964 DVDD.n7377 DVDD.n7376 0.019716
R38965 DVDD.n7382 DVDD.n7073 0.019716
R38966 DVDD.n7382 DVDD.n7381 0.019716
R38967 DVDD.n7388 DVDD.n7072 0.019716
R38968 DVDD.n7389 DVDD.n7388 0.019716
R38969 DVDD.n7394 DVDD.n7071 0.019716
R38970 DVDD.n7394 DVDD.n7393 0.019716
R38971 DVDD.n7401 DVDD.n7070 0.019716
R38972 DVDD.n7402 DVDD.n7401 0.019716
R38973 DVDD.n15059 DVDD.n7455 0.019716
R38974 DVDD.n7561 DVDD.n7499 0.019716
R38975 DVDD.n7561 DVDD.n7453 0.019716
R38976 DVDD.n14877 DVDD.n7498 0.019716
R38977 DVDD.n14877 DVDD.n7452 0.019716
R38978 DVDD.n7558 DVDD.n7497 0.019716
R38979 DVDD.n7558 DVDD.n7451 0.019716
R38980 DVDD.n14886 DVDD.n7496 0.019716
R38981 DVDD.n14886 DVDD.n7450 0.019716
R38982 DVDD.n7555 DVDD.n7495 0.019716
R38983 DVDD.n7555 DVDD.n7449 0.019716
R38984 DVDD.n14895 DVDD.n7494 0.019716
R38985 DVDD.n14895 DVDD.n7448 0.019716
R38986 DVDD.n7552 DVDD.n7493 0.019716
R38987 DVDD.n7552 DVDD.n7447 0.019716
R38988 DVDD.n14904 DVDD.n7492 0.019716
R38989 DVDD.n14904 DVDD.n7446 0.019716
R38990 DVDD.n7549 DVDD.n7491 0.019716
R38991 DVDD.n7549 DVDD.n7445 0.019716
R38992 DVDD.n14913 DVDD.n7490 0.019716
R38993 DVDD.n14913 DVDD.n7444 0.019716
R38994 DVDD.n7546 DVDD.n7489 0.019716
R38995 DVDD.n7546 DVDD.n7443 0.019716
R38996 DVDD.n14922 DVDD.n7488 0.019716
R38997 DVDD.n14922 DVDD.n7442 0.019716
R38998 DVDD.n7543 DVDD.n7487 0.019716
R38999 DVDD.n7543 DVDD.n7441 0.019716
R39000 DVDD.n14931 DVDD.n7486 0.019716
R39001 DVDD.n14931 DVDD.n7440 0.019716
R39002 DVDD.n7540 DVDD.n7485 0.019716
R39003 DVDD.n7540 DVDD.n7439 0.019716
R39004 DVDD.n14940 DVDD.n7484 0.019716
R39005 DVDD.n14940 DVDD.n7438 0.019716
R39006 DVDD.n7537 DVDD.n7483 0.019716
R39007 DVDD.n7537 DVDD.n7437 0.019716
R39008 DVDD.n14949 DVDD.n7482 0.019716
R39009 DVDD.n14949 DVDD.n7436 0.019716
R39010 DVDD.n7534 DVDD.n7481 0.019716
R39011 DVDD.n7534 DVDD.n7435 0.019716
R39012 DVDD.n14958 DVDD.n7480 0.019716
R39013 DVDD.n14958 DVDD.n7434 0.019716
R39014 DVDD.n7531 DVDD.n7479 0.019716
R39015 DVDD.n7531 DVDD.n7433 0.019716
R39016 DVDD.n14967 DVDD.n7478 0.019716
R39017 DVDD.n14967 DVDD.n7432 0.019716
R39018 DVDD.n7528 DVDD.n7477 0.019716
R39019 DVDD.n7528 DVDD.n7431 0.019716
R39020 DVDD.n14976 DVDD.n7476 0.019716
R39021 DVDD.n14976 DVDD.n7430 0.019716
R39022 DVDD.n7525 DVDD.n7475 0.019716
R39023 DVDD.n7525 DVDD.n7429 0.019716
R39024 DVDD.n14985 DVDD.n7474 0.019716
R39025 DVDD.n14985 DVDD.n7428 0.019716
R39026 DVDD.n7522 DVDD.n7473 0.019716
R39027 DVDD.n7522 DVDD.n7427 0.019716
R39028 DVDD.n14994 DVDD.n7472 0.019716
R39029 DVDD.n14994 DVDD.n7426 0.019716
R39030 DVDD.n7519 DVDD.n7471 0.019716
R39031 DVDD.n7519 DVDD.n7425 0.019716
R39032 DVDD.n15003 DVDD.n7470 0.019716
R39033 DVDD.n15003 DVDD.n7424 0.019716
R39034 DVDD.n7516 DVDD.n7469 0.019716
R39035 DVDD.n7516 DVDD.n7423 0.019716
R39036 DVDD.n15012 DVDD.n7468 0.019716
R39037 DVDD.n15012 DVDD.n7422 0.019716
R39038 DVDD.n7513 DVDD.n7467 0.019716
R39039 DVDD.n7513 DVDD.n7421 0.019716
R39040 DVDD.n15021 DVDD.n7466 0.019716
R39041 DVDD.n15021 DVDD.n7420 0.019716
R39042 DVDD.n7510 DVDD.n7465 0.019716
R39043 DVDD.n7510 DVDD.n7419 0.019716
R39044 DVDD.n15030 DVDD.n7464 0.019716
R39045 DVDD.n15030 DVDD.n7418 0.019716
R39046 DVDD.n7507 DVDD.n7463 0.019716
R39047 DVDD.n7507 DVDD.n7417 0.019716
R39048 DVDD.n15039 DVDD.n7462 0.019716
R39049 DVDD.n15039 DVDD.n7416 0.019716
R39050 DVDD.n7504 DVDD.n7461 0.019716
R39051 DVDD.n7504 DVDD.n7415 0.019716
R39052 DVDD.n15048 DVDD.n7460 0.019716
R39053 DVDD.n15048 DVDD.n7414 0.019716
R39054 DVDD.n7501 DVDD.n7459 0.019716
R39055 DVDD.n7501 DVDD.n7413 0.019716
R39056 DVDD.n14862 DVDD.n7612 0.019716
R39057 DVDD.n9214 DVDD.n7656 0.019716
R39058 DVDD.n9214 DVDD.n7610 0.019716
R39059 DVDD.n8976 DVDD.n7655 0.019716
R39060 DVDD.n8976 DVDD.n7609 0.019716
R39061 DVDD.n9205 DVDD.n7654 0.019716
R39062 DVDD.n9205 DVDD.n7608 0.019716
R39063 DVDD.n8979 DVDD.n7653 0.019716
R39064 DVDD.n8979 DVDD.n7607 0.019716
R39065 DVDD.n9196 DVDD.n7652 0.019716
R39066 DVDD.n9196 DVDD.n7606 0.019716
R39067 DVDD.n8982 DVDD.n7651 0.019716
R39068 DVDD.n8982 DVDD.n7605 0.019716
R39069 DVDD.n9187 DVDD.n7650 0.019716
R39070 DVDD.n9187 DVDD.n7604 0.019716
R39071 DVDD.n8985 DVDD.n7649 0.019716
R39072 DVDD.n8985 DVDD.n7603 0.019716
R39073 DVDD.n9178 DVDD.n7648 0.019716
R39074 DVDD.n9178 DVDD.n7602 0.019716
R39075 DVDD.n8988 DVDD.n7647 0.019716
R39076 DVDD.n8988 DVDD.n7601 0.019716
R39077 DVDD.n9169 DVDD.n7646 0.019716
R39078 DVDD.n9169 DVDD.n7600 0.019716
R39079 DVDD.n8991 DVDD.n7645 0.019716
R39080 DVDD.n8991 DVDD.n7599 0.019716
R39081 DVDD.n9160 DVDD.n7644 0.019716
R39082 DVDD.n9160 DVDD.n7598 0.019716
R39083 DVDD.n8994 DVDD.n7643 0.019716
R39084 DVDD.n8994 DVDD.n7597 0.019716
R39085 DVDD.n9151 DVDD.n7642 0.019716
R39086 DVDD.n9151 DVDD.n7596 0.019716
R39087 DVDD.n8997 DVDD.n7641 0.019716
R39088 DVDD.n8997 DVDD.n7595 0.019716
R39089 DVDD.n9142 DVDD.n7640 0.019716
R39090 DVDD.n9142 DVDD.n7594 0.019716
R39091 DVDD.n9000 DVDD.n7639 0.019716
R39092 DVDD.n9000 DVDD.n7593 0.019716
R39093 DVDD.n9133 DVDD.n7638 0.019716
R39094 DVDD.n9133 DVDD.n7592 0.019716
R39095 DVDD.n9003 DVDD.n7637 0.019716
R39096 DVDD.n9003 DVDD.n7591 0.019716
R39097 DVDD.n9124 DVDD.n7636 0.019716
R39098 DVDD.n9124 DVDD.n7590 0.019716
R39099 DVDD.n9006 DVDD.n7635 0.019716
R39100 DVDD.n9006 DVDD.n7589 0.019716
R39101 DVDD.n9115 DVDD.n7634 0.019716
R39102 DVDD.n9115 DVDD.n7588 0.019716
R39103 DVDD.n9009 DVDD.n7633 0.019716
R39104 DVDD.n9009 DVDD.n7587 0.019716
R39105 DVDD.n9106 DVDD.n7632 0.019716
R39106 DVDD.n9106 DVDD.n7586 0.019716
R39107 DVDD.n9012 DVDD.n7631 0.019716
R39108 DVDD.n9012 DVDD.n7585 0.019716
R39109 DVDD.n9097 DVDD.n7630 0.019716
R39110 DVDD.n9097 DVDD.n7584 0.019716
R39111 DVDD.n9015 DVDD.n7629 0.019716
R39112 DVDD.n9015 DVDD.n7583 0.019716
R39113 DVDD.n9088 DVDD.n7628 0.019716
R39114 DVDD.n9088 DVDD.n7582 0.019716
R39115 DVDD.n9018 DVDD.n7627 0.019716
R39116 DVDD.n9018 DVDD.n7581 0.019716
R39117 DVDD.n9079 DVDD.n7626 0.019716
R39118 DVDD.n9079 DVDD.n7580 0.019716
R39119 DVDD.n9021 DVDD.n7625 0.019716
R39120 DVDD.n9021 DVDD.n7579 0.019716
R39121 DVDD.n9070 DVDD.n7624 0.019716
R39122 DVDD.n9070 DVDD.n7578 0.019716
R39123 DVDD.n9024 DVDD.n7623 0.019716
R39124 DVDD.n9024 DVDD.n7577 0.019716
R39125 DVDD.n9061 DVDD.n7622 0.019716
R39126 DVDD.n9061 DVDD.n7576 0.019716
R39127 DVDD.n9027 DVDD.n7621 0.019716
R39128 DVDD.n9027 DVDD.n7575 0.019716
R39129 DVDD.n9052 DVDD.n7620 0.019716
R39130 DVDD.n9052 DVDD.n7574 0.019716
R39131 DVDD.n9030 DVDD.n7619 0.019716
R39132 DVDD.n9030 DVDD.n7573 0.019716
R39133 DVDD.n9043 DVDD.n7618 0.019716
R39134 DVDD.n9043 DVDD.n7572 0.019716
R39135 DVDD.n9033 DVDD.n7617 0.019716
R39136 DVDD.n9033 DVDD.n7571 0.019716
R39137 DVDD.n7659 DVDD.n7616 0.019716
R39138 DVDD.n7659 DVDD.n7570 0.019716
R39139 DVDD.n9557 DVDD.n9264 0.019716
R39140 DVDD.n9267 DVDD.n9266 0.019716
R39141 DVDD.n9267 DVDD.n9263 0.019716
R39142 DVDD.n9548 DVDD.n9547 0.019716
R39143 DVDD.n9547 DVDD.n9262 0.019716
R39144 DVDD.n9543 DVDD.n9542 0.019716
R39145 DVDD.n9542 DVDD.n9261 0.019716
R39146 DVDD.n9536 DVDD.n9535 0.019716
R39147 DVDD.n9535 DVDD.n9260 0.019716
R39148 DVDD.n9531 DVDD.n9530 0.019716
R39149 DVDD.n9530 DVDD.n9259 0.019716
R39150 DVDD.n9524 DVDD.n9523 0.019716
R39151 DVDD.n9523 DVDD.n9258 0.019716
R39152 DVDD.n9519 DVDD.n9518 0.019716
R39153 DVDD.n9518 DVDD.n9257 0.019716
R39154 DVDD.n9512 DVDD.n9511 0.019716
R39155 DVDD.n9511 DVDD.n9256 0.019716
R39156 DVDD.n9507 DVDD.n9506 0.019716
R39157 DVDD.n9506 DVDD.n9255 0.019716
R39158 DVDD.n9500 DVDD.n9499 0.019716
R39159 DVDD.n9499 DVDD.n9254 0.019716
R39160 DVDD.n9495 DVDD.n9494 0.019716
R39161 DVDD.n9494 DVDD.n9253 0.019716
R39162 DVDD.n9488 DVDD.n9487 0.019716
R39163 DVDD.n9487 DVDD.n9252 0.019716
R39164 DVDD.n9483 DVDD.n9482 0.019716
R39165 DVDD.n9482 DVDD.n9251 0.019716
R39166 DVDD.n9476 DVDD.n9475 0.019716
R39167 DVDD.n9475 DVDD.n9250 0.019716
R39168 DVDD.n9471 DVDD.n9470 0.019716
R39169 DVDD.n9470 DVDD.n9249 0.019716
R39170 DVDD.n9464 DVDD.n9463 0.019716
R39171 DVDD.n9463 DVDD.n9248 0.019716
R39172 DVDD.n9459 DVDD.n9458 0.019716
R39173 DVDD.n9458 DVDD.n9247 0.019716
R39174 DVDD.n9452 DVDD.n9451 0.019716
R39175 DVDD.n9451 DVDD.n9246 0.019716
R39176 DVDD.n9447 DVDD.n9446 0.019716
R39177 DVDD.n9446 DVDD.n9245 0.019716
R39178 DVDD.n9440 DVDD.n9439 0.019716
R39179 DVDD.n9439 DVDD.n9244 0.019716
R39180 DVDD.n9435 DVDD.n9434 0.019716
R39181 DVDD.n9434 DVDD.n9243 0.019716
R39182 DVDD.n9428 DVDD.n9427 0.019716
R39183 DVDD.n9427 DVDD.n9242 0.019716
R39184 DVDD.n9423 DVDD.n9422 0.019716
R39185 DVDD.n9422 DVDD.n9241 0.019716
R39186 DVDD.n9416 DVDD.n9415 0.019716
R39187 DVDD.n9415 DVDD.n9240 0.019716
R39188 DVDD.n9411 DVDD.n9410 0.019716
R39189 DVDD.n9410 DVDD.n9239 0.019716
R39190 DVDD.n9404 DVDD.n9403 0.019716
R39191 DVDD.n9403 DVDD.n9238 0.019716
R39192 DVDD.n9399 DVDD.n9398 0.019716
R39193 DVDD.n9398 DVDD.n9237 0.019716
R39194 DVDD.n9392 DVDD.n9391 0.019716
R39195 DVDD.n9391 DVDD.n9236 0.019716
R39196 DVDD.n9387 DVDD.n9386 0.019716
R39197 DVDD.n9386 DVDD.n9235 0.019716
R39198 DVDD.n9380 DVDD.n9379 0.019716
R39199 DVDD.n9379 DVDD.n9234 0.019716
R39200 DVDD.n9375 DVDD.n9374 0.019716
R39201 DVDD.n9374 DVDD.n9233 0.019716
R39202 DVDD.n9368 DVDD.n9367 0.019716
R39203 DVDD.n9367 DVDD.n9232 0.019716
R39204 DVDD.n9363 DVDD.n9362 0.019716
R39205 DVDD.n9362 DVDD.n9231 0.019716
R39206 DVDD.n9356 DVDD.n9355 0.019716
R39207 DVDD.n9355 DVDD.n9230 0.019716
R39208 DVDD.n9351 DVDD.n9350 0.019716
R39209 DVDD.n9350 DVDD.n9229 0.019716
R39210 DVDD.n9344 DVDD.n9343 0.019716
R39211 DVDD.n9343 DVDD.n9228 0.019716
R39212 DVDD.n9339 DVDD.n9338 0.019716
R39213 DVDD.n9338 DVDD.n9227 0.019716
R39214 DVDD.n9332 DVDD.n9331 0.019716
R39215 DVDD.n9331 DVDD.n9226 0.019716
R39216 DVDD.n9327 DVDD.n9326 0.019716
R39217 DVDD.n9326 DVDD.n9225 0.019716
R39218 DVDD.n9320 DVDD.n9319 0.019716
R39219 DVDD.n9319 DVDD.n9224 0.019716
R39220 DVDD.n9315 DVDD.n9314 0.019716
R39221 DVDD.n9314 DVDD.n9223 0.019716
R39222 DVDD.n14839 DVDD.n7731 0.019716
R39223 DVDD.n7837 DVDD.n7774 0.019716
R39224 DVDD.n7837 DVDD.n7729 0.019716
R39225 DVDD.n7846 DVDD.n7773 0.019716
R39226 DVDD.n7846 DVDD.n7728 0.019716
R39227 DVDD.n7834 DVDD.n7772 0.019716
R39228 DVDD.n7834 DVDD.n7727 0.019716
R39229 DVDD.n7855 DVDD.n7771 0.019716
R39230 DVDD.n7855 DVDD.n7726 0.019716
R39231 DVDD.n7831 DVDD.n7770 0.019716
R39232 DVDD.n7831 DVDD.n7725 0.019716
R39233 DVDD.n7864 DVDD.n7769 0.019716
R39234 DVDD.n7864 DVDD.n7724 0.019716
R39235 DVDD.n7828 DVDD.n7768 0.019716
R39236 DVDD.n7828 DVDD.n7723 0.019716
R39237 DVDD.n7873 DVDD.n7767 0.019716
R39238 DVDD.n7873 DVDD.n7722 0.019716
R39239 DVDD.n7825 DVDD.n7766 0.019716
R39240 DVDD.n7825 DVDD.n7721 0.019716
R39241 DVDD.n7882 DVDD.n7765 0.019716
R39242 DVDD.n7882 DVDD.n7720 0.019716
R39243 DVDD.n7822 DVDD.n7764 0.019716
R39244 DVDD.n7822 DVDD.n7719 0.019716
R39245 DVDD.n7891 DVDD.n7763 0.019716
R39246 DVDD.n7891 DVDD.n7718 0.019716
R39247 DVDD.n7819 DVDD.n7762 0.019716
R39248 DVDD.n7819 DVDD.n7717 0.019716
R39249 DVDD.n7900 DVDD.n7761 0.019716
R39250 DVDD.n7900 DVDD.n7716 0.019716
R39251 DVDD.n7816 DVDD.n7760 0.019716
R39252 DVDD.n7816 DVDD.n7715 0.019716
R39253 DVDD.n7909 DVDD.n7759 0.019716
R39254 DVDD.n7909 DVDD.n7714 0.019716
R39255 DVDD.n7813 DVDD.n7758 0.019716
R39256 DVDD.n7813 DVDD.n7713 0.019716
R39257 DVDD.n7918 DVDD.n7757 0.019716
R39258 DVDD.n7918 DVDD.n7712 0.019716
R39259 DVDD.n7810 DVDD.n7756 0.019716
R39260 DVDD.n7810 DVDD.n7711 0.019716
R39261 DVDD.n7927 DVDD.n7755 0.019716
R39262 DVDD.n7927 DVDD.n7710 0.019716
R39263 DVDD.n7807 DVDD.n7754 0.019716
R39264 DVDD.n7807 DVDD.n7709 0.019716
R39265 DVDD.n7936 DVDD.n7753 0.019716
R39266 DVDD.n7936 DVDD.n7708 0.019716
R39267 DVDD.n7804 DVDD.n7752 0.019716
R39268 DVDD.n7804 DVDD.n7707 0.019716
R39269 DVDD.n7945 DVDD.n7751 0.019716
R39270 DVDD.n7945 DVDD.n7706 0.019716
R39271 DVDD.n7801 DVDD.n7750 0.019716
R39272 DVDD.n7801 DVDD.n7705 0.019716
R39273 DVDD.n7954 DVDD.n7749 0.019716
R39274 DVDD.n7954 DVDD.n7704 0.019716
R39275 DVDD.n7798 DVDD.n7748 0.019716
R39276 DVDD.n7798 DVDD.n7703 0.019716
R39277 DVDD.n7963 DVDD.n7747 0.019716
R39278 DVDD.n7963 DVDD.n7702 0.019716
R39279 DVDD.n7795 DVDD.n7746 0.019716
R39280 DVDD.n7795 DVDD.n7701 0.019716
R39281 DVDD.n7972 DVDD.n7745 0.019716
R39282 DVDD.n7972 DVDD.n7700 0.019716
R39283 DVDD.n7792 DVDD.n7744 0.019716
R39284 DVDD.n7792 DVDD.n7699 0.019716
R39285 DVDD.n7981 DVDD.n7743 0.019716
R39286 DVDD.n7981 DVDD.n7698 0.019716
R39287 DVDD.n7789 DVDD.n7742 0.019716
R39288 DVDD.n7789 DVDD.n7697 0.019716
R39289 DVDD.n7990 DVDD.n7741 0.019716
R39290 DVDD.n7990 DVDD.n7696 0.019716
R39291 DVDD.n7786 DVDD.n7740 0.019716
R39292 DVDD.n7786 DVDD.n7695 0.019716
R39293 DVDD.n7999 DVDD.n7739 0.019716
R39294 DVDD.n7999 DVDD.n7694 0.019716
R39295 DVDD.n7783 DVDD.n7738 0.019716
R39296 DVDD.n7783 DVDD.n7693 0.019716
R39297 DVDD.n8008 DVDD.n7737 0.019716
R39298 DVDD.n8008 DVDD.n7692 0.019716
R39299 DVDD.n7780 DVDD.n7736 0.019716
R39300 DVDD.n7780 DVDD.n7691 0.019716
R39301 DVDD.n8017 DVDD.n7735 0.019716
R39302 DVDD.n8017 DVDD.n7690 0.019716
R39303 DVDD.n7777 DVDD.n7734 0.019716
R39304 DVDD.n7777 DVDD.n7689 0.019716
R39305 DVDD.n8131 DVDD.n8130 0.019716
R39306 DVDD.n14582 DVDD.n8085 0.019716
R39307 DVDD.n14583 DVDD.n14582 0.019716
R39308 DVDD.n14588 DVDD.n8084 0.019716
R39309 DVDD.n14588 DVDD.n14587 0.019716
R39310 DVDD.n14594 DVDD.n8083 0.019716
R39311 DVDD.n14595 DVDD.n14594 0.019716
R39312 DVDD.n14600 DVDD.n8082 0.019716
R39313 DVDD.n14600 DVDD.n14599 0.019716
R39314 DVDD.n14606 DVDD.n8081 0.019716
R39315 DVDD.n14607 DVDD.n14606 0.019716
R39316 DVDD.n14612 DVDD.n8080 0.019716
R39317 DVDD.n14612 DVDD.n14611 0.019716
R39318 DVDD.n14618 DVDD.n8079 0.019716
R39319 DVDD.n14619 DVDD.n14618 0.019716
R39320 DVDD.n14624 DVDD.n8078 0.019716
R39321 DVDD.n14624 DVDD.n14623 0.019716
R39322 DVDD.n14630 DVDD.n8077 0.019716
R39323 DVDD.n14631 DVDD.n14630 0.019716
R39324 DVDD.n14636 DVDD.n8076 0.019716
R39325 DVDD.n14636 DVDD.n14635 0.019716
R39326 DVDD.n14642 DVDD.n8075 0.019716
R39327 DVDD.n14643 DVDD.n14642 0.019716
R39328 DVDD.n14648 DVDD.n8074 0.019716
R39329 DVDD.n14648 DVDD.n14647 0.019716
R39330 DVDD.n14654 DVDD.n8073 0.019716
R39331 DVDD.n14655 DVDD.n14654 0.019716
R39332 DVDD.n14660 DVDD.n8072 0.019716
R39333 DVDD.n14660 DVDD.n14659 0.019716
R39334 DVDD.n14666 DVDD.n8071 0.019716
R39335 DVDD.n14667 DVDD.n14666 0.019716
R39336 DVDD.n14672 DVDD.n8070 0.019716
R39337 DVDD.n14672 DVDD.n14671 0.019716
R39338 DVDD.n14678 DVDD.n8069 0.019716
R39339 DVDD.n14679 DVDD.n14678 0.019716
R39340 DVDD.n14684 DVDD.n8068 0.019716
R39341 DVDD.n14684 DVDD.n14683 0.019716
R39342 DVDD.n14690 DVDD.n8067 0.019716
R39343 DVDD.n14691 DVDD.n14690 0.019716
R39344 DVDD.n14696 DVDD.n8066 0.019716
R39345 DVDD.n14696 DVDD.n14695 0.019716
R39346 DVDD.n14702 DVDD.n8065 0.019716
R39347 DVDD.n14703 DVDD.n14702 0.019716
R39348 DVDD.n14708 DVDD.n8064 0.019716
R39349 DVDD.n14708 DVDD.n14707 0.019716
R39350 DVDD.n14714 DVDD.n8063 0.019716
R39351 DVDD.n14715 DVDD.n14714 0.019716
R39352 DVDD.n14720 DVDD.n8062 0.019716
R39353 DVDD.n14720 DVDD.n14719 0.019716
R39354 DVDD.n14726 DVDD.n8061 0.019716
R39355 DVDD.n14727 DVDD.n14726 0.019716
R39356 DVDD.n14732 DVDD.n8060 0.019716
R39357 DVDD.n14732 DVDD.n14731 0.019716
R39358 DVDD.n14738 DVDD.n8059 0.019716
R39359 DVDD.n14739 DVDD.n14738 0.019716
R39360 DVDD.n14744 DVDD.n8058 0.019716
R39361 DVDD.n14744 DVDD.n14743 0.019716
R39362 DVDD.n14750 DVDD.n8057 0.019716
R39363 DVDD.n14751 DVDD.n14750 0.019716
R39364 DVDD.n14756 DVDD.n8056 0.019716
R39365 DVDD.n14756 DVDD.n14755 0.019716
R39366 DVDD.n14762 DVDD.n8055 0.019716
R39367 DVDD.n14763 DVDD.n14762 0.019716
R39368 DVDD.n14768 DVDD.n8054 0.019716
R39369 DVDD.n14768 DVDD.n14767 0.019716
R39370 DVDD.n14774 DVDD.n8053 0.019716
R39371 DVDD.n14775 DVDD.n14774 0.019716
R39372 DVDD.n14780 DVDD.n8052 0.019716
R39373 DVDD.n14780 DVDD.n14779 0.019716
R39374 DVDD.n14786 DVDD.n8051 0.019716
R39375 DVDD.n14787 DVDD.n14786 0.019716
R39376 DVDD.n14792 DVDD.n8050 0.019716
R39377 DVDD.n14792 DVDD.n14791 0.019716
R39378 DVDD.n14798 DVDD.n8049 0.019716
R39379 DVDD.n14799 DVDD.n14798 0.019716
R39380 DVDD.n14804 DVDD.n8048 0.019716
R39381 DVDD.n14804 DVDD.n14803 0.019716
R39382 DVDD.n14810 DVDD.n8047 0.019716
R39383 DVDD.n14811 DVDD.n14810 0.019716
R39384 DVDD.n14816 DVDD.n8046 0.019716
R39385 DVDD.n14816 DVDD.n14815 0.019716
R39386 DVDD.n14822 DVDD.n8045 0.019716
R39387 DVDD.n14823 DVDD.n14822 0.019716
R39388 DVDD.n8248 DVDD.n8247 0.019716
R39389 DVDD.n14316 DVDD.n8203 0.019716
R39390 DVDD.n14317 DVDD.n14316 0.019716
R39391 DVDD.n14322 DVDD.n8202 0.019716
R39392 DVDD.n14322 DVDD.n14321 0.019716
R39393 DVDD.n14328 DVDD.n8201 0.019716
R39394 DVDD.n14329 DVDD.n14328 0.019716
R39395 DVDD.n14334 DVDD.n8200 0.019716
R39396 DVDD.n14334 DVDD.n14333 0.019716
R39397 DVDD.n14340 DVDD.n8199 0.019716
R39398 DVDD.n14341 DVDD.n14340 0.019716
R39399 DVDD.n14346 DVDD.n8198 0.019716
R39400 DVDD.n14346 DVDD.n14345 0.019716
R39401 DVDD.n14352 DVDD.n8197 0.019716
R39402 DVDD.n14353 DVDD.n14352 0.019716
R39403 DVDD.n14358 DVDD.n8196 0.019716
R39404 DVDD.n14358 DVDD.n14357 0.019716
R39405 DVDD.n14364 DVDD.n8195 0.019716
R39406 DVDD.n14365 DVDD.n14364 0.019716
R39407 DVDD.n14370 DVDD.n8194 0.019716
R39408 DVDD.n14370 DVDD.n14369 0.019716
R39409 DVDD.n14376 DVDD.n8193 0.019716
R39410 DVDD.n14377 DVDD.n14376 0.019716
R39411 DVDD.n14382 DVDD.n8192 0.019716
R39412 DVDD.n14382 DVDD.n14381 0.019716
R39413 DVDD.n14388 DVDD.n8191 0.019716
R39414 DVDD.n14389 DVDD.n14388 0.019716
R39415 DVDD.n14394 DVDD.n8190 0.019716
R39416 DVDD.n14394 DVDD.n14393 0.019716
R39417 DVDD.n14400 DVDD.n8189 0.019716
R39418 DVDD.n14401 DVDD.n14400 0.019716
R39419 DVDD.n14406 DVDD.n8188 0.019716
R39420 DVDD.n14406 DVDD.n14405 0.019716
R39421 DVDD.n14412 DVDD.n8187 0.019716
R39422 DVDD.n14413 DVDD.n14412 0.019716
R39423 DVDD.n14418 DVDD.n8186 0.019716
R39424 DVDD.n14418 DVDD.n14417 0.019716
R39425 DVDD.n14424 DVDD.n8185 0.019716
R39426 DVDD.n14425 DVDD.n14424 0.019716
R39427 DVDD.n14430 DVDD.n8184 0.019716
R39428 DVDD.n14430 DVDD.n14429 0.019716
R39429 DVDD.n14436 DVDD.n8183 0.019716
R39430 DVDD.n14437 DVDD.n14436 0.019716
R39431 DVDD.n14442 DVDD.n8182 0.019716
R39432 DVDD.n14442 DVDD.n14441 0.019716
R39433 DVDD.n14448 DVDD.n8181 0.019716
R39434 DVDD.n14449 DVDD.n14448 0.019716
R39435 DVDD.n14454 DVDD.n8180 0.019716
R39436 DVDD.n14454 DVDD.n14453 0.019716
R39437 DVDD.n14460 DVDD.n8179 0.019716
R39438 DVDD.n14461 DVDD.n14460 0.019716
R39439 DVDD.n14466 DVDD.n8178 0.019716
R39440 DVDD.n14466 DVDD.n14465 0.019716
R39441 DVDD.n14472 DVDD.n8177 0.019716
R39442 DVDD.n14473 DVDD.n14472 0.019716
R39443 DVDD.n14478 DVDD.n8176 0.019716
R39444 DVDD.n14478 DVDD.n14477 0.019716
R39445 DVDD.n14484 DVDD.n8175 0.019716
R39446 DVDD.n14485 DVDD.n14484 0.019716
R39447 DVDD.n14490 DVDD.n8174 0.019716
R39448 DVDD.n14490 DVDD.n14489 0.019716
R39449 DVDD.n14496 DVDD.n8173 0.019716
R39450 DVDD.n14497 DVDD.n14496 0.019716
R39451 DVDD.n14502 DVDD.n8172 0.019716
R39452 DVDD.n14502 DVDD.n14501 0.019716
R39453 DVDD.n14508 DVDD.n8171 0.019716
R39454 DVDD.n14509 DVDD.n14508 0.019716
R39455 DVDD.n14514 DVDD.n8170 0.019716
R39456 DVDD.n14514 DVDD.n14513 0.019716
R39457 DVDD.n14520 DVDD.n8169 0.019716
R39458 DVDD.n14521 DVDD.n14520 0.019716
R39459 DVDD.n14526 DVDD.n8168 0.019716
R39460 DVDD.n14526 DVDD.n14525 0.019716
R39461 DVDD.n14532 DVDD.n8167 0.019716
R39462 DVDD.n14533 DVDD.n14532 0.019716
R39463 DVDD.n14538 DVDD.n8166 0.019716
R39464 DVDD.n14538 DVDD.n14537 0.019716
R39465 DVDD.n14544 DVDD.n8165 0.019716
R39466 DVDD.n14545 DVDD.n14544 0.019716
R39467 DVDD.n14550 DVDD.n8164 0.019716
R39468 DVDD.n14550 DVDD.n14549 0.019716
R39469 DVDD.n14556 DVDD.n8163 0.019716
R39470 DVDD.n14557 DVDD.n14556 0.019716
R39471 DVDD.n8351 DVDD.n8350 0.019716
R39472 DVDD.n8355 DVDD.n8352 0.019716
R39473 DVDD.n8355 DVDD.n8354 0.019716
R39474 DVDD.n8361 DVDD.n8343 0.019716
R39475 DVDD.n8362 DVDD.n8361 0.019716
R39476 DVDD.n8367 DVDD.n8364 0.019716
R39477 DVDD.n8367 DVDD.n8366 0.019716
R39478 DVDD.n8373 DVDD.n8339 0.019716
R39479 DVDD.n8374 DVDD.n8373 0.019716
R39480 DVDD.n8379 DVDD.n8376 0.019716
R39481 DVDD.n8379 DVDD.n8378 0.019716
R39482 DVDD.n8385 DVDD.n8335 0.019716
R39483 DVDD.n8386 DVDD.n8385 0.019716
R39484 DVDD.n8391 DVDD.n8388 0.019716
R39485 DVDD.n8391 DVDD.n8390 0.019716
R39486 DVDD.n8397 DVDD.n8331 0.019716
R39487 DVDD.n8398 DVDD.n8397 0.019716
R39488 DVDD.n8403 DVDD.n8400 0.019716
R39489 DVDD.n8403 DVDD.n8402 0.019716
R39490 DVDD.n8409 DVDD.n8327 0.019716
R39491 DVDD.n8410 DVDD.n8409 0.019716
R39492 DVDD.n8415 DVDD.n8412 0.019716
R39493 DVDD.n8415 DVDD.n8414 0.019716
R39494 DVDD.n8421 DVDD.n8323 0.019716
R39495 DVDD.n8422 DVDD.n8421 0.019716
R39496 DVDD.n8427 DVDD.n8424 0.019716
R39497 DVDD.n8427 DVDD.n8426 0.019716
R39498 DVDD.n8433 DVDD.n8319 0.019716
R39499 DVDD.n8434 DVDD.n8433 0.019716
R39500 DVDD.n8439 DVDD.n8436 0.019716
R39501 DVDD.n8439 DVDD.n8438 0.019716
R39502 DVDD.n8445 DVDD.n8315 0.019716
R39503 DVDD.n8446 DVDD.n8445 0.019716
R39504 DVDD.n8451 DVDD.n8448 0.019716
R39505 DVDD.n8451 DVDD.n8450 0.019716
R39506 DVDD.n8457 DVDD.n8311 0.019716
R39507 DVDD.n8458 DVDD.n8457 0.019716
R39508 DVDD.n8463 DVDD.n8460 0.019716
R39509 DVDD.n8463 DVDD.n8462 0.019716
R39510 DVDD.n8469 DVDD.n8307 0.019716
R39511 DVDD.n8470 DVDD.n8469 0.019716
R39512 DVDD.n8475 DVDD.n8472 0.019716
R39513 DVDD.n8475 DVDD.n8474 0.019716
R39514 DVDD.n8481 DVDD.n8303 0.019716
R39515 DVDD.n8482 DVDD.n8481 0.019716
R39516 DVDD.n8487 DVDD.n8484 0.019716
R39517 DVDD.n8487 DVDD.n8486 0.019716
R39518 DVDD.n8493 DVDD.n8299 0.019716
R39519 DVDD.n8494 DVDD.n8493 0.019716
R39520 DVDD.n8499 DVDD.n8496 0.019716
R39521 DVDD.n8499 DVDD.n8498 0.019716
R39522 DVDD.n8505 DVDD.n8295 0.019716
R39523 DVDD.n8506 DVDD.n8505 0.019716
R39524 DVDD.n8511 DVDD.n8508 0.019716
R39525 DVDD.n8511 DVDD.n8510 0.019716
R39526 DVDD.n8517 DVDD.n8291 0.019716
R39527 DVDD.n8518 DVDD.n8517 0.019716
R39528 DVDD.n8523 DVDD.n8520 0.019716
R39529 DVDD.n8523 DVDD.n8522 0.019716
R39530 DVDD.n8529 DVDD.n8287 0.019716
R39531 DVDD.n8530 DVDD.n8529 0.019716
R39532 DVDD.n8535 DVDD.n8532 0.019716
R39533 DVDD.n8535 DVDD.n8534 0.019716
R39534 DVDD.n8541 DVDD.n8283 0.019716
R39535 DVDD.n8542 DVDD.n8541 0.019716
R39536 DVDD.n8547 DVDD.n8544 0.019716
R39537 DVDD.n8547 DVDD.n8546 0.019716
R39538 DVDD.n8553 DVDD.n8279 0.019716
R39539 DVDD.n8554 DVDD.n8553 0.019716
R39540 DVDD.n8559 DVDD.n8556 0.019716
R39541 DVDD.n8559 DVDD.n8558 0.019716
R39542 DVDD.n8565 DVDD.n8275 0.019716
R39543 DVDD.n8566 DVDD.n8565 0.019716
R39544 DVDD.n8571 DVDD.n8568 0.019716
R39545 DVDD.n8571 DVDD.n8570 0.019716
R39546 DVDD.n8577 DVDD.n8271 0.019716
R39547 DVDD.n8578 DVDD.n8577 0.019716
R39548 DVDD.n8583 DVDD.n8580 0.019716
R39549 DVDD.n8583 DVDD.n8582 0.019716
R39550 DVDD.n8590 DVDD.n8267 0.019716
R39551 DVDD.n8591 DVDD.n8590 0.019716
R39552 DVDD.n8594 DVDD.n8593 0.019716
R39553 DVDD.n8595 DVDD.n8594 0.019716
R39554 DVDD.n8946 DVDD.n8945 0.019716
R39555 DVDD.n8944 DVDD.n8943 0.019716
R39556 DVDD.n8943 DVDD.n8617 0.019716
R39557 DVDD.n8937 DVDD.n8622 0.019716
R39558 DVDD.n8937 DVDD.n8936 0.019716
R39559 DVDD.n8934 DVDD.n8933 0.019716
R39560 DVDD.n8933 DVDD.n8623 0.019716
R39561 DVDD.n8927 DVDD.n8628 0.019716
R39562 DVDD.n8927 DVDD.n8926 0.019716
R39563 DVDD.n8924 DVDD.n8923 0.019716
R39564 DVDD.n8923 DVDD.n8629 0.019716
R39565 DVDD.n8917 DVDD.n8634 0.019716
R39566 DVDD.n8917 DVDD.n8916 0.019716
R39567 DVDD.n8914 DVDD.n8913 0.019716
R39568 DVDD.n8913 DVDD.n8635 0.019716
R39569 DVDD.n8907 DVDD.n8640 0.019716
R39570 DVDD.n8907 DVDD.n8906 0.019716
R39571 DVDD.n8904 DVDD.n8903 0.019716
R39572 DVDD.n8903 DVDD.n8641 0.019716
R39573 DVDD.n8897 DVDD.n8646 0.019716
R39574 DVDD.n8897 DVDD.n8896 0.019716
R39575 DVDD.n8894 DVDD.n8893 0.019716
R39576 DVDD.n8893 DVDD.n8647 0.019716
R39577 DVDD.n8887 DVDD.n8652 0.019716
R39578 DVDD.n8887 DVDD.n8886 0.019716
R39579 DVDD.n8884 DVDD.n8883 0.019716
R39580 DVDD.n8883 DVDD.n8653 0.019716
R39581 DVDD.n8877 DVDD.n8658 0.019716
R39582 DVDD.n8877 DVDD.n8876 0.019716
R39583 DVDD.n8874 DVDD.n8873 0.019716
R39584 DVDD.n8873 DVDD.n8659 0.019716
R39585 DVDD.n8867 DVDD.n8664 0.019716
R39586 DVDD.n8867 DVDD.n8866 0.019716
R39587 DVDD.n8864 DVDD.n8863 0.019716
R39588 DVDD.n8863 DVDD.n8665 0.019716
R39589 DVDD.n8857 DVDD.n8670 0.019716
R39590 DVDD.n8857 DVDD.n8856 0.019716
R39591 DVDD.n8854 DVDD.n8853 0.019716
R39592 DVDD.n8853 DVDD.n8671 0.019716
R39593 DVDD.n8847 DVDD.n8676 0.019716
R39594 DVDD.n8847 DVDD.n8846 0.019716
R39595 DVDD.n8844 DVDD.n8843 0.019716
R39596 DVDD.n8843 DVDD.n8677 0.019716
R39597 DVDD.n8837 DVDD.n8682 0.019716
R39598 DVDD.n8837 DVDD.n8836 0.019716
R39599 DVDD.n8834 DVDD.n8833 0.019716
R39600 DVDD.n8833 DVDD.n8683 0.019716
R39601 DVDD.n8827 DVDD.n8688 0.019716
R39602 DVDD.n8827 DVDD.n8826 0.019716
R39603 DVDD.n8824 DVDD.n8823 0.019716
R39604 DVDD.n8823 DVDD.n8689 0.019716
R39605 DVDD.n8817 DVDD.n8694 0.019716
R39606 DVDD.n8817 DVDD.n8816 0.019716
R39607 DVDD.n8814 DVDD.n8813 0.019716
R39608 DVDD.n8813 DVDD.n8695 0.019716
R39609 DVDD.n8807 DVDD.n8700 0.019716
R39610 DVDD.n8807 DVDD.n8806 0.019716
R39611 DVDD.n8804 DVDD.n8803 0.019716
R39612 DVDD.n8803 DVDD.n8701 0.019716
R39613 DVDD.n8797 DVDD.n8706 0.019716
R39614 DVDD.n8797 DVDD.n8796 0.019716
R39615 DVDD.n8794 DVDD.n8793 0.019716
R39616 DVDD.n8793 DVDD.n8707 0.019716
R39617 DVDD.n8787 DVDD.n8712 0.019716
R39618 DVDD.n8787 DVDD.n8786 0.019716
R39619 DVDD.n8784 DVDD.n8783 0.019716
R39620 DVDD.n8783 DVDD.n8713 0.019716
R39621 DVDD.n8777 DVDD.n8718 0.019716
R39622 DVDD.n8777 DVDD.n8776 0.019716
R39623 DVDD.n8774 DVDD.n8773 0.019716
R39624 DVDD.n8773 DVDD.n8719 0.019716
R39625 DVDD.n8767 DVDD.n8724 0.019716
R39626 DVDD.n8767 DVDD.n8766 0.019716
R39627 DVDD.n8764 DVDD.n8763 0.019716
R39628 DVDD.n8763 DVDD.n8725 0.019716
R39629 DVDD.n8757 DVDD.n8730 0.019716
R39630 DVDD.n8757 DVDD.n8756 0.019716
R39631 DVDD.n8754 DVDD.n8753 0.019716
R39632 DVDD.n8753 DVDD.n8731 0.019716
R39633 DVDD.n8747 DVDD.n8736 0.019716
R39634 DVDD.n8747 DVDD.n8746 0.019716
R39635 DVDD.n8744 DVDD.n8743 0.019716
R39636 DVDD.n8743 DVDD.n8737 0.019716
R39637 DVDD.n14283 DVDD.n10284 0.019716
R39638 DVDD.n10390 DVDD.n10327 0.019716
R39639 DVDD.n10390 DVDD.n10282 0.019716
R39640 DVDD.n10399 DVDD.n10326 0.019716
R39641 DVDD.n10399 DVDD.n10281 0.019716
R39642 DVDD.n10387 DVDD.n10325 0.019716
R39643 DVDD.n10387 DVDD.n10280 0.019716
R39644 DVDD.n10408 DVDD.n10324 0.019716
R39645 DVDD.n10408 DVDD.n10279 0.019716
R39646 DVDD.n10384 DVDD.n10323 0.019716
R39647 DVDD.n10384 DVDD.n10278 0.019716
R39648 DVDD.n10417 DVDD.n10322 0.019716
R39649 DVDD.n10417 DVDD.n10277 0.019716
R39650 DVDD.n10381 DVDD.n10321 0.019716
R39651 DVDD.n10381 DVDD.n10276 0.019716
R39652 DVDD.n10426 DVDD.n10320 0.019716
R39653 DVDD.n10426 DVDD.n10275 0.019716
R39654 DVDD.n10378 DVDD.n10319 0.019716
R39655 DVDD.n10378 DVDD.n10274 0.019716
R39656 DVDD.n10435 DVDD.n10318 0.019716
R39657 DVDD.n10435 DVDD.n10273 0.019716
R39658 DVDD.n10375 DVDD.n10317 0.019716
R39659 DVDD.n10375 DVDD.n10272 0.019716
R39660 DVDD.n10444 DVDD.n10316 0.019716
R39661 DVDD.n10444 DVDD.n10271 0.019716
R39662 DVDD.n10372 DVDD.n10315 0.019716
R39663 DVDD.n10372 DVDD.n10270 0.019716
R39664 DVDD.n10453 DVDD.n10314 0.019716
R39665 DVDD.n10453 DVDD.n10269 0.019716
R39666 DVDD.n10369 DVDD.n10313 0.019716
R39667 DVDD.n10369 DVDD.n10268 0.019716
R39668 DVDD.n10462 DVDD.n10312 0.019716
R39669 DVDD.n10462 DVDD.n10267 0.019716
R39670 DVDD.n10366 DVDD.n10311 0.019716
R39671 DVDD.n10366 DVDD.n10266 0.019716
R39672 DVDD.n10471 DVDD.n10310 0.019716
R39673 DVDD.n10471 DVDD.n10265 0.019716
R39674 DVDD.n10363 DVDD.n10309 0.019716
R39675 DVDD.n10363 DVDD.n10264 0.019716
R39676 DVDD.n10480 DVDD.n10308 0.019716
R39677 DVDD.n10480 DVDD.n10263 0.019716
R39678 DVDD.n10360 DVDD.n10307 0.019716
R39679 DVDD.n10360 DVDD.n10262 0.019716
R39680 DVDD.n10489 DVDD.n10306 0.019716
R39681 DVDD.n10489 DVDD.n10261 0.019716
R39682 DVDD.n10357 DVDD.n10305 0.019716
R39683 DVDD.n10357 DVDD.n10260 0.019716
R39684 DVDD.n10498 DVDD.n10304 0.019716
R39685 DVDD.n10498 DVDD.n10259 0.019716
R39686 DVDD.n10354 DVDD.n10303 0.019716
R39687 DVDD.n10354 DVDD.n10258 0.019716
R39688 DVDD.n10507 DVDD.n10302 0.019716
R39689 DVDD.n10507 DVDD.n10257 0.019716
R39690 DVDD.n10351 DVDD.n10301 0.019716
R39691 DVDD.n10351 DVDD.n10256 0.019716
R39692 DVDD.n10516 DVDD.n10300 0.019716
R39693 DVDD.n10516 DVDD.n10255 0.019716
R39694 DVDD.n10348 DVDD.n10299 0.019716
R39695 DVDD.n10348 DVDD.n10254 0.019716
R39696 DVDD.n10525 DVDD.n10298 0.019716
R39697 DVDD.n10525 DVDD.n10253 0.019716
R39698 DVDD.n10345 DVDD.n10297 0.019716
R39699 DVDD.n10345 DVDD.n10252 0.019716
R39700 DVDD.n10534 DVDD.n10296 0.019716
R39701 DVDD.n10534 DVDD.n10251 0.019716
R39702 DVDD.n10342 DVDD.n10295 0.019716
R39703 DVDD.n10342 DVDD.n10250 0.019716
R39704 DVDD.n10543 DVDD.n10294 0.019716
R39705 DVDD.n10543 DVDD.n10249 0.019716
R39706 DVDD.n10339 DVDD.n10293 0.019716
R39707 DVDD.n10339 DVDD.n10248 0.019716
R39708 DVDD.n10552 DVDD.n10292 0.019716
R39709 DVDD.n10552 DVDD.n10247 0.019716
R39710 DVDD.n10336 DVDD.n10291 0.019716
R39711 DVDD.n10336 DVDD.n10246 0.019716
R39712 DVDD.n10561 DVDD.n10290 0.019716
R39713 DVDD.n10561 DVDD.n10245 0.019716
R39714 DVDD.n10333 DVDD.n10289 0.019716
R39715 DVDD.n10333 DVDD.n10244 0.019716
R39716 DVDD.n10570 DVDD.n10288 0.019716
R39717 DVDD.n10570 DVDD.n10243 0.019716
R39718 DVDD.n10330 DVDD.n10287 0.019716
R39719 DVDD.n10330 DVDD.n10242 0.019716
R39720 DVDD.n10684 DVDD.n10683 0.019716
R39721 DVDD.n14026 DVDD.n10638 0.019716
R39722 DVDD.n14027 DVDD.n14026 0.019716
R39723 DVDD.n14032 DVDD.n10637 0.019716
R39724 DVDD.n14032 DVDD.n14031 0.019716
R39725 DVDD.n14038 DVDD.n10636 0.019716
R39726 DVDD.n14039 DVDD.n14038 0.019716
R39727 DVDD.n14044 DVDD.n10635 0.019716
R39728 DVDD.n14044 DVDD.n14043 0.019716
R39729 DVDD.n14050 DVDD.n10634 0.019716
R39730 DVDD.n14051 DVDD.n14050 0.019716
R39731 DVDD.n14056 DVDD.n10633 0.019716
R39732 DVDD.n14056 DVDD.n14055 0.019716
R39733 DVDD.n14062 DVDD.n10632 0.019716
R39734 DVDD.n14063 DVDD.n14062 0.019716
R39735 DVDD.n14068 DVDD.n10631 0.019716
R39736 DVDD.n14068 DVDD.n14067 0.019716
R39737 DVDD.n14074 DVDD.n10630 0.019716
R39738 DVDD.n14075 DVDD.n14074 0.019716
R39739 DVDD.n14080 DVDD.n10629 0.019716
R39740 DVDD.n14080 DVDD.n14079 0.019716
R39741 DVDD.n14086 DVDD.n10628 0.019716
R39742 DVDD.n14087 DVDD.n14086 0.019716
R39743 DVDD.n14092 DVDD.n10627 0.019716
R39744 DVDD.n14092 DVDD.n14091 0.019716
R39745 DVDD.n14098 DVDD.n10626 0.019716
R39746 DVDD.n14099 DVDD.n14098 0.019716
R39747 DVDD.n14104 DVDD.n10625 0.019716
R39748 DVDD.n14104 DVDD.n14103 0.019716
R39749 DVDD.n14110 DVDD.n10624 0.019716
R39750 DVDD.n14111 DVDD.n14110 0.019716
R39751 DVDD.n14116 DVDD.n10623 0.019716
R39752 DVDD.n14116 DVDD.n14115 0.019716
R39753 DVDD.n14122 DVDD.n10622 0.019716
R39754 DVDD.n14123 DVDD.n14122 0.019716
R39755 DVDD.n14128 DVDD.n10621 0.019716
R39756 DVDD.n14128 DVDD.n14127 0.019716
R39757 DVDD.n14134 DVDD.n10620 0.019716
R39758 DVDD.n14135 DVDD.n14134 0.019716
R39759 DVDD.n14140 DVDD.n10619 0.019716
R39760 DVDD.n14140 DVDD.n14139 0.019716
R39761 DVDD.n14146 DVDD.n10618 0.019716
R39762 DVDD.n14147 DVDD.n14146 0.019716
R39763 DVDD.n14152 DVDD.n10617 0.019716
R39764 DVDD.n14152 DVDD.n14151 0.019716
R39765 DVDD.n14158 DVDD.n10616 0.019716
R39766 DVDD.n14159 DVDD.n14158 0.019716
R39767 DVDD.n14164 DVDD.n10615 0.019716
R39768 DVDD.n14164 DVDD.n14163 0.019716
R39769 DVDD.n14170 DVDD.n10614 0.019716
R39770 DVDD.n14171 DVDD.n14170 0.019716
R39771 DVDD.n14176 DVDD.n10613 0.019716
R39772 DVDD.n14176 DVDD.n14175 0.019716
R39773 DVDD.n14182 DVDD.n10612 0.019716
R39774 DVDD.n14183 DVDD.n14182 0.019716
R39775 DVDD.n14188 DVDD.n10611 0.019716
R39776 DVDD.n14188 DVDD.n14187 0.019716
R39777 DVDD.n14194 DVDD.n10610 0.019716
R39778 DVDD.n14195 DVDD.n14194 0.019716
R39779 DVDD.n14200 DVDD.n10609 0.019716
R39780 DVDD.n14200 DVDD.n14199 0.019716
R39781 DVDD.n14206 DVDD.n10608 0.019716
R39782 DVDD.n14207 DVDD.n14206 0.019716
R39783 DVDD.n14212 DVDD.n10607 0.019716
R39784 DVDD.n14212 DVDD.n14211 0.019716
R39785 DVDD.n14218 DVDD.n10606 0.019716
R39786 DVDD.n14219 DVDD.n14218 0.019716
R39787 DVDD.n14224 DVDD.n10605 0.019716
R39788 DVDD.n14224 DVDD.n14223 0.019716
R39789 DVDD.n14230 DVDD.n10604 0.019716
R39790 DVDD.n14231 DVDD.n14230 0.019716
R39791 DVDD.n14236 DVDD.n10603 0.019716
R39792 DVDD.n14236 DVDD.n14235 0.019716
R39793 DVDD.n14242 DVDD.n10602 0.019716
R39794 DVDD.n14243 DVDD.n14242 0.019716
R39795 DVDD.n14248 DVDD.n10601 0.019716
R39796 DVDD.n14248 DVDD.n14247 0.019716
R39797 DVDD.n14254 DVDD.n10600 0.019716
R39798 DVDD.n14255 DVDD.n14254 0.019716
R39799 DVDD.n14260 DVDD.n10599 0.019716
R39800 DVDD.n14260 DVDD.n14259 0.019716
R39801 DVDD.n14266 DVDD.n10598 0.019716
R39802 DVDD.n14267 DVDD.n14266 0.019716
R39803 DVDD.n10803 DVDD.n10802 0.019716
R39804 DVDD.n10807 DVDD.n10804 0.019716
R39805 DVDD.n10807 DVDD.n10806 0.019716
R39806 DVDD.n10813 DVDD.n10795 0.019716
R39807 DVDD.n10814 DVDD.n10813 0.019716
R39808 DVDD.n10819 DVDD.n10816 0.019716
R39809 DVDD.n10819 DVDD.n10818 0.019716
R39810 DVDD.n10825 DVDD.n10791 0.019716
R39811 DVDD.n10826 DVDD.n10825 0.019716
R39812 DVDD.n10831 DVDD.n10828 0.019716
R39813 DVDD.n10831 DVDD.n10830 0.019716
R39814 DVDD.n10837 DVDD.n10787 0.019716
R39815 DVDD.n10838 DVDD.n10837 0.019716
R39816 DVDD.n10843 DVDD.n10840 0.019716
R39817 DVDD.n10843 DVDD.n10842 0.019716
R39818 DVDD.n10849 DVDD.n10783 0.019716
R39819 DVDD.n10850 DVDD.n10849 0.019716
R39820 DVDD.n10855 DVDD.n10852 0.019716
R39821 DVDD.n10855 DVDD.n10854 0.019716
R39822 DVDD.n10861 DVDD.n10779 0.019716
R39823 DVDD.n10862 DVDD.n10861 0.019716
R39824 DVDD.n10867 DVDD.n10864 0.019716
R39825 DVDD.n10867 DVDD.n10866 0.019716
R39826 DVDD.n10873 DVDD.n10775 0.019716
R39827 DVDD.n10874 DVDD.n10873 0.019716
R39828 DVDD.n10879 DVDD.n10876 0.019716
R39829 DVDD.n10879 DVDD.n10878 0.019716
R39830 DVDD.n10885 DVDD.n10771 0.019716
R39831 DVDD.n10886 DVDD.n10885 0.019716
R39832 DVDD.n10891 DVDD.n10888 0.019716
R39833 DVDD.n10891 DVDD.n10890 0.019716
R39834 DVDD.n10897 DVDD.n10767 0.019716
R39835 DVDD.n10898 DVDD.n10897 0.019716
R39836 DVDD.n10903 DVDD.n10900 0.019716
R39837 DVDD.n10903 DVDD.n10902 0.019716
R39838 DVDD.n10909 DVDD.n10763 0.019716
R39839 DVDD.n10910 DVDD.n10909 0.019716
R39840 DVDD.n10915 DVDD.n10912 0.019716
R39841 DVDD.n10915 DVDD.n10914 0.019716
R39842 DVDD.n10921 DVDD.n10759 0.019716
R39843 DVDD.n10922 DVDD.n10921 0.019716
R39844 DVDD.n10927 DVDD.n10924 0.019716
R39845 DVDD.n10927 DVDD.n10926 0.019716
R39846 DVDD.n10933 DVDD.n10755 0.019716
R39847 DVDD.n10934 DVDD.n10933 0.019716
R39848 DVDD.n10939 DVDD.n10936 0.019716
R39849 DVDD.n10939 DVDD.n10938 0.019716
R39850 DVDD.n10945 DVDD.n10751 0.019716
R39851 DVDD.n10946 DVDD.n10945 0.019716
R39852 DVDD.n10951 DVDD.n10948 0.019716
R39853 DVDD.n10951 DVDD.n10950 0.019716
R39854 DVDD.n10957 DVDD.n10747 0.019716
R39855 DVDD.n10958 DVDD.n10957 0.019716
R39856 DVDD.n10963 DVDD.n10960 0.019716
R39857 DVDD.n10963 DVDD.n10962 0.019716
R39858 DVDD.n10969 DVDD.n10743 0.019716
R39859 DVDD.n10970 DVDD.n10969 0.019716
R39860 DVDD.n10975 DVDD.n10972 0.019716
R39861 DVDD.n10975 DVDD.n10974 0.019716
R39862 DVDD.n10981 DVDD.n10739 0.019716
R39863 DVDD.n10982 DVDD.n10981 0.019716
R39864 DVDD.n10987 DVDD.n10984 0.019716
R39865 DVDD.n10987 DVDD.n10986 0.019716
R39866 DVDD.n10993 DVDD.n10735 0.019716
R39867 DVDD.n10994 DVDD.n10993 0.019716
R39868 DVDD.n10999 DVDD.n10996 0.019716
R39869 DVDD.n10999 DVDD.n10998 0.019716
R39870 DVDD.n11005 DVDD.n10731 0.019716
R39871 DVDD.n11006 DVDD.n11005 0.019716
R39872 DVDD.n11011 DVDD.n11008 0.019716
R39873 DVDD.n11011 DVDD.n11010 0.019716
R39874 DVDD.n11017 DVDD.n10727 0.019716
R39875 DVDD.n11018 DVDD.n11017 0.019716
R39876 DVDD.n11023 DVDD.n11020 0.019716
R39877 DVDD.n11023 DVDD.n11022 0.019716
R39878 DVDD.n11029 DVDD.n10723 0.019716
R39879 DVDD.n11030 DVDD.n11029 0.019716
R39880 DVDD.n11035 DVDD.n11032 0.019716
R39881 DVDD.n11035 DVDD.n11034 0.019716
R39882 DVDD.n11042 DVDD.n10719 0.019716
R39883 DVDD.n11043 DVDD.n11042 0.019716
R39884 DVDD.n11046 DVDD.n11045 0.019716
R39885 DVDD.n11047 DVDD.n11046 0.019716
R39886 DVDD.n14002 DVDD.n11104 0.019716
R39887 DVDD.n11210 DVDD.n11148 0.019716
R39888 DVDD.n11210 DVDD.n11102 0.019716
R39889 DVDD.n13820 DVDD.n11147 0.019716
R39890 DVDD.n13820 DVDD.n11101 0.019716
R39891 DVDD.n11207 DVDD.n11146 0.019716
R39892 DVDD.n11207 DVDD.n11100 0.019716
R39893 DVDD.n13829 DVDD.n11145 0.019716
R39894 DVDD.n13829 DVDD.n11099 0.019716
R39895 DVDD.n11204 DVDD.n11144 0.019716
R39896 DVDD.n11204 DVDD.n11098 0.019716
R39897 DVDD.n13838 DVDD.n11143 0.019716
R39898 DVDD.n13838 DVDD.n11097 0.019716
R39899 DVDD.n11201 DVDD.n11142 0.019716
R39900 DVDD.n11201 DVDD.n11096 0.019716
R39901 DVDD.n13847 DVDD.n11141 0.019716
R39902 DVDD.n13847 DVDD.n11095 0.019716
R39903 DVDD.n11198 DVDD.n11140 0.019716
R39904 DVDD.n11198 DVDD.n11094 0.019716
R39905 DVDD.n13856 DVDD.n11139 0.019716
R39906 DVDD.n13856 DVDD.n11093 0.019716
R39907 DVDD.n11195 DVDD.n11138 0.019716
R39908 DVDD.n11195 DVDD.n11092 0.019716
R39909 DVDD.n13865 DVDD.n11137 0.019716
R39910 DVDD.n13865 DVDD.n11091 0.019716
R39911 DVDD.n11192 DVDD.n11136 0.019716
R39912 DVDD.n11192 DVDD.n11090 0.019716
R39913 DVDD.n13874 DVDD.n11135 0.019716
R39914 DVDD.n13874 DVDD.n11089 0.019716
R39915 DVDD.n11189 DVDD.n11134 0.019716
R39916 DVDD.n11189 DVDD.n11088 0.019716
R39917 DVDD.n13883 DVDD.n11133 0.019716
R39918 DVDD.n13883 DVDD.n11087 0.019716
R39919 DVDD.n11186 DVDD.n11132 0.019716
R39920 DVDD.n11186 DVDD.n11086 0.019716
R39921 DVDD.n13892 DVDD.n11131 0.019716
R39922 DVDD.n13892 DVDD.n11085 0.019716
R39923 DVDD.n11183 DVDD.n11130 0.019716
R39924 DVDD.n11183 DVDD.n11084 0.019716
R39925 DVDD.n13901 DVDD.n11129 0.019716
R39926 DVDD.n13901 DVDD.n11083 0.019716
R39927 DVDD.n11180 DVDD.n11128 0.019716
R39928 DVDD.n11180 DVDD.n11082 0.019716
R39929 DVDD.n13910 DVDD.n11127 0.019716
R39930 DVDD.n13910 DVDD.n11081 0.019716
R39931 DVDD.n11177 DVDD.n11126 0.019716
R39932 DVDD.n11177 DVDD.n11080 0.019716
R39933 DVDD.n13919 DVDD.n11125 0.019716
R39934 DVDD.n13919 DVDD.n11079 0.019716
R39935 DVDD.n11174 DVDD.n11124 0.019716
R39936 DVDD.n11174 DVDD.n11078 0.019716
R39937 DVDD.n13928 DVDD.n11123 0.019716
R39938 DVDD.n13928 DVDD.n11077 0.019716
R39939 DVDD.n11171 DVDD.n11122 0.019716
R39940 DVDD.n11171 DVDD.n11076 0.019716
R39941 DVDD.n13937 DVDD.n11121 0.019716
R39942 DVDD.n13937 DVDD.n11075 0.019716
R39943 DVDD.n11168 DVDD.n11120 0.019716
R39944 DVDD.n11168 DVDD.n11074 0.019716
R39945 DVDD.n13946 DVDD.n11119 0.019716
R39946 DVDD.n13946 DVDD.n11073 0.019716
R39947 DVDD.n11165 DVDD.n11118 0.019716
R39948 DVDD.n11165 DVDD.n11072 0.019716
R39949 DVDD.n13955 DVDD.n11117 0.019716
R39950 DVDD.n13955 DVDD.n11071 0.019716
R39951 DVDD.n11162 DVDD.n11116 0.019716
R39952 DVDD.n11162 DVDD.n11070 0.019716
R39953 DVDD.n13964 DVDD.n11115 0.019716
R39954 DVDD.n13964 DVDD.n11069 0.019716
R39955 DVDD.n11159 DVDD.n11114 0.019716
R39956 DVDD.n11159 DVDD.n11068 0.019716
R39957 DVDD.n13973 DVDD.n11113 0.019716
R39958 DVDD.n13973 DVDD.n11067 0.019716
R39959 DVDD.n11156 DVDD.n11112 0.019716
R39960 DVDD.n11156 DVDD.n11066 0.019716
R39961 DVDD.n13982 DVDD.n11111 0.019716
R39962 DVDD.n13982 DVDD.n11065 0.019716
R39963 DVDD.n11153 DVDD.n11110 0.019716
R39964 DVDD.n11153 DVDD.n11064 0.019716
R39965 DVDD.n13991 DVDD.n11109 0.019716
R39966 DVDD.n13991 DVDD.n11063 0.019716
R39967 DVDD.n11150 DVDD.n11108 0.019716
R39968 DVDD.n11150 DVDD.n11062 0.019716
R39969 DVDD.n11322 DVDD.n11321 0.019716
R39970 DVDD.n11327 DVDD.n11274 0.019716
R39971 DVDD.n11328 DVDD.n11327 0.019716
R39972 DVDD.n11333 DVDD.n11273 0.019716
R39973 DVDD.n11333 DVDD.n11332 0.019716
R39974 DVDD.n11339 DVDD.n11272 0.019716
R39975 DVDD.n11340 DVDD.n11339 0.019716
R39976 DVDD.n11345 DVDD.n11271 0.019716
R39977 DVDD.n11345 DVDD.n11344 0.019716
R39978 DVDD.n11351 DVDD.n11270 0.019716
R39979 DVDD.n11352 DVDD.n11351 0.019716
R39980 DVDD.n11357 DVDD.n11269 0.019716
R39981 DVDD.n11357 DVDD.n11356 0.019716
R39982 DVDD.n11363 DVDD.n11268 0.019716
R39983 DVDD.n11364 DVDD.n11363 0.019716
R39984 DVDD.n11369 DVDD.n11267 0.019716
R39985 DVDD.n11369 DVDD.n11368 0.019716
R39986 DVDD.n11375 DVDD.n11266 0.019716
R39987 DVDD.n11376 DVDD.n11375 0.019716
R39988 DVDD.n11381 DVDD.n11265 0.019716
R39989 DVDD.n11381 DVDD.n11380 0.019716
R39990 DVDD.n11387 DVDD.n11264 0.019716
R39991 DVDD.n11388 DVDD.n11387 0.019716
R39992 DVDD.n11393 DVDD.n11263 0.019716
R39993 DVDD.n11393 DVDD.n11392 0.019716
R39994 DVDD.n11399 DVDD.n11262 0.019716
R39995 DVDD.n11400 DVDD.n11399 0.019716
R39996 DVDD.n11405 DVDD.n11261 0.019716
R39997 DVDD.n11405 DVDD.n11404 0.019716
R39998 DVDD.n11411 DVDD.n11260 0.019716
R39999 DVDD.n11412 DVDD.n11411 0.019716
R40000 DVDD.n11417 DVDD.n11259 0.019716
R40001 DVDD.n11417 DVDD.n11416 0.019716
R40002 DVDD.n11423 DVDD.n11258 0.019716
R40003 DVDD.n11424 DVDD.n11423 0.019716
R40004 DVDD.n11429 DVDD.n11257 0.019716
R40005 DVDD.n11429 DVDD.n11428 0.019716
R40006 DVDD.n11435 DVDD.n11256 0.019716
R40007 DVDD.n11436 DVDD.n11435 0.019716
R40008 DVDD.n11441 DVDD.n11255 0.019716
R40009 DVDD.n11441 DVDD.n11440 0.019716
R40010 DVDD.n11447 DVDD.n11254 0.019716
R40011 DVDD.n11448 DVDD.n11447 0.019716
R40012 DVDD.n11453 DVDD.n11253 0.019716
R40013 DVDD.n11453 DVDD.n11452 0.019716
R40014 DVDD.n11459 DVDD.n11252 0.019716
R40015 DVDD.n11460 DVDD.n11459 0.019716
R40016 DVDD.n11465 DVDD.n11251 0.019716
R40017 DVDD.n11465 DVDD.n11464 0.019716
R40018 DVDD.n11471 DVDD.n11250 0.019716
R40019 DVDD.n11472 DVDD.n11471 0.019716
R40020 DVDD.n11477 DVDD.n11249 0.019716
R40021 DVDD.n11477 DVDD.n11476 0.019716
R40022 DVDD.n11483 DVDD.n11248 0.019716
R40023 DVDD.n11484 DVDD.n11483 0.019716
R40024 DVDD.n11489 DVDD.n11247 0.019716
R40025 DVDD.n11489 DVDD.n11488 0.019716
R40026 DVDD.n11495 DVDD.n11246 0.019716
R40027 DVDD.n11496 DVDD.n11495 0.019716
R40028 DVDD.n11501 DVDD.n11245 0.019716
R40029 DVDD.n11501 DVDD.n11500 0.019716
R40030 DVDD.n11507 DVDD.n11244 0.019716
R40031 DVDD.n11508 DVDD.n11507 0.019716
R40032 DVDD.n11513 DVDD.n11243 0.019716
R40033 DVDD.n11513 DVDD.n11512 0.019716
R40034 DVDD.n11519 DVDD.n11242 0.019716
R40035 DVDD.n11520 DVDD.n11519 0.019716
R40036 DVDD.n11525 DVDD.n11241 0.019716
R40037 DVDD.n11525 DVDD.n11524 0.019716
R40038 DVDD.n11531 DVDD.n11240 0.019716
R40039 DVDD.n11532 DVDD.n11531 0.019716
R40040 DVDD.n11537 DVDD.n11239 0.019716
R40041 DVDD.n11537 DVDD.n11536 0.019716
R40042 DVDD.n11543 DVDD.n11238 0.019716
R40043 DVDD.n11544 DVDD.n11543 0.019716
R40044 DVDD.n11549 DVDD.n11237 0.019716
R40045 DVDD.n11549 DVDD.n11548 0.019716
R40046 DVDD.n11555 DVDD.n11236 0.019716
R40047 DVDD.n11556 DVDD.n11555 0.019716
R40048 DVDD.n11561 DVDD.n11235 0.019716
R40049 DVDD.n11561 DVDD.n11560 0.019716
R40050 DVDD.n13796 DVDD.n11234 0.019716
R40051 DVDD.n13797 DVDD.n13796 0.019716
R40052 DVDD.n11676 DVDD.n11675 0.019716
R40053 DVDD.n11681 DVDD.n11629 0.019716
R40054 DVDD.n11682 DVDD.n11681 0.019716
R40055 DVDD.n11687 DVDD.n11628 0.019716
R40056 DVDD.n11687 DVDD.n11686 0.019716
R40057 DVDD.n11693 DVDD.n11627 0.019716
R40058 DVDD.n11694 DVDD.n11693 0.019716
R40059 DVDD.n11699 DVDD.n11626 0.019716
R40060 DVDD.n11699 DVDD.n11698 0.019716
R40061 DVDD.n11705 DVDD.n11625 0.019716
R40062 DVDD.n11706 DVDD.n11705 0.019716
R40063 DVDD.n11711 DVDD.n11624 0.019716
R40064 DVDD.n11711 DVDD.n11710 0.019716
R40065 DVDD.n11717 DVDD.n11623 0.019716
R40066 DVDD.n11718 DVDD.n11717 0.019716
R40067 DVDD.n11723 DVDD.n11622 0.019716
R40068 DVDD.n11723 DVDD.n11722 0.019716
R40069 DVDD.n11729 DVDD.n11621 0.019716
R40070 DVDD.n11730 DVDD.n11729 0.019716
R40071 DVDD.n11735 DVDD.n11620 0.019716
R40072 DVDD.n11735 DVDD.n11734 0.019716
R40073 DVDD.n11741 DVDD.n11619 0.019716
R40074 DVDD.n11742 DVDD.n11741 0.019716
R40075 DVDD.n11747 DVDD.n11618 0.019716
R40076 DVDD.n11747 DVDD.n11746 0.019716
R40077 DVDD.n11753 DVDD.n11617 0.019716
R40078 DVDD.n11754 DVDD.n11753 0.019716
R40079 DVDD.n11759 DVDD.n11616 0.019716
R40080 DVDD.n11759 DVDD.n11758 0.019716
R40081 DVDD.n11765 DVDD.n11615 0.019716
R40082 DVDD.n11766 DVDD.n11765 0.019716
R40083 DVDD.n11771 DVDD.n11614 0.019716
R40084 DVDD.n11771 DVDD.n11770 0.019716
R40085 DVDD.n11777 DVDD.n11613 0.019716
R40086 DVDD.n11778 DVDD.n11777 0.019716
R40087 DVDD.n11783 DVDD.n11612 0.019716
R40088 DVDD.n11783 DVDD.n11782 0.019716
R40089 DVDD.n11789 DVDD.n11611 0.019716
R40090 DVDD.n11790 DVDD.n11789 0.019716
R40091 DVDD.n11795 DVDD.n11610 0.019716
R40092 DVDD.n11795 DVDD.n11794 0.019716
R40093 DVDD.n11801 DVDD.n11609 0.019716
R40094 DVDD.n11802 DVDD.n11801 0.019716
R40095 DVDD.n11807 DVDD.n11608 0.019716
R40096 DVDD.n11807 DVDD.n11806 0.019716
R40097 DVDD.n11813 DVDD.n11607 0.019716
R40098 DVDD.n11814 DVDD.n11813 0.019716
R40099 DVDD.n11819 DVDD.n11606 0.019716
R40100 DVDD.n11819 DVDD.n11818 0.019716
R40101 DVDD.n11825 DVDD.n11605 0.019716
R40102 DVDD.n11826 DVDD.n11825 0.019716
R40103 DVDD.n11831 DVDD.n11604 0.019716
R40104 DVDD.n11831 DVDD.n11830 0.019716
R40105 DVDD.n11837 DVDD.n11603 0.019716
R40106 DVDD.n11838 DVDD.n11837 0.019716
R40107 DVDD.n11843 DVDD.n11602 0.019716
R40108 DVDD.n11843 DVDD.n11842 0.019716
R40109 DVDD.n11849 DVDD.n11601 0.019716
R40110 DVDD.n11850 DVDD.n11849 0.019716
R40111 DVDD.n11855 DVDD.n11600 0.019716
R40112 DVDD.n11855 DVDD.n11854 0.019716
R40113 DVDD.n11861 DVDD.n11599 0.019716
R40114 DVDD.n11862 DVDD.n11861 0.019716
R40115 DVDD.n11867 DVDD.n11598 0.019716
R40116 DVDD.n11867 DVDD.n11866 0.019716
R40117 DVDD.n11873 DVDD.n11597 0.019716
R40118 DVDD.n11874 DVDD.n11873 0.019716
R40119 DVDD.n11879 DVDD.n11596 0.019716
R40120 DVDD.n11879 DVDD.n11878 0.019716
R40121 DVDD.n11885 DVDD.n11595 0.019716
R40122 DVDD.n11886 DVDD.n11885 0.019716
R40123 DVDD.n11891 DVDD.n11594 0.019716
R40124 DVDD.n11891 DVDD.n11890 0.019716
R40125 DVDD.n11897 DVDD.n11593 0.019716
R40126 DVDD.n11898 DVDD.n11897 0.019716
R40127 DVDD.n11903 DVDD.n11592 0.019716
R40128 DVDD.n11903 DVDD.n11902 0.019716
R40129 DVDD.n11909 DVDD.n11591 0.019716
R40130 DVDD.n11910 DVDD.n11909 0.019716
R40131 DVDD.n11915 DVDD.n11590 0.019716
R40132 DVDD.n11915 DVDD.n11914 0.019716
R40133 DVDD.n13774 DVDD.n11589 0.019716
R40134 DVDD.n13775 DVDD.n13774 0.019716
R40135 DVDD.n12030 DVDD.n12029 0.019716
R40136 DVDD.n12034 DVDD.n12031 0.019716
R40137 DVDD.n12034 DVDD.n12033 0.019716
R40138 DVDD.n12040 DVDD.n12023 0.019716
R40139 DVDD.n12041 DVDD.n12040 0.019716
R40140 DVDD.n12046 DVDD.n12043 0.019716
R40141 DVDD.n12046 DVDD.n12045 0.019716
R40142 DVDD.n12052 DVDD.n12019 0.019716
R40143 DVDD.n12053 DVDD.n12052 0.019716
R40144 DVDD.n12058 DVDD.n12055 0.019716
R40145 DVDD.n12058 DVDD.n12057 0.019716
R40146 DVDD.n12064 DVDD.n12015 0.019716
R40147 DVDD.n12065 DVDD.n12064 0.019716
R40148 DVDD.n12070 DVDD.n12067 0.019716
R40149 DVDD.n12070 DVDD.n12069 0.019716
R40150 DVDD.n12076 DVDD.n12011 0.019716
R40151 DVDD.n12077 DVDD.n12076 0.019716
R40152 DVDD.n12082 DVDD.n12079 0.019716
R40153 DVDD.n12082 DVDD.n12081 0.019716
R40154 DVDD.n12088 DVDD.n12007 0.019716
R40155 DVDD.n12089 DVDD.n12088 0.019716
R40156 DVDD.n12094 DVDD.n12091 0.019716
R40157 DVDD.n12094 DVDD.n12093 0.019716
R40158 DVDD.n12100 DVDD.n12003 0.019716
R40159 DVDD.n12101 DVDD.n12100 0.019716
R40160 DVDD.n12106 DVDD.n12103 0.019716
R40161 DVDD.n12106 DVDD.n12105 0.019716
R40162 DVDD.n12112 DVDD.n11999 0.019716
R40163 DVDD.n12113 DVDD.n12112 0.019716
R40164 DVDD.n12118 DVDD.n12115 0.019716
R40165 DVDD.n12118 DVDD.n12117 0.019716
R40166 DVDD.n12124 DVDD.n11995 0.019716
R40167 DVDD.n12125 DVDD.n12124 0.019716
R40168 DVDD.n12130 DVDD.n12127 0.019716
R40169 DVDD.n12130 DVDD.n12129 0.019716
R40170 DVDD.n12136 DVDD.n11991 0.019716
R40171 DVDD.n12137 DVDD.n12136 0.019716
R40172 DVDD.n12142 DVDD.n12139 0.019716
R40173 DVDD.n12142 DVDD.n12141 0.019716
R40174 DVDD.n12148 DVDD.n11987 0.019716
R40175 DVDD.n12149 DVDD.n12148 0.019716
R40176 DVDD.n12154 DVDD.n12151 0.019716
R40177 DVDD.n12154 DVDD.n12153 0.019716
R40178 DVDD.n12160 DVDD.n11983 0.019716
R40179 DVDD.n12161 DVDD.n12160 0.019716
R40180 DVDD.n12166 DVDD.n12163 0.019716
R40181 DVDD.n12166 DVDD.n12165 0.019716
R40182 DVDD.n12172 DVDD.n11979 0.019716
R40183 DVDD.n12173 DVDD.n12172 0.019716
R40184 DVDD.n12178 DVDD.n12175 0.019716
R40185 DVDD.n12178 DVDD.n12177 0.019716
R40186 DVDD.n12184 DVDD.n11975 0.019716
R40187 DVDD.n12185 DVDD.n12184 0.019716
R40188 DVDD.n12190 DVDD.n12187 0.019716
R40189 DVDD.n12190 DVDD.n12189 0.019716
R40190 DVDD.n12196 DVDD.n11971 0.019716
R40191 DVDD.n12197 DVDD.n12196 0.019716
R40192 DVDD.n12202 DVDD.n12199 0.019716
R40193 DVDD.n12202 DVDD.n12201 0.019716
R40194 DVDD.n12208 DVDD.n11967 0.019716
R40195 DVDD.n12209 DVDD.n12208 0.019716
R40196 DVDD.n12214 DVDD.n12211 0.019716
R40197 DVDD.n12214 DVDD.n12213 0.019716
R40198 DVDD.n12220 DVDD.n11963 0.019716
R40199 DVDD.n12221 DVDD.n12220 0.019716
R40200 DVDD.n12226 DVDD.n12223 0.019716
R40201 DVDD.n12226 DVDD.n12225 0.019716
R40202 DVDD.n12232 DVDD.n11959 0.019716
R40203 DVDD.n12233 DVDD.n12232 0.019716
R40204 DVDD.n12238 DVDD.n12235 0.019716
R40205 DVDD.n12238 DVDD.n12237 0.019716
R40206 DVDD.n12244 DVDD.n11955 0.019716
R40207 DVDD.n12245 DVDD.n12244 0.019716
R40208 DVDD.n12250 DVDD.n12247 0.019716
R40209 DVDD.n12250 DVDD.n12249 0.019716
R40210 DVDD.n12256 DVDD.n11951 0.019716
R40211 DVDD.n12257 DVDD.n12256 0.019716
R40212 DVDD.n12262 DVDD.n12259 0.019716
R40213 DVDD.n12262 DVDD.n12261 0.019716
R40214 DVDD.n12269 DVDD.n11947 0.019716
R40215 DVDD.n12270 DVDD.n12269 0.019716
R40216 DVDD.n12273 DVDD.n12272 0.019716
R40217 DVDD.n12274 DVDD.n12273 0.019716
R40218 DVDD.n12375 DVDD.n12374 0.019716
R40219 DVDD.n13501 DVDD.n12328 0.019716
R40220 DVDD.n13502 DVDD.n13501 0.019716
R40221 DVDD.n13507 DVDD.n12327 0.019716
R40222 DVDD.n13507 DVDD.n13506 0.019716
R40223 DVDD.n13513 DVDD.n12326 0.019716
R40224 DVDD.n13514 DVDD.n13513 0.019716
R40225 DVDD.n13519 DVDD.n12325 0.019716
R40226 DVDD.n13519 DVDD.n13518 0.019716
R40227 DVDD.n13525 DVDD.n12324 0.019716
R40228 DVDD.n13526 DVDD.n13525 0.019716
R40229 DVDD.n13531 DVDD.n12323 0.019716
R40230 DVDD.n13531 DVDD.n13530 0.019716
R40231 DVDD.n13537 DVDD.n12322 0.019716
R40232 DVDD.n13538 DVDD.n13537 0.019716
R40233 DVDD.n13543 DVDD.n12321 0.019716
R40234 DVDD.n13543 DVDD.n13542 0.019716
R40235 DVDD.n13549 DVDD.n12320 0.019716
R40236 DVDD.n13550 DVDD.n13549 0.019716
R40237 DVDD.n13555 DVDD.n12319 0.019716
R40238 DVDD.n13555 DVDD.n13554 0.019716
R40239 DVDD.n13561 DVDD.n12318 0.019716
R40240 DVDD.n13562 DVDD.n13561 0.019716
R40241 DVDD.n13567 DVDD.n12317 0.019716
R40242 DVDD.n13567 DVDD.n13566 0.019716
R40243 DVDD.n13573 DVDD.n12316 0.019716
R40244 DVDD.n13574 DVDD.n13573 0.019716
R40245 DVDD.n13579 DVDD.n12315 0.019716
R40246 DVDD.n13579 DVDD.n13578 0.019716
R40247 DVDD.n13585 DVDD.n12314 0.019716
R40248 DVDD.n13586 DVDD.n13585 0.019716
R40249 DVDD.n13591 DVDD.n12313 0.019716
R40250 DVDD.n13591 DVDD.n13590 0.019716
R40251 DVDD.n13597 DVDD.n12312 0.019716
R40252 DVDD.n13598 DVDD.n13597 0.019716
R40253 DVDD.n13603 DVDD.n12311 0.019716
R40254 DVDD.n13603 DVDD.n13602 0.019716
R40255 DVDD.n13609 DVDD.n12310 0.019716
R40256 DVDD.n13610 DVDD.n13609 0.019716
R40257 DVDD.n13615 DVDD.n12309 0.019716
R40258 DVDD.n13615 DVDD.n13614 0.019716
R40259 DVDD.n13621 DVDD.n12308 0.019716
R40260 DVDD.n13622 DVDD.n13621 0.019716
R40261 DVDD.n13627 DVDD.n12307 0.019716
R40262 DVDD.n13627 DVDD.n13626 0.019716
R40263 DVDD.n13633 DVDD.n12306 0.019716
R40264 DVDD.n13634 DVDD.n13633 0.019716
R40265 DVDD.n13639 DVDD.n12305 0.019716
R40266 DVDD.n13639 DVDD.n13638 0.019716
R40267 DVDD.n13645 DVDD.n12304 0.019716
R40268 DVDD.n13646 DVDD.n13645 0.019716
R40269 DVDD.n13651 DVDD.n12303 0.019716
R40270 DVDD.n13651 DVDD.n13650 0.019716
R40271 DVDD.n13657 DVDD.n12302 0.019716
R40272 DVDD.n13658 DVDD.n13657 0.019716
R40273 DVDD.n13663 DVDD.n12301 0.019716
R40274 DVDD.n13663 DVDD.n13662 0.019716
R40275 DVDD.n13669 DVDD.n12300 0.019716
R40276 DVDD.n13670 DVDD.n13669 0.019716
R40277 DVDD.n13675 DVDD.n12299 0.019716
R40278 DVDD.n13675 DVDD.n13674 0.019716
R40279 DVDD.n13681 DVDD.n12298 0.019716
R40280 DVDD.n13682 DVDD.n13681 0.019716
R40281 DVDD.n13687 DVDD.n12297 0.019716
R40282 DVDD.n13687 DVDD.n13686 0.019716
R40283 DVDD.n13693 DVDD.n12296 0.019716
R40284 DVDD.n13694 DVDD.n13693 0.019716
R40285 DVDD.n13699 DVDD.n12295 0.019716
R40286 DVDD.n13699 DVDD.n13698 0.019716
R40287 DVDD.n13705 DVDD.n12294 0.019716
R40288 DVDD.n13706 DVDD.n13705 0.019716
R40289 DVDD.n13711 DVDD.n12293 0.019716
R40290 DVDD.n13711 DVDD.n13710 0.019716
R40291 DVDD.n13717 DVDD.n12292 0.019716
R40292 DVDD.n13718 DVDD.n13717 0.019716
R40293 DVDD.n13723 DVDD.n12291 0.019716
R40294 DVDD.n13723 DVDD.n13722 0.019716
R40295 DVDD.n13729 DVDD.n12290 0.019716
R40296 DVDD.n13730 DVDD.n13729 0.019716
R40297 DVDD.n13735 DVDD.n12289 0.019716
R40298 DVDD.n13735 DVDD.n13734 0.019716
R40299 DVDD.n13741 DVDD.n12288 0.019716
R40300 DVDD.n13742 DVDD.n13741 0.019716
R40301 DVDD.n13486 DVDD.n12433 0.019716
R40302 DVDD.n12539 DVDD.n12476 0.019716
R40303 DVDD.n12539 DVDD.n12431 0.019716
R40304 DVDD.n12548 DVDD.n12475 0.019716
R40305 DVDD.n12548 DVDD.n12430 0.019716
R40306 DVDD.n12536 DVDD.n12474 0.019716
R40307 DVDD.n12536 DVDD.n12429 0.019716
R40308 DVDD.n12557 DVDD.n12473 0.019716
R40309 DVDD.n12557 DVDD.n12428 0.019716
R40310 DVDD.n12533 DVDD.n12472 0.019716
R40311 DVDD.n12533 DVDD.n12427 0.019716
R40312 DVDD.n12566 DVDD.n12471 0.019716
R40313 DVDD.n12566 DVDD.n12426 0.019716
R40314 DVDD.n12530 DVDD.n12470 0.019716
R40315 DVDD.n12530 DVDD.n12425 0.019716
R40316 DVDD.n12575 DVDD.n12469 0.019716
R40317 DVDD.n12575 DVDD.n12424 0.019716
R40318 DVDD.n12527 DVDD.n12468 0.019716
R40319 DVDD.n12527 DVDD.n12423 0.019716
R40320 DVDD.n12584 DVDD.n12467 0.019716
R40321 DVDD.n12584 DVDD.n12422 0.019716
R40322 DVDD.n12524 DVDD.n12466 0.019716
R40323 DVDD.n12524 DVDD.n12421 0.019716
R40324 DVDD.n12593 DVDD.n12465 0.019716
R40325 DVDD.n12593 DVDD.n12420 0.019716
R40326 DVDD.n12521 DVDD.n12464 0.019716
R40327 DVDD.n12521 DVDD.n12419 0.019716
R40328 DVDD.n12602 DVDD.n12463 0.019716
R40329 DVDD.n12602 DVDD.n12418 0.019716
R40330 DVDD.n12518 DVDD.n12462 0.019716
R40331 DVDD.n12518 DVDD.n12417 0.019716
R40332 DVDD.n12611 DVDD.n12461 0.019716
R40333 DVDD.n12611 DVDD.n12416 0.019716
R40334 DVDD.n12515 DVDD.n12460 0.019716
R40335 DVDD.n12515 DVDD.n12415 0.019716
R40336 DVDD.n12620 DVDD.n12459 0.019716
R40337 DVDD.n12620 DVDD.n12414 0.019716
R40338 DVDD.n12512 DVDD.n12458 0.019716
R40339 DVDD.n12512 DVDD.n12413 0.019716
R40340 DVDD.n12629 DVDD.n12457 0.019716
R40341 DVDD.n12629 DVDD.n12412 0.019716
R40342 DVDD.n12509 DVDD.n12456 0.019716
R40343 DVDD.n12509 DVDD.n12411 0.019716
R40344 DVDD.n12638 DVDD.n12455 0.019716
R40345 DVDD.n12638 DVDD.n12410 0.019716
R40346 DVDD.n12506 DVDD.n12454 0.019716
R40347 DVDD.n12506 DVDD.n12409 0.019716
R40348 DVDD.n12647 DVDD.n12453 0.019716
R40349 DVDD.n12647 DVDD.n12408 0.019716
R40350 DVDD.n12503 DVDD.n12452 0.019716
R40351 DVDD.n12503 DVDD.n12407 0.019716
R40352 DVDD.n12656 DVDD.n12451 0.019716
R40353 DVDD.n12656 DVDD.n12406 0.019716
R40354 DVDD.n12500 DVDD.n12450 0.019716
R40355 DVDD.n12500 DVDD.n12405 0.019716
R40356 DVDD.n12665 DVDD.n12449 0.019716
R40357 DVDD.n12665 DVDD.n12404 0.019716
R40358 DVDD.n12497 DVDD.n12448 0.019716
R40359 DVDD.n12497 DVDD.n12403 0.019716
R40360 DVDD.n12674 DVDD.n12447 0.019716
R40361 DVDD.n12674 DVDD.n12402 0.019716
R40362 DVDD.n12494 DVDD.n12446 0.019716
R40363 DVDD.n12494 DVDD.n12401 0.019716
R40364 DVDD.n12683 DVDD.n12445 0.019716
R40365 DVDD.n12683 DVDD.n12400 0.019716
R40366 DVDD.n12491 DVDD.n12444 0.019716
R40367 DVDD.n12491 DVDD.n12399 0.019716
R40368 DVDD.n12692 DVDD.n12443 0.019716
R40369 DVDD.n12692 DVDD.n12398 0.019716
R40370 DVDD.n12488 DVDD.n12442 0.019716
R40371 DVDD.n12488 DVDD.n12397 0.019716
R40372 DVDD.n12701 DVDD.n12441 0.019716
R40373 DVDD.n12701 DVDD.n12396 0.019716
R40374 DVDD.n12485 DVDD.n12440 0.019716
R40375 DVDD.n12485 DVDD.n12395 0.019716
R40376 DVDD.n12710 DVDD.n12439 0.019716
R40377 DVDD.n12710 DVDD.n12394 0.019716
R40378 DVDD.n12482 DVDD.n12438 0.019716
R40379 DVDD.n12482 DVDD.n12393 0.019716
R40380 DVDD.n12719 DVDD.n12437 0.019716
R40381 DVDD.n12719 DVDD.n12392 0.019716
R40382 DVDD.n12479 DVDD.n12436 0.019716
R40383 DVDD.n12479 DVDD.n12391 0.019716
R40384 DVDD.n13472 DVDD.n12780 0.019716
R40385 DVDD.n12886 DVDD.n12824 0.019716
R40386 DVDD.n12886 DVDD.n12778 0.019716
R40387 DVDD.n13290 DVDD.n12823 0.019716
R40388 DVDD.n13290 DVDD.n12777 0.019716
R40389 DVDD.n12883 DVDD.n12822 0.019716
R40390 DVDD.n12883 DVDD.n12776 0.019716
R40391 DVDD.n13299 DVDD.n12821 0.019716
R40392 DVDD.n13299 DVDD.n12775 0.019716
R40393 DVDD.n12880 DVDD.n12820 0.019716
R40394 DVDD.n12880 DVDD.n12774 0.019716
R40395 DVDD.n13308 DVDD.n12819 0.019716
R40396 DVDD.n13308 DVDD.n12773 0.019716
R40397 DVDD.n12877 DVDD.n12818 0.019716
R40398 DVDD.n12877 DVDD.n12772 0.019716
R40399 DVDD.n13317 DVDD.n12817 0.019716
R40400 DVDD.n13317 DVDD.n12771 0.019716
R40401 DVDD.n12874 DVDD.n12816 0.019716
R40402 DVDD.n12874 DVDD.n12770 0.019716
R40403 DVDD.n13326 DVDD.n12815 0.019716
R40404 DVDD.n13326 DVDD.n12769 0.019716
R40405 DVDD.n12871 DVDD.n12814 0.019716
R40406 DVDD.n12871 DVDD.n12768 0.019716
R40407 DVDD.n13335 DVDD.n12813 0.019716
R40408 DVDD.n13335 DVDD.n12767 0.019716
R40409 DVDD.n12868 DVDD.n12812 0.019716
R40410 DVDD.n12868 DVDD.n12766 0.019716
R40411 DVDD.n13344 DVDD.n12811 0.019716
R40412 DVDD.n13344 DVDD.n12765 0.019716
R40413 DVDD.n12865 DVDD.n12810 0.019716
R40414 DVDD.n12865 DVDD.n12764 0.019716
R40415 DVDD.n13353 DVDD.n12809 0.019716
R40416 DVDD.n13353 DVDD.n12763 0.019716
R40417 DVDD.n12862 DVDD.n12808 0.019716
R40418 DVDD.n12862 DVDD.n12762 0.019716
R40419 DVDD.n13362 DVDD.n12807 0.019716
R40420 DVDD.n13362 DVDD.n12761 0.019716
R40421 DVDD.n12859 DVDD.n12806 0.019716
R40422 DVDD.n12859 DVDD.n12760 0.019716
R40423 DVDD.n13371 DVDD.n12805 0.019716
R40424 DVDD.n13371 DVDD.n12759 0.019716
R40425 DVDD.n12856 DVDD.n12804 0.019716
R40426 DVDD.n12856 DVDD.n12758 0.019716
R40427 DVDD.n13380 DVDD.n12803 0.019716
R40428 DVDD.n13380 DVDD.n12757 0.019716
R40429 DVDD.n12853 DVDD.n12802 0.019716
R40430 DVDD.n12853 DVDD.n12756 0.019716
R40431 DVDD.n13389 DVDD.n12801 0.019716
R40432 DVDD.n13389 DVDD.n12755 0.019716
R40433 DVDD.n12850 DVDD.n12800 0.019716
R40434 DVDD.n12850 DVDD.n12754 0.019716
R40435 DVDD.n13398 DVDD.n12799 0.019716
R40436 DVDD.n13398 DVDD.n12753 0.019716
R40437 DVDD.n12847 DVDD.n12798 0.019716
R40438 DVDD.n12847 DVDD.n12752 0.019716
R40439 DVDD.n13407 DVDD.n12797 0.019716
R40440 DVDD.n13407 DVDD.n12751 0.019716
R40441 DVDD.n12844 DVDD.n12796 0.019716
R40442 DVDD.n12844 DVDD.n12750 0.019716
R40443 DVDD.n13416 DVDD.n12795 0.019716
R40444 DVDD.n13416 DVDD.n12749 0.019716
R40445 DVDD.n12841 DVDD.n12794 0.019716
R40446 DVDD.n12841 DVDD.n12748 0.019716
R40447 DVDD.n13425 DVDD.n12793 0.019716
R40448 DVDD.n13425 DVDD.n12747 0.019716
R40449 DVDD.n12838 DVDD.n12792 0.019716
R40450 DVDD.n12838 DVDD.n12746 0.019716
R40451 DVDD.n13434 DVDD.n12791 0.019716
R40452 DVDD.n13434 DVDD.n12745 0.019716
R40453 DVDD.n12835 DVDD.n12790 0.019716
R40454 DVDD.n12835 DVDD.n12744 0.019716
R40455 DVDD.n13443 DVDD.n12789 0.019716
R40456 DVDD.n13443 DVDD.n12743 0.019716
R40457 DVDD.n12832 DVDD.n12788 0.019716
R40458 DVDD.n12832 DVDD.n12742 0.019716
R40459 DVDD.n13452 DVDD.n12787 0.019716
R40460 DVDD.n13452 DVDD.n12741 0.019716
R40461 DVDD.n12829 DVDD.n12786 0.019716
R40462 DVDD.n12829 DVDD.n12740 0.019716
R40463 DVDD.n13461 DVDD.n12785 0.019716
R40464 DVDD.n13461 DVDD.n12739 0.019716
R40465 DVDD.n12826 DVDD.n12784 0.019716
R40466 DVDD.n12826 DVDD.n12738 0.019716
R40467 DVDD.n13255 DVDD.n12964 0.019716
R40468 DVDD.n12966 DVDD.n12965 0.019716
R40469 DVDD.n12966 DVDD.n12963 0.019716
R40470 DVDD.n13246 DVDD.n13245 0.019716
R40471 DVDD.n13245 DVDD.n12962 0.019716
R40472 DVDD.n13241 DVDD.n13240 0.019716
R40473 DVDD.n13240 DVDD.n12961 0.019716
R40474 DVDD.n13234 DVDD.n13233 0.019716
R40475 DVDD.n13233 DVDD.n12960 0.019716
R40476 DVDD.n13229 DVDD.n13228 0.019716
R40477 DVDD.n13228 DVDD.n12959 0.019716
R40478 DVDD.n13222 DVDD.n13221 0.019716
R40479 DVDD.n13221 DVDD.n12958 0.019716
R40480 DVDD.n13217 DVDD.n13216 0.019716
R40481 DVDD.n13216 DVDD.n12957 0.019716
R40482 DVDD.n13210 DVDD.n13209 0.019716
R40483 DVDD.n13209 DVDD.n12956 0.019716
R40484 DVDD.n13205 DVDD.n13204 0.019716
R40485 DVDD.n13204 DVDD.n12955 0.019716
R40486 DVDD.n13198 DVDD.n13197 0.019716
R40487 DVDD.n13197 DVDD.n12954 0.019716
R40488 DVDD.n13193 DVDD.n13192 0.019716
R40489 DVDD.n13192 DVDD.n12953 0.019716
R40490 DVDD.n13186 DVDD.n13185 0.019716
R40491 DVDD.n13185 DVDD.n12952 0.019716
R40492 DVDD.n13181 DVDD.n13180 0.019716
R40493 DVDD.n13180 DVDD.n12951 0.019716
R40494 DVDD.n13174 DVDD.n13173 0.019716
R40495 DVDD.n13173 DVDD.n12950 0.019716
R40496 DVDD.n13169 DVDD.n13168 0.019716
R40497 DVDD.n13168 DVDD.n12949 0.019716
R40498 DVDD.n13162 DVDD.n13161 0.019716
R40499 DVDD.n13161 DVDD.n12948 0.019716
R40500 DVDD.n13157 DVDD.n13156 0.019716
R40501 DVDD.n13156 DVDD.n12947 0.019716
R40502 DVDD.n13150 DVDD.n13149 0.019716
R40503 DVDD.n13149 DVDD.n12946 0.019716
R40504 DVDD.n13145 DVDD.n13144 0.019716
R40505 DVDD.n13144 DVDD.n12945 0.019716
R40506 DVDD.n13138 DVDD.n13137 0.019716
R40507 DVDD.n13137 DVDD.n12944 0.019716
R40508 DVDD.n13133 DVDD.n13132 0.019716
R40509 DVDD.n13132 DVDD.n12943 0.019716
R40510 DVDD.n13126 DVDD.n13125 0.019716
R40511 DVDD.n13125 DVDD.n12942 0.019716
R40512 DVDD.n13121 DVDD.n13120 0.019716
R40513 DVDD.n13120 DVDD.n12941 0.019716
R40514 DVDD.n13114 DVDD.n13113 0.019716
R40515 DVDD.n13113 DVDD.n12940 0.019716
R40516 DVDD.n13109 DVDD.n13108 0.019716
R40517 DVDD.n13108 DVDD.n12939 0.019716
R40518 DVDD.n13102 DVDD.n13101 0.019716
R40519 DVDD.n13101 DVDD.n12938 0.019716
R40520 DVDD.n13097 DVDD.n13096 0.019716
R40521 DVDD.n13096 DVDD.n12937 0.019716
R40522 DVDD.n13090 DVDD.n13089 0.019716
R40523 DVDD.n13089 DVDD.n12936 0.019716
R40524 DVDD.n13085 DVDD.n13084 0.019716
R40525 DVDD.n13084 DVDD.n12935 0.019716
R40526 DVDD.n13078 DVDD.n13077 0.019716
R40527 DVDD.n13077 DVDD.n12934 0.019716
R40528 DVDD.n13073 DVDD.n13072 0.019716
R40529 DVDD.n13072 DVDD.n12933 0.019716
R40530 DVDD.n13066 DVDD.n13065 0.019716
R40531 DVDD.n13065 DVDD.n12932 0.019716
R40532 DVDD.n13061 DVDD.n13060 0.019716
R40533 DVDD.n13060 DVDD.n12931 0.019716
R40534 DVDD.n13054 DVDD.n13053 0.019716
R40535 DVDD.n13053 DVDD.n12930 0.019716
R40536 DVDD.n13049 DVDD.n13048 0.019716
R40537 DVDD.n13048 DVDD.n12929 0.019716
R40538 DVDD.n13042 DVDD.n13041 0.019716
R40539 DVDD.n13041 DVDD.n12928 0.019716
R40540 DVDD.n13037 DVDD.n13036 0.019716
R40541 DVDD.n13036 DVDD.n12927 0.019716
R40542 DVDD.n13030 DVDD.n13029 0.019716
R40543 DVDD.n13029 DVDD.n12926 0.019716
R40544 DVDD.n13025 DVDD.n13024 0.019716
R40545 DVDD.n13024 DVDD.n12925 0.019716
R40546 DVDD.n13018 DVDD.n13017 0.019716
R40547 DVDD.n13017 DVDD.n12924 0.019716
R40548 DVDD.n13013 DVDD.n13012 0.019716
R40549 DVDD.n13012 DVDD.n12923 0.019716
R40550 DVDD.n2252 DVDD.n2251 0.019716
R40551 DVDD.n16461 DVDD.n2206 0.019716
R40552 DVDD.n16462 DVDD.n16461 0.019716
R40553 DVDD.n16467 DVDD.n2205 0.019716
R40554 DVDD.n16467 DVDD.n16466 0.019716
R40555 DVDD.n16473 DVDD.n2204 0.019716
R40556 DVDD.n16474 DVDD.n16473 0.019716
R40557 DVDD.n16479 DVDD.n2203 0.019716
R40558 DVDD.n16479 DVDD.n16478 0.019716
R40559 DVDD.n16485 DVDD.n2202 0.019716
R40560 DVDD.n16486 DVDD.n16485 0.019716
R40561 DVDD.n16491 DVDD.n2201 0.019716
R40562 DVDD.n16491 DVDD.n16490 0.019716
R40563 DVDD.n16497 DVDD.n2200 0.019716
R40564 DVDD.n16498 DVDD.n16497 0.019716
R40565 DVDD.n16503 DVDD.n2199 0.019716
R40566 DVDD.n16503 DVDD.n16502 0.019716
R40567 DVDD.n16509 DVDD.n2198 0.019716
R40568 DVDD.n16510 DVDD.n16509 0.019716
R40569 DVDD.n16515 DVDD.n2197 0.019716
R40570 DVDD.n16515 DVDD.n16514 0.019716
R40571 DVDD.n16521 DVDD.n2196 0.019716
R40572 DVDD.n16522 DVDD.n16521 0.019716
R40573 DVDD.n16527 DVDD.n2195 0.019716
R40574 DVDD.n16527 DVDD.n16526 0.019716
R40575 DVDD.n16533 DVDD.n2194 0.019716
R40576 DVDD.n16534 DVDD.n16533 0.019716
R40577 DVDD.n16539 DVDD.n2193 0.019716
R40578 DVDD.n16539 DVDD.n16538 0.019716
R40579 DVDD.n16545 DVDD.n2192 0.019716
R40580 DVDD.n16546 DVDD.n16545 0.019716
R40581 DVDD.n16551 DVDD.n2191 0.019716
R40582 DVDD.n16551 DVDD.n16550 0.019716
R40583 DVDD.n16557 DVDD.n2190 0.019716
R40584 DVDD.n16558 DVDD.n16557 0.019716
R40585 DVDD.n16563 DVDD.n2189 0.019716
R40586 DVDD.n16563 DVDD.n16562 0.019716
R40587 DVDD.n16569 DVDD.n2188 0.019716
R40588 DVDD.n16570 DVDD.n16569 0.019716
R40589 DVDD.n16575 DVDD.n2187 0.019716
R40590 DVDD.n16575 DVDD.n16574 0.019716
R40591 DVDD.n16581 DVDD.n2186 0.019716
R40592 DVDD.n16582 DVDD.n16581 0.019716
R40593 DVDD.n16587 DVDD.n2185 0.019716
R40594 DVDD.n16587 DVDD.n16586 0.019716
R40595 DVDD.n16593 DVDD.n2184 0.019716
R40596 DVDD.n16594 DVDD.n16593 0.019716
R40597 DVDD.n16599 DVDD.n2183 0.019716
R40598 DVDD.n16599 DVDD.n16598 0.019716
R40599 DVDD.n16605 DVDD.n2182 0.019716
R40600 DVDD.n16606 DVDD.n16605 0.019716
R40601 DVDD.n16611 DVDD.n2181 0.019716
R40602 DVDD.n16611 DVDD.n16610 0.019716
R40603 DVDD.n16617 DVDD.n2180 0.019716
R40604 DVDD.n16618 DVDD.n16617 0.019716
R40605 DVDD.n16623 DVDD.n2179 0.019716
R40606 DVDD.n16623 DVDD.n16622 0.019716
R40607 DVDD.n16629 DVDD.n2178 0.019716
R40608 DVDD.n16630 DVDD.n16629 0.019716
R40609 DVDD.n16635 DVDD.n2177 0.019716
R40610 DVDD.n16635 DVDD.n16634 0.019716
R40611 DVDD.n16641 DVDD.n2176 0.019716
R40612 DVDD.n16642 DVDD.n16641 0.019716
R40613 DVDD.n16647 DVDD.n2175 0.019716
R40614 DVDD.n16647 DVDD.n16646 0.019716
R40615 DVDD.n16653 DVDD.n2174 0.019716
R40616 DVDD.n16654 DVDD.n16653 0.019716
R40617 DVDD.n16659 DVDD.n2173 0.019716
R40618 DVDD.n16659 DVDD.n16658 0.019716
R40619 DVDD.n16665 DVDD.n2172 0.019716
R40620 DVDD.n16666 DVDD.n16665 0.019716
R40621 DVDD.n16671 DVDD.n2171 0.019716
R40622 DVDD.n16671 DVDD.n16670 0.019716
R40623 DVDD.n16677 DVDD.n2170 0.019716
R40624 DVDD.n16678 DVDD.n16677 0.019716
R40625 DVDD.n16683 DVDD.n2169 0.019716
R40626 DVDD.n16683 DVDD.n16682 0.019716
R40627 DVDD.n16689 DVDD.n2168 0.019716
R40628 DVDD.n16690 DVDD.n16689 0.019716
R40629 DVDD.n16695 DVDD.n2167 0.019716
R40630 DVDD.n16695 DVDD.n16694 0.019716
R40631 DVDD.n16701 DVDD.n2166 0.019716
R40632 DVDD.n16702 DVDD.n16701 0.019716
R40633 DVDD.n2155 DVDD.n1863 0.019716
R40634 DVDD.n1865 DVDD.n1864 0.019716
R40635 DVDD.n1865 DVDD.n1862 0.019716
R40636 DVDD.n2146 DVDD.n2145 0.019716
R40637 DVDD.n2145 DVDD.n1861 0.019716
R40638 DVDD.n2141 DVDD.n2140 0.019716
R40639 DVDD.n2140 DVDD.n1860 0.019716
R40640 DVDD.n2134 DVDD.n2133 0.019716
R40641 DVDD.n2133 DVDD.n1859 0.019716
R40642 DVDD.n2129 DVDD.n2128 0.019716
R40643 DVDD.n2128 DVDD.n1858 0.019716
R40644 DVDD.n2122 DVDD.n2121 0.019716
R40645 DVDD.n2121 DVDD.n1857 0.019716
R40646 DVDD.n2117 DVDD.n2116 0.019716
R40647 DVDD.n2116 DVDD.n1856 0.019716
R40648 DVDD.n2110 DVDD.n2109 0.019716
R40649 DVDD.n2109 DVDD.n1855 0.019716
R40650 DVDD.n2105 DVDD.n2104 0.019716
R40651 DVDD.n2104 DVDD.n1854 0.019716
R40652 DVDD.n2098 DVDD.n2097 0.019716
R40653 DVDD.n2097 DVDD.n1853 0.019716
R40654 DVDD.n2093 DVDD.n2092 0.019716
R40655 DVDD.n2092 DVDD.n1852 0.019716
R40656 DVDD.n2086 DVDD.n2085 0.019716
R40657 DVDD.n2085 DVDD.n1851 0.019716
R40658 DVDD.n2081 DVDD.n2080 0.019716
R40659 DVDD.n2080 DVDD.n1850 0.019716
R40660 DVDD.n2074 DVDD.n2073 0.019716
R40661 DVDD.n2073 DVDD.n1849 0.019716
R40662 DVDD.n2069 DVDD.n2068 0.019716
R40663 DVDD.n2068 DVDD.n1848 0.019716
R40664 DVDD.n2062 DVDD.n2061 0.019716
R40665 DVDD.n2061 DVDD.n1847 0.019716
R40666 DVDD.n2057 DVDD.n2056 0.019716
R40667 DVDD.n2056 DVDD.n1846 0.019716
R40668 DVDD.n2050 DVDD.n2049 0.019716
R40669 DVDD.n2049 DVDD.n1845 0.019716
R40670 DVDD.n2045 DVDD.n2044 0.019716
R40671 DVDD.n2044 DVDD.n1844 0.019716
R40672 DVDD.n2038 DVDD.n2037 0.019716
R40673 DVDD.n2037 DVDD.n1843 0.019716
R40674 DVDD.n2033 DVDD.n2032 0.019716
R40675 DVDD.n2032 DVDD.n1842 0.019716
R40676 DVDD.n2026 DVDD.n2025 0.019716
R40677 DVDD.n2025 DVDD.n1841 0.019716
R40678 DVDD.n2021 DVDD.n2020 0.019716
R40679 DVDD.n2020 DVDD.n1840 0.019716
R40680 DVDD.n2014 DVDD.n2013 0.019716
R40681 DVDD.n2013 DVDD.n1839 0.019716
R40682 DVDD.n2009 DVDD.n2008 0.019716
R40683 DVDD.n2008 DVDD.n1838 0.019716
R40684 DVDD.n2002 DVDD.n2001 0.019716
R40685 DVDD.n2001 DVDD.n1837 0.019716
R40686 DVDD.n1997 DVDD.n1996 0.019716
R40687 DVDD.n1996 DVDD.n1836 0.019716
R40688 DVDD.n1990 DVDD.n1989 0.019716
R40689 DVDD.n1989 DVDD.n1835 0.019716
R40690 DVDD.n1985 DVDD.n1984 0.019716
R40691 DVDD.n1984 DVDD.n1834 0.019716
R40692 DVDD.n1978 DVDD.n1977 0.019716
R40693 DVDD.n1977 DVDD.n1833 0.019716
R40694 DVDD.n1973 DVDD.n1972 0.019716
R40695 DVDD.n1972 DVDD.n1832 0.019716
R40696 DVDD.n1966 DVDD.n1965 0.019716
R40697 DVDD.n1965 DVDD.n1831 0.019716
R40698 DVDD.n1961 DVDD.n1960 0.019716
R40699 DVDD.n1960 DVDD.n1830 0.019716
R40700 DVDD.n1954 DVDD.n1953 0.019716
R40701 DVDD.n1953 DVDD.n1829 0.019716
R40702 DVDD.n1949 DVDD.n1948 0.019716
R40703 DVDD.n1948 DVDD.n1828 0.019716
R40704 DVDD.n1942 DVDD.n1941 0.019716
R40705 DVDD.n1941 DVDD.n1827 0.019716
R40706 DVDD.n1937 DVDD.n1936 0.019716
R40707 DVDD.n1936 DVDD.n1826 0.019716
R40708 DVDD.n1930 DVDD.n1929 0.019716
R40709 DVDD.n1929 DVDD.n1825 0.019716
R40710 DVDD.n1925 DVDD.n1924 0.019716
R40711 DVDD.n1924 DVDD.n1824 0.019716
R40712 DVDD.n1918 DVDD.n1917 0.019716
R40713 DVDD.n1917 DVDD.n1823 0.019716
R40714 DVDD.n1913 DVDD.n1912 0.019716
R40715 DVDD.n1912 DVDD.n1822 0.019716
R40716 DVDD.n1799 DVDD.n1798 0.019716
R40717 DVDD.n16750 DVDD.n1753 0.019716
R40718 DVDD.n16751 DVDD.n16750 0.019716
R40719 DVDD.n16756 DVDD.n1752 0.019716
R40720 DVDD.n16756 DVDD.n16755 0.019716
R40721 DVDD.n16762 DVDD.n1751 0.019716
R40722 DVDD.n16763 DVDD.n16762 0.019716
R40723 DVDD.n16768 DVDD.n1750 0.019716
R40724 DVDD.n16768 DVDD.n16767 0.019716
R40725 DVDD.n16774 DVDD.n1749 0.019716
R40726 DVDD.n16775 DVDD.n16774 0.019716
R40727 DVDD.n16780 DVDD.n1748 0.019716
R40728 DVDD.n16780 DVDD.n16779 0.019716
R40729 DVDD.n16786 DVDD.n1747 0.019716
R40730 DVDD.n16787 DVDD.n16786 0.019716
R40731 DVDD.n16792 DVDD.n1746 0.019716
R40732 DVDD.n16792 DVDD.n16791 0.019716
R40733 DVDD.n16798 DVDD.n1745 0.019716
R40734 DVDD.n16799 DVDD.n16798 0.019716
R40735 DVDD.n16804 DVDD.n1744 0.019716
R40736 DVDD.n16804 DVDD.n16803 0.019716
R40737 DVDD.n16810 DVDD.n1743 0.019716
R40738 DVDD.n16811 DVDD.n16810 0.019716
R40739 DVDD.n16816 DVDD.n1742 0.019716
R40740 DVDD.n16816 DVDD.n16815 0.019716
R40741 DVDD.n16822 DVDD.n1741 0.019716
R40742 DVDD.n16823 DVDD.n16822 0.019716
R40743 DVDD.n16828 DVDD.n1740 0.019716
R40744 DVDD.n16828 DVDD.n16827 0.019716
R40745 DVDD.n16834 DVDD.n1739 0.019716
R40746 DVDD.n16835 DVDD.n16834 0.019716
R40747 DVDD.n16840 DVDD.n1738 0.019716
R40748 DVDD.n16840 DVDD.n16839 0.019716
R40749 DVDD.n16846 DVDD.n1737 0.019716
R40750 DVDD.n16847 DVDD.n16846 0.019716
R40751 DVDD.n16852 DVDD.n1736 0.019716
R40752 DVDD.n16852 DVDD.n16851 0.019716
R40753 DVDD.n16858 DVDD.n1735 0.019716
R40754 DVDD.n16859 DVDD.n16858 0.019716
R40755 DVDD.n16864 DVDD.n1734 0.019716
R40756 DVDD.n16864 DVDD.n16863 0.019716
R40757 DVDD.n16870 DVDD.n1733 0.019716
R40758 DVDD.n16871 DVDD.n16870 0.019716
R40759 DVDD.n16876 DVDD.n1732 0.019716
R40760 DVDD.n16876 DVDD.n16875 0.019716
R40761 DVDD.n16882 DVDD.n1731 0.019716
R40762 DVDD.n16883 DVDD.n16882 0.019716
R40763 DVDD.n16888 DVDD.n1730 0.019716
R40764 DVDD.n16888 DVDD.n16887 0.019716
R40765 DVDD.n16894 DVDD.n1729 0.019716
R40766 DVDD.n16895 DVDD.n16894 0.019716
R40767 DVDD.n16900 DVDD.n1728 0.019716
R40768 DVDD.n16900 DVDD.n16899 0.019716
R40769 DVDD.n16906 DVDD.n1727 0.019716
R40770 DVDD.n16907 DVDD.n16906 0.019716
R40771 DVDD.n16912 DVDD.n1726 0.019716
R40772 DVDD.n16912 DVDD.n16911 0.019716
R40773 DVDD.n16918 DVDD.n1725 0.019716
R40774 DVDD.n16919 DVDD.n16918 0.019716
R40775 DVDD.n16924 DVDD.n1724 0.019716
R40776 DVDD.n16924 DVDD.n16923 0.019716
R40777 DVDD.n16930 DVDD.n1723 0.019716
R40778 DVDD.n16931 DVDD.n16930 0.019716
R40779 DVDD.n16936 DVDD.n1722 0.019716
R40780 DVDD.n16936 DVDD.n16935 0.019716
R40781 DVDD.n16942 DVDD.n1721 0.019716
R40782 DVDD.n16943 DVDD.n16942 0.019716
R40783 DVDD.n16948 DVDD.n1720 0.019716
R40784 DVDD.n16948 DVDD.n16947 0.019716
R40785 DVDD.n16954 DVDD.n1719 0.019716
R40786 DVDD.n16955 DVDD.n16954 0.019716
R40787 DVDD.n16960 DVDD.n1718 0.019716
R40788 DVDD.n16960 DVDD.n16959 0.019716
R40789 DVDD.n16966 DVDD.n1717 0.019716
R40790 DVDD.n16967 DVDD.n16966 0.019716
R40791 DVDD.n16972 DVDD.n1716 0.019716
R40792 DVDD.n16972 DVDD.n16971 0.019716
R40793 DVDD.n16978 DVDD.n1715 0.019716
R40794 DVDD.n16979 DVDD.n16978 0.019716
R40795 DVDD.n16984 DVDD.n1714 0.019716
R40796 DVDD.n16984 DVDD.n16983 0.019716
R40797 DVDD.n16991 DVDD.n1713 0.019716
R40798 DVDD.n16992 DVDD.n16991 0.019716
R40799 DVDD.n1700 DVDD.n1699 0.019716
R40800 DVDD.n17018 DVDD.n1652 0.019716
R40801 DVDD.n17019 DVDD.n17018 0.019716
R40802 DVDD.n17024 DVDD.n1651 0.019716
R40803 DVDD.n17024 DVDD.n17023 0.019716
R40804 DVDD.n17030 DVDD.n1650 0.019716
R40805 DVDD.n17031 DVDD.n17030 0.019716
R40806 DVDD.n17036 DVDD.n1649 0.019716
R40807 DVDD.n17036 DVDD.n17035 0.019716
R40808 DVDD.n17042 DVDD.n1648 0.019716
R40809 DVDD.n17043 DVDD.n17042 0.019716
R40810 DVDD.n17048 DVDD.n1647 0.019716
R40811 DVDD.n17048 DVDD.n17047 0.019716
R40812 DVDD.n17054 DVDD.n1646 0.019716
R40813 DVDD.n17055 DVDD.n17054 0.019716
R40814 DVDD.n17060 DVDD.n1645 0.019716
R40815 DVDD.n17060 DVDD.n17059 0.019716
R40816 DVDD.n17066 DVDD.n1644 0.019716
R40817 DVDD.n17067 DVDD.n17066 0.019716
R40818 DVDD.n17072 DVDD.n1643 0.019716
R40819 DVDD.n17072 DVDD.n17071 0.019716
R40820 DVDD.n17078 DVDD.n1642 0.019716
R40821 DVDD.n17079 DVDD.n17078 0.019716
R40822 DVDD.n17084 DVDD.n1641 0.019716
R40823 DVDD.n17084 DVDD.n17083 0.019716
R40824 DVDD.n17090 DVDD.n1640 0.019716
R40825 DVDD.n17091 DVDD.n17090 0.019716
R40826 DVDD.n17096 DVDD.n1639 0.019716
R40827 DVDD.n17096 DVDD.n17095 0.019716
R40828 DVDD.n17102 DVDD.n1638 0.019716
R40829 DVDD.n17103 DVDD.n17102 0.019716
R40830 DVDD.n17108 DVDD.n1637 0.019716
R40831 DVDD.n17108 DVDD.n17107 0.019716
R40832 DVDD.n17114 DVDD.n1636 0.019716
R40833 DVDD.n17115 DVDD.n17114 0.019716
R40834 DVDD.n17120 DVDD.n1635 0.019716
R40835 DVDD.n17120 DVDD.n17119 0.019716
R40836 DVDD.n17126 DVDD.n1634 0.019716
R40837 DVDD.n17127 DVDD.n17126 0.019716
R40838 DVDD.n17132 DVDD.n1633 0.019716
R40839 DVDD.n17132 DVDD.n17131 0.019716
R40840 DVDD.n17138 DVDD.n1632 0.019716
R40841 DVDD.n17139 DVDD.n17138 0.019716
R40842 DVDD.n17144 DVDD.n1631 0.019716
R40843 DVDD.n17144 DVDD.n17143 0.019716
R40844 DVDD.n17150 DVDD.n1630 0.019716
R40845 DVDD.n17151 DVDD.n17150 0.019716
R40846 DVDD.n17156 DVDD.n1629 0.019716
R40847 DVDD.n17156 DVDD.n17155 0.019716
R40848 DVDD.n17162 DVDD.n1628 0.019716
R40849 DVDD.n17163 DVDD.n17162 0.019716
R40850 DVDD.n17168 DVDD.n1627 0.019716
R40851 DVDD.n17168 DVDD.n17167 0.019716
R40852 DVDD.n17174 DVDD.n1626 0.019716
R40853 DVDD.n17175 DVDD.n17174 0.019716
R40854 DVDD.n17180 DVDD.n1625 0.019716
R40855 DVDD.n17180 DVDD.n17179 0.019716
R40856 DVDD.n17186 DVDD.n1624 0.019716
R40857 DVDD.n17187 DVDD.n17186 0.019716
R40858 DVDD.n17192 DVDD.n1623 0.019716
R40859 DVDD.n17192 DVDD.n17191 0.019716
R40860 DVDD.n17198 DVDD.n1622 0.019716
R40861 DVDD.n17199 DVDD.n17198 0.019716
R40862 DVDD.n17204 DVDD.n1621 0.019716
R40863 DVDD.n17204 DVDD.n17203 0.019716
R40864 DVDD.n17210 DVDD.n1620 0.019716
R40865 DVDD.n17211 DVDD.n17210 0.019716
R40866 DVDD.n17216 DVDD.n1619 0.019716
R40867 DVDD.n17216 DVDD.n17215 0.019716
R40868 DVDD.n17222 DVDD.n1618 0.019716
R40869 DVDD.n17223 DVDD.n17222 0.019716
R40870 DVDD.n17228 DVDD.n1617 0.019716
R40871 DVDD.n17228 DVDD.n17227 0.019716
R40872 DVDD.n17234 DVDD.n1616 0.019716
R40873 DVDD.n17235 DVDD.n17234 0.019716
R40874 DVDD.n17240 DVDD.n1615 0.019716
R40875 DVDD.n17240 DVDD.n17239 0.019716
R40876 DVDD.n17246 DVDD.n1614 0.019716
R40877 DVDD.n17247 DVDD.n17246 0.019716
R40878 DVDD.n17252 DVDD.n1613 0.019716
R40879 DVDD.n17252 DVDD.n17251 0.019716
R40880 DVDD.n17259 DVDD.n1612 0.019716
R40881 DVDD.n17260 DVDD.n17259 0.019716
R40882 DVDD.n1604 DVDD.n1312 0.019716
R40883 DVDD.n1314 DVDD.n1313 0.019716
R40884 DVDD.n1314 DVDD.n1311 0.019716
R40885 DVDD.n1595 DVDD.n1594 0.019716
R40886 DVDD.n1594 DVDD.n1310 0.019716
R40887 DVDD.n1590 DVDD.n1589 0.019716
R40888 DVDD.n1589 DVDD.n1309 0.019716
R40889 DVDD.n1583 DVDD.n1582 0.019716
R40890 DVDD.n1582 DVDD.n1308 0.019716
R40891 DVDD.n1578 DVDD.n1577 0.019716
R40892 DVDD.n1577 DVDD.n1307 0.019716
R40893 DVDD.n1571 DVDD.n1570 0.019716
R40894 DVDD.n1570 DVDD.n1306 0.019716
R40895 DVDD.n1566 DVDD.n1565 0.019716
R40896 DVDD.n1565 DVDD.n1305 0.019716
R40897 DVDD.n1559 DVDD.n1558 0.019716
R40898 DVDD.n1558 DVDD.n1304 0.019716
R40899 DVDD.n1554 DVDD.n1553 0.019716
R40900 DVDD.n1553 DVDD.n1303 0.019716
R40901 DVDD.n1547 DVDD.n1546 0.019716
R40902 DVDD.n1546 DVDD.n1302 0.019716
R40903 DVDD.n1542 DVDD.n1541 0.019716
R40904 DVDD.n1541 DVDD.n1301 0.019716
R40905 DVDD.n1535 DVDD.n1534 0.019716
R40906 DVDD.n1534 DVDD.n1300 0.019716
R40907 DVDD.n1530 DVDD.n1529 0.019716
R40908 DVDD.n1529 DVDD.n1299 0.019716
R40909 DVDD.n1523 DVDD.n1522 0.019716
R40910 DVDD.n1522 DVDD.n1298 0.019716
R40911 DVDD.n1518 DVDD.n1517 0.019716
R40912 DVDD.n1517 DVDD.n1297 0.019716
R40913 DVDD.n1511 DVDD.n1510 0.019716
R40914 DVDD.n1510 DVDD.n1296 0.019716
R40915 DVDD.n1506 DVDD.n1505 0.019716
R40916 DVDD.n1505 DVDD.n1295 0.019716
R40917 DVDD.n1499 DVDD.n1498 0.019716
R40918 DVDD.n1498 DVDD.n1294 0.019716
R40919 DVDD.n1494 DVDD.n1493 0.019716
R40920 DVDD.n1493 DVDD.n1293 0.019716
R40921 DVDD.n1487 DVDD.n1486 0.019716
R40922 DVDD.n1486 DVDD.n1292 0.019716
R40923 DVDD.n1482 DVDD.n1481 0.019716
R40924 DVDD.n1481 DVDD.n1291 0.019716
R40925 DVDD.n1475 DVDD.n1474 0.019716
R40926 DVDD.n1474 DVDD.n1290 0.019716
R40927 DVDD.n1470 DVDD.n1469 0.019716
R40928 DVDD.n1469 DVDD.n1289 0.019716
R40929 DVDD.n1463 DVDD.n1462 0.019716
R40930 DVDD.n1462 DVDD.n1288 0.019716
R40931 DVDD.n1458 DVDD.n1457 0.019716
R40932 DVDD.n1457 DVDD.n1287 0.019716
R40933 DVDD.n1451 DVDD.n1450 0.019716
R40934 DVDD.n1450 DVDD.n1286 0.019716
R40935 DVDD.n1446 DVDD.n1445 0.019716
R40936 DVDD.n1445 DVDD.n1285 0.019716
R40937 DVDD.n1439 DVDD.n1438 0.019716
R40938 DVDD.n1438 DVDD.n1284 0.019716
R40939 DVDD.n1434 DVDD.n1433 0.019716
R40940 DVDD.n1433 DVDD.n1283 0.019716
R40941 DVDD.n1427 DVDD.n1426 0.019716
R40942 DVDD.n1426 DVDD.n1282 0.019716
R40943 DVDD.n1422 DVDD.n1421 0.019716
R40944 DVDD.n1421 DVDD.n1281 0.019716
R40945 DVDD.n1415 DVDD.n1414 0.019716
R40946 DVDD.n1414 DVDD.n1280 0.019716
R40947 DVDD.n1410 DVDD.n1409 0.019716
R40948 DVDD.n1409 DVDD.n1279 0.019716
R40949 DVDD.n1403 DVDD.n1402 0.019716
R40950 DVDD.n1402 DVDD.n1278 0.019716
R40951 DVDD.n1398 DVDD.n1397 0.019716
R40952 DVDD.n1397 DVDD.n1277 0.019716
R40953 DVDD.n1391 DVDD.n1390 0.019716
R40954 DVDD.n1390 DVDD.n1276 0.019716
R40955 DVDD.n1386 DVDD.n1385 0.019716
R40956 DVDD.n1385 DVDD.n1275 0.019716
R40957 DVDD.n1379 DVDD.n1378 0.019716
R40958 DVDD.n1378 DVDD.n1274 0.019716
R40959 DVDD.n1374 DVDD.n1373 0.019716
R40960 DVDD.n1373 DVDD.n1273 0.019716
R40961 DVDD.n1367 DVDD.n1366 0.019716
R40962 DVDD.n1366 DVDD.n1272 0.019716
R40963 DVDD.n1362 DVDD.n1361 0.019716
R40964 DVDD.n1361 DVDD.n1271 0.019716
R40965 DVDD.n1604 DVDD.n1603 0.019716
R40966 DVDD.n1313 DVDD.n1312 0.019716
R40967 DVDD.n1596 DVDD.n1595 0.019716
R40968 DVDD.n1596 DVDD.n1311 0.019716
R40969 DVDD.n1591 DVDD.n1590 0.019716
R40970 DVDD.n1591 DVDD.n1310 0.019716
R40971 DVDD.n1584 DVDD.n1583 0.019716
R40972 DVDD.n1584 DVDD.n1309 0.019716
R40973 DVDD.n1579 DVDD.n1578 0.019716
R40974 DVDD.n1579 DVDD.n1308 0.019716
R40975 DVDD.n1572 DVDD.n1571 0.019716
R40976 DVDD.n1572 DVDD.n1307 0.019716
R40977 DVDD.n1567 DVDD.n1566 0.019716
R40978 DVDD.n1567 DVDD.n1306 0.019716
R40979 DVDD.n1560 DVDD.n1559 0.019716
R40980 DVDD.n1560 DVDD.n1305 0.019716
R40981 DVDD.n1555 DVDD.n1554 0.019716
R40982 DVDD.n1555 DVDD.n1304 0.019716
R40983 DVDD.n1548 DVDD.n1547 0.019716
R40984 DVDD.n1548 DVDD.n1303 0.019716
R40985 DVDD.n1543 DVDD.n1542 0.019716
R40986 DVDD.n1543 DVDD.n1302 0.019716
R40987 DVDD.n1536 DVDD.n1535 0.019716
R40988 DVDD.n1536 DVDD.n1301 0.019716
R40989 DVDD.n1531 DVDD.n1530 0.019716
R40990 DVDD.n1531 DVDD.n1300 0.019716
R40991 DVDD.n1524 DVDD.n1523 0.019716
R40992 DVDD.n1524 DVDD.n1299 0.019716
R40993 DVDD.n1519 DVDD.n1518 0.019716
R40994 DVDD.n1519 DVDD.n1298 0.019716
R40995 DVDD.n1512 DVDD.n1511 0.019716
R40996 DVDD.n1512 DVDD.n1297 0.019716
R40997 DVDD.n1507 DVDD.n1506 0.019716
R40998 DVDD.n1507 DVDD.n1296 0.019716
R40999 DVDD.n1500 DVDD.n1499 0.019716
R41000 DVDD.n1500 DVDD.n1295 0.019716
R41001 DVDD.n1495 DVDD.n1494 0.019716
R41002 DVDD.n1495 DVDD.n1294 0.019716
R41003 DVDD.n1488 DVDD.n1487 0.019716
R41004 DVDD.n1488 DVDD.n1293 0.019716
R41005 DVDD.n1483 DVDD.n1482 0.019716
R41006 DVDD.n1483 DVDD.n1292 0.019716
R41007 DVDD.n1476 DVDD.n1475 0.019716
R41008 DVDD.n1476 DVDD.n1291 0.019716
R41009 DVDD.n1471 DVDD.n1470 0.019716
R41010 DVDD.n1471 DVDD.n1290 0.019716
R41011 DVDD.n1464 DVDD.n1463 0.019716
R41012 DVDD.n1464 DVDD.n1289 0.019716
R41013 DVDD.n1459 DVDD.n1458 0.019716
R41014 DVDD.n1459 DVDD.n1288 0.019716
R41015 DVDD.n1452 DVDD.n1451 0.019716
R41016 DVDD.n1452 DVDD.n1287 0.019716
R41017 DVDD.n1447 DVDD.n1446 0.019716
R41018 DVDD.n1447 DVDD.n1286 0.019716
R41019 DVDD.n1440 DVDD.n1439 0.019716
R41020 DVDD.n1440 DVDD.n1285 0.019716
R41021 DVDD.n1435 DVDD.n1434 0.019716
R41022 DVDD.n1435 DVDD.n1284 0.019716
R41023 DVDD.n1428 DVDD.n1427 0.019716
R41024 DVDD.n1428 DVDD.n1283 0.019716
R41025 DVDD.n1423 DVDD.n1422 0.019716
R41026 DVDD.n1423 DVDD.n1282 0.019716
R41027 DVDD.n1416 DVDD.n1415 0.019716
R41028 DVDD.n1416 DVDD.n1281 0.019716
R41029 DVDD.n1411 DVDD.n1410 0.019716
R41030 DVDD.n1411 DVDD.n1280 0.019716
R41031 DVDD.n1404 DVDD.n1403 0.019716
R41032 DVDD.n1404 DVDD.n1279 0.019716
R41033 DVDD.n1399 DVDD.n1398 0.019716
R41034 DVDD.n1399 DVDD.n1278 0.019716
R41035 DVDD.n1392 DVDD.n1391 0.019716
R41036 DVDD.n1392 DVDD.n1277 0.019716
R41037 DVDD.n1387 DVDD.n1386 0.019716
R41038 DVDD.n1387 DVDD.n1276 0.019716
R41039 DVDD.n1380 DVDD.n1379 0.019716
R41040 DVDD.n1380 DVDD.n1275 0.019716
R41041 DVDD.n1375 DVDD.n1374 0.019716
R41042 DVDD.n1375 DVDD.n1274 0.019716
R41043 DVDD.n1368 DVDD.n1367 0.019716
R41044 DVDD.n1368 DVDD.n1273 0.019716
R41045 DVDD.n1363 DVDD.n1362 0.019716
R41046 DVDD.n1363 DVDD.n1272 0.019716
R41047 DVDD.n1356 DVDD.n1271 0.019716
R41048 DVDD.n1699 DVDD.n1653 0.019716
R41049 DVDD.n1700 DVDD.n1652 0.019716
R41050 DVDD.n17020 DVDD.n1651 0.019716
R41051 DVDD.n17020 DVDD.n17019 0.019716
R41052 DVDD.n17022 DVDD.n1650 0.019716
R41053 DVDD.n17023 DVDD.n17022 0.019716
R41054 DVDD.n17032 DVDD.n1649 0.019716
R41055 DVDD.n17032 DVDD.n17031 0.019716
R41056 DVDD.n17034 DVDD.n1648 0.019716
R41057 DVDD.n17035 DVDD.n17034 0.019716
R41058 DVDD.n17044 DVDD.n1647 0.019716
R41059 DVDD.n17044 DVDD.n17043 0.019716
R41060 DVDD.n17046 DVDD.n1646 0.019716
R41061 DVDD.n17047 DVDD.n17046 0.019716
R41062 DVDD.n17056 DVDD.n1645 0.019716
R41063 DVDD.n17056 DVDD.n17055 0.019716
R41064 DVDD.n17058 DVDD.n1644 0.019716
R41065 DVDD.n17059 DVDD.n17058 0.019716
R41066 DVDD.n17068 DVDD.n1643 0.019716
R41067 DVDD.n17068 DVDD.n17067 0.019716
R41068 DVDD.n17070 DVDD.n1642 0.019716
R41069 DVDD.n17071 DVDD.n17070 0.019716
R41070 DVDD.n17080 DVDD.n1641 0.019716
R41071 DVDD.n17080 DVDD.n17079 0.019716
R41072 DVDD.n17082 DVDD.n1640 0.019716
R41073 DVDD.n17083 DVDD.n17082 0.019716
R41074 DVDD.n17092 DVDD.n1639 0.019716
R41075 DVDD.n17092 DVDD.n17091 0.019716
R41076 DVDD.n17094 DVDD.n1638 0.019716
R41077 DVDD.n17095 DVDD.n17094 0.019716
R41078 DVDD.n17104 DVDD.n1637 0.019716
R41079 DVDD.n17104 DVDD.n17103 0.019716
R41080 DVDD.n17106 DVDD.n1636 0.019716
R41081 DVDD.n17107 DVDD.n17106 0.019716
R41082 DVDD.n17116 DVDD.n1635 0.019716
R41083 DVDD.n17116 DVDD.n17115 0.019716
R41084 DVDD.n17118 DVDD.n1634 0.019716
R41085 DVDD.n17119 DVDD.n17118 0.019716
R41086 DVDD.n17128 DVDD.n1633 0.019716
R41087 DVDD.n17128 DVDD.n17127 0.019716
R41088 DVDD.n17130 DVDD.n1632 0.019716
R41089 DVDD.n17131 DVDD.n17130 0.019716
R41090 DVDD.n17140 DVDD.n1631 0.019716
R41091 DVDD.n17140 DVDD.n17139 0.019716
R41092 DVDD.n17142 DVDD.n1630 0.019716
R41093 DVDD.n17143 DVDD.n17142 0.019716
R41094 DVDD.n17152 DVDD.n1629 0.019716
R41095 DVDD.n17152 DVDD.n17151 0.019716
R41096 DVDD.n17154 DVDD.n1628 0.019716
R41097 DVDD.n17155 DVDD.n17154 0.019716
R41098 DVDD.n17164 DVDD.n1627 0.019716
R41099 DVDD.n17164 DVDD.n17163 0.019716
R41100 DVDD.n17166 DVDD.n1626 0.019716
R41101 DVDD.n17167 DVDD.n17166 0.019716
R41102 DVDD.n17176 DVDD.n1625 0.019716
R41103 DVDD.n17176 DVDD.n17175 0.019716
R41104 DVDD.n17178 DVDD.n1624 0.019716
R41105 DVDD.n17179 DVDD.n17178 0.019716
R41106 DVDD.n17188 DVDD.n1623 0.019716
R41107 DVDD.n17188 DVDD.n17187 0.019716
R41108 DVDD.n17190 DVDD.n1622 0.019716
R41109 DVDD.n17191 DVDD.n17190 0.019716
R41110 DVDD.n17200 DVDD.n1621 0.019716
R41111 DVDD.n17200 DVDD.n17199 0.019716
R41112 DVDD.n17202 DVDD.n1620 0.019716
R41113 DVDD.n17203 DVDD.n17202 0.019716
R41114 DVDD.n17212 DVDD.n1619 0.019716
R41115 DVDD.n17212 DVDD.n17211 0.019716
R41116 DVDD.n17214 DVDD.n1618 0.019716
R41117 DVDD.n17215 DVDD.n17214 0.019716
R41118 DVDD.n17224 DVDD.n1617 0.019716
R41119 DVDD.n17224 DVDD.n17223 0.019716
R41120 DVDD.n17226 DVDD.n1616 0.019716
R41121 DVDD.n17227 DVDD.n17226 0.019716
R41122 DVDD.n17236 DVDD.n1615 0.019716
R41123 DVDD.n17236 DVDD.n17235 0.019716
R41124 DVDD.n17238 DVDD.n1614 0.019716
R41125 DVDD.n17239 DVDD.n17238 0.019716
R41126 DVDD.n17248 DVDD.n1613 0.019716
R41127 DVDD.n17248 DVDD.n17247 0.019716
R41128 DVDD.n17250 DVDD.n1612 0.019716
R41129 DVDD.n17251 DVDD.n17250 0.019716
R41130 DVDD.n17261 DVDD.n17260 0.019716
R41131 DVDD.n1798 DVDD.n1754 0.019716
R41132 DVDD.n1799 DVDD.n1753 0.019716
R41133 DVDD.n16752 DVDD.n1752 0.019716
R41134 DVDD.n16752 DVDD.n16751 0.019716
R41135 DVDD.n16754 DVDD.n1751 0.019716
R41136 DVDD.n16755 DVDD.n16754 0.019716
R41137 DVDD.n16764 DVDD.n1750 0.019716
R41138 DVDD.n16764 DVDD.n16763 0.019716
R41139 DVDD.n16766 DVDD.n1749 0.019716
R41140 DVDD.n16767 DVDD.n16766 0.019716
R41141 DVDD.n16776 DVDD.n1748 0.019716
R41142 DVDD.n16776 DVDD.n16775 0.019716
R41143 DVDD.n16778 DVDD.n1747 0.019716
R41144 DVDD.n16779 DVDD.n16778 0.019716
R41145 DVDD.n16788 DVDD.n1746 0.019716
R41146 DVDD.n16788 DVDD.n16787 0.019716
R41147 DVDD.n16790 DVDD.n1745 0.019716
R41148 DVDD.n16791 DVDD.n16790 0.019716
R41149 DVDD.n16800 DVDD.n1744 0.019716
R41150 DVDD.n16800 DVDD.n16799 0.019716
R41151 DVDD.n16802 DVDD.n1743 0.019716
R41152 DVDD.n16803 DVDD.n16802 0.019716
R41153 DVDD.n16812 DVDD.n1742 0.019716
R41154 DVDD.n16812 DVDD.n16811 0.019716
R41155 DVDD.n16814 DVDD.n1741 0.019716
R41156 DVDD.n16815 DVDD.n16814 0.019716
R41157 DVDD.n16824 DVDD.n1740 0.019716
R41158 DVDD.n16824 DVDD.n16823 0.019716
R41159 DVDD.n16826 DVDD.n1739 0.019716
R41160 DVDD.n16827 DVDD.n16826 0.019716
R41161 DVDD.n16836 DVDD.n1738 0.019716
R41162 DVDD.n16836 DVDD.n16835 0.019716
R41163 DVDD.n16838 DVDD.n1737 0.019716
R41164 DVDD.n16839 DVDD.n16838 0.019716
R41165 DVDD.n16848 DVDD.n1736 0.019716
R41166 DVDD.n16848 DVDD.n16847 0.019716
R41167 DVDD.n16850 DVDD.n1735 0.019716
R41168 DVDD.n16851 DVDD.n16850 0.019716
R41169 DVDD.n16860 DVDD.n1734 0.019716
R41170 DVDD.n16860 DVDD.n16859 0.019716
R41171 DVDD.n16862 DVDD.n1733 0.019716
R41172 DVDD.n16863 DVDD.n16862 0.019716
R41173 DVDD.n16872 DVDD.n1732 0.019716
R41174 DVDD.n16872 DVDD.n16871 0.019716
R41175 DVDD.n16874 DVDD.n1731 0.019716
R41176 DVDD.n16875 DVDD.n16874 0.019716
R41177 DVDD.n16884 DVDD.n1730 0.019716
R41178 DVDD.n16884 DVDD.n16883 0.019716
R41179 DVDD.n16886 DVDD.n1729 0.019716
R41180 DVDD.n16887 DVDD.n16886 0.019716
R41181 DVDD.n16896 DVDD.n1728 0.019716
R41182 DVDD.n16896 DVDD.n16895 0.019716
R41183 DVDD.n16898 DVDD.n1727 0.019716
R41184 DVDD.n16899 DVDD.n16898 0.019716
R41185 DVDD.n16908 DVDD.n1726 0.019716
R41186 DVDD.n16908 DVDD.n16907 0.019716
R41187 DVDD.n16910 DVDD.n1725 0.019716
R41188 DVDD.n16911 DVDD.n16910 0.019716
R41189 DVDD.n16920 DVDD.n1724 0.019716
R41190 DVDD.n16920 DVDD.n16919 0.019716
R41191 DVDD.n16922 DVDD.n1723 0.019716
R41192 DVDD.n16923 DVDD.n16922 0.019716
R41193 DVDD.n16932 DVDD.n1722 0.019716
R41194 DVDD.n16932 DVDD.n16931 0.019716
R41195 DVDD.n16934 DVDD.n1721 0.019716
R41196 DVDD.n16935 DVDD.n16934 0.019716
R41197 DVDD.n16944 DVDD.n1720 0.019716
R41198 DVDD.n16944 DVDD.n16943 0.019716
R41199 DVDD.n16946 DVDD.n1719 0.019716
R41200 DVDD.n16947 DVDD.n16946 0.019716
R41201 DVDD.n16956 DVDD.n1718 0.019716
R41202 DVDD.n16956 DVDD.n16955 0.019716
R41203 DVDD.n16958 DVDD.n1717 0.019716
R41204 DVDD.n16959 DVDD.n16958 0.019716
R41205 DVDD.n16968 DVDD.n1716 0.019716
R41206 DVDD.n16968 DVDD.n16967 0.019716
R41207 DVDD.n16970 DVDD.n1715 0.019716
R41208 DVDD.n16971 DVDD.n16970 0.019716
R41209 DVDD.n16980 DVDD.n1714 0.019716
R41210 DVDD.n16980 DVDD.n16979 0.019716
R41211 DVDD.n16982 DVDD.n1713 0.019716
R41212 DVDD.n16983 DVDD.n16982 0.019716
R41213 DVDD.n16993 DVDD.n16992 0.019716
R41214 DVDD.n2155 DVDD.n2154 0.019716
R41215 DVDD.n1864 DVDD.n1863 0.019716
R41216 DVDD.n2147 DVDD.n2146 0.019716
R41217 DVDD.n2147 DVDD.n1862 0.019716
R41218 DVDD.n2142 DVDD.n2141 0.019716
R41219 DVDD.n2142 DVDD.n1861 0.019716
R41220 DVDD.n2135 DVDD.n2134 0.019716
R41221 DVDD.n2135 DVDD.n1860 0.019716
R41222 DVDD.n2130 DVDD.n2129 0.019716
R41223 DVDD.n2130 DVDD.n1859 0.019716
R41224 DVDD.n2123 DVDD.n2122 0.019716
R41225 DVDD.n2123 DVDD.n1858 0.019716
R41226 DVDD.n2118 DVDD.n2117 0.019716
R41227 DVDD.n2118 DVDD.n1857 0.019716
R41228 DVDD.n2111 DVDD.n2110 0.019716
R41229 DVDD.n2111 DVDD.n1856 0.019716
R41230 DVDD.n2106 DVDD.n2105 0.019716
R41231 DVDD.n2106 DVDD.n1855 0.019716
R41232 DVDD.n2099 DVDD.n2098 0.019716
R41233 DVDD.n2099 DVDD.n1854 0.019716
R41234 DVDD.n2094 DVDD.n2093 0.019716
R41235 DVDD.n2094 DVDD.n1853 0.019716
R41236 DVDD.n2087 DVDD.n2086 0.019716
R41237 DVDD.n2087 DVDD.n1852 0.019716
R41238 DVDD.n2082 DVDD.n2081 0.019716
R41239 DVDD.n2082 DVDD.n1851 0.019716
R41240 DVDD.n2075 DVDD.n2074 0.019716
R41241 DVDD.n2075 DVDD.n1850 0.019716
R41242 DVDD.n2070 DVDD.n2069 0.019716
R41243 DVDD.n2070 DVDD.n1849 0.019716
R41244 DVDD.n2063 DVDD.n2062 0.019716
R41245 DVDD.n2063 DVDD.n1848 0.019716
R41246 DVDD.n2058 DVDD.n2057 0.019716
R41247 DVDD.n2058 DVDD.n1847 0.019716
R41248 DVDD.n2051 DVDD.n2050 0.019716
R41249 DVDD.n2051 DVDD.n1846 0.019716
R41250 DVDD.n2046 DVDD.n2045 0.019716
R41251 DVDD.n2046 DVDD.n1845 0.019716
R41252 DVDD.n2039 DVDD.n2038 0.019716
R41253 DVDD.n2039 DVDD.n1844 0.019716
R41254 DVDD.n2034 DVDD.n2033 0.019716
R41255 DVDD.n2034 DVDD.n1843 0.019716
R41256 DVDD.n2027 DVDD.n2026 0.019716
R41257 DVDD.n2027 DVDD.n1842 0.019716
R41258 DVDD.n2022 DVDD.n2021 0.019716
R41259 DVDD.n2022 DVDD.n1841 0.019716
R41260 DVDD.n2015 DVDD.n2014 0.019716
R41261 DVDD.n2015 DVDD.n1840 0.019716
R41262 DVDD.n2010 DVDD.n2009 0.019716
R41263 DVDD.n2010 DVDD.n1839 0.019716
R41264 DVDD.n2003 DVDD.n2002 0.019716
R41265 DVDD.n2003 DVDD.n1838 0.019716
R41266 DVDD.n1998 DVDD.n1997 0.019716
R41267 DVDD.n1998 DVDD.n1837 0.019716
R41268 DVDD.n1991 DVDD.n1990 0.019716
R41269 DVDD.n1991 DVDD.n1836 0.019716
R41270 DVDD.n1986 DVDD.n1985 0.019716
R41271 DVDD.n1986 DVDD.n1835 0.019716
R41272 DVDD.n1979 DVDD.n1978 0.019716
R41273 DVDD.n1979 DVDD.n1834 0.019716
R41274 DVDD.n1974 DVDD.n1973 0.019716
R41275 DVDD.n1974 DVDD.n1833 0.019716
R41276 DVDD.n1967 DVDD.n1966 0.019716
R41277 DVDD.n1967 DVDD.n1832 0.019716
R41278 DVDD.n1962 DVDD.n1961 0.019716
R41279 DVDD.n1962 DVDD.n1831 0.019716
R41280 DVDD.n1955 DVDD.n1954 0.019716
R41281 DVDD.n1955 DVDD.n1830 0.019716
R41282 DVDD.n1950 DVDD.n1949 0.019716
R41283 DVDD.n1950 DVDD.n1829 0.019716
R41284 DVDD.n1943 DVDD.n1942 0.019716
R41285 DVDD.n1943 DVDD.n1828 0.019716
R41286 DVDD.n1938 DVDD.n1937 0.019716
R41287 DVDD.n1938 DVDD.n1827 0.019716
R41288 DVDD.n1931 DVDD.n1930 0.019716
R41289 DVDD.n1931 DVDD.n1826 0.019716
R41290 DVDD.n1926 DVDD.n1925 0.019716
R41291 DVDD.n1926 DVDD.n1825 0.019716
R41292 DVDD.n1919 DVDD.n1918 0.019716
R41293 DVDD.n1919 DVDD.n1824 0.019716
R41294 DVDD.n1914 DVDD.n1913 0.019716
R41295 DVDD.n1914 DVDD.n1823 0.019716
R41296 DVDD.n1907 DVDD.n1822 0.019716
R41297 DVDD.n2251 DVDD.n2207 0.019716
R41298 DVDD.n2252 DVDD.n2206 0.019716
R41299 DVDD.n16463 DVDD.n2205 0.019716
R41300 DVDD.n16463 DVDD.n16462 0.019716
R41301 DVDD.n16465 DVDD.n2204 0.019716
R41302 DVDD.n16466 DVDD.n16465 0.019716
R41303 DVDD.n16475 DVDD.n2203 0.019716
R41304 DVDD.n16475 DVDD.n16474 0.019716
R41305 DVDD.n16477 DVDD.n2202 0.019716
R41306 DVDD.n16478 DVDD.n16477 0.019716
R41307 DVDD.n16487 DVDD.n2201 0.019716
R41308 DVDD.n16487 DVDD.n16486 0.019716
R41309 DVDD.n16489 DVDD.n2200 0.019716
R41310 DVDD.n16490 DVDD.n16489 0.019716
R41311 DVDD.n16499 DVDD.n2199 0.019716
R41312 DVDD.n16499 DVDD.n16498 0.019716
R41313 DVDD.n16501 DVDD.n2198 0.019716
R41314 DVDD.n16502 DVDD.n16501 0.019716
R41315 DVDD.n16511 DVDD.n2197 0.019716
R41316 DVDD.n16511 DVDD.n16510 0.019716
R41317 DVDD.n16513 DVDD.n2196 0.019716
R41318 DVDD.n16514 DVDD.n16513 0.019716
R41319 DVDD.n16523 DVDD.n2195 0.019716
R41320 DVDD.n16523 DVDD.n16522 0.019716
R41321 DVDD.n16525 DVDD.n2194 0.019716
R41322 DVDD.n16526 DVDD.n16525 0.019716
R41323 DVDD.n16535 DVDD.n2193 0.019716
R41324 DVDD.n16535 DVDD.n16534 0.019716
R41325 DVDD.n16537 DVDD.n2192 0.019716
R41326 DVDD.n16538 DVDD.n16537 0.019716
R41327 DVDD.n16547 DVDD.n2191 0.019716
R41328 DVDD.n16547 DVDD.n16546 0.019716
R41329 DVDD.n16549 DVDD.n2190 0.019716
R41330 DVDD.n16550 DVDD.n16549 0.019716
R41331 DVDD.n16559 DVDD.n2189 0.019716
R41332 DVDD.n16559 DVDD.n16558 0.019716
R41333 DVDD.n16561 DVDD.n2188 0.019716
R41334 DVDD.n16562 DVDD.n16561 0.019716
R41335 DVDD.n16571 DVDD.n2187 0.019716
R41336 DVDD.n16571 DVDD.n16570 0.019716
R41337 DVDD.n16573 DVDD.n2186 0.019716
R41338 DVDD.n16574 DVDD.n16573 0.019716
R41339 DVDD.n16583 DVDD.n2185 0.019716
R41340 DVDD.n16583 DVDD.n16582 0.019716
R41341 DVDD.n16585 DVDD.n2184 0.019716
R41342 DVDD.n16586 DVDD.n16585 0.019716
R41343 DVDD.n16595 DVDD.n2183 0.019716
R41344 DVDD.n16595 DVDD.n16594 0.019716
R41345 DVDD.n16597 DVDD.n2182 0.019716
R41346 DVDD.n16598 DVDD.n16597 0.019716
R41347 DVDD.n16607 DVDD.n2181 0.019716
R41348 DVDD.n16607 DVDD.n16606 0.019716
R41349 DVDD.n16609 DVDD.n2180 0.019716
R41350 DVDD.n16610 DVDD.n16609 0.019716
R41351 DVDD.n16619 DVDD.n2179 0.019716
R41352 DVDD.n16619 DVDD.n16618 0.019716
R41353 DVDD.n16621 DVDD.n2178 0.019716
R41354 DVDD.n16622 DVDD.n16621 0.019716
R41355 DVDD.n16631 DVDD.n2177 0.019716
R41356 DVDD.n16631 DVDD.n16630 0.019716
R41357 DVDD.n16633 DVDD.n2176 0.019716
R41358 DVDD.n16634 DVDD.n16633 0.019716
R41359 DVDD.n16643 DVDD.n2175 0.019716
R41360 DVDD.n16643 DVDD.n16642 0.019716
R41361 DVDD.n16645 DVDD.n2174 0.019716
R41362 DVDD.n16646 DVDD.n16645 0.019716
R41363 DVDD.n16655 DVDD.n2173 0.019716
R41364 DVDD.n16655 DVDD.n16654 0.019716
R41365 DVDD.n16657 DVDD.n2172 0.019716
R41366 DVDD.n16658 DVDD.n16657 0.019716
R41367 DVDD.n16667 DVDD.n2171 0.019716
R41368 DVDD.n16667 DVDD.n16666 0.019716
R41369 DVDD.n16669 DVDD.n2170 0.019716
R41370 DVDD.n16670 DVDD.n16669 0.019716
R41371 DVDD.n16679 DVDD.n2169 0.019716
R41372 DVDD.n16679 DVDD.n16678 0.019716
R41373 DVDD.n16681 DVDD.n2168 0.019716
R41374 DVDD.n16682 DVDD.n16681 0.019716
R41375 DVDD.n16691 DVDD.n2167 0.019716
R41376 DVDD.n16691 DVDD.n16690 0.019716
R41377 DVDD.n16693 DVDD.n2166 0.019716
R41378 DVDD.n16694 DVDD.n16693 0.019716
R41379 DVDD.n16703 DVDD.n16702 0.019716
R41380 DVDD.n13255 DVDD.n13254 0.019716
R41381 DVDD.n12965 DVDD.n12964 0.019716
R41382 DVDD.n13247 DVDD.n13246 0.019716
R41383 DVDD.n13247 DVDD.n12963 0.019716
R41384 DVDD.n13242 DVDD.n13241 0.019716
R41385 DVDD.n13242 DVDD.n12962 0.019716
R41386 DVDD.n13235 DVDD.n13234 0.019716
R41387 DVDD.n13235 DVDD.n12961 0.019716
R41388 DVDD.n13230 DVDD.n13229 0.019716
R41389 DVDD.n13230 DVDD.n12960 0.019716
R41390 DVDD.n13223 DVDD.n13222 0.019716
R41391 DVDD.n13223 DVDD.n12959 0.019716
R41392 DVDD.n13218 DVDD.n13217 0.019716
R41393 DVDD.n13218 DVDD.n12958 0.019716
R41394 DVDD.n13211 DVDD.n13210 0.019716
R41395 DVDD.n13211 DVDD.n12957 0.019716
R41396 DVDD.n13206 DVDD.n13205 0.019716
R41397 DVDD.n13206 DVDD.n12956 0.019716
R41398 DVDD.n13199 DVDD.n13198 0.019716
R41399 DVDD.n13199 DVDD.n12955 0.019716
R41400 DVDD.n13194 DVDD.n13193 0.019716
R41401 DVDD.n13194 DVDD.n12954 0.019716
R41402 DVDD.n13187 DVDD.n13186 0.019716
R41403 DVDD.n13187 DVDD.n12953 0.019716
R41404 DVDD.n13182 DVDD.n13181 0.019716
R41405 DVDD.n13182 DVDD.n12952 0.019716
R41406 DVDD.n13175 DVDD.n13174 0.019716
R41407 DVDD.n13175 DVDD.n12951 0.019716
R41408 DVDD.n13170 DVDD.n13169 0.019716
R41409 DVDD.n13170 DVDD.n12950 0.019716
R41410 DVDD.n13163 DVDD.n13162 0.019716
R41411 DVDD.n13163 DVDD.n12949 0.019716
R41412 DVDD.n13158 DVDD.n13157 0.019716
R41413 DVDD.n13158 DVDD.n12948 0.019716
R41414 DVDD.n13151 DVDD.n13150 0.019716
R41415 DVDD.n13151 DVDD.n12947 0.019716
R41416 DVDD.n13146 DVDD.n13145 0.019716
R41417 DVDD.n13146 DVDD.n12946 0.019716
R41418 DVDD.n13139 DVDD.n13138 0.019716
R41419 DVDD.n13139 DVDD.n12945 0.019716
R41420 DVDD.n13134 DVDD.n13133 0.019716
R41421 DVDD.n13134 DVDD.n12944 0.019716
R41422 DVDD.n13127 DVDD.n13126 0.019716
R41423 DVDD.n13127 DVDD.n12943 0.019716
R41424 DVDD.n13122 DVDD.n13121 0.019716
R41425 DVDD.n13122 DVDD.n12942 0.019716
R41426 DVDD.n13115 DVDD.n13114 0.019716
R41427 DVDD.n13115 DVDD.n12941 0.019716
R41428 DVDD.n13110 DVDD.n13109 0.019716
R41429 DVDD.n13110 DVDD.n12940 0.019716
R41430 DVDD.n13103 DVDD.n13102 0.019716
R41431 DVDD.n13103 DVDD.n12939 0.019716
R41432 DVDD.n13098 DVDD.n13097 0.019716
R41433 DVDD.n13098 DVDD.n12938 0.019716
R41434 DVDD.n13091 DVDD.n13090 0.019716
R41435 DVDD.n13091 DVDD.n12937 0.019716
R41436 DVDD.n13086 DVDD.n13085 0.019716
R41437 DVDD.n13086 DVDD.n12936 0.019716
R41438 DVDD.n13079 DVDD.n13078 0.019716
R41439 DVDD.n13079 DVDD.n12935 0.019716
R41440 DVDD.n13074 DVDD.n13073 0.019716
R41441 DVDD.n13074 DVDD.n12934 0.019716
R41442 DVDD.n13067 DVDD.n13066 0.019716
R41443 DVDD.n13067 DVDD.n12933 0.019716
R41444 DVDD.n13062 DVDD.n13061 0.019716
R41445 DVDD.n13062 DVDD.n12932 0.019716
R41446 DVDD.n13055 DVDD.n13054 0.019716
R41447 DVDD.n13055 DVDD.n12931 0.019716
R41448 DVDD.n13050 DVDD.n13049 0.019716
R41449 DVDD.n13050 DVDD.n12930 0.019716
R41450 DVDD.n13043 DVDD.n13042 0.019716
R41451 DVDD.n13043 DVDD.n12929 0.019716
R41452 DVDD.n13038 DVDD.n13037 0.019716
R41453 DVDD.n13038 DVDD.n12928 0.019716
R41454 DVDD.n13031 DVDD.n13030 0.019716
R41455 DVDD.n13031 DVDD.n12927 0.019716
R41456 DVDD.n13026 DVDD.n13025 0.019716
R41457 DVDD.n13026 DVDD.n12926 0.019716
R41458 DVDD.n13019 DVDD.n13018 0.019716
R41459 DVDD.n13019 DVDD.n12925 0.019716
R41460 DVDD.n13014 DVDD.n13013 0.019716
R41461 DVDD.n13014 DVDD.n12924 0.019716
R41462 DVDD.n13007 DVDD.n12923 0.019716
R41463 DVDD.n13472 DVDD.n13471 0.019716
R41464 DVDD.n12824 DVDD.n12780 0.019716
R41465 DVDD.n13288 DVDD.n12823 0.019716
R41466 DVDD.n13288 DVDD.n12778 0.019716
R41467 DVDD.n13292 DVDD.n12822 0.019716
R41468 DVDD.n13292 DVDD.n12777 0.019716
R41469 DVDD.n13297 DVDD.n12821 0.019716
R41470 DVDD.n13297 DVDD.n12776 0.019716
R41471 DVDD.n13301 DVDD.n12820 0.019716
R41472 DVDD.n13301 DVDD.n12775 0.019716
R41473 DVDD.n13306 DVDD.n12819 0.019716
R41474 DVDD.n13306 DVDD.n12774 0.019716
R41475 DVDD.n13310 DVDD.n12818 0.019716
R41476 DVDD.n13310 DVDD.n12773 0.019716
R41477 DVDD.n13315 DVDD.n12817 0.019716
R41478 DVDD.n13315 DVDD.n12772 0.019716
R41479 DVDD.n13319 DVDD.n12816 0.019716
R41480 DVDD.n13319 DVDD.n12771 0.019716
R41481 DVDD.n13324 DVDD.n12815 0.019716
R41482 DVDD.n13324 DVDD.n12770 0.019716
R41483 DVDD.n13328 DVDD.n12814 0.019716
R41484 DVDD.n13328 DVDD.n12769 0.019716
R41485 DVDD.n13333 DVDD.n12813 0.019716
R41486 DVDD.n13333 DVDD.n12768 0.019716
R41487 DVDD.n13337 DVDD.n12812 0.019716
R41488 DVDD.n13337 DVDD.n12767 0.019716
R41489 DVDD.n13342 DVDD.n12811 0.019716
R41490 DVDD.n13342 DVDD.n12766 0.019716
R41491 DVDD.n13346 DVDD.n12810 0.019716
R41492 DVDD.n13346 DVDD.n12765 0.019716
R41493 DVDD.n13351 DVDD.n12809 0.019716
R41494 DVDD.n13351 DVDD.n12764 0.019716
R41495 DVDD.n13355 DVDD.n12808 0.019716
R41496 DVDD.n13355 DVDD.n12763 0.019716
R41497 DVDD.n13360 DVDD.n12807 0.019716
R41498 DVDD.n13360 DVDD.n12762 0.019716
R41499 DVDD.n13364 DVDD.n12806 0.019716
R41500 DVDD.n13364 DVDD.n12761 0.019716
R41501 DVDD.n13369 DVDD.n12805 0.019716
R41502 DVDD.n13369 DVDD.n12760 0.019716
R41503 DVDD.n13373 DVDD.n12804 0.019716
R41504 DVDD.n13373 DVDD.n12759 0.019716
R41505 DVDD.n13378 DVDD.n12803 0.019716
R41506 DVDD.n13378 DVDD.n12758 0.019716
R41507 DVDD.n13382 DVDD.n12802 0.019716
R41508 DVDD.n13382 DVDD.n12757 0.019716
R41509 DVDD.n13387 DVDD.n12801 0.019716
R41510 DVDD.n13387 DVDD.n12756 0.019716
R41511 DVDD.n13391 DVDD.n12800 0.019716
R41512 DVDD.n13391 DVDD.n12755 0.019716
R41513 DVDD.n13396 DVDD.n12799 0.019716
R41514 DVDD.n13396 DVDD.n12754 0.019716
R41515 DVDD.n13400 DVDD.n12798 0.019716
R41516 DVDD.n13400 DVDD.n12753 0.019716
R41517 DVDD.n13405 DVDD.n12797 0.019716
R41518 DVDD.n13405 DVDD.n12752 0.019716
R41519 DVDD.n13409 DVDD.n12796 0.019716
R41520 DVDD.n13409 DVDD.n12751 0.019716
R41521 DVDD.n13414 DVDD.n12795 0.019716
R41522 DVDD.n13414 DVDD.n12750 0.019716
R41523 DVDD.n13418 DVDD.n12794 0.019716
R41524 DVDD.n13418 DVDD.n12749 0.019716
R41525 DVDD.n13423 DVDD.n12793 0.019716
R41526 DVDD.n13423 DVDD.n12748 0.019716
R41527 DVDD.n13427 DVDD.n12792 0.019716
R41528 DVDD.n13427 DVDD.n12747 0.019716
R41529 DVDD.n13432 DVDD.n12791 0.019716
R41530 DVDD.n13432 DVDD.n12746 0.019716
R41531 DVDD.n13436 DVDD.n12790 0.019716
R41532 DVDD.n13436 DVDD.n12745 0.019716
R41533 DVDD.n13441 DVDD.n12789 0.019716
R41534 DVDD.n13441 DVDD.n12744 0.019716
R41535 DVDD.n13445 DVDD.n12788 0.019716
R41536 DVDD.n13445 DVDD.n12743 0.019716
R41537 DVDD.n13450 DVDD.n12787 0.019716
R41538 DVDD.n13450 DVDD.n12742 0.019716
R41539 DVDD.n13454 DVDD.n12786 0.019716
R41540 DVDD.n13454 DVDD.n12741 0.019716
R41541 DVDD.n13459 DVDD.n12785 0.019716
R41542 DVDD.n13459 DVDD.n12740 0.019716
R41543 DVDD.n13463 DVDD.n12784 0.019716
R41544 DVDD.n13463 DVDD.n12739 0.019716
R41545 DVDD.n13469 DVDD.n12738 0.019716
R41546 DVDD.n13486 DVDD.n13485 0.019716
R41547 DVDD.n12476 DVDD.n12433 0.019716
R41548 DVDD.n12546 DVDD.n12475 0.019716
R41549 DVDD.n12546 DVDD.n12431 0.019716
R41550 DVDD.n12550 DVDD.n12474 0.019716
R41551 DVDD.n12550 DVDD.n12430 0.019716
R41552 DVDD.n12555 DVDD.n12473 0.019716
R41553 DVDD.n12555 DVDD.n12429 0.019716
R41554 DVDD.n12559 DVDD.n12472 0.019716
R41555 DVDD.n12559 DVDD.n12428 0.019716
R41556 DVDD.n12564 DVDD.n12471 0.019716
R41557 DVDD.n12564 DVDD.n12427 0.019716
R41558 DVDD.n12568 DVDD.n12470 0.019716
R41559 DVDD.n12568 DVDD.n12426 0.019716
R41560 DVDD.n12573 DVDD.n12469 0.019716
R41561 DVDD.n12573 DVDD.n12425 0.019716
R41562 DVDD.n12577 DVDD.n12468 0.019716
R41563 DVDD.n12577 DVDD.n12424 0.019716
R41564 DVDD.n12582 DVDD.n12467 0.019716
R41565 DVDD.n12582 DVDD.n12423 0.019716
R41566 DVDD.n12586 DVDD.n12466 0.019716
R41567 DVDD.n12586 DVDD.n12422 0.019716
R41568 DVDD.n12591 DVDD.n12465 0.019716
R41569 DVDD.n12591 DVDD.n12421 0.019716
R41570 DVDD.n12595 DVDD.n12464 0.019716
R41571 DVDD.n12595 DVDD.n12420 0.019716
R41572 DVDD.n12600 DVDD.n12463 0.019716
R41573 DVDD.n12600 DVDD.n12419 0.019716
R41574 DVDD.n12604 DVDD.n12462 0.019716
R41575 DVDD.n12604 DVDD.n12418 0.019716
R41576 DVDD.n12609 DVDD.n12461 0.019716
R41577 DVDD.n12609 DVDD.n12417 0.019716
R41578 DVDD.n12613 DVDD.n12460 0.019716
R41579 DVDD.n12613 DVDD.n12416 0.019716
R41580 DVDD.n12618 DVDD.n12459 0.019716
R41581 DVDD.n12618 DVDD.n12415 0.019716
R41582 DVDD.n12622 DVDD.n12458 0.019716
R41583 DVDD.n12622 DVDD.n12414 0.019716
R41584 DVDD.n12627 DVDD.n12457 0.019716
R41585 DVDD.n12627 DVDD.n12413 0.019716
R41586 DVDD.n12631 DVDD.n12456 0.019716
R41587 DVDD.n12631 DVDD.n12412 0.019716
R41588 DVDD.n12636 DVDD.n12455 0.019716
R41589 DVDD.n12636 DVDD.n12411 0.019716
R41590 DVDD.n12640 DVDD.n12454 0.019716
R41591 DVDD.n12640 DVDD.n12410 0.019716
R41592 DVDD.n12645 DVDD.n12453 0.019716
R41593 DVDD.n12645 DVDD.n12409 0.019716
R41594 DVDD.n12649 DVDD.n12452 0.019716
R41595 DVDD.n12649 DVDD.n12408 0.019716
R41596 DVDD.n12654 DVDD.n12451 0.019716
R41597 DVDD.n12654 DVDD.n12407 0.019716
R41598 DVDD.n12658 DVDD.n12450 0.019716
R41599 DVDD.n12658 DVDD.n12406 0.019716
R41600 DVDD.n12663 DVDD.n12449 0.019716
R41601 DVDD.n12663 DVDD.n12405 0.019716
R41602 DVDD.n12667 DVDD.n12448 0.019716
R41603 DVDD.n12667 DVDD.n12404 0.019716
R41604 DVDD.n12672 DVDD.n12447 0.019716
R41605 DVDD.n12672 DVDD.n12403 0.019716
R41606 DVDD.n12676 DVDD.n12446 0.019716
R41607 DVDD.n12676 DVDD.n12402 0.019716
R41608 DVDD.n12681 DVDD.n12445 0.019716
R41609 DVDD.n12681 DVDD.n12401 0.019716
R41610 DVDD.n12685 DVDD.n12444 0.019716
R41611 DVDD.n12685 DVDD.n12400 0.019716
R41612 DVDD.n12690 DVDD.n12443 0.019716
R41613 DVDD.n12690 DVDD.n12399 0.019716
R41614 DVDD.n12694 DVDD.n12442 0.019716
R41615 DVDD.n12694 DVDD.n12398 0.019716
R41616 DVDD.n12699 DVDD.n12441 0.019716
R41617 DVDD.n12699 DVDD.n12397 0.019716
R41618 DVDD.n12703 DVDD.n12440 0.019716
R41619 DVDD.n12703 DVDD.n12396 0.019716
R41620 DVDD.n12708 DVDD.n12439 0.019716
R41621 DVDD.n12708 DVDD.n12395 0.019716
R41622 DVDD.n12712 DVDD.n12438 0.019716
R41623 DVDD.n12712 DVDD.n12394 0.019716
R41624 DVDD.n12717 DVDD.n12437 0.019716
R41625 DVDD.n12717 DVDD.n12393 0.019716
R41626 DVDD.n12721 DVDD.n12436 0.019716
R41627 DVDD.n12721 DVDD.n12392 0.019716
R41628 DVDD.n13483 DVDD.n12391 0.019716
R41629 DVDD.n12374 DVDD.n12329 0.019716
R41630 DVDD.n12375 DVDD.n12328 0.019716
R41631 DVDD.n13503 DVDD.n12327 0.019716
R41632 DVDD.n13503 DVDD.n13502 0.019716
R41633 DVDD.n13505 DVDD.n12326 0.019716
R41634 DVDD.n13506 DVDD.n13505 0.019716
R41635 DVDD.n13515 DVDD.n12325 0.019716
R41636 DVDD.n13515 DVDD.n13514 0.019716
R41637 DVDD.n13517 DVDD.n12324 0.019716
R41638 DVDD.n13518 DVDD.n13517 0.019716
R41639 DVDD.n13527 DVDD.n12323 0.019716
R41640 DVDD.n13527 DVDD.n13526 0.019716
R41641 DVDD.n13529 DVDD.n12322 0.019716
R41642 DVDD.n13530 DVDD.n13529 0.019716
R41643 DVDD.n13539 DVDD.n12321 0.019716
R41644 DVDD.n13539 DVDD.n13538 0.019716
R41645 DVDD.n13541 DVDD.n12320 0.019716
R41646 DVDD.n13542 DVDD.n13541 0.019716
R41647 DVDD.n13551 DVDD.n12319 0.019716
R41648 DVDD.n13551 DVDD.n13550 0.019716
R41649 DVDD.n13553 DVDD.n12318 0.019716
R41650 DVDD.n13554 DVDD.n13553 0.019716
R41651 DVDD.n13563 DVDD.n12317 0.019716
R41652 DVDD.n13563 DVDD.n13562 0.019716
R41653 DVDD.n13565 DVDD.n12316 0.019716
R41654 DVDD.n13566 DVDD.n13565 0.019716
R41655 DVDD.n13575 DVDD.n12315 0.019716
R41656 DVDD.n13575 DVDD.n13574 0.019716
R41657 DVDD.n13577 DVDD.n12314 0.019716
R41658 DVDD.n13578 DVDD.n13577 0.019716
R41659 DVDD.n13587 DVDD.n12313 0.019716
R41660 DVDD.n13587 DVDD.n13586 0.019716
R41661 DVDD.n13589 DVDD.n12312 0.019716
R41662 DVDD.n13590 DVDD.n13589 0.019716
R41663 DVDD.n13599 DVDD.n12311 0.019716
R41664 DVDD.n13599 DVDD.n13598 0.019716
R41665 DVDD.n13601 DVDD.n12310 0.019716
R41666 DVDD.n13602 DVDD.n13601 0.019716
R41667 DVDD.n13611 DVDD.n12309 0.019716
R41668 DVDD.n13611 DVDD.n13610 0.019716
R41669 DVDD.n13613 DVDD.n12308 0.019716
R41670 DVDD.n13614 DVDD.n13613 0.019716
R41671 DVDD.n13623 DVDD.n12307 0.019716
R41672 DVDD.n13623 DVDD.n13622 0.019716
R41673 DVDD.n13625 DVDD.n12306 0.019716
R41674 DVDD.n13626 DVDD.n13625 0.019716
R41675 DVDD.n13635 DVDD.n12305 0.019716
R41676 DVDD.n13635 DVDD.n13634 0.019716
R41677 DVDD.n13637 DVDD.n12304 0.019716
R41678 DVDD.n13638 DVDD.n13637 0.019716
R41679 DVDD.n13647 DVDD.n12303 0.019716
R41680 DVDD.n13647 DVDD.n13646 0.019716
R41681 DVDD.n13649 DVDD.n12302 0.019716
R41682 DVDD.n13650 DVDD.n13649 0.019716
R41683 DVDD.n13659 DVDD.n12301 0.019716
R41684 DVDD.n13659 DVDD.n13658 0.019716
R41685 DVDD.n13661 DVDD.n12300 0.019716
R41686 DVDD.n13662 DVDD.n13661 0.019716
R41687 DVDD.n13671 DVDD.n12299 0.019716
R41688 DVDD.n13671 DVDD.n13670 0.019716
R41689 DVDD.n13673 DVDD.n12298 0.019716
R41690 DVDD.n13674 DVDD.n13673 0.019716
R41691 DVDD.n13683 DVDD.n12297 0.019716
R41692 DVDD.n13683 DVDD.n13682 0.019716
R41693 DVDD.n13685 DVDD.n12296 0.019716
R41694 DVDD.n13686 DVDD.n13685 0.019716
R41695 DVDD.n13695 DVDD.n12295 0.019716
R41696 DVDD.n13695 DVDD.n13694 0.019716
R41697 DVDD.n13697 DVDD.n12294 0.019716
R41698 DVDD.n13698 DVDD.n13697 0.019716
R41699 DVDD.n13707 DVDD.n12293 0.019716
R41700 DVDD.n13707 DVDD.n13706 0.019716
R41701 DVDD.n13709 DVDD.n12292 0.019716
R41702 DVDD.n13710 DVDD.n13709 0.019716
R41703 DVDD.n13719 DVDD.n12291 0.019716
R41704 DVDD.n13719 DVDD.n13718 0.019716
R41705 DVDD.n13721 DVDD.n12290 0.019716
R41706 DVDD.n13722 DVDD.n13721 0.019716
R41707 DVDD.n13731 DVDD.n12289 0.019716
R41708 DVDD.n13731 DVDD.n13730 0.019716
R41709 DVDD.n13733 DVDD.n12288 0.019716
R41710 DVDD.n13734 DVDD.n13733 0.019716
R41711 DVDD.n13743 DVDD.n13742 0.019716
R41712 DVDD.n12029 DVDD.n12028 0.019716
R41713 DVDD.n12031 DVDD.n12030 0.019716
R41714 DVDD.n12032 DVDD.n12023 0.019716
R41715 DVDD.n12033 DVDD.n12032 0.019716
R41716 DVDD.n12043 DVDD.n12042 0.019716
R41717 DVDD.n12042 DVDD.n12041 0.019716
R41718 DVDD.n12044 DVDD.n12019 0.019716
R41719 DVDD.n12045 DVDD.n12044 0.019716
R41720 DVDD.n12055 DVDD.n12054 0.019716
R41721 DVDD.n12054 DVDD.n12053 0.019716
R41722 DVDD.n12056 DVDD.n12015 0.019716
R41723 DVDD.n12057 DVDD.n12056 0.019716
R41724 DVDD.n12067 DVDD.n12066 0.019716
R41725 DVDD.n12066 DVDD.n12065 0.019716
R41726 DVDD.n12068 DVDD.n12011 0.019716
R41727 DVDD.n12069 DVDD.n12068 0.019716
R41728 DVDD.n12079 DVDD.n12078 0.019716
R41729 DVDD.n12078 DVDD.n12077 0.019716
R41730 DVDD.n12080 DVDD.n12007 0.019716
R41731 DVDD.n12081 DVDD.n12080 0.019716
R41732 DVDD.n12091 DVDD.n12090 0.019716
R41733 DVDD.n12090 DVDD.n12089 0.019716
R41734 DVDD.n12092 DVDD.n12003 0.019716
R41735 DVDD.n12093 DVDD.n12092 0.019716
R41736 DVDD.n12103 DVDD.n12102 0.019716
R41737 DVDD.n12102 DVDD.n12101 0.019716
R41738 DVDD.n12104 DVDD.n11999 0.019716
R41739 DVDD.n12105 DVDD.n12104 0.019716
R41740 DVDD.n12115 DVDD.n12114 0.019716
R41741 DVDD.n12114 DVDD.n12113 0.019716
R41742 DVDD.n12116 DVDD.n11995 0.019716
R41743 DVDD.n12117 DVDD.n12116 0.019716
R41744 DVDD.n12127 DVDD.n12126 0.019716
R41745 DVDD.n12126 DVDD.n12125 0.019716
R41746 DVDD.n12128 DVDD.n11991 0.019716
R41747 DVDD.n12129 DVDD.n12128 0.019716
R41748 DVDD.n12139 DVDD.n12138 0.019716
R41749 DVDD.n12138 DVDD.n12137 0.019716
R41750 DVDD.n12140 DVDD.n11987 0.019716
R41751 DVDD.n12141 DVDD.n12140 0.019716
R41752 DVDD.n12151 DVDD.n12150 0.019716
R41753 DVDD.n12150 DVDD.n12149 0.019716
R41754 DVDD.n12152 DVDD.n11983 0.019716
R41755 DVDD.n12153 DVDD.n12152 0.019716
R41756 DVDD.n12163 DVDD.n12162 0.019716
R41757 DVDD.n12162 DVDD.n12161 0.019716
R41758 DVDD.n12164 DVDD.n11979 0.019716
R41759 DVDD.n12165 DVDD.n12164 0.019716
R41760 DVDD.n12175 DVDD.n12174 0.019716
R41761 DVDD.n12174 DVDD.n12173 0.019716
R41762 DVDD.n12176 DVDD.n11975 0.019716
R41763 DVDD.n12177 DVDD.n12176 0.019716
R41764 DVDD.n12187 DVDD.n12186 0.019716
R41765 DVDD.n12186 DVDD.n12185 0.019716
R41766 DVDD.n12188 DVDD.n11971 0.019716
R41767 DVDD.n12189 DVDD.n12188 0.019716
R41768 DVDD.n12199 DVDD.n12198 0.019716
R41769 DVDD.n12198 DVDD.n12197 0.019716
R41770 DVDD.n12200 DVDD.n11967 0.019716
R41771 DVDD.n12201 DVDD.n12200 0.019716
R41772 DVDD.n12211 DVDD.n12210 0.019716
R41773 DVDD.n12210 DVDD.n12209 0.019716
R41774 DVDD.n12212 DVDD.n11963 0.019716
R41775 DVDD.n12213 DVDD.n12212 0.019716
R41776 DVDD.n12223 DVDD.n12222 0.019716
R41777 DVDD.n12222 DVDD.n12221 0.019716
R41778 DVDD.n12224 DVDD.n11959 0.019716
R41779 DVDD.n12225 DVDD.n12224 0.019716
R41780 DVDD.n12235 DVDD.n12234 0.019716
R41781 DVDD.n12234 DVDD.n12233 0.019716
R41782 DVDD.n12236 DVDD.n11955 0.019716
R41783 DVDD.n12237 DVDD.n12236 0.019716
R41784 DVDD.n12247 DVDD.n12246 0.019716
R41785 DVDD.n12246 DVDD.n12245 0.019716
R41786 DVDD.n12248 DVDD.n11951 0.019716
R41787 DVDD.n12249 DVDD.n12248 0.019716
R41788 DVDD.n12259 DVDD.n12258 0.019716
R41789 DVDD.n12258 DVDD.n12257 0.019716
R41790 DVDD.n12260 DVDD.n11947 0.019716
R41791 DVDD.n12261 DVDD.n12260 0.019716
R41792 DVDD.n12272 DVDD.n12271 0.019716
R41793 DVDD.n12271 DVDD.n12270 0.019716
R41794 DVDD.n12275 DVDD.n12274 0.019716
R41795 DVDD.n11675 DVDD.n11630 0.019716
R41796 DVDD.n11676 DVDD.n11629 0.019716
R41797 DVDD.n11683 DVDD.n11628 0.019716
R41798 DVDD.n11683 DVDD.n11682 0.019716
R41799 DVDD.n11685 DVDD.n11627 0.019716
R41800 DVDD.n11686 DVDD.n11685 0.019716
R41801 DVDD.n11695 DVDD.n11626 0.019716
R41802 DVDD.n11695 DVDD.n11694 0.019716
R41803 DVDD.n11697 DVDD.n11625 0.019716
R41804 DVDD.n11698 DVDD.n11697 0.019716
R41805 DVDD.n11707 DVDD.n11624 0.019716
R41806 DVDD.n11707 DVDD.n11706 0.019716
R41807 DVDD.n11709 DVDD.n11623 0.019716
R41808 DVDD.n11710 DVDD.n11709 0.019716
R41809 DVDD.n11719 DVDD.n11622 0.019716
R41810 DVDD.n11719 DVDD.n11718 0.019716
R41811 DVDD.n11721 DVDD.n11621 0.019716
R41812 DVDD.n11722 DVDD.n11721 0.019716
R41813 DVDD.n11731 DVDD.n11620 0.019716
R41814 DVDD.n11731 DVDD.n11730 0.019716
R41815 DVDD.n11733 DVDD.n11619 0.019716
R41816 DVDD.n11734 DVDD.n11733 0.019716
R41817 DVDD.n11743 DVDD.n11618 0.019716
R41818 DVDD.n11743 DVDD.n11742 0.019716
R41819 DVDD.n11745 DVDD.n11617 0.019716
R41820 DVDD.n11746 DVDD.n11745 0.019716
R41821 DVDD.n11755 DVDD.n11616 0.019716
R41822 DVDD.n11755 DVDD.n11754 0.019716
R41823 DVDD.n11757 DVDD.n11615 0.019716
R41824 DVDD.n11758 DVDD.n11757 0.019716
R41825 DVDD.n11767 DVDD.n11614 0.019716
R41826 DVDD.n11767 DVDD.n11766 0.019716
R41827 DVDD.n11769 DVDD.n11613 0.019716
R41828 DVDD.n11770 DVDD.n11769 0.019716
R41829 DVDD.n11779 DVDD.n11612 0.019716
R41830 DVDD.n11779 DVDD.n11778 0.019716
R41831 DVDD.n11781 DVDD.n11611 0.019716
R41832 DVDD.n11782 DVDD.n11781 0.019716
R41833 DVDD.n11791 DVDD.n11610 0.019716
R41834 DVDD.n11791 DVDD.n11790 0.019716
R41835 DVDD.n11793 DVDD.n11609 0.019716
R41836 DVDD.n11794 DVDD.n11793 0.019716
R41837 DVDD.n11803 DVDD.n11608 0.019716
R41838 DVDD.n11803 DVDD.n11802 0.019716
R41839 DVDD.n11805 DVDD.n11607 0.019716
R41840 DVDD.n11806 DVDD.n11805 0.019716
R41841 DVDD.n11815 DVDD.n11606 0.019716
R41842 DVDD.n11815 DVDD.n11814 0.019716
R41843 DVDD.n11817 DVDD.n11605 0.019716
R41844 DVDD.n11818 DVDD.n11817 0.019716
R41845 DVDD.n11827 DVDD.n11604 0.019716
R41846 DVDD.n11827 DVDD.n11826 0.019716
R41847 DVDD.n11829 DVDD.n11603 0.019716
R41848 DVDD.n11830 DVDD.n11829 0.019716
R41849 DVDD.n11839 DVDD.n11602 0.019716
R41850 DVDD.n11839 DVDD.n11838 0.019716
R41851 DVDD.n11841 DVDD.n11601 0.019716
R41852 DVDD.n11842 DVDD.n11841 0.019716
R41853 DVDD.n11851 DVDD.n11600 0.019716
R41854 DVDD.n11851 DVDD.n11850 0.019716
R41855 DVDD.n11853 DVDD.n11599 0.019716
R41856 DVDD.n11854 DVDD.n11853 0.019716
R41857 DVDD.n11863 DVDD.n11598 0.019716
R41858 DVDD.n11863 DVDD.n11862 0.019716
R41859 DVDD.n11865 DVDD.n11597 0.019716
R41860 DVDD.n11866 DVDD.n11865 0.019716
R41861 DVDD.n11875 DVDD.n11596 0.019716
R41862 DVDD.n11875 DVDD.n11874 0.019716
R41863 DVDD.n11877 DVDD.n11595 0.019716
R41864 DVDD.n11878 DVDD.n11877 0.019716
R41865 DVDD.n11887 DVDD.n11594 0.019716
R41866 DVDD.n11887 DVDD.n11886 0.019716
R41867 DVDD.n11889 DVDD.n11593 0.019716
R41868 DVDD.n11890 DVDD.n11889 0.019716
R41869 DVDD.n11899 DVDD.n11592 0.019716
R41870 DVDD.n11899 DVDD.n11898 0.019716
R41871 DVDD.n11901 DVDD.n11591 0.019716
R41872 DVDD.n11902 DVDD.n11901 0.019716
R41873 DVDD.n11911 DVDD.n11590 0.019716
R41874 DVDD.n11911 DVDD.n11910 0.019716
R41875 DVDD.n11913 DVDD.n11589 0.019716
R41876 DVDD.n11914 DVDD.n11913 0.019716
R41877 DVDD.n13776 DVDD.n13775 0.019716
R41878 DVDD.n11321 DVDD.n11275 0.019716
R41879 DVDD.n11322 DVDD.n11274 0.019716
R41880 DVDD.n11329 DVDD.n11273 0.019716
R41881 DVDD.n11329 DVDD.n11328 0.019716
R41882 DVDD.n11331 DVDD.n11272 0.019716
R41883 DVDD.n11332 DVDD.n11331 0.019716
R41884 DVDD.n11341 DVDD.n11271 0.019716
R41885 DVDD.n11341 DVDD.n11340 0.019716
R41886 DVDD.n11343 DVDD.n11270 0.019716
R41887 DVDD.n11344 DVDD.n11343 0.019716
R41888 DVDD.n11353 DVDD.n11269 0.019716
R41889 DVDD.n11353 DVDD.n11352 0.019716
R41890 DVDD.n11355 DVDD.n11268 0.019716
R41891 DVDD.n11356 DVDD.n11355 0.019716
R41892 DVDD.n11365 DVDD.n11267 0.019716
R41893 DVDD.n11365 DVDD.n11364 0.019716
R41894 DVDD.n11367 DVDD.n11266 0.019716
R41895 DVDD.n11368 DVDD.n11367 0.019716
R41896 DVDD.n11377 DVDD.n11265 0.019716
R41897 DVDD.n11377 DVDD.n11376 0.019716
R41898 DVDD.n11379 DVDD.n11264 0.019716
R41899 DVDD.n11380 DVDD.n11379 0.019716
R41900 DVDD.n11389 DVDD.n11263 0.019716
R41901 DVDD.n11389 DVDD.n11388 0.019716
R41902 DVDD.n11391 DVDD.n11262 0.019716
R41903 DVDD.n11392 DVDD.n11391 0.019716
R41904 DVDD.n11401 DVDD.n11261 0.019716
R41905 DVDD.n11401 DVDD.n11400 0.019716
R41906 DVDD.n11403 DVDD.n11260 0.019716
R41907 DVDD.n11404 DVDD.n11403 0.019716
R41908 DVDD.n11413 DVDD.n11259 0.019716
R41909 DVDD.n11413 DVDD.n11412 0.019716
R41910 DVDD.n11415 DVDD.n11258 0.019716
R41911 DVDD.n11416 DVDD.n11415 0.019716
R41912 DVDD.n11425 DVDD.n11257 0.019716
R41913 DVDD.n11425 DVDD.n11424 0.019716
R41914 DVDD.n11427 DVDD.n11256 0.019716
R41915 DVDD.n11428 DVDD.n11427 0.019716
R41916 DVDD.n11437 DVDD.n11255 0.019716
R41917 DVDD.n11437 DVDD.n11436 0.019716
R41918 DVDD.n11439 DVDD.n11254 0.019716
R41919 DVDD.n11440 DVDD.n11439 0.019716
R41920 DVDD.n11449 DVDD.n11253 0.019716
R41921 DVDD.n11449 DVDD.n11448 0.019716
R41922 DVDD.n11451 DVDD.n11252 0.019716
R41923 DVDD.n11452 DVDD.n11451 0.019716
R41924 DVDD.n11461 DVDD.n11251 0.019716
R41925 DVDD.n11461 DVDD.n11460 0.019716
R41926 DVDD.n11463 DVDD.n11250 0.019716
R41927 DVDD.n11464 DVDD.n11463 0.019716
R41928 DVDD.n11473 DVDD.n11249 0.019716
R41929 DVDD.n11473 DVDD.n11472 0.019716
R41930 DVDD.n11475 DVDD.n11248 0.019716
R41931 DVDD.n11476 DVDD.n11475 0.019716
R41932 DVDD.n11485 DVDD.n11247 0.019716
R41933 DVDD.n11485 DVDD.n11484 0.019716
R41934 DVDD.n11487 DVDD.n11246 0.019716
R41935 DVDD.n11488 DVDD.n11487 0.019716
R41936 DVDD.n11497 DVDD.n11245 0.019716
R41937 DVDD.n11497 DVDD.n11496 0.019716
R41938 DVDD.n11499 DVDD.n11244 0.019716
R41939 DVDD.n11500 DVDD.n11499 0.019716
R41940 DVDD.n11509 DVDD.n11243 0.019716
R41941 DVDD.n11509 DVDD.n11508 0.019716
R41942 DVDD.n11511 DVDD.n11242 0.019716
R41943 DVDD.n11512 DVDD.n11511 0.019716
R41944 DVDD.n11521 DVDD.n11241 0.019716
R41945 DVDD.n11521 DVDD.n11520 0.019716
R41946 DVDD.n11523 DVDD.n11240 0.019716
R41947 DVDD.n11524 DVDD.n11523 0.019716
R41948 DVDD.n11533 DVDD.n11239 0.019716
R41949 DVDD.n11533 DVDD.n11532 0.019716
R41950 DVDD.n11535 DVDD.n11238 0.019716
R41951 DVDD.n11536 DVDD.n11535 0.019716
R41952 DVDD.n11545 DVDD.n11237 0.019716
R41953 DVDD.n11545 DVDD.n11544 0.019716
R41954 DVDD.n11547 DVDD.n11236 0.019716
R41955 DVDD.n11548 DVDD.n11547 0.019716
R41956 DVDD.n11557 DVDD.n11235 0.019716
R41957 DVDD.n11557 DVDD.n11556 0.019716
R41958 DVDD.n11559 DVDD.n11234 0.019716
R41959 DVDD.n11560 DVDD.n11559 0.019716
R41960 DVDD.n13798 DVDD.n13797 0.019716
R41961 DVDD.n14002 DVDD.n14001 0.019716
R41962 DVDD.n11148 DVDD.n11104 0.019716
R41963 DVDD.n13818 DVDD.n11147 0.019716
R41964 DVDD.n13818 DVDD.n11102 0.019716
R41965 DVDD.n13822 DVDD.n11146 0.019716
R41966 DVDD.n13822 DVDD.n11101 0.019716
R41967 DVDD.n13827 DVDD.n11145 0.019716
R41968 DVDD.n13827 DVDD.n11100 0.019716
R41969 DVDD.n13831 DVDD.n11144 0.019716
R41970 DVDD.n13831 DVDD.n11099 0.019716
R41971 DVDD.n13836 DVDD.n11143 0.019716
R41972 DVDD.n13836 DVDD.n11098 0.019716
R41973 DVDD.n13840 DVDD.n11142 0.019716
R41974 DVDD.n13840 DVDD.n11097 0.019716
R41975 DVDD.n13845 DVDD.n11141 0.019716
R41976 DVDD.n13845 DVDD.n11096 0.019716
R41977 DVDD.n13849 DVDD.n11140 0.019716
R41978 DVDD.n13849 DVDD.n11095 0.019716
R41979 DVDD.n13854 DVDD.n11139 0.019716
R41980 DVDD.n13854 DVDD.n11094 0.019716
R41981 DVDD.n13858 DVDD.n11138 0.019716
R41982 DVDD.n13858 DVDD.n11093 0.019716
R41983 DVDD.n13863 DVDD.n11137 0.019716
R41984 DVDD.n13863 DVDD.n11092 0.019716
R41985 DVDD.n13867 DVDD.n11136 0.019716
R41986 DVDD.n13867 DVDD.n11091 0.019716
R41987 DVDD.n13872 DVDD.n11135 0.019716
R41988 DVDD.n13872 DVDD.n11090 0.019716
R41989 DVDD.n13876 DVDD.n11134 0.019716
R41990 DVDD.n13876 DVDD.n11089 0.019716
R41991 DVDD.n13881 DVDD.n11133 0.019716
R41992 DVDD.n13881 DVDD.n11088 0.019716
R41993 DVDD.n13885 DVDD.n11132 0.019716
R41994 DVDD.n13885 DVDD.n11087 0.019716
R41995 DVDD.n13890 DVDD.n11131 0.019716
R41996 DVDD.n13890 DVDD.n11086 0.019716
R41997 DVDD.n13894 DVDD.n11130 0.019716
R41998 DVDD.n13894 DVDD.n11085 0.019716
R41999 DVDD.n13899 DVDD.n11129 0.019716
R42000 DVDD.n13899 DVDD.n11084 0.019716
R42001 DVDD.n13903 DVDD.n11128 0.019716
R42002 DVDD.n13903 DVDD.n11083 0.019716
R42003 DVDD.n13908 DVDD.n11127 0.019716
R42004 DVDD.n13908 DVDD.n11082 0.019716
R42005 DVDD.n13912 DVDD.n11126 0.019716
R42006 DVDD.n13912 DVDD.n11081 0.019716
R42007 DVDD.n13917 DVDD.n11125 0.019716
R42008 DVDD.n13917 DVDD.n11080 0.019716
R42009 DVDD.n13921 DVDD.n11124 0.019716
R42010 DVDD.n13921 DVDD.n11079 0.019716
R42011 DVDD.n13926 DVDD.n11123 0.019716
R42012 DVDD.n13926 DVDD.n11078 0.019716
R42013 DVDD.n13930 DVDD.n11122 0.019716
R42014 DVDD.n13930 DVDD.n11077 0.019716
R42015 DVDD.n13935 DVDD.n11121 0.019716
R42016 DVDD.n13935 DVDD.n11076 0.019716
R42017 DVDD.n13939 DVDD.n11120 0.019716
R42018 DVDD.n13939 DVDD.n11075 0.019716
R42019 DVDD.n13944 DVDD.n11119 0.019716
R42020 DVDD.n13944 DVDD.n11074 0.019716
R42021 DVDD.n13948 DVDD.n11118 0.019716
R42022 DVDD.n13948 DVDD.n11073 0.019716
R42023 DVDD.n13953 DVDD.n11117 0.019716
R42024 DVDD.n13953 DVDD.n11072 0.019716
R42025 DVDD.n13957 DVDD.n11116 0.019716
R42026 DVDD.n13957 DVDD.n11071 0.019716
R42027 DVDD.n13962 DVDD.n11115 0.019716
R42028 DVDD.n13962 DVDD.n11070 0.019716
R42029 DVDD.n13966 DVDD.n11114 0.019716
R42030 DVDD.n13966 DVDD.n11069 0.019716
R42031 DVDD.n13971 DVDD.n11113 0.019716
R42032 DVDD.n13971 DVDD.n11068 0.019716
R42033 DVDD.n13975 DVDD.n11112 0.019716
R42034 DVDD.n13975 DVDD.n11067 0.019716
R42035 DVDD.n13980 DVDD.n11111 0.019716
R42036 DVDD.n13980 DVDD.n11066 0.019716
R42037 DVDD.n13984 DVDD.n11110 0.019716
R42038 DVDD.n13984 DVDD.n11065 0.019716
R42039 DVDD.n13989 DVDD.n11109 0.019716
R42040 DVDD.n13989 DVDD.n11064 0.019716
R42041 DVDD.n13993 DVDD.n11108 0.019716
R42042 DVDD.n13993 DVDD.n11063 0.019716
R42043 DVDD.n13999 DVDD.n11062 0.019716
R42044 DVDD.n10802 DVDD.n10801 0.019716
R42045 DVDD.n10804 DVDD.n10803 0.019716
R42046 DVDD.n10805 DVDD.n10795 0.019716
R42047 DVDD.n10806 DVDD.n10805 0.019716
R42048 DVDD.n10816 DVDD.n10815 0.019716
R42049 DVDD.n10815 DVDD.n10814 0.019716
R42050 DVDD.n10817 DVDD.n10791 0.019716
R42051 DVDD.n10818 DVDD.n10817 0.019716
R42052 DVDD.n10828 DVDD.n10827 0.019716
R42053 DVDD.n10827 DVDD.n10826 0.019716
R42054 DVDD.n10829 DVDD.n10787 0.019716
R42055 DVDD.n10830 DVDD.n10829 0.019716
R42056 DVDD.n10840 DVDD.n10839 0.019716
R42057 DVDD.n10839 DVDD.n10838 0.019716
R42058 DVDD.n10841 DVDD.n10783 0.019716
R42059 DVDD.n10842 DVDD.n10841 0.019716
R42060 DVDD.n10852 DVDD.n10851 0.019716
R42061 DVDD.n10851 DVDD.n10850 0.019716
R42062 DVDD.n10853 DVDD.n10779 0.019716
R42063 DVDD.n10854 DVDD.n10853 0.019716
R42064 DVDD.n10864 DVDD.n10863 0.019716
R42065 DVDD.n10863 DVDD.n10862 0.019716
R42066 DVDD.n10865 DVDD.n10775 0.019716
R42067 DVDD.n10866 DVDD.n10865 0.019716
R42068 DVDD.n10876 DVDD.n10875 0.019716
R42069 DVDD.n10875 DVDD.n10874 0.019716
R42070 DVDD.n10877 DVDD.n10771 0.019716
R42071 DVDD.n10878 DVDD.n10877 0.019716
R42072 DVDD.n10888 DVDD.n10887 0.019716
R42073 DVDD.n10887 DVDD.n10886 0.019716
R42074 DVDD.n10889 DVDD.n10767 0.019716
R42075 DVDD.n10890 DVDD.n10889 0.019716
R42076 DVDD.n10900 DVDD.n10899 0.019716
R42077 DVDD.n10899 DVDD.n10898 0.019716
R42078 DVDD.n10901 DVDD.n10763 0.019716
R42079 DVDD.n10902 DVDD.n10901 0.019716
R42080 DVDD.n10912 DVDD.n10911 0.019716
R42081 DVDD.n10911 DVDD.n10910 0.019716
R42082 DVDD.n10913 DVDD.n10759 0.019716
R42083 DVDD.n10914 DVDD.n10913 0.019716
R42084 DVDD.n10924 DVDD.n10923 0.019716
R42085 DVDD.n10923 DVDD.n10922 0.019716
R42086 DVDD.n10925 DVDD.n10755 0.019716
R42087 DVDD.n10926 DVDD.n10925 0.019716
R42088 DVDD.n10936 DVDD.n10935 0.019716
R42089 DVDD.n10935 DVDD.n10934 0.019716
R42090 DVDD.n10937 DVDD.n10751 0.019716
R42091 DVDD.n10938 DVDD.n10937 0.019716
R42092 DVDD.n10948 DVDD.n10947 0.019716
R42093 DVDD.n10947 DVDD.n10946 0.019716
R42094 DVDD.n10949 DVDD.n10747 0.019716
R42095 DVDD.n10950 DVDD.n10949 0.019716
R42096 DVDD.n10960 DVDD.n10959 0.019716
R42097 DVDD.n10959 DVDD.n10958 0.019716
R42098 DVDD.n10961 DVDD.n10743 0.019716
R42099 DVDD.n10962 DVDD.n10961 0.019716
R42100 DVDD.n10972 DVDD.n10971 0.019716
R42101 DVDD.n10971 DVDD.n10970 0.019716
R42102 DVDD.n10973 DVDD.n10739 0.019716
R42103 DVDD.n10974 DVDD.n10973 0.019716
R42104 DVDD.n10984 DVDD.n10983 0.019716
R42105 DVDD.n10983 DVDD.n10982 0.019716
R42106 DVDD.n10985 DVDD.n10735 0.019716
R42107 DVDD.n10986 DVDD.n10985 0.019716
R42108 DVDD.n10996 DVDD.n10995 0.019716
R42109 DVDD.n10995 DVDD.n10994 0.019716
R42110 DVDD.n10997 DVDD.n10731 0.019716
R42111 DVDD.n10998 DVDD.n10997 0.019716
R42112 DVDD.n11008 DVDD.n11007 0.019716
R42113 DVDD.n11007 DVDD.n11006 0.019716
R42114 DVDD.n11009 DVDD.n10727 0.019716
R42115 DVDD.n11010 DVDD.n11009 0.019716
R42116 DVDD.n11020 DVDD.n11019 0.019716
R42117 DVDD.n11019 DVDD.n11018 0.019716
R42118 DVDD.n11021 DVDD.n10723 0.019716
R42119 DVDD.n11022 DVDD.n11021 0.019716
R42120 DVDD.n11032 DVDD.n11031 0.019716
R42121 DVDD.n11031 DVDD.n11030 0.019716
R42122 DVDD.n11033 DVDD.n10719 0.019716
R42123 DVDD.n11034 DVDD.n11033 0.019716
R42124 DVDD.n11045 DVDD.n11044 0.019716
R42125 DVDD.n11044 DVDD.n11043 0.019716
R42126 DVDD.n11048 DVDD.n11047 0.019716
R42127 DVDD.n10683 DVDD.n10639 0.019716
R42128 DVDD.n10684 DVDD.n10638 0.019716
R42129 DVDD.n14028 DVDD.n10637 0.019716
R42130 DVDD.n14028 DVDD.n14027 0.019716
R42131 DVDD.n14030 DVDD.n10636 0.019716
R42132 DVDD.n14031 DVDD.n14030 0.019716
R42133 DVDD.n14040 DVDD.n10635 0.019716
R42134 DVDD.n14040 DVDD.n14039 0.019716
R42135 DVDD.n14042 DVDD.n10634 0.019716
R42136 DVDD.n14043 DVDD.n14042 0.019716
R42137 DVDD.n14052 DVDD.n10633 0.019716
R42138 DVDD.n14052 DVDD.n14051 0.019716
R42139 DVDD.n14054 DVDD.n10632 0.019716
R42140 DVDD.n14055 DVDD.n14054 0.019716
R42141 DVDD.n14064 DVDD.n10631 0.019716
R42142 DVDD.n14064 DVDD.n14063 0.019716
R42143 DVDD.n14066 DVDD.n10630 0.019716
R42144 DVDD.n14067 DVDD.n14066 0.019716
R42145 DVDD.n14076 DVDD.n10629 0.019716
R42146 DVDD.n14076 DVDD.n14075 0.019716
R42147 DVDD.n14078 DVDD.n10628 0.019716
R42148 DVDD.n14079 DVDD.n14078 0.019716
R42149 DVDD.n14088 DVDD.n10627 0.019716
R42150 DVDD.n14088 DVDD.n14087 0.019716
R42151 DVDD.n14090 DVDD.n10626 0.019716
R42152 DVDD.n14091 DVDD.n14090 0.019716
R42153 DVDD.n14100 DVDD.n10625 0.019716
R42154 DVDD.n14100 DVDD.n14099 0.019716
R42155 DVDD.n14102 DVDD.n10624 0.019716
R42156 DVDD.n14103 DVDD.n14102 0.019716
R42157 DVDD.n14112 DVDD.n10623 0.019716
R42158 DVDD.n14112 DVDD.n14111 0.019716
R42159 DVDD.n14114 DVDD.n10622 0.019716
R42160 DVDD.n14115 DVDD.n14114 0.019716
R42161 DVDD.n14124 DVDD.n10621 0.019716
R42162 DVDD.n14124 DVDD.n14123 0.019716
R42163 DVDD.n14126 DVDD.n10620 0.019716
R42164 DVDD.n14127 DVDD.n14126 0.019716
R42165 DVDD.n14136 DVDD.n10619 0.019716
R42166 DVDD.n14136 DVDD.n14135 0.019716
R42167 DVDD.n14138 DVDD.n10618 0.019716
R42168 DVDD.n14139 DVDD.n14138 0.019716
R42169 DVDD.n14148 DVDD.n10617 0.019716
R42170 DVDD.n14148 DVDD.n14147 0.019716
R42171 DVDD.n14150 DVDD.n10616 0.019716
R42172 DVDD.n14151 DVDD.n14150 0.019716
R42173 DVDD.n14160 DVDD.n10615 0.019716
R42174 DVDD.n14160 DVDD.n14159 0.019716
R42175 DVDD.n14162 DVDD.n10614 0.019716
R42176 DVDD.n14163 DVDD.n14162 0.019716
R42177 DVDD.n14172 DVDD.n10613 0.019716
R42178 DVDD.n14172 DVDD.n14171 0.019716
R42179 DVDD.n14174 DVDD.n10612 0.019716
R42180 DVDD.n14175 DVDD.n14174 0.019716
R42181 DVDD.n14184 DVDD.n10611 0.019716
R42182 DVDD.n14184 DVDD.n14183 0.019716
R42183 DVDD.n14186 DVDD.n10610 0.019716
R42184 DVDD.n14187 DVDD.n14186 0.019716
R42185 DVDD.n14196 DVDD.n10609 0.019716
R42186 DVDD.n14196 DVDD.n14195 0.019716
R42187 DVDD.n14198 DVDD.n10608 0.019716
R42188 DVDD.n14199 DVDD.n14198 0.019716
R42189 DVDD.n14208 DVDD.n10607 0.019716
R42190 DVDD.n14208 DVDD.n14207 0.019716
R42191 DVDD.n14210 DVDD.n10606 0.019716
R42192 DVDD.n14211 DVDD.n14210 0.019716
R42193 DVDD.n14220 DVDD.n10605 0.019716
R42194 DVDD.n14220 DVDD.n14219 0.019716
R42195 DVDD.n14222 DVDD.n10604 0.019716
R42196 DVDD.n14223 DVDD.n14222 0.019716
R42197 DVDD.n14232 DVDD.n10603 0.019716
R42198 DVDD.n14232 DVDD.n14231 0.019716
R42199 DVDD.n14234 DVDD.n10602 0.019716
R42200 DVDD.n14235 DVDD.n14234 0.019716
R42201 DVDD.n14244 DVDD.n10601 0.019716
R42202 DVDD.n14244 DVDD.n14243 0.019716
R42203 DVDD.n14246 DVDD.n10600 0.019716
R42204 DVDD.n14247 DVDD.n14246 0.019716
R42205 DVDD.n14256 DVDD.n10599 0.019716
R42206 DVDD.n14256 DVDD.n14255 0.019716
R42207 DVDD.n14258 DVDD.n10598 0.019716
R42208 DVDD.n14259 DVDD.n14258 0.019716
R42209 DVDD.n14268 DVDD.n14267 0.019716
R42210 DVDD.n14283 DVDD.n14282 0.019716
R42211 DVDD.n10327 DVDD.n10284 0.019716
R42212 DVDD.n10397 DVDD.n10326 0.019716
R42213 DVDD.n10397 DVDD.n10282 0.019716
R42214 DVDD.n10401 DVDD.n10325 0.019716
R42215 DVDD.n10401 DVDD.n10281 0.019716
R42216 DVDD.n10406 DVDD.n10324 0.019716
R42217 DVDD.n10406 DVDD.n10280 0.019716
R42218 DVDD.n10410 DVDD.n10323 0.019716
R42219 DVDD.n10410 DVDD.n10279 0.019716
R42220 DVDD.n10415 DVDD.n10322 0.019716
R42221 DVDD.n10415 DVDD.n10278 0.019716
R42222 DVDD.n10419 DVDD.n10321 0.019716
R42223 DVDD.n10419 DVDD.n10277 0.019716
R42224 DVDD.n10424 DVDD.n10320 0.019716
R42225 DVDD.n10424 DVDD.n10276 0.019716
R42226 DVDD.n10428 DVDD.n10319 0.019716
R42227 DVDD.n10428 DVDD.n10275 0.019716
R42228 DVDD.n10433 DVDD.n10318 0.019716
R42229 DVDD.n10433 DVDD.n10274 0.019716
R42230 DVDD.n10437 DVDD.n10317 0.019716
R42231 DVDD.n10437 DVDD.n10273 0.019716
R42232 DVDD.n10442 DVDD.n10316 0.019716
R42233 DVDD.n10442 DVDD.n10272 0.019716
R42234 DVDD.n10446 DVDD.n10315 0.019716
R42235 DVDD.n10446 DVDD.n10271 0.019716
R42236 DVDD.n10451 DVDD.n10314 0.019716
R42237 DVDD.n10451 DVDD.n10270 0.019716
R42238 DVDD.n10455 DVDD.n10313 0.019716
R42239 DVDD.n10455 DVDD.n10269 0.019716
R42240 DVDD.n10460 DVDD.n10312 0.019716
R42241 DVDD.n10460 DVDD.n10268 0.019716
R42242 DVDD.n10464 DVDD.n10311 0.019716
R42243 DVDD.n10464 DVDD.n10267 0.019716
R42244 DVDD.n10469 DVDD.n10310 0.019716
R42245 DVDD.n10469 DVDD.n10266 0.019716
R42246 DVDD.n10473 DVDD.n10309 0.019716
R42247 DVDD.n10473 DVDD.n10265 0.019716
R42248 DVDD.n10478 DVDD.n10308 0.019716
R42249 DVDD.n10478 DVDD.n10264 0.019716
R42250 DVDD.n10482 DVDD.n10307 0.019716
R42251 DVDD.n10482 DVDD.n10263 0.019716
R42252 DVDD.n10487 DVDD.n10306 0.019716
R42253 DVDD.n10487 DVDD.n10262 0.019716
R42254 DVDD.n10491 DVDD.n10305 0.019716
R42255 DVDD.n10491 DVDD.n10261 0.019716
R42256 DVDD.n10496 DVDD.n10304 0.019716
R42257 DVDD.n10496 DVDD.n10260 0.019716
R42258 DVDD.n10500 DVDD.n10303 0.019716
R42259 DVDD.n10500 DVDD.n10259 0.019716
R42260 DVDD.n10505 DVDD.n10302 0.019716
R42261 DVDD.n10505 DVDD.n10258 0.019716
R42262 DVDD.n10509 DVDD.n10301 0.019716
R42263 DVDD.n10509 DVDD.n10257 0.019716
R42264 DVDD.n10514 DVDD.n10300 0.019716
R42265 DVDD.n10514 DVDD.n10256 0.019716
R42266 DVDD.n10518 DVDD.n10299 0.019716
R42267 DVDD.n10518 DVDD.n10255 0.019716
R42268 DVDD.n10523 DVDD.n10298 0.019716
R42269 DVDD.n10523 DVDD.n10254 0.019716
R42270 DVDD.n10527 DVDD.n10297 0.019716
R42271 DVDD.n10527 DVDD.n10253 0.019716
R42272 DVDD.n10532 DVDD.n10296 0.019716
R42273 DVDD.n10532 DVDD.n10252 0.019716
R42274 DVDD.n10536 DVDD.n10295 0.019716
R42275 DVDD.n10536 DVDD.n10251 0.019716
R42276 DVDD.n10541 DVDD.n10294 0.019716
R42277 DVDD.n10541 DVDD.n10250 0.019716
R42278 DVDD.n10545 DVDD.n10293 0.019716
R42279 DVDD.n10545 DVDD.n10249 0.019716
R42280 DVDD.n10550 DVDD.n10292 0.019716
R42281 DVDD.n10550 DVDD.n10248 0.019716
R42282 DVDD.n10554 DVDD.n10291 0.019716
R42283 DVDD.n10554 DVDD.n10247 0.019716
R42284 DVDD.n10559 DVDD.n10290 0.019716
R42285 DVDD.n10559 DVDD.n10246 0.019716
R42286 DVDD.n10563 DVDD.n10289 0.019716
R42287 DVDD.n10563 DVDD.n10245 0.019716
R42288 DVDD.n10568 DVDD.n10288 0.019716
R42289 DVDD.n10568 DVDD.n10244 0.019716
R42290 DVDD.n10572 DVDD.n10287 0.019716
R42291 DVDD.n10572 DVDD.n10243 0.019716
R42292 DVDD.n14280 DVDD.n10242 0.019716
R42293 DVDD.n8947 DVDD.n8946 0.019716
R42294 DVDD.n8945 DVDD.n8944 0.019716
R42295 DVDD.n8622 DVDD.n8621 0.019716
R42296 DVDD.n8621 DVDD.n8617 0.019716
R42297 DVDD.n8935 DVDD.n8934 0.019716
R42298 DVDD.n8936 DVDD.n8935 0.019716
R42299 DVDD.n8628 DVDD.n8627 0.019716
R42300 DVDD.n8627 DVDD.n8623 0.019716
R42301 DVDD.n8925 DVDD.n8924 0.019716
R42302 DVDD.n8926 DVDD.n8925 0.019716
R42303 DVDD.n8634 DVDD.n8633 0.019716
R42304 DVDD.n8633 DVDD.n8629 0.019716
R42305 DVDD.n8915 DVDD.n8914 0.019716
R42306 DVDD.n8916 DVDD.n8915 0.019716
R42307 DVDD.n8640 DVDD.n8639 0.019716
R42308 DVDD.n8639 DVDD.n8635 0.019716
R42309 DVDD.n8905 DVDD.n8904 0.019716
R42310 DVDD.n8906 DVDD.n8905 0.019716
R42311 DVDD.n8646 DVDD.n8645 0.019716
R42312 DVDD.n8645 DVDD.n8641 0.019716
R42313 DVDD.n8895 DVDD.n8894 0.019716
R42314 DVDD.n8896 DVDD.n8895 0.019716
R42315 DVDD.n8652 DVDD.n8651 0.019716
R42316 DVDD.n8651 DVDD.n8647 0.019716
R42317 DVDD.n8885 DVDD.n8884 0.019716
R42318 DVDD.n8886 DVDD.n8885 0.019716
R42319 DVDD.n8658 DVDD.n8657 0.019716
R42320 DVDD.n8657 DVDD.n8653 0.019716
R42321 DVDD.n8875 DVDD.n8874 0.019716
R42322 DVDD.n8876 DVDD.n8875 0.019716
R42323 DVDD.n8664 DVDD.n8663 0.019716
R42324 DVDD.n8663 DVDD.n8659 0.019716
R42325 DVDD.n8865 DVDD.n8864 0.019716
R42326 DVDD.n8866 DVDD.n8865 0.019716
R42327 DVDD.n8670 DVDD.n8669 0.019716
R42328 DVDD.n8669 DVDD.n8665 0.019716
R42329 DVDD.n8855 DVDD.n8854 0.019716
R42330 DVDD.n8856 DVDD.n8855 0.019716
R42331 DVDD.n8676 DVDD.n8675 0.019716
R42332 DVDD.n8675 DVDD.n8671 0.019716
R42333 DVDD.n8845 DVDD.n8844 0.019716
R42334 DVDD.n8846 DVDD.n8845 0.019716
R42335 DVDD.n8682 DVDD.n8681 0.019716
R42336 DVDD.n8681 DVDD.n8677 0.019716
R42337 DVDD.n8835 DVDD.n8834 0.019716
R42338 DVDD.n8836 DVDD.n8835 0.019716
R42339 DVDD.n8688 DVDD.n8687 0.019716
R42340 DVDD.n8687 DVDD.n8683 0.019716
R42341 DVDD.n8825 DVDD.n8824 0.019716
R42342 DVDD.n8826 DVDD.n8825 0.019716
R42343 DVDD.n8694 DVDD.n8693 0.019716
R42344 DVDD.n8693 DVDD.n8689 0.019716
R42345 DVDD.n8815 DVDD.n8814 0.019716
R42346 DVDD.n8816 DVDD.n8815 0.019716
R42347 DVDD.n8700 DVDD.n8699 0.019716
R42348 DVDD.n8699 DVDD.n8695 0.019716
R42349 DVDD.n8805 DVDD.n8804 0.019716
R42350 DVDD.n8806 DVDD.n8805 0.019716
R42351 DVDD.n8706 DVDD.n8705 0.019716
R42352 DVDD.n8705 DVDD.n8701 0.019716
R42353 DVDD.n8795 DVDD.n8794 0.019716
R42354 DVDD.n8796 DVDD.n8795 0.019716
R42355 DVDD.n8712 DVDD.n8711 0.019716
R42356 DVDD.n8711 DVDD.n8707 0.019716
R42357 DVDD.n8785 DVDD.n8784 0.019716
R42358 DVDD.n8786 DVDD.n8785 0.019716
R42359 DVDD.n8718 DVDD.n8717 0.019716
R42360 DVDD.n8717 DVDD.n8713 0.019716
R42361 DVDD.n8775 DVDD.n8774 0.019716
R42362 DVDD.n8776 DVDD.n8775 0.019716
R42363 DVDD.n8724 DVDD.n8723 0.019716
R42364 DVDD.n8723 DVDD.n8719 0.019716
R42365 DVDD.n8765 DVDD.n8764 0.019716
R42366 DVDD.n8766 DVDD.n8765 0.019716
R42367 DVDD.n8730 DVDD.n8729 0.019716
R42368 DVDD.n8729 DVDD.n8725 0.019716
R42369 DVDD.n8755 DVDD.n8754 0.019716
R42370 DVDD.n8756 DVDD.n8755 0.019716
R42371 DVDD.n8736 DVDD.n8735 0.019716
R42372 DVDD.n8735 DVDD.n8731 0.019716
R42373 DVDD.n8745 DVDD.n8744 0.019716
R42374 DVDD.n8746 DVDD.n8745 0.019716
R42375 DVDD.n8738 DVDD.n8737 0.019716
R42376 DVDD.n8350 DVDD.n8349 0.019716
R42377 DVDD.n8352 DVDD.n8351 0.019716
R42378 DVDD.n8353 DVDD.n8343 0.019716
R42379 DVDD.n8354 DVDD.n8353 0.019716
R42380 DVDD.n8364 DVDD.n8363 0.019716
R42381 DVDD.n8363 DVDD.n8362 0.019716
R42382 DVDD.n8365 DVDD.n8339 0.019716
R42383 DVDD.n8366 DVDD.n8365 0.019716
R42384 DVDD.n8376 DVDD.n8375 0.019716
R42385 DVDD.n8375 DVDD.n8374 0.019716
R42386 DVDD.n8377 DVDD.n8335 0.019716
R42387 DVDD.n8378 DVDD.n8377 0.019716
R42388 DVDD.n8388 DVDD.n8387 0.019716
R42389 DVDD.n8387 DVDD.n8386 0.019716
R42390 DVDD.n8389 DVDD.n8331 0.019716
R42391 DVDD.n8390 DVDD.n8389 0.019716
R42392 DVDD.n8400 DVDD.n8399 0.019716
R42393 DVDD.n8399 DVDD.n8398 0.019716
R42394 DVDD.n8401 DVDD.n8327 0.019716
R42395 DVDD.n8402 DVDD.n8401 0.019716
R42396 DVDD.n8412 DVDD.n8411 0.019716
R42397 DVDD.n8411 DVDD.n8410 0.019716
R42398 DVDD.n8413 DVDD.n8323 0.019716
R42399 DVDD.n8414 DVDD.n8413 0.019716
R42400 DVDD.n8424 DVDD.n8423 0.019716
R42401 DVDD.n8423 DVDD.n8422 0.019716
R42402 DVDD.n8425 DVDD.n8319 0.019716
R42403 DVDD.n8426 DVDD.n8425 0.019716
R42404 DVDD.n8436 DVDD.n8435 0.019716
R42405 DVDD.n8435 DVDD.n8434 0.019716
R42406 DVDD.n8437 DVDD.n8315 0.019716
R42407 DVDD.n8438 DVDD.n8437 0.019716
R42408 DVDD.n8448 DVDD.n8447 0.019716
R42409 DVDD.n8447 DVDD.n8446 0.019716
R42410 DVDD.n8449 DVDD.n8311 0.019716
R42411 DVDD.n8450 DVDD.n8449 0.019716
R42412 DVDD.n8460 DVDD.n8459 0.019716
R42413 DVDD.n8459 DVDD.n8458 0.019716
R42414 DVDD.n8461 DVDD.n8307 0.019716
R42415 DVDD.n8462 DVDD.n8461 0.019716
R42416 DVDD.n8472 DVDD.n8471 0.019716
R42417 DVDD.n8471 DVDD.n8470 0.019716
R42418 DVDD.n8473 DVDD.n8303 0.019716
R42419 DVDD.n8474 DVDD.n8473 0.019716
R42420 DVDD.n8484 DVDD.n8483 0.019716
R42421 DVDD.n8483 DVDD.n8482 0.019716
R42422 DVDD.n8485 DVDD.n8299 0.019716
R42423 DVDD.n8486 DVDD.n8485 0.019716
R42424 DVDD.n8496 DVDD.n8495 0.019716
R42425 DVDD.n8495 DVDD.n8494 0.019716
R42426 DVDD.n8497 DVDD.n8295 0.019716
R42427 DVDD.n8498 DVDD.n8497 0.019716
R42428 DVDD.n8508 DVDD.n8507 0.019716
R42429 DVDD.n8507 DVDD.n8506 0.019716
R42430 DVDD.n8509 DVDD.n8291 0.019716
R42431 DVDD.n8510 DVDD.n8509 0.019716
R42432 DVDD.n8520 DVDD.n8519 0.019716
R42433 DVDD.n8519 DVDD.n8518 0.019716
R42434 DVDD.n8521 DVDD.n8287 0.019716
R42435 DVDD.n8522 DVDD.n8521 0.019716
R42436 DVDD.n8532 DVDD.n8531 0.019716
R42437 DVDD.n8531 DVDD.n8530 0.019716
R42438 DVDD.n8533 DVDD.n8283 0.019716
R42439 DVDD.n8534 DVDD.n8533 0.019716
R42440 DVDD.n8544 DVDD.n8543 0.019716
R42441 DVDD.n8543 DVDD.n8542 0.019716
R42442 DVDD.n8545 DVDD.n8279 0.019716
R42443 DVDD.n8546 DVDD.n8545 0.019716
R42444 DVDD.n8556 DVDD.n8555 0.019716
R42445 DVDD.n8555 DVDD.n8554 0.019716
R42446 DVDD.n8557 DVDD.n8275 0.019716
R42447 DVDD.n8558 DVDD.n8557 0.019716
R42448 DVDD.n8568 DVDD.n8567 0.019716
R42449 DVDD.n8567 DVDD.n8566 0.019716
R42450 DVDD.n8569 DVDD.n8271 0.019716
R42451 DVDD.n8570 DVDD.n8569 0.019716
R42452 DVDD.n8580 DVDD.n8579 0.019716
R42453 DVDD.n8579 DVDD.n8578 0.019716
R42454 DVDD.n8581 DVDD.n8267 0.019716
R42455 DVDD.n8582 DVDD.n8581 0.019716
R42456 DVDD.n8593 DVDD.n8592 0.019716
R42457 DVDD.n8592 DVDD.n8591 0.019716
R42458 DVDD.n8596 DVDD.n8595 0.019716
R42459 DVDD.n8247 DVDD.n8204 0.019716
R42460 DVDD.n8248 DVDD.n8203 0.019716
R42461 DVDD.n14318 DVDD.n8202 0.019716
R42462 DVDD.n14318 DVDD.n14317 0.019716
R42463 DVDD.n14320 DVDD.n8201 0.019716
R42464 DVDD.n14321 DVDD.n14320 0.019716
R42465 DVDD.n14330 DVDD.n8200 0.019716
R42466 DVDD.n14330 DVDD.n14329 0.019716
R42467 DVDD.n14332 DVDD.n8199 0.019716
R42468 DVDD.n14333 DVDD.n14332 0.019716
R42469 DVDD.n14342 DVDD.n8198 0.019716
R42470 DVDD.n14342 DVDD.n14341 0.019716
R42471 DVDD.n14344 DVDD.n8197 0.019716
R42472 DVDD.n14345 DVDD.n14344 0.019716
R42473 DVDD.n14354 DVDD.n8196 0.019716
R42474 DVDD.n14354 DVDD.n14353 0.019716
R42475 DVDD.n14356 DVDD.n8195 0.019716
R42476 DVDD.n14357 DVDD.n14356 0.019716
R42477 DVDD.n14366 DVDD.n8194 0.019716
R42478 DVDD.n14366 DVDD.n14365 0.019716
R42479 DVDD.n14368 DVDD.n8193 0.019716
R42480 DVDD.n14369 DVDD.n14368 0.019716
R42481 DVDD.n14378 DVDD.n8192 0.019716
R42482 DVDD.n14378 DVDD.n14377 0.019716
R42483 DVDD.n14380 DVDD.n8191 0.019716
R42484 DVDD.n14381 DVDD.n14380 0.019716
R42485 DVDD.n14390 DVDD.n8190 0.019716
R42486 DVDD.n14390 DVDD.n14389 0.019716
R42487 DVDD.n14392 DVDD.n8189 0.019716
R42488 DVDD.n14393 DVDD.n14392 0.019716
R42489 DVDD.n14402 DVDD.n8188 0.019716
R42490 DVDD.n14402 DVDD.n14401 0.019716
R42491 DVDD.n14404 DVDD.n8187 0.019716
R42492 DVDD.n14405 DVDD.n14404 0.019716
R42493 DVDD.n14414 DVDD.n8186 0.019716
R42494 DVDD.n14414 DVDD.n14413 0.019716
R42495 DVDD.n14416 DVDD.n8185 0.019716
R42496 DVDD.n14417 DVDD.n14416 0.019716
R42497 DVDD.n14426 DVDD.n8184 0.019716
R42498 DVDD.n14426 DVDD.n14425 0.019716
R42499 DVDD.n14428 DVDD.n8183 0.019716
R42500 DVDD.n14429 DVDD.n14428 0.019716
R42501 DVDD.n14438 DVDD.n8182 0.019716
R42502 DVDD.n14438 DVDD.n14437 0.019716
R42503 DVDD.n14440 DVDD.n8181 0.019716
R42504 DVDD.n14441 DVDD.n14440 0.019716
R42505 DVDD.n14450 DVDD.n8180 0.019716
R42506 DVDD.n14450 DVDD.n14449 0.019716
R42507 DVDD.n14452 DVDD.n8179 0.019716
R42508 DVDD.n14453 DVDD.n14452 0.019716
R42509 DVDD.n14462 DVDD.n8178 0.019716
R42510 DVDD.n14462 DVDD.n14461 0.019716
R42511 DVDD.n14464 DVDD.n8177 0.019716
R42512 DVDD.n14465 DVDD.n14464 0.019716
R42513 DVDD.n14474 DVDD.n8176 0.019716
R42514 DVDD.n14474 DVDD.n14473 0.019716
R42515 DVDD.n14476 DVDD.n8175 0.019716
R42516 DVDD.n14477 DVDD.n14476 0.019716
R42517 DVDD.n14486 DVDD.n8174 0.019716
R42518 DVDD.n14486 DVDD.n14485 0.019716
R42519 DVDD.n14488 DVDD.n8173 0.019716
R42520 DVDD.n14489 DVDD.n14488 0.019716
R42521 DVDD.n14498 DVDD.n8172 0.019716
R42522 DVDD.n14498 DVDD.n14497 0.019716
R42523 DVDD.n14500 DVDD.n8171 0.019716
R42524 DVDD.n14501 DVDD.n14500 0.019716
R42525 DVDD.n14510 DVDD.n8170 0.019716
R42526 DVDD.n14510 DVDD.n14509 0.019716
R42527 DVDD.n14512 DVDD.n8169 0.019716
R42528 DVDD.n14513 DVDD.n14512 0.019716
R42529 DVDD.n14522 DVDD.n8168 0.019716
R42530 DVDD.n14522 DVDD.n14521 0.019716
R42531 DVDD.n14524 DVDD.n8167 0.019716
R42532 DVDD.n14525 DVDD.n14524 0.019716
R42533 DVDD.n14534 DVDD.n8166 0.019716
R42534 DVDD.n14534 DVDD.n14533 0.019716
R42535 DVDD.n14536 DVDD.n8165 0.019716
R42536 DVDD.n14537 DVDD.n14536 0.019716
R42537 DVDD.n14546 DVDD.n8164 0.019716
R42538 DVDD.n14546 DVDD.n14545 0.019716
R42539 DVDD.n14548 DVDD.n8163 0.019716
R42540 DVDD.n14549 DVDD.n14548 0.019716
R42541 DVDD.n14558 DVDD.n14557 0.019716
R42542 DVDD.n8130 DVDD.n8086 0.019716
R42543 DVDD.n8131 DVDD.n8085 0.019716
R42544 DVDD.n14584 DVDD.n8084 0.019716
R42545 DVDD.n14584 DVDD.n14583 0.019716
R42546 DVDD.n14586 DVDD.n8083 0.019716
R42547 DVDD.n14587 DVDD.n14586 0.019716
R42548 DVDD.n14596 DVDD.n8082 0.019716
R42549 DVDD.n14596 DVDD.n14595 0.019716
R42550 DVDD.n14598 DVDD.n8081 0.019716
R42551 DVDD.n14599 DVDD.n14598 0.019716
R42552 DVDD.n14608 DVDD.n8080 0.019716
R42553 DVDD.n14608 DVDD.n14607 0.019716
R42554 DVDD.n14610 DVDD.n8079 0.019716
R42555 DVDD.n14611 DVDD.n14610 0.019716
R42556 DVDD.n14620 DVDD.n8078 0.019716
R42557 DVDD.n14620 DVDD.n14619 0.019716
R42558 DVDD.n14622 DVDD.n8077 0.019716
R42559 DVDD.n14623 DVDD.n14622 0.019716
R42560 DVDD.n14632 DVDD.n8076 0.019716
R42561 DVDD.n14632 DVDD.n14631 0.019716
R42562 DVDD.n14634 DVDD.n8075 0.019716
R42563 DVDD.n14635 DVDD.n14634 0.019716
R42564 DVDD.n14644 DVDD.n8074 0.019716
R42565 DVDD.n14644 DVDD.n14643 0.019716
R42566 DVDD.n14646 DVDD.n8073 0.019716
R42567 DVDD.n14647 DVDD.n14646 0.019716
R42568 DVDD.n14656 DVDD.n8072 0.019716
R42569 DVDD.n14656 DVDD.n14655 0.019716
R42570 DVDD.n14658 DVDD.n8071 0.019716
R42571 DVDD.n14659 DVDD.n14658 0.019716
R42572 DVDD.n14668 DVDD.n8070 0.019716
R42573 DVDD.n14668 DVDD.n14667 0.019716
R42574 DVDD.n14670 DVDD.n8069 0.019716
R42575 DVDD.n14671 DVDD.n14670 0.019716
R42576 DVDD.n14680 DVDD.n8068 0.019716
R42577 DVDD.n14680 DVDD.n14679 0.019716
R42578 DVDD.n14682 DVDD.n8067 0.019716
R42579 DVDD.n14683 DVDD.n14682 0.019716
R42580 DVDD.n14692 DVDD.n8066 0.019716
R42581 DVDD.n14692 DVDD.n14691 0.019716
R42582 DVDD.n14694 DVDD.n8065 0.019716
R42583 DVDD.n14695 DVDD.n14694 0.019716
R42584 DVDD.n14704 DVDD.n8064 0.019716
R42585 DVDD.n14704 DVDD.n14703 0.019716
R42586 DVDD.n14706 DVDD.n8063 0.019716
R42587 DVDD.n14707 DVDD.n14706 0.019716
R42588 DVDD.n14716 DVDD.n8062 0.019716
R42589 DVDD.n14716 DVDD.n14715 0.019716
R42590 DVDD.n14718 DVDD.n8061 0.019716
R42591 DVDD.n14719 DVDD.n14718 0.019716
R42592 DVDD.n14728 DVDD.n8060 0.019716
R42593 DVDD.n14728 DVDD.n14727 0.019716
R42594 DVDD.n14730 DVDD.n8059 0.019716
R42595 DVDD.n14731 DVDD.n14730 0.019716
R42596 DVDD.n14740 DVDD.n8058 0.019716
R42597 DVDD.n14740 DVDD.n14739 0.019716
R42598 DVDD.n14742 DVDD.n8057 0.019716
R42599 DVDD.n14743 DVDD.n14742 0.019716
R42600 DVDD.n14752 DVDD.n8056 0.019716
R42601 DVDD.n14752 DVDD.n14751 0.019716
R42602 DVDD.n14754 DVDD.n8055 0.019716
R42603 DVDD.n14755 DVDD.n14754 0.019716
R42604 DVDD.n14764 DVDD.n8054 0.019716
R42605 DVDD.n14764 DVDD.n14763 0.019716
R42606 DVDD.n14766 DVDD.n8053 0.019716
R42607 DVDD.n14767 DVDD.n14766 0.019716
R42608 DVDD.n14776 DVDD.n8052 0.019716
R42609 DVDD.n14776 DVDD.n14775 0.019716
R42610 DVDD.n14778 DVDD.n8051 0.019716
R42611 DVDD.n14779 DVDD.n14778 0.019716
R42612 DVDD.n14788 DVDD.n8050 0.019716
R42613 DVDD.n14788 DVDD.n14787 0.019716
R42614 DVDD.n14790 DVDD.n8049 0.019716
R42615 DVDD.n14791 DVDD.n14790 0.019716
R42616 DVDD.n14800 DVDD.n8048 0.019716
R42617 DVDD.n14800 DVDD.n14799 0.019716
R42618 DVDD.n14802 DVDD.n8047 0.019716
R42619 DVDD.n14803 DVDD.n14802 0.019716
R42620 DVDD.n14812 DVDD.n8046 0.019716
R42621 DVDD.n14812 DVDD.n14811 0.019716
R42622 DVDD.n14814 DVDD.n8045 0.019716
R42623 DVDD.n14815 DVDD.n14814 0.019716
R42624 DVDD.n14824 DVDD.n14823 0.019716
R42625 DVDD.n14839 DVDD.n14838 0.019716
R42626 DVDD.n7774 DVDD.n7731 0.019716
R42627 DVDD.n7844 DVDD.n7773 0.019716
R42628 DVDD.n7844 DVDD.n7729 0.019716
R42629 DVDD.n7848 DVDD.n7772 0.019716
R42630 DVDD.n7848 DVDD.n7728 0.019716
R42631 DVDD.n7853 DVDD.n7771 0.019716
R42632 DVDD.n7853 DVDD.n7727 0.019716
R42633 DVDD.n7857 DVDD.n7770 0.019716
R42634 DVDD.n7857 DVDD.n7726 0.019716
R42635 DVDD.n7862 DVDD.n7769 0.019716
R42636 DVDD.n7862 DVDD.n7725 0.019716
R42637 DVDD.n7866 DVDD.n7768 0.019716
R42638 DVDD.n7866 DVDD.n7724 0.019716
R42639 DVDD.n7871 DVDD.n7767 0.019716
R42640 DVDD.n7871 DVDD.n7723 0.019716
R42641 DVDD.n7875 DVDD.n7766 0.019716
R42642 DVDD.n7875 DVDD.n7722 0.019716
R42643 DVDD.n7880 DVDD.n7765 0.019716
R42644 DVDD.n7880 DVDD.n7721 0.019716
R42645 DVDD.n7884 DVDD.n7764 0.019716
R42646 DVDD.n7884 DVDD.n7720 0.019716
R42647 DVDD.n7889 DVDD.n7763 0.019716
R42648 DVDD.n7889 DVDD.n7719 0.019716
R42649 DVDD.n7893 DVDD.n7762 0.019716
R42650 DVDD.n7893 DVDD.n7718 0.019716
R42651 DVDD.n7898 DVDD.n7761 0.019716
R42652 DVDD.n7898 DVDD.n7717 0.019716
R42653 DVDD.n7902 DVDD.n7760 0.019716
R42654 DVDD.n7902 DVDD.n7716 0.019716
R42655 DVDD.n7907 DVDD.n7759 0.019716
R42656 DVDD.n7907 DVDD.n7715 0.019716
R42657 DVDD.n7911 DVDD.n7758 0.019716
R42658 DVDD.n7911 DVDD.n7714 0.019716
R42659 DVDD.n7916 DVDD.n7757 0.019716
R42660 DVDD.n7916 DVDD.n7713 0.019716
R42661 DVDD.n7920 DVDD.n7756 0.019716
R42662 DVDD.n7920 DVDD.n7712 0.019716
R42663 DVDD.n7925 DVDD.n7755 0.019716
R42664 DVDD.n7925 DVDD.n7711 0.019716
R42665 DVDD.n7929 DVDD.n7754 0.019716
R42666 DVDD.n7929 DVDD.n7710 0.019716
R42667 DVDD.n7934 DVDD.n7753 0.019716
R42668 DVDD.n7934 DVDD.n7709 0.019716
R42669 DVDD.n7938 DVDD.n7752 0.019716
R42670 DVDD.n7938 DVDD.n7708 0.019716
R42671 DVDD.n7943 DVDD.n7751 0.019716
R42672 DVDD.n7943 DVDD.n7707 0.019716
R42673 DVDD.n7947 DVDD.n7750 0.019716
R42674 DVDD.n7947 DVDD.n7706 0.019716
R42675 DVDD.n7952 DVDD.n7749 0.019716
R42676 DVDD.n7952 DVDD.n7705 0.019716
R42677 DVDD.n7956 DVDD.n7748 0.019716
R42678 DVDD.n7956 DVDD.n7704 0.019716
R42679 DVDD.n7961 DVDD.n7747 0.019716
R42680 DVDD.n7961 DVDD.n7703 0.019716
R42681 DVDD.n7965 DVDD.n7746 0.019716
R42682 DVDD.n7965 DVDD.n7702 0.019716
R42683 DVDD.n7970 DVDD.n7745 0.019716
R42684 DVDD.n7970 DVDD.n7701 0.019716
R42685 DVDD.n7974 DVDD.n7744 0.019716
R42686 DVDD.n7974 DVDD.n7700 0.019716
R42687 DVDD.n7979 DVDD.n7743 0.019716
R42688 DVDD.n7979 DVDD.n7699 0.019716
R42689 DVDD.n7983 DVDD.n7742 0.019716
R42690 DVDD.n7983 DVDD.n7698 0.019716
R42691 DVDD.n7988 DVDD.n7741 0.019716
R42692 DVDD.n7988 DVDD.n7697 0.019716
R42693 DVDD.n7992 DVDD.n7740 0.019716
R42694 DVDD.n7992 DVDD.n7696 0.019716
R42695 DVDD.n7997 DVDD.n7739 0.019716
R42696 DVDD.n7997 DVDD.n7695 0.019716
R42697 DVDD.n8001 DVDD.n7738 0.019716
R42698 DVDD.n8001 DVDD.n7694 0.019716
R42699 DVDD.n8006 DVDD.n7737 0.019716
R42700 DVDD.n8006 DVDD.n7693 0.019716
R42701 DVDD.n8010 DVDD.n7736 0.019716
R42702 DVDD.n8010 DVDD.n7692 0.019716
R42703 DVDD.n8015 DVDD.n7735 0.019716
R42704 DVDD.n8015 DVDD.n7691 0.019716
R42705 DVDD.n8019 DVDD.n7734 0.019716
R42706 DVDD.n8019 DVDD.n7690 0.019716
R42707 DVDD.n14836 DVDD.n7689 0.019716
R42708 DVDD.n9557 DVDD.n9556 0.019716
R42709 DVDD.n9266 DVDD.n9264 0.019716
R42710 DVDD.n9549 DVDD.n9548 0.019716
R42711 DVDD.n9549 DVDD.n9263 0.019716
R42712 DVDD.n9544 DVDD.n9543 0.019716
R42713 DVDD.n9544 DVDD.n9262 0.019716
R42714 DVDD.n9537 DVDD.n9536 0.019716
R42715 DVDD.n9537 DVDD.n9261 0.019716
R42716 DVDD.n9532 DVDD.n9531 0.019716
R42717 DVDD.n9532 DVDD.n9260 0.019716
R42718 DVDD.n9525 DVDD.n9524 0.019716
R42719 DVDD.n9525 DVDD.n9259 0.019716
R42720 DVDD.n9520 DVDD.n9519 0.019716
R42721 DVDD.n9520 DVDD.n9258 0.019716
R42722 DVDD.n9513 DVDD.n9512 0.019716
R42723 DVDD.n9513 DVDD.n9257 0.019716
R42724 DVDD.n9508 DVDD.n9507 0.019716
R42725 DVDD.n9508 DVDD.n9256 0.019716
R42726 DVDD.n9501 DVDD.n9500 0.019716
R42727 DVDD.n9501 DVDD.n9255 0.019716
R42728 DVDD.n9496 DVDD.n9495 0.019716
R42729 DVDD.n9496 DVDD.n9254 0.019716
R42730 DVDD.n9489 DVDD.n9488 0.019716
R42731 DVDD.n9489 DVDD.n9253 0.019716
R42732 DVDD.n9484 DVDD.n9483 0.019716
R42733 DVDD.n9484 DVDD.n9252 0.019716
R42734 DVDD.n9477 DVDD.n9476 0.019716
R42735 DVDD.n9477 DVDD.n9251 0.019716
R42736 DVDD.n9472 DVDD.n9471 0.019716
R42737 DVDD.n9472 DVDD.n9250 0.019716
R42738 DVDD.n9465 DVDD.n9464 0.019716
R42739 DVDD.n9465 DVDD.n9249 0.019716
R42740 DVDD.n9460 DVDD.n9459 0.019716
R42741 DVDD.n9460 DVDD.n9248 0.019716
R42742 DVDD.n9453 DVDD.n9452 0.019716
R42743 DVDD.n9453 DVDD.n9247 0.019716
R42744 DVDD.n9448 DVDD.n9447 0.019716
R42745 DVDD.n9448 DVDD.n9246 0.019716
R42746 DVDD.n9441 DVDD.n9440 0.019716
R42747 DVDD.n9441 DVDD.n9245 0.019716
R42748 DVDD.n9436 DVDD.n9435 0.019716
R42749 DVDD.n9436 DVDD.n9244 0.019716
R42750 DVDD.n9429 DVDD.n9428 0.019716
R42751 DVDD.n9429 DVDD.n9243 0.019716
R42752 DVDD.n9424 DVDD.n9423 0.019716
R42753 DVDD.n9424 DVDD.n9242 0.019716
R42754 DVDD.n9417 DVDD.n9416 0.019716
R42755 DVDD.n9417 DVDD.n9241 0.019716
R42756 DVDD.n9412 DVDD.n9411 0.019716
R42757 DVDD.n9412 DVDD.n9240 0.019716
R42758 DVDD.n9405 DVDD.n9404 0.019716
R42759 DVDD.n9405 DVDD.n9239 0.019716
R42760 DVDD.n9400 DVDD.n9399 0.019716
R42761 DVDD.n9400 DVDD.n9238 0.019716
R42762 DVDD.n9393 DVDD.n9392 0.019716
R42763 DVDD.n9393 DVDD.n9237 0.019716
R42764 DVDD.n9388 DVDD.n9387 0.019716
R42765 DVDD.n9388 DVDD.n9236 0.019716
R42766 DVDD.n9381 DVDD.n9380 0.019716
R42767 DVDD.n9381 DVDD.n9235 0.019716
R42768 DVDD.n9376 DVDD.n9375 0.019716
R42769 DVDD.n9376 DVDD.n9234 0.019716
R42770 DVDD.n9369 DVDD.n9368 0.019716
R42771 DVDD.n9369 DVDD.n9233 0.019716
R42772 DVDD.n9364 DVDD.n9363 0.019716
R42773 DVDD.n9364 DVDD.n9232 0.019716
R42774 DVDD.n9357 DVDD.n9356 0.019716
R42775 DVDD.n9357 DVDD.n9231 0.019716
R42776 DVDD.n9352 DVDD.n9351 0.019716
R42777 DVDD.n9352 DVDD.n9230 0.019716
R42778 DVDD.n9345 DVDD.n9344 0.019716
R42779 DVDD.n9345 DVDD.n9229 0.019716
R42780 DVDD.n9340 DVDD.n9339 0.019716
R42781 DVDD.n9340 DVDD.n9228 0.019716
R42782 DVDD.n9333 DVDD.n9332 0.019716
R42783 DVDD.n9333 DVDD.n9227 0.019716
R42784 DVDD.n9328 DVDD.n9327 0.019716
R42785 DVDD.n9328 DVDD.n9226 0.019716
R42786 DVDD.n9321 DVDD.n9320 0.019716
R42787 DVDD.n9321 DVDD.n9225 0.019716
R42788 DVDD.n9316 DVDD.n9315 0.019716
R42789 DVDD.n9316 DVDD.n9224 0.019716
R42790 DVDD.n9309 DVDD.n9223 0.019716
R42791 DVDD.n14862 DVDD.n14861 0.019716
R42792 DVDD.n7656 DVDD.n7612 0.019716
R42793 DVDD.n9212 DVDD.n7655 0.019716
R42794 DVDD.n9212 DVDD.n7610 0.019716
R42795 DVDD.n9207 DVDD.n7654 0.019716
R42796 DVDD.n9207 DVDD.n7609 0.019716
R42797 DVDD.n9203 DVDD.n7653 0.019716
R42798 DVDD.n9203 DVDD.n7608 0.019716
R42799 DVDD.n9198 DVDD.n7652 0.019716
R42800 DVDD.n9198 DVDD.n7607 0.019716
R42801 DVDD.n9194 DVDD.n7651 0.019716
R42802 DVDD.n9194 DVDD.n7606 0.019716
R42803 DVDD.n9189 DVDD.n7650 0.019716
R42804 DVDD.n9189 DVDD.n7605 0.019716
R42805 DVDD.n9185 DVDD.n7649 0.019716
R42806 DVDD.n9185 DVDD.n7604 0.019716
R42807 DVDD.n9180 DVDD.n7648 0.019716
R42808 DVDD.n9180 DVDD.n7603 0.019716
R42809 DVDD.n9176 DVDD.n7647 0.019716
R42810 DVDD.n9176 DVDD.n7602 0.019716
R42811 DVDD.n9171 DVDD.n7646 0.019716
R42812 DVDD.n9171 DVDD.n7601 0.019716
R42813 DVDD.n9167 DVDD.n7645 0.019716
R42814 DVDD.n9167 DVDD.n7600 0.019716
R42815 DVDD.n9162 DVDD.n7644 0.019716
R42816 DVDD.n9162 DVDD.n7599 0.019716
R42817 DVDD.n9158 DVDD.n7643 0.019716
R42818 DVDD.n9158 DVDD.n7598 0.019716
R42819 DVDD.n9153 DVDD.n7642 0.019716
R42820 DVDD.n9153 DVDD.n7597 0.019716
R42821 DVDD.n9149 DVDD.n7641 0.019716
R42822 DVDD.n9149 DVDD.n7596 0.019716
R42823 DVDD.n9144 DVDD.n7640 0.019716
R42824 DVDD.n9144 DVDD.n7595 0.019716
R42825 DVDD.n9140 DVDD.n7639 0.019716
R42826 DVDD.n9140 DVDD.n7594 0.019716
R42827 DVDD.n9135 DVDD.n7638 0.019716
R42828 DVDD.n9135 DVDD.n7593 0.019716
R42829 DVDD.n9131 DVDD.n7637 0.019716
R42830 DVDD.n9131 DVDD.n7592 0.019716
R42831 DVDD.n9126 DVDD.n7636 0.019716
R42832 DVDD.n9126 DVDD.n7591 0.019716
R42833 DVDD.n9122 DVDD.n7635 0.019716
R42834 DVDD.n9122 DVDD.n7590 0.019716
R42835 DVDD.n9117 DVDD.n7634 0.019716
R42836 DVDD.n9117 DVDD.n7589 0.019716
R42837 DVDD.n9113 DVDD.n7633 0.019716
R42838 DVDD.n9113 DVDD.n7588 0.019716
R42839 DVDD.n9108 DVDD.n7632 0.019716
R42840 DVDD.n9108 DVDD.n7587 0.019716
R42841 DVDD.n9104 DVDD.n7631 0.019716
R42842 DVDD.n9104 DVDD.n7586 0.019716
R42843 DVDD.n9099 DVDD.n7630 0.019716
R42844 DVDD.n9099 DVDD.n7585 0.019716
R42845 DVDD.n9095 DVDD.n7629 0.019716
R42846 DVDD.n9095 DVDD.n7584 0.019716
R42847 DVDD.n9090 DVDD.n7628 0.019716
R42848 DVDD.n9090 DVDD.n7583 0.019716
R42849 DVDD.n9086 DVDD.n7627 0.019716
R42850 DVDD.n9086 DVDD.n7582 0.019716
R42851 DVDD.n9081 DVDD.n7626 0.019716
R42852 DVDD.n9081 DVDD.n7581 0.019716
R42853 DVDD.n9077 DVDD.n7625 0.019716
R42854 DVDD.n9077 DVDD.n7580 0.019716
R42855 DVDD.n9072 DVDD.n7624 0.019716
R42856 DVDD.n9072 DVDD.n7579 0.019716
R42857 DVDD.n9068 DVDD.n7623 0.019716
R42858 DVDD.n9068 DVDD.n7578 0.019716
R42859 DVDD.n9063 DVDD.n7622 0.019716
R42860 DVDD.n9063 DVDD.n7577 0.019716
R42861 DVDD.n9059 DVDD.n7621 0.019716
R42862 DVDD.n9059 DVDD.n7576 0.019716
R42863 DVDD.n9054 DVDD.n7620 0.019716
R42864 DVDD.n9054 DVDD.n7575 0.019716
R42865 DVDD.n9050 DVDD.n7619 0.019716
R42866 DVDD.n9050 DVDD.n7574 0.019716
R42867 DVDD.n9045 DVDD.n7618 0.019716
R42868 DVDD.n9045 DVDD.n7573 0.019716
R42869 DVDD.n9041 DVDD.n7617 0.019716
R42870 DVDD.n9041 DVDD.n7572 0.019716
R42871 DVDD.n9036 DVDD.n7616 0.019716
R42872 DVDD.n9036 DVDD.n7571 0.019716
R42873 DVDD.n14859 DVDD.n7570 0.019716
R42874 DVDD.n15059 DVDD.n15058 0.019716
R42875 DVDD.n7499 DVDD.n7455 0.019716
R42876 DVDD.n14875 DVDD.n7498 0.019716
R42877 DVDD.n14875 DVDD.n7453 0.019716
R42878 DVDD.n14879 DVDD.n7497 0.019716
R42879 DVDD.n14879 DVDD.n7452 0.019716
R42880 DVDD.n14884 DVDD.n7496 0.019716
R42881 DVDD.n14884 DVDD.n7451 0.019716
R42882 DVDD.n14888 DVDD.n7495 0.019716
R42883 DVDD.n14888 DVDD.n7450 0.019716
R42884 DVDD.n14893 DVDD.n7494 0.019716
R42885 DVDD.n14893 DVDD.n7449 0.019716
R42886 DVDD.n14897 DVDD.n7493 0.019716
R42887 DVDD.n14897 DVDD.n7448 0.019716
R42888 DVDD.n14902 DVDD.n7492 0.019716
R42889 DVDD.n14902 DVDD.n7447 0.019716
R42890 DVDD.n14906 DVDD.n7491 0.019716
R42891 DVDD.n14906 DVDD.n7446 0.019716
R42892 DVDD.n14911 DVDD.n7490 0.019716
R42893 DVDD.n14911 DVDD.n7445 0.019716
R42894 DVDD.n14915 DVDD.n7489 0.019716
R42895 DVDD.n14915 DVDD.n7444 0.019716
R42896 DVDD.n14920 DVDD.n7488 0.019716
R42897 DVDD.n14920 DVDD.n7443 0.019716
R42898 DVDD.n14924 DVDD.n7487 0.019716
R42899 DVDD.n14924 DVDD.n7442 0.019716
R42900 DVDD.n14929 DVDD.n7486 0.019716
R42901 DVDD.n14929 DVDD.n7441 0.019716
R42902 DVDD.n14933 DVDD.n7485 0.019716
R42903 DVDD.n14933 DVDD.n7440 0.019716
R42904 DVDD.n14938 DVDD.n7484 0.019716
R42905 DVDD.n14938 DVDD.n7439 0.019716
R42906 DVDD.n14942 DVDD.n7483 0.019716
R42907 DVDD.n14942 DVDD.n7438 0.019716
R42908 DVDD.n14947 DVDD.n7482 0.019716
R42909 DVDD.n14947 DVDD.n7437 0.019716
R42910 DVDD.n14951 DVDD.n7481 0.019716
R42911 DVDD.n14951 DVDD.n7436 0.019716
R42912 DVDD.n14956 DVDD.n7480 0.019716
R42913 DVDD.n14956 DVDD.n7435 0.019716
R42914 DVDD.n14960 DVDD.n7479 0.019716
R42915 DVDD.n14960 DVDD.n7434 0.019716
R42916 DVDD.n14965 DVDD.n7478 0.019716
R42917 DVDD.n14965 DVDD.n7433 0.019716
R42918 DVDD.n14969 DVDD.n7477 0.019716
R42919 DVDD.n14969 DVDD.n7432 0.019716
R42920 DVDD.n14974 DVDD.n7476 0.019716
R42921 DVDD.n14974 DVDD.n7431 0.019716
R42922 DVDD.n14978 DVDD.n7475 0.019716
R42923 DVDD.n14978 DVDD.n7430 0.019716
R42924 DVDD.n14983 DVDD.n7474 0.019716
R42925 DVDD.n14983 DVDD.n7429 0.019716
R42926 DVDD.n14987 DVDD.n7473 0.019716
R42927 DVDD.n14987 DVDD.n7428 0.019716
R42928 DVDD.n14992 DVDD.n7472 0.019716
R42929 DVDD.n14992 DVDD.n7427 0.019716
R42930 DVDD.n14996 DVDD.n7471 0.019716
R42931 DVDD.n14996 DVDD.n7426 0.019716
R42932 DVDD.n15001 DVDD.n7470 0.019716
R42933 DVDD.n15001 DVDD.n7425 0.019716
R42934 DVDD.n15005 DVDD.n7469 0.019716
R42935 DVDD.n15005 DVDD.n7424 0.019716
R42936 DVDD.n15010 DVDD.n7468 0.019716
R42937 DVDD.n15010 DVDD.n7423 0.019716
R42938 DVDD.n15014 DVDD.n7467 0.019716
R42939 DVDD.n15014 DVDD.n7422 0.019716
R42940 DVDD.n15019 DVDD.n7466 0.019716
R42941 DVDD.n15019 DVDD.n7421 0.019716
R42942 DVDD.n15023 DVDD.n7465 0.019716
R42943 DVDD.n15023 DVDD.n7420 0.019716
R42944 DVDD.n15028 DVDD.n7464 0.019716
R42945 DVDD.n15028 DVDD.n7419 0.019716
R42946 DVDD.n15032 DVDD.n7463 0.019716
R42947 DVDD.n15032 DVDD.n7418 0.019716
R42948 DVDD.n15037 DVDD.n7462 0.019716
R42949 DVDD.n15037 DVDD.n7417 0.019716
R42950 DVDD.n15041 DVDD.n7461 0.019716
R42951 DVDD.n15041 DVDD.n7416 0.019716
R42952 DVDD.n15046 DVDD.n7460 0.019716
R42953 DVDD.n15046 DVDD.n7415 0.019716
R42954 DVDD.n15050 DVDD.n7459 0.019716
R42955 DVDD.n15050 DVDD.n7414 0.019716
R42956 DVDD.n15056 DVDD.n7413 0.019716
R42957 DVDD.n7154 DVDD.n7111 0.019716
R42958 DVDD.n7155 DVDD.n7110 0.019716
R42959 DVDD.n7162 DVDD.n7109 0.019716
R42960 DVDD.n7162 DVDD.n7161 0.019716
R42961 DVDD.n7164 DVDD.n7108 0.019716
R42962 DVDD.n7165 DVDD.n7164 0.019716
R42963 DVDD.n7174 DVDD.n7107 0.019716
R42964 DVDD.n7174 DVDD.n7173 0.019716
R42965 DVDD.n7176 DVDD.n7106 0.019716
R42966 DVDD.n7177 DVDD.n7176 0.019716
R42967 DVDD.n7186 DVDD.n7105 0.019716
R42968 DVDD.n7186 DVDD.n7185 0.019716
R42969 DVDD.n7188 DVDD.n7104 0.019716
R42970 DVDD.n7189 DVDD.n7188 0.019716
R42971 DVDD.n7198 DVDD.n7103 0.019716
R42972 DVDD.n7198 DVDD.n7197 0.019716
R42973 DVDD.n7200 DVDD.n7102 0.019716
R42974 DVDD.n7201 DVDD.n7200 0.019716
R42975 DVDD.n7210 DVDD.n7101 0.019716
R42976 DVDD.n7210 DVDD.n7209 0.019716
R42977 DVDD.n7212 DVDD.n7100 0.019716
R42978 DVDD.n7213 DVDD.n7212 0.019716
R42979 DVDD.n7222 DVDD.n7099 0.019716
R42980 DVDD.n7222 DVDD.n7221 0.019716
R42981 DVDD.n7224 DVDD.n7098 0.019716
R42982 DVDD.n7225 DVDD.n7224 0.019716
R42983 DVDD.n7234 DVDD.n7097 0.019716
R42984 DVDD.n7234 DVDD.n7233 0.019716
R42985 DVDD.n7236 DVDD.n7096 0.019716
R42986 DVDD.n7237 DVDD.n7236 0.019716
R42987 DVDD.n7246 DVDD.n7095 0.019716
R42988 DVDD.n7246 DVDD.n7245 0.019716
R42989 DVDD.n7248 DVDD.n7094 0.019716
R42990 DVDD.n7249 DVDD.n7248 0.019716
R42991 DVDD.n7258 DVDD.n7093 0.019716
R42992 DVDD.n7258 DVDD.n7257 0.019716
R42993 DVDD.n7260 DVDD.n7092 0.019716
R42994 DVDD.n7261 DVDD.n7260 0.019716
R42995 DVDD.n7270 DVDD.n7091 0.019716
R42996 DVDD.n7270 DVDD.n7269 0.019716
R42997 DVDD.n7272 DVDD.n7090 0.019716
R42998 DVDD.n7273 DVDD.n7272 0.019716
R42999 DVDD.n7282 DVDD.n7089 0.019716
R43000 DVDD.n7282 DVDD.n7281 0.019716
R43001 DVDD.n7284 DVDD.n7088 0.019716
R43002 DVDD.n7285 DVDD.n7284 0.019716
R43003 DVDD.n7294 DVDD.n7087 0.019716
R43004 DVDD.n7294 DVDD.n7293 0.019716
R43005 DVDD.n7296 DVDD.n7086 0.019716
R43006 DVDD.n7297 DVDD.n7296 0.019716
R43007 DVDD.n7306 DVDD.n7085 0.019716
R43008 DVDD.n7306 DVDD.n7305 0.019716
R43009 DVDD.n7308 DVDD.n7084 0.019716
R43010 DVDD.n7309 DVDD.n7308 0.019716
R43011 DVDD.n7318 DVDD.n7083 0.019716
R43012 DVDD.n7318 DVDD.n7317 0.019716
R43013 DVDD.n7320 DVDD.n7082 0.019716
R43014 DVDD.n7321 DVDD.n7320 0.019716
R43015 DVDD.n7330 DVDD.n7081 0.019716
R43016 DVDD.n7330 DVDD.n7329 0.019716
R43017 DVDD.n7332 DVDD.n7080 0.019716
R43018 DVDD.n7333 DVDD.n7332 0.019716
R43019 DVDD.n7342 DVDD.n7079 0.019716
R43020 DVDD.n7342 DVDD.n7341 0.019716
R43021 DVDD.n7344 DVDD.n7078 0.019716
R43022 DVDD.n7345 DVDD.n7344 0.019716
R43023 DVDD.n7354 DVDD.n7077 0.019716
R43024 DVDD.n7354 DVDD.n7353 0.019716
R43025 DVDD.n7356 DVDD.n7076 0.019716
R43026 DVDD.n7357 DVDD.n7356 0.019716
R43027 DVDD.n7366 DVDD.n7075 0.019716
R43028 DVDD.n7366 DVDD.n7365 0.019716
R43029 DVDD.n7368 DVDD.n7074 0.019716
R43030 DVDD.n7369 DVDD.n7368 0.019716
R43031 DVDD.n7378 DVDD.n7073 0.019716
R43032 DVDD.n7378 DVDD.n7377 0.019716
R43033 DVDD.n7380 DVDD.n7072 0.019716
R43034 DVDD.n7381 DVDD.n7380 0.019716
R43035 DVDD.n7390 DVDD.n7071 0.019716
R43036 DVDD.n7390 DVDD.n7389 0.019716
R43037 DVDD.n7392 DVDD.n7070 0.019716
R43038 DVDD.n7393 DVDD.n7392 0.019716
R43039 DVDD.n7403 DVDD.n7402 0.019716
R43040 DVDD.n15091 DVDD.n15090 0.019716
R43041 DVDD.n6793 DVDD.n6750 0.019716
R43042 DVDD.n6863 DVDD.n6792 0.019716
R43043 DVDD.n6863 DVDD.n6748 0.019716
R43044 DVDD.n6867 DVDD.n6791 0.019716
R43045 DVDD.n6867 DVDD.n6747 0.019716
R43046 DVDD.n6872 DVDD.n6790 0.019716
R43047 DVDD.n6872 DVDD.n6746 0.019716
R43048 DVDD.n6876 DVDD.n6789 0.019716
R43049 DVDD.n6876 DVDD.n6745 0.019716
R43050 DVDD.n6881 DVDD.n6788 0.019716
R43051 DVDD.n6881 DVDD.n6744 0.019716
R43052 DVDD.n6885 DVDD.n6787 0.019716
R43053 DVDD.n6885 DVDD.n6743 0.019716
R43054 DVDD.n6890 DVDD.n6786 0.019716
R43055 DVDD.n6890 DVDD.n6742 0.019716
R43056 DVDD.n6894 DVDD.n6785 0.019716
R43057 DVDD.n6894 DVDD.n6741 0.019716
R43058 DVDD.n6899 DVDD.n6784 0.019716
R43059 DVDD.n6899 DVDD.n6740 0.019716
R43060 DVDD.n6903 DVDD.n6783 0.019716
R43061 DVDD.n6903 DVDD.n6739 0.019716
R43062 DVDD.n6908 DVDD.n6782 0.019716
R43063 DVDD.n6908 DVDD.n6738 0.019716
R43064 DVDD.n6912 DVDD.n6781 0.019716
R43065 DVDD.n6912 DVDD.n6737 0.019716
R43066 DVDD.n6917 DVDD.n6780 0.019716
R43067 DVDD.n6917 DVDD.n6736 0.019716
R43068 DVDD.n6921 DVDD.n6779 0.019716
R43069 DVDD.n6921 DVDD.n6735 0.019716
R43070 DVDD.n6926 DVDD.n6778 0.019716
R43071 DVDD.n6926 DVDD.n6734 0.019716
R43072 DVDD.n6930 DVDD.n6777 0.019716
R43073 DVDD.n6930 DVDD.n6733 0.019716
R43074 DVDD.n6935 DVDD.n6776 0.019716
R43075 DVDD.n6935 DVDD.n6732 0.019716
R43076 DVDD.n6939 DVDD.n6775 0.019716
R43077 DVDD.n6939 DVDD.n6731 0.019716
R43078 DVDD.n6944 DVDD.n6774 0.019716
R43079 DVDD.n6944 DVDD.n6730 0.019716
R43080 DVDD.n6948 DVDD.n6773 0.019716
R43081 DVDD.n6948 DVDD.n6729 0.019716
R43082 DVDD.n6953 DVDD.n6772 0.019716
R43083 DVDD.n6953 DVDD.n6728 0.019716
R43084 DVDD.n6957 DVDD.n6771 0.019716
R43085 DVDD.n6957 DVDD.n6727 0.019716
R43086 DVDD.n6962 DVDD.n6770 0.019716
R43087 DVDD.n6962 DVDD.n6726 0.019716
R43088 DVDD.n6966 DVDD.n6769 0.019716
R43089 DVDD.n6966 DVDD.n6725 0.019716
R43090 DVDD.n6971 DVDD.n6768 0.019716
R43091 DVDD.n6971 DVDD.n6724 0.019716
R43092 DVDD.n6975 DVDD.n6767 0.019716
R43093 DVDD.n6975 DVDD.n6723 0.019716
R43094 DVDD.n6980 DVDD.n6766 0.019716
R43095 DVDD.n6980 DVDD.n6722 0.019716
R43096 DVDD.n6984 DVDD.n6765 0.019716
R43097 DVDD.n6984 DVDD.n6721 0.019716
R43098 DVDD.n6989 DVDD.n6764 0.019716
R43099 DVDD.n6989 DVDD.n6720 0.019716
R43100 DVDD.n6993 DVDD.n6763 0.019716
R43101 DVDD.n6993 DVDD.n6719 0.019716
R43102 DVDD.n6998 DVDD.n6762 0.019716
R43103 DVDD.n6998 DVDD.n6718 0.019716
R43104 DVDD.n7002 DVDD.n6761 0.019716
R43105 DVDD.n7002 DVDD.n6717 0.019716
R43106 DVDD.n7007 DVDD.n6760 0.019716
R43107 DVDD.n7007 DVDD.n6716 0.019716
R43108 DVDD.n7011 DVDD.n6759 0.019716
R43109 DVDD.n7011 DVDD.n6715 0.019716
R43110 DVDD.n7016 DVDD.n6758 0.019716
R43111 DVDD.n7016 DVDD.n6714 0.019716
R43112 DVDD.n7020 DVDD.n6757 0.019716
R43113 DVDD.n7020 DVDD.n6713 0.019716
R43114 DVDD.n7025 DVDD.n6756 0.019716
R43115 DVDD.n7025 DVDD.n6712 0.019716
R43116 DVDD.n7029 DVDD.n6755 0.019716
R43117 DVDD.n7029 DVDD.n6711 0.019716
R43118 DVDD.n7034 DVDD.n6754 0.019716
R43119 DVDD.n7034 DVDD.n6710 0.019716
R43120 DVDD.n7038 DVDD.n6753 0.019716
R43121 DVDD.n7038 DVDD.n6709 0.019716
R43122 DVDD.n15088 DVDD.n6708 0.019716
R43123 DVDD.n6509 DVDD.n6390 0.019716
R43124 DVDD.n6509 DVDD.n6405 0.019716
R43125 DVDD.n6514 DVDD.n6389 0.019716
R43126 DVDD.n6514 DVDD.n6406 0.019716
R43127 DVDD.n6518 DVDD.n6388 0.019716
R43128 DVDD.n6518 DVDD.n6407 0.019716
R43129 DVDD.n6523 DVDD.n6387 0.019716
R43130 DVDD.n6523 DVDD.n6408 0.019716
R43131 DVDD.n6527 DVDD.n6386 0.019716
R43132 DVDD.n6527 DVDD.n6409 0.019716
R43133 DVDD.n6532 DVDD.n6385 0.019716
R43134 DVDD.n6532 DVDD.n6410 0.019716
R43135 DVDD.n6536 DVDD.n6384 0.019716
R43136 DVDD.n6536 DVDD.n6411 0.019716
R43137 DVDD.n6541 DVDD.n6383 0.019716
R43138 DVDD.n6541 DVDD.n6412 0.019716
R43139 DVDD.n6545 DVDD.n6382 0.019716
R43140 DVDD.n6545 DVDD.n6413 0.019716
R43141 DVDD.n6550 DVDD.n6381 0.019716
R43142 DVDD.n6550 DVDD.n6414 0.019716
R43143 DVDD.n6554 DVDD.n6380 0.019716
R43144 DVDD.n6554 DVDD.n6415 0.019716
R43145 DVDD.n6559 DVDD.n6379 0.019716
R43146 DVDD.n6559 DVDD.n6416 0.019716
R43147 DVDD.n6563 DVDD.n6378 0.019716
R43148 DVDD.n6563 DVDD.n6417 0.019716
R43149 DVDD.n6568 DVDD.n6377 0.019716
R43150 DVDD.n6568 DVDD.n6418 0.019716
R43151 DVDD.n6572 DVDD.n6376 0.019716
R43152 DVDD.n6572 DVDD.n6419 0.019716
R43153 DVDD.n6577 DVDD.n6375 0.019716
R43154 DVDD.n6577 DVDD.n6420 0.019716
R43155 DVDD.n6581 DVDD.n6374 0.019716
R43156 DVDD.n6581 DVDD.n6421 0.019716
R43157 DVDD.n6586 DVDD.n6373 0.019716
R43158 DVDD.n6586 DVDD.n6422 0.019716
R43159 DVDD.n6590 DVDD.n6372 0.019716
R43160 DVDD.n6590 DVDD.n6423 0.019716
R43161 DVDD.n6595 DVDD.n6371 0.019716
R43162 DVDD.n6595 DVDD.n6424 0.019716
R43163 DVDD.n6599 DVDD.n6370 0.019716
R43164 DVDD.n6599 DVDD.n6425 0.019716
R43165 DVDD.n6604 DVDD.n6369 0.019716
R43166 DVDD.n6604 DVDD.n6426 0.019716
R43167 DVDD.n6608 DVDD.n6368 0.019716
R43168 DVDD.n6608 DVDD.n6427 0.019716
R43169 DVDD.n6613 DVDD.n6367 0.019716
R43170 DVDD.n6613 DVDD.n6428 0.019716
R43171 DVDD.n6617 DVDD.n6366 0.019716
R43172 DVDD.n6617 DVDD.n6429 0.019716
R43173 DVDD.n6622 DVDD.n6365 0.019716
R43174 DVDD.n6622 DVDD.n6430 0.019716
R43175 DVDD.n6626 DVDD.n6364 0.019716
R43176 DVDD.n6626 DVDD.n6431 0.019716
R43177 DVDD.n6631 DVDD.n6363 0.019716
R43178 DVDD.n6631 DVDD.n6432 0.019716
R43179 DVDD.n6635 DVDD.n6362 0.019716
R43180 DVDD.n6635 DVDD.n6433 0.019716
R43181 DVDD.n6640 DVDD.n6361 0.019716
R43182 DVDD.n6640 DVDD.n6434 0.019716
R43183 DVDD.n6644 DVDD.n6360 0.019716
R43184 DVDD.n6644 DVDD.n6435 0.019716
R43185 DVDD.n6649 DVDD.n6359 0.019716
R43186 DVDD.n6649 DVDD.n6436 0.019716
R43187 DVDD.n6653 DVDD.n6358 0.019716
R43188 DVDD.n6653 DVDD.n6437 0.019716
R43189 DVDD.n6658 DVDD.n6357 0.019716
R43190 DVDD.n6658 DVDD.n6438 0.019716
R43191 DVDD.n6662 DVDD.n6356 0.019716
R43192 DVDD.n6662 DVDD.n6439 0.019716
R43193 DVDD.n6667 DVDD.n6355 0.019716
R43194 DVDD.n6667 DVDD.n6440 0.019716
R43195 DVDD.n6671 DVDD.n6354 0.019716
R43196 DVDD.n6671 DVDD.n6441 0.019716
R43197 DVDD.n6676 DVDD.n6353 0.019716
R43198 DVDD.n6676 DVDD.n6442 0.019716
R43199 DVDD.n6680 DVDD.n6352 0.019716
R43200 DVDD.n6680 DVDD.n6443 0.019716
R43201 DVDD.n6685 DVDD.n6351 0.019716
R43202 DVDD.n6685 DVDD.n6444 0.019716
R43203 DVDD.n6689 DVDD.n6350 0.019716
R43204 DVDD.n6689 DVDD.n6445 0.019716
R43205 DVDD.n6695 DVDD.n6349 0.019716
R43206 DVDD.n6404 DVDD.n6390 0.019716
R43207 DVDD.n6506 DVDD.n6389 0.019716
R43208 DVDD.n6506 DVDD.n6405 0.019716
R43209 DVDD.n6516 DVDD.n6388 0.019716
R43210 DVDD.n6516 DVDD.n6406 0.019716
R43211 DVDD.n6503 DVDD.n6387 0.019716
R43212 DVDD.n6503 DVDD.n6407 0.019716
R43213 DVDD.n6525 DVDD.n6386 0.019716
R43214 DVDD.n6525 DVDD.n6408 0.019716
R43215 DVDD.n6500 DVDD.n6385 0.019716
R43216 DVDD.n6500 DVDD.n6409 0.019716
R43217 DVDD.n6534 DVDD.n6384 0.019716
R43218 DVDD.n6534 DVDD.n6410 0.019716
R43219 DVDD.n6497 DVDD.n6383 0.019716
R43220 DVDD.n6497 DVDD.n6411 0.019716
R43221 DVDD.n6543 DVDD.n6382 0.019716
R43222 DVDD.n6543 DVDD.n6412 0.019716
R43223 DVDD.n6494 DVDD.n6381 0.019716
R43224 DVDD.n6494 DVDD.n6413 0.019716
R43225 DVDD.n6552 DVDD.n6380 0.019716
R43226 DVDD.n6552 DVDD.n6414 0.019716
R43227 DVDD.n6491 DVDD.n6379 0.019716
R43228 DVDD.n6491 DVDD.n6415 0.019716
R43229 DVDD.n6561 DVDD.n6378 0.019716
R43230 DVDD.n6561 DVDD.n6416 0.019716
R43231 DVDD.n6488 DVDD.n6377 0.019716
R43232 DVDD.n6488 DVDD.n6417 0.019716
R43233 DVDD.n6570 DVDD.n6376 0.019716
R43234 DVDD.n6570 DVDD.n6418 0.019716
R43235 DVDD.n6485 DVDD.n6375 0.019716
R43236 DVDD.n6485 DVDD.n6419 0.019716
R43237 DVDD.n6579 DVDD.n6374 0.019716
R43238 DVDD.n6579 DVDD.n6420 0.019716
R43239 DVDD.n6482 DVDD.n6373 0.019716
R43240 DVDD.n6482 DVDD.n6421 0.019716
R43241 DVDD.n6588 DVDD.n6372 0.019716
R43242 DVDD.n6588 DVDD.n6422 0.019716
R43243 DVDD.n6479 DVDD.n6371 0.019716
R43244 DVDD.n6479 DVDD.n6423 0.019716
R43245 DVDD.n6597 DVDD.n6370 0.019716
R43246 DVDD.n6597 DVDD.n6424 0.019716
R43247 DVDD.n6476 DVDD.n6369 0.019716
R43248 DVDD.n6476 DVDD.n6425 0.019716
R43249 DVDD.n6606 DVDD.n6368 0.019716
R43250 DVDD.n6606 DVDD.n6426 0.019716
R43251 DVDD.n6473 DVDD.n6367 0.019716
R43252 DVDD.n6473 DVDD.n6427 0.019716
R43253 DVDD.n6615 DVDD.n6366 0.019716
R43254 DVDD.n6615 DVDD.n6428 0.019716
R43255 DVDD.n6470 DVDD.n6365 0.019716
R43256 DVDD.n6470 DVDD.n6429 0.019716
R43257 DVDD.n6624 DVDD.n6364 0.019716
R43258 DVDD.n6624 DVDD.n6430 0.019716
R43259 DVDD.n6467 DVDD.n6363 0.019716
R43260 DVDD.n6467 DVDD.n6431 0.019716
R43261 DVDD.n6633 DVDD.n6362 0.019716
R43262 DVDD.n6633 DVDD.n6432 0.019716
R43263 DVDD.n6464 DVDD.n6361 0.019716
R43264 DVDD.n6464 DVDD.n6433 0.019716
R43265 DVDD.n6642 DVDD.n6360 0.019716
R43266 DVDD.n6642 DVDD.n6434 0.019716
R43267 DVDD.n6461 DVDD.n6359 0.019716
R43268 DVDD.n6461 DVDD.n6435 0.019716
R43269 DVDD.n6651 DVDD.n6358 0.019716
R43270 DVDD.n6651 DVDD.n6436 0.019716
R43271 DVDD.n6458 DVDD.n6357 0.019716
R43272 DVDD.n6458 DVDD.n6437 0.019716
R43273 DVDD.n6660 DVDD.n6356 0.019716
R43274 DVDD.n6660 DVDD.n6438 0.019716
R43275 DVDD.n6455 DVDD.n6355 0.019716
R43276 DVDD.n6455 DVDD.n6439 0.019716
R43277 DVDD.n6669 DVDD.n6354 0.019716
R43278 DVDD.n6669 DVDD.n6440 0.019716
R43279 DVDD.n6452 DVDD.n6353 0.019716
R43280 DVDD.n6452 DVDD.n6441 0.019716
R43281 DVDD.n6678 DVDD.n6352 0.019716
R43282 DVDD.n6678 DVDD.n6442 0.019716
R43283 DVDD.n6449 DVDD.n6351 0.019716
R43284 DVDD.n6449 DVDD.n6443 0.019716
R43285 DVDD.n6687 DVDD.n6350 0.019716
R43286 DVDD.n6687 DVDD.n6444 0.019716
R43287 DVDD.n6446 DVDD.n6349 0.019716
R43288 DVDD.n6446 DVDD.n6445 0.019716
R43289 DVDD.n1255 DVDD.n963 0.019716
R43290 DVDD.n966 DVDD.n964 0.019716
R43291 DVDD.n966 DVDD.n962 0.019716
R43292 DVDD.n1247 DVDD.n1246 0.019716
R43293 DVDD.n1246 DVDD.n961 0.019716
R43294 DVDD.n971 DVDD.n970 0.019716
R43295 DVDD.n970 DVDD.n960 0.019716
R43296 DVDD.n1238 DVDD.n1237 0.019716
R43297 DVDD.n1237 DVDD.n959 0.019716
R43298 DVDD.n976 DVDD.n975 0.019716
R43299 DVDD.n975 DVDD.n958 0.019716
R43300 DVDD.n1229 DVDD.n1228 0.019716
R43301 DVDD.n1228 DVDD.n957 0.019716
R43302 DVDD.n981 DVDD.n980 0.019716
R43303 DVDD.n980 DVDD.n956 0.019716
R43304 DVDD.n1220 DVDD.n1219 0.019716
R43305 DVDD.n1219 DVDD.n955 0.019716
R43306 DVDD.n986 DVDD.n985 0.019716
R43307 DVDD.n985 DVDD.n954 0.019716
R43308 DVDD.n1211 DVDD.n1210 0.019716
R43309 DVDD.n1210 DVDD.n953 0.019716
R43310 DVDD.n991 DVDD.n990 0.019716
R43311 DVDD.n990 DVDD.n952 0.019716
R43312 DVDD.n1202 DVDD.n1201 0.019716
R43313 DVDD.n1201 DVDD.n951 0.019716
R43314 DVDD.n996 DVDD.n995 0.019716
R43315 DVDD.n995 DVDD.n950 0.019716
R43316 DVDD.n1193 DVDD.n1192 0.019716
R43317 DVDD.n1192 DVDD.n949 0.019716
R43318 DVDD.n1001 DVDD.n1000 0.019716
R43319 DVDD.n1000 DVDD.n948 0.019716
R43320 DVDD.n1184 DVDD.n1183 0.019716
R43321 DVDD.n1183 DVDD.n947 0.019716
R43322 DVDD.n1006 DVDD.n1005 0.019716
R43323 DVDD.n1005 DVDD.n946 0.019716
R43324 DVDD.n1175 DVDD.n1174 0.019716
R43325 DVDD.n1174 DVDD.n945 0.019716
R43326 DVDD.n1011 DVDD.n1010 0.019716
R43327 DVDD.n1010 DVDD.n944 0.019716
R43328 DVDD.n1166 DVDD.n1165 0.019716
R43329 DVDD.n1165 DVDD.n943 0.019716
R43330 DVDD.n1016 DVDD.n1015 0.019716
R43331 DVDD.n1015 DVDD.n942 0.019716
R43332 DVDD.n1157 DVDD.n1156 0.019716
R43333 DVDD.n1156 DVDD.n941 0.019716
R43334 DVDD.n1021 DVDD.n1020 0.019716
R43335 DVDD.n1020 DVDD.n940 0.019716
R43336 DVDD.n1148 DVDD.n1147 0.019716
R43337 DVDD.n1147 DVDD.n939 0.019716
R43338 DVDD.n1026 DVDD.n1025 0.019716
R43339 DVDD.n1025 DVDD.n938 0.019716
R43340 DVDD.n1139 DVDD.n1138 0.019716
R43341 DVDD.n1138 DVDD.n937 0.019716
R43342 DVDD.n1031 DVDD.n1030 0.019716
R43343 DVDD.n1030 DVDD.n936 0.019716
R43344 DVDD.n1130 DVDD.n1129 0.019716
R43345 DVDD.n1129 DVDD.n935 0.019716
R43346 DVDD.n1036 DVDD.n1035 0.019716
R43347 DVDD.n1035 DVDD.n934 0.019716
R43348 DVDD.n1121 DVDD.n1120 0.019716
R43349 DVDD.n1120 DVDD.n933 0.019716
R43350 DVDD.n1041 DVDD.n1040 0.019716
R43351 DVDD.n1040 DVDD.n932 0.019716
R43352 DVDD.n1112 DVDD.n1111 0.019716
R43353 DVDD.n1111 DVDD.n931 0.019716
R43354 DVDD.n1046 DVDD.n1045 0.019716
R43355 DVDD.n1045 DVDD.n930 0.019716
R43356 DVDD.n1103 DVDD.n1102 0.019716
R43357 DVDD.n1102 DVDD.n929 0.019716
R43358 DVDD.n1051 DVDD.n1050 0.019716
R43359 DVDD.n1050 DVDD.n928 0.019716
R43360 DVDD.n1094 DVDD.n1093 0.019716
R43361 DVDD.n1093 DVDD.n927 0.019716
R43362 DVDD.n1056 DVDD.n1055 0.019716
R43363 DVDD.n1055 DVDD.n926 0.019716
R43364 DVDD.n1085 DVDD.n1084 0.019716
R43365 DVDD.n1084 DVDD.n925 0.019716
R43366 DVDD.n1061 DVDD.n1060 0.019716
R43367 DVDD.n1060 DVDD.n924 0.019716
R43368 DVDD.n1076 DVDD.n1075 0.019716
R43369 DVDD.n1075 DVDD.n923 0.019716
R43370 DVDD.n1066 DVDD.n1065 0.019716
R43371 DVDD.n1065 DVDD.n922 0.019716
R43372 DVDD.n1254 DVDD.n964 0.019716
R43373 DVDD.n1255 DVDD.n1254 0.019716
R43374 DVDD.n1248 DVDD.n1247 0.019716
R43375 DVDD.n1248 DVDD.n962 0.019716
R43376 DVDD.n972 DVDD.n971 0.019716
R43377 DVDD.n972 DVDD.n961 0.019716
R43378 DVDD.n1239 DVDD.n1238 0.019716
R43379 DVDD.n1239 DVDD.n960 0.019716
R43380 DVDD.n977 DVDD.n976 0.019716
R43381 DVDD.n977 DVDD.n959 0.019716
R43382 DVDD.n1230 DVDD.n1229 0.019716
R43383 DVDD.n1230 DVDD.n958 0.019716
R43384 DVDD.n982 DVDD.n981 0.019716
R43385 DVDD.n982 DVDD.n957 0.019716
R43386 DVDD.n1221 DVDD.n1220 0.019716
R43387 DVDD.n1221 DVDD.n956 0.019716
R43388 DVDD.n987 DVDD.n986 0.019716
R43389 DVDD.n987 DVDD.n955 0.019716
R43390 DVDD.n1212 DVDD.n1211 0.019716
R43391 DVDD.n1212 DVDD.n954 0.019716
R43392 DVDD.n992 DVDD.n991 0.019716
R43393 DVDD.n992 DVDD.n953 0.019716
R43394 DVDD.n1203 DVDD.n1202 0.019716
R43395 DVDD.n1203 DVDD.n952 0.019716
R43396 DVDD.n997 DVDD.n996 0.019716
R43397 DVDD.n997 DVDD.n951 0.019716
R43398 DVDD.n1194 DVDD.n1193 0.019716
R43399 DVDD.n1194 DVDD.n950 0.019716
R43400 DVDD.n1002 DVDD.n1001 0.019716
R43401 DVDD.n1002 DVDD.n949 0.019716
R43402 DVDD.n1185 DVDD.n1184 0.019716
R43403 DVDD.n1185 DVDD.n948 0.019716
R43404 DVDD.n1007 DVDD.n1006 0.019716
R43405 DVDD.n1007 DVDD.n947 0.019716
R43406 DVDD.n1176 DVDD.n1175 0.019716
R43407 DVDD.n1176 DVDD.n946 0.019716
R43408 DVDD.n1012 DVDD.n1011 0.019716
R43409 DVDD.n1012 DVDD.n945 0.019716
R43410 DVDD.n1167 DVDD.n1166 0.019716
R43411 DVDD.n1167 DVDD.n944 0.019716
R43412 DVDD.n1017 DVDD.n1016 0.019716
R43413 DVDD.n1017 DVDD.n943 0.019716
R43414 DVDD.n1158 DVDD.n1157 0.019716
R43415 DVDD.n1158 DVDD.n942 0.019716
R43416 DVDD.n1022 DVDD.n1021 0.019716
R43417 DVDD.n1022 DVDD.n941 0.019716
R43418 DVDD.n1149 DVDD.n1148 0.019716
R43419 DVDD.n1149 DVDD.n940 0.019716
R43420 DVDD.n1027 DVDD.n1026 0.019716
R43421 DVDD.n1027 DVDD.n939 0.019716
R43422 DVDD.n1140 DVDD.n1139 0.019716
R43423 DVDD.n1140 DVDD.n938 0.019716
R43424 DVDD.n1032 DVDD.n1031 0.019716
R43425 DVDD.n1032 DVDD.n937 0.019716
R43426 DVDD.n1131 DVDD.n1130 0.019716
R43427 DVDD.n1131 DVDD.n936 0.019716
R43428 DVDD.n1037 DVDD.n1036 0.019716
R43429 DVDD.n1037 DVDD.n935 0.019716
R43430 DVDD.n1122 DVDD.n1121 0.019716
R43431 DVDD.n1122 DVDD.n934 0.019716
R43432 DVDD.n1042 DVDD.n1041 0.019716
R43433 DVDD.n1042 DVDD.n933 0.019716
R43434 DVDD.n1113 DVDD.n1112 0.019716
R43435 DVDD.n1113 DVDD.n932 0.019716
R43436 DVDD.n1047 DVDD.n1046 0.019716
R43437 DVDD.n1047 DVDD.n931 0.019716
R43438 DVDD.n1104 DVDD.n1103 0.019716
R43439 DVDD.n1104 DVDD.n930 0.019716
R43440 DVDD.n1052 DVDD.n1051 0.019716
R43441 DVDD.n1052 DVDD.n929 0.019716
R43442 DVDD.n1095 DVDD.n1094 0.019716
R43443 DVDD.n1095 DVDD.n928 0.019716
R43444 DVDD.n1057 DVDD.n1056 0.019716
R43445 DVDD.n1057 DVDD.n927 0.019716
R43446 DVDD.n1086 DVDD.n1085 0.019716
R43447 DVDD.n1086 DVDD.n926 0.019716
R43448 DVDD.n1062 DVDD.n1061 0.019716
R43449 DVDD.n1062 DVDD.n925 0.019716
R43450 DVDD.n1077 DVDD.n1076 0.019716
R43451 DVDD.n1077 DVDD.n924 0.019716
R43452 DVDD.n1067 DVDD.n1066 0.019716
R43453 DVDD.n1067 DVDD.n923 0.019716
R43454 DVDD.n1068 DVDD.n922 0.019716
R43455 DVDD.n6330 DVDD.n6042 0.019716
R43456 DVDD.n6092 DVDD.n6041 0.019716
R43457 DVDD.n6092 DVDD.n6090 0.019716
R43458 DVDD.n6321 DVDD.n6040 0.019716
R43459 DVDD.n6321 DVDD.n6089 0.019716
R43460 DVDD.n6096 DVDD.n6039 0.019716
R43461 DVDD.n6096 DVDD.n6088 0.019716
R43462 DVDD.n6312 DVDD.n6038 0.019716
R43463 DVDD.n6312 DVDD.n6087 0.019716
R43464 DVDD.n6099 DVDD.n6037 0.019716
R43465 DVDD.n6099 DVDD.n6086 0.019716
R43466 DVDD.n6303 DVDD.n6036 0.019716
R43467 DVDD.n6303 DVDD.n6085 0.019716
R43468 DVDD.n6102 DVDD.n6035 0.019716
R43469 DVDD.n6102 DVDD.n6084 0.019716
R43470 DVDD.n6294 DVDD.n6034 0.019716
R43471 DVDD.n6294 DVDD.n6083 0.019716
R43472 DVDD.n6105 DVDD.n6033 0.019716
R43473 DVDD.n6105 DVDD.n6082 0.019716
R43474 DVDD.n6285 DVDD.n6032 0.019716
R43475 DVDD.n6285 DVDD.n6081 0.019716
R43476 DVDD.n6108 DVDD.n6031 0.019716
R43477 DVDD.n6108 DVDD.n6080 0.019716
R43478 DVDD.n6276 DVDD.n6030 0.019716
R43479 DVDD.n6276 DVDD.n6079 0.019716
R43480 DVDD.n6111 DVDD.n6029 0.019716
R43481 DVDD.n6111 DVDD.n6078 0.019716
R43482 DVDD.n6267 DVDD.n6028 0.019716
R43483 DVDD.n6267 DVDD.n6077 0.019716
R43484 DVDD.n6114 DVDD.n6027 0.019716
R43485 DVDD.n6114 DVDD.n6076 0.019716
R43486 DVDD.n6258 DVDD.n6026 0.019716
R43487 DVDD.n6258 DVDD.n6075 0.019716
R43488 DVDD.n6117 DVDD.n6025 0.019716
R43489 DVDD.n6117 DVDD.n6074 0.019716
R43490 DVDD.n6249 DVDD.n6024 0.019716
R43491 DVDD.n6249 DVDD.n6073 0.019716
R43492 DVDD.n6120 DVDD.n6023 0.019716
R43493 DVDD.n6120 DVDD.n6072 0.019716
R43494 DVDD.n6240 DVDD.n6022 0.019716
R43495 DVDD.n6240 DVDD.n6071 0.019716
R43496 DVDD.n6123 DVDD.n6021 0.019716
R43497 DVDD.n6123 DVDD.n6070 0.019716
R43498 DVDD.n6231 DVDD.n6020 0.019716
R43499 DVDD.n6231 DVDD.n6069 0.019716
R43500 DVDD.n6126 DVDD.n6019 0.019716
R43501 DVDD.n6126 DVDD.n6068 0.019716
R43502 DVDD.n6222 DVDD.n6018 0.019716
R43503 DVDD.n6222 DVDD.n6067 0.019716
R43504 DVDD.n6129 DVDD.n6017 0.019716
R43505 DVDD.n6129 DVDD.n6066 0.019716
R43506 DVDD.n6213 DVDD.n6016 0.019716
R43507 DVDD.n6213 DVDD.n6065 0.019716
R43508 DVDD.n6132 DVDD.n6015 0.019716
R43509 DVDD.n6132 DVDD.n6064 0.019716
R43510 DVDD.n6204 DVDD.n6014 0.019716
R43511 DVDD.n6204 DVDD.n6063 0.019716
R43512 DVDD.n6135 DVDD.n6013 0.019716
R43513 DVDD.n6135 DVDD.n6062 0.019716
R43514 DVDD.n6195 DVDD.n6012 0.019716
R43515 DVDD.n6195 DVDD.n6061 0.019716
R43516 DVDD.n6138 DVDD.n6011 0.019716
R43517 DVDD.n6138 DVDD.n6060 0.019716
R43518 DVDD.n6186 DVDD.n6010 0.019716
R43519 DVDD.n6186 DVDD.n6059 0.019716
R43520 DVDD.n6141 DVDD.n6009 0.019716
R43521 DVDD.n6141 DVDD.n6058 0.019716
R43522 DVDD.n6177 DVDD.n6008 0.019716
R43523 DVDD.n6177 DVDD.n6057 0.019716
R43524 DVDD.n6144 DVDD.n6007 0.019716
R43525 DVDD.n6144 DVDD.n6056 0.019716
R43526 DVDD.n6168 DVDD.n6006 0.019716
R43527 DVDD.n6168 DVDD.n6055 0.019716
R43528 DVDD.n6147 DVDD.n6005 0.019716
R43529 DVDD.n6147 DVDD.n6054 0.019716
R43530 DVDD.n6159 DVDD.n6004 0.019716
R43531 DVDD.n6159 DVDD.n6053 0.019716
R43532 DVDD.n6150 DVDD.n6003 0.019716
R43533 DVDD.n6150 DVDD.n6052 0.019716
R43534 DVDD.n6050 DVDD.n6002 0.019716
R43535 DVDD.n6332 DVDD.n6050 0.019716
R43536 DVDD.n6046 DVDD.n6001 0.019716
R43537 DVDD.n6046 DVDD.n6045 0.019716
R43538 DVDD.n6329 DVDD.n6041 0.019716
R43539 DVDD.n6330 DVDD.n6329 0.019716
R43540 DVDD.n6323 DVDD.n6040 0.019716
R43541 DVDD.n6323 DVDD.n6090 0.019716
R43542 DVDD.n6319 DVDD.n6039 0.019716
R43543 DVDD.n6319 DVDD.n6089 0.019716
R43544 DVDD.n6314 DVDD.n6038 0.019716
R43545 DVDD.n6314 DVDD.n6088 0.019716
R43546 DVDD.n6310 DVDD.n6037 0.019716
R43547 DVDD.n6310 DVDD.n6087 0.019716
R43548 DVDD.n6305 DVDD.n6036 0.019716
R43549 DVDD.n6305 DVDD.n6086 0.019716
R43550 DVDD.n6301 DVDD.n6035 0.019716
R43551 DVDD.n6301 DVDD.n6085 0.019716
R43552 DVDD.n6296 DVDD.n6034 0.019716
R43553 DVDD.n6296 DVDD.n6084 0.019716
R43554 DVDD.n6292 DVDD.n6033 0.019716
R43555 DVDD.n6292 DVDD.n6083 0.019716
R43556 DVDD.n6287 DVDD.n6032 0.019716
R43557 DVDD.n6287 DVDD.n6082 0.019716
R43558 DVDD.n6283 DVDD.n6031 0.019716
R43559 DVDD.n6283 DVDD.n6081 0.019716
R43560 DVDD.n6278 DVDD.n6030 0.019716
R43561 DVDD.n6278 DVDD.n6080 0.019716
R43562 DVDD.n6274 DVDD.n6029 0.019716
R43563 DVDD.n6274 DVDD.n6079 0.019716
R43564 DVDD.n6269 DVDD.n6028 0.019716
R43565 DVDD.n6269 DVDD.n6078 0.019716
R43566 DVDD.n6265 DVDD.n6027 0.019716
R43567 DVDD.n6265 DVDD.n6077 0.019716
R43568 DVDD.n6260 DVDD.n6026 0.019716
R43569 DVDD.n6260 DVDD.n6076 0.019716
R43570 DVDD.n6256 DVDD.n6025 0.019716
R43571 DVDD.n6256 DVDD.n6075 0.019716
R43572 DVDD.n6251 DVDD.n6024 0.019716
R43573 DVDD.n6251 DVDD.n6074 0.019716
R43574 DVDD.n6247 DVDD.n6023 0.019716
R43575 DVDD.n6247 DVDD.n6073 0.019716
R43576 DVDD.n6242 DVDD.n6022 0.019716
R43577 DVDD.n6242 DVDD.n6072 0.019716
R43578 DVDD.n6238 DVDD.n6021 0.019716
R43579 DVDD.n6238 DVDD.n6071 0.019716
R43580 DVDD.n6233 DVDD.n6020 0.019716
R43581 DVDD.n6233 DVDD.n6070 0.019716
R43582 DVDD.n6229 DVDD.n6019 0.019716
R43583 DVDD.n6229 DVDD.n6069 0.019716
R43584 DVDD.n6224 DVDD.n6018 0.019716
R43585 DVDD.n6224 DVDD.n6068 0.019716
R43586 DVDD.n6220 DVDD.n6017 0.019716
R43587 DVDD.n6220 DVDD.n6067 0.019716
R43588 DVDD.n6215 DVDD.n6016 0.019716
R43589 DVDD.n6215 DVDD.n6066 0.019716
R43590 DVDD.n6211 DVDD.n6015 0.019716
R43591 DVDD.n6211 DVDD.n6065 0.019716
R43592 DVDD.n6206 DVDD.n6014 0.019716
R43593 DVDD.n6206 DVDD.n6064 0.019716
R43594 DVDD.n6202 DVDD.n6013 0.019716
R43595 DVDD.n6202 DVDD.n6063 0.019716
R43596 DVDD.n6197 DVDD.n6012 0.019716
R43597 DVDD.n6197 DVDD.n6062 0.019716
R43598 DVDD.n6193 DVDD.n6011 0.019716
R43599 DVDD.n6193 DVDD.n6061 0.019716
R43600 DVDD.n6188 DVDD.n6010 0.019716
R43601 DVDD.n6188 DVDD.n6060 0.019716
R43602 DVDD.n6184 DVDD.n6009 0.019716
R43603 DVDD.n6184 DVDD.n6059 0.019716
R43604 DVDD.n6179 DVDD.n6008 0.019716
R43605 DVDD.n6179 DVDD.n6058 0.019716
R43606 DVDD.n6175 DVDD.n6007 0.019716
R43607 DVDD.n6175 DVDD.n6057 0.019716
R43608 DVDD.n6170 DVDD.n6006 0.019716
R43609 DVDD.n6170 DVDD.n6056 0.019716
R43610 DVDD.n6166 DVDD.n6005 0.019716
R43611 DVDD.n6166 DVDD.n6055 0.019716
R43612 DVDD.n6161 DVDD.n6004 0.019716
R43613 DVDD.n6161 DVDD.n6054 0.019716
R43614 DVDD.n6157 DVDD.n6003 0.019716
R43615 DVDD.n6157 DVDD.n6053 0.019716
R43616 DVDD.n6152 DVDD.n6002 0.019716
R43617 DVDD.n6152 DVDD.n6052 0.019716
R43618 DVDD.n6333 DVDD.n6001 0.019716
R43619 DVDD.n6333 DVDD.n6332 0.019716
R43620 DVDD.n15111 DVDD.n6045 0.019716
R43621 DVDD.n18414 DVDD.n18401 0.019625
R43622 DVDD.n22015 DVDD.n21985 0.019625
R43623 DVDD.n21353 DVDD.n21352 0.019625
R43624 DVDD.n21703 DVDD.n21702 0.019625
R43625 DVDD.n18251 DVDD.n18229 0.019625
R43626 DVDD.n18436 DVDD.n161 0.019625
R43627 DVDD.n4290 DVDD.n4283 0.019625
R43628 DVDD.n3692 DVDD.n3691 0.019625
R43629 DVDD.n14007 DVDD.n11058 0.019625
R43630 DVDD.n17284 DVDD.n1259 0.019625
R43631 DVDD.n12726 DVDD.n12478 0.0195611
R43632 DVDD.n13265 DVDD.n12913 0.0195611
R43633 DVDD.n13481 DVDD.n12727 0.0195611
R43634 DVDD.n13264 DVDD.n12914 0.0195611
R43635 DVDD.n13792 DVDD.n13791 0.019175
R43636 DVDD.n17000 DVDD.n1608 0.019175
R43637 DVDD.n10584 DVDD.n8608 0.0191681
R43638 DVDD.n10581 DVDD.n8607 0.0191681
R43639 DVDD.n6341 DVDD.n6044 0.0187751
R43640 DVDD.n15109 DVDD.n15108 0.0187751
R43641 DVDD.n14855 DVDD.n7673 0.018725
R43642 DVDD.n9668 DVDD.n9608 0.0177098
R43643 DVDD.n9741 DVDD.n9740 0.0177098
R43644 DVDD.n10095 DVDD.n10094 0.0177098
R43645 DVDD.n10097 DVDD.n9610 0.0177098
R43646 DVDD.n15062 DVDD.n7409 0.0175961
R43647 DVDD.n15063 DVDD.n7408 0.0175961
R43648 DVDD.n21684 DVDD.n18533 0.0175526
R43649 DVDD.n18364 DVDD.n18315 0.0175526
R43650 DVDD.n3916 DVDD.n229 0.0175526
R43651 DVDD.n21769 DVDD.n18392 0.0175526
R43652 DVDD.n21931 DVDD.n21930 0.0175526
R43653 DVDD.n22121 DVDD.n22069 0.0175526
R43654 DVDD.n21944 DVDD.n18380 0.017375
R43655 DVDD.n22209 DVDD.n182 0.017375
R43656 DVDD.n22039 DVDD.n18246 0.017375
R43657 DVDD.n18277 DVDD.n223 0.017375
R43658 DVDD.n22229 DVDD.n141 0.017375
R43659 DVDD.n21239 DVDD.n18432 0.017375
R43660 DVDD.n21944 DVDD.n18304 0.017375
R43661 DVDD.n22209 DVDD.n192 0.017375
R43662 DVDD.n22039 DVDD.n18250 0.017375
R43663 DVDD.n21820 DVDD.n223 0.017375
R43664 DVDD.n22229 DVDD.n153 0.017375
R43665 DVDD.n18468 DVDD.n18432 0.017375
R43666 DVDD.n4574 DVDD.n4314 0.017375
R43667 DVDD.n4313 DVDD.n4282 0.017375
R43668 DVDD.n3709 DVDD.n3708 0.017375
R43669 DVDD.n4759 DVDD.n3675 0.017375
R43670 DVDD.n15139 DVDD.n15138 0.017282
R43671 DVDD.n15118 DVDD.n5582 0.017282
R43672 DVDD.n15118 DVDD.n15117 0.017282
R43673 DVDD.n15117 DVDD.n15116 0.017282
R43674 DVDD.n6399 DVDD.n6397 0.017282
R43675 DVDD.n6701 DVDD.n6397 0.017282
R43676 DVDD.n15097 DVDD.n15096 0.017282
R43677 DVDD.n15096 DVDD.n15095 0.017282
R43678 DVDD.n7065 DVDD.n7064 0.017282
R43679 DVDD.n15075 DVDD.n7065 0.017282
R43680 DVDD.n15073 DVDD.n7067 0.017282
R43681 DVDD.n7563 DVDD.n7067 0.017282
R43682 DVDD.n14869 DVDD.n7563 0.017282
R43683 DVDD.n14869 DVDD.n7564 0.017282
R43684 DVDD.n8974 DVDD.n7564 0.017282
R43685 DVDD.n9566 DVDD.n9565 0.017282
R43686 DVDD.n9565 DVDD.n9564 0.017282
R43687 DVDD.n14846 DVDD.n14845 0.017282
R43688 DVDD.n14845 DVDD.n14844 0.017282
R43689 DVDD.n8140 DVDD.n8138 0.017282
R43690 DVDD.n8140 DVDD.n8139 0.017282
R43691 DVDD.n14574 DVDD.n14573 0.017282
R43692 DVDD.n14573 DVDD.n14572 0.017282
R43693 DVDD.n14572 DVDD.n8150 0.017282
R43694 DVDD.n14308 DVDD.n14307 0.017282
R43695 DVDD.n14307 DVDD.n14306 0.017282
R43696 DVDD.n10227 DVDD.n10226 0.017282
R43697 DVDD.n14290 DVDD.n14289 0.017282
R43698 DVDD.n14289 DVDD.n14288 0.017282
R43699 DVDD.n10698 DVDD.n10697 0.017282
R43700 DVDD.n10700 DVDD.n10698 0.017282
R43701 DVDD.n10700 DVDD.n10699 0.017282
R43702 DVDD.n14018 DVDD.n14017 0.017282
R43703 DVDD.n14017 DVDD.n14016 0.017282
R43704 DVDD.n11218 DVDD.n11217 0.017282
R43705 DVDD.n11217 DVDD.n11212 0.017282
R43706 DVDD.n13811 DVDD.n11213 0.017282
R43707 DVDD.n13805 DVDD.n11213 0.017282
R43708 DVDD.n13803 DVDD.n11230 0.017282
R43709 DVDD.n13783 DVDD.n11230 0.017282
R43710 DVDD.n13781 DVDD.n11585 0.017282
R43711 DVDD.n13761 DVDD.n13760 0.017282
R43712 DVDD.n13758 DVDD.n11931 0.017282
R43713 DVDD.n12378 DVDD.n11931 0.017282
R43714 DVDD.n13493 DVDD.n13492 0.017282
R43715 DVDD.n13492 DVDD.n13491 0.017282
R43716 DVDD.n12892 DVDD.n12891 0.017282
R43717 DVDD.n12891 DVDD.n12888 0.017282
R43718 DVDD.n13281 DVDD.n12889 0.017282
R43719 DVDD.n13275 DVDD.n12889 0.017282
R43720 DVDD.n13275 DVDD.n13274 0.017282
R43721 DVDD.n13272 DVDD.n12905 0.017282
R43722 DVDD.n12905 DVDD.n12904 0.017282
R43723 DVDD.n16719 DVDD.n1818 0.017282
R43724 DVDD.n16723 DVDD.n16722 0.017282
R43725 DVDD.n16722 DVDD.n16721 0.017282
R43726 DVDD.n16742 DVDD.n16741 0.017282
R43727 DVDD.n16741 DVDD.n16740 0.017282
R43728 DVDD.n17010 DVDD.n17009 0.017282
R43729 DVDD.n17009 DVDD.n1268 0.017282
R43730 DVDD.n17275 DVDD.n1268 0.017282
R43731 DVDD.n17277 DVDD.n919 0.017282
R43732 DVDD.n17293 DVDD.n919 0.017282
R43733 DVDD.n17295 DVDD.n901 0.017282
R43734 DVDD.n17721 DVDD.n901 0.017282
R43735 DVDD.n17724 DVDD.n17721 0.017282
R43736 DVDD.n17724 DVDD.n17723 0.017282
R43737 DVDD.n17723 DVDD.n890 0.017282
R43738 DVDD.n4845 DVDD.n4839 0.0172684
R43739 DVDD.n18125 DVDD.n474 0.0172684
R43740 DVDD.n14005 DVDD.n11060 0.0172031
R43741 DVDD.n17282 DVDD.n1261 0.0172031
R43742 DVDD.n14006 DVDD.n11059 0.0172031
R43743 DVDD.n17283 DVDD.n1260 0.0172031
R43744 DVDD.n21969 DVDD.n18275 0.0170221
R43745 DVDD.n21697 DVDD.n21696 0.0170221
R43746 DVDD.n21822 DVDD.n21818 0.0170221
R43747 DVDD.n18420 DVDD.n18412 0.0170221
R43748 DVDD.n4802 DVDD.n3565 0.0169834
R43749 DVDD.n8605 DVDD.n8604 0.016925
R43750 DVDD.n13789 DVDD.n11277 0.01681
R43751 DVDD.n17002 DVDD.n1610 0.01681
R43752 DVDD.n13790 DVDD.n11577 0.01681
R43753 DVDD.n17001 DVDD.n1609 0.01681
R43754 DVDD.n14018 DVDD.n10686 0.0167406
R43755 DVDD.n16740 DVDD.n1702 0.0167406
R43756 DVDD.n22020 DVDD.n22019 0.0166964
R43757 DVDD.n21348 DVDD.n21347 0.0166964
R43758 DVDD.n21244 DVDD.n21218 0.0166964
R43759 DVDD.n21957 DVDD.n21956 0.0166964
R43760 DVDD.n18258 DVDD.n18257 0.0166964
R43761 DVDD.n21854 DVDD.n21853 0.0166964
R43762 DVDD.n18442 DVDD.n18441 0.0166964
R43763 DVDD.n18470 DVDD.n18466 0.0166964
R43764 DVDD.n4286 DVDD.n4285 0.0166964
R43765 DVDD.n4308 DVDD.n4301 0.0166964
R43766 DVDD.n3686 DVDD.n3685 0.0166964
R43767 DVDD.n3702 DVDD.n3701 0.0166964
R43768 DVDD.n13477 DVDD.n12732 0.016475
R43769 DVDD.n12918 DVDD.n12732 0.016475
R43770 DVDD.n15138 DVDD.n15136 0.0164699
R43771 DVDD.n7664 DVDD.n7658 0.016417
R43772 DVDD.n14857 DVDD.n14856 0.016417
R43773 DVDD.n18409 DVDD.n18403 0.0163049
R43774 DVDD.n21858 DVDD.n21809 0.0163049
R43775 DVDD.n22157 DVDD.n315 0.0163049
R43776 DVDD.n21737 DVDD.n18424 0.0163049
R43777 DVDD.n21901 DVDD.n21811 0.0163049
R43778 DVDD.n22139 DVDD.n366 0.0163049
R43779 DVDD.n21647 DVDD.n18529 0.0163049
R43780 DVDD.n21965 DVDD.n21964 0.0163049
R43781 DVDD.n22183 DVDD.n22182 0.0163049
R43782 DVDD.n21686 DVDD.n18530 0.0163049
R43783 DVDD.n21967 DVDD.n18280 0.0163049
R43784 DVDD.n22185 DVDD.n231 0.0163049
R43785 DVDD.n15142 DVDD.n5577 0.0161992
R43786 DVDD.n13783 DVDD.n13782 0.0161992
R43787 DVDD.n13273 DVDD.n13272 0.0161992
R43788 DVDD.n20496 DVDD.n20495 0.0161121
R43789 DVDD.n20518 DVDD.n20517 0.0161121
R43790 DVDD.n20503 DVDD.n20497 0.0161121
R43791 DVDD.n20503 DVDD.n20494 0.0161121
R43792 DVDD.n20504 DVDD.n20502 0.0161121
R43793 DVDD.n20502 DVDD.n20493 0.0161121
R43794 DVDD.n20506 DVDD.n20501 0.0161121
R43795 DVDD.n20501 DVDD.n20492 0.0161121
R43796 DVDD.n20508 DVDD.n20500 0.0161121
R43797 DVDD.n20500 DVDD.n20491 0.0161121
R43798 DVDD.n20510 DVDD.n20499 0.0161121
R43799 DVDD.n20499 DVDD.n20490 0.0161121
R43800 DVDD.n20512 DVDD.n20498 0.0161121
R43801 DVDD.n20498 DVDD.n20489 0.0161121
R43802 DVDD.n20514 DVDD.n20488 0.0161121
R43803 DVDD.n19787 DVDD.n19773 0.0161121
R43804 DVDD.n19796 DVDD.n19772 0.0161121
R43805 DVDD.n19786 DVDD.n19772 0.0161121
R43806 DVDD.n19795 DVDD.n19771 0.0161121
R43807 DVDD.n19785 DVDD.n19771 0.0161121
R43808 DVDD.n19794 DVDD.n19770 0.0161121
R43809 DVDD.n19784 DVDD.n19770 0.0161121
R43810 DVDD.n19793 DVDD.n19769 0.0161121
R43811 DVDD.n19783 DVDD.n19769 0.0161121
R43812 DVDD.n19792 DVDD.n19768 0.0161121
R43813 DVDD.n19782 DVDD.n19768 0.0161121
R43814 DVDD.n20536 DVDD.n19791 0.0161121
R43815 DVDD.n20537 DVDD.n19780 0.0161121
R43816 DVDD.n20449 DVDD.n19817 0.0161121
R43817 DVDD.n20448 DVDD.n19816 0.0161121
R43818 DVDD.n20451 DVDD.n20448 0.0161121
R43819 DVDD.n20447 DVDD.n19815 0.0161121
R43820 DVDD.n20453 DVDD.n20447 0.0161121
R43821 DVDD.n20446 DVDD.n19814 0.0161121
R43822 DVDD.n20455 DVDD.n20446 0.0161121
R43823 DVDD.n20445 DVDD.n19813 0.0161121
R43824 DVDD.n20457 DVDD.n20445 0.0161121
R43825 DVDD.n20444 DVDD.n19812 0.0161121
R43826 DVDD.n20459 DVDD.n20444 0.0161121
R43827 DVDD.n20442 DVDD.n19811 0.0161121
R43828 DVDD.n20461 DVDD.n19818 0.0161121
R43829 DVDD.n20908 DVDD.n20907 0.0161121
R43830 DVDD.n20908 DVDD.n18910 0.0161121
R43831 DVDD.n20910 DVDD.n20909 0.0161121
R43832 DVDD.n20910 DVDD.n18911 0.0161121
R43833 DVDD.n20912 DVDD.n20911 0.0161121
R43834 DVDD.n20912 DVDD.n18912 0.0161121
R43835 DVDD.n20914 DVDD.n20913 0.0161121
R43836 DVDD.n20914 DVDD.n18913 0.0161121
R43837 DVDD.n20916 DVDD.n20915 0.0161121
R43838 DVDD.n20916 DVDD.n18914 0.0161121
R43839 DVDD.n20918 DVDD.n20917 0.0161121
R43840 DVDD.n20918 DVDD.n18915 0.0161121
R43841 DVDD.n20920 DVDD.n18918 0.0161121
R43842 DVDD.n20921 DVDD.n20920 0.0161121
R43843 DVDD.n18916 DVDD.n18820 0.0161121
R43844 DVDD.n21011 DVDD.n18823 0.0161121
R43845 DVDD.n21010 DVDD.n20991 0.0161121
R43846 DVDD.n20990 DVDD.n20989 0.0161121
R43847 DVDD.n20993 DVDD.n20989 0.0161121
R43848 DVDD.n20992 DVDD.n20988 0.0161121
R43849 DVDD.n20996 DVDD.n20988 0.0161121
R43850 DVDD.n20995 DVDD.n20987 0.0161121
R43851 DVDD.n20999 DVDD.n20987 0.0161121
R43852 DVDD.n20998 DVDD.n20986 0.0161121
R43853 DVDD.n21002 DVDD.n20986 0.0161121
R43854 DVDD.n21001 DVDD.n20985 0.0161121
R43855 DVDD.n21005 DVDD.n20985 0.0161121
R43856 DVDD.n21004 DVDD.n20984 0.0161121
R43857 DVDD.n21008 DVDD.n20984 0.0161121
R43858 DVDD.n21007 DVDD.n20983 0.0161121
R43859 DVDD.n21067 DVDD.n18751 0.0161121
R43860 DVDD.n21066 DVDD.n18750 0.0161121
R43861 DVDD.n21069 DVDD.n21066 0.0161121
R43862 DVDD.n21065 DVDD.n18749 0.0161121
R43863 DVDD.n21071 DVDD.n21065 0.0161121
R43864 DVDD.n21064 DVDD.n18748 0.0161121
R43865 DVDD.n21073 DVDD.n21064 0.0161121
R43866 DVDD.n21063 DVDD.n18747 0.0161121
R43867 DVDD.n21075 DVDD.n21063 0.0161121
R43868 DVDD.n21062 DVDD.n18746 0.0161121
R43869 DVDD.n21077 DVDD.n21062 0.0161121
R43870 DVDD.n21061 DVDD.n18745 0.0161121
R43871 DVDD.n21079 DVDD.n21061 0.0161121
R43872 DVDD.n18752 DVDD.n18744 0.0161121
R43873 DVDD.n18800 DVDD.n18799 0.0161121
R43874 DVDD.n18798 DVDD.n18797 0.0161121
R43875 DVDD.n18797 DVDD.n18795 0.0161121
R43876 DVDD.n18793 DVDD.n18792 0.0161121
R43877 DVDD.n18802 DVDD.n18792 0.0161121
R43878 DVDD.n18803 DVDD.n18791 0.0161121
R43879 DVDD.n18805 DVDD.n18791 0.0161121
R43880 DVDD.n18806 DVDD.n18790 0.0161121
R43881 DVDD.n18808 DVDD.n18790 0.0161121
R43882 DVDD.n18809 DVDD.n18789 0.0161121
R43883 DVDD.n18811 DVDD.n18789 0.0161121
R43884 DVDD.n18812 DVDD.n18788 0.0161121
R43885 DVDD.n18814 DVDD.n18788 0.0161121
R43886 DVDD.n18815 DVDD.n18787 0.0161121
R43887 DVDD.n18817 DVDD.n18787 0.0161121
R43888 DVDD.n21027 DVDD.n18818 0.0161121
R43889 DVDD.n21027 DVDD.n21026 0.0161121
R43890 DVDD.n21030 DVDD.n21028 0.0161121
R43891 DVDD.n21030 DVDD.n21029 0.0161121
R43892 DVDD.n21033 DVDD.n21031 0.0161121
R43893 DVDD.n21033 DVDD.n21032 0.0161121
R43894 DVDD.n21036 DVDD.n21034 0.0161121
R43895 DVDD.n21036 DVDD.n21035 0.0161121
R43896 DVDD.n21039 DVDD.n21037 0.0161121
R43897 DVDD.n21039 DVDD.n21038 0.0161121
R43898 DVDD.n21042 DVDD.n21040 0.0161121
R43899 DVDD.n21042 DVDD.n21041 0.0161121
R43900 DVDD.n21044 DVDD.n21043 0.0161121
R43901 DVDD.n21046 DVDD.n21044 0.0161121
R43902 DVDD.n21045 DVDD.n21019 0.0161121
R43903 DVDD.n18801 DVDD.n18800 0.0161121
R43904 DVDD.n18794 DVDD.n18793 0.0161121
R43905 DVDD.n18804 DVDD.n18803 0.0161121
R43906 DVDD.n18807 DVDD.n18806 0.0161121
R43907 DVDD.n18810 DVDD.n18809 0.0161121
R43908 DVDD.n18813 DVDD.n18812 0.0161121
R43909 DVDD.n18816 DVDD.n18815 0.0161121
R43910 DVDD.n18801 DVDD.n18798 0.0161121
R43911 DVDD.n18804 DVDD.n18802 0.0161121
R43912 DVDD.n18807 DVDD.n18805 0.0161121
R43913 DVDD.n18810 DVDD.n18808 0.0161121
R43914 DVDD.n18813 DVDD.n18811 0.0161121
R43915 DVDD.n18816 DVDD.n18814 0.0161121
R43916 DVDD.n21050 DVDD.n18817 0.0161121
R43917 DVDD.n18795 DVDD.n18794 0.0161121
R43918 DVDD.n20450 DVDD.n19816 0.0161121
R43919 DVDD.n20452 DVDD.n19815 0.0161121
R43920 DVDD.n20454 DVDD.n19814 0.0161121
R43921 DVDD.n20456 DVDD.n19813 0.0161121
R43922 DVDD.n20458 DVDD.n19812 0.0161121
R43923 DVDD.n20460 DVDD.n19811 0.0161121
R43924 DVDD.n20450 DVDD.n20449 0.0161121
R43925 DVDD.n20452 DVDD.n20451 0.0161121
R43926 DVDD.n20454 DVDD.n20453 0.0161121
R43927 DVDD.n20456 DVDD.n20455 0.0161121
R43928 DVDD.n20458 DVDD.n20457 0.0161121
R43929 DVDD.n20460 DVDD.n20459 0.0161121
R43930 DVDD.n20461 DVDD.n19819 0.0161121
R43931 DVDD.n21026 DVDD.n21025 0.0161121
R43932 DVDD.n21029 DVDD.n21024 0.0161121
R43933 DVDD.n21032 DVDD.n21023 0.0161121
R43934 DVDD.n21035 DVDD.n21022 0.0161121
R43935 DVDD.n21038 DVDD.n21021 0.0161121
R43936 DVDD.n21041 DVDD.n21020 0.0161121
R43937 DVDD.n21049 DVDD.n18818 0.0161121
R43938 DVDD.n21028 DVDD.n21025 0.0161121
R43939 DVDD.n21031 DVDD.n21024 0.0161121
R43940 DVDD.n21034 DVDD.n21023 0.0161121
R43941 DVDD.n21037 DVDD.n21022 0.0161121
R43942 DVDD.n21040 DVDD.n21021 0.0161121
R43943 DVDD.n21043 DVDD.n21020 0.0161121
R43944 DVDD.n20906 DVDD.n18910 0.0161121
R43945 DVDD.n20905 DVDD.n18911 0.0161121
R43946 DVDD.n20904 DVDD.n18912 0.0161121
R43947 DVDD.n20903 DVDD.n18913 0.0161121
R43948 DVDD.n20902 DVDD.n18914 0.0161121
R43949 DVDD.n20901 DVDD.n18915 0.0161121
R43950 DVDD.n20907 DVDD.n18909 0.0161121
R43951 DVDD.n20909 DVDD.n20906 0.0161121
R43952 DVDD.n20911 DVDD.n20905 0.0161121
R43953 DVDD.n20913 DVDD.n20904 0.0161121
R43954 DVDD.n20915 DVDD.n20903 0.0161121
R43955 DVDD.n20917 DVDD.n20902 0.0161121
R43956 DVDD.n20901 DVDD.n18918 0.0161121
R43957 DVDD.n21047 DVDD.n21046 0.0161121
R43958 DVDD.n21047 DVDD.n21045 0.0161121
R43959 DVDD.n20921 DVDD.n18917 0.0161121
R43960 DVDD.n18917 DVDD.n18916 0.0161121
R43961 DVDD.n21068 DVDD.n18750 0.0161121
R43962 DVDD.n21070 DVDD.n18749 0.0161121
R43963 DVDD.n21072 DVDD.n18748 0.0161121
R43964 DVDD.n21074 DVDD.n18747 0.0161121
R43965 DVDD.n21076 DVDD.n18746 0.0161121
R43966 DVDD.n21078 DVDD.n18745 0.0161121
R43967 DVDD.n21080 DVDD.n18744 0.0161121
R43968 DVDD.n21068 DVDD.n21067 0.0161121
R43969 DVDD.n21070 DVDD.n21069 0.0161121
R43970 DVDD.n21072 DVDD.n21071 0.0161121
R43971 DVDD.n21074 DVDD.n21073 0.0161121
R43972 DVDD.n21076 DVDD.n21075 0.0161121
R43973 DVDD.n21078 DVDD.n21077 0.0161121
R43974 DVDD.n21080 DVDD.n21079 0.0161121
R43975 DVDD.n19796 DVDD.n19774 0.0161121
R43976 DVDD.n19795 DVDD.n19775 0.0161121
R43977 DVDD.n19794 DVDD.n19776 0.0161121
R43978 DVDD.n19793 DVDD.n19777 0.0161121
R43979 DVDD.n19792 DVDD.n19778 0.0161121
R43980 DVDD.n19791 DVDD.n19779 0.0161121
R43981 DVDD.n19787 DVDD.n19774 0.0161121
R43982 DVDD.n19786 DVDD.n19775 0.0161121
R43983 DVDD.n19785 DVDD.n19776 0.0161121
R43984 DVDD.n19784 DVDD.n19777 0.0161121
R43985 DVDD.n19783 DVDD.n19778 0.0161121
R43986 DVDD.n19782 DVDD.n19779 0.0161121
R43987 DVDD.n19781 DVDD.n19780 0.0161121
R43988 DVDD.n20994 DVDD.n20993 0.0161121
R43989 DVDD.n20997 DVDD.n20996 0.0161121
R43990 DVDD.n21000 DVDD.n20999 0.0161121
R43991 DVDD.n21003 DVDD.n21002 0.0161121
R43992 DVDD.n21006 DVDD.n21005 0.0161121
R43993 DVDD.n21009 DVDD.n21008 0.0161121
R43994 DVDD.n21013 DVDD.n18823 0.0161121
R43995 DVDD.n20991 DVDD.n20990 0.0161121
R43996 DVDD.n20994 DVDD.n20992 0.0161121
R43997 DVDD.n20997 DVDD.n20995 0.0161121
R43998 DVDD.n21000 DVDD.n20998 0.0161121
R43999 DVDD.n21003 DVDD.n21001 0.0161121
R44000 DVDD.n21006 DVDD.n21004 0.0161121
R44001 DVDD.n21009 DVDD.n21007 0.0161121
R44002 DVDD.n20505 DVDD.n20494 0.0161121
R44003 DVDD.n20507 DVDD.n20493 0.0161121
R44004 DVDD.n20509 DVDD.n20492 0.0161121
R44005 DVDD.n20511 DVDD.n20491 0.0161121
R44006 DVDD.n20513 DVDD.n20490 0.0161121
R44007 DVDD.n20515 DVDD.n20489 0.0161121
R44008 DVDD.n20495 DVDD.n18822 0.0161121
R44009 DVDD.n20517 DVDD.n20497 0.0161121
R44010 DVDD.n20505 DVDD.n20504 0.0161121
R44011 DVDD.n20507 DVDD.n20506 0.0161121
R44012 DVDD.n20509 DVDD.n20508 0.0161121
R44013 DVDD.n20511 DVDD.n20510 0.0161121
R44014 DVDD.n20513 DVDD.n20512 0.0161121
R44015 DVDD.n20515 DVDD.n20514 0.0161121
R44016 DVDD.n20518 DVDD.n20496 0.0161121
R44017 DVDD.n21011 DVDD.n21010 0.0161121
R44018 DVDD.n4602 DVDD.n4601 0.0160415
R44019 DVDD.n3783 DVDD.n3729 0.0160415
R44020 DVDD.n3839 DVDD.n3648 0.0160415
R44021 DVDD.n14299 DVDD.n8605 0.016025
R44022 DVDD.n16269 DVDD.n2361 0.015778
R44023 DVDD.n2997 DVDD.n2769 0.015778
R44024 DVDD.n16313 DVDD.n2485 0.015778
R44025 DVDD.n2926 DVDD.n2791 0.015778
R44026 DVDD.n15908 DVDD.n3260 0.015778
R44027 DVDD.n3161 DVDD.n3059 0.015778
R44028 DVDD.n15679 DVDD.n3431 0.015778
R44029 DVDD.n5158 DVDD.n3107 0.015778
R44030 DVDD.n6399 DVDD.n5997 0.0156579
R44031 DVDD.n8139 DVDD.n8133 0.0156579
R44032 DVDD.n21944 DVDD.n18379 0.015575
R44033 DVDD.n22209 DVDD.n178 0.015575
R44034 DVDD.n22039 DVDD.n18247 0.015575
R44035 DVDD.n22013 DVDD.n223 0.015575
R44036 DVDD.n22229 DVDD.n140 0.015575
R44037 DVDD.n21341 DVDD.n18432 0.015575
R44038 DVDD.n21944 DVDD.n18305 0.015575
R44039 DVDD.n22209 DVDD.n191 0.015575
R44040 DVDD.n22039 DVDD.n18263 0.015575
R44041 DVDD.n18262 DVDD.n223 0.015575
R44042 DVDD.n22229 DVDD.n152 0.015575
R44043 DVDD.n18446 DVDD.n18432 0.015575
R44044 DVDD.n4574 DVDD.n4298 0.015575
R44045 DVDD.n4297 DVDD.n4282 0.015575
R44046 DVDD.n3709 DVDD.n3693 0.015575
R44047 DVDD.n4759 DVDD.n3674 0.015575
R44048 DVDD.n15120 DVDD.n5994 0.0154799
R44049 DVDD.n15114 DVDD.n5994 0.0154799
R44050 DVDD.n6698 DVDD.n6401 0.0154799
R44051 DVDD.n6699 DVDD.n6698 0.0154799
R44052 DVDD.n15099 DVDD.n6393 0.0154799
R44053 DVDD.n15093 DVDD.n6393 0.0154799
R44054 DVDD.n7062 DVDD.n7058 0.0154799
R44055 DVDD.n15077 DVDD.n7058 0.0154799
R44056 DVDD.n15071 DVDD.n7069 0.0154799
R44057 DVDD.n7565 DVDD.n7069 0.0154799
R44058 DVDD.n7565 DVDD.n7456 0.0154799
R44059 DVDD.n14866 DVDD.n7456 0.0154799
R44060 DVDD.n14866 DVDD.n14865 0.0154799
R44061 DVDD.n14865 DVDD.n7568 0.0154799
R44062 DVDD.n9561 DVDD.n9221 0.0154799
R44063 DVDD.n9562 DVDD.n9561 0.0154799
R44064 DVDD.n14848 DVDD.n7681 0.0154799
R44065 DVDD.n14842 DVDD.n7681 0.0154799
R44066 DVDD.n8142 DVDD.n8136 0.0154799
R44067 DVDD.n8147 DVDD.n8142 0.0154799
R44068 DVDD.n8152 DVDD.n8149 0.0154799
R44069 DVDD.n14570 DVDD.n8152 0.0154799
R44070 DVDD.n14570 DVDD.n8153 0.0154799
R44071 DVDD.n8256 DVDD.n8253 0.0154799
R44072 DVDD.n14304 DVDD.n8256 0.0154799
R44073 DVDD.n10229 DVDD.n10225 0.0154799
R44074 DVDD.n10234 DVDD.n10225 0.0154799
R44075 DVDD.n14292 DVDD.n8612 0.0154799
R44076 DVDD.n14286 DVDD.n8612 0.0154799
R44077 DVDD.n10695 DVDD.n10689 0.0154799
R44078 DVDD.n10702 DVDD.n10689 0.0154799
R44079 DVDD.n10703 DVDD.n10702 0.0154799
R44080 DVDD.n10708 DVDD.n10705 0.0154799
R44081 DVDD.n14014 DVDD.n10708 0.0154799
R44082 DVDD.n11221 DVDD.n11220 0.0154799
R44083 DVDD.n11222 DVDD.n11221 0.0154799
R44084 DVDD.n13809 DVDD.n13808 0.0154799
R44085 DVDD.n13808 DVDD.n13807 0.0154799
R44086 DVDD.n13801 DVDD.n11232 0.0154799
R44087 DVDD.n13785 DVDD.n11232 0.0154799
R44088 DVDD.n13779 DVDD.n11587 0.0154799
R44089 DVDD.n13763 DVDD.n11587 0.0154799
R44090 DVDD.n13763 DVDD.n11927 0.0154799
R44091 DVDD.n13756 DVDD.n11935 0.0154799
R44092 DVDD.n12381 DVDD.n11935 0.0154799
R44093 DVDD.n12386 DVDD.n12383 0.0154799
R44094 DVDD.n13489 DVDD.n12386 0.0154799
R44095 DVDD.n12895 DVDD.n12894 0.0154799
R44096 DVDD.n12896 DVDD.n12895 0.0154799
R44097 DVDD.n13279 DVDD.n13278 0.0154799
R44098 DVDD.n13278 DVDD.n13277 0.0154799
R44099 DVDD.n13277 DVDD.n12900 0.0154799
R44100 DVDD.n13270 DVDD.n12911 0.0154799
R44101 DVDD.n12911 DVDD.n12910 0.0154799
R44102 DVDD.n16716 DVDD.n1820 0.0154799
R44103 DVDD.n16717 DVDD.n16716 0.0154799
R44104 DVDD.n16725 DVDD.n1804 0.0154799
R44105 DVDD.n16737 DVDD.n1804 0.0154799
R44106 DVDD.n16739 DVDD.n1705 0.0154799
R44107 DVDD.n17005 DVDD.n1705 0.0154799
R44108 DVDD.n17008 DVDD.n17007 0.0154799
R44109 DVDD.n17007 DVDD.n1270 0.0154799
R44110 DVDD.n17273 DVDD.n1270 0.0154799
R44111 DVDD.n17279 DVDD.n921 0.0154799
R44112 DVDD.n17291 DVDD.n921 0.0154799
R44113 DVDD.n17297 DVDD.n904 0.0154799
R44114 DVDD.n17719 DVDD.n904 0.0154799
R44115 DVDD.n15119 DVDD.n5996 0.0154799
R44116 DVDD.n15115 DVDD.n5996 0.0154799
R44117 DVDD.n6400 DVDD.n6398 0.0154799
R44118 DVDD.n6700 DVDD.n6398 0.0154799
R44119 DVDD.n15098 DVDD.n6395 0.0154799
R44120 DVDD.n15094 DVDD.n6395 0.0154799
R44121 DVDD.n7063 DVDD.n7060 0.0154799
R44122 DVDD.n15076 DVDD.n7060 0.0154799
R44123 DVDD.n15072 DVDD.n7068 0.0154799
R44124 DVDD.n7566 DVDD.n7068 0.0154799
R44125 DVDD.n14868 DVDD.n7566 0.0154799
R44126 DVDD.n14868 DVDD.n14867 0.0154799
R44127 DVDD.n14867 DVDD.n7567 0.0154799
R44128 DVDD.n9569 DVDD.n7567 0.0154799
R44129 DVDD.n9567 DVDD.n9220 0.0154799
R44130 DVDD.n9563 DVDD.n9220 0.0154799
R44131 DVDD.n14847 DVDD.n7683 0.0154799
R44132 DVDD.n14843 DVDD.n7683 0.0154799
R44133 DVDD.n8141 DVDD.n8137 0.0154799
R44134 DVDD.n8141 DVDD.n8134 0.0154799
R44135 DVDD.n14575 DVDD.n8135 0.0154799
R44136 DVDD.n14571 DVDD.n8135 0.0154799
R44137 DVDD.n14571 DVDD.n8151 0.0154799
R44138 DVDD.n14309 DVDD.n8251 0.0154799
R44139 DVDD.n14305 DVDD.n8251 0.0154799
R44140 DVDD.n10228 DVDD.n10224 0.0154799
R44141 DVDD.n10235 DVDD.n10224 0.0154799
R44142 DVDD.n14291 DVDD.n8614 0.0154799
R44143 DVDD.n14287 DVDD.n8614 0.0154799
R44144 DVDD.n10696 DVDD.n10694 0.0154799
R44145 DVDD.n10701 DVDD.n10694 0.0154799
R44146 DVDD.n10701 DVDD.n10687 0.0154799
R44147 DVDD.n14019 DVDD.n10688 0.0154799
R44148 DVDD.n14015 DVDD.n10688 0.0154799
R44149 DVDD.n11219 DVDD.n11214 0.0154799
R44150 DVDD.n11223 DVDD.n11214 0.0154799
R44151 DVDD.n13810 DVDD.n11225 0.0154799
R44152 DVDD.n13806 DVDD.n11225 0.0154799
R44153 DVDD.n13802 DVDD.n11231 0.0154799
R44154 DVDD.n13784 DVDD.n11231 0.0154799
R44155 DVDD.n13780 DVDD.n11586 0.0154799
R44156 DVDD.n13762 DVDD.n11586 0.0154799
R44157 DVDD.n13762 DVDD.n11928 0.0154799
R44158 DVDD.n13757 DVDD.n11933 0.0154799
R44159 DVDD.n12379 DVDD.n11933 0.0154799
R44160 DVDD.n13494 DVDD.n12380 0.0154799
R44161 DVDD.n13490 DVDD.n12380 0.0154799
R44162 DVDD.n12893 DVDD.n12890 0.0154799
R44163 DVDD.n12897 DVDD.n12890 0.0154799
R44164 DVDD.n13280 DVDD.n12899 0.0154799
R44165 DVDD.n13276 DVDD.n12899 0.0154799
R44166 DVDD.n13276 DVDD.n12902 0.0154799
R44167 DVDD.n13271 DVDD.n12907 0.0154799
R44168 DVDD.n12907 DVDD.n2255 0.0154799
R44169 DVDD.n16454 DVDD.n1819 0.0154799
R44170 DVDD.n16718 DVDD.n1819 0.0154799
R44171 DVDD.n16724 DVDD.n1816 0.0154799
R44172 DVDD.n1816 DVDD.n1802 0.0154799
R44173 DVDD.n16743 DVDD.n1803 0.0154799
R44174 DVDD.n1803 DVDD.n1703 0.0154799
R44175 DVDD.n17011 DVDD.n1704 0.0154799
R44176 DVDD.n1704 DVDD.n1269 0.0154799
R44177 DVDD.n17274 DVDD.n1269 0.0154799
R44178 DVDD.n17278 DVDD.n920 0.0154799
R44179 DVDD.n17292 DVDD.n920 0.0154799
R44180 DVDD.n17296 DVDD.n902 0.0154799
R44181 DVDD.n17720 DVDD.n902 0.0154799
R44182 DVDD.n21680 DVDD.n21679 0.0153088
R44183 DVDD.n21679 DVDD.n21675 0.0153088
R44184 DVDD.n21675 DVDD.n183 0.0153088
R44185 DVDD.n18372 DVDD.n184 0.0153088
R44186 DVDD.n18372 DVDD.n18309 0.0153088
R44187 DVDD.n18368 DVDD.n18309 0.0153088
R44188 DVDD.n18343 DVDD.n18335 0.0153088
R44189 DVDD.n18347 DVDD.n18335 0.0153088
R44190 DVDD.n18347 DVDD.n18336 0.0153088
R44191 DVDD.n22001 DVDD.n21996 0.0153088
R44192 DVDD.n22001 DVDD.n21994 0.0153088
R44193 DVDD.n22005 DVDD.n21994 0.0153088
R44194 DVDD.n21268 DVDD.n21267 0.0153088
R44195 DVDD.n21267 DVDD.n21264 0.0153088
R44196 DVDD.n21264 DVDD.n21263 0.0153088
R44197 DVDD.n21337 DVDD.n21336 0.0153088
R44198 DVDD.n21364 DVDD.n21337 0.0153088
R44199 DVDD.n21364 DVDD.n21334 0.0153088
R44200 DVDD.n4849 DVDD.n3548 0.0153088
R44201 DVDD.n4849 DVDD.n3544 0.0153088
R44202 DVDD.n4859 DVDD.n3544 0.0153088
R44203 DVDD.n4863 DVDD.n3535 0.0153088
R44204 DVDD.n4876 DVDD.n3535 0.0153088
R44205 DVDD.n4876 DVDD.n3533 0.0153088
R44206 DVDD.n14308 DVDD.n8250 0.0151165
R44207 DVDD.n10705 DVDD.n10704 0.0149966
R44208 DVDD.n17006 DVDD.n17005 0.0149966
R44209 DVDD.n14020 DVDD.n14019 0.0149966
R44210 DVDD.n17012 DVDD.n1703 0.0149966
R44211 DVDD.n8602 DVDD.n8260 0.014845
R44212 DVDD.n8603 DVDD.n8262 0.014845
R44213 DVDD.n17719 DVDD.n905 0.014755
R44214 DVDD.n17720 DVDD.n903 0.014755
R44215 DVDD.n18614 DVDD.n18611 0.0147105
R44216 DVDD.n13759 DVDD.n13758 0.0145752
R44217 DVDD.n13282 DVDD.n12888 0.0145752
R44218 DVDD.n9788 DVDD.n9663 0.0145488
R44219 DVDD.n9786 DVDD.n9734 0.0145488
R44220 DVDD.n9793 DVDD.n9628 0.0145488
R44221 DVDD.n9796 DVDD.n9795 0.0145488
R44222 DVDD.n13785 DVDD.n11582 0.0145134
R44223 DVDD.n13270 DVDD.n12908 0.0145134
R44224 DVDD.n13784 DVDD.n11583 0.0145134
R44225 DVDD.n13271 DVDD.n12906 0.0145134
R44226 DVDD.n13475 DVDD.n12735 0.014452
R44227 DVDD.n12920 DVDD.n12735 0.014452
R44228 DVDD.n13476 DVDD.n12733 0.014452
R44229 DVDD.n12919 DVDD.n12733 0.014452
R44230 DVDD.n17516 DVDD.n17515 0.01445
R44231 DVDD.n17517 DVDD.n17516 0.01445
R44232 DVDD.n17518 DVDD.n17517 0.01445
R44233 DVDD.n17519 DVDD.n17518 0.01445
R44234 DVDD.n17520 DVDD.n17519 0.01445
R44235 DVDD.n17521 DVDD.n17520 0.01445
R44236 DVDD.n17522 DVDD.n17521 0.01445
R44237 DVDD.n17523 DVDD.n17522 0.01445
R44238 DVDD.n17524 DVDD.n17523 0.01445
R44239 DVDD.n17525 DVDD.n17524 0.01445
R44240 DVDD.n17526 DVDD.n17525 0.01445
R44241 DVDD.n17527 DVDD.n17526 0.01445
R44242 DVDD.n17528 DVDD.n17527 0.01445
R44243 DVDD.n17529 DVDD.n17528 0.01445
R44244 DVDD.n17530 DVDD.n17529 0.01445
R44245 DVDD.n17531 DVDD.n17530 0.01445
R44246 DVDD.n17532 DVDD.n17531 0.01445
R44247 DVDD.n17533 DVDD.n17532 0.01445
R44248 DVDD.n17534 DVDD.n17533 0.01445
R44249 DVDD.n17535 DVDD.n17534 0.01445
R44250 DVDD.n17536 DVDD.n17535 0.01445
R44251 DVDD.n17537 DVDD.n17536 0.01445
R44252 DVDD.n17538 DVDD.n17537 0.01445
R44253 DVDD.n17539 DVDD.n17538 0.01445
R44254 DVDD.n17540 DVDD.n17539 0.01445
R44255 DVDD.n17541 DVDD.n17540 0.01445
R44256 DVDD.n17542 DVDD.n17541 0.01445
R44257 DVDD.n17543 DVDD.n17542 0.01445
R44258 DVDD.n17544 DVDD.n17543 0.01445
R44259 DVDD.n17545 DVDD.n17544 0.01445
R44260 DVDD.n17546 DVDD.n17545 0.01445
R44261 DVDD.n17547 DVDD.n17546 0.01445
R44262 DVDD.n17548 DVDD.n17547 0.01445
R44263 DVDD.n17549 DVDD.n17548 0.01445
R44264 DVDD.n17550 DVDD.n17549 0.01445
R44265 DVDD.n17551 DVDD.n17550 0.01445
R44266 DVDD.n17552 DVDD.n17551 0.01445
R44267 DVDD.n17553 DVDD.n17552 0.01445
R44268 DVDD.n17554 DVDD.n17553 0.01445
R44269 DVDD.n17555 DVDD.n17554 0.01445
R44270 DVDD.n17556 DVDD.n17555 0.01445
R44271 DVDD.n17557 DVDD.n17556 0.01445
R44272 DVDD.n17558 DVDD.n17557 0.01445
R44273 DVDD.n17559 DVDD.n17558 0.01445
R44274 DVDD.n17560 DVDD.n17559 0.01445
R44275 DVDD.n17561 DVDD.n17560 0.01445
R44276 DVDD.n17562 DVDD.n17561 0.01445
R44277 DVDD.n17563 DVDD.n17562 0.01445
R44278 DVDD.n17564 DVDD.n17563 0.01445
R44279 DVDD.n17565 DVDD.n17564 0.01445
R44280 DVDD.n17566 DVDD.n17565 0.01445
R44281 DVDD.n17567 DVDD.n17566 0.01445
R44282 DVDD.n17568 DVDD.n17567 0.01445
R44283 DVDD.n17569 DVDD.n17568 0.01445
R44284 DVDD.n17570 DVDD.n17569 0.01445
R44285 DVDD.n17571 DVDD.n17570 0.01445
R44286 DVDD.n17572 DVDD.n17571 0.01445
R44287 DVDD.n17573 DVDD.n17572 0.01445
R44288 DVDD.n17574 DVDD.n17573 0.01445
R44289 DVDD.n17575 DVDD.n17574 0.01445
R44290 DVDD.n17576 DVDD.n17575 0.01445
R44291 DVDD.n17577 DVDD.n17576 0.01445
R44292 DVDD.n17578 DVDD.n17577 0.01445
R44293 DVDD.n17579 DVDD.n17578 0.01445
R44294 DVDD.n17580 DVDD.n17579 0.01445
R44295 DVDD.n17581 DVDD.n17580 0.01445
R44296 DVDD.n17582 DVDD.n17581 0.01445
R44297 DVDD.n17583 DVDD.n17582 0.01445
R44298 DVDD.n17584 DVDD.n17583 0.01445
R44299 DVDD.n17585 DVDD.n17584 0.01445
R44300 DVDD.n17586 DVDD.n17585 0.01445
R44301 DVDD.n17587 DVDD.n17586 0.01445
R44302 DVDD.n17588 DVDD.n17587 0.01445
R44303 DVDD.n17589 DVDD.n17588 0.01445
R44304 DVDD.n17590 DVDD.n17589 0.01445
R44305 DVDD.n17591 DVDD.n17590 0.01445
R44306 DVDD.n17592 DVDD.n17591 0.01445
R44307 DVDD.n17593 DVDD.n17592 0.01445
R44308 DVDD.n17594 DVDD.n17593 0.01445
R44309 DVDD.n17595 DVDD.n17594 0.01445
R44310 DVDD.n17596 DVDD.n17595 0.01445
R44311 DVDD.n17597 DVDD.n17596 0.01445
R44312 DVDD.n17598 DVDD.n17597 0.01445
R44313 DVDD.n17599 DVDD.n17598 0.01445
R44314 DVDD.n17600 DVDD.n17599 0.01445
R44315 DVDD.n17601 DVDD.n17600 0.01445
R44316 DVDD.n17602 DVDD.n17601 0.01445
R44317 DVDD.n17603 DVDD.n17602 0.01445
R44318 DVDD.n17604 DVDD.n17603 0.01445
R44319 DVDD.n17605 DVDD.n17604 0.01445
R44320 DVDD.n17606 DVDD.n17605 0.01445
R44321 DVDD.n17607 DVDD.n17606 0.01445
R44322 DVDD.n17608 DVDD.n17607 0.01445
R44323 DVDD.n17609 DVDD.n17608 0.01445
R44324 DVDD.n17610 DVDD.n17609 0.01445
R44325 DVDD.n17611 DVDD.n17610 0.01445
R44326 DVDD.n17611 DVDD.n17305 0.01445
R44327 DVDD.n17708 DVDD.n897 0.01445
R44328 DVDD.n17708 DVDD.n17707 0.01445
R44329 DVDD.n17707 DVDD.n17706 0.01445
R44330 DVDD.n17706 DVDD.n17705 0.01445
R44331 DVDD.n17705 DVDD.n17704 0.01445
R44332 DVDD.n17704 DVDD.n17703 0.01445
R44333 DVDD.n17703 DVDD.n17702 0.01445
R44334 DVDD.n17702 DVDD.n17701 0.01445
R44335 DVDD.n17701 DVDD.n17700 0.01445
R44336 DVDD.n17700 DVDD.n17699 0.01445
R44337 DVDD.n17699 DVDD.n17698 0.01445
R44338 DVDD.n17698 DVDD.n17697 0.01445
R44339 DVDD.n17697 DVDD.n17696 0.01445
R44340 DVDD.n17696 DVDD.n17695 0.01445
R44341 DVDD.n17695 DVDD.n17694 0.01445
R44342 DVDD.n17694 DVDD.n17693 0.01445
R44343 DVDD.n17693 DVDD.n17692 0.01445
R44344 DVDD.n17692 DVDD.n17691 0.01445
R44345 DVDD.n17691 DVDD.n17690 0.01445
R44346 DVDD.n17690 DVDD.n17689 0.01445
R44347 DVDD.n17689 DVDD.n17688 0.01445
R44348 DVDD.n17688 DVDD.n17687 0.01445
R44349 DVDD.n17687 DVDD.n17686 0.01445
R44350 DVDD.n17686 DVDD.n17685 0.01445
R44351 DVDD.n17685 DVDD.n17684 0.01445
R44352 DVDD.n17684 DVDD.n17683 0.01445
R44353 DVDD.n17683 DVDD.n17682 0.01445
R44354 DVDD.n17682 DVDD.n17681 0.01445
R44355 DVDD.n17681 DVDD.n17680 0.01445
R44356 DVDD.n17680 DVDD.n17679 0.01445
R44357 DVDD.n17679 DVDD.n17678 0.01445
R44358 DVDD.n17678 DVDD.n17677 0.01445
R44359 DVDD.n17677 DVDD.n17676 0.01445
R44360 DVDD.n17676 DVDD.n17675 0.01445
R44361 DVDD.n17675 DVDD.n17674 0.01445
R44362 DVDD.n17674 DVDD.n17673 0.01445
R44363 DVDD.n17673 DVDD.n17672 0.01445
R44364 DVDD.n17672 DVDD.n17671 0.01445
R44365 DVDD.n17671 DVDD.n17670 0.01445
R44366 DVDD.n17670 DVDD.n17669 0.01445
R44367 DVDD.n17669 DVDD.n17668 0.01445
R44368 DVDD.n17668 DVDD.n17667 0.01445
R44369 DVDD.n17667 DVDD.n17666 0.01445
R44370 DVDD.n17666 DVDD.n17665 0.01445
R44371 DVDD.n17665 DVDD.n17664 0.01445
R44372 DVDD.n17664 DVDD.n17663 0.01445
R44373 DVDD.n17663 DVDD.n17662 0.01445
R44374 DVDD.n17662 DVDD.n17661 0.01445
R44375 DVDD.n17661 DVDD.n17660 0.01445
R44376 DVDD.n17660 DVDD.n17659 0.01445
R44377 DVDD.n17659 DVDD.n17658 0.01445
R44378 DVDD.n17658 DVDD.n17657 0.01445
R44379 DVDD.n17657 DVDD.n17656 0.01445
R44380 DVDD.n17656 DVDD.n17655 0.01445
R44381 DVDD.n17655 DVDD.n17654 0.01445
R44382 DVDD.n17654 DVDD.n17653 0.01445
R44383 DVDD.n17653 DVDD.n17652 0.01445
R44384 DVDD.n17652 DVDD.n17651 0.01445
R44385 DVDD.n17651 DVDD.n17650 0.01445
R44386 DVDD.n17650 DVDD.n17649 0.01445
R44387 DVDD.n17649 DVDD.n17648 0.01445
R44388 DVDD.n17648 DVDD.n17647 0.01445
R44389 DVDD.n17647 DVDD.n17646 0.01445
R44390 DVDD.n17646 DVDD.n17645 0.01445
R44391 DVDD.n17645 DVDD.n17644 0.01445
R44392 DVDD.n17644 DVDD.n17643 0.01445
R44393 DVDD.n17643 DVDD.n17642 0.01445
R44394 DVDD.n17642 DVDD.n17641 0.01445
R44395 DVDD.n17641 DVDD.n17640 0.01445
R44396 DVDD.n17640 DVDD.n17639 0.01445
R44397 DVDD.n17639 DVDD.n17638 0.01445
R44398 DVDD.n17638 DVDD.n17637 0.01445
R44399 DVDD.n17637 DVDD.n17636 0.01445
R44400 DVDD.n17636 DVDD.n17635 0.01445
R44401 DVDD.n17635 DVDD.n17634 0.01445
R44402 DVDD.n17634 DVDD.n17633 0.01445
R44403 DVDD.n17633 DVDD.n17632 0.01445
R44404 DVDD.n17632 DVDD.n17631 0.01445
R44405 DVDD.n17631 DVDD.n17630 0.01445
R44406 DVDD.n17630 DVDD.n17629 0.01445
R44407 DVDD.n17629 DVDD.n17628 0.01445
R44408 DVDD.n17628 DVDD.n17627 0.01445
R44409 DVDD.n17627 DVDD.n17626 0.01445
R44410 DVDD.n17626 DVDD.n17625 0.01445
R44411 DVDD.n17625 DVDD.n17624 0.01445
R44412 DVDD.n17624 DVDD.n17623 0.01445
R44413 DVDD.n17623 DVDD.n17622 0.01445
R44414 DVDD.n17622 DVDD.n17621 0.01445
R44415 DVDD.n17621 DVDD.n17620 0.01445
R44416 DVDD.n17620 DVDD.n17619 0.01445
R44417 DVDD.n17619 DVDD.n17618 0.01445
R44418 DVDD.n17618 DVDD.n17617 0.01445
R44419 DVDD.n17617 DVDD.n17616 0.01445
R44420 DVDD.n17616 DVDD.n17615 0.01445
R44421 DVDD.n17615 DVDD.n17614 0.01445
R44422 DVDD.n17614 DVDD.n17613 0.01445
R44423 DVDD.n17613 DVDD.n17612 0.01445
R44424 DVDD.n15133 DVDD.n5583 0.01445
R44425 DVDD.n15133 DVDD.n5589 0.01445
R44426 DVDD.n5790 DVDD.n5589 0.01445
R44427 DVDD.n5790 DVDD.n5789 0.01445
R44428 DVDD.n5794 DVDD.n5789 0.01445
R44429 DVDD.n5795 DVDD.n5794 0.01445
R44430 DVDD.n5796 DVDD.n5795 0.01445
R44431 DVDD.n5796 DVDD.n5787 0.01445
R44432 DVDD.n5800 DVDD.n5787 0.01445
R44433 DVDD.n5801 DVDD.n5800 0.01445
R44434 DVDD.n5802 DVDD.n5801 0.01445
R44435 DVDD.n5802 DVDD.n5785 0.01445
R44436 DVDD.n5806 DVDD.n5785 0.01445
R44437 DVDD.n5807 DVDD.n5806 0.01445
R44438 DVDD.n5808 DVDD.n5807 0.01445
R44439 DVDD.n5808 DVDD.n5783 0.01445
R44440 DVDD.n5812 DVDD.n5783 0.01445
R44441 DVDD.n5813 DVDD.n5812 0.01445
R44442 DVDD.n5814 DVDD.n5813 0.01445
R44443 DVDD.n5814 DVDD.n5781 0.01445
R44444 DVDD.n5818 DVDD.n5781 0.01445
R44445 DVDD.n5819 DVDD.n5818 0.01445
R44446 DVDD.n5820 DVDD.n5819 0.01445
R44447 DVDD.n5820 DVDD.n5779 0.01445
R44448 DVDD.n5824 DVDD.n5779 0.01445
R44449 DVDD.n5825 DVDD.n5824 0.01445
R44450 DVDD.n5826 DVDD.n5825 0.01445
R44451 DVDD.n5826 DVDD.n5777 0.01445
R44452 DVDD.n5830 DVDD.n5777 0.01445
R44453 DVDD.n5831 DVDD.n5830 0.01445
R44454 DVDD.n5832 DVDD.n5831 0.01445
R44455 DVDD.n5832 DVDD.n5775 0.01445
R44456 DVDD.n5836 DVDD.n5775 0.01445
R44457 DVDD.n5837 DVDD.n5836 0.01445
R44458 DVDD.n5838 DVDD.n5837 0.01445
R44459 DVDD.n5838 DVDD.n5773 0.01445
R44460 DVDD.n5842 DVDD.n5773 0.01445
R44461 DVDD.n5843 DVDD.n5842 0.01445
R44462 DVDD.n5844 DVDD.n5843 0.01445
R44463 DVDD.n5844 DVDD.n5771 0.01445
R44464 DVDD.n5848 DVDD.n5771 0.01445
R44465 DVDD.n5849 DVDD.n5848 0.01445
R44466 DVDD.n5850 DVDD.n5849 0.01445
R44467 DVDD.n5850 DVDD.n5769 0.01445
R44468 DVDD.n5854 DVDD.n5769 0.01445
R44469 DVDD.n5855 DVDD.n5854 0.01445
R44470 DVDD.n5856 DVDD.n5855 0.01445
R44471 DVDD.n5856 DVDD.n5767 0.01445
R44472 DVDD.n5860 DVDD.n5767 0.01445
R44473 DVDD.n5861 DVDD.n5860 0.01445
R44474 DVDD.n5862 DVDD.n5861 0.01445
R44475 DVDD.n5862 DVDD.n5765 0.01445
R44476 DVDD.n5866 DVDD.n5765 0.01445
R44477 DVDD.n5867 DVDD.n5866 0.01445
R44478 DVDD.n5868 DVDD.n5867 0.01445
R44479 DVDD.n5868 DVDD.n5763 0.01445
R44480 DVDD.n5872 DVDD.n5763 0.01445
R44481 DVDD.n5873 DVDD.n5872 0.01445
R44482 DVDD.n5874 DVDD.n5873 0.01445
R44483 DVDD.n5874 DVDD.n5761 0.01445
R44484 DVDD.n5878 DVDD.n5761 0.01445
R44485 DVDD.n5879 DVDD.n5878 0.01445
R44486 DVDD.n5880 DVDD.n5879 0.01445
R44487 DVDD.n5880 DVDD.n5759 0.01445
R44488 DVDD.n5884 DVDD.n5759 0.01445
R44489 DVDD.n5885 DVDD.n5884 0.01445
R44490 DVDD.n5886 DVDD.n5885 0.01445
R44491 DVDD.n5886 DVDD.n5757 0.01445
R44492 DVDD.n5890 DVDD.n5757 0.01445
R44493 DVDD.n5891 DVDD.n5890 0.01445
R44494 DVDD.n5892 DVDD.n5891 0.01445
R44495 DVDD.n5892 DVDD.n5755 0.01445
R44496 DVDD.n5896 DVDD.n5755 0.01445
R44497 DVDD.n5897 DVDD.n5896 0.01445
R44498 DVDD.n5898 DVDD.n5897 0.01445
R44499 DVDD.n5898 DVDD.n5753 0.01445
R44500 DVDD.n5902 DVDD.n5753 0.01445
R44501 DVDD.n5903 DVDD.n5902 0.01445
R44502 DVDD.n5904 DVDD.n5903 0.01445
R44503 DVDD.n5904 DVDD.n5751 0.01445
R44504 DVDD.n5908 DVDD.n5751 0.01445
R44505 DVDD.n5909 DVDD.n5908 0.01445
R44506 DVDD.n5910 DVDD.n5909 0.01445
R44507 DVDD.n5910 DVDD.n5749 0.01445
R44508 DVDD.n5914 DVDD.n5749 0.01445
R44509 DVDD.n5915 DVDD.n5914 0.01445
R44510 DVDD.n5916 DVDD.n5915 0.01445
R44511 DVDD.n5916 DVDD.n5747 0.01445
R44512 DVDD.n5920 DVDD.n5747 0.01445
R44513 DVDD.n5921 DVDD.n5920 0.01445
R44514 DVDD.n5922 DVDD.n5921 0.01445
R44515 DVDD.n5922 DVDD.n5745 0.01445
R44516 DVDD.n5926 DVDD.n5745 0.01445
R44517 DVDD.n5927 DVDD.n5926 0.01445
R44518 DVDD.n5928 DVDD.n5927 0.01445
R44519 DVDD.n5928 DVDD.n5742 0.01445
R44520 DVDD.n15129 DVDD.n5742 0.01445
R44521 DVDD.n15135 DVDD.n15134 0.01445
R44522 DVDD.n15134 DVDD.n5588 0.01445
R44523 DVDD.n5791 DVDD.n5588 0.01445
R44524 DVDD.n5792 DVDD.n5791 0.01445
R44525 DVDD.n5793 DVDD.n5792 0.01445
R44526 DVDD.n5793 DVDD.n5788 0.01445
R44527 DVDD.n5797 DVDD.n5788 0.01445
R44528 DVDD.n5798 DVDD.n5797 0.01445
R44529 DVDD.n5799 DVDD.n5798 0.01445
R44530 DVDD.n5799 DVDD.n5786 0.01445
R44531 DVDD.n5803 DVDD.n5786 0.01445
R44532 DVDD.n5804 DVDD.n5803 0.01445
R44533 DVDD.n5805 DVDD.n5804 0.01445
R44534 DVDD.n5805 DVDD.n5784 0.01445
R44535 DVDD.n5809 DVDD.n5784 0.01445
R44536 DVDD.n5810 DVDD.n5809 0.01445
R44537 DVDD.n5811 DVDD.n5810 0.01445
R44538 DVDD.n5811 DVDD.n5782 0.01445
R44539 DVDD.n5815 DVDD.n5782 0.01445
R44540 DVDD.n5816 DVDD.n5815 0.01445
R44541 DVDD.n5817 DVDD.n5816 0.01445
R44542 DVDD.n5817 DVDD.n5780 0.01445
R44543 DVDD.n5821 DVDD.n5780 0.01445
R44544 DVDD.n5822 DVDD.n5821 0.01445
R44545 DVDD.n5823 DVDD.n5822 0.01445
R44546 DVDD.n5823 DVDD.n5778 0.01445
R44547 DVDD.n5827 DVDD.n5778 0.01445
R44548 DVDD.n5828 DVDD.n5827 0.01445
R44549 DVDD.n5829 DVDD.n5828 0.01445
R44550 DVDD.n5829 DVDD.n5776 0.01445
R44551 DVDD.n5833 DVDD.n5776 0.01445
R44552 DVDD.n5834 DVDD.n5833 0.01445
R44553 DVDD.n5835 DVDD.n5834 0.01445
R44554 DVDD.n5835 DVDD.n5774 0.01445
R44555 DVDD.n5839 DVDD.n5774 0.01445
R44556 DVDD.n5840 DVDD.n5839 0.01445
R44557 DVDD.n5841 DVDD.n5840 0.01445
R44558 DVDD.n5841 DVDD.n5772 0.01445
R44559 DVDD.n5845 DVDD.n5772 0.01445
R44560 DVDD.n5846 DVDD.n5845 0.01445
R44561 DVDD.n5847 DVDD.n5846 0.01445
R44562 DVDD.n5847 DVDD.n5770 0.01445
R44563 DVDD.n5851 DVDD.n5770 0.01445
R44564 DVDD.n5852 DVDD.n5851 0.01445
R44565 DVDD.n5853 DVDD.n5852 0.01445
R44566 DVDD.n5853 DVDD.n5768 0.01445
R44567 DVDD.n5857 DVDD.n5768 0.01445
R44568 DVDD.n5858 DVDD.n5857 0.01445
R44569 DVDD.n5859 DVDD.n5858 0.01445
R44570 DVDD.n5859 DVDD.n5766 0.01445
R44571 DVDD.n5863 DVDD.n5766 0.01445
R44572 DVDD.n5864 DVDD.n5863 0.01445
R44573 DVDD.n5865 DVDD.n5864 0.01445
R44574 DVDD.n5865 DVDD.n5764 0.01445
R44575 DVDD.n5869 DVDD.n5764 0.01445
R44576 DVDD.n5870 DVDD.n5869 0.01445
R44577 DVDD.n5871 DVDD.n5870 0.01445
R44578 DVDD.n5871 DVDD.n5762 0.01445
R44579 DVDD.n5875 DVDD.n5762 0.01445
R44580 DVDD.n5876 DVDD.n5875 0.01445
R44581 DVDD.n5877 DVDD.n5876 0.01445
R44582 DVDD.n5877 DVDD.n5760 0.01445
R44583 DVDD.n5881 DVDD.n5760 0.01445
R44584 DVDD.n5882 DVDD.n5881 0.01445
R44585 DVDD.n5883 DVDD.n5882 0.01445
R44586 DVDD.n5883 DVDD.n5758 0.01445
R44587 DVDD.n5887 DVDD.n5758 0.01445
R44588 DVDD.n5888 DVDD.n5887 0.01445
R44589 DVDD.n5889 DVDD.n5888 0.01445
R44590 DVDD.n5889 DVDD.n5756 0.01445
R44591 DVDD.n5893 DVDD.n5756 0.01445
R44592 DVDD.n5894 DVDD.n5893 0.01445
R44593 DVDD.n5895 DVDD.n5894 0.01445
R44594 DVDD.n5895 DVDD.n5754 0.01445
R44595 DVDD.n5899 DVDD.n5754 0.01445
R44596 DVDD.n5900 DVDD.n5899 0.01445
R44597 DVDD.n5901 DVDD.n5900 0.01445
R44598 DVDD.n5901 DVDD.n5752 0.01445
R44599 DVDD.n5905 DVDD.n5752 0.01445
R44600 DVDD.n5906 DVDD.n5905 0.01445
R44601 DVDD.n5907 DVDD.n5906 0.01445
R44602 DVDD.n5907 DVDD.n5750 0.01445
R44603 DVDD.n5911 DVDD.n5750 0.01445
R44604 DVDD.n5912 DVDD.n5911 0.01445
R44605 DVDD.n5913 DVDD.n5912 0.01445
R44606 DVDD.n5913 DVDD.n5748 0.01445
R44607 DVDD.n5917 DVDD.n5748 0.01445
R44608 DVDD.n5918 DVDD.n5917 0.01445
R44609 DVDD.n5919 DVDD.n5918 0.01445
R44610 DVDD.n5919 DVDD.n5746 0.01445
R44611 DVDD.n5923 DVDD.n5746 0.01445
R44612 DVDD.n5924 DVDD.n5923 0.01445
R44613 DVDD.n5925 DVDD.n5924 0.01445
R44614 DVDD.n5925 DVDD.n5744 0.01445
R44615 DVDD.n5929 DVDD.n5744 0.01445
R44616 DVDD.n5930 DVDD.n5929 0.01445
R44617 DVDD.n15128 DVDD.n5930 0.01445
R44618 DVDD.n900 DVDD.n893 0.0143045
R44619 DVDD.n7673 DVDD.n7672 0.014225
R44620 DVDD.n4994 DVDD.n4906 0.0141679
R44621 DVDD.n4991 DVDD.n4985 0.0141679
R44622 DVDD.n4989 DVDD.n4986 0.0141679
R44623 DVDD.n4989 DVDD.n4984 0.0141679
R44624 DVDD.n4993 DVDD.n4988 0.0141679
R44625 DVDD.n4988 DVDD.n4983 0.0141679
R44626 DVDD.n4998 DVDD.n4982 0.0141679
R44627 DVDD.n4916 DVDD.n4907 0.0141679
R44628 DVDD.n4917 DVDD.n4916 0.0141679
R44629 DVDD.n4918 DVDD.n4915 0.0141679
R44630 DVDD.n4920 DVDD.n4915 0.0141679
R44631 DVDD.n4921 DVDD.n4914 0.0141679
R44632 DVDD.n4923 DVDD.n4914 0.0141679
R44633 DVDD.n4924 DVDD.n4913 0.0141679
R44634 DVDD.n4926 DVDD.n4913 0.0141679
R44635 DVDD.n4927 DVDD.n4912 0.0141679
R44636 DVDD.n4929 DVDD.n4912 0.0141679
R44637 DVDD.n4930 DVDD.n4911 0.0141679
R44638 DVDD.n4932 DVDD.n4911 0.0141679
R44639 DVDD.n4933 DVDD.n4910 0.0141679
R44640 DVDD.n4935 DVDD.n4910 0.0141679
R44641 DVDD.n4936 DVDD.n4909 0.0141679
R44642 DVDD.n4938 DVDD.n4909 0.0141679
R44643 DVDD.n4939 DVDD.n4908 0.0141679
R44644 DVDD.n4941 DVDD.n4908 0.0141679
R44645 DVDD.n4952 DVDD.n4942 0.0141679
R44646 DVDD.n4955 DVDD.n4953 0.0141679
R44647 DVDD.n4954 DVDD.n4951 0.0141679
R44648 DVDD.n4958 DVDD.n4956 0.0141679
R44649 DVDD.n4957 DVDD.n4950 0.0141679
R44650 DVDD.n4961 DVDD.n4959 0.0141679
R44651 DVDD.n4960 DVDD.n4949 0.0141679
R44652 DVDD.n4964 DVDD.n4962 0.0141679
R44653 DVDD.n4963 DVDD.n4948 0.0141679
R44654 DVDD.n4967 DVDD.n4965 0.0141679
R44655 DVDD.n4966 DVDD.n4947 0.0141679
R44656 DVDD.n4970 DVDD.n4968 0.0141679
R44657 DVDD.n4969 DVDD.n4946 0.0141679
R44658 DVDD.n4973 DVDD.n4971 0.0141679
R44659 DVDD.n4972 DVDD.n4945 0.0141679
R44660 DVDD.n4976 DVDD.n4974 0.0141679
R44661 DVDD.n4975 DVDD.n4944 0.0141679
R44662 DVDD.n4943 DVDD.n2293 0.0141679
R44663 DVDD.n2305 DVDD.n2295 0.0141679
R44664 DVDD.n2307 DVDD.n2305 0.0141679
R44665 DVDD.n2333 DVDD.n2304 0.0141679
R44666 DVDD.n2309 DVDD.n2304 0.0141679
R44667 DVDD.n2332 DVDD.n2303 0.0141679
R44668 DVDD.n2311 DVDD.n2303 0.0141679
R44669 DVDD.n2331 DVDD.n2302 0.0141679
R44670 DVDD.n2313 DVDD.n2302 0.0141679
R44671 DVDD.n2330 DVDD.n2301 0.0141679
R44672 DVDD.n2315 DVDD.n2301 0.0141679
R44673 DVDD.n2329 DVDD.n2300 0.0141679
R44674 DVDD.n2317 DVDD.n2300 0.0141679
R44675 DVDD.n2328 DVDD.n2299 0.0141679
R44676 DVDD.n2319 DVDD.n2299 0.0141679
R44677 DVDD.n2327 DVDD.n2298 0.0141679
R44678 DVDD.n2321 DVDD.n2298 0.0141679
R44679 DVDD.n2326 DVDD.n2297 0.0141679
R44680 DVDD.n2323 DVDD.n2297 0.0141679
R44681 DVDD.n2456 DVDD.n2446 0.0141679
R44682 DVDD.n2457 DVDD.n2456 0.0141679
R44683 DVDD.n2455 DVDD.n2445 0.0141679
R44684 DVDD.n2459 DVDD.n2455 0.0141679
R44685 DVDD.n2454 DVDD.n2444 0.0141679
R44686 DVDD.n2461 DVDD.n2454 0.0141679
R44687 DVDD.n2453 DVDD.n2443 0.0141679
R44688 DVDD.n2463 DVDD.n2453 0.0141679
R44689 DVDD.n2452 DVDD.n2442 0.0141679
R44690 DVDD.n2465 DVDD.n2452 0.0141679
R44691 DVDD.n2451 DVDD.n2441 0.0141679
R44692 DVDD.n2467 DVDD.n2451 0.0141679
R44693 DVDD.n2450 DVDD.n2440 0.0141679
R44694 DVDD.n2469 DVDD.n2450 0.0141679
R44695 DVDD.n2449 DVDD.n2439 0.0141679
R44696 DVDD.n2471 DVDD.n2449 0.0141679
R44697 DVDD.n2448 DVDD.n2438 0.0141679
R44698 DVDD.n2448 DVDD.n2447 0.0141679
R44699 DVDD.n18025 DVDD.n547 0.0141679
R44700 DVDD.n18026 DVDD.n18025 0.0141679
R44701 DVDD.n18028 DVDD.n548 0.0141679
R44702 DVDD.n18029 DVDD.n18028 0.0141679
R44703 DVDD.n18031 DVDD.n549 0.0141679
R44704 DVDD.n18033 DVDD.n542 0.0141679
R44705 DVDD.n545 DVDD.n542 0.0141679
R44706 DVDD.n4953 DVDD.n4952 0.0141679
R44707 DVDD.n4956 DVDD.n4951 0.0141679
R44708 DVDD.n4959 DVDD.n4950 0.0141679
R44709 DVDD.n4962 DVDD.n4949 0.0141679
R44710 DVDD.n4965 DVDD.n4948 0.0141679
R44711 DVDD.n4968 DVDD.n4947 0.0141679
R44712 DVDD.n4971 DVDD.n4946 0.0141679
R44713 DVDD.n4974 DVDD.n4945 0.0141679
R44714 DVDD.n4944 DVDD.n4943 0.0141679
R44715 DVDD.n16399 DVDD.n2295 0.0141679
R44716 DVDD.n2333 DVDD.n2308 0.0141679
R44717 DVDD.n2332 DVDD.n2310 0.0141679
R44718 DVDD.n2331 DVDD.n2312 0.0141679
R44719 DVDD.n2330 DVDD.n2314 0.0141679
R44720 DVDD.n2329 DVDD.n2316 0.0141679
R44721 DVDD.n2328 DVDD.n2318 0.0141679
R44722 DVDD.n2327 DVDD.n2320 0.0141679
R44723 DVDD.n2326 DVDD.n2322 0.0141679
R44724 DVDD.n2446 DVDD.n2324 0.0141679
R44725 DVDD.n2458 DVDD.n2445 0.0141679
R44726 DVDD.n2460 DVDD.n2444 0.0141679
R44727 DVDD.n2462 DVDD.n2443 0.0141679
R44728 DVDD.n2464 DVDD.n2442 0.0141679
R44729 DVDD.n2466 DVDD.n2441 0.0141679
R44730 DVDD.n2468 DVDD.n2440 0.0141679
R44731 DVDD.n2470 DVDD.n2439 0.0141679
R44732 DVDD.n2472 DVDD.n2438 0.0141679
R44733 DVDD.n4978 DVDD.n4942 0.0141679
R44734 DVDD.n4955 DVDD.n4954 0.0141679
R44735 DVDD.n4958 DVDD.n4957 0.0141679
R44736 DVDD.n4961 DVDD.n4960 0.0141679
R44737 DVDD.n4964 DVDD.n4963 0.0141679
R44738 DVDD.n4967 DVDD.n4966 0.0141679
R44739 DVDD.n4970 DVDD.n4969 0.0141679
R44740 DVDD.n4973 DVDD.n4972 0.0141679
R44741 DVDD.n4976 DVDD.n4975 0.0141679
R44742 DVDD.n2308 DVDD.n2307 0.0141679
R44743 DVDD.n2310 DVDD.n2309 0.0141679
R44744 DVDD.n2312 DVDD.n2311 0.0141679
R44745 DVDD.n2314 DVDD.n2313 0.0141679
R44746 DVDD.n2316 DVDD.n2315 0.0141679
R44747 DVDD.n2318 DVDD.n2317 0.0141679
R44748 DVDD.n2320 DVDD.n2319 0.0141679
R44749 DVDD.n2322 DVDD.n2321 0.0141679
R44750 DVDD.n16397 DVDD.n2323 0.0141679
R44751 DVDD.n2458 DVDD.n2457 0.0141679
R44752 DVDD.n2460 DVDD.n2459 0.0141679
R44753 DVDD.n2462 DVDD.n2461 0.0141679
R44754 DVDD.n2464 DVDD.n2463 0.0141679
R44755 DVDD.n2466 DVDD.n2465 0.0141679
R44756 DVDD.n2468 DVDD.n2467 0.0141679
R44757 DVDD.n2470 DVDD.n2469 0.0141679
R44758 DVDD.n2472 DVDD.n2471 0.0141679
R44759 DVDD.n2474 DVDD.n2447 0.0141679
R44760 DVDD.n4990 DVDD.n4984 0.0141679
R44761 DVDD.n4999 DVDD.n4983 0.0141679
R44762 DVDD.n4991 DVDD.n4906 0.0141679
R44763 DVDD.n4993 DVDD.n4990 0.0141679
R44764 DVDD.n4999 DVDD.n4998 0.0141679
R44765 DVDD.n4995 DVDD.n4994 0.0141679
R44766 DVDD.n5001 DVDD.n4986 0.0141679
R44767 DVDD.n15148 DVDD.n5561 0.0141679
R44768 DVDD.n15146 DVDD.n5562 0.0141679
R44769 DVDD.n5575 DVDD.n5567 0.0141679
R44770 DVDD.n5576 DVDD.n5575 0.0141679
R44771 DVDD.n5573 DVDD.n5572 0.0141679
R44772 DVDD.n5572 DVDD.n5571 0.0141679
R44773 DVDD.n5569 DVDD.n5568 0.0141679
R44774 DVDD.n10176 DVDD.n10175 0.0141679
R44775 DVDD.n10178 DVDD.n10175 0.0141679
R44776 DVDD.n10179 DVDD.n10174 0.0141679
R44777 DVDD.n10181 DVDD.n10174 0.0141679
R44778 DVDD.n10182 DVDD.n10173 0.0141679
R44779 DVDD.n10184 DVDD.n10173 0.0141679
R44780 DVDD.n10185 DVDD.n10172 0.0141679
R44781 DVDD.n10187 DVDD.n10172 0.0141679
R44782 DVDD.n10188 DVDD.n10171 0.0141679
R44783 DVDD.n10190 DVDD.n10171 0.0141679
R44784 DVDD.n10191 DVDD.n10170 0.0141679
R44785 DVDD.n10193 DVDD.n10170 0.0141679
R44786 DVDD.n10194 DVDD.n10169 0.0141679
R44787 DVDD.n10196 DVDD.n10169 0.0141679
R44788 DVDD.n10199 DVDD.n10198 0.0141679
R44789 DVDD.n10201 DVDD.n10200 0.0141679
R44790 DVDD.n8970 DVDD.n8958 0.0141679
R44791 DVDD.n10205 DVDD.n8970 0.0141679
R44792 DVDD.n8969 DVDD.n8957 0.0141679
R44793 DVDD.n10207 DVDD.n8969 0.0141679
R44794 DVDD.n8968 DVDD.n8956 0.0141679
R44795 DVDD.n10209 DVDD.n8968 0.0141679
R44796 DVDD.n8967 DVDD.n8955 0.0141679
R44797 DVDD.n10211 DVDD.n8967 0.0141679
R44798 DVDD.n8966 DVDD.n8954 0.0141679
R44799 DVDD.n10213 DVDD.n8966 0.0141679
R44800 DVDD.n8965 DVDD.n8953 0.0141679
R44801 DVDD.n10215 DVDD.n8965 0.0141679
R44802 DVDD.n8964 DVDD.n8952 0.0141679
R44803 DVDD.n10217 DVDD.n8964 0.0141679
R44804 DVDD.n8959 DVDD.n8951 0.0141679
R44805 DVDD.n10221 DVDD.n10220 0.0141679
R44806 DVDD.n16405 DVDD.n2290 0.0141679
R44807 DVDD.n16407 DVDD.n2290 0.0141679
R44808 DVDD.n16408 DVDD.n2289 0.0141679
R44809 DVDD.n16410 DVDD.n2289 0.0141679
R44810 DVDD.n16411 DVDD.n2288 0.0141679
R44811 DVDD.n16413 DVDD.n2288 0.0141679
R44812 DVDD.n16414 DVDD.n2287 0.0141679
R44813 DVDD.n16416 DVDD.n2287 0.0141679
R44814 DVDD.n16417 DVDD.n2286 0.0141679
R44815 DVDD.n16419 DVDD.n2286 0.0141679
R44816 DVDD.n16420 DVDD.n2285 0.0141679
R44817 DVDD.n16422 DVDD.n2285 0.0141679
R44818 DVDD.n16423 DVDD.n2284 0.0141679
R44819 DVDD.n16425 DVDD.n2284 0.0141679
R44820 DVDD.n16428 DVDD.n16427 0.0141679
R44821 DVDD.n16430 DVDD.n16429 0.0141679
R44822 DVDD.n2277 DVDD.n2264 0.0141679
R44823 DVDD.n16434 DVDD.n2277 0.0141679
R44824 DVDD.n2276 DVDD.n2263 0.0141679
R44825 DVDD.n16436 DVDD.n2276 0.0141679
R44826 DVDD.n2275 DVDD.n2262 0.0141679
R44827 DVDD.n16438 DVDD.n2275 0.0141679
R44828 DVDD.n2274 DVDD.n2261 0.0141679
R44829 DVDD.n16440 DVDD.n2274 0.0141679
R44830 DVDD.n2273 DVDD.n2260 0.0141679
R44831 DVDD.n16442 DVDD.n2273 0.0141679
R44832 DVDD.n2272 DVDD.n2259 0.0141679
R44833 DVDD.n16444 DVDD.n2272 0.0141679
R44834 DVDD.n2271 DVDD.n2258 0.0141679
R44835 DVDD.n16446 DVDD.n2271 0.0141679
R44836 DVDD.n2269 DVDD.n2257 0.0141679
R44837 DVDD.n16448 DVDD.n2265 0.0141679
R44838 DVDD.n17733 DVDD.n881 0.0141679
R44839 DVDD.n17732 DVDD.n879 0.0141679
R44840 DVDD.n887 DVDD.n879 0.0141679
R44841 DVDD.n883 DVDD.n878 0.0141679
R44842 DVDD.n17735 DVDD.n878 0.0141679
R44843 DVDD.n17728 DVDD.n889 0.0141679
R44844 DVDD.n17729 DVDD.n17728 0.0141679
R44845 DVDD.n15148 DVDD.n5562 0.0141679
R44846 DVDD.n5576 DVDD.n5574 0.0141679
R44847 DVDD.n5571 DVDD.n5570 0.0141679
R44848 DVDD.n10204 DVDD.n8958 0.0141679
R44849 DVDD.n10206 DVDD.n8957 0.0141679
R44850 DVDD.n10208 DVDD.n8956 0.0141679
R44851 DVDD.n10210 DVDD.n8955 0.0141679
R44852 DVDD.n10212 DVDD.n8954 0.0141679
R44853 DVDD.n10214 DVDD.n8953 0.0141679
R44854 DVDD.n10216 DVDD.n8952 0.0141679
R44855 DVDD.n10218 DVDD.n8951 0.0141679
R44856 DVDD.n16406 DVDD.n16405 0.0141679
R44857 DVDD.n16409 DVDD.n16408 0.0141679
R44858 DVDD.n16412 DVDD.n16411 0.0141679
R44859 DVDD.n16415 DVDD.n16414 0.0141679
R44860 DVDD.n16418 DVDD.n16417 0.0141679
R44861 DVDD.n16421 DVDD.n16420 0.0141679
R44862 DVDD.n16424 DVDD.n16423 0.0141679
R44863 DVDD.n16427 DVDD.n16426 0.0141679
R44864 DVDD.n16433 DVDD.n2264 0.0141679
R44865 DVDD.n16435 DVDD.n2263 0.0141679
R44866 DVDD.n16437 DVDD.n2262 0.0141679
R44867 DVDD.n16439 DVDD.n2261 0.0141679
R44868 DVDD.n16441 DVDD.n2260 0.0141679
R44869 DVDD.n16443 DVDD.n2259 0.0141679
R44870 DVDD.n16445 DVDD.n2258 0.0141679
R44871 DVDD.n16447 DVDD.n2257 0.0141679
R44872 DVDD.n5565 DVDD.n5561 0.0141679
R44873 DVDD.n5574 DVDD.n5573 0.0141679
R44874 DVDD.n5570 DVDD.n5569 0.0141679
R44875 DVDD.n10206 DVDD.n10205 0.0141679
R44876 DVDD.n10208 DVDD.n10207 0.0141679
R44877 DVDD.n10210 DVDD.n10209 0.0141679
R44878 DVDD.n10212 DVDD.n10211 0.0141679
R44879 DVDD.n10214 DVDD.n10213 0.0141679
R44880 DVDD.n10216 DVDD.n10215 0.0141679
R44881 DVDD.n10218 DVDD.n10217 0.0141679
R44882 DVDD.n16409 DVDD.n16407 0.0141679
R44883 DVDD.n16412 DVDD.n16410 0.0141679
R44884 DVDD.n16415 DVDD.n16413 0.0141679
R44885 DVDD.n16418 DVDD.n16416 0.0141679
R44886 DVDD.n16421 DVDD.n16419 0.0141679
R44887 DVDD.n16424 DVDD.n16422 0.0141679
R44888 DVDD.n16426 DVDD.n16425 0.0141679
R44889 DVDD.n16435 DVDD.n16434 0.0141679
R44890 DVDD.n16437 DVDD.n16436 0.0141679
R44891 DVDD.n16439 DVDD.n16438 0.0141679
R44892 DVDD.n16441 DVDD.n16440 0.0141679
R44893 DVDD.n16443 DVDD.n16442 0.0141679
R44894 DVDD.n16445 DVDD.n16444 0.0141679
R44895 DVDD.n16447 DVDD.n16446 0.0141679
R44896 DVDD.n10220 DVDD.n8961 0.0141679
R44897 DVDD.n16430 DVDD.n2278 0.0141679
R44898 DVDD.n16448 DVDD.n2266 0.0141679
R44899 DVDD.n15145 DVDD.n5567 0.0141679
R44900 DVDD.n887 DVDD.n882 0.0141679
R44901 DVDD.n889 DVDD.n885 0.0141679
R44902 DVDD.n17733 DVDD.n17732 0.0141679
R44903 DVDD.n883 DVDD.n882 0.0141679
R44904 DVDD.n17730 DVDD.n17729 0.0141679
R44905 DVDD.n888 DVDD.n881 0.0141679
R44906 DVDD.n18026 DVDD.n18024 0.0141679
R44907 DVDD.n18030 DVDD.n18029 0.0141679
R44908 DVDD.n18033 DVDD.n544 0.0141679
R44909 DVDD.n550 DVDD.n547 0.0141679
R44910 DVDD.n18024 DVDD.n548 0.0141679
R44911 DVDD.n18031 DVDD.n18030 0.0141679
R44912 DVDD.n18035 DVDD.n545 0.0141679
R44913 DVDD.n17736 DVDD.n17735 0.0141679
R44914 DVDD.n10177 DVDD.n10176 0.0141679
R44915 DVDD.n10180 DVDD.n10179 0.0141679
R44916 DVDD.n10183 DVDD.n10182 0.0141679
R44917 DVDD.n10186 DVDD.n10185 0.0141679
R44918 DVDD.n10189 DVDD.n10188 0.0141679
R44919 DVDD.n10192 DVDD.n10191 0.0141679
R44920 DVDD.n10195 DVDD.n10194 0.0141679
R44921 DVDD.n10198 DVDD.n10197 0.0141679
R44922 DVDD.n10180 DVDD.n10178 0.0141679
R44923 DVDD.n10183 DVDD.n10181 0.0141679
R44924 DVDD.n10186 DVDD.n10184 0.0141679
R44925 DVDD.n10189 DVDD.n10187 0.0141679
R44926 DVDD.n10192 DVDD.n10190 0.0141679
R44927 DVDD.n10195 DVDD.n10193 0.0141679
R44928 DVDD.n10197 DVDD.n10196 0.0141679
R44929 DVDD.n10201 DVDD.n8971 0.0141679
R44930 DVDD.n4981 DVDD.n4907 0.0141679
R44931 DVDD.n4919 DVDD.n4918 0.0141679
R44932 DVDD.n4922 DVDD.n4921 0.0141679
R44933 DVDD.n4925 DVDD.n4924 0.0141679
R44934 DVDD.n4928 DVDD.n4927 0.0141679
R44935 DVDD.n4931 DVDD.n4930 0.0141679
R44936 DVDD.n4934 DVDD.n4933 0.0141679
R44937 DVDD.n4937 DVDD.n4936 0.0141679
R44938 DVDD.n4940 DVDD.n4939 0.0141679
R44939 DVDD.n4919 DVDD.n4917 0.0141679
R44940 DVDD.n4922 DVDD.n4920 0.0141679
R44941 DVDD.n4925 DVDD.n4923 0.0141679
R44942 DVDD.n4928 DVDD.n4926 0.0141679
R44943 DVDD.n4931 DVDD.n4929 0.0141679
R44944 DVDD.n4934 DVDD.n4932 0.0141679
R44945 DVDD.n4937 DVDD.n4935 0.0141679
R44946 DVDD.n4940 DVDD.n4938 0.0141679
R44947 DVDD.n4979 DVDD.n4941 0.0141679
R44948 DVDD.n22236 DVDD.n22235 0.0141393
R44949 DVDD.n22235 DVDD.n132 0.0141393
R44950 DVDD.n22231 DVDD.n132 0.0141393
R44951 DVDD.n21724 DVDD.n21723 0.0141393
R44952 DVDD.n21729 DVDD.n21724 0.0141393
R44953 DVDD.n21729 DVDD.n18430 0.0141393
R44954 DVDD.n21927 DVDD.n21926 0.0141393
R44955 DVDD.n21926 DVDD.n21794 0.0141393
R44956 DVDD.n21922 DVDD.n21794 0.0141393
R44957 DVDD.n22040 DVDD.n18209 0.0141393
R44958 DVDD.n22065 DVDD.n18209 0.0141393
R44959 DVDD.n22065 DVDD.n18207 0.0141393
R44960 DVDD.n18390 DVDD.n18389 0.0141393
R44961 DVDD.n21775 DVDD.n18389 0.0141393
R44962 DVDD.n21775 DVDD.n180 0.0141393
R44963 DVDD.n21939 DVDD.n21782 0.0141393
R44964 DVDD.n21935 DVDD.n21782 0.0141393
R44965 DVDD.n18121 DVDD.n18120 0.0141393
R44966 DVDD.n18120 DVDD.n18066 0.0141393
R44967 DVDD.n18116 DVDD.n18066 0.0141393
R44968 DVDD.n18112 DVDD.n18098 0.0141393
R44969 DVDD.n18108 DVDD.n18098 0.0141393
R44970 DVDD.n18108 DVDD.n18100 0.0141393
R44971 DVDD.n14301 DVDD.n8260 0.014059
R44972 DVDD.n14300 DVDD.n8262 0.014059
R44973 DVDD.n14288 DVDD.n10238 0.0140338
R44974 DVDD.n17277 DVDD.n17276 0.0140338
R44975 DVDD.n17727 DVDD.n17726 0.0140338
R44976 DVDD.n6401 DVDD.n5999 0.0140302
R44977 DVDD.n8148 DVDD.n8147 0.0140302
R44978 DVDD.n6400 DVDD.n5998 0.0140302
R44979 DVDD.n14576 DVDD.n8134 0.0140302
R44980 DVDD.n13792 DVDD.n11565 0.013775
R44981 DVDD.n17266 DVDD.n1608 0.013775
R44982 DVDD.n779 DVDD.n777 0.0137065
R44983 DVDD.n17895 DVDD.n779 0.0137065
R44984 DVDD.n15308 DVDD.n15307 0.0137065
R44985 DVDD.n15307 DVDD.n15306 0.0137065
R44986 DVDD.n8253 DVDD.n8252 0.013547
R44987 DVDD.n14310 DVDD.n14309 0.013547
R44988 DVDD.n15075 DVDD.n15074 0.0134925
R44989 DVDD.n9566 DVDD.n9219 0.0134925
R44990 DVDD.n21683 DVDD.n21682 0.0134316
R44991 DVDD.n18366 DVDD.n18313 0.0134316
R44992 DVDD.n21221 DVDD.n18657 0.0134316
R44993 DVDD.n21368 DVDD.n21367 0.0134316
R44994 DVDD.n18341 DVDD.n18338 0.0134316
R44995 DVDD.n21995 DVDD.n21993 0.0134316
R44996 DVDD.n4846 DVDD.n3550 0.0134316
R44997 DVDD.n4874 DVDD.n3537 0.0134316
R44998 DVDD.n18401 DVDD.n18379 0.013325
R44999 DVDD.n21985 DVDD.n18247 0.013325
R45000 DVDD.n21353 DVDD.n140 0.013325
R45001 DVDD.n21703 DVDD.n18305 0.013325
R45002 DVDD.n18263 DVDD.n18229 0.013325
R45003 DVDD.n161 DVDD.n152 0.013325
R45004 DVDD.n4298 DVDD.n4283 0.013325
R45005 DVDD.n3693 DVDD.n3692 0.013325
R45006 DVDD.n11570 DVDD.n11058 0.013325
R45007 DVDD.n17268 DVDD.n1259 0.013325
R45008 DVDD.n21681 DVDD.n18536 0.0131188
R45009 DVDD.n21362 DVDD.n21333 0.0131188
R45010 DVDD.n22007 DVDD.n22006 0.0131188
R45011 DVDD.n3549 DVDD.n3547 0.0131188
R45012 DVDD.n13756 DVDD.n11934 0.0130638
R45013 DVDD.n12896 DVDD.n12781 0.0130638
R45014 DVDD.n13757 DVDD.n11932 0.0130638
R45015 DVDD.n12898 DVDD.n12897 0.0130638
R45016 DVDD.n11218 DVDD.n10706 0.0129511
R45017 DVDD.n16721 DVDD.n1801 0.0129511
R45018 DVDD.n18367 DVDD.n18311 0.0129102
R45019 DVDD.n21270 DVDD.n21269 0.0129102
R45020 DVDD.n18342 DVDD.n18337 0.0129102
R45021 DVDD.n4879 DVDD.n3532 0.0129102
R45022 DVDD.n7665 DVDD.n7407 0.012875
R45023 DVDD.n15120 DVDD.n5993 0.0128221
R45024 DVDD.n15119 DVDD.n5995 0.0128221
R45025 DVDD.n14286 DVDD.n10240 0.0125805
R45026 DVDD.n17279 DVDD.n1265 0.0125805
R45027 DVDD.n14287 DVDD.n10239 0.0125805
R45028 DVDD.n17278 DVDD.n1266 0.0125805
R45029 DVDD.n7668 DVDD.n7658 0.0124869
R45030 DVDD.n14857 DVDD.n7662 0.0124869
R45031 DVDD.n21770 DVDD.n18391 0.0124104
R45032 DVDD.n21933 DVDD.n21786 0.0124104
R45033 DVDD.n18481 DVDD.n131 0.0124104
R45034 DVDD.n21733 DVDD.n21732 0.0124104
R45035 DVDD.n21896 DVDD.n21793 0.0124104
R45036 DVDD.n22068 DVDD.n18206 0.0124104
R45037 DVDD.n18124 DVDD.n18123 0.0124104
R45038 DVDD.n18106 DVDD.n18105 0.0124104
R45039 DVDD.n13805 DVDD.n13804 0.0124098
R45040 DVDD.n16453 DVDD.n2254 0.0124098
R45041 DVDD.n903 DVDD.n894 0.0123125
R45042 DVDD.n17361 DVDD.n905 0.0123125
R45043 DVDD.n5995 DVDD.n5580 0.0123125
R45044 DVDD.n5993 DVDD.n5936 0.0123125
R45045 DVDD.n16402 DVDD.n779 0.01221
R45046 DVDD.n15307 DVDD.n2292 0.01221
R45047 DVDD.n21766 DVDD.n21764 0.0121222
R45048 DVDD.n21727 DVDD.n18429 0.0121222
R45049 DVDD.n22063 DVDD.n18211 0.0121222
R45050 DVDD.n18122 DVDD.n18065 0.0121222
R45051 DVDD.n15077 DVDD.n7059 0.0120973
R45052 DVDD.n9221 DVDD.n7613 0.0120973
R45053 DVDD.n15076 DVDD.n7061 0.0120973
R45054 DVDD.n9568 DVDD.n9567 0.0120973
R45055 DVDD.n11575 DVDD.n11277 0.0120939
R45056 DVDD.n17264 DVDD.n1610 0.0120939
R45057 DVDD.n11577 DVDD.n11576 0.0120939
R45058 DVDD.n17265 DVDD.n1609 0.0120939
R45059 DVDD.n18312 DVDD.n18308 0.0120759
R45060 DVDD.n18659 DVDD.n18658 0.0120759
R45061 DVDD.n18349 DVDD.n18333 0.0120759
R45062 DVDD.n4875 DVDD.n3536 0.0120759
R45063 DVDD.n17713 DVDD.n17305 0.011975
R45064 DVDD.n15128 DVDD.n15127 0.011975
R45065 DVDD.n21934 DVDD.n21784 0.0119301
R45066 DVDD.n22238 DVDD.n22237 0.0119301
R45067 DVDD.n21929 DVDD.n21928 0.0119301
R45068 DVDD.n18104 DVDD.n18103 0.0119301
R45069 DVDD.n15097 DVDD.n6702 0.0118684
R45070 DVDD.n14844 DVDD.n7685 0.0118684
R45071 DVDD.n22193 DVDD.n209 0.01175
R45072 DVDD.n21721 DVDD.n18503 0.01175
R45073 DVDD.n18290 DVDD.n196 0.01175
R45074 DVDD.n22193 DVDD.n216 0.01175
R45075 DVDD.n21847 DVDD.n196 0.01175
R45076 DVDD.n21721 DVDD.n18448 0.01175
R45077 DVDD.n4312 DVDD.n4281 0.01175
R45078 DVDD.n3697 DVDD.n3673 0.01175
R45079 DVDD.n11572 DVDD.n11060 0.0117009
R45080 DVDD.n17270 DVDD.n1261 0.0117009
R45081 DVDD.n11571 DVDD.n11059 0.0117009
R45082 DVDD.n17269 DVDD.n1260 0.0117009
R45083 DVDD.n20594 DVDD.n19712 0.01166
R45084 DVDD.n20588 DVDD.n19712 0.01166
R45085 DVDD.n20588 DVDD.n20587 0.01166
R45086 DVDD.n20587 DVDD.n20586 0.01166
R45087 DVDD.n20586 DVDD.n19716 0.01166
R45088 DVDD.n20580 DVDD.n19716 0.01166
R45089 DVDD.n20580 DVDD.n20579 0.01166
R45090 DVDD.n20579 DVDD.n20578 0.01166
R45091 DVDD.n20578 DVDD.n19720 0.01166
R45092 DVDD.n19752 DVDD.n19720 0.01166
R45093 DVDD.n19753 DVDD.n19752 0.01166
R45094 DVDD.n19754 DVDD.n19753 0.01166
R45095 DVDD.n20566 DVDD.n19754 0.01166
R45096 DVDD.n20566 DVDD.n20565 0.01166
R45097 DVDD.n20565 DVDD.n20563 0.01166
R45098 DVDD.n20563 DVDD.n19757 0.01166
R45099 DVDD.n20556 DVDD.n19757 0.01166
R45100 DVDD.n20556 DVDD.n20555 0.01166
R45101 DVDD.n20555 DVDD.n19759 0.01166
R45102 DVDD.n19763 DVDD.n19759 0.01166
R45103 DVDD.n20548 DVDD.n19763 0.01166
R45104 DVDD.n20548 DVDD.n20547 0.01166
R45105 DVDD.n20547 DVDD.n20546 0.01166
R45106 DVDD.n20546 DVDD.n19710 0.01166
R45107 DVDD.n20080 DVDD.n19711 0.01166
R45108 DVDD.n20084 DVDD.n20080 0.01166
R45109 DVDD.n20085 DVDD.n20084 0.01166
R45110 DVDD.n20086 DVDD.n20085 0.01166
R45111 DVDD.n20086 DVDD.n20078 0.01166
R45112 DVDD.n20090 DVDD.n20078 0.01166
R45113 DVDD.n20091 DVDD.n20090 0.01166
R45114 DVDD.n20120 DVDD.n20091 0.01166
R45115 DVDD.n20120 DVDD.n20119 0.01166
R45116 DVDD.n20119 DVDD.n20117 0.01166
R45117 DVDD.n20117 DVDD.n20115 0.01166
R45118 DVDD.n20115 DVDD.n20113 0.01166
R45119 DVDD.n20113 DVDD.n20111 0.01166
R45120 DVDD.n20111 DVDD.n20109 0.01166
R45121 DVDD.n20109 DVDD.n20107 0.01166
R45122 DVDD.n20107 DVDD.n20105 0.01166
R45123 DVDD.n20105 DVDD.n20103 0.01166
R45124 DVDD.n20103 DVDD.n20101 0.01166
R45125 DVDD.n20101 DVDD.n20092 0.01166
R45126 DVDD.n20097 DVDD.n20092 0.01166
R45127 DVDD.n20097 DVDD.n20096 0.01166
R45128 DVDD.n20096 DVDD.n20095 0.01166
R45129 DVDD.n20095 DVDD.n19709 0.01166
R45130 DVDD.n20595 DVDD.n19709 0.01166
R45131 DVDD.n20592 DVDD.n20591 0.01166
R45132 DVDD.n20591 DVDD.n20590 0.01166
R45133 DVDD.n20590 DVDD.n19714 0.01166
R45134 DVDD.n20584 DVDD.n19714 0.01166
R45135 DVDD.n20584 DVDD.n20583 0.01166
R45136 DVDD.n20583 DVDD.n20582 0.01166
R45137 DVDD.n20582 DVDD.n19718 0.01166
R45138 DVDD.n20576 DVDD.n19718 0.01166
R45139 DVDD.n20576 DVDD.n20575 0.01166
R45140 DVDD.n20575 DVDD.n19723 0.01166
R45141 DVDD.n19755 DVDD.n19723 0.01166
R45142 DVDD.n20569 DVDD.n19755 0.01166
R45143 DVDD.n20569 DVDD.n20568 0.01166
R45144 DVDD.n20568 DVDD.n19756 0.01166
R45145 DVDD.n20561 DVDD.n19756 0.01166
R45146 DVDD.n20561 DVDD.n20560 0.01166
R45147 DVDD.n20560 DVDD.n20558 0.01166
R45148 DVDD.n20558 DVDD.n19758 0.01166
R45149 DVDD.n20552 DVDD.n19758 0.01166
R45150 DVDD.n20552 DVDD.n20551 0.01166
R45151 DVDD.n20551 DVDD.n20550 0.01166
R45152 DVDD.n20550 DVDD.n19761 0.01166
R45153 DVDD.n20544 DVDD.n19761 0.01166
R45154 DVDD.n20544 DVDD.n20543 0.01166
R45155 DVDD.n19981 DVDD.n19980 0.01166
R45156 DVDD.n19985 DVDD.n19980 0.01166
R45157 DVDD.n19986 DVDD.n19985 0.01166
R45158 DVDD.n19987 DVDD.n19986 0.01166
R45159 DVDD.n19987 DVDD.n19978 0.01166
R45160 DVDD.n19991 DVDD.n19978 0.01166
R45161 DVDD.n19992 DVDD.n19991 0.01166
R45162 DVDD.n20021 DVDD.n19992 0.01166
R45163 DVDD.n20021 DVDD.n20020 0.01166
R45164 DVDD.n20020 DVDD.n20018 0.01166
R45165 DVDD.n20018 DVDD.n20016 0.01166
R45166 DVDD.n20016 DVDD.n20014 0.01166
R45167 DVDD.n20014 DVDD.n20012 0.01166
R45168 DVDD.n20012 DVDD.n20010 0.01166
R45169 DVDD.n20010 DVDD.n20008 0.01166
R45170 DVDD.n20008 DVDD.n20006 0.01166
R45171 DVDD.n20006 DVDD.n20004 0.01166
R45172 DVDD.n20004 DVDD.n20002 0.01166
R45173 DVDD.n20002 DVDD.n19993 0.01166
R45174 DVDD.n19998 DVDD.n19993 0.01166
R45175 DVDD.n19998 DVDD.n19997 0.01166
R45176 DVDD.n19997 DVDD.n19996 0.01166
R45177 DVDD.n19996 DVDD.n19765 0.01166
R45178 DVDD.n20542 DVDD.n19765 0.01166
R45179 DVDD.n20898 DVDD.n18924 0.01166
R45180 DVDD.n20894 DVDD.n18924 0.01166
R45181 DVDD.n20894 DVDD.n20893 0.01166
R45182 DVDD.n20893 DVDD.n20892 0.01166
R45183 DVDD.n20892 DVDD.n18926 0.01166
R45184 DVDD.n20888 DVDD.n18926 0.01166
R45185 DVDD.n20888 DVDD.n20887 0.01166
R45186 DVDD.n20887 DVDD.n20886 0.01166
R45187 DVDD.n20886 DVDD.n18928 0.01166
R45188 DVDD.n20880 DVDD.n18928 0.01166
R45189 DVDD.n20880 DVDD.n20879 0.01166
R45190 DVDD.n20879 DVDD.n20877 0.01166
R45191 DVDD.n20877 DVDD.n20875 0.01166
R45192 DVDD.n20875 DVDD.n20873 0.01166
R45193 DVDD.n20873 DVDD.n20871 0.01166
R45194 DVDD.n20871 DVDD.n20869 0.01166
R45195 DVDD.n20869 DVDD.n20867 0.01166
R45196 DVDD.n20867 DVDD.n20865 0.01166
R45197 DVDD.n20865 DVDD.n18957 0.01166
R45198 DVDD.n20861 DVDD.n18957 0.01166
R45199 DVDD.n20861 DVDD.n20860 0.01166
R45200 DVDD.n20860 DVDD.n20859 0.01166
R45201 DVDD.n20859 DVDD.n18959 0.01166
R45202 DVDD.n18959 DVDD.n18922 0.01166
R45203 DVDD.n20436 DVDD.n18923 0.01166
R45204 DVDD.n20436 DVDD.n20435 0.01166
R45205 DVDD.n20435 DVDD.n20434 0.01166
R45206 DVDD.n20434 DVDD.n19826 0.01166
R45207 DVDD.n20428 DVDD.n19826 0.01166
R45208 DVDD.n20428 DVDD.n20427 0.01166
R45209 DVDD.n20427 DVDD.n20426 0.01166
R45210 DVDD.n20426 DVDD.n19831 0.01166
R45211 DVDD.n20379 DVDD.n19831 0.01166
R45212 DVDD.n20417 DVDD.n20379 0.01166
R45213 DVDD.n20417 DVDD.n20416 0.01166
R45214 DVDD.n20416 DVDD.n20380 0.01166
R45215 DVDD.n20409 DVDD.n20380 0.01166
R45216 DVDD.n20409 DVDD.n20408 0.01166
R45217 DVDD.n20408 DVDD.n20406 0.01166
R45218 DVDD.n20406 DVDD.n20382 0.01166
R45219 DVDD.n20399 DVDD.n20382 0.01166
R45220 DVDD.n20399 DVDD.n20398 0.01166
R45221 DVDD.n20398 DVDD.n20384 0.01166
R45222 DVDD.n20389 DVDD.n20384 0.01166
R45223 DVDD.n20391 DVDD.n20389 0.01166
R45224 DVDD.n20391 DVDD.n20390 0.01166
R45225 DVDD.n20390 DVDD.n18921 0.01166
R45226 DVDD.n20899 DVDD.n18921 0.01166
R45227 DVDD.n20439 DVDD.n19824 0.01166
R45228 DVDD.n19828 DVDD.n19824 0.01166
R45229 DVDD.n20432 DVDD.n19828 0.01166
R45230 DVDD.n20432 DVDD.n20431 0.01166
R45231 DVDD.n20431 DVDD.n20430 0.01166
R45232 DVDD.n20430 DVDD.n19829 0.01166
R45233 DVDD.n20424 DVDD.n19829 0.01166
R45234 DVDD.n20424 DVDD.n20423 0.01166
R45235 DVDD.n20423 DVDD.n19833 0.01166
R45236 DVDD.n20378 DVDD.n19833 0.01166
R45237 DVDD.n20414 DVDD.n20378 0.01166
R45238 DVDD.n20414 DVDD.n20413 0.01166
R45239 DVDD.n20413 DVDD.n20411 0.01166
R45240 DVDD.n20411 DVDD.n20381 0.01166
R45241 DVDD.n20404 DVDD.n20381 0.01166
R45242 DVDD.n20404 DVDD.n20403 0.01166
R45243 DVDD.n20403 DVDD.n20401 0.01166
R45244 DVDD.n20401 DVDD.n20383 0.01166
R45245 DVDD.n20395 DVDD.n20383 0.01166
R45246 DVDD.n20395 DVDD.n20394 0.01166
R45247 DVDD.n20394 DVDD.n20393 0.01166
R45248 DVDD.n20393 DVDD.n20387 0.01166
R45249 DVDD.n20387 DVDD.n20386 0.01166
R45250 DVDD.n20386 DVDD.n18920 0.01166
R45251 DVDD.n19894 DVDD.n19823 0.01166
R45252 DVDD.n19898 DVDD.n19894 0.01166
R45253 DVDD.n19899 DVDD.n19898 0.01166
R45254 DVDD.n19900 DVDD.n19899 0.01166
R45255 DVDD.n19900 DVDD.n19892 0.01166
R45256 DVDD.n19904 DVDD.n19892 0.01166
R45257 DVDD.n19905 DVDD.n19904 0.01166
R45258 DVDD.n19934 DVDD.n19905 0.01166
R45259 DVDD.n19934 DVDD.n19933 0.01166
R45260 DVDD.n19933 DVDD.n19931 0.01166
R45261 DVDD.n19931 DVDD.n19929 0.01166
R45262 DVDD.n19929 DVDD.n19927 0.01166
R45263 DVDD.n19927 DVDD.n19925 0.01166
R45264 DVDD.n19925 DVDD.n19923 0.01166
R45265 DVDD.n19923 DVDD.n19921 0.01166
R45266 DVDD.n19921 DVDD.n19919 0.01166
R45267 DVDD.n19919 DVDD.n19917 0.01166
R45268 DVDD.n19917 DVDD.n19915 0.01166
R45269 DVDD.n19915 DVDD.n19906 0.01166
R45270 DVDD.n19911 DVDD.n19906 0.01166
R45271 DVDD.n19911 DVDD.n19910 0.01166
R45272 DVDD.n19910 DVDD.n19909 0.01166
R45273 DVDD.n19909 DVDD.n19822 0.01166
R45274 DVDD.n20440 DVDD.n19822 0.01166
R45275 DVDD.n11220 DVDD.n10709 0.0116141
R45276 DVDD.n16738 DVDD.n16737 0.0116141
R45277 DVDD.n11219 DVDD.n10707 0.0116141
R45278 DVDD.n16744 DVDD.n1802 0.0116141
R45279 DVDD.n21848 DVDD.n18380 0.011525
R45280 DVDD.n18268 DVDD.n18246 0.011525
R45281 DVDD.n18663 DVDD.n141 0.011525
R45282 DVDD.n18304 DVDD.n18291 0.011525
R45283 DVDD.n21801 DVDD.n18250 0.011525
R45284 DVDD.n18459 DVDD.n153 0.011525
R45285 DVDD.n4314 DVDD.n4299 0.011525
R45286 DVDD.n3708 DVDD.n3707 0.011525
R45287 DVDD.n6343 DVDD.n6342 0.011525
R45288 DVDD.n10226 DVDD.n10223 0.0114624
R45289 DVDD.n10227 DVDD.n8254 0.0113271
R45290 DVDD.n7667 DVDD.n7409 0.0113079
R45291 DVDD.n7666 DVDD.n7408 0.0113079
R45292 DVDD.n18538 DVDD.n18537 0.0112416
R45293 DVDD.n21363 DVDD.n21361 0.0112416
R45294 DVDD.n21999 DVDD.n21992 0.0112416
R45295 DVDD.n4851 DVDD.n4850 0.0112416
R45296 DVDD.n21785 DVDD.n21781 0.0111617
R45297 DVDD.n18479 DVDD.n133 0.0111617
R45298 DVDD.n21797 DVDD.n21795 0.0111617
R45299 DVDD.n18107 DVDD.n18102 0.0111617
R45300 DVDD.n18162 DVDD.n18161 0.0111596
R45301 DVDD.n13807 DVDD.n11226 0.0111309
R45302 DVDD.n12909 DVDD.n1820 0.0111309
R45303 DVDD.n13806 DVDD.n11228 0.0111309
R45304 DVDD.n16455 DVDD.n16454 0.0111309
R45305 DVDD.n14297 DVDD.n8606 0.011075
R45306 DVDD.n13493 DVDD.n12377 0.0107857
R45307 DVDD.n13491 DVDD.n12384 0.0107857
R45308 DVDD.n15099 DVDD.n6392 0.0106477
R45309 DVDD.n14842 DVDD.n7687 0.0106477
R45310 DVDD.n15098 DVDD.n6394 0.0106477
R45311 DVDD.n14843 DVDD.n7686 0.0106477
R45312 DVDD.n13479 DVDD.n12731 0.010625
R45313 DVDD.n13262 DVDD.n13261 0.010625
R45314 DVDD.n6751 DVDD.n6704 0.0105588
R45315 DVDD.n15087 DVDD.n15086 0.0105588
R45316 DVDD.n15090 DVDD.n6705 0.0105588
R45317 DVDD.n15088 DVDD.n6795 0.0105588
R45318 DVDD.n7153 DVDD.n7061 0.0105588
R45319 DVDD.n7112 DVDD.n7053 0.0105588
R45320 DVDD.n7111 DVDD.n7059 0.0105588
R45321 DVDD.n7403 DVDD.n7055 0.0105588
R45322 DVDD.n14868 DVDD.n7457 0.0105588
R45323 DVDD.n15055 DVDD.n7408 0.0105588
R45324 DVDD.n15058 DVDD.n7456 0.0105588
R45325 DVDD.n15056 DVDD.n7409 0.0105588
R45326 DVDD.n9568 DVDD.n7614 0.0105588
R45327 DVDD.n14858 DVDD.n14857 0.0105588
R45328 DVDD.n14861 DVDD.n7613 0.0105588
R45329 DVDD.n14859 DVDD.n7658 0.0105588
R45330 DVDD.n9555 DVDD.n7682 0.0105588
R45331 DVDD.n9310 DVDD.n7675 0.0105588
R45332 DVDD.n9556 DVDD.n7680 0.0105588
R45333 DVDD.n9309 DVDD.n7677 0.0105588
R45334 DVDD.n7732 DVDD.n7686 0.0105588
R45335 DVDD.n14835 DVDD.n14834 0.0105588
R45336 DVDD.n14838 DVDD.n7687 0.0105588
R45337 DVDD.n14836 DVDD.n7776 0.0105588
R45338 DVDD.n14577 DVDD.n14576 0.0105588
R45339 DVDD.n8088 DVDD.n8040 0.0105588
R45340 DVDD.n8148 DVDD.n8086 0.0105588
R45341 DVDD.n14824 DVDD.n8042 0.0105588
R45342 DVDD.n14311 DVDD.n14310 0.0105588
R45343 DVDD.n8206 DVDD.n8157 0.0105588
R45344 DVDD.n8252 DVDD.n8204 0.0105588
R45345 DVDD.n14558 DVDD.n8156 0.0105588
R45346 DVDD.n8348 DVDD.n8255 0.0105588
R45347 DVDD.n8597 DVDD.n8262 0.0105588
R45348 DVDD.n8349 DVDD.n8257 0.0105588
R45349 DVDD.n8596 DVDD.n8260 0.0105588
R45350 DVDD.n8948 DVDD.n8613 0.0105588
R45351 DVDD.n8739 DVDD.n8607 0.0105588
R45352 DVDD.n8947 DVDD.n8611 0.0105588
R45353 DVDD.n8738 DVDD.n8608 0.0105588
R45354 DVDD.n10285 DVDD.n10239 0.0105588
R45355 DVDD.n14279 DVDD.n14278 0.0105588
R45356 DVDD.n14282 DVDD.n10240 0.0105588
R45357 DVDD.n14280 DVDD.n10329 0.0105588
R45358 DVDD.n14021 DVDD.n14020 0.0105588
R45359 DVDD.n10641 DVDD.n10593 0.0105588
R45360 DVDD.n10704 DVDD.n10639 0.0105588
R45361 DVDD.n14268 DVDD.n10595 0.0105588
R45362 DVDD.n10800 DVDD.n10707 0.0105588
R45363 DVDD.n11049 DVDD.n10714 0.0105588
R45364 DVDD.n10801 DVDD.n10709 0.0105588
R45365 DVDD.n11048 DVDD.n10712 0.0105588
R45366 DVDD.n11224 DVDD.n11106 0.0105588
R45367 DVDD.n13998 DVDD.n11059 0.0105588
R45368 DVDD.n14001 DVDD.n11105 0.0105588
R45369 DVDD.n13999 DVDD.n11060 0.0105588
R45370 DVDD.n11320 DVDD.n11228 0.0105588
R45371 DVDD.n11577 DVDD.n11278 0.0105588
R45372 DVDD.n11275 DVDD.n11226 0.0105588
R45373 DVDD.n13798 DVDD.n11277 0.0105588
R45374 DVDD.n11674 DVDD.n11583 0.0105588
R45375 DVDD.n11922 DVDD.n11633 0.0105588
R45376 DVDD.n11630 DVDD.n11582 0.0105588
R45377 DVDD.n13776 DVDD.n11632 0.0105588
R45378 DVDD.n12027 DVDD.n11932 0.0105588
R45379 DVDD.n12276 DVDD.n11942 0.0105588
R45380 DVDD.n12028 DVDD.n11934 0.0105588
R45381 DVDD.n12275 DVDD.n11940 0.0105588
R45382 DVDD.n13496 DVDD.n13495 0.0105588
R45383 DVDD.n12331 DVDD.n12283 0.0105588
R45384 DVDD.n12382 DVDD.n12329 0.0105588
R45385 DVDD.n13743 DVDD.n12285 0.0105588
R45386 DVDD.n12434 DVDD.n12385 0.0105588
R45387 DVDD.n13482 DVDD.n13481 0.0105588
R45388 DVDD.n13485 DVDD.n12387 0.0105588
R45389 DVDD.n13483 DVDD.n12478 0.0105588
R45390 DVDD.n12898 DVDD.n12782 0.0105588
R45391 DVDD.n13468 DVDD.n12733 0.0105588
R45392 DVDD.n13471 DVDD.n12781 0.0105588
R45393 DVDD.n13469 DVDD.n12735 0.0105588
R45394 DVDD.n13253 DVDD.n12906 0.0105588
R45395 DVDD.n13008 DVDD.n12914 0.0105588
R45396 DVDD.n13254 DVDD.n12908 0.0105588
R45397 DVDD.n13007 DVDD.n12913 0.0105588
R45398 DVDD.n16456 DVDD.n16455 0.0105588
R45399 DVDD.n2209 DVDD.n2162 0.0105588
R45400 DVDD.n12909 DVDD.n2207 0.0105588
R45401 DVDD.n16703 DVDD.n2164 0.0105588
R45402 DVDD.n2153 DVDD.n1815 0.0105588
R45403 DVDD.n1908 DVDD.n1809 0.0105588
R45404 DVDD.n2154 DVDD.n1814 0.0105588
R45405 DVDD.n1907 DVDD.n1810 0.0105588
R45406 DVDD.n16745 DVDD.n16744 0.0105588
R45407 DVDD.n1756 DVDD.n1710 0.0105588
R45408 DVDD.n16738 DVDD.n1754 0.0105588
R45409 DVDD.n16993 DVDD.n1711 0.0105588
R45410 DVDD.n17013 DVDD.n17012 0.0105588
R45411 DVDD.n1657 DVDD.n1609 0.0105588
R45412 DVDD.n17006 DVDD.n1653 0.0105588
R45413 DVDD.n17261 DVDD.n1610 0.0105588
R45414 DVDD.n1603 DVDD.n1265 0.0105588
R45415 DVDD.n1356 DVDD.n1261 0.0105588
R45416 DVDD.n6508 DVDD.n6394 0.0105588
R45417 DVDD.n6694 DVDD.n6345 0.0105588
R45418 DVDD.n6404 DVDD.n6392 0.0105588
R45419 DVDD.n6695 DVDD.n6347 0.0105588
R45420 DVDD.n963 DVDD.n916 0.0105588
R45421 DVDD.n1068 DVDD.n914 0.0105588
R45422 DVDD.n6042 DVDD.n5999 0.0105588
R45423 DVDD.n15111 DVDD.n6044 0.0105588
R45424 DVDD.n6091 DVDD.n5998 0.0105588
R45425 DVDD.n15110 DVDD.n15109 0.0105588
R45426 DVDD.n1602 DVDD.n1266 0.0105588
R45427 DVDD.n1357 DVDD.n1260 0.0105588
R45428 DVDD.n965 DVDD.n917 0.0105588
R45429 DVDD.n1069 DVDD.n913 0.0105588
R45430 DVDD.n22193 DVDD.n220 0.01055
R45431 DVDD.n21721 DVDD.n18506 0.01055
R45432 DVDD.n21699 DVDD.n196 0.01055
R45433 DVDD.n22193 DVDD.n212 0.01055
R45434 DVDD.n18416 DVDD.n196 0.01055
R45435 DVDD.n21721 DVDD.n18447 0.01055
R45436 DVDD.n4296 DVDD.n4281 0.01055
R45437 DVDD.n3688 DVDD.n3673 0.01055
R45438 DVDD.n172 DVDD.n171 0.0104
R45439 DVDD.n18514 DVDD.n18513 0.0104
R45440 DVDD.n18544 DVDD.n18531 0.0104
R45441 DVDD.n21661 DVDD.n21660 0.0104
R45442 DVDD.n21713 DVDD.n21712 0.0104
R45443 DVDD.n22217 DVDD.n22216 0.0104
R45444 DVDD.n21741 DVDD.n18405 0.0104
R45445 DVDD.n21740 DVDD.n21739 0.0104
R45446 DVDD.n21765 DVDD.n18388 0.0103933
R45447 DVDD.n21728 DVDD.n21726 0.0103933
R45448 DVDD.n22064 DVDD.n18210 0.0103933
R45449 DVDD.n18093 DVDD.n18067 0.0103933
R45450 DVDD.n16453 DVDD.n16452 0.0103797
R45451 DVDD.n21678 DVDD.n21677 0.0103725
R45452 DVDD.n21677 DVDD.n21676 0.0103725
R45453 DVDD.n18371 DVDD.n18310 0.0103725
R45454 DVDD.n18371 DVDD.n18370 0.0103725
R45455 DVDD.n18346 DVDD.n18345 0.0103725
R45456 DVDD.n18346 DVDD.n207 0.0103725
R45457 DVDD.n22002 DVDD.n208 0.0103725
R45458 DVDD.n22003 DVDD.n22002 0.0103725
R45459 DVDD.n21266 DVDD.n21265 0.0103725
R45460 DVDD.n21265 DVDD.n18433 0.0103725
R45461 DVDD.n21335 DVDD.n18434 0.0103725
R45462 DVDD.n21365 DVDD.n21335 0.0103725
R45463 DVDD.n4848 DVDD.n3543 0.0103725
R45464 DVDD.n4860 DVDD.n3543 0.0103725
R45465 DVDD.n4862 DVDD.n3534 0.0103725
R45466 DVDD.n4877 DVDD.n3534 0.0103725
R45467 DVDD.n10237 DVDD.n10236 0.0102444
R45468 DVDD.n17295 DVDD.n17294 0.0102444
R45469 DVDD.n18374 DVDD.n18373 0.0101987
R45470 DVDD.n21262 DVDD.n21261 0.0101987
R45471 DVDD.n18348 DVDD.n18334 0.0101987
R45472 DVDD.n4866 DVDD.n4865 0.0101987
R45473 DVDD.n14564 DVDD.n14563 0.010175
R45474 DVDD.n17714 DVDD.n17713 0.010175
R45475 DVDD.n10229 DVDD.n8257 0.0101644
R45476 DVDD.n10228 DVDD.n8255 0.0101644
R45477 DVDD.n6338 DVDD.n6044 0.0101288
R45478 DVDD.n15109 DVDD.n6339 0.0101288
R45479 DVDD.n21888 DVDD.n21887 0.00992
R45480 DVDD.n18282 DVDD.n200 0.00992
R45481 DVDD.n18362 DVDD.n18317 0.00992
R45482 DVDD.n18361 DVDD.n18319 0.00992
R45483 DVDD.n22202 DVDD.n201 0.00992
R45484 DVDD.n21889 DVDD.n21886 0.00992
R45485 DVDD.n21904 DVDD.n21807 0.00992
R45486 DVDD.n21903 DVDD.n21808 0.00992
R45487 DVDD.n14295 DVDD.n8608 0.00973581
R45488 DVDD.n14296 DVDD.n8607 0.00973581
R45489 DVDD.n15095 DVDD.n6703 0.00970301
R45490 DVDD.n14846 DVDD.n7684 0.00970301
R45491 DVDD.n12383 DVDD.n12382 0.00968121
R45492 DVDD.n13489 DVDD.n12387 0.00968121
R45493 DVDD.n13495 DVDD.n13494 0.00968121
R45494 DVDD.n13490 DVDD.n12385 0.00968121
R45495 DVDD.n20139 DVDD.n20137 0.00962857
R45496 DVDD.n20144 DVDD.n20137 0.00962857
R45497 DVDD.n20146 DVDD.n20144 0.00962857
R45498 DVDD.n20148 DVDD.n20146 0.00962857
R45499 DVDD.n20148 DVDD.n20134 0.00962857
R45500 DVDD.n20153 DVDD.n20134 0.00962857
R45501 DVDD.n20155 DVDD.n20153 0.00962857
R45502 DVDD.n20157 DVDD.n20155 0.00962857
R45503 DVDD.n20157 DVDD.n20131 0.00962857
R45504 DVDD.n20161 DVDD.n20131 0.00962857
R45505 DVDD.n20161 DVDD.n20058 0.00962857
R45506 DVDD.n20167 DVDD.n20058 0.00962857
R45507 DVDD.n20167 DVDD.n20056 0.00962857
R45508 DVDD.n20172 DVDD.n20056 0.00962857
R45509 DVDD.n20172 DVDD.n20054 0.00962857
R45510 DVDD.n20176 DVDD.n20054 0.00962857
R45511 DVDD.n20178 DVDD.n20176 0.00962857
R45512 DVDD.n20178 DVDD.n20052 0.00962857
R45513 DVDD.n20183 DVDD.n20052 0.00962857
R45514 DVDD.n20185 DVDD.n20183 0.00962857
R45515 DVDD.n20187 DVDD.n20185 0.00962857
R45516 DVDD.n20187 DVDD.n20049 0.00962857
R45517 DVDD.n20192 DVDD.n20049 0.00962857
R45518 DVDD.n20194 DVDD.n20192 0.00962857
R45519 DVDD.n20196 DVDD.n20194 0.00962857
R45520 DVDD.n20196 DVDD.n20046 0.00962857
R45521 DVDD.n20201 DVDD.n20046 0.00962857
R45522 DVDD.n20203 DVDD.n20201 0.00962857
R45523 DVDD.n20204 DVDD.n20203 0.00962857
R45524 DVDD.n20204 DVDD.n20043 0.00962857
R45525 DVDD.n20209 DVDD.n20043 0.00962857
R45526 DVDD.n20209 DVDD.n20041 0.00962857
R45527 DVDD.n20213 DVDD.n20041 0.00962857
R45528 DVDD.n20215 DVDD.n20213 0.00962857
R45529 DVDD.n20217 DVDD.n20215 0.00962857
R45530 DVDD.n20217 DVDD.n20039 0.00962857
R45531 DVDD.n20222 DVDD.n20039 0.00962857
R45532 DVDD.n20224 DVDD.n20222 0.00962857
R45533 DVDD.n20226 DVDD.n20224 0.00962857
R45534 DVDD.n20226 DVDD.n20036 0.00962857
R45535 DVDD.n20231 DVDD.n20036 0.00962857
R45536 DVDD.n20233 DVDD.n20231 0.00962857
R45537 DVDD.n20235 DVDD.n20233 0.00962857
R45538 DVDD.n20235 DVDD.n20032 0.00962857
R45539 DVDD.n20240 DVDD.n20032 0.00962857
R45540 DVDD.n20240 DVDD.n20033 0.00962857
R45541 DVDD.n20033 DVDD.n19957 0.00962857
R45542 DVDD.n20247 DVDD.n19957 0.00962857
R45543 DVDD.n20247 DVDD.n19955 0.00962857
R45544 DVDD.n20252 DVDD.n19955 0.00962857
R45545 DVDD.n20252 DVDD.n19953 0.00962857
R45546 DVDD.n20256 DVDD.n19953 0.00962857
R45547 DVDD.n20258 DVDD.n20256 0.00962857
R45548 DVDD.n20258 DVDD.n19951 0.00962857
R45549 DVDD.n20263 DVDD.n19951 0.00962857
R45550 DVDD.n20265 DVDD.n20263 0.00962857
R45551 DVDD.n20267 DVDD.n20265 0.00962857
R45552 DVDD.n20267 DVDD.n19948 0.00962857
R45553 DVDD.n20272 DVDD.n19948 0.00962857
R45554 DVDD.n20274 DVDD.n20272 0.00962857
R45555 DVDD.n20276 DVDD.n20274 0.00962857
R45556 DVDD.n20276 DVDD.n19945 0.00962857
R45557 DVDD.n20280 DVDD.n19945 0.00962857
R45558 DVDD.n20280 DVDD.n19872 0.00962857
R45559 DVDD.n20287 DVDD.n19872 0.00962857
R45560 DVDD.n20287 DVDD.n19870 0.00962857
R45561 DVDD.n20291 DVDD.n19870 0.00962857
R45562 DVDD.n20291 DVDD.n19868 0.00962857
R45563 DVDD.n20295 DVDD.n19868 0.00962857
R45564 DVDD.n20295 DVDD.n19866 0.00962857
R45565 DVDD.n20300 DVDD.n19866 0.00962857
R45566 DVDD.n20302 DVDD.n20300 0.00962857
R45567 DVDD.n20304 DVDD.n20302 0.00962857
R45568 DVDD.n20304 DVDD.n19863 0.00962857
R45569 DVDD.n20309 DVDD.n19863 0.00962857
R45570 DVDD.n20311 DVDD.n20309 0.00962857
R45571 DVDD.n20313 DVDD.n20311 0.00962857
R45572 DVDD.n20313 DVDD.n19860 0.00962857
R45573 DVDD.n20318 DVDD.n19860 0.00962857
R45574 DVDD.n20320 DVDD.n20318 0.00962857
R45575 DVDD.n20322 DVDD.n20320 0.00962857
R45576 DVDD.n20322 DVDD.n19856 0.00962857
R45577 DVDD.n20370 DVDD.n19856 0.00962857
R45578 DVDD.n20370 DVDD.n19857 0.00962857
R45579 DVDD.n20366 DVDD.n19857 0.00962857
R45580 DVDD.n20366 DVDD.n20326 0.00962857
R45581 DVDD.n20362 DVDD.n20326 0.00962857
R45582 DVDD.n20362 DVDD.n20328 0.00962857
R45583 DVDD.n20358 DVDD.n20328 0.00962857
R45584 DVDD.n20358 DVDD.n20356 0.00962857
R45585 DVDD.n20356 DVDD.n20354 0.00962857
R45586 DVDD.n20354 DVDD.n20331 0.00962857
R45587 DVDD.n20349 DVDD.n20331 0.00962857
R45588 DVDD.n20349 DVDD.n20347 0.00962857
R45589 DVDD.n20347 DVDD.n20345 0.00962857
R45590 DVDD.n20345 DVDD.n20334 0.00962857
R45591 DVDD.n20340 DVDD.n20338 0.00962857
R45592 DVDD.n20338 DVDD.n20335 0.00962857
R45593 DVDD.n20166 DVDD.n20055 0.00962857
R45594 DVDD.n20173 DVDD.n20055 0.00962857
R45595 DVDD.n20174 DVDD.n20173 0.00962857
R45596 DVDD.n20175 DVDD.n20174 0.00962857
R45597 DVDD.n20210 DVDD.n19745 0.00962857
R45598 DVDD.n20211 DVDD.n20210 0.00962857
R45599 DVDD.n20212 DVDD.n20211 0.00962857
R45600 DVDD.n20246 DVDD.n20245 0.00962857
R45601 DVDD.n20246 DVDD.n19954 0.00962857
R45602 DVDD.n20253 DVDD.n19954 0.00962857
R45603 DVDD.n20254 DVDD.n20253 0.00962857
R45604 DVDD.n20255 DVDD.n20254 0.00962857
R45605 DVDD.n20292 DVDD.n19869 0.00962857
R45606 DVDD.n20293 DVDD.n20292 0.00962857
R45607 DVDD.n20294 DVDD.n20293 0.00962857
R45608 DVDD.n20371 DVDD.n19855 0.00962857
R45609 DVDD.n20365 DVDD.n19855 0.00962857
R45610 DVDD.n20365 DVDD.n20364 0.00962857
R45611 DVDD.n20364 DVDD.n20363 0.00962857
R45612 DVDD.n20626 DVDD.n20624 0.00962857
R45613 DVDD.n20631 DVDD.n20624 0.00962857
R45614 DVDD.n20633 DVDD.n20631 0.00962857
R45615 DVDD.n20635 DVDD.n20633 0.00962857
R45616 DVDD.n20635 DVDD.n20621 0.00962857
R45617 DVDD.n20640 DVDD.n20621 0.00962857
R45618 DVDD.n20642 DVDD.n20640 0.00962857
R45619 DVDD.n20649 DVDD.n20642 0.00962857
R45620 DVDD.n20649 DVDD.n20618 0.00962857
R45621 DVDD.n20653 DVDD.n20618 0.00962857
R45622 DVDD.n20653 DVDD.n19180 0.00962857
R45623 DVDD.n20659 DVDD.n19180 0.00962857
R45624 DVDD.n20659 DVDD.n19178 0.00962857
R45625 DVDD.n20664 DVDD.n19178 0.00962857
R45626 DVDD.n20664 DVDD.n19176 0.00962857
R45627 DVDD.n20668 DVDD.n19176 0.00962857
R45628 DVDD.n20670 DVDD.n20668 0.00962857
R45629 DVDD.n20670 DVDD.n19174 0.00962857
R45630 DVDD.n20675 DVDD.n19174 0.00962857
R45631 DVDD.n20677 DVDD.n20675 0.00962857
R45632 DVDD.n20679 DVDD.n20677 0.00962857
R45633 DVDD.n20679 DVDD.n19171 0.00962857
R45634 DVDD.n20684 DVDD.n19171 0.00962857
R45635 DVDD.n20686 DVDD.n20684 0.00962857
R45636 DVDD.n20688 DVDD.n20686 0.00962857
R45637 DVDD.n20688 DVDD.n19168 0.00962857
R45638 DVDD.n20693 DVDD.n19168 0.00962857
R45639 DVDD.n20695 DVDD.n20693 0.00962857
R45640 DVDD.n20696 DVDD.n20695 0.00962857
R45641 DVDD.n20696 DVDD.n19165 0.00962857
R45642 DVDD.n20701 DVDD.n19165 0.00962857
R45643 DVDD.n20701 DVDD.n19163 0.00962857
R45644 DVDD.n20705 DVDD.n19163 0.00962857
R45645 DVDD.n20707 DVDD.n20705 0.00962857
R45646 DVDD.n20709 DVDD.n20707 0.00962857
R45647 DVDD.n20709 DVDD.n19161 0.00962857
R45648 DVDD.n20714 DVDD.n19161 0.00962857
R45649 DVDD.n20716 DVDD.n20714 0.00962857
R45650 DVDD.n20718 DVDD.n20716 0.00962857
R45651 DVDD.n20718 DVDD.n19158 0.00962857
R45652 DVDD.n20723 DVDD.n19158 0.00962857
R45653 DVDD.n20725 DVDD.n20723 0.00962857
R45654 DVDD.n20727 DVDD.n20725 0.00962857
R45655 DVDD.n20727 DVDD.n19154 0.00962857
R45656 DVDD.n20732 DVDD.n19154 0.00962857
R45657 DVDD.n20732 DVDD.n19155 0.00962857
R45658 DVDD.n19155 DVDD.n19072 0.00962857
R45659 DVDD.n20739 DVDD.n19072 0.00962857
R45660 DVDD.n20739 DVDD.n19070 0.00962857
R45661 DVDD.n20744 DVDD.n19070 0.00962857
R45662 DVDD.n20744 DVDD.n19067 0.00962857
R45663 DVDD.n20748 DVDD.n19067 0.00962857
R45664 DVDD.n20750 DVDD.n20748 0.00962857
R45665 DVDD.n20752 DVDD.n20750 0.00962857
R45666 DVDD.n20752 DVDD.n19065 0.00962857
R45667 DVDD.n20757 DVDD.n19065 0.00962857
R45668 DVDD.n20759 DVDD.n20757 0.00962857
R45669 DVDD.n20761 DVDD.n20759 0.00962857
R45670 DVDD.n20761 DVDD.n19062 0.00962857
R45671 DVDD.n20766 DVDD.n19062 0.00962857
R45672 DVDD.n20768 DVDD.n20766 0.00962857
R45673 DVDD.n20770 DVDD.n20768 0.00962857
R45674 DVDD.n20770 DVDD.n19058 0.00962857
R45675 DVDD.n20775 DVDD.n19058 0.00962857
R45676 DVDD.n20775 DVDD.n19059 0.00962857
R45677 DVDD.n19059 DVDD.n19021 0.00962857
R45678 DVDD.n20783 DVDD.n19021 0.00962857
R45679 DVDD.n20783 DVDD.n19019 0.00962857
R45680 DVDD.n20787 DVDD.n19019 0.00962857
R45681 DVDD.n20788 DVDD.n20787 0.00962857
R45682 DVDD.n20790 DVDD.n20788 0.00962857
R45683 DVDD.n20790 DVDD.n19017 0.00962857
R45684 DVDD.n20795 DVDD.n19017 0.00962857
R45685 DVDD.n20797 DVDD.n20795 0.00962857
R45686 DVDD.n20799 DVDD.n20797 0.00962857
R45687 DVDD.n20799 DVDD.n19014 0.00962857
R45688 DVDD.n20804 DVDD.n19014 0.00962857
R45689 DVDD.n20806 DVDD.n20804 0.00962857
R45690 DVDD.n20808 DVDD.n20806 0.00962857
R45691 DVDD.n20808 DVDD.n19011 0.00962857
R45692 DVDD.n20813 DVDD.n19011 0.00962857
R45693 DVDD.n20815 DVDD.n20813 0.00962857
R45694 DVDD.n20817 DVDD.n20815 0.00962857
R45695 DVDD.n20817 DVDD.n19008 0.00962857
R45696 DVDD.n20822 DVDD.n19008 0.00962857
R45697 DVDD.n20822 DVDD.n19006 0.00962857
R45698 DVDD.n20826 DVDD.n19006 0.00962857
R45699 DVDD.n20828 DVDD.n20826 0.00962857
R45700 DVDD.n20828 DVDD.n19004 0.00962857
R45701 DVDD.n20833 DVDD.n19004 0.00962857
R45702 DVDD.n20835 DVDD.n20833 0.00962857
R45703 DVDD.n20837 DVDD.n20835 0.00962857
R45704 DVDD.n20837 DVDD.n19001 0.00962857
R45705 DVDD.n20842 DVDD.n19001 0.00962857
R45706 DVDD.n20844 DVDD.n20842 0.00962857
R45707 DVDD.n20846 DVDD.n20844 0.00962857
R45708 DVDD.n20850 DVDD.n18997 0.00962857
R45709 DVDD.n20850 DVDD.n18998 0.00962857
R45710 DVDD.n20658 DVDD.n19177 0.00962857
R45711 DVDD.n20665 DVDD.n19177 0.00962857
R45712 DVDD.n20666 DVDD.n20665 0.00962857
R45713 DVDD.n20667 DVDD.n20666 0.00962857
R45714 DVDD.n20702 DVDD.n18853 0.00962857
R45715 DVDD.n20703 DVDD.n20702 0.00962857
R45716 DVDD.n20704 DVDD.n20703 0.00962857
R45717 DVDD.n20738 DVDD.n20737 0.00962857
R45718 DVDD.n20738 DVDD.n19069 0.00962857
R45719 DVDD.n20745 DVDD.n19069 0.00962857
R45720 DVDD.n20746 DVDD.n20745 0.00962857
R45721 DVDD.n20747 DVDD.n20746 0.00962857
R45722 DVDD.n20782 DVDD.n20780 0.00962857
R45723 DVDD.n20782 DVDD.n20781 0.00962857
R45724 DVDD.n20781 DVDD.n18887 0.00962857
R45725 DVDD.n20816 DVDD.n19007 0.00962857
R45726 DVDD.n20823 DVDD.n19007 0.00962857
R45727 DVDD.n20824 DVDD.n20823 0.00962857
R45728 DVDD.n20825 DVDD.n20824 0.00962857
R45729 DVDD.n3974 DVDD.n3973 0.00962857
R45730 DVDD.n3973 DVDD.n3941 0.00962857
R45731 DVDD.n3961 DVDD.n3941 0.00962857
R45732 DVDD.n3961 DVDD.n3959 0.00962857
R45733 DVDD.n3959 DVDD.n3957 0.00962857
R45734 DVDD.n3957 DVDD.n3944 0.00962857
R45735 DVDD.n3952 DVDD.n3944 0.00962857
R45736 DVDD.n3952 DVDD.n3950 0.00962857
R45737 DVDD.n3950 DVDD.n3948 0.00962857
R45738 DVDD.n3948 DVDD.n3909 0.00962857
R45739 DVDD.n3980 DVDD.n3909 0.00962857
R45740 DVDD.n3980 DVDD.n3907 0.00962857
R45741 DVDD.n3984 DVDD.n3907 0.00962857
R45742 DVDD.n3984 DVDD.n3905 0.00962857
R45743 DVDD.n3989 DVDD.n3905 0.00962857
R45744 DVDD.n3989 DVDD.n3903 0.00962857
R45745 DVDD.n3994 DVDD.n3903 0.00962857
R45746 DVDD.n3996 DVDD.n3994 0.00962857
R45747 DVDD.n3998 DVDD.n3996 0.00962857
R45748 DVDD.n3998 DVDD.n3899 0.00962857
R45749 DVDD.n4061 DVDD.n3899 0.00962857
R45750 DVDD.n4061 DVDD.n3901 0.00962857
R45751 DVDD.n4057 DVDD.n3901 0.00962857
R45752 DVDD.n4057 DVDD.n4055 0.00962857
R45753 DVDD.n4055 DVDD.n4053 0.00962857
R45754 DVDD.n4053 DVDD.n4003 0.00962857
R45755 DVDD.n4048 DVDD.n4003 0.00962857
R45756 DVDD.n4048 DVDD.n4046 0.00962857
R45757 DVDD.n4046 DVDD.n4044 0.00962857
R45758 DVDD.n4044 DVDD.n4005 0.00962857
R45759 DVDD.n4040 DVDD.n4005 0.00962857
R45760 DVDD.n4040 DVDD.n4007 0.00962857
R45761 DVDD.n4036 DVDD.n4007 0.00962857
R45762 DVDD.n4036 DVDD.n4009 0.00962857
R45763 DVDD.n4032 DVDD.n4009 0.00962857
R45764 DVDD.n4032 DVDD.n4030 0.00962857
R45765 DVDD.n4030 DVDD.n4028 0.00962857
R45766 DVDD.n4028 DVDD.n4012 0.00962857
R45767 DVDD.n4023 DVDD.n4012 0.00962857
R45768 DVDD.n4023 DVDD.n4021 0.00962857
R45769 DVDD.n4021 DVDD.n4019 0.00962857
R45770 DVDD.n4019 DVDD.n4015 0.00962857
R45771 DVDD.n4015 DVDD.n273 0.00962857
R45772 DVDD.n22176 DVDD.n273 0.00962857
R45773 DVDD.n22176 DVDD.n275 0.00962857
R45774 DVDD.n22172 DVDD.n275 0.00962857
R45775 DVDD.n22172 DVDD.n22171 0.00962857
R45776 DVDD.n22171 DVDD.n22170 0.00962857
R45777 DVDD.n22170 DVDD.n278 0.00962857
R45778 DVDD.n22166 DVDD.n278 0.00962857
R45779 DVDD.n22166 DVDD.n281 0.00962857
R45780 DVDD.n22162 DVDD.n281 0.00962857
R45781 DVDD.n22162 DVDD.n284 0.00962857
R45782 DVDD.n334 DVDD.n284 0.00962857
R45783 DVDD.n336 DVDD.n334 0.00962857
R45784 DVDD.n338 DVDD.n336 0.00962857
R45785 DVDD.n338 DVDD.n330 0.00962857
R45786 DVDD.n343 DVDD.n330 0.00962857
R45787 DVDD.n345 DVDD.n343 0.00962857
R45788 DVDD.n347 DVDD.n345 0.00962857
R45789 DVDD.n347 DVDD.n325 0.00962857
R45790 DVDD.n22154 DVDD.n325 0.00962857
R45791 DVDD.n22154 DVDD.n327 0.00962857
R45792 DVDD.n22150 DVDD.n327 0.00962857
R45793 DVDD.n22150 DVDD.n22148 0.00962857
R45794 DVDD.n22148 DVDD.n22147 0.00962857
R45795 DVDD.n22147 DVDD.n351 0.00962857
R45796 DVDD.n22143 DVDD.n351 0.00962857
R45797 DVDD.n22143 DVDD.n353 0.00962857
R45798 DVDD.n399 DVDD.n353 0.00962857
R45799 DVDD.n403 DVDD.n399 0.00962857
R45800 DVDD.n405 DVDD.n403 0.00962857
R45801 DVDD.n407 DVDD.n405 0.00962857
R45802 DVDD.n407 DVDD.n397 0.00962857
R45803 DVDD.n412 DVDD.n397 0.00962857
R45804 DVDD.n414 DVDD.n412 0.00962857
R45805 DVDD.n416 DVDD.n414 0.00962857
R45806 DVDD.n416 DVDD.n394 0.00962857
R45807 DVDD.n420 DVDD.n394 0.00962857
R45808 DVDD.n428 DVDD.n420 0.00962857
R45809 DVDD.n430 DVDD.n428 0.00962857
R45810 DVDD.n430 DVDD.n390 0.00962857
R45811 DVDD.n22136 DVDD.n390 0.00962857
R45812 DVDD.n22136 DVDD.n391 0.00962857
R45813 DVDD.n22132 DVDD.n391 0.00962857
R45814 DVDD.n22132 DVDD.n434 0.00962857
R45815 DVDD.n22128 DVDD.n434 0.00962857
R45816 DVDD.n22128 DVDD.n436 0.00962857
R45817 DVDD.n22124 DVDD.n436 0.00962857
R45818 DVDD.n22124 DVDD.n438 0.00962857
R45819 DVDD.n22094 DVDD.n438 0.00962857
R45820 DVDD.n22096 DVDD.n22094 0.00962857
R45821 DVDD.n22096 DVDD.n22091 0.00962857
R45822 DVDD.n22101 DVDD.n22091 0.00962857
R45823 DVDD.n22103 DVDD.n22101 0.00962857
R45824 DVDD.n22105 DVDD.n22103 0.00962857
R45825 DVDD.n22117 DVDD.n22108 0.00962857
R45826 DVDD.n22118 DVDD.n22117 0.00962857
R45827 DVDD.n3985 DVDD.n3906 0.00962857
R45828 DVDD.n3986 DVDD.n3985 0.00962857
R45829 DVDD.n3988 DVDD.n3986 0.00962857
R45830 DVDD.n3988 DVDD.n3987 0.00962857
R45831 DVDD.n4039 DVDD.n3883 0.00962857
R45832 DVDD.n4039 DVDD.n4038 0.00962857
R45833 DVDD.n4038 DVDD.n4037 0.00962857
R45834 DVDD.n22169 DVDD.n257 0.00962857
R45835 DVDD.n22169 DVDD.n22168 0.00962857
R45836 DVDD.n22168 DVDD.n22167 0.00962857
R45837 DVDD.n22167 DVDD.n280 0.00962857
R45838 DVDD.n22161 DVDD.n280 0.00962857
R45839 DVDD.n354 DVDD.n310 0.00962857
R45840 DVDD.n22142 DVDD.n354 0.00962857
R45841 DVDD.n22142 DVDD.n22141 0.00962857
R45842 DVDD.n22137 DVDD.n389 0.00962857
R45843 DVDD.n22131 DVDD.n389 0.00962857
R45844 DVDD.n22131 DVDD.n22130 0.00962857
R45845 DVDD.n22130 DVDD.n22129 0.00962857
R45846 DVDD.n9839 DVDD.n9837 0.00962857
R45847 DVDD.n9843 DVDD.n9839 0.00962857
R45848 DVDD.n9845 DVDD.n9843 0.00962857
R45849 DVDD.n9847 DVDD.n9845 0.00962857
R45850 DVDD.n9847 DVDD.n9835 0.00962857
R45851 DVDD.n9852 DVDD.n9835 0.00962857
R45852 DVDD.n9854 DVDD.n9852 0.00962857
R45853 DVDD.n9856 DVDD.n9854 0.00962857
R45854 DVDD.n9856 DVDD.n9832 0.00962857
R45855 DVDD.n9861 DVDD.n9832 0.00962857
R45856 DVDD.n9863 DVDD.n9861 0.00962857
R45857 DVDD.n9865 DVDD.n9863 0.00962857
R45858 DVDD.n9865 DVDD.n9829 0.00962857
R45859 DVDD.n9870 DVDD.n9829 0.00962857
R45860 DVDD.n9870 DVDD.n9826 0.00962857
R45861 DVDD.n9874 DVDD.n9826 0.00962857
R45862 DVDD.n9876 DVDD.n9874 0.00962857
R45863 DVDD.n9878 DVDD.n9876 0.00962857
R45864 DVDD.n9878 DVDD.n9824 0.00962857
R45865 DVDD.n9883 DVDD.n9824 0.00962857
R45866 DVDD.n9885 DVDD.n9883 0.00962857
R45867 DVDD.n9887 DVDD.n9885 0.00962857
R45868 DVDD.n9887 DVDD.n9821 0.00962857
R45869 DVDD.n9892 DVDD.n9821 0.00962857
R45870 DVDD.n9894 DVDD.n9892 0.00962857
R45871 DVDD.n9896 DVDD.n9894 0.00962857
R45872 DVDD.n9896 DVDD.n9817 0.00962857
R45873 DVDD.n9936 DVDD.n9817 0.00962857
R45874 DVDD.n9936 DVDD.n9818 0.00962857
R45875 DVDD.n9932 DVDD.n9818 0.00962857
R45876 DVDD.n9932 DVDD.n9931 0.00962857
R45877 DVDD.n9931 DVDD.n9900 0.00962857
R45878 DVDD.n9927 DVDD.n9900 0.00962857
R45879 DVDD.n9927 DVDD.n9902 0.00962857
R45880 DVDD.n9923 DVDD.n9902 0.00962857
R45881 DVDD.n9923 DVDD.n9921 0.00962857
R45882 DVDD.n9921 DVDD.n9919 0.00962857
R45883 DVDD.n9919 DVDD.n9906 0.00962857
R45884 DVDD.n9914 DVDD.n9906 0.00962857
R45885 DVDD.n9914 DVDD.n9912 0.00962857
R45886 DVDD.n9912 DVDD.n9910 0.00962857
R45887 DVDD.n9910 DVDD.n9644 0.00962857
R45888 DVDD.n10089 DVDD.n9644 0.00962857
R45889 DVDD.n10089 DVDD.n9650 0.00962857
R45890 DVDD.n10085 DVDD.n9650 0.00962857
R45891 DVDD.n10085 DVDD.n10083 0.00962857
R45892 DVDD.n10083 DVDD.n10082 0.00962857
R45893 DVDD.n10082 DVDD.n9653 0.00962857
R45894 DVDD.n10078 DVDD.n9653 0.00962857
R45895 DVDD.n10078 DVDD.n9655 0.00962857
R45896 DVDD.n10074 DVDD.n9655 0.00962857
R45897 DVDD.n10074 DVDD.n9658 0.00962857
R45898 DVDD.n10070 DVDD.n9658 0.00962857
R45899 DVDD.n10070 DVDD.n9660 0.00962857
R45900 DVDD.n9708 DVDD.n9660 0.00962857
R45901 DVDD.n9710 DVDD.n9708 0.00962857
R45902 DVDD.n9710 DVDD.n9705 0.00962857
R45903 DVDD.n9715 DVDD.n9705 0.00962857
R45904 DVDD.n9717 DVDD.n9715 0.00962857
R45905 DVDD.n9719 DVDD.n9717 0.00962857
R45906 DVDD.n9719 DVDD.n9702 0.00962857
R45907 DVDD.n9724 DVDD.n9702 0.00962857
R45908 DVDD.n9726 DVDD.n9724 0.00962857
R45909 DVDD.n9728 DVDD.n9726 0.00962857
R45910 DVDD.n9728 DVDD.n9698 0.00962857
R45911 DVDD.n10064 DVDD.n9698 0.00962857
R45912 DVDD.n10064 DVDD.n9699 0.00962857
R45913 DVDD.n10060 DVDD.n9699 0.00962857
R45914 DVDD.n10060 DVDD.n9732 0.00962857
R45915 DVDD.n9975 DVDD.n9732 0.00962857
R45916 DVDD.n9979 DVDD.n9975 0.00962857
R45917 DVDD.n9981 DVDD.n9979 0.00962857
R45918 DVDD.n9983 DVDD.n9981 0.00962857
R45919 DVDD.n9983 DVDD.n9973 0.00962857
R45920 DVDD.n9988 DVDD.n9973 0.00962857
R45921 DVDD.n9990 DVDD.n9988 0.00962857
R45922 DVDD.n9992 DVDD.n9990 0.00962857
R45923 DVDD.n9992 DVDD.n9970 0.00962857
R45924 DVDD.n9996 DVDD.n9970 0.00962857
R45925 DVDD.n10003 DVDD.n9996 0.00962857
R45926 DVDD.n10005 DVDD.n10003 0.00962857
R45927 DVDD.n10005 DVDD.n9966 0.00962857
R45928 DVDD.n10053 DVDD.n9966 0.00962857
R45929 DVDD.n10053 DVDD.n9967 0.00962857
R45930 DVDD.n10049 DVDD.n9967 0.00962857
R45931 DVDD.n10049 DVDD.n10046 0.00962857
R45932 DVDD.n10046 DVDD.n10045 0.00962857
R45933 DVDD.n10045 DVDD.n10009 0.00962857
R45934 DVDD.n10041 DVDD.n10009 0.00962857
R45935 DVDD.n10041 DVDD.n10039 0.00962857
R45936 DVDD.n10039 DVDD.n10037 0.00962857
R45937 DVDD.n10037 DVDD.n10012 0.00962857
R45938 DVDD.n10032 DVDD.n10012 0.00962857
R45939 DVDD.n10032 DVDD.n10030 0.00962857
R45940 DVDD.n10030 DVDD.n10028 0.00962857
R45941 DVDD.n10028 DVDD.n10015 0.00962857
R45942 DVDD.n10023 DVDD.n10021 0.00962857
R45943 DVDD.n10021 DVDD.n10017 0.00962857
R45944 DVDD.n9864 DVDD.n9828 0.00962857
R45945 DVDD.n9871 DVDD.n9828 0.00962857
R45946 DVDD.n9872 DVDD.n9871 0.00962857
R45947 DVDD.n9873 DVDD.n9872 0.00962857
R45948 DVDD.n9930 DVDD.n9807 0.00962857
R45949 DVDD.n9930 DVDD.n9929 0.00962857
R45950 DVDD.n9929 DVDD.n9928 0.00962857
R45951 DVDD.n9656 DVDD.n9632 0.00962857
R45952 DVDD.n10077 DVDD.n9656 0.00962857
R45953 DVDD.n10077 DVDD.n10076 0.00962857
R45954 DVDD.n10076 DVDD.n10075 0.00962857
R45955 DVDD.n10075 DVDD.n9657 0.00962857
R45956 DVDD.n10065 DVDD.n9697 0.00962857
R45957 DVDD.n10059 DVDD.n9697 0.00962857
R45958 DVDD.n10059 DVDD.n10058 0.00962857
R45959 DVDD.n10054 DVDD.n9965 0.00962857
R45960 DVDD.n10048 DVDD.n9965 0.00962857
R45961 DVDD.n10048 DVDD.n10047 0.00962857
R45962 DVDD.n10047 DVDD.n800 0.00962857
R45963 DVDD.n19689 DVDD.n19207 0.00962857
R45964 DVDD.n19689 DVDD.n19688 0.00962857
R45965 DVDD.n19688 DVDD.n19687 0.00962857
R45966 DVDD.n19687 DVDD.n18685 0.00962857
R45967 DVDD.n18723 DVDD.n18720 0.00962857
R45968 DVDD.n21188 DVDD.n18723 0.00962857
R45969 DVDD.n21188 DVDD.n21187 0.00962857
R45970 DVDD.n21159 DVDD.n21158 0.00962857
R45971 DVDD.n21158 DVDD.n21157 0.00962857
R45972 DVDD.n21157 DVDD.n21117 0.00962857
R45973 DVDD.n21151 DVDD.n21117 0.00962857
R45974 DVDD.n21151 DVDD.n112 0.00962857
R45975 DVDD.n22261 DVDD.n22260 0.00962857
R45976 DVDD.n22262 DVDD.n22261 0.00962857
R45977 DVDD.n22262 DVDD.n79 0.00962857
R45978 DVDD.n22306 DVDD.n38 0.00962857
R45979 DVDD.n22307 DVDD.n22306 0.00962857
R45980 DVDD.n22308 DVDD.n22307 0.00962857
R45981 DVDD.n22308 DVDD.n27 0.00962857
R45982 DVDD.n19649 DVDD.n19647 0.00962857
R45983 DVDD.n19654 DVDD.n19647 0.00962857
R45984 DVDD.n19656 DVDD.n19654 0.00962857
R45985 DVDD.n19658 DVDD.n19656 0.00962857
R45986 DVDD.n19658 DVDD.n19643 0.00962857
R45987 DVDD.n19662 DVDD.n19643 0.00962857
R45988 DVDD.n19664 DVDD.n19662 0.00962857
R45989 DVDD.n19666 DVDD.n19664 0.00962857
R45990 DVDD.n19666 DVDD.n19639 0.00962857
R45991 DVDD.n19695 DVDD.n19639 0.00962857
R45992 DVDD.n19695 DVDD.n19640 0.00962857
R45993 DVDD.n19691 DVDD.n19640 0.00962857
R45994 DVDD.n19691 DVDD.n19690 0.00962857
R45995 DVDD.n19690 DVDD.n19670 0.00962857
R45996 DVDD.n19686 DVDD.n19670 0.00962857
R45997 DVDD.n19686 DVDD.n19671 0.00962857
R45998 DVDD.n19682 DVDD.n19671 0.00962857
R45999 DVDD.n19682 DVDD.n19681 0.00962857
R46000 DVDD.n19681 DVDD.n19679 0.00962857
R46001 DVDD.n19679 DVDD.n19675 0.00962857
R46002 DVDD.n19675 DVDD.n18710 0.00962857
R46003 DVDD.n21209 DVDD.n18710 0.00962857
R46004 DVDD.n21209 DVDD.n18712 0.00962857
R46005 DVDD.n21205 DVDD.n18712 0.00962857
R46006 DVDD.n21205 DVDD.n21203 0.00962857
R46007 DVDD.n21203 DVDD.n21201 0.00962857
R46008 DVDD.n21201 DVDD.n18716 0.00962857
R46009 DVDD.n21197 DVDD.n18716 0.00962857
R46010 DVDD.n21197 DVDD.n21195 0.00962857
R46011 DVDD.n21195 DVDD.n21193 0.00962857
R46012 DVDD.n21193 DVDD.n18719 0.00962857
R46013 DVDD.n21189 DVDD.n18719 0.00962857
R46014 DVDD.n21189 DVDD.n18722 0.00962857
R46015 DVDD.n21104 DVDD.n18722 0.00962857
R46016 DVDD.n21104 DVDD.n21101 0.00962857
R46017 DVDD.n21182 DVDD.n21101 0.00962857
R46018 DVDD.n21182 DVDD.n21103 0.00962857
R46019 DVDD.n21178 DVDD.n21103 0.00962857
R46020 DVDD.n21178 DVDD.n21176 0.00962857
R46021 DVDD.n21176 DVDD.n21174 0.00962857
R46022 DVDD.n21174 DVDD.n21109 0.00962857
R46023 DVDD.n21170 DVDD.n21109 0.00962857
R46024 DVDD.n21170 DVDD.n21168 0.00962857
R46025 DVDD.n21168 DVDD.n21166 0.00962857
R46026 DVDD.n21166 DVDD.n21113 0.00962857
R46027 DVDD.n21162 DVDD.n21113 0.00962857
R46028 DVDD.n21162 DVDD.n21160 0.00962857
R46029 DVDD.n21160 DVDD.n21116 0.00962857
R46030 DVDD.n21156 DVDD.n21116 0.00962857
R46031 DVDD.n21156 DVDD.n21118 0.00962857
R46032 DVDD.n21152 DVDD.n21118 0.00962857
R46033 DVDD.n21152 DVDD.n21150 0.00962857
R46034 DVDD.n21150 DVDD.n21149 0.00962857
R46035 DVDD.n21149 DVDD.n21122 0.00962857
R46036 DVDD.n21145 DVDD.n21122 0.00962857
R46037 DVDD.n21145 DVDD.n21143 0.00962857
R46038 DVDD.n21143 DVDD.n21141 0.00962857
R46039 DVDD.n21141 DVDD.n21125 0.00962857
R46040 DVDD.n21137 DVDD.n21125 0.00962857
R46041 DVDD.n21137 DVDD.n21135 0.00962857
R46042 DVDD.n21135 DVDD.n21133 0.00962857
R46043 DVDD.n21133 DVDD.n21129 0.00962857
R46044 DVDD.n21129 DVDD.n88 0.00962857
R46045 DVDD.n22255 DVDD.n88 0.00962857
R46046 DVDD.n22255 DVDD.n86 0.00962857
R46047 DVDD.n22259 DVDD.n86 0.00962857
R46048 DVDD.n22259 DVDD.n84 0.00962857
R46049 DVDD.n22263 DVDD.n84 0.00962857
R46050 DVDD.n22263 DVDD.n80 0.00962857
R46051 DVDD.n22295 DVDD.n80 0.00962857
R46052 DVDD.n22295 DVDD.n82 0.00962857
R46053 DVDD.n22291 DVDD.n82 0.00962857
R46054 DVDD.n22291 DVDD.n22289 0.00962857
R46055 DVDD.n22289 DVDD.n22287 0.00962857
R46056 DVDD.n22287 DVDD.n22268 0.00962857
R46057 DVDD.n22283 DVDD.n22268 0.00962857
R46058 DVDD.n22283 DVDD.n22281 0.00962857
R46059 DVDD.n22281 DVDD.n22279 0.00962857
R46060 DVDD.n22279 DVDD.n22272 0.00962857
R46061 DVDD.n22275 DVDD.n22272 0.00962857
R46062 DVDD.n22275 DVDD.n41 0.00962857
R46063 DVDD.n22301 DVDD.n41 0.00962857
R46064 DVDD.n22301 DVDD.n39 0.00962857
R46065 DVDD.n22305 DVDD.n39 0.00962857
R46066 DVDD.n22305 DVDD.n37 0.00962857
R46067 DVDD.n22309 DVDD.n37 0.00962857
R46068 DVDD.n22309 DVDD.n33 0.00962857
R46069 DVDD.n22334 DVDD.n33 0.00962857
R46070 DVDD.n22334 DVDD.n35 0.00962857
R46071 DVDD.n22330 DVDD.n35 0.00962857
R46072 DVDD.n22330 DVDD.n22328 0.00962857
R46073 DVDD.n22328 DVDD.n22326 0.00962857
R46074 DVDD.n22326 DVDD.n22314 0.00962857
R46075 DVDD.n22322 DVDD.n22314 0.00962857
R46076 DVDD.n22322 DVDD.n22320 0.00962857
R46077 DVDD.n22320 DVDD.n22318 0.00962857
R46078 DVDD.n22350 DVDD.n2 0.00962857
R46079 DVDD.n22346 DVDD.n2 0.00962857
R46080 DVDD.n22234 DVDD.n22233 0.00959285
R46081 DVDD.n22233 DVDD.n22232 0.00959285
R46082 DVDD.n21722 DVDD.n18431 0.00959285
R46083 DVDD.n21730 DVDD.n18431 0.00959285
R46084 DVDD.n21925 DVDD.n21924 0.00959285
R46085 DVDD.n21924 DVDD.n21923 0.00959285
R46086 DVDD.n18208 DVDD.n213 0.00959285
R46087 DVDD.n22066 DVDD.n18208 0.00959285
R46088 DVDD.n21774 DVDD.n21772 0.00959285
R46089 DVDD.n21774 DVDD.n21773 0.00959285
R46090 DVDD.n21938 DVDD.n21937 0.00959285
R46091 DVDD.n18119 DVDD.n18118 0.00959285
R46092 DVDD.n18118 DVDD.n18117 0.00959285
R46093 DVDD.n18111 DVDD.n18110 0.00959285
R46094 DVDD.n18110 DVDD.n18109 0.00959285
R46095 DVDD.n9571 DVDD.n8974 0.00956767
R46096 DVDD.n21927 DVDD.n21792 0.00956522
R46097 DVDD.n21771 DVDD.n18390 0.00956522
R46098 DVDD.n18478 DVDD.n134 0.00943276
R46099 DVDD.n21920 DVDD.n21796 0.00943276
R46100 DVDD.n18101 DVDD.n18097 0.00943276
R46101 DVDD.n15141 DVDD.n5579 0.00937536
R46102 DVDD.n5585 DVDD.n5582 0.00937536
R46103 DVDD.n899 DVDD.n896 0.00937536
R46104 DVDD.n900 DVDD.n899 0.00937536
R46105 DVDD.n5586 DVDD.n5579 0.00937536
R46106 DVDD.n5586 DVDD.n5585 0.00937536
R46107 DVDD.n21674 DVDD.n21673 0.00936443
R46108 DVDD.n21358 DVDD.n21338 0.00936443
R46109 DVDD.n22000 DVDD.n21998 0.00936443
R46110 DVDD.n4857 DVDD.n3545 0.00936443
R46111 DVDD.n12729 DVDD.n12478 0.00934279
R46112 DVDD.n13259 DVDD.n12913 0.00934279
R46113 DVDD.n13481 DVDD.n13480 0.00934279
R46114 DVDD.n13260 DVDD.n12914 0.00934279
R46115 DVDD.n13761 DVDD.n11929 0.00929699
R46116 DVDD.n18414 DVDD.n18399 0.009275
R46117 DVDD.n22015 DVDD.n22014 0.009275
R46118 DVDD.n21352 DVDD.n21340 0.009275
R46119 DVDD.n21702 DVDD.n18521 0.009275
R46120 DVDD.n18252 DVDD.n18251 0.009275
R46121 DVDD.n18436 DVDD.n163 0.009275
R46122 DVDD.n4291 DVDD.n4290 0.009275
R46123 DVDD.n3691 DVDD.n3678 0.009275
R46124 DVDD.n10234 DVDD.n8611 0.00919799
R46125 DVDD.n17297 DVDD.n916 0.00919799
R46126 DVDD.n10235 DVDD.n8613 0.00919799
R46127 DVDD.n17296 DVDD.n917 0.00919799
R46128 DVDD.n13812 DVDD.n13811 0.00916165
R46129 DVDD.n16720 DVDD.n16719 0.00916165
R46130 DVDD.n2734 DVDD.n2656 0.00901707
R46131 DVDD.n2804 DVDD.n2583 0.00901707
R46132 DVDD.n3247 DVDD.n3174 0.00901707
R46133 DVDD.n15534 DVDD.n15533 0.00901707
R46134 DVDD.n14561 DVDD.n8156 0.00894978
R46135 DVDD.n17716 DVDD.n909 0.00894978
R46136 DVDD.n14562 DVDD.n8157 0.00894978
R46137 DVDD.n17715 DVDD.n911 0.00894978
R46138 DVDD.n22347 DVDD.n22346 0.00881417
R46139 DVDD.n19650 DVDD.n19649 0.00881417
R46140 DVDD.n20140 DVDD.n20139 0.00880519
R46141 DVDD.n20335 DVDD.n18950 0.00880519
R46142 DVDD.n20627 DVDD.n20626 0.00880519
R46143 DVDD.n18998 DVDD.n18979 0.00880519
R46144 DVDD.n3974 DVDD.n3934 0.00880519
R46145 DVDD.n22119 DVDD.n22118 0.00880519
R46146 DVDD.n9837 DVDD.n5486 0.00880519
R46147 DVDD.n10018 DVDD.n10017 0.00880519
R46148 DVDD DVDD.n21940 0.00876041
R46149 DVDD.n21939 DVDD 0.00876041
R46150 DVDD.n4557 DVDD.n4388 0.00875734
R46151 DVDD.n4531 DVDD.n4388 0.00875734
R46152 DVDD.n15093 DVDD.n6705 0.00871477
R46153 DVDD.n14848 DVDD.n7680 0.00871477
R46154 DVDD.n15094 DVDD.n6704 0.00871477
R46155 DVDD.n14847 DVDD.n7682 0.00871477
R46156 DVDD.n17612 DVDD.n911 0.0087125
R46157 DVDD.n17371 DVDD.n909 0.0087125
R46158 DVDD.n15129 DVDD.n5743 0.0087125
R46159 DVDD.n15130 DVDD.n5741 0.0087125
R46160 DVDD.n21777 DVDD.n21776 0.00866435
R46161 DVDD.n21725 DVDD.n159 0.00866435
R46162 DVDD.n22043 DVDD.n22042 0.00866435
R46163 DVDD.n18095 DVDD.n18094 0.00866435
R46164 DVDD.n13812 DVDD.n11212 0.0086203
R46165 DVDD.n16723 DVDD.n16720 0.0086203
R46166 DVDD.n18344 DVDD.n18343 0.00859753
R46167 DVDD.n4847 DVDD.n3548 0.00859753
R46168 DVDD.n4751 DVDD.n4750 0.0084875
R46169 DVDD.n4750 DVDD.n3718 0.0084875
R46170 DVDD.n4744 DVDD.n3718 0.0084875
R46171 DVDD.n3633 DVDD.n3603 0.0084875
R46172 DVDD.n4778 DVDD.n4777 0.0084875
R46173 DVDD.n4777 DVDD.n4776 0.0084875
R46174 DVDD.n4590 DVDD.n4589 0.0084875
R46175 DVDD.n4589 DVDD.n488 0.0084875
R46176 DVDD.n18133 DVDD.n489 0.0084875
R46177 DVDD.n4576 DVDD.n4279 0.0084875
R46178 DVDD.n4580 DVDD.n4279 0.0084875
R46179 DVDD.n4581 DVDD.n4580 0.0084875
R46180 DVDD.n4582 DVDD.n4581 0.0084875
R46181 DVDD.n4582 DVDD.n4274 0.0084875
R46182 DVDD.n4595 DVDD.n4274 0.0084875
R46183 DVDD.n4595 DVDD.n4276 0.0084875
R46184 DVDD.n4591 DVDD.n4276 0.0084875
R46185 DVDD.n4591 DVDD.n4588 0.0084875
R46186 DVDD.n4588 DVDD.n4587 0.0084875
R46187 DVDD.n18132 DVDD.n491 0.0084875
R46188 DVDD.n18128 DVDD.n491 0.0084875
R46189 DVDD.n18128 DVDD.n495 0.0084875
R46190 DVDD.n18073 DVDD.n495 0.0084875
R46191 DVDD.n18077 DVDD.n18073 0.0084875
R46192 DVDD.n18079 DVDD.n18077 0.0084875
R46193 DVDD.n18087 DVDD.n18079 0.0084875
R46194 DVDD.n18087 DVDD.n18069 0.0084875
R46195 DVDD.n18091 DVDD.n18069 0.0084875
R46196 DVDD.n3615 DVDD.n3612 0.0084875
R46197 DVDD.n3617 DVDD.n3615 0.0084875
R46198 DVDD.n3619 DVDD.n3617 0.0084875
R46199 DVDD.n3619 DVDD.n3608 0.0084875
R46200 DVDD.n3623 DVDD.n3608 0.0084875
R46201 DVDD.n3625 DVDD.n3623 0.0084875
R46202 DVDD.n3627 DVDD.n3625 0.0084875
R46203 DVDD.n3627 DVDD.n3605 0.0084875
R46204 DVDD.n3631 DVDD.n3605 0.0084875
R46205 DVDD.n3632 DVDD.n3631 0.0084875
R46206 DVDD.n4779 DVDD.n3602 0.0084875
R46207 DVDD.n4775 DVDD.n3602 0.0084875
R46208 DVDD.n4775 DVDD.n3636 0.0084875
R46209 DVDD.n4771 DVDD.n3636 0.0084875
R46210 DVDD.n4771 DVDD.n3638 0.0084875
R46211 DVDD.n3669 DVDD.n3638 0.0084875
R46212 DVDD.n4765 DVDD.n3669 0.0084875
R46213 DVDD.n4765 DVDD.n3671 0.0084875
R46214 DVDD.n4761 DVDD.n3671 0.0084875
R46215 DVDD.n4455 DVDD.n4412 0.0084875
R46216 DVDD.n4553 DVDD.n4412 0.0084875
R46217 DVDD.n4553 DVDD.n4414 0.0084875
R46218 DVDD.n4549 DVDD.n4414 0.0084875
R46219 DVDD.n4549 DVDD.n4547 0.0084875
R46220 DVDD.n4547 DVDD.n4545 0.0084875
R46221 DVDD.n4545 DVDD.n4460 0.0084875
R46222 DVDD.n4540 DVDD.n4460 0.0084875
R46223 DVDD.n4540 DVDD.n4538 0.0084875
R46224 DVDD.n4538 DVDD.n4536 0.0084875
R46225 DVDD.n4477 DVDD.n4476 0.0084875
R46226 DVDD.n4476 DVDD.n4322 0.0084875
R46227 DVDD.n4560 DVDD.n4322 0.0084875
R46228 DVDD.n4560 DVDD.n4320 0.0084875
R46229 DVDD.n4564 DVDD.n4320 0.0084875
R46230 DVDD.n4564 DVDD.n4318 0.0084875
R46231 DVDD.n4568 DVDD.n4318 0.0084875
R46232 DVDD.n4568 DVDD.n4316 0.0084875
R46233 DVDD.n4572 DVDD.n4316 0.0084875
R46234 DVDD.n4758 DVDD.n3676 0.0084875
R46235 DVDD.n4754 DVDD.n3676 0.0084875
R46236 DVDD.n4754 DVDD.n3715 0.0084875
R46237 DVDD.n4749 DVDD.n3715 0.0084875
R46238 DVDD.n4749 DVDD.n3719 0.0084875
R46239 DVDD.n4745 DVDD.n3719 0.0084875
R46240 DVDD.n4745 DVDD.n3721 0.0084875
R46241 DVDD.n3754 DVDD.n3721 0.0084875
R46242 DVDD.n4739 DVDD.n3754 0.0084875
R46243 DVDD.n4739 DVDD.n3755 0.0084875
R46244 DVDD.n4431 DVDD.n4428 0.0084875
R46245 DVDD.n4433 DVDD.n4431 0.0084875
R46246 DVDD.n4435 DVDD.n4433 0.0084875
R46247 DVDD.n4435 DVDD.n4424 0.0084875
R46248 DVDD.n4439 DVDD.n4424 0.0084875
R46249 DVDD.n4443 DVDD.n4439 0.0084875
R46250 DVDD.n4445 DVDD.n4443 0.0084875
R46251 DVDD.n4445 DVDD.n4421 0.0084875
R46252 DVDD.n4449 DVDD.n4421 0.0084875
R46253 DVDD.n4454 DVDD.n4407 0.0084875
R46254 DVDD.n4565 DVDD.n4319 0.0084875
R46255 DVDD.n4566 DVDD.n4565 0.0084875
R46256 DVDD.n4567 DVDD.n4566 0.0084875
R46257 DVDD.n11929 DVDD.n11585 0.00848496
R46258 DVDD.n17515 DVDD.n893 0.008375
R46259 DVDD.n14853 DVDD.n7674 0.008375
R46260 DVDD.n15136 DVDD.n15135 0.008375
R46261 DVDD.n20048 DVDD.n19736 0.00834286
R46262 DVDD.n20264 DVDD.n19939 0.00834286
R46263 DVDD.n19170 DVDD.n18843 0.00834286
R46264 DVDD.n20756 DVDD.n19049 0.00834286
R46265 DVDD.n3900 DVDD.n3872 0.00834286
R46266 DVDD.n337 DVDD.n300 0.00834286
R46267 DVDD.n9886 DVDD.n9768 0.00834286
R46268 DVDD.n9709 DVDD.n9690 0.00834286
R46269 DVDD.n21210 DVDD.n18679 0.00834286
R46270 DVDD.n21142 DVDD.n100 0.00834286
R46271 DVDD.n21944 DVDD.n18302 0.00832155
R46272 DVDD.n22209 DVDD.n184 0.00832155
R46273 DVDD.n22229 DVDD.n143 0.00832155
R46274 DVDD.n22039 DVDD.n18245 0.00832155
R46275 DVDD.n18336 DVDD.n223 0.00832155
R46276 DVDD.n21263 DVDD.n18432 0.00832155
R46277 DVDD.n4864 DVDD.n3540 0.00832155
R46278 DVDD.n4863 DVDD.n3541 0.00832155
R46279 DVDD.n21680 DVDD.n18535 0.00830425
R46280 DVDD.n18369 DVDD.n18368 0.00830425
R46281 DVDD.n22005 DVDD.n22004 0.00830425
R46282 DVDD.n21366 DVDD.n21334 0.00830425
R46283 DVDD.n21268 DVDD.n18656 0.00830425
R46284 DVDD.n4878 DVDD.n3533 0.00830425
R46285 DVDD.n20330 DVDD.n18941 0.00827857
R46286 DVDD.n20836 DVDD.n18969 0.00827857
R46287 DVDD.n22095 DVDD.n22077 0.00827857
R46288 DVDD.n10011 DVDD.n797 0.00827857
R46289 DVDD.n22315 DVDD.n24 0.00827857
R46290 DVDD.n13809 DVDD.n11105 0.00823154
R46291 DVDD.n16717 DVDD.n1814 0.00823154
R46292 DVDD.n13810 DVDD.n11224 0.00823154
R46293 DVDD.n16718 DVDD.n1815 0.00823154
R46294 DVDD.n20572 DVDD.n19740 0.00821429
R46295 DVDD.n20283 DVDD.n20281 0.00821429
R46296 DVDD.n20970 DVDD.n18847 0.00821429
R46297 DVDD.n20777 DVDD.n19054 0.00821429
R46298 DVDD.n4065 DVDD.n3876 0.00821429
R46299 DVDD.n326 DVDD.n303 0.00821429
R46300 DVDD.n9948 DVDD.n9773 0.00821429
R46301 DVDD.n9725 DVDD.n9695 0.00821429
R46302 DVDD.n9571 DVDD.n9570 0.00821429
R46303 DVDD.n21194 DVDD.n18702 0.00821429
R46304 DVDD.n105 DVDD.n89 0.00821429
R46305 DVDD.n20883 DVDD.n18945 0.00815
R46306 DVDD.n20854 DVDD.n18973 0.00815
R46307 DVDD.n22120 DVDD.n22087 0.00815
R46308 DVDD.n10016 DVDD.n796 0.00815
R46309 DVDD.n22345 DVDD.n4 0.00815
R46310 DVDD.n20234 DVDD.n19972 0.00808571
R46311 DVDD.n20312 DVDD.n19837 0.00808571
R46312 DVDD.n20726 DVDD.n19135 0.00808571
R46313 DVDD.n20803 DVDD.n18883 0.00808571
R46314 DVDD.n272 DVDD.n238 0.00808571
R46315 DVDD.n415 DVDD.n375 0.00808571
R46316 DVDD.n10090 DVDD.n9615 0.00808571
R46317 DVDD.n9991 DVDD.n9752 0.00808571
R46318 DVDD.n21167 DVDD.n21095 0.00808571
R46319 DVDD.n22280 DVDD.n74 0.00808571
R46320 DVDD.n7064 DVDD.n6703 0.00807895
R46321 DVDD.n9564 DVDD.n7684 0.00807895
R46322 DVDD.n20154 DVDD.n20127 0.00802143
R46323 DVDD.n20641 DVDD.n20614 0.00802143
R46324 DVDD.n3951 DVDD.n3930 0.00802143
R46325 DVDD.n9853 DVDD.n5481 0.00802143
R46326 DVDD.n19663 DVDD.n19198 0.00802143
R46327 DVDD.n18121 DVDD.n18064 0.0080019
R46328 DVDD.n17722 DVDD.n894 0.00796421
R46329 DVDD.n17725 DVDD.n895 0.00796421
R46330 DVDD.n17365 DVDD.n17361 0.00796421
R46331 DVDD.n17363 DVDD.n898 0.00796421
R46332 DVDD.n17709 DVDD.n17513 0.00796421
R46333 DVDD.n17514 DVDD.n17313 0.00796421
R46334 DVDD.n17512 DVDD.n17510 0.00796421
R46335 DVDD.n17511 DVDD.n17314 0.00796421
R46336 DVDD.n17509 DVDD.n17507 0.00796421
R46337 DVDD.n17508 DVDD.n17315 0.00796421
R46338 DVDD.n17506 DVDD.n17504 0.00796421
R46339 DVDD.n17505 DVDD.n17316 0.00796421
R46340 DVDD.n17503 DVDD.n17501 0.00796421
R46341 DVDD.n17502 DVDD.n17317 0.00796421
R46342 DVDD.n17500 DVDD.n17498 0.00796421
R46343 DVDD.n17499 DVDD.n17318 0.00796421
R46344 DVDD.n17497 DVDD.n17495 0.00796421
R46345 DVDD.n17496 DVDD.n17319 0.00796421
R46346 DVDD.n17494 DVDD.n17492 0.00796421
R46347 DVDD.n17493 DVDD.n17320 0.00796421
R46348 DVDD.n17491 DVDD.n17489 0.00796421
R46349 DVDD.n17490 DVDD.n17321 0.00796421
R46350 DVDD.n17488 DVDD.n17486 0.00796421
R46351 DVDD.n17487 DVDD.n17322 0.00796421
R46352 DVDD.n17485 DVDD.n17483 0.00796421
R46353 DVDD.n17484 DVDD.n17323 0.00796421
R46354 DVDD.n17482 DVDD.n17480 0.00796421
R46355 DVDD.n17481 DVDD.n17324 0.00796421
R46356 DVDD.n17479 DVDD.n17477 0.00796421
R46357 DVDD.n17478 DVDD.n17325 0.00796421
R46358 DVDD.n17476 DVDD.n17474 0.00796421
R46359 DVDD.n17475 DVDD.n17326 0.00796421
R46360 DVDD.n17473 DVDD.n17471 0.00796421
R46361 DVDD.n17472 DVDD.n17327 0.00796421
R46362 DVDD.n17470 DVDD.n17468 0.00796421
R46363 DVDD.n17469 DVDD.n17328 0.00796421
R46364 DVDD.n17467 DVDD.n17465 0.00796421
R46365 DVDD.n17466 DVDD.n17329 0.00796421
R46366 DVDD.n17464 DVDD.n17462 0.00796421
R46367 DVDD.n17463 DVDD.n17330 0.00796421
R46368 DVDD.n17461 DVDD.n17459 0.00796421
R46369 DVDD.n17460 DVDD.n17331 0.00796421
R46370 DVDD.n17458 DVDD.n17456 0.00796421
R46371 DVDD.n17457 DVDD.n17332 0.00796421
R46372 DVDD.n17455 DVDD.n17453 0.00796421
R46373 DVDD.n17454 DVDD.n17333 0.00796421
R46374 DVDD.n17452 DVDD.n17450 0.00796421
R46375 DVDD.n17451 DVDD.n17334 0.00796421
R46376 DVDD.n17449 DVDD.n17447 0.00796421
R46377 DVDD.n17448 DVDD.n17335 0.00796421
R46378 DVDD.n17446 DVDD.n17444 0.00796421
R46379 DVDD.n17445 DVDD.n17336 0.00796421
R46380 DVDD.n17443 DVDD.n17441 0.00796421
R46381 DVDD.n17442 DVDD.n17337 0.00796421
R46382 DVDD.n17440 DVDD.n17438 0.00796421
R46383 DVDD.n17439 DVDD.n17338 0.00796421
R46384 DVDD.n17437 DVDD.n17435 0.00796421
R46385 DVDD.n17436 DVDD.n17339 0.00796421
R46386 DVDD.n17434 DVDD.n17432 0.00796421
R46387 DVDD.n17433 DVDD.n17340 0.00796421
R46388 DVDD.n17431 DVDD.n17429 0.00796421
R46389 DVDD.n17430 DVDD.n17341 0.00796421
R46390 DVDD.n17428 DVDD.n17426 0.00796421
R46391 DVDD.n17427 DVDD.n17342 0.00796421
R46392 DVDD.n17425 DVDD.n17423 0.00796421
R46393 DVDD.n17424 DVDD.n17343 0.00796421
R46394 DVDD.n17422 DVDD.n17420 0.00796421
R46395 DVDD.n17421 DVDD.n17344 0.00796421
R46396 DVDD.n17419 DVDD.n17417 0.00796421
R46397 DVDD.n17418 DVDD.n17345 0.00796421
R46398 DVDD.n17416 DVDD.n17414 0.00796421
R46399 DVDD.n17415 DVDD.n17346 0.00796421
R46400 DVDD.n17413 DVDD.n17411 0.00796421
R46401 DVDD.n17412 DVDD.n17347 0.00796421
R46402 DVDD.n17410 DVDD.n17408 0.00796421
R46403 DVDD.n17409 DVDD.n17348 0.00796421
R46404 DVDD.n17407 DVDD.n17405 0.00796421
R46405 DVDD.n17406 DVDD.n17349 0.00796421
R46406 DVDD.n17404 DVDD.n17402 0.00796421
R46407 DVDD.n17403 DVDD.n17350 0.00796421
R46408 DVDD.n17401 DVDD.n17399 0.00796421
R46409 DVDD.n17400 DVDD.n17351 0.00796421
R46410 DVDD.n17398 DVDD.n17396 0.00796421
R46411 DVDD.n17397 DVDD.n17352 0.00796421
R46412 DVDD.n17395 DVDD.n17393 0.00796421
R46413 DVDD.n17394 DVDD.n17353 0.00796421
R46414 DVDD.n17392 DVDD.n17390 0.00796421
R46415 DVDD.n17391 DVDD.n17354 0.00796421
R46416 DVDD.n17389 DVDD.n17387 0.00796421
R46417 DVDD.n17388 DVDD.n17355 0.00796421
R46418 DVDD.n17386 DVDD.n17384 0.00796421
R46419 DVDD.n17385 DVDD.n17356 0.00796421
R46420 DVDD.n17383 DVDD.n17381 0.00796421
R46421 DVDD.n17382 DVDD.n17357 0.00796421
R46422 DVDD.n17380 DVDD.n17378 0.00796421
R46423 DVDD.n17379 DVDD.n17358 0.00796421
R46424 DVDD.n17377 DVDD.n17375 0.00796421
R46425 DVDD.n17376 DVDD.n17359 0.00796421
R46426 DVDD.n17374 DVDD.n17372 0.00796421
R46427 DVDD.n17373 DVDD.n17360 0.00796421
R46428 DVDD.n17371 DVDD.n17370 0.00796421
R46429 DVDD.n15137 DVDD.n5580 0.00796421
R46430 DVDD.n15140 DVDD.n5581 0.00796421
R46431 DVDD.n5989 DVDD.n5936 0.00796421
R46432 DVDD.n5937 DVDD.n5584 0.00796421
R46433 DVDD.n15132 DVDD.n5590 0.00796421
R46434 DVDD.n5645 DVDD.n5591 0.00796421
R46435 DVDD.n5985 DVDD.n5640 0.00796421
R46436 DVDD.n5694 DVDD.n5646 0.00796421
R46437 DVDD.n5984 DVDD.n5639 0.00796421
R46438 DVDD.n5695 DVDD.n5647 0.00796421
R46439 DVDD.n5983 DVDD.n5638 0.00796421
R46440 DVDD.n5696 DVDD.n5648 0.00796421
R46441 DVDD.n5982 DVDD.n5637 0.00796421
R46442 DVDD.n5697 DVDD.n5649 0.00796421
R46443 DVDD.n5981 DVDD.n5636 0.00796421
R46444 DVDD.n5698 DVDD.n5650 0.00796421
R46445 DVDD.n5980 DVDD.n5635 0.00796421
R46446 DVDD.n5699 DVDD.n5651 0.00796421
R46447 DVDD.n5979 DVDD.n5634 0.00796421
R46448 DVDD.n5700 DVDD.n5652 0.00796421
R46449 DVDD.n5978 DVDD.n5633 0.00796421
R46450 DVDD.n5701 DVDD.n5653 0.00796421
R46451 DVDD.n5977 DVDD.n5632 0.00796421
R46452 DVDD.n5702 DVDD.n5654 0.00796421
R46453 DVDD.n5976 DVDD.n5631 0.00796421
R46454 DVDD.n5703 DVDD.n5655 0.00796421
R46455 DVDD.n5975 DVDD.n5630 0.00796421
R46456 DVDD.n5704 DVDD.n5656 0.00796421
R46457 DVDD.n5974 DVDD.n5629 0.00796421
R46458 DVDD.n5705 DVDD.n5657 0.00796421
R46459 DVDD.n5973 DVDD.n5628 0.00796421
R46460 DVDD.n5706 DVDD.n5658 0.00796421
R46461 DVDD.n5972 DVDD.n5627 0.00796421
R46462 DVDD.n5707 DVDD.n5659 0.00796421
R46463 DVDD.n5971 DVDD.n5626 0.00796421
R46464 DVDD.n5708 DVDD.n5660 0.00796421
R46465 DVDD.n5970 DVDD.n5625 0.00796421
R46466 DVDD.n5709 DVDD.n5661 0.00796421
R46467 DVDD.n5969 DVDD.n5624 0.00796421
R46468 DVDD.n5710 DVDD.n5662 0.00796421
R46469 DVDD.n5968 DVDD.n5623 0.00796421
R46470 DVDD.n5711 DVDD.n5663 0.00796421
R46471 DVDD.n5967 DVDD.n5622 0.00796421
R46472 DVDD.n5712 DVDD.n5664 0.00796421
R46473 DVDD.n5966 DVDD.n5621 0.00796421
R46474 DVDD.n5713 DVDD.n5665 0.00796421
R46475 DVDD.n5965 DVDD.n5620 0.00796421
R46476 DVDD.n5714 DVDD.n5666 0.00796421
R46477 DVDD.n5964 DVDD.n5619 0.00796421
R46478 DVDD.n5715 DVDD.n5667 0.00796421
R46479 DVDD.n5963 DVDD.n5618 0.00796421
R46480 DVDD.n5716 DVDD.n5668 0.00796421
R46481 DVDD.n5962 DVDD.n5617 0.00796421
R46482 DVDD.n5717 DVDD.n5669 0.00796421
R46483 DVDD.n5961 DVDD.n5616 0.00796421
R46484 DVDD.n5718 DVDD.n5670 0.00796421
R46485 DVDD.n5960 DVDD.n5615 0.00796421
R46486 DVDD.n5719 DVDD.n5671 0.00796421
R46487 DVDD.n5959 DVDD.n5614 0.00796421
R46488 DVDD.n5720 DVDD.n5672 0.00796421
R46489 DVDD.n5958 DVDD.n5613 0.00796421
R46490 DVDD.n5721 DVDD.n5673 0.00796421
R46491 DVDD.n5957 DVDD.n5612 0.00796421
R46492 DVDD.n5722 DVDD.n5674 0.00796421
R46493 DVDD.n5956 DVDD.n5611 0.00796421
R46494 DVDD.n5723 DVDD.n5675 0.00796421
R46495 DVDD.n5955 DVDD.n5610 0.00796421
R46496 DVDD.n5724 DVDD.n5676 0.00796421
R46497 DVDD.n5954 DVDD.n5609 0.00796421
R46498 DVDD.n5725 DVDD.n5677 0.00796421
R46499 DVDD.n5953 DVDD.n5608 0.00796421
R46500 DVDD.n5726 DVDD.n5678 0.00796421
R46501 DVDD.n5952 DVDD.n5607 0.00796421
R46502 DVDD.n5727 DVDD.n5679 0.00796421
R46503 DVDD.n5951 DVDD.n5606 0.00796421
R46504 DVDD.n5728 DVDD.n5680 0.00796421
R46505 DVDD.n5950 DVDD.n5605 0.00796421
R46506 DVDD.n5729 DVDD.n5681 0.00796421
R46507 DVDD.n5949 DVDD.n5604 0.00796421
R46508 DVDD.n5730 DVDD.n5682 0.00796421
R46509 DVDD.n5948 DVDD.n5603 0.00796421
R46510 DVDD.n5731 DVDD.n5683 0.00796421
R46511 DVDD.n5947 DVDD.n5602 0.00796421
R46512 DVDD.n5732 DVDD.n5684 0.00796421
R46513 DVDD.n5946 DVDD.n5601 0.00796421
R46514 DVDD.n5733 DVDD.n5685 0.00796421
R46515 DVDD.n5945 DVDD.n5600 0.00796421
R46516 DVDD.n5734 DVDD.n5686 0.00796421
R46517 DVDD.n5944 DVDD.n5599 0.00796421
R46518 DVDD.n5735 DVDD.n5687 0.00796421
R46519 DVDD.n5943 DVDD.n5598 0.00796421
R46520 DVDD.n5736 DVDD.n5688 0.00796421
R46521 DVDD.n5942 DVDD.n5597 0.00796421
R46522 DVDD.n5737 DVDD.n5689 0.00796421
R46523 DVDD.n5941 DVDD.n5596 0.00796421
R46524 DVDD.n5738 DVDD.n5690 0.00796421
R46525 DVDD.n5940 DVDD.n5595 0.00796421
R46526 DVDD.n5739 DVDD.n5691 0.00796421
R46527 DVDD.n5939 DVDD.n5594 0.00796421
R46528 DVDD.n5693 DVDD.n5641 0.00796421
R46529 DVDD.n15130 DVDD.n5692 0.00796421
R46530 DVDD.n5692 DVDD.n5641 0.00796421
R46531 DVDD.n17370 DVDD.n17360 0.00796421
R46532 DVDD.n17374 DVDD.n17373 0.00796421
R46533 DVDD.n17372 DVDD.n17359 0.00796421
R46534 DVDD.n17377 DVDD.n17376 0.00796421
R46535 DVDD.n17375 DVDD.n17358 0.00796421
R46536 DVDD.n17380 DVDD.n17379 0.00796421
R46537 DVDD.n17378 DVDD.n17357 0.00796421
R46538 DVDD.n17383 DVDD.n17382 0.00796421
R46539 DVDD.n17381 DVDD.n17356 0.00796421
R46540 DVDD.n17386 DVDD.n17385 0.00796421
R46541 DVDD.n17384 DVDD.n17355 0.00796421
R46542 DVDD.n17389 DVDD.n17388 0.00796421
R46543 DVDD.n17387 DVDD.n17354 0.00796421
R46544 DVDD.n17392 DVDD.n17391 0.00796421
R46545 DVDD.n17390 DVDD.n17353 0.00796421
R46546 DVDD.n17395 DVDD.n17394 0.00796421
R46547 DVDD.n17393 DVDD.n17352 0.00796421
R46548 DVDD.n17398 DVDD.n17397 0.00796421
R46549 DVDD.n17396 DVDD.n17351 0.00796421
R46550 DVDD.n17401 DVDD.n17400 0.00796421
R46551 DVDD.n17399 DVDD.n17350 0.00796421
R46552 DVDD.n17404 DVDD.n17403 0.00796421
R46553 DVDD.n17402 DVDD.n17349 0.00796421
R46554 DVDD.n17407 DVDD.n17406 0.00796421
R46555 DVDD.n17405 DVDD.n17348 0.00796421
R46556 DVDD.n17410 DVDD.n17409 0.00796421
R46557 DVDD.n17408 DVDD.n17347 0.00796421
R46558 DVDD.n17413 DVDD.n17412 0.00796421
R46559 DVDD.n17411 DVDD.n17346 0.00796421
R46560 DVDD.n17416 DVDD.n17415 0.00796421
R46561 DVDD.n17414 DVDD.n17345 0.00796421
R46562 DVDD.n17419 DVDD.n17418 0.00796421
R46563 DVDD.n17417 DVDD.n17344 0.00796421
R46564 DVDD.n17422 DVDD.n17421 0.00796421
R46565 DVDD.n17420 DVDD.n17343 0.00796421
R46566 DVDD.n17425 DVDD.n17424 0.00796421
R46567 DVDD.n17423 DVDD.n17342 0.00796421
R46568 DVDD.n17428 DVDD.n17427 0.00796421
R46569 DVDD.n17426 DVDD.n17341 0.00796421
R46570 DVDD.n17431 DVDD.n17430 0.00796421
R46571 DVDD.n17429 DVDD.n17340 0.00796421
R46572 DVDD.n17434 DVDD.n17433 0.00796421
R46573 DVDD.n17432 DVDD.n17339 0.00796421
R46574 DVDD.n17437 DVDD.n17436 0.00796421
R46575 DVDD.n17435 DVDD.n17338 0.00796421
R46576 DVDD.n17440 DVDD.n17439 0.00796421
R46577 DVDD.n17438 DVDD.n17337 0.00796421
R46578 DVDD.n17443 DVDD.n17442 0.00796421
R46579 DVDD.n17441 DVDD.n17336 0.00796421
R46580 DVDD.n17446 DVDD.n17445 0.00796421
R46581 DVDD.n17444 DVDD.n17335 0.00796421
R46582 DVDD.n17449 DVDD.n17448 0.00796421
R46583 DVDD.n17447 DVDD.n17334 0.00796421
R46584 DVDD.n17452 DVDD.n17451 0.00796421
R46585 DVDD.n17450 DVDD.n17333 0.00796421
R46586 DVDD.n17455 DVDD.n17454 0.00796421
R46587 DVDD.n17453 DVDD.n17332 0.00796421
R46588 DVDD.n17458 DVDD.n17457 0.00796421
R46589 DVDD.n17456 DVDD.n17331 0.00796421
R46590 DVDD.n17461 DVDD.n17460 0.00796421
R46591 DVDD.n17459 DVDD.n17330 0.00796421
R46592 DVDD.n17464 DVDD.n17463 0.00796421
R46593 DVDD.n17462 DVDD.n17329 0.00796421
R46594 DVDD.n17467 DVDD.n17466 0.00796421
R46595 DVDD.n17465 DVDD.n17328 0.00796421
R46596 DVDD.n17470 DVDD.n17469 0.00796421
R46597 DVDD.n17468 DVDD.n17327 0.00796421
R46598 DVDD.n17473 DVDD.n17472 0.00796421
R46599 DVDD.n17471 DVDD.n17326 0.00796421
R46600 DVDD.n17476 DVDD.n17475 0.00796421
R46601 DVDD.n17474 DVDD.n17325 0.00796421
R46602 DVDD.n17479 DVDD.n17478 0.00796421
R46603 DVDD.n17477 DVDD.n17324 0.00796421
R46604 DVDD.n17482 DVDD.n17481 0.00796421
R46605 DVDD.n17480 DVDD.n17323 0.00796421
R46606 DVDD.n17485 DVDD.n17484 0.00796421
R46607 DVDD.n17483 DVDD.n17322 0.00796421
R46608 DVDD.n17488 DVDD.n17487 0.00796421
R46609 DVDD.n17486 DVDD.n17321 0.00796421
R46610 DVDD.n17491 DVDD.n17490 0.00796421
R46611 DVDD.n17489 DVDD.n17320 0.00796421
R46612 DVDD.n17494 DVDD.n17493 0.00796421
R46613 DVDD.n17492 DVDD.n17319 0.00796421
R46614 DVDD.n17497 DVDD.n17496 0.00796421
R46615 DVDD.n17495 DVDD.n17318 0.00796421
R46616 DVDD.n17500 DVDD.n17499 0.00796421
R46617 DVDD.n17498 DVDD.n17317 0.00796421
R46618 DVDD.n17503 DVDD.n17502 0.00796421
R46619 DVDD.n17501 DVDD.n17316 0.00796421
R46620 DVDD.n17506 DVDD.n17505 0.00796421
R46621 DVDD.n17504 DVDD.n17315 0.00796421
R46622 DVDD.n17509 DVDD.n17508 0.00796421
R46623 DVDD.n17507 DVDD.n17314 0.00796421
R46624 DVDD.n17512 DVDD.n17511 0.00796421
R46625 DVDD.n17510 DVDD.n17313 0.00796421
R46626 DVDD.n17709 DVDD.n17514 0.00796421
R46627 DVDD.n17513 DVDD.n17312 0.00796421
R46628 DVDD.n5992 DVDD.n5937 0.00796421
R46629 DVDD.n17363 DVDD.n17362 0.00796421
R46630 DVDD.n5990 DVDD.n5989 0.00796421
R46631 DVDD.n17368 DVDD.n17365 0.00796421
R46632 DVDD.n5644 DVDD.n5590 0.00796421
R46633 DVDD.n15132 DVDD.n5591 0.00796421
R46634 DVDD.n5985 DVDD.n5645 0.00796421
R46635 DVDD.n5694 DVDD.n5640 0.00796421
R46636 DVDD.n5984 DVDD.n5646 0.00796421
R46637 DVDD.n5695 DVDD.n5639 0.00796421
R46638 DVDD.n5983 DVDD.n5647 0.00796421
R46639 DVDD.n5696 DVDD.n5638 0.00796421
R46640 DVDD.n5982 DVDD.n5648 0.00796421
R46641 DVDD.n5697 DVDD.n5637 0.00796421
R46642 DVDD.n5981 DVDD.n5649 0.00796421
R46643 DVDD.n5698 DVDD.n5636 0.00796421
R46644 DVDD.n5980 DVDD.n5650 0.00796421
R46645 DVDD.n5699 DVDD.n5635 0.00796421
R46646 DVDD.n5979 DVDD.n5651 0.00796421
R46647 DVDD.n5700 DVDD.n5634 0.00796421
R46648 DVDD.n5978 DVDD.n5652 0.00796421
R46649 DVDD.n5701 DVDD.n5633 0.00796421
R46650 DVDD.n5977 DVDD.n5653 0.00796421
R46651 DVDD.n5702 DVDD.n5632 0.00796421
R46652 DVDD.n5976 DVDD.n5654 0.00796421
R46653 DVDD.n5703 DVDD.n5631 0.00796421
R46654 DVDD.n5975 DVDD.n5655 0.00796421
R46655 DVDD.n5704 DVDD.n5630 0.00796421
R46656 DVDD.n5974 DVDD.n5656 0.00796421
R46657 DVDD.n5705 DVDD.n5629 0.00796421
R46658 DVDD.n5973 DVDD.n5657 0.00796421
R46659 DVDD.n5706 DVDD.n5628 0.00796421
R46660 DVDD.n5972 DVDD.n5658 0.00796421
R46661 DVDD.n5707 DVDD.n5627 0.00796421
R46662 DVDD.n5971 DVDD.n5659 0.00796421
R46663 DVDD.n5708 DVDD.n5626 0.00796421
R46664 DVDD.n5970 DVDD.n5660 0.00796421
R46665 DVDD.n5709 DVDD.n5625 0.00796421
R46666 DVDD.n5969 DVDD.n5661 0.00796421
R46667 DVDD.n5710 DVDD.n5624 0.00796421
R46668 DVDD.n5968 DVDD.n5662 0.00796421
R46669 DVDD.n5711 DVDD.n5623 0.00796421
R46670 DVDD.n5967 DVDD.n5663 0.00796421
R46671 DVDD.n5712 DVDD.n5622 0.00796421
R46672 DVDD.n5966 DVDD.n5664 0.00796421
R46673 DVDD.n5713 DVDD.n5621 0.00796421
R46674 DVDD.n5965 DVDD.n5665 0.00796421
R46675 DVDD.n5714 DVDD.n5620 0.00796421
R46676 DVDD.n5964 DVDD.n5666 0.00796421
R46677 DVDD.n5715 DVDD.n5619 0.00796421
R46678 DVDD.n5963 DVDD.n5667 0.00796421
R46679 DVDD.n5716 DVDD.n5618 0.00796421
R46680 DVDD.n5962 DVDD.n5668 0.00796421
R46681 DVDD.n5717 DVDD.n5617 0.00796421
R46682 DVDD.n5961 DVDD.n5669 0.00796421
R46683 DVDD.n5718 DVDD.n5616 0.00796421
R46684 DVDD.n5960 DVDD.n5670 0.00796421
R46685 DVDD.n5719 DVDD.n5615 0.00796421
R46686 DVDD.n5959 DVDD.n5671 0.00796421
R46687 DVDD.n5720 DVDD.n5614 0.00796421
R46688 DVDD.n5958 DVDD.n5672 0.00796421
R46689 DVDD.n5721 DVDD.n5613 0.00796421
R46690 DVDD.n5957 DVDD.n5673 0.00796421
R46691 DVDD.n5722 DVDD.n5612 0.00796421
R46692 DVDD.n5956 DVDD.n5674 0.00796421
R46693 DVDD.n5723 DVDD.n5611 0.00796421
R46694 DVDD.n5955 DVDD.n5675 0.00796421
R46695 DVDD.n5724 DVDD.n5610 0.00796421
R46696 DVDD.n5954 DVDD.n5676 0.00796421
R46697 DVDD.n5725 DVDD.n5609 0.00796421
R46698 DVDD.n5953 DVDD.n5677 0.00796421
R46699 DVDD.n5726 DVDD.n5608 0.00796421
R46700 DVDD.n5952 DVDD.n5678 0.00796421
R46701 DVDD.n5727 DVDD.n5607 0.00796421
R46702 DVDD.n5951 DVDD.n5679 0.00796421
R46703 DVDD.n5728 DVDD.n5606 0.00796421
R46704 DVDD.n5950 DVDD.n5680 0.00796421
R46705 DVDD.n5729 DVDD.n5605 0.00796421
R46706 DVDD.n5949 DVDD.n5681 0.00796421
R46707 DVDD.n5730 DVDD.n5604 0.00796421
R46708 DVDD.n5948 DVDD.n5682 0.00796421
R46709 DVDD.n5731 DVDD.n5603 0.00796421
R46710 DVDD.n5947 DVDD.n5683 0.00796421
R46711 DVDD.n5732 DVDD.n5602 0.00796421
R46712 DVDD.n5946 DVDD.n5684 0.00796421
R46713 DVDD.n5733 DVDD.n5601 0.00796421
R46714 DVDD.n5945 DVDD.n5685 0.00796421
R46715 DVDD.n5734 DVDD.n5600 0.00796421
R46716 DVDD.n5944 DVDD.n5686 0.00796421
R46717 DVDD.n5735 DVDD.n5599 0.00796421
R46718 DVDD.n5943 DVDD.n5687 0.00796421
R46719 DVDD.n5736 DVDD.n5598 0.00796421
R46720 DVDD.n5942 DVDD.n5688 0.00796421
R46721 DVDD.n5737 DVDD.n5597 0.00796421
R46722 DVDD.n5941 DVDD.n5689 0.00796421
R46723 DVDD.n5738 DVDD.n5596 0.00796421
R46724 DVDD.n5940 DVDD.n5690 0.00796421
R46725 DVDD.n5739 DVDD.n5595 0.00796421
R46726 DVDD.n5939 DVDD.n5691 0.00796421
R46727 DVDD.n5693 DVDD.n5594 0.00796421
R46728 DVDD.n17722 DVDD.n892 0.00796421
R46729 DVDD.n15137 DVDD.n5587 0.00796421
R46730 DVDD.n895 DVDD.n891 0.00796421
R46731 DVDD.n5581 DVDD.n5578 0.00796421
R46732 DVDD.n20038 DVDD.n19976 0.00795714
R46733 DVDD.n19865 DVDD.n19841 0.00795714
R46734 DVDD.n19160 DVDD.n19139 0.00795714
R46735 DVDD.n20929 DVDD.n18893 0.00795714
R46736 DVDD.n4029 DVDD.n242 0.00795714
R46737 DVDD.n22140 DVDD.n360 0.00795714
R46738 DVDD.n9920 DVDD.n9619 0.00795714
R46739 DVDD.n10057 DVDD.n9738 0.00795714
R46740 DVDD.n21184 DVDD.n21183 0.00795714
R46741 DVDD.n22297 DVDD.n22296 0.00795714
R46742 DVDD.n13770 DVDD.n11919 0.007925
R46743 DVDD.n16998 DVDD.n1709 0.007925
R46744 DVDD.n20138 DVDD.n20122 0.00789286
R46745 DVDD.n20136 DVDD.n20076 0.00789286
R46746 DVDD.n20625 DVDD.n20609 0.00789286
R46747 DVDD.n20623 DVDD.n20607 0.00789286
R46748 DVDD.n3976 DVDD.n3975 0.00789286
R46749 DVDD.n3972 DVDD.n3971 0.00789286
R46750 DVDD.n15285 DVDD.n5491 0.00789286
R46751 DVDD.n9838 DVDD.n5470 0.00789286
R46752 DVDD.n19648 DVDD.n19194 0.00789286
R46753 DVDD.n19646 DVDD.n19192 0.00789286
R46754 DVDD DVDD.n20334 0.00782857
R46755 DVDD.n20221 DVDD.n20026 0.00782857
R46756 DVDD.n20299 DVDD.n19844 0.00782857
R46757 DVDD.n20846 DVDD 0.00782857
R46758 DVDD.n20713 DVDD.n19144 0.00782857
R46759 DVDD.n20789 DVDD.n18873 0.00782857
R46760 DVDD.n22105 DVDD 0.00782857
R46761 DVDD.n4027 DVDD.n246 0.00782857
R46762 DVDD.n402 DVDD.n381 0.00782857
R46763 DVDD DVDD.n10015 0.00782857
R46764 DVDD.n9918 DVDD.n9622 0.00782857
R46765 DVDD.n9978 DVDD.n9957 0.00782857
R46766 DVDD.n21102 DVDD.n18738 0.00782857
R46767 DVDD.n81 DVDD.n59 0.00782857
R46768 DVDD.n22318 DVDD 0.00782857
R46769 DVDD.n20156 DVDD.n20072 0.00776429
R46770 DVDD.n20648 DVDD.n20647 0.00776429
R46771 DVDD.n3949 DVDD.n3925 0.00776429
R46772 DVDD.n9855 DVDD.n5474 0.00776429
R46773 DVDD.n19665 DVDD.n19188 0.00776429
R46774 DVDD.n11222 DVDD.n11105 0.00774832
R46775 DVDD.n16725 DVDD.n1814 0.00774832
R46776 DVDD.n11224 DVDD.n11223 0.00774832
R46777 DVDD.n16724 DVDD.n1815 0.00774832
R46778 DVDD.n21731 DVDD.n18430 0.00771783
R46779 DVDD.n22236 DVDD.n130 0.00771783
R46780 DVDD.n22067 DVDD.n18207 0.00771783
R46781 DVDD.n21936 DVDD.n21935 0.00771783
R46782 DVDD.n18100 DVDD.n18099 0.00771783
R46783 DVDD.n21944 DVDD.n18385 0.00770384
R46784 DVDD.n22209 DVDD.n179 0.00770384
R46785 DVDD.n20242 DVDD.n20031 0.0077
R46786 DVDD.n19859 DVDD.n19848 0.0077
R46787 DVDD.n20734 DVDD.n19149 0.0077
R46788 DVDD.n20805 DVDD.n18878 0.0077
R46789 DVDD.n22177 DVDD.n250 0.0077
R46790 DVDD.n393 DVDD.n386 0.0077
R46791 DVDD.n4761 DVDD.n4759 0.0077
R46792 DVDD.n9649 DVDD.n9625 0.0077
R46793 DVDD.n9969 DVDD.n9962 0.0077
R46794 DVDD.n21114 DVDD.n18742 0.0077
R46795 DVDD.n22273 DVDD.n63 0.0077
R46796 DVDD.n20337 DVDD.n18931 0.00763571
R46797 DVDD.n20851 DVDD.n18995 0.00763571
R46798 DVDD.n22116 DVDD.n22114 0.00763571
R46799 DVDD.n10020 DVDD.n790 0.00763571
R46800 DVDD.n20 DVDD.n1 0.00763571
R46801 DVDD.n20202 DVDD.n19725 0.00757143
R46802 DVDD.n19944 DVDD.n19886 0.00757143
R46803 DVDD.n20694 DVDD.n18832 0.00757143
R46804 DVDD.n20769 DVDD.n19036 0.00757143
R46805 DVDD.n4045 DVDD.n3863 0.00757143
R46806 DVDD.n22155 DVDD.n293 0.00757143
R46807 DVDD.n9939 DVDD.n9937 0.00757143
R46808 DVDD.n9723 DVDD.n9682 0.00757143
R46809 DVDD.n21196 DVDD.n18674 0.00757143
R46810 DVDD.n21128 DVDD.n107 0.00757143
R46811 DVDD.n14290 DVDD.n10237 0.00753759
R46812 DVDD.n17294 DVDD.n17293 0.00753759
R46813 DVDD.n20353 DVDD.n18935 0.00750714
R46814 DVDD.n20834 DVDD.n18964 0.00750714
R46815 DVDD.n22093 DVDD.n22074 0.00750714
R46816 DVDD.n10036 DVDD.n786 0.00750714
R46817 DVDD.n22327 DVDD.n15 0.00750714
R46818 DVDD.n21944 DVDD.n18378 0.00748725
R46819 DVDD.n22209 DVDD.n183 0.00748725
R46820 DVDD.n22229 DVDD.n138 0.00748725
R46821 DVDD.n22039 DVDD.n18244 0.00748725
R46822 DVDD.n21996 DVDD.n223 0.00748725
R46823 DVDD.n21336 DVDD.n18432 0.00748725
R46824 DVDD.n4858 DVDD.n3540 0.00748725
R46825 DVDD.n4859 DVDD.n3541 0.00748725
R46826 DVDD.n21849 DVDD.n21840 0.007475
R46827 DVDD.n18276 DVDD.n18274 0.007475
R46828 DVDD.n21238 DVDD.n21237 0.007475
R46829 DVDD.n21952 DVDD.n21951 0.007475
R46830 DVDD.n21819 DVDD.n21816 0.007475
R46831 DVDD.n18467 DVDD.n18464 0.007475
R46832 DVDD.n4303 DVDD.n4302 0.007475
R46833 DVDD.n3706 DVDD.n3694 0.007475
R46834 DVDD.n14009 DVDD.n11057 0.007475
R46835 DVDD.n17286 DVDD.n912 0.007475
R46836 DVDD.n20186 DVDD.n19729 0.00744286
R46837 DVDD.n20262 DVDD.n19890 0.00744286
R46838 DVDD.n20678 DVDD.n18836 0.00744286
R46839 DVDD.n19064 DVDD.n19040 0.00744286
R46840 DVDD.n4062 DVDD.n3867 0.00744286
R46841 DVDD.n335 DVDD.n297 0.00744286
R46842 DVDD.n9884 DVDD.n9761 0.00744286
R46843 DVDD.n9707 DVDD.n9686 0.00744286
R46844 DVDD.n18709 DVDD.n18681 0.00744286
R46845 DVDD.n21144 DVDD.n111 0.00744286
R46846 DVDD.n16452 DVDD.n1818 0.00740226
R46847 DVDD.n14851 DVDD.n7677 0.00737773
R46848 DVDD.n14852 DVDD.n7675 0.00737773
R46849 DVDD.n3670 DVDD.n3654 0.0073625
R46850 DVDD.n4546 DVDD.n4391 0.0073625
R46851 DVDD.n20175 DVDD.n19731 0.00731429
R46852 DVDD.n20667 DVDD.n18838 0.00731429
R46853 DVDD.n3987 DVDD.n3869 0.00731429
R46854 DVDD.n9873 DVDD.n9763 0.00731429
R46855 DVDD.n21213 DVDD.n18685 0.00731429
R46856 DVDD.n18078 DVDD.n18062 0.00730625
R46857 DVDD.n7062 DVDD.n6705 0.0072651
R46858 DVDD.n9562 DVDD.n7680 0.0072651
R46859 DVDD.n7063 DVDD.n6704 0.0072651
R46860 DVDD.n9563 DVDD.n7682 0.0072651
R46861 DVDD.n16256 DVDD.n2734 0.00726098
R46862 DVDD.n9785 DVDD.n3007 0.00726098
R46863 DVDD.n16247 DVDD.n2804 0.00726098
R46864 DVDD.n9781 DVDD.n2936 0.00726098
R46865 DVDD.n15988 DVDD.n3174 0.00726098
R46866 DVDD.n9779 DVDD.n9778 0.00726098
R46867 DVDD.n15533 DVDD.n15529 0.00726098
R46868 DVDD.n9782 DVDD.n3136 0.00726098
R46869 DVDD.n4753 DVDD.n4752 0.00725
R46870 DVDD.n4453 DVDD.n4450 0.00725
R46871 DVDD.n4449 DVDD.n4416 0.00725
R46872 DVDD.n4475 DVDD.n4399 0.00725
R46873 DVDD.n20191 DVDD.n19727 0.00718571
R46874 DVDD.n20266 DVDD.n19888 0.00718571
R46875 DVDD.n20683 DVDD.n18834 0.00718571
R46876 DVDD.n20758 DVDD.n19038 0.00718571
R46877 DVDD.n4056 DVDD.n3865 0.00718571
R46878 DVDD.n329 DVDD.n295 0.00718571
R46879 DVDD.n9820 DVDD.n9759 0.00718571
R46880 DVDD.n9704 DVDD.n9684 0.00718571
R46881 DVDD.n18711 DVDD.n18678 0.00718571
R46882 DVDD.n21126 DVDD.n109 0.00718571
R46883 DVDD.n4425 DVDD.n3748 0.0071375
R46884 DVDD.n4280 DVDD.n4241 0.0071375
R46885 DVDD.n18134 DVDD.n18133 0.0071375
R46886 DVDD.n18132 DVDD.n490 0.0071375
R46887 DVDD.n20348 DVDD.n18933 0.00712143
R46888 DVDD.n19000 DVDD.n18962 0.00712143
R46889 DVDD.n22090 DVDD.n22072 0.00712143
R46890 DVDD.n10031 DVDD.n788 0.00712143
R46891 DVDD.n22313 DVDD.n17 0.00712143
R46892 DVDD.n21714 DVDD.n18512 0.0071
R46893 DVDD.n21659 DVDD.n18542 0.0071
R46894 DVDD.n22218 DVDD.n170 0.0071
R46895 DVDD.n21743 DVDD.n21742 0.0071
R46896 DVDD.n3607 DVDD.n3530 0.00708125
R46897 DVDD.n20282 DVDD.n19873 0.00705714
R46898 DVDD.n20420 DVDD.n20371 0.00705714
R46899 DVDD.n20776 DVDD.n19057 0.00705714
R46900 DVDD.n20816 DVDD.n18876 0.00705714
R46901 DVDD.n22149 DVDD.n320 0.00705714
R46902 DVDD.n22138 DVDD.n22137 0.00705714
R46903 DVDD.n9727 DVDD.n9680 0.00705714
R46904 DVDD.n10055 DVDD.n10054 0.00705714
R46905 DVDD.n22254 DVDD.n22253 0.00705714
R46906 DVDD.n22299 DVDD.n38 0.00705714
R46907 DVDD.n4741 DVDD.n4740 0.007025
R46908 DVDD.n4315 DVDD.n4244 0.007025
R46909 DVDD.n15127 DVDD.n15125 0.007025
R46910 DVDD.n15066 DVDD.n7052 0.007025
R46911 DVDD.n12378 DVDD.n12377 0.00699624
R46912 DVDD.n12892 DVDD.n12384 0.00699624
R46913 DVDD.n11632 DVDD.n11579 0.00698472
R46914 DVDD.n16996 DVDD.n1711 0.00698472
R46915 DVDD.n11922 DVDD.n11921 0.00698472
R46916 DVDD.n16997 DVDD.n1710 0.00698472
R46917 DVDD.n21944 DVDD.n18297 0.00693543
R46918 DVDD.n22229 DVDD.n155 0.00693543
R46919 DVDD.n21723 DVDD.n18432 0.00693543
R46920 DVDD.n22041 DVDD.n22039 0.00693543
R46921 DVDD.n22040 DVDD.n223 0.00693543
R46922 DVDD.n22209 DVDD.n180 0.00693543
R46923 DVDD.n18115 DVDD.n18114 0.00693543
R46924 DVDD.n18116 DVDD.n18092 0.00693543
R46925 DVDD.n20232 DVDD.n20028 0.00692857
R46926 DVDD.n20310 DVDD.n19846 0.00692857
R46927 DVDD.n20724 DVDD.n19146 0.00692857
R46928 DVDD.n19013 DVDD.n18875 0.00692857
R46929 DVDD.n4014 DVDD.n248 0.00692857
R46930 DVDD.n413 DVDD.n383 0.00692857
R46931 DVDD.n9643 DVDD.n9624 0.00692857
R46932 DVDD.n9989 DVDD.n9959 0.00692857
R46933 DVDD.n21169 DVDD.n18740 0.00692857
R46934 DVDD.n22282 DVDD.n61 0.00692857
R46935 DVDD.n20152 DVDD.n20074 0.00686429
R46936 DVDD.n20639 DVDD.n20605 0.00686429
R46937 DVDD.n3943 DVDD.n3923 0.00686429
R46938 DVDD.n9851 DVDD.n5472 0.00686429
R46939 DVDD.n19644 DVDD.n19190 0.00686429
R46940 DVDD.n3609 DVDD.n3525 0.00685625
R46941 DVDD.n20216 DVDD.n20023 0.0068
R46942 DVDD.n20708 DVDD.n19141 0.0068
R46943 DVDD.n4031 DVDD.n244 0.0068
R46944 DVDD.n4442 DVDD.n3739 0.0068
R46945 DVDD.n4600 DVDD.n4252 0.0068
R46946 DVDD.n4572 DVDD.n4282 0.0068
R46947 DVDD.n4574 DVDD.n4573 0.0068
R46948 DVDD.n9922 DVDD.n9621 0.0068
R46949 DVDD.n21100 DVDD.n18736 0.0068
R46950 DVDD.n14292 DVDD.n8611 0.00678188
R46951 DVDD.n17291 DVDD.n916 0.00678188
R46952 DVDD.n14291 DVDD.n8613 0.00678188
R46953 DVDD.n17292 DVDD.n917 0.00678188
R46954 DVDD.n22201 DVDD.n22200 0.00678
R46955 DVDD.n18360 DVDD.n18359 0.00678
R46956 DVDD.n21890 DVDD.n21834 0.00678
R46957 DVDD.n21905 DVDD.n21806 0.00678
R46958 DVDD.n20143 DVDD.n20125 0.00673571
R46959 DVDD.n20630 DVDD.n20612 0.00673571
R46960 DVDD.n3966 DVDD.n3932 0.00673571
R46961 DVDD.n9842 DVDD.n5483 0.00673571
R46962 DVDD.n19653 DVDD.n19196 0.00673571
R46963 DVDD.n3712 DVDD.n3711 0.0066875
R46964 DVDD.n4477 DVDD.n4202 0.0066875
R46965 DVDD.n4534 DVDD.n4478 0.0066875
R46966 DVDD.n20223 DVDD.n19974 0.00667143
R46967 DVDD.n20301 DVDD.n19839 0.00667143
R46968 DVDD.n20715 DVDD.n19137 0.00667143
R46969 DVDD.n19016 DVDD.n18885 0.00667143
R46970 DVDD.n4011 DVDD.n240 0.00667143
R46971 DVDD.n404 DVDD.n377 0.00667143
R46972 DVDD.n9905 DVDD.n9617 0.00667143
R46973 DVDD.n9980 DVDD.n9754 0.00667143
R46974 DVDD.n21177 DVDD.n21097 0.00667143
R46975 DVDD.n22290 DVDD.n76 0.00667143
R46976 DVDD.n18074 DVDD.n18058 0.00663125
R46977 DVDD.n20163 DVDD.n20130 0.00660714
R46978 DVDD.n20655 DVDD.n20617 0.00660714
R46979 DVDD.n3947 DVDD.n3927 0.00660714
R46980 DVDD.n9831 DVDD.n5478 0.00660714
R46981 DVDD.n19638 DVDD.n19200 0.00660714
R46982 DVDD.n14011 DVDD.n10712 0.0065917
R46983 DVDD.n17288 DVDD.n914 0.0065917
R46984 DVDD.n14010 DVDD.n10714 0.0065917
R46985 DVDD.n17287 DVDD.n913 0.0065917
R46986 DVDD.n19652 DVDD.n19651 0.00658571
R46987 DVDD.n19652 DVDD.n19645 0.00658571
R46988 DVDD.n19659 DVDD.n19645 0.00658571
R46989 DVDD.n19660 DVDD.n19659 0.00658571
R46990 DVDD.n19661 DVDD.n19660 0.00658571
R46991 DVDD.n19661 DVDD.n19641 0.00658571
R46992 DVDD.n19667 DVDD.n19641 0.00658571
R46993 DVDD.n19668 DVDD.n19667 0.00658571
R46994 DVDD.n19694 DVDD.n19668 0.00658571
R46995 DVDD.n19694 DVDD.n19693 0.00658571
R46996 DVDD.n19693 DVDD.n19692 0.00658571
R46997 DVDD.n19692 DVDD.n19669 0.00658571
R46998 DVDD.n19672 DVDD.n19669 0.00658571
R46999 DVDD.n19685 DVDD.n19672 0.00658571
R47000 DVDD.n19685 DVDD.n19684 0.00658571
R47001 DVDD.n19684 DVDD.n19683 0.00658571
R47002 DVDD.n19683 DVDD.n19673 0.00658571
R47003 DVDD.n19678 DVDD.n19673 0.00658571
R47004 DVDD.n19678 DVDD.n19677 0.00658571
R47005 DVDD.n19677 DVDD.n18713 0.00658571
R47006 DVDD.n21208 DVDD.n18713 0.00658571
R47007 DVDD.n21208 DVDD.n21207 0.00658571
R47008 DVDD.n21207 DVDD.n21206 0.00658571
R47009 DVDD.n21206 DVDD.n18714 0.00658571
R47010 DVDD.n21200 DVDD.n18714 0.00658571
R47011 DVDD.n21200 DVDD.n21199 0.00658571
R47012 DVDD.n21199 DVDD.n21198 0.00658571
R47013 DVDD.n21198 DVDD.n18718 0.00658571
R47014 DVDD.n21192 DVDD.n18718 0.00658571
R47015 DVDD.n21192 DVDD.n21191 0.00658571
R47016 DVDD.n21191 DVDD.n21190 0.00658571
R47017 DVDD.n21190 DVDD.n18721 0.00658571
R47018 DVDD.n21105 DVDD.n18721 0.00658571
R47019 DVDD.n21106 DVDD.n21105 0.00658571
R47020 DVDD.n21181 DVDD.n21106 0.00658571
R47021 DVDD.n21181 DVDD.n21180 0.00658571
R47022 DVDD.n21180 DVDD.n21179 0.00658571
R47023 DVDD.n21179 DVDD.n21107 0.00658571
R47024 DVDD.n21173 DVDD.n21107 0.00658571
R47025 DVDD.n21173 DVDD.n21172 0.00658571
R47026 DVDD.n21172 DVDD.n21171 0.00658571
R47027 DVDD.n21171 DVDD.n21111 0.00658571
R47028 DVDD.n21165 DVDD.n21111 0.00658571
R47029 DVDD.n21165 DVDD.n21164 0.00658571
R47030 DVDD.n21164 DVDD.n21163 0.00658571
R47031 DVDD.n21163 DVDD.n21115 0.00658571
R47032 DVDD.n21119 DVDD.n21115 0.00658571
R47033 DVDD.n21155 DVDD.n21119 0.00658571
R47034 DVDD.n21155 DVDD.n21154 0.00658571
R47035 DVDD.n21154 DVDD.n21153 0.00658571
R47036 DVDD.n21153 DVDD.n21120 0.00658571
R47037 DVDD.n21148 DVDD.n21120 0.00658571
R47038 DVDD.n21148 DVDD.n21147 0.00658571
R47039 DVDD.n21147 DVDD.n21146 0.00658571
R47040 DVDD.n21146 DVDD.n21123 0.00658571
R47041 DVDD.n21140 DVDD.n21123 0.00658571
R47042 DVDD.n21140 DVDD.n21139 0.00658571
R47043 DVDD.n21139 DVDD.n21138 0.00658571
R47044 DVDD.n21138 DVDD.n21127 0.00658571
R47045 DVDD.n21132 DVDD.n21127 0.00658571
R47046 DVDD.n21132 DVDD.n21131 0.00658571
R47047 DVDD.n21131 DVDD.n87 0.00658571
R47048 DVDD.n22256 DVDD.n87 0.00658571
R47049 DVDD.n22257 DVDD.n22256 0.00658571
R47050 DVDD.n22258 DVDD.n22257 0.00658571
R47051 DVDD.n22258 DVDD.n83 0.00658571
R47052 DVDD.n22264 DVDD.n83 0.00658571
R47053 DVDD.n22265 DVDD.n22264 0.00658571
R47054 DVDD.n22294 DVDD.n22265 0.00658571
R47055 DVDD.n22294 DVDD.n22293 0.00658571
R47056 DVDD.n22293 DVDD.n22292 0.00658571
R47057 DVDD.n22292 DVDD.n22266 0.00658571
R47058 DVDD.n22286 DVDD.n22266 0.00658571
R47059 DVDD.n22286 DVDD.n22285 0.00658571
R47060 DVDD.n22285 DVDD.n22284 0.00658571
R47061 DVDD.n22284 DVDD.n22270 0.00658571
R47062 DVDD.n22278 DVDD.n22270 0.00658571
R47063 DVDD.n22278 DVDD.n22277 0.00658571
R47064 DVDD.n22277 DVDD.n22276 0.00658571
R47065 DVDD.n22276 DVDD.n40 0.00658571
R47066 DVDD.n22302 DVDD.n40 0.00658571
R47067 DVDD.n22303 DVDD.n22302 0.00658571
R47068 DVDD.n22304 DVDD.n22303 0.00658571
R47069 DVDD.n22304 DVDD.n36 0.00658571
R47070 DVDD.n22310 DVDD.n36 0.00658571
R47071 DVDD.n22311 DVDD.n22310 0.00658571
R47072 DVDD.n22333 DVDD.n22311 0.00658571
R47073 DVDD.n22333 DVDD.n22332 0.00658571
R47074 DVDD.n22332 DVDD.n22331 0.00658571
R47075 DVDD.n22331 DVDD.n22312 0.00658571
R47076 DVDD.n22325 DVDD.n22312 0.00658571
R47077 DVDD.n22325 DVDD.n22324 0.00658571
R47078 DVDD.n22324 DVDD.n22323 0.00658571
R47079 DVDD.n22323 DVDD.n22316 0.00658571
R47080 DVDD.n22316 DVDD.n3 0.00658571
R47081 DVDD.n22349 DVDD.n3 0.00658571
R47082 DVDD.n20142 DVDD.n20141 0.00658571
R47083 DVDD.n20142 DVDD.n20135 0.00658571
R47084 DVDD.n20149 DVDD.n20135 0.00658571
R47085 DVDD.n20150 DVDD.n20149 0.00658571
R47086 DVDD.n20151 DVDD.n20150 0.00658571
R47087 DVDD.n20151 DVDD.n20132 0.00658571
R47088 DVDD.n20158 DVDD.n20132 0.00658571
R47089 DVDD.n20159 DVDD.n20158 0.00658571
R47090 DVDD.n20160 DVDD.n20159 0.00658571
R47091 DVDD.n20160 DVDD.n20057 0.00658571
R47092 DVDD.n20168 DVDD.n20057 0.00658571
R47093 DVDD.n20169 DVDD.n20168 0.00658571
R47094 DVDD.n20171 DVDD.n20169 0.00658571
R47095 DVDD.n20171 DVDD.n20170 0.00658571
R47096 DVDD.n20170 DVDD.n20053 0.00658571
R47097 DVDD.n20179 DVDD.n20053 0.00658571
R47098 DVDD.n20180 DVDD.n20179 0.00658571
R47099 DVDD.n20181 DVDD.n20180 0.00658571
R47100 DVDD.n20181 DVDD.n20050 0.00658571
R47101 DVDD.n20188 DVDD.n20050 0.00658571
R47102 DVDD.n20189 DVDD.n20188 0.00658571
R47103 DVDD.n20190 DVDD.n20189 0.00658571
R47104 DVDD.n20190 DVDD.n20047 0.00658571
R47105 DVDD.n20197 DVDD.n20047 0.00658571
R47106 DVDD.n20198 DVDD.n20197 0.00658571
R47107 DVDD.n20199 DVDD.n20198 0.00658571
R47108 DVDD.n20199 DVDD.n20044 0.00658571
R47109 DVDD.n20205 DVDD.n20044 0.00658571
R47110 DVDD.n20206 DVDD.n20205 0.00658571
R47111 DVDD.n20208 DVDD.n20206 0.00658571
R47112 DVDD.n20208 DVDD.n20207 0.00658571
R47113 DVDD.n20207 DVDD.n20042 0.00658571
R47114 DVDD.n20042 DVDD.n20040 0.00658571
R47115 DVDD.n20218 DVDD.n20040 0.00658571
R47116 DVDD.n20219 DVDD.n20218 0.00658571
R47117 DVDD.n20220 DVDD.n20219 0.00658571
R47118 DVDD.n20220 DVDD.n20037 0.00658571
R47119 DVDD.n20227 DVDD.n20037 0.00658571
R47120 DVDD.n20228 DVDD.n20227 0.00658571
R47121 DVDD.n20229 DVDD.n20228 0.00658571
R47122 DVDD.n20229 DVDD.n20034 0.00658571
R47123 DVDD.n20236 DVDD.n20034 0.00658571
R47124 DVDD.n20237 DVDD.n20236 0.00658571
R47125 DVDD.n20239 DVDD.n20237 0.00658571
R47126 DVDD.n20239 DVDD.n20238 0.00658571
R47127 DVDD.n20238 DVDD.n19956 0.00658571
R47128 DVDD.n20248 DVDD.n19956 0.00658571
R47129 DVDD.n20249 DVDD.n20248 0.00658571
R47130 DVDD.n20251 DVDD.n20249 0.00658571
R47131 DVDD.n20251 DVDD.n20250 0.00658571
R47132 DVDD.n20250 DVDD.n19952 0.00658571
R47133 DVDD.n20259 DVDD.n19952 0.00658571
R47134 DVDD.n20260 DVDD.n20259 0.00658571
R47135 DVDD.n20261 DVDD.n20260 0.00658571
R47136 DVDD.n20261 DVDD.n19949 0.00658571
R47137 DVDD.n20268 DVDD.n19949 0.00658571
R47138 DVDD.n20269 DVDD.n20268 0.00658571
R47139 DVDD.n20270 DVDD.n20269 0.00658571
R47140 DVDD.n20270 DVDD.n19946 0.00658571
R47141 DVDD.n20277 DVDD.n19946 0.00658571
R47142 DVDD.n20278 DVDD.n20277 0.00658571
R47143 DVDD.n20279 DVDD.n20278 0.00658571
R47144 DVDD.n20279 DVDD.n19871 0.00658571
R47145 DVDD.n20288 DVDD.n19871 0.00658571
R47146 DVDD.n20289 DVDD.n20288 0.00658571
R47147 DVDD.n20290 DVDD.n20289 0.00658571
R47148 DVDD.n20290 DVDD.n19867 0.00658571
R47149 DVDD.n20296 DVDD.n19867 0.00658571
R47150 DVDD.n20297 DVDD.n20296 0.00658571
R47151 DVDD.n20298 DVDD.n20297 0.00658571
R47152 DVDD.n20298 DVDD.n19864 0.00658571
R47153 DVDD.n20305 DVDD.n19864 0.00658571
R47154 DVDD.n20306 DVDD.n20305 0.00658571
R47155 DVDD.n20307 DVDD.n20306 0.00658571
R47156 DVDD.n20307 DVDD.n19861 0.00658571
R47157 DVDD.n20314 DVDD.n19861 0.00658571
R47158 DVDD.n20315 DVDD.n20314 0.00658571
R47159 DVDD.n20316 DVDD.n20315 0.00658571
R47160 DVDD.n20316 DVDD.n19858 0.00658571
R47161 DVDD.n20323 DVDD.n19858 0.00658571
R47162 DVDD.n20324 DVDD.n20323 0.00658571
R47163 DVDD.n20369 DVDD.n20324 0.00658571
R47164 DVDD.n20369 DVDD.n20368 0.00658571
R47165 DVDD.n20368 DVDD.n20367 0.00658571
R47166 DVDD.n20367 DVDD.n20325 0.00658571
R47167 DVDD.n20361 DVDD.n20325 0.00658571
R47168 DVDD.n20361 DVDD.n20360 0.00658571
R47169 DVDD.n20360 DVDD.n20359 0.00658571
R47170 DVDD.n20359 DVDD.n20329 0.00658571
R47171 DVDD.n20352 DVDD.n20329 0.00658571
R47172 DVDD.n20352 DVDD.n20351 0.00658571
R47173 DVDD.n20351 DVDD.n20350 0.00658571
R47174 DVDD.n20350 DVDD.n20332 0.00658571
R47175 DVDD.n20343 DVDD.n20332 0.00658571
R47176 DVDD.n20343 DVDD.n20342 0.00658571
R47177 DVDD.n20342 DVDD.n20341 0.00658571
R47178 DVDD.n20629 DVDD.n20628 0.00658571
R47179 DVDD.n20629 DVDD.n20622 0.00658571
R47180 DVDD.n20636 DVDD.n20622 0.00658571
R47181 DVDD.n20637 DVDD.n20636 0.00658571
R47182 DVDD.n20638 DVDD.n20637 0.00658571
R47183 DVDD.n20638 DVDD.n20619 0.00658571
R47184 DVDD.n20650 DVDD.n20619 0.00658571
R47185 DVDD.n20651 DVDD.n20650 0.00658571
R47186 DVDD.n20652 DVDD.n20651 0.00658571
R47187 DVDD.n20652 DVDD.n19179 0.00658571
R47188 DVDD.n20660 DVDD.n19179 0.00658571
R47189 DVDD.n20661 DVDD.n20660 0.00658571
R47190 DVDD.n20663 DVDD.n20661 0.00658571
R47191 DVDD.n20663 DVDD.n20662 0.00658571
R47192 DVDD.n20662 DVDD.n19175 0.00658571
R47193 DVDD.n20671 DVDD.n19175 0.00658571
R47194 DVDD.n20672 DVDD.n20671 0.00658571
R47195 DVDD.n20673 DVDD.n20672 0.00658571
R47196 DVDD.n20673 DVDD.n19172 0.00658571
R47197 DVDD.n20680 DVDD.n19172 0.00658571
R47198 DVDD.n20681 DVDD.n20680 0.00658571
R47199 DVDD.n20682 DVDD.n20681 0.00658571
R47200 DVDD.n20682 DVDD.n19169 0.00658571
R47201 DVDD.n20689 DVDD.n19169 0.00658571
R47202 DVDD.n20690 DVDD.n20689 0.00658571
R47203 DVDD.n20691 DVDD.n20690 0.00658571
R47204 DVDD.n20691 DVDD.n19166 0.00658571
R47205 DVDD.n20697 DVDD.n19166 0.00658571
R47206 DVDD.n20698 DVDD.n20697 0.00658571
R47207 DVDD.n20700 DVDD.n20698 0.00658571
R47208 DVDD.n20700 DVDD.n20699 0.00658571
R47209 DVDD.n20699 DVDD.n19164 0.00658571
R47210 DVDD.n19164 DVDD.n19162 0.00658571
R47211 DVDD.n20710 DVDD.n19162 0.00658571
R47212 DVDD.n20711 DVDD.n20710 0.00658571
R47213 DVDD.n20712 DVDD.n20711 0.00658571
R47214 DVDD.n20712 DVDD.n19159 0.00658571
R47215 DVDD.n20719 DVDD.n19159 0.00658571
R47216 DVDD.n20720 DVDD.n20719 0.00658571
R47217 DVDD.n20721 DVDD.n20720 0.00658571
R47218 DVDD.n20721 DVDD.n19156 0.00658571
R47219 DVDD.n20728 DVDD.n19156 0.00658571
R47220 DVDD.n20729 DVDD.n20728 0.00658571
R47221 DVDD.n20731 DVDD.n20729 0.00658571
R47222 DVDD.n20731 DVDD.n20730 0.00658571
R47223 DVDD.n20730 DVDD.n19071 0.00658571
R47224 DVDD.n20740 DVDD.n19071 0.00658571
R47225 DVDD.n20741 DVDD.n20740 0.00658571
R47226 DVDD.n20743 DVDD.n20741 0.00658571
R47227 DVDD.n20743 DVDD.n20742 0.00658571
R47228 DVDD.n20742 DVDD.n19068 0.00658571
R47229 DVDD.n19068 DVDD.n19066 0.00658571
R47230 DVDD.n20753 DVDD.n19066 0.00658571
R47231 DVDD.n20754 DVDD.n20753 0.00658571
R47232 DVDD.n20755 DVDD.n20754 0.00658571
R47233 DVDD.n20755 DVDD.n19063 0.00658571
R47234 DVDD.n20762 DVDD.n19063 0.00658571
R47235 DVDD.n20763 DVDD.n20762 0.00658571
R47236 DVDD.n20764 DVDD.n20763 0.00658571
R47237 DVDD.n20764 DVDD.n19060 0.00658571
R47238 DVDD.n20771 DVDD.n19060 0.00658571
R47239 DVDD.n20772 DVDD.n20771 0.00658571
R47240 DVDD.n20774 DVDD.n20772 0.00658571
R47241 DVDD.n20774 DVDD.n20773 0.00658571
R47242 DVDD.n20773 DVDD.n19020 0.00658571
R47243 DVDD.n20784 DVDD.n19020 0.00658571
R47244 DVDD.n20785 DVDD.n20784 0.00658571
R47245 DVDD.n20786 DVDD.n20785 0.00658571
R47246 DVDD.n20786 DVDD.n19018 0.00658571
R47247 DVDD.n20791 DVDD.n19018 0.00658571
R47248 DVDD.n20792 DVDD.n20791 0.00658571
R47249 DVDD.n20793 DVDD.n20792 0.00658571
R47250 DVDD.n20793 DVDD.n19015 0.00658571
R47251 DVDD.n20800 DVDD.n19015 0.00658571
R47252 DVDD.n20801 DVDD.n20800 0.00658571
R47253 DVDD.n20802 DVDD.n20801 0.00658571
R47254 DVDD.n20802 DVDD.n19012 0.00658571
R47255 DVDD.n20809 DVDD.n19012 0.00658571
R47256 DVDD.n20810 DVDD.n20809 0.00658571
R47257 DVDD.n20811 DVDD.n20810 0.00658571
R47258 DVDD.n20811 DVDD.n19009 0.00658571
R47259 DVDD.n20818 DVDD.n19009 0.00658571
R47260 DVDD.n20819 DVDD.n20818 0.00658571
R47261 DVDD.n20821 DVDD.n20819 0.00658571
R47262 DVDD.n20821 DVDD.n20820 0.00658571
R47263 DVDD.n20820 DVDD.n19005 0.00658571
R47264 DVDD.n20829 DVDD.n19005 0.00658571
R47265 DVDD.n20830 DVDD.n20829 0.00658571
R47266 DVDD.n20831 DVDD.n20830 0.00658571
R47267 DVDD.n20831 DVDD.n19002 0.00658571
R47268 DVDD.n20838 DVDD.n19002 0.00658571
R47269 DVDD.n20839 DVDD.n20838 0.00658571
R47270 DVDD.n20840 DVDD.n20839 0.00658571
R47271 DVDD.n20840 DVDD.n18999 0.00658571
R47272 DVDD.n20847 DVDD.n18999 0.00658571
R47273 DVDD.n20848 DVDD.n20847 0.00658571
R47274 DVDD.n3964 DVDD.n3963 0.00658571
R47275 DVDD.n3963 DVDD.n3962 0.00658571
R47276 DVDD.n3962 DVDD.n3942 0.00658571
R47277 DVDD.n3955 DVDD.n3942 0.00658571
R47278 DVDD.n3955 DVDD.n3954 0.00658571
R47279 DVDD.n3954 DVDD.n3953 0.00658571
R47280 DVDD.n3953 DVDD.n3945 0.00658571
R47281 DVDD.n3946 DVDD.n3945 0.00658571
R47282 DVDD.n3946 DVDD.n3908 0.00658571
R47283 DVDD.n3981 DVDD.n3908 0.00658571
R47284 DVDD.n3982 DVDD.n3981 0.00658571
R47285 DVDD.n3983 DVDD.n3982 0.00658571
R47286 DVDD.n3983 DVDD.n3904 0.00658571
R47287 DVDD.n3990 DVDD.n3904 0.00658571
R47288 DVDD.n3991 DVDD.n3990 0.00658571
R47289 DVDD.n3992 DVDD.n3991 0.00658571
R47290 DVDD.n3992 DVDD.n3902 0.00658571
R47291 DVDD.n3999 DVDD.n3902 0.00658571
R47292 DVDD.n4000 DVDD.n3999 0.00658571
R47293 DVDD.n4060 DVDD.n4000 0.00658571
R47294 DVDD.n4060 DVDD.n4059 0.00658571
R47295 DVDD.n4059 DVDD.n4058 0.00658571
R47296 DVDD.n4058 DVDD.n4001 0.00658571
R47297 DVDD.n4051 DVDD.n4001 0.00658571
R47298 DVDD.n4051 DVDD.n4050 0.00658571
R47299 DVDD.n4050 DVDD.n4049 0.00658571
R47300 DVDD.n4049 DVDD.n4004 0.00658571
R47301 DVDD.n4043 DVDD.n4004 0.00658571
R47302 DVDD.n4043 DVDD.n4042 0.00658571
R47303 DVDD.n4042 DVDD.n4041 0.00658571
R47304 DVDD.n4041 DVDD.n4006 0.00658571
R47305 DVDD.n4035 DVDD.n4006 0.00658571
R47306 DVDD.n4035 DVDD.n4034 0.00658571
R47307 DVDD.n4034 DVDD.n4033 0.00658571
R47308 DVDD.n4033 DVDD.n4010 0.00658571
R47309 DVDD.n4026 DVDD.n4010 0.00658571
R47310 DVDD.n4026 DVDD.n4025 0.00658571
R47311 DVDD.n4025 DVDD.n4024 0.00658571
R47312 DVDD.n4024 DVDD.n4013 0.00658571
R47313 DVDD.n4017 DVDD.n4013 0.00658571
R47314 DVDD.n4017 DVDD.n4016 0.00658571
R47315 DVDD.n4016 DVDD.n276 0.00658571
R47316 DVDD.n22175 DVDD.n276 0.00658571
R47317 DVDD.n22175 DVDD.n22174 0.00658571
R47318 DVDD.n22174 DVDD.n22173 0.00658571
R47319 DVDD.n22173 DVDD.n277 0.00658571
R47320 DVDD.n279 DVDD.n277 0.00658571
R47321 DVDD.n282 DVDD.n279 0.00658571
R47322 DVDD.n22165 DVDD.n282 0.00658571
R47323 DVDD.n22165 DVDD.n22164 0.00658571
R47324 DVDD.n22164 DVDD.n22163 0.00658571
R47325 DVDD.n22163 DVDD.n283 0.00658571
R47326 DVDD.n332 DVDD.n283 0.00658571
R47327 DVDD.n332 DVDD.n331 0.00658571
R47328 DVDD.n339 DVDD.n331 0.00658571
R47329 DVDD.n340 DVDD.n339 0.00658571
R47330 DVDD.n341 DVDD.n340 0.00658571
R47331 DVDD.n341 DVDD.n328 0.00658571
R47332 DVDD.n348 DVDD.n328 0.00658571
R47333 DVDD.n349 DVDD.n348 0.00658571
R47334 DVDD.n22153 DVDD.n349 0.00658571
R47335 DVDD.n22153 DVDD.n22152 0.00658571
R47336 DVDD.n22152 DVDD.n22151 0.00658571
R47337 DVDD.n22151 DVDD.n350 0.00658571
R47338 DVDD.n22146 DVDD.n350 0.00658571
R47339 DVDD.n22146 DVDD.n22145 0.00658571
R47340 DVDD.n22145 DVDD.n22144 0.00658571
R47341 DVDD.n22144 DVDD.n352 0.00658571
R47342 DVDD.n400 DVDD.n352 0.00658571
R47343 DVDD.n401 DVDD.n400 0.00658571
R47344 DVDD.n401 DVDD.n398 0.00658571
R47345 DVDD.n408 DVDD.n398 0.00658571
R47346 DVDD.n409 DVDD.n408 0.00658571
R47347 DVDD.n410 DVDD.n409 0.00658571
R47348 DVDD.n410 DVDD.n395 0.00658571
R47349 DVDD.n417 DVDD.n395 0.00658571
R47350 DVDD.n418 DVDD.n417 0.00658571
R47351 DVDD.n419 DVDD.n418 0.00658571
R47352 DVDD.n419 DVDD.n392 0.00658571
R47353 DVDD.n431 DVDD.n392 0.00658571
R47354 DVDD.n432 DVDD.n431 0.00658571
R47355 DVDD.n22135 DVDD.n432 0.00658571
R47356 DVDD.n22135 DVDD.n22134 0.00658571
R47357 DVDD.n22134 DVDD.n22133 0.00658571
R47358 DVDD.n22133 DVDD.n433 0.00658571
R47359 DVDD.n22127 DVDD.n433 0.00658571
R47360 DVDD.n22127 DVDD.n22126 0.00658571
R47361 DVDD.n22126 DVDD.n22125 0.00658571
R47362 DVDD.n22125 DVDD.n437 0.00658571
R47363 DVDD.n22092 DVDD.n437 0.00658571
R47364 DVDD.n22097 DVDD.n22092 0.00658571
R47365 DVDD.n22098 DVDD.n22097 0.00658571
R47366 DVDD.n22099 DVDD.n22098 0.00658571
R47367 DVDD.n22099 DVDD.n22089 0.00658571
R47368 DVDD.n22106 DVDD.n22089 0.00658571
R47369 DVDD.n22107 DVDD.n22106 0.00658571
R47370 DVDD.n9841 DVDD.n9840 0.00658571
R47371 DVDD.n9841 DVDD.n9836 0.00658571
R47372 DVDD.n9848 DVDD.n9836 0.00658571
R47373 DVDD.n9849 DVDD.n9848 0.00658571
R47374 DVDD.n9850 DVDD.n9849 0.00658571
R47375 DVDD.n9850 DVDD.n9833 0.00658571
R47376 DVDD.n9857 DVDD.n9833 0.00658571
R47377 DVDD.n9858 DVDD.n9857 0.00658571
R47378 DVDD.n9859 DVDD.n9858 0.00658571
R47379 DVDD.n9859 DVDD.n9830 0.00658571
R47380 DVDD.n9866 DVDD.n9830 0.00658571
R47381 DVDD.n9867 DVDD.n9866 0.00658571
R47382 DVDD.n9869 DVDD.n9867 0.00658571
R47383 DVDD.n9869 DVDD.n9868 0.00658571
R47384 DVDD.n9868 DVDD.n9827 0.00658571
R47385 DVDD.n9827 DVDD.n9825 0.00658571
R47386 DVDD.n9879 DVDD.n9825 0.00658571
R47387 DVDD.n9880 DVDD.n9879 0.00658571
R47388 DVDD.n9881 DVDD.n9880 0.00658571
R47389 DVDD.n9881 DVDD.n9822 0.00658571
R47390 DVDD.n9888 DVDD.n9822 0.00658571
R47391 DVDD.n9889 DVDD.n9888 0.00658571
R47392 DVDD.n9890 DVDD.n9889 0.00658571
R47393 DVDD.n9890 DVDD.n9819 0.00658571
R47394 DVDD.n9897 DVDD.n9819 0.00658571
R47395 DVDD.n9898 DVDD.n9897 0.00658571
R47396 DVDD.n9935 DVDD.n9898 0.00658571
R47397 DVDD.n9935 DVDD.n9934 0.00658571
R47398 DVDD.n9934 DVDD.n9933 0.00658571
R47399 DVDD.n9933 DVDD.n9899 0.00658571
R47400 DVDD.n9903 DVDD.n9899 0.00658571
R47401 DVDD.n9926 DVDD.n9903 0.00658571
R47402 DVDD.n9926 DVDD.n9925 0.00658571
R47403 DVDD.n9925 DVDD.n9924 0.00658571
R47404 DVDD.n9924 DVDD.n9904 0.00658571
R47405 DVDD.n9917 DVDD.n9904 0.00658571
R47406 DVDD.n9917 DVDD.n9916 0.00658571
R47407 DVDD.n9916 DVDD.n9915 0.00658571
R47408 DVDD.n9915 DVDD.n9907 0.00658571
R47409 DVDD.n9908 DVDD.n9907 0.00658571
R47410 DVDD.n9908 DVDD.n9651 0.00658571
R47411 DVDD.n10088 DVDD.n9651 0.00658571
R47412 DVDD.n10088 DVDD.n10087 0.00658571
R47413 DVDD.n10087 DVDD.n10086 0.00658571
R47414 DVDD.n10086 DVDD.n9652 0.00658571
R47415 DVDD.n10081 DVDD.n9652 0.00658571
R47416 DVDD.n10081 DVDD.n10080 0.00658571
R47417 DVDD.n10080 DVDD.n10079 0.00658571
R47418 DVDD.n10079 DVDD.n9654 0.00658571
R47419 DVDD.n10073 DVDD.n9654 0.00658571
R47420 DVDD.n10073 DVDD.n10072 0.00658571
R47421 DVDD.n10072 DVDD.n10071 0.00658571
R47422 DVDD.n10071 DVDD.n9659 0.00658571
R47423 DVDD.n9706 DVDD.n9659 0.00658571
R47424 DVDD.n9711 DVDD.n9706 0.00658571
R47425 DVDD.n9712 DVDD.n9711 0.00658571
R47426 DVDD.n9713 DVDD.n9712 0.00658571
R47427 DVDD.n9713 DVDD.n9703 0.00658571
R47428 DVDD.n9720 DVDD.n9703 0.00658571
R47429 DVDD.n9721 DVDD.n9720 0.00658571
R47430 DVDD.n9722 DVDD.n9721 0.00658571
R47431 DVDD.n9722 DVDD.n9700 0.00658571
R47432 DVDD.n9729 DVDD.n9700 0.00658571
R47433 DVDD.n9730 DVDD.n9729 0.00658571
R47434 DVDD.n10063 DVDD.n9730 0.00658571
R47435 DVDD.n10063 DVDD.n10062 0.00658571
R47436 DVDD.n10062 DVDD.n10061 0.00658571
R47437 DVDD.n10061 DVDD.n9731 0.00658571
R47438 DVDD.n9976 DVDD.n9731 0.00658571
R47439 DVDD.n9977 DVDD.n9976 0.00658571
R47440 DVDD.n9977 DVDD.n9974 0.00658571
R47441 DVDD.n9984 DVDD.n9974 0.00658571
R47442 DVDD.n9985 DVDD.n9984 0.00658571
R47443 DVDD.n9986 DVDD.n9985 0.00658571
R47444 DVDD.n9986 DVDD.n9971 0.00658571
R47445 DVDD.n9993 DVDD.n9971 0.00658571
R47446 DVDD.n9994 DVDD.n9993 0.00658571
R47447 DVDD.n9995 DVDD.n9994 0.00658571
R47448 DVDD.n9995 DVDD.n9968 0.00658571
R47449 DVDD.n10006 DVDD.n9968 0.00658571
R47450 DVDD.n10007 DVDD.n10006 0.00658571
R47451 DVDD.n10052 DVDD.n10007 0.00658571
R47452 DVDD.n10052 DVDD.n10051 0.00658571
R47453 DVDD.n10051 DVDD.n10050 0.00658571
R47454 DVDD.n10050 DVDD.n10008 0.00658571
R47455 DVDD.n10044 DVDD.n10008 0.00658571
R47456 DVDD.n10044 DVDD.n10043 0.00658571
R47457 DVDD.n10043 DVDD.n10042 0.00658571
R47458 DVDD.n10042 DVDD.n10010 0.00658571
R47459 DVDD.n10035 DVDD.n10010 0.00658571
R47460 DVDD.n10035 DVDD.n10034 0.00658571
R47461 DVDD.n10034 DVDD.n10033 0.00658571
R47462 DVDD.n10033 DVDD.n10013 0.00658571
R47463 DVDD.n10026 DVDD.n10013 0.00658571
R47464 DVDD.n10026 DVDD.n10025 0.00658571
R47465 DVDD.n10025 DVDD.n10024 0.00658571
R47466 DVDD.n4767 DVDD.n4766 0.006575
R47467 DVDD.n4548 DVDD.n4406 0.006575
R47468 DVDD DVDD.n18113 0.00655123
R47469 DVDD.n18112 DVDD 0.00655123
R47470 DVDD.n20241 DVDD.n19970 0.00654286
R47471 DVDD.n20317 DVDD.n19835 0.00654286
R47472 DVDD.n20733 DVDD.n19153 0.00654286
R47473 DVDD.n20807 DVDD.n18881 0.00654286
R47474 DVDD.n274 DVDD.n236 0.00654286
R47475 DVDD.n426 DVDD.n421 0.00654286
R47476 DVDD.n10084 DVDD.n9613 0.00654286
R47477 DVDD.n10001 DVDD.n9997 0.00654286
R47478 DVDD.n21112 DVDD.n21088 0.00654286
R47479 DVDD.n22271 DVDD.n71 0.00654286
R47480 DVDD.n2686 DVDD.n2336 0.0065
R47481 DVDD.n2710 DVDD.n2686 0.0065
R47482 DVDD.n3027 DVDD.n2710 0.0065
R47483 DVDD.n15395 DVDD.n5111 0.0065
R47484 DVDD.n15686 DVDD.n5111 0.0065
R47485 DVDD.n15912 DVDD.n3231 0.0065
R47486 DVDD.n15879 DVDD.n15878 0.0065
R47487 DVDD.n5225 DVDD.n5113 0.0065
R47488 DVDD.n15913 DVDD.n15912 0.0065
R47489 DVDD.n15348 DVDD.n5225 0.0065
R47490 DVDD.n15913 DVDD.n3147 0.0065
R47491 DVDD.n16240 DVDD.n16199 0.0065
R47492 DVDD.n15879 DVDD.n2708 0.0065
R47493 DVDD.n16134 DVDD.n2708 0.0065
R47494 DVDD.n2527 DVDD.n2523 0.0065
R47495 DVDD.n16240 DVDD.n2527 0.0065
R47496 DVDD.n5113 DVDD.n3506 0.0065
R47497 DVDD.n15813 DVDD.n3148 0.0065
R47498 DVDD.n15686 DVDD.n3505 0.0065
R47499 DVDD.n16362 DVDD.n16361 0.0065
R47500 DVDD.n16361 DVDD.n2525 0.0065
R47501 DVDD.n15990 DVDD.n3148 0.0065
R47502 DVDD.n15991 DVDD.n15990 0.0065
R47503 DVDD.n16195 DVDD.n2525 0.0065
R47504 DVDD.n4776 DVDD.n3635 0.0064625
R47505 DVDD.n14306 DVDD.n8254 0.00645489
R47506 DVDD.n21673 DVDD.n18378 0.00644438
R47507 DVDD.n21358 DVDD.n138 0.00644438
R47508 DVDD.n21998 DVDD.n18244 0.00644438
R47509 DVDD.n4858 DVDD.n4857 0.00644438
R47510 DVDD DVDD.n22348 0.00641429
R47511 DVDD.n20336 DVDD 0.00641429
R47512 DVDD.n20200 DVDD.n19738 0.00641429
R47513 DVDD.n20275 DVDD.n19941 0.00641429
R47514 DVDD.n20849 DVDD 0.00641429
R47515 DVDD.n20692 DVDD.n18845 0.00641429
R47516 DVDD.n20767 DVDD.n19051 0.00641429
R47517 DVDD DVDD.n22088 0.00641429
R47518 DVDD.n4047 DVDD.n3874 0.00641429
R47519 DVDD.n324 DVDD.n302 0.00641429
R47520 DVDD.n10019 DVDD 0.00641429
R47521 DVDD.n9814 DVDD.n9770 0.00641429
R47522 DVDD.n9701 DVDD.n9692 0.00641429
R47523 DVDD.n18715 DVDD.n18675 0.00641429
R47524 DVDD.n21130 DVDD.n102 0.00641429
R47525 DVDD.n20082 DVDD.n20081 0.00637368
R47526 DVDD.n20083 DVDD.n20082 0.00637368
R47527 DVDD.n20083 DVDD.n20079 0.00637368
R47528 DVDD.n20087 DVDD.n20079 0.00637368
R47529 DVDD.n20088 DVDD.n20087 0.00637368
R47530 DVDD.n20089 DVDD.n20088 0.00637368
R47531 DVDD.n20089 DVDD.n20070 0.00637368
R47532 DVDD.n20100 DVDD.n20099 0.00637368
R47533 DVDD.n20099 DVDD.n20098 0.00637368
R47534 DVDD.n20098 DVDD.n20093 0.00637368
R47535 DVDD.n20094 DVDD.n20093 0.00637368
R47536 DVDD.n20094 DVDD.n19708 0.00637368
R47537 DVDD.n20596 DVDD.n19708 0.00637368
R47538 DVDD.n21271 DVDD.n18654 0.00637368
R47539 DVDD.n21222 DVDD.n18654 0.00637368
R47540 DVDD.n21222 DVDD.n18660 0.00637368
R47541 DVDD.n21260 DVDD.n18660 0.00637368
R47542 DVDD.n21260 DVDD.n137 0.00637368
R47543 DVDD.n21359 DVDD.n137 0.00637368
R47544 DVDD.n21360 DVDD.n21359 0.00637368
R47545 DVDD.n21360 DVDD.n18549 0.00637368
R47546 DVDD.n21369 DVDD.n18549 0.00637368
R47547 DVDD.n21684 DVDD.n18534 0.00637368
R47548 DVDD.n18539 DVDD.n18534 0.00637368
R47549 DVDD.n21671 DVDD.n18539 0.00637368
R47550 DVDD.n21672 DVDD.n21671 0.00637368
R47551 DVDD.n21672 DVDD.n18301 0.00637368
R47552 DVDD.n18375 DVDD.n18301 0.00637368
R47553 DVDD.n18375 DVDD.n18307 0.00637368
R47554 DVDD.n18314 DVDD.n18307 0.00637368
R47555 DVDD.n18365 DVDD.n18314 0.00637368
R47556 DVDD.n18365 DVDD.n18364 0.00637368
R47557 DVDD.n18340 DVDD.n18315 0.00637368
R47558 DVDD.n18340 DVDD.n18331 0.00637368
R47559 DVDD.n18350 DVDD.n18331 0.00637368
R47560 DVDD.n18350 DVDD.n18332 0.00637368
R47561 DVDD.n18332 DVDD.n18243 0.00637368
R47562 DVDD.n21997 DVDD.n18243 0.00637368
R47563 DVDD.n21997 DVDD.n21990 0.00637368
R47564 DVDD.n22008 DVDD.n21990 0.00637368
R47565 DVDD.n22008 DVDD.n21991 0.00637368
R47566 DVDD.n21991 DVDD.n229 0.00637368
R47567 DVDD.n20897 DVDD.n20896 0.00637368
R47568 DVDD.n20896 DVDD.n20895 0.00637368
R47569 DVDD.n20895 DVDD.n18925 0.00637368
R47570 DVDD.n20891 DVDD.n18925 0.00637368
R47571 DVDD.n20891 DVDD.n20890 0.00637368
R47572 DVDD.n20890 DVDD.n20889 0.00637368
R47573 DVDD.n20889 DVDD.n18927 0.00637368
R47574 DVDD.n20864 DVDD.n20863 0.00637368
R47575 DVDD.n20863 DVDD.n20862 0.00637368
R47576 DVDD.n20862 DVDD.n18958 0.00637368
R47577 DVDD.n20858 DVDD.n18958 0.00637368
R47578 DVDD.n20858 DVDD.n20857 0.00637368
R47579 DVDD.n20857 DVDD.n20856 0.00637368
R47580 DVDD.n22239 DVDD.n129 0.00637368
R47581 DVDD.n18482 DVDD.n129 0.00637368
R47582 DVDD.n18482 DVDD.n18480 0.00637368
R47583 DVDD.n18480 DVDD.n157 0.00637368
R47584 DVDD.n22228 DVDD.n157 0.00637368
R47585 DVDD.n22228 DVDD.n22227 0.00637368
R47586 DVDD.n22227 DVDD.n158 0.00637368
R47587 DVDD.n18427 DVDD.n158 0.00637368
R47588 DVDD.n21734 DVDD.n18427 0.00637368
R47589 DVDD.n21769 DVDD.n21768 0.00637368
R47590 DVDD.n21768 DVDD.n21767 0.00637368
R47591 DVDD.n21767 DVDD.n18386 0.00637368
R47592 DVDD.n21778 DVDD.n18386 0.00637368
R47593 DVDD.n21943 DVDD.n21778 0.00637368
R47594 DVDD.n21943 DVDD.n21942 0.00637368
R47595 DVDD.n21942 DVDD.n21780 0.00637368
R47596 DVDD.n21787 DVDD.n21780 0.00637368
R47597 DVDD.n21932 DVDD.n21787 0.00637368
R47598 DVDD.n21932 DVDD.n21931 0.00637368
R47599 DVDD.n21930 DVDD.n21791 0.00637368
R47600 DVDD.n21897 DVDD.n21791 0.00637368
R47601 DVDD.n21897 DVDD.n21798 0.00637368
R47602 DVDD.n21919 DVDD.n21798 0.00637368
R47603 DVDD.n21919 DVDD.n18240 0.00637368
R47604 DVDD.n22044 DVDD.n18240 0.00637368
R47605 DVDD.n22044 DVDD.n18212 0.00637368
R47606 DVDD.n22062 DVDD.n18212 0.00637368
R47607 DVDD.n22062 DVDD.n18204 0.00637368
R47608 DVDD.n22069 DVDD.n18204 0.00637368
R47609 DVDD.n20355 DVDD.n18939 0.00635
R47610 DVDD.n20832 DVDD.n18967 0.00635
R47611 DVDD.n22122 DVDD.n446 0.00635
R47612 DVDD.n4760 DVDD.n3665 0.00635
R47613 DVDD.n18092 DVDD.n18091 0.00635
R47614 DVDD.n4544 DVDD.n4403 0.00635
R47615 DVDD.n10038 DVDD.n799 0.00635
R47616 DVDD.n22329 DVDD.n26 0.00635
R47617 DVDD.n10236 DVDD.n10223 0.00631955
R47618 DVDD.n12382 DVDD.n12381 0.00629866
R47619 DVDD.n12894 DVDD.n12387 0.00629866
R47620 DVDD.n13495 DVDD.n12379 0.00629866
R47621 DVDD.n12893 DVDD.n12385 0.00629866
R47622 DVDD.n18086 DVDD.n18085 0.00629375
R47623 DVDD.n20184 DVDD.n19734 0.00628571
R47624 DVDD.n19950 DVDD.n19936 0.00628571
R47625 DVDD.n20676 DVDD.n18840 0.00628571
R47626 DVDD.n20751 DVDD.n19046 0.00628571
R47627 DVDD.n3898 DVDD.n3871 0.00628571
R47628 DVDD.n333 DVDD.n299 0.00628571
R47629 DVDD.n9882 DVDD.n9765 0.00628571
R47630 DVDD.n10068 DVDD.n9667 0.00628571
R47631 DVDD.n19674 DVDD.n18682 0.00628571
R47632 DVDD.n21121 DVDD.n98 0.00628571
R47633 DVDD.n4590 DVDD.n4248 0.0062375
R47634 DVDD.n4428 DVDD.n3760 0.0062375
R47635 DVDD.n4398 DVDD.n4323 0.0062375
R47636 DVDD.n17712 DVDD.n911 0.0062375
R47637 DVDD.n17711 DVDD.n909 0.0062375
R47638 DVDD.n15126 DVDD.n5743 0.0062375
R47639 DVDD.n5741 DVDD.n5643 0.0062375
R47640 DVDD.n15123 DVDD.n5741 0.00619869
R47641 DVDD.n15068 DVDD.n7055 0.00619869
R47642 DVDD.n15124 DVDD.n5743 0.00619869
R47643 DVDD.n15067 DVDD.n7053 0.00619869
R47644 DVDD.n20177 DVDD.n19733 0.00615714
R47645 DVDD.n20669 DVDD.n18839 0.00615714
R47646 DVDD.n3993 DVDD.n3870 0.00615714
R47647 DVDD.n9875 DVDD.n9764 0.00615714
R47648 DVDD.n18691 DVDD.n18684 0.00615714
R47649 DVDD.n4423 DVDD.n3737 0.006125
R47650 DVDD.n4278 DVDD.n4250 0.006125
R47651 DVDD.n20363 DVDD.n18938 0.00609286
R47652 DVDD.n20825 DVDD.n18966 0.00609286
R47653 DVDD.n22129 DVDD.n435 0.00609286
R47654 DVDD.n17877 DVDD.n800 0.00609286
R47655 DVDD.n22342 DVDD.n27 0.00609286
R47656 DVDD.n3618 DVDD.n3538 0.00606875
R47657 DVDD.n20193 DVDD.n19737 0.00602857
R47658 DVDD.n19947 DVDD.n19940 0.00602857
R47659 DVDD.n20685 DVDD.n18844 0.00602857
R47660 DVDD.n20760 DVDD.n19050 0.00602857
R47661 DVDD.n4054 DVDD.n3873 0.00602857
R47662 DVDD.n342 DVDD.n301 0.00602857
R47663 DVDD.n9891 DVDD.n9769 0.00602857
R47664 DVDD.n9714 DVDD.n9691 0.00602857
R47665 DVDD.n21204 DVDD.n18677 0.00602857
R47666 DVDD.n21124 DVDD.n101 0.00602857
R47667 DVDD.n3753 DVDD.n3733 0.0060125
R47668 DVDD.n21938 DVDD 0.00600694
R47669 DVDD.n21777 DVDD.n18297 0.00597492
R47670 DVDD.n159 DVDD.n155 0.00597492
R47671 DVDD.n22043 DVDD.n22041 0.00597492
R47672 DVDD.n18115 DVDD.n18095 0.00597492
R47673 DVDD.n20346 DVDD.n18942 0.00596429
R47674 DVDD.n20841 DVDD.n18970 0.00596429
R47675 DVDD.n22100 DVDD.n22078 0.00596429
R47676 DVDD.n10029 DVDD.n793 0.00596429
R47677 DVDD.n22321 DVDD.n23 0.00596429
R47678 DVDD.n19896 DVDD.n19895 0.0059439
R47679 DVDD.n19897 DVDD.n19896 0.0059439
R47680 DVDD.n19897 DVDD.n19893 0.0059439
R47681 DVDD.n19901 DVDD.n19893 0.0059439
R47682 DVDD.n19902 DVDD.n19901 0.0059439
R47683 DVDD.n19903 DVDD.n19902 0.0059439
R47684 DVDD.n19903 DVDD.n19884 0.0059439
R47685 DVDD.n19914 DVDD.n19913 0.0059439
R47686 DVDD.n19913 DVDD.n19912 0.0059439
R47687 DVDD.n19912 DVDD.n19907 0.0059439
R47688 DVDD.n19908 DVDD.n19907 0.0059439
R47689 DVDD.n19908 DVDD.n19821 0.0059439
R47690 DVDD.n20441 DVDD.n19821 0.0059439
R47691 DVDD.n22243 DVDD.n121 0.0059439
R47692 DVDD.n18461 DVDD.n121 0.0059439
R47693 DVDD.n18494 DVDD.n18461 0.0059439
R47694 DVDD.n18495 DVDD.n18494 0.0059439
R47695 DVDD.n18495 DVDD.n150 0.0059439
R47696 DVDD.n21582 DVDD.n150 0.0059439
R47697 DVDD.n21583 DVDD.n21582 0.0059439
R47698 DVDD.n21593 DVDD.n21583 0.0059439
R47699 DVDD.n21594 DVDD.n21593 0.0059439
R47700 DVDD.n21754 DVDD.n18403 0.0059439
R47701 DVDD.n21755 DVDD.n21754 0.0059439
R47702 DVDD.n21756 DVDD.n21755 0.0059439
R47703 DVDD.n21757 DVDD.n21756 0.0059439
R47704 DVDD.n21757 DVDD.n18382 0.0059439
R47705 DVDD.n21865 DVDD.n18382 0.0059439
R47706 DVDD.n21865 DVDD.n21864 0.0059439
R47707 DVDD.n21864 DVDD.n21863 0.0059439
R47708 DVDD.n21863 DVDD.n21857 0.0059439
R47709 DVDD.n21858 DVDD.n21857 0.0059439
R47710 DVDD.n21814 DVDD.n21809 0.0059439
R47711 DVDD.n21814 DVDD.n21803 0.0059439
R47712 DVDD.n21914 DVDD.n21803 0.0059439
R47713 DVDD.n21915 DVDD.n21914 0.0059439
R47714 DVDD.n21915 DVDD.n18225 0.0059439
R47715 DVDD.n22048 DVDD.n18225 0.0059439
R47716 DVDD.n22050 DVDD.n22048 0.0059439
R47717 DVDD.n22050 DVDD.n22049 0.0059439
R47718 DVDD.n22049 DVDD.n18220 0.0059439
R47719 DVDD.n18220 DVDD.n315 0.0059439
R47720 DVDD.n20438 DVDD.n20437 0.0059439
R47721 DVDD.n20437 DVDD.n19825 0.0059439
R47722 DVDD.n20433 DVDD.n19825 0.0059439
R47723 DVDD.n20433 DVDD.n19827 0.0059439
R47724 DVDD.n20429 DVDD.n19827 0.0059439
R47725 DVDD.n20429 DVDD.n19830 0.0059439
R47726 DVDD.n20425 DVDD.n19830 0.0059439
R47727 DVDD.n20397 DVDD.n20396 0.0059439
R47728 DVDD.n20396 DVDD.n20385 0.0059439
R47729 DVDD.n20392 DVDD.n20385 0.0059439
R47730 DVDD.n20392 DVDD.n20388 0.0059439
R47731 DVDD.n20388 DVDD.n18919 0.0059439
R47732 DVDD.n20900 DVDD.n18919 0.0059439
R47733 DVDD.n20919 DVDD.n18908 0.0059439
R47734 DVDD.n20922 DVDD.n18908 0.0059439
R47735 DVDD.n21048 DVDD.n57 0.0059439
R47736 DVDD.n22241 DVDD.n125 0.0059439
R47737 DVDD.n18484 DVDD.n125 0.0059439
R47738 DVDD.n18484 DVDD.n18458 0.0059439
R47739 DVDD.n18497 DVDD.n18458 0.0059439
R47740 DVDD.n18497 DVDD.n156 0.0059439
R47741 DVDD.n22225 DVDD.n156 0.0059439
R47742 DVDD.n22225 DVDD.n22224 0.0059439
R47743 DVDD.n22224 DVDD.n165 0.0059439
R47744 DVDD.n18426 DVDD.n165 0.0059439
R47745 DVDD.n18424 DVDD.n18396 0.0059439
R47746 DVDD.n21762 DVDD.n18396 0.0059439
R47747 DVDD.n21762 DVDD.n21761 0.0059439
R47748 DVDD.n21761 DVDD.n21759 0.0059439
R47749 DVDD.n21759 DVDD.n18298 0.0059439
R47750 DVDD.n21839 DVDD.n18298 0.0059439
R47751 DVDD.n21878 DVDD.n21839 0.0059439
R47752 DVDD.n21878 DVDD.n21877 0.0059439
R47753 DVDD.n21877 DVDD.n21875 0.0059439
R47754 DVDD.n21875 DVDD.n21811 0.0059439
R47755 DVDD.n21901 DVDD.n21900 0.0059439
R47756 DVDD.n21900 DVDD.n21828 0.0059439
R47757 DVDD.n21828 DVDD.n21800 0.0059439
R47758 DVDD.n21917 DVDD.n21800 0.0059439
R47759 DVDD.n21917 DVDD.n18228 0.0059439
R47760 DVDD.n22046 DVDD.n18228 0.0059439
R47761 DVDD.n22046 DVDD.n18215 0.0059439
R47762 DVDD.n22060 DVDD.n18215 0.0059439
R47763 DVDD.n22060 DVDD.n22059 0.0059439
R47764 DVDD.n22059 DVDD.n366 0.0059439
R47765 DVDD.n19983 DVDD.n19982 0.0059439
R47766 DVDD.n19984 DVDD.n19983 0.0059439
R47767 DVDD.n19984 DVDD.n19979 0.0059439
R47768 DVDD.n19988 DVDD.n19979 0.0059439
R47769 DVDD.n19989 DVDD.n19988 0.0059439
R47770 DVDD.n19990 DVDD.n19989 0.0059439
R47771 DVDD.n19990 DVDD.n19969 0.0059439
R47772 DVDD.n20001 DVDD.n20000 0.0059439
R47773 DVDD.n20000 DVDD.n19999 0.0059439
R47774 DVDD.n19999 DVDD.n19994 0.0059439
R47775 DVDD.n19995 DVDD.n19994 0.0059439
R47776 DVDD.n19995 DVDD.n19766 0.0059439
R47777 DVDD.n20541 DVDD.n19766 0.0059439
R47778 DVDD.n21215 DVDD.n18671 0.0059439
R47779 DVDD.n21215 DVDD.n18665 0.0059439
R47780 DVDD.n21255 DVDD.n18665 0.0059439
R47781 DVDD.n21256 DVDD.n21255 0.0059439
R47782 DVDD.n21256 DVDD.n136 0.0059439
R47783 DVDD.n21354 DVDD.n136 0.0059439
R47784 DVDD.n21354 DVDD.n18556 0.0059439
R47785 DVDD.n21651 DVDD.n18556 0.0059439
R47786 DVDD.n21651 DVDD.n21650 0.0059439
R47787 DVDD.n21689 DVDD.n18529 0.0059439
R47788 DVDD.n21691 DVDD.n21689 0.0059439
R47789 DVDD.n21691 DVDD.n21690 0.0059439
R47790 DVDD.n21690 DVDD.n18296 0.0059439
R47791 DVDD.n21945 DVDD.n18296 0.0059439
R47792 DVDD.n21947 DVDD.n21945 0.0059439
R47793 DVDD.n21948 DVDD.n21947 0.0059439
R47794 DVDD.n21948 DVDD.n18283 0.0059439
R47795 DVDD.n21962 DVDD.n18283 0.0059439
R47796 DVDD.n21964 DVDD.n21962 0.0059439
R47797 DVDD.n21965 DVDD.n18269 0.0059439
R47798 DVDD.n21977 DVDD.n18269 0.0059439
R47799 DVDD.n21979 DVDD.n21977 0.0059439
R47800 DVDD.n21980 DVDD.n21979 0.0059439
R47801 DVDD.n21980 DVDD.n18265 0.0059439
R47802 DVDD.n22035 DVDD.n18265 0.0059439
R47803 DVDD.n22035 DVDD.n22034 0.0059439
R47804 DVDD.n22034 DVDD.n21987 0.0059439
R47805 DVDD.n21987 DVDD.n235 0.0059439
R47806 DVDD.n22183 DVDD.n235 0.0059439
R47807 DVDD.n20593 DVDD.n19713 0.0059439
R47808 DVDD.n20589 DVDD.n19713 0.0059439
R47809 DVDD.n20589 DVDD.n19715 0.0059439
R47810 DVDD.n20585 DVDD.n19715 0.0059439
R47811 DVDD.n20585 DVDD.n19717 0.0059439
R47812 DVDD.n20581 DVDD.n19717 0.0059439
R47813 DVDD.n20581 DVDD.n19719 0.0059439
R47814 DVDD.n20554 DVDD.n20553 0.0059439
R47815 DVDD.n20553 DVDD.n19760 0.0059439
R47816 DVDD.n20549 DVDD.n19760 0.0059439
R47817 DVDD.n20549 DVDD.n19762 0.0059439
R47818 DVDD.n20545 DVDD.n19762 0.0059439
R47819 DVDD.n20545 DVDD.n19764 0.0059439
R47820 DVDD.n20516 DVDD.n20487 0.0059439
R47821 DVDD.n20519 DVDD.n20487 0.0059439
R47822 DVDD.n21012 DVDD.n18699 0.0059439
R47823 DVDD.n21247 DVDD.n21217 0.0059439
R47824 DVDD.n21234 DVDD.n21217 0.0059439
R47825 DVDD.n21234 DVDD.n18662 0.0059439
R47826 DVDD.n21258 DVDD.n18662 0.0059439
R47827 DVDD.n21258 DVDD.n145 0.0059439
R47828 DVDD.n21356 DVDD.n145 0.0059439
R47829 DVDD.n21356 DVDD.n18551 0.0059439
R47830 DVDD.n21653 DVDD.n18551 0.0059439
R47831 DVDD.n21653 DVDD.n18552 0.0059439
R47832 DVDD.n21686 DVDD.n18526 0.0059439
R47833 DVDD.n21693 DVDD.n18526 0.0059439
R47834 DVDD.n21693 DVDD.n18519 0.0059439
R47835 DVDD.n21704 DVDD.n18519 0.0059439
R47836 DVDD.n21704 DVDD.n18384 0.0059439
R47837 DVDD.n18384 DVDD.n18293 0.0059439
R47838 DVDD.n21950 DVDD.n18293 0.0059439
R47839 DVDD.n21950 DVDD.n18285 0.0059439
R47840 DVDD.n21960 DVDD.n18285 0.0059439
R47841 DVDD.n21960 DVDD.n18280 0.0059439
R47842 DVDD.n21967 DVDD.n18271 0.0059439
R47843 DVDD.n21975 DVDD.n18271 0.0059439
R47844 DVDD.n21975 DVDD.n18266 0.0059439
R47845 DVDD.n21982 DVDD.n18266 0.0059439
R47846 DVDD.n22038 DVDD.n21982 0.0059439
R47847 DVDD.n22038 DVDD.n22037 0.0059439
R47848 DVDD.n22037 DVDD.n21984 0.0059439
R47849 DVDD.n22023 DVDD.n21984 0.0059439
R47850 DVDD.n22023 DVDD.n230 0.0059439
R47851 DVDD.n22185 DVDD.n230 0.0059439
R47852 DVDD.n6702 DVDD.n6701 0.00591353
R47853 DVDD.n8138 DVDD.n7685 0.00591353
R47854 DVDD.n20286 DVDD.n20285 0.0059
R47855 DVDD.n19850 DVDD.n19834 0.0059
R47856 DVDD.n20779 DVDD.n19022 0.0059
R47857 DVDD.n20814 DVDD.n18882 0.0059
R47858 DVDD.n22158 DVDD.n304 0.0059
R47859 DVDD.n388 DVDD.n372 0.0059
R47860 DVDD.n4427 DVDD.n3750 0.0059
R47861 DVDD.n10066 DVDD.n9696 0.0059
R47862 DVDD.n9964 DVDD.n9750 0.0059
R47863 DVDD.n93 DVDD.n85 0.0059
R47864 DVDD.n22300 DVDD.n42 0.0059
R47865 DVDD DVDD.n179 0.00587887
R47866 DVDD.n3624 DVDD.n3528 0.00584375
R47867 DVDD.n20166 DVDD.n20165 0.00583571
R47868 DVDD.n20658 DVDD.n20657 0.00583571
R47869 DVDD.n3978 DVDD.n3906 0.00583571
R47870 DVDD.n9864 DVDD.n5477 0.00583571
R47871 DVDD.n19701 DVDD.n19207 0.00583571
R47872 DVDD.n4578 DVDD.n4577 0.005825
R47873 DVDD.n4579 DVDD.n4578 0.005825
R47874 DVDD.n4579 DVDD.n4277 0.005825
R47875 DVDD.n4583 DVDD.n4277 0.005825
R47876 DVDD.n4584 DVDD.n4583 0.005825
R47877 DVDD.n4594 DVDD.n4584 0.005825
R47878 DVDD.n4594 DVDD.n4593 0.005825
R47879 DVDD.n4593 DVDD.n4592 0.005825
R47880 DVDD.n4592 DVDD.n4585 0.005825
R47881 DVDD.n4586 DVDD.n4585 0.005825
R47882 DVDD.n18131 DVDD.n18130 0.005825
R47883 DVDD.n18130 DVDD.n18129 0.005825
R47884 DVDD.n18129 DVDD.n494 0.005825
R47885 DVDD.n18075 DVDD.n494 0.005825
R47886 DVDD.n18076 DVDD.n18075 0.005825
R47887 DVDD.n18076 DVDD.n18071 0.005825
R47888 DVDD.n18088 DVDD.n18071 0.005825
R47889 DVDD.n18089 DVDD.n18088 0.005825
R47890 DVDD.n18090 DVDD.n18089 0.005825
R47891 DVDD.n4457 DVDD.n4456 0.005825
R47892 DVDD.n4552 DVDD.n4457 0.005825
R47893 DVDD.n4552 DVDD.n4551 0.005825
R47894 DVDD.n4551 DVDD.n4550 0.005825
R47895 DVDD.n4550 DVDD.n4458 0.005825
R47896 DVDD.n4543 DVDD.n4458 0.005825
R47897 DVDD.n4543 DVDD.n4542 0.005825
R47898 DVDD.n4542 DVDD.n4541 0.005825
R47899 DVDD.n4541 DVDD.n4461 0.005825
R47900 DVDD.n4461 DVDD.n4199 0.005825
R47901 DVDD.n4474 DVDD.n4200 0.005825
R47902 DVDD.n4474 DVDD.n4321 0.005825
R47903 DVDD.n4561 DVDD.n4321 0.005825
R47904 DVDD.n4562 DVDD.n4561 0.005825
R47905 DVDD.n4563 DVDD.n4562 0.005825
R47906 DVDD.n4563 DVDD.n4317 0.005825
R47907 DVDD.n4569 DVDD.n4317 0.005825
R47908 DVDD.n4570 DVDD.n4569 0.005825
R47909 DVDD.n4571 DVDD.n4570 0.005825
R47910 DVDD.n4757 DVDD.n4756 0.005825
R47911 DVDD.n4756 DVDD.n4755 0.005825
R47912 DVDD.n4755 DVDD.n3714 0.005825
R47913 DVDD.n4748 DVDD.n3714 0.005825
R47914 DVDD.n4748 DVDD.n4747 0.005825
R47915 DVDD.n4747 DVDD.n4746 0.005825
R47916 DVDD.n4746 DVDD.n3720 0.005825
R47917 DVDD.n3756 DVDD.n3720 0.005825
R47918 DVDD.n4738 DVDD.n3756 0.005825
R47919 DVDD.n4738 DVDD.n4737 0.005825
R47920 DVDD.n4430 DVDD.n3757 0.005825
R47921 DVDD.n4430 DVDD.n4426 0.005825
R47922 DVDD.n4436 DVDD.n4426 0.005825
R47923 DVDD.n4437 DVDD.n4436 0.005825
R47924 DVDD.n4438 DVDD.n4437 0.005825
R47925 DVDD.n4438 DVDD.n4422 0.005825
R47926 DVDD.n4446 DVDD.n4422 0.005825
R47927 DVDD.n4447 DVDD.n4446 0.005825
R47928 DVDD.n4448 DVDD.n4447 0.005825
R47929 DVDD.n3614 DVDD.n3542 0.005825
R47930 DVDD.n3614 DVDD.n3610 0.005825
R47931 DVDD.n3620 DVDD.n3610 0.005825
R47932 DVDD.n3621 DVDD.n3620 0.005825
R47933 DVDD.n3622 DVDD.n3621 0.005825
R47934 DVDD.n3622 DVDD.n3606 0.005825
R47935 DVDD.n3628 DVDD.n3606 0.005825
R47936 DVDD.n3629 DVDD.n3628 0.005825
R47937 DVDD.n3630 DVDD.n3629 0.005825
R47938 DVDD.n3630 DVDD.n3600 0.005825
R47939 DVDD.n4780 DVDD.n3601 0.005825
R47940 DVDD.n4774 DVDD.n3601 0.005825
R47941 DVDD.n4774 DVDD.n4773 0.005825
R47942 DVDD.n4773 DVDD.n4772 0.005825
R47943 DVDD.n4772 DVDD.n3637 0.005825
R47944 DVDD.n3672 DVDD.n3637 0.005825
R47945 DVDD.n4764 DVDD.n3672 0.005825
R47946 DVDD.n4764 DVDD.n4763 0.005825
R47947 DVDD.n4763 DVDD.n4762 0.005825
R47948 DVDD.n14304 DVDD.n8257 0.00581544
R47949 DVDD.n14305 DVDD.n8255 0.00581544
R47950 DVDD.n4444 DVDD.n3746 0.0057875
R47951 DVDD.n4778 DVDD.n3634 0.0057875
R47952 DVDD.n4258 DVDD.n4246 0.0057875
R47953 DVDD.n4779 DVDD.n3598 0.0057875
R47954 DVDD.n20230 DVDD.n19973 0.00577143
R47955 DVDD.n20308 DVDD.n19838 0.00577143
R47956 DVDD.n20722 DVDD.n19136 0.00577143
R47957 DVDD.n20798 DVDD.n18884 0.00577143
R47958 DVDD.n4018 DVDD.n239 0.00577143
R47959 DVDD.n411 DVDD.n376 0.00577143
R47960 DVDD.n9909 DVDD.n9616 0.00577143
R47961 DVDD.n9987 DVDD.n9753 0.00577143
R47962 DVDD.n21108 DVDD.n21096 0.00577143
R47963 DVDD.n22267 DVDD.n75 0.00577143
R47964 DVDD.n19024 DVDD.n18868 0.00572439
R47965 DVDD.n19031 DVDD.n18869 0.00572439
R47966 DVDD.n20931 DVDD.n20930 0.00572439
R47967 DVDD.n18904 DVDD.n18870 0.00572439
R47968 DVDD.n19075 DVDD.n18866 0.00572439
R47969 DVDD.n19127 DVDD.n18867 0.00572439
R47970 DVDD.n20969 DVDD.n18860 0.00572439
R47971 DVDD.n20968 DVDD.n18858 0.00572439
R47972 DVDD.n18310 DVDD.n196 0.00571437
R47973 DVDD.n22193 DVDD.n207 0.00571437
R47974 DVDD.n21721 DVDD.n18433 0.00571437
R47975 DVDD.n4862 DVDD.n4861 0.00571437
R47976 DVDD.n20133 DVDD.n20126 0.00570714
R47977 DVDD.n20620 DVDD.n20613 0.00570714
R47978 DVDD.n3956 DVDD.n3931 0.00570714
R47979 DVDD.n9834 DVDD.n5482 0.00570714
R47980 DVDD.n19642 DVDD.n19197 0.00570714
R47981 DVDD.n22252 DVDD.n97 0.00568049
R47982 DVDD.n104 DVDD.n90 0.00568049
R47983 DVDD.n3456 DVDD.n2369 0.00568049
R47984 DVDD.n16269 DVDD.n2692 0.00568049
R47985 DVDD.n22298 DVDD.n57 0.00568049
R47986 DVDD.n66 DVDD.n43 0.00568049
R47987 DVDD.n3455 DVDD.n2406 0.00568049
R47988 DVDD.n16313 DVDD.n2620 0.00568049
R47989 DVDD.n21185 DVDD.n18735 0.00568049
R47990 DVDD.n21083 DVDD.n18724 0.00568049
R47991 DVDD.n3458 DVDD.n3363 0.00568049
R47992 DVDD.n15908 DVDD.n3286 0.00568049
R47993 DVDD.n21212 DVDD.n18699 0.00568049
R47994 DVDD.n18703 DVDD.n18686 0.00568049
R47995 DVDD.n3461 DVDD.n3460 0.00568049
R47996 DVDD.n15679 DVDD.n15609 0.00568049
R47997 DVDD.n4535 DVDD.n4393 0.005675
R47998 DVDD.n15105 DVDD.n6344 0.005675
R47999 DVDD.n21370 DVDD.n21369 0.00566316
R48000 DVDD.n21734 DVDD.n18428 0.00566316
R48001 DVDD.n20214 DVDD.n19977 0.00564286
R48002 DVDD.n20706 DVDD.n19140 0.00564286
R48003 DVDD.n4008 DVDD.n243 0.00564286
R48004 DVDD.n9901 DVDD.n9620 0.00564286
R48005 DVDD.n21186 DVDD.n18729 0.00564286
R48006 DVDD.n18072 DVDD.n18059 0.00561875
R48007 DVDD.n5017 DVDD.n5016 0.00561579
R48008 DVDD.n5029 DVDD.n4891 0.00561579
R48009 DVDD.n5032 DVDD.n4891 0.00561579
R48010 DVDD.n15706 DVDD.n4905 0.00561579
R48011 DVDD.n15702 DVDD.n4905 0.00561579
R48012 DVDD.n5264 DVDD.n5263 0.00561579
R48013 DVDD.n5276 DVDD.n5061 0.00561579
R48014 DVDD.n5279 DVDD.n5061 0.00561579
R48015 DVDD.n5293 DVDD.n5292 0.00561579
R48016 DVDD.n5309 DVDD.n5308 0.00561579
R48017 DVDD.n5314 DVDD.n5080 0.00561579
R48018 DVDD.n5315 DVDD.n5314 0.00561579
R48019 DVDD.n5325 DVDD.n5324 0.00561579
R48020 DVDD.n5341 DVDD.n5340 0.00561579
R48021 DVDD.n5357 DVDD.n5356 0.00561579
R48022 DVDD.n15415 DVDD.n5261 0.00561579
R48023 DVDD.n15411 DVDD.n5261 0.00561579
R48024 DVDD.n15411 DVDD.n15410 0.00561579
R48025 DVDD.n5423 DVDD.n5422 0.00561579
R48026 DVDD.n5435 DVDD.n5401 0.00561579
R48027 DVDD.n5438 DVDD.n5401 0.00561579
R48028 DVDD.n5452 DVDD.n5451 0.00561579
R48029 DVDD.n15316 DVDD.n5409 0.00561579
R48030 DVDD.n15312 DVDD.n5409 0.00561579
R48031 DVDD.n15312 DVDD.n15311 0.00561579
R48032 DVDD.n15311 DVDD.n15310 0.00561579
R48033 DVDD.n15310 DVDD.n5460 0.00561579
R48034 DVDD.n15305 DVDD.n5460 0.00561579
R48035 DVDD.n15305 DVDD.n15304 0.00561579
R48036 DVDD.n15304 DVDD.n15303 0.00561579
R48037 DVDD.n15303 DVDD.n5462 0.00561579
R48038 DVDD.n15299 DVDD.n5462 0.00561579
R48039 DVDD.n15299 DVDD.n15298 0.00561579
R48040 DVDD.n15298 DVDD.n15297 0.00561579
R48041 DVDD.n15297 DVDD.n5464 0.00561579
R48042 DVDD.n15293 DVDD.n5464 0.00561579
R48043 DVDD.n15293 DVDD.n15292 0.00561579
R48044 DVDD.n15292 DVDD.n15291 0.00561579
R48045 DVDD.n15291 DVDD.n5466 0.00561579
R48046 DVDD.n5500 DVDD.n5499 0.00561579
R48047 DVDD.n5514 DVDD.n5496 0.00561579
R48048 DVDD.n15283 DVDD.n5497 0.00561579
R48049 DVDD.n15279 DVDD.n5497 0.00561579
R48050 DVDD.n15279 DVDD.n15278 0.00561579
R48051 DVDD.n15278 DVDD.n15277 0.00561579
R48052 DVDD.n15277 DVDD.n5518 0.00561579
R48053 DVDD.n15273 DVDD.n5518 0.00561579
R48054 DVDD.n15273 DVDD.n15272 0.00561579
R48055 DVDD.n15272 DVDD.n15271 0.00561579
R48056 DVDD.n15271 DVDD.n5520 0.00561579
R48057 DVDD.n15267 DVDD.n5520 0.00561579
R48058 DVDD.n15267 DVDD.n15266 0.00561579
R48059 DVDD.n15266 DVDD.n15265 0.00561579
R48060 DVDD.n15265 DVDD.n5522 0.00561579
R48061 DVDD.n15261 DVDD.n5522 0.00561579
R48062 DVDD.n15261 DVDD.n15260 0.00561579
R48063 DVDD.n15260 DVDD.n15259 0.00561579
R48064 DVDD.n15259 DVDD.n5524 0.00561579
R48065 DVDD.n15255 DVDD.n5524 0.00561579
R48066 DVDD.n15255 DVDD.n15254 0.00561579
R48067 DVDD.n15254 DVDD.n15253 0.00561579
R48068 DVDD.n15253 DVDD.n5526 0.00561579
R48069 DVDD.n15249 DVDD.n5526 0.00561579
R48070 DVDD.n15249 DVDD.n15248 0.00561579
R48071 DVDD.n15248 DVDD.n15247 0.00561579
R48072 DVDD.n15247 DVDD.n5528 0.00561579
R48073 DVDD.n15243 DVDD.n5528 0.00561579
R48074 DVDD.n15243 DVDD.n15242 0.00561579
R48075 DVDD.n15242 DVDD.n15241 0.00561579
R48076 DVDD.n15241 DVDD.n5530 0.00561579
R48077 DVDD.n15237 DVDD.n5530 0.00561579
R48078 DVDD.n15237 DVDD.n15236 0.00561579
R48079 DVDD.n15236 DVDD.n15235 0.00561579
R48080 DVDD.n15235 DVDD.n5532 0.00561579
R48081 DVDD.n15231 DVDD.n5532 0.00561579
R48082 DVDD.n15231 DVDD.n15230 0.00561579
R48083 DVDD.n15230 DVDD.n15229 0.00561579
R48084 DVDD.n15229 DVDD.n5534 0.00561579
R48085 DVDD.n15225 DVDD.n5534 0.00561579
R48086 DVDD.n15225 DVDD.n15224 0.00561579
R48087 DVDD.n15224 DVDD.n15223 0.00561579
R48088 DVDD.n15223 DVDD.n5536 0.00561579
R48089 DVDD.n15219 DVDD.n5536 0.00561579
R48090 DVDD.n15219 DVDD.n15218 0.00561579
R48091 DVDD.n15218 DVDD.n15217 0.00561579
R48092 DVDD.n15217 DVDD.n5538 0.00561579
R48093 DVDD.n15213 DVDD.n5538 0.00561579
R48094 DVDD.n15213 DVDD.n15212 0.00561579
R48095 DVDD.n15212 DVDD.n15211 0.00561579
R48096 DVDD.n15211 DVDD.n5540 0.00561579
R48097 DVDD.n15207 DVDD.n5540 0.00561579
R48098 DVDD.n15207 DVDD.n15206 0.00561579
R48099 DVDD.n15206 DVDD.n15205 0.00561579
R48100 DVDD.n15205 DVDD.n5542 0.00561579
R48101 DVDD.n15201 DVDD.n5542 0.00561579
R48102 DVDD.n15201 DVDD.n15200 0.00561579
R48103 DVDD.n15200 DVDD.n15199 0.00561579
R48104 DVDD.n15199 DVDD.n5544 0.00561579
R48105 DVDD.n15195 DVDD.n5544 0.00561579
R48106 DVDD.n15195 DVDD.n15194 0.00561579
R48107 DVDD.n15194 DVDD.n15193 0.00561579
R48108 DVDD.n15193 DVDD.n5546 0.00561579
R48109 DVDD.n15189 DVDD.n5546 0.00561579
R48110 DVDD.n15189 DVDD.n15188 0.00561579
R48111 DVDD.n15188 DVDD.n15187 0.00561579
R48112 DVDD.n15187 DVDD.n5548 0.00561579
R48113 DVDD.n15183 DVDD.n5548 0.00561579
R48114 DVDD.n15183 DVDD.n15182 0.00561579
R48115 DVDD.n15182 DVDD.n15181 0.00561579
R48116 DVDD.n15181 DVDD.n5550 0.00561579
R48117 DVDD.n15177 DVDD.n5550 0.00561579
R48118 DVDD.n15177 DVDD.n15176 0.00561579
R48119 DVDD.n15176 DVDD.n15175 0.00561579
R48120 DVDD.n15175 DVDD.n5552 0.00561579
R48121 DVDD.n15171 DVDD.n5552 0.00561579
R48122 DVDD.n15171 DVDD.n15170 0.00561579
R48123 DVDD.n15170 DVDD.n15169 0.00561579
R48124 DVDD.n15169 DVDD.n5554 0.00561579
R48125 DVDD.n15165 DVDD.n5554 0.00561579
R48126 DVDD.n15165 DVDD.n15164 0.00561579
R48127 DVDD.n15164 DVDD.n15163 0.00561579
R48128 DVDD.n15163 DVDD.n5556 0.00561579
R48129 DVDD.n15159 DVDD.n5556 0.00561579
R48130 DVDD.n15159 DVDD.n15158 0.00561579
R48131 DVDD.n15158 DVDD.n15157 0.00561579
R48132 DVDD.n15157 DVDD.n5558 0.00561579
R48133 DVDD.n15153 DVDD.n5558 0.00561579
R48134 DVDD.n15153 DVDD.n15152 0.00561579
R48135 DVDD.n15152 DVDD.n15151 0.00561579
R48136 DVDD.n15151 DVDD.n5560 0.00561579
R48137 DVDD.n18010 DVDD.n18009 0.00561579
R48138 DVDD.n17996 DVDD.n527 0.00561579
R48139 DVDD.n17993 DVDD.n527 0.00561579
R48140 DVDD.n17985 DVDD.n17984 0.00561579
R48141 DVDD.n17984 DVDD.n17983 0.00561579
R48142 DVDD.n596 DVDD.n561 0.00561579
R48143 DVDD.n608 DVDD.n588 0.00561579
R48144 DVDD.n611 DVDD.n588 0.00561579
R48145 DVDD.n625 DVDD.n624 0.00561579
R48146 DVDD.n17976 DVDD.n595 0.00561579
R48147 DVDD.n17970 DVDD.n17969 0.00561579
R48148 DVDD.n17969 DVDD.n17968 0.00561579
R48149 DVDD.n687 DVDD.n686 0.00561579
R48150 DVDD.n703 DVDD.n702 0.00561579
R48151 DVDD.n719 DVDD.n718 0.00561579
R48152 DVDD.n17961 DVDD.n682 0.00561579
R48153 DVDD.n17957 DVDD.n682 0.00561579
R48154 DVDD.n17957 DVDD.n17956 0.00561579
R48155 DVDD.n17943 DVDD.n17942 0.00561579
R48156 DVDD.n17929 DVDD.n753 0.00561579
R48157 DVDD.n17926 DVDD.n753 0.00561579
R48158 DVDD.n17914 DVDD.n17913 0.00561579
R48159 DVDD.n17904 DVDD.n17903 0.00561579
R48160 DVDD.n17903 DVDD.n17902 0.00561579
R48161 DVDD.n17902 DVDD.n776 0.00561579
R48162 DVDD.n17898 DVDD.n776 0.00561579
R48163 DVDD.n17898 DVDD.n17897 0.00561579
R48164 DVDD.n17897 DVDD.n17896 0.00561579
R48165 DVDD.n17896 DVDD.n778 0.00561579
R48166 DVDD.n17892 DVDD.n778 0.00561579
R48167 DVDD.n17892 DVDD.n17891 0.00561579
R48168 DVDD.n17891 DVDD.n17890 0.00561579
R48169 DVDD.n17890 DVDD.n781 0.00561579
R48170 DVDD.n17886 DVDD.n781 0.00561579
R48171 DVDD.n17886 DVDD.n17885 0.00561579
R48172 DVDD.n17885 DVDD.n17884 0.00561579
R48173 DVDD.n17884 DVDD.n783 0.00561579
R48174 DVDD.n17880 DVDD.n783 0.00561579
R48175 DVDD.n17880 DVDD.n17879 0.00561579
R48176 DVDD.n820 DVDD.n819 0.00561579
R48177 DVDD.n17875 DVDD.n814 0.00561579
R48178 DVDD.n17871 DVDD.n17870 0.00561579
R48179 DVDD.n17870 DVDD.n17869 0.00561579
R48180 DVDD.n17869 DVDD.n834 0.00561579
R48181 DVDD.n17865 DVDD.n834 0.00561579
R48182 DVDD.n17865 DVDD.n17864 0.00561579
R48183 DVDD.n17864 DVDD.n17863 0.00561579
R48184 DVDD.n17863 DVDD.n836 0.00561579
R48185 DVDD.n17859 DVDD.n836 0.00561579
R48186 DVDD.n17859 DVDD.n17858 0.00561579
R48187 DVDD.n17858 DVDD.n17857 0.00561579
R48188 DVDD.n17857 DVDD.n838 0.00561579
R48189 DVDD.n17853 DVDD.n838 0.00561579
R48190 DVDD.n17853 DVDD.n17852 0.00561579
R48191 DVDD.n17852 DVDD.n17851 0.00561579
R48192 DVDD.n17851 DVDD.n840 0.00561579
R48193 DVDD.n17847 DVDD.n840 0.00561579
R48194 DVDD.n17847 DVDD.n17846 0.00561579
R48195 DVDD.n17846 DVDD.n17845 0.00561579
R48196 DVDD.n17845 DVDD.n842 0.00561579
R48197 DVDD.n17841 DVDD.n842 0.00561579
R48198 DVDD.n17841 DVDD.n17840 0.00561579
R48199 DVDD.n17840 DVDD.n17839 0.00561579
R48200 DVDD.n17839 DVDD.n844 0.00561579
R48201 DVDD.n17835 DVDD.n844 0.00561579
R48202 DVDD.n17835 DVDD.n17834 0.00561579
R48203 DVDD.n17834 DVDD.n17833 0.00561579
R48204 DVDD.n17833 DVDD.n846 0.00561579
R48205 DVDD.n17829 DVDD.n846 0.00561579
R48206 DVDD.n17829 DVDD.n17828 0.00561579
R48207 DVDD.n17828 DVDD.n17827 0.00561579
R48208 DVDD.n17827 DVDD.n848 0.00561579
R48209 DVDD.n17823 DVDD.n848 0.00561579
R48210 DVDD.n17823 DVDD.n17822 0.00561579
R48211 DVDD.n17822 DVDD.n17821 0.00561579
R48212 DVDD.n17821 DVDD.n850 0.00561579
R48213 DVDD.n17817 DVDD.n850 0.00561579
R48214 DVDD.n17817 DVDD.n17816 0.00561579
R48215 DVDD.n17816 DVDD.n17815 0.00561579
R48216 DVDD.n17815 DVDD.n852 0.00561579
R48217 DVDD.n17811 DVDD.n852 0.00561579
R48218 DVDD.n17811 DVDD.n17810 0.00561579
R48219 DVDD.n17810 DVDD.n17809 0.00561579
R48220 DVDD.n17809 DVDD.n854 0.00561579
R48221 DVDD.n17805 DVDD.n854 0.00561579
R48222 DVDD.n17805 DVDD.n17804 0.00561579
R48223 DVDD.n17804 DVDD.n17803 0.00561579
R48224 DVDD.n17803 DVDD.n856 0.00561579
R48225 DVDD.n17799 DVDD.n856 0.00561579
R48226 DVDD.n17799 DVDD.n17798 0.00561579
R48227 DVDD.n17798 DVDD.n17797 0.00561579
R48228 DVDD.n17797 DVDD.n858 0.00561579
R48229 DVDD.n17793 DVDD.n858 0.00561579
R48230 DVDD.n17793 DVDD.n17792 0.00561579
R48231 DVDD.n17792 DVDD.n17791 0.00561579
R48232 DVDD.n17791 DVDD.n860 0.00561579
R48233 DVDD.n17787 DVDD.n860 0.00561579
R48234 DVDD.n17787 DVDD.n17786 0.00561579
R48235 DVDD.n17786 DVDD.n17785 0.00561579
R48236 DVDD.n17785 DVDD.n862 0.00561579
R48237 DVDD.n17781 DVDD.n862 0.00561579
R48238 DVDD.n17781 DVDD.n17780 0.00561579
R48239 DVDD.n17780 DVDD.n17779 0.00561579
R48240 DVDD.n17779 DVDD.n864 0.00561579
R48241 DVDD.n17775 DVDD.n864 0.00561579
R48242 DVDD.n17775 DVDD.n17774 0.00561579
R48243 DVDD.n17774 DVDD.n17773 0.00561579
R48244 DVDD.n17773 DVDD.n866 0.00561579
R48245 DVDD.n17769 DVDD.n866 0.00561579
R48246 DVDD.n17769 DVDD.n17768 0.00561579
R48247 DVDD.n17768 DVDD.n17767 0.00561579
R48248 DVDD.n17767 DVDD.n868 0.00561579
R48249 DVDD.n17763 DVDD.n868 0.00561579
R48250 DVDD.n17763 DVDD.n17762 0.00561579
R48251 DVDD.n17762 DVDD.n17761 0.00561579
R48252 DVDD.n17761 DVDD.n870 0.00561579
R48253 DVDD.n17757 DVDD.n870 0.00561579
R48254 DVDD.n17757 DVDD.n17756 0.00561579
R48255 DVDD.n17756 DVDD.n17755 0.00561579
R48256 DVDD.n17755 DVDD.n872 0.00561579
R48257 DVDD.n17751 DVDD.n872 0.00561579
R48258 DVDD.n17751 DVDD.n17750 0.00561579
R48259 DVDD.n17750 DVDD.n17749 0.00561579
R48260 DVDD.n17749 DVDD.n874 0.00561579
R48261 DVDD.n17745 DVDD.n874 0.00561579
R48262 DVDD.n17745 DVDD.n17744 0.00561579
R48263 DVDD.n17744 DVDD.n17743 0.00561579
R48264 DVDD.n17743 DVDD.n876 0.00561579
R48265 DVDD.n17739 DVDD.n876 0.00561579
R48266 DVDD.n17739 DVDD.n17738 0.00561579
R48267 DVDD.n18374 DVDD.n18302 0.00561008
R48268 DVDD.n21261 DVDD.n143 0.00561008
R48269 DVDD.n18334 DVDD.n18245 0.00561008
R48270 DVDD.n4866 DVDD.n4864 0.00561008
R48271 DVDD.n20145 DVDD.n20075 0.00557857
R48272 DVDD.n20632 DVDD.n20606 0.00557857
R48273 DVDD.n3960 DVDD.n3922 0.00557857
R48274 DVDD.n9844 DVDD.n5471 0.00557857
R48275 DVDD.n19655 DVDD.n19191 0.00557857
R48276 DVDD.n3668 DVDD.n3652 0.0055625
R48277 DVDD.n4413 DVDD.n4389 0.0055625
R48278 DVDD.n5502 DVDD.n5490 0.00552105
R48279 DVDD.n822 DVDD.n810 0.00552105
R48280 DVDD.n20225 DVDD.n20027 0.00551429
R48281 DVDD.n20303 DVDD.n19845 0.00551429
R48282 DVDD.n20717 DVDD.n19145 0.00551429
R48283 DVDD.n20794 DVDD.n18874 0.00551429
R48284 DVDD.n4022 DVDD.n247 0.00551429
R48285 DVDD.n406 DVDD.n382 0.00551429
R48286 DVDD.n9913 DVDD.n9623 0.00551429
R48287 DVDD.n9982 DVDD.n9958 0.00551429
R48288 DVDD.n21175 DVDD.n18739 0.00551429
R48289 DVDD.n22288 DVDD.n60 0.00551429
R48290 DVDD.n20162 DVDD.n20071 0.00545
R48291 DVDD.n20654 DVDD.n20602 0.00545
R48292 DVDD.n3926 DVDD.n3910 0.00545
R48293 DVDD.n3640 DVDD.n3639 0.00545
R48294 DVDD.n9860 DVDD.n5475 0.00545
R48295 DVDD.n19699 DVDD.n19696 0.00545
R48296 DVDD.n5013 DVDD.n3516 0.00542632
R48297 DVDD.n5066 DVDD.n5047 0.00542632
R48298 DVDD.n5295 DVDD.n5073 0.00542632
R48299 DVDD.n5327 DVDD.n5239 0.00542632
R48300 DVDD.n5353 DVDD.n5250 0.00542632
R48301 DVDD.n5419 DVDD.n5391 0.00542632
R48302 DVDD.n5454 DVDD.n5384 0.00542632
R48303 DVDD.n18012 DVDD.n537 0.00542632
R48304 DVDD.n17980 DVDD.n17979 0.00542632
R48305 DVDD.n627 DVDD.n586 0.00542632
R48306 DVDD.n689 DVDD.n675 0.00542632
R48307 DVDD.n715 DVDD.n658 0.00542632
R48308 DVDD.n17945 DVDD.n770 0.00542632
R48309 DVDD.n17910 DVDD.n763 0.00542632
R48310 DVDD.n496 DVDD.n489 0.00539375
R48311 DVDD.n20244 DVDD.n19958 0.00538571
R48312 DVDD.n20319 DVDD.n19849 0.00538571
R48313 DVDD.n20736 DVDD.n19073 0.00538571
R48314 DVDD.n19010 DVDD.n18877 0.00538571
R48315 DVDD.n22181 DVDD.n251 0.00538571
R48316 DVDD.n427 DVDD.n387 0.00538571
R48317 DVDD.n10093 DVDD.n9626 0.00538571
R48318 DVDD.n10002 DVDD.n9963 0.00538571
R48319 DVDD.n21161 DVDD.n18743 0.00538571
R48320 DVDD.n22274 DVDD.n65 0.00538571
R48321 DVDD.n13804 DVDD.n13803 0.00537218
R48322 DVDD.n12904 DVDD.n2254 0.00537218
R48323 DVDD.n4459 DVDD.n4392 0.0053375
R48324 DVDD.n6699 DVDD.n6392 0.00533221
R48325 DVDD.n8136 DVDD.n7687 0.00533221
R48326 DVDD.n6700 DVDD.n6394 0.00533221
R48327 DVDD.n8137 DVDD.n7686 0.00533221
R48328 DVDD.n15284 DVDD.n15283 0.00533158
R48329 DVDD.n17871 DVDD.n808 0.00533158
R48330 DVDD.n3445 DVDD.n2366 0.00532927
R48331 DVDD.n15574 DVDD.n2676 0.00532927
R48332 DVDD.n3444 DVDD.n2404 0.00532927
R48333 DVDD.n15573 DVDD.n2593 0.00532927
R48334 DVDD.n3448 DVDD.n3361 0.00532927
R48335 DVDD.n15577 DVDD.n3258 0.00532927
R48336 DVDD.n3451 DVDD.n3450 0.00532927
R48337 DVDD.n15580 DVDD.n15579 0.00532927
R48338 DVDD.n20333 DVDD.n18932 0.00532143
R48339 DVDD.n20845 DVDD.n18961 0.00532143
R48340 DVDD.n22104 DVDD.n22071 0.00532143
R48341 DVDD.n10014 DVDD.n791 0.00532143
R48342 DVDD.n22317 DVDD.n18 0.00532143
R48343 DVDD.n21783 DVDD.n196 0.00530256
R48344 DVDD.n4762 DVDD.n3673 0.0053
R48345 DVDD.n21595 DVDD.n21594 0.00528537
R48346 DVDD.n18426 DVDD.n18410 0.00528537
R48347 DVDD.n21650 DVDD.n21646 0.00528537
R48348 DVDD.n21441 DVDD.n18552 0.00528537
R48349 DVDD.n18084 DVDD.n18063 0.00528125
R48350 DVDD.n20045 DVDD.n19726 0.00525714
R48351 DVDD.n20273 DVDD.n19887 0.00525714
R48352 DVDD.n19167 DVDD.n18833 0.00525714
R48353 DVDD.n20765 DVDD.n19037 0.00525714
R48354 DVDD.n4002 DVDD.n3864 0.00525714
R48355 DVDD.n346 DVDD.n294 0.00525714
R48356 DVDD.n9895 DVDD.n9758 0.00525714
R48357 DVDD.n9718 DVDD.n9683 0.00525714
R48358 DVDD.n18717 DVDD.n18676 0.00525714
R48359 DVDD.n21134 DVDD.n108 0.00525714
R48360 DVDD.n16396 DVDD.n16395 0.00524146
R48361 DVDD.n2475 DVDD.n2393 0.00524146
R48362 DVDD.n3396 DVDD.n3351 0.00524146
R48363 DVDD.n3488 DVDD.n3423 0.00524146
R48364 DVDD.n5305 DVDD.n5076 0.00523684
R48365 DVDD.n5077 DVDD.n5054 0.00523684
R48366 DVDD.n5337 DVDD.n5236 0.00523684
R48367 DVDD.n5343 DVDD.n5247 0.00523684
R48368 DVDD.n15409 DVDD.n5376 0.00523684
R48369 DVDD.n17977 DVDD.n594 0.00523684
R48370 DVDD.n17972 DVDD.n584 0.00523684
R48371 DVDD.n699 DVDD.n660 0.00523684
R48372 DVDD.n705 DVDD.n673 0.00523684
R48373 DVDD.n17955 DVDD.n738 0.00523684
R48374 DVDD.n18413 DVDD.n18397 0.005225
R48375 DVDD.n22022 DVDD.n22010 0.005225
R48376 DVDD.n21342 DVDD.n18553 0.005225
R48377 DVDD.n21694 DVDD.n18525 0.005225
R48378 DVDD.n18253 DVDD.n18216 0.005225
R48379 DVDD.n18438 DVDD.n18437 0.005225
R48380 DVDD.n4275 DVDD.n4245 0.005225
R48381 DVDD.n4292 DVDD.n4289 0.005225
R48382 DVDD.n3683 DVDD.n3682 0.005225
R48383 DVDD.n4559 DVDD.n4558 0.005225
R48384 DVDD.n10590 DVDD.n10589 0.005225
R48385 DVDD.n21941 DVDD.n18385 0.00520651
R48386 DVDD.n22230 DVDD.n134 0.00520651
R48387 DVDD.n21921 DVDD.n21920 0.00520651
R48388 DVDD.n18113 DVDD.n18097 0.00520651
R48389 DVDD.n20357 DVDD.n18936 0.00519286
R48390 DVDD.n19003 DVDD.n18965 0.00519286
R48391 DVDD.n22123 DVDD.n440 0.00519286
R48392 DVDD.n10040 DVDD.n785 0.00519286
R48393 DVDD.n34 DVDD.n14 0.00519286
R48394 DVDD.n3603 DVDD.n3527 0.00516875
R48395 DVDD.n21676 DVDD.n196 0.00515817
R48396 DVDD.n22193 DVDD.n208 0.00515817
R48397 DVDD.n21721 DVDD.n18434 0.00515817
R48398 DVDD.n4861 DVDD.n4860 0.00515817
R48399 DVDD.n5512 DVDD.n5487 0.00514211
R48400 DVDD.n17876 DVDD.n813 0.00514211
R48401 DVDD.n20182 DVDD.n19730 0.00512857
R48402 DVDD.n20257 DVDD.n19891 0.00512857
R48403 DVDD.n20674 DVDD.n18837 0.00512857
R48404 DVDD.n20749 DVDD.n19045 0.00512857
R48405 DVDD.n3997 DVDD.n3868 0.00512857
R48406 DVDD.n22160 DVDD.n290 0.00512857
R48407 DVDD.n9823 DVDD.n9762 0.00512857
R48408 DVDD.n10069 DVDD.n9661 0.00512857
R48409 DVDD.n19676 DVDD.n18683 0.00512857
R48410 DVDD.n22251 DVDD.n118 0.00512857
R48411 DVDD.n4434 DVDD.n3749 0.0051125
R48412 DVDD.n3616 DVDD.n3531 0.00505625
R48413 DVDD.n5019 DVDD.n4888 0.00504737
R48414 DVDD.n5266 DVDD.n5064 0.00504737
R48415 DVDD.n5289 DVDD.n5058 0.00504737
R48416 DVDD.n5321 DVDD.n5243 0.00504737
R48417 DVDD.n5359 DVDD.n5232 0.00504737
R48418 DVDD.n5425 DVDD.n5398 0.00504737
R48419 DVDD.n5448 DVDD.n5404 0.00504737
R48420 DVDD.n18006 DVDD.n524 0.00504737
R48421 DVDD.n598 DVDD.n574 0.00504737
R48422 DVDD.n621 DVDD.n571 0.00504737
R48423 DVDD.n683 DVDD.n676 0.00504737
R48424 DVDD.n721 DVDD.n666 0.00504737
R48425 DVDD.n17939 DVDD.n750 0.00504737
R48426 DVDD.n17916 DVDD.n756 0.00504737
R48427 DVDD.n15103 DVDD.n6347 0.00501965
R48428 DVDD.n15104 DVDD.n6345 0.00501965
R48429 DVDD.n20051 DVDD.n19730 0.005
R48430 DVDD.n20255 DVDD.n19891 0.005
R48431 DVDD.n19173 DVDD.n18837 0.005
R48432 DVDD.n20747 DVDD.n19045 0.005
R48433 DVDD.n3995 DVDD.n3868 0.005
R48434 DVDD.n22161 DVDD.n22160 0.005
R48435 DVDD.n4743 DVDD.n3727 0.005
R48436 DVDD.n4448 DVDD.n4415 0.005
R48437 DVDD.n9877 DVDD.n9762 0.005
R48438 DVDD.n9661 DVDD.n9657 0.005
R48439 DVDD.n19680 DVDD.n18683 0.005
R48440 DVDD.n22251 DVDD.n112 0.005
R48441 DVDD.n20123 DVDD.n20077 0.00498219
R48442 DVDD.n20128 DVDD.n20073 0.00498219
R48443 DVDD.n19747 DVDD.n19728 0.00498219
R48444 DVDD.n19746 DVDD.n19724 0.00498219
R48445 DVDD.n20024 DVDD.n19975 0.00498219
R48446 DVDD.n20029 DVDD.n19971 0.00498219
R48447 DVDD.n19937 DVDD.n19889 0.00498219
R48448 DVDD.n19942 DVDD.n19885 0.00498219
R48449 DVDD.n20373 DVDD.n19840 0.00498219
R48450 DVDD.n20372 DVDD.n19836 0.00498219
R48451 DVDD.n18952 DVDD.n18934 0.00498219
R48452 DVDD.n18951 DVDD.n18930 0.00498219
R48453 DVDD.n20610 DVDD.n20608 0.00498219
R48454 DVDD.n20615 DVDD.n20604 0.00498219
R48455 DVDD.n18841 DVDD.n18835 0.00498219
R48456 DVDD.n18865 DVDD.n18861 0.00498219
R48457 DVDD.n19142 DVDD.n19138 0.00498219
R48458 DVDD.n19147 DVDD.n19134 0.00498219
R48459 DVDD.n19047 DVDD.n19039 0.00498219
R48460 DVDD.n19052 DVDD.n19035 0.00498219
R48461 DVDD.n18895 DVDD.n18886 0.00498219
R48462 DVDD.n18894 DVDD.n18880 0.00498219
R48463 DVDD.n18980 DVDD.n18963 0.00498219
R48464 DVDD.n20852 DVDD.n18972 0.00498219
R48465 DVDD.n3965 DVDD.n3933 0.00498219
R48466 DVDD.n3928 DVDD.n3924 0.00498219
R48467 DVDD.n3897 DVDD.n3866 0.00498219
R48468 DVDD.n3893 DVDD.n3875 0.00498219
R48469 DVDD.n259 DVDD.n241 0.00498219
R48470 DVDD.n22178 DVDD.n268 0.00498219
R48471 DVDD.n322 DVDD.n296 0.00498219
R48472 DVDD.n321 DVDD.n292 0.00498219
R48473 DVDD.n379 DVDD.n378 0.00498219
R48474 DVDD.n384 DVDD.n374 0.00498219
R48475 DVDD.n22075 DVDD.n22073 0.00498219
R48476 DVDD.n22115 DVDD.n22080 0.00498219
R48477 DVDD.n5484 DVDD.n5469 0.00498219
R48478 DVDD.n5479 DVDD.n5473 0.00498219
R48479 DVDD.n9766 DVDD.n9760 0.00498219
R48480 DVDD.n9771 DVDD.n9757 0.00498219
R48481 DVDD.n9641 DVDD.n9618 0.00498219
R48482 DVDD.n9648 DVDD.n9614 0.00498219
R48483 DVDD.n9688 DVDD.n9685 0.00498219
R48484 DVDD.n9693 DVDD.n9681 0.00498219
R48485 DVDD.n9955 DVDD.n9755 0.00498219
R48486 DVDD.n9960 DVDD.n9751 0.00498219
R48487 DVDD.n807 DVDD.n787 0.00498219
R48488 DVDD.n806 DVDD.n789 0.00498219
R48489 DVDD.n9689 DVDD.n9688 0.00498219
R48490 DVDD.n9694 DVDD.n9693 0.00498219
R48491 DVDD.n323 DVDD.n296 0.00498219
R48492 DVDD.n22156 DVDD.n292 0.00498219
R48493 DVDD.n19048 DVDD.n19047 0.00498219
R48494 DVDD.n19053 DVDD.n19052 0.00498219
R48495 DVDD.n19938 DVDD.n19937 0.00498219
R48496 DVDD.n19943 DVDD.n19942 0.00498219
R48497 DVDD.n9956 DVDD.n9955 0.00498219
R48498 DVDD.n9961 DVDD.n9960 0.00498219
R48499 DVDD.n380 DVDD.n379 0.00498219
R48500 DVDD.n385 DVDD.n384 0.00498219
R48501 DVDD.n18895 DVDD.n18872 0.00498219
R48502 DVDD.n18894 DVDD.n18879 0.00498219
R48503 DVDD.n20373 DVDD.n19843 0.00498219
R48504 DVDD.n20372 DVDD.n19847 0.00498219
R48505 DVDD.n9642 DVDD.n9618 0.00498219
R48506 DVDD.n10091 DVDD.n9614 0.00498219
R48507 DVDD.n259 DVDD.n245 0.00498219
R48508 DVDD.n268 DVDD.n249 0.00498219
R48509 DVDD.n19143 DVDD.n19142 0.00498219
R48510 DVDD.n19148 DVDD.n19147 0.00498219
R48511 DVDD.n20025 DVDD.n20024 0.00498219
R48512 DVDD.n20030 DVDD.n20029 0.00498219
R48513 DVDD.n3929 DVDD.n3928 0.00498219
R48514 DVDD.n3940 DVDD.n3933 0.00498219
R48515 DVDD.n5480 DVDD.n5479 0.00498219
R48516 DVDD.n5485 DVDD.n5484 0.00498219
R48517 DVDD.n20611 DVDD.n20610 0.00498219
R48518 DVDD.n20616 DVDD.n20615 0.00498219
R48519 DVDD.n20124 DVDD.n20123 0.00498219
R48520 DVDD.n20129 DVDD.n20128 0.00498219
R48521 DVDD.n807 DVDD.n798 0.00498219
R48522 DVDD.n806 DVDD.n795 0.00498219
R48523 DVDD.n22076 DVDD.n22075 0.00498219
R48524 DVDD.n22086 DVDD.n22080 0.00498219
R48525 DVDD.n18980 DVDD.n18968 0.00498219
R48526 DVDD.n18989 DVDD.n18972 0.00498219
R48527 DVDD.n18952 DVDD.n18940 0.00498219
R48528 DVDD.n18951 DVDD.n18944 0.00498219
R48529 DVDD.n9767 DVDD.n9766 0.00498219
R48530 DVDD.n9772 DVDD.n9771 0.00498219
R48531 DVDD.n4063 DVDD.n3866 0.00498219
R48532 DVDD.n3894 DVDD.n3893 0.00498219
R48533 DVDD.n18842 DVDD.n18841 0.00498219
R48534 DVDD.n18861 DVDD.n18846 0.00498219
R48535 DVDD.n19747 DVDD.n19735 0.00498219
R48536 DVDD.n19746 DVDD.n19739 0.00498219
R48537 DVDD.n19209 DVDD.n19193 0.00498219
R48538 DVDD.n19208 DVDD.n19189 0.00498219
R48539 DVDD.n21211 DVDD.n18680 0.00498219
R48540 DVDD.n18708 DVDD.n18673 0.00498219
R48541 DVDD.n21099 DVDD.n21098 0.00498219
R48542 DVDD.n21094 DVDD.n21089 0.00498219
R48543 DVDD.n120 DVDD.n110 0.00498219
R48544 DVDD.n119 DVDD.n106 0.00498219
R48545 DVDD.n78 DVDD.n77 0.00498219
R48546 DVDD.n73 DVDD.n72 0.00498219
R48547 DVDD.n22336 DVDD.n16 0.00498219
R48548 DVDD.n22344 DVDD.n5 0.00498219
R48549 DVDD.n18700 DVDD.n18680 0.00498219
R48550 DVDD.n18701 DVDD.n18673 0.00498219
R48551 DVDD.n21098 DVDD.n18737 0.00498219
R48552 DVDD.n21089 DVDD.n18741 0.00498219
R48553 DVDD.n120 DVDD.n99 0.00498219
R48554 DVDD.n119 DVDD.n103 0.00498219
R48555 DVDD.n77 DVDD.n58 0.00498219
R48556 DVDD.n72 DVDD.n62 0.00498219
R48557 DVDD.n22 DVDD.n5 0.00498219
R48558 DVDD.n22336 DVDD.n25 0.00498219
R48559 DVDD.n19209 DVDD.n19195 0.00498219
R48560 DVDD.n19208 DVDD.n19199 0.00498219
R48561 DVDD.n3434 DVDD.n2363 0.00497805
R48562 DVDD.n15565 DVDD.n2672 0.00497805
R48563 DVDD.n3433 DVDD.n2402 0.00497805
R48564 DVDD.n15564 DVDD.n2591 0.00497805
R48565 DVDD.n3437 DVDD.n3359 0.00497805
R48566 DVDD.n15568 DVDD.n3256 0.00497805
R48567 DVDD.n3440 DVDD.n3439 0.00497805
R48568 DVDD.n15571 DVDD.n15570 0.00497805
R48569 DVDD.n5492 DVDD.n5476 0.00495263
R48570 DVDD.n816 DVDD.n802 0.00495263
R48571 DVDD.n3611 DVDD.n3523 0.00494375
R48572 DVDD.n20327 DVDD.n18936 0.00493571
R48573 DVDD.n20827 DVDD.n18965 0.00493571
R48574 DVDD.n440 DVDD.n439 0.00493571
R48575 DVDD.n805 DVDD.n785 0.00493571
R48576 DVDD.n22335 DVDD.n14 0.00493571
R48577 DVDD.n18131 DVDD.n493 0.004925
R48578 DVDD.n2896 DVDD.n761 0.00488868
R48579 DVDD.n15326 DVDD.n15324 0.00488868
R48580 DVDD.n15457 DVDD.n15424 0.00488868
R48581 DVDD.n16215 DVDD.n16213 0.00488868
R48582 DVDD.n5088 DVDD.n5053 0.00488868
R48583 DVDD.n16336 DVDD.n16334 0.00488868
R48584 DVDD.n15748 DVDD.n15715 0.00488868
R48585 DVDD.n2540 DVDD.n530 0.00488868
R48586 DVDD.n4429 DVDD.n3736 0.0048875
R48587 DVDD.n20195 DVDD.n19726 0.00487143
R48588 DVDD.n20271 DVDD.n19887 0.00487143
R48589 DVDD.n20687 DVDD.n18833 0.00487143
R48590 DVDD.n19061 DVDD.n19037 0.00487143
R48591 DVDD.n4052 DVDD.n3864 0.00487143
R48592 DVDD.n344 DVDD.n294 0.00487143
R48593 DVDD.n9893 DVDD.n9758 0.00487143
R48594 DVDD.n9716 DVDD.n9683 0.00487143
R48595 DVDD.n21202 DVDD.n18676 0.00487143
R48596 DVDD.n21136 DVDD.n108 0.00487143
R48597 DVDD.n5027 DVDD.n3513 0.00485789
R48598 DVDD.n5034 DVDD.n3512 0.00485789
R48599 DVDD.n5274 DVDD.n5069 0.00485789
R48600 DVDD.n5281 DVDD.n5070 0.00485789
R48601 DVDD.n15460 DVDD.n5253 0.00485789
R48602 DVDD.n5433 DVDD.n5388 0.00485789
R48603 DVDD.n5440 DVDD.n5387 0.00485789
R48604 DVDD.n17998 DVDD.n534 0.00485789
R48605 DVDD.n17991 DVDD.n533 0.00485789
R48606 DVDD.n606 DVDD.n591 0.00485789
R48607 DVDD.n613 DVDD.n576 0.00485789
R48608 DVDD.n17962 DVDD.n681 0.00485789
R48609 DVDD.n17931 DVDD.n767 0.00485789
R48610 DVDD.n17924 DVDD.n766 0.00485789
R48611 DVDD.n13801 DVDD.n11226 0.00484899
R48612 DVDD.n12910 DVDD.n12909 0.00484899
R48613 DVDD.n13802 DVDD.n11228 0.00484899
R48614 DVDD.n16455 DVDD.n2255 0.00484899
R48615 DVDD.n3626 DVDD.n3526 0.00483125
R48616 DVDD.n14016 DVDD.n10706 0.00483083
R48617 DVDD.n16742 DVDD.n1801 0.00483083
R48618 DVDD.n20344 DVDD.n18932 0.00480714
R48619 DVDD.n20843 DVDD.n18961 0.00480714
R48620 DVDD.n22102 DVDD.n22071 0.00480714
R48621 DVDD.n10027 DVDD.n791 0.00480714
R48622 DVDD.n22319 DVDD.n18 0.00480714
R48623 DVDD.n21722 DVDD.n21721 0.00479029
R48624 DVDD.n22193 DVDD.n213 0.00479029
R48625 DVDD.n21773 DVDD.n196 0.00479029
R48626 DVDD.n18117 DVDD.n18068 0.00479029
R48627 DVDD.n4420 DVDD.n4419 0.004775
R48628 DVDD.n4597 DVDD.n4271 0.004775
R48629 DVDD.n13749 DVDD.n13748 0.004775
R48630 DVDD.n16709 DVDD.n16708 0.004775
R48631 DVDD.n5504 DVDD.n5493 0.00476316
R48632 DVDD.n824 DVDD.n803 0.00476316
R48633 DVDD.n21231 DVDD.n21225 0.00476
R48634 DVDD.n21231 DVDD.n21227 0.00476
R48635 DVDD.n21227 DVDD.n21226 0.00476
R48636 DVDD.n18547 DVDD.n18546 0.00476
R48637 DVDD.n21656 DVDD.n18547 0.00476
R48638 DVDD.n21656 DVDD.n18543 0.00476
R48639 DVDD.n21660 DVDD.n18543 0.00476
R48640 DVDD.n21663 DVDD.n21661 0.00476
R48641 DVDD.n21663 DVDD.n18541 0.00476
R48642 DVDD.n21668 DVDD.n18541 0.00476
R48643 DVDD.n21668 DVDD.n185 0.00476
R48644 DVDD.n18322 DVDD.n186 0.00476
R48645 DVDD.n18325 DVDD.n18322 0.00476
R48646 DVDD.n18325 DVDD.n18318 0.00476
R48647 DVDD.n18361 DVDD.n18318 0.00476
R48648 DVDD.n18357 DVDD.n18319 0.00476
R48649 DVDD.n18357 DVDD.n18356 0.00476
R48650 DVDD.n18356 DVDD.n18355 0.00476
R48651 DVDD.n18355 DVDD.n18353 0.00476
R48652 DVDD.n22191 DVDD.n22190 0.00476
R48653 DVDD.n22190 DVDD.n22189 0.00476
R48654 DVDD.n22189 DVDD.n227 0.00476
R48655 DVDD.n21252 DVDD.n18667 0.00476
R48656 DVDD.n21252 DVDD.n18669 0.00476
R48657 DVDD.n18669 DVDD.n18668 0.00476
R48658 DVDD.n21719 DVDD.n21718 0.00476
R48659 DVDD.n21718 DVDD.n21717 0.00476
R48660 DVDD.n21717 DVDD.n18511 0.00476
R48661 DVDD.n21713 DVDD.n18511 0.00476
R48662 DVDD.n21712 DVDD.n21711 0.00476
R48663 DVDD.n21711 DVDD.n18516 0.00476
R48664 DVDD.n21707 DVDD.n18516 0.00476
R48665 DVDD.n21707 DVDD.n193 0.00476
R48666 DVDD.n22208 DVDD.n195 0.00476
R48667 DVDD.n22204 DVDD.n195 0.00476
R48668 DVDD.n22204 DVDD.n22203 0.00476
R48669 DVDD.n22203 DVDD.n22202 0.00476
R48670 DVDD.n22198 DVDD.n201 0.00476
R48671 DVDD.n22198 DVDD.n22197 0.00476
R48672 DVDD.n22197 DVDD.n22196 0.00476
R48673 DVDD.n22196 DVDD.n206 0.00476
R48674 DVDD.n22026 DVDD.n22025 0.00476
R48675 DVDD.n22031 DVDD.n22026 0.00476
R48676 DVDD.n22031 DVDD.n22028 0.00476
R48677 DVDD.n18456 DVDD.n18454 0.00476
R48678 DVDD.n18500 DVDD.n18456 0.00476
R48679 DVDD.n18501 DVDD.n18500 0.00476
R48680 DVDD.n18451 DVDD.n167 0.00476
R48681 DVDD.n22221 DVDD.n167 0.00476
R48682 DVDD.n22221 DVDD.n168 0.00476
R48683 DVDD.n22217 DVDD.n168 0.00476
R48684 DVDD.n22216 DVDD.n22215 0.00476
R48685 DVDD.n22215 DVDD.n174 0.00476
R48686 DVDD.n22211 DVDD.n174 0.00476
R48687 DVDD.n22211 DVDD.n22210 0.00476
R48688 DVDD.n21881 DVDD.n181 0.00476
R48689 DVDD.n21881 DVDD.n21835 0.00476
R48690 DVDD.n21885 DVDD.n21835 0.00476
R48691 DVDD.n21886 DVDD.n21885 0.00476
R48692 DVDD.n21889 DVDD.n21831 0.00476
R48693 DVDD.n21894 DVDD.n21831 0.00476
R48694 DVDD.n21894 DVDD.n21833 0.00476
R48695 DVDD.n21833 DVDD.n21832 0.00476
R48696 DVDD.n18238 DVDD.n18232 0.00476
R48697 DVDD.n18238 DVDD.n18233 0.00476
R48698 DVDD.n18234 DVDD.n18233 0.00476
R48699 DVDD.n18491 DVDD.n18486 0.00476
R48700 DVDD.n18491 DVDD.n18490 0.00476
R48701 DVDD.n18490 DVDD.n18489 0.00476
R48702 DVDD.n21586 DVDD.n21584 0.00476
R48703 DVDD.n21589 DVDD.n21586 0.00476
R48704 DVDD.n21589 DVDD.n18407 0.00476
R48705 DVDD.n21741 DVDD.n18407 0.00476
R48706 DVDD.n21751 DVDD.n18405 0.00476
R48707 DVDD.n21751 DVDD.n21750 0.00476
R48708 DVDD.n21750 DVDD.n21748 0.00476
R48709 DVDD.n21748 DVDD.n189 0.00476
R48710 DVDD.n21868 DVDD.n188 0.00476
R48711 DVDD.n21868 DVDD.n21861 0.00476
R48712 DVDD.n21872 DVDD.n21861 0.00476
R48713 DVDD.n21872 DVDD.n21807 0.00476
R48714 DVDD.n21904 DVDD.n21805 0.00476
R48715 DVDD.n21911 DVDD.n21805 0.00476
R48716 DVDD.n21911 DVDD.n21910 0.00476
R48717 DVDD.n21910 DVDD.n21909 0.00476
R48718 DVDD.n18226 DVDD.n18223 0.00476
R48719 DVDD.n22053 DVDD.n18223 0.00476
R48720 DVDD.n22053 DVDD.n18221 0.00476
R48721 DVDD.n3597 DVDD.n3596 0.00476
R48722 DVDD.n4107 DVDD.n4106 0.00476
R48723 DVDD.n4108 DVDD.n4107 0.00476
R48724 DVDD.n4145 DVDD.n3823 0.00476
R48725 DVDD.n4146 DVDD.n4145 0.00476
R48726 DVDD.n4147 DVDD.n4146 0.00476
R48727 DVDD.n4181 DVDD.n4180 0.00476
R48728 DVDD.n4184 DVDD.n4181 0.00476
R48729 DVDD.n4185 DVDD.n4184 0.00476
R48730 DVDD.n4186 DVDD.n4185 0.00476
R48731 DVDD.n4187 DVDD.n4186 0.00476
R48732 DVDD.n4209 DVDD.n4208 0.00476
R48733 DVDD.n4210 DVDD.n4209 0.00476
R48734 DVDD.n4632 DVDD.n4210 0.00476
R48735 DVDD.n4661 DVDD.n4660 0.00476
R48736 DVDD.n4661 DVDD.n487 0.00476
R48737 DVDD.n18136 DVDD.n18135 0.00476
R48738 DVDD.n4802 DVDD.n4801 0.00476
R48739 DVDD.n4801 DVDD.n3581 0.00476
R48740 DVDD.n4797 DVDD.n3581 0.00476
R48741 DVDD.n4797 DVDD.n4796 0.00476
R48742 DVDD.n4796 DVDD.n4795 0.00476
R48743 DVDD.n4795 DVDD.n3587 0.00476
R48744 DVDD.n4791 DVDD.n3587 0.00476
R48745 DVDD.n4791 DVDD.n4790 0.00476
R48746 DVDD.n4790 DVDD.n4789 0.00476
R48747 DVDD.n4789 DVDD.n3593 0.00476
R48748 DVDD.n4785 DVDD.n3593 0.00476
R48749 DVDD.n4785 DVDD.n4784 0.00476
R48750 DVDD.n4784 DVDD.n4783 0.00476
R48751 DVDD.n4105 DVDD.n4104 0.00476
R48752 DVDD.n4109 DVDD.n4104 0.00476
R48753 DVDD.n4111 DVDD.n4109 0.00476
R48754 DVDD.n4111 DVDD.n4100 0.00476
R48755 DVDD.n4115 DVDD.n4100 0.00476
R48756 DVDD.n4117 DVDD.n4115 0.00476
R48757 DVDD.n4119 DVDD.n4117 0.00476
R48758 DVDD.n4119 DVDD.n4096 0.00476
R48759 DVDD.n4123 DVDD.n4096 0.00476
R48760 DVDD.n4125 DVDD.n4123 0.00476
R48761 DVDD.n4127 DVDD.n4125 0.00476
R48762 DVDD.n4127 DVDD.n4093 0.00476
R48763 DVDD.n4131 DVDD.n4093 0.00476
R48764 DVDD.n4131 DVDD.n3826 0.00476
R48765 DVDD.n4139 DVDD.n3826 0.00476
R48766 DVDD.n4139 DVDD.n3824 0.00476
R48767 DVDD.n4144 DVDD.n3824 0.00476
R48768 DVDD.n4144 DVDD.n3822 0.00476
R48769 DVDD.n4148 DVDD.n3822 0.00476
R48770 DVDD.n4150 DVDD.n4148 0.00476
R48771 DVDD.n4150 DVDD.n3819 0.00476
R48772 DVDD.n4154 DVDD.n3819 0.00476
R48773 DVDD.n4155 DVDD.n4154 0.00476
R48774 DVDD.n4734 DVDD.n4733 0.00476
R48775 DVDD.n4733 DVDD.n4732 0.00476
R48776 DVDD.n4732 DVDD.n3764 0.00476
R48777 DVDD.n4728 DVDD.n3764 0.00476
R48778 DVDD.n4728 DVDD.n4727 0.00476
R48779 DVDD.n4727 DVDD.n4726 0.00476
R48780 DVDD.n4726 DVDD.n3769 0.00476
R48781 DVDD.n4722 DVDD.n3769 0.00476
R48782 DVDD.n4722 DVDD.n4721 0.00476
R48783 DVDD.n4721 DVDD.n4720 0.00476
R48784 DVDD.n4720 DVDD.n4182 0.00476
R48785 DVDD.n4716 DVDD.n4182 0.00476
R48786 DVDD.n4716 DVDD.n4715 0.00476
R48787 DVDD.n4715 DVDD.n4714 0.00476
R48788 DVDD.n4714 DVDD.n4188 0.00476
R48789 DVDD.n4710 DVDD.n4188 0.00476
R48790 DVDD.n4710 DVDD.n4709 0.00476
R48791 DVDD.n4709 DVDD.n4708 0.00476
R48792 DVDD.n4708 DVDD.n4193 0.00476
R48793 DVDD.n4704 DVDD.n4193 0.00476
R48794 DVDD.n4704 DVDD.n4703 0.00476
R48795 DVDD.n4703 DVDD.n4702 0.00476
R48796 DVDD.n4702 DVDD.n4198 0.00476
R48797 DVDD.n4697 DVDD.n4696 0.00476
R48798 DVDD.n4696 DVDD.n4695 0.00476
R48799 DVDD.n4695 DVDD.n4206 0.00476
R48800 DVDD.n4691 DVDD.n4206 0.00476
R48801 DVDD.n4691 DVDD.n4690 0.00476
R48802 DVDD.n4690 DVDD.n4689 0.00476
R48803 DVDD.n4689 DVDD.n4211 0.00476
R48804 DVDD.n4685 DVDD.n4211 0.00476
R48805 DVDD.n4685 DVDD.n4684 0.00476
R48806 DVDD.n4684 DVDD.n4683 0.00476
R48807 DVDD.n4683 DVDD.n4216 0.00476
R48808 DVDD.n4679 DVDD.n4216 0.00476
R48809 DVDD.n4679 DVDD.n4678 0.00476
R48810 DVDD.n4678 DVDD.n4677 0.00476
R48811 DVDD.n4677 DVDD.n4221 0.00476
R48812 DVDD.n4673 DVDD.n4221 0.00476
R48813 DVDD.n4673 DVDD.n4672 0.00476
R48814 DVDD.n4672 DVDD.n4671 0.00476
R48815 DVDD.n4671 DVDD.n4226 0.00476
R48816 DVDD.n4667 DVDD.n4226 0.00476
R48817 DVDD.n4667 DVDD.n4666 0.00476
R48818 DVDD.n4666 DVDD.n4665 0.00476
R48819 DVDD.n4665 DVDD.n4662 0.00476
R48820 DVDD.n18137 DVDD.n486 0.00476
R48821 DVDD.n18139 DVDD.n18137 0.00476
R48822 DVDD.n18139 DVDD.n483 0.00476
R48823 DVDD.n18143 DVDD.n483 0.00476
R48824 DVDD.n18145 DVDD.n18143 0.00476
R48825 DVDD.n18147 DVDD.n18145 0.00476
R48826 DVDD.n18147 DVDD.n479 0.00476
R48827 DVDD.n18151 DVDD.n479 0.00476
R48828 DVDD.n18153 DVDD.n18151 0.00476
R48829 DVDD.n18155 DVDD.n18153 0.00476
R48830 DVDD.n18160 DVDD.n18158 0.00476
R48831 DVDD.n18161 DVDD.n18160 0.00476
R48832 DVDD.n15328 DVDD.n15326 0.00476
R48833 DVDD.n15330 DVDD.n15328 0.00476
R48834 DVDD.n15330 DVDD.n15322 0.00476
R48835 DVDD.n15335 DVDD.n15322 0.00476
R48836 DVDD.n15337 DVDD.n15335 0.00476
R48837 DVDD.n15339 DVDD.n15337 0.00476
R48838 DVDD.n15339 DVDD.n15319 0.00476
R48839 DVDD.n15404 DVDD.n15319 0.00476
R48840 DVDD.n15404 DVDD.n15403 0.00476
R48841 DVDD.n15403 DVDD.n15401 0.00476
R48842 DVDD.n15401 DVDD.n15399 0.00476
R48843 DVDD.n15399 DVDD.n15398 0.00476
R48844 DVDD.n15398 DVDD.n15397 0.00476
R48845 DVDD.n15393 DVDD.n15392 0.00476
R48846 DVDD.n15392 DVDD.n15391 0.00476
R48847 DVDD.n15391 DVDD.n15389 0.00476
R48848 DVDD.n15389 DVDD.n15387 0.00476
R48849 DVDD.n15387 DVDD.n15385 0.00476
R48850 DVDD.n15385 DVDD.n15383 0.00476
R48851 DVDD.n15383 DVDD.n15381 0.00476
R48852 DVDD.n15381 DVDD.n15379 0.00476
R48853 DVDD.n15379 DVDD.n15377 0.00476
R48854 DVDD.n15377 DVDD.n15375 0.00476
R48855 DVDD.n15375 DVDD.n15373 0.00476
R48856 DVDD.n15373 DVDD.n15371 0.00476
R48857 DVDD.n15371 DVDD.n15369 0.00476
R48858 DVDD.n15369 DVDD.n15367 0.00476
R48859 DVDD.n15367 DVDD.n3138 0.00476
R48860 DVDD.n16005 DVDD.n3138 0.00476
R48861 DVDD.n16005 DVDD.n16004 0.00476
R48862 DVDD.n16004 DVDD.n16003 0.00476
R48863 DVDD.n16003 DVDD.n16000 0.00476
R48864 DVDD.n16000 DVDD.n15999 0.00476
R48865 DVDD.n15999 DVDD.n15997 0.00476
R48866 DVDD.n15997 DVDD.n15995 0.00476
R48867 DVDD.n15995 DVDD.n15993 0.00476
R48868 DVDD.n3224 DVDD.n3222 0.00476
R48869 DVDD.n3222 DVDD.n3220 0.00476
R48870 DVDD.n3220 DVDD.n3218 0.00476
R48871 DVDD.n3218 DVDD.n3216 0.00476
R48872 DVDD.n3216 DVDD.n3214 0.00476
R48873 DVDD.n3214 DVDD.n3056 0.00476
R48874 DVDD.n16087 DVDD.n3056 0.00476
R48875 DVDD.n16087 DVDD.n3054 0.00476
R48876 DVDD.n16091 DVDD.n3054 0.00476
R48877 DVDD.n16091 DVDD.n3052 0.00476
R48878 DVDD.n16095 DVDD.n3052 0.00476
R48879 DVDD.n16095 DVDD.n3050 0.00476
R48880 DVDD.n16100 DVDD.n3050 0.00476
R48881 DVDD.n16100 DVDD.n3047 0.00476
R48882 DVDD.n16115 DVDD.n3047 0.00476
R48883 DVDD.n16117 DVDD.n16115 0.00476
R48884 DVDD.n16119 DVDD.n16117 0.00476
R48885 DVDD.n16119 DVDD.n3045 0.00476
R48886 DVDD.n16124 DVDD.n3045 0.00476
R48887 DVDD.n16126 DVDD.n16124 0.00476
R48888 DVDD.n16128 DVDD.n16126 0.00476
R48889 DVDD.n16128 DVDD.n3042 0.00476
R48890 DVDD.n16133 DVDD.n3042 0.00476
R48891 DVDD.n16139 DVDD.n16136 0.00476
R48892 DVDD.n16139 DVDD.n2994 0.00476
R48893 DVDD.n16146 DVDD.n2994 0.00476
R48894 DVDD.n16146 DVDD.n2992 0.00476
R48895 DVDD.n16151 DVDD.n2992 0.00476
R48896 DVDD.n16151 DVDD.n2990 0.00476
R48897 DVDD.n16155 DVDD.n2990 0.00476
R48898 DVDD.n16157 DVDD.n16155 0.00476
R48899 DVDD.n16157 DVDD.n2988 0.00476
R48900 DVDD.n16162 DVDD.n2988 0.00476
R48901 DVDD.n16164 DVDD.n16162 0.00476
R48902 DVDD.n16166 DVDD.n16164 0.00476
R48903 DVDD.n16166 DVDD.n2985 0.00476
R48904 DVDD.n16171 DVDD.n2985 0.00476
R48905 DVDD.n16173 DVDD.n16171 0.00476
R48906 DVDD.n16175 DVDD.n16173 0.00476
R48907 DVDD.n16175 DVDD.n2982 0.00476
R48908 DVDD.n16179 DVDD.n2982 0.00476
R48909 DVDD.n16179 DVDD.n2923 0.00476
R48910 DVDD.n16186 DVDD.n2923 0.00476
R48911 DVDD.n16186 DVDD.n2921 0.00476
R48912 DVDD.n16192 DVDD.n2921 0.00476
R48913 DVDD.n16192 DVDD.n2882 0.00476
R48914 DVDD.n16198 DVDD.n2919 0.00476
R48915 DVDD.n2919 DVDD.n2918 0.00476
R48916 DVDD.n2918 DVDD.n2916 0.00476
R48917 DVDD.n2916 DVDD.n2914 0.00476
R48918 DVDD.n2914 DVDD.n2912 0.00476
R48919 DVDD.n2912 DVDD.n2910 0.00476
R48920 DVDD.n2910 DVDD.n2908 0.00476
R48921 DVDD.n2908 DVDD.n2906 0.00476
R48922 DVDD.n2906 DVDD.n2904 0.00476
R48923 DVDD.n2904 DVDD.n2902 0.00476
R48924 DVDD.n2900 DVDD.n2898 0.00476
R48925 DVDD.n2898 DVDD.n2896 0.00476
R48926 DVDD.n15457 DVDD.n15456 0.00476
R48927 DVDD.n15456 DVDD.n15454 0.00476
R48928 DVDD.n15454 DVDD.n15452 0.00476
R48929 DVDD.n15452 DVDD.n15450 0.00476
R48930 DVDD.n15450 DVDD.n15448 0.00476
R48931 DVDD.n15448 DVDD.n15446 0.00476
R48932 DVDD.n15446 DVDD.n15444 0.00476
R48933 DVDD.n15444 DVDD.n15442 0.00476
R48934 DVDD.n15442 DVDD.n15440 0.00476
R48935 DVDD.n15440 DVDD.n15438 0.00476
R48936 DVDD.n15438 DVDD.n15436 0.00476
R48937 DVDD.n15436 DVDD.n5228 0.00476
R48938 DVDD.n15464 DVDD.n5228 0.00476
R48939 DVDD.n15469 DVDD.n5223 0.00476
R48940 DVDD.n15473 DVDD.n5223 0.00476
R48941 DVDD.n15475 DVDD.n15473 0.00476
R48942 DVDD.n15477 DVDD.n15475 0.00476
R48943 DVDD.n15477 DVDD.n5221 0.00476
R48944 DVDD.n15482 DVDD.n5221 0.00476
R48945 DVDD.n15484 DVDD.n15482 0.00476
R48946 DVDD.n15486 DVDD.n15484 0.00476
R48947 DVDD.n15486 DVDD.n5218 0.00476
R48948 DVDD.n15491 DVDD.n5218 0.00476
R48949 DVDD.n15493 DVDD.n15491 0.00476
R48950 DVDD.n15495 DVDD.n15493 0.00476
R48951 DVDD.n15495 DVDD.n5215 0.00476
R48952 DVDD.n15518 DVDD.n5215 0.00476
R48953 DVDD.n15518 DVDD.n15517 0.00476
R48954 DVDD.n15517 DVDD.n15516 0.00476
R48955 DVDD.n15516 DVDD.n15515 0.00476
R48956 DVDD.n15515 DVDD.n15502 0.00476
R48957 DVDD.n15511 DVDD.n15502 0.00476
R48958 DVDD.n15511 DVDD.n15510 0.00476
R48959 DVDD.n15510 DVDD.n15508 0.00476
R48960 DVDD.n15508 DVDD.n3230 0.00476
R48961 DVDD.n15914 DVDD.n3230 0.00476
R48962 DVDD.n15920 DVDD.n3208 0.00476
R48963 DVDD.n15922 DVDD.n15920 0.00476
R48964 DVDD.n15924 DVDD.n15922 0.00476
R48965 DVDD.n15924 DVDD.n3206 0.00476
R48966 DVDD.n15929 DVDD.n3206 0.00476
R48967 DVDD.n15939 DVDD.n15929 0.00476
R48968 DVDD.n15941 DVDD.n15939 0.00476
R48969 DVDD.n15941 DVDD.n3203 0.00476
R48970 DVDD.n15985 DVDD.n3203 0.00476
R48971 DVDD.n15985 DVDD.n15984 0.00476
R48972 DVDD.n15984 DVDD.n15983 0.00476
R48973 DVDD.n15983 DVDD.n15947 0.00476
R48974 DVDD.n15979 DVDD.n15947 0.00476
R48975 DVDD.n15979 DVDD.n15978 0.00476
R48976 DVDD.n15978 DVDD.n15977 0.00476
R48977 DVDD.n15977 DVDD.n15975 0.00476
R48978 DVDD.n15975 DVDD.n15973 0.00476
R48979 DVDD.n15973 DVDD.n15971 0.00476
R48980 DVDD.n15971 DVDD.n15969 0.00476
R48981 DVDD.n15969 DVDD.n15967 0.00476
R48982 DVDD.n15967 DVDD.n15965 0.00476
R48983 DVDD.n15965 DVDD.n15963 0.00476
R48984 DVDD.n15963 DVDD.n15961 0.00476
R48985 DVDD.n16259 DVDD.n2709 0.00476
R48986 DVDD.n2773 DVDD.n2709 0.00476
R48987 DVDD.n2773 DVDD.n2771 0.00476
R48988 DVDD.n16253 DVDD.n2771 0.00476
R48989 DVDD.n16253 DVDD.n16252 0.00476
R48990 DVDD.n16252 DVDD.n16251 0.00476
R48991 DVDD.n16251 DVDD.n2779 0.00476
R48992 DVDD.n2842 DVDD.n2779 0.00476
R48993 DVDD.n2847 DVDD.n2842 0.00476
R48994 DVDD.n2849 DVDD.n2847 0.00476
R48995 DVDD.n2851 DVDD.n2849 0.00476
R48996 DVDD.n2851 DVDD.n2840 0.00476
R48997 DVDD.n2856 DVDD.n2840 0.00476
R48998 DVDD.n2858 DVDD.n2856 0.00476
R48999 DVDD.n2860 DVDD.n2858 0.00476
R49000 DVDD.n2860 DVDD.n2837 0.00476
R49001 DVDD.n2864 DVDD.n2837 0.00476
R49002 DVDD.n2874 DVDD.n2864 0.00476
R49003 DVDD.n2876 DVDD.n2874 0.00476
R49004 DVDD.n2876 DVDD.n2834 0.00476
R49005 DVDD.n16244 DVDD.n2834 0.00476
R49006 DVDD.n16244 DVDD.n16243 0.00476
R49007 DVDD.n16243 DVDD.n16242 0.00476
R49008 DVDD.n16239 DVDD.n16237 0.00476
R49009 DVDD.n16237 DVDD.n16236 0.00476
R49010 DVDD.n16236 DVDD.n16235 0.00476
R49011 DVDD.n16235 DVDD.n16233 0.00476
R49012 DVDD.n16233 DVDD.n16231 0.00476
R49013 DVDD.n16231 DVDD.n16229 0.00476
R49014 DVDD.n16229 DVDD.n16227 0.00476
R49015 DVDD.n16227 DVDD.n16225 0.00476
R49016 DVDD.n16225 DVDD.n16223 0.00476
R49017 DVDD.n16223 DVDD.n16221 0.00476
R49018 DVDD.n16219 DVDD.n16217 0.00476
R49019 DVDD.n16217 DVDD.n16215 0.00476
R49020 DVDD.n5090 DVDD.n5088 0.00476
R49021 DVDD.n5092 DVDD.n5090 0.00476
R49022 DVDD.n5092 DVDD.n5086 0.00476
R49023 DVDD.n5097 DVDD.n5086 0.00476
R49024 DVDD.n5099 DVDD.n5097 0.00476
R49025 DVDD.n5101 DVDD.n5099 0.00476
R49026 DVDD.n5101 DVDD.n5083 0.00476
R49027 DVDD.n15696 DVDD.n5083 0.00476
R49028 DVDD.n15696 DVDD.n15695 0.00476
R49029 DVDD.n15695 DVDD.n15693 0.00476
R49030 DVDD.n15693 DVDD.n15691 0.00476
R49031 DVDD.n15691 DVDD.n15689 0.00476
R49032 DVDD.n15689 DVDD.n5110 0.00476
R49033 DVDD.n15684 DVDD.n15683 0.00476
R49034 DVDD.n15683 DVDD.n15682 0.00476
R49035 DVDD.n15682 DVDD.n5117 0.00476
R49036 DVDD.n15632 DVDD.n5117 0.00476
R49037 DVDD.n15634 DVDD.n15632 0.00476
R49038 DVDD.n15636 DVDD.n15634 0.00476
R49039 DVDD.n15636 DVDD.n15627 0.00476
R49040 DVDD.n15641 DVDD.n15627 0.00476
R49041 DVDD.n15643 DVDD.n15641 0.00476
R49042 DVDD.n15645 DVDD.n15643 0.00476
R49043 DVDD.n15645 DVDD.n15624 0.00476
R49044 DVDD.n15650 DVDD.n15624 0.00476
R49045 DVDD.n15652 DVDD.n15650 0.00476
R49046 DVDD.n15654 DVDD.n15652 0.00476
R49047 DVDD.n15654 DVDD.n15621 0.00476
R49048 DVDD.n15676 DVDD.n15621 0.00476
R49049 DVDD.n15676 DVDD.n15675 0.00476
R49050 DVDD.n15675 DVDD.n15674 0.00476
R49051 DVDD.n15674 DVDD.n15671 0.00476
R49052 DVDD.n15671 DVDD.n15670 0.00476
R49053 DVDD.n15670 DVDD.n15668 0.00476
R49054 DVDD.n15668 DVDD.n15666 0.00476
R49055 DVDD.n15666 DVDD.n3232 0.00476
R49056 DVDD.n15911 DVDD.n3234 0.00476
R49057 DVDD.n3304 DVDD.n3234 0.00476
R49058 DVDD.n3306 DVDD.n3304 0.00476
R49059 DVDD.n3306 DVDD.n3300 0.00476
R49060 DVDD.n3311 DVDD.n3300 0.00476
R49061 DVDD.n3313 DVDD.n3311 0.00476
R49062 DVDD.n3315 DVDD.n3313 0.00476
R49063 DVDD.n3315 DVDD.n3297 0.00476
R49064 DVDD.n15905 DVDD.n3297 0.00476
R49065 DVDD.n15905 DVDD.n15904 0.00476
R49066 DVDD.n15904 DVDD.n15903 0.00476
R49067 DVDD.n15903 DVDD.n3321 0.00476
R49068 DVDD.n15899 DVDD.n3321 0.00476
R49069 DVDD.n15899 DVDD.n15898 0.00476
R49070 DVDD.n15898 DVDD.n15897 0.00476
R49071 DVDD.n15897 DVDD.n15895 0.00476
R49072 DVDD.n15895 DVDD.n15893 0.00476
R49073 DVDD.n15893 DVDD.n15891 0.00476
R49074 DVDD.n15891 DVDD.n15889 0.00476
R49075 DVDD.n15889 DVDD.n15887 0.00476
R49076 DVDD.n15887 DVDD.n15885 0.00476
R49077 DVDD.n15885 DVDD.n15883 0.00476
R49078 DVDD.n15883 DVDD.n15881 0.00476
R49079 DVDD.n16265 DVDD.n2702 0.00476
R49080 DVDD.n16265 DVDD.n2643 0.00476
R49081 DVDD.n16272 DVDD.n2643 0.00476
R49082 DVDD.n16272 DVDD.n2641 0.00476
R49083 DVDD.n16277 DVDD.n2641 0.00476
R49084 DVDD.n16277 DVDD.n2638 0.00476
R49085 DVDD.n16281 DVDD.n2638 0.00476
R49086 DVDD.n16283 DVDD.n16281 0.00476
R49087 DVDD.n16285 DVDD.n16283 0.00476
R49088 DVDD.n16285 DVDD.n2636 0.00476
R49089 DVDD.n16290 DVDD.n2636 0.00476
R49090 DVDD.n16292 DVDD.n16290 0.00476
R49091 DVDD.n16294 DVDD.n16292 0.00476
R49092 DVDD.n16294 DVDD.n2633 0.00476
R49093 DVDD.n16299 DVDD.n2633 0.00476
R49094 DVDD.n16301 DVDD.n16299 0.00476
R49095 DVDD.n16303 DVDD.n16301 0.00476
R49096 DVDD.n16303 DVDD.n2630 0.00476
R49097 DVDD.n16310 DVDD.n2630 0.00476
R49098 DVDD.n16310 DVDD.n16309 0.00476
R49099 DVDD.n16309 DVDD.n2570 0.00476
R49100 DVDD.n16317 DVDD.n2570 0.00476
R49101 DVDD.n16318 DVDD.n16317 0.00476
R49102 DVDD.n16359 DVDD.n16358 0.00476
R49103 DVDD.n16358 DVDD.n16357 0.00476
R49104 DVDD.n16357 DVDD.n16356 0.00476
R49105 DVDD.n16356 DVDD.n16354 0.00476
R49106 DVDD.n16354 DVDD.n16352 0.00476
R49107 DVDD.n16352 DVDD.n16350 0.00476
R49108 DVDD.n16350 DVDD.n16348 0.00476
R49109 DVDD.n16348 DVDD.n16346 0.00476
R49110 DVDD.n16346 DVDD.n16344 0.00476
R49111 DVDD.n16344 DVDD.n16342 0.00476
R49112 DVDD.n16340 DVDD.n16338 0.00476
R49113 DVDD.n16338 DVDD.n16336 0.00476
R49114 DVDD.n15748 DVDD.n15747 0.00476
R49115 DVDD.n15747 DVDD.n15745 0.00476
R49116 DVDD.n15745 DVDD.n15743 0.00476
R49117 DVDD.n15743 DVDD.n15741 0.00476
R49118 DVDD.n15741 DVDD.n15739 0.00476
R49119 DVDD.n15739 DVDD.n15737 0.00476
R49120 DVDD.n15737 DVDD.n15735 0.00476
R49121 DVDD.n15735 DVDD.n15733 0.00476
R49122 DVDD.n15733 DVDD.n15731 0.00476
R49123 DVDD.n15731 DVDD.n15729 0.00476
R49124 DVDD.n15729 DVDD.n15727 0.00476
R49125 DVDD.n15727 DVDD.n3509 0.00476
R49126 DVDD.n15755 DVDD.n3509 0.00476
R49127 DVDD.n15760 DVDD.n3504 0.00476
R49128 DVDD.n15764 DVDD.n3504 0.00476
R49129 DVDD.n15766 DVDD.n15764 0.00476
R49130 DVDD.n15766 DVDD.n3502 0.00476
R49131 DVDD.n15771 DVDD.n3502 0.00476
R49132 DVDD.n15773 DVDD.n15771 0.00476
R49133 DVDD.n15775 DVDD.n15773 0.00476
R49134 DVDD.n15775 DVDD.n3499 0.00476
R49135 DVDD.n15780 DVDD.n3499 0.00476
R49136 DVDD.n15782 DVDD.n15780 0.00476
R49137 DVDD.n15784 DVDD.n15782 0.00476
R49138 DVDD.n15784 DVDD.n3496 0.00476
R49139 DVDD.n15788 DVDD.n3496 0.00476
R49140 DVDD.n15788 DVDD.n3418 0.00476
R49141 DVDD.n15797 DVDD.n3418 0.00476
R49142 DVDD.n15797 DVDD.n3416 0.00476
R49143 DVDD.n15801 DVDD.n3416 0.00476
R49144 DVDD.n15801 DVDD.n3414 0.00476
R49145 DVDD.n15805 DVDD.n3414 0.00476
R49146 DVDD.n15805 DVDD.n3412 0.00476
R49147 DVDD.n15810 DVDD.n3412 0.00476
R49148 DVDD.n15812 DVDD.n15810 0.00476
R49149 DVDD.n15815 DVDD.n15812 0.00476
R49150 DVDD.n15822 DVDD.n15820 0.00476
R49151 DVDD.n15822 DVDD.n3409 0.00476
R49152 DVDD.n15827 DVDD.n3409 0.00476
R49153 DVDD.n15829 DVDD.n15827 0.00476
R49154 DVDD.n15831 DVDD.n15829 0.00476
R49155 DVDD.n15831 DVDD.n3406 0.00476
R49156 DVDD.n15835 DVDD.n3406 0.00476
R49157 DVDD.n15835 DVDD.n3346 0.00476
R49158 DVDD.n15841 DVDD.n3346 0.00476
R49159 DVDD.n15841 DVDD.n3344 0.00476
R49160 DVDD.n15845 DVDD.n3344 0.00476
R49161 DVDD.n15845 DVDD.n3342 0.00476
R49162 DVDD.n15850 DVDD.n3342 0.00476
R49163 DVDD.n15850 DVDD.n3340 0.00476
R49164 DVDD.n15855 DVDD.n3340 0.00476
R49165 DVDD.n15857 DVDD.n15855 0.00476
R49166 DVDD.n15859 DVDD.n15857 0.00476
R49167 DVDD.n15859 DVDD.n3338 0.00476
R49168 DVDD.n15864 DVDD.n3338 0.00476
R49169 DVDD.n15866 DVDD.n15864 0.00476
R49170 DVDD.n15868 DVDD.n15866 0.00476
R49171 DVDD.n15868 DVDD.n3335 0.00476
R49172 DVDD.n15873 DVDD.n3335 0.00476
R49173 DVDD.n15877 DVDD.n2379 0.00476
R49174 DVDD.n16380 DVDD.n2379 0.00476
R49175 DVDD.n16380 DVDD.n16379 0.00476
R49176 DVDD.n16379 DVDD.n16378 0.00476
R49177 DVDD.n16378 DVDD.n16377 0.00476
R49178 DVDD.n16377 DVDD.n2384 0.00476
R49179 DVDD.n16373 DVDD.n2384 0.00476
R49180 DVDD.n16373 DVDD.n16372 0.00476
R49181 DVDD.n16372 DVDD.n2389 0.00476
R49182 DVDD.n2497 DVDD.n2389 0.00476
R49183 DVDD.n2499 DVDD.n2497 0.00476
R49184 DVDD.n2499 DVDD.n2493 0.00476
R49185 DVDD.n2504 DVDD.n2493 0.00476
R49186 DVDD.n2506 DVDD.n2504 0.00476
R49187 DVDD.n2508 DVDD.n2506 0.00476
R49188 DVDD.n2508 DVDD.n2490 0.00476
R49189 DVDD.n2513 DVDD.n2490 0.00476
R49190 DVDD.n2515 DVDD.n2513 0.00476
R49191 DVDD.n2517 DVDD.n2515 0.00476
R49192 DVDD.n2517 DVDD.n2487 0.00476
R49193 DVDD.n16366 DVDD.n2487 0.00476
R49194 DVDD.n16366 DVDD.n16365 0.00476
R49195 DVDD.n16365 DVDD.n16364 0.00476
R49196 DVDD.n2565 DVDD.n2564 0.00476
R49197 DVDD.n2564 DVDD.n2562 0.00476
R49198 DVDD.n2562 DVDD.n2560 0.00476
R49199 DVDD.n2560 DVDD.n2558 0.00476
R49200 DVDD.n2558 DVDD.n2556 0.00476
R49201 DVDD.n2556 DVDD.n2554 0.00476
R49202 DVDD.n2554 DVDD.n2552 0.00476
R49203 DVDD.n2552 DVDD.n2550 0.00476
R49204 DVDD.n2550 DVDD.n2548 0.00476
R49205 DVDD.n2548 DVDD.n2546 0.00476
R49206 DVDD.n2544 DVDD.n2542 0.00476
R49207 DVDD.n2542 DVDD.n2540 0.00476
R49208 DVDD.n15754 DVDD.n15753 0.00476
R49209 DVDD.n15762 DVDD.n15761 0.00476
R49210 DVDD.n15763 DVDD.n15762 0.00476
R49211 DVDD.n15802 DVDD.n3415 0.00476
R49212 DVDD.n15803 DVDD.n15802 0.00476
R49213 DVDD.n15804 DVDD.n15803 0.00476
R49214 DVDD.n15840 DVDD.n3343 0.00476
R49215 DVDD.n15846 DVDD.n3343 0.00476
R49216 DVDD.n15847 DVDD.n15846 0.00476
R49217 DVDD.n15849 DVDD.n15847 0.00476
R49218 DVDD.n15849 DVDD.n15848 0.00476
R49219 DVDD.n16376 DVDD.n2362 0.00476
R49220 DVDD.n16376 DVDD.n16375 0.00476
R49221 DVDD.n16375 DVDD.n16374 0.00476
R49222 DVDD.n16367 DVDD.n2486 0.00476
R49223 DVDD.n16363 DVDD.n2486 0.00476
R49224 DVDD.n2563 DVDD.n2524 0.00476
R49225 DVDD.n15688 DVDD.n15687 0.00476
R49226 DVDD.n15685 DVDD.n5112 0.00476
R49227 DVDD.n15681 DVDD.n5112 0.00476
R49228 DVDD.n15677 DVDD.n15620 0.00476
R49229 DVDD.n15673 DVDD.n15620 0.00476
R49230 DVDD.n15673 DVDD.n15672 0.00476
R49231 DVDD.n15906 DVDD.n3296 0.00476
R49232 DVDD.n15902 DVDD.n3296 0.00476
R49233 DVDD.n15902 DVDD.n15901 0.00476
R49234 DVDD.n15901 DVDD.n15900 0.00476
R49235 DVDD.n15900 DVDD.n3322 0.00476
R49236 DVDD.n16278 DVDD.n2640 0.00476
R49237 DVDD.n16279 DVDD.n16278 0.00476
R49238 DVDD.n16280 DVDD.n16279 0.00476
R49239 DVDD.n16316 DVDD.n16315 0.00476
R49240 DVDD.n16316 DVDD.n2526 0.00476
R49241 DVDD.n16360 DVDD.n569 0.00476
R49242 DVDD.n15463 DVDD.n15462 0.00476
R49243 DVDD.n15471 DVDD.n15470 0.00476
R49244 DVDD.n15472 DVDD.n15471 0.00476
R49245 DVDD.n15514 DVDD.n5159 0.00476
R49246 DVDD.n15514 DVDD.n15513 0.00476
R49247 DVDD.n15513 DVDD.n15512 0.00476
R49248 DVDD.n15986 DVDD.n3202 0.00476
R49249 DVDD.n15982 DVDD.n3202 0.00476
R49250 DVDD.n15982 DVDD.n15981 0.00476
R49251 DVDD.n15981 DVDD.n15980 0.00476
R49252 DVDD.n15980 DVDD.n15948 0.00476
R49253 DVDD.n16254 DVDD.n2770 0.00476
R49254 DVDD.n16250 DVDD.n2770 0.00476
R49255 DVDD.n16250 DVDD.n16249 0.00476
R49256 DVDD.n16245 DVDD.n2833 0.00476
R49257 DVDD.n16241 DVDD.n2833 0.00476
R49258 DVDD.n16238 DVDD.n656 0.00476
R49259 DVDD.n15396 DVDD.n5394 0.00476
R49260 DVDD.n15394 DVDD.n15349 0.00476
R49261 DVDD.n15390 DVDD.n15349 0.00476
R49262 DVDD.n16006 DVDD.n3137 0.00476
R49263 DVDD.n16002 DVDD.n3137 0.00476
R49264 DVDD.n16002 DVDD.n16001 0.00476
R49265 DVDD.n16093 DVDD.n16092 0.00476
R49266 DVDD.n16094 DVDD.n16093 0.00476
R49267 DVDD.n16094 DVDD.n3049 0.00476
R49268 DVDD.n16101 DVDD.n3049 0.00476
R49269 DVDD.n16102 DVDD.n16101 0.00476
R49270 DVDD.n16152 DVDD.n2991 0.00476
R49271 DVDD.n16153 DVDD.n16152 0.00476
R49272 DVDD.n16154 DVDD.n16153 0.00476
R49273 DVDD.n16193 DVDD.n2920 0.00476
R49274 DVDD.n16194 DVDD.n16193 0.00476
R49275 DVDD.n16197 DVDD.n16196 0.00476
R49276 DVDD.n20245 DVDD.n20244 0.00474286
R49277 DVDD.n20321 DVDD.n19849 0.00474286
R49278 DVDD.n20737 DVDD.n20736 0.00474286
R49279 DVDD.n20812 DVDD.n18877 0.00474286
R49280 DVDD.n22181 DVDD.n257 0.00474286
R49281 DVDD.n429 DVDD.n387 0.00474286
R49282 DVDD.n10093 DVDD.n9632 0.00474286
R49283 DVDD.n10004 DVDD.n9963 0.00474286
R49284 DVDD.n21159 DVDD.n18743 0.00474286
R49285 DVDD.n65 DVDD.n64 0.00474286
R49286 DVDD.n9687 DVDD.n9668 0.00471463
R49287 DVDD.n9954 DVDD.n9741 0.00471463
R49288 DVDD.n10094 DVDD.n9612 0.00471463
R49289 DVDD.n9950 DVDD.n9610 0.00471463
R49290 DVDD.n4571 DVDD.n4281 0.0047
R49291 DVDD.n20071 DVDD.n20059 0.00467857
R49292 DVDD DVDD.n18943 0.00467857
R49293 DVDD.n20602 DVDD.n19181 0.00467857
R49294 DVDD DVDD.n18971 0.00467857
R49295 DVDD.n3979 DVDD.n3910 0.00467857
R49296 DVDD DVDD.n22079 0.00467857
R49297 DVDD.n9862 DVDD.n5475 0.00467857
R49298 DVDD DVDD.n794 0.00467857
R49299 DVDD.n19699 DVDD.n19201 0.00467857
R49300 DVDD DVDD.n0 0.00467857
R49301 DVDD.n5011 DVDD.n4887 0.00466842
R49302 DVDD.n15702 DVDD.n15701 0.00466842
R49303 DVDD.n5297 DVDD.n5057 0.00466842
R49304 DVDD.n5329 DVDD.n5244 0.00466842
R49305 DVDD.n5351 DVDD.n5233 0.00466842
R49306 DVDD.n5417 DVDD.n5397 0.00466842
R49307 DVDD.n5456 DVDD.n5405 0.00466842
R49308 DVDD.n18014 DVDD.n523 0.00466842
R49309 DVDD.n17983 DVDD.n552 0.00466842
R49310 DVDD.n629 DVDD.n578 0.00466842
R49311 DVDD.n691 DVDD.n663 0.00466842
R49312 DVDD.n713 DVDD.n679 0.00466842
R49313 DVDD.n17947 DVDD.n749 0.00466842
R49314 DVDD.n17908 DVDD.n757 0.00466842
R49315 DVDD.n4157 DVDD.n3735 0.0046625
R49316 DVDD.n4537 DVDD.n4402 0.0046625
R49317 DVDD.n15556 DVDD.n2668 0.00462683
R49318 DVDD.n15555 DVDD.n2589 0.00462683
R49319 DVDD.n15559 DVDD.n3254 0.00462683
R49320 DVDD.n15562 DVDD.n15561 0.00462683
R49321 DVDD.n10585 DVDD.n10329 0.00462664
R49322 DVDD.n14278 DVDD.n10577 0.00462664
R49323 DVDD.n4699 DVDD.n4200 0.004625
R49324 DVDD.n20035 DVDD.n20027 0.00461429
R49325 DVDD.n19862 DVDD.n19845 0.00461429
R49326 DVDD.n19157 DVDD.n19145 0.00461429
R49327 DVDD.n20796 DVDD.n18874 0.00461429
R49328 DVDD.n4020 DVDD.n247 0.00461429
R49329 DVDD.n396 DVDD.n382 0.00461429
R49330 DVDD.n9911 DVDD.n9623 0.00461429
R49331 DVDD.n9972 DVDD.n9958 0.00461429
R49332 DVDD.n21110 DVDD.n18739 0.00461429
R49333 DVDD.n22269 DVDD.n60 0.00461429
R49334 DVDD.n18126 DVDD.n502 0.00460625
R49335 DVDD.n21674 DVDD.n18538 0.00456721
R49336 DVDD.n21361 DVDD.n21338 0.00456721
R49337 DVDD.n22000 DVDD.n21999 0.00456721
R49338 DVDD.n4851 DVDD.n3545 0.00456721
R49339 DVDD.n20147 DVDD.n20075 0.00455
R49340 DVDD.n20634 DVDD.n20606 0.00455
R49341 DVDD.n3958 DVDD.n3922 0.00455
R49342 DVDD.n4769 DVDD.n3646 0.00455
R49343 DVDD.n4555 DVDD.n4554 0.00455
R49344 DVDD.n9846 DVDD.n5471 0.00455
R49345 DVDD.n19657 DVDD.n19191 0.00455
R49346 DVDD.n2325 DVDD.n2294 0.00453902
R49347 DVDD.n16369 DVDD.n2413 0.00453902
R49348 DVDD.n15838 DVDD.n3370 0.00453902
R49349 DVDD.n15794 DVDD.n3473 0.00453902
R49350 DVDD.n18111 DVDD 0.00453415
R49351 DVDD.n15466 DVDD.n5226 0.0045
R49352 DVDD.n15916 DVDD.n3226 0.0045
R49353 DVDD.n15466 DVDD.n3507 0.0045
R49354 DVDD.n15916 DVDD.n3227 0.0045
R49355 DVDD.n16262 DVDD.n2703 0.0045
R49356 DVDD.n15817 DVDD.n3227 0.0045
R49357 DVDD.n15757 DVDD.n3507 0.0045
R49358 DVDD.n16320 DVDD.n2567 0.0045
R49359 DVDD.n16320 DVDD.n2568 0.0045
R49360 DVDD.n16262 DVDD.n16261 0.0045
R49361 DVDD.n16261 DVDD.n2705 0.0045
R49362 DVDD.n16189 DVDD.n2568 0.0045
R49363 DVDD.n20212 DVDD.n19977 0.00448571
R49364 DVDD.n20704 DVDD.n19140 0.00448571
R49365 DVDD.n4037 DVDD.n243 0.00448571
R49366 DVDD.n9928 DVDD.n9620 0.00448571
R49367 DVDD.n21187 DVDD.n21186 0.00448571
R49368 DVDD.n3663 DVDD.n3658 0.0044848
R49369 DVDD.n3752 DVDD.n3751 0.0044848
R49370 DVDD.n4441 DVDD.n4440 0.0044848
R49371 DVDD.n4844 DVDD.n3524 0.0044848
R49372 DVDD.n3667 DVDD.n3666 0.0044848
R49373 DVDD.n4260 DVDD.n4240 0.0044848
R49374 DVDD.n18060 DVDD.n18057 0.0044848
R49375 DVDD.n4405 DVDD.n4404 0.0044848
R49376 DVDD.n4401 DVDD.n4400 0.0044848
R49377 DVDD.n4261 DVDD.n4243 0.0044848
R49378 DVDD.n4404 DVDD.n4390 0.0044848
R49379 DVDD.n4400 DVDD.n4394 0.0044848
R49380 DVDD.n4261 DVDD.n4249 0.0044848
R49381 DVDD.n4260 DVDD.n4251 0.0044848
R49382 DVDD.n3751 DVDD.n3734 0.0044848
R49383 DVDD.n4440 DVDD.n3738 0.0044848
R49384 DVDD.n4844 DVDD.n3529 0.0044848
R49385 DVDD.n18061 DVDD.n18060 0.0044848
R49386 DVDD.n3666 DVDD.n3653 0.0044848
R49387 DVDD.n3658 DVDD.n3656 0.0044848
R49388 DVDD.n4997 DVDD.n4996 0.00447895
R49389 DVDD.n5003 DVDD.n5002 0.00447895
R49390 DVDD.n5005 DVDD.n4885 0.00447895
R49391 DVDD.n5303 DVDD.n5055 0.00447895
R49392 DVDD.n15699 DVDD.n5080 0.00447895
R49393 DVDD.n5335 DVDD.n5246 0.00447895
R49394 DVDD.n5345 DVDD.n5235 0.00447895
R49395 DVDD.n5411 DVDD.n5395 0.00447895
R49396 DVDD.n5563 DVDD.n5560 0.00447895
R49397 DVDD.n15147 DVDD.n5564 0.00447895
R49398 DVDD.n15144 DVDD.n5566 0.00447895
R49399 DVDD.n18034 DVDD.n18032 0.00447895
R49400 DVDD.n18027 DVDD.n18023 0.00447895
R49401 DVDD.n18020 DVDD.n521 0.00447895
R49402 DVDD.n635 DVDD.n570 0.00447895
R49403 DVDD.n17970 DVDD.n582 0.00447895
R49404 DVDD.n697 DVDD.n677 0.00447895
R49405 DVDD.n707 DVDD.n665 0.00447895
R49406 DVDD.n772 DVDD.n747 0.00447895
R49407 DVDD.n17738 DVDD.n17737 0.00447895
R49408 DVDD.n884 DVDD.n880 0.00447895
R49409 DVDD.n17734 DVDD.n886 0.00447895
R49410 DVDD.n22230 DVDD 0.0044381
R49411 DVDD.n22231 DVDD 0.0044381
R49412 DVDD.n21921 DVDD 0.0044381
R49413 DVDD.n21922 DVDD 0.0044381
R49414 DVDD.n4770 DVDD.n4769 0.0044375
R49415 DVDD.n4555 DVDD.n4407 0.0044375
R49416 DVDD.n20147 DVDD.n20126 0.00442143
R49417 DVDD.n20634 DVDD.n20613 0.00442143
R49418 DVDD.n3958 DVDD.n3931 0.00442143
R49419 DVDD.n9846 DVDD.n5482 0.00442143
R49420 DVDD.n19657 DVDD.n19197 0.00442143
R49421 DVDD.n18090 DVDD.n18068 0.0044
R49422 DVDD.n5510 DVDD.n5495 0.00438421
R49423 DVDD.n830 DVDD.n801 0.00438421
R49424 DVDD.n18127 DVDD.n18126 0.00438125
R49425 DVDD.n14014 DVDD.n10709 0.00436577
R49426 DVDD.n16739 DVDD.n16738 0.00436577
R49427 DVDD.n14015 DVDD.n10707 0.00436577
R49428 DVDD.n16744 DVDD.n16743 0.00436577
R49429 DVDD.n9799 DVDD.n9665 0.00436341
R49430 DVDD.n9798 DVDD.n9736 0.00436341
R49431 DVDD.n9802 DVDD.n9630 0.00436341
R49432 DVDD.n9805 DVDD.n9804 0.00436341
R49433 DVDD.n20035 DVDD.n19973 0.00435714
R49434 DVDD.n19862 DVDD.n19838 0.00435714
R49435 DVDD.n19157 DVDD.n19136 0.00435714
R49436 DVDD.n20796 DVDD.n18884 0.00435714
R49437 DVDD.n4020 DVDD.n239 0.00435714
R49438 DVDD.n396 DVDD.n376 0.00435714
R49439 DVDD.n9911 DVDD.n9616 0.00435714
R49440 DVDD.n9972 DVDD.n9753 0.00435714
R49441 DVDD.n21110 DVDD.n21096 0.00435714
R49442 DVDD.n22269 DVDD.n75 0.00435714
R49443 DVDD.n4736 DVDD.n3757 0.004325
R49444 DVDD.n4539 DVDD.n4402 0.004325
R49445 DVDD.n14830 DVDD.n14829 0.004325
R49446 DVDD.n20165 DVDD.n20059 0.00429286
R49447 DVDD.n20657 DVDD.n19181 0.00429286
R49448 DVDD.n3979 DVDD.n3978 0.00429286
R49449 DVDD.n9862 DVDD.n5477 0.00429286
R49450 DVDD.n19701 DVDD.n19201 0.00429286
R49451 DVDD.n5021 DVDD.n3515 0.00428947
R49452 DVDD.n5268 DVDD.n5067 0.00428947
R49453 DVDD.n5287 DVDD.n5072 0.00428947
R49454 DVDD.n5319 DVDD.n5240 0.00428947
R49455 DVDD.n5361 DVDD.n5251 0.00428947
R49456 DVDD.n5427 DVDD.n5390 0.00428947
R49457 DVDD.n5446 DVDD.n5385 0.00428947
R49458 DVDD.n18004 DVDD.n536 0.00428947
R49459 DVDD.n600 DVDD.n589 0.00428947
R49460 DVDD.n619 DVDD.n592 0.00428947
R49461 DVDD.n662 DVDD.n648 0.00428947
R49462 DVDD.n723 DVDD.n671 0.00428947
R49463 DVDD.n17937 DVDD.n769 0.00428947
R49464 DVDD.n17918 DVDD.n764 0.00428947
R49465 DVDD.n15074 DVDD.n15073 0.00428947
R49466 DVDD.n9570 DVDD.n9219 0.00428947
R49467 DVDD.n15547 DVDD.n2664 0.00427561
R49468 DVDD.n15522 DVDD.n2733 0.00427561
R49469 DVDD.n5195 DVDD.n2729 0.00427561
R49470 DVDD.n3032 DVDD.n3006 0.00427561
R49471 DVDD.n15546 DVDD.n2587 0.00427561
R49472 DVDD.n15521 DVDD.n2803 0.00427561
R49473 DVDD.n5194 DVDD.n2799 0.00427561
R49474 DVDD.n2963 DVDD.n2935 0.00427561
R49475 DVDD.n15550 DVDD.n3252 0.00427561
R49476 DVDD.n15524 DVDD.n3173 0.00427561
R49477 DVDD.n5197 DVDD.n3169 0.00427561
R49478 DVDD.n3081 DVDD.n3066 0.00427561
R49479 DVDD.n15553 DVDD.n15552 0.00427561
R49480 DVDD.n15527 DVDD.n15526 0.00427561
R49481 DVDD.n5200 DVDD.n5199 0.00427561
R49482 DVDD.n16065 DVDD.n3134 0.00427561
R49483 DVDD.n18070 DVDD.n18054 0.00426875
R49484 DVDD.n21776 DVDD.n18388 0.004246
R49485 DVDD.n21726 DVDD.n21725 0.004246
R49486 DVDD.n22042 DVDD.n18210 0.004246
R49487 DVDD.n18094 DVDD.n18093 0.004246
R49488 DVDD.n13746 DVDD.n12285 0.00423362
R49489 DVDD.n16706 DVDD.n2164 0.00423362
R49490 DVDD.n13747 DVDD.n12283 0.00423362
R49491 DVDD.n16707 DVDD.n2162 0.00423362
R49492 DVDD.n20285 DVDD.n19869 0.00422857
R49493 DVDD.n20321 DVDD.n19834 0.00422857
R49494 DVDD.n20780 DVDD.n20779 0.00422857
R49495 DVDD.n20812 DVDD.n18882 0.00422857
R49496 DVDD.n22158 DVDD.n310 0.00422857
R49497 DVDD.n429 DVDD.n372 0.00422857
R49498 DVDD.n10066 DVDD.n10065 0.00422857
R49499 DVDD.n10004 DVDD.n9750 0.00422857
R49500 DVDD.n22260 DVDD.n85 0.00422857
R49501 DVDD.n64 DVDD.n42 0.00422857
R49502 DVDD.n18483 DVDD.n18476 0.00422
R49503 DVDD.n21736 DVDD.n21735 0.00422
R49504 DVDD.n18394 DVDD.n18393 0.00422
R49505 DVDD.n21876 DVDD.n21788 0.00422
R49506 DVDD.n21899 DVDD.n21898 0.00422
R49507 DVDD.n22058 DVDD.n18205 0.00422
R49508 DVDD.n21216 DVDD.n18666 0.00422
R49509 DVDD.n21649 DVDD.n21648 0.00422
R49510 DVDD.n21688 DVDD.n21687 0.00422
R49511 DVDD.n21961 DVDD.n18284 0.00422
R49512 DVDD.n21976 DVDD.n18270 0.00422
R49513 DVDD.n22184 DVDD.n233 0.00422
R49514 DVDD.n21233 DVDD.n21220 0.00422
R49515 DVDD.n21332 DVDD.n21331 0.00422
R49516 DVDD.n21685 DVDD.n18532 0.00422
R49517 DVDD.n18323 DVDD.n18286 0.00422
R49518 DVDD.n18339 DVDD.n18272 0.00422
R49519 DVDD.n22186 DVDD.n228 0.00422
R49520 DVDD.n18485 DVDD.n18462 0.00422
R49521 DVDD.n21738 DVDD.n18408 0.00422
R49522 DVDD.n21753 DVDD.n18404 0.00422
R49523 DVDD.n21874 DVDD.n21843 0.00422
R49524 DVDD.n21815 DVDD.n21804 0.00422
R49525 DVDD.n22057 DVDD.n22056 0.00422
R49526 DVDD.n4834 DVDD.n3564 0.00422
R49527 DVDD.n4135 DVDD.n3827 0.00422
R49528 DVDD.n18194 DVDD.n460 0.00422
R49529 DVDD.n4450 DVDD.n4419 0.0042125
R49530 DVDD.n4597 DVDD.n4596 0.0042125
R49531 DVDD.n15287 DVDD.n15286 0.00419474
R49532 DVDD.n811 DVDD.n792 0.00419474
R49533 DVDD.n20344 DVDD.n18942 0.00416429
R49534 DVDD.n20843 DVDD.n18970 0.00416429
R49535 DVDD.n22102 DVDD.n22078 0.00416429
R49536 DVDD.n10027 DVDD.n793 0.00416429
R49537 DVDD.n22319 DVDD.n23 0.00416429
R49538 DVDD.n4095 DVDD.n4090 0.00416
R49539 DVDD.n4500 DVDD.n4192 0.00416
R49540 DVDD.n3498 DVDD.n3493 0.00416
R49541 DVDD.n3337 DVDD.n2344 0.00416
R49542 DVDD.n15640 DVDD.n15614 0.00416
R49543 DVDD.n15890 DVDD.n2696 0.00416
R49544 DVDD.n15485 DVDD.n5140 0.00416
R49545 DVDD.n15970 DVDD.n2755 0.00416
R49546 DVDD.n15378 DVDD.n3119 0.00416
R49547 DVDD.n3044 DVDD.n3036 0.00416
R49548 DVDD.n3604 DVDD.n3526 0.00415625
R49549 DVDD.n18425 DVDD.n166 0.00413
R49550 DVDD.n21763 DVDD.n173 0.00413
R49551 DVDD.n22061 DVDD.n18214 0.00413
R49552 DVDD.n21652 DVDD.n18554 0.00413
R49553 DVDD.n21692 DVDD.n18515 0.00413
R49554 DVDD.n22027 DVDD.n22024 0.00413
R49555 DVDD.n21654 DVDD.n18550 0.00413
R49556 DVDD.n21662 DVDD.n18527 0.00413
R49557 DVDD.n22009 DVDD.n21988 0.00413
R49558 DVDD.n21592 DVDD.n21591 0.00413
R49559 DVDD.n21752 DVDD.n18398 0.00413
R49560 DVDD.n18219 DVDD.n18217 0.00413
R49561 DVDD.n18146 DVDD.n457 0.00413
R49562 DVDD.n2553 DVDD.n513 0.00413
R49563 DVDD.n16349 DVDD.n566 0.00413
R49564 DVDD.n16228 DVDD.n653 0.00413
R49565 DVDD.n2909 DVDD.n742 0.00413
R49566 DVDD.n20195 DVDD.n19737 0.0041
R49567 DVDD.n20271 DVDD.n19940 0.0041
R49568 DVDD.n20687 DVDD.n18844 0.0041
R49569 DVDD.n19061 DVDD.n19050 0.0041
R49570 DVDD.n4052 DVDD.n3873 0.0041
R49571 DVDD.n344 DVDD.n301 0.0041
R49572 DVDD.n4432 DVDD.n3736 0.0041
R49573 DVDD.n4138 DVDD.n4137 0.0041
R49574 DVDD.n4504 DVDD.n4204 0.0041
R49575 DVDD.n15796 DVDD.n15795 0.0041
R49576 DVDD.n2378 DVDD.n2348 0.0041
R49577 DVDD.n15678 DVDD.n15619 0.0041
R49578 DVDD.n16268 DVDD.n16266 0.0041
R49579 DVDD.n15528 DVDD.n5144 0.0041
R49580 DVDD.n2766 DVDD.n2765 0.0041
R49581 DVDD.n16067 DVDD.n3123 0.0041
R49582 DVDD.n16142 DVDD.n16140 0.0041
R49583 DVDD.n9893 DVDD.n9769 0.0041
R49584 DVDD.n9716 DVDD.n9691 0.0041
R49585 DVDD.n5000 DVDD.n4884 0.0041
R49586 DVDD.n5025 DVDD.n4890 0.0041
R49587 DVDD.n5036 DVDD.n4892 0.0041
R49588 DVDD.n5272 DVDD.n5062 0.0041
R49589 DVDD.n5283 DVDD.n5060 0.0041
R49590 DVDD.n5365 DVDD.n5230 0.0041
R49591 DVDD.n5431 DVDD.n5400 0.0041
R49592 DVDD.n5442 DVDD.n5402 0.0041
R49593 DVDD.n543 DVDD.n520 0.0041
R49594 DVDD.n18000 DVDD.n526 0.0041
R49595 DVDD.n17989 DVDD.n528 0.0041
R49596 DVDD.n604 DVDD.n573 0.0041
R49597 DVDD.n615 DVDD.n587 0.0041
R49598 DVDD.n727 DVDD.n657 0.0041
R49599 DVDD.n17933 DVDD.n752 0.0041
R49600 DVDD.n17922 DVDD.n754 0.0041
R49601 DVDD.n21202 DVDD.n18677 0.0041
R49602 DVDD.n21136 DVDD.n101 0.0041
R49603 DVDD DVDD.n21783 0.00408591
R49604 DVDD.n22240 DVDD.n127 0.00407
R49605 DVDD.n21836 DVDD.n21789 0.00407
R49606 DVDD.n21829 DVDD.n21790 0.00407
R49607 DVDD.n21248 DVDD.n18670 0.00407
R49608 DVDD.n21963 DVDD.n199 0.00407
R49609 DVDD.n21966 DVDD.n203 0.00407
R49610 DVDD.n21224 DVDD.n18655 0.00407
R49611 DVDD.n18363 DVDD.n18316 0.00407
R49612 DVDD.n18329 DVDD.n18281 0.00407
R49613 DVDD.n22242 DVDD.n123 0.00407
R49614 DVDD.n21873 DVDD.n21859 0.00407
R49615 DVDD.n21902 DVDD.n21810 0.00407
R49616 DVDD.n18197 DVDD.n461 0.00407
R49617 DVDD.n18043 DVDD.n517 0.00407
R49618 DVDD.n16335 DVDD.n565 0.00407
R49619 DVDD.n16214 DVDD.n652 0.00407
R49620 DVDD.n17954 DVDD.n746 0.00407
R49621 DVDD.n3613 DVDD.n3523 0.00404375
R49622 DVDD.n3808 DVDD.n3767 0.00404
R49623 DVDD.n4640 DVDD.n4628 0.00404
R49624 DVDD.n18135 DVDD.n18134 0.00404
R49625 DVDD.n490 DVDD.n486 0.00404
R49626 DVDD.n16199 DVDD.n16198 0.00404
R49627 DVDD.n16240 DVDD.n16239 0.00404
R49628 DVDD.n16359 DVDD.n2527 0.00404
R49629 DVDD.n2565 DVDD.n2523 0.00404
R49630 DVDD.n15830 DVDD.n3390 0.00404
R49631 DVDD.n2507 DVDD.n2434 0.00404
R49632 DVDD.n16362 DVDD.n2524 0.00404
R49633 DVDD.n3310 DVDD.n3280 0.00404
R49634 DVDD.n16298 DVDD.n2615 0.00404
R49635 DVDD.n16361 DVDD.n16360 0.00404
R49636 DVDD.n15928 DVDD.n3188 0.00404
R49637 DVDD.n2859 DVDD.n2819 0.00404
R49638 DVDD.n16238 DVDD.n2525 0.00404
R49639 DVDD.n3087 DVDD.n3075 0.00404
R49640 DVDD.n16172 DVDD.n2958 0.00404
R49641 DVDD.n16197 DVDD.n16195 0.00404
R49642 DVDD.n20327 DVDD.n18938 0.00403571
R49643 DVDD.n20827 DVDD.n18966 0.00403571
R49644 DVDD.n439 DVDD.n435 0.00403571
R49645 DVDD.n17877 DVDD.n805 0.00403571
R49646 DVDD.n22342 DVDD.n22335 0.00403571
R49647 DVDD.n4781 DVDD.n4780 0.004025
R49648 DVDD.n9941 DVDD.n9674 0.0040122
R49649 DVDD.n9940 DVDD.n9744 0.0040122
R49650 DVDD.n9944 DVDD.n9637 0.0040122
R49651 DVDD.n9946 DVDD.n9812 0.0040122
R49652 DVDD.n3589 DVDD.n3561 0.00401
R49653 DVDD.n15734 DVDD.n15710 0.00401
R49654 DVDD.n5082 DVDD.n5050 0.00401
R49655 DVDD.n15443 DVDD.n15419 0.00401
R49656 DVDD.n15318 DVDD.n5380 0.00401
R49657 DVDD.n5506 DVDD.n5489 0.00400526
R49658 DVDD.n826 DVDD.n809 0.00400526
R49659 DVDD.n4744 DVDD.n4743 0.0039875
R49660 DVDD.n3820 DVDD.n3812 0.00398
R49661 DVDD.n4633 DVDD.n4213 0.00398
R49662 DVDD.n15811 DVDD.n3394 0.00398
R49663 DVDD.n16371 DVDD.n2385 0.00398
R49664 DVDD.n15665 DVDD.n3284 0.00398
R49665 DVDD.n16282 DVDD.n2619 0.00398
R49666 DVDD.n3229 DVDD.n3192 0.00398
R49667 DVDD.n16248 DVDD.n2792 0.00398
R49668 DVDD.n15994 DVDD.n3079 0.00398
R49669 DVDD.n16156 DVDD.n2962 0.00398
R49670 DVDD.n20051 DVDD.n19733 0.00397143
R49671 DVDD.n19173 DVDD.n18839 0.00397143
R49672 DVDD.n3995 DVDD.n3870 0.00397143
R49673 DVDD.n9877 DVDD.n9764 0.00397143
R49674 DVDD.n19680 DVDD.n18684 0.00397143
R49675 DVDD.n4838 DVDD.n4803 0.00395
R49676 DVDD.n3579 DVDD.n3552 0.00395
R49677 DVDD.n15750 DVDD.n15749 0.00395
R49678 DVDD.n15746 DVDD.n4899 0.00395
R49679 DVDD.n15700 DVDD.n5065 0.00395
R49680 DVDD.n5089 DVDD.n5041 0.00395
R49681 DVDD.n15459 DVDD.n15458 0.00395
R49682 DVDD.n15455 DVDD.n5255 0.00395
R49683 DVDD.n15325 DVDD.n5379 0.00395
R49684 DVDD.n15327 DVDD.n5374 0.00395
R49685 DVDD.n20603 DVDD.n19182 0.00393493
R49686 DVDD.n20601 DVDD.n19707 0.00393493
R49687 DVDD.n20643 DVDD.n19183 0.00393493
R49688 DVDD.n20600 DVDD.n19706 0.00393493
R49689 DVDD.n20644 DVDD.n19184 0.00393493
R49690 DVDD.n20599 DVDD.n19705 0.00393493
R49691 DVDD.n20645 DVDD.n19185 0.00393493
R49692 DVDD.n20598 DVDD.n19704 0.00393493
R49693 DVDD.n20646 DVDD.n19186 0.00393493
R49694 DVDD.n20597 DVDD.n19703 0.00393493
R49695 DVDD.n19214 DVDD.n19187 0.00393493
R49696 DVDD.n19213 DVDD.n19205 0.00393493
R49697 DVDD.n19698 DVDD.n19212 0.00393493
R49698 DVDD.n19211 DVDD.n19206 0.00393493
R49699 DVDD.n19697 DVDD.n19210 0.00393493
R49700 DVDD.n3939 DVDD.n3915 0.00393493
R49701 DVDD.n3967 DVDD.n3917 0.00393493
R49702 DVDD.n3938 DVDD.n3914 0.00393493
R49703 DVDD.n3968 DVDD.n3918 0.00393493
R49704 DVDD.n3937 DVDD.n3913 0.00393493
R49705 DVDD.n3969 DVDD.n3919 0.00393493
R49706 DVDD.n3936 DVDD.n3912 0.00393493
R49707 DVDD.n3970 DVDD.n3920 0.00393493
R49708 DVDD.n3935 DVDD.n3911 0.00393493
R49709 DVDD.n3977 DVDD.n3921 0.00393493
R49710 DVDD.n4824 DVDD.n4805 0.00393493
R49711 DVDD.n4804 DVDD.n3576 0.00393493
R49712 DVDD.n4825 DVDD.n4807 0.00393493
R49713 DVDD.n4806 DVDD.n3575 0.00393493
R49714 DVDD.n4826 DVDD.n4809 0.00393493
R49715 DVDD.n4808 DVDD.n3574 0.00393493
R49716 DVDD.n4827 DVDD.n4811 0.00393493
R49717 DVDD.n4810 DVDD.n3573 0.00393493
R49718 DVDD.n4828 DVDD.n4813 0.00393493
R49719 DVDD.n4812 DVDD.n3572 0.00393493
R49720 DVDD.n4829 DVDD.n4815 0.00393493
R49721 DVDD.n4814 DVDD.n3571 0.00393493
R49722 DVDD.n4830 DVDD.n4817 0.00393493
R49723 DVDD.n4816 DVDD.n3570 0.00393493
R49724 DVDD.n4831 DVDD.n4819 0.00393493
R49725 DVDD.n4818 DVDD.n3569 0.00393493
R49726 DVDD.n4832 DVDD.n4821 0.00393493
R49727 DVDD.n4820 DVDD.n3568 0.00393493
R49728 DVDD.n4833 DVDD.n4823 0.00393493
R49729 DVDD.n4822 DVDD.n3567 0.00393493
R49730 DVDD.n4837 DVDD.n4835 0.00393493
R49731 DVDD.n4836 DVDD.n3566 0.00393493
R49732 DVDD.n4839 DVDD.n3551 0.00393493
R49733 DVDD.n4843 DVDD.n4842 0.00393493
R49734 DVDD.n4841 DVDD.n4840 0.00393493
R49735 DVDD.n4852 DVDD.n3546 0.00393493
R49736 DVDD.n4856 DVDD.n4853 0.00393493
R49737 DVDD.n4855 DVDD.n4854 0.00393493
R49738 DVDD.n4867 DVDD.n3539 0.00393493
R49739 DVDD.n4869 DVDD.n4868 0.00393493
R49740 DVDD.n4873 DVDD.n4870 0.00393493
R49741 DVDD.n4872 DVDD.n4871 0.00393493
R49742 DVDD.n4880 DVDD.n3522 0.00393493
R49743 DVDD.n4894 DVDD.n4882 0.00393493
R49744 DVDD.n4898 DVDD.n3521 0.00393493
R49745 DVDD.n4895 DVDD.n4883 0.00393493
R49746 DVDD.n4897 DVDD.n3520 0.00393493
R49747 DVDD.n3939 DVDD.n3916 0.00393493
R49748 DVDD.n3967 DVDD.n3915 0.00393493
R49749 DVDD.n3938 DVDD.n3917 0.00393493
R49750 DVDD.n3968 DVDD.n3914 0.00393493
R49751 DVDD.n3937 DVDD.n3918 0.00393493
R49752 DVDD.n3969 DVDD.n3913 0.00393493
R49753 DVDD.n3936 DVDD.n3919 0.00393493
R49754 DVDD.n3970 DVDD.n3912 0.00393493
R49755 DVDD.n3935 DVDD.n3920 0.00393493
R49756 DVDD.n3921 DVDD.n3911 0.00393493
R49757 DVDD.n4824 DVDD.n3578 0.00393493
R49758 DVDD.n4805 DVDD.n4804 0.00393493
R49759 DVDD.n4825 DVDD.n3576 0.00393493
R49760 DVDD.n4807 DVDD.n4806 0.00393493
R49761 DVDD.n4826 DVDD.n3575 0.00393493
R49762 DVDD.n4809 DVDD.n4808 0.00393493
R49763 DVDD.n4827 DVDD.n3574 0.00393493
R49764 DVDD.n4811 DVDD.n4810 0.00393493
R49765 DVDD.n4828 DVDD.n3573 0.00393493
R49766 DVDD.n4813 DVDD.n4812 0.00393493
R49767 DVDD.n4829 DVDD.n3572 0.00393493
R49768 DVDD.n4815 DVDD.n4814 0.00393493
R49769 DVDD.n4830 DVDD.n3571 0.00393493
R49770 DVDD.n4817 DVDD.n4816 0.00393493
R49771 DVDD.n4831 DVDD.n3570 0.00393493
R49772 DVDD.n4819 DVDD.n4818 0.00393493
R49773 DVDD.n4832 DVDD.n3569 0.00393493
R49774 DVDD.n4821 DVDD.n4820 0.00393493
R49775 DVDD.n4833 DVDD.n3568 0.00393493
R49776 DVDD.n4823 DVDD.n4822 0.00393493
R49777 DVDD.n4835 DVDD.n3567 0.00393493
R49778 DVDD.n4837 DVDD.n4836 0.00393493
R49779 DVDD.n3566 DVDD.n3551 0.00393493
R49780 DVDD.n4845 DVDD.n4843 0.00393493
R49781 DVDD.n4842 DVDD.n4841 0.00393493
R49782 DVDD.n4840 DVDD.n3546 0.00393493
R49783 DVDD.n4853 DVDD.n4852 0.00393493
R49784 DVDD.n4856 DVDD.n4855 0.00393493
R49785 DVDD.n4854 DVDD.n3539 0.00393493
R49786 DVDD.n4868 DVDD.n4867 0.00393493
R49787 DVDD.n4870 DVDD.n4869 0.00393493
R49788 DVDD.n4873 DVDD.n4872 0.00393493
R49789 DVDD.n4871 DVDD.n3522 0.00393493
R49790 DVDD.n4894 DVDD.n4881 0.00393493
R49791 DVDD.n4898 DVDD.n4882 0.00393493
R49792 DVDD.n4895 DVDD.n3521 0.00393493
R49793 DVDD.n4897 DVDD.n4883 0.00393493
R49794 DVDD.n20597 DVDD.n19186 0.00393493
R49795 DVDD.n20646 DVDD.n19704 0.00393493
R49796 DVDD.n20598 DVDD.n19185 0.00393493
R49797 DVDD.n20645 DVDD.n19705 0.00393493
R49798 DVDD.n20599 DVDD.n19184 0.00393493
R49799 DVDD.n20644 DVDD.n19706 0.00393493
R49800 DVDD.n20600 DVDD.n19183 0.00393493
R49801 DVDD.n20643 DVDD.n19707 0.00393493
R49802 DVDD.n20601 DVDD.n19182 0.00393493
R49803 DVDD.n20656 DVDD.n20603 0.00393493
R49804 DVDD.n18974 DVDD.n18960 0.00393493
R49805 DVDD.n20853 DVDD.n18990 0.00393493
R49806 DVDD.n18991 DVDD.n18975 0.00393493
R49807 DVDD.n18988 DVDD.n18984 0.00393493
R49808 DVDD.n18992 DVDD.n18976 0.00393493
R49809 DVDD.n18987 DVDD.n18983 0.00393493
R49810 DVDD.n18993 DVDD.n18977 0.00393493
R49811 DVDD.n18986 DVDD.n18982 0.00393493
R49812 DVDD.n18994 DVDD.n18978 0.00393493
R49813 DVDD.n18985 DVDD.n18981 0.00393493
R49814 DVDD.n22341 DVDD.n6 0.00393493
R49815 DVDD.n22340 DVDD.n31 0.00393493
R49816 DVDD.n22339 DVDD.n7 0.00393493
R49817 DVDD.n22338 DVDD.n32 0.00393493
R49818 DVDD.n22337 DVDD.n8 0.00393493
R49819 DVDD.n22070 DVDD.n441 0.00393493
R49820 DVDD.n22085 DVDD.n18203 0.00393493
R49821 DVDD.n22110 DVDD.n442 0.00393493
R49822 DVDD.n22084 DVDD.n18202 0.00393493
R49823 DVDD.n22111 DVDD.n443 0.00393493
R49824 DVDD.n22083 DVDD.n18201 0.00393493
R49825 DVDD.n22112 DVDD.n444 0.00393493
R49826 DVDD.n22082 DVDD.n18200 0.00393493
R49827 DVDD.n22113 DVDD.n445 0.00393493
R49828 DVDD.n22081 DVDD.n18199 0.00393493
R49829 DVDD.n462 DVDD.n447 0.00393493
R49830 DVDD.n18196 DVDD.n18183 0.00393493
R49831 DVDD.n18195 DVDD.n463 0.00393493
R49832 DVDD.n18182 DVDD.n18181 0.00393493
R49833 DVDD.n18184 DVDD.n464 0.00393493
R49834 DVDD.n18180 DVDD.n18179 0.00393493
R49835 DVDD.n18185 DVDD.n465 0.00393493
R49836 DVDD.n18178 DVDD.n18177 0.00393493
R49837 DVDD.n18186 DVDD.n466 0.00393493
R49838 DVDD.n18176 DVDD.n18175 0.00393493
R49839 DVDD.n18187 DVDD.n467 0.00393493
R49840 DVDD.n18174 DVDD.n18173 0.00393493
R49841 DVDD.n18188 DVDD.n468 0.00393493
R49842 DVDD.n18172 DVDD.n18171 0.00393493
R49843 DVDD.n18189 DVDD.n469 0.00393493
R49844 DVDD.n18170 DVDD.n18169 0.00393493
R49845 DVDD.n18190 DVDD.n470 0.00393493
R49846 DVDD.n18168 DVDD.n18167 0.00393493
R49847 DVDD.n18191 DVDD.n471 0.00393493
R49848 DVDD.n18166 DVDD.n18165 0.00393493
R49849 DVDD.n18192 DVDD.n472 0.00393493
R49850 DVDD.n18164 DVDD.n18163 0.00393493
R49851 DVDD.n18193 DVDD.n474 0.00393493
R49852 DVDD.n18055 DVDD.n497 0.00393493
R49853 DVDD.n18053 DVDD.n18049 0.00393493
R49854 DVDD.n18080 DVDD.n498 0.00393493
R49855 DVDD.n18052 DVDD.n18048 0.00393493
R49856 DVDD.n18081 DVDD.n499 0.00393493
R49857 DVDD.n18056 DVDD.n18047 0.00393493
R49858 DVDD.n18082 DVDD.n500 0.00393493
R49859 DVDD.n18051 DVDD.n18046 0.00393493
R49860 DVDD.n18083 DVDD.n501 0.00393493
R49861 DVDD.n18050 DVDD.n18045 0.00393493
R49862 DVDD.n518 DVDD.n503 0.00393493
R49863 DVDD.n18042 DVDD.n18038 0.00393493
R49864 DVDD.n18041 DVDD.n519 0.00393493
R49865 DVDD.n18037 DVDD.n541 0.00393493
R49866 DVDD.n541 DVDD.n519 0.00393493
R49867 DVDD.n18042 DVDD.n18041 0.00393493
R49868 DVDD.n18038 DVDD.n518 0.00393493
R49869 DVDD.n18044 DVDD.n503 0.00393493
R49870 DVDD.n18050 DVDD.n501 0.00393493
R49871 DVDD.n18083 DVDD.n18046 0.00393493
R49872 DVDD.n18051 DVDD.n500 0.00393493
R49873 DVDD.n18082 DVDD.n18047 0.00393493
R49874 DVDD.n18056 DVDD.n499 0.00393493
R49875 DVDD.n18081 DVDD.n18048 0.00393493
R49876 DVDD.n18052 DVDD.n498 0.00393493
R49877 DVDD.n18080 DVDD.n18049 0.00393493
R49878 DVDD.n18053 DVDD.n497 0.00393493
R49879 DVDD.n18125 DVDD.n18055 0.00393493
R49880 DVDD.n18193 DVDD.n18164 0.00393493
R49881 DVDD.n18163 DVDD.n472 0.00393493
R49882 DVDD.n18192 DVDD.n18166 0.00393493
R49883 DVDD.n18165 DVDD.n471 0.00393493
R49884 DVDD.n18191 DVDD.n18168 0.00393493
R49885 DVDD.n18167 DVDD.n470 0.00393493
R49886 DVDD.n18190 DVDD.n18170 0.00393493
R49887 DVDD.n18169 DVDD.n469 0.00393493
R49888 DVDD.n18189 DVDD.n18172 0.00393493
R49889 DVDD.n18171 DVDD.n468 0.00393493
R49890 DVDD.n18188 DVDD.n18174 0.00393493
R49891 DVDD.n18173 DVDD.n467 0.00393493
R49892 DVDD.n18187 DVDD.n18176 0.00393493
R49893 DVDD.n18175 DVDD.n466 0.00393493
R49894 DVDD.n18186 DVDD.n18178 0.00393493
R49895 DVDD.n18177 DVDD.n465 0.00393493
R49896 DVDD.n18185 DVDD.n18180 0.00393493
R49897 DVDD.n18179 DVDD.n464 0.00393493
R49898 DVDD.n18184 DVDD.n18182 0.00393493
R49899 DVDD.n18181 DVDD.n463 0.00393493
R49900 DVDD.n18196 DVDD.n18195 0.00393493
R49901 DVDD.n18183 DVDD.n462 0.00393493
R49902 DVDD.n18198 DVDD.n447 0.00393493
R49903 DVDD.n22081 DVDD.n445 0.00393493
R49904 DVDD.n22113 DVDD.n18200 0.00393493
R49905 DVDD.n22082 DVDD.n444 0.00393493
R49906 DVDD.n22112 DVDD.n18201 0.00393493
R49907 DVDD.n22083 DVDD.n443 0.00393493
R49908 DVDD.n22111 DVDD.n18202 0.00393493
R49909 DVDD.n22084 DVDD.n442 0.00393493
R49910 DVDD.n22110 DVDD.n18203 0.00393493
R49911 DVDD.n22085 DVDD.n441 0.00393493
R49912 DVDD.n22121 DVDD.n22070 0.00393493
R49913 DVDD.n18985 DVDD.n18978 0.00393493
R49914 DVDD.n18994 DVDD.n18982 0.00393493
R49915 DVDD.n18986 DVDD.n18977 0.00393493
R49916 DVDD.n18993 DVDD.n18983 0.00393493
R49917 DVDD.n18987 DVDD.n18976 0.00393493
R49918 DVDD.n18992 DVDD.n18984 0.00393493
R49919 DVDD.n18988 DVDD.n18975 0.00393493
R49920 DVDD.n20853 DVDD.n18991 0.00393493
R49921 DVDD.n18990 DVDD.n18974 0.00393493
R49922 DVDD.n20855 DVDD.n18960 0.00393493
R49923 DVDD.n32 DVDD.n8 0.00393493
R49924 DVDD.n22339 DVDD.n22338 0.00393493
R49925 DVDD.n31 DVDD.n7 0.00393493
R49926 DVDD.n22341 DVDD.n22340 0.00393493
R49927 DVDD.n30 DVDD.n6 0.00393493
R49928 DVDD.n19697 DVDD.n19206 0.00393493
R49929 DVDD.n19212 DVDD.n19211 0.00393493
R49930 DVDD.n19698 DVDD.n19205 0.00393493
R49931 DVDD.n19214 DVDD.n19213 0.00393493
R49932 DVDD.n19702 DVDD.n19187 0.00393493
R49933 DVDD.n19634 DVDD.n19204 0.00393493
R49934 DVDD.n19637 DVDD.n19204 0.00393493
R49935 DVDD.n19636 DVDD.n19203 0.00393493
R49936 DVDD.n19203 DVDD.n19202 0.00393493
R49937 DVDD.n29 DVDD.n19 0.00393493
R49938 DVDD.n29 DVDD.n28 0.00393493
R49939 DVDD.n21 DVDD.n9 0.00393493
R49940 DVDD.n10 DVDD.n9 0.00393493
R49941 DVDD.n11 DVDD.n10 0.00393493
R49942 DVDD.n28 DVDD.n12 0.00393493
R49943 DVDD.n21 DVDD.n12 0.00393493
R49944 DVDD.n22343 DVDD.n19 0.00393493
R49945 DVDD.n19202 DVDD.n18653 0.00393493
R49946 DVDD.n19700 DVDD.n19637 0.00393493
R49947 DVDD.n19700 DVDD.n19636 0.00393493
R49948 DVDD.n19635 DVDD.n19634 0.00393493
R49949 DVDD.n3613 DVDD.n3531 0.00393125
R49950 DVDD.n15538 DVDD.n2660 0.00392439
R49951 DVDD.n5184 DVDD.n2727 0.00392439
R49952 DVDD.n3104 DVDD.n2997 0.00392439
R49953 DVDD.n16011 DVDD.n3012 0.00392439
R49954 DVDD.n15537 DVDD.n2585 0.00392439
R49955 DVDD.n5183 DVDD.n2797 0.00392439
R49956 DVDD.n3103 DVDD.n2926 0.00392439
R49957 DVDD.n16010 DVDD.n2941 0.00392439
R49958 DVDD.n15541 DVDD.n3250 0.00392439
R49959 DVDD.n5187 DVDD.n3167 0.00392439
R49960 DVDD.n16071 DVDD.n3059 0.00392439
R49961 DVDD.n16014 DVDD.n3070 0.00392439
R49962 DVDD.n15544 DVDD.n15543 0.00392439
R49963 DVDD.n5190 DVDD.n5189 0.00392439
R49964 DVDD.n16069 DVDD.n3107 0.00392439
R49965 DVDD.n16018 DVDD.n16016 0.00392439
R49966 DVDD.n4636 DVDD.n4214 0.00392
R49967 DVDD.n18155 DVDD 0.00392
R49968 DVDD.n2902 DVDD 0.00392
R49969 DVDD.n16221 DVDD 0.00392
R49970 DVDD.n16342 DVDD 0.00392
R49971 DVDD.n2546 DVDD 0.00392
R49972 DVDD.n2477 DVDD.n2476 0.00392
R49973 DVDD.n16284 DVDD.n2623 0.00392
R49974 DVDD.n2846 DVDD.n2825 0.00392
R49975 DVDD.n2987 DVDD.n2966 0.00392
R49976 DVDD.n5009 DVDD.n3517 0.00391053
R49977 DVDD.n5299 DVDD.n5074 0.00391053
R49978 DVDD.n5331 DVDD.n5238 0.00391053
R49979 DVDD.n5349 DVDD.n5249 0.00391053
R49980 DVDD.n5415 DVDD.n5392 0.00391053
R49981 DVDD.n5406 DVDD.n5383 0.00391053
R49982 DVDD.n18016 DVDD.n538 0.00391053
R49983 DVDD.n631 DVDD.n585 0.00391053
R49984 DVDD.n693 DVDD.n674 0.00391053
R49985 DVDD.n711 DVDD.n659 0.00391053
R49986 DVDD.n17949 DVDD.n771 0.00391053
R49987 DVDD.n17906 DVDD.n762 0.00391053
R49988 DVDD.n3590 DVDD.n3556 0.00389
R49989 DVDD.n15732 DVDD.n4903 0.00389
R49990 DVDD.n15697 DVDD.n5045 0.00389
R49991 DVDD.n15441 DVDD.n5259 0.00389
R49992 DVDD.n15405 DVDD.n5370 0.00389
R49993 DVDD.n15071 DVDD.n7059 0.00388255
R49994 DVDD.n7613 DVDD.n7568 0.00388255
R49995 DVDD.n15072 DVDD.n7061 0.00388255
R49996 DVDD.n9569 DVDD.n9568 0.00388255
R49997 DVDD.n4432 DVDD.n3749 0.003875
R49998 DVDD.n4177 DVDD.n3768 0.00386
R49999 DVDD.n4643 DVDD.n4223 0.00386
R50000 DVDD.n15837 DVDD.n3405 0.00386
R50001 DVDD.n2489 DVDD.n2481 0.00386
R50002 DVDD.n3312 DVDD.n3294 0.00386
R50003 DVDD.n16300 DVDD.n2628 0.00386
R50004 DVDD.n15938 DVDD.n3200 0.00386
R50005 DVDD.n2836 DVDD.n2830 0.00386
R50006 DVDD.n16075 DVDD.n3057 0.00386
R50007 DVDD.n16174 DVDD.n2971 0.00386
R50008 DVDD.n20182 DVDD.n19734 0.00384286
R50009 DVDD.n20257 DVDD.n19936 0.00384286
R50010 DVDD.n20674 DVDD.n18840 0.00384286
R50011 DVDD.n20749 DVDD.n19046 0.00384286
R50012 DVDD.n3997 DVDD.n3871 0.00384286
R50013 DVDD.n299 DVDD.n290 0.00384286
R50014 DVDD.n9823 DVDD.n9765 0.00384286
R50015 DVDD.n10069 DVDD.n10068 0.00384286
R50016 DVDD.n19676 DVDD.n18682 0.00384286
R50017 DVDD.n118 DVDD.n98 0.00384286
R50018 DVDD.n14827 DVDD.n8042 0.00384061
R50019 DVDD.n14828 DVDD.n8040 0.00384061
R50020 DVDD.n16398 DVDD.n2306 0.00383659
R50021 DVDD.n2473 DVDD.n2390 0.00383659
R50022 DVDD.n4977 DVDD.n3348 0.00383659
R50023 DVDD.n4980 DVDD.n3420 0.00383659
R50024 DVDD.n18477 DVDD.n18457 0.00383
R50025 DVDD.n21879 DVDD.n21838 0.00383
R50026 DVDD.n21895 DVDD.n21830 0.00383
R50027 DVDD.n21254 DVDD.n21253 0.00383
R50028 DVDD.n21949 DVDD.n198 0.00383
R50029 DVDD.n21978 DVDD.n204 0.00383
R50030 DVDD.n21232 DVDD.n21223 0.00383
R50031 DVDD.n18324 DVDD.n18294 0.00383
R50032 DVDD.n18351 DVDD.n18330 0.00383
R50033 DVDD.n18493 DVDD.n18492 0.00383
R50034 DVDD.n21860 DVDD.n21841 0.00383
R50035 DVDD.n21913 DVDD.n21912 0.00383
R50036 DVDD.n18159 DVDD.n448 0.00383
R50037 DVDD.n2541 DVDD.n504 0.00383
R50038 DVDD.n16337 DVDD.n559 0.00383
R50039 DVDD.n16216 DVDD.n646 0.00383
R50040 DVDD.n2897 DVDD.n732 0.00383
R50041 DVDD.n3604 DVDD.n3527 0.00381875
R50042 DVDD.n4134 DVDD.n4079 0.0038
R50043 DVDD.n4534 DVDD.n4203 0.0038
R50044 DVDD.n4697 DVDD.n4202 0.0038
R50045 DVDD.n16136 DVDD.n16134 0.0038
R50046 DVDD.n16259 DVDD.n2708 0.0038
R50047 DVDD.n15879 DVDD.n2702 0.0038
R50048 DVDD.n15878 DVDD.n15877 0.0038
R50049 DVDD.n15791 DVDD.n3481 0.0038
R50050 DVDD.n15876 DVDD.n2336 0.0038
R50051 DVDD.n15653 DVDD.n15600 0.0038
R50052 DVDD.n2701 DVDD.n2686 0.0038
R50053 DVDD.n15520 DVDD.n15519 0.0038
R50054 DVDD.n16258 DVDD.n2710 0.0038
R50055 DVDD.n15366 DVDD.n3109 0.0038
R50056 DVDD.n16135 DVDD.n3027 0.0038
R50057 DVDD.n20357 DVDD.n18939 0.00377857
R50058 DVDD.n19003 DVDD.n18967 0.00377857
R50059 DVDD.n22123 DVDD.n22122 0.00377857
R50060 DVDD.n10040 DVDD.n799 0.00377857
R50061 DVDD.n34 DVDD.n26 0.00377857
R50062 DVDD.n18144 DVDD.n452 0.00377
R50063 DVDD.n2555 DVDD.n508 0.00377
R50064 DVDD.n16351 DVDD.n555 0.00377
R50065 DVDD.n16230 DVDD.n642 0.00377
R50066 DVDD.n2911 DVDD.n736 0.00377
R50067 DVDD.n20164 DVDD.n20121 0.00376842
R50068 DVDD.n20118 DVDD.n20060 0.00376842
R50069 DVDD.n20116 DVDD.n20069 0.00376842
R50070 DVDD.n20114 DVDD.n20061 0.00376842
R50071 DVDD.n20112 DVDD.n20068 0.00376842
R50072 DVDD.n20110 DVDD.n20062 0.00376842
R50073 DVDD.n20108 DVDD.n20067 0.00376842
R50074 DVDD.n20106 DVDD.n20063 0.00376842
R50075 DVDD.n20104 DVDD.n20066 0.00376842
R50076 DVDD.n20102 DVDD.n20064 0.00376842
R50077 DVDD.n20100 DVDD.n20065 0.00376842
R50078 DVDD.n20885 DVDD.n18929 0.00376842
R50079 DVDD.n20884 DVDD.n18937 0.00376842
R50080 DVDD.n20882 DVDD.n20881 0.00376842
R50081 DVDD.n20878 DVDD.n18946 0.00376842
R50082 DVDD.n20876 DVDD.n18956 0.00376842
R50083 DVDD.n20874 DVDD.n18947 0.00376842
R50084 DVDD.n20872 DVDD.n18955 0.00376842
R50085 DVDD.n20870 DVDD.n18948 0.00376842
R50086 DVDD.n20868 DVDD.n18954 0.00376842
R50087 DVDD.n20866 DVDD.n18949 0.00376842
R50088 DVDD.n20864 DVDD.n18953 0.00376842
R50089 DVDD DVDD.n22229 0.00376574
R50090 DVDD.n18432 DVDD 0.00376574
R50091 DVDD.n22039 DVDD 0.00376574
R50092 DVDD DVDD.n223 0.00376574
R50093 DVDD.n4596 DVDD.n4245 0.0037625
R50094 DVDD.n4558 DVDD.n4319 0.0037625
R50095 DVDD.n4385 DVDD.n4325 0.00374878
R50096 DVDD.n4351 DVDD.n4255 0.00374878
R50097 DVDD.n4362 DVDD.n3724 0.00374878
R50098 DVDD.n4371 DVDD.n3643 0.00374878
R50099 DVDD.n10697 DVDD.n10238 0.00374812
R50100 DVDD.n17276 DVDD.n17275 0.00374812
R50101 DVDD.n17727 DVDD.n890 0.00374812
R50102 DVDD.n4118 DVDD.n4083 0.00374
R50103 DVDD.n4494 DVDD.n4191 0.00374
R50104 DVDD.n15774 DVDD.n3485 0.00374
R50105 DVDD.n15858 DVDD.n2340 0.00374
R50106 DVDD.n15626 DVDD.n15604 0.00374
R50107 DVDD.n15892 DVDD.n2690 0.00374
R50108 DVDD.n15483 DVDD.n5134 0.00374
R50109 DVDD.n15972 DVDD.n2751 0.00374
R50110 DVDD.n15380 DVDD.n3113 0.00374
R50111 DVDD.n16118 DVDD.n3031 0.00374
R50112 DVDD.n18373 DVDD.n18308 0.00373291
R50113 DVDD.n21262 DVDD.n18659 0.00373291
R50114 DVDD.n18349 DVDD.n18348 0.00373291
R50115 DVDD.n4865 DVDD.n3536 0.00373291
R50116 DVDD.n5007 DVDD.n3518 0.00372105
R50117 DVDD.n5301 DVDD.n5075 0.00372105
R50118 DVDD.n5333 DVDD.n5237 0.00372105
R50119 DVDD.n5347 DVDD.n5248 0.00372105
R50120 DVDD.n5413 DVDD.n5393 0.00372105
R50121 DVDD.n18018 DVDD.n539 0.00372105
R50122 DVDD.n633 DVDD.n593 0.00372105
R50123 DVDD.n695 DVDD.n661 0.00372105
R50124 DVDD.n709 DVDD.n672 0.00372105
R50125 DVDD.n17953 DVDD.n17952 0.00372105
R50126 DVDD.n20443 DVDD.n19820 0.00372031
R50127 DVDD.n20464 DVDD.n19810 0.00372031
R50128 DVDD.n20480 DVDD.n19033 0.00372031
R50129 DVDD.n19034 DVDD.n19023 0.00372031
R50130 DVDD.n19056 DVDD.n19030 0.00372031
R50131 DVDD.n19055 DVDD.n19029 0.00372031
R50132 DVDD.n21052 DVDD.n18772 0.00372031
R50133 DVDD.n22250 DVDD.n22249 0.00372031
R50134 DVDD.n113 DVDD.n91 0.00372031
R50135 DVDD.n22248 DVDD.n22247 0.00372031
R50136 DVDD.n114 DVDD.n92 0.00372031
R50137 DVDD.n116 DVDD.n115 0.00372031
R50138 DVDD.n22246 DVDD.n95 0.00372031
R50139 DVDD.n22245 DVDD.n117 0.00372031
R50140 DVDD.n22244 DVDD.n94 0.00372031
R50141 DVDD.n319 DVDD.n314 0.00372031
R50142 DVDD.n318 DVDD.n313 0.00372031
R50143 DVDD.n317 DVDD.n312 0.00372031
R50144 DVDD.n316 DVDD.n311 0.00372031
R50145 DVDD.n22159 DVDD.n291 0.00372031
R50146 DVDD.n4506 DVDD.n4463 0.00372031
R50147 DVDD.n4533 DVDD.n4489 0.00372031
R50148 DVDD.n4490 DVDD.n4464 0.00372031
R50149 DVDD.n4527 DVDD.n4488 0.00372031
R50150 DVDD.n4507 DVDD.n4465 0.00372031
R50151 DVDD.n4526 DVDD.n4487 0.00372031
R50152 DVDD.n4508 DVDD.n4466 0.00372031
R50153 DVDD.n4525 DVDD.n4486 0.00372031
R50154 DVDD.n4509 DVDD.n4467 0.00372031
R50155 DVDD.n4524 DVDD.n4485 0.00372031
R50156 DVDD.n4510 DVDD.n4468 0.00372031
R50157 DVDD.n4523 DVDD.n4484 0.00372031
R50158 DVDD.n4511 DVDD.n4469 0.00372031
R50159 DVDD.n4522 DVDD.n4483 0.00372031
R50160 DVDD.n4512 DVDD.n4470 0.00372031
R50161 DVDD.n4521 DVDD.n4482 0.00372031
R50162 DVDD.n4513 DVDD.n4471 0.00372031
R50163 DVDD.n4520 DVDD.n4481 0.00372031
R50164 DVDD.n4514 DVDD.n4472 0.00372031
R50165 DVDD.n4519 DVDD.n4480 0.00372031
R50166 DVDD.n4515 DVDD.n4473 0.00372031
R50167 DVDD.n4518 DVDD.n4479 0.00372031
R50168 DVDD.n4531 DVDD.n4517 0.00372031
R50169 DVDD.n4330 DVDD.n4328 0.00372031
R50170 DVDD.n16393 DVDD.n16391 0.00372031
R50171 DVDD.n16392 DVDD.n2351 0.00372031
R50172 DVDD.n16389 DVDD.n2377 0.00372031
R50173 DVDD.n2376 DVDD.n2296 0.00372031
R50174 DVDD.n2375 DVDD.n2334 0.00372031
R50175 DVDD.n2374 DVDD.n2352 0.00372031
R50176 DVDD.n16388 DVDD.n2373 0.00372031
R50177 DVDD.n2372 DVDD.n2353 0.00372031
R50178 DVDD.n16387 DVDD.n2371 0.00372031
R50179 DVDD.n2370 DVDD.n2354 0.00372031
R50180 DVDD.n16386 DVDD.n2369 0.00372031
R50181 DVDD.n16385 DVDD.n2368 0.00372031
R50182 DVDD.n2367 DVDD.n2356 0.00372031
R50183 DVDD.n16384 DVDD.n2366 0.00372031
R50184 DVDD.n16383 DVDD.n2365 0.00372031
R50185 DVDD.n2364 DVDD.n2358 0.00372031
R50186 DVDD.n16382 DVDD.n2363 0.00372031
R50187 DVDD.n2678 DVDD.n2677 0.00372031
R50188 DVDD.n2679 DVDD.n2646 0.00372031
R50189 DVDD.n2676 DVDD.n2675 0.00372031
R50190 DVDD.n2674 DVDD.n2673 0.00372031
R50191 DVDD.n2680 DVDD.n2648 0.00372031
R50192 DVDD.n2672 DVDD.n2671 0.00372031
R50193 DVDD.n2670 DVDD.n2669 0.00372031
R50194 DVDD.n2681 DVDD.n2650 0.00372031
R50195 DVDD.n2668 DVDD.n2667 0.00372031
R50196 DVDD.n2666 DVDD.n2665 0.00372031
R50197 DVDD.n2682 DVDD.n2652 0.00372031
R50198 DVDD.n2664 DVDD.n2663 0.00372031
R50199 DVDD.n2662 DVDD.n2661 0.00372031
R50200 DVDD.n2683 DVDD.n2654 0.00372031
R50201 DVDD.n2660 DVDD.n2659 0.00372031
R50202 DVDD.n2684 DVDD.n2658 0.00372031
R50203 DVDD.n2657 DVDD.n2656 0.00372031
R50204 DVDD.n2747 DVDD.n2711 0.00372031
R50205 DVDD.n2745 DVDD.n2733 0.00372031
R50206 DVDD.n2744 DVDD.n2732 0.00372031
R50207 DVDD.n2758 DVDD.n2713 0.00372031
R50208 DVDD.n2743 DVDD.n2731 0.00372031
R50209 DVDD.n2759 DVDD.n2714 0.00372031
R50210 DVDD.n2742 DVDD.n2730 0.00372031
R50211 DVDD.n2760 DVDD.n2715 0.00372031
R50212 DVDD.n2741 DVDD.n2729 0.00372031
R50213 DVDD.n2740 DVDD.n2728 0.00372031
R50214 DVDD.n2761 DVDD.n2717 0.00372031
R50215 DVDD.n2739 DVDD.n2727 0.00372031
R50216 DVDD.n2738 DVDD.n2726 0.00372031
R50217 DVDD.n2762 DVDD.n2719 0.00372031
R50218 DVDD.n2737 DVDD.n2725 0.00372031
R50219 DVDD.n2736 DVDD.n2724 0.00372031
R50220 DVDD.n2763 DVDD.n2721 0.00372031
R50221 DVDD.n2735 DVDD.n2723 0.00372031
R50222 DVDD.n3022 DVDD.n3021 0.00372031
R50223 DVDD.n3019 DVDD.n3018 0.00372031
R50224 DVDD.n3016 DVDD.n3015 0.00372031
R50225 DVDD.n3013 DVDD.n3004 0.00372031
R50226 DVDD.n3011 DVDD.n3010 0.00372031
R50227 DVDD.n3008 DVDD.n3007 0.00372031
R50228 DVDD.n9679 DVDD.n9672 0.00372031
R50229 DVDD.n9678 DVDD.n9666 0.00372031
R50230 DVDD.n18772 DVDD.n18770 0.00372031
R50231 DVDD.n20480 DVDD.n20465 0.00372031
R50232 DVDD.n19820 DVDD.n19810 0.00372031
R50233 DVDD.n20462 DVDD.n20443 0.00372031
R50234 DVDD.n9678 DVDD.n9670 0.00372031
R50235 DVDD.n9679 DVDD.n9664 0.00372031
R50236 DVDD.n3009 DVDD.n3008 0.00372031
R50237 DVDD.n3010 DVDD.n3005 0.00372031
R50238 DVDD.n3014 DVDD.n3013 0.00372031
R50239 DVDD.n3015 DVDD.n3002 0.00372031
R50240 DVDD.n3018 DVDD.n3000 0.00372031
R50241 DVDD.n3021 DVDD.n2998 0.00372031
R50242 DVDD.n2735 DVDD.n2721 0.00372031
R50243 DVDD.n2763 DVDD.n2724 0.00372031
R50244 DVDD.n2736 DVDD.n2720 0.00372031
R50245 DVDD.n2737 DVDD.n2719 0.00372031
R50246 DVDD.n2762 DVDD.n2726 0.00372031
R50247 DVDD.n2738 DVDD.n2718 0.00372031
R50248 DVDD.n2739 DVDD.n2717 0.00372031
R50249 DVDD.n2761 DVDD.n2728 0.00372031
R50250 DVDD.n2740 DVDD.n2716 0.00372031
R50251 DVDD.n2741 DVDD.n2715 0.00372031
R50252 DVDD.n2760 DVDD.n2730 0.00372031
R50253 DVDD.n2742 DVDD.n2714 0.00372031
R50254 DVDD.n2759 DVDD.n2731 0.00372031
R50255 DVDD.n2743 DVDD.n2713 0.00372031
R50256 DVDD.n2758 DVDD.n2732 0.00372031
R50257 DVDD.n2744 DVDD.n2712 0.00372031
R50258 DVDD.n2745 DVDD.n2711 0.00372031
R50259 DVDD.n16256 DVDD.n2747 0.00372031
R50260 DVDD.n2658 DVDD.n2657 0.00372031
R50261 DVDD.n2684 DVDD.n2655 0.00372031
R50262 DVDD.n2659 DVDD.n2654 0.00372031
R50263 DVDD.n2683 DVDD.n2662 0.00372031
R50264 DVDD.n2661 DVDD.n2653 0.00372031
R50265 DVDD.n2663 DVDD.n2652 0.00372031
R50266 DVDD.n2682 DVDD.n2666 0.00372031
R50267 DVDD.n2665 DVDD.n2651 0.00372031
R50268 DVDD.n2667 DVDD.n2650 0.00372031
R50269 DVDD.n2681 DVDD.n2670 0.00372031
R50270 DVDD.n2669 DVDD.n2649 0.00372031
R50271 DVDD.n2671 DVDD.n2648 0.00372031
R50272 DVDD.n2680 DVDD.n2674 0.00372031
R50273 DVDD.n2673 DVDD.n2647 0.00372031
R50274 DVDD.n2675 DVDD.n2646 0.00372031
R50275 DVDD.n2679 DVDD.n2678 0.00372031
R50276 DVDD.n2677 DVDD.n2645 0.00372031
R50277 DVDD.n16382 DVDD.n2358 0.00372031
R50278 DVDD.n2365 DVDD.n2364 0.00372031
R50279 DVDD.n16383 DVDD.n2357 0.00372031
R50280 DVDD.n16384 DVDD.n2356 0.00372031
R50281 DVDD.n2368 DVDD.n2367 0.00372031
R50282 DVDD.n16385 DVDD.n2355 0.00372031
R50283 DVDD.n16386 DVDD.n2354 0.00372031
R50284 DVDD.n2371 DVDD.n2370 0.00372031
R50285 DVDD.n16387 DVDD.n2353 0.00372031
R50286 DVDD.n2373 DVDD.n2372 0.00372031
R50287 DVDD.n16388 DVDD.n2352 0.00372031
R50288 DVDD.n2375 DVDD.n2374 0.00372031
R50289 DVDD.n16395 DVDD.n2334 0.00372031
R50290 DVDD.n2377 DVDD.n2376 0.00372031
R50291 DVDD.n16389 DVDD.n2351 0.00372031
R50292 DVDD.n16393 DVDD.n16392 0.00372031
R50293 DVDD.n16391 DVDD.n2350 0.00372031
R50294 DVDD.n4331 DVDD.n4330 0.00372031
R50295 DVDD.n4517 DVDD.n4479 0.00372031
R50296 DVDD.n4518 DVDD.n4473 0.00372031
R50297 DVDD.n4515 DVDD.n4480 0.00372031
R50298 DVDD.n4519 DVDD.n4472 0.00372031
R50299 DVDD.n4514 DVDD.n4481 0.00372031
R50300 DVDD.n4520 DVDD.n4471 0.00372031
R50301 DVDD.n4513 DVDD.n4482 0.00372031
R50302 DVDD.n4521 DVDD.n4470 0.00372031
R50303 DVDD.n4512 DVDD.n4483 0.00372031
R50304 DVDD.n4522 DVDD.n4469 0.00372031
R50305 DVDD.n4511 DVDD.n4484 0.00372031
R50306 DVDD.n4523 DVDD.n4468 0.00372031
R50307 DVDD.n4510 DVDD.n4485 0.00372031
R50308 DVDD.n4524 DVDD.n4467 0.00372031
R50309 DVDD.n4509 DVDD.n4486 0.00372031
R50310 DVDD.n4525 DVDD.n4466 0.00372031
R50311 DVDD.n4508 DVDD.n4487 0.00372031
R50312 DVDD.n4526 DVDD.n4465 0.00372031
R50313 DVDD.n4507 DVDD.n4488 0.00372031
R50314 DVDD.n4527 DVDD.n4464 0.00372031
R50315 DVDD.n4533 DVDD.n4490 0.00372031
R50316 DVDD.n4489 DVDD.n4463 0.00372031
R50317 DVDD.n4506 DVDD.n298 0.00372031
R50318 DVDD.n309 DVDD.n291 0.00372031
R50319 DVDD.n316 DVDD.n308 0.00372031
R50320 DVDD.n317 DVDD.n307 0.00372031
R50321 DVDD.n318 DVDD.n306 0.00372031
R50322 DVDD.n319 DVDD.n305 0.00372031
R50323 DVDD.n19055 DVDD.n19026 0.00372031
R50324 DVDD.n19056 DVDD.n19025 0.00372031
R50325 DVDD.n20778 DVDD.n19034 0.00372031
R50326 DVDD.n20926 DVDD.n18905 0.00372031
R50327 DVDD.n20927 DVDD.n18889 0.00372031
R50328 DVDD.n18888 DVDD.n18871 0.00372031
R50329 DVDD.n18903 DVDD.n18890 0.00372031
R50330 DVDD.n18902 DVDD.n18900 0.00372031
R50331 DVDD.n18901 DVDD.n18891 0.00372031
R50332 DVDD.n18899 DVDD.n18897 0.00372031
R50333 DVDD.n18898 DVDD.n18892 0.00372031
R50334 DVDD.n19096 DVDD.n18819 0.00372031
R50335 DVDD.n70 DVDD.n56 0.00372031
R50336 DVDD.n55 DVDD.n44 0.00372031
R50337 DVDD.n69 DVDD.n54 0.00372031
R50338 DVDD.n53 DVDD.n45 0.00372031
R50339 DVDD.n67 DVDD.n46 0.00372031
R50340 DVDD.n51 DVDD.n50 0.00372031
R50341 DVDD.n68 DVDD.n47 0.00372031
R50342 DVDD.n49 DVDD.n48 0.00372031
R50343 DVDD.n373 DVDD.n355 0.00372031
R50344 DVDD.n371 DVDD.n365 0.00372031
R50345 DVDD.n422 DVDD.n356 0.00372031
R50346 DVDD.n370 DVDD.n364 0.00372031
R50347 DVDD.n423 DVDD.n357 0.00372031
R50348 DVDD.n369 DVDD.n363 0.00372031
R50349 DVDD.n424 DVDD.n358 0.00372031
R50350 DVDD.n368 DVDD.n362 0.00372031
R50351 DVDD.n425 DVDD.n359 0.00372031
R50352 DVDD.n367 DVDD.n361 0.00372031
R50353 DVDD.n4614 DVDD.n4229 0.00372031
R50354 DVDD.n4625 DVDD.n4613 0.00372031
R50355 DVDD.n4644 DVDD.n4230 0.00372031
R50356 DVDD.n4624 DVDD.n4612 0.00372031
R50357 DVDD.n4645 DVDD.n4231 0.00372031
R50358 DVDD.n4623 DVDD.n4611 0.00372031
R50359 DVDD.n4646 DVDD.n4232 0.00372031
R50360 DVDD.n4622 DVDD.n4610 0.00372031
R50361 DVDD.n4647 DVDD.n4233 0.00372031
R50362 DVDD.n4621 DVDD.n4609 0.00372031
R50363 DVDD.n4648 DVDD.n4234 0.00372031
R50364 DVDD.n4620 DVDD.n4608 0.00372031
R50365 DVDD.n4649 DVDD.n4235 0.00372031
R50366 DVDD.n4619 DVDD.n4607 0.00372031
R50367 DVDD.n4650 DVDD.n4236 0.00372031
R50368 DVDD.n4618 DVDD.n4606 0.00372031
R50369 DVDD.n4651 DVDD.n4237 0.00372031
R50370 DVDD.n4617 DVDD.n4605 0.00372031
R50371 DVDD.n4652 DVDD.n4238 0.00372031
R50372 DVDD.n4616 DVDD.n4604 0.00372031
R50373 DVDD.n4653 DVDD.n4239 0.00372031
R50374 DVDD.n4615 DVDD.n4603 0.00372031
R50375 DVDD.n4654 DVDD.n4602 0.00372031
R50376 DVDD.n4270 DVDD.n4257 0.00372031
R50377 DVDD.n4262 DVDD.n4259 0.00372031
R50378 DVDD.n2423 DVDD.n2411 0.00372031
R50379 DVDD.n2425 DVDD.n2392 0.00372031
R50380 DVDD.n2422 DVDD.n2410 0.00372031
R50381 DVDD.n2431 DVDD.n2412 0.00372031
R50382 DVDD.n2421 DVDD.n2409 0.00372031
R50383 DVDD.n2426 DVDD.n2394 0.00372031
R50384 DVDD.n2420 DVDD.n2408 0.00372031
R50385 DVDD.n2427 DVDD.n2395 0.00372031
R50386 DVDD.n2419 DVDD.n2407 0.00372031
R50387 DVDD.n2428 DVDD.n2396 0.00372031
R50388 DVDD.n2418 DVDD.n2406 0.00372031
R50389 DVDD.n2417 DVDD.n2405 0.00372031
R50390 DVDD.n2429 DVDD.n2398 0.00372031
R50391 DVDD.n2416 DVDD.n2404 0.00372031
R50392 DVDD.n2415 DVDD.n2403 0.00372031
R50393 DVDD.n2430 DVDD.n2400 0.00372031
R50394 DVDD.n2414 DVDD.n2402 0.00372031
R50395 DVDD.n2605 DVDD.n2594 0.00372031
R50396 DVDD.n2607 DVDD.n2573 0.00372031
R50397 DVDD.n2604 DVDD.n2593 0.00372031
R50398 DVDD.n2603 DVDD.n2592 0.00372031
R50399 DVDD.n2608 DVDD.n2575 0.00372031
R50400 DVDD.n2602 DVDD.n2591 0.00372031
R50401 DVDD.n2601 DVDD.n2590 0.00372031
R50402 DVDD.n2609 DVDD.n2577 0.00372031
R50403 DVDD.n2600 DVDD.n2589 0.00372031
R50404 DVDD.n2599 DVDD.n2588 0.00372031
R50405 DVDD.n2610 DVDD.n2579 0.00372031
R50406 DVDD.n2598 DVDD.n2587 0.00372031
R50407 DVDD.n2597 DVDD.n2586 0.00372031
R50408 DVDD.n2611 DVDD.n2581 0.00372031
R50409 DVDD.n2596 DVDD.n2585 0.00372031
R50410 DVDD.n2612 DVDD.n2584 0.00372031
R50411 DVDD.n2595 DVDD.n2583 0.00372031
R50412 DVDD.n2817 DVDD.n2780 0.00372031
R50413 DVDD.n2815 DVDD.n2803 0.00372031
R50414 DVDD.n2814 DVDD.n2802 0.00372031
R50415 DVDD.n2866 DVDD.n2782 0.00372031
R50416 DVDD.n2813 DVDD.n2801 0.00372031
R50417 DVDD.n2867 DVDD.n2783 0.00372031
R50418 DVDD.n2812 DVDD.n2800 0.00372031
R50419 DVDD.n2868 DVDD.n2784 0.00372031
R50420 DVDD.n2811 DVDD.n2799 0.00372031
R50421 DVDD.n2810 DVDD.n2798 0.00372031
R50422 DVDD.n2869 DVDD.n2786 0.00372031
R50423 DVDD.n2809 DVDD.n2797 0.00372031
R50424 DVDD.n2808 DVDD.n2796 0.00372031
R50425 DVDD.n2870 DVDD.n2788 0.00372031
R50426 DVDD.n2807 DVDD.n2795 0.00372031
R50427 DVDD.n2806 DVDD.n2794 0.00372031
R50428 DVDD.n2871 DVDD.n2790 0.00372031
R50429 DVDD.n2805 DVDD.n2793 0.00372031
R50430 DVDD.n2953 DVDD.n2927 0.00372031
R50431 DVDD.n2978 DVDD.n2952 0.00372031
R50432 DVDD.n2951 DVDD.n2928 0.00372031
R50433 DVDD.n2949 DVDD.n2929 0.00372031
R50434 DVDD.n2977 DVDD.n2948 0.00372031
R50435 DVDD.n2947 DVDD.n2930 0.00372031
R50436 DVDD.n2973 DVDD.n2931 0.00372031
R50437 DVDD.n2945 DVDD.n2944 0.00372031
R50438 DVDD.n2979 DVDD.n2955 0.00372031
R50439 DVDD.n2976 DVDD.n2943 0.00372031
R50440 DVDD.n2942 DVDD.n2933 0.00372031
R50441 DVDD.n2972 DVDD.n2925 0.00372031
R50442 DVDD.n2974 DVDD.n2934 0.00372031
R50443 DVDD.n2940 DVDD.n2939 0.00372031
R50444 DVDD.n16183 DVDD.n2956 0.00372031
R50445 DVDD.n2975 DVDD.n2938 0.00372031
R50446 DVDD.n2937 DVDD.n2936 0.00372031
R50447 DVDD.n9749 DVDD.n9745 0.00372031
R50448 DVDD.n9999 DVDD.n9735 0.00372031
R50449 DVDD.n9748 DVDD.n9743 0.00372031
R50450 DVDD.n9998 DVDD.n9733 0.00372031
R50451 DVDD.n10000 DVDD.n9742 0.00372031
R50452 DVDD.n9747 DVDD.n9737 0.00372031
R50453 DVDD.n10056 DVDD.n9746 0.00372031
R50454 DVDD.n19101 DVDD.n19096 0.00372031
R50455 DVDD.n20923 DVDD.n18905 0.00372031
R50456 DVDD.n9746 DVDD.n9737 0.00372031
R50457 DVDD.n9747 DVDD.n9742 0.00372031
R50458 DVDD.n10000 DVDD.n9736 0.00372031
R50459 DVDD.n9998 DVDD.n9743 0.00372031
R50460 DVDD.n9748 DVDD.n9735 0.00372031
R50461 DVDD.n9999 DVDD.n9744 0.00372031
R50462 DVDD.n9749 DVDD.n9734 0.00372031
R50463 DVDD.n2938 DVDD.n2937 0.00372031
R50464 DVDD.n2975 DVDD.n2935 0.00372031
R50465 DVDD.n2956 DVDD.n2940 0.00372031
R50466 DVDD.n2939 DVDD.n2934 0.00372031
R50467 DVDD.n2974 DVDD.n2941 0.00372031
R50468 DVDD.n2972 DVDD.n2933 0.00372031
R50469 DVDD.n2943 DVDD.n2942 0.00372031
R50470 DVDD.n2976 DVDD.n2932 0.00372031
R50471 DVDD.n2979 DVDD.n2945 0.00372031
R50472 DVDD.n2944 DVDD.n2931 0.00372031
R50473 DVDD.n2973 DVDD.n2946 0.00372031
R50474 DVDD.n2948 DVDD.n2947 0.00372031
R50475 DVDD.n2977 DVDD.n2929 0.00372031
R50476 DVDD.n2950 DVDD.n2949 0.00372031
R50477 DVDD.n2952 DVDD.n2951 0.00372031
R50478 DVDD.n2978 DVDD.n2927 0.00372031
R50479 DVDD.n2954 DVDD.n2953 0.00372031
R50480 DVDD.n2805 DVDD.n2790 0.00372031
R50481 DVDD.n2871 DVDD.n2794 0.00372031
R50482 DVDD.n2806 DVDD.n2789 0.00372031
R50483 DVDD.n2807 DVDD.n2788 0.00372031
R50484 DVDD.n2870 DVDD.n2796 0.00372031
R50485 DVDD.n2808 DVDD.n2787 0.00372031
R50486 DVDD.n2809 DVDD.n2786 0.00372031
R50487 DVDD.n2869 DVDD.n2798 0.00372031
R50488 DVDD.n2810 DVDD.n2785 0.00372031
R50489 DVDD.n2811 DVDD.n2784 0.00372031
R50490 DVDD.n2868 DVDD.n2800 0.00372031
R50491 DVDD.n2812 DVDD.n2783 0.00372031
R50492 DVDD.n2867 DVDD.n2801 0.00372031
R50493 DVDD.n2813 DVDD.n2782 0.00372031
R50494 DVDD.n2866 DVDD.n2802 0.00372031
R50495 DVDD.n2814 DVDD.n2781 0.00372031
R50496 DVDD.n2815 DVDD.n2780 0.00372031
R50497 DVDD.n16247 DVDD.n2817 0.00372031
R50498 DVDD.n2595 DVDD.n2584 0.00372031
R50499 DVDD.n2612 DVDD.n2582 0.00372031
R50500 DVDD.n2596 DVDD.n2581 0.00372031
R50501 DVDD.n2611 DVDD.n2586 0.00372031
R50502 DVDD.n2597 DVDD.n2580 0.00372031
R50503 DVDD.n2598 DVDD.n2579 0.00372031
R50504 DVDD.n2610 DVDD.n2588 0.00372031
R50505 DVDD.n2599 DVDD.n2578 0.00372031
R50506 DVDD.n2600 DVDD.n2577 0.00372031
R50507 DVDD.n2609 DVDD.n2590 0.00372031
R50508 DVDD.n2601 DVDD.n2576 0.00372031
R50509 DVDD.n2602 DVDD.n2575 0.00372031
R50510 DVDD.n2608 DVDD.n2592 0.00372031
R50511 DVDD.n2603 DVDD.n2574 0.00372031
R50512 DVDD.n2604 DVDD.n2573 0.00372031
R50513 DVDD.n2607 DVDD.n2594 0.00372031
R50514 DVDD.n2605 DVDD.n2572 0.00372031
R50515 DVDD.n2414 DVDD.n2400 0.00372031
R50516 DVDD.n2430 DVDD.n2403 0.00372031
R50517 DVDD.n2415 DVDD.n2399 0.00372031
R50518 DVDD.n2416 DVDD.n2398 0.00372031
R50519 DVDD.n2429 DVDD.n2405 0.00372031
R50520 DVDD.n2417 DVDD.n2397 0.00372031
R50521 DVDD.n2418 DVDD.n2396 0.00372031
R50522 DVDD.n2428 DVDD.n2407 0.00372031
R50523 DVDD.n2419 DVDD.n2395 0.00372031
R50524 DVDD.n2427 DVDD.n2408 0.00372031
R50525 DVDD.n2420 DVDD.n2394 0.00372031
R50526 DVDD.n2426 DVDD.n2409 0.00372031
R50527 DVDD.n2421 DVDD.n2393 0.00372031
R50528 DVDD.n2431 DVDD.n2410 0.00372031
R50529 DVDD.n2422 DVDD.n2392 0.00372031
R50530 DVDD.n2425 DVDD.n2411 0.00372031
R50531 DVDD.n2423 DVDD.n2391 0.00372031
R50532 DVDD.n4259 DVDD.n4257 0.00372031
R50533 DVDD.n4599 DVDD.n4270 0.00372031
R50534 DVDD.n4654 DVDD.n4603 0.00372031
R50535 DVDD.n4615 DVDD.n4239 0.00372031
R50536 DVDD.n4653 DVDD.n4604 0.00372031
R50537 DVDD.n4616 DVDD.n4238 0.00372031
R50538 DVDD.n4652 DVDD.n4605 0.00372031
R50539 DVDD.n4617 DVDD.n4237 0.00372031
R50540 DVDD.n4651 DVDD.n4606 0.00372031
R50541 DVDD.n4618 DVDD.n4236 0.00372031
R50542 DVDD.n4650 DVDD.n4607 0.00372031
R50543 DVDD.n4619 DVDD.n4235 0.00372031
R50544 DVDD.n4649 DVDD.n4608 0.00372031
R50545 DVDD.n4620 DVDD.n4234 0.00372031
R50546 DVDD.n4648 DVDD.n4609 0.00372031
R50547 DVDD.n4621 DVDD.n4233 0.00372031
R50548 DVDD.n4647 DVDD.n4610 0.00372031
R50549 DVDD.n4622 DVDD.n4232 0.00372031
R50550 DVDD.n4646 DVDD.n4611 0.00372031
R50551 DVDD.n4623 DVDD.n4231 0.00372031
R50552 DVDD.n4645 DVDD.n4612 0.00372031
R50553 DVDD.n4624 DVDD.n4230 0.00372031
R50554 DVDD.n4644 DVDD.n4613 0.00372031
R50555 DVDD.n4625 DVDD.n4229 0.00372031
R50556 DVDD.n4658 DVDD.n4614 0.00372031
R50557 DVDD.n367 DVDD.n359 0.00372031
R50558 DVDD.n425 DVDD.n362 0.00372031
R50559 DVDD.n368 DVDD.n358 0.00372031
R50560 DVDD.n424 DVDD.n363 0.00372031
R50561 DVDD.n369 DVDD.n357 0.00372031
R50562 DVDD.n423 DVDD.n364 0.00372031
R50563 DVDD.n370 DVDD.n356 0.00372031
R50564 DVDD.n422 DVDD.n365 0.00372031
R50565 DVDD.n371 DVDD.n355 0.00372031
R50566 DVDD.n22139 DVDD.n373 0.00372031
R50567 DVDD.n18899 DVDD.n18898 0.00372031
R50568 DVDD.n18897 DVDD.n18891 0.00372031
R50569 DVDD.n18902 DVDD.n18901 0.00372031
R50570 DVDD.n18900 DVDD.n18890 0.00372031
R50571 DVDD.n18904 DVDD.n18903 0.00372031
R50572 DVDD.n18889 DVDD.n18888 0.00372031
R50573 DVDD.n20928 DVDD.n20927 0.00372031
R50574 DVDD.n19788 DVDD.n19767 0.00372031
R50575 DVDD.n20538 DVDD.n19790 0.00372031
R50576 DVDD.n19797 DVDD.n19129 0.00372031
R50577 DVDD.n19130 DVDD.n19074 0.00372031
R50578 DVDD.n19131 DVDD.n19128 0.00372031
R50579 DVDD.n19150 DVDD.n19076 0.00372031
R50580 DVDD.n19133 DVDD.n19126 0.00372031
R50581 DVDD.n19151 DVDD.n19077 0.00372031
R50582 DVDD.n19132 DVDD.n19125 0.00372031
R50583 DVDD.n19152 DVDD.n19078 0.00372031
R50584 DVDD.n21059 DVDD.n18754 0.00372031
R50585 DVDD.n21060 DVDD.n18735 0.00372031
R50586 DVDD.n21093 DVDD.n18734 0.00372031
R50587 DVDD.n21084 DVDD.n18725 0.00372031
R50588 DVDD.n21092 DVDD.n18733 0.00372031
R50589 DVDD.n21085 DVDD.n18726 0.00372031
R50590 DVDD.n21090 DVDD.n18727 0.00372031
R50591 DVDD.n21087 DVDD.n18731 0.00372031
R50592 DVDD.n21091 DVDD.n18728 0.00372031
R50593 DVDD.n21086 DVDD.n18730 0.00372031
R50594 DVDD.n252 DVDD.n237 0.00372031
R50595 DVDD.n22180 DVDD.n267 0.00372031
R50596 DVDD.n22179 DVDD.n253 0.00372031
R50597 DVDD.n266 DVDD.n265 0.00372031
R50598 DVDD.n269 DVDD.n254 0.00372031
R50599 DVDD.n264 DVDD.n263 0.00372031
R50600 DVDD.n270 DVDD.n255 0.00372031
R50601 DVDD.n262 DVDD.n261 0.00372031
R50602 DVDD.n271 DVDD.n256 0.00372031
R50603 DVDD.n260 DVDD.n258 0.00372031
R50604 DVDD.n3795 DVDD.n3772 0.00372031
R50605 DVDD.n3806 DVDD.n3794 0.00372031
R50606 DVDD.n4164 DVDD.n3773 0.00372031
R50607 DVDD.n3805 DVDD.n3793 0.00372031
R50608 DVDD.n4165 DVDD.n3774 0.00372031
R50609 DVDD.n3804 DVDD.n3792 0.00372031
R50610 DVDD.n4166 DVDD.n3775 0.00372031
R50611 DVDD.n3803 DVDD.n3791 0.00372031
R50612 DVDD.n4167 DVDD.n3776 0.00372031
R50613 DVDD.n3802 DVDD.n3790 0.00372031
R50614 DVDD.n4168 DVDD.n3777 0.00372031
R50615 DVDD.n3801 DVDD.n3789 0.00372031
R50616 DVDD.n4169 DVDD.n3778 0.00372031
R50617 DVDD.n3800 DVDD.n3788 0.00372031
R50618 DVDD.n4170 DVDD.n3779 0.00372031
R50619 DVDD.n3799 DVDD.n3787 0.00372031
R50620 DVDD.n4171 DVDD.n3780 0.00372031
R50621 DVDD.n3798 DVDD.n3786 0.00372031
R50622 DVDD.n4172 DVDD.n3781 0.00372031
R50623 DVDD.n3797 DVDD.n3785 0.00372031
R50624 DVDD.n4173 DVDD.n3782 0.00372031
R50625 DVDD.n3796 DVDD.n3784 0.00372031
R50626 DVDD.n4174 DVDD.n3783 0.00372031
R50627 DVDD.n3747 DVDD.n3726 0.00372031
R50628 DVDD.n3745 DVDD.n3728 0.00372031
R50629 DVDD.n3380 DVDD.n3368 0.00372031
R50630 DVDD.n3382 DVDD.n3350 0.00372031
R50631 DVDD.n3379 DVDD.n3367 0.00372031
R50632 DVDD.n3388 DVDD.n3369 0.00372031
R50633 DVDD.n3378 DVDD.n3366 0.00372031
R50634 DVDD.n3383 DVDD.n3352 0.00372031
R50635 DVDD.n3377 DVDD.n3365 0.00372031
R50636 DVDD.n3384 DVDD.n3353 0.00372031
R50637 DVDD.n3376 DVDD.n3364 0.00372031
R50638 DVDD.n3385 DVDD.n3354 0.00372031
R50639 DVDD.n3375 DVDD.n3363 0.00372031
R50640 DVDD.n3374 DVDD.n3362 0.00372031
R50641 DVDD.n3386 DVDD.n3356 0.00372031
R50642 DVDD.n3373 DVDD.n3361 0.00372031
R50643 DVDD.n3372 DVDD.n3360 0.00372031
R50644 DVDD.n3387 DVDD.n3358 0.00372031
R50645 DVDD.n3371 DVDD.n3359 0.00372031
R50646 DVDD.n3271 DVDD.n3259 0.00372031
R50647 DVDD.n3273 DVDD.n3237 0.00372031
R50648 DVDD.n3270 DVDD.n3258 0.00372031
R50649 DVDD.n3269 DVDD.n3257 0.00372031
R50650 DVDD.n3274 DVDD.n3239 0.00372031
R50651 DVDD.n3268 DVDD.n3256 0.00372031
R50652 DVDD.n3267 DVDD.n3255 0.00372031
R50653 DVDD.n3275 DVDD.n3241 0.00372031
R50654 DVDD.n3266 DVDD.n3254 0.00372031
R50655 DVDD.n3265 DVDD.n3253 0.00372031
R50656 DVDD.n3276 DVDD.n3243 0.00372031
R50657 DVDD.n3264 DVDD.n3252 0.00372031
R50658 DVDD.n3263 DVDD.n3251 0.00372031
R50659 DVDD.n3277 DVDD.n3245 0.00372031
R50660 DVDD.n3262 DVDD.n3250 0.00372031
R50661 DVDD.n3278 DVDD.n3249 0.00372031
R50662 DVDD.n3261 DVDD.n3247 0.00372031
R50663 DVDD.n3187 DVDD.n3150 0.00372031
R50664 DVDD.n3185 DVDD.n3173 0.00372031
R50665 DVDD.n3184 DVDD.n3172 0.00372031
R50666 DVDD.n15931 DVDD.n3152 0.00372031
R50667 DVDD.n3183 DVDD.n3171 0.00372031
R50668 DVDD.n15932 DVDD.n3153 0.00372031
R50669 DVDD.n3182 DVDD.n3170 0.00372031
R50670 DVDD.n15933 DVDD.n3154 0.00372031
R50671 DVDD.n3181 DVDD.n3169 0.00372031
R50672 DVDD.n3180 DVDD.n3168 0.00372031
R50673 DVDD.n15934 DVDD.n3156 0.00372031
R50674 DVDD.n3179 DVDD.n3167 0.00372031
R50675 DVDD.n3178 DVDD.n3166 0.00372031
R50676 DVDD.n15935 DVDD.n3158 0.00372031
R50677 DVDD.n3177 DVDD.n3165 0.00372031
R50678 DVDD.n3176 DVDD.n3164 0.00372031
R50679 DVDD.n15936 DVDD.n3160 0.00372031
R50680 DVDD.n3175 DVDD.n3163 0.00372031
R50681 DVDD.n3088 DVDD.n3060 0.00372031
R50682 DVDD.n16079 DVDD.n3102 0.00372031
R50683 DVDD.n3089 DVDD.n3061 0.00372031
R50684 DVDD.n3090 DVDD.n3062 0.00372031
R50685 DVDD.n16078 DVDD.n3100 0.00372031
R50686 DVDD.n3091 DVDD.n3063 0.00372031
R50687 DVDD.n16073 DVDD.n3092 0.00372031
R50688 DVDD.n3099 DVDD.n3071 0.00372031
R50689 DVDD.n16080 DVDD.n3073 0.00372031
R50690 DVDD.n16077 DVDD.n3098 0.00372031
R50691 DVDD.n3093 DVDD.n3065 0.00372031
R50692 DVDD.n16072 DVDD.n3058 0.00372031
R50693 DVDD.n16074 DVDD.n3094 0.00372031
R50694 DVDD.n3097 DVDD.n3069 0.00372031
R50695 DVDD.n16084 DVDD.n3074 0.00372031
R50696 DVDD.n16076 DVDD.n3096 0.00372031
R50697 DVDD.n9778 DVDD.n3067 0.00372031
R50698 DVDD.n9639 DVDD.n9638 0.00372031
R50699 DVDD.n9646 DVDD.n9629 0.00372031
R50700 DVDD.n9636 DVDD.n9635 0.00372031
R50701 DVDD.n9645 DVDD.n9627 0.00372031
R50702 DVDD.n9647 DVDD.n9634 0.00372031
R50703 DVDD.n9633 DVDD.n9631 0.00372031
R50704 DVDD.n10092 DVDD.n9640 0.00372031
R50705 DVDD.n21081 DVDD.n21060 0.00372031
R50706 DVDD.n21055 DVDD.n18754 0.00372031
R50707 DVDD.n20535 DVDD.n19797 0.00372031
R50708 DVDD.n19790 DVDD.n19788 0.00372031
R50709 DVDD.n20540 DVDD.n19767 0.00372031
R50710 DVDD.n9640 DVDD.n9631 0.00372031
R50711 DVDD.n9634 DVDD.n9633 0.00372031
R50712 DVDD.n9647 DVDD.n9630 0.00372031
R50713 DVDD.n9645 DVDD.n9636 0.00372031
R50714 DVDD.n9635 DVDD.n9629 0.00372031
R50715 DVDD.n9646 DVDD.n9637 0.00372031
R50716 DVDD.n9638 DVDD.n9628 0.00372031
R50717 DVDD.n3096 DVDD.n3067 0.00372031
R50718 DVDD.n16076 DVDD.n3066 0.00372031
R50719 DVDD.n3097 DVDD.n3074 0.00372031
R50720 DVDD.n3094 DVDD.n3069 0.00372031
R50721 DVDD.n16074 DVDD.n3070 0.00372031
R50722 DVDD.n16072 DVDD.n3093 0.00372031
R50723 DVDD.n3098 DVDD.n3065 0.00372031
R50724 DVDD.n16077 DVDD.n3064 0.00372031
R50725 DVDD.n16080 DVDD.n3099 0.00372031
R50726 DVDD.n3092 DVDD.n3071 0.00372031
R50727 DVDD.n16073 DVDD.n3072 0.00372031
R50728 DVDD.n3100 DVDD.n3063 0.00372031
R50729 DVDD.n16078 DVDD.n3090 0.00372031
R50730 DVDD.n3101 DVDD.n3062 0.00372031
R50731 DVDD.n3102 DVDD.n3061 0.00372031
R50732 DVDD.n16079 DVDD.n3088 0.00372031
R50733 DVDD.n16082 DVDD.n3060 0.00372031
R50734 DVDD.n3175 DVDD.n3160 0.00372031
R50735 DVDD.n15936 DVDD.n3164 0.00372031
R50736 DVDD.n3176 DVDD.n3159 0.00372031
R50737 DVDD.n3177 DVDD.n3158 0.00372031
R50738 DVDD.n15935 DVDD.n3166 0.00372031
R50739 DVDD.n3178 DVDD.n3157 0.00372031
R50740 DVDD.n3179 DVDD.n3156 0.00372031
R50741 DVDD.n15934 DVDD.n3168 0.00372031
R50742 DVDD.n3180 DVDD.n3155 0.00372031
R50743 DVDD.n3181 DVDD.n3154 0.00372031
R50744 DVDD.n15933 DVDD.n3170 0.00372031
R50745 DVDD.n3182 DVDD.n3153 0.00372031
R50746 DVDD.n15932 DVDD.n3171 0.00372031
R50747 DVDD.n3183 DVDD.n3152 0.00372031
R50748 DVDD.n15931 DVDD.n3172 0.00372031
R50749 DVDD.n3184 DVDD.n3151 0.00372031
R50750 DVDD.n3185 DVDD.n3150 0.00372031
R50751 DVDD.n15988 DVDD.n3187 0.00372031
R50752 DVDD.n3261 DVDD.n3249 0.00372031
R50753 DVDD.n3278 DVDD.n3246 0.00372031
R50754 DVDD.n3262 DVDD.n3245 0.00372031
R50755 DVDD.n3277 DVDD.n3251 0.00372031
R50756 DVDD.n3263 DVDD.n3244 0.00372031
R50757 DVDD.n3264 DVDD.n3243 0.00372031
R50758 DVDD.n3276 DVDD.n3253 0.00372031
R50759 DVDD.n3265 DVDD.n3242 0.00372031
R50760 DVDD.n3266 DVDD.n3241 0.00372031
R50761 DVDD.n3275 DVDD.n3255 0.00372031
R50762 DVDD.n3267 DVDD.n3240 0.00372031
R50763 DVDD.n3268 DVDD.n3239 0.00372031
R50764 DVDD.n3274 DVDD.n3257 0.00372031
R50765 DVDD.n3269 DVDD.n3238 0.00372031
R50766 DVDD.n3270 DVDD.n3237 0.00372031
R50767 DVDD.n3273 DVDD.n3259 0.00372031
R50768 DVDD.n3271 DVDD.n3236 0.00372031
R50769 DVDD.n3371 DVDD.n3358 0.00372031
R50770 DVDD.n3387 DVDD.n3360 0.00372031
R50771 DVDD.n3372 DVDD.n3357 0.00372031
R50772 DVDD.n3373 DVDD.n3356 0.00372031
R50773 DVDD.n3386 DVDD.n3362 0.00372031
R50774 DVDD.n3374 DVDD.n3355 0.00372031
R50775 DVDD.n3375 DVDD.n3354 0.00372031
R50776 DVDD.n3385 DVDD.n3364 0.00372031
R50777 DVDD.n3376 DVDD.n3353 0.00372031
R50778 DVDD.n3384 DVDD.n3365 0.00372031
R50779 DVDD.n3377 DVDD.n3352 0.00372031
R50780 DVDD.n3383 DVDD.n3366 0.00372031
R50781 DVDD.n3378 DVDD.n3351 0.00372031
R50782 DVDD.n3388 DVDD.n3367 0.00372031
R50783 DVDD.n3379 DVDD.n3350 0.00372031
R50784 DVDD.n3382 DVDD.n3368 0.00372031
R50785 DVDD.n3380 DVDD.n3349 0.00372031
R50786 DVDD.n3745 DVDD.n3726 0.00372031
R50787 DVDD.n4174 DVDD.n3784 0.00372031
R50788 DVDD.n3796 DVDD.n3782 0.00372031
R50789 DVDD.n4173 DVDD.n3785 0.00372031
R50790 DVDD.n3797 DVDD.n3781 0.00372031
R50791 DVDD.n4172 DVDD.n3786 0.00372031
R50792 DVDD.n3798 DVDD.n3780 0.00372031
R50793 DVDD.n4171 DVDD.n3787 0.00372031
R50794 DVDD.n3799 DVDD.n3779 0.00372031
R50795 DVDD.n4170 DVDD.n3788 0.00372031
R50796 DVDD.n3800 DVDD.n3778 0.00372031
R50797 DVDD.n4169 DVDD.n3789 0.00372031
R50798 DVDD.n3801 DVDD.n3777 0.00372031
R50799 DVDD.n4168 DVDD.n3790 0.00372031
R50800 DVDD.n3802 DVDD.n3776 0.00372031
R50801 DVDD.n4167 DVDD.n3791 0.00372031
R50802 DVDD.n3803 DVDD.n3775 0.00372031
R50803 DVDD.n4166 DVDD.n3792 0.00372031
R50804 DVDD.n3804 DVDD.n3774 0.00372031
R50805 DVDD.n4165 DVDD.n3793 0.00372031
R50806 DVDD.n3805 DVDD.n3773 0.00372031
R50807 DVDD.n4164 DVDD.n3794 0.00372031
R50808 DVDD.n3806 DVDD.n3772 0.00372031
R50809 DVDD.n4178 DVDD.n3795 0.00372031
R50810 DVDD.n258 DVDD.n256 0.00372031
R50811 DVDD.n271 DVDD.n262 0.00372031
R50812 DVDD.n261 DVDD.n255 0.00372031
R50813 DVDD.n270 DVDD.n264 0.00372031
R50814 DVDD.n263 DVDD.n254 0.00372031
R50815 DVDD.n269 DVDD.n266 0.00372031
R50816 DVDD.n265 DVDD.n253 0.00372031
R50817 DVDD.n22180 DVDD.n22179 0.00372031
R50818 DVDD.n267 DVDD.n252 0.00372031
R50819 DVDD.n22182 DVDD.n237 0.00372031
R50820 DVDD.n19152 DVDD.n19125 0.00372031
R50821 DVDD.n19132 DVDD.n19077 0.00372031
R50822 DVDD.n19151 DVDD.n19126 0.00372031
R50823 DVDD.n19133 DVDD.n19076 0.00372031
R50824 DVDD.n19150 DVDD.n19127 0.00372031
R50825 DVDD.n19131 DVDD.n19074 0.00372031
R50826 DVDD.n20735 DVDD.n19130 0.00372031
R50827 DVDD.n4742 DVDD.n3747 0.00372031
R50828 DVDD.n20529 DVDD.n20520 0.00372031
R50829 DVDD.n18862 DVDD.n18850 0.00372031
R50830 DVDD.n18849 DVDD.n18848 0.00372031
R50831 DVDD.n18863 DVDD.n18851 0.00372031
R50832 DVDD.n18857 DVDD.n18856 0.00372031
R50833 DVDD.n18864 DVDD.n18852 0.00372031
R50834 DVDD.n18855 DVDD.n18854 0.00372031
R50835 DVDD.n20971 DVDD.n18831 0.00372031
R50836 DVDD.n20982 DVDD.n18824 0.00372031
R50837 DVDD.n18698 DVDD.n18697 0.00372031
R50838 DVDD.n18704 DVDD.n18687 0.00372031
R50839 DVDD.n18696 DVDD.n18695 0.00372031
R50840 DVDD.n18705 DVDD.n18688 0.00372031
R50841 DVDD.n18706 DVDD.n18689 0.00372031
R50842 DVDD.n18693 DVDD.n18692 0.00372031
R50843 DVDD.n18707 DVDD.n18690 0.00372031
R50844 DVDD.n21214 DVDD.n18672 0.00372031
R50845 DVDD.n3878 DVDD.n3877 0.00372031
R50846 DVDD.n4064 DVDD.n3895 0.00372031
R50847 DVDD.n3896 DVDD.n3879 0.00372031
R50848 DVDD.n3892 DVDD.n3889 0.00372031
R50849 DVDD.n3888 DVDD.n3880 0.00372031
R50850 DVDD.n3891 DVDD.n3887 0.00372031
R50851 DVDD.n3886 DVDD.n3881 0.00372031
R50852 DVDD.n3890 DVDD.n3885 0.00372031
R50853 DVDD.n3884 DVDD.n3882 0.00372031
R50854 DVDD.n4066 DVDD.n3862 0.00372031
R50855 DVDD.n4067 DVDD.n3828 0.00372031
R50856 DVDD.n4078 DVDD.n3861 0.00372031
R50857 DVDD.n3860 DVDD.n3829 0.00372031
R50858 DVDD.n4077 DVDD.n3859 0.00372031
R50859 DVDD.n3858 DVDD.n3830 0.00372031
R50860 DVDD.n4076 DVDD.n3857 0.00372031
R50861 DVDD.n3856 DVDD.n3831 0.00372031
R50862 DVDD.n4075 DVDD.n3855 0.00372031
R50863 DVDD.n3854 DVDD.n3832 0.00372031
R50864 DVDD.n4074 DVDD.n3853 0.00372031
R50865 DVDD.n3852 DVDD.n3833 0.00372031
R50866 DVDD.n4073 DVDD.n3851 0.00372031
R50867 DVDD.n3850 DVDD.n3834 0.00372031
R50868 DVDD.n4072 DVDD.n3849 0.00372031
R50869 DVDD.n3848 DVDD.n3835 0.00372031
R50870 DVDD.n4071 DVDD.n3847 0.00372031
R50871 DVDD.n3846 DVDD.n3836 0.00372031
R50872 DVDD.n4070 DVDD.n3845 0.00372031
R50873 DVDD.n3844 DVDD.n3837 0.00372031
R50874 DVDD.n4069 DVDD.n3843 0.00372031
R50875 DVDD.n3842 DVDD.n3838 0.00372031
R50876 DVDD.n4068 DVDD.n3841 0.00372031
R50877 DVDD.n3840 DVDD.n3839 0.00372031
R50878 DVDD.n3664 DVDD.n3645 0.00372031
R50879 DVDD.n3662 DVDD.n3647 0.00372031
R50880 DVDD.n3471 DVDD.n3470 0.00372031
R50881 DVDD.n3474 DVDD.n3422 0.00372031
R50882 DVDD.n3469 DVDD.n3468 0.00372031
R50883 DVDD.n3480 DVDD.n3472 0.00372031
R50884 DVDD.n3467 DVDD.n3466 0.00372031
R50885 DVDD.n3475 DVDD.n3424 0.00372031
R50886 DVDD.n3465 DVDD.n3464 0.00372031
R50887 DVDD.n3476 DVDD.n3425 0.00372031
R50888 DVDD.n3463 DVDD.n3462 0.00372031
R50889 DVDD.n3477 DVDD.n3426 0.00372031
R50890 DVDD.n3461 DVDD.n3454 0.00372031
R50891 DVDD.n3453 DVDD.n3452 0.00372031
R50892 DVDD.n3478 DVDD.n3428 0.00372031
R50893 DVDD.n3451 DVDD.n3443 0.00372031
R50894 DVDD.n3442 DVDD.n3441 0.00372031
R50895 DVDD.n3479 DVDD.n3430 0.00372031
R50896 DVDD.n3440 DVDD.n3432 0.00372031
R50897 DVDD.n15592 DVDD.n15581 0.00372031
R50898 DVDD.n15594 DVDD.n5119 0.00372031
R50899 DVDD.n15591 DVDD.n15580 0.00372031
R50900 DVDD.n15590 DVDD.n15572 0.00372031
R50901 DVDD.n15595 DVDD.n5121 0.00372031
R50902 DVDD.n15589 DVDD.n15571 0.00372031
R50903 DVDD.n15588 DVDD.n15563 0.00372031
R50904 DVDD.n15596 DVDD.n5123 0.00372031
R50905 DVDD.n15587 DVDD.n15562 0.00372031
R50906 DVDD.n15586 DVDD.n15554 0.00372031
R50907 DVDD.n15597 DVDD.n5125 0.00372031
R50908 DVDD.n15585 DVDD.n15553 0.00372031
R50909 DVDD.n15584 DVDD.n15545 0.00372031
R50910 DVDD.n15598 DVDD.n5127 0.00372031
R50911 DVDD.n15583 DVDD.n15544 0.00372031
R50912 DVDD.n15599 DVDD.n15536 0.00372031
R50913 DVDD.n15582 DVDD.n15534 0.00372031
R50914 DVDD.n5145 DVDD.n5130 0.00372031
R50915 DVDD.n15527 DVDD.n5207 0.00372031
R50916 DVDD.n5206 DVDD.n5205 0.00372031
R50917 DVDD.n5209 DVDD.n5147 0.00372031
R50918 DVDD.n5204 DVDD.n5203 0.00372031
R50919 DVDD.n5210 DVDD.n5148 0.00372031
R50920 DVDD.n5202 DVDD.n5201 0.00372031
R50921 DVDD.n5211 DVDD.n5149 0.00372031
R50922 DVDD.n5200 DVDD.n5193 0.00372031
R50923 DVDD.n5192 DVDD.n5191 0.00372031
R50924 DVDD.n5212 DVDD.n5151 0.00372031
R50925 DVDD.n5190 DVDD.n5182 0.00372031
R50926 DVDD.n5181 DVDD.n5180 0.00372031
R50927 DVDD.n5213 DVDD.n5153 0.00372031
R50928 DVDD.n5179 DVDD.n5171 0.00372031
R50929 DVDD.n5170 DVDD.n5169 0.00372031
R50930 DVDD.n5214 DVDD.n5155 0.00372031
R50931 DVDD.n5168 DVDD.n5160 0.00372031
R50932 DVDD.n3125 DVDD.n3108 0.00372031
R50933 DVDD.n16042 DVDD.n16041 0.00372031
R50934 DVDD.n16054 DVDD.n3126 0.00372031
R50935 DVDD.n16055 DVDD.n3127 0.00372031
R50936 DVDD.n16032 DVDD.n16031 0.00372031
R50937 DVDD.n16056 DVDD.n3128 0.00372031
R50938 DVDD.n16029 DVDD.n3129 0.00372031
R50939 DVDD.n16060 DVDD.n16021 0.00372031
R50940 DVDD.n16051 DVDD.n16043 0.00372031
R50941 DVDD.n16020 DVDD.n16019 0.00372031
R50942 DVDD.n16057 DVDD.n3132 0.00372031
R50943 DVDD.n3131 DVDD.n3124 0.00372031
R50944 DVDD.n16017 DVDD.n3133 0.00372031
R50945 DVDD.n16059 DVDD.n16009 0.00372031
R50946 DVDD.n16066 DVDD.n16052 0.00372031
R50947 DVDD.n16008 DVDD.n16007 0.00372031
R50948 DVDD.n16058 DVDD.n3136 0.00372031
R50949 DVDD.n9947 DVDD.n9813 0.00372031
R50950 DVDD.n9816 DVDD.n9797 0.00372031
R50951 DVDD.n9811 DVDD.n9810 0.00372031
R50952 DVDD.n9815 DVDD.n9774 0.00372031
R50953 DVDD.n9938 DVDD.n9809 0.00372031
R50954 DVDD.n9808 DVDD.n9806 0.00372031
R50955 DVDD.n9949 DVDD.n9756 0.00372031
R50956 DVDD.n20978 DVDD.n18824 0.00372031
R50957 DVDD.n20531 DVDD.n20520 0.00372031
R50958 DVDD.n9806 DVDD.n9756 0.00372031
R50959 DVDD.n9809 DVDD.n9808 0.00372031
R50960 DVDD.n9938 DVDD.n9805 0.00372031
R50961 DVDD.n9815 DVDD.n9811 0.00372031
R50962 DVDD.n9810 DVDD.n9797 0.00372031
R50963 DVDD.n9816 DVDD.n9812 0.00372031
R50964 DVDD.n9813 DVDD.n9796 0.00372031
R50965 DVDD.n16058 DVDD.n16008 0.00372031
R50966 DVDD.n16007 DVDD.n3134 0.00372031
R50967 DVDD.n16052 DVDD.n16009 0.00372031
R50968 DVDD.n16059 DVDD.n3133 0.00372031
R50969 DVDD.n16018 DVDD.n16017 0.00372031
R50970 DVDD.n3132 DVDD.n3131 0.00372031
R50971 DVDD.n16057 DVDD.n16020 0.00372031
R50972 DVDD.n16019 DVDD.n3130 0.00372031
R50973 DVDD.n16043 DVDD.n16021 0.00372031
R50974 DVDD.n16060 DVDD.n3129 0.00372031
R50975 DVDD.n16030 DVDD.n16029 0.00372031
R50976 DVDD.n16056 DVDD.n16032 0.00372031
R50977 DVDD.n16031 DVDD.n3127 0.00372031
R50978 DVDD.n16055 DVDD.n16040 0.00372031
R50979 DVDD.n16054 DVDD.n16042 0.00372031
R50980 DVDD.n16041 DVDD.n3125 0.00372031
R50981 DVDD.n16068 DVDD.n3108 0.00372031
R50982 DVDD.n5160 DVDD.n5155 0.00372031
R50983 DVDD.n5214 DVDD.n5170 0.00372031
R50984 DVDD.n5169 DVDD.n5154 0.00372031
R50985 DVDD.n5171 DVDD.n5153 0.00372031
R50986 DVDD.n5213 DVDD.n5181 0.00372031
R50987 DVDD.n5180 DVDD.n5152 0.00372031
R50988 DVDD.n5182 DVDD.n5151 0.00372031
R50989 DVDD.n5212 DVDD.n5192 0.00372031
R50990 DVDD.n5191 DVDD.n5150 0.00372031
R50991 DVDD.n5193 DVDD.n5149 0.00372031
R50992 DVDD.n5211 DVDD.n5202 0.00372031
R50993 DVDD.n5201 DVDD.n5148 0.00372031
R50994 DVDD.n5210 DVDD.n5204 0.00372031
R50995 DVDD.n5203 DVDD.n5147 0.00372031
R50996 DVDD.n5209 DVDD.n5206 0.00372031
R50997 DVDD.n5205 DVDD.n5146 0.00372031
R50998 DVDD.n5207 DVDD.n5145 0.00372031
R50999 DVDD.n15529 DVDD.n5130 0.00372031
R51000 DVDD.n15582 DVDD.n15536 0.00372031
R51001 DVDD.n15599 DVDD.n5128 0.00372031
R51002 DVDD.n15583 DVDD.n5127 0.00372031
R51003 DVDD.n15598 DVDD.n15545 0.00372031
R51004 DVDD.n15584 DVDD.n5126 0.00372031
R51005 DVDD.n15585 DVDD.n5125 0.00372031
R51006 DVDD.n15597 DVDD.n15554 0.00372031
R51007 DVDD.n15586 DVDD.n5124 0.00372031
R51008 DVDD.n15587 DVDD.n5123 0.00372031
R51009 DVDD.n15596 DVDD.n15563 0.00372031
R51010 DVDD.n15588 DVDD.n5122 0.00372031
R51011 DVDD.n15589 DVDD.n5121 0.00372031
R51012 DVDD.n15595 DVDD.n15572 0.00372031
R51013 DVDD.n15590 DVDD.n5120 0.00372031
R51014 DVDD.n15591 DVDD.n5119 0.00372031
R51015 DVDD.n15594 DVDD.n15581 0.00372031
R51016 DVDD.n15592 DVDD.n5118 0.00372031
R51017 DVDD.n3432 DVDD.n3430 0.00372031
R51018 DVDD.n3479 DVDD.n3442 0.00372031
R51019 DVDD.n3441 DVDD.n3429 0.00372031
R51020 DVDD.n3443 DVDD.n3428 0.00372031
R51021 DVDD.n3478 DVDD.n3453 0.00372031
R51022 DVDD.n3452 DVDD.n3427 0.00372031
R51023 DVDD.n3454 DVDD.n3426 0.00372031
R51024 DVDD.n3477 DVDD.n3463 0.00372031
R51025 DVDD.n3462 DVDD.n3425 0.00372031
R51026 DVDD.n3476 DVDD.n3465 0.00372031
R51027 DVDD.n3464 DVDD.n3424 0.00372031
R51028 DVDD.n3475 DVDD.n3467 0.00372031
R51029 DVDD.n3466 DVDD.n3423 0.00372031
R51030 DVDD.n3480 DVDD.n3469 0.00372031
R51031 DVDD.n3468 DVDD.n3422 0.00372031
R51032 DVDD.n3474 DVDD.n3471 0.00372031
R51033 DVDD.n3470 DVDD.n3421 0.00372031
R51034 DVDD.n3662 DVDD.n3645 0.00372031
R51035 DVDD.n3841 DVDD.n3840 0.00372031
R51036 DVDD.n4068 DVDD.n3838 0.00372031
R51037 DVDD.n3843 DVDD.n3842 0.00372031
R51038 DVDD.n4069 DVDD.n3837 0.00372031
R51039 DVDD.n3845 DVDD.n3844 0.00372031
R51040 DVDD.n4070 DVDD.n3836 0.00372031
R51041 DVDD.n3847 DVDD.n3846 0.00372031
R51042 DVDD.n4071 DVDD.n3835 0.00372031
R51043 DVDD.n3849 DVDD.n3848 0.00372031
R51044 DVDD.n4072 DVDD.n3834 0.00372031
R51045 DVDD.n3851 DVDD.n3850 0.00372031
R51046 DVDD.n4073 DVDD.n3833 0.00372031
R51047 DVDD.n3853 DVDD.n3852 0.00372031
R51048 DVDD.n4074 DVDD.n3832 0.00372031
R51049 DVDD.n3855 DVDD.n3854 0.00372031
R51050 DVDD.n4075 DVDD.n3831 0.00372031
R51051 DVDD.n3857 DVDD.n3856 0.00372031
R51052 DVDD.n4076 DVDD.n3830 0.00372031
R51053 DVDD.n3859 DVDD.n3858 0.00372031
R51054 DVDD.n4077 DVDD.n3829 0.00372031
R51055 DVDD.n3861 DVDD.n3860 0.00372031
R51056 DVDD.n4078 DVDD.n3828 0.00372031
R51057 DVDD.n4136 DVDD.n4067 0.00372031
R51058 DVDD.n3882 DVDD.n3862 0.00372031
R51059 DVDD.n3885 DVDD.n3884 0.00372031
R51060 DVDD.n3890 DVDD.n3881 0.00372031
R51061 DVDD.n3887 DVDD.n3886 0.00372031
R51062 DVDD.n3891 DVDD.n3880 0.00372031
R51063 DVDD.n3889 DVDD.n3888 0.00372031
R51064 DVDD.n3892 DVDD.n3879 0.00372031
R51065 DVDD.n4064 DVDD.n3896 0.00372031
R51066 DVDD.n3895 DVDD.n3878 0.00372031
R51067 DVDD.n3877 DVDD.n231 0.00372031
R51068 DVDD.n18855 DVDD.n18831 0.00372031
R51069 DVDD.n18854 DVDD.n18852 0.00372031
R51070 DVDD.n18864 DVDD.n18857 0.00372031
R51071 DVDD.n18856 DVDD.n18851 0.00372031
R51072 DVDD.n18863 DVDD.n18858 0.00372031
R51073 DVDD.n18850 DVDD.n18849 0.00372031
R51074 DVDD.n18862 DVDD.n18859 0.00372031
R51075 DVDD.n4768 DVDD.n3664 0.00372031
R51076 DVDD.n18690 DVDD.n18672 0.00372031
R51077 DVDD.n18707 DVDD.n18693 0.00372031
R51078 DVDD.n18692 DVDD.n18689 0.00372031
R51079 DVDD.n18706 DVDD.n18694 0.00372031
R51080 DVDD.n18705 DVDD.n18696 0.00372031
R51081 DVDD.n18695 DVDD.n18687 0.00372031
R51082 DVDD.n18704 DVDD.n18698 0.00372031
R51083 DVDD.n18697 DVDD.n18686 0.00372031
R51084 DVDD.n21086 DVDD.n18728 0.00372031
R51085 DVDD.n21091 DVDD.n18731 0.00372031
R51086 DVDD.n21087 DVDD.n18727 0.00372031
R51087 DVDD.n21090 DVDD.n18732 0.00372031
R51088 DVDD.n21085 DVDD.n18733 0.00372031
R51089 DVDD.n21092 DVDD.n18725 0.00372031
R51090 DVDD.n21084 DVDD.n18734 0.00372031
R51091 DVDD.n21093 DVDD.n18724 0.00372031
R51092 DVDD.n117 DVDD.n94 0.00372031
R51093 DVDD.n22246 DVDD.n22245 0.00372031
R51094 DVDD.n116 DVDD.n95 0.00372031
R51095 DVDD.n115 DVDD.n96 0.00372031
R51096 DVDD.n22248 DVDD.n92 0.00372031
R51097 DVDD.n22247 DVDD.n113 0.00372031
R51098 DVDD.n22250 DVDD.n91 0.00372031
R51099 DVDD.n22249 DVDD.n90 0.00372031
R51100 DVDD.n48 DVDD.n47 0.00372031
R51101 DVDD.n68 DVDD.n51 0.00372031
R51102 DVDD.n50 DVDD.n46 0.00372031
R51103 DVDD.n67 DVDD.n52 0.00372031
R51104 DVDD.n54 DVDD.n53 0.00372031
R51105 DVDD.n69 DVDD.n44 0.00372031
R51106 DVDD.n56 DVDD.n55 0.00372031
R51107 DVDD.n70 DVDD.n43 0.00372031
R51108 DVDD.n19041 DVDD.n19032 0.00372031
R51109 DVDD.n19042 DVDD.n19031 0.00372031
R51110 DVDD.n19043 DVDD.n19030 0.00372031
R51111 DVDD.n19044 DVDD.n19029 0.00372031
R51112 DVDD.n21051 DVDD.n18796 0.00372031
R51113 DVDD.n22157 DVDD.n285 0.00372031
R51114 DVDD.n314 DVDD.n286 0.00372031
R51115 DVDD.n313 DVDD.n287 0.00372031
R51116 DVDD.n312 DVDD.n288 0.00372031
R51117 DVDD.n311 DVDD.n289 0.00372031
R51118 DVDD.n4556 DVDD.n4324 0.00372031
R51119 DVDD.n4395 DVDD.n4324 0.00372031
R51120 DVDD.n4410 DVDD.n4325 0.00372031
R51121 DVDD.n4396 DVDD.n4326 0.00372031
R51122 DVDD.n4409 DVDD.n4332 0.00372031
R51123 DVDD.n4397 DVDD.n4327 0.00372031
R51124 DVDD.n4408 DVDD.n4331 0.00372031
R51125 DVDD.n4411 DVDD.n4328 0.00372031
R51126 DVDD.n16105 DVDD.n3023 0.00372031
R51127 DVDD.n16106 DVDD.n3022 0.00372031
R51128 DVDD.n16107 DVDD.n3020 0.00372031
R51129 DVDD.n16108 DVDD.n3019 0.00372031
R51130 DVDD.n16109 DVDD.n3017 0.00372031
R51131 DVDD.n16104 DVDD.n3024 0.00372031
R51132 DVDD.n16110 DVDD.n3003 0.00372031
R51133 DVDD.n16103 DVDD.n2996 0.00372031
R51134 DVDD.n16111 DVDD.n3012 0.00372031
R51135 DVDD.n16143 DVDD.n3025 0.00372031
R51136 DVDD.n16112 DVDD.n3006 0.00372031
R51137 DVDD.n9676 DVDD.n9675 0.00372031
R51138 DVDD.n9674 DVDD.n9673 0.00372031
R51139 DVDD.n9671 DVDD.n9662 0.00372031
R51140 DVDD.n9669 DVDD.n9665 0.00372031
R51141 DVDD.n10067 DVDD.n9677 0.00372031
R51142 DVDD.n18796 DVDD.n97 0.00372031
R51143 DVDD.n9677 DVDD.n9666 0.00372031
R51144 DVDD.n9670 DVDD.n9669 0.00372031
R51145 DVDD.n9672 DVDD.n9671 0.00372031
R51146 DVDD.n9673 DVDD.n9664 0.00372031
R51147 DVDD.n9675 DVDD.n9663 0.00372031
R51148 DVDD.n16112 DVDD.n3009 0.00372031
R51149 DVDD.n3025 DVDD.n3011 0.00372031
R51150 DVDD.n16111 DVDD.n3005 0.00372031
R51151 DVDD.n16103 DVDD.n3004 0.00372031
R51152 DVDD.n16110 DVDD.n3014 0.00372031
R51153 DVDD.n16104 DVDD.n3016 0.00372031
R51154 DVDD.n16109 DVDD.n3002 0.00372031
R51155 DVDD.n16108 DVDD.n3001 0.00372031
R51156 DVDD.n16107 DVDD.n3000 0.00372031
R51157 DVDD.n16106 DVDD.n2999 0.00372031
R51158 DVDD.n16105 DVDD.n2998 0.00372031
R51159 DVDD.n4411 DVDD.n4329 0.00372031
R51160 DVDD.n4397 DVDD.n4332 0.00372031
R51161 DVDD.n4396 DVDD.n4386 0.00372031
R51162 DVDD.n4395 DVDD.n4387 0.00372031
R51163 DVDD.n309 DVDD.n289 0.00372031
R51164 DVDD.n308 DVDD.n288 0.00372031
R51165 DVDD.n307 DVDD.n287 0.00372031
R51166 DVDD.n306 DVDD.n286 0.00372031
R51167 DVDD.n305 DVDD.n285 0.00372031
R51168 DVDD.n19044 DVDD.n19027 0.00372031
R51169 DVDD.n19043 DVDD.n19026 0.00372031
R51170 DVDD.n19042 DVDD.n19025 0.00372031
R51171 DVDD.n19041 DVDD.n19023 0.00372031
R51172 DVDD.n4557 DVDD.n4556 0.00372031
R51173 DVDD.n4410 DVDD.n4387 0.00372031
R51174 DVDD.n4409 DVDD.n4326 0.00372031
R51175 DVDD.n4408 DVDD.n4327 0.00372031
R51176 DVDD.n4256 DVDD.n4247 0.00372031
R51177 DVDD.n4263 DVDD.n4256 0.00372031
R51178 DVDD.n4272 DVDD.n4255 0.00372031
R51179 DVDD.n4273 DVDD.n4254 0.00372031
R51180 DVDD.n4267 DVDD.n4254 0.00372031
R51181 DVDD.n4266 DVDD.n4253 0.00372031
R51182 DVDD.n4598 DVDD.n4253 0.00372031
R51183 DVDD.n4599 DVDD.n4598 0.00372031
R51184 DVDD.n4268 DVDD.n4267 0.00372031
R51185 DVDD.n4268 DVDD.n4266 0.00372031
R51186 DVDD.n4273 DVDD.n4265 0.00372031
R51187 DVDD.n4264 DVDD.n4263 0.00372031
R51188 DVDD.n4272 DVDD.n4264 0.00372031
R51189 DVDD.n4601 DVDD.n4247 0.00372031
R51190 DVDD.n3744 DVDD.n3725 0.00372031
R51191 DVDD.n4417 DVDD.n3725 0.00372031
R51192 DVDD.n3743 DVDD.n3724 0.00372031
R51193 DVDD.n3742 DVDD.n3723 0.00372031
R51194 DVDD.n4418 DVDD.n3723 0.00372031
R51195 DVDD.n3741 DVDD.n3722 0.00372031
R51196 DVDD.n3740 DVDD.n3722 0.00372031
R51197 DVDD.n4742 DVDD.n3740 0.00372031
R51198 DVDD.n4418 DVDD.n3732 0.00372031
R51199 DVDD.n4417 DVDD.n3730 0.00372031
R51200 DVDD.n3744 DVDD.n3729 0.00372031
R51201 DVDD.n3743 DVDD.n3730 0.00372031
R51202 DVDD.n3742 DVDD.n3731 0.00372031
R51203 DVDD.n3741 DVDD.n3732 0.00372031
R51204 DVDD.n3661 DVDD.n3644 0.00372031
R51205 DVDD.n3716 DVDD.n3644 0.00372031
R51206 DVDD.n3660 DVDD.n3643 0.00372031
R51207 DVDD.n3659 DVDD.n3642 0.00372031
R51208 DVDD.n3717 DVDD.n3642 0.00372031
R51209 DVDD.n3710 DVDD.n3641 0.00372031
R51210 DVDD.n3657 DVDD.n3641 0.00372031
R51211 DVDD.n4768 DVDD.n3657 0.00372031
R51212 DVDD.n3717 DVDD.n3651 0.00372031
R51213 DVDD.n3716 DVDD.n3649 0.00372031
R51214 DVDD.n3661 DVDD.n3648 0.00372031
R51215 DVDD.n3660 DVDD.n3649 0.00372031
R51216 DVDD.n3659 DVDD.n3650 0.00372031
R51217 DVDD.n3710 DVDD.n3651 0.00372031
R51218 DVDD.n20045 DVDD.n19738 0.00371429
R51219 DVDD.n20273 DVDD.n19941 0.00371429
R51220 DVDD.n19167 DVDD.n18845 0.00371429
R51221 DVDD.n20765 DVDD.n19051 0.00371429
R51222 DVDD.n4002 DVDD.n3874 0.00371429
R51223 DVDD.n346 DVDD.n302 0.00371429
R51224 DVDD.n9895 DVDD.n9770 0.00371429
R51225 DVDD.n9718 DVDD.n9692 0.00371429
R51226 DVDD.n18717 DVDD.n18675 0.00371429
R51227 DVDD.n21134 DVDD.n102 0.00371429
R51228 DVDD.n18070 DVDD.n18063 0.00370625
R51229 DVDD.n4108 DVDD.n4085 0.00368
R51230 DVDD.n15763 DVDD.n3487 0.00368
R51231 DVDD.n15681 DVDD.n15680 0.00368
R51232 DVDD.n15472 DVDD.n5136 0.00368
R51233 DVDD.n15390 DVDD.n3115 0.00368
R51234 DVDD.n20333 DVDD.n18943 0.00365
R51235 DVDD.n20845 DVDD.n18971 0.00365
R51236 DVDD.n22104 DVDD.n22079 0.00365
R51237 DVDD.n4575 DVDD.n4574 0.00365
R51238 DVDD.n4576 DVDD.n4282 0.00365
R51239 DVDD.n4539 DVDD.n4392 0.00365
R51240 DVDD.n10014 DVDD.n794 0.00365
R51241 DVDD.n22317 DVDD.n0 0.00365
R51242 DVDD.n5508 DVDD.n5488 0.00362632
R51243 DVDD.n828 DVDD.n812 0.00362632
R51244 DVDD.n4097 DVDD.n4081 0.00362
R51245 DVDD.n4499 DVDD.n4492 0.00362
R51246 DVDD.n15779 DVDD.n3483 0.00362
R51247 DVDD.n15863 DVDD.n2338 0.00362
R51248 DVDD.n15642 DVDD.n15602 0.00362
R51249 DVDD.n15888 DVDD.n2688 0.00362
R51250 DVDD.n5217 DVDD.n5132 0.00362
R51251 DVDD.n15968 DVDD.n2749 0.00362
R51252 DVDD.n15376 DVDD.n3111 0.00362
R51253 DVDD.n16123 DVDD.n3029 0.00362
R51254 DVDD.n19094 DVDD.n19027 0.00361707
R51255 DVDD.n19095 DVDD.n19028 0.00361707
R51256 DVDD.n19103 DVDD.n18892 0.00361707
R51257 DVDD.n19102 DVDD.n18896 0.00361707
R51258 DVDD.n19123 DVDD.n19078 0.00361707
R51259 DVDD.n19124 DVDD.n18763 0.00361707
R51260 DVDD.n20972 DVDD.n20971 0.00361707
R51261 DVDD.n20974 DVDD.n18829 0.00361707
R51262 DVDD.n18127 DVDD.n496 0.00359375
R51263 DVDD.n22223 DVDD.n22222 0.00359
R51264 DVDD.n21760 DVDD.n18395 0.00359
R51265 DVDD.n18231 DVDD.n18213 0.00359
R51266 DVDD.n18555 DVDD.n18510 0.00359
R51267 DVDD.n18528 DVDD.n18518 0.00359
R51268 DVDD.n22033 DVDD.n22032 0.00359
R51269 DVDD.n21655 DVDD.n18548 0.00359
R51270 DVDD.n21670 DVDD.n18540 0.00359
R51271 DVDD.n21989 DVDD.n226 0.00359
R51272 DVDD.n21590 DVDD.n164 0.00359
R51273 DVDD.n21749 DVDD.n18400 0.00359
R51274 DVDD.n22052 DVDD.n22051 0.00359
R51275 DVDD.n478 DVDD.n450 0.00359
R51276 DVDD.n2551 DVDD.n506 0.00359
R51277 DVDD.n16347 DVDD.n557 0.00359
R51278 DVDD.n16226 DVDD.n644 0.00359
R51279 DVDD.n2907 DVDD.n734 0.00359
R51280 DVDD.n19970 DVDD.n19958 0.00358571
R51281 DVDD.n20319 DVDD.n19835 0.00358571
R51282 DVDD.n19153 DVDD.n19073 0.00358571
R51283 DVDD.n19010 DVDD.n18881 0.00358571
R51284 DVDD.n251 DVDD.n236 0.00358571
R51285 DVDD.n427 DVDD.n426 0.00358571
R51286 DVDD.n9626 DVDD.n9613 0.00358571
R51287 DVDD.n10002 DVDD.n10001 0.00358571
R51288 DVDD.n21161 DVDD.n21088 0.00358571
R51289 DVDD.n22274 DVDD.n71 0.00358571
R51290 DVDD.n19633 DVDD.n19210 0.00357895
R51291 DVDD.n22337 DVDD.n13 0.00357895
R51292 DVDD.n5173 DVDD.n2725 0.00357317
R51293 DVDD.n16034 DVDD.n2999 0.00357317
R51294 DVDD.n16045 DVDD.n3003 0.00357317
R51295 DVDD.n5172 DVDD.n2795 0.00357317
R51296 DVDD.n16033 DVDD.n2928 0.00357317
R51297 DVDD.n16044 DVDD.n2932 0.00357317
R51298 DVDD.n5176 DVDD.n3165 0.00357317
R51299 DVDD.n16037 DVDD.n3089 0.00357317
R51300 DVDD.n16048 DVDD.n3064 0.00357317
R51301 DVDD.n5179 DVDD.n5178 0.00357317
R51302 DVDD.n16039 DVDD.n3126 0.00357317
R51303 DVDD.n16050 DVDD.n3130 0.00357317
R51304 DVDD.n4516 DVDD.n4205 0.00356
R51305 DVDD.n4660 DVDD.n4659 0.00356
R51306 DVDD.n4734 DVDD.n3760 0.00356
R51307 DVDD.n3224 DVDD.n3147 0.00356
R51308 DVDD.n15913 DVDD.n3208 0.00356
R51309 DVDD.n15912 DVDD.n15911 0.00356
R51310 DVDD.n15820 DVDD.n3231 0.00356
R51311 DVDD.n16390 DVDD.n16381 0.00356
R51312 DVDD.n16368 DVDD.n16367 0.00356
R51313 DVDD.n16267 DVDD.n2644 0.00356
R51314 DVDD.n16315 DVDD.n16314 0.00356
R51315 DVDD.n2772 DVDD.n2746 0.00356
R51316 DVDD.n16246 DVDD.n16245 0.00356
R51317 DVDD.n16141 DVDD.n2995 0.00356
R51318 DVDD.n16184 DVDD.n2920 0.00356
R51319 DVDD.n4770 DVDD.n3640 0.0035375
R51320 DVDD.n5023 DVDD.n4889 0.00353158
R51321 DVDD.n15751 DVDD.n4893 0.00353158
R51322 DVDD.n5270 DVDD.n5063 0.00353158
R51323 DVDD.n5285 DVDD.n5059 0.00353158
R51324 DVDD.n5317 DVDD.n5242 0.00353158
R51325 DVDD.n5363 DVDD.n5231 0.00353158
R51326 DVDD.n5429 DVDD.n5399 0.00353158
R51327 DVDD.n5444 DVDD.n5403 0.00353158
R51328 DVDD.n18002 DVDD.n525 0.00353158
R51329 DVDD.n17987 DVDD.n529 0.00353158
R51330 DVDD.n602 DVDD.n575 0.00353158
R51331 DVDD.n617 DVDD.n572 0.00353158
R51332 DVDD.n17965 DVDD.n17964 0.00353158
R51333 DVDD.n725 DVDD.n669 0.00353158
R51334 DVDD.n17935 DVDD.n751 0.00353158
R51335 DVDD.n17920 DVDD.n755 0.00353158
R51336 DVDD.n20284 DVDD.n19935 0.00352927
R51337 DVDD.n19932 DVDD.n19874 0.00352927
R51338 DVDD.n19930 DVDD.n19883 0.00352927
R51339 DVDD.n19928 DVDD.n19875 0.00352927
R51340 DVDD.n19926 DVDD.n19882 0.00352927
R51341 DVDD.n19924 DVDD.n19876 0.00352927
R51342 DVDD.n19922 DVDD.n19881 0.00352927
R51343 DVDD.n19920 DVDD.n19877 0.00352927
R51344 DVDD.n19918 DVDD.n19880 0.00352927
R51345 DVDD.n19916 DVDD.n19878 0.00352927
R51346 DVDD.n19914 DVDD.n19879 0.00352927
R51347 DVDD.n20422 DVDD.n19832 0.00352927
R51348 DVDD.n20421 DVDD.n19842 0.00352927
R51349 DVDD.n20419 DVDD.n20418 0.00352927
R51350 DVDD.n20415 DVDD.n19851 0.00352927
R51351 DVDD.n20412 DVDD.n20377 0.00352927
R51352 DVDD.n20410 DVDD.n19852 0.00352927
R51353 DVDD.n20407 DVDD.n20376 0.00352927
R51354 DVDD.n20405 DVDD.n19853 0.00352927
R51355 DVDD.n20402 DVDD.n20375 0.00352927
R51356 DVDD.n20400 DVDD.n19854 0.00352927
R51357 DVDD.n20397 DVDD.n20374 0.00352927
R51358 DVDD.n20243 DVDD.n20022 0.00352927
R51359 DVDD.n20019 DVDD.n19959 0.00352927
R51360 DVDD.n20017 DVDD.n19968 0.00352927
R51361 DVDD.n20015 DVDD.n19960 0.00352927
R51362 DVDD.n20013 DVDD.n19967 0.00352927
R51363 DVDD.n20011 DVDD.n19961 0.00352927
R51364 DVDD.n20009 DVDD.n19966 0.00352927
R51365 DVDD.n20007 DVDD.n19962 0.00352927
R51366 DVDD.n20005 DVDD.n19965 0.00352927
R51367 DVDD.n20003 DVDD.n19963 0.00352927
R51368 DVDD.n20001 DVDD.n19964 0.00352927
R51369 DVDD.n20577 DVDD.n19721 0.00352927
R51370 DVDD.n20574 DVDD.n19722 0.00352927
R51371 DVDD.n20573 DVDD.n19732 0.00352927
R51372 DVDD.n19751 DVDD.n19741 0.00352927
R51373 DVDD.n20571 DVDD.n20570 0.00352927
R51374 DVDD.n20567 DVDD.n19742 0.00352927
R51375 DVDD.n20564 DVDD.n19750 0.00352927
R51376 DVDD.n20562 DVDD.n19743 0.00352927
R51377 DVDD.n20559 DVDD.n19749 0.00352927
R51378 DVDD.n20557 DVDD.n19744 0.00352927
R51379 DVDD.n20554 DVDD.n19748 0.00352927
R51380 DVDD.n20163 DVDD.n20162 0.00352143
R51381 DVDD.n20655 DVDD.n20654 0.00352143
R51382 DVDD.n3927 DVDD.n3926 0.00352143
R51383 DVDD.n9860 DVDD.n5478 0.00352143
R51384 DVDD.n19696 DVDD.n19200 0.00352143
R51385 DVDD.n4161 DVDD.n3766 0.0035
R51386 DVDD.n4639 DVDD.n4220 0.0035
R51387 DVDD.n15828 DVDD.n3402 0.0035
R51388 DVDD.n2505 DVDD.n2479 0.0035
R51389 DVDD.n3299 DVDD.n3291 0.0035
R51390 DVDD.n2632 DVDD.n2625 0.0035
R51391 DVDD.n3205 DVDD.n3198 0.0035
R51392 DVDD.n2857 DVDD.n2827 0.0035
R51393 DVDD.n3215 DVDD.n3086 0.0035
R51394 DVDD.n16170 DVDD.n2968 0.0035
R51395 DVDD.n21940 DVDD.n21781 0.00347759
R51396 DVDD.n18479 DVDD.n18478 0.00347759
R51397 DVDD.n21797 DVDD.n21796 0.00347759
R51398 DVDD.n18102 DVDD.n18101 0.00347759
R51399 DVDD.n17726 DVDD.n893 0.00347744
R51400 DVDD.n3586 DVDD.n3554 0.00347
R51401 DVDD.n15736 DVDD.n4901 0.00347
R51402 DVDD.n5100 DVDD.n5043 0.00347
R51403 DVDD.n15445 DVDD.n5257 0.00347
R51404 DVDD.n15338 DVDD.n5372 0.00347
R51405 DVDD.n20225 DVDD.n19974 0.00345714
R51406 DVDD.n20303 DVDD.n19839 0.00345714
R51407 DVDD.n20717 DVDD.n19137 0.00345714
R51408 DVDD.n20794 DVDD.n18885 0.00345714
R51409 DVDD.n4022 DVDD.n240 0.00345714
R51410 DVDD.n406 DVDD.n377 0.00345714
R51411 DVDD.n9913 DVDD.n9617 0.00345714
R51412 DVDD.n9982 DVDD.n9754 0.00345714
R51413 DVDD.n21175 DVDD.n21097 0.00345714
R51414 DVDD.n22288 DVDD.n76 0.00345714
R51415 DVDD.n3818 DVDD.n3814 0.00344
R51416 DVDD.n15809 DVDD.n3397 0.00344
R51417 DVDD.n15667 DVDD.n3287 0.00344
R51418 DVDD.n15507 DVDD.n3194 0.00344
R51419 DVDD.n15996 DVDD.n3082 0.00344
R51420 DVDD.n5468 DVDD.n5466 0.00343684
R51421 DVDD.n17879 DVDD.n17878 0.00343684
R51422 DVDD.n21845 DVDD.n21842 0.003425
R51423 DVDD.n21974 DVDD.n21973 0.003425
R51424 DVDD.n21236 DVDD.n21235 0.003425
R51425 DVDD.n18292 DVDD.n18287 0.003425
R51426 DVDD.n21827 DVDD.n21826 0.003425
R51427 DVDD.n18475 DVDD.n18474 0.003425
R51428 DVDD.n3652 DVDD.n3646 0.003425
R51429 DVDD.n4304 DVDD.n4269 0.003425
R51430 DVDD.n3695 DVDD.n3655 0.003425
R51431 DVDD.n4554 DVDD.n4389 0.003425
R51432 DVDD.n3580 DVDD.n3563 0.00341
R51433 DVDD.n15744 DVDD.n15712 0.00341
R51434 DVDD.n5091 DVDD.n5052 0.00341
R51435 DVDD.n15453 DVDD.n15421 0.00341
R51436 DVDD.n15329 DVDD.n5378 0.00341
R51437 DVDD.n10695 DVDD.n10240 0.00339933
R51438 DVDD.n17273 DVDD.n1265 0.00339933
R51439 DVDD.n10696 DVDD.n10239 0.00339933
R51440 DVDD.n17274 DVDD.n1266 0.00339933
R51441 DVDD.n20145 DVDD.n20125 0.00339286
R51442 DVDD.n20632 DVDD.n20612 0.00339286
R51443 DVDD.n3960 DVDD.n3932 0.00339286
R51444 DVDD.n9844 DVDD.n5483 0.00339286
R51445 DVDD.n19655 DVDD.n19196 0.00339286
R51446 DVDD.n3810 DVDD.n3761 0.00338
R51447 DVDD.n4630 DVDD.n4215 0.00338
R51448 DVDD.n15819 DVDD.n3392 0.00338
R51449 DVDD.n2496 DVDD.n2436 0.00338
R51450 DVDD.n15910 DVDD.n15909 0.00338
R51451 DVDD.n2635 DVDD.n2617 0.00338
R51452 DVDD.n3190 DVDD.n3162 0.00338
R51453 DVDD.n2848 DVDD.n2821 0.00338
R51454 DVDD.n3223 DVDD.n3077 0.00338
R51455 DVDD.n16161 DVDD.n2960 0.00338
R51456 DVDD.n2283 DVDD.n2279 0.00336948
R51457 DVDD.n2281 DVDD.n2280 0.00336948
R51458 DVDD.n2270 DVDD.n2267 0.00336948
R51459 DVDD.n16451 DVDD.n2256 0.00336948
R51460 DVDD.n8963 DVDD.n8960 0.00336948
R51461 DVDD.n10222 DVDD.n8950 0.00336948
R51462 DVDD.n8960 DVDD.n8950 0.00336948
R51463 DVDD.n2280 DVDD.n2279 0.00336948
R51464 DVDD.n2267 DVDD.n2256 0.00336948
R51465 DVDD.n10219 DVDD.n8963 0.00336948
R51466 DVDD.n16431 DVDD.n2283 0.00336948
R51467 DVDD.n16449 DVDD.n2270 0.00336948
R51468 DVDD.n10168 DVDD.n8972 0.00336948
R51469 DVDD.n9572 DVDD.n8973 0.00336948
R51470 DVDD.n8973 DVDD.n8972 0.00336948
R51471 DVDD.n10202 DVDD.n10168 0.00336948
R51472 DVDD.n18059 DVDD.n502 0.00336875
R51473 DVDD.n19503 DVDD.n114 0.00335366
R51474 DVDD.n19288 DVDD.n45 0.00335366
R51475 DVDD.n19553 DVDD.n18726 0.00335366
R51476 DVDD.n19235 DVDD.n18688 0.00335366
R51477 DVDD.n3591 DVDD.n3559 0.00335
R51478 DVDD.n15730 DVDD.n15707 0.00335
R51479 DVDD.n15694 DVDD.n5049 0.00335
R51480 DVDD.n15439 DVDD.n15416 0.00335
R51481 DVDD.n15402 DVDD.n5381 0.00335
R51482 DVDD.n5023 DVDD.n3514 0.00334211
R51483 DVDD.n4893 DVDD.n3511 0.00334211
R51484 DVDD.n5270 DVDD.n5068 0.00334211
R51485 DVDD.n5285 DVDD.n5071 0.00334211
R51486 DVDD.n5317 DVDD.n5241 0.00334211
R51487 DVDD.n5363 DVDD.n5252 0.00334211
R51488 DVDD.n5429 DVDD.n5389 0.00334211
R51489 DVDD.n5444 DVDD.n5386 0.00334211
R51490 DVDD.n18002 DVDD.n535 0.00334211
R51491 DVDD.n17987 DVDD.n532 0.00334211
R51492 DVDD.n602 DVDD.n590 0.00334211
R51493 DVDD.n617 DVDD.n577 0.00334211
R51494 DVDD.n17965 DVDD.n639 0.00334211
R51495 DVDD.n725 DVDD.n680 0.00334211
R51496 DVDD.n17935 DVDD.n768 0.00334211
R51497 DVDD.n17920 DVDD.n765 0.00334211
R51498 DVDD.n21251 DVDD.n21250 0.00334
R51499 DVDD.n21250 DVDD.n18507 0.00334
R51500 DVDD.n21720 DVDD.n18508 0.00334
R51501 DVDD.n21716 DVDD.n18508 0.00334
R51502 DVDD.n21716 DVDD.n21715 0.00334
R51503 DVDD.n21715 DVDD.n21714 0.00334
R51504 DVDD.n21710 DVDD.n18512 0.00334
R51505 DVDD.n21710 DVDD.n21709 0.00334
R51506 DVDD.n21709 DVDD.n21708 0.00334
R51507 DVDD.n21708 DVDD.n18517 0.00334
R51508 DVDD.n22207 DVDD.n22206 0.00334
R51509 DVDD.n22206 DVDD.n22205 0.00334
R51510 DVDD.n22205 DVDD.n197 0.00334
R51511 DVDD.n22201 DVDD.n197 0.00334
R51512 DVDD.n22200 DVDD.n22199 0.00334
R51513 DVDD.n22199 DVDD.n202 0.00334
R51514 DVDD.n22195 DVDD.n202 0.00334
R51515 DVDD.n22195 DVDD.n22194 0.00334
R51516 DVDD.n22029 DVDD.n219 0.00334
R51517 DVDD.n22030 DVDD.n22029 0.00334
R51518 DVDD.n21230 DVDD.n21229 0.00334
R51519 DVDD.n21229 DVDD.n18505 0.00334
R51520 DVDD.n18545 DVDD.n18504 0.00334
R51521 DVDD.n21657 DVDD.n18545 0.00334
R51522 DVDD.n21658 DVDD.n21657 0.00334
R51523 DVDD.n21659 DVDD.n21658 0.00334
R51524 DVDD.n21664 DVDD.n18542 0.00334
R51525 DVDD.n21665 DVDD.n21664 0.00334
R51526 DVDD.n21667 DVDD.n21665 0.00334
R51527 DVDD.n21667 DVDD.n21666 0.00334
R51528 DVDD.n18321 DVDD.n18320 0.00334
R51529 DVDD.n18326 DVDD.n18321 0.00334
R51530 DVDD.n18327 DVDD.n18326 0.00334
R51531 DVDD.n18360 DVDD.n18327 0.00334
R51532 DVDD.n18359 DVDD.n18358 0.00334
R51533 DVDD.n18358 DVDD.n18328 0.00334
R51534 DVDD.n18354 DVDD.n18328 0.00334
R51535 DVDD.n18354 DVDD.n221 0.00334
R51536 DVDD.n22192 DVDD.n222 0.00334
R51537 DVDD.n22188 DVDD.n222 0.00334
R51538 DVDD.n18455 DVDD.n18453 0.00334
R51539 DVDD.n18502 DVDD.n18453 0.00334
R51540 DVDD.n18452 DVDD.n169 0.00334
R51541 DVDD.n22220 DVDD.n169 0.00334
R51542 DVDD.n22220 DVDD.n22219 0.00334
R51543 DVDD.n22219 DVDD.n22218 0.00334
R51544 DVDD.n22214 DVDD.n170 0.00334
R51545 DVDD.n22214 DVDD.n22213 0.00334
R51546 DVDD.n22213 DVDD.n22212 0.00334
R51547 DVDD.n22212 DVDD.n175 0.00334
R51548 DVDD.n21882 DVDD.n21837 0.00334
R51549 DVDD.n21883 DVDD.n21882 0.00334
R51550 DVDD.n21884 DVDD.n21883 0.00334
R51551 DVDD.n21884 DVDD.n21834 0.00334
R51552 DVDD.n21891 DVDD.n21890 0.00334
R51553 DVDD.n21893 DVDD.n21891 0.00334
R51554 DVDD.n21893 DVDD.n21892 0.00334
R51555 DVDD.n21892 DVDD.n214 0.00334
R51556 DVDD.n18237 DVDD.n215 0.00334
R51557 DVDD.n18237 DVDD.n18236 0.00334
R51558 DVDD.n18488 DVDD.n18487 0.00334
R51559 DVDD.n18488 DVDD.n18450 0.00334
R51560 DVDD.n21587 DVDD.n18449 0.00334
R51561 DVDD.n21588 DVDD.n21587 0.00334
R51562 DVDD.n21588 DVDD.n18406 0.00334
R51563 DVDD.n21742 DVDD.n18406 0.00334
R51564 DVDD.n21744 DVDD.n21743 0.00334
R51565 DVDD.n21745 DVDD.n21744 0.00334
R51566 DVDD.n21747 DVDD.n21745 0.00334
R51567 DVDD.n21747 DVDD.n21746 0.00334
R51568 DVDD.n21869 DVDD.n21862 0.00334
R51569 DVDD.n21870 DVDD.n21869 0.00334
R51570 DVDD.n21871 DVDD.n21870 0.00334
R51571 DVDD.n21871 DVDD.n21806 0.00334
R51572 DVDD.n21906 DVDD.n21905 0.00334
R51573 DVDD.n21907 DVDD.n21906 0.00334
R51574 DVDD.n21908 DVDD.n21907 0.00334
R51575 DVDD.n21908 DVDD.n211 0.00334
R51576 DVDD.n18222 DVDD.n210 0.00334
R51577 DVDD.n22054 DVDD.n18222 0.00334
R51578 DVDD.n4800 DVDD.n4799 0.00334
R51579 DVDD.n4799 DVDD.n4798 0.00334
R51580 DVDD.n4798 DVDD.n3582 0.00334
R51581 DVDD.n4794 DVDD.n3582 0.00334
R51582 DVDD.n4794 DVDD.n4793 0.00334
R51583 DVDD.n4793 DVDD.n4792 0.00334
R51584 DVDD.n4792 DVDD.n3588 0.00334
R51585 DVDD.n4788 DVDD.n3588 0.00334
R51586 DVDD.n4788 DVDD.n4787 0.00334
R51587 DVDD.n4787 DVDD.n4786 0.00334
R51588 DVDD.n4786 DVDD.n3594 0.00334
R51589 DVDD.n4782 DVDD.n3594 0.00334
R51590 DVDD.n4103 DVDD.n3599 0.00334
R51591 DVDD.n4103 DVDD.n4102 0.00334
R51592 DVDD.n4112 DVDD.n4102 0.00334
R51593 DVDD.n4113 DVDD.n4112 0.00334
R51594 DVDD.n4114 DVDD.n4113 0.00334
R51595 DVDD.n4114 DVDD.n4098 0.00334
R51596 DVDD.n4120 DVDD.n4098 0.00334
R51597 DVDD.n4121 DVDD.n4120 0.00334
R51598 DVDD.n4122 DVDD.n4121 0.00334
R51599 DVDD.n4122 DVDD.n4094 0.00334
R51600 DVDD.n4128 DVDD.n4094 0.00334
R51601 DVDD.n4129 DVDD.n4128 0.00334
R51602 DVDD.n4130 DVDD.n4129 0.00334
R51603 DVDD.n4130 DVDD.n3825 0.00334
R51604 DVDD.n4140 DVDD.n3825 0.00334
R51605 DVDD.n4141 DVDD.n4140 0.00334
R51606 DVDD.n4143 DVDD.n4141 0.00334
R51607 DVDD.n4143 DVDD.n4142 0.00334
R51608 DVDD.n4142 DVDD.n3821 0.00334
R51609 DVDD.n4151 DVDD.n3821 0.00334
R51610 DVDD.n4152 DVDD.n4151 0.00334
R51611 DVDD.n4153 DVDD.n4152 0.00334
R51612 DVDD.n4153 DVDD.n3758 0.00334
R51613 DVDD.n4735 DVDD.n3759 0.00334
R51614 DVDD.n4731 DVDD.n3759 0.00334
R51615 DVDD.n4731 DVDD.n4730 0.00334
R51616 DVDD.n4730 DVDD.n4729 0.00334
R51617 DVDD.n4729 DVDD.n3765 0.00334
R51618 DVDD.n4725 DVDD.n3765 0.00334
R51619 DVDD.n4725 DVDD.n4724 0.00334
R51620 DVDD.n4724 DVDD.n4723 0.00334
R51621 DVDD.n4723 DVDD.n3770 0.00334
R51622 DVDD.n4719 DVDD.n3770 0.00334
R51623 DVDD.n4719 DVDD.n4718 0.00334
R51624 DVDD.n4718 DVDD.n4717 0.00334
R51625 DVDD.n4717 DVDD.n4183 0.00334
R51626 DVDD.n4713 DVDD.n4183 0.00334
R51627 DVDD.n4713 DVDD.n4712 0.00334
R51628 DVDD.n4712 DVDD.n4711 0.00334
R51629 DVDD.n4711 DVDD.n4189 0.00334
R51630 DVDD.n4707 DVDD.n4189 0.00334
R51631 DVDD.n4707 DVDD.n4706 0.00334
R51632 DVDD.n4706 DVDD.n4705 0.00334
R51633 DVDD.n4705 DVDD.n4194 0.00334
R51634 DVDD.n4701 DVDD.n4194 0.00334
R51635 DVDD.n4701 DVDD.n4700 0.00334
R51636 DVDD.n4698 DVDD.n4201 0.00334
R51637 DVDD.n4694 DVDD.n4201 0.00334
R51638 DVDD.n4694 DVDD.n4693 0.00334
R51639 DVDD.n4693 DVDD.n4692 0.00334
R51640 DVDD.n4692 DVDD.n4207 0.00334
R51641 DVDD.n4688 DVDD.n4207 0.00334
R51642 DVDD.n4688 DVDD.n4687 0.00334
R51643 DVDD.n4687 DVDD.n4686 0.00334
R51644 DVDD.n4686 DVDD.n4212 0.00334
R51645 DVDD.n4682 DVDD.n4212 0.00334
R51646 DVDD.n4682 DVDD.n4681 0.00334
R51647 DVDD.n4681 DVDD.n4680 0.00334
R51648 DVDD.n4680 DVDD.n4217 0.00334
R51649 DVDD.n4676 DVDD.n4217 0.00334
R51650 DVDD.n4676 DVDD.n4675 0.00334
R51651 DVDD.n4675 DVDD.n4674 0.00334
R51652 DVDD.n4674 DVDD.n4222 0.00334
R51653 DVDD.n4670 DVDD.n4222 0.00334
R51654 DVDD.n4670 DVDD.n4669 0.00334
R51655 DVDD.n4669 DVDD.n4668 0.00334
R51656 DVDD.n4668 DVDD.n4227 0.00334
R51657 DVDD.n4664 DVDD.n4227 0.00334
R51658 DVDD.n4664 DVDD.n4663 0.00334
R51659 DVDD.n492 DVDD.n485 0.00334
R51660 DVDD.n18140 DVDD.n485 0.00334
R51661 DVDD.n18141 DVDD.n18140 0.00334
R51662 DVDD.n18142 DVDD.n18141 0.00334
R51663 DVDD.n18142 DVDD.n481 0.00334
R51664 DVDD.n18148 DVDD.n481 0.00334
R51665 DVDD.n18149 DVDD.n18148 0.00334
R51666 DVDD.n18150 DVDD.n18149 0.00334
R51667 DVDD.n18150 DVDD.n477 0.00334
R51668 DVDD.n18156 DVDD.n477 0.00334
R51669 DVDD.n15717 DVDD.n15716 0.00334
R51670 DVDD.n15718 DVDD.n15717 0.00334
R51671 DVDD.n15719 DVDD.n15718 0.00334
R51672 DVDD.n15720 DVDD.n15719 0.00334
R51673 DVDD.n15721 DVDD.n15720 0.00334
R51674 DVDD.n15722 DVDD.n15721 0.00334
R51675 DVDD.n15723 DVDD.n15722 0.00334
R51676 DVDD.n15724 DVDD.n15723 0.00334
R51677 DVDD.n15725 DVDD.n15724 0.00334
R51678 DVDD.n15726 DVDD.n15725 0.00334
R51679 DVDD.n15726 DVDD.n3508 0.00334
R51680 DVDD.n15756 DVDD.n3508 0.00334
R51681 DVDD.n15759 DVDD.n15758 0.00334
R51682 DVDD.n15758 DVDD.n3503 0.00334
R51683 DVDD.n15767 DVDD.n3503 0.00334
R51684 DVDD.n15768 DVDD.n15767 0.00334
R51685 DVDD.n15769 DVDD.n15768 0.00334
R51686 DVDD.n15769 DVDD.n3500 0.00334
R51687 DVDD.n15776 DVDD.n3500 0.00334
R51688 DVDD.n15777 DVDD.n15776 0.00334
R51689 DVDD.n15778 DVDD.n15777 0.00334
R51690 DVDD.n15778 DVDD.n3497 0.00334
R51691 DVDD.n15785 DVDD.n3497 0.00334
R51692 DVDD.n15786 DVDD.n15785 0.00334
R51693 DVDD.n15787 DVDD.n15786 0.00334
R51694 DVDD.n15787 DVDD.n3417 0.00334
R51695 DVDD.n15798 DVDD.n3417 0.00334
R51696 DVDD.n15799 DVDD.n15798 0.00334
R51697 DVDD.n15800 DVDD.n15799 0.00334
R51698 DVDD.n15800 DVDD.n3413 0.00334
R51699 DVDD.n15806 DVDD.n3413 0.00334
R51700 DVDD.n15807 DVDD.n15806 0.00334
R51701 DVDD.n15808 DVDD.n15807 0.00334
R51702 DVDD.n15808 DVDD.n3410 0.00334
R51703 DVDD.n15816 DVDD.n3410 0.00334
R51704 DVDD.n15823 DVDD.n15818 0.00334
R51705 DVDD.n15824 DVDD.n15823 0.00334
R51706 DVDD.n15825 DVDD.n15824 0.00334
R51707 DVDD.n15825 DVDD.n3407 0.00334
R51708 DVDD.n15832 DVDD.n3407 0.00334
R51709 DVDD.n15833 DVDD.n15832 0.00334
R51710 DVDD.n15834 DVDD.n15833 0.00334
R51711 DVDD.n15834 DVDD.n3345 0.00334
R51712 DVDD.n15842 DVDD.n3345 0.00334
R51713 DVDD.n15843 DVDD.n15842 0.00334
R51714 DVDD.n15844 DVDD.n15843 0.00334
R51715 DVDD.n15844 DVDD.n3341 0.00334
R51716 DVDD.n15851 DVDD.n3341 0.00334
R51717 DVDD.n15852 DVDD.n15851 0.00334
R51718 DVDD.n15853 DVDD.n15852 0.00334
R51719 DVDD.n15853 DVDD.n3339 0.00334
R51720 DVDD.n15860 DVDD.n3339 0.00334
R51721 DVDD.n15861 DVDD.n15860 0.00334
R51722 DVDD.n15862 DVDD.n15861 0.00334
R51723 DVDD.n15862 DVDD.n3336 0.00334
R51724 DVDD.n15869 DVDD.n3336 0.00334
R51725 DVDD.n15870 DVDD.n15869 0.00334
R51726 DVDD.n15871 DVDD.n15870 0.00334
R51727 DVDD.n15875 DVDD.n15874 0.00334
R51728 DVDD.n15874 DVDD.n2380 0.00334
R51729 DVDD.n2381 DVDD.n2380 0.00334
R51730 DVDD.n2382 DVDD.n2381 0.00334
R51731 DVDD.n2383 DVDD.n2382 0.00334
R51732 DVDD.n2386 DVDD.n2383 0.00334
R51733 DVDD.n2387 DVDD.n2386 0.00334
R51734 DVDD.n2388 DVDD.n2387 0.00334
R51735 DVDD.n2494 DVDD.n2388 0.00334
R51736 DVDD.n2495 DVDD.n2494 0.00334
R51737 DVDD.n2500 DVDD.n2495 0.00334
R51738 DVDD.n2501 DVDD.n2500 0.00334
R51739 DVDD.n2502 DVDD.n2501 0.00334
R51740 DVDD.n2502 DVDD.n2491 0.00334
R51741 DVDD.n2509 DVDD.n2491 0.00334
R51742 DVDD.n2510 DVDD.n2509 0.00334
R51743 DVDD.n2511 DVDD.n2510 0.00334
R51744 DVDD.n2511 DVDD.n2488 0.00334
R51745 DVDD.n2518 DVDD.n2488 0.00334
R51746 DVDD.n2519 DVDD.n2518 0.00334
R51747 DVDD.n2520 DVDD.n2519 0.00334
R51748 DVDD.n2521 DVDD.n2520 0.00334
R51749 DVDD.n2522 DVDD.n2521 0.00334
R51750 DVDD.n2566 DVDD.n2528 0.00334
R51751 DVDD.n2529 DVDD.n2528 0.00334
R51752 DVDD.n2530 DVDD.n2529 0.00334
R51753 DVDD.n2531 DVDD.n2530 0.00334
R51754 DVDD.n2532 DVDD.n2531 0.00334
R51755 DVDD.n2533 DVDD.n2532 0.00334
R51756 DVDD.n2534 DVDD.n2533 0.00334
R51757 DVDD.n2535 DVDD.n2534 0.00334
R51758 DVDD.n2536 DVDD.n2535 0.00334
R51759 DVDD.n2537 DVDD.n2536 0.00334
R51760 DVDD.n5093 DVDD.n5087 0.00334
R51761 DVDD.n5094 DVDD.n5093 0.00334
R51762 DVDD.n5095 DVDD.n5094 0.00334
R51763 DVDD.n5095 DVDD.n5084 0.00334
R51764 DVDD.n5102 DVDD.n5084 0.00334
R51765 DVDD.n5103 DVDD.n5102 0.00334
R51766 DVDD.n5104 DVDD.n5103 0.00334
R51767 DVDD.n5105 DVDD.n5104 0.00334
R51768 DVDD.n5106 DVDD.n5105 0.00334
R51769 DVDD.n5107 DVDD.n5106 0.00334
R51770 DVDD.n5108 DVDD.n5107 0.00334
R51771 DVDD.n5109 DVDD.n5108 0.00334
R51772 DVDD.n5115 DVDD.n5114 0.00334
R51773 DVDD.n5116 DVDD.n5115 0.00334
R51774 DVDD.n15629 DVDD.n5116 0.00334
R51775 DVDD.n15630 DVDD.n15629 0.00334
R51776 DVDD.n15630 DVDD.n15628 0.00334
R51777 DVDD.n15637 DVDD.n15628 0.00334
R51778 DVDD.n15638 DVDD.n15637 0.00334
R51779 DVDD.n15639 DVDD.n15638 0.00334
R51780 DVDD.n15639 DVDD.n15625 0.00334
R51781 DVDD.n15646 DVDD.n15625 0.00334
R51782 DVDD.n15647 DVDD.n15646 0.00334
R51783 DVDD.n15648 DVDD.n15647 0.00334
R51784 DVDD.n15648 DVDD.n15622 0.00334
R51785 DVDD.n15655 DVDD.n15622 0.00334
R51786 DVDD.n15656 DVDD.n15655 0.00334
R51787 DVDD.n15657 DVDD.n15656 0.00334
R51788 DVDD.n15658 DVDD.n15657 0.00334
R51789 DVDD.n15659 DVDD.n15658 0.00334
R51790 DVDD.n15660 DVDD.n15659 0.00334
R51791 DVDD.n15661 DVDD.n15660 0.00334
R51792 DVDD.n15662 DVDD.n15661 0.00334
R51793 DVDD.n15664 DVDD.n15662 0.00334
R51794 DVDD.n15664 DVDD.n15663 0.00334
R51795 DVDD.n3301 DVDD.n3233 0.00334
R51796 DVDD.n3302 DVDD.n3301 0.00334
R51797 DVDD.n3307 DVDD.n3302 0.00334
R51798 DVDD.n3308 DVDD.n3307 0.00334
R51799 DVDD.n3309 DVDD.n3308 0.00334
R51800 DVDD.n3309 DVDD.n3298 0.00334
R51801 DVDD.n3316 DVDD.n3298 0.00334
R51802 DVDD.n3317 DVDD.n3316 0.00334
R51803 DVDD.n3318 DVDD.n3317 0.00334
R51804 DVDD.n3319 DVDD.n3318 0.00334
R51805 DVDD.n3320 DVDD.n3319 0.00334
R51806 DVDD.n3323 DVDD.n3320 0.00334
R51807 DVDD.n3324 DVDD.n3323 0.00334
R51808 DVDD.n3325 DVDD.n3324 0.00334
R51809 DVDD.n3326 DVDD.n3325 0.00334
R51810 DVDD.n3327 DVDD.n3326 0.00334
R51811 DVDD.n3328 DVDD.n3327 0.00334
R51812 DVDD.n3329 DVDD.n3328 0.00334
R51813 DVDD.n3330 DVDD.n3329 0.00334
R51814 DVDD.n3331 DVDD.n3330 0.00334
R51815 DVDD.n3332 DVDD.n3331 0.00334
R51816 DVDD.n3333 DVDD.n3332 0.00334
R51817 DVDD.n3333 DVDD.n2704 0.00334
R51818 DVDD.n16264 DVDD.n16263 0.00334
R51819 DVDD.n16264 DVDD.n2642 0.00334
R51820 DVDD.n16273 DVDD.n2642 0.00334
R51821 DVDD.n16274 DVDD.n16273 0.00334
R51822 DVDD.n16276 DVDD.n16274 0.00334
R51823 DVDD.n16276 DVDD.n16275 0.00334
R51824 DVDD.n16275 DVDD.n2639 0.00334
R51825 DVDD.n2639 DVDD.n2637 0.00334
R51826 DVDD.n16286 DVDD.n2637 0.00334
R51827 DVDD.n16287 DVDD.n16286 0.00334
R51828 DVDD.n16288 DVDD.n16287 0.00334
R51829 DVDD.n16288 DVDD.n2634 0.00334
R51830 DVDD.n16295 DVDD.n2634 0.00334
R51831 DVDD.n16296 DVDD.n16295 0.00334
R51832 DVDD.n16297 DVDD.n16296 0.00334
R51833 DVDD.n16297 DVDD.n2631 0.00334
R51834 DVDD.n16304 DVDD.n2631 0.00334
R51835 DVDD.n16305 DVDD.n16304 0.00334
R51836 DVDD.n16306 DVDD.n16305 0.00334
R51837 DVDD.n16308 DVDD.n16306 0.00334
R51838 DVDD.n16308 DVDD.n16307 0.00334
R51839 DVDD.n16307 DVDD.n2569 0.00334
R51840 DVDD.n16319 DVDD.n2569 0.00334
R51841 DVDD.n16322 DVDD.n16321 0.00334
R51842 DVDD.n16323 DVDD.n16322 0.00334
R51843 DVDD.n16324 DVDD.n16323 0.00334
R51844 DVDD.n16325 DVDD.n16324 0.00334
R51845 DVDD.n16326 DVDD.n16325 0.00334
R51846 DVDD.n16327 DVDD.n16326 0.00334
R51847 DVDD.n16328 DVDD.n16327 0.00334
R51848 DVDD.n16329 DVDD.n16328 0.00334
R51849 DVDD.n16330 DVDD.n16329 0.00334
R51850 DVDD.n16331 DVDD.n16330 0.00334
R51851 DVDD.n16332 DVDD.n16331 0.00334
R51852 DVDD.n15426 DVDD.n15425 0.00334
R51853 DVDD.n15427 DVDD.n15426 0.00334
R51854 DVDD.n15428 DVDD.n15427 0.00334
R51855 DVDD.n15429 DVDD.n15428 0.00334
R51856 DVDD.n15430 DVDD.n15429 0.00334
R51857 DVDD.n15431 DVDD.n15430 0.00334
R51858 DVDD.n15432 DVDD.n15431 0.00334
R51859 DVDD.n15433 DVDD.n15432 0.00334
R51860 DVDD.n15434 DVDD.n15433 0.00334
R51861 DVDD.n15435 DVDD.n15434 0.00334
R51862 DVDD.n15435 DVDD.n5227 0.00334
R51863 DVDD.n15465 DVDD.n5227 0.00334
R51864 DVDD.n15468 DVDD.n15467 0.00334
R51865 DVDD.n15467 DVDD.n5224 0.00334
R51866 DVDD.n5224 DVDD.n5222 0.00334
R51867 DVDD.n15478 DVDD.n5222 0.00334
R51868 DVDD.n15479 DVDD.n15478 0.00334
R51869 DVDD.n15480 DVDD.n15479 0.00334
R51870 DVDD.n15480 DVDD.n5219 0.00334
R51871 DVDD.n15487 DVDD.n5219 0.00334
R51872 DVDD.n15488 DVDD.n15487 0.00334
R51873 DVDD.n15489 DVDD.n15488 0.00334
R51874 DVDD.n15489 DVDD.n5216 0.00334
R51875 DVDD.n15496 DVDD.n5216 0.00334
R51876 DVDD.n15497 DVDD.n15496 0.00334
R51877 DVDD.n15498 DVDD.n15497 0.00334
R51878 DVDD.n15499 DVDD.n15498 0.00334
R51879 DVDD.n15500 DVDD.n15499 0.00334
R51880 DVDD.n15501 DVDD.n15500 0.00334
R51881 DVDD.n15503 DVDD.n15501 0.00334
R51882 DVDD.n15504 DVDD.n15503 0.00334
R51883 DVDD.n15505 DVDD.n15504 0.00334
R51884 DVDD.n15506 DVDD.n15505 0.00334
R51885 DVDD.n15506 DVDD.n3228 0.00334
R51886 DVDD.n15915 DVDD.n3228 0.00334
R51887 DVDD.n15918 DVDD.n15917 0.00334
R51888 DVDD.n15918 DVDD.n3207 0.00334
R51889 DVDD.n15925 DVDD.n3207 0.00334
R51890 DVDD.n15926 DVDD.n15925 0.00334
R51891 DVDD.n15927 DVDD.n15926 0.00334
R51892 DVDD.n15927 DVDD.n3204 0.00334
R51893 DVDD.n15942 DVDD.n3204 0.00334
R51894 DVDD.n15943 DVDD.n15942 0.00334
R51895 DVDD.n15944 DVDD.n15943 0.00334
R51896 DVDD.n15945 DVDD.n15944 0.00334
R51897 DVDD.n15946 DVDD.n15945 0.00334
R51898 DVDD.n15949 DVDD.n15946 0.00334
R51899 DVDD.n15950 DVDD.n15949 0.00334
R51900 DVDD.n15951 DVDD.n15950 0.00334
R51901 DVDD.n15952 DVDD.n15951 0.00334
R51902 DVDD.n15953 DVDD.n15952 0.00334
R51903 DVDD.n15954 DVDD.n15953 0.00334
R51904 DVDD.n15955 DVDD.n15954 0.00334
R51905 DVDD.n15956 DVDD.n15955 0.00334
R51906 DVDD.n15957 DVDD.n15956 0.00334
R51907 DVDD.n15958 DVDD.n15957 0.00334
R51908 DVDD.n15959 DVDD.n15958 0.00334
R51909 DVDD.n15959 DVDD.n2706 0.00334
R51910 DVDD.n16260 DVDD.n2707 0.00334
R51911 DVDD.n2774 DVDD.n2707 0.00334
R51912 DVDD.n2775 DVDD.n2774 0.00334
R51913 DVDD.n2776 DVDD.n2775 0.00334
R51914 DVDD.n2777 DVDD.n2776 0.00334
R51915 DVDD.n2778 DVDD.n2777 0.00334
R51916 DVDD.n2843 DVDD.n2778 0.00334
R51917 DVDD.n2844 DVDD.n2843 0.00334
R51918 DVDD.n2845 DVDD.n2844 0.00334
R51919 DVDD.n2845 DVDD.n2841 0.00334
R51920 DVDD.n2852 DVDD.n2841 0.00334
R51921 DVDD.n2853 DVDD.n2852 0.00334
R51922 DVDD.n2854 DVDD.n2853 0.00334
R51923 DVDD.n2854 DVDD.n2838 0.00334
R51924 DVDD.n2861 DVDD.n2838 0.00334
R51925 DVDD.n2862 DVDD.n2861 0.00334
R51926 DVDD.n2863 DVDD.n2862 0.00334
R51927 DVDD.n2863 DVDD.n2835 0.00334
R51928 DVDD.n2877 DVDD.n2835 0.00334
R51929 DVDD.n2878 DVDD.n2877 0.00334
R51930 DVDD.n2879 DVDD.n2878 0.00334
R51931 DVDD.n2880 DVDD.n2879 0.00334
R51932 DVDD.n2881 DVDD.n2880 0.00334
R51933 DVDD.n16201 DVDD.n16200 0.00334
R51934 DVDD.n16202 DVDD.n16201 0.00334
R51935 DVDD.n16203 DVDD.n16202 0.00334
R51936 DVDD.n16204 DVDD.n16203 0.00334
R51937 DVDD.n16205 DVDD.n16204 0.00334
R51938 DVDD.n16206 DVDD.n16205 0.00334
R51939 DVDD.n16207 DVDD.n16206 0.00334
R51940 DVDD.n16208 DVDD.n16207 0.00334
R51941 DVDD.n16209 DVDD.n16208 0.00334
R51942 DVDD.n16210 DVDD.n16209 0.00334
R51943 DVDD.n15331 DVDD.n15323 0.00334
R51944 DVDD.n15332 DVDD.n15331 0.00334
R51945 DVDD.n15333 DVDD.n15332 0.00334
R51946 DVDD.n15333 DVDD.n15320 0.00334
R51947 DVDD.n15340 DVDD.n15320 0.00334
R51948 DVDD.n15341 DVDD.n15340 0.00334
R51949 DVDD.n15342 DVDD.n15341 0.00334
R51950 DVDD.n15343 DVDD.n15342 0.00334
R51951 DVDD.n15344 DVDD.n15343 0.00334
R51952 DVDD.n15345 DVDD.n15344 0.00334
R51953 DVDD.n15346 DVDD.n15345 0.00334
R51954 DVDD.n15347 DVDD.n15346 0.00334
R51955 DVDD.n15351 DVDD.n15350 0.00334
R51956 DVDD.n15352 DVDD.n15351 0.00334
R51957 DVDD.n15353 DVDD.n15352 0.00334
R51958 DVDD.n15354 DVDD.n15353 0.00334
R51959 DVDD.n15355 DVDD.n15354 0.00334
R51960 DVDD.n15356 DVDD.n15355 0.00334
R51961 DVDD.n15357 DVDD.n15356 0.00334
R51962 DVDD.n15358 DVDD.n15357 0.00334
R51963 DVDD.n15359 DVDD.n15358 0.00334
R51964 DVDD.n15360 DVDD.n15359 0.00334
R51965 DVDD.n15361 DVDD.n15360 0.00334
R51966 DVDD.n15362 DVDD.n15361 0.00334
R51967 DVDD.n15363 DVDD.n15362 0.00334
R51968 DVDD.n15365 DVDD.n15363 0.00334
R51969 DVDD.n15365 DVDD.n15364 0.00334
R51970 DVDD.n15364 DVDD.n3139 0.00334
R51971 DVDD.n3140 DVDD.n3139 0.00334
R51972 DVDD.n3141 DVDD.n3140 0.00334
R51973 DVDD.n3142 DVDD.n3141 0.00334
R51974 DVDD.n3143 DVDD.n3142 0.00334
R51975 DVDD.n3144 DVDD.n3143 0.00334
R51976 DVDD.n3145 DVDD.n3144 0.00334
R51977 DVDD.n3146 DVDD.n3145 0.00334
R51978 DVDD.n3225 DVDD.n3209 0.00334
R51979 DVDD.n3210 DVDD.n3209 0.00334
R51980 DVDD.n3211 DVDD.n3210 0.00334
R51981 DVDD.n3212 DVDD.n3211 0.00334
R51982 DVDD.n3213 DVDD.n3212 0.00334
R51983 DVDD.n3213 DVDD.n3055 0.00334
R51984 DVDD.n16088 DVDD.n3055 0.00334
R51985 DVDD.n16089 DVDD.n16088 0.00334
R51986 DVDD.n16090 DVDD.n16089 0.00334
R51987 DVDD.n16090 DVDD.n3051 0.00334
R51988 DVDD.n16096 DVDD.n3051 0.00334
R51989 DVDD.n16097 DVDD.n16096 0.00334
R51990 DVDD.n16099 DVDD.n16097 0.00334
R51991 DVDD.n16099 DVDD.n16098 0.00334
R51992 DVDD.n16098 DVDD.n3048 0.00334
R51993 DVDD.n3048 DVDD.n3046 0.00334
R51994 DVDD.n16120 DVDD.n3046 0.00334
R51995 DVDD.n16121 DVDD.n16120 0.00334
R51996 DVDD.n16122 DVDD.n16121 0.00334
R51997 DVDD.n16122 DVDD.n3043 0.00334
R51998 DVDD.n16129 DVDD.n3043 0.00334
R51999 DVDD.n16130 DVDD.n16129 0.00334
R52000 DVDD.n16131 DVDD.n16130 0.00334
R52001 DVDD.n16138 DVDD.n16137 0.00334
R52002 DVDD.n16138 DVDD.n2993 0.00334
R52003 DVDD.n16147 DVDD.n2993 0.00334
R52004 DVDD.n16148 DVDD.n16147 0.00334
R52005 DVDD.n16150 DVDD.n16148 0.00334
R52006 DVDD.n16150 DVDD.n16149 0.00334
R52007 DVDD.n16149 DVDD.n2989 0.00334
R52008 DVDD.n16158 DVDD.n2989 0.00334
R52009 DVDD.n16159 DVDD.n16158 0.00334
R52010 DVDD.n16160 DVDD.n16159 0.00334
R52011 DVDD.n16160 DVDD.n2986 0.00334
R52012 DVDD.n16167 DVDD.n2986 0.00334
R52013 DVDD.n16168 DVDD.n16167 0.00334
R52014 DVDD.n16169 DVDD.n16168 0.00334
R52015 DVDD.n16169 DVDD.n2983 0.00334
R52016 DVDD.n16176 DVDD.n2983 0.00334
R52017 DVDD.n16177 DVDD.n16176 0.00334
R52018 DVDD.n16178 DVDD.n16177 0.00334
R52019 DVDD.n16178 DVDD.n2922 0.00334
R52020 DVDD.n16187 DVDD.n2922 0.00334
R52021 DVDD.n16188 DVDD.n16187 0.00334
R52022 DVDD.n16191 DVDD.n16188 0.00334
R52023 DVDD.n16191 DVDD.n16190 0.00334
R52024 DVDD.n2884 DVDD.n2883 0.00334
R52025 DVDD.n2885 DVDD.n2884 0.00334
R52026 DVDD.n2886 DVDD.n2885 0.00334
R52027 DVDD.n2887 DVDD.n2886 0.00334
R52028 DVDD.n2888 DVDD.n2887 0.00334
R52029 DVDD.n2889 DVDD.n2888 0.00334
R52030 DVDD.n2890 DVDD.n2889 0.00334
R52031 DVDD.n2891 DVDD.n2890 0.00334
R52032 DVDD.n2892 DVDD.n2891 0.00334
R52033 DVDD.n2893 DVDD.n2892 0.00334
R52034 DVDD.n20214 DVDD.n20023 0.00332857
R52035 DVDD.n20706 DVDD.n19141 0.00332857
R52036 DVDD.n4008 DVDD.n244 0.00332857
R52037 DVDD.n9901 DVDD.n9621 0.00332857
R52038 DVDD.n18736 DVDD.n18729 0.00332857
R52039 DVDD.n4106 DVDD.n3634 0.00332
R52040 DVDD.n4176 DVDD.n4175 0.00332
R52041 DVDD.n4626 DVDD.n4224 0.00332
R52042 DVDD.n4105 DVDD.n3598 0.00332
R52043 DVDD.n15393 DVDD.n15348 0.00332
R52044 DVDD.n15469 DVDD.n5225 0.00332
R52045 DVDD.n15684 DVDD.n5113 0.00332
R52046 DVDD.n15760 DVDD.n3506 0.00332
R52047 DVDD.n15761 DVDD.n3505 0.00332
R52048 DVDD.n15836 DVDD.n3381 0.00332
R52049 DVDD.n2512 DVDD.n2432 0.00332
R52050 DVDD.n15686 DVDD.n15685 0.00332
R52051 DVDD.n3314 DVDD.n3272 0.00332
R52052 DVDD.n16302 DVDD.n2613 0.00332
R52053 DVDD.n15470 DVDD.n5111 0.00332
R52054 DVDD.n15940 DVDD.n3186 0.00332
R52055 DVDD.n2872 DVDD.n2865 0.00332
R52056 DVDD.n15395 DVDD.n15394 0.00332
R52057 DVDD.n16086 DVDD.n16085 0.00332
R52058 DVDD.n2981 DVDD.n2980 0.00332
R52059 DVDD.n4537 DVDD.n4393 0.0033125
R52060 DVDD.n19635 DVDD.n19633 0.00329474
R52061 DVDD.n22343 DVDD.n13 0.00329474
R52062 DVDD.n18499 DVDD.n18498 0.00329
R52063 DVDD.n21880 DVDD.n21779 0.00329
R52064 DVDD.n21918 DVDD.n21799 0.00329
R52065 DVDD.n21257 DVDD.n18664 0.00329
R52066 DVDD.n21946 DVDD.n18295 0.00329
R52067 DVDD.n21981 DVDD.n205 0.00329
R52068 DVDD.n21259 DVDD.n18661 0.00329
R52069 DVDD.n18376 DVDD.n18306 0.00329
R52070 DVDD.n18352 DVDD.n18267 0.00329
R52071 DVDD.n18496 DVDD.n18460 0.00329
R52072 DVDD.n21867 DVDD.n21866 0.00329
R52073 DVDD.n21916 DVDD.n21802 0.00329
R52074 DVDD.n20133 DVDD.n20074 0.00326429
R52075 DVDD.n20620 DVDD.n20605 0.00326429
R52076 DVDD.n3956 DVDD.n3923 0.00326429
R52077 DVDD.n9834 DVDD.n5472 0.00326429
R52078 DVDD.n19642 DVDD.n19190 0.00326429
R52079 DVDD.n4133 DVDD.n4132 0.00326
R52080 DVDD.n4502 DVDD.n4462 0.00326
R52081 DVDD DVDD.n475 0.00326
R52082 DVDD.n2539 DVDD 0.00326
R52083 DVDD.n16333 DVDD 0.00326
R52084 DVDD.n16212 DVDD 0.00326
R52085 DVDD.n2895 DVDD 0.00326
R52086 DVDD.n15790 DVDD.n15789 0.00326
R52087 DVDD.n15872 DVDD.n2346 0.00326
R52088 DVDD.n15651 DVDD.n15616 0.00326
R52089 DVDD.n15880 DVDD.n2698 0.00326
R52090 DVDD.n5208 DVDD.n5142 0.00326
R52091 DVDD.n15960 DVDD.n2757 0.00326
R52092 DVDD.n15368 DVDD.n3121 0.00326
R52093 DVDD.n16132 DVDD.n3038 0.00326
R52094 DVDD.n5508 DVDD.n5494 0.00324737
R52095 DVDD.n828 DVDD.n804 0.00324737
R52096 DVDD.n484 DVDD.n455 0.00323
R52097 DVDD.n2557 DVDD.n511 0.00323
R52098 DVDD.n16353 DVDD.n568 0.00323
R52099 DVDD.n16232 DVDD.n655 0.00323
R52100 DVDD.n2913 DVDD.n740 0.00323
R52101 DVDD.n5162 DVDD.n2723 0.00322195
R52102 DVDD.n5162 DVDD.n2769 0.00322195
R52103 DVDD.n16023 DVDD.n3001 0.00322195
R52104 DVDD.n16023 DVDD.n3017 0.00322195
R52105 DVDD.n5161 DVDD.n2793 0.00322195
R52106 DVDD.n5161 DVDD.n2791 0.00322195
R52107 DVDD.n16022 DVDD.n2930 0.00322195
R52108 DVDD.n16022 DVDD.n2946 0.00322195
R52109 DVDD.n5165 DVDD.n3163 0.00322195
R52110 DVDD.n5165 DVDD.n3161 0.00322195
R52111 DVDD.n16026 DVDD.n3091 0.00322195
R52112 DVDD.n16026 DVDD.n3072 0.00322195
R52113 DVDD.n5168 DVDD.n5167 0.00322195
R52114 DVDD.n5167 DVDD.n5158 0.00322195
R52115 DVDD.n16028 DVDD.n3128 0.00322195
R52116 DVDD.n16030 DVDD.n16028 0.00322195
R52117 DVDD.n13760 DVDD.n13759 0.00320677
R52118 DVDD.n13282 DVDD.n13281 0.00320677
R52119 DVDD.n20230 DVDD.n20028 0.0032
R52120 DVDD.n20308 DVDD.n19846 0.0032
R52121 DVDD.n20722 DVDD.n19146 0.0032
R52122 DVDD.n20798 DVDD.n18875 0.0032
R52123 DVDD.n4018 DVDD.n248 0.0032
R52124 DVDD.n411 DVDD.n383 0.0032
R52125 DVDD.n4420 DVDD.n3746 0.0032
R52126 DVDD.n3634 DVDD.n3633 0.0032
R52127 DVDD.n4116 DVDD.n4087 0.0032
R52128 DVDD.n4497 DVDD.n4190 0.0032
R52129 DVDD.n4271 DVDD.n4246 0.0032
R52130 DVDD.n3632 DVDD.n3598 0.0032
R52131 DVDD.n4455 DVDD.n4416 0.0032
R52132 DVDD.n4454 DVDD.n4453 0.0032
R52133 DVDD.n15772 DVDD.n3490 0.0032
R52134 DVDD.n15856 DVDD.n2342 0.0032
R52135 DVDD.n15635 DVDD.n15611 0.0032
R52136 DVDD.n15894 DVDD.n2693 0.0032
R52137 DVDD.n15481 DVDD.n5138 0.0032
R52138 DVDD.n15974 DVDD.n2753 0.0032
R52139 DVDD.n15382 DVDD.n3117 0.0032
R52140 DVDD.n16116 DVDD.n3033 0.0032
R52141 DVDD.n9909 DVDD.n9624 0.0032
R52142 DVDD.n9987 DVDD.n9959 0.0032
R52143 DVDD.n21108 DVDD.n18740 0.0032
R52144 DVDD.n22267 DVDD.n61 0.0032
R52145 DVDD.n5007 DVDD.n4886 0.00315263
R52146 DVDD.n5301 DVDD.n5056 0.00315263
R52147 DVDD.n5333 DVDD.n5245 0.00315263
R52148 DVDD.n5347 DVDD.n5234 0.00315263
R52149 DVDD.n5413 DVDD.n5396 0.00315263
R52150 DVDD.n15407 DVDD.n15316 0.00315263
R52151 DVDD.n18018 DVDD.n522 0.00315263
R52152 DVDD.n633 DVDD.n579 0.00315263
R52153 DVDD.n695 DVDD.n664 0.00315263
R52154 DVDD.n709 DVDD.n678 0.00315263
R52155 DVDD.n17952 DVDD.n748 0.00315263
R52156 DVDD.n17904 DVDD.n760 0.00315263
R52157 DVDD.n3626 DVDD.n3528 0.00314375
R52158 DVDD.n4110 DVDD.n4086 0.00314
R52159 DVDD.n15765 DVDD.n3489 0.00314
R52160 DVDD.n15610 DVDD.n15535 0.00314
R52161 DVDD.n15474 DVDD.n5137 0.00314
R52162 DVDD.n15388 DVDD.n3116 0.00314
R52163 DVDD.n22232 DVDD 0.0031254
R52164 DVDD.n21923 DVDD 0.0031254
R52165 DVDD.n18136 DVDD.n454 0.00311
R52166 DVDD.n2563 DVDD.n510 0.00311
R52167 DVDD.n17978 DVDD.n569 0.00311
R52168 DVDD.n17963 DVDD.n656 0.00311
R52169 DVDD.n16196 DVDD.n739 0.00311
R52170 DVDD.n20164 DVDD.n20070 0.00310526
R52171 DVDD.n20121 DVDD.n20060 0.00310526
R52172 DVDD.n20118 DVDD.n20069 0.00310526
R52173 DVDD.n20116 DVDD.n20061 0.00310526
R52174 DVDD.n20114 DVDD.n20068 0.00310526
R52175 DVDD.n20112 DVDD.n20062 0.00310526
R52176 DVDD.n20110 DVDD.n20067 0.00310526
R52177 DVDD.n20108 DVDD.n20063 0.00310526
R52178 DVDD.n20106 DVDD.n20066 0.00310526
R52179 DVDD.n20104 DVDD.n20064 0.00310526
R52180 DVDD.n20102 DVDD.n20065 0.00310526
R52181 DVDD.n18929 DVDD.n18927 0.00310526
R52182 DVDD.n20885 DVDD.n20884 0.00310526
R52183 DVDD.n20882 DVDD.n18937 0.00310526
R52184 DVDD.n20881 DVDD.n18946 0.00310526
R52185 DVDD.n20878 DVDD.n18956 0.00310526
R52186 DVDD.n20876 DVDD.n18947 0.00310526
R52187 DVDD.n20874 DVDD.n18955 0.00310526
R52188 DVDD.n20872 DVDD.n18948 0.00310526
R52189 DVDD.n20870 DVDD.n18954 0.00310526
R52190 DVDD.n20868 DVDD.n18949 0.00310526
R52191 DVDD.n20866 DVDD.n18953 0.00310526
R52192 DVDD.n21228 DVDD.n21225 0.00309529
R52193 DVDD.n22187 DVDD.n227 0.00309529
R52194 DVDD.n21249 DVDD.n18667 0.00309529
R52195 DVDD.n22028 DVDD.n234 0.00309529
R52196 DVDD.n18454 DVDD.n126 0.00309529
R52197 DVDD.n18235 DVDD.n18234 0.00309529
R52198 DVDD.n18486 DVDD.n122 0.00309529
R52199 DVDD.n22055 DVDD.n18221 0.00309529
R52200 DVDD.n19503 DVDD.n96 0.00309024
R52201 DVDD.n19288 DVDD.n52 0.00309024
R52202 DVDD.n19553 DVDD.n18732 0.00309024
R52203 DVDD.n19235 DVDD.n18694 0.00309024
R52204 DVDD.n4429 DVDD.n3750 0.0030875
R52205 DVDD.n4124 DVDD.n4091 0.00308
R52206 DVDD.n4501 DVDD.n4195 0.00308
R52207 DVDD.n15781 DVDD.n3494 0.00308
R52208 DVDD.n15865 DVDD.n2345 0.00308
R52209 DVDD.n15644 DVDD.n15615 0.00308
R52210 DVDD.n15886 DVDD.n2697 0.00308
R52211 DVDD.n15490 DVDD.n5141 0.00308
R52212 DVDD.n15966 DVDD.n2756 0.00308
R52213 DVDD.n15374 DVDD.n3120 0.00308
R52214 DVDD.n16125 DVDD.n3037 0.00308
R52215 DVDD.n20286 DVDD.n19873 0.00307143
R52216 DVDD.n20420 DVDD.n19850 0.00307143
R52217 DVDD.n19057 DVDD.n19022 0.00307143
R52218 DVDD.n20814 DVDD.n18876 0.00307143
R52219 DVDD.n320 DVDD.n304 0.00307143
R52220 DVDD.n22138 DVDD.n388 0.00307143
R52221 DVDD.n9696 DVDD.n9680 0.00307143
R52222 DVDD.n10055 DVDD.n9964 0.00307143
R52223 DVDD.n22253 DVDD.n93 0.00307143
R52224 DVDD.n22300 DVDD.n22299 0.00307143
R52225 DVDD.n22226 DVDD.n160 0.00305
R52226 DVDD.n18387 DVDD.n176 0.00305
R52227 DVDD.n22045 DVDD.n18239 0.00305
R52228 DVDD.n21355 DVDD.n18509 0.00305
R52229 DVDD.n21706 DVDD.n21705 0.00305
R52230 DVDD.n22036 DVDD.n21986 0.00305
R52231 DVDD.n21357 DVDD.n21339 0.00305
R52232 DVDD.n21669 DVDD.n18520 0.00305
R52233 DVDD.n21983 DVDD.n225 0.00305
R52234 DVDD.n21585 DVDD.n162 0.00305
R52235 DVDD.n21758 DVDD.n18402 0.00305
R52236 DVDD.n22047 DVDD.n18224 0.00305
R52237 DVDD.n480 DVDD.n458 0.00305
R52238 DVDD.n2549 DVDD.n514 0.00305
R52239 DVDD.n16345 DVDD.n562 0.00305
R52240 DVDD.n16224 DVDD.n649 0.00305
R52241 DVDD.n2905 DVDD.n743 0.00305
R52242 DVDD.n4532 DVDD.n4505 0.00302
R52243 DVDD.n4655 DVDD.n4228 0.00302
R52244 DVDD.n16394 DVDD.n2349 0.00302
R52245 DVDD.n2483 DVDD.n2424 0.00302
R52246 DVDD.n16271 DVDD.n16270 0.00302
R52247 DVDD.n2606 DVDD.n2571 0.00302
R52248 DVDD.n16255 DVDD.n2767 0.00302
R52249 DVDD.n2832 DVDD.n2816 0.00302
R52250 DVDD.n16145 DVDD.n16144 0.00302
R52251 DVDD.n16185 DVDD.n2924 0.00302
R52252 DVDD.n20346 DVDD.n18933 0.00300714
R52253 DVDD.n20841 DVDD.n18962 0.00300714
R52254 DVDD.n22100 DVDD.n22072 0.00300714
R52255 DVDD.n10029 DVDD.n788 0.00300714
R52256 DVDD.n22321 DVDD.n17 0.00300714
R52257 DVDD.n3596 DVDD.n3558 0.00299
R52258 DVDD.n15753 DVDD.n15752 0.00299
R52259 DVDD.n15688 DVDD.n5048 0.00299
R52260 DVDD.n15462 DVDD.n15461 0.00299
R52261 DVDD.n15408 DVDD.n5394 0.00299
R52262 DVDD.n3733 DVDD.n3727 0.002975
R52263 DVDD.n5009 DVDD.n4886 0.00296316
R52264 DVDD.n5299 DVDD.n5056 0.00296316
R52265 DVDD.n5331 DVDD.n5245 0.00296316
R52266 DVDD.n5349 DVDD.n5234 0.00296316
R52267 DVDD.n5415 DVDD.n5396 0.00296316
R52268 DVDD.n15407 DVDD.n5406 0.00296316
R52269 DVDD.n18016 DVDD.n522 0.00296316
R52270 DVDD.n631 DVDD.n579 0.00296316
R52271 DVDD.n693 DVDD.n664 0.00296316
R52272 DVDD.n711 DVDD.n678 0.00296316
R52273 DVDD.n17949 DVDD.n748 0.00296316
R52274 DVDD.n17906 DVDD.n760 0.00296316
R52275 DVDD.n4160 DVDD.n3809 0.00296
R52276 DVDD.n4629 DVDD.n4219 0.00296
R52277 DVDD.n15826 DVDD.n3391 0.00296
R52278 DVDD.n2503 DVDD.n2435 0.00296
R52279 DVDD.n3305 DVDD.n3281 0.00296
R52280 DVDD.n16293 DVDD.n2616 0.00296
R52281 DVDD.n15923 DVDD.n3189 0.00296
R52282 DVDD.n2855 DVDD.n2820 0.00296
R52283 DVDD.n3217 DVDD.n3076 0.00296
R52284 DVDD.n2984 DVDD.n2959 0.00296
R52285 DVDD.n20193 DVDD.n19727 0.00294286
R52286 DVDD.n19947 DVDD.n19888 0.00294286
R52287 DVDD.n20685 DVDD.n18834 0.00294286
R52288 DVDD.n20760 DVDD.n19038 0.00294286
R52289 DVDD.n4054 DVDD.n3865 0.00294286
R52290 DVDD.n342 DVDD.n295 0.00294286
R52291 DVDD.n9891 DVDD.n9759 0.00294286
R52292 DVDD.n9714 DVDD.n9684 0.00294286
R52293 DVDD.n21204 DVDD.n18678 0.00294286
R52294 DVDD.n21124 DVDD.n109 0.00294286
R52295 DVDD.n3585 DVDD.n3562 0.00293
R52296 DVDD.n15738 DVDD.n15711 0.00293
R52297 DVDD.n5098 DVDD.n5051 0.00293
R52298 DVDD.n15447 DVDD.n15420 0.00293
R52299 DVDD.n15336 DVDD.n5377 0.00293
R52300 DVDD.n3616 DVDD.n3538 0.00291875
R52301 DVDD.n11934 DVDD.n11927 0.00291611
R52302 DVDD.n13279 DVDD.n12781 0.00291611
R52303 DVDD.n11932 DVDD.n11928 0.00291611
R52304 DVDD.n13280 DVDD.n12898 0.00291611
R52305 DVDD.n20284 DVDD.n19884 0.00291463
R52306 DVDD.n19935 DVDD.n19874 0.00291463
R52307 DVDD.n19932 DVDD.n19883 0.00291463
R52308 DVDD.n19930 DVDD.n19875 0.00291463
R52309 DVDD.n19928 DVDD.n19882 0.00291463
R52310 DVDD.n19926 DVDD.n19876 0.00291463
R52311 DVDD.n19924 DVDD.n19881 0.00291463
R52312 DVDD.n19922 DVDD.n19877 0.00291463
R52313 DVDD.n19920 DVDD.n19880 0.00291463
R52314 DVDD.n19918 DVDD.n19878 0.00291463
R52315 DVDD.n19916 DVDD.n19879 0.00291463
R52316 DVDD.n20425 DVDD.n19832 0.00291463
R52317 DVDD.n20422 DVDD.n20421 0.00291463
R52318 DVDD.n20419 DVDD.n19842 0.00291463
R52319 DVDD.n20418 DVDD.n19851 0.00291463
R52320 DVDD.n20415 DVDD.n20377 0.00291463
R52321 DVDD.n20412 DVDD.n19852 0.00291463
R52322 DVDD.n20410 DVDD.n20376 0.00291463
R52323 DVDD.n20407 DVDD.n19853 0.00291463
R52324 DVDD.n20405 DVDD.n20375 0.00291463
R52325 DVDD.n20402 DVDD.n19854 0.00291463
R52326 DVDD.n20400 DVDD.n20374 0.00291463
R52327 DVDD.n20243 DVDD.n19969 0.00291463
R52328 DVDD.n20022 DVDD.n19959 0.00291463
R52329 DVDD.n20019 DVDD.n19968 0.00291463
R52330 DVDD.n20017 DVDD.n19960 0.00291463
R52331 DVDD.n20015 DVDD.n19967 0.00291463
R52332 DVDD.n20013 DVDD.n19961 0.00291463
R52333 DVDD.n20011 DVDD.n19966 0.00291463
R52334 DVDD.n20009 DVDD.n19962 0.00291463
R52335 DVDD.n20007 DVDD.n19965 0.00291463
R52336 DVDD.n20005 DVDD.n19963 0.00291463
R52337 DVDD.n20003 DVDD.n19964 0.00291463
R52338 DVDD.n19721 DVDD.n19719 0.00291463
R52339 DVDD.n20577 DVDD.n19722 0.00291463
R52340 DVDD.n20574 DVDD.n20573 0.00291463
R52341 DVDD.n19741 DVDD.n19732 0.00291463
R52342 DVDD.n20571 DVDD.n19751 0.00291463
R52343 DVDD.n20570 DVDD.n19742 0.00291463
R52344 DVDD.n20567 DVDD.n19750 0.00291463
R52345 DVDD.n20564 DVDD.n19743 0.00291463
R52346 DVDD.n20562 DVDD.n19749 0.00291463
R52347 DVDD.n20559 DVDD.n19744 0.00291463
R52348 DVDD.n20557 DVDD.n19748 0.00291463
R52349 DVDD.n4149 DVDD.n3813 0.0029
R52350 DVDD.n3411 DVDD.n3395 0.0029
R52351 DVDD.n15669 DVDD.n3285 0.0029
R52352 DVDD.n15509 DVDD.n3193 0.0029
R52353 DVDD.n15998 DVDD.n3080 0.0029
R52354 DVDD.n5173 DVDD.n2720 0.00287073
R52355 DVDD.n16034 DVDD.n3020 0.00287073
R52356 DVDD.n16045 DVDD.n3024 0.00287073
R52357 DVDD.n5172 DVDD.n2789 0.00287073
R52358 DVDD.n16033 DVDD.n2950 0.00287073
R52359 DVDD.n16044 DVDD.n2955 0.00287073
R52360 DVDD.n5176 DVDD.n3159 0.00287073
R52361 DVDD.n16037 DVDD.n3101 0.00287073
R52362 DVDD.n16048 DVDD.n3073 0.00287073
R52363 DVDD.n5178 DVDD.n5154 0.00287073
R52364 DVDD.n16040 DVDD.n16039 0.00287073
R52365 DVDD.n16051 DVDD.n16050 0.00287073
R52366 DVDD.n3583 DVDD.n3553 0.00287
R52367 DVDD.n15742 DVDD.n4900 0.00287
R52368 DVDD.n5085 DVDD.n5042 0.00287
R52369 DVDD.n15451 DVDD.n5256 0.00287
R52370 DVDD.n15321 DVDD.n5375 0.00287
R52371 DVDD.n5506 DVDD.n5494 0.00286842
R52372 DVDD.n826 DVDD.n804 0.00286842
R52373 DVDD.n4434 DVDD.n3737 0.0028625
R52374 DVDD.n4575 DVDD.n4250 0.0028625
R52375 DVDD.n493 DVDD.n492 0.00286
R52376 DVDD.n2567 DVDD.n2566 0.00286
R52377 DVDD.n16321 DVDD.n16320 0.00286
R52378 DVDD.n16200 DVDD.n2568 0.00286
R52379 DVDD.n16189 DVDD.n2883 0.00286
R52380 DVDD.n3577 DVDD.n3555 0.00285923
R52381 DVDD.n4088 DVDD.n4082 0.00285923
R52382 DVDD.n3815 DVDD.n3811 0.00285923
R52383 DVDD.n4162 DVDD.n3807 0.00285923
R52384 DVDD.n4530 DVDD.n4493 0.00285923
R52385 DVDD.n4529 DVDD.n4528 0.00285923
R52386 DVDD.n4634 DVDD.n4631 0.00285923
R52387 DVDD.n4641 DVDD.n4627 0.00285923
R52388 DVDD.n473 DVDD.n451 0.00285923
R52389 DVDD.n15713 DVDD.n4896 0.00285923
R52390 DVDD.n15708 DVDD.n4902 0.00285923
R52391 DVDD.n3491 DVDD.n3484 0.00285923
R52392 DVDD.n15792 DVDD.n3419 0.00285923
R52393 DVDD.n3398 DVDD.n3393 0.00285923
R52394 DVDD.n3403 DVDD.n3389 0.00285923
R52395 DVDD.n2360 DVDD.n2339 0.00285923
R52396 DVDD.n2359 DVDD.n2335 0.00285923
R52397 DVDD.n2437 DVDD.n2401 0.00285923
R52398 DVDD.n2484 DVDD.n2433 0.00285923
R52399 DVDD.n531 DVDD.n507 0.00285923
R52400 DVDD.n18040 DVDD.n18039 0.00285923
R52401 DVDD.n5079 DVDD.n5040 0.00285923
R52402 DVDD.n5078 DVDD.n5044 0.00285923
R52403 DVDD.n15612 DVDD.n15603 0.00285923
R52404 DVDD.n15617 DVDD.n15593 0.00285923
R52405 DVDD.n3288 DVDD.n3283 0.00285923
R52406 DVDD.n3292 DVDD.n3279 0.00285923
R52407 DVDD.n2694 DVDD.n2689 0.00285923
R52408 DVDD.n2699 DVDD.n2685 0.00285923
R52409 DVDD.n2621 DVDD.n2618 0.00285923
R52410 DVDD.n2626 DVDD.n2614 0.00285923
R52411 DVDD.n581 DVDD.n556 0.00285923
R52412 DVDD.n580 DVDD.n558 0.00285923
R52413 DVDD.n15422 DVDD.n5254 0.00285923
R52414 DVDD.n15417 DVDD.n5258 0.00285923
R52415 DVDD.n5157 DVDD.n5133 0.00285923
R52416 DVDD.n5156 DVDD.n5129 0.00285923
R52417 DVDD.n3195 DVDD.n3191 0.00285923
R52418 DVDD.n15937 DVDD.n15930 0.00285923
R52419 DVDD.n2768 DVDD.n2750 0.00285923
R52420 DVDD.n2764 DVDD.n2722 0.00285923
R52421 DVDD.n2823 DVDD.n2822 0.00285923
R52422 DVDD.n2828 DVDD.n2818 0.00285923
R52423 DVDD.n668 DVDD.n643 0.00285923
R52424 DVDD.n667 DVDD.n645 0.00285923
R52425 DVDD.n5408 DVDD.n5373 0.00285923
R52426 DVDD.n5407 DVDD.n5371 0.00285923
R52427 DVDD.n3135 DVDD.n3112 0.00285923
R52428 DVDD.n16061 DVDD.n16053 0.00285923
R52429 DVDD.n9777 DVDD.n3078 0.00285923
R52430 DVDD.n16081 DVDD.n3095 0.00285923
R52431 DVDD.n3034 DVDD.n3030 0.00285923
R52432 DVDD.n3039 DVDD.n3026 0.00285923
R52433 DVDD.n2964 DVDD.n2961 0.00285923
R52434 DVDD.n2969 DVDD.n2957 0.00285923
R52435 DVDD.n759 DVDD.n735 0.00285923
R52436 DVDD.n758 DVDD.n731 0.00285923
R52437 DVDD.n3035 DVDD.n3034 0.00285923
R52438 DVDD.n3040 DVDD.n3039 0.00285923
R52439 DVDD.n2768 DVDD.n2754 0.00285923
R52440 DVDD.n16257 DVDD.n2722 0.00285923
R52441 DVDD.n2695 DVDD.n2694 0.00285923
R52442 DVDD.n2700 DVDD.n2699 0.00285923
R52443 DVDD.n2360 DVDD.n2343 0.00285923
R52444 DVDD.n2359 DVDD.n2347 0.00285923
R52445 DVDD.n4530 DVDD.n4498 0.00285923
R52446 DVDD.n4529 DVDD.n4503 0.00285923
R52447 DVDD.n2965 DVDD.n2964 0.00285923
R52448 DVDD.n2970 DVDD.n2969 0.00285923
R52449 DVDD.n2824 DVDD.n2823 0.00285923
R52450 DVDD.n2829 DVDD.n2828 0.00285923
R52451 DVDD.n2622 DVDD.n2621 0.00285923
R52452 DVDD.n2627 DVDD.n2626 0.00285923
R52453 DVDD.n16370 DVDD.n2401 0.00285923
R52454 DVDD.n2484 DVDD.n2480 0.00285923
R52455 DVDD.n4635 DVDD.n4634 0.00285923
R52456 DVDD.n4642 DVDD.n4641 0.00285923
R52457 DVDD.n9777 DVDD.n3083 0.00285923
R52458 DVDD.n16083 DVDD.n3095 0.00285923
R52459 DVDD.n3196 DVDD.n3195 0.00285923
R52460 DVDD.n15930 DVDD.n3199 0.00285923
R52461 DVDD.n3289 DVDD.n3288 0.00285923
R52462 DVDD.n3293 DVDD.n3292 0.00285923
R52463 DVDD.n3399 DVDD.n3398 0.00285923
R52464 DVDD.n3404 DVDD.n3403 0.00285923
R52465 DVDD.n3816 DVDD.n3815 0.00285923
R52466 DVDD.n4163 DVDD.n4162 0.00285923
R52467 DVDD.n3577 DVDD.n3560 0.00285923
R52468 DVDD.n15709 DVDD.n15708 0.00285923
R52469 DVDD.n15714 DVDD.n15713 0.00285923
R52470 DVDD.n15698 DVDD.n5044 0.00285923
R52471 DVDD.n5081 DVDD.n5040 0.00285923
R52472 DVDD.n15423 DVDD.n15422 0.00285923
R52473 DVDD.n15418 DVDD.n15417 0.00285923
R52474 DVDD.n15317 DVDD.n5373 0.00285923
R52475 DVDD.n15406 DVDD.n5371 0.00285923
R52476 DVDD.n759 DVDD.n741 0.00285923
R52477 DVDD.n758 DVDD.n745 0.00285923
R52478 DVDD.n668 DVDD.n654 0.00285923
R52479 DVDD.n667 DVDD.n651 0.00285923
R52480 DVDD.n581 DVDD.n567 0.00285923
R52481 DVDD.n580 DVDD.n564 0.00285923
R52482 DVDD.n531 DVDD.n512 0.00285923
R52483 DVDD.n18039 DVDD.n516 0.00285923
R52484 DVDD.n473 DVDD.n456 0.00285923
R52485 DVDD.n3135 DVDD.n3118 0.00285923
R52486 DVDD.n16053 DVDD.n3122 0.00285923
R52487 DVDD.n5157 DVDD.n5139 0.00285923
R52488 DVDD.n5156 DVDD.n5143 0.00285923
R52489 DVDD.n15613 DVDD.n15612 0.00285923
R52490 DVDD.n15618 DVDD.n15617 0.00285923
R52491 DVDD.n3492 DVDD.n3491 0.00285923
R52492 DVDD.n15793 DVDD.n15792 0.00285923
R52493 DVDD.n4089 DVDD.n4088 0.00285923
R52494 DVDD.n4159 DVDD.n3762 0.00284
R52495 DVDD.n4638 DVDD.n4637 0.00284
R52496 DVDD.n15821 DVDD.n3401 0.00284
R52497 DVDD.n2498 DVDD.n2478 0.00284
R52498 DVDD.n3290 DVDD.n3248 0.00284
R52499 DVDD.n16289 DVDD.n2624 0.00284
R52500 DVDD.n15919 DVDD.n3197 0.00284
R52501 DVDD.n2850 DVDD.n2826 0.00284
R52502 DVDD.n3221 DVDD.n3085 0.00284
R52503 DVDD.n16163 DVDD.n2967 0.00284
R52504 DVDD.n19094 DVDD.n19028 0.00282683
R52505 DVDD.n19103 DVDD.n18896 0.00282683
R52506 DVDD.n19124 DVDD.n19123 0.00282683
R52507 DVDD.n20972 DVDD.n18829 0.00282683
R52508 DVDD.n20177 DVDD.n19731 0.00281429
R52509 DVDD.n20669 DVDD.n18838 0.00281429
R52510 DVDD.n3993 DVDD.n3869 0.00281429
R52511 DVDD.n9875 DVDD.n9763 0.00281429
R52512 DVDD.n21213 DVDD.n18691 0.00281429
R52513 DVDD.n3592 DVDD.n3557 0.00281
R52514 DVDD.n15728 DVDD.n4904 0.00281
R52515 DVDD.n15692 DVDD.n5046 0.00281
R52516 DVDD.n15437 DVDD.n5260 0.00281
R52517 DVDD.n15400 DVDD.n5369 0.00281
R52518 DVDD.n4179 DVDD.n3771 0.00278
R52519 DVDD.n4657 DVDD.n4225 0.00278
R52520 DVDD DVDD.n18156 0.00278
R52521 DVDD DVDD.n2537 0.00278
R52522 DVDD DVDD.n16210 0.00278
R52523 DVDD DVDD.n2893 0.00278
R52524 DVDD.n15839 DVDD.n3347 0.00278
R52525 DVDD.n2514 DVDD.n2482 0.00278
R52526 DVDD.n15907 DVDD.n3295 0.00278
R52527 DVDD.n16312 DVDD.n2629 0.00278
R52528 DVDD.n15987 DVDD.n3201 0.00278
R52529 DVDD.n2873 DVDD.n2831 0.00278
R52530 DVDD.n3068 DVDD.n3053 0.00278
R52531 DVDD.n16182 DVDD.n16180 0.00278
R52532 DVDD.n5025 DVDD.n3514 0.00277368
R52533 DVDD.n5036 DVDD.n3511 0.00277368
R52534 DVDD.n5272 DVDD.n5068 0.00277368
R52535 DVDD.n5283 DVDD.n5071 0.00277368
R52536 DVDD.n5315 DVDD.n5241 0.00277368
R52537 DVDD.n5365 DVDD.n5252 0.00277368
R52538 DVDD.n5431 DVDD.n5389 0.00277368
R52539 DVDD.n5442 DVDD.n5386 0.00277368
R52540 DVDD.n18000 DVDD.n535 0.00277368
R52541 DVDD.n17989 DVDD.n532 0.00277368
R52542 DVDD.n604 DVDD.n590 0.00277368
R52543 DVDD.n615 DVDD.n577 0.00277368
R52544 DVDD.n17968 DVDD.n639 0.00277368
R52545 DVDD.n727 DVDD.n680 0.00277368
R52546 DVDD.n17933 DVDD.n768 0.00277368
R52547 DVDD.n17922 DVDD.n765 0.00277368
R52548 DVDD.n22229 DVDD.n148 0.00275
R52549 DVDD.n21944 DVDD.n18299 0.00275
R52550 DVDD.n22039 DVDD.n18241 0.00275
R52551 DVDD.n22229 DVDD.n146 0.00275
R52552 DVDD.n21944 DVDD.n194 0.00275
R52553 DVDD.n22039 DVDD.n18242 0.00275
R52554 DVDD.n22229 DVDD.n139 0.00275
R52555 DVDD.n21944 DVDD.n18377 0.00275
R52556 DVDD.n22039 DVDD.n18248 0.00275
R52557 DVDD.n21226 DVDD.n18432 0.00275
R52558 DVDD.n22209 DVDD.n186 0.00275
R52559 DVDD.n18353 DVDD.n223 0.00275
R52560 DVDD.n18668 DVDD.n18432 0.00275
R52561 DVDD.n22209 DVDD.n22208 0.00275
R52562 DVDD.n223 DVDD.n206 0.00275
R52563 DVDD.n18501 DVDD.n18432 0.00275
R52564 DVDD.n22209 DVDD.n181 0.00275
R52565 DVDD.n21832 DVDD.n223 0.00275
R52566 DVDD.n18489 DVDD.n18432 0.00275
R52567 DVDD.n22209 DVDD.n188 0.00275
R52568 DVDD.n21909 DVDD.n223 0.00275
R52569 DVDD.n22229 DVDD.n151 0.00275
R52570 DVDD.n21944 DVDD.n18383 0.00275
R52571 DVDD.n22039 DVDD.n18264 0.00275
R52572 DVDD.n3713 DVDD.n3709 0.00275
R52573 DVDD.n4157 DVDD.n3817 0.00275
R52574 DVDD.n18154 DVDD.n449 0.00275
R52575 DVDD.n4275 DVDD.n4248 0.00275
R52576 DVDD.n4759 DVDD.n4758 0.00275
R52577 DVDD.n3760 DVDD.n3755 0.00275
R52578 DVDD.n4559 DVDD.n4323 0.00275
R52579 DVDD.n2545 DVDD.n505 0.00275
R52580 DVDD.n16341 DVDD.n560 0.00275
R52581 DVDD.n16220 DVDD.n647 0.00275
R52582 DVDD.n2901 DVDD.n733 0.00275
R52583 DVDD.n18096 DVDD.n18054 0.00273371
R52584 DVDD.n4092 DVDD.n4080 0.00272
R52585 DVDD.n4158 DVDD.n4157 0.00272
R52586 DVDD.n4491 DVDD.n4197 0.00272
R52587 DVDD.n3495 DVDD.n3482 0.00272
R52588 DVDD.n15813 DVDD.n3400 0.00272
R52589 DVDD.n3334 DVDD.n2337 0.00272
R52590 DVDD.n15649 DVDD.n15601 0.00272
R52591 DVDD.n3235 DVDD.n3148 0.00272
R52592 DVDD.n15882 DVDD.n2687 0.00272
R52593 DVDD.n15494 DVDD.n5131 0.00272
R52594 DVDD.n15990 DVDD.n15989 0.00272
R52595 DVDD.n15962 DVDD.n2748 0.00272
R52596 DVDD.n15370 DVDD.n3110 0.00272
R52597 DVDD.n15991 DVDD.n3084 0.00272
R52598 DVDD.n3041 DVDD.n3028 0.00272
R52599 DVDD.n4699 DVDD.n4698 0.0027
R52600 DVDD.n15875 DVDD.n2703 0.0027
R52601 DVDD.n16263 DVDD.n16262 0.0027
R52602 DVDD.n16261 DVDD.n16260 0.0027
R52603 DVDD.n16137 DVDD.n2705 0.0027
R52604 DVDD.n4386 DVDD.n4385 0.00269512
R52605 DVDD.n4362 DVDD.n3731 0.00269512
R52606 DVDD.n4371 DVDD.n3650 0.00269512
R52607 DVDD.n18085 DVDD.n18084 0.00269375
R52608 DVDD.n18537 DVDD.n18536 0.00269003
R52609 DVDD.n21363 DVDD.n21362 0.00269003
R52610 DVDD.n22007 DVDD.n21992 0.00269003
R52611 DVDD.n4850 DVDD.n3547 0.00269003
R52612 DVDD.n482 DVDD.n453 0.00269
R52613 DVDD.n2559 DVDD.n509 0.00269
R52614 DVDD.n16355 DVDD.n554 0.00269
R52615 DVDD.n16234 DVDD.n641 0.00269
R52616 DVDD.n2915 DVDD.n737 0.00269
R52617 DVDD.n20184 DVDD.n19729 0.00268571
R52618 DVDD.n19950 DVDD.n19890 0.00268571
R52619 DVDD.n20676 DVDD.n18836 0.00268571
R52620 DVDD.n20751 DVDD.n19040 0.00268571
R52621 DVDD.n3898 DVDD.n3867 0.00268571
R52622 DVDD.n333 DVDD.n297 0.00268571
R52623 DVDD.n9882 DVDD.n9761 0.00268571
R52624 DVDD.n9686 DVDD.n9667 0.00268571
R52625 DVDD.n19674 DVDD.n18681 0.00268571
R52626 DVDD.n21121 DVDD.n111 0.00268571
R52627 DVDD.n15287 DVDD.n5468 0.00267895
R52628 DVDD.n17878 DVDD.n792 0.00267895
R52629 DVDD.n21721 DVDD 0.00267716
R52630 DVDD.n22193 DVDD 0.00267716
R52631 DVDD.n8250 DVDD.n8150 0.00266541
R52632 DVDD.n4101 DVDD.n4084 0.00266
R52633 DVDD.n4496 DVDD.n4495 0.00266
R52634 DVDD.n15770 DVDD.n3486 0.00266
R52635 DVDD.n15854 DVDD.n2341 0.00266
R52636 DVDD.n15633 DVDD.n15605 0.00266
R52637 DVDD.n15896 DVDD.n2691 0.00266
R52638 DVDD.n5220 DVDD.n5135 0.00266
R52639 DVDD.n15976 DVDD.n2752 0.00266
R52640 DVDD.n15384 DVDD.n3114 0.00266
R52641 DVDD.n16114 DVDD.n16113 0.00266
R52642 DVDD.n4459 DVDD.n4403 0.0026375
R52643 DVDD.n903 DVDD.n891 0.0026375
R52644 DVDD.n17362 DVDD.n905 0.0026375
R52645 DVDD.n5995 DVDD.n5578 0.0026375
R52646 DVDD.n5993 DVDD.n5992 0.0026375
R52647 DVDD.n20355 DVDD.n18935 0.00262143
R52648 DVDD.n20832 DVDD.n18964 0.00262143
R52649 DVDD.n22074 DVDD.n446 0.00262143
R52650 DVDD.n10038 DVDD.n786 0.00262143
R52651 DVDD.n22329 DVDD.n15 0.00262143
R52652 DVDD.n16398 DVDD.n2296 0.00260732
R52653 DVDD.n2473 DVDD.n2412 0.00260732
R52654 DVDD.n4977 DVDD.n3369 0.00260732
R52655 DVDD.n4980 DVDD.n3472 0.00260732
R52656 DVDD.n4099 DVDD.n4084 0.0026
R52657 DVDD.n4495 DVDD.n4187 0.0026
R52658 DVDD.n4577 DVDD.n4281 0.0026
R52659 DVDD.n3501 DVDD.n3486 0.0026
R52660 DVDD.n15848 DVDD.n2341 0.0026
R52661 DVDD.n15631 DVDD.n15605 0.0026
R52662 DVDD.n3322 DVDD.n2691 0.0026
R52663 DVDD.n15476 DVDD.n5135 0.0026
R52664 DVDD.n15948 DVDD.n2752 0.0026
R52665 DVDD.n15386 DVDD.n3114 0.0026
R52666 DVDD.n16113 DVDD.n16102 0.0026
R52667 DVDD.n5021 DVDD.n4889 0.00258421
R52668 DVDD.n15751 DVDD.n15706 0.00258421
R52669 DVDD.n5268 DVDD.n5063 0.00258421
R52670 DVDD.n5287 DVDD.n5059 0.00258421
R52671 DVDD.n5319 DVDD.n5242 0.00258421
R52672 DVDD.n5361 DVDD.n5231 0.00258421
R52673 DVDD.n5427 DVDD.n5399 0.00258421
R52674 DVDD.n5446 DVDD.n5403 0.00258421
R52675 DVDD.n18004 DVDD.n525 0.00258421
R52676 DVDD.n17985 DVDD.n529 0.00258421
R52677 DVDD.n600 DVDD.n575 0.00258421
R52678 DVDD.n619 DVDD.n572 0.00258421
R52679 DVDD.n17964 DVDD.n648 0.00258421
R52680 DVDD.n723 DVDD.n669 0.00258421
R52681 DVDD.n17937 DVDD.n751 0.00258421
R52682 DVDD.n17918 DVDD.n755 0.00258421
R52683 DVDD.n18138 DVDD.n453 0.00257
R52684 DVDD.n2561 DVDD.n509 0.00257
R52685 DVDD.n583 DVDD.n554 0.00257
R52686 DVDD.n670 DVDD.n641 0.00257
R52687 DVDD.n2917 DVDD.n737 0.00257
R52688 DVDD.n20200 DVDD.n19725 0.00255714
R52689 DVDD.n20275 DVDD.n19886 0.00255714
R52690 DVDD.n20692 DVDD.n18832 0.00255714
R52691 DVDD.n20767 DVDD.n19036 0.00255714
R52692 DVDD.n4047 DVDD.n3863 0.00255714
R52693 DVDD.n324 DVDD.n293 0.00255714
R52694 DVDD.n9939 DVDD.n9814 0.00255714
R52695 DVDD.n9701 DVDD.n9682 0.00255714
R52696 DVDD.n18715 DVDD.n18674 0.00255714
R52697 DVDD.n21130 DVDD.n107 0.00255714
R52698 DVDD.n4126 DVDD.n4080 0.00254
R52699 DVDD.n4491 DVDD.n4196 0.00254
R52700 DVDD.n4736 DVDD.n4735 0.00254
R52701 DVDD.n15818 DVDD.n15817 0.00254
R52702 DVDD.n3233 DVDD.n3227 0.00254
R52703 DVDD.n15917 DVDD.n15916 0.00254
R52704 DVDD.n3226 DVDD.n3225 0.00254
R52705 DVDD.n15783 DVDD.n3482 0.00254
R52706 DVDD.n15867 DVDD.n2337 0.00254
R52707 DVDD.n15623 DVDD.n15601 0.00254
R52708 DVDD.n15884 DVDD.n2687 0.00254
R52709 DVDD.n15492 DVDD.n5131 0.00254
R52710 DVDD.n15964 DVDD.n2748 0.00254
R52711 DVDD.n15372 DVDD.n3110 0.00254
R52712 DVDD.n16127 DVDD.n3028 0.00254
R52713 DVDD.n3639 DVDD.n3635 0.002525
R52714 DVDD.n8037 DVDD.n8036 0.002525
R52715 DVDD.n15538 DVDD.n2655 0.00251951
R52716 DVDD.n5184 DVDD.n2718 0.00251951
R52717 DVDD.n3104 DVDD.n3023 0.00251951
R52718 DVDD.n16011 DVDD.n2996 0.00251951
R52719 DVDD.n15537 DVDD.n2582 0.00251951
R52720 DVDD.n5183 DVDD.n2787 0.00251951
R52721 DVDD.n3103 DVDD.n2954 0.00251951
R52722 DVDD.n16010 DVDD.n2925 0.00251951
R52723 DVDD.n15541 DVDD.n3246 0.00251951
R52724 DVDD.n5187 DVDD.n3157 0.00251951
R52725 DVDD.n16082 DVDD.n16071 0.00251951
R52726 DVDD.n16014 DVDD.n3058 0.00251951
R52727 DVDD.n15543 DVDD.n5128 0.00251951
R52728 DVDD.n5189 DVDD.n5152 0.00251951
R52729 DVDD.n16069 DVDD.n16068 0.00251951
R52730 DVDD.n16016 DVDD.n3124 0.00251951
R52731 DVDD.n21766 DVDD.n21765 0.00251708
R52732 DVDD.n21728 DVDD.n21727 0.00251708
R52733 DVDD.n22064 DVDD.n22063 0.00251708
R52734 DVDD.n18067 DVDD.n18065 0.00251708
R52735 DVDD.n22229 DVDD.n154 0.00251
R52736 DVDD.n21944 DVDD.n177 0.00251
R52737 DVDD.n22039 DVDD.n18230 0.00251
R52738 DVDD.n22229 DVDD.n144 0.00251
R52739 DVDD.n21944 DVDD.n18300 0.00251
R52740 DVDD.n22039 DVDD.n18249 0.00251
R52741 DVDD.n22229 DVDD.n142 0.00251
R52742 DVDD.n21944 DVDD.n18303 0.00251
R52743 DVDD.n22039 DVDD.n224 0.00251
R52744 DVDD.n18546 DVDD.n18432 0.00251
R52745 DVDD.n22209 DVDD.n185 0.00251
R52746 DVDD.n22191 DVDD.n223 0.00251
R52747 DVDD.n21719 DVDD.n18432 0.00251
R52748 DVDD.n22209 DVDD.n193 0.00251
R52749 DVDD.n22025 DVDD.n223 0.00251
R52750 DVDD.n18451 DVDD.n18432 0.00251
R52751 DVDD.n22210 DVDD.n22209 0.00251
R52752 DVDD.n18232 DVDD.n223 0.00251
R52753 DVDD.n21584 DVDD.n18432 0.00251
R52754 DVDD.n22209 DVDD.n189 0.00251
R52755 DVDD.n18226 DVDD.n223 0.00251
R52756 DVDD.n22229 DVDD.n149 0.00251
R52757 DVDD.n21944 DVDD.n18381 0.00251
R52758 DVDD.n22039 DVDD.n18227 0.00251
R52759 DVDD.n18152 DVDD.n449 0.00251
R52760 DVDD.n2547 DVDD.n505 0.00251
R52761 DVDD.n16343 DVDD.n560 0.00251
R52762 DVDD.n16222 DVDD.n647 0.00251
R52763 DVDD.n2903 DVDD.n733 0.00251
R52764 DVDD.n20339 DVDD.n18931 0.00249286
R52765 DVDD.n18996 DVDD.n18995 0.00249286
R52766 DVDD.n22114 DVDD.n22109 0.00249286
R52767 DVDD.n10022 DVDD.n790 0.00249286
R52768 DVDD.n22351 DVDD.n1 0.00249286
R52769 DVDD.n5510 DVDD.n5488 0.00248947
R52770 DVDD.n830 DVDD.n812 0.00248947
R52771 DVDD.n4180 DVDD.n4179 0.00248
R52772 DVDD.n4657 DVDD.n4656 0.00248
R52773 DVDD.n15840 DVDD.n15839 0.00248
R52774 DVDD.n2516 DVDD.n2482 0.00248
R52775 DVDD.n15907 DVDD.n15906 0.00248
R52776 DVDD.n16312 DVDD.n16311 0.00248
R52777 DVDD.n15987 DVDD.n15986 0.00248
R52778 DVDD.n2875 DVDD.n2831 0.00248
R52779 DVDD.n16092 DVDD.n3053 0.00248
R52780 DVDD.n16182 DVDD.n16181 0.00248
R52781 DVDD.n18022 DVDD.n542 0.00245652
R52782 DVDD.n17728 DVDD.n877 0.00245652
R52783 DVDD.n5004 DVDD.n4906 0.00245652
R52784 DVDD.n15149 DVDD.n15148 0.00245652
R52785 DVDD.n3595 DVDD.n3557 0.00245
R52786 DVDD DVDD.n459 0.00245
R52787 DVDD.n4904 DVDD.n3510 0.00245
R52788 DVDD DVDD.n515 0.00245
R52789 DVDD.n15690 DVDD.n5046 0.00245
R52790 DVDD DVDD.n563 0.00245
R52791 DVDD.n5260 DVDD.n5229 0.00245
R52792 DVDD DVDD.n650 0.00245
R52793 DVDD.n5382 DVDD.n5369 0.00245
R52794 DVDD DVDD.n744 0.00245
R52795 DVDD.n8252 DVDD.n8153 0.00243289
R52796 DVDD.n14310 DVDD.n8151 0.00243289
R52797 DVDD.n9941 DVDD.n9676 0.00243171
R52798 DVDD.n9940 DVDD.n9745 0.00243171
R52799 DVDD.n9944 DVDD.n9639 0.00243171
R52800 DVDD.n9947 DVDD.n9946 0.00243171
R52801 DVDD.n20242 DVDD.n20241 0.00242857
R52802 DVDD.n20317 DVDD.n19848 0.00242857
R52803 DVDD.n20734 DVDD.n20733 0.00242857
R52804 DVDD.n20807 DVDD.n18878 0.00242857
R52805 DVDD.n274 DVDD.n250 0.00242857
R52806 DVDD.n421 DVDD.n386 0.00242857
R52807 DVDD.n10084 DVDD.n9625 0.00242857
R52808 DVDD.n9997 DVDD.n9962 0.00242857
R52809 DVDD.n21112 DVDD.n18742 0.00242857
R52810 DVDD.n22271 DVDD.n63 0.00242857
R52811 DVDD.n4159 DVDD.n3763 0.00242
R52812 DVDD.n4638 DVDD.n4218 0.00242
R52813 DVDD.n3408 DVDD.n3401 0.00242
R52814 DVDD.n2492 DVDD.n2478 0.00242
R52815 DVDD.n3303 DVDD.n3290 0.00242
R52816 DVDD.n16291 DVDD.n2624 0.00242
R52817 DVDD.n15921 DVDD.n3197 0.00242
R52818 DVDD.n2839 DVDD.n2826 0.00242
R52819 DVDD.n3219 DVDD.n3085 0.00242
R52820 DVDD.n16165 DVDD.n2967 0.00242
R52821 DVDD.n4767 DVDD.n3668 0.0024125
R52822 DVDD.n4413 DVDD.n4406 0.0024125
R52823 DVDD.n5005 DVDD.n3518 0.00239474
R52824 DVDD.n5303 DVDD.n5075 0.00239474
R52825 DVDD.n5335 DVDD.n5237 0.00239474
R52826 DVDD.n5345 DVDD.n5248 0.00239474
R52827 DVDD.n5411 DVDD.n5393 0.00239474
R52828 DVDD.n18020 DVDD.n539 0.00239474
R52829 DVDD.n635 DVDD.n593 0.00239474
R52830 DVDD.n697 DVDD.n661 0.00239474
R52831 DVDD.n707 DVDD.n672 0.00239474
R52832 DVDD.n17953 DVDD.n772 0.00239474
R52833 DVDD.n3584 DVDD.n3553 0.00239
R52834 DVDD.n15740 DVDD.n4900 0.00239
R52835 DVDD.n5096 DVDD.n5042 0.00239
R52836 DVDD.n15449 DVDD.n5256 0.00239
R52837 DVDD.n15334 DVDD.n5375 0.00239
R52838 DVDD.n4781 DVDD.n3599 0.00238
R52839 DVDD.n15759 DVDD.n15757 0.00238
R52840 DVDD.n5114 DVDD.n3507 0.00238
R52841 DVDD.n15468 DVDD.n15466 0.00238
R52842 DVDD.n15350 DVDD.n5226 0.00238
R52843 DVDD.n20130 DVDD.n20072 0.00236429
R52844 DVDD.n20647 DVDD.n20617 0.00236429
R52845 DVDD.n3947 DVDD.n3925 0.00236429
R52846 DVDD.n9831 DVDD.n5474 0.00236429
R52847 DVDD.n19638 DVDD.n19188 0.00236429
R52848 DVDD.n4147 DVDD.n3813 0.00236
R52849 DVDD.n15804 DVDD.n3395 0.00236
R52850 DVDD.n15672 DVDD.n3285 0.00236
R52851 DVDD.n15512 DVDD.n3193 0.00236
R52852 DVDD.n16001 DVDD.n3080 0.00236
R52853 DVDD.n18072 DVDD.n18058 0.00235625
R52854 DVDD.n3584 DVDD.n3562 0.00233
R52855 DVDD.n15740 DVDD.n15711 0.00233
R52856 DVDD.n5096 DVDD.n5051 0.00233
R52857 DVDD.n15449 DVDD.n15420 0.00233
R52858 DVDD.n15334 DVDD.n5377 0.00233
R52859 DVDD.n20340 DVDD 0.0023
R52860 DVDD.n20223 DVDD.n20026 0.0023
R52861 DVDD.n20301 DVDD.n19844 0.0023
R52862 DVDD.n20339 DVDD 0.0023
R52863 DVDD DVDD.n18997 0.0023
R52864 DVDD.n20715 DVDD.n19144 0.0023
R52865 DVDD.n19016 DVDD.n18873 0.0023
R52866 DVDD.n18996 DVDD 0.0023
R52867 DVDD.n22108 DVDD 0.0023
R52868 DVDD.n4011 DVDD.n246 0.0023
R52869 DVDD.n404 DVDD.n381 0.0023
R52870 DVDD.n22109 DVDD 0.0023
R52871 DVDD.n3713 DVDD.n3712 0.0023
R52872 DVDD.n3611 DVDD.n3540 0.0023
R52873 DVDD.n3809 DVDD.n3763 0.0023
R52874 DVDD.n4629 DVDD.n4218 0.0023
R52875 DVDD.n4456 DVDD.n4415 0.0023
R52876 DVDD.n4781 DVDD.n3600 0.0023
R52877 DVDD.n3612 DVDD.n3541 0.0023
R52878 DVDD.n4536 DVDD.n4202 0.0023
R52879 DVDD.n4535 DVDD.n4534 0.0023
R52880 DVDD.n3408 DVDD.n3391 0.0023
R52881 DVDD.n2492 DVDD.n2435 0.0023
R52882 DVDD.n3303 DVDD.n3281 0.0023
R52883 DVDD.n16291 DVDD.n2616 0.0023
R52884 DVDD.n15921 DVDD.n3189 0.0023
R52885 DVDD.n2839 DVDD.n2820 0.0023
R52886 DVDD.n3219 DVDD.n3076 0.0023
R52887 DVDD.n16165 DVDD.n2959 0.0023
R52888 DVDD.n10023 DVDD 0.0023
R52889 DVDD.n9905 DVDD.n9622 0.0023
R52890 DVDD.n9980 DVDD.n9957 0.0023
R52891 DVDD.n10022 DVDD 0.0023
R52892 DVDD.n21177 DVDD.n18738 0.0023
R52893 DVDD.n22290 DVDD.n59 0.0023
R52894 DVDD DVDD.n22351 0.0023
R52895 DVDD.n22350 DVDD 0.0023
R52896 DVDD.n3595 DVDD.n3558 0.00227
R52897 DVDD.n15752 DVDD.n3510 0.00227
R52898 DVDD.n15690 DVDD.n5048 0.00227
R52899 DVDD.n15461 DVDD.n5229 0.00227
R52900 DVDD.n15408 DVDD.n5382 0.00227
R52901 DVDD.n8032 DVDD.n7776 0.00226856
R52902 DVDD.n14834 DVDD.n8024 0.00226856
R52903 DVDD.n4532 DVDD.n4208 0.00224
R52904 DVDD.n4656 DVDD.n4655 0.00224
R52905 DVDD.n16394 DVDD.n2362 0.00224
R52906 DVDD.n2516 DVDD.n2424 0.00224
R52907 DVDD.n16270 DVDD.n2640 0.00224
R52908 DVDD.n16311 DVDD.n2606 0.00224
R52909 DVDD.n16255 DVDD.n16254 0.00224
R52910 DVDD.n2875 DVDD.n2816 0.00224
R52911 DVDD.n16144 DVDD.n2991 0.00224
R52912 DVDD.n16181 DVDD.n2924 0.00224
R52913 DVDD.n20143 DVDD.n20076 0.00223571
R52914 DVDD.n20630 DVDD.n20607 0.00223571
R52915 DVDD.n3971 DVDD.n3966 0.00223571
R52916 DVDD.n9842 DVDD.n5470 0.00223571
R52917 DVDD.n19653 DVDD.n19192 0.00223571
R52918 DVDD.n22226 DVDD.n154 0.00221
R52919 DVDD.n18387 DVDD.n177 0.00221
R52920 DVDD.n22045 DVDD.n18230 0.00221
R52921 DVDD.n21355 DVDD.n144 0.00221
R52922 DVDD.n21705 DVDD.n18300 0.00221
R52923 DVDD.n22036 DVDD.n18249 0.00221
R52924 DVDD.n21357 DVDD.n142 0.00221
R52925 DVDD.n18520 DVDD.n18303 0.00221
R52926 DVDD.n21983 DVDD.n224 0.00221
R52927 DVDD.n162 DVDD.n149 0.00221
R52928 DVDD.n21758 DVDD.n18381 0.00221
R52929 DVDD.n22047 DVDD.n18227 0.00221
R52930 DVDD.n18152 DVDD.n458 0.00221
R52931 DVDD.n2547 DVDD.n514 0.00221
R52932 DVDD.n16343 DVDD.n562 0.00221
R52933 DVDD.n16222 DVDD.n649 0.00221
R52934 DVDD.n2903 DVDD.n743 0.00221
R52935 DVDD.n5011 DVDD.n3517 0.00220526
R52936 DVDD.n5297 DVDD.n5074 0.00220526
R52937 DVDD.n5329 DVDD.n5238 0.00220526
R52938 DVDD.n5351 DVDD.n5249 0.00220526
R52939 DVDD.n5417 DVDD.n5392 0.00220526
R52940 DVDD.n5456 DVDD.n5383 0.00220526
R52941 DVDD.n18014 DVDD.n538 0.00220526
R52942 DVDD.n629 DVDD.n585 0.00220526
R52943 DVDD.n691 DVDD.n674 0.00220526
R52944 DVDD.n713 DVDD.n659 0.00220526
R52945 DVDD.n17947 DVDD.n771 0.00220526
R52946 DVDD.n17908 DVDD.n762 0.00220526
R52947 DVDD.n4444 DVDD.n3739 0.0021875
R52948 DVDD.n4600 DVDD.n4258 0.0021875
R52949 DVDD.n4126 DVDD.n4091 0.00218
R52950 DVDD.n4501 DVDD.n4196 0.00218
R52951 DVDD.n15783 DVDD.n3494 0.00218
R52952 DVDD.n15867 DVDD.n2345 0.00218
R52953 DVDD.n15623 DVDD.n15615 0.00218
R52954 DVDD.n15884 DVDD.n2697 0.00218
R52955 DVDD.n15492 DVDD.n5141 0.00218
R52956 DVDD.n15964 DVDD.n2756 0.00218
R52957 DVDD.n15372 DVDD.n3120 0.00218
R52958 DVDD.n16127 DVDD.n3037 0.00218
R52959 DVDD.n20216 DVDD.n19976 0.00217143
R52960 DVDD.n20294 DVDD.n19841 0.00217143
R52961 DVDD.n20708 DVDD.n19139 0.00217143
R52962 DVDD.n20929 DVDD.n18887 0.00217143
R52963 DVDD.n4031 DVDD.n242 0.00217143
R52964 DVDD.n22141 DVDD.n22140 0.00217143
R52965 DVDD.n9922 DVDD.n9619 0.00217143
R52966 DVDD.n10058 DVDD.n10057 0.00217143
R52967 DVDD.n21184 DVDD.n21100 0.00217143
R52968 DVDD.n22297 DVDD.n79 0.00217143
R52969 DVDD.n15547 DVDD.n2653 0.00216829
R52970 DVDD.n15522 DVDD.n2712 0.00216829
R52971 DVDD.n5195 DVDD.n2716 0.00216829
R52972 DVDD.n16143 DVDD.n3032 0.00216829
R52973 DVDD.n15546 DVDD.n2580 0.00216829
R52974 DVDD.n15521 DVDD.n2781 0.00216829
R52975 DVDD.n5194 DVDD.n2785 0.00216829
R52976 DVDD.n16183 DVDD.n2963 0.00216829
R52977 DVDD.n15550 DVDD.n3244 0.00216829
R52978 DVDD.n15524 DVDD.n3151 0.00216829
R52979 DVDD.n5197 DVDD.n3155 0.00216829
R52980 DVDD.n16084 DVDD.n3081 0.00216829
R52981 DVDD.n15552 DVDD.n5126 0.00216829
R52982 DVDD.n15526 DVDD.n5146 0.00216829
R52983 DVDD.n5199 DVDD.n5150 0.00216829
R52984 DVDD.n16066 DVDD.n16065 0.00216829
R52985 DVDD.n18138 DVDD.n454 0.00215
R52986 DVDD.n2561 DVDD.n510 0.00215
R52987 DVDD.n17978 DVDD.n583 0.00215
R52988 DVDD.n17963 DVDD.n670 0.00215
R52989 DVDD.n2917 DVDD.n739 0.00215
R52990 DVDD.n3624 DVDD.n3525 0.00213125
R52991 DVDD.n15116 DVDD.n5997 0.00212406
R52992 DVDD.n14574 DVDD.n8133 0.00212406
R52993 DVDD.n4099 DVDD.n4086 0.00212
R52994 DVDD.n3501 DVDD.n3489 0.00212
R52995 DVDD.n15631 DVDD.n15610 0.00212
R52996 DVDD.n15476 DVDD.n5137 0.00212
R52997 DVDD.n15386 DVDD.n3116 0.00212
R52998 DVDD.n5504 DVDD.n5489 0.00211053
R52999 DVDD.n824 DVDD.n809 0.00211053
R53000 DVDD.n20152 DVDD.n20127 0.00210714
R53001 DVDD.n20639 DVDD.n20614 0.00210714
R53002 DVDD.n3943 DVDD.n3930 0.00210714
R53003 DVDD.n9851 DVDD.n5481 0.00210714
R53004 DVDD.n19644 DVDD.n19198 0.00210714
R53005 DVDD.n9799 DVDD.n9662 0.00208049
R53006 DVDD.n9798 DVDD.n9733 0.00208049
R53007 DVDD.n9802 DVDD.n9627 0.00208049
R53008 DVDD.n9804 DVDD.n9774 0.00208049
R53009 DVDD.n4427 DVDD.n3735 0.002075
R53010 DVDD.n12280 DVDD.n12279 0.002075
R53011 DVDD.n16730 DVDD.n1808 0.002075
R53012 DVDD.n4101 DVDD.n4087 0.00206
R53013 DVDD.n4497 DVDD.n4496 0.00206
R53014 DVDD.n15770 DVDD.n3490 0.00206
R53015 DVDD.n15854 DVDD.n2342 0.00206
R53016 DVDD.n15633 DVDD.n15611 0.00206
R53017 DVDD.n15896 DVDD.n2693 0.00206
R53018 DVDD.n5220 DVDD.n5138 0.00206
R53019 DVDD.n15976 DVDD.n2753 0.00206
R53020 DVDD.n15384 DVDD.n3117 0.00206
R53021 DVDD.n16114 DVDD.n3033 0.00206
R53022 DVDD.n20232 DVDD.n19972 0.00204286
R53023 DVDD.n20310 DVDD.n19837 0.00204286
R53024 DVDD.n20724 DVDD.n19135 0.00204286
R53025 DVDD.n19013 DVDD.n18883 0.00204286
R53026 DVDD.n4014 DVDD.n238 0.00204286
R53027 DVDD.n413 DVDD.n375 0.00204286
R53028 DVDD.n9643 DVDD.n9615 0.00204286
R53029 DVDD.n9989 DVDD.n9752 0.00204286
R53030 DVDD.n21169 DVDD.n21095 0.00204286
R53031 DVDD.n22282 DVDD.n74 0.00204286
R53032 DVDD.n482 DVDD.n455 0.00203
R53033 DVDD.n2559 DVDD.n511 0.00203
R53034 DVDD.n16355 DVDD.n568 0.00203
R53035 DVDD.n16234 DVDD.n655 0.00203
R53036 DVDD.n2915 DVDD.n740 0.00203
R53037 DVDD.n5027 DVDD.n4890 0.00201579
R53038 DVDD.n5034 DVDD.n4892 0.00201579
R53039 DVDD.n5274 DVDD.n5062 0.00201579
R53040 DVDD.n5281 DVDD.n5060 0.00201579
R53041 DVDD.n5253 DVDD.n5230 0.00201579
R53042 DVDD.n5433 DVDD.n5400 0.00201579
R53043 DVDD.n5440 DVDD.n5402 0.00201579
R53044 DVDD.n17998 DVDD.n526 0.00201579
R53045 DVDD.n17991 DVDD.n528 0.00201579
R53046 DVDD.n606 DVDD.n573 0.00201579
R53047 DVDD.n613 DVDD.n587 0.00201579
R53048 DVDD.n681 DVDD.n657 0.00201579
R53049 DVDD.n17931 DVDD.n752 0.00201579
R53050 DVDD.n17924 DVDD.n754 0.00201579
R53051 DVDD.n3677 DVDD.n3665 0.00201227
R53052 DVDD.n21721 DVDD.n18507 0.002
R53053 DVDD.n22207 DVDD.n196 0.002
R53054 DVDD.n22194 DVDD.n22193 0.002
R53055 DVDD.n21721 DVDD.n18505 0.002
R53056 DVDD.n18320 DVDD.n196 0.002
R53057 DVDD.n22193 DVDD.n221 0.002
R53058 DVDD.n21721 DVDD.n18502 0.002
R53059 DVDD.n21837 DVDD.n196 0.002
R53060 DVDD.n22193 DVDD.n214 0.002
R53061 DVDD.n21721 DVDD.n18450 0.002
R53062 DVDD.n21862 DVDD.n196 0.002
R53063 DVDD.n22193 DVDD.n211 0.002
R53064 DVDD.n4133 DVDD.n4092 0.002
R53065 DVDD.n4502 DVDD.n4197 0.002
R53066 DVDD.n4757 DVDD.n3673 0.002
R53067 DVDD.n4737 DVDD.n4736 0.002
R53068 DVDD.n15790 DVDD.n3495 0.002
R53069 DVDD.n3334 DVDD.n2346 0.002
R53070 DVDD.n15649 DVDD.n15616 0.002
R53071 DVDD.n15882 DVDD.n2698 0.002
R53072 DVDD.n15494 DVDD.n5142 0.002
R53073 DVDD.n15962 DVDD.n2757 0.002
R53074 DVDD.n15370 DVDD.n3121 0.002
R53075 DVDD.n3041 DVDD.n3038 0.002
R53076 DVDD.n4352 DVDD.n4265 0.00199268
R53077 DVDD.n18498 DVDD.n148 0.00197
R53078 DVDD.n21779 DVDD.n18299 0.00197
R53079 DVDD.n21918 DVDD.n18241 0.00197
R53080 DVDD.n21257 DVDD.n146 0.00197
R53081 DVDD.n21946 DVDD.n194 0.00197
R53082 DVDD.n21981 DVDD.n18242 0.00197
R53083 DVDD.n21259 DVDD.n139 0.00197
R53084 DVDD.n18377 DVDD.n18376 0.00197
R53085 DVDD.n18267 DVDD.n18248 0.00197
R53086 DVDD.n18496 DVDD.n151 0.00197
R53087 DVDD.n21866 DVDD.n18383 0.00197
R53088 DVDD.n21916 DVDD.n18264 0.00197
R53089 DVDD.n18154 DVDD.n459 0.00197
R53090 DVDD.n2545 DVDD.n515 0.00197
R53091 DVDD.n16341 DVDD.n563 0.00197
R53092 DVDD.n16220 DVDD.n650 0.00197
R53093 DVDD.n2901 DVDD.n744 0.00197
R53094 DVDD.n4741 DVDD.n3753 0.0019625
R53095 DVDD.n4567 DVDD.n4244 0.0019625
R53096 DVDD.n15114 DVDD.n5999 0.00194966
R53097 DVDD.n8149 DVDD.n8148 0.00194966
R53098 DVDD.n15115 DVDD.n5998 0.00194966
R53099 DVDD.n14576 DVDD.n14575 0.00194966
R53100 DVDD.n3634 DVDD.n3597 0.00194
R53101 DVDD.n4175 DVDD.n3771 0.00194
R53102 DVDD.n4626 DVDD.n4225 0.00194
R53103 DVDD.n4783 DVDD.n3598 0.00194
R53104 DVDD.n15397 DVDD.n15348 0.00194
R53105 DVDD.n15464 DVDD.n5225 0.00194
R53106 DVDD.n5113 DVDD.n5110 0.00194
R53107 DVDD.n15755 DVDD.n3506 0.00194
R53108 DVDD.n15754 DVDD.n3505 0.00194
R53109 DVDD.n3381 DVDD.n3347 0.00194
R53110 DVDD.n2514 DVDD.n2432 0.00194
R53111 DVDD.n15687 DVDD.n15686 0.00194
R53112 DVDD.n3295 DVDD.n3272 0.00194
R53113 DVDD.n2629 DVDD.n2613 0.00194
R53114 DVDD.n15463 DVDD.n5111 0.00194
R53115 DVDD.n3201 DVDD.n3186 0.00194
R53116 DVDD.n2873 DVDD.n2872 0.00194
R53117 DVDD.n15396 DVDD.n15395 0.00194
R53118 DVDD.n16085 DVDD.n3068 0.00194
R53119 DVDD.n16180 DVDD.n2980 0.00194
R53120 DVDD.n15286 DVDD.n5476 0.00192105
R53121 DVDD.n816 DVDD.n811 0.00192105
R53122 DVDD.n20572 DVDD.n19745 0.00191429
R53123 DVDD.n20283 DVDD.n20282 0.00191429
R53124 DVDD.n20970 DVDD.n18853 0.00191429
R53125 DVDD.n20777 DVDD.n20776 0.00191429
R53126 DVDD.n4065 DVDD.n3883 0.00191429
R53127 DVDD.n22149 DVDD.n303 0.00191429
R53128 DVDD.n9948 DVDD.n9807 0.00191429
R53129 DVDD.n9727 DVDD.n9695 0.00191429
R53130 DVDD.n18720 DVDD.n18702 0.00191429
R53131 DVDD.n22254 DVDD.n89 0.00191429
R53132 DVDD.n3592 DVDD.n3559 0.00191
R53133 DVDD.n15728 DVDD.n15707 0.00191
R53134 DVDD.n15692 DVDD.n5049 0.00191
R53135 DVDD.n15437 DVDD.n15416 0.00191
R53136 DVDD.n15400 DVDD.n5381 0.00191
R53137 DVDD.n3618 DVDD.n3530 0.00190625
R53138 DVDD.n2306 DVDD.n2294 0.00190488
R53139 DVDD.n2413 DVDD.n2390 0.00190488
R53140 DVDD.n3370 DVDD.n3348 0.00190488
R53141 DVDD.n3473 DVDD.n3420 0.00190488
R53142 DVDD.n3810 DVDD.n3762 0.00188
R53143 DVDD.n4637 DVDD.n4630 0.00188
R53144 DVDD.n15821 DVDD.n3392 0.00188
R53145 DVDD.n2498 DVDD.n2436 0.00188
R53146 DVDD.n15909 DVDD.n3248 0.00188
R53147 DVDD.n16289 DVDD.n2617 0.00188
R53148 DVDD.n15919 DVDD.n3190 0.00188
R53149 DVDD.n2850 DVDD.n2821 0.00188
R53150 DVDD.n3221 DVDD.n3077 0.00188
R53151 DVDD.n16163 DVDD.n2960 0.00188
R53152 DVDD.n11940 DVDD.n11924 0.00187555
R53153 DVDD.n16728 DVDD.n1810 0.00187555
R53154 DVDD.n12278 DVDD.n11942 0.00187555
R53155 DVDD.n16729 DVDD.n1809 0.00187555
R53156 DVDD.n18313 DVDD.n18312 0.00185574
R53157 DVDD.n21221 DVDD.n18658 0.00185574
R53158 DVDD.n18338 DVDD.n18333 0.00185574
R53159 DVDD.n4875 DVDD.n4874 0.00185574
R53160 DVDD.n20348 DVDD.n18941 0.00185
R53161 DVDD.n19000 DVDD.n18969 0.00185
R53162 DVDD.n22090 DVDD.n22077 0.00185
R53163 DVDD.n4423 DVDD.n3748 0.00185
R53164 DVDD.n3583 DVDD.n3563 0.00185
R53165 DVDD.n4278 DVDD.n4241 0.00185
R53166 DVDD.n18134 DVDD.n488 0.00185
R53167 DVDD.n4587 DVDD.n490 0.00185
R53168 DVDD.n15742 DVDD.n15712 0.00185
R53169 DVDD.n5085 DVDD.n5052 0.00185
R53170 DVDD.n15451 DVDD.n15421 0.00185
R53171 DVDD.n15321 DVDD.n5378 0.00185
R53172 DVDD.n10031 DVDD.n797 0.00185
R53173 DVDD.n22313 DVDD.n24 0.00185
R53174 DVDD.n21721 DVDD.n21720 0.00184
R53175 DVDD.n18517 DVDD.n196 0.00184
R53176 DVDD.n22193 DVDD.n219 0.00184
R53177 DVDD.n21721 DVDD.n18504 0.00184
R53178 DVDD.n21666 DVDD.n196 0.00184
R53179 DVDD.n22193 DVDD.n22192 0.00184
R53180 DVDD.n21721 DVDD.n18452 0.00184
R53181 DVDD.n196 DVDD.n175 0.00184
R53182 DVDD.n22193 DVDD.n215 0.00184
R53183 DVDD.n21721 DVDD.n18449 0.00184
R53184 DVDD.n21746 DVDD.n196 0.00184
R53185 DVDD.n22193 DVDD.n210 0.00184
R53186 DVDD.n5019 DVDD.n3515 0.00182632
R53187 DVDD.n5266 DVDD.n5067 0.00182632
R53188 DVDD.n5289 DVDD.n5072 0.00182632
R53189 DVDD.n5321 DVDD.n5240 0.00182632
R53190 DVDD.n5359 DVDD.n5251 0.00182632
R53191 DVDD.n5425 DVDD.n5390 0.00182632
R53192 DVDD.n5448 DVDD.n5385 0.00182632
R53193 DVDD.n18006 DVDD.n536 0.00182632
R53194 DVDD.n598 DVDD.n589 0.00182632
R53195 DVDD.n621 DVDD.n592 0.00182632
R53196 DVDD.n683 DVDD.n662 0.00182632
R53197 DVDD.n721 DVDD.n671 0.00182632
R53198 DVDD.n17939 DVDD.n769 0.00182632
R53199 DVDD.n17916 DVDD.n764 0.00182632
R53200 DVDD.n4149 DVDD.n3814 0.00182
R53201 DVDD.n3411 DVDD.n3397 0.00182
R53202 DVDD.n15669 DVDD.n3287 0.00182
R53203 DVDD.n15509 DVDD.n3194 0.00182
R53204 DVDD.n15998 DVDD.n3082 0.00182
R53205 DVDD.n15556 DVDD.n2651 0.00181707
R53206 DVDD.n15555 DVDD.n2578 0.00181707
R53207 DVDD.n15559 DVDD.n3242 0.00181707
R53208 DVDD.n15561 DVDD.n5124 0.00181707
R53209 DVDD.n3585 DVDD.n3554 0.00179
R53210 DVDD.n15738 DVDD.n4901 0.00179
R53211 DVDD.n5098 DVDD.n5043 0.00179
R53212 DVDD.n15447 DVDD.n5257 0.00179
R53213 DVDD.n15336 DVDD.n5372 0.00179
R53214 DVDD.n20191 DVDD.n19736 0.00178571
R53215 DVDD.n20266 DVDD.n19939 0.00178571
R53216 DVDD.n20683 DVDD.n18843 0.00178571
R53217 DVDD.n20758 DVDD.n19049 0.00178571
R53218 DVDD.n4056 DVDD.n3872 0.00178571
R53219 DVDD.n329 DVDD.n300 0.00178571
R53220 DVDD.n9820 DVDD.n9768 0.00178571
R53221 DVDD.n9704 DVDD.n9690 0.00178571
R53222 DVDD.n18711 DVDD.n18679 0.00178571
R53223 DVDD.n21126 DVDD.n100 0.00178571
R53224 DVDD.n4161 DVDD.n4160 0.00176
R53225 DVDD.n4639 DVDD.n4219 0.00176
R53226 DVDD.n15826 DVDD.n3402 0.00176
R53227 DVDD.n2503 DVDD.n2479 0.00176
R53228 DVDD.n3305 DVDD.n3291 0.00176
R53229 DVDD.n16293 DVDD.n2625 0.00176
R53230 DVDD.n15923 DVDD.n3198 0.00176
R53231 DVDD.n2855 DVDD.n2827 0.00176
R53232 DVDD.n3217 DVDD.n3086 0.00176
R53233 DVDD.n2984 DVDD.n2968 0.00176
R53234 DVDD.n21786 DVDD.n21785 0.00174867
R53235 DVDD.n18481 DVDD.n133 0.00174867
R53236 DVDD.n21896 DVDD.n21795 0.00174867
R53237 DVDD.n18107 DVDD.n18106 0.00174867
R53238 DVDD.n4752 DVDD.n4751 0.0017375
R53239 DVDD.n4399 DVDD.n4398 0.0017375
R53240 DVDD.n5512 DVDD.n5495 0.00173158
R53241 DVDD.n813 DVDD.n801 0.00173158
R53242 DVDD.n10067 DVDD.n9687 0.00172927
R53243 DVDD.n10056 DVDD.n9954 0.00172927
R53244 DVDD.n10092 DVDD.n9612 0.00172927
R53245 DVDD.n9950 DVDD.n9949 0.00172927
R53246 DVDD.n4157 DVDD.n4156 0.0017
R53247 DVDD.n4516 DVDD.n4505 0.0017
R53248 DVDD.n4659 DVDD.n4228 0.0017
R53249 DVDD.n4699 DVDD.n4199 0.0017
R53250 DVDD.n4861 DVDD.n3542 0.0017
R53251 DVDD.n4155 DVDD.n3760 0.0017
R53252 DVDD.n15993 DVDD.n3147 0.0017
R53253 DVDD.n15914 DVDD.n15913 0.0017
R53254 DVDD.n15912 DVDD.n3232 0.0017
R53255 DVDD.n15815 DVDD.n3231 0.0017
R53256 DVDD.n15814 DVDD.n15813 0.0017
R53257 DVDD.n16390 DVDD.n2349 0.0017
R53258 DVDD.n16368 DVDD.n2483 0.0017
R53259 DVDD.n3282 DVDD.n3148 0.0017
R53260 DVDD.n16271 DVDD.n2644 0.0017
R53261 DVDD.n16314 DVDD.n2571 0.0017
R53262 DVDD.n15990 DVDD.n3149 0.0017
R53263 DVDD.n2767 DVDD.n2746 0.0017
R53264 DVDD.n16246 DVDD.n2832 0.0017
R53265 DVDD.n15992 DVDD.n15991 0.0017
R53266 DVDD.n16145 DVDD.n2995 0.0017
R53267 DVDD.n16185 DVDD.n16184 0.0017
R53268 DVDD.n21645 DVDD.n21644 0.00168421
R53269 DVDD.n21597 DVDD.n21596 0.00168421
R53270 DVDD.n19554 DVDD.n19552 0.00168421
R53271 DVDD.n19505 DVDD.n19504 0.00168421
R53272 DVDD.n18086 DVDD.n18062 0.00168125
R53273 DVDD.n22223 DVDD.n160 0.00167
R53274 DVDD.n21760 DVDD.n176 0.00167
R53275 DVDD.n18239 DVDD.n18231 0.00167
R53276 DVDD.n18555 DVDD.n18509 0.00167
R53277 DVDD.n21706 DVDD.n18518 0.00167
R53278 DVDD.n22033 DVDD.n21986 0.00167
R53279 DVDD.n21339 DVDD.n18548 0.00167
R53280 DVDD.n21670 DVDD.n21669 0.00167
R53281 DVDD.n21989 DVDD.n225 0.00167
R53282 DVDD.n21585 DVDD.n164 0.00167
R53283 DVDD.n18402 DVDD.n18400 0.00167
R53284 DVDD.n22051 DVDD.n18224 0.00167
R53285 DVDD.n480 DVDD.n450 0.00167
R53286 DVDD.n2549 DVDD.n506 0.00167
R53287 DVDD.n16345 DVDD.n557 0.00167
R53288 DVDD.n16224 DVDD.n644 0.00167
R53289 DVDD.n2905 DVDD.n734 0.00167
R53290 DVDD.n18114 DVDD 0.00165261
R53291 DVDD DVDD.n18092 0.00165261
R53292 DVDD.n4124 DVDD.n4081 0.00164
R53293 DVDD.n4492 DVDD.n4195 0.00164
R53294 DVDD.n15781 DVDD.n3483 0.00164
R53295 DVDD.n15865 DVDD.n2338 0.00164
R53296 DVDD.n15644 DVDD.n15602 0.00164
R53297 DVDD.n15886 DVDD.n2688 0.00164
R53298 DVDD.n15490 DVDD.n5132 0.00164
R53299 DVDD.n15966 DVDD.n2749 0.00164
R53300 DVDD.n15374 DVDD.n3111 0.00164
R53301 DVDD.n16125 DVDD.n3029 0.00164
R53302 DVDD.n4987 DVDD.n3520 0.00163684
R53303 DVDD.n5000 DVDD.n4987 0.00163684
R53304 DVDD.n4997 DVDD.n4992 0.00163684
R53305 DVDD.n5003 DVDD.n4885 0.00163684
R53306 DVDD.n5305 DVDD.n5055 0.00163684
R53307 DVDD.n15699 DVDD.n5077 0.00163684
R53308 DVDD.n5337 DVDD.n5246 0.00163684
R53309 DVDD.n5343 DVDD.n5235 0.00163684
R53310 DVDD.n5395 DVDD.n5376 0.00163684
R53311 DVDD.n15147 DVDD.n5563 0.00163684
R53312 DVDD.n5566 DVDD.n5564 0.00163684
R53313 DVDD.n15144 DVDD.n15143 0.00163684
R53314 DVDD.n18037 DVDD.n18036 0.00163684
R53315 DVDD.n18036 DVDD.n543 0.00163684
R53316 DVDD.n18032 DVDD.n546 0.00163684
R53317 DVDD.n18023 DVDD.n521 0.00163684
R53318 DVDD.n594 DVDD.n570 0.00163684
R53319 DVDD.n17972 DVDD.n582 0.00163684
R53320 DVDD.n699 DVDD.n677 0.00163684
R53321 DVDD.n705 DVDD.n665 0.00163684
R53322 DVDD.n747 DVDD.n738 0.00163684
R53323 DVDD.n17737 DVDD.n880 0.00163684
R53324 DVDD.n886 DVDD.n884 0.00163684
R53325 DVDD.n17734 DVDD.n17731 0.00163684
R53326 DVDD.n21856 DVDD.n21855 0.001625
R53327 DVDD.n18279 DVDD.n18273 0.001625
R53328 DVDD.n21245 DVDD.n21219 0.001625
R53329 DVDD.n21959 DVDD.n21958 0.001625
R53330 DVDD.n21817 DVDD.n21813 0.001625
R53331 DVDD.n18465 DVDD.n18463 0.001625
R53332 DVDD.n4760 DVDD.n3654 0.001625
R53333 DVDD.n4307 DVDD.n4305 0.001625
R53334 DVDD.n3700 DVDD.n3699 0.001625
R53335 DVDD.n4544 DVDD.n4391 0.001625
R53336 DVDD.n14274 DVDD.n14273 0.001625
R53337 DVDD.n15142 DVDD.n15141 0.00158271
R53338 DVDD.n13782 DVDD.n13781 0.00158271
R53339 DVDD.n13274 DVDD.n13273 0.00158271
R53340 DVDD.n4110 DVDD.n4085 0.00158
R53341 DVDD.n15765 DVDD.n3487 0.00158
R53342 DVDD.n15680 DVDD.n15535 0.00158
R53343 DVDD.n15474 DVDD.n5136 0.00158
R53344 DVDD.n15388 DVDD.n3115 0.00158
R53345 DVDD.n20186 DVDD.n19735 0.00152857
R53346 DVDD.n20262 DVDD.n19938 0.00152857
R53347 DVDD.n20678 DVDD.n18842 0.00152857
R53348 DVDD.n19064 DVDD.n19048 0.00152857
R53349 DVDD.n4063 DVDD.n4062 0.00152857
R53350 DVDD.n335 DVDD.n323 0.00152857
R53351 DVDD.n9884 DVDD.n9767 0.00152857
R53352 DVDD.n9707 DVDD.n9689 0.00152857
R53353 DVDD.n18709 DVDD.n18700 0.00152857
R53354 DVDD.n21144 DVDD.n99 0.00152857
R53355 DVDD.n4116 DVDD.n4083 0.00152
R53356 DVDD.n4494 DVDD.n4190 0.00152
R53357 DVDD.n15772 DVDD.n3485 0.00152
R53358 DVDD.n15856 DVDD.n2340 0.00152
R53359 DVDD.n15635 DVDD.n15604 0.00152
R53360 DVDD.n15894 DVDD.n2690 0.00152
R53361 DVDD.n15481 DVDD.n5134 0.00152
R53362 DVDD.n15974 DVDD.n2751 0.00152
R53363 DVDD.n15382 DVDD.n3113 0.00152
R53364 DVDD.n16116 DVDD.n3031 0.00152
R53365 DVDD.n484 DVDD.n452 0.00149
R53366 DVDD.n2557 DVDD.n508 0.00149
R53367 DVDD.n16353 DVDD.n555 0.00149
R53368 DVDD.n16232 DVDD.n642 0.00149
R53369 DVDD.n2913 DVDD.n736 0.00149
R53370 DVDD.n14271 DVDD.n10595 0.00148253
R53371 DVDD.n14272 DVDD.n10593 0.00148253
R53372 DVDD.n13779 DVDD.n11582 0.00146644
R53373 DVDD.n12908 DVDD.n12900 0.00146644
R53374 DVDD.n13780 DVDD.n11583 0.00146644
R53375 DVDD.n12906 DVDD.n12902 0.00146644
R53376 DVDD.n3434 DVDD.n2361 0.00146585
R53377 DVDD.n15565 DVDD.n2649 0.00146585
R53378 DVDD.n3433 DVDD.n2485 0.00146585
R53379 DVDD.n15564 DVDD.n2576 0.00146585
R53380 DVDD.n3437 DVDD.n3260 0.00146585
R53381 DVDD.n15568 DVDD.n3240 0.00146585
R53382 DVDD.n3439 DVDD.n3431 0.00146585
R53383 DVDD.n15570 DVDD.n5122 0.00146585
R53384 DVDD.n20353 DVDD.n18940 0.00146429
R53385 DVDD.n20834 DVDD.n18968 0.00146429
R53386 DVDD.n22093 DVDD.n22076 0.00146429
R53387 DVDD.n10036 DVDD.n798 0.00146429
R53388 DVDD.n22327 DVDD.n25 0.00146429
R53389 DVDD.n4132 DVDD.n4079 0.00146
R53390 DVDD.n4534 DVDD.n4462 0.00146
R53391 DVDD.n4782 DVDD.n4781 0.00146
R53392 DVDD.n4202 DVDD.n4198 0.00146
R53393 DVDD.n15757 DVDD.n15756 0.00146
R53394 DVDD.n5109 DVDD.n3507 0.00146
R53395 DVDD.n15466 DVDD.n15465 0.00146
R53396 DVDD.n15347 DVDD.n5226 0.00146
R53397 DVDD.n16134 DVDD.n16133 0.00146
R53398 DVDD.n15961 DVDD.n2708 0.00146
R53399 DVDD.n15881 DVDD.n15879 0.00146
R53400 DVDD.n15878 DVDD.n15873 0.00146
R53401 DVDD.n15789 DVDD.n3481 0.00146
R53402 DVDD.n15872 DVDD.n2336 0.00146
R53403 DVDD.n15651 DVDD.n15600 0.00146
R53404 DVDD.n15880 DVDD.n2686 0.00146
R53405 DVDD.n15520 DVDD.n5208 0.00146
R53406 DVDD.n15960 DVDD.n2710 0.00146
R53407 DVDD.n15368 DVDD.n3109 0.00146
R53408 DVDD.n16132 DVDD.n3027 0.00146
R53409 DVDD.n5013 DVDD.n4887 0.00144737
R53410 DVDD.n15701 DVDD.n5047 0.00144737
R53411 DVDD.n5295 DVDD.n5057 0.00144737
R53412 DVDD.n5327 DVDD.n5244 0.00144737
R53413 DVDD.n5353 DVDD.n5233 0.00144737
R53414 DVDD.n5419 DVDD.n5397 0.00144737
R53415 DVDD.n5454 DVDD.n5405 0.00144737
R53416 DVDD.n18012 DVDD.n523 0.00144737
R53417 DVDD.n17980 DVDD.n552 0.00144737
R53418 DVDD.n627 DVDD.n578 0.00144737
R53419 DVDD.n689 DVDD.n663 0.00144737
R53420 DVDD.n715 DVDD.n679 0.00144737
R53421 DVDD.n17945 DVDD.n749 0.00144737
R53422 DVDD.n17910 DVDD.n757 0.00144737
R53423 DVDD.n18499 DVDD.n18457 0.00143
R53424 DVDD.n21880 DVDD.n21879 0.00143
R53425 DVDD.n21830 DVDD.n21799 0.00143
R53426 DVDD.n21254 DVDD.n18664 0.00143
R53427 DVDD.n21949 DVDD.n18295 0.00143
R53428 DVDD.n21978 DVDD.n205 0.00143
R53429 DVDD.n21223 DVDD.n18661 0.00143
R53430 DVDD.n18306 DVDD.n18294 0.00143
R53431 DVDD.n18352 DVDD.n18351 0.00143
R53432 DVDD.n18493 DVDD.n18460 0.00143
R53433 DVDD.n21867 DVDD.n21841 0.00143
R53434 DVDD.n21913 DVDD.n21802 0.00143
R53435 DVDD.n476 DVDD.n448 0.00143
R53436 DVDD.n2543 DVDD.n504 0.00143
R53437 DVDD.n16339 DVDD.n559 0.00143
R53438 DVDD.n16218 DVDD.n646 0.00143
R53439 DVDD.n2899 DVDD.n732 0.00143
R53440 DVDD.n20202 DVDD.n19739 0.0014
R53441 DVDD.n19944 DVDD.n19943 0.0014
R53442 DVDD.n20694 DVDD.n18846 0.0014
R53443 DVDD.n20769 DVDD.n19053 0.0014
R53444 DVDD.n4045 DVDD.n3875 0.0014
R53445 DVDD.n22156 DVDD.n22155 0.0014
R53446 DVDD.n4766 DVDD.n3653 0.0014
R53447 DVDD.n4177 DVDD.n4176 0.0014
R53448 DVDD.n4643 DVDD.n4224 0.0014
R53449 DVDD.n4586 DVDD.n493 0.0014
R53450 DVDD.n4548 DVDD.n4390 0.0014
R53451 DVDD.n15837 DVDD.n15836 0.0014
R53452 DVDD.n2512 DVDD.n2481 0.0014
R53453 DVDD.n3314 DVDD.n3294 0.0014
R53454 DVDD.n16302 DVDD.n2628 0.0014
R53455 DVDD.n15940 DVDD.n3200 0.0014
R53456 DVDD.n2865 DVDD.n2830 0.0014
R53457 DVDD.n16086 DVDD.n3057 0.0014
R53458 DVDD.n2981 DVDD.n2971 0.0014
R53459 DVDD.n9937 DVDD.n9772 0.0014
R53460 DVDD.n9723 DVDD.n9694 0.0014
R53461 DVDD.n21196 DVDD.n18701 0.0014
R53462 DVDD.n21128 DVDD.n103 0.0014
R53463 DVDD.n3591 DVDD.n3556 0.00137
R53464 DVDD.n15730 DVDD.n4903 0.00137
R53465 DVDD.n15694 DVDD.n5045 0.00137
R53466 DVDD.n15439 DVDD.n5259 0.00137
R53467 DVDD.n15402 DVDD.n5370 0.00137
R53468 DVDD.n5502 DVDD.n5493 0.00135263
R53469 DVDD.n822 DVDD.n803 0.00135263
R53470 DVDD.n18114 DVDD.n18096 0.00134674
R53471 DVDD.n18074 DVDD.n18061 0.00134375
R53472 DVDD.n4158 DVDD.n3761 0.00134
R53473 DVDD.n4636 DVDD.n4215 0.00134
R53474 DVDD.n476 DVDD 0.00134
R53475 DVDD.n18158 DVDD 0.00134
R53476 DVDD DVDD.n2900 0.00134
R53477 DVDD DVDD.n16219 0.00134
R53478 DVDD DVDD.n16340 0.00134
R53479 DVDD DVDD.n2544 0.00134
R53480 DVDD.n15819 DVDD.n3400 0.00134
R53481 DVDD.n2496 DVDD.n2477 0.00134
R53482 DVDD.n2543 DVDD 0.00134
R53483 DVDD.n15910 DVDD.n3235 0.00134
R53484 DVDD.n2635 DVDD.n2623 0.00134
R53485 DVDD.n16339 DVDD 0.00134
R53486 DVDD.n15989 DVDD.n3162 0.00134
R53487 DVDD.n2848 DVDD.n2825 0.00134
R53488 DVDD.n16218 DVDD 0.00134
R53489 DVDD.n3223 DVDD.n3084 0.00134
R53490 DVDD.n16161 DVDD.n2966 0.00134
R53491 DVDD.n2899 DVDD 0.00134
R53492 DVDD.n3709 DVDD.n3677 0.00133742
R53493 DVDD.n20337 DVDD.n18944 0.00133571
R53494 DVDD.n20852 DVDD.n20851 0.00133571
R53495 DVDD.n22116 DVDD.n22115 0.00133571
R53496 DVDD.n10020 DVDD.n795 0.00133571
R53497 DVDD.n22 DVDD.n20 0.00133571
R53498 DVDD.n15136 DVDD.n5577 0.00131203
R53499 DVDD.n3580 DVDD.n3552 0.00131
R53500 DVDD.n15744 DVDD.n4899 0.00131
R53501 DVDD.n5091 DVDD.n5041 0.00131
R53502 DVDD.n15453 DVDD.n5255 0.00131
R53503 DVDD.n15329 DVDD.n5374 0.00131
R53504 DVDD.n4736 DVDD.n3758 0.0013
R53505 DVDD.n15817 DVDD.n15816 0.0013
R53506 DVDD.n15663 DVDD.n3227 0.0013
R53507 DVDD.n15916 DVDD.n15915 0.0013
R53508 DVDD.n3226 DVDD.n3146 0.0013
R53509 DVDD.n3711 DVDD.n3656 0.0012875
R53510 DVDD.n4478 DVDD.n4394 0.0012875
R53511 DVDD.n17310 DVDD.n907 0.00128471
R53512 DVDD.n17311 DVDD.n17310 0.00128471
R53513 DVDD.n3818 DVDD.n3812 0.00128
R53514 DVDD.n4633 DVDD.n4632 0.00128
R53515 DVDD.n15809 DVDD.n3394 0.00128
R53516 DVDD.n16374 DVDD.n2385 0.00128
R53517 DVDD.n15667 DVDD.n3284 0.00128
R53518 DVDD.n16280 DVDD.n2619 0.00128
R53519 DVDD.n15507 DVDD.n3192 0.00128
R53520 DVDD.n16249 DVDD.n16248 0.00128
R53521 DVDD.n15996 DVDD.n3079 0.00128
R53522 DVDD.n16154 DVDD.n2962 0.00128
R53523 DVDD.n20031 DVDD.n19971 0.00127143
R53524 DVDD.n19859 DVDD.n19836 0.00127143
R53525 DVDD.n19149 DVDD.n19134 0.00127143
R53526 DVDD.n20805 DVDD.n18880 0.00127143
R53527 DVDD.n22178 DVDD.n22177 0.00127143
R53528 DVDD.n393 DVDD.n374 0.00127143
R53529 DVDD.n9649 DVDD.n9648 0.00127143
R53530 DVDD.n9969 DVDD.n9751 0.00127143
R53531 DVDD.n21114 DVDD.n21094 0.00127143
R53532 DVDD.n22273 DVDD.n73 0.00127143
R53533 DVDD DVDD.n18068 0.00126841
R53534 DVDD.n5002 DVDD.n3519 0.00125789
R53535 DVDD.n5029 DVDD.n3513 0.00125789
R53536 DVDD.n5032 DVDD.n3512 0.00125789
R53537 DVDD.n5276 DVDD.n5069 0.00125789
R53538 DVDD.n5279 DVDD.n5070 0.00125789
R53539 DVDD.n15460 DVDD.n15415 0.00125789
R53540 DVDD.n5435 DVDD.n5388 0.00125789
R53541 DVDD.n5438 DVDD.n5387 0.00125789
R53542 DVDD.n18027 DVDD.n540 0.00125789
R53543 DVDD.n17996 DVDD.n534 0.00125789
R53544 DVDD.n17993 DVDD.n533 0.00125789
R53545 DVDD.n608 DVDD.n591 0.00125789
R53546 DVDD.n611 DVDD.n576 0.00125789
R53547 DVDD.n17962 DVDD.n17961 0.00125789
R53548 DVDD.n17929 DVDD.n767 0.00125789
R53549 DVDD.n17926 DVDD.n766 0.00125789
R53550 DVDD.n3586 DVDD.n3561 0.00125
R53551 DVDD.n15736 DVDD.n15710 0.00125
R53552 DVDD.n5100 DVDD.n5050 0.00125
R53553 DVDD.n15445 DVDD.n15419 0.00125
R53554 DVDD.n15338 DVDD.n5380 0.00125
R53555 DVDD.n3808 DVDD.n3766 0.00122
R53556 DVDD.n4628 DVDD.n4220 0.00122
R53557 DVDD.n18134 DVDD.n487 0.00122
R53558 DVDD.n4662 DVDD.n490 0.00122
R53559 DVDD.n16199 DVDD.n2882 0.00122
R53560 DVDD.n16242 DVDD.n16240 0.00122
R53561 DVDD.n16318 DVDD.n2527 0.00122
R53562 DVDD.n16364 DVDD.n2523 0.00122
R53563 DVDD.n15828 DVDD.n3390 0.00122
R53564 DVDD.n2505 DVDD.n2434 0.00122
R53565 DVDD.n16363 DVDD.n16362 0.00122
R53566 DVDD.n3299 DVDD.n3280 0.00122
R53567 DVDD.n2632 DVDD.n2615 0.00122
R53568 DVDD.n16361 DVDD.n2526 0.00122
R53569 DVDD.n3205 DVDD.n3188 0.00122
R53570 DVDD.n2857 DVDD.n2819 0.00122
R53571 DVDD.n16241 DVDD.n2525 0.00122
R53572 DVDD.n3215 DVDD.n3075 0.00122
R53573 DVDD.n16170 DVDD.n2958 0.00122
R53574 DVDD.n16195 DVDD.n16194 0.00122
R53575 DVDD.n21370 DVDD.n18533 0.00121053
R53576 DVDD.n18428 DVDD.n18392 0.00121053
R53577 DVDD.n20156 DVDD.n20129 0.00120714
R53578 DVDD.n20648 DVDD.n20616 0.00120714
R53579 DVDD.n3949 DVDD.n3929 0.00120714
R53580 DVDD.n9855 DVDD.n5480 0.00120714
R53581 DVDD.n19665 DVDD.n19199 0.00120714
R53582 DVDD.n16396 DVDD.n2325 0.00120244
R53583 DVDD.n4352 DVDD.n4351 0.00120244
R53584 DVDD.n16369 DVDD.n2475 0.00120244
R53585 DVDD.n15838 DVDD.n3396 0.00120244
R53586 DVDD.n15794 DVDD.n3488 0.00120244
R53587 DVDD.n21887 DVDD.n21789 0.00119
R53588 DVDD.n21888 DVDD.n21790 0.00119
R53589 DVDD.n21963 DVDD.n200 0.00119
R53590 DVDD.n21966 DVDD.n18282 0.00119
R53591 DVDD.n18363 DVDD.n18362 0.00119
R53592 DVDD.n18317 DVDD.n18281 0.00119
R53593 DVDD.n21859 DVDD.n21808 0.00119
R53594 DVDD.n21903 DVDD.n21902 0.00119
R53595 DVDD.n18422 DVDD.n18421 0.001175
R53596 DVDD.n22021 DVDD.n22011 0.001175
R53597 DVDD.n21346 DVDD.n21345 0.001175
R53598 DVDD.n21695 DVDD.n18524 0.001175
R53599 DVDD.n18256 DVDD.n18218 0.001175
R53600 DVDD.n18440 DVDD.n18439 0.001175
R53601 DVDD.n4442 DVDD.n4441 0.001175
R53602 DVDD.n4252 DVDD.n4240 0.001175
R53603 DVDD.n4288 DVDD.n4287 0.001175
R53604 DVDD.n3684 DVDD.n3681 0.001175
R53605 DVDD.n15084 DVDD.n7051 0.001175
R53606 DVDD.n21941 DVDD 0.00117236
R53607 DVDD.n5499 DVDD.n5492 0.00116316
R53608 DVDD.n819 DVDD.n802 0.00116316
R53609 DVDD.n4137 DVDD.n3823 0.00116
R53610 DVDD.n4504 DVDD.n4205 0.00116
R53611 DVDD.n15795 DVDD.n3415 0.00116
R53612 DVDD.n16381 DVDD.n2348 0.00116
R53613 DVDD.n15678 DVDD.n15677 0.00116
R53614 DVDD.n16268 DVDD.n16267 0.00116
R53615 DVDD.n15528 DVDD.n5159 0.00116
R53616 DVDD.n2772 DVDD.n2766 0.00116
R53617 DVDD.n16067 DVDD.n16006 0.00116
R53618 DVDD.n16142 DVDD.n16141 0.00116
R53619 DVDD.n21595 DVDD.n18409 0.00115854
R53620 DVDD.n21737 DVDD.n18410 0.00115854
R53621 DVDD.n21647 DVDD.n21646 0.00115854
R53622 DVDD.n21441 DVDD.n18530 0.00115854
R53623 DVDD.n20221 DVDD.n19975 0.00114286
R53624 DVDD.n20299 DVDD.n19840 0.00114286
R53625 DVDD.n20713 DVDD.n19138 0.00114286
R53626 DVDD.n20789 DVDD.n18886 0.00114286
R53627 DVDD.n4027 DVDD.n241 0.00114286
R53628 DVDD.n402 DVDD.n378 0.00114286
R53629 DVDD.n9918 DVDD.n9641 0.00114286
R53630 DVDD.n9978 DVDD.n9755 0.00114286
R53631 DVDD.n21102 DVDD.n21099 0.00114286
R53632 DVDD.n81 DVDD.n78 0.00114286
R53633 DVDD.n4700 DVDD.n4699 0.00114
R53634 DVDD.n15871 DVDD.n2703 0.00114
R53635 DVDD.n16262 DVDD.n2704 0.00114
R53636 DVDD.n16261 DVDD.n2706 0.00114
R53637 DVDD.n16131 DVDD.n2705 0.00114
R53638 DVDD.n22222 DVDD.n166 0.00113
R53639 DVDD.n21763 DVDD.n18395 0.00113
R53640 DVDD.n22061 DVDD.n18213 0.00113
R53641 DVDD.n21652 DVDD.n18510 0.00113
R53642 DVDD.n21692 DVDD.n18528 0.00113
R53643 DVDD.n22032 DVDD.n22024 0.00113
R53644 DVDD.n21655 DVDD.n21654 0.00113
R53645 DVDD.n18540 DVDD.n18527 0.00113
R53646 DVDD.n22009 DVDD.n226 0.00113
R53647 DVDD.n21592 DVDD.n21590 0.00113
R53648 DVDD.n21749 DVDD.n18398 0.00113
R53649 DVDD.n22052 DVDD.n18217 0.00113
R53650 DVDD.n478 DVDD.n457 0.00113
R53651 DVDD.n2551 DVDD.n513 0.00113
R53652 DVDD.n16347 DVDD.n566 0.00113
R53653 DVDD.n16226 DVDD.n653 0.00113
R53654 DVDD.n2907 DVDD.n742 0.00113
R53655 DVDD.n3609 DVDD.n3529 0.00111875
R53656 DVDD.n3445 DVDD.n2357 0.00111463
R53657 DVDD.n15574 DVDD.n2647 0.00111463
R53658 DVDD.n3444 DVDD.n2399 0.00111463
R53659 DVDD.n15573 DVDD.n2574 0.00111463
R53660 DVDD.n3448 DVDD.n3357 0.00111463
R53661 DVDD.n15577 DVDD.n3238 0.00111463
R53662 DVDD.n3450 DVDD.n3429 0.00111463
R53663 DVDD.n15579 DVDD.n5120 0.00111463
R53664 DVDD.n4097 DVDD.n4090 0.0011
R53665 DVDD.n4500 DVDD.n4499 0.0011
R53666 DVDD.n15779 DVDD.n3493 0.0011
R53667 DVDD.n15863 DVDD.n2344 0.0011
R53668 DVDD.n15642 DVDD.n15614 0.0011
R53669 DVDD.n15888 DVDD.n2696 0.0011
R53670 DVDD.n5217 DVDD.n5140 0.0011
R53671 DVDD.n15968 DVDD.n2755 0.0011
R53672 DVDD.n15376 DVDD.n3119 0.0011
R53673 DVDD.n16123 DVDD.n3036 0.0011
R53674 DVDD.n7045 DVDD.n6795 0.00108952
R53675 DVDD.n15086 DVDD.n15085 0.00108952
R53676 DVDD.n20138 DVDD.n20077 0.00107857
R53677 DVDD.n20136 DVDD.n20124 0.00107857
R53678 DVDD.n20625 DVDD.n20608 0.00107857
R53679 DVDD.n20623 DVDD.n20611 0.00107857
R53680 DVDD.n3975 DVDD.n3940 0.00107857
R53681 DVDD.n3972 DVDD.n3965 0.00107857
R53682 DVDD.n5491 DVDD.n5469 0.00107857
R53683 DVDD.n9838 DVDD.n5485 0.00107857
R53684 DVDD.n19648 DVDD.n19193 0.00107857
R53685 DVDD.n19646 DVDD.n19195 0.00107857
R53686 DVDD.n5988 DVDD.n5934 0.00106946
R53687 DVDD.n9560 DVDD.n9222 0.00106946
R53688 DVDD.n10231 DVDD.n10230 0.00106946
R53689 DVDD.n17280 DVDD.n1264 0.00106946
R53690 DVDD.n5017 DVDD.n4888 0.00106842
R53691 DVDD.n5264 DVDD.n5064 0.00106842
R53692 DVDD.n5292 DVDD.n5058 0.00106842
R53693 DVDD.n5324 DVDD.n5243 0.00106842
R53694 DVDD.n5357 DVDD.n5232 0.00106842
R53695 DVDD.n5423 DVDD.n5398 0.00106842
R53696 DVDD.n5451 DVDD.n5404 0.00106842
R53697 DVDD.n18009 DVDD.n524 0.00106842
R53698 DVDD.n596 DVDD.n574 0.00106842
R53699 DVDD.n624 DVDD.n571 0.00106842
R53700 DVDD.n686 DVDD.n676 0.00106842
R53701 DVDD.n719 DVDD.n666 0.00106842
R53702 DVDD.n17942 DVDD.n750 0.00106842
R53703 DVDD.n17914 DVDD.n756 0.00106842
R53704 DVDD.n6403 DVDD.n6402 0.00106487
R53705 DVDD.n13269 DVDD.n13268 0.00106487
R53706 DVDD.n3817 DVDD.n3752 0.0010625
R53707 DVDD.n4573 DVDD.n4243 0.0010625
R53708 DVDD.n18157 DVDD 0.00106
R53709 DVDD.n2538 DVDD 0.00106
R53710 DVDD.n16211 DVDD 0.00106
R53711 DVDD.n2894 DVDD 0.00106
R53712 DVDD.n13765 DVDD.n11925 0.0010465
R53713 DVDD.n10699 DVDD.n10686 0.00104135
R53714 DVDD.n17010 DVDD.n1702 0.00104135
R53715 DVDD.n10233 DVDD.n10232 0.00103731
R53716 DVDD.n11568 DVDD.n11103 0.00103731
R53717 DVDD.n5986 DVDD.n5642 0.00103272
R53718 DVDD.n5987 DVDD.n5593 0.00103272
R53719 DVDD.n5938 DVDD.n5740 0.00103272
R53720 DVDD.n5991 DVDD.n5592 0.00103272
R53721 DVDD.n10692 DVDD.n10690 0.00102813
R53722 DVDD.n14000 DVDD.n11149 0.00102813
R53723 DVDD.n18367 DVDD.n18366 0.00102144
R53724 DVDD.n21269 DVDD.n18657 0.00102144
R53725 DVDD.n18342 DVDD.n18341 0.00102144
R53726 DVDD.n3537 DVDD.n3532 0.00102144
R53727 DVDD.n14303 DVDD.n14302 0.00101894
R53728 DVDD.n11573 DVDD.n11227 0.00101894
R53729 DVDD.n20038 DVDD.n20025 0.00101429
R53730 DVDD.n19865 DVDD.n19843 0.00101429
R53731 DVDD.n19160 DVDD.n19143 0.00101429
R53732 DVDD.n18893 DVDD.n18872 0.00101429
R53733 DVDD.n4029 DVDD.n245 0.00101429
R53734 DVDD.n380 DVDD.n360 0.00101429
R53735 DVDD.n9920 DVDD.n9642 0.00101429
R53736 DVDD.n9956 DVDD.n9738 0.00101429
R53737 DVDD.n21183 DVDD.n18737 0.00101429
R53738 DVDD.n22296 DVDD.n58 0.00101429
R53739 DVDD.n8145 DVDD.n8143 0.00100976
R53740 DVDD.n13487 DVDD.n12432 0.00100517
R53741 DVDD.n12737 DVDD.n12736 0.00100057
R53742 DVDD.n15079 DVDD.n7056 0.000991389
R53743 DVDD.n9559 DVDD.n9558 0.000991389
R53744 DVDD.n16735 DVDD.n1805 0.000991389
R53745 DVDD.n10704 DVDD.n10703 0.000983221
R53746 DVDD.n17008 DVDD.n17006 0.000983221
R53747 DVDD.n14020 DVDD.n10687 0.000983221
R53748 DVDD.n17012 DVDD.n17011 0.000983221
R53749 DVDD.n7412 DVDD.n7411 0.000982204
R53750 DVDD.n17004 DVDD.n1706 0.000982204
R53751 DVDD.n21934 DVDD.n21933 0.000980256
R53752 DVDD.n22237 DVDD.n131 0.000980256
R53753 DVDD.n21928 DVDD.n21793 0.000980256
R53754 DVDD.n18105 DVDD.n18104 0.000980256
R53755 DVDD.n4118 DVDD.n4089 0.00098
R53756 DVDD.n4498 DVDD.n4191 0.00098
R53757 DVDD.n4663 DVDD.n493 0.00098
R53758 DVDD.n2567 DVDD.n2522 0.00098
R53759 DVDD.n16320 DVDD.n16319 0.00098
R53760 DVDD.n2881 DVDD.n2568 0.00098
R53761 DVDD.n16190 DVDD.n16189 0.00098
R53762 DVDD.n15774 DVDD.n3492 0.00098
R53763 DVDD.n15858 DVDD.n2343 0.00098
R53764 DVDD.n15626 DVDD.n15613 0.00098
R53765 DVDD.n15892 DVDD.n2695 0.00098
R53766 DVDD.n15483 DVDD.n5139 0.00098
R53767 DVDD.n15972 DVDD.n2754 0.00098
R53768 DVDD.n15380 DVDD.n3118 0.00098
R53769 DVDD.n16118 DVDD.n3035 0.00098
R53770 DVDD.n14860 DVDD.n7615 0.000977612
R53771 DVDD.n5514 DVDD.n5487 0.000973684
R53772 DVDD.n17876 DVDD.n17875 0.000973684
R53773 DVDD.n14850 DVDD.n14849 0.00097302
R53774 DVDD.n12390 DVDD.n12389 0.00097302
R53775 DVDD.n1757 DVDD.n1712 0.00097302
R53776 DVDD.n14569 DVDD.n8154 0.000963835
R53777 DVDD.n1263 DVDD.n1256 0.000959242
R53778 DVDD.n17289 DVDD.n915 0.000959242
R53779 DVDD.n14294 DVDD.n14293 0.00095465
R53780 DVDD.n14004 DVDD.n11061 0.00095465
R53781 DVDD.n20154 DVDD.n20073 0.00095
R53782 DVDD.n20641 DVDD.n20604 0.00095
R53783 DVDD.n21736 DVDD.n171 0.00095
R53784 DVDD.n18393 DVDD.n172 0.00095
R53785 DVDD.n21648 DVDD.n18513 0.00095
R53786 DVDD.n21687 DVDD.n18514 0.00095
R53787 DVDD.n21331 DVDD.n18544 0.00095
R53788 DVDD.n21685 DVDD.n18531 0.00095
R53789 DVDD.n21740 DVDD.n21738 0.00095
R53790 DVDD.n21739 DVDD.n18404 0.00095
R53791 DVDD.n3951 DVDD.n3924 0.00095
R53792 DVDD.n4740 DVDD.n3734 0.00095
R53793 DVDD.n18144 DVDD.n456 0.00095
R53794 DVDD.n4315 DVDD.n4249 0.00095
R53795 DVDD.n2555 DVDD.n512 0.00095
R53796 DVDD.n16351 DVDD.n567 0.00095
R53797 DVDD.n16230 DVDD.n654 0.00095
R53798 DVDD.n2911 DVDD.n741 0.00095
R53799 DVDD.n9853 DVDD.n5473 0.00095
R53800 DVDD.n19663 DVDD.n19189 0.00095
R53801 DVDD.n15102 DVDD.n15101 0.000945465
R53802 DVDD.n6697 DVDD.n6696 0.000940873
R53803 DVDD.n8601 DVDD.n8600 0.00093628
R53804 DVDD.n13800 DVDD.n11233 0.00093628
R53805 DVDD.n13484 DVDD.n12477 0.00093628
R53806 DVDD.n13754 DVDD.n11939 0.000927095
R53807 DVDD.n17272 DVDD.n1262 0.000922503
R53808 DVDD.n17710 DVDD.n17369 0.000922503
R53809 DVDD.n17366 DVDD.n17306 0.000922503
R53810 DVDD.n17364 DVDD.n17309 0.000922503
R53811 DVDD.n17367 DVDD.n17307 0.000922503
R53812 DVDD.n4135 DVDD.n4134 0.00092
R53813 DVDD.n4503 DVDD.n4203 0.00092
R53814 DVDD.n15793 DVDD.n15791 0.00092
R53815 DVDD.n15876 DVDD.n2347 0.00092
R53816 DVDD.n15653 DVDD.n15618 0.00092
R53817 DVDD.n2701 DVDD.n2700 0.00092
R53818 DVDD.n15519 DVDD.n5143 0.00092
R53819 DVDD.n16258 DVDD.n16257 0.00092
R53820 DVDD.n15366 DVDD.n3122 0.00092
R53821 DVDD.n16135 DVDD.n3040 0.00092
R53822 DVDD.n15070 DVDD.n7057 0.00091791
R53823 DVDD.n6706 DVDD.n6391 0.000908726
R53824 DVDD.n16705 DVDD.n16704 0.000908726
R53825 DVDD.n16715 DVDD.n1821 0.000908726
R53826 DVDD.n13473 DVDD.n12779 0.000904133
R53827 DVDD.n13267 DVDD.n2210 0.000904133
R53828 DVDD.n14864 DVDD.n14863 0.000894948
R53829 DVDD.n11052 DVDD 0.000894948
R53830 DVDD.n3607 DVDD.n3524 0.00089375
R53831 DVDD.n8030 DVDD.n8029 0.000890356
R53832 DVDD.n12388 DVDD.n12330 0.000890356
R53833 DVDD.n16994 DVDD.n1755 0.000890356
R53834 DVDD.n17300 DVDD.n17299 0.000890356
R53835 DVDD.n18483 DVDD.n18477 0.00089
R53836 DVDD.n21876 DVDD.n21838 0.00089
R53837 DVDD.n21898 DVDD.n21895 0.00089
R53838 DVDD.n21253 DVDD.n18666 0.00089
R53839 DVDD.n18284 DVDD.n198 0.00089
R53840 DVDD.n21976 DVDD.n204 0.00089
R53841 DVDD.n21233 DVDD.n21232 0.00089
R53842 DVDD.n18324 DVDD.n18323 0.00089
R53843 DVDD.n18330 DVDD.n18272 0.00089
R53844 DVDD.n18492 DVDD.n18485 0.00089
R53845 DVDD.n21860 DVDD.n21843 0.00089
R53846 DVDD.n21912 DVDD.n21804 0.00089
R53847 DVDD.n18159 DVDD.n460 0.00089
R53848 DVDD.n2541 DVDD.n516 0.00089
R53849 DVDD.n16337 DVDD.n564 0.00089
R53850 DVDD.n16216 DVDD.n651 0.00089
R53851 DVDD.n2897 DVDD.n745 0.00089
R53852 DVDD.n20234 DVDD.n20030 0.000885714
R53853 DVDD.n20312 DVDD.n19847 0.000885714
R53854 DVDD.n20726 DVDD.n19148 0.000885714
R53855 DVDD.n20803 DVDD.n18879 0.000885714
R53856 DVDD.n272 DVDD.n249 0.000885714
R53857 DVDD.n415 DVDD.n385 0.000885714
R53858 DVDD.n10091 DVDD.n10090 0.000885714
R53859 DVDD.n9991 DVDD.n9961 0.000885714
R53860 DVDD.n21167 DVDD.n18741 0.000885714
R53861 DVDD.n22280 DVDD.n62 0.000885714
R53862 DVDD.n4992 DVDD.n4884 0.000878947
R53863 DVDD.n4996 DVDD.n3519 0.000878947
R53864 DVDD.n5308 DVDD.n5076 0.000878947
R53865 DVDD.n5309 DVDD.n5054 0.000878947
R53866 DVDD.n5340 DVDD.n5236 0.000878947
R53867 DVDD.n5341 DVDD.n5247 0.000878947
R53868 DVDD.n15410 DVDD.n15409 0.000878947
R53869 DVDD.n546 DVDD.n520 0.000878947
R53870 DVDD.n18034 DVDD.n540 0.000878947
R53871 DVDD.n17977 DVDD.n17976 0.000878947
R53872 DVDD.n595 DVDD.n584 0.000878947
R53873 DVDD.n702 DVDD.n660 0.000878947
R53874 DVDD.n703 DVDD.n673 0.000878947
R53875 DVDD.n17956 DVDD.n17955 0.000878947
R53876 DVDD.n13257 DVDD.n12912 0.000876579
R53877 DVDD.n15113 DVDD.n15112 0.000871986
R53878 DVDD.n8089 DVDD.n8044 0.000871986
R53879 DVDD.n10583 DVDD.n10582 0.000871986
R53880 DVDD.n11216 DVDD.n11215 0.000871986
R53881 DVDD.n11938 DVDD.n11937 0.000862801
R53882 DVDD.n3807 DVDD.n3768 0.00086
R53883 DVDD.n4627 DVDD.n4223 0.00086
R53884 DVDD.n3405 DVDD.n3389 0.00086
R53885 DVDD.n2489 DVDD.n2433 0.00086
R53886 DVDD.n3312 DVDD.n3279 0.00086
R53887 DVDD.n16300 DVDD.n2614 0.00086
R53888 DVDD.n15938 DVDD.n15937 0.00086
R53889 DVDD.n2836 DVDD.n2818 0.00086
R53890 DVDD.n16081 DVDD.n16075 0.00086
R53891 DVDD.n16174 DVDD.n2957 0.00086
R53892 DVDD.n1658 DVDD.n1611 0.000858209
R53893 DVDD.n8599 DVDD.n8205 0.000853617
R53894 DVDD.n11580 DVDD.n11276 0.000853617
R53895 DVDD.n1813 DVDD.n1812 0.000844432
R53896 DVDD.n17718 DVDD.n17717 0.000844432
R53897 DVDD.n13764 DVDD.n11926 0.000839839
R53898 DVDD.n1654 DVDD.n1605 0.000839839
R53899 DVDD.n4425 DVDD.n3738 0.0008375
R53900 DVDD.n4280 DVDD.n4251 0.0008375
R53901 DVDD.n15122 DVDD.n15121 0.000835247
R53902 DVDD.n7410 DVDD.n7404 0.000835247
R53903 DVDD.n7569 DVDD.n7500 0.000835247
R53904 DVDD.n1656 DVDD.n1655 0.000835247
R53905 DVDD.n3590 DVDD.n3560 0.00083
R53906 DVDD.n15732 DVDD.n15709 0.00083
R53907 DVDD.n15698 DVDD.n15697 0.00083
R53908 DVDD.n15441 DVDD.n15418 0.00083
R53909 DVDD.n15406 DVDD.n15405 0.00083
R53910 DVDD.n15092 DVDD.n6707 0.000826062
R53911 DVDD.n15092 DVDD.n6749 0.000826062
R53912 DVDD.n15089 DVDD.n6794 0.000826062
R53913 DVDD.n16727 DVDD.n1811 0.000826062
R53914 DVDD.n10642 DVDD.n10597 0.00082147
R53915 DVDD.n13470 DVDD.n12825 0.00082147
R53916 DVDD.n18945 DVDD.n18930 0.000821429
R53917 DVDD.n18989 DVDD.n18973 0.000821429
R53918 DVDD.n22087 DVDD.n22086 0.000821429
R53919 DVDD.n10016 DVDD.n789 0.000821429
R53920 DVDD.n22345 DVDD.n22344 0.000821429
R53921 DVDD.n15121 DVDD.n5935 0.000816877
R53922 DVDD.n12921 DVDD.n12825 0.000816877
R53923 DVDD.n21682 DVDD.n21681 0.000812862
R53924 DVDD.n21368 DVDD.n21333 0.000812862
R53925 DVDD.n22006 DVDD.n21993 0.000812862
R53926 DVDD.n3550 DVDD.n3549 0.000812862
R53927 DVDD.n14841 DVDD.n7688 0.000807692
R53928 DVDD.n13745 DVDD.n12287 0.000807692
R53929 DVDD.n16714 DVDD.n2156 0.000807692
R53930 DVDD.n17718 DVDD.n906 0.000807692
R53931 DVDD.n15060 DVDD.n7454 0.0008031
R53932 DVDD.n4156 DVDD.n3811 0.0008
R53933 DVDD.n4631 DVDD.n4214 0.0008
R53934 DVDD.n15814 DVDD.n3393 0.0008
R53935 DVDD.n2476 DVDD.n2437 0.0008
R53936 DVDD.n3283 DVDD.n3282 0.0008
R53937 DVDD.n16284 DVDD.n2618 0.0008
R53938 DVDD.n3191 DVDD.n3149 0.0008
R53939 DVDD.n2846 DVDD.n2822 0.0008
R53940 DVDD.n15992 DVDD.n3078 0.0008
R53941 DVDD.n2987 DVDD.n2961 0.0008
R53942 DVDD.n13787 DVDD.n11580 0.000798507
R53943 DVDD.n13256 DVDD.n12901 0.000793915
R53944 DVDD.n6331 DVDD.n6051 0.000789323
R53945 DVDD.n14825 DVDD.n8087 0.000789323
R53946 DVDD.n14285 DVDD.n10241 0.000789323
R53947 DVDD.n14270 DVDD.n14269 0.000789323
R53948 DVDD.n14013 DVDD.n14012 0.000789323
R53949 DVDD.n21764 DVDD.n18391 0.000788154
R53950 DVDD.n21733 DVDD.n18429 0.000788154
R53951 DVDD.n18211 DVDD.n18206 0.000788154
R53952 DVDD.n18123 DVDD.n18122 0.000788154
R53953 DVDD.n15284 DVDD.n5496 0.000784211
R53954 DVDD.n814 DVDD.n808 0.000784211
R53955 DVDD.n10582 DVDD.n10241 0.000780138
R53956 DVDD.n17262 DVDD.n1656 0.000775545
R53957 DVDD.n14560 DVDD.n8162 0.000770953
R53958 DVDD.n13787 DVDD.n13786 0.000770953
R53959 DVDD.n13778 DVDD.n13777 0.000770953
R53960 DVDD.n4834 DVDD.n4803 0.00077
R53961 DVDD.n3579 DVDD.n3564 0.00077
R53962 DVDD.n15749 DVDD.n4896 0.00077
R53963 DVDD.n15746 DVDD.n15714 0.00077
R53964 DVDD.n5079 DVDD.n5065 0.00077
R53965 DVDD.n5089 DVDD.n5081 0.00077
R53966 DVDD.n15458 DVDD.n5254 0.00077
R53967 DVDD.n15455 DVDD.n15423 0.00077
R53968 DVDD.n15325 DVDD.n5408 0.00077
R53969 DVDD.n15327 DVDD.n15317 0.00077
R53970 DVDD.n22252 DVDD.n104 0.000763415
R53971 DVDD.n3456 DVDD.n2355 0.000763415
R53972 DVDD.n2692 DVDD.n2645 0.000763415
R53973 DVDD.n22298 DVDD.n66 0.000763415
R53974 DVDD.n3455 DVDD.n2397 0.000763415
R53975 DVDD.n2620 DVDD.n2572 0.000763415
R53976 DVDD.n21185 DVDD.n21083 0.000763415
R53977 DVDD.n3458 DVDD.n3355 0.000763415
R53978 DVDD.n3286 DVDD.n3236 0.000763415
R53979 DVDD.n21212 DVDD.n18703 0.000763415
R53980 DVDD.n3460 DVDD.n3427 0.000763415
R53981 DVDD.n15609 DVDD.n5118 0.000763415
R53982 DVDD.n8029 DVDD.n7688 0.000761768
R53983 DVDD.n14840 DVDD.n7730 0.000761768
R53984 DVDD.n14837 DVDD.n7775 0.000761768
R53985 DVDD.n17299 DVDD.n906 0.000761768
R53986 DVDD.n14826 DVDD.n14825 0.000757176
R53987 DVDD.n8162 DVDD.n8155 0.000757176
R53988 DVDD.n14284 DVDD.n10283 0.000757176
R53989 DVDD.n14281 DVDD.n10328 0.000757176
R53990 DVDD.n19740 DVDD.n19724 0.000757143
R53991 DVDD.n20281 DVDD.n19885 0.000757143
R53992 DVDD.n18865 DVDD.n18847 0.000757143
R53993 DVDD.n19054 DVDD.n19035 0.000757143
R53994 DVDD.n3894 DVDD.n3876 0.000757143
R53995 DVDD.n326 DVDD.n321 0.000757143
R53996 DVDD.n9773 DVDD.n9757 0.000757143
R53997 DVDD.n9725 DVDD.n9681 0.000757143
R53998 DVDD.n21194 DVDD.n18708 0.000757143
R53999 DVDD.n106 DVDD.n105 0.000757143
R54000 DVDD.n6051 DVDD.n5935 0.000752583
R54001 DVDD.n7458 DVDD.n7454 0.000752583
R54002 DVDD.n12921 DVDD.n12901 0.000752583
R54003 DVDD.n17263 DVDD.n1611 0.000752583
R54004 DVDD.n10693 DVDD.n10642 0.000747991
R54005 DVDD.n6707 DVDD.n6706 0.000743398
R54006 DVDD.n6752 DVDD.n6749 0.000743398
R54007 DVDD.n12333 DVDD.n12332 0.000743398
R54008 DVDD.n13745 DVDD.n13744 0.000743398
R54009 DVDD.n16715 DVDD.n16714 0.000743398
R54010 DVDD.n16727 DVDD.n16726 0.000743398
R54011 DVDD.n3820 DVDD.n3816 0.00074
R54012 DVDD.n4635 DVDD.n4213 0.00074
R54013 DVDD.n15811 DVDD.n3399 0.00074
R54014 DVDD.n16371 DVDD.n16370 0.00074
R54015 DVDD.n15665 DVDD.n3289 0.00074
R54016 DVDD.n16282 DVDD.n2622 0.00074
R54017 DVDD.n3229 DVDD.n3196 0.00074
R54018 DVDD.n2824 DVDD.n2792 0.00074
R54019 DVDD.n15994 DVDD.n3083 0.00074
R54020 DVDD.n16156 DVDD.n2965 0.00074
R54021 DVDD.n14269 DVDD.n10640 0.000738806
R54022 DVDD.n15122 DVDD.n5934 0.000734214
R54023 DVDD.n14864 DVDD.n7569 0.000734214
R54024 DVDD.n12783 DVDD.n12779 0.000734214
R54025 DVDD.n1655 DVDD.n1654 0.000734214
R54026 DVDD.n15069 DVDD.n7404 0.000729621
R54027 DVDD.n11936 DVDD.n11926 0.000729621
R54028 DVDD.n7733 DVDD.n7730 0.000725029
R54029 DVDD.n12332 DVDD.n11939 0.000725029
R54030 DVDD.n17717 DVDD.n907 0.000725029
R54031 DVDD.n4753 DVDD.n3663 0.000725
R54032 DVDD.n4475 DVDD.n4401 0.000725
R54033 DVDD.n15057 DVDD.n7500 0.000720436
R54034 DVDD.n19032 DVDD.n18868 0.000719512
R54035 DVDD.n19024 DVDD.n18869 0.000719512
R54036 DVDD.n20931 DVDD.n18871 0.000719512
R54037 DVDD.n20930 DVDD.n18870 0.000719512
R54038 DVDD.n19128 DVDD.n18866 0.000719512
R54039 DVDD.n19075 DVDD.n18867 0.000719512
R54040 DVDD.n18860 DVDD.n18848 0.000719512
R54041 DVDD.n20969 DVDD.n20968 0.000719512
R54042 DVDD.n8600 DVDD.n8599 0.000715844
R54043 DVDD.n3589 DVDD.n3555 0.00071
R54044 DVDD.n15734 DVDD.n4902 0.00071
R54045 DVDD.n5082 DVDD.n5078 0.00071
R54046 DVDD.n15443 DVDD.n5258 0.00071
R54047 DVDD.n15318 DVDD.n5407 0.00071
R54048 DVDD.n10286 DVDD.n10283 0.000706659
R54049 DVDD.n11053 DVDD.n11052 0.000706659
R54050 DVDD.n8146 DVDD.n8089 0.000697474
R54051 DVDD.n11215 DVDD.n11061 0.000697474
R54052 DVDD.n11588 DVDD.n11581 0.000692882
R54053 DVDD.n13777 DVDD.n11631 0.000692882
R54054 DVDD.n20330 DVDD.n18934 0.000692857
R54055 DVDD.n20836 DVDD.n18963 0.000692857
R54056 DVDD.n22095 DVDD.n22073 0.000692857
R54057 DVDD.n10011 DVDD.n787 0.000692857
R54058 DVDD.n22315 DVDD.n16 0.000692857
R54059 DVDD.n5016 DVDD.n3516 0.000689474
R54060 DVDD.n5263 DVDD.n5066 0.000689474
R54061 DVDD.n5293 DVDD.n5073 0.000689474
R54062 DVDD.n5325 DVDD.n5239 0.000689474
R54063 DVDD.n5356 DVDD.n5250 0.000689474
R54064 DVDD.n5422 DVDD.n5391 0.000689474
R54065 DVDD.n5452 DVDD.n5384 0.000689474
R54066 DVDD.n18010 DVDD.n537 0.000689474
R54067 DVDD.n17979 DVDD.n561 0.000689474
R54068 DVDD.n625 DVDD.n586 0.000689474
R54069 DVDD.n687 DVDD.n675 0.000689474
R54070 DVDD.n718 DVDD.n658 0.000689474
R54071 DVDD.n17943 DVDD.n770 0.000689474
R54072 DVDD.n17913 DVDD.n763 0.000689474
R54073 DVDD.n14569 DVDD.n14568 0.000688289
R54074 DVDD.n14281 DVDD.n10286 0.000688289
R54075 DVDD.n13786 DVDD.n11581 0.000688289
R54076 DVDD.n13778 DVDD.n11588 0.000688289
R54077 DVDD.n14013 DVDD.n10710 0.000683697
R54078 DVDD.n4163 DVDD.n3767 0.00068
R54079 DVDD.n4642 DVDD.n4640 0.00068
R54080 DVDD.n15830 DVDD.n3404 0.00068
R54081 DVDD.n2507 DVDD.n2480 0.00068
R54082 DVDD.n3310 DVDD.n3293 0.00068
R54083 DVDD.n16298 DVDD.n2627 0.00068
R54084 DVDD.n15928 DVDD.n3199 0.00068
R54085 DVDD.n2859 DVDD.n2829 0.00068
R54086 DVDD.n16083 DVDD.n3087 0.00068
R54087 DVDD.n16172 DVDD.n2970 0.00068
R54088 DVDD.n11053 DVDD.n10710 0.000679104
R54089 DVDD.n14012 DVDD.n10711 0.000679104
R54090 DVDD.n12389 DVDD.n12388 0.000679104
R54091 DVDD.n17300 DVDD.n17298 0.000679104
R54092 DVDD.n14559 DVDD.n8205 0.000674512
R54093 DVDD.n16995 DVDD.n16994 0.000674512
R54094 DVDD.n22349 DVDD 0.000671429
R54095 DVDD.n20341 DVDD 0.000671429
R54096 DVDD DVDD.n20848 0.000671429
R54097 DVDD.n22107 DVDD 0.000671429
R54098 DVDD.n10024 DVDD 0.000671429
R54099 DVDD.n15113 DVDD.n6000 0.00066992
R54100 DVDD.n15061 DVDD.n7412 0.00066992
R54101 DVDD.n13258 DVDD.n13257 0.00066992
R54102 DVDD.n17004 DVDD.n17003 0.00066992
R54103 DVDD.n18078 DVDD.n18057 0.00066875
R54104 DVDD.n14837 DVDD.n7733 0.000665327
R54105 DVDD.n2210 DVDD.n2165 0.000665327
R54106 DVDD.n15100 DVDD.n6391 0.000660735
R54107 DVDD.n7056 DVDD.n6794 0.000660735
R54108 DVDD.n8030 DVDD.n7679 0.000660735
R54109 DVDD.n2208 DVDD.n1821 0.000660735
R54110 DVDD.n1812 DVDD.n1805 0.000660735
R54111 DVDD.n13800 DVDD.n13799 0.000656142
R54112 DVDD.n15078 DVDD.n7057 0.00065155
R54113 DVDD.n7615 DVDD.n7611 0.00065155
R54114 DVDD.n13474 DVDD.n12737 0.00065155
R54115 DVDD.n17272 DVDD.n17271 0.00065155
R54116 DVDD.n18476 DVDD.n127 0.00065
R54117 DVDD.n21836 DVDD.n21788 0.00065
R54118 DVDD.n21899 DVDD.n21829 0.00065
R54119 DVDD.n21216 DVDD.n18670 0.00065
R54120 DVDD.n21961 DVDD.n199 0.00065
R54121 DVDD.n18270 DVDD.n203 0.00065
R54122 DVDD.n21224 DVDD.n21220 0.00065
R54123 DVDD.n18316 DVDD.n18286 0.00065
R54124 DVDD.n18339 DVDD.n18329 0.00065
R54125 DVDD.n18462 DVDD.n123 0.00065
R54126 DVDD.n21874 DVDD.n21873 0.00065
R54127 DVDD.n21815 DVDD.n21810 0.00065
R54128 DVDD.n18194 DVDD.n461 0.00065
R54129 DVDD.n18040 DVDD.n517 0.00065
R54130 DVDD.n16335 DVDD.n558 0.00065
R54131 DVDD.n16214 DVDD.n645 0.00065
R54132 DVDD.n746 DVDD.n731 0.00065
R54133 DVDD.n13755 DVDD.n11938 0.000646958
R54134 DVDD.n17710 DVDD.n17311 0.000646958
R54135 DVDD.n17369 DVDD.n17306 0.000646958
R54136 DVDD.n17366 DVDD.n17309 0.000646958
R54137 DVDD.n17364 DVDD.n17307 0.000646958
R54138 DVDD.n17367 DVDD.n17308 0.000646958
R54139 DVDD.n8143 DVDD.n7775 0.000642365
R54140 DVDD.n13755 DVDD.n13754 0.000642365
R54141 DVDD.n13484 DVDD.n12435 0.00063318
R54142 DVDD.n6696 DVDD.n6348 0.000628588
R54143 DVDD.n14303 DVDD.n8258 0.000628588
R54144 DVDD.n20048 DVDD.n19728 0.000628571
R54145 DVDD.n20264 DVDD.n19889 0.000628571
R54146 DVDD.n19170 DVDD.n18835 0.000628571
R54147 DVDD.n20756 DVDD.n19039 0.000628571
R54148 DVDD.n3900 DVDD.n3897 0.000628571
R54149 DVDD.n337 DVDD.n322 0.000628571
R54150 DVDD.n9886 DVDD.n9760 0.000628571
R54151 DVDD.n9709 DVDD.n9685 0.000628571
R54152 DVDD.n21211 DVDD.n21210 0.000628571
R54153 DVDD.n21142 DVDD.n110 0.000628571
R54154 DVDD.n14568 DVDD.n8155 0.000623995
R54155 DVDD.n14560 DVDD.n14559 0.000623995
R54156 DVDD.n10690 DVDD.n10328 0.000623995
R54157 DVDD.n11051 DVDD.n10640 0.000623995
R54158 DVDD.n4138 DVDD.n3827 0.00062
R54159 DVDD.n4528 DVDD.n4204 0.00062
R54160 DVDD.n15796 DVDD.n3419 0.00062
R54161 DVDD.n2378 DVDD.n2335 0.00062
R54162 DVDD.n15619 DVDD.n15593 0.00062
R54163 DVDD.n16266 DVDD.n2685 0.00062
R54164 DVDD.n5144 DVDD.n5129 0.00062
R54165 DVDD.n2765 DVDD.n2764 0.00062
R54166 DVDD.n16061 DVDD.n3123 0.00062
R54167 DVDD.n16140 DVDD.n3026 0.00062
R54168 DVDD.n3670 DVDD.n3667 0.0006125
R54169 DVDD.n4546 DVDD.n4405 0.0006125
R54170 DVDD.n6331 DVDD.n6000 0.000610218
R54171 DVDD.n15112 DVDD.n6043 0.000610218
R54172 DVDD.n14294 DVDD.n8609 0.000610218
R54173 DVDD.n10583 DVDD.n8610 0.000610218
R54174 DVDD.n8154 DVDD.n8087 0.000605626
R54175 DVDD.n14285 DVDD.n14284 0.000605626
R54176 DVDD.n11925 DVDD.n11631 0.000605626
R54177 DVDD.n13258 DVDD.n13256 0.000605626
R54178 DVDD.n13266 DVDD.n12912 0.000605626
R54179 DVDD.n11216 DVDD.n10711 0.000601033
R54180 DVDD.n12333 DVDD.n12287 0.000601033
R54181 DVDD.n15061 DVDD.n15060 0.000596441
R54182 DVDD.n15057 DVDD.n7458 0.000596441
R54183 DVDD.n14850 DVDD.n7678 0.000596441
R54184 DVDD.n13488 DVDD.n12390 0.000596441
R54185 DVDD.n16736 DVDD.n1757 0.000596441
R54186 DVDD.n17290 DVDD.n1256 0.000596441
R54187 DVDD.n17290 DVDD.n17289 0.000596441
R54188 DVDD.n5500 DVDD.n5490 0.000594737
R54189 DVDD.n820 DVDD.n810 0.000594737
R54190 DVDD.n21735 DVDD.n18425 0.00059
R54191 DVDD.n18394 DVDD.n173 0.00059
R54192 DVDD.n22058 DVDD.n18214 0.00059
R54193 DVDD.n21649 DVDD.n18554 0.00059
R54194 DVDD.n21688 DVDD.n18515 0.00059
R54195 DVDD.n22027 DVDD.n233 0.00059
R54196 DVDD.n21332 DVDD.n18550 0.00059
R54197 DVDD.n21662 DVDD.n18532 0.00059
R54198 DVDD.n21988 DVDD.n228 0.00059
R54199 DVDD.n21591 DVDD.n18408 0.00059
R54200 DVDD.n21753 DVDD.n21752 0.00059
R54201 DVDD.n22057 DVDD.n18219 0.00059
R54202 DVDD.n18146 DVDD.n451 0.00059
R54203 DVDD.n2553 DVDD.n507 0.00059
R54204 DVDD.n16349 DVDD.n556 0.00059
R54205 DVDD.n16228 DVDD.n643 0.00059
R54206 DVDD.n2909 DVDD.n735 0.00059
R54207 DVDD.n6402 DVDD.n6043 0.000587256
R54208 DVDD.n7411 DVDD.n7410 0.000587256
R54209 DVDD.n14293 DVDD.n8610 0.000587256
R54210 DVDD.n13269 DVDD.n13266 0.000587256
R54211 DVDD.n1755 DVDD.n1706 0.000587256
R54212 DVDD.n15089 DVDD.n6752 0.000582664
R54213 DVDD.n14841 DVDD.n14840 0.000582664
R54214 DVDD.n16704 DVDD.n2208 0.000582664
R54215 DVDD.n18157 DVDD 0.00058
R54216 DVDD DVDD.n2538 0.00058
R54217 DVDD DVDD.n16332 0.00058
R54218 DVDD DVDD.n16211 0.00058
R54219 DVDD DVDD.n2894 0.00058
R54220 DVDD.n15102 DVDD.n6348 0.000578071
R54221 DVDD.n15079 DVDD.n15078 0.000578071
R54222 DVDD.n16705 DVDD.n2165 0.000578071
R54223 DVDD.n16736 DVDD.n16735 0.000578071
R54224 DVDD.n17271 DVDD.n1605 0.000578071
R54225 DVDD.n17281 DVDD.n1262 0.000578071
R54226 DVDD.n14004 DVDD.n14003 0.000573479
R54227 DVDD.n11279 DVDD.n11227 0.000573479
R54228 DVDD.n9222 DVDD.n7657 0.000568886
R54229 DVDD.n12736 DVDD.n12477 0.000568886
R54230 DVDD.n17281 DVDD.n17280 0.000568886
R54231 DVDD.n9558 DVDD.n7678 0.000564294
R54232 DVDD.n16726 DVDD.n1813 0.000564294
R54233 DVDD.n4095 DVDD.n4082 0.00056
R54234 DVDD.n4493 DVDD.n4192 0.00056
R54235 DVDD.n3498 DVDD.n3484 0.00056
R54236 DVDD.n3337 DVDD.n2339 0.00056
R54237 DVDD.n15640 DVDD.n15603 0.00056
R54238 DVDD.n15890 DVDD.n2689 0.00056
R54239 DVDD.n15485 DVDD.n5133 0.00056
R54240 DVDD.n15970 DVDD.n2750 0.00056
R54241 DVDD.n15378 DVDD.n3112 0.00056
R54242 DVDD.n3044 DVDD.n3030 0.00056
R54243 DVDD.n8146 DVDD.n8145 0.000559702
R54244 DVDD.n11279 DVDD.n11233 0.000559702
R54245 DVDD.n13799 DVDD.n11276 0.000559702
R54246 DVDD.n11937 DVDD.n11936 0.000559702
R54247 DVDD DVDD.n11051 0.000550517
R54248 DVDD.n11573 DVDD.n11149 0.000550517
R54249 DVDD.n13488 DVDD.n13487 0.000550517
R54250 DVDD.n15101 DVDD.n15100 0.000545924
R54251 DVDD.n10230 DVDD.n8259 0.000545924
R54252 DVDD.n10693 DVDD.n10692 0.000541332
R54253 DVDD.n14270 DVDD.n10597 0.000541332
R54254 DVDD.n14003 DVDD.n11103 0.000541332
R54255 DVDD.n14000 DVDD.n11107 0.000541332
R54256 DVDD.n17003 DVDD.n1658 0.000541332
R54257 DVDD.n17263 DVDD.n17262 0.000541332
R54258 DVDD.n15131 DVDD.n5642 0.000536739
R54259 DVDD.n5987 DVDD.n5986 0.000536739
R54260 DVDD.n5938 DVDD.n5593 0.000536739
R54261 DVDD.n5991 DVDD.n5740 0.000536739
R54262 DVDD.n5988 DVDD.n5592 0.000536739
R54263 DVDD.n10232 DVDD.n10231 0.000532147
R54264 DVDD.n11568 DVDD.n11107 0.000532147
R54265 DVDD.n14863 DVDD.n7611 0.000522962
R54266 DVDD.n14860 DVDD.n7657 0.000522962
R54267 DVDD.n14826 DVDD.n8044 0.000522962
R54268 DVDD.n13765 DVDD.n13764 0.000522962
R54269 DVDD.n14849 DVDD.n7679 0.00051837
R54270 DVDD.n13744 DVDD.n12330 0.00051837
R54271 DVDD.n2156 DVDD.n1811 0.00051837
R54272 DVDD.n9560 DVDD.n9559 0.000513777
R54273 DVDD.n12435 DVDD.n12432 0.000513777
R54274 DVDD.n13474 DVDD.n13473 0.000513777
R54275 DVDD.n13470 DVDD.n12783 0.000513777
R54276 DVDD.n1264 DVDD.n1263 0.000513777
R54277 DVDD.n17298 DVDD.n915 0.000513777
R54278 DVDD.n6697 DVDD.n6403 0.000504592
R54279 DVDD.n15070 DVDD.n15069 0.000504592
R54280 DVDD.n8601 DVDD.n8258 0.000504592
R54281 DVDD.n14302 DVDD.n8259 0.000504592
R54282 DVDD.n10233 DVDD.n8609 0.000504592
R54283 DVDD.n13268 DVDD.n13267 0.000504592
R54284 DVDD.n16995 DVDD.n1712 0.000504592
R54285 DVSS.n3087 DVSS.n2135 82387.9
R54286 DVSS.n5670 DVSS.n1275 69392.3
R54287 DVSS.n1281 DVSS.n1275 69376.4
R54288 DVSS.n2135 DVSS.n1520 20752.5
R54289 DVSS.n3088 DVSS.n3087 20730.8
R54290 DVSS.n5671 DVSS.n5670 16226.6
R54291 DVSS.n5663 DVSS.n1281 16226.6
R54292 DVSS.n3518 DVSS.n2134 4180.28
R54293 DVSS.n3071 DVSS.n3070 4158.32
R54294 DVSS.n3087 DVSS.n3086 3610.1
R54295 DVSS.n3517 DVSS.n2135 3610.1
R54296 DVSS.n4956 DVSS.t24 3372.16
R54297 DVSS.n4979 DVSS.t24 3372.16
R54298 DVSS.n3086 DVSS.n3071 3351.4
R54299 DVSS.n3518 DVSS.n3517 3351.4
R54300 DVSS.t6 DVSS.n5672 2629.04
R54301 DVSS.n5667 DVSS.n1278 2402.48
R54302 DVSS.n5667 DVSS.n5666 2401.2
R54303 DVSS.n5665 DVSS.n1278 2400.01
R54304 DVSS.n5666 DVSS.n5665 2398.73
R54305 DVSS.n5662 DVSS.n1282 1820
R54306 DVSS.n5671 DVSS.n1274 1409.58
R54307 DVSS.n5664 DVSS.n5663 1409.58
R54308 DVSS.n1520 DVSS.n1274 1327.85
R54309 DVSS.n5664 DVSS.n1280 1327.85
R54310 DVSS.n1291 DVSS.n1282 1096.7
R54311 DVSS.n5673 DVSS.n1273 864.362
R54312 DVSS.t14 DVSS.n1291 843.617
R54313 DVSS.n3071 DVSS.n3069 551.231
R54314 DVSS.n3519 DVSS.n3518 551.231
R54315 DVSS.n5673 DVSS.t6 425.957
R54316 DVSS.t12 DVSS.t14 337.447
R54317 DVSS.t18 DVSS.t16 337.447
R54318 DVSS.t22 DVSS.t20 337.447
R54319 DVSS.t20 DVSS.t197 337.447
R54320 DVSS.t197 DVSS.t195 337.447
R54321 DVSS.t195 DVSS.t191 337.447
R54322 DVSS.t191 DVSS.t189 337.447
R54323 DVSS.t189 DVSS.t193 337.447
R54324 DVSS.t193 DVSS.t10 337.447
R54325 DVSS.n4744 DVSS.n1272 290.034
R54326 DVSS.n4744 DVSS.n1283 266.233
R54327 DVSS.n5661 DVSS.n1283 233.644
R54328 DVSS.n5674 DVSS.n1272 227.811
R54329 DVSS.n5674 DVSS.n1271 201.056
R54330 DVSS.t127 DVSS.n5684 196.893
R54331 DVSS.t147 DVSS.n146 196.893
R54332 DVSS.n1293 DVSS.t12 192.234
R54333 DVSS.t10 DVSS.n1273 178.405
R54334 DVSS.n5361 DVSS.n1520 177.477
R54335 DVSS.n4318 DVSS.n1280 177.222
R54336 DVSS.n5663 DVSS.n5662 177.022
R54337 DVSS.n5672 DVSS.n5671 177.022
R54338 DVSS.n1292 DVSS.t22 170.107
R54339 DVSS.n5685 DVSS.t41 168.048
R54340 DVSS.n5685 DVSS.t161 168.048
R54341 DVSS.n6428 DVSS.t83 168.048
R54342 DVSS.n6428 DVSS.t37 168.048
R54343 DVSS.n504 DVSS.t71 168.048
R54344 DVSS.n504 DVSS.t81 168.048
R54345 DVSS.t16 DVSS.n1292 167.34
R54346 DVSS.n5661 DVSS.n1284 158.357
R54347 DVSS.n1293 DVSS.t18 145.214
R54348 DVSS.n1294 DVSS.n1284 138.911
R54349 DVSS.n4980 DVSS.n1762 130.275
R54350 DVSS.n1785 DVSS.n1762 130.275
R54351 DVSS.n4955 DVSS.n1766 130.275
R54352 DVSS.n4978 DVSS.n1766 130.275
R54353 DVSS.n4956 DVSS.n1780 123.9
R54354 DVSS.n4979 DVSS.n1764 123.9
R54355 DVSS.n1784 DVSS.n1783 75.1538
R54356 DVSS.n1783 DVSS.n1760 75.1538
R54357 DVSS.n4960 DVSS.n4958 75.1538
R54358 DVSS.n4960 DVSS.n4959 75.1538
R54359 DVSS.n2417 DVSS.n1781 75.1538
R54360 DVSS.n2417 DVSS.n1767 75.1538
R54361 DVSS.t97 DVSS.t127 66.3492
R54362 DVSS.t149 DVSS.t97 66.3492
R54363 DVSS.t117 DVSS.t149 66.3492
R54364 DVSS.t35 DVSS.t117 66.3492
R54365 DVSS.t87 DVSS.t35 66.3492
R54366 DVSS.t63 DVSS.t87 66.3492
R54367 DVSS.t107 DVSS.t63 66.3492
R54368 DVSS.t77 DVSS.t107 66.3492
R54369 DVSS.t119 DVSS.t77 66.3492
R54370 DVSS.t49 DVSS.t119 66.3492
R54371 DVSS.t141 DVSS.t49 66.3492
R54372 DVSS.t65 DVSS.t141 66.3492
R54373 DVSS.t29 DVSS.t65 66.3492
R54374 DVSS.t91 DVSS.t29 66.3492
R54375 DVSS.t163 DVSS.t91 66.3492
R54376 DVSS.t99 DVSS.t163 66.3492
R54377 DVSS.t173 DVSS.t99 66.3492
R54378 DVSS.t121 DVSS.t173 66.3492
R54379 DVSS.t41 DVSS.t121 66.3492
R54380 DVSS.t161 DVSS.t47 66.3492
R54381 DVSS.t47 DVSS.t133 66.3492
R54382 DVSS.t133 DVSS.t69 66.3492
R54383 DVSS.t69 DVSS.t151 66.3492
R54384 DVSS.t151 DVSS.t85 66.3492
R54385 DVSS.t85 DVSS.t101 66.3492
R54386 DVSS.t101 DVSS.t177 66.3492
R54387 DVSS.t177 DVSS.t111 66.3492
R54388 DVSS.t111 DVSS.t31 66.3492
R54389 DVSS.t31 DVSS.t131 66.3492
R54390 DVSS.t131 DVSS.t53 66.3492
R54391 DVSS.t53 DVSS.t103 66.3492
R54392 DVSS.t103 DVSS.t73 66.3492
R54393 DVSS.t73 DVSS.t123 66.3492
R54394 DVSS.t123 DVSS.t93 66.3492
R54395 DVSS.t93 DVSS.t167 66.3492
R54396 DVSS.t167 DVSS.t59 66.3492
R54397 DVSS.t59 DVSS.t183 66.3492
R54398 DVSS.t183 DVSS.t83 66.3492
R54399 DVSS.t89 DVSS.t37 66.3492
R54400 DVSS.t51 DVSS.t89 66.3492
R54401 DVSS.t143 DVSS.t51 66.3492
R54402 DVSS.t187 DVSS.t143 66.3492
R54403 DVSS.t155 DVSS.t187 66.3492
R54404 DVSS.t39 DVSS.t155 66.3492
R54405 DVSS.t175 DVSS.t39 66.3492
R54406 DVSS.t67 DVSS.t175 66.3492
R54407 DVSS.t145 DVSS.t67 66.3492
R54408 DVSS.t79 DVSS.t145 66.3492
R54409 DVSS.t165 DVSS.t79 66.3492
R54410 DVSS.t135 DVSS.t165 66.3492
R54411 DVSS.t179 DVSS.t135 66.3492
R54412 DVSS.t105 DVSS.t179 66.3492
R54413 DVSS.t43 DVSS.t105 66.3492
R54414 DVSS.t125 DVSS.t43 66.3492
R54415 DVSS.t55 DVSS.t125 66.3492
R54416 DVSS.t137 DVSS.t55 66.3492
R54417 DVSS.t71 DVSS.t137 66.3492
R54418 DVSS.t81 DVSS.t157 66.3492
R54419 DVSS.t157 DVSS.t95 66.3492
R54420 DVSS.t95 DVSS.t181 66.3492
R54421 DVSS.t181 DVSS.t113 66.3492
R54422 DVSS.t113 DVSS.t33 66.3492
R54423 DVSS.t33 DVSS.t115 66.3492
R54424 DVSS.t115 DVSS.t57 66.3492
R54425 DVSS.t57 DVSS.t139 66.3492
R54426 DVSS.t139 DVSS.t75 66.3492
R54427 DVSS.t75 DVSS.t153 66.3492
R54428 DVSS.t153 DVSS.t45 66.3492
R54429 DVSS.t45 DVSS.t169 66.3492
R54430 DVSS.t169 DVSS.t61 66.3492
R54431 DVSS.t61 DVSS.t185 66.3492
R54432 DVSS.t185 DVSS.t109 66.3492
R54433 DVSS.t109 DVSS.t159 66.3492
R54434 DVSS.t159 DVSS.t129 66.3492
R54435 DVSS.t129 DVSS.t171 66.3492
R54436 DVSS.t171 DVSS.t147 66.3492
R54437 DVSS.n4005 DVSS.n3890 39.3263
R54438 DVSS.n5503 DVSS.n1375 39.3263
R54439 DVSS.n1294 DVSS.n1271 36.5561
R54440 DVSS.n4427 DVSS.n3890 29.1118
R54441 DVSS.n4427 DVSS.n3891 29.1118
R54442 DVSS.n4421 DVSS.n3891 29.1118
R54443 DVSS.n4421 DVSS.n3958 29.1118
R54444 DVSS.n4415 DVSS.n3958 29.1118
R54445 DVSS.n4415 DVSS.n3963 29.1118
R54446 DVSS.n4409 DVSS.n3963 29.1118
R54447 DVSS.n4409 DVSS.n3968 29.1118
R54448 DVSS.n4403 DVSS.n3968 29.1118
R54449 DVSS.n4403 DVSS.n3973 29.1118
R54450 DVSS.n4397 DVSS.n3973 29.1118
R54451 DVSS.n4397 DVSS.n3978 29.1118
R54452 DVSS.n4391 DVSS.n3978 29.1118
R54453 DVSS.n4391 DVSS.n3983 29.1118
R54454 DVSS.n4385 DVSS.n3983 29.1118
R54455 DVSS.n4385 DVSS.n3988 29.1118
R54456 DVSS.n4379 DVSS.n3988 29.1118
R54457 DVSS.n4379 DVSS.n3993 29.1118
R54458 DVSS.n4373 DVSS.n3993 29.1118
R54459 DVSS.n4373 DVSS.n3999 29.1118
R54460 DVSS.n3999 DVSS.n1808 29.1118
R54461 DVSS.n4909 DVSS.n1808 29.1118
R54462 DVSS.n4909 DVSS.n1809 29.1118
R54463 DVSS.n4903 DVSS.n1809 29.1118
R54464 DVSS.n4903 DVSS.n1816 29.1118
R54465 DVSS.n4897 DVSS.n1816 29.1118
R54466 DVSS.n4897 DVSS.n1823 29.1118
R54467 DVSS.n4891 DVSS.n1823 29.1118
R54468 DVSS.n4891 DVSS.n1828 29.1118
R54469 DVSS.n4885 DVSS.n1828 29.1118
R54470 DVSS.n4885 DVSS.n1833 29.1118
R54471 DVSS.n4879 DVSS.n1833 29.1118
R54472 DVSS.n4879 DVSS.n1838 29.1118
R54473 DVSS.n4873 DVSS.n1838 29.1118
R54474 DVSS.n4873 DVSS.n1843 29.1118
R54475 DVSS.n4867 DVSS.n1843 29.1118
R54476 DVSS.n4867 DVSS.n1848 29.1118
R54477 DVSS.n4861 DVSS.n1848 29.1118
R54478 DVSS.n4861 DVSS.n1853 29.1118
R54479 DVSS.n4855 DVSS.n1853 29.1118
R54480 DVSS.n4855 DVSS.n1858 29.1118
R54481 DVSS.n1962 DVSS.n1858 29.1118
R54482 DVSS.n4751 DVSS.n1962 29.1118
R54483 DVSS.n4751 DVSS.n1878 29.1118
R54484 DVSS.n4846 DVSS.n1878 29.1118
R54485 DVSS.n4846 DVSS.n1879 29.1118
R54486 DVSS.n4840 DVSS.n1879 29.1118
R54487 DVSS.n4840 DVSS.n1886 29.1118
R54488 DVSS.n4834 DVSS.n1886 29.1118
R54489 DVSS.n4834 DVSS.n1892 29.1118
R54490 DVSS.n4828 DVSS.n1892 29.1118
R54491 DVSS.n4828 DVSS.n1897 29.1118
R54492 DVSS.n4822 DVSS.n1897 29.1118
R54493 DVSS.n4822 DVSS.n1902 29.1118
R54494 DVSS.n4816 DVSS.n1902 29.1118
R54495 DVSS.n4816 DVSS.n1907 29.1118
R54496 DVSS.n4810 DVSS.n1907 29.1118
R54497 DVSS.n4810 DVSS.n1912 29.1118
R54498 DVSS.n4804 DVSS.n1912 29.1118
R54499 DVSS.n4804 DVSS.n1917 29.1118
R54500 DVSS.n4798 DVSS.n1917 29.1118
R54501 DVSS.n4798 DVSS.n1922 29.1118
R54502 DVSS.n4792 DVSS.n1922 29.1118
R54503 DVSS.n4792 DVSS.n1927 29.1118
R54504 DVSS.n1927 DVSS.n1596 29.1118
R54505 DVSS.n5257 DVSS.n1596 29.1118
R54506 DVSS.n5257 DVSS.n1597 29.1118
R54507 DVSS.n5251 DVSS.n1597 29.1118
R54508 DVSS.n5251 DVSS.n1604 29.1118
R54509 DVSS.n5245 DVSS.n1604 29.1118
R54510 DVSS.n5245 DVSS.n1609 29.1118
R54511 DVSS.n5239 DVSS.n1609 29.1118
R54512 DVSS.n5239 DVSS.n1614 29.1118
R54513 DVSS.n5233 DVSS.n1614 29.1118
R54514 DVSS.n5233 DVSS.n1619 29.1118
R54515 DVSS.n5227 DVSS.n1619 29.1118
R54516 DVSS.n5227 DVSS.n1624 29.1118
R54517 DVSS.n5221 DVSS.n1624 29.1118
R54518 DVSS.n5221 DVSS.n1629 29.1118
R54519 DVSS.n5215 DVSS.n1629 29.1118
R54520 DVSS.n5215 DVSS.n1634 29.1118
R54521 DVSS.n5209 DVSS.n1634 29.1118
R54522 DVSS.n5209 DVSS.n1639 29.1118
R54523 DVSS.n5203 DVSS.n1639 29.1118
R54524 DVSS.n5203 DVSS.n1645 29.1118
R54525 DVSS.n1645 DVSS.n1374 29.1118
R54526 DVSS.n5503 DVSS.n1374 29.1118
R54527 DVSS.n5361 DVSS.n1375 29.1118
R54528 DVSS.n3088 DVSS.n1280 21.9617
R54529 DVSS.n3070 DVSS.n2134 21.96
R54530 DVSS.n3328 DVSS.n3327 17.2463
R54531 DVSS.n3510 DVSS.n3509 7.85992
R54532 DVSS.n3509 DVSS.n3508 7.82456
R54533 DVSS.n4980 DVSS.n1760 7.68902
R54534 DVSS.n4958 DVSS.n1779 7.68902
R54535 DVSS.n1784 DVSS.n1779 7.68902
R54536 DVSS.n1785 DVSS.n1784 7.68902
R54537 DVSS.n1767 DVSS.n1763 7.68902
R54538 DVSS.n4959 DVSS.n1763 7.68902
R54539 DVSS.n4959 DVSS.n1765 7.68902
R54540 DVSS.n1765 DVSS.n1760 7.68902
R54541 DVSS.n4955 DVSS.n1781 7.68902
R54542 DVSS.n4957 DVSS.n1781 7.68902
R54543 DVSS.n4958 DVSS.n4957 7.68902
R54544 DVSS.n4978 DVSS.n1767 7.68902
R54545 DVSS.n5669 DVSS.n1276 6.84065
R54546 DVSS.n2379 DVSS.n1276 6.80529
R54547 DVSS.n5504 DVSS.n1373 5.28481
R54548 DVSS.n5502 DVSS.n1378 5.28481
R54549 DVSS.n5351 DVSS.n1376 5.28481
R54550 DVSS.n4329 DVSS.n4003 5.2005
R54551 DVSS.n4005 DVSS.n4003 5.2005
R54552 DVSS.n4327 DVSS.n4003 5.2005
R54553 DVSS.n4329 DVSS.n4328 5.2005
R54554 DVSS.n4328 DVSS.n4327 5.2005
R54555 DVSS.n4182 DVSS.n4037 5.2005
R54556 DVSS.n4318 DVSS.n4037 5.2005
R54557 DVSS.n4182 DVSS.n4061 5.2005
R54558 DVSS.n4318 DVSS.n4061 5.2005
R54559 DVSS.n4182 DVSS.n4036 5.2005
R54560 DVSS.n4318 DVSS.n4036 5.2005
R54561 DVSS.n4182 DVSS.n4063 5.2005
R54562 DVSS.n4318 DVSS.n4063 5.2005
R54563 DVSS.n4182 DVSS.n4035 5.2005
R54564 DVSS.n4318 DVSS.n4035 5.2005
R54565 DVSS.n4182 DVSS.n4064 5.2005
R54566 DVSS.n4318 DVSS.n4064 5.2005
R54567 DVSS.n4315 DVSS.n4009 5.2005
R54568 DVSS.n4318 DVSS.n4009 5.2005
R54569 DVSS.n4316 DVSS.n4315 5.2005
R54570 DVSS.n1522 DVSS.n1375 5.2005
R54571 DVSS.n1518 DVSS.n1375 5.2005
R54572 DVSS.n1411 DVSS.n1375 5.2005
R54573 DVSS.n5499 DVSS.n1384 5.2005
R54574 DVSS.n1384 DVSS.n1375 5.2005
R54575 DVSS.n5499 DVSS.n1383 5.2005
R54576 DVSS.n1383 DVSS.n1375 5.2005
R54577 DVSS.n5355 DVSS.n1375 5.2005
R54578 DVSS.n5359 DVSS.n5358 5.2005
R54579 DVSS.n5361 DVSS.n5359 5.2005
R54580 DVSS.n5499 DVSS.n1378 5.2005
R54581 DVSS.n1378 DVSS.n1375 5.2005
R54582 DVSS.n5358 DVSS.n1386 5.2005
R54583 DVSS.n5499 DVSS.n1386 5.2005
R54584 DVSS.n1386 DVSS.n1375 5.2005
R54585 DVSS.n5499 DVSS.n1382 5.2005
R54586 DVSS.n1382 DVSS.n1375 5.2005
R54587 DVSS.n5499 DVSS.n5498 5.2005
R54588 DVSS.n5498 DVSS.n1375 5.2005
R54589 DVSS.n5393 DVSS.n1375 5.2005
R54590 DVSS.n6442 DVSS.n180 5.02526
R54591 DVSS.n6404 DVSS.n6402 5.02526
R54592 DVSS.n269 DVSS.n268 5.02526
R54593 DVSS.n6392 DVSS.n6391 5.02526
R54594 DVSS.n6380 DVSS.n6379 5.02526
R54595 DVSS.n6497 DVSS.n6496 5.02526
R54596 DVSS.n376 DVSS.n368 5.02526
R54597 DVSS.n6289 DVSS.n6285 5.02526
R54598 DVSS.n6282 DVSS.n6274 5.02526
R54599 DVSS.n6271 DVSS.n6263 5.02526
R54600 DVSS.n6248 DVSS.n392 5.02526
R54601 DVSS.n6220 DVSS.n458 5.02526
R54602 DVSS.n6208 DVSS.n460 5.02526
R54603 DVSS.n1117 DVSS.n1109 5.02526
R54604 DVSS.n1106 DVSS.n1098 5.02526
R54605 DVSS.n6123 DVSS.n6122 5.02526
R54606 DVSS.n6115 DVSS.n1095 5.02526
R54607 DVSS.n6112 DVSS.n1138 5.02526
R54608 DVSS.n5783 DVSS.n5782 5.02526
R54609 DVSS.n6055 DVSS.n5799 5.02526
R54610 DVSS.n6068 DVSS.n6067 5.02526
R54611 DVSS.n5770 DVSS.n1197 5.02526
R54612 DVSS.n5767 DVSS.n1202 5.02526
R54613 DVSS.n1213 DVSS.n1212 5.02526
R54614 DVSS.n5750 DVSS.n1214 5.02526
R54615 DVSS.n5747 DVSS.n1216 5.02526
R54616 DVSS.n1226 DVSS.n1225 5.02526
R54617 DVSS.n5733 DVSS.n1227 5.02526
R54618 DVSS.n5730 DVSS.n1229 5.02526
R54619 DVSS.n5694 DVSS.n5693 5.02526
R54620 DVSS.n5696 DVSS.n1245 5.02526
R54621 DVSS.n5706 DVSS.n1241 5.02526
R54622 DVSS.n5641 DVSS.n5640 5.02526
R54623 DVSS.n5639 DVSS.n5638 5.02526
R54624 DVSS.n5630 DVSS.n1322 5.02526
R54625 DVSS.n5627 DVSS.n5623 5.02526
R54626 DVSS.n5622 DVSS.n5621 5.02526
R54627 DVSS.n5613 DVSS.n1327 5.02526
R54628 DVSS.n5610 DVSS.n5606 5.02526
R54629 DVSS.n5605 DVSS.n5604 5.02526
R54630 DVSS.n1313 DVSS.n1301 5.02426
R54631 DVSS.n1314 DVSS.n1302 5.02426
R54632 DVSS.n1315 DVSS.n1303 5.02426
R54633 DVSS.n1316 DVSS.n1304 5.02426
R54634 DVSS.n1317 DVSS.n1305 5.02426
R54635 DVSS.n1318 DVSS.n1306 5.02426
R54636 DVSS.n1320 DVSS.n1319 5.02426
R54637 DVSS.n5644 DVSS.n1237 5.02426
R54638 DVSS.n5711 DVSS.n5710 5.02426
R54639 DVSS.n5717 DVSS.n5716 5.02426
R54640 DVSS.n5724 DVSS.n5723 5.02426
R54641 DVSS.n5726 DVSS.n5725 5.02426
R54642 DVSS.n5737 DVSS.n1217 5.02426
R54643 DVSS.n5741 DVSS.n5740 5.02426
R54644 DVSS.n5743 DVSS.n5742 5.02426
R54645 DVSS.n5754 DVSS.n1204 5.02426
R54646 DVSS.n5758 DVSS.n5757 5.02426
R54647 DVSS.n5763 DVSS.n5762 5.02426
R54648 DVSS.n5761 DVSS.n5760 5.02426
R54649 DVSS.n6063 DVSS.n1166 5.02426
R54650 DVSS.n6096 DVSS.n6095 5.02426
R54651 DVSS.n6106 DVSS.n6105 5.02426
R54652 DVSS.n6108 DVSS.n6107 5.02426
R54653 DVSS.n1135 DVSS.n424 5.02426
R54654 DVSS.n6236 DVSS.n6235 5.02426
R54655 DVSS.n1102 DVSS.n1101 5.02426
R54656 DVSS.n1113 DVSS.n1112 5.02426
R54657 DVSS.n6204 DVSS.n6203 5.02426
R54658 DVSS.n6225 DVSS.n6224 5.02426
R54659 DVSS.n6244 DVSS.n6243 5.02426
R54660 DVSS.n6267 DVSS.n6266 5.02426
R54661 DVSS.n6278 DVSS.n6277 5.02426
R54662 DVSS.n6483 DVSS.n6482 5.02426
R54663 DVSS.n372 DVSS.n371 5.02426
R54664 DVSS.n6492 DVSS.n6491 5.02426
R54665 DVSS.n107 DVSS.n64 5.02426
R54666 DVSS.n6387 DVSS.n6386 5.02426
R54667 DVSS.n264 DVSS.n263 5.02426
R54668 DVSS.n6410 DVSS.n6409 5.02426
R54669 DVSS.n6415 DVSS.n6414 5.02426
R54670 DVSS.n3094 DVSS.n2368 4.7928
R54671 DVSS.n3516 DVSS.n2136 4.72792
R54672 DVSS.n3283 DVSS.n2136 4.60071
R54673 DVSS.n3078 DVSS.n3077 4.60071
R54674 DVSS.n6071 DVSS.n1194 4.5005
R54675 DVSS.n6071 DVSS.n1191 4.5005
R54676 DVSS.n6071 DVSS.n1196 4.5005
R54677 DVSS.n6071 DVSS.n1186 4.5005
R54678 DVSS.n6072 DVSS.n1183 4.5005
R54679 DVSS.n6072 DVSS.n6071 4.5005
R54680 DVSS.n6071 DVSS.n1182 4.5005
R54681 DVSS.n6071 DVSS.n6070 4.5005
R54682 DVSS.n5552 DVSS.n1333 4.5005
R54683 DVSS.n5509 DVSS.n5508 4.5005
R54684 DVSS.n1525 DVSS.n1369 4.5005
R54685 DVSS.n5346 DVSS.n1525 4.5005
R54686 DVSS.n5131 DVSS.n1524 4.5005
R54687 DVSS.n5088 DVSS.n5087 4.5005
R54688 DVSS.n5086 DVSS.n5085 4.5005
R54689 DVSS.n2878 DVSS.n1696 4.5005
R54690 DVSS.n2880 DVSS.n2879 4.5005
R54691 DVSS.n2883 DVSS.n2132 4.5005
R54692 DVSS.n2883 DVSS.n2131 4.5005
R54693 DVSS.n2883 DVSS.n2614 4.5005
R54694 DVSS.n2883 DVSS.n2610 4.5005
R54695 DVSS.n2884 DVSS.n2883 4.5005
R54696 DVSS.n2885 DVSS.n2599 4.5005
R54697 DVSS.n2927 DVSS.n2600 4.5005
R54698 DVSS.n2926 DVSS.n2599 4.5005
R54699 DVSS.n2927 DVSS.n2926 4.5005
R54700 DVSS.n2880 DVSS.n2614 4.5005
R54701 DVSS.n2880 DVSS.n2131 4.5005
R54702 DVSS.n3522 DVSS.n2129 4.5005
R54703 DVSS.n3520 DVSS.n2129 4.5005
R54704 DVSS.n3522 DVSS.n3521 4.5005
R54705 DVSS.n3521 DVSS.n3520 4.5005
R54706 DVSS.n3505 DVSS.n2141 4.5005
R54707 DVSS.n3507 DVSS.n3506 4.5005
R54708 DVSS.n3511 DVSS.n2139 4.5005
R54709 DVSS.n3513 DVSS.n3512 4.5005
R54710 DVSS.n3285 DVSS.n3283 4.5005
R54711 DVSS.n3287 DVSS.n3286 4.5005
R54712 DVSS.n3289 DVSS.n3288 4.5005
R54713 DVSS.n3290 DVSS.n3281 4.5005
R54714 DVSS.n3292 DVSS.n3291 4.5005
R54715 DVSS.n3076 DVSS.n3075 4.5005
R54716 DVSS.n3077 DVSS.n3074 4.5005
R54717 DVSS.n3040 DVSS.n3037 4.5005
R54718 DVSS.n3040 DVSS.n1768 4.5005
R54719 DVSS.n4985 DVSS.n1756 4.5005
R54720 DVSS.n4983 DVSS.n1756 4.5005
R54721 DVSS.n4971 DVSS.n4970 4.5005
R54722 DVSS.n4975 DVSS.n1771 4.5005
R54723 DVSS.n4972 DVSS.n1770 4.5005
R54724 DVSS.n4968 DVSS.n4966 4.5005
R54725 DVSS.n4984 DVSS.n4983 4.5005
R54726 DVSS.n4985 DVSS.n4984 4.5005
R54727 DVSS.n5005 DVSS.n1730 4.5005
R54728 DVSS.n5005 DVSS.n5004 4.5005
R54729 DVSS.n3527 DVSS.n2125 4.5005
R54730 DVSS.n3525 DVSS.n2125 4.5005
R54731 DVSS.n3527 DVSS.n3526 4.5005
R54732 DVSS.n3526 DVSS.n3525 4.5005
R54733 DVSS.n6052 DVSS.n5805 4.5005
R54734 DVSS.n6053 DVSS.n6052 4.5005
R54735 DVSS.n6049 DVSS.n6048 4.5005
R54736 DVSS.n6049 DVSS.n1180 4.5005
R54737 DVSS.n6052 DVSS.n1180 4.5005
R54738 DVSS.n6052 DVSS.n1179 4.5005
R54739 DVSS.n6052 DVSS.n6051 4.5005
R54740 DVSS.n5586 DVSS.n5585 4.5005
R54741 DVSS.n4703 DVSS.n4702 4.5005
R54742 DVSS.n5262 DVSS.n1564 4.5005
R54743 DVSS.n5166 DVSS.n1564 4.5005
R54744 DVSS.n5165 DVSS.n5164 4.5005
R54745 DVSS.n3756 DVSS.n3755 4.5005
R54746 DVSS.n3754 DVSS.n1713 4.5005
R54747 DVSS.n1731 DVSS.n1713 4.5005
R54748 DVSS.n5006 DVSS.n1713 4.5005
R54749 DVSS.n5007 DVSS.n1727 4.5005
R54750 DVSS.n5007 DVSS.n1719 4.5005
R54751 DVSS.n1719 DVSS.n1713 4.5005
R54752 DVSS.n5007 DVSS.n1728 4.5005
R54753 DVSS.n1728 DVSS.n1713 4.5005
R54754 DVSS.n3044 DVSS.n3041 4.5005
R54755 DVSS.n2401 DVSS.n2128 4.5005
R54756 DVSS.n3044 DVSS.n2127 4.5005
R54757 DVSS.n3044 DVSS.n3043 4.5005
R54758 DVSS.n3051 DVSS.n2401 4.5005
R54759 DVSS.n3052 DVSS.n2400 4.5005
R54760 DVSS.n3061 DVSS.n2399 4.5005
R54761 DVSS.n2399 DVSS.n2398 4.5005
R54762 DVSS.n2400 DVSS.n2398 4.5005
R54763 DVSS.n3045 DVSS.n2401 4.5005
R54764 DVSS.n3043 DVSS.n2401 4.5005
R54765 DVSS.n2401 DVSS.n2127 4.5005
R54766 DVSS.n5007 DVSS.n1718 4.5005
R54767 DVSS.n5007 DVSS.n5006 4.5005
R54768 DVSS.n6049 DVSS.n5800 4.5005
R54769 DVSS.n5701 DVSS.n1246 4.5005
R54770 DVSS.n5698 DVSS.n5695 4.5005
R54771 DVSS.n5703 DVSS.n1246 4.5005
R54772 DVSS.n5698 DVSS.n5697 4.5005
R54773 DVSS.n5689 DVSS.n1234 4.5005
R54774 DVSS.n5689 DVSS.n5688 4.5005
R54775 DVSS.n5687 DVSS.n5686 4.5005
R54776 DVSS.n5688 DVSS.n5687 4.5005
R54777 DVSS.n3036 DVSS.n2407 4.5005
R54778 DVSS.n1754 DVSS.n1748 4.5005
R54779 DVSS.n4992 DVSS.n1748 4.5005
R54780 DVSS.n4990 DVSS.n1748 4.5005
R54781 DVSS.n4986 DVSS.n1748 4.5005
R54782 DVSS.n4964 DVSS.n4963 4.5005
R54783 DVSS.n4965 DVSS.n4964 4.5005
R54784 DVSS.n4965 DVSS.n1774 4.5005
R54785 DVSS.n2421 DVSS.n2420 4.5005
R54786 DVSS.n2422 DVSS.n2421 4.5005
R54787 DVSS.n2423 DVSS.n2422 4.5005
R54788 DVSS.n3036 DVSS.n3035 4.5005
R54789 DVSS.n3035 DVSS.n2410 4.5005
R54790 DVSS.n3035 DVSS.n3034 4.5005
R54791 DVSS.n2420 DVSS.n2419 4.5005
R54792 DVSS.n4963 DVSS.n4962 4.5005
R54793 DVSS.n4991 DVSS.n4986 4.5005
R54794 DVSS.n4991 DVSS.n4990 4.5005
R54795 DVSS.n4992 DVSS.n4991 4.5005
R54796 DVSS.n4991 DVSS.n1754 4.5005
R54797 DVSS.n5002 DVSS.n5001 4.5005
R54798 DVSS.n5001 DVSS.n1736 4.5005
R54799 DVSS.n5001 DVSS.n1734 4.5005
R54800 DVSS.n5001 DVSS.n5000 4.5005
R54801 DVSS.n3530 DVSS.n2121 4.5005
R54802 DVSS.n3528 DVSS.n2121 4.5005
R54803 DVSS.n3530 DVSS.n2116 4.5005
R54804 DVSS.n3528 DVSS.n2116 4.5005
R54805 DVSS.n3530 DVSS.n3529 4.5005
R54806 DVSS.n3529 DVSS.n3528 4.5005
R54807 DVSS.n5787 DVSS.n5775 4.5005
R54808 DVSS.n5787 DVSS.n5776 4.5005
R54809 DVSS.n6060 DVSS.n5787 4.5005
R54810 DVSS.n5780 DVSS.n5775 4.5005
R54811 DVSS.n5780 DVSS.n5776 4.5005
R54812 DVSS.n6060 DVSS.n5780 4.5005
R54813 DVSS.n5788 DVSS.n5776 4.5005
R54814 DVSS.n6060 DVSS.n5788 4.5005
R54815 DVSS.n5779 DVSS.n5776 4.5005
R54816 DVSS.n6060 DVSS.n5779 4.5005
R54817 DVSS.n5790 DVSS.n5776 4.5005
R54818 DVSS.n6060 DVSS.n5790 4.5005
R54819 DVSS.n5778 DVSS.n5776 4.5005
R54820 DVSS.n6060 DVSS.n5778 4.5005
R54821 DVSS.n6060 DVSS.n5792 4.5005
R54822 DVSS.n5775 DVSS.n1176 4.5005
R54823 DVSS.n5776 DVSS.n1176 4.5005
R54824 DVSS.n5798 DVSS.n1176 4.5005
R54825 DVSS.n6060 DVSS.n1176 4.5005
R54826 DVSS.n5775 DVSS.n1174 4.5005
R54827 DVSS.n5776 DVSS.n1174 4.5005
R54828 DVSS.n6060 DVSS.n1174 4.5005
R54829 DVSS.n6061 DVSS.n5775 4.5005
R54830 DVSS.n6061 DVSS.n5776 4.5005
R54831 DVSS.n6061 DVSS.n6060 4.5005
R54832 DVSS.n1994 DVSS.n1261 4.5005
R54833 DVSS.n4740 DVSS.n1261 4.5005
R54834 DVSS.n4742 DVSS.n1261 4.5005
R54835 DVSS.n4740 DVSS.n1979 4.5005
R54836 DVSS.n4742 DVSS.n1979 4.5005
R54837 DVSS.n4740 DVSS.n1981 4.5005
R54838 DVSS.n4742 DVSS.n1981 4.5005
R54839 DVSS.n4740 DVSS.n1978 4.5005
R54840 DVSS.n4742 DVSS.n1978 4.5005
R54841 DVSS.n4740 DVSS.n1982 4.5005
R54842 DVSS.n4742 DVSS.n1982 4.5005
R54843 DVSS.n4740 DVSS.n1977 4.5005
R54844 DVSS.n4742 DVSS.n1977 4.5005
R54845 DVSS.n4740 DVSS.n1983 4.5005
R54846 DVSS.n4742 DVSS.n1983 4.5005
R54847 DVSS.n4740 DVSS.n1976 4.5005
R54848 DVSS.n4742 DVSS.n1976 4.5005
R54849 DVSS.n4741 DVSS.n4740 4.5005
R54850 DVSS.n4742 DVSS.n4741 4.5005
R54851 DVSS.n4740 DVSS.n1975 4.5005
R54852 DVSS.n4742 DVSS.n1975 4.5005
R54853 DVSS.n4743 DVSS.n4742 4.5005
R54854 DVSS.n4501 DVSS.n1971 4.5005
R54855 DVSS.n4596 DVSS.n1971 4.5005
R54856 DVSS.n4594 DVSS.n1971 4.5005
R54857 DVSS.n4596 DVSS.n4518 4.5005
R54858 DVSS.n4594 DVSS.n4518 4.5005
R54859 DVSS.n4596 DVSS.n4516 4.5005
R54860 DVSS.n4594 DVSS.n4516 4.5005
R54861 DVSS.n4596 DVSS.n4520 4.5005
R54862 DVSS.n4594 DVSS.n4520 4.5005
R54863 DVSS.n4596 DVSS.n4515 4.5005
R54864 DVSS.n4594 DVSS.n4515 4.5005
R54865 DVSS.n4596 DVSS.n4522 4.5005
R54866 DVSS.n4594 DVSS.n4522 4.5005
R54867 DVSS.n4596 DVSS.n4514 4.5005
R54868 DVSS.n4594 DVSS.n4514 4.5005
R54869 DVSS.n4596 DVSS.n4524 4.5005
R54870 DVSS.n4594 DVSS.n4524 4.5005
R54871 DVSS.n4596 DVSS.n4513 4.5005
R54872 DVSS.n4594 DVSS.n4513 4.5005
R54873 DVSS.n4596 DVSS.n4526 4.5005
R54874 DVSS.n4594 DVSS.n4526 4.5005
R54875 DVSS.n4596 DVSS.n4512 4.5005
R54876 DVSS.n4594 DVSS.n4512 4.5005
R54877 DVSS.n4596 DVSS.n4528 4.5005
R54878 DVSS.n4594 DVSS.n4528 4.5005
R54879 DVSS.n4596 DVSS.n4511 4.5005
R54880 DVSS.n4594 DVSS.n4511 4.5005
R54881 DVSS.n4596 DVSS.n4530 4.5005
R54882 DVSS.n4594 DVSS.n4530 4.5005
R54883 DVSS.n4596 DVSS.n4510 4.5005
R54884 DVSS.n4594 DVSS.n4510 4.5005
R54885 DVSS.n4596 DVSS.n4532 4.5005
R54886 DVSS.n4594 DVSS.n4532 4.5005
R54887 DVSS.n4596 DVSS.n4509 4.5005
R54888 DVSS.n4594 DVSS.n4509 4.5005
R54889 DVSS.n4596 DVSS.n4534 4.5005
R54890 DVSS.n4594 DVSS.n4534 4.5005
R54891 DVSS.n4596 DVSS.n4508 4.5005
R54892 DVSS.n4594 DVSS.n4508 4.5005
R54893 DVSS.n4596 DVSS.n4536 4.5005
R54894 DVSS.n4594 DVSS.n4536 4.5005
R54895 DVSS.n4596 DVSS.n4507 4.5005
R54896 DVSS.n4594 DVSS.n4507 4.5005
R54897 DVSS.n4596 DVSS.n4595 4.5005
R54898 DVSS.n4595 DVSS.n4594 4.5005
R54899 DVSS.n4594 DVSS.n1873 4.5005
R54900 DVSS.n4594 DVSS.n1867 4.5005
R54901 DVSS.n3791 DVSS.n3726 4.5005
R54902 DVSS.n3807 DVSS.n3791 4.5005
R54903 DVSS.n3810 DVSS.n3791 4.5005
R54904 DVSS.n3807 DVSS.n3735 4.5005
R54905 DVSS.n3810 DVSS.n3735 4.5005
R54906 DVSS.n3807 DVSS.n3794 4.5005
R54907 DVSS.n3810 DVSS.n3794 4.5005
R54908 DVSS.n3807 DVSS.n3734 4.5005
R54909 DVSS.n3810 DVSS.n3734 4.5005
R54910 DVSS.n3807 DVSS.n3797 4.5005
R54911 DVSS.n3810 DVSS.n3797 4.5005
R54912 DVSS.n3807 DVSS.n3733 4.5005
R54913 DVSS.n3810 DVSS.n3733 4.5005
R54914 DVSS.n3807 DVSS.n3800 4.5005
R54915 DVSS.n3810 DVSS.n3800 4.5005
R54916 DVSS.n3807 DVSS.n3732 4.5005
R54917 DVSS.n3810 DVSS.n3732 4.5005
R54918 DVSS.n3807 DVSS.n3803 4.5005
R54919 DVSS.n3810 DVSS.n3803 4.5005
R54920 DVSS.n3807 DVSS.n3731 4.5005
R54921 DVSS.n3810 DVSS.n3731 4.5005
R54922 DVSS.n3810 DVSS.n3809 4.5005
R54923 DVSS.n3804 DVSS.n1752 4.5005
R54924 DVSS.n3804 DVSS.n1739 4.5005
R54925 DVSS.n3804 DVSS.n1740 4.5005
R54926 DVSS.n1752 DVSS.n1735 4.5005
R54927 DVSS.n1739 DVSS.n1735 4.5005
R54928 DVSS.n1740 DVSS.n1735 4.5005
R54929 DVSS.n1740 DVSS.n1733 4.5005
R54930 DVSS.n4997 DVSS.n1740 4.5005
R54931 DVSS.n1745 DVSS.n1739 4.5005
R54932 DVSS.n1745 DVSS.n1740 4.5005
R54933 DVSS.n1750 DVSS.n1739 4.5005
R54934 DVSS.n1750 DVSS.n1740 4.5005
R54935 DVSS.n1749 DVSS.n1739 4.5005
R54936 DVSS.n1749 DVSS.n1740 4.5005
R54937 DVSS.n4987 DVSS.n1739 4.5005
R54938 DVSS.n4987 DVSS.n1740 4.5005
R54939 DVSS.n4989 DVSS.n1740 4.5005
R54940 DVSS.n1752 DVSS.n1742 4.5005
R54941 DVSS.n1742 DVSS.n1739 4.5005
R54942 DVSS.n4996 DVSS.n1742 4.5005
R54943 DVSS.n1742 DVSS.n1740 4.5005
R54944 DVSS.n4995 DVSS.n1752 4.5005
R54945 DVSS.n4995 DVSS.n1739 4.5005
R54946 DVSS.n4996 DVSS.n4995 4.5005
R54947 DVSS.n4995 DVSS.n1740 4.5005
R54948 DVSS.n2752 DVSS.n2745 4.5005
R54949 DVSS.n2765 DVSS.n2752 4.5005
R54950 DVSS.n2752 DVSS.n2647 4.5005
R54951 DVSS.n2765 DVSS.n2751 4.5005
R54952 DVSS.n2751 DVSS.n2647 4.5005
R54953 DVSS.n2647 DVSS.n2124 4.5005
R54954 DVSS.n2765 DVSS.n2749 4.5005
R54955 DVSS.n2749 DVSS.n2647 4.5005
R54956 DVSS.n2765 DVSS.n2755 4.5005
R54957 DVSS.n2755 DVSS.n2647 4.5005
R54958 DVSS.n2765 DVSS.n2748 4.5005
R54959 DVSS.n2748 DVSS.n2647 4.5005
R54960 DVSS.n2765 DVSS.n2757 4.5005
R54961 DVSS.n2757 DVSS.n2647 4.5005
R54962 DVSS.n2765 DVSS.n2747 4.5005
R54963 DVSS.n2763 DVSS.n2747 4.5005
R54964 DVSS.n2747 DVSS.n2647 4.5005
R54965 DVSS.n2534 DVSS.n2525 4.5005
R54966 DVSS.n2983 DVSS.n2534 4.5005
R54967 DVSS.n2981 DVSS.n2534 4.5005
R54968 DVSS.n2983 DVSS.n2536 4.5005
R54969 DVSS.n2981 DVSS.n2536 4.5005
R54970 DVSS.n2983 DVSS.n2533 4.5005
R54971 DVSS.n2981 DVSS.n2533 4.5005
R54972 DVSS.n2983 DVSS.n2538 4.5005
R54973 DVSS.n2981 DVSS.n2538 4.5005
R54974 DVSS.n2983 DVSS.n2532 4.5005
R54975 DVSS.n2981 DVSS.n2532 4.5005
R54976 DVSS.n2983 DVSS.n2540 4.5005
R54977 DVSS.n2981 DVSS.n2540 4.5005
R54978 DVSS.n2983 DVSS.n2531 4.5005
R54979 DVSS.n2981 DVSS.n2531 4.5005
R54980 DVSS.n2983 DVSS.n2982 4.5005
R54981 DVSS.n2982 DVSS.n2981 4.5005
R54982 DVSS.n2981 DVSS.n2397 4.5005
R54983 DVSS.n2525 DVSS.n2396 4.5005
R54984 DVSS.n2983 DVSS.n2396 4.5005
R54985 DVSS.n2546 DVSS.n2396 4.5005
R54986 DVSS.n2981 DVSS.n2396 4.5005
R54987 DVSS.n2765 DVSS.n2764 4.5005
R54988 DVSS.n2764 DVSS.n2763 4.5005
R54989 DVSS.n2764 DVSS.n2647 4.5005
R54990 DVSS.n2746 DVSS.n2745 4.5005
R54991 DVSS.n2765 DVSS.n2746 4.5005
R54992 DVSS.n2763 DVSS.n2746 4.5005
R54993 DVSS.n2746 DVSS.n2647 4.5005
R54994 DVSS.n2745 DVSS.n2122 4.5005
R54995 DVSS.n2765 DVSS.n2122 4.5005
R54996 DVSS.n2763 DVSS.n2122 4.5005
R54997 DVSS.n2647 DVSS.n2122 4.5005
R54998 DVSS.n4997 DVSS.n4996 4.5005
R54999 DVSS.n4997 DVSS.n1739 4.5005
R55000 DVSS.n4996 DVSS.n1733 4.5005
R55001 DVSS.n1739 DVSS.n1733 4.5005
R55002 DVSS.n1752 DVSS.n1733 4.5005
R55003 DVSS.n4549 DVSS.n1867 4.5005
R55004 DVSS.n4596 DVSS.n1867 4.5005
R55005 DVSS.n4501 DVSS.n1867 4.5005
R55006 DVSS.n6059 DVSS.n5776 4.5005
R55007 DVSS.n6059 DVSS.n5798 4.5005
R55008 DVSS.n6060 DVSS.n6059 4.5005
R55009 DVSS.n1872 DVSS.n1863 4.5005
R55010 DVSS.n4849 DVSS.n1863 4.5005
R55011 DVSS.n4851 DVSS.n1863 4.5005
R55012 DVSS.n4849 DVSS.n1865 4.5005
R55013 DVSS.n4851 DVSS.n1865 4.5005
R55014 DVSS.n4849 DVSS.n1862 4.5005
R55015 DVSS.n4851 DVSS.n1862 4.5005
R55016 DVSS.n4851 DVSS.n1866 4.5005
R55017 DVSS.n1872 DVSS.n1866 4.5005
R55018 DVSS.n1872 DVSS.n1861 4.5005
R55019 DVSS.n1870 DVSS.n1861 4.5005
R55020 DVSS.n4851 DVSS.n1861 4.5005
R55021 DVSS.n4850 DVSS.n1872 4.5005
R55022 DVSS.n4850 DVSS.n4849 4.5005
R55023 DVSS.n4850 DVSS.n1870 4.5005
R55024 DVSS.n4851 DVSS.n4850 4.5005
R55025 DVSS.n6081 DVSS.n1172 4.5005
R55026 DVSS.n6079 DVSS.n6078 4.5005
R55027 DVSS.n6077 DVSS.n6076 4.5005
R55028 DVSS.n6076 DVSS.n6075 4.5005
R55029 DVSS.n6074 DVSS.n6073 4.5005
R55030 DVSS.n6073 DVSS.n214 4.5005
R55031 DVSS.n6084 DVSS.n6083 4.5005
R55032 DVSS.n6083 DVSS.n6082 4.5005
R55033 DVSS.n5721 DVSS.n5720 4.5005
R55034 DVSS.n5720 DVSS.n5719 4.5005
R55035 DVSS.n3032 DVSS.n3028 4.5005
R55036 DVSS.n4946 DVSS.n1793 4.5005
R55037 DVSS.n4946 DVSS.n4945 4.5005
R55038 DVSS.n4950 DVSS.n4949 4.5005
R55039 DVSS.n3030 DVSS.n1787 4.5005
R55040 DVSS.n3032 DVSS.n3031 4.5005
R55041 DVSS.n4952 DVSS.n4951 4.5005
R55042 DVSS.n4947 DVSS.n1791 4.5005
R55043 DVSS.n4945 DVSS.n4944 4.5005
R55044 DVSS.n4944 DVSS.n1793 4.5005
R55045 DVSS.n4934 DVSS.n1737 4.5005
R55046 DVSS.n4934 DVSS.n4933 4.5005
R55047 DVSS.n3533 DVSS.n2112 4.5005
R55048 DVSS.n3531 DVSS.n2112 4.5005
R55049 DVSS.n3533 DVSS.n3532 4.5005
R55050 DVSS.n3532 DVSS.n3531 4.5005
R55051 DVSS.n6103 DVSS.n6102 4.5005
R55052 DVSS.n6102 DVSS.n1146 4.5005
R55053 DVSS.n6099 DVSS.n1155 4.5005
R55054 DVSS.n6099 DVSS.n1150 4.5005
R55055 DVSS.n6102 DVSS.n1150 4.5005
R55056 DVSS.n6102 DVSS.n1144 4.5005
R55057 DVSS.n6102 DVSS.n6101 4.5005
R55058 DVSS.n2011 DVSS.n1298 4.5005
R55059 DVSS.n4645 DVSS.n4644 4.5005
R55060 DVSS.n4640 DVSS.n4639 4.5005
R55061 DVSS.n4639 DVSS.n4638 4.5005
R55062 DVSS.n4914 DVSS.n1802 4.5005
R55063 DVSS.n4925 DVSS.n1801 4.5005
R55064 DVSS.n4926 DVSS.n1799 4.5005
R55065 DVSS.n4928 DVSS.n1799 4.5005
R55066 DVSS.n4935 DVSS.n1799 4.5005
R55067 DVSS.n4943 DVSS.n1798 4.5005
R55068 DVSS.n1798 DVSS.n1797 4.5005
R55069 DVSS.n1799 DVSS.n1797 4.5005
R55070 DVSS.n1798 DVSS.n1794 4.5005
R55071 DVSS.n1799 DVSS.n1794 4.5005
R55072 DVSS.n3027 DVSS.n3026 4.5005
R55073 DVSS.n3023 DVSS.n2115 4.5005
R55074 DVSS.n3026 DVSS.n2114 4.5005
R55075 DVSS.n3026 DVSS.n2431 4.5005
R55076 DVSS.n3023 DVSS.n3021 4.5005
R55077 DVSS.n3020 DVSS.n3019 4.5005
R55078 DVSS.n3017 DVSS.n3013 4.5005
R55079 DVSS.n3018 DVSS.n3017 4.5005
R55080 DVSS.n3019 DVSS.n3018 4.5005
R55081 DVSS.n3023 DVSS.n2432 4.5005
R55082 DVSS.n3023 DVSS.n2431 4.5005
R55083 DVSS.n3023 DVSS.n2114 4.5005
R55084 DVSS.n4937 DVSS.n1798 4.5005
R55085 DVSS.n4935 DVSS.n1798 4.5005
R55086 DVSS.n6099 DVSS.n6098 4.5005
R55087 DVSS.n498 DVSS.n496 4.5005
R55088 DVSS.n506 DVSS.n505 4.5005
R55089 DVSS.n507 DVSS.n506 4.5005
R55090 DVSS.n6258 DVSS.n6257 4.5005
R55091 DVSS.n1072 DVSS.n213 4.5005
R55092 DVSS.n497 DVSS.n496 4.5005
R55093 DVSS.n508 DVSS.n501 4.5005
R55094 DVSS.n508 DVSS.n507 4.5005
R55095 DVSS.n6257 DVSS.n6256 4.5005
R55096 DVSS.n1074 DVSS.n213 4.5005
R55097 DVSS.n5653 DVSS.n1300 4.5005
R55098 DVSS.n5684 DVSS.n1254 4.5005
R55099 DVSS.n5682 DVSS.n1254 4.5005
R55100 DVSS.n5588 DVSS.n5587 4.5005
R55101 DVSS.n5599 DVSS.n5598 4.5005
R55102 DVSS.n5683 DVSS.n1258 4.5005
R55103 DVSS.n5684 DVSS.n5683 4.5005
R55104 DVSS.n5683 DVSS.n5682 4.5005
R55105 DVSS.n5656 DVSS.n1299 4.5005
R55106 DVSS.n5681 DVSS.n1258 4.5005
R55107 DVSS.n5682 DVSS.n5681 4.5005
R55108 DVSS.n5591 DVSS.n1260 4.5005
R55109 DVSS.n5596 DVSS.n1332 4.5005
R55110 DVSS.n6463 DVSS.n6462 4.5005
R55111 DVSS.n138 DVSS.n123 4.5005
R55112 DVSS.n6467 DVSS.n123 4.5005
R55113 DVSS.n6465 DVSS.n139 4.5005
R55114 DVSS.n208 DVSS.n148 4.5005
R55115 DVSS.n6435 DVSS.n208 4.5005
R55116 DVSS.n6433 DVSS.n209 4.5005
R55117 DVSS.n6431 DVSS.n209 4.5005
R55118 DVSS.n6468 DVSS.n138 4.5005
R55119 DVSS.n6468 DVSS.n6467 4.5005
R55120 DVSS.n6465 DVSS.n6464 4.5005
R55121 DVSS.n6464 DVSS.n143 4.5005
R55122 DVSS.n6464 DVSS.n146 4.5005
R55123 DVSS.n6464 DVSS.n142 4.5005
R55124 DVSS.n6464 DVSS.n6463 4.5005
R55125 DVSS.n6434 DVSS.n148 4.5005
R55126 DVSS.n6435 DVSS.n6434 4.5005
R55127 DVSS.n6433 DVSS.n6432 4.5005
R55128 DVSS.n6432 DVSS.n6431 4.5005
R55129 DVSS.n6425 DVSS.n6424 4.5005
R55130 DVSS.n6424 DVSS.n6423 4.5005
R55131 DVSS.n6425 DVSS.n221 4.5005
R55132 DVSS.n6423 DVSS.n221 4.5005
R55133 DVSS.n1312 DVSS.n1311 4.5005
R55134 DVSS.n1309 DVSS.n1308 4.5005
R55135 DVSS.n495 DVSS.n492 4.5005
R55136 DVSS.n5714 DVSS.n1230 4.5005
R55137 DVSS.n5715 DVSS.n5714 4.5005
R55138 DVSS.n6085 DVSS.n217 4.5005
R55139 DVSS.n6086 DVSS.n6085 4.5005
R55140 DVSS.n495 DVSS.n494 4.5005
R55141 DVSS.n2110 DVSS.n2109 4.5005
R55142 DVSS.n3537 DVSS.n2110 4.5005
R55143 DVSS.n3538 DVSS.n2109 4.5005
R55144 DVSS.n3538 DVSS.n3537 4.5005
R55145 DVSS.n6093 DVSS.n1140 4.5005
R55146 DVSS.n6094 DVSS.n6093 4.5005
R55147 DVSS.n6090 DVSS.n6089 4.5005
R55148 DVSS.n6090 DVSS.n1165 4.5005
R55149 DVSS.n6093 DVSS.n1165 4.5005
R55150 DVSS.n6093 DVSS.n1160 4.5005
R55151 DVSS.n6093 DVSS.n6092 4.5005
R55152 DVSS.n3942 DVSS.n3941 4.5005
R55153 DVSS.n3953 DVSS.n3895 4.5005
R55154 DVSS.n4448 DVSS.n2057 4.5005
R55155 DVSS.n4448 DVSS.n4447 4.5005
R55156 DVSS.n3884 DVSS.n3883 4.5005
R55157 DVSS.n3695 DVSS.n3694 4.5005
R55158 DVSS.n3693 DVSS.n3692 4.5005
R55159 DVSS.n3546 DVSS.n3545 4.5005
R55160 DVSS.n3544 DVSS.n3543 4.5005
R55161 DVSS.n3540 DVSS.n3539 4.5005
R55162 DVSS.n3543 DVSS.n2101 4.5005
R55163 DVSS.n3543 DVSS.n2104 4.5005
R55164 DVSS.n3540 DVSS.n2107 4.5005
R55165 DVSS.n2472 DVSS.n2458 4.5005
R55166 DVSS.n2470 DVSS.n2465 4.5005
R55167 DVSS.n2471 DVSS.n2470 4.5005
R55168 DVSS.n2472 DVSS.n2471 4.5005
R55169 DVSS.n3540 DVSS.n2105 4.5005
R55170 DVSS.n3540 DVSS.n2104 4.5005
R55171 DVSS.n3540 DVSS.n2101 4.5005
R55172 DVSS.n6090 DVSS.n1157 4.5005
R55173 DVSS.n6421 DVSS.n240 4.5005
R55174 DVSS.n6421 DVSS.n243 4.5005
R55175 DVSS.n6421 DVSS.n239 4.5005
R55176 DVSS.n6421 DVSS.n245 4.5005
R55177 DVSS.n6421 DVSS.n236 4.5005
R55178 DVSS.n6421 DVSS.n6412 4.5005
R55179 DVSS.n6421 DVSS.n233 4.5005
R55180 DVSS.n6421 DVSS.n6417 4.5005
R55181 DVSS.n6421 DVSS.n230 4.5005
R55182 DVSS.n6421 DVSS.n6420 4.5005
R55183 DVSS.n225 DVSS.n223 4.5005
R55184 DVSS.n6421 DVSS.n225 4.5005
R55185 DVSS.n223 DVSS.n222 4.5005
R55186 DVSS.n6421 DVSS.n222 4.5005
R55187 DVSS.n6473 DVSS.n6472 4.5005
R55188 DVSS.n6472 DVSS.n118 4.5005
R55189 DVSS.n6470 DVSS.n133 4.5005
R55190 DVSS.n6470 DVSS.n135 4.5005
R55191 DVSS.n6470 DVSS.n131 4.5005
R55192 DVSS.n6470 DVSS.n136 4.5005
R55193 DVSS.n6470 DVSS.n129 4.5005
R55194 DVSS.n6470 DVSS.n137 4.5005
R55195 DVSS.n6470 DVSS.n127 4.5005
R55196 DVSS.n6470 DVSS.n6469 4.5005
R55197 DVSS.n6472 DVSS.n111 4.5005
R55198 DVSS.n6470 DVSS.n111 4.5005
R55199 DVSS.n6472 DVSS.n6471 4.5005
R55200 DVSS.n6471 DVSS.n6470 4.5005
R55201 DVSS.n165 DVSS.n152 4.5005
R55202 DVSS.n165 DVSS.n153 4.5005
R55203 DVSS.n6460 DVSS.n165 4.5005
R55204 DVSS.n167 DVSS.n152 4.5005
R55205 DVSS.n167 DVSS.n153 4.5005
R55206 DVSS.n6460 DVSS.n167 4.5005
R55207 DVSS.n6460 DVSS.n164 4.5005
R55208 DVSS.n6456 DVSS.n164 4.5005
R55209 DVSS.n164 DVSS.n152 4.5005
R55210 DVSS.n169 DVSS.n152 4.5005
R55211 DVSS.n6460 DVSS.n169 4.5005
R55212 DVSS.n163 DVSS.n153 4.5005
R55213 DVSS.n6460 DVSS.n163 4.5005
R55214 DVSS.n6460 DVSS.n171 4.5005
R55215 DVSS.n6460 DVSS.n162 4.5005
R55216 DVSS.n6456 DVSS.n162 4.5005
R55217 DVSS.n162 DVSS.n152 4.5005
R55218 DVSS.n173 DVSS.n152 4.5005
R55219 DVSS.n6460 DVSS.n173 4.5005
R55220 DVSS.n161 DVSS.n153 4.5005
R55221 DVSS.n6460 DVSS.n161 4.5005
R55222 DVSS.n175 DVSS.n153 4.5005
R55223 DVSS.n6456 DVSS.n175 4.5005
R55224 DVSS.n6460 DVSS.n175 4.5005
R55225 DVSS.n6460 DVSS.n160 4.5005
R55226 DVSS.n6456 DVSS.n160 4.5005
R55227 DVSS.n160 DVSS.n152 4.5005
R55228 DVSS.n177 DVSS.n152 4.5005
R55229 DVSS.n6460 DVSS.n177 4.5005
R55230 DVSS.n159 DVSS.n153 4.5005
R55231 DVSS.n6460 DVSS.n159 4.5005
R55232 DVSS.n6446 DVSS.n153 4.5005
R55233 DVSS.n6456 DVSS.n6446 4.5005
R55234 DVSS.n6460 DVSS.n6446 4.5005
R55235 DVSS.n6460 DVSS.n158 4.5005
R55236 DVSS.n6456 DVSS.n158 4.5005
R55237 DVSS.n158 DVSS.n152 4.5005
R55238 DVSS.n6448 DVSS.n152 4.5005
R55239 DVSS.n6460 DVSS.n6448 4.5005
R55240 DVSS.n157 DVSS.n153 4.5005
R55241 DVSS.n6460 DVSS.n157 4.5005
R55242 DVSS.n6458 DVSS.n153 4.5005
R55243 DVSS.n6460 DVSS.n6458 4.5005
R55244 DVSS.n156 DVSS.n153 4.5005
R55245 DVSS.n6460 DVSS.n156 4.5005
R55246 DVSS.n153 DVSS.n141 4.5005
R55247 DVSS.n6456 DVSS.n141 4.5005
R55248 DVSS.n6460 DVSS.n141 4.5005
R55249 DVSS.n6460 DVSS.n144 4.5005
R55250 DVSS.n6456 DVSS.n144 4.5005
R55251 DVSS.n153 DVSS.n144 4.5005
R55252 DVSS.n152 DVSS.n144 4.5005
R55253 DVSS.n6460 DVSS.n149 4.5005
R55254 DVSS.n6456 DVSS.n149 4.5005
R55255 DVSS.n153 DVSS.n149 4.5005
R55256 DVSS.n152 DVSS.n149 4.5005
R55257 DVSS.n6461 DVSS.n152 4.5005
R55258 DVSS.n6461 DVSS.n153 4.5005
R55259 DVSS.n6461 DVSS.n6460 4.5005
R55260 DVSS.n6459 DVSS.n152 4.5005
R55261 DVSS.n6459 DVSS.n153 4.5005
R55262 DVSS.n6460 DVSS.n6459 4.5005
R55263 DVSS.n280 DVSS.n207 4.5005
R55264 DVSS.n6382 DVSS.n207 4.5005
R55265 DVSS.n6439 DVSS.n192 4.5005
R55266 DVSS.n6439 DVSS.n195 4.5005
R55267 DVSS.n6439 DVSS.n190 4.5005
R55268 DVSS.n6439 DVSS.n196 4.5005
R55269 DVSS.n6439 DVSS.n188 4.5005
R55270 DVSS.n6439 DVSS.n181 4.5005
R55271 DVSS.n6440 DVSS.n6439 4.5005
R55272 DVSS.n6439 DVSS.n197 4.5005
R55273 DVSS.n207 DVSS.n184 4.5005
R55274 DVSS.n6439 DVSS.n184 4.5005
R55275 DVSS.n207 DVSS.n198 4.5005
R55276 DVSS.n6439 DVSS.n198 4.5005
R55277 DVSS.n6397 DVSS.n6381 4.5005
R55278 DVSS.n6397 DVSS.n6393 4.5005
R55279 DVSS.n6400 DVSS.n257 4.5005
R55280 DVSS.n6400 DVSS.n270 4.5005
R55281 DVSS.n6400 DVSS.n255 4.5005
R55282 DVSS.n6400 DVSS.n247 4.5005
R55283 DVSS.n6401 DVSS.n6400 4.5005
R55284 DVSS.n6400 DVSS.n271 4.5005
R55285 DVSS.n6400 DVSS.n252 4.5005
R55286 DVSS.n6400 DVSS.n211 4.5005
R55287 DVSS.n6397 DVSS.n212 4.5005
R55288 DVSS.n6400 DVSS.n212 4.5005
R55289 DVSS.n6397 DVSS.n272 4.5005
R55290 DVSS.n6400 DVSS.n272 4.5005
R55291 DVSS.n6486 DVSS.n72 4.5005
R55292 DVSS.n6489 DVSS.n59 4.5005
R55293 DVSS.n6486 DVSS.n75 4.5005
R55294 DVSS.n6486 DVSS.n70 4.5005
R55295 DVSS.n6486 DVSS.n76 4.5005
R55296 DVSS.n6486 DVSS.n68 4.5005
R55297 DVSS.n6486 DVSS.n6484 4.5005
R55298 DVSS.n6489 DVSS.n63 4.5005
R55299 DVSS.n6489 DVSS.n53 4.5005
R55300 DVSS.n6489 DVSS.n48 4.5005
R55301 DVSS.n6490 DVSS.n6489 4.5005
R55302 DVSS.n6489 DVSS.n6488 4.5005
R55303 DVSS.n6479 DVSS.n87 4.5005
R55304 DVSS.n6476 DVSS.n101 4.5005
R55305 DVSS.n6479 DVSS.n91 4.5005
R55306 DVSS.n6479 DVSS.n85 4.5005
R55307 DVSS.n6479 DVSS.n92 4.5005
R55308 DVSS.n6479 DVSS.n78 4.5005
R55309 DVSS.n6480 DVSS.n6479 4.5005
R55310 DVSS.n6476 DVSS.n105 4.5005
R55311 DVSS.n6476 DVSS.n96 4.5005
R55312 DVSS.n6476 DVSS.n106 4.5005
R55313 DVSS.n6477 DVSS.n6476 4.5005
R55314 DVSS.n6476 DVSS.n6475 4.5005
R55315 DVSS.n6371 DVSS.n298 4.5005
R55316 DVSS.n298 DVSS.n284 4.5005
R55317 DVSS.n6373 DVSS.n298 4.5005
R55318 DVSS.n301 DVSS.n284 4.5005
R55319 DVSS.n6373 DVSS.n301 4.5005
R55320 DVSS.n297 DVSS.n284 4.5005
R55321 DVSS.n6373 DVSS.n297 4.5005
R55322 DVSS.n303 DVSS.n284 4.5005
R55323 DVSS.n6373 DVSS.n303 4.5005
R55324 DVSS.n6373 DVSS.n296 4.5005
R55325 DVSS.n6371 DVSS.n305 4.5005
R55326 DVSS.n305 DVSS.n284 4.5005
R55327 DVSS.n6373 DVSS.n305 4.5005
R55328 DVSS.n294 DVSS.n284 4.5005
R55329 DVSS.n6373 DVSS.n294 4.5005
R55330 DVSS.n307 DVSS.n284 4.5005
R55331 DVSS.n6373 DVSS.n307 4.5005
R55332 DVSS.n6371 DVSS.n293 4.5005
R55333 DVSS.n293 DVSS.n284 4.5005
R55334 DVSS.n6373 DVSS.n293 4.5005
R55335 DVSS.n6371 DVSS.n309 4.5005
R55336 DVSS.n309 DVSS.n284 4.5005
R55337 DVSS.n6373 DVSS.n309 4.5005
R55338 DVSS.n292 DVSS.n284 4.5005
R55339 DVSS.n6373 DVSS.n292 4.5005
R55340 DVSS.n311 DVSS.n284 4.5005
R55341 DVSS.n6373 DVSS.n311 4.5005
R55342 DVSS.n6371 DVSS.n291 4.5005
R55343 DVSS.n291 DVSS.n284 4.5005
R55344 DVSS.n6373 DVSS.n291 4.5005
R55345 DVSS.n6371 DVSS.n313 4.5005
R55346 DVSS.n313 DVSS.n284 4.5005
R55347 DVSS.n6373 DVSS.n313 4.5005
R55348 DVSS.n290 DVSS.n284 4.5005
R55349 DVSS.n6373 DVSS.n290 4.5005
R55350 DVSS.n314 DVSS.n284 4.5005
R55351 DVSS.n314 DVSS.n283 4.5005
R55352 DVSS.n6373 DVSS.n314 4.5005
R55353 DVSS.n6373 DVSS.n289 4.5005
R55354 DVSS.n289 DVSS.n283 4.5005
R55355 DVSS.n6371 DVSS.n289 4.5005
R55356 DVSS.n6371 DVSS.n317 4.5005
R55357 DVSS.n6373 DVSS.n317 4.5005
R55358 DVSS.n288 DVSS.n284 4.5005
R55359 DVSS.n6373 DVSS.n288 4.5005
R55360 DVSS.n318 DVSS.n284 4.5005
R55361 DVSS.n318 DVSS.n283 4.5005
R55362 DVSS.n6373 DVSS.n318 4.5005
R55363 DVSS.n6373 DVSS.n287 4.5005
R55364 DVSS.n287 DVSS.n283 4.5005
R55365 DVSS.n6371 DVSS.n287 4.5005
R55366 DVSS.n6372 DVSS.n6371 4.5005
R55367 DVSS.n6373 DVSS.n6372 4.5005
R55368 DVSS.n286 DVSS.n284 4.5005
R55369 DVSS.n6373 DVSS.n286 4.5005
R55370 DVSS.n6374 DVSS.n284 4.5005
R55371 DVSS.n6374 DVSS.n283 4.5005
R55372 DVSS.n6374 DVSS.n6373 4.5005
R55373 DVSS.n6294 DVSS.n6259 4.5005
R55374 DVSS.n6297 DVSS.n363 4.5005
R55375 DVSS.n6294 DVSS.n6273 4.5005
R55376 DVSS.n6294 DVSS.n384 4.5005
R55377 DVSS.n6294 DVSS.n6284 4.5005
R55378 DVSS.n6294 DVSS.n382 4.5005
R55379 DVSS.n6294 DVSS.n6291 4.5005
R55380 DVSS.n6297 DVSS.n378 4.5005
R55381 DVSS.n6297 DVSS.n357 4.5005
R55382 DVSS.n6297 DVSS.n379 4.5005
R55383 DVSS.n6297 DVSS.n355 4.5005
R55384 DVSS.n6297 DVSS.n6296 4.5005
R55385 DVSS.n6500 DVSS.n29 4.5005
R55386 DVSS.n6262 DVSS.n15 4.5005
R55387 DVSS.n6500 DVSS.n36 4.5005
R55388 DVSS.n6500 DVSS.n26 4.5005
R55389 DVSS.n6500 DVSS.n38 4.5005
R55390 DVSS.n6500 DVSS.n23 4.5005
R55391 DVSS.n6500 DVSS.n40 4.5005
R55392 DVSS.n366 DVSS.n15 4.5005
R55393 DVSS.n367 DVSS.n15 4.5005
R55394 DVSS.n44 DVSS.n15 4.5005
R55395 DVSS.n6498 DVSS.n15 4.5005
R55396 DVSS.n279 DVSS.n15 4.5005
R55397 DVSS.n6241 DVSS.n403 4.5005
R55398 DVSS.n6241 DVSS.n407 4.5005
R55399 DVSS.n6241 DVSS.n401 4.5005
R55400 DVSS.n6241 DVSS.n409 4.5005
R55401 DVSS.n6238 DVSS.n6237 4.5005
R55402 DVSS.n6241 DVSS.n399 4.5005
R55403 DVSS.n6241 DVSS.n410 4.5005
R55404 DVSS.n6241 DVSS.n398 4.5005
R55405 DVSS.n6241 DVSS.n411 4.5005
R55406 DVSS.n6242 DVSS.n6241 4.5005
R55407 DVSS.n6238 DVSS.n413 4.5005
R55408 DVSS.n6241 DVSS.n395 4.5005
R55409 DVSS.n6229 DVSS.n448 4.5005
R55410 DVSS.n6229 DVSS.n451 4.5005
R55411 DVSS.n6229 DVSS.n446 4.5005
R55412 DVSS.n6229 DVSS.n453 4.5005
R55413 DVSS.n6233 DVSS.n6232 4.5005
R55414 DVSS.n6229 DVSS.n445 4.5005
R55415 DVSS.n6229 DVSS.n454 4.5005
R55416 DVSS.n6229 DVSS.n444 4.5005
R55417 DVSS.n6229 DVSS.n6227 4.5005
R55418 DVSS.n6229 DVSS.n443 4.5005
R55419 DVSS.n6232 DVSS.n429 4.5005
R55420 DVSS.n6229 DVSS.n6228 4.5005
R55421 DVSS.n474 DVSS.n465 4.5005
R55422 DVSS.n6199 DVSS.n474 4.5005
R55423 DVSS.n477 DVSS.n465 4.5005
R55424 DVSS.n6199 DVSS.n477 4.5005
R55425 DVSS.n6199 DVSS.n457 4.5005
R55426 DVSS.n479 DVSS.n465 4.5005
R55427 DVSS.n6199 DVSS.n479 4.5005
R55428 DVSS.n473 DVSS.n465 4.5005
R55429 DVSS.n6199 DVSS.n473 4.5005
R55430 DVSS.n6200 DVSS.n465 4.5005
R55431 DVSS.n6200 DVSS.n462 4.5005
R55432 DVSS.n6200 DVSS.n6199 4.5005
R55433 DVSS.n472 DVSS.n465 4.5005
R55434 DVSS.n6199 DVSS.n472 4.5005
R55435 DVSS.n481 DVSS.n465 4.5005
R55436 DVSS.n6199 DVSS.n481 4.5005
R55437 DVSS.n471 DVSS.n465 4.5005
R55438 DVSS.n471 DVSS.n462 4.5005
R55439 DVSS.n6199 DVSS.n471 4.5005
R55440 DVSS.n483 DVSS.n465 4.5005
R55441 DVSS.n6199 DVSS.n483 4.5005
R55442 DVSS.n470 DVSS.n465 4.5005
R55443 DVSS.n6199 DVSS.n470 4.5005
R55444 DVSS.n484 DVSS.n465 4.5005
R55445 DVSS.n484 DVSS.n462 4.5005
R55446 DVSS.n6199 DVSS.n484 4.5005
R55447 DVSS.n469 DVSS.n465 4.5005
R55448 DVSS.n6199 DVSS.n469 4.5005
R55449 DVSS.n6196 DVSS.n486 4.5005
R55450 DVSS.n486 DVSS.n465 4.5005
R55451 DVSS.n6199 DVSS.n486 4.5005
R55452 DVSS.n468 DVSS.n465 4.5005
R55453 DVSS.n468 DVSS.n462 4.5005
R55454 DVSS.n6199 DVSS.n468 4.5005
R55455 DVSS.n487 DVSS.n465 4.5005
R55456 DVSS.n487 DVSS.n462 4.5005
R55457 DVSS.n6199 DVSS.n487 4.5005
R55458 DVSS.n465 DVSS.n461 4.5005
R55459 DVSS.n462 DVSS.n461 4.5005
R55460 DVSS.n6199 DVSS.n461 4.5005
R55461 DVSS.n465 DVSS.n456 4.5005
R55462 DVSS.n462 DVSS.n456 4.5005
R55463 DVSS.n6199 DVSS.n456 4.5005
R55464 DVSS.n467 DVSS.n462 4.5005
R55465 DVSS.n6199 DVSS.n467 4.5005
R55466 DVSS.n6199 DVSS.n488 4.5005
R55467 DVSS.n488 DVSS.n462 4.5005
R55468 DVSS.n6196 DVSS.n488 4.5005
R55469 DVSS.n6194 DVSS.n462 4.5005
R55470 DVSS.n6196 DVSS.n6194 4.5005
R55471 DVSS.n512 DVSS.n462 4.5005
R55472 DVSS.n6196 DVSS.n512 4.5005
R55473 DVSS.n6197 DVSS.n462 4.5005
R55474 DVSS.n6197 DVSS.n6196 4.5005
R55475 DVSS.n509 DVSS.n462 4.5005
R55476 DVSS.n509 DVSS.n465 4.5005
R55477 DVSS.n6196 DVSS.n509 4.5005
R55478 DVSS.n467 DVSS.n465 4.5005
R55479 DVSS.n6218 DVSS.n390 4.5005
R55480 DVSS.n6210 DVSS.n390 4.5005
R55481 DVSS.n1121 DVSS.n390 4.5005
R55482 DVSS.n1127 DVSS.n390 4.5005
R55483 DVSS.n1132 DVSS.n389 4.5005
R55484 DVSS.n1129 DVSS.n390 4.5005
R55485 DVSS.n1123 DVSS.n390 4.5005
R55486 DVSS.n459 DVSS.n390 4.5005
R55487 DVSS.n6214 DVSS.n390 4.5005
R55488 DVSS.n6250 DVSS.n390 4.5005
R55489 DVSS.n6255 DVSS.n389 4.5005
R55490 DVSS.n391 DVSS.n390 4.5005
R55491 DVSS.n1085 DVSS.n1071 4.5005
R55492 DVSS.n1088 DVSS.n1071 4.5005
R55493 DVSS.n1108 DVSS.n1071 4.5005
R55494 DVSS.n1097 DVSS.n1071 4.5005
R55495 DVSS.n6131 DVSS.n6125 4.5005
R55496 DVSS.n1096 DVSS.n1071 4.5005
R55497 DVSS.n1107 DVSS.n1071 4.5005
R55498 DVSS.n1078 DVSS.n1071 4.5005
R55499 DVSS.n1080 DVSS.n1071 4.5005
R55500 DVSS.n6126 DVSS.n1071 4.5005
R55501 DVSS.n6131 DVSS.n1075 4.5005
R55502 DVSS.n1082 DVSS.n1071 4.5005
R55503 DVSS.n3085 DVSS.n3084 4.17693
R55504 DVSS.n4426 DVSS.n3893 3.91226
R55505 DVSS.n4426 DVSS.n3894 3.91226
R55506 DVSS.n4422 DVSS.n3894 3.91226
R55507 DVSS.n4422 DVSS.n3957 3.91226
R55508 DVSS.n4414 DVSS.n3957 3.91226
R55509 DVSS.n4414 DVSS.n3965 3.91226
R55510 DVSS.n4410 DVSS.n3965 3.91226
R55511 DVSS.n4410 DVSS.n3967 3.91226
R55512 DVSS.n4402 DVSS.n3967 3.91226
R55513 DVSS.n4402 DVSS.n3975 3.91226
R55514 DVSS.n4398 DVSS.n3975 3.91226
R55515 DVSS.n4398 DVSS.n3977 3.91226
R55516 DVSS.n4390 DVSS.n3977 3.91226
R55517 DVSS.n4390 DVSS.n3985 3.91226
R55518 DVSS.n4386 DVSS.n3985 3.91226
R55519 DVSS.n4386 DVSS.n3987 3.91226
R55520 DVSS.n4378 DVSS.n3987 3.91226
R55521 DVSS.n4378 DVSS.n3995 3.91226
R55522 DVSS.n4374 DVSS.n3995 3.91226
R55523 DVSS.n4374 DVSS.n3998 3.91226
R55524 DVSS.n3998 DVSS.n1811 3.91226
R55525 DVSS.n4908 DVSS.n1811 3.91226
R55526 DVSS.n4908 DVSS.n1812 3.91226
R55527 DVSS.n4904 DVSS.n1812 3.91226
R55528 DVSS.n4904 DVSS.n1815 3.91226
R55529 DVSS.n4896 DVSS.n1815 3.91226
R55530 DVSS.n4896 DVSS.n1825 3.91226
R55531 DVSS.n4892 DVSS.n1825 3.91226
R55532 DVSS.n4892 DVSS.n1827 3.91226
R55533 DVSS.n4884 DVSS.n1827 3.91226
R55534 DVSS.n4884 DVSS.n1835 3.91226
R55535 DVSS.n4880 DVSS.n1835 3.91226
R55536 DVSS.n4880 DVSS.n1837 3.91226
R55537 DVSS.n4872 DVSS.n1837 3.91226
R55538 DVSS.n4872 DVSS.n1845 3.91226
R55539 DVSS.n4868 DVSS.n1845 3.91226
R55540 DVSS.n4868 DVSS.n1847 3.91226
R55541 DVSS.n4860 DVSS.n1847 3.91226
R55542 DVSS.n4860 DVSS.n1855 3.91226
R55543 DVSS.n4856 DVSS.n1855 3.91226
R55544 DVSS.n4856 DVSS.n1857 3.91226
R55545 DVSS.n1969 DVSS.n1857 3.91226
R55546 DVSS.n4750 DVSS.n1969 3.91226
R55547 DVSS.n4750 DVSS.n1881 3.91226
R55548 DVSS.n4845 DVSS.n1881 3.91226
R55549 DVSS.n4845 DVSS.n1882 3.91226
R55550 DVSS.n4841 DVSS.n1882 3.91226
R55551 DVSS.n4841 DVSS.n1885 3.91226
R55552 DVSS.n4833 DVSS.n1885 3.91226
R55553 DVSS.n4833 DVSS.n1894 3.91226
R55554 DVSS.n4829 DVSS.n1894 3.91226
R55555 DVSS.n4829 DVSS.n1896 3.91226
R55556 DVSS.n4821 DVSS.n1896 3.91226
R55557 DVSS.n4821 DVSS.n1904 3.91226
R55558 DVSS.n4817 DVSS.n1904 3.91226
R55559 DVSS.n4817 DVSS.n1906 3.91226
R55560 DVSS.n4809 DVSS.n1906 3.91226
R55561 DVSS.n4809 DVSS.n1914 3.91226
R55562 DVSS.n4805 DVSS.n1914 3.91226
R55563 DVSS.n4805 DVSS.n1916 3.91226
R55564 DVSS.n4797 DVSS.n1916 3.91226
R55565 DVSS.n4797 DVSS.n1924 3.91226
R55566 DVSS.n4793 DVSS.n1924 3.91226
R55567 DVSS.n4793 DVSS.n1926 3.91226
R55568 DVSS.n1926 DVSS.n1594 3.91226
R55569 DVSS.n5258 DVSS.n1594 3.91226
R55570 DVSS.n5258 DVSS.n1595 3.91226
R55571 DVSS.n5250 DVSS.n1595 3.91226
R55572 DVSS.n5250 DVSS.n1606 3.91226
R55573 DVSS.n5246 DVSS.n1606 3.91226
R55574 DVSS.n5246 DVSS.n1608 3.91226
R55575 DVSS.n5238 DVSS.n1608 3.91226
R55576 DVSS.n5238 DVSS.n1616 3.91226
R55577 DVSS.n5234 DVSS.n1616 3.91226
R55578 DVSS.n5234 DVSS.n1618 3.91226
R55579 DVSS.n5226 DVSS.n1618 3.91226
R55580 DVSS.n5226 DVSS.n1626 3.91226
R55581 DVSS.n5222 DVSS.n1626 3.91226
R55582 DVSS.n5222 DVSS.n1628 3.91226
R55583 DVSS.n5214 DVSS.n1628 3.91226
R55584 DVSS.n5214 DVSS.n1636 3.91226
R55585 DVSS.n5210 DVSS.n1636 3.91226
R55586 DVSS.n5210 DVSS.n1638 3.91226
R55587 DVSS.n5202 DVSS.n1638 3.91226
R55588 DVSS.n5202 DVSS.n5199 3.91226
R55589 DVSS.n5199 DVSS.n1372 3.91226
R55590 DVSS.n5504 DVSS.n1372 3.91226
R55591 DVSS.n4428 DVSS.n3888 3.91226
R55592 DVSS.n4428 DVSS.n3889 3.91226
R55593 DVSS.n4420 DVSS.n3889 3.91226
R55594 DVSS.n4420 DVSS.n3960 3.91226
R55595 DVSS.n4416 DVSS.n3960 3.91226
R55596 DVSS.n4416 DVSS.n3962 3.91226
R55597 DVSS.n4408 DVSS.n3962 3.91226
R55598 DVSS.n4408 DVSS.n3970 3.91226
R55599 DVSS.n4404 DVSS.n3970 3.91226
R55600 DVSS.n4404 DVSS.n3972 3.91226
R55601 DVSS.n4396 DVSS.n3972 3.91226
R55602 DVSS.n4396 DVSS.n3980 3.91226
R55603 DVSS.n4392 DVSS.n3980 3.91226
R55604 DVSS.n4392 DVSS.n3982 3.91226
R55605 DVSS.n4384 DVSS.n3982 3.91226
R55606 DVSS.n4384 DVSS.n3990 3.91226
R55607 DVSS.n4380 DVSS.n3990 3.91226
R55608 DVSS.n4380 DVSS.n3992 3.91226
R55609 DVSS.n4372 DVSS.n3992 3.91226
R55610 DVSS.n4372 DVSS.n4362 3.91226
R55611 DVSS.n4368 DVSS.n4362 3.91226
R55612 DVSS.n4368 DVSS.n1810 3.91226
R55613 DVSS.n1818 DVSS.n1810 3.91226
R55614 DVSS.n4902 DVSS.n1818 3.91226
R55615 DVSS.n4902 DVSS.n1819 3.91226
R55616 DVSS.n4898 DVSS.n1819 3.91226
R55617 DVSS.n4898 DVSS.n1822 3.91226
R55618 DVSS.n4890 DVSS.n1822 3.91226
R55619 DVSS.n4890 DVSS.n1830 3.91226
R55620 DVSS.n4886 DVSS.n1830 3.91226
R55621 DVSS.n4886 DVSS.n1832 3.91226
R55622 DVSS.n4878 DVSS.n1832 3.91226
R55623 DVSS.n4878 DVSS.n1840 3.91226
R55624 DVSS.n4874 DVSS.n1840 3.91226
R55625 DVSS.n4874 DVSS.n1842 3.91226
R55626 DVSS.n4866 DVSS.n1842 3.91226
R55627 DVSS.n4866 DVSS.n1850 3.91226
R55628 DVSS.n4862 DVSS.n1850 3.91226
R55629 DVSS.n4862 DVSS.n1852 3.91226
R55630 DVSS.n4854 DVSS.n1852 3.91226
R55631 DVSS.n4854 DVSS.n1860 3.91226
R55632 DVSS.n1963 DVSS.n1860 3.91226
R55633 DVSS.n1968 DVSS.n1963 3.91226
R55634 DVSS.n1968 DVSS.n1876 3.91226
R55635 DVSS.n4847 DVSS.n1876 3.91226
R55636 DVSS.n4847 DVSS.n1877 3.91226
R55637 DVSS.n4839 DVSS.n1877 3.91226
R55638 DVSS.n4839 DVSS.n1888 3.91226
R55639 DVSS.n4835 DVSS.n1888 3.91226
R55640 DVSS.n4835 DVSS.n1891 3.91226
R55641 DVSS.n4827 DVSS.n1891 3.91226
R55642 DVSS.n4827 DVSS.n1899 3.91226
R55643 DVSS.n4823 DVSS.n1899 3.91226
R55644 DVSS.n4823 DVSS.n1901 3.91226
R55645 DVSS.n4815 DVSS.n1901 3.91226
R55646 DVSS.n4815 DVSS.n1909 3.91226
R55647 DVSS.n4811 DVSS.n1909 3.91226
R55648 DVSS.n4811 DVSS.n1911 3.91226
R55649 DVSS.n4803 DVSS.n1911 3.91226
R55650 DVSS.n4803 DVSS.n1919 3.91226
R55651 DVSS.n4799 DVSS.n1919 3.91226
R55652 DVSS.n4799 DVSS.n1921 3.91226
R55653 DVSS.n4791 DVSS.n1921 3.91226
R55654 DVSS.n4791 DVSS.n4784 3.91226
R55655 DVSS.n4784 DVSS.n1599 3.91226
R55656 DVSS.n5256 DVSS.n1599 3.91226
R55657 DVSS.n5256 DVSS.n1600 3.91226
R55658 DVSS.n5252 DVSS.n1600 3.91226
R55659 DVSS.n5252 DVSS.n1603 3.91226
R55660 DVSS.n5244 DVSS.n1603 3.91226
R55661 DVSS.n5244 DVSS.n1611 3.91226
R55662 DVSS.n5240 DVSS.n1611 3.91226
R55663 DVSS.n5240 DVSS.n1613 3.91226
R55664 DVSS.n5232 DVSS.n1613 3.91226
R55665 DVSS.n5232 DVSS.n1621 3.91226
R55666 DVSS.n5228 DVSS.n1621 3.91226
R55667 DVSS.n5228 DVSS.n1623 3.91226
R55668 DVSS.n5220 DVSS.n1623 3.91226
R55669 DVSS.n5220 DVSS.n1631 3.91226
R55670 DVSS.n5216 DVSS.n1631 3.91226
R55671 DVSS.n5216 DVSS.n1633 3.91226
R55672 DVSS.n5208 DVSS.n1633 3.91226
R55673 DVSS.n5208 DVSS.n1641 3.91226
R55674 DVSS.n5204 DVSS.n1641 3.91226
R55675 DVSS.n5204 DVSS.n1644 3.91226
R55676 DVSS.n1644 DVSS.n1377 3.91226
R55677 DVSS.n5502 DVSS.n1377 3.91226
R55678 DVSS.n4330 DVSS.n3892 3.91226
R55679 DVSS.n4334 DVSS.n3892 3.91226
R55680 DVSS.n4334 DVSS.n3959 3.91226
R55681 DVSS.n4337 DVSS.n3959 3.91226
R55682 DVSS.n4337 DVSS.n3964 3.91226
R55683 DVSS.n4340 DVSS.n3964 3.91226
R55684 DVSS.n4340 DVSS.n3969 3.91226
R55685 DVSS.n4343 DVSS.n3969 3.91226
R55686 DVSS.n4343 DVSS.n3974 3.91226
R55687 DVSS.n4346 DVSS.n3974 3.91226
R55688 DVSS.n4346 DVSS.n3979 3.91226
R55689 DVSS.n4349 DVSS.n3979 3.91226
R55690 DVSS.n4349 DVSS.n3984 3.91226
R55691 DVSS.n4352 DVSS.n3984 3.91226
R55692 DVSS.n4352 DVSS.n3989 3.91226
R55693 DVSS.n4355 DVSS.n3989 3.91226
R55694 DVSS.n4355 DVSS.n3994 3.91226
R55695 DVSS.n4000 DVSS.n3994 3.91226
R55696 DVSS.n4361 DVSS.n4000 3.91226
R55697 DVSS.n4361 DVSS.n4001 3.91226
R55698 DVSS.n4001 DVSS.n1806 3.91226
R55699 DVSS.n4910 DVSS.n1806 3.91226
R55700 DVSS.n4910 DVSS.n1807 3.91226
R55701 DVSS.n1817 DVSS.n1807 3.91226
R55702 DVSS.n1934 DVSS.n1817 3.91226
R55703 DVSS.n1934 DVSS.n1824 3.91226
R55704 DVSS.n1937 DVSS.n1824 3.91226
R55705 DVSS.n1937 DVSS.n1829 3.91226
R55706 DVSS.n1940 DVSS.n1829 3.91226
R55707 DVSS.n1940 DVSS.n1834 3.91226
R55708 DVSS.n1943 DVSS.n1834 3.91226
R55709 DVSS.n1943 DVSS.n1839 3.91226
R55710 DVSS.n1946 DVSS.n1839 3.91226
R55711 DVSS.n1946 DVSS.n1844 3.91226
R55712 DVSS.n1949 DVSS.n1844 3.91226
R55713 DVSS.n1949 DVSS.n1849 3.91226
R55714 DVSS.n1952 DVSS.n1849 3.91226
R55715 DVSS.n1952 DVSS.n1854 3.91226
R55716 DVSS.n1955 DVSS.n1854 3.91226
R55717 DVSS.n1955 DVSS.n1859 3.91226
R55718 DVSS.n1958 DVSS.n1859 3.91226
R55719 DVSS.n1958 DVSS.n1932 3.91226
R55720 DVSS.n4752 DVSS.n1932 3.91226
R55721 DVSS.n4753 DVSS.n4752 3.91226
R55722 DVSS.n4753 DVSS.n1880 3.91226
R55723 DVSS.n4756 DVSS.n1880 3.91226
R55724 DVSS.n4756 DVSS.n1887 3.91226
R55725 DVSS.n4759 DVSS.n1887 3.91226
R55726 DVSS.n4759 DVSS.n1893 3.91226
R55727 DVSS.n4762 DVSS.n1893 3.91226
R55728 DVSS.n4762 DVSS.n1898 3.91226
R55729 DVSS.n4765 DVSS.n1898 3.91226
R55730 DVSS.n4765 DVSS.n1903 3.91226
R55731 DVSS.n4768 DVSS.n1903 3.91226
R55732 DVSS.n4768 DVSS.n1908 3.91226
R55733 DVSS.n4771 DVSS.n1908 3.91226
R55734 DVSS.n4771 DVSS.n1913 3.91226
R55735 DVSS.n4774 DVSS.n1913 3.91226
R55736 DVSS.n4774 DVSS.n1918 3.91226
R55737 DVSS.n4777 DVSS.n1918 3.91226
R55738 DVSS.n4777 DVSS.n1923 3.91226
R55739 DVSS.n1928 DVSS.n1923 3.91226
R55740 DVSS.n4783 DVSS.n1928 3.91226
R55741 DVSS.n4783 DVSS.n1930 3.91226
R55742 DVSS.n1930 DVSS.n1929 3.91226
R55743 DVSS.n1929 DVSS.n1598 3.91226
R55744 DVSS.n5171 DVSS.n1598 3.91226
R55745 DVSS.n5171 DVSS.n1605 3.91226
R55746 DVSS.n5174 DVSS.n1605 3.91226
R55747 DVSS.n5174 DVSS.n1610 3.91226
R55748 DVSS.n5177 DVSS.n1610 3.91226
R55749 DVSS.n5177 DVSS.n1615 3.91226
R55750 DVSS.n5180 DVSS.n1615 3.91226
R55751 DVSS.n5180 DVSS.n1620 3.91226
R55752 DVSS.n5183 DVSS.n1620 3.91226
R55753 DVSS.n5183 DVSS.n1625 3.91226
R55754 DVSS.n5186 DVSS.n1625 3.91226
R55755 DVSS.n5186 DVSS.n1630 3.91226
R55756 DVSS.n5189 DVSS.n1630 3.91226
R55757 DVSS.n5189 DVSS.n1635 3.91226
R55758 DVSS.n5192 DVSS.n1635 3.91226
R55759 DVSS.n5192 DVSS.n1640 3.91226
R55760 DVSS.n1646 DVSS.n1640 3.91226
R55761 DVSS.n5198 DVSS.n1646 3.91226
R55762 DVSS.n5198 DVSS.n1648 3.91226
R55763 DVSS.n1648 DVSS.n1647 3.91226
R55764 DVSS.n1647 DVSS.n1376 3.91226
R55765 DVSS.n4317 DVSS.n4005 3.83228
R55766 DVSS.n4318 DVSS.n4317 3.83228
R55767 DVSS.n4745 DVSS.n1591 3.81164
R55768 DVSS.n3519 DVSS.n2133 3.70786
R55769 DVSS.n3069 DVSS.n3068 3.70786
R55770 DVSS.n5394 DVSS.n5393 3.39586
R55771 DVSS.n5395 DVSS.n5394 3.39586
R55772 DVSS.n3067 DVSS.n3066 3.1804
R55773 DVSS.n4746 DVSS.n4745 3.14175
R55774 DVSS.n1519 DVSS.n1518 3.12476
R55775 DVSS.n1522 DVSS.n1519 3.12476
R55776 DVSS.n3064 DVSS.n3063 3.11878
R55777 DVSS.n3068 DVSS.n3067 3.11084
R55778 DVSS.n3063 DVSS.n2133 3.11084
R55779 DVSS.n5595 DVSS.n5594 3.10905
R55780 DVSS.n5660 DVSS.n1285 3.10905
R55781 DVSS.n4642 DVSS.n1283 2.99652
R55782 DVSS.n5604 DVSS.n5603 2.87501
R55783 DVSS.n5610 DVSS.n5609 2.87501
R55784 DVSS.n5615 DVSS.n5613 2.87501
R55785 DVSS.n5621 DVSS.n5620 2.87501
R55786 DVSS.n5627 DVSS.n5626 2.87501
R55787 DVSS.n5632 DVSS.n5630 2.87501
R55788 DVSS.n5638 DVSS.n5637 2.87501
R55789 DVSS.n5642 DVSS.n5641 2.87501
R55790 DVSS.n5707 DVSS.n5706 2.87501
R55791 DVSS.n1245 DVSS.n1244 2.87501
R55792 DVSS.n5693 DVSS.n5692 2.87501
R55793 DVSS.n5730 DVSS.n5729 2.87501
R55794 DVSS.n5734 DVSS.n5733 2.87501
R55795 DVSS.n1225 DVSS.n1224 2.87501
R55796 DVSS.n5747 DVSS.n5746 2.87501
R55797 DVSS.n5751 DVSS.n5750 2.87501
R55798 DVSS.n1212 DVSS.n1211 2.87501
R55799 DVSS.n5767 DVSS.n5766 2.87501
R55800 DVSS.n5772 DVSS.n5770 2.87501
R55801 DVSS.n6067 DVSS.n6066 2.87501
R55802 DVSS.n6057 DVSS.n6055 2.87501
R55803 DVSS.n5785 DVSS.n5783 2.87501
R55804 DVSS.n6112 DVSS.n6111 2.87501
R55805 DVSS.n6117 DVSS.n6115 2.87501
R55806 DVSS.n6122 DVSS.n6121 2.87501
R55807 DVSS.n1106 DVSS.n1105 2.87501
R55808 DVSS.n1117 DVSS.n1116 2.87501
R55809 DVSS.n6208 DVSS.n6207 2.87501
R55810 DVSS.n6221 DVSS.n6220 2.87501
R55811 DVSS.n6248 DVSS.n6247 2.87501
R55812 DVSS.n6271 DVSS.n6270 2.87501
R55813 DVSS.n6282 DVSS.n6281 2.87501
R55814 DVSS.n6289 DVSS.n6288 2.87501
R55815 DVSS.n376 DVSS.n375 2.87501
R55816 DVSS.n6496 DVSS.n6495 2.87501
R55817 DVSS.n6379 DVSS.n6378 2.87501
R55818 DVSS.n6391 DVSS.n6390 2.87501
R55819 DVSS.n268 DVSS.n267 2.87501
R55820 DVSS.n6405 DVSS.n6404 2.87501
R55821 DVSS.n6444 DVSS.n6442 2.87501
R55822 DVSS.n5601 DVSS.n1301 2.81339
R55823 DVSS.n5607 DVSS.n1302 2.81339
R55824 DVSS.n1329 DVSS.n1303 2.81339
R55825 DVSS.n5618 DVSS.n1304 2.81339
R55826 DVSS.n5624 DVSS.n1305 2.81339
R55827 DVSS.n1325 DVSS.n1306 2.81339
R55828 DVSS.n5635 DVSS.n1320 2.81339
R55829 DVSS.n5644 DVSS.n5643 2.81339
R55830 DVSS.n5710 DVSS.n5709 2.81339
R55831 DVSS.n5717 DVSS.n1236 2.81339
R55832 DVSS.n5723 DVSS.n1231 2.81339
R55833 DVSS.n5727 DVSS.n5726 2.81339
R55834 DVSS.n5737 DVSS.n5736 2.81339
R55835 DVSS.n5740 DVSS.n1218 2.81339
R55836 DVSS.n5744 DVSS.n5743 2.81339
R55837 DVSS.n5754 DVSS.n5753 2.81339
R55838 DVSS.n5757 DVSS.n1205 2.81339
R55839 DVSS.n5764 DVSS.n5763 2.81339
R55840 DVSS.n5760 DVSS.n1200 2.81339
R55841 DVSS.n6064 DVSS.n6063 2.81339
R55842 DVSS.n6096 DVSS.n1156 2.81339
R55843 DVSS.n6105 DVSS.n1141 2.81339
R55844 DVSS.n6109 DVSS.n6108 2.81339
R55845 DVSS.n1136 DVSS.n1135 2.81339
R55846 DVSS.n6235 DVSS.n425 2.81339
R55847 DVSS.n1103 DVSS.n1102 2.81339
R55848 DVSS.n1114 DVSS.n1113 2.81339
R55849 DVSS.n6205 DVSS.n6204 2.81339
R55850 DVSS.n6225 DVSS.n6223 2.81339
R55851 DVSS.n6245 DVSS.n6244 2.81339
R55852 DVSS.n6268 DVSS.n6267 2.81339
R55853 DVSS.n6279 DVSS.n6278 2.81339
R55854 DVSS.n6482 DVSS.n77 2.81339
R55855 DVSS.n373 DVSS.n372 2.81339
R55856 DVSS.n6493 DVSS.n6492 2.81339
R55857 DVSS.n6376 DVSS.n107 2.81339
R55858 DVSS.n6388 DVSS.n6387 2.81339
R55859 DVSS.n265 DVSS.n264 2.81339
R55860 DVSS.n6409 DVSS.n6407 2.81339
R55861 DVSS.n6414 DVSS.n179 2.81339
R55862 DVSS.n5348 DVSS.n5347 2.69735
R55863 DVSS.n5168 DVSS.n5167 2.69735
R55864 DVSS.n4913 DVSS.n1803 2.69735
R55865 DVSS.n4431 DVSS.n3885 2.69735
R55866 DVSS.n5391 DVSS.n5390 2.62838
R55867 DVSS.n5354 DVSS.n5353 2.62838
R55868 DVSS.n5353 DVSS.n1522 2.62235
R55869 DVSS.n5398 DVSS.n5395 2.61801
R55870 DVSS.n5393 DVSS.n5390 2.61724
R55871 DVSS.n4325 DVSS.n4324 2.6005
R55872 DVSS.n4323 DVSS.n4322 2.6005
R55873 DVSS.n4320 DVSS.n4007 2.6005
R55874 DVSS.n4069 DVSS.n4008 2.6005
R55875 DVSS.n4072 DVSS.n4071 2.6005
R55876 DVSS.n4074 DVSS.n4073 2.6005
R55877 DVSS.n4077 DVSS.n4076 2.6005
R55878 DVSS.n4079 DVSS.n4078 2.6005
R55879 DVSS.n4082 DVSS.n4081 2.6005
R55880 DVSS.n4084 DVSS.n4083 2.6005
R55881 DVSS.n4087 DVSS.n4086 2.6005
R55882 DVSS.n4089 DVSS.n4088 2.6005
R55883 DVSS.n4092 DVSS.n4091 2.6005
R55884 DVSS.n4094 DVSS.n4093 2.6005
R55885 DVSS.n4097 DVSS.n4096 2.6005
R55886 DVSS.n4099 DVSS.n4098 2.6005
R55887 DVSS.n4102 DVSS.n4101 2.6005
R55888 DVSS.n4104 DVSS.n4103 2.6005
R55889 DVSS.n4107 DVSS.n4106 2.6005
R55890 DVSS.n4109 DVSS.n4108 2.6005
R55891 DVSS.n4112 DVSS.n4111 2.6005
R55892 DVSS.n4114 DVSS.n4113 2.6005
R55893 DVSS.n4117 DVSS.n4116 2.6005
R55894 DVSS.n4119 DVSS.n4118 2.6005
R55895 DVSS.n4122 DVSS.n4121 2.6005
R55896 DVSS.n4125 DVSS.n4124 2.6005
R55897 DVSS.n4128 DVSS.n4127 2.6005
R55898 DVSS.n4130 DVSS.n4129 2.6005
R55899 DVSS.n4133 DVSS.n4132 2.6005
R55900 DVSS.n4135 DVSS.n4134 2.6005
R55901 DVSS.n4138 DVSS.n4137 2.6005
R55902 DVSS.n4140 DVSS.n4139 2.6005
R55903 DVSS.n4143 DVSS.n4142 2.6005
R55904 DVSS.n4145 DVSS.n4144 2.6005
R55905 DVSS.n4148 DVSS.n4147 2.6005
R55906 DVSS.n4150 DVSS.n4149 2.6005
R55907 DVSS.n4153 DVSS.n4152 2.6005
R55908 DVSS.n4155 DVSS.n4154 2.6005
R55909 DVSS.n4158 DVSS.n4157 2.6005
R55910 DVSS.n4160 DVSS.n4159 2.6005
R55911 DVSS.n4163 DVSS.n4162 2.6005
R55912 DVSS.n4165 DVSS.n4164 2.6005
R55913 DVSS.n4168 DVSS.n4167 2.6005
R55914 DVSS.n4170 DVSS.n4169 2.6005
R55915 DVSS.n4173 DVSS.n4172 2.6005
R55916 DVSS.n4175 DVSS.n4174 2.6005
R55917 DVSS.n4178 DVSS.n4177 2.6005
R55918 DVSS.n4181 DVSS.n4180 2.6005
R55919 DVSS.n4192 DVSS.n4191 2.6005
R55920 DVSS.n4195 DVSS.n4194 2.6005
R55921 DVSS.n4197 DVSS.n4196 2.6005
R55922 DVSS.n4200 DVSS.n4199 2.6005
R55923 DVSS.n4202 DVSS.n4201 2.6005
R55924 DVSS.n4205 DVSS.n4204 2.6005
R55925 DVSS.n4207 DVSS.n4206 2.6005
R55926 DVSS.n4210 DVSS.n4209 2.6005
R55927 DVSS.n4212 DVSS.n4211 2.6005
R55928 DVSS.n4215 DVSS.n4214 2.6005
R55929 DVSS.n4217 DVSS.n4216 2.6005
R55930 DVSS.n4220 DVSS.n4219 2.6005
R55931 DVSS.n4222 DVSS.n4221 2.6005
R55932 DVSS.n4225 DVSS.n4224 2.6005
R55933 DVSS.n4227 DVSS.n4226 2.6005
R55934 DVSS.n4230 DVSS.n4229 2.6005
R55935 DVSS.n4232 DVSS.n4231 2.6005
R55936 DVSS.n4235 DVSS.n4234 2.6005
R55937 DVSS.n4237 DVSS.n4236 2.6005
R55938 DVSS.n4240 DVSS.n4239 2.6005
R55939 DVSS.n4242 DVSS.n4241 2.6005
R55940 DVSS.n4245 DVSS.n4244 2.6005
R55941 DVSS.n4247 DVSS.n4246 2.6005
R55942 DVSS.n4250 DVSS.n4249 2.6005
R55943 DVSS.n4252 DVSS.n4251 2.6005
R55944 DVSS.n4255 DVSS.n4254 2.6005
R55945 DVSS.n4257 DVSS.n4256 2.6005
R55946 DVSS.n4260 DVSS.n4259 2.6005
R55947 DVSS.n4262 DVSS.n4261 2.6005
R55948 DVSS.n4265 DVSS.n4264 2.6005
R55949 DVSS.n4267 DVSS.n4266 2.6005
R55950 DVSS.n4270 DVSS.n4269 2.6005
R55951 DVSS.n4272 DVSS.n4271 2.6005
R55952 DVSS.n4275 DVSS.n4274 2.6005
R55953 DVSS.n4277 DVSS.n4276 2.6005
R55954 DVSS.n4280 DVSS.n4279 2.6005
R55955 DVSS.n4282 DVSS.n4281 2.6005
R55956 DVSS.n4285 DVSS.n4284 2.6005
R55957 DVSS.n4287 DVSS.n4286 2.6005
R55958 DVSS.n4290 DVSS.n4289 2.6005
R55959 DVSS.n4292 DVSS.n4291 2.6005
R55960 DVSS.n4295 DVSS.n4294 2.6005
R55961 DVSS.n4297 DVSS.n4296 2.6005
R55962 DVSS.n4300 DVSS.n4299 2.6005
R55963 DVSS.n4302 DVSS.n4301 2.6005
R55964 DVSS.n4305 DVSS.n4304 2.6005
R55965 DVSS.n4307 DVSS.n4306 2.6005
R55966 DVSS.n4310 DVSS.n4309 2.6005
R55967 DVSS.n4313 DVSS.n4312 2.6005
R55968 DVSS.n5361 DVSS.n5354 2.6005
R55969 DVSS.n5352 DVSS.n5351 2.6005
R55970 DVSS.n5351 DVSS.n1375 2.6005
R55971 DVSS.n5350 DVSS.n1376 2.6005
R55972 DVSS.n5503 DVSS.n1376 2.6005
R55973 DVSS.n1647 DVSS.n1523 2.6005
R55974 DVSS.n1647 DVSS.n1374 2.6005
R55975 DVSS.n5196 DVSS.n1648 2.6005
R55976 DVSS.n1648 DVSS.n1645 2.6005
R55977 DVSS.n5198 DVSS.n5197 2.6005
R55978 DVSS.n5203 DVSS.n5198 2.6005
R55979 DVSS.n5195 DVSS.n1646 2.6005
R55980 DVSS.n1646 DVSS.n1639 2.6005
R55981 DVSS.n5194 DVSS.n1640 2.6005
R55982 DVSS.n5209 DVSS.n1640 2.6005
R55983 DVSS.n5193 DVSS.n5192 2.6005
R55984 DVSS.n5192 DVSS.n1634 2.6005
R55985 DVSS.n5191 DVSS.n1635 2.6005
R55986 DVSS.n5215 DVSS.n1635 2.6005
R55987 DVSS.n5190 DVSS.n5189 2.6005
R55988 DVSS.n5189 DVSS.n1629 2.6005
R55989 DVSS.n5188 DVSS.n1630 2.6005
R55990 DVSS.n5221 DVSS.n1630 2.6005
R55991 DVSS.n5187 DVSS.n5186 2.6005
R55992 DVSS.n5186 DVSS.n1624 2.6005
R55993 DVSS.n5185 DVSS.n1625 2.6005
R55994 DVSS.n5227 DVSS.n1625 2.6005
R55995 DVSS.n5184 DVSS.n5183 2.6005
R55996 DVSS.n5183 DVSS.n1619 2.6005
R55997 DVSS.n5182 DVSS.n1620 2.6005
R55998 DVSS.n5233 DVSS.n1620 2.6005
R55999 DVSS.n5181 DVSS.n5180 2.6005
R56000 DVSS.n5180 DVSS.n1614 2.6005
R56001 DVSS.n5179 DVSS.n1615 2.6005
R56002 DVSS.n5239 DVSS.n1615 2.6005
R56003 DVSS.n5178 DVSS.n5177 2.6005
R56004 DVSS.n5177 DVSS.n1609 2.6005
R56005 DVSS.n5176 DVSS.n1610 2.6005
R56006 DVSS.n5245 DVSS.n1610 2.6005
R56007 DVSS.n5175 DVSS.n5174 2.6005
R56008 DVSS.n5174 DVSS.n1604 2.6005
R56009 DVSS.n5173 DVSS.n1605 2.6005
R56010 DVSS.n5251 DVSS.n1605 2.6005
R56011 DVSS.n5172 DVSS.n5171 2.6005
R56012 DVSS.n5171 DVSS.n1597 2.6005
R56013 DVSS.n5170 DVSS.n1598 2.6005
R56014 DVSS.n5257 DVSS.n1598 2.6005
R56015 DVSS.n1929 DVSS.n1649 2.6005
R56016 DVSS.n1929 DVSS.n1596 2.6005
R56017 DVSS.n4781 DVSS.n1930 2.6005
R56018 DVSS.n1930 DVSS.n1927 2.6005
R56019 DVSS.n4783 DVSS.n4782 2.6005
R56020 DVSS.n4792 DVSS.n4783 2.6005
R56021 DVSS.n4780 DVSS.n1928 2.6005
R56022 DVSS.n1928 DVSS.n1922 2.6005
R56023 DVSS.n4779 DVSS.n1923 2.6005
R56024 DVSS.n4798 DVSS.n1923 2.6005
R56025 DVSS.n4778 DVSS.n4777 2.6005
R56026 DVSS.n4777 DVSS.n1917 2.6005
R56027 DVSS.n4776 DVSS.n1918 2.6005
R56028 DVSS.n4804 DVSS.n1918 2.6005
R56029 DVSS.n4775 DVSS.n4774 2.6005
R56030 DVSS.n4774 DVSS.n1912 2.6005
R56031 DVSS.n4773 DVSS.n1913 2.6005
R56032 DVSS.n4810 DVSS.n1913 2.6005
R56033 DVSS.n4772 DVSS.n4771 2.6005
R56034 DVSS.n4771 DVSS.n1907 2.6005
R56035 DVSS.n4770 DVSS.n1908 2.6005
R56036 DVSS.n4816 DVSS.n1908 2.6005
R56037 DVSS.n4769 DVSS.n4768 2.6005
R56038 DVSS.n4768 DVSS.n1902 2.6005
R56039 DVSS.n4767 DVSS.n1903 2.6005
R56040 DVSS.n4822 DVSS.n1903 2.6005
R56041 DVSS.n4766 DVSS.n4765 2.6005
R56042 DVSS.n4765 DVSS.n1897 2.6005
R56043 DVSS.n4764 DVSS.n1898 2.6005
R56044 DVSS.n4828 DVSS.n1898 2.6005
R56045 DVSS.n4763 DVSS.n4762 2.6005
R56046 DVSS.n4762 DVSS.n1892 2.6005
R56047 DVSS.n4761 DVSS.n1893 2.6005
R56048 DVSS.n4834 DVSS.n1893 2.6005
R56049 DVSS.n4760 DVSS.n4759 2.6005
R56050 DVSS.n4759 DVSS.n1886 2.6005
R56051 DVSS.n4758 DVSS.n1887 2.6005
R56052 DVSS.n4840 DVSS.n1887 2.6005
R56053 DVSS.n4757 DVSS.n4756 2.6005
R56054 DVSS.n4756 DVSS.n1879 2.6005
R56055 DVSS.n4755 DVSS.n1880 2.6005
R56056 DVSS.n4846 DVSS.n1880 2.6005
R56057 DVSS.n4754 DVSS.n4753 2.6005
R56058 DVSS.n4753 DVSS.n1878 2.6005
R56059 DVSS.n4752 DVSS.n1961 2.6005
R56060 DVSS.n4752 DVSS.n4751 2.6005
R56061 DVSS.n1960 DVSS.n1932 2.6005
R56062 DVSS.n1962 DVSS.n1932 2.6005
R56063 DVSS.n1959 DVSS.n1958 2.6005
R56064 DVSS.n1958 DVSS.n1858 2.6005
R56065 DVSS.n1957 DVSS.n1859 2.6005
R56066 DVSS.n4855 DVSS.n1859 2.6005
R56067 DVSS.n1956 DVSS.n1955 2.6005
R56068 DVSS.n1955 DVSS.n1853 2.6005
R56069 DVSS.n1954 DVSS.n1854 2.6005
R56070 DVSS.n4861 DVSS.n1854 2.6005
R56071 DVSS.n1953 DVSS.n1952 2.6005
R56072 DVSS.n1952 DVSS.n1848 2.6005
R56073 DVSS.n1951 DVSS.n1849 2.6005
R56074 DVSS.n4867 DVSS.n1849 2.6005
R56075 DVSS.n1950 DVSS.n1949 2.6005
R56076 DVSS.n1949 DVSS.n1843 2.6005
R56077 DVSS.n1948 DVSS.n1844 2.6005
R56078 DVSS.n4873 DVSS.n1844 2.6005
R56079 DVSS.n1947 DVSS.n1946 2.6005
R56080 DVSS.n1946 DVSS.n1838 2.6005
R56081 DVSS.n1945 DVSS.n1839 2.6005
R56082 DVSS.n4879 DVSS.n1839 2.6005
R56083 DVSS.n1944 DVSS.n1943 2.6005
R56084 DVSS.n1943 DVSS.n1833 2.6005
R56085 DVSS.n1942 DVSS.n1834 2.6005
R56086 DVSS.n4885 DVSS.n1834 2.6005
R56087 DVSS.n1941 DVSS.n1940 2.6005
R56088 DVSS.n1940 DVSS.n1828 2.6005
R56089 DVSS.n1939 DVSS.n1829 2.6005
R56090 DVSS.n4891 DVSS.n1829 2.6005
R56091 DVSS.n1938 DVSS.n1937 2.6005
R56092 DVSS.n1937 DVSS.n1823 2.6005
R56093 DVSS.n1936 DVSS.n1824 2.6005
R56094 DVSS.n4897 DVSS.n1824 2.6005
R56095 DVSS.n1935 DVSS.n1934 2.6005
R56096 DVSS.n1934 DVSS.n1816 2.6005
R56097 DVSS.n1933 DVSS.n1817 2.6005
R56098 DVSS.n4903 DVSS.n1817 2.6005
R56099 DVSS.n1807 DVSS.n1805 2.6005
R56100 DVSS.n1809 DVSS.n1807 2.6005
R56101 DVSS.n4911 DVSS.n4910 2.6005
R56102 DVSS.n4910 DVSS.n4909 2.6005
R56103 DVSS.n1806 DVSS.n1804 2.6005
R56104 DVSS.n1808 DVSS.n1806 2.6005
R56105 DVSS.n4359 DVSS.n4001 2.6005
R56106 DVSS.n4001 DVSS.n3999 2.6005
R56107 DVSS.n4361 DVSS.n4360 2.6005
R56108 DVSS.n4373 DVSS.n4361 2.6005
R56109 DVSS.n4358 DVSS.n4000 2.6005
R56110 DVSS.n4000 DVSS.n3993 2.6005
R56111 DVSS.n4357 DVSS.n3994 2.6005
R56112 DVSS.n4379 DVSS.n3994 2.6005
R56113 DVSS.n4356 DVSS.n4355 2.6005
R56114 DVSS.n4355 DVSS.n3988 2.6005
R56115 DVSS.n4354 DVSS.n3989 2.6005
R56116 DVSS.n4385 DVSS.n3989 2.6005
R56117 DVSS.n4353 DVSS.n4352 2.6005
R56118 DVSS.n4352 DVSS.n3983 2.6005
R56119 DVSS.n4351 DVSS.n3984 2.6005
R56120 DVSS.n4391 DVSS.n3984 2.6005
R56121 DVSS.n4350 DVSS.n4349 2.6005
R56122 DVSS.n4349 DVSS.n3978 2.6005
R56123 DVSS.n4348 DVSS.n3979 2.6005
R56124 DVSS.n4397 DVSS.n3979 2.6005
R56125 DVSS.n4347 DVSS.n4346 2.6005
R56126 DVSS.n4346 DVSS.n3973 2.6005
R56127 DVSS.n4345 DVSS.n3974 2.6005
R56128 DVSS.n4403 DVSS.n3974 2.6005
R56129 DVSS.n4344 DVSS.n4343 2.6005
R56130 DVSS.n4343 DVSS.n3968 2.6005
R56131 DVSS.n4342 DVSS.n3969 2.6005
R56132 DVSS.n4409 DVSS.n3969 2.6005
R56133 DVSS.n4341 DVSS.n4340 2.6005
R56134 DVSS.n4340 DVSS.n3963 2.6005
R56135 DVSS.n4339 DVSS.n3964 2.6005
R56136 DVSS.n4415 DVSS.n3964 2.6005
R56137 DVSS.n4338 DVSS.n4337 2.6005
R56138 DVSS.n4337 DVSS.n3958 2.6005
R56139 DVSS.n4336 DVSS.n3959 2.6005
R56140 DVSS.n4421 DVSS.n3959 2.6005
R56141 DVSS.n4335 DVSS.n4334 2.6005
R56142 DVSS.n4334 DVSS.n3891 2.6005
R56143 DVSS.n4333 DVSS.n3892 2.6005
R56144 DVSS.n4427 DVSS.n3892 2.6005
R56145 DVSS.n4331 DVSS.n4330 2.6005
R56146 DVSS.n4330 DVSS.n3890 2.6005
R56147 DVSS.n1516 DVSS.n1515 2.6005
R56148 DVSS.n1513 DVSS.n1512 2.6005
R56149 DVSS.n1511 DVSS.n1510 2.6005
R56150 DVSS.n1508 DVSS.n1507 2.6005
R56151 DVSS.n1506 DVSS.n1505 2.6005
R56152 DVSS.n1503 DVSS.n1502 2.6005
R56153 DVSS.n1501 DVSS.n1500 2.6005
R56154 DVSS.n1498 DVSS.n1497 2.6005
R56155 DVSS.n1496 DVSS.n1495 2.6005
R56156 DVSS.n1493 DVSS.n1492 2.6005
R56157 DVSS.n1491 DVSS.n1490 2.6005
R56158 DVSS.n1488 DVSS.n1487 2.6005
R56159 DVSS.n1486 DVSS.n1485 2.6005
R56160 DVSS.n1483 DVSS.n1482 2.6005
R56161 DVSS.n1481 DVSS.n1480 2.6005
R56162 DVSS.n1478 DVSS.n1477 2.6005
R56163 DVSS.n1476 DVSS.n1475 2.6005
R56164 DVSS.n1473 DVSS.n1472 2.6005
R56165 DVSS.n1471 DVSS.n1470 2.6005
R56166 DVSS.n1468 DVSS.n1467 2.6005
R56167 DVSS.n1466 DVSS.n1465 2.6005
R56168 DVSS.n1463 DVSS.n1462 2.6005
R56169 DVSS.n1461 DVSS.n1460 2.6005
R56170 DVSS.n1458 DVSS.n1457 2.6005
R56171 DVSS.n1456 DVSS.n1455 2.6005
R56172 DVSS.n1453 DVSS.n1452 2.6005
R56173 DVSS.n1451 DVSS.n1450 2.6005
R56174 DVSS.n1448 DVSS.n1447 2.6005
R56175 DVSS.n1446 DVSS.n1445 2.6005
R56176 DVSS.n1443 DVSS.n1442 2.6005
R56177 DVSS.n1441 DVSS.n1440 2.6005
R56178 DVSS.n1438 DVSS.n1437 2.6005
R56179 DVSS.n1436 DVSS.n1435 2.6005
R56180 DVSS.n1433 DVSS.n1432 2.6005
R56181 DVSS.n1431 DVSS.n1430 2.6005
R56182 DVSS.n1428 DVSS.n1427 2.6005
R56183 DVSS.n1426 DVSS.n1425 2.6005
R56184 DVSS.n1423 DVSS.n1422 2.6005
R56185 DVSS.n1421 DVSS.n1420 2.6005
R56186 DVSS.n1418 DVSS.n1417 2.6005
R56187 DVSS.n1416 DVSS.n1415 2.6005
R56188 DVSS.n1413 DVSS.n1380 2.6005
R56189 DVSS.n5502 DVSS.n5501 2.6005
R56190 DVSS.n5503 DVSS.n5502 2.6005
R56191 DVSS.n1642 DVSS.n1377 2.6005
R56192 DVSS.n1377 DVSS.n1374 2.6005
R56193 DVSS.n1644 DVSS.n1643 2.6005
R56194 DVSS.n1645 DVSS.n1644 2.6005
R56195 DVSS.n5205 DVSS.n5204 2.6005
R56196 DVSS.n5204 DVSS.n5203 2.6005
R56197 DVSS.n5206 DVSS.n1641 2.6005
R56198 DVSS.n1641 DVSS.n1639 2.6005
R56199 DVSS.n5208 DVSS.n5207 2.6005
R56200 DVSS.n5209 DVSS.n5208 2.6005
R56201 DVSS.n1633 DVSS.n1632 2.6005
R56202 DVSS.n1634 DVSS.n1633 2.6005
R56203 DVSS.n5217 DVSS.n5216 2.6005
R56204 DVSS.n5216 DVSS.n5215 2.6005
R56205 DVSS.n5218 DVSS.n1631 2.6005
R56206 DVSS.n1631 DVSS.n1629 2.6005
R56207 DVSS.n5220 DVSS.n5219 2.6005
R56208 DVSS.n5221 DVSS.n5220 2.6005
R56209 DVSS.n1623 DVSS.n1622 2.6005
R56210 DVSS.n1624 DVSS.n1623 2.6005
R56211 DVSS.n5229 DVSS.n5228 2.6005
R56212 DVSS.n5228 DVSS.n5227 2.6005
R56213 DVSS.n5230 DVSS.n1621 2.6005
R56214 DVSS.n1621 DVSS.n1619 2.6005
R56215 DVSS.n5232 DVSS.n5231 2.6005
R56216 DVSS.n5233 DVSS.n5232 2.6005
R56217 DVSS.n1613 DVSS.n1612 2.6005
R56218 DVSS.n1614 DVSS.n1613 2.6005
R56219 DVSS.n5241 DVSS.n5240 2.6005
R56220 DVSS.n5240 DVSS.n5239 2.6005
R56221 DVSS.n5242 DVSS.n1611 2.6005
R56222 DVSS.n1611 DVSS.n1609 2.6005
R56223 DVSS.n5244 DVSS.n5243 2.6005
R56224 DVSS.n5245 DVSS.n5244 2.6005
R56225 DVSS.n1603 DVSS.n1602 2.6005
R56226 DVSS.n1604 DVSS.n1603 2.6005
R56227 DVSS.n5253 DVSS.n5252 2.6005
R56228 DVSS.n5252 DVSS.n5251 2.6005
R56229 DVSS.n5254 DVSS.n1600 2.6005
R56230 DVSS.n1600 DVSS.n1597 2.6005
R56231 DVSS.n5256 DVSS.n5255 2.6005
R56232 DVSS.n5257 DVSS.n5256 2.6005
R56233 DVSS.n4787 DVSS.n1599 2.6005
R56234 DVSS.n1599 DVSS.n1596 2.6005
R56235 DVSS.n4789 DVSS.n4784 2.6005
R56236 DVSS.n4784 DVSS.n1927 2.6005
R56237 DVSS.n4791 DVSS.n4790 2.6005
R56238 DVSS.n4792 DVSS.n4791 2.6005
R56239 DVSS.n1921 DVSS.n1920 2.6005
R56240 DVSS.n1922 DVSS.n1921 2.6005
R56241 DVSS.n4800 DVSS.n4799 2.6005
R56242 DVSS.n4799 DVSS.n4798 2.6005
R56243 DVSS.n4801 DVSS.n1919 2.6005
R56244 DVSS.n1919 DVSS.n1917 2.6005
R56245 DVSS.n4803 DVSS.n4802 2.6005
R56246 DVSS.n4804 DVSS.n4803 2.6005
R56247 DVSS.n1911 DVSS.n1910 2.6005
R56248 DVSS.n1912 DVSS.n1911 2.6005
R56249 DVSS.n4812 DVSS.n4811 2.6005
R56250 DVSS.n4811 DVSS.n4810 2.6005
R56251 DVSS.n4813 DVSS.n1909 2.6005
R56252 DVSS.n1909 DVSS.n1907 2.6005
R56253 DVSS.n4815 DVSS.n4814 2.6005
R56254 DVSS.n4816 DVSS.n4815 2.6005
R56255 DVSS.n1901 DVSS.n1900 2.6005
R56256 DVSS.n1902 DVSS.n1901 2.6005
R56257 DVSS.n4824 DVSS.n4823 2.6005
R56258 DVSS.n4823 DVSS.n4822 2.6005
R56259 DVSS.n4825 DVSS.n1899 2.6005
R56260 DVSS.n1899 DVSS.n1897 2.6005
R56261 DVSS.n4827 DVSS.n4826 2.6005
R56262 DVSS.n4828 DVSS.n4827 2.6005
R56263 DVSS.n1891 DVSS.n1890 2.6005
R56264 DVSS.n1892 DVSS.n1891 2.6005
R56265 DVSS.n4836 DVSS.n4835 2.6005
R56266 DVSS.n4835 DVSS.n4834 2.6005
R56267 DVSS.n4837 DVSS.n1888 2.6005
R56268 DVSS.n1888 DVSS.n1886 2.6005
R56269 DVSS.n4839 DVSS.n4838 2.6005
R56270 DVSS.n4840 DVSS.n4839 2.6005
R56271 DVSS.n1889 DVSS.n1877 2.6005
R56272 DVSS.n1879 DVSS.n1877 2.6005
R56273 DVSS.n4848 DVSS.n4847 2.6005
R56274 DVSS.n4847 DVSS.n4846 2.6005
R56275 DVSS.n1876 DVSS.n1874 2.6005
R56276 DVSS.n1878 DVSS.n1876 2.6005
R56277 DVSS.n1968 DVSS.n1967 2.6005
R56278 DVSS.n4751 DVSS.n1968 2.6005
R56279 DVSS.n1963 DVSS.n1864 2.6005
R56280 DVSS.n1963 DVSS.n1962 2.6005
R56281 DVSS.n4852 DVSS.n1860 2.6005
R56282 DVSS.n1860 DVSS.n1858 2.6005
R56283 DVSS.n4854 DVSS.n4853 2.6005
R56284 DVSS.n4855 DVSS.n4854 2.6005
R56285 DVSS.n1852 DVSS.n1851 2.6005
R56286 DVSS.n1853 DVSS.n1852 2.6005
R56287 DVSS.n4863 DVSS.n4862 2.6005
R56288 DVSS.n4862 DVSS.n4861 2.6005
R56289 DVSS.n4864 DVSS.n1850 2.6005
R56290 DVSS.n1850 DVSS.n1848 2.6005
R56291 DVSS.n4866 DVSS.n4865 2.6005
R56292 DVSS.n4867 DVSS.n4866 2.6005
R56293 DVSS.n1842 DVSS.n1841 2.6005
R56294 DVSS.n1843 DVSS.n1842 2.6005
R56295 DVSS.n4875 DVSS.n4874 2.6005
R56296 DVSS.n4874 DVSS.n4873 2.6005
R56297 DVSS.n4876 DVSS.n1840 2.6005
R56298 DVSS.n1840 DVSS.n1838 2.6005
R56299 DVSS.n4878 DVSS.n4877 2.6005
R56300 DVSS.n4879 DVSS.n4878 2.6005
R56301 DVSS.n1832 DVSS.n1831 2.6005
R56302 DVSS.n1833 DVSS.n1832 2.6005
R56303 DVSS.n4887 DVSS.n4886 2.6005
R56304 DVSS.n4886 DVSS.n4885 2.6005
R56305 DVSS.n4888 DVSS.n1830 2.6005
R56306 DVSS.n1830 DVSS.n1828 2.6005
R56307 DVSS.n4890 DVSS.n4889 2.6005
R56308 DVSS.n4891 DVSS.n4890 2.6005
R56309 DVSS.n1822 DVSS.n1821 2.6005
R56310 DVSS.n1823 DVSS.n1822 2.6005
R56311 DVSS.n4899 DVSS.n4898 2.6005
R56312 DVSS.n4898 DVSS.n4897 2.6005
R56313 DVSS.n4900 DVSS.n1819 2.6005
R56314 DVSS.n1819 DVSS.n1816 2.6005
R56315 DVSS.n4902 DVSS.n4901 2.6005
R56316 DVSS.n4903 DVSS.n4902 2.6005
R56317 DVSS.n1820 DVSS.n1818 2.6005
R56318 DVSS.n1818 DVSS.n1809 2.6005
R56319 DVSS.n4366 DVSS.n1810 2.6005
R56320 DVSS.n4909 DVSS.n1810 2.6005
R56321 DVSS.n4369 DVSS.n4368 2.6005
R56322 DVSS.n4368 DVSS.n1808 2.6005
R56323 DVSS.n4370 DVSS.n4362 2.6005
R56324 DVSS.n4362 DVSS.n3999 2.6005
R56325 DVSS.n4372 DVSS.n4371 2.6005
R56326 DVSS.n4373 DVSS.n4372 2.6005
R56327 DVSS.n3992 DVSS.n3991 2.6005
R56328 DVSS.n3993 DVSS.n3992 2.6005
R56329 DVSS.n4381 DVSS.n4380 2.6005
R56330 DVSS.n4380 DVSS.n4379 2.6005
R56331 DVSS.n4382 DVSS.n3990 2.6005
R56332 DVSS.n3990 DVSS.n3988 2.6005
R56333 DVSS.n4384 DVSS.n4383 2.6005
R56334 DVSS.n4385 DVSS.n4384 2.6005
R56335 DVSS.n3982 DVSS.n3981 2.6005
R56336 DVSS.n3983 DVSS.n3982 2.6005
R56337 DVSS.n4393 DVSS.n4392 2.6005
R56338 DVSS.n4392 DVSS.n4391 2.6005
R56339 DVSS.n4394 DVSS.n3980 2.6005
R56340 DVSS.n3980 DVSS.n3978 2.6005
R56341 DVSS.n4396 DVSS.n4395 2.6005
R56342 DVSS.n4397 DVSS.n4396 2.6005
R56343 DVSS.n3972 DVSS.n3971 2.6005
R56344 DVSS.n3973 DVSS.n3972 2.6005
R56345 DVSS.n4405 DVSS.n4404 2.6005
R56346 DVSS.n4404 DVSS.n4403 2.6005
R56347 DVSS.n4406 DVSS.n3970 2.6005
R56348 DVSS.n3970 DVSS.n3968 2.6005
R56349 DVSS.n4408 DVSS.n4407 2.6005
R56350 DVSS.n4409 DVSS.n4408 2.6005
R56351 DVSS.n3962 DVSS.n3961 2.6005
R56352 DVSS.n3963 DVSS.n3962 2.6005
R56353 DVSS.n4417 DVSS.n4416 2.6005
R56354 DVSS.n4416 DVSS.n4415 2.6005
R56355 DVSS.n4418 DVSS.n3960 2.6005
R56356 DVSS.n3960 DVSS.n3958 2.6005
R56357 DVSS.n4420 DVSS.n4419 2.6005
R56358 DVSS.n4421 DVSS.n4420 2.6005
R56359 DVSS.n3889 DVSS.n3887 2.6005
R56360 DVSS.n3891 DVSS.n3889 2.6005
R56361 DVSS.n4429 DVSS.n4428 2.6005
R56362 DVSS.n4428 DVSS.n4427 2.6005
R56363 DVSS.n3888 DVSS.n3886 2.6005
R56364 DVSS.n3890 DVSS.n3888 2.6005
R56365 DVSS.n5496 DVSS.n1381 2.6005
R56366 DVSS.n5494 DVSS.n5493 2.6005
R56367 DVSS.n5492 DVSS.n5491 2.6005
R56368 DVSS.n5489 DVSS.n5363 2.6005
R56369 DVSS.n5487 DVSS.n5486 2.6005
R56370 DVSS.n5485 DVSS.n5484 2.6005
R56371 DVSS.n5482 DVSS.n5365 2.6005
R56372 DVSS.n5480 DVSS.n5479 2.6005
R56373 DVSS.n5478 DVSS.n5477 2.6005
R56374 DVSS.n5475 DVSS.n5367 2.6005
R56375 DVSS.n5473 DVSS.n5472 2.6005
R56376 DVSS.n5471 DVSS.n5470 2.6005
R56377 DVSS.n5468 DVSS.n5369 2.6005
R56378 DVSS.n5466 DVSS.n5465 2.6005
R56379 DVSS.n5464 DVSS.n5463 2.6005
R56380 DVSS.n5461 DVSS.n5371 2.6005
R56381 DVSS.n5459 DVSS.n5458 2.6005
R56382 DVSS.n5457 DVSS.n5456 2.6005
R56383 DVSS.n5454 DVSS.n5373 2.6005
R56384 DVSS.n5452 DVSS.n5451 2.6005
R56385 DVSS.n5450 DVSS.n5449 2.6005
R56386 DVSS.n5447 DVSS.n5446 2.6005
R56387 DVSS.n5445 DVSS.n5444 2.6005
R56388 DVSS.n5442 DVSS.n5441 2.6005
R56389 DVSS.n5440 DVSS.n5439 2.6005
R56390 DVSS.n5437 DVSS.n5378 2.6005
R56391 DVSS.n5435 DVSS.n5434 2.6005
R56392 DVSS.n5433 DVSS.n5432 2.6005
R56393 DVSS.n5430 DVSS.n5380 2.6005
R56394 DVSS.n5428 DVSS.n5427 2.6005
R56395 DVSS.n5426 DVSS.n5425 2.6005
R56396 DVSS.n5423 DVSS.n5382 2.6005
R56397 DVSS.n5421 DVSS.n5420 2.6005
R56398 DVSS.n5419 DVSS.n5418 2.6005
R56399 DVSS.n5416 DVSS.n5384 2.6005
R56400 DVSS.n5414 DVSS.n5413 2.6005
R56401 DVSS.n5412 DVSS.n5411 2.6005
R56402 DVSS.n5409 DVSS.n5386 2.6005
R56403 DVSS.n5407 DVSS.n5406 2.6005
R56404 DVSS.n5405 DVSS.n5404 2.6005
R56405 DVSS.n5402 DVSS.n5388 2.6005
R56406 DVSS.n5400 DVSS.n5399 2.6005
R56407 DVSS.n5398 DVSS.n5397 2.6005
R56408 DVSS.n5391 DVSS.n5361 2.6005
R56409 DVSS.n1373 DVSS.n1371 2.6005
R56410 DVSS.n1375 DVSS.n1373 2.6005
R56411 DVSS.n5505 DVSS.n5504 2.6005
R56412 DVSS.n5504 DVSS.n5503 2.6005
R56413 DVSS.n1372 DVSS.n1370 2.6005
R56414 DVSS.n1374 DVSS.n1372 2.6005
R56415 DVSS.n5200 DVSS.n5199 2.6005
R56416 DVSS.n5199 DVSS.n1645 2.6005
R56417 DVSS.n5202 DVSS.n5201 2.6005
R56418 DVSS.n5203 DVSS.n5202 2.6005
R56419 DVSS.n1638 DVSS.n1637 2.6005
R56420 DVSS.n1639 DVSS.n1638 2.6005
R56421 DVSS.n5211 DVSS.n5210 2.6005
R56422 DVSS.n5210 DVSS.n5209 2.6005
R56423 DVSS.n5212 DVSS.n1636 2.6005
R56424 DVSS.n1636 DVSS.n1634 2.6005
R56425 DVSS.n5214 DVSS.n5213 2.6005
R56426 DVSS.n5215 DVSS.n5214 2.6005
R56427 DVSS.n1628 DVSS.n1627 2.6005
R56428 DVSS.n1629 DVSS.n1628 2.6005
R56429 DVSS.n5223 DVSS.n5222 2.6005
R56430 DVSS.n5222 DVSS.n5221 2.6005
R56431 DVSS.n5224 DVSS.n1626 2.6005
R56432 DVSS.n1626 DVSS.n1624 2.6005
R56433 DVSS.n5226 DVSS.n5225 2.6005
R56434 DVSS.n5227 DVSS.n5226 2.6005
R56435 DVSS.n1618 DVSS.n1617 2.6005
R56436 DVSS.n1619 DVSS.n1618 2.6005
R56437 DVSS.n5235 DVSS.n5234 2.6005
R56438 DVSS.n5234 DVSS.n5233 2.6005
R56439 DVSS.n5236 DVSS.n1616 2.6005
R56440 DVSS.n1616 DVSS.n1614 2.6005
R56441 DVSS.n5238 DVSS.n5237 2.6005
R56442 DVSS.n5239 DVSS.n5238 2.6005
R56443 DVSS.n1608 DVSS.n1607 2.6005
R56444 DVSS.n1609 DVSS.n1608 2.6005
R56445 DVSS.n5247 DVSS.n5246 2.6005
R56446 DVSS.n5246 DVSS.n5245 2.6005
R56447 DVSS.n5248 DVSS.n1606 2.6005
R56448 DVSS.n1606 DVSS.n1604 2.6005
R56449 DVSS.n5250 DVSS.n5249 2.6005
R56450 DVSS.n5251 DVSS.n5250 2.6005
R56451 DVSS.n1595 DVSS.n1593 2.6005
R56452 DVSS.n1597 DVSS.n1595 2.6005
R56453 DVSS.n5259 DVSS.n5258 2.6005
R56454 DVSS.n5258 DVSS.n5257 2.6005
R56455 DVSS.n1594 DVSS.n1592 2.6005
R56456 DVSS.n1596 DVSS.n1594 2.6005
R56457 DVSS.n1926 DVSS.n1925 2.6005
R56458 DVSS.n1927 DVSS.n1926 2.6005
R56459 DVSS.n4794 DVSS.n4793 2.6005
R56460 DVSS.n4793 DVSS.n4792 2.6005
R56461 DVSS.n4795 DVSS.n1924 2.6005
R56462 DVSS.n1924 DVSS.n1922 2.6005
R56463 DVSS.n4797 DVSS.n4796 2.6005
R56464 DVSS.n4798 DVSS.n4797 2.6005
R56465 DVSS.n1916 DVSS.n1915 2.6005
R56466 DVSS.n1917 DVSS.n1916 2.6005
R56467 DVSS.n4806 DVSS.n4805 2.6005
R56468 DVSS.n4805 DVSS.n4804 2.6005
R56469 DVSS.n4807 DVSS.n1914 2.6005
R56470 DVSS.n1914 DVSS.n1912 2.6005
R56471 DVSS.n4809 DVSS.n4808 2.6005
R56472 DVSS.n4810 DVSS.n4809 2.6005
R56473 DVSS.n1906 DVSS.n1905 2.6005
R56474 DVSS.n1907 DVSS.n1906 2.6005
R56475 DVSS.n4818 DVSS.n4817 2.6005
R56476 DVSS.n4817 DVSS.n4816 2.6005
R56477 DVSS.n4819 DVSS.n1904 2.6005
R56478 DVSS.n1904 DVSS.n1902 2.6005
R56479 DVSS.n4821 DVSS.n4820 2.6005
R56480 DVSS.n4822 DVSS.n4821 2.6005
R56481 DVSS.n1896 DVSS.n1895 2.6005
R56482 DVSS.n1897 DVSS.n1896 2.6005
R56483 DVSS.n4830 DVSS.n4829 2.6005
R56484 DVSS.n4829 DVSS.n4828 2.6005
R56485 DVSS.n4831 DVSS.n1894 2.6005
R56486 DVSS.n1894 DVSS.n1892 2.6005
R56487 DVSS.n4833 DVSS.n4832 2.6005
R56488 DVSS.n4834 DVSS.n4833 2.6005
R56489 DVSS.n1885 DVSS.n1884 2.6005
R56490 DVSS.n1886 DVSS.n1885 2.6005
R56491 DVSS.n4842 DVSS.n4841 2.6005
R56492 DVSS.n4841 DVSS.n4840 2.6005
R56493 DVSS.n4843 DVSS.n1882 2.6005
R56494 DVSS.n1882 DVSS.n1879 2.6005
R56495 DVSS.n4845 DVSS.n4844 2.6005
R56496 DVSS.n4846 DVSS.n4845 2.6005
R56497 DVSS.n1883 DVSS.n1881 2.6005
R56498 DVSS.n1881 DVSS.n1878 2.6005
R56499 DVSS.n4750 DVSS.n4749 2.6005
R56500 DVSS.n4751 DVSS.n4750 2.6005
R56501 DVSS.n1970 DVSS.n1969 2.6005
R56502 DVSS.n1969 DVSS.n1962 2.6005
R56503 DVSS.n1857 DVSS.n1856 2.6005
R56504 DVSS.n1858 DVSS.n1857 2.6005
R56505 DVSS.n4857 DVSS.n4856 2.6005
R56506 DVSS.n4856 DVSS.n4855 2.6005
R56507 DVSS.n4858 DVSS.n1855 2.6005
R56508 DVSS.n1855 DVSS.n1853 2.6005
R56509 DVSS.n4860 DVSS.n4859 2.6005
R56510 DVSS.n4861 DVSS.n4860 2.6005
R56511 DVSS.n1847 DVSS.n1846 2.6005
R56512 DVSS.n1848 DVSS.n1847 2.6005
R56513 DVSS.n4869 DVSS.n4868 2.6005
R56514 DVSS.n4868 DVSS.n4867 2.6005
R56515 DVSS.n4870 DVSS.n1845 2.6005
R56516 DVSS.n1845 DVSS.n1843 2.6005
R56517 DVSS.n4872 DVSS.n4871 2.6005
R56518 DVSS.n4873 DVSS.n4872 2.6005
R56519 DVSS.n1837 DVSS.n1836 2.6005
R56520 DVSS.n1838 DVSS.n1837 2.6005
R56521 DVSS.n4881 DVSS.n4880 2.6005
R56522 DVSS.n4880 DVSS.n4879 2.6005
R56523 DVSS.n4882 DVSS.n1835 2.6005
R56524 DVSS.n1835 DVSS.n1833 2.6005
R56525 DVSS.n4884 DVSS.n4883 2.6005
R56526 DVSS.n4885 DVSS.n4884 2.6005
R56527 DVSS.n1827 DVSS.n1826 2.6005
R56528 DVSS.n1828 DVSS.n1827 2.6005
R56529 DVSS.n4893 DVSS.n4892 2.6005
R56530 DVSS.n4892 DVSS.n4891 2.6005
R56531 DVSS.n4894 DVSS.n1825 2.6005
R56532 DVSS.n1825 DVSS.n1823 2.6005
R56533 DVSS.n4896 DVSS.n4895 2.6005
R56534 DVSS.n4897 DVSS.n4896 2.6005
R56535 DVSS.n1815 DVSS.n1814 2.6005
R56536 DVSS.n1816 DVSS.n1815 2.6005
R56537 DVSS.n4905 DVSS.n4904 2.6005
R56538 DVSS.n4904 DVSS.n4903 2.6005
R56539 DVSS.n4906 DVSS.n1812 2.6005
R56540 DVSS.n1812 DVSS.n1809 2.6005
R56541 DVSS.n4908 DVSS.n4907 2.6005
R56542 DVSS.n4909 DVSS.n4908 2.6005
R56543 DVSS.n3996 DVSS.n1811 2.6005
R56544 DVSS.n1811 DVSS.n1808 2.6005
R56545 DVSS.n3998 DVSS.n3997 2.6005
R56546 DVSS.n3999 DVSS.n3998 2.6005
R56547 DVSS.n4375 DVSS.n4374 2.6005
R56548 DVSS.n4374 DVSS.n4373 2.6005
R56549 DVSS.n4376 DVSS.n3995 2.6005
R56550 DVSS.n3995 DVSS.n3993 2.6005
R56551 DVSS.n4378 DVSS.n4377 2.6005
R56552 DVSS.n4379 DVSS.n4378 2.6005
R56553 DVSS.n3987 DVSS.n3986 2.6005
R56554 DVSS.n3988 DVSS.n3987 2.6005
R56555 DVSS.n4387 DVSS.n4386 2.6005
R56556 DVSS.n4386 DVSS.n4385 2.6005
R56557 DVSS.n4388 DVSS.n3985 2.6005
R56558 DVSS.n3985 DVSS.n3983 2.6005
R56559 DVSS.n4390 DVSS.n4389 2.6005
R56560 DVSS.n4391 DVSS.n4390 2.6005
R56561 DVSS.n3977 DVSS.n3976 2.6005
R56562 DVSS.n3978 DVSS.n3977 2.6005
R56563 DVSS.n4399 DVSS.n4398 2.6005
R56564 DVSS.n4398 DVSS.n4397 2.6005
R56565 DVSS.n4400 DVSS.n3975 2.6005
R56566 DVSS.n3975 DVSS.n3973 2.6005
R56567 DVSS.n4402 DVSS.n4401 2.6005
R56568 DVSS.n4403 DVSS.n4402 2.6005
R56569 DVSS.n3967 DVSS.n3966 2.6005
R56570 DVSS.n3968 DVSS.n3967 2.6005
R56571 DVSS.n4411 DVSS.n4410 2.6005
R56572 DVSS.n4410 DVSS.n4409 2.6005
R56573 DVSS.n4412 DVSS.n3965 2.6005
R56574 DVSS.n3965 DVSS.n3963 2.6005
R56575 DVSS.n4414 DVSS.n4413 2.6005
R56576 DVSS.n4415 DVSS.n4414 2.6005
R56577 DVSS.n3957 DVSS.n3956 2.6005
R56578 DVSS.n3958 DVSS.n3957 2.6005
R56579 DVSS.n4423 DVSS.n4422 2.6005
R56580 DVSS.n4422 DVSS.n4421 2.6005
R56581 DVSS.n4424 DVSS.n3894 2.6005
R56582 DVSS.n3894 DVSS.n3891 2.6005
R56583 DVSS.n4426 DVSS.n4425 2.6005
R56584 DVSS.n4427 DVSS.n4426 2.6005
R56585 DVSS.n4066 DVSS.n3893 2.6005
R56586 DVSS.n3893 DVSS.n3890 2.6005
R56587 DVSS.n4185 DVSS.n4184 2.5974
R56588 DVSS.n5355 DVSS.n1385 2.5974
R56589 DVSS.n5393 DVSS.n5392 2.36815
R56590 DVSS.n1522 DVSS.n1521 2.36815
R56591 DVSS.n6422 DVSS.n6421 2.25175
R56592 DVSS.n6470 DVSS.n110 2.25175
R56593 DVSS.n6439 DVSS.n6438 2.25175
R56594 DVSS.n6400 DVSS.n6399 2.25175
R56595 DVSS.n6422 DVSS.n223 2.251
R56596 DVSS.n6472 DVSS.n110 2.251
R56597 DVSS.n6438 DVSS.n207 2.251
R56598 DVSS.n6399 DVSS.n6397 2.251
R56599 DVSS.n5593 DVSS.n5592 2.2505
R56600 DVSS.n5658 DVSS.n5657 2.2505
R56601 DVSS.n4506 DVSS.n1873 2.25007
R56602 DVSS.n6454 DVSS.n171 2.25007
R56603 DVSS.n296 DVSS.n295 2.25007
R56604 DVSS.n464 DVSS.n457 2.25007
R56605 DVSS.n4743 DVSS.n1973 2.24901
R56606 DVSS.n3809 DVSS.n3808 2.24901
R56607 DVSS.n5794 DVSS.n5792 2.24901
R56608 DVSS.n4989 DVSS.n1741 2.24901
R56609 DVSS.n2753 DVSS.n2124 2.24901
R56610 DVSS.n2530 DVSS.n2397 2.24882
R56611 DVSS.n1250 DVSS.n1248 2.24648
R56612 DVSS.n502 DVSS.n490 2.24648
R56613 DVSS.n1259 DVSS.n1256 2.24648
R56614 DVSS.n1255 DVSS.n1252 2.24648
R56615 DVSS.n1778 DVSS.n1775 2.24581
R56616 DVSS.n2416 DVSS.n2411 2.24581
R56617 DVSS.n2408 DVSS.n2406 2.24581
R56618 DVSS.n2415 DVSS.n2414 2.24581
R56619 DVSS.n1792 DVSS.n1776 2.24581
R56620 DVSS.n5798 DVSS.n5795 2.24581
R56621 DVSS.n5798 DVSS.n5796 2.24581
R56622 DVSS.n5789 DVSS.n5775 2.24581
R56623 DVSS.n5798 DVSS.n5797 2.24581
R56624 DVSS.n5791 DVSS.n5775 2.24581
R56625 DVSS.n5798 DVSS.n5774 2.24581
R56626 DVSS.n1988 DVSS.n1984 2.24581
R56627 DVSS.n1994 DVSS.n1993 2.24581
R56628 DVSS.n1988 DVSS.n1985 2.24581
R56629 DVSS.n1994 DVSS.n1992 2.24581
R56630 DVSS.n1988 DVSS.n1986 2.24581
R56631 DVSS.n1994 DVSS.n1991 2.24581
R56632 DVSS.n1988 DVSS.n1987 2.24581
R56633 DVSS.n1994 DVSS.n1990 2.24581
R56634 DVSS.n1989 DVSS.n1988 2.24581
R56635 DVSS.n1994 DVSS.n1972 2.24581
R56636 DVSS.n4549 DVSS.n4548 2.24581
R56637 DVSS.n4517 DVSS.n4501 2.24581
R56638 DVSS.n4549 DVSS.n4547 2.24581
R56639 DVSS.n4519 DVSS.n4501 2.24581
R56640 DVSS.n4549 DVSS.n4546 2.24581
R56641 DVSS.n4521 DVSS.n4501 2.24581
R56642 DVSS.n4549 DVSS.n4545 2.24581
R56643 DVSS.n4523 DVSS.n4501 2.24581
R56644 DVSS.n4549 DVSS.n4544 2.24581
R56645 DVSS.n4525 DVSS.n4501 2.24581
R56646 DVSS.n4549 DVSS.n4543 2.24581
R56647 DVSS.n4527 DVSS.n4501 2.24581
R56648 DVSS.n4549 DVSS.n4542 2.24581
R56649 DVSS.n4529 DVSS.n4501 2.24581
R56650 DVSS.n4549 DVSS.n4541 2.24581
R56651 DVSS.n4531 DVSS.n4501 2.24581
R56652 DVSS.n4549 DVSS.n4540 2.24581
R56653 DVSS.n4533 DVSS.n4501 2.24581
R56654 DVSS.n4549 DVSS.n4539 2.24581
R56655 DVSS.n4535 DVSS.n4501 2.24581
R56656 DVSS.n4549 DVSS.n4538 2.24581
R56657 DVSS.n4537 DVSS.n4501 2.24581
R56658 DVSS.n3789 DVSS.n3730 2.24581
R56659 DVSS.n3793 DVSS.n3726 2.24581
R56660 DVSS.n3792 DVSS.n3730 2.24581
R56661 DVSS.n3796 DVSS.n3726 2.24581
R56662 DVSS.n3795 DVSS.n3730 2.24581
R56663 DVSS.n3799 DVSS.n3726 2.24581
R56664 DVSS.n3798 DVSS.n3730 2.24581
R56665 DVSS.n3802 DVSS.n3726 2.24581
R56666 DVSS.n3801 DVSS.n3730 2.24581
R56667 DVSS.n3805 DVSS.n3726 2.24581
R56668 DVSS.n4996 DVSS.n1744 2.24581
R56669 DVSS.n4996 DVSS.n1746 2.24581
R56670 DVSS.n1752 DVSS.n1751 2.24581
R56671 DVSS.n4996 DVSS.n1747 2.24581
R56672 DVSS.n4988 DVSS.n1752 2.24581
R56673 DVSS.n2763 DVSS.n2762 2.24581
R56674 DVSS.n2750 DVSS.n2745 2.24581
R56675 DVSS.n2763 DVSS.n2760 2.24581
R56676 DVSS.n2754 DVSS.n2745 2.24581
R56677 DVSS.n2763 DVSS.n2759 2.24581
R56678 DVSS.n2756 DVSS.n2745 2.24581
R56679 DVSS.n2546 DVSS.n2545 2.24581
R56680 DVSS.n2535 DVSS.n2525 2.24581
R56681 DVSS.n2546 DVSS.n2544 2.24581
R56682 DVSS.n2537 DVSS.n2525 2.24581
R56683 DVSS.n2546 DVSS.n2543 2.24581
R56684 DVSS.n2539 DVSS.n2525 2.24581
R56685 DVSS.n2546 DVSS.n2542 2.24581
R56686 DVSS.n2541 DVSS.n2525 2.24581
R56687 DVSS.n2758 DVSS.n2745 2.24581
R56688 DVSS.n1752 DVSS.n1738 2.24581
R56689 DVSS.n5793 DVSS.n5775 2.24581
R56690 DVSS.n1870 DVSS.n1868 2.24581
R56691 DVSS.n1872 DVSS.n1871 2.24581
R56692 DVSS.n1870 DVSS.n1869 2.24581
R56693 DVSS.n4849 DVSS.n1875 2.24581
R56694 DVSS.n6456 DVSS.n6455 2.24581
R56695 DVSS.n168 DVSS.n153 2.24581
R56696 DVSS.n6456 DVSS.n6453 2.24581
R56697 DVSS.n170 DVSS.n152 2.24581
R56698 DVSS.n172 DVSS.n153 2.24581
R56699 DVSS.n6456 DVSS.n6452 2.24581
R56700 DVSS.n174 DVSS.n152 2.24581
R56701 DVSS.n176 DVSS.n153 2.24581
R56702 DVSS.n6456 DVSS.n6451 2.24581
R56703 DVSS.n178 DVSS.n152 2.24581
R56704 DVSS.n6447 DVSS.n153 2.24581
R56705 DVSS.n6456 DVSS.n6450 2.24581
R56706 DVSS.n6449 DVSS.n152 2.24581
R56707 DVSS.n6457 DVSS.n6456 2.24581
R56708 DVSS.n155 DVSS.n152 2.24581
R56709 DVSS.n6456 DVSS.n151 2.24581
R56710 DVSS.n300 DVSS.n283 2.24581
R56711 DVSS.n6371 DVSS.n323 2.24581
R56712 DVSS.n302 DVSS.n283 2.24581
R56713 DVSS.n6371 DVSS.n322 2.24581
R56714 DVSS.n304 DVSS.n283 2.24581
R56715 DVSS.n6371 DVSS.n6367 2.24581
R56716 DVSS.n306 DVSS.n283 2.24581
R56717 DVSS.n308 DVSS.n283 2.24581
R56718 DVSS.n6371 DVSS.n6368 2.24581
R56719 DVSS.n310 DVSS.n283 2.24581
R56720 DVSS.n312 DVSS.n283 2.24581
R56721 DVSS.n6371 DVSS.n6369 2.24581
R56722 DVSS.n315 DVSS.n284 2.24581
R56723 DVSS.n316 DVSS.n283 2.24581
R56724 DVSS.n6371 DVSS.n6370 2.24581
R56725 DVSS.n319 DVSS.n284 2.24581
R56726 DVSS.n320 DVSS.n283 2.24581
R56727 DVSS.n6371 DVSS.n282 2.24581
R56728 DVSS.n476 DVSS.n462 2.24581
R56729 DVSS.n6196 DVSS.n6189 2.24581
R56730 DVSS.n478 DVSS.n462 2.24581
R56731 DVSS.n6196 DVSS.n463 2.24581
R56732 DVSS.n480 DVSS.n462 2.24581
R56733 DVSS.n6196 DVSS.n6190 2.24581
R56734 DVSS.n482 DVSS.n462 2.24581
R56735 DVSS.n6196 DVSS.n515 2.24581
R56736 DVSS.n485 DVSS.n462 2.24581
R56737 DVSS.n6196 DVSS.n514 2.24581
R56738 DVSS.n6196 DVSS.n6191 2.24581
R56739 DVSS.n6196 DVSS.n513 2.24581
R56740 DVSS.n6196 DVSS.n6192 2.24581
R56741 DVSS.n6193 DVSS.n465 2.24581
R56742 DVSS.n6199 DVSS.n489 2.24581
R56743 DVSS.n510 DVSS.n465 2.24581
R56744 DVSS.n6199 DVSS.n6198 2.24581
R56745 DVSS.n6196 DVSS.n6195 2.24581
R56746 DVSS.n1257 DVSS.n1254 2.24442
R56747 DVSS.n5681 DVSS.n1253 2.24442
R56748 DVSS.n6466 DVSS.n124 2.24442
R56749 DVSS.n6462 DVSS.n140 2.24442
R56750 DVSS.n6462 DVSS.n150 2.24442
R56751 DVSS.n6437 DVSS.n6436 2.24442
R56752 DVSS.n6398 DVSS.n210 2.24442
R56753 DVSS.n145 DVSS.n139 2.24442
R56754 DVSS.n147 DVSS.n139 2.24442
R56755 DVSS.n6418 DVSS.n220 2.24442
R56756 DVSS.n1758 DVSS.n1757 2.2436
R56757 DVSS.n4994 DVSS.n4993 2.2436
R56758 DVSS.n4994 DVSS.n1753 2.2436
R56759 DVSS.n1777 DVSS.n1774 2.2436
R56760 DVSS.n2423 DVSS.n2412 2.2436
R56761 DVSS.n2419 DVSS.n2413 2.2436
R56762 DVSS.n4962 DVSS.n1773 2.2436
R56763 DVSS.n1796 DVSS.n1795 2.2436
R56764 DVSS.n2613 DVSS.n2130 2.24321
R56765 DVSS.n3042 DVSS.n2126 2.24321
R56766 DVSS.n2430 DVSS.n2113 2.24321
R56767 DVSS.n3536 DVSS.n3535 2.24321
R56768 DVSS.n5702 DVSS.n5700 2.23892
R56769 DVSS.n5699 DVSS.n1247 2.23892
R56770 DVSS.n1233 DVSS.n1232 2.23892
R56771 DVSS.n500 DVSS.n499 2.23892
R56772 DVSS.n387 DVSS.n386 2.23892
R56773 DVSS.n1073 DVSS.n388 2.23892
R56774 DVSS.n5654 DVSS.n1299 2.23892
R56775 DVSS.n5589 DVSS.n1260 2.23892
R56776 DVSS.n1332 DVSS.n1331 2.23892
R56777 DVSS.n5655 DVSS.n1300 2.23892
R56778 DVSS.n5590 DVSS.n5587 2.23892
R56779 DVSS.n5598 DVSS.n5597 2.23892
R56780 DVSS.n1308 DVSS.n1307 2.23892
R56781 DVSS.n1311 DVSS.n1310 2.23892
R56782 DVSS.n493 DVSS.n219 2.23892
R56783 DVSS.n5713 DVSS.n5712 2.23892
R56784 DVSS.n5003 DVSS.n1729 2.2385
R56785 DVSS.n3039 DVSS.n3038 2.2385
R56786 DVSS.n3033 DVSS.n2407 2.2385
R56787 DVSS.n4999 DVSS.n4998 2.2385
R56788 DVSS.n4998 DVSS.n1732 2.2385
R56789 DVSS.n4936 DVSS.n1800 2.2385
R56790 DVSS.n5689 DVSS.n1249 2.23787
R56791 DVSS.n5687 DVSS.n1251 2.23787
R56792 DVSS.n1173 DVSS.n1172 2.23787
R56793 DVSS.n1177 DVSS.n1172 2.23787
R56794 DVSS.n6047 DVSS.n1178 2.23787
R56795 DVSS.n1184 DVSS.n1181 2.23787
R56796 DVSS.n6080 DVSS.n6079 2.23787
R56797 DVSS.n6079 DVSS.n1175 2.23787
R56798 DVSS.n1171 DVSS.n1170 2.23787
R56799 DVSS.n506 DVSS.n503 2.23787
R56800 DVSS.n508 DVSS.n491 2.23787
R56801 DVSS.n6088 DVSS.n6087 2.23787
R56802 DVSS.n1193 DVSS.n1183 2.23714
R56803 DVSS.n6071 DVSS.n1190 2.23714
R56804 DVSS.n1189 DVSS.n1183 2.23714
R56805 DVSS.n6071 DVSS.n1188 2.23714
R56806 DVSS.n1187 DVSS.n1183 2.23714
R56807 DVSS.n6069 DVSS.n1183 2.23714
R56808 DVSS.n5509 DVSS.n1364 2.23714
R56809 DVSS.n5552 DVSS.n1363 2.23714
R56810 DVSS.n5509 DVSS.n1365 2.23714
R56811 DVSS.n5552 DVSS.n1362 2.23714
R56812 DVSS.n5509 DVSS.n1366 2.23714
R56813 DVSS.n5552 DVSS.n1361 2.23714
R56814 DVSS.n5509 DVSS.n1367 2.23714
R56815 DVSS.n5552 DVSS.n1360 2.23714
R56816 DVSS.n5509 DVSS.n1368 2.23714
R56817 DVSS.n5552 DVSS.n1359 2.23714
R56818 DVSS.n5344 DVSS.n1548 2.23714
R56819 DVSS.n1547 DVSS.n1525 2.23714
R56820 DVSS.n5344 DVSS.n1546 2.23714
R56821 DVSS.n1545 DVSS.n1525 2.23714
R56822 DVSS.n5344 DVSS.n1544 2.23714
R56823 DVSS.n1543 DVSS.n1525 2.23714
R56824 DVSS.n5344 DVSS.n1542 2.23714
R56825 DVSS.n1541 DVSS.n1525 2.23714
R56826 DVSS.n5344 DVSS.n1540 2.23714
R56827 DVSS.n1539 DVSS.n1525 2.23714
R56828 DVSS.n5344 DVSS.n1538 2.23714
R56829 DVSS.n1537 DVSS.n1525 2.23714
R56830 DVSS.n5344 DVSS.n1536 2.23714
R56831 DVSS.n1535 DVSS.n1525 2.23714
R56832 DVSS.n5344 DVSS.n1534 2.23714
R56833 DVSS.n1533 DVSS.n1525 2.23714
R56834 DVSS.n5344 DVSS.n1532 2.23714
R56835 DVSS.n1531 DVSS.n1525 2.23714
R56836 DVSS.n5344 DVSS.n1530 2.23714
R56837 DVSS.n1529 DVSS.n1525 2.23714
R56838 DVSS.n5344 DVSS.n1528 2.23714
R56839 DVSS.n1526 DVSS.n1525 2.23714
R56840 DVSS.n5088 DVSS.n1680 2.23714
R56841 DVSS.n5131 DVSS.n1679 2.23714
R56842 DVSS.n5088 DVSS.n1681 2.23714
R56843 DVSS.n5131 DVSS.n1678 2.23714
R56844 DVSS.n5088 DVSS.n1682 2.23714
R56845 DVSS.n5131 DVSS.n1677 2.23714
R56846 DVSS.n5088 DVSS.n1683 2.23714
R56847 DVSS.n5131 DVSS.n1676 2.23714
R56848 DVSS.n5088 DVSS.n1684 2.23714
R56849 DVSS.n5131 DVSS.n1675 2.23714
R56850 DVSS.n1696 DVSS.n1685 2.23714
R56851 DVSS.n5085 DVSS.n1691 2.23714
R56852 DVSS.n1696 DVSS.n1692 2.23714
R56853 DVSS.n5085 DVSS.n1690 2.23714
R56854 DVSS.n1696 DVSS.n1693 2.23714
R56855 DVSS.n5085 DVSS.n1689 2.23714
R56856 DVSS.n1696 DVSS.n1694 2.23714
R56857 DVSS.n5085 DVSS.n1688 2.23714
R56858 DVSS.n1696 DVSS.n1695 2.23714
R56859 DVSS.n5085 DVSS.n1687 2.23714
R56860 DVSS.n2883 DVSS.n2612 2.23714
R56861 DVSS.n2880 DVSS.n2877 2.23714
R56862 DVSS.n2883 DVSS.n2615 2.23714
R56863 DVSS.n2881 DVSS.n2880 2.23714
R56864 DVSS.n2883 DVSS.n2882 2.23714
R56865 DVSS.n2880 DVSS.n2608 2.23714
R56866 DVSS.n2927 DVSS.n2886 2.23714
R56867 DVSS.n2607 DVSS.n2599 2.23714
R56868 DVSS.n2927 DVSS.n2606 2.23714
R56869 DVSS.n2605 DVSS.n2599 2.23714
R56870 DVSS.n2927 DVSS.n2604 2.23714
R56871 DVSS.n2603 DVSS.n2599 2.23714
R56872 DVSS.n2927 DVSS.n2602 2.23714
R56873 DVSS.n2601 DVSS.n2599 2.23714
R56874 DVSS.n2880 DVSS.n2876 2.23714
R56875 DVSS.n5345 DVSS.n5344 2.23714
R56876 DVSS.n1195 DVSS.n1183 2.23714
R56877 DVSS.n4966 DVSS.n1772 2.23714
R56878 DVSS.n4970 DVSS.n4969 2.23714
R56879 DVSS.n4973 DVSS.n1770 2.23714
R56880 DVSS.n4975 DVSS.n4974 2.23714
R56881 DVSS.n6049 DVSS.n5801 2.23714
R56882 DVSS.n6049 DVSS.n6045 2.23714
R56883 DVSS.n6052 DVSS.n5803 2.23714
R56884 DVSS.n6052 DVSS.n5806 2.23714
R56885 DVSS.n6049 DVSS.n6046 2.23714
R56886 DVSS.n6052 DVSS.n5807 2.23714
R56887 DVSS.n6050 DVSS.n6049 2.23714
R56888 DVSS.n4703 DVSS.n1334 2.23714
R56889 DVSS.n5585 DVSS.n1340 2.23714
R56890 DVSS.n4703 DVSS.n4698 2.23714
R56891 DVSS.n5585 DVSS.n1339 2.23714
R56892 DVSS.n4703 DVSS.n4699 2.23714
R56893 DVSS.n5585 DVSS.n1338 2.23714
R56894 DVSS.n4703 DVSS.n4700 2.23714
R56895 DVSS.n5585 DVSS.n1337 2.23714
R56896 DVSS.n4703 DVSS.n4701 2.23714
R56897 DVSS.n5585 DVSS.n1336 2.23714
R56898 DVSS.n5265 DVSS.n5263 2.23714
R56899 DVSS.n1590 DVSS.n1564 2.23714
R56900 DVSS.n5265 DVSS.n1589 2.23714
R56901 DVSS.n1588 DVSS.n1564 2.23714
R56902 DVSS.n5265 DVSS.n1587 2.23714
R56903 DVSS.n1586 DVSS.n1564 2.23714
R56904 DVSS.n5265 DVSS.n1585 2.23714
R56905 DVSS.n1584 DVSS.n1564 2.23714
R56906 DVSS.n5265 DVSS.n1583 2.23714
R56907 DVSS.n1582 DVSS.n1564 2.23714
R56908 DVSS.n5265 DVSS.n1581 2.23714
R56909 DVSS.n1580 DVSS.n1564 2.23714
R56910 DVSS.n5265 DVSS.n1579 2.23714
R56911 DVSS.n1578 DVSS.n1564 2.23714
R56912 DVSS.n5265 DVSS.n1577 2.23714
R56913 DVSS.n1576 DVSS.n1564 2.23714
R56914 DVSS.n5265 DVSS.n1575 2.23714
R56915 DVSS.n1574 DVSS.n1564 2.23714
R56916 DVSS.n5265 DVSS.n1573 2.23714
R56917 DVSS.n1572 DVSS.n1564 2.23714
R56918 DVSS.n5265 DVSS.n1571 2.23714
R56919 DVSS.n1570 DVSS.n1564 2.23714
R56920 DVSS.n5265 DVSS.n1569 2.23714
R56921 DVSS.n3756 DVSS.n1650 2.23714
R56922 DVSS.n5164 DVSS.n1656 2.23714
R56923 DVSS.n3756 DVSS.n3750 2.23714
R56924 DVSS.n5164 DVSS.n1655 2.23714
R56925 DVSS.n3756 DVSS.n3751 2.23714
R56926 DVSS.n5164 DVSS.n1654 2.23714
R56927 DVSS.n3756 DVSS.n3752 2.23714
R56928 DVSS.n5164 DVSS.n1653 2.23714
R56929 DVSS.n3756 DVSS.n3753 2.23714
R56930 DVSS.n5164 DVSS.n1652 2.23714
R56931 DVSS.n5007 DVSS.n1721 2.23714
R56932 DVSS.n5007 DVSS.n1723 2.23714
R56933 DVSS.n1722 DVSS.n1713 2.23714
R56934 DVSS.n1724 DVSS.n1713 2.23714
R56935 DVSS.n5007 DVSS.n1725 2.23714
R56936 DVSS.n1726 DVSS.n1713 2.23714
R56937 DVSS.n2405 DVSS.n2401 2.23714
R56938 DVSS.n3044 DVSS.n2403 2.23714
R56939 DVSS.n3047 DVSS.n2401 2.23714
R56940 DVSS.n3046 DVSS.n3044 2.23714
R56941 DVSS.n3048 DVSS.n3044 2.23714
R56942 DVSS.n3049 DVSS.n2401 2.23714
R56943 DVSS.n3050 DVSS.n3044 2.23714
R56944 DVSS.n3053 DVSS.n2399 2.23714
R56945 DVSS.n3054 DVSS.n2400 2.23714
R56946 DVSS.n3055 DVSS.n2399 2.23714
R56947 DVSS.n3056 DVSS.n2400 2.23714
R56948 DVSS.n3057 DVSS.n2399 2.23714
R56949 DVSS.n3058 DVSS.n2400 2.23714
R56950 DVSS.n3059 DVSS.n2399 2.23714
R56951 DVSS.n3060 DVSS.n2400 2.23714
R56952 DVSS.n1791 DVSS.n1790 2.23714
R56953 DVSS.n4949 DVSS.n4948 2.23714
R56954 DVSS.n4952 DVSS.n1788 2.23714
R56955 DVSS.n1789 DVSS.n1787 2.23714
R56956 DVSS.n3029 DVSS.n1786 2.23714
R56957 DVSS.n6099 DVSS.n1142 2.23714
R56958 DVSS.n6099 DVSS.n1153 2.23714
R56959 DVSS.n6102 DVSS.n1145 2.23714
R56960 DVSS.n6102 DVSS.n1148 2.23714
R56961 DVSS.n6099 DVSS.n1154 2.23714
R56962 DVSS.n6102 DVSS.n1149 2.23714
R56963 DVSS.n6100 DVSS.n6099 2.23714
R56964 DVSS.n4645 DVSS.n2017 2.23714
R56965 DVSS.n2018 DVSS.n2011 2.23714
R56966 DVSS.n4645 DVSS.n2019 2.23714
R56967 DVSS.n2020 DVSS.n2011 2.23714
R56968 DVSS.n4645 DVSS.n2021 2.23714
R56969 DVSS.n2022 DVSS.n2011 2.23714
R56970 DVSS.n4645 DVSS.n2023 2.23714
R56971 DVSS.n2024 DVSS.n2011 2.23714
R56972 DVSS.n4645 DVSS.n2025 2.23714
R56973 DVSS.n4643 DVSS.n2011 2.23714
R56974 DVSS.n4636 DVSS.n2026 2.23714
R56975 DVSS.n4639 DVSS.n2029 2.23714
R56976 DVSS.n4636 DVSS.n4635 2.23714
R56977 DVSS.n4639 DVSS.n2030 2.23714
R56978 DVSS.n4636 DVSS.n4634 2.23714
R56979 DVSS.n4639 DVSS.n2031 2.23714
R56980 DVSS.n4636 DVSS.n4633 2.23714
R56981 DVSS.n4639 DVSS.n2032 2.23714
R56982 DVSS.n4636 DVSS.n4632 2.23714
R56983 DVSS.n4639 DVSS.n2033 2.23714
R56984 DVSS.n4636 DVSS.n4631 2.23714
R56985 DVSS.n4639 DVSS.n2034 2.23714
R56986 DVSS.n4636 DVSS.n4630 2.23714
R56987 DVSS.n4639 DVSS.n2035 2.23714
R56988 DVSS.n4636 DVSS.n4629 2.23714
R56989 DVSS.n4639 DVSS.n2036 2.23714
R56990 DVSS.n4636 DVSS.n4628 2.23714
R56991 DVSS.n4639 DVSS.n2037 2.23714
R56992 DVSS.n4636 DVSS.n4627 2.23714
R56993 DVSS.n4639 DVSS.n2038 2.23714
R56994 DVSS.n4636 DVSS.n4626 2.23714
R56995 DVSS.n4639 DVSS.n2039 2.23714
R56996 DVSS.n4637 DVSS.n4636 2.23714
R56997 DVSS.n4915 DVSS.n1801 2.23714
R56998 DVSS.n4916 DVSS.n1802 2.23714
R56999 DVSS.n4917 DVSS.n1801 2.23714
R57000 DVSS.n4918 DVSS.n1802 2.23714
R57001 DVSS.n4919 DVSS.n1801 2.23714
R57002 DVSS.n4920 DVSS.n1802 2.23714
R57003 DVSS.n4921 DVSS.n1801 2.23714
R57004 DVSS.n4922 DVSS.n1802 2.23714
R57005 DVSS.n4923 DVSS.n1801 2.23714
R57006 DVSS.n4924 DVSS.n1802 2.23714
R57007 DVSS.n4927 DVSS.n1798 2.23714
R57008 DVSS.n4939 DVSS.n1798 2.23714
R57009 DVSS.n4938 DVSS.n1799 2.23714
R57010 DVSS.n4940 DVSS.n1799 2.23714
R57011 DVSS.n4941 DVSS.n1798 2.23714
R57012 DVSS.n4942 DVSS.n1799 2.23714
R57013 DVSS.n3023 DVSS.n2424 2.23714
R57014 DVSS.n3026 DVSS.n2428 2.23714
R57015 DVSS.n3024 DVSS.n3023 2.23714
R57016 DVSS.n3026 DVSS.n3025 2.23714
R57017 DVSS.n3026 DVSS.n2427 2.23714
R57018 DVSS.n3023 DVSS.n3022 2.23714
R57019 DVSS.n3026 DVSS.n2426 2.23714
R57020 DVSS.n3017 DVSS.n2434 2.23714
R57021 DVSS.n3019 DVSS.n2437 2.23714
R57022 DVSS.n3017 DVSS.n3016 2.23714
R57023 DVSS.n3019 DVSS.n2438 2.23714
R57024 DVSS.n3017 DVSS.n3015 2.23714
R57025 DVSS.n3019 DVSS.n2439 2.23714
R57026 DVSS.n3017 DVSS.n3014 2.23714
R57027 DVSS.n3019 DVSS.n2440 2.23714
R57028 DVSS.n6090 DVSS.n1158 2.23714
R57029 DVSS.n6090 DVSS.n1168 2.23714
R57030 DVSS.n6093 DVSS.n1161 2.23714
R57031 DVSS.n6093 DVSS.n1163 2.23714
R57032 DVSS.n6090 DVSS.n1169 2.23714
R57033 DVSS.n6093 DVSS.n1164 2.23714
R57034 DVSS.n6091 DVSS.n6090 2.23714
R57035 DVSS.n3943 DVSS.n3895 2.23714
R57036 DVSS.n3944 DVSS.n3941 2.23714
R57037 DVSS.n3945 DVSS.n3895 2.23714
R57038 DVSS.n3946 DVSS.n3941 2.23714
R57039 DVSS.n3947 DVSS.n3895 2.23714
R57040 DVSS.n3948 DVSS.n3941 2.23714
R57041 DVSS.n3949 DVSS.n3895 2.23714
R57042 DVSS.n3950 DVSS.n3941 2.23714
R57043 DVSS.n3951 DVSS.n3895 2.23714
R57044 DVSS.n3952 DVSS.n3941 2.23714
R57045 DVSS.n4445 DVSS.n4444 2.23714
R57046 DVSS.n4448 DVSS.n2058 2.23714
R57047 DVSS.n4445 DVSS.n4443 2.23714
R57048 DVSS.n4448 DVSS.n2059 2.23714
R57049 DVSS.n4445 DVSS.n4442 2.23714
R57050 DVSS.n4448 DVSS.n2060 2.23714
R57051 DVSS.n4445 DVSS.n4441 2.23714
R57052 DVSS.n4448 DVSS.n2061 2.23714
R57053 DVSS.n4445 DVSS.n4440 2.23714
R57054 DVSS.n4448 DVSS.n2062 2.23714
R57055 DVSS.n4445 DVSS.n4439 2.23714
R57056 DVSS.n4448 DVSS.n2063 2.23714
R57057 DVSS.n4445 DVSS.n4438 2.23714
R57058 DVSS.n4448 DVSS.n2064 2.23714
R57059 DVSS.n4445 DVSS.n4437 2.23714
R57060 DVSS.n4448 DVSS.n2065 2.23714
R57061 DVSS.n4445 DVSS.n4436 2.23714
R57062 DVSS.n4448 DVSS.n2066 2.23714
R57063 DVSS.n4445 DVSS.n4435 2.23714
R57064 DVSS.n4448 DVSS.n2067 2.23714
R57065 DVSS.n4445 DVSS.n4434 2.23714
R57066 DVSS.n4448 DVSS.n2068 2.23714
R57067 DVSS.n4446 DVSS.n4445 2.23714
R57068 DVSS.n3695 DVSS.n2069 2.23714
R57069 DVSS.n3883 DVSS.n2075 2.23714
R57070 DVSS.n3695 DVSS.n2079 2.23714
R57071 DVSS.n3883 DVSS.n2074 2.23714
R57072 DVSS.n3695 DVSS.n2080 2.23714
R57073 DVSS.n3883 DVSS.n2073 2.23714
R57074 DVSS.n3695 DVSS.n2081 2.23714
R57075 DVSS.n3883 DVSS.n2072 2.23714
R57076 DVSS.n3695 DVSS.n2082 2.23714
R57077 DVSS.n3883 DVSS.n2071 2.23714
R57078 DVSS.n3546 DVSS.n2083 2.23714
R57079 DVSS.n3692 DVSS.n2089 2.23714
R57080 DVSS.n3546 DVSS.n2093 2.23714
R57081 DVSS.n3692 DVSS.n2088 2.23714
R57082 DVSS.n3546 DVSS.n2094 2.23714
R57083 DVSS.n3692 DVSS.n2087 2.23714
R57084 DVSS.n3546 DVSS.n2095 2.23714
R57085 DVSS.n3692 DVSS.n2086 2.23714
R57086 DVSS.n3546 DVSS.n2096 2.23714
R57087 DVSS.n3692 DVSS.n2085 2.23714
R57088 DVSS.n3540 DVSS.n2097 2.23714
R57089 DVSS.n3543 DVSS.n2102 2.23714
R57090 DVSS.n3541 DVSS.n3540 2.23714
R57091 DVSS.n3543 DVSS.n3542 2.23714
R57092 DVSS.n3543 DVSS.n2100 2.23714
R57093 DVSS.n3540 DVSS.n2108 2.23714
R57094 DVSS.n3543 DVSS.n2099 2.23714
R57095 DVSS.n2470 DVSS.n2469 2.23714
R57096 DVSS.n2472 DVSS.n2459 2.23714
R57097 DVSS.n2470 DVSS.n2468 2.23714
R57098 DVSS.n2472 DVSS.n2460 2.23714
R57099 DVSS.n2470 DVSS.n2467 2.23714
R57100 DVSS.n2472 DVSS.n2461 2.23714
R57101 DVSS.n2470 DVSS.n2466 2.23714
R57102 DVSS.n2472 DVSS.n2462 2.23714
R57103 DVSS.n242 DVSS.n223 2.23714
R57104 DVSS.n238 DVSS.n223 2.23714
R57105 DVSS.n6421 DVSS.n237 2.23714
R57106 DVSS.n244 DVSS.n223 2.23714
R57107 DVSS.n235 DVSS.n223 2.23714
R57108 DVSS.n6421 DVSS.n234 2.23714
R57109 DVSS.n6411 DVSS.n223 2.23714
R57110 DVSS.n232 DVSS.n223 2.23714
R57111 DVSS.n6421 DVSS.n231 2.23714
R57112 DVSS.n6416 DVSS.n223 2.23714
R57113 DVSS.n229 DVSS.n223 2.23714
R57114 DVSS.n6421 DVSS.n228 2.23714
R57115 DVSS.n227 DVSS.n223 2.23714
R57116 DVSS.n6421 DVSS.n226 2.23714
R57117 DVSS.n6419 DVSS.n223 2.23714
R57118 DVSS.n6470 DVSS.n108 2.23714
R57119 DVSS.n6472 DVSS.n119 2.23714
R57120 DVSS.n6470 DVSS.n132 2.23714
R57121 DVSS.n6472 DVSS.n116 2.23714
R57122 DVSS.n6472 DVSS.n120 2.23714
R57123 DVSS.n6470 DVSS.n130 2.23714
R57124 DVSS.n6472 DVSS.n115 2.23714
R57125 DVSS.n6472 DVSS.n121 2.23714
R57126 DVSS.n6470 DVSS.n128 2.23714
R57127 DVSS.n6472 DVSS.n114 2.23714
R57128 DVSS.n6472 DVSS.n122 2.23714
R57129 DVSS.n6470 DVSS.n126 2.23714
R57130 DVSS.n6472 DVSS.n113 2.23714
R57131 DVSS.n6470 DVSS.n125 2.23714
R57132 DVSS.n6472 DVSS.n112 2.23714
R57133 DVSS.n6439 DVSS.n194 2.23714
R57134 DVSS.n207 DVSS.n204 2.23714
R57135 DVSS.n6439 DVSS.n191 2.23714
R57136 DVSS.n207 DVSS.n203 2.23714
R57137 DVSS.n207 DVSS.n205 2.23714
R57138 DVSS.n6439 DVSS.n189 2.23714
R57139 DVSS.n207 DVSS.n202 2.23714
R57140 DVSS.n207 DVSS.n206 2.23714
R57141 DVSS.n6439 DVSS.n187 2.23714
R57142 DVSS.n207 DVSS.n201 2.23714
R57143 DVSS.n207 DVSS.n182 2.23714
R57144 DVSS.n6439 DVSS.n186 2.23714
R57145 DVSS.n207 DVSS.n200 2.23714
R57146 DVSS.n6439 DVSS.n185 2.23714
R57147 DVSS.n207 DVSS.n199 2.23714
R57148 DVSS.n6400 DVSS.n259 2.23714
R57149 DVSS.n6397 DVSS.n6394 2.23714
R57150 DVSS.n6400 DVSS.n256 2.23714
R57151 DVSS.n6397 DVSS.n278 2.23714
R57152 DVSS.n6397 DVSS.n6395 2.23714
R57153 DVSS.n6400 DVSS.n254 2.23714
R57154 DVSS.n6397 DVSS.n277 2.23714
R57155 DVSS.n6397 DVSS.n248 2.23714
R57156 DVSS.n6400 DVSS.n253 2.23714
R57157 DVSS.n6397 DVSS.n276 2.23714
R57158 DVSS.n6397 DVSS.n6396 2.23714
R57159 DVSS.n6400 DVSS.n251 2.23714
R57160 DVSS.n6397 DVSS.n275 2.23714
R57161 DVSS.n6400 DVSS.n250 2.23714
R57162 DVSS.n6397 DVSS.n274 2.23714
R57163 DVSS.n6489 DVSS.n61 2.23714
R57164 DVSS.n6486 DVSS.n73 2.23714
R57165 DVSS.n6489 DVSS.n62 2.23714
R57166 DVSS.n6486 DVSS.n74 2.23714
R57167 DVSS.n6489 DVSS.n58 2.23714
R57168 DVSS.n6486 DVSS.n71 2.23714
R57169 DVSS.n6489 DVSS.n57 2.23714
R57170 DVSS.n6489 DVSS.n56 2.23714
R57171 DVSS.n6486 DVSS.n69 2.23714
R57172 DVSS.n6489 DVSS.n55 2.23714
R57173 DVSS.n6489 DVSS.n54 2.23714
R57174 DVSS.n6486 DVSS.n67 2.23714
R57175 DVSS.n6486 DVSS.n6485 2.23714
R57176 DVSS.n6489 DVSS.n52 2.23714
R57177 DVSS.n6486 DVSS.n66 2.23714
R57178 DVSS.n6486 DVSS.n49 2.23714
R57179 DVSS.n6489 DVSS.n51 2.23714
R57180 DVSS.n6487 DVSS.n6486 2.23714
R57181 DVSS.n6476 DVSS.n103 2.23714
R57182 DVSS.n6479 DVSS.n89 2.23714
R57183 DVSS.n6476 DVSS.n104 2.23714
R57184 DVSS.n6479 DVSS.n90 2.23714
R57185 DVSS.n6476 DVSS.n100 2.23714
R57186 DVSS.n6479 DVSS.n86 2.23714
R57187 DVSS.n6476 DVSS.n99 2.23714
R57188 DVSS.n6476 DVSS.n98 2.23714
R57189 DVSS.n6479 DVSS.n84 2.23714
R57190 DVSS.n6476 DVSS.n97 2.23714
R57191 DVSS.n6476 DVSS.n79 2.23714
R57192 DVSS.n6479 DVSS.n83 2.23714
R57193 DVSS.n6479 DVSS.n93 2.23714
R57194 DVSS.n6476 DVSS.n95 2.23714
R57195 DVSS.n6479 DVSS.n82 2.23714
R57196 DVSS.n6479 DVSS.n6478 2.23714
R57197 DVSS.n6476 DVSS.n94 2.23714
R57198 DVSS.n6479 DVSS.n81 2.23714
R57199 DVSS.n6297 DVSS.n364 2.23714
R57200 DVSS.n6294 DVSS.n6260 2.23714
R57201 DVSS.n6297 DVSS.n365 2.23714
R57202 DVSS.n6294 DVSS.n6261 2.23714
R57203 DVSS.n6297 DVSS.n362 2.23714
R57204 DVSS.n6294 DVSS.n385 2.23714
R57205 DVSS.n6297 DVSS.n361 2.23714
R57206 DVSS.n6297 DVSS.n360 2.23714
R57207 DVSS.n6294 DVSS.n383 2.23714
R57208 DVSS.n6297 DVSS.n359 2.23714
R57209 DVSS.n6297 DVSS.n358 2.23714
R57210 DVSS.n6294 DVSS.n381 2.23714
R57211 DVSS.n6294 DVSS.n6292 2.23714
R57212 DVSS.n6297 DVSS.n356 2.23714
R57213 DVSS.n6294 DVSS.n380 2.23714
R57214 DVSS.n6294 DVSS.n6293 2.23714
R57215 DVSS.n6297 DVSS.n354 2.23714
R57216 DVSS.n6295 DVSS.n6294 2.23714
R57217 DVSS.n31 DVSS.n15 2.23714
R57218 DVSS.n6500 DVSS.n32 2.23714
R57219 DVSS.n33 DVSS.n15 2.23714
R57220 DVSS.n6500 DVSS.n34 2.23714
R57221 DVSS.n35 DVSS.n15 2.23714
R57222 DVSS.n6500 DVSS.n28 2.23714
R57223 DVSS.n27 DVSS.n15 2.23714
R57224 DVSS.n37 DVSS.n15 2.23714
R57225 DVSS.n6500 DVSS.n25 2.23714
R57226 DVSS.n24 DVSS.n15 2.23714
R57227 DVSS.n39 DVSS.n15 2.23714
R57228 DVSS.n6500 DVSS.n22 2.23714
R57229 DVSS.n6500 DVSS.n42 2.23714
R57230 DVSS.n41 DVSS.n15 2.23714
R57231 DVSS.n6500 DVSS.n21 2.23714
R57232 DVSS.n6500 DVSS.n6499 2.23714
R57233 DVSS.n43 DVSS.n15 2.23714
R57234 DVSS.n6500 DVSS.n20 2.23714
R57235 DVSS.n6241 DVSS.n404 2.23714
R57236 DVSS.n6238 DVSS.n418 2.23714
R57237 DVSS.n6238 DVSS.n420 2.23714
R57238 DVSS.n6241 DVSS.n406 2.23714
R57239 DVSS.n6238 DVSS.n417 2.23714
R57240 DVSS.n6238 DVSS.n421 2.23714
R57241 DVSS.n6241 DVSS.n402 2.23714
R57242 DVSS.n6238 DVSS.n416 2.23714
R57243 DVSS.n6238 DVSS.n422 2.23714
R57244 DVSS.n6241 DVSS.n408 2.23714
R57245 DVSS.n6238 DVSS.n415 2.23714
R57246 DVSS.n6238 DVSS.n423 2.23714
R57247 DVSS.n6241 DVSS.n400 2.23714
R57248 DVSS.n6238 DVSS.n414 2.23714
R57249 DVSS.n6238 DVSS.n396 2.23714
R57250 DVSS.n6241 DVSS.n412 2.23714
R57251 DVSS.n6239 DVSS.n6238 2.23714
R57252 DVSS.n6241 DVSS.n6240 2.23714
R57253 DVSS.n6229 DVSS.n449 2.23714
R57254 DVSS.n6232 DVSS.n434 2.23714
R57255 DVSS.n6232 DVSS.n436 2.23714
R57256 DVSS.n6229 DVSS.n450 2.23714
R57257 DVSS.n6232 DVSS.n433 2.23714
R57258 DVSS.n6232 DVSS.n437 2.23714
R57259 DVSS.n6229 DVSS.n447 2.23714
R57260 DVSS.n6232 DVSS.n432 2.23714
R57261 DVSS.n6232 DVSS.n438 2.23714
R57262 DVSS.n6229 DVSS.n452 2.23714
R57263 DVSS.n6232 DVSS.n431 2.23714
R57264 DVSS.n6232 DVSS.n439 2.23714
R57265 DVSS.n6229 DVSS.n427 2.23714
R57266 DVSS.n6232 DVSS.n430 2.23714
R57267 DVSS.n6232 DVSS.n440 2.23714
R57268 DVSS.n6230 DVSS.n6229 2.23714
R57269 DVSS.n6232 DVSS.n6231 2.23714
R57270 DVSS.n6229 DVSS.n441 2.23714
R57271 DVSS.n6216 DVSS.n390 2.23714
R57272 DVSS.n6215 DVSS.n389 2.23714
R57273 DVSS.n6217 DVSS.n389 2.23714
R57274 DVSS.n6212 DVSS.n390 2.23714
R57275 DVSS.n6213 DVSS.n389 2.23714
R57276 DVSS.n6211 DVSS.n389 2.23714
R57277 DVSS.n1119 DVSS.n390 2.23714
R57278 DVSS.n1118 DVSS.n389 2.23714
R57279 DVSS.n1120 DVSS.n389 2.23714
R57280 DVSS.n1125 DVSS.n390 2.23714
R57281 DVSS.n1124 DVSS.n389 2.23714
R57282 DVSS.n1126 DVSS.n389 2.23714
R57283 DVSS.n1131 DVSS.n390 2.23714
R57284 DVSS.n1130 DVSS.n389 2.23714
R57285 DVSS.n6251 DVSS.n389 2.23714
R57286 DVSS.n6252 DVSS.n390 2.23714
R57287 DVSS.n6253 DVSS.n389 2.23714
R57288 DVSS.n6254 DVSS.n390 2.23714
R57289 DVSS.n1086 DVSS.n1071 2.23714
R57290 DVSS.n6131 DVSS.n1083 2.23714
R57291 DVSS.n6131 DVSS.n1087 2.23714
R57292 DVSS.n1089 DVSS.n1071 2.23714
R57293 DVSS.n6131 DVSS.n1081 2.23714
R57294 DVSS.n6131 DVSS.n1090 2.23714
R57295 DVSS.n1091 DVSS.n1071 2.23714
R57296 DVSS.n6131 DVSS.n1079 2.23714
R57297 DVSS.n6131 DVSS.n1092 2.23714
R57298 DVSS.n1093 DVSS.n1071 2.23714
R57299 DVSS.n6131 DVSS.n1077 2.23714
R57300 DVSS.n6131 DVSS.n1094 2.23714
R57301 DVSS.n6124 DVSS.n1071 2.23714
R57302 DVSS.n6131 DVSS.n1076 2.23714
R57303 DVSS.n6131 DVSS.n6127 2.23714
R57304 DVSS.n6129 DVSS.n1071 2.23714
R57305 DVSS.n6131 DVSS.n6130 2.23714
R57306 DVSS.n6128 DVSS.n1071 2.23714
R57307 DVSS.n2925 DVSS.n2133 2.21947
R57308 DVSS.n3063 DVSS.n3062 2.21947
R57309 DVSS.n6442 DVSS.n6441 2.21947
R57310 DVSS.n6404 DVSS.n6403 2.21947
R57311 DVSS.n268 DVSS.n260 2.21947
R57312 DVSS.n6391 DVSS.n6383 2.21947
R57313 DVSS.n6379 DVSS.n281 2.21947
R57314 DVSS.n6496 DVSS.n45 2.21947
R57315 DVSS.n377 DVSS.n376 2.21947
R57316 DVSS.n6290 DVSS.n6289 2.21947
R57317 DVSS.n6283 DVSS.n6282 2.21947
R57318 DVSS.n6272 DVSS.n6271 2.21947
R57319 DVSS.n6249 DVSS.n6248 2.21947
R57320 DVSS.n6220 DVSS.n6219 2.21947
R57321 DVSS.n6209 DVSS.n6208 2.21947
R57322 DVSS.n1122 DVSS.n1117 2.21947
R57323 DVSS.n1128 DVSS.n1106 2.21947
R57324 DVSS.n6122 DVSS.n1133 2.21947
R57325 DVSS.n6115 DVSS.n6114 2.21947
R57326 DVSS.n6113 DVSS.n6112 2.21947
R57327 DVSS.n5783 DVSS.n1137 2.21947
R57328 DVSS.n6055 DVSS.n6054 2.21947
R57329 DVSS.n6067 DVSS.n1198 2.21947
R57330 DVSS.n5770 DVSS.n5769 2.21947
R57331 DVSS.n5768 DVSS.n5767 2.21947
R57332 DVSS.n1212 DVSS.n1201 2.21947
R57333 DVSS.n5750 DVSS.n5749 2.21947
R57334 DVSS.n5748 DVSS.n5747 2.21947
R57335 DVSS.n1225 DVSS.n1215 2.21947
R57336 DVSS.n5733 DVSS.n5732 2.21947
R57337 DVSS.n5731 DVSS.n5730 2.21947
R57338 DVSS.n5693 DVSS.n1228 2.21947
R57339 DVSS.n5704 DVSS.n1245 2.21947
R57340 DVSS.n5706 DVSS.n5705 2.21947
R57341 DVSS.n5641 DVSS.n1242 2.21947
R57342 DVSS.n5638 DVSS.n1323 2.21947
R57343 DVSS.n5630 DVSS.n5629 2.21947
R57344 DVSS.n5628 DVSS.n5627 2.21947
R57345 DVSS.n5621 DVSS.n1326 2.21947
R57346 DVSS.n5613 DVSS.n5612 2.21947
R57347 DVSS.n5611 DVSS.n5610 2.21947
R57348 DVSS.n5604 DVSS.n1330 2.21947
R57349 DVSS.n3065 DVSS.n3064 2.21947
R57350 DVSS.n6445 DVSS.n179 2.21947
R57351 DVSS.n6407 DVSS.n6406 2.21947
R57352 DVSS.n265 DVSS.n261 2.21947
R57353 DVSS.n6388 DVSS.n6384 2.21947
R57354 DVSS.n6376 DVSS.n6375 2.21947
R57355 DVSS.n6493 DVSS.n46 2.21947
R57356 DVSS.n373 DVSS.n369 2.21947
R57357 DVSS.n6286 DVSS.n77 2.21947
R57358 DVSS.n6279 DVSS.n6275 2.21947
R57359 DVSS.n6268 DVSS.n6264 2.21947
R57360 DVSS.n6245 DVSS.n393 2.21947
R57361 DVSS.n6223 DVSS.n6222 2.21947
R57362 DVSS.n6205 DVSS.n6201 2.21947
R57363 DVSS.n1114 DVSS.n1110 2.21947
R57364 DVSS.n1103 DVSS.n1099 2.21947
R57365 DVSS.n6119 DVSS.n425 2.21947
R57366 DVSS.n6118 DVSS.n1136 2.21947
R57367 DVSS.n6109 DVSS.n1134 2.21947
R57368 DVSS.n5786 DVSS.n1141 2.21947
R57369 DVSS.n6058 DVSS.n1156 2.21947
R57370 DVSS.n6064 DVSS.n6062 2.21947
R57371 DVSS.n5773 DVSS.n1200 2.21947
R57372 DVSS.n5764 DVSS.n1199 2.21947
R57373 DVSS.n1209 DVSS.n1205 2.21947
R57374 DVSS.n5753 DVSS.n5752 2.21947
R57375 DVSS.n5744 DVSS.n1208 2.21947
R57376 DVSS.n1222 DVSS.n1218 2.21947
R57377 DVSS.n5736 DVSS.n5735 2.21947
R57378 DVSS.n5727 DVSS.n1221 2.21947
R57379 DVSS.n5690 DVSS.n1231 2.21947
R57380 DVSS.n1240 DVSS.n1236 2.21947
R57381 DVSS.n5709 DVSS.n5708 2.21947
R57382 DVSS.n5643 DVSS.n1239 2.21947
R57383 DVSS.n5635 DVSS.n5634 2.21947
R57384 DVSS.n5633 DVSS.n1325 2.21947
R57385 DVSS.n5624 DVSS.n1324 2.21947
R57386 DVSS.n5618 DVSS.n5617 2.21947
R57387 DVSS.n5616 DVSS.n1329 2.21947
R57388 DVSS.n5607 DVSS.n1328 2.21947
R57389 DVSS.n5601 DVSS.n5600 2.21947
R57390 DVSS.n3067 DVSS.n2394 2.21947
R57391 DVSS.n6414 DVSS.n6413 2.21947
R57392 DVSS.n6409 DVSS.n6408 2.21947
R57393 DVSS.n264 DVSS.n262 2.21947
R57394 DVSS.n6387 DVSS.n6385 2.21947
R57395 DVSS.n6474 DVSS.n107 2.21947
R57396 DVSS.n6492 DVSS.n47 2.21947
R57397 DVSS.n372 DVSS.n370 2.21947
R57398 DVSS.n6482 DVSS.n6481 2.21947
R57399 DVSS.n6278 DVSS.n6276 2.21947
R57400 DVSS.n6267 DVSS.n6265 2.21947
R57401 DVSS.n6244 DVSS.n394 2.21947
R57402 DVSS.n6226 DVSS.n6225 2.21947
R57403 DVSS.n6204 DVSS.n6202 2.21947
R57404 DVSS.n1113 DVSS.n1111 2.21947
R57405 DVSS.n1102 DVSS.n1100 2.21947
R57406 DVSS.n6235 DVSS.n6234 2.21947
R57407 DVSS.n1135 DVSS.n426 2.21947
R57408 DVSS.n6108 DVSS.n1139 2.21947
R57409 DVSS.n6105 DVSS.n6104 2.21947
R57410 DVSS.n6097 DVSS.n6096 2.21947
R57411 DVSS.n6063 DVSS.n1151 2.21947
R57412 DVSS.n5760 DVSS.n5759 2.21947
R57413 DVSS.n5763 DVSS.n1203 2.21947
R57414 DVSS.n5757 DVSS.n5756 2.21947
R57415 DVSS.n5755 DVSS.n5754 2.21947
R57416 DVSS.n5743 DVSS.n1206 2.21947
R57417 DVSS.n5740 DVSS.n5739 2.21947
R57418 DVSS.n5738 DVSS.n5737 2.21947
R57419 DVSS.n5726 DVSS.n1219 2.21947
R57420 DVSS.n5723 DVSS.n5722 2.21947
R57421 DVSS.n5718 DVSS.n5717 2.21947
R57422 DVSS.n5710 DVSS.n1235 2.21947
R57423 DVSS.n5645 DVSS.n5644 2.21947
R57424 DVSS.n5646 DVSS.n1320 2.21947
R57425 DVSS.n5647 DVSS.n1306 2.21947
R57426 DVSS.n5648 DVSS.n1305 2.21947
R57427 DVSS.n5649 DVSS.n1304 2.21947
R57428 DVSS.n5650 DVSS.n1303 2.21947
R57429 DVSS.n5651 DVSS.n1302 2.21947
R57430 DVSS.n5652 DVSS.n1301 2.21947
R57431 DVSS.n3068 DVSS.n2393 2.21947
R57432 DVSS.n5594 DVSS.n5593 2.16043
R57433 DVSS.n5392 DVSS.n1373 1.95638
R57434 DVSS.n5392 DVSS.n5391 1.95638
R57435 DVSS.n5356 DVSS.n1378 1.95638
R57436 DVSS.n5359 DVSS.n5356 1.95638
R57437 DVSS.n5351 DVSS.n1521 1.95638
R57438 DVSS.n5354 DVSS.n1521 1.95638
R57439 DVSS.n4318 DVSS.n4004 1.89035
R57440 DVSS.n4326 DVSS.n4005 1.89035
R57441 DVSS.n4318 DVSS.n4006 1.89035
R57442 DVSS.n4321 DVSS.n4005 1.89035
R57443 DVSS.n4319 DVSS.n4318 1.89035
R57444 DVSS.n4070 DVSS.n4005 1.89035
R57445 DVSS.n4318 DVSS.n4059 1.89035
R57446 DVSS.n4075 DVSS.n4005 1.89035
R57447 DVSS.n4318 DVSS.n4058 1.89035
R57448 DVSS.n4080 DVSS.n4005 1.89035
R57449 DVSS.n4318 DVSS.n4057 1.89035
R57450 DVSS.n4085 DVSS.n4005 1.89035
R57451 DVSS.n4318 DVSS.n4056 1.89035
R57452 DVSS.n4090 DVSS.n4005 1.89035
R57453 DVSS.n4318 DVSS.n4055 1.89035
R57454 DVSS.n4095 DVSS.n4005 1.89035
R57455 DVSS.n4318 DVSS.n4054 1.89035
R57456 DVSS.n4100 DVSS.n4005 1.89035
R57457 DVSS.n4318 DVSS.n4053 1.89035
R57458 DVSS.n4105 DVSS.n4005 1.89035
R57459 DVSS.n4318 DVSS.n4052 1.89035
R57460 DVSS.n4110 DVSS.n4005 1.89035
R57461 DVSS.n4318 DVSS.n4051 1.89035
R57462 DVSS.n4115 DVSS.n4005 1.89035
R57463 DVSS.n4318 DVSS.n4050 1.89035
R57464 DVSS.n4120 DVSS.n4005 1.89035
R57465 DVSS.n4318 DVSS.n4049 1.89035
R57466 DVSS.n4126 DVSS.n4005 1.89035
R57467 DVSS.n4318 DVSS.n4048 1.89035
R57468 DVSS.n4131 DVSS.n4005 1.89035
R57469 DVSS.n4318 DVSS.n4047 1.89035
R57470 DVSS.n4136 DVSS.n4005 1.89035
R57471 DVSS.n4318 DVSS.n4046 1.89035
R57472 DVSS.n4141 DVSS.n4005 1.89035
R57473 DVSS.n4318 DVSS.n4045 1.89035
R57474 DVSS.n4146 DVSS.n4005 1.89035
R57475 DVSS.n4318 DVSS.n4044 1.89035
R57476 DVSS.n4151 DVSS.n4005 1.89035
R57477 DVSS.n4318 DVSS.n4043 1.89035
R57478 DVSS.n4156 DVSS.n4005 1.89035
R57479 DVSS.n4318 DVSS.n4042 1.89035
R57480 DVSS.n4161 DVSS.n4005 1.89035
R57481 DVSS.n4318 DVSS.n4041 1.89035
R57482 DVSS.n4166 DVSS.n4005 1.89035
R57483 DVSS.n4318 DVSS.n4040 1.89035
R57484 DVSS.n4171 DVSS.n4005 1.89035
R57485 DVSS.n4318 DVSS.n4039 1.89035
R57486 DVSS.n4176 DVSS.n4005 1.89035
R57487 DVSS.n4318 DVSS.n4038 1.89035
R57488 DVSS.n4179 DVSS.n4005 1.89035
R57489 DVSS.n4189 DVSS.n4188 1.89035
R57490 DVSS.n4060 DVSS.n4005 1.89035
R57491 DVSS.n4189 DVSS.n4187 1.89035
R57492 DVSS.n4062 DVSS.n4005 1.89035
R57493 DVSS.n4189 DVSS.n4186 1.89035
R57494 DVSS.n4183 DVSS.n4005 1.89035
R57495 DVSS.n4318 DVSS.n4034 1.89035
R57496 DVSS.n4193 DVSS.n4005 1.89035
R57497 DVSS.n4318 DVSS.n4033 1.89035
R57498 DVSS.n4198 DVSS.n4005 1.89035
R57499 DVSS.n4318 DVSS.n4032 1.89035
R57500 DVSS.n4203 DVSS.n4005 1.89035
R57501 DVSS.n4318 DVSS.n4031 1.89035
R57502 DVSS.n4208 DVSS.n4005 1.89035
R57503 DVSS.n4318 DVSS.n4030 1.89035
R57504 DVSS.n4213 DVSS.n4005 1.89035
R57505 DVSS.n4318 DVSS.n4029 1.89035
R57506 DVSS.n4218 DVSS.n4005 1.89035
R57507 DVSS.n4318 DVSS.n4028 1.89035
R57508 DVSS.n4223 DVSS.n4005 1.89035
R57509 DVSS.n4318 DVSS.n4027 1.89035
R57510 DVSS.n4228 DVSS.n4005 1.89035
R57511 DVSS.n4318 DVSS.n4026 1.89035
R57512 DVSS.n4233 DVSS.n4005 1.89035
R57513 DVSS.n4318 DVSS.n4025 1.89035
R57514 DVSS.n4238 DVSS.n4005 1.89035
R57515 DVSS.n4318 DVSS.n4024 1.89035
R57516 DVSS.n4243 DVSS.n4005 1.89035
R57517 DVSS.n4318 DVSS.n4023 1.89035
R57518 DVSS.n4248 DVSS.n4005 1.89035
R57519 DVSS.n4318 DVSS.n4022 1.89035
R57520 DVSS.n4253 DVSS.n4005 1.89035
R57521 DVSS.n4318 DVSS.n4021 1.89035
R57522 DVSS.n4258 DVSS.n4005 1.89035
R57523 DVSS.n4318 DVSS.n4020 1.89035
R57524 DVSS.n4263 DVSS.n4005 1.89035
R57525 DVSS.n4318 DVSS.n4019 1.89035
R57526 DVSS.n4268 DVSS.n4005 1.89035
R57527 DVSS.n4318 DVSS.n4018 1.89035
R57528 DVSS.n4273 DVSS.n4005 1.89035
R57529 DVSS.n4318 DVSS.n4017 1.89035
R57530 DVSS.n4278 DVSS.n4005 1.89035
R57531 DVSS.n4318 DVSS.n4016 1.89035
R57532 DVSS.n4283 DVSS.n4005 1.89035
R57533 DVSS.n4318 DVSS.n4015 1.89035
R57534 DVSS.n4288 DVSS.n4005 1.89035
R57535 DVSS.n4318 DVSS.n4014 1.89035
R57536 DVSS.n4293 DVSS.n4005 1.89035
R57537 DVSS.n4318 DVSS.n4013 1.89035
R57538 DVSS.n4298 DVSS.n4005 1.89035
R57539 DVSS.n4318 DVSS.n4012 1.89035
R57540 DVSS.n4303 DVSS.n4005 1.89035
R57541 DVSS.n4318 DVSS.n4011 1.89035
R57542 DVSS.n4308 DVSS.n4005 1.89035
R57543 DVSS.n4318 DVSS.n4010 1.89035
R57544 DVSS.n4311 DVSS.n4005 1.89035
R57545 DVSS.n4067 DVSS.n4065 1.89035
R57546 DVSS.n5361 DVSS.n1410 1.89035
R57547 DVSS.n1514 DVSS.n1375 1.89035
R57548 DVSS.n5361 DVSS.n1409 1.89035
R57549 DVSS.n1509 DVSS.n1375 1.89035
R57550 DVSS.n5361 DVSS.n1408 1.89035
R57551 DVSS.n1504 DVSS.n1375 1.89035
R57552 DVSS.n5361 DVSS.n1407 1.89035
R57553 DVSS.n1499 DVSS.n1375 1.89035
R57554 DVSS.n5361 DVSS.n1406 1.89035
R57555 DVSS.n1494 DVSS.n1375 1.89035
R57556 DVSS.n5361 DVSS.n1405 1.89035
R57557 DVSS.n1489 DVSS.n1375 1.89035
R57558 DVSS.n5361 DVSS.n1404 1.89035
R57559 DVSS.n1484 DVSS.n1375 1.89035
R57560 DVSS.n5361 DVSS.n1403 1.89035
R57561 DVSS.n1479 DVSS.n1375 1.89035
R57562 DVSS.n5361 DVSS.n1402 1.89035
R57563 DVSS.n1474 DVSS.n1375 1.89035
R57564 DVSS.n5361 DVSS.n1401 1.89035
R57565 DVSS.n1469 DVSS.n1375 1.89035
R57566 DVSS.n5361 DVSS.n1400 1.89035
R57567 DVSS.n1464 DVSS.n1375 1.89035
R57568 DVSS.n5361 DVSS.n1399 1.89035
R57569 DVSS.n1459 DVSS.n1375 1.89035
R57570 DVSS.n5361 DVSS.n1398 1.89035
R57571 DVSS.n1454 DVSS.n1375 1.89035
R57572 DVSS.n5361 DVSS.n1397 1.89035
R57573 DVSS.n1449 DVSS.n1375 1.89035
R57574 DVSS.n5361 DVSS.n1396 1.89035
R57575 DVSS.n1444 DVSS.n1375 1.89035
R57576 DVSS.n5361 DVSS.n1395 1.89035
R57577 DVSS.n1439 DVSS.n1375 1.89035
R57578 DVSS.n5361 DVSS.n1394 1.89035
R57579 DVSS.n1434 DVSS.n1375 1.89035
R57580 DVSS.n5361 DVSS.n1393 1.89035
R57581 DVSS.n1429 DVSS.n1375 1.89035
R57582 DVSS.n5361 DVSS.n1392 1.89035
R57583 DVSS.n1424 DVSS.n1375 1.89035
R57584 DVSS.n5361 DVSS.n1391 1.89035
R57585 DVSS.n1419 DVSS.n1375 1.89035
R57586 DVSS.n5361 DVSS.n1390 1.89035
R57587 DVSS.n1414 DVSS.n1375 1.89035
R57588 DVSS.n5361 DVSS.n1389 1.89035
R57589 DVSS.n5358 DVSS.n5357 1.89035
R57590 DVSS.n5361 DVSS.n1388 1.89035
R57591 DVSS.n5361 DVSS.n5360 1.89035
R57592 DVSS.n5358 DVSS.n1387 1.89035
R57593 DVSS.n5497 DVSS.n5361 1.89035
R57594 DVSS.n5495 DVSS.n1375 1.89035
R57595 DVSS.n5362 DVSS.n5361 1.89035
R57596 DVSS.n5490 DVSS.n1375 1.89035
R57597 DVSS.n5488 DVSS.n5361 1.89035
R57598 DVSS.n5364 DVSS.n1375 1.89035
R57599 DVSS.n5483 DVSS.n5361 1.89035
R57600 DVSS.n5481 DVSS.n1375 1.89035
R57601 DVSS.n5366 DVSS.n5361 1.89035
R57602 DVSS.n5476 DVSS.n1375 1.89035
R57603 DVSS.n5474 DVSS.n5361 1.89035
R57604 DVSS.n5368 DVSS.n1375 1.89035
R57605 DVSS.n5469 DVSS.n5361 1.89035
R57606 DVSS.n5467 DVSS.n1375 1.89035
R57607 DVSS.n5370 DVSS.n5361 1.89035
R57608 DVSS.n5462 DVSS.n1375 1.89035
R57609 DVSS.n5460 DVSS.n5361 1.89035
R57610 DVSS.n5372 DVSS.n1375 1.89035
R57611 DVSS.n5455 DVSS.n5361 1.89035
R57612 DVSS.n5453 DVSS.n1375 1.89035
R57613 DVSS.n5374 DVSS.n5361 1.89035
R57614 DVSS.n5448 DVSS.n1375 1.89035
R57615 DVSS.n5375 DVSS.n5361 1.89035
R57616 DVSS.n5443 DVSS.n1375 1.89035
R57617 DVSS.n5377 DVSS.n5361 1.89035
R57618 DVSS.n5438 DVSS.n1375 1.89035
R57619 DVSS.n5436 DVSS.n5361 1.89035
R57620 DVSS.n5379 DVSS.n1375 1.89035
R57621 DVSS.n5431 DVSS.n5361 1.89035
R57622 DVSS.n5429 DVSS.n1375 1.89035
R57623 DVSS.n5381 DVSS.n5361 1.89035
R57624 DVSS.n5424 DVSS.n1375 1.89035
R57625 DVSS.n5422 DVSS.n5361 1.89035
R57626 DVSS.n5383 DVSS.n1375 1.89035
R57627 DVSS.n5417 DVSS.n5361 1.89035
R57628 DVSS.n5415 DVSS.n1375 1.89035
R57629 DVSS.n5385 DVSS.n5361 1.89035
R57630 DVSS.n5410 DVSS.n1375 1.89035
R57631 DVSS.n5408 DVSS.n5361 1.89035
R57632 DVSS.n5387 DVSS.n1375 1.89035
R57633 DVSS.n5403 DVSS.n5361 1.89035
R57634 DVSS.n5401 DVSS.n1375 1.89035
R57635 DVSS.n5389 DVSS.n5361 1.89035
R57636 DVSS.n5396 DVSS.n1375 1.89035
R57637 DVSS.n5660 DVSS.n5659 1.73753
R57638 DVSS.n1288 DVSS.n1271 1.73383
R57639 DVSS.n1292 DVSS.n1271 1.73383
R57640 DVSS.n1295 DVSS.n1294 1.73383
R57641 DVSS.n1294 DVSS.n1293 1.73383
R57642 DVSS.n2879 DVSS.n2878 1.6025
R57643 DVSS.n3545 DVSS.n3544 1.6025
R57644 DVSS.n5598 DVSS.n215 1.59898
R57645 DVSS.n6431 DVSS.n6430 1.59898
R57646 DVSS.n1308 DVSS.n218 1.59898
R57647 DVSS.n6426 DVSS.n6425 1.59898
R57648 DVSS.n2121 DVSS.n2120 1.5005
R57649 DVSS.n2119 DVSS.n2116 1.5005
R57650 DVSS.n3529 DVSS.n2123 1.5005
R57651 DVSS.n3066 DVSS.n3065 1.44597
R57652 DVSS.n6445 DVSS.n6444 1.44597
R57653 DVSS.n6406 DVSS.n6405 1.44597
R57654 DVSS.n267 DVSS.n261 1.44597
R57655 DVSS.n6390 DVSS.n6384 1.44597
R57656 DVSS.n6378 DVSS.n6375 1.44597
R57657 DVSS.n6495 DVSS.n46 1.44597
R57658 DVSS.n375 DVSS.n369 1.44597
R57659 DVSS.n6288 DVSS.n6286 1.44597
R57660 DVSS.n6281 DVSS.n6275 1.44597
R57661 DVSS.n6270 DVSS.n6264 1.44597
R57662 DVSS.n6247 DVSS.n393 1.44597
R57663 DVSS.n6222 DVSS.n6221 1.44597
R57664 DVSS.n6207 DVSS.n6201 1.44597
R57665 DVSS.n1116 DVSS.n1110 1.44597
R57666 DVSS.n1105 DVSS.n1099 1.44597
R57667 DVSS.n6121 DVSS.n6119 1.44597
R57668 DVSS.n6118 DVSS.n6117 1.44597
R57669 DVSS.n6111 DVSS.n1134 1.44597
R57670 DVSS.n5786 DVSS.n5785 1.44597
R57671 DVSS.n6058 DVSS.n6057 1.44597
R57672 DVSS.n6066 DVSS.n6062 1.44597
R57673 DVSS.n5773 DVSS.n5772 1.44597
R57674 DVSS.n5766 DVSS.n1199 1.44597
R57675 DVSS.n1211 DVSS.n1209 1.44597
R57676 DVSS.n5752 DVSS.n5751 1.44597
R57677 DVSS.n5746 DVSS.n1208 1.44597
R57678 DVSS.n1224 DVSS.n1222 1.44597
R57679 DVSS.n5735 DVSS.n5734 1.44597
R57680 DVSS.n5729 DVSS.n1221 1.44597
R57681 DVSS.n5692 DVSS.n5690 1.44597
R57682 DVSS.n1244 DVSS.n1240 1.44597
R57683 DVSS.n5708 DVSS.n5707 1.44597
R57684 DVSS.n5642 DVSS.n1239 1.44597
R57685 DVSS.n5637 DVSS.n5634 1.44597
R57686 DVSS.n5633 DVSS.n5632 1.44597
R57687 DVSS.n5626 DVSS.n1324 1.44597
R57688 DVSS.n5620 DVSS.n5617 1.44597
R57689 DVSS.n5616 DVSS.n5615 1.44597
R57690 DVSS.n5609 DVSS.n1328 1.44597
R57691 DVSS.n5603 DVSS.n5600 1.44597
R57692 DVSS.n6429 DVSS.n215 1.43659
R57693 DVSS.n6430 DVSS.n6429 1.43659
R57694 DVSS.n6427 DVSS.n218 1.43659
R57695 DVSS.n6427 DVSS.n6426 1.43659
R57696 DVSS.n5360 DVSS.n1382 1.42229
R57697 DVSS.n5498 DVSS.n1387 1.42229
R57698 DVSS.n5497 DVSS.n5496 1.42229
R57699 DVSS.n5496 DVSS.n5495 1.42229
R57700 DVSS.n5491 DVSS.n5362 1.42229
R57701 DVSS.n5491 DVSS.n5490 1.42229
R57702 DVSS.n5488 DVSS.n5487 1.42229
R57703 DVSS.n5487 DVSS.n5364 1.42229
R57704 DVSS.n5483 DVSS.n5482 1.42229
R57705 DVSS.n5482 DVSS.n5481 1.42229
R57706 DVSS.n5477 DVSS.n5366 1.42229
R57707 DVSS.n5477 DVSS.n5476 1.42229
R57708 DVSS.n5474 DVSS.n5473 1.42229
R57709 DVSS.n5473 DVSS.n5368 1.42229
R57710 DVSS.n5469 DVSS.n5468 1.42229
R57711 DVSS.n5468 DVSS.n5467 1.42229
R57712 DVSS.n5463 DVSS.n5370 1.42229
R57713 DVSS.n5463 DVSS.n5462 1.42229
R57714 DVSS.n5460 DVSS.n5459 1.42229
R57715 DVSS.n5459 DVSS.n5372 1.42229
R57716 DVSS.n5455 DVSS.n5454 1.42229
R57717 DVSS.n5454 DVSS.n5453 1.42229
R57718 DVSS.n5449 DVSS.n5374 1.42229
R57719 DVSS.n5449 DVSS.n5448 1.42229
R57720 DVSS.n5444 DVSS.n5375 1.42229
R57721 DVSS.n5444 DVSS.n5443 1.42229
R57722 DVSS.n5439 DVSS.n5377 1.42229
R57723 DVSS.n5439 DVSS.n5438 1.42229
R57724 DVSS.n5436 DVSS.n5435 1.42229
R57725 DVSS.n5435 DVSS.n5379 1.42229
R57726 DVSS.n5431 DVSS.n5430 1.42229
R57727 DVSS.n5430 DVSS.n5429 1.42229
R57728 DVSS.n5425 DVSS.n5381 1.42229
R57729 DVSS.n5425 DVSS.n5424 1.42229
R57730 DVSS.n5422 DVSS.n5421 1.42229
R57731 DVSS.n5421 DVSS.n5383 1.42229
R57732 DVSS.n5417 DVSS.n5416 1.42229
R57733 DVSS.n5416 DVSS.n5415 1.42229
R57734 DVSS.n5411 DVSS.n5385 1.42229
R57735 DVSS.n5411 DVSS.n5410 1.42229
R57736 DVSS.n5408 DVSS.n5407 1.42229
R57737 DVSS.n5407 DVSS.n5387 1.42229
R57738 DVSS.n5403 DVSS.n5402 1.42229
R57739 DVSS.n5402 DVSS.n5401 1.42229
R57740 DVSS.n5397 DVSS.n5389 1.42229
R57741 DVSS.n5397 DVSS.n5396 1.42229
R57742 DVSS.n1515 DVSS.n1410 1.42229
R57743 DVSS.n1515 DVSS.n1514 1.42229
R57744 DVSS.n1510 DVSS.n1409 1.42229
R57745 DVSS.n1510 DVSS.n1509 1.42229
R57746 DVSS.n1505 DVSS.n1408 1.42229
R57747 DVSS.n1505 DVSS.n1504 1.42229
R57748 DVSS.n1500 DVSS.n1407 1.42229
R57749 DVSS.n1500 DVSS.n1499 1.42229
R57750 DVSS.n1495 DVSS.n1406 1.42229
R57751 DVSS.n1495 DVSS.n1494 1.42229
R57752 DVSS.n1490 DVSS.n1405 1.42229
R57753 DVSS.n1490 DVSS.n1489 1.42229
R57754 DVSS.n1485 DVSS.n1404 1.42229
R57755 DVSS.n1485 DVSS.n1484 1.42229
R57756 DVSS.n1480 DVSS.n1403 1.42229
R57757 DVSS.n1480 DVSS.n1479 1.42229
R57758 DVSS.n1475 DVSS.n1402 1.42229
R57759 DVSS.n1475 DVSS.n1474 1.42229
R57760 DVSS.n1470 DVSS.n1401 1.42229
R57761 DVSS.n1470 DVSS.n1469 1.42229
R57762 DVSS.n1465 DVSS.n1400 1.42229
R57763 DVSS.n1465 DVSS.n1464 1.42229
R57764 DVSS.n1460 DVSS.n1399 1.42229
R57765 DVSS.n1460 DVSS.n1459 1.42229
R57766 DVSS.n1455 DVSS.n1398 1.42229
R57767 DVSS.n1455 DVSS.n1454 1.42229
R57768 DVSS.n1450 DVSS.n1397 1.42229
R57769 DVSS.n1450 DVSS.n1449 1.42229
R57770 DVSS.n1445 DVSS.n1396 1.42229
R57771 DVSS.n1445 DVSS.n1444 1.42229
R57772 DVSS.n1440 DVSS.n1395 1.42229
R57773 DVSS.n1440 DVSS.n1439 1.42229
R57774 DVSS.n1435 DVSS.n1394 1.42229
R57775 DVSS.n1435 DVSS.n1434 1.42229
R57776 DVSS.n1430 DVSS.n1393 1.42229
R57777 DVSS.n1430 DVSS.n1429 1.42229
R57778 DVSS.n1425 DVSS.n1392 1.42229
R57779 DVSS.n1425 DVSS.n1424 1.42229
R57780 DVSS.n1420 DVSS.n1391 1.42229
R57781 DVSS.n1420 DVSS.n1419 1.42229
R57782 DVSS.n1415 DVSS.n1390 1.42229
R57783 DVSS.n1415 DVSS.n1414 1.42229
R57784 DVSS.n1389 DVSS.n1384 1.42229
R57785 DVSS.n5357 DVSS.n1383 1.42229
R57786 DVSS.n5355 DVSS.n1388 1.42229
R57787 DVSS.n4328 DVSS.n4004 1.42229
R57788 DVSS.n4326 DVSS.n4325 1.42229
R57789 DVSS.n4325 DVSS.n4006 1.42229
R57790 DVSS.n4321 DVSS.n4320 1.42229
R57791 DVSS.n4320 DVSS.n4319 1.42229
R57792 DVSS.n4071 DVSS.n4070 1.42229
R57793 DVSS.n4071 DVSS.n4059 1.42229
R57794 DVSS.n4076 DVSS.n4075 1.42229
R57795 DVSS.n4076 DVSS.n4058 1.42229
R57796 DVSS.n4081 DVSS.n4080 1.42229
R57797 DVSS.n4081 DVSS.n4057 1.42229
R57798 DVSS.n4086 DVSS.n4085 1.42229
R57799 DVSS.n4086 DVSS.n4056 1.42229
R57800 DVSS.n4091 DVSS.n4090 1.42229
R57801 DVSS.n4091 DVSS.n4055 1.42229
R57802 DVSS.n4096 DVSS.n4095 1.42229
R57803 DVSS.n4096 DVSS.n4054 1.42229
R57804 DVSS.n4101 DVSS.n4100 1.42229
R57805 DVSS.n4101 DVSS.n4053 1.42229
R57806 DVSS.n4106 DVSS.n4105 1.42229
R57807 DVSS.n4106 DVSS.n4052 1.42229
R57808 DVSS.n4111 DVSS.n4110 1.42229
R57809 DVSS.n4111 DVSS.n4051 1.42229
R57810 DVSS.n4116 DVSS.n4115 1.42229
R57811 DVSS.n4116 DVSS.n4050 1.42229
R57812 DVSS.n4121 DVSS.n4120 1.42229
R57813 DVSS.n4121 DVSS.n4049 1.42229
R57814 DVSS.n4127 DVSS.n4126 1.42229
R57815 DVSS.n4127 DVSS.n4048 1.42229
R57816 DVSS.n4132 DVSS.n4131 1.42229
R57817 DVSS.n4132 DVSS.n4047 1.42229
R57818 DVSS.n4137 DVSS.n4136 1.42229
R57819 DVSS.n4137 DVSS.n4046 1.42229
R57820 DVSS.n4142 DVSS.n4141 1.42229
R57821 DVSS.n4142 DVSS.n4045 1.42229
R57822 DVSS.n4147 DVSS.n4146 1.42229
R57823 DVSS.n4147 DVSS.n4044 1.42229
R57824 DVSS.n4152 DVSS.n4151 1.42229
R57825 DVSS.n4152 DVSS.n4043 1.42229
R57826 DVSS.n4157 DVSS.n4156 1.42229
R57827 DVSS.n4157 DVSS.n4042 1.42229
R57828 DVSS.n4162 DVSS.n4161 1.42229
R57829 DVSS.n4162 DVSS.n4041 1.42229
R57830 DVSS.n4167 DVSS.n4166 1.42229
R57831 DVSS.n4167 DVSS.n4040 1.42229
R57832 DVSS.n4172 DVSS.n4171 1.42229
R57833 DVSS.n4172 DVSS.n4039 1.42229
R57834 DVSS.n4177 DVSS.n4176 1.42229
R57835 DVSS.n4177 DVSS.n4038 1.42229
R57836 DVSS.n4179 DVSS.n4037 1.42229
R57837 DVSS.n4188 DVSS.n4061 1.42229
R57838 DVSS.n4060 DVSS.n4036 1.42229
R57839 DVSS.n4187 DVSS.n4063 1.42229
R57840 DVSS.n4062 DVSS.n4035 1.42229
R57841 DVSS.n4186 DVSS.n4064 1.42229
R57842 DVSS.n4184 DVSS.n4183 1.42229
R57843 DVSS.n4184 DVSS.n4034 1.42229
R57844 DVSS.n4194 DVSS.n4193 1.42229
R57845 DVSS.n4194 DVSS.n4033 1.42229
R57846 DVSS.n4199 DVSS.n4198 1.42229
R57847 DVSS.n4199 DVSS.n4032 1.42229
R57848 DVSS.n4204 DVSS.n4203 1.42229
R57849 DVSS.n4204 DVSS.n4031 1.42229
R57850 DVSS.n4209 DVSS.n4208 1.42229
R57851 DVSS.n4209 DVSS.n4030 1.42229
R57852 DVSS.n4214 DVSS.n4213 1.42229
R57853 DVSS.n4214 DVSS.n4029 1.42229
R57854 DVSS.n4219 DVSS.n4218 1.42229
R57855 DVSS.n4219 DVSS.n4028 1.42229
R57856 DVSS.n4224 DVSS.n4223 1.42229
R57857 DVSS.n4224 DVSS.n4027 1.42229
R57858 DVSS.n4229 DVSS.n4228 1.42229
R57859 DVSS.n4229 DVSS.n4026 1.42229
R57860 DVSS.n4234 DVSS.n4233 1.42229
R57861 DVSS.n4234 DVSS.n4025 1.42229
R57862 DVSS.n4239 DVSS.n4238 1.42229
R57863 DVSS.n4239 DVSS.n4024 1.42229
R57864 DVSS.n4244 DVSS.n4243 1.42229
R57865 DVSS.n4244 DVSS.n4023 1.42229
R57866 DVSS.n4249 DVSS.n4248 1.42229
R57867 DVSS.n4249 DVSS.n4022 1.42229
R57868 DVSS.n4254 DVSS.n4253 1.42229
R57869 DVSS.n4254 DVSS.n4021 1.42229
R57870 DVSS.n4259 DVSS.n4258 1.42229
R57871 DVSS.n4259 DVSS.n4020 1.42229
R57872 DVSS.n4264 DVSS.n4263 1.42229
R57873 DVSS.n4264 DVSS.n4019 1.42229
R57874 DVSS.n4269 DVSS.n4268 1.42229
R57875 DVSS.n4269 DVSS.n4018 1.42229
R57876 DVSS.n4274 DVSS.n4273 1.42229
R57877 DVSS.n4274 DVSS.n4017 1.42229
R57878 DVSS.n4279 DVSS.n4278 1.42229
R57879 DVSS.n4279 DVSS.n4016 1.42229
R57880 DVSS.n4284 DVSS.n4283 1.42229
R57881 DVSS.n4284 DVSS.n4015 1.42229
R57882 DVSS.n4289 DVSS.n4288 1.42229
R57883 DVSS.n4289 DVSS.n4014 1.42229
R57884 DVSS.n4294 DVSS.n4293 1.42229
R57885 DVSS.n4294 DVSS.n4013 1.42229
R57886 DVSS.n4299 DVSS.n4298 1.42229
R57887 DVSS.n4299 DVSS.n4012 1.42229
R57888 DVSS.n4304 DVSS.n4303 1.42229
R57889 DVSS.n4304 DVSS.n4011 1.42229
R57890 DVSS.n4309 DVSS.n4308 1.42229
R57891 DVSS.n4309 DVSS.n4010 1.42229
R57892 DVSS.n4311 DVSS.n4009 1.42229
R57893 DVSS.n4316 DVSS.n4065 1.42229
R57894 DVSS.n4004 DVSS.n4003 1.42229
R57895 DVSS.n4328 DVSS.n4326 1.42229
R57896 DVSS.n4322 DVSS.n4321 1.42229
R57897 DVSS.n4322 DVSS.n4006 1.42229
R57898 DVSS.n4070 DVSS.n4008 1.42229
R57899 DVSS.n4319 DVSS.n4008 1.42229
R57900 DVSS.n4075 DVSS.n4074 1.42229
R57901 DVSS.n4074 DVSS.n4059 1.42229
R57902 DVSS.n4080 DVSS.n4079 1.42229
R57903 DVSS.n4079 DVSS.n4058 1.42229
R57904 DVSS.n4085 DVSS.n4084 1.42229
R57905 DVSS.n4084 DVSS.n4057 1.42229
R57906 DVSS.n4090 DVSS.n4089 1.42229
R57907 DVSS.n4089 DVSS.n4056 1.42229
R57908 DVSS.n4095 DVSS.n4094 1.42229
R57909 DVSS.n4094 DVSS.n4055 1.42229
R57910 DVSS.n4100 DVSS.n4099 1.42229
R57911 DVSS.n4099 DVSS.n4054 1.42229
R57912 DVSS.n4105 DVSS.n4104 1.42229
R57913 DVSS.n4104 DVSS.n4053 1.42229
R57914 DVSS.n4110 DVSS.n4109 1.42229
R57915 DVSS.n4109 DVSS.n4052 1.42229
R57916 DVSS.n4115 DVSS.n4114 1.42229
R57917 DVSS.n4114 DVSS.n4051 1.42229
R57918 DVSS.n4120 DVSS.n4119 1.42229
R57919 DVSS.n4119 DVSS.n4050 1.42229
R57920 DVSS.n4126 DVSS.n4125 1.42229
R57921 DVSS.n4125 DVSS.n4049 1.42229
R57922 DVSS.n4131 DVSS.n4130 1.42229
R57923 DVSS.n4130 DVSS.n4048 1.42229
R57924 DVSS.n4136 DVSS.n4135 1.42229
R57925 DVSS.n4135 DVSS.n4047 1.42229
R57926 DVSS.n4141 DVSS.n4140 1.42229
R57927 DVSS.n4140 DVSS.n4046 1.42229
R57928 DVSS.n4146 DVSS.n4145 1.42229
R57929 DVSS.n4145 DVSS.n4045 1.42229
R57930 DVSS.n4151 DVSS.n4150 1.42229
R57931 DVSS.n4150 DVSS.n4044 1.42229
R57932 DVSS.n4156 DVSS.n4155 1.42229
R57933 DVSS.n4155 DVSS.n4043 1.42229
R57934 DVSS.n4161 DVSS.n4160 1.42229
R57935 DVSS.n4160 DVSS.n4042 1.42229
R57936 DVSS.n4166 DVSS.n4165 1.42229
R57937 DVSS.n4165 DVSS.n4041 1.42229
R57938 DVSS.n4171 DVSS.n4170 1.42229
R57939 DVSS.n4170 DVSS.n4040 1.42229
R57940 DVSS.n4176 DVSS.n4175 1.42229
R57941 DVSS.n4175 DVSS.n4039 1.42229
R57942 DVSS.n4180 DVSS.n4179 1.42229
R57943 DVSS.n4180 DVSS.n4038 1.42229
R57944 DVSS.n4188 DVSS.n4037 1.42229
R57945 DVSS.n4061 DVSS.n4060 1.42229
R57946 DVSS.n4187 DVSS.n4036 1.42229
R57947 DVSS.n4063 DVSS.n4062 1.42229
R57948 DVSS.n4186 DVSS.n4035 1.42229
R57949 DVSS.n4183 DVSS.n4064 1.42229
R57950 DVSS.n4193 DVSS.n4192 1.42229
R57951 DVSS.n4192 DVSS.n4034 1.42229
R57952 DVSS.n4198 DVSS.n4197 1.42229
R57953 DVSS.n4197 DVSS.n4033 1.42229
R57954 DVSS.n4203 DVSS.n4202 1.42229
R57955 DVSS.n4202 DVSS.n4032 1.42229
R57956 DVSS.n4208 DVSS.n4207 1.42229
R57957 DVSS.n4207 DVSS.n4031 1.42229
R57958 DVSS.n4213 DVSS.n4212 1.42229
R57959 DVSS.n4212 DVSS.n4030 1.42229
R57960 DVSS.n4218 DVSS.n4217 1.42229
R57961 DVSS.n4217 DVSS.n4029 1.42229
R57962 DVSS.n4223 DVSS.n4222 1.42229
R57963 DVSS.n4222 DVSS.n4028 1.42229
R57964 DVSS.n4228 DVSS.n4227 1.42229
R57965 DVSS.n4227 DVSS.n4027 1.42229
R57966 DVSS.n4233 DVSS.n4232 1.42229
R57967 DVSS.n4232 DVSS.n4026 1.42229
R57968 DVSS.n4238 DVSS.n4237 1.42229
R57969 DVSS.n4237 DVSS.n4025 1.42229
R57970 DVSS.n4243 DVSS.n4242 1.42229
R57971 DVSS.n4242 DVSS.n4024 1.42229
R57972 DVSS.n4248 DVSS.n4247 1.42229
R57973 DVSS.n4247 DVSS.n4023 1.42229
R57974 DVSS.n4253 DVSS.n4252 1.42229
R57975 DVSS.n4252 DVSS.n4022 1.42229
R57976 DVSS.n4258 DVSS.n4257 1.42229
R57977 DVSS.n4257 DVSS.n4021 1.42229
R57978 DVSS.n4263 DVSS.n4262 1.42229
R57979 DVSS.n4262 DVSS.n4020 1.42229
R57980 DVSS.n4268 DVSS.n4267 1.42229
R57981 DVSS.n4267 DVSS.n4019 1.42229
R57982 DVSS.n4273 DVSS.n4272 1.42229
R57983 DVSS.n4272 DVSS.n4018 1.42229
R57984 DVSS.n4278 DVSS.n4277 1.42229
R57985 DVSS.n4277 DVSS.n4017 1.42229
R57986 DVSS.n4283 DVSS.n4282 1.42229
R57987 DVSS.n4282 DVSS.n4016 1.42229
R57988 DVSS.n4288 DVSS.n4287 1.42229
R57989 DVSS.n4287 DVSS.n4015 1.42229
R57990 DVSS.n4293 DVSS.n4292 1.42229
R57991 DVSS.n4292 DVSS.n4014 1.42229
R57992 DVSS.n4298 DVSS.n4297 1.42229
R57993 DVSS.n4297 DVSS.n4013 1.42229
R57994 DVSS.n4303 DVSS.n4302 1.42229
R57995 DVSS.n4302 DVSS.n4012 1.42229
R57996 DVSS.n4308 DVSS.n4307 1.42229
R57997 DVSS.n4307 DVSS.n4011 1.42229
R57998 DVSS.n4312 DVSS.n4311 1.42229
R57999 DVSS.n4312 DVSS.n4010 1.42229
R58000 DVSS.n4065 DVSS.n4009 1.42229
R58001 DVSS.n1411 DVSS.n1410 1.42229
R58002 DVSS.n1513 DVSS.n1409 1.42229
R58003 DVSS.n1514 DVSS.n1513 1.42229
R58004 DVSS.n1508 DVSS.n1408 1.42229
R58005 DVSS.n1509 DVSS.n1508 1.42229
R58006 DVSS.n1503 DVSS.n1407 1.42229
R58007 DVSS.n1504 DVSS.n1503 1.42229
R58008 DVSS.n1498 DVSS.n1406 1.42229
R58009 DVSS.n1499 DVSS.n1498 1.42229
R58010 DVSS.n1493 DVSS.n1405 1.42229
R58011 DVSS.n1494 DVSS.n1493 1.42229
R58012 DVSS.n1488 DVSS.n1404 1.42229
R58013 DVSS.n1489 DVSS.n1488 1.42229
R58014 DVSS.n1483 DVSS.n1403 1.42229
R58015 DVSS.n1484 DVSS.n1483 1.42229
R58016 DVSS.n1478 DVSS.n1402 1.42229
R58017 DVSS.n1479 DVSS.n1478 1.42229
R58018 DVSS.n1473 DVSS.n1401 1.42229
R58019 DVSS.n1474 DVSS.n1473 1.42229
R58020 DVSS.n1468 DVSS.n1400 1.42229
R58021 DVSS.n1469 DVSS.n1468 1.42229
R58022 DVSS.n1463 DVSS.n1399 1.42229
R58023 DVSS.n1464 DVSS.n1463 1.42229
R58024 DVSS.n1458 DVSS.n1398 1.42229
R58025 DVSS.n1459 DVSS.n1458 1.42229
R58026 DVSS.n1453 DVSS.n1397 1.42229
R58027 DVSS.n1454 DVSS.n1453 1.42229
R58028 DVSS.n1448 DVSS.n1396 1.42229
R58029 DVSS.n1449 DVSS.n1448 1.42229
R58030 DVSS.n1443 DVSS.n1395 1.42229
R58031 DVSS.n1444 DVSS.n1443 1.42229
R58032 DVSS.n1438 DVSS.n1394 1.42229
R58033 DVSS.n1439 DVSS.n1438 1.42229
R58034 DVSS.n1433 DVSS.n1393 1.42229
R58035 DVSS.n1434 DVSS.n1433 1.42229
R58036 DVSS.n1428 DVSS.n1392 1.42229
R58037 DVSS.n1429 DVSS.n1428 1.42229
R58038 DVSS.n1423 DVSS.n1391 1.42229
R58039 DVSS.n1424 DVSS.n1423 1.42229
R58040 DVSS.n1418 DVSS.n1390 1.42229
R58041 DVSS.n1419 DVSS.n1418 1.42229
R58042 DVSS.n1413 DVSS.n1389 1.42229
R58043 DVSS.n1414 DVSS.n1413 1.42229
R58044 DVSS.n5357 DVSS.n1384 1.42229
R58045 DVSS.n1388 DVSS.n1383 1.42229
R58046 DVSS.n5360 DVSS.n1386 1.42229
R58047 DVSS.n1387 DVSS.n1382 1.42229
R58048 DVSS.n5498 DVSS.n5497 1.42229
R58049 DVSS.n5494 DVSS.n5362 1.42229
R58050 DVSS.n5495 DVSS.n5494 1.42229
R58051 DVSS.n5489 DVSS.n5488 1.42229
R58052 DVSS.n5490 DVSS.n5489 1.42229
R58053 DVSS.n5484 DVSS.n5483 1.42229
R58054 DVSS.n5484 DVSS.n5364 1.42229
R58055 DVSS.n5480 DVSS.n5366 1.42229
R58056 DVSS.n5481 DVSS.n5480 1.42229
R58057 DVSS.n5475 DVSS.n5474 1.42229
R58058 DVSS.n5476 DVSS.n5475 1.42229
R58059 DVSS.n5470 DVSS.n5469 1.42229
R58060 DVSS.n5470 DVSS.n5368 1.42229
R58061 DVSS.n5466 DVSS.n5370 1.42229
R58062 DVSS.n5467 DVSS.n5466 1.42229
R58063 DVSS.n5461 DVSS.n5460 1.42229
R58064 DVSS.n5462 DVSS.n5461 1.42229
R58065 DVSS.n5456 DVSS.n5455 1.42229
R58066 DVSS.n5456 DVSS.n5372 1.42229
R58067 DVSS.n5452 DVSS.n5374 1.42229
R58068 DVSS.n5453 DVSS.n5452 1.42229
R58069 DVSS.n5447 DVSS.n5375 1.42229
R58070 DVSS.n5448 DVSS.n5447 1.42229
R58071 DVSS.n5442 DVSS.n5377 1.42229
R58072 DVSS.n5443 DVSS.n5442 1.42229
R58073 DVSS.n5437 DVSS.n5436 1.42229
R58074 DVSS.n5438 DVSS.n5437 1.42229
R58075 DVSS.n5432 DVSS.n5431 1.42229
R58076 DVSS.n5432 DVSS.n5379 1.42229
R58077 DVSS.n5428 DVSS.n5381 1.42229
R58078 DVSS.n5429 DVSS.n5428 1.42229
R58079 DVSS.n5423 DVSS.n5422 1.42229
R58080 DVSS.n5424 DVSS.n5423 1.42229
R58081 DVSS.n5418 DVSS.n5417 1.42229
R58082 DVSS.n5418 DVSS.n5383 1.42229
R58083 DVSS.n5414 DVSS.n5385 1.42229
R58084 DVSS.n5415 DVSS.n5414 1.42229
R58085 DVSS.n5409 DVSS.n5408 1.42229
R58086 DVSS.n5410 DVSS.n5409 1.42229
R58087 DVSS.n5404 DVSS.n5403 1.42229
R58088 DVSS.n5404 DVSS.n5387 1.42229
R58089 DVSS.n5400 DVSS.n5389 1.42229
R58090 DVSS.n5401 DVSS.n5400 1.42229
R58091 DVSS.n5396 DVSS.n5395 1.42229
R58092 DVSS.n4958 DVSS.n1780 1.35477
R58093 DVSS.n4959 DVSS.n1764 1.35477
R58094 DVSS.n5507 DVSS.n1369 1.3307
R58095 DVSS.n5262 DVSS.n5261 1.3307
R58096 DVSS.n4641 DVSS.n4640 1.3307
R58097 DVSS.n3954 DVSS.n2057 1.3307
R58098 DVSS.n5594 DVSS.n1272 1.32884
R58099 DVSS.n5661 DVSS.n5660 1.32884
R58100 DVSS.n3511 DVSS.n3510 1.29118
R58101 DVSS.n3508 DVSS.n3507 1.29118
R58102 DVSS.n5658 DVSS.n1297 1.19767
R58103 DVSS.n5349 DVSS.n5348 1.1255
R58104 DVSS.n5507 DVSS.n5506 1.1255
R58105 DVSS.n5169 DVSS.n5168 1.1255
R58106 DVSS.n5261 DVSS.n5260 1.1255
R58107 DVSS.n4913 DVSS.n4912 1.1255
R58108 DVSS.n4641 DVSS.n1813 1.1255
R58109 DVSS.n4332 DVSS.n3885 1.1255
R58110 DVSS.n3955 DVSS.n3954 1.1255
R58111 DVSS.n1518 DVSS.n1517 1.12321
R58112 DVSS.n1517 DVSS.n1411 1.11525
R58113 DVSS.n5720 DVSS.n1234 1.10985
R58114 DVSS.n5688 DVSS.n1246 1.10985
R58115 DVSS.n6082 DVSS.n6081 1.10985
R58116 DVSS.n6078 DVSS.n6077 1.10985
R58117 DVSS.n501 DVSS.n500 1.10985
R58118 DVSS.n507 DVSS.n387 1.10985
R58119 DVSS.n5714 DVSS.n1233 1.10691
R58120 DVSS.n5700 DVSS.n5699 1.10691
R58121 DVSS.n6086 DVSS.n6084 1.10691
R58122 DVSS.n6075 DVSS.n6074 1.10691
R58123 DVSS.n496 DVSS.n495 1.10691
R58124 DVSS.n6257 DVSS.n388 1.10691
R58125 DVSS.n3093 DVSS.n2367 1.06594
R58126 DVSS.n5361 DVSS.n1519 1.03912
R58127 DVSS.n5668 DVSS.n1277 1.00453
R58128 DVSS.n5508 DVSS.n5507 0.9896
R58129 DVSS.n3954 DVSS.n3953 0.9896
R58130 DVSS.n3790 DVSS.n1863 0.954735
R58131 DVSS.n5261 DVSS.n1591 0.95135
R58132 DVSS.n4642 DVSS.n4641 0.95135
R58133 DVSS.n5348 DVSS.n1524 0.9356
R58134 DVSS.n5168 DVSS.n5165 0.9356
R58135 DVSS.n4914 DVSS.n4913 0.9356
R58136 DVSS.n3885 DVSS.n3884 0.9356
R58137 DVSS.n5000 DVSS.n1737 0.928878
R58138 DVSS.n5004 DVSS.n5002 0.928878
R58139 DVSS.n3034 DVSS.n3032 0.928878
R58140 DVSS.n3037 DVSS.n3036 0.928878
R58141 DVSS.n1296 DVSS.t15 0.913226
R58142 DVSS.n1268 DVSS.t11 0.913226
R58143 DVSS.n1269 DVSS.t7 0.913226
R58144 DVSS.n5394 DVSS.n5361 0.903572
R58145 DVSS.n5669 DVSS.n5668 0.902201
R58146 DVSS.n5680 DVSS.n5679 0.9005
R58147 DVSS.n2885 DVSS.n2884 0.88295
R58148 DVSS.n3052 DVSS.n3051 0.88295
R58149 DVSS.n3021 DVSS.n3020 0.88295
R58150 DVSS.n2458 DVSS.n2107 0.88295
R58151 DVSS.n5087 DVSS.n5086 0.8825
R58152 DVSS.n3755 DVSS.n3754 0.8825
R58153 DVSS.n4926 DVSS.n4925 0.8825
R58154 DVSS.n3694 DVSS.n3693 0.8825
R58155 DVSS.n3094 DVSS.n3093 0.825923
R58156 DVSS.n3293 DVSS.n1277 0.800919
R58157 DVSS.n4933 DVSS.n4932 0.791851
R58158 DVSS.n4981 DVSS.n1730 0.791851
R58159 DVSS.n4977 DVSS.n1768 0.791851
R58160 DVSS.n4954 DVSS.n1786 0.791851
R58161 DVSS.n5676 DVSS.n5675 0.786676
R58162 DVSS.n5679 DVSS.n1263 0.785781
R58163 DVSS.n1517 DVSS.n1516 0.764199
R58164 DVSS.n3504 DVSS.n3503 0.763161
R58165 DVSS.n3514 DVSS.n2138 0.763161
R58166 DVSS.n4981 DVSS.n4980 0.743357
R58167 DVSS.n4980 DVSS.n4979 0.743357
R58168 DVSS.n4930 DVSS.n1779 0.743357
R58169 DVSS.n4956 DVSS.n1779 0.743357
R58170 DVSS.n4932 DVSS.n1785 0.743357
R58171 DVSS.n4956 DVSS.n1785 0.743357
R58172 DVSS.n1765 DVSS.n1759 0.743357
R58173 DVSS.n4979 DVSS.n1765 0.743357
R58174 DVSS.n4957 DVSS.n1782 0.743357
R58175 DVSS.n4957 DVSS.n4956 0.743357
R58176 DVSS.n4978 DVSS.n4977 0.743357
R58177 DVSS.n4979 DVSS.n4978 0.743357
R58178 DVSS.n1769 DVSS.n1763 0.743357
R58179 DVSS.n4979 DVSS.n1763 0.743357
R58180 DVSS.n4955 DVSS.n4954 0.743357
R58181 DVSS.n4956 DVSS.n4955 0.743357
R58182 DVSS.n1288 DVSS.n1287 0.691044
R58183 DVSS.n1295 DVSS.n1290 0.691044
R58184 DVSS.n5678 DVSS.n1265 0.691044
R58185 DVSS.n5677 DVSS.n1267 0.691044
R58186 DVSS.n1297 DVSS.n1296 0.690906
R58187 DVSS.n5676 DVSS.n1268 0.690906
R58188 DVSS.n5356 DVSS.n5355 0.686775
R58189 DVSS.n4317 DVSS.n4316 0.685361
R58190 DVSS.n2380 DVSS.n2379 0.66902
R58191 DVSS.n1270 DVSS.n1269 0.641169
R58192 DVSS.n1287 DVSS.n1286 0.585514
R58193 DVSS.n1290 DVSS.n1289 0.585514
R58194 DVSS.n1263 DVSS.n1262 0.585514
R58195 DVSS.n1265 DVSS.n1264 0.585514
R58196 DVSS.n1267 DVSS.n1266 0.585514
R58197 DVSS.n5675 DVSS.n1270 0.564324
R58198 DVSS.n4365 DVSS 0.557375
R58199 DVSS.n4365 DVSS 0.557375
R58200 DVSS.n1966 DVSS 0.557375
R58201 DVSS.n1966 DVSS 0.557375
R58202 DVSS.n4788 DVSS 0.557375
R58203 DVSS.n4788 DVSS 0.557375
R58204 DVSS.n1300 DVSS.n1258 0.555174
R58205 DVSS.n5682 DVSS.n1260 0.555174
R58206 DVSS.n6467 DVSS.n6465 0.555174
R58207 DVSS.n6463 DVSS.n148 0.555174
R58208 DVSS.n1311 DVSS.n1299 0.553707
R58209 DVSS.n5587 DVSS.n1332 0.553707
R58210 DVSS.n6423 DVSS.n138 0.553707
R58211 DVSS.n6435 DVSS.n6433 0.553707
R58212 DVSS.n4949 DVSS.n1792 0.548638
R58213 DVSS.n4966 DVSS.n4965 0.548638
R58214 DVSS.n4945 DVSS.n1754 0.548638
R58215 DVSS.n4986 DVSS.n4985 0.548638
R58216 DVSS.n2414 DVSS.n1787 0.548638
R58217 DVSS.n2422 DVSS.n1770 0.548638
R58218 DVSS.n1295 DVSS.n1288 0.545794
R58219 DVSS.n1297 DVSS.n1295 0.545794
R58220 DVSS.n5678 DVSS.n5677 0.545794
R58221 DVSS.n5677 DVSS.n5676 0.545794
R58222 DVSS.n5596 DVSS.n5595 0.5072
R58223 DVSS.n5592 DVSS.n5591 0.5072
R58224 DVSS.n5657 DVSS.n5656 0.5072
R58225 DVSS.n1309 DVSS.n1285 0.5072
R58226 DVSS.n2905 DVSS.n2904 0.5005
R58227 DVSS.n2908 DVSS.n2903 0.5005
R58228 DVSS.n2909 DVSS.n2902 0.5005
R58229 DVSS.n2910 DVSS.n2901 0.5005
R58230 DVSS.n2900 DVSS.n2898 0.5005
R58231 DVSS.n2914 DVSS.n2897 0.5005
R58232 DVSS.n2915 DVSS.n2896 0.5005
R58233 DVSS.n2916 DVSS.n2895 0.5005
R58234 DVSS.n2894 DVSS.n2892 0.5005
R58235 DVSS.n2920 DVSS.n2891 0.5005
R58236 DVSS.n2921 DVSS.n2890 0.5005
R58237 DVSS.n2922 DVSS.n2889 0.5005
R58238 DVSS.n2888 DVSS.n2598 0.5005
R58239 DVSS.n2456 DVSS.n2455 0.5005
R58240 DVSS.n2476 DVSS.n2475 0.5005
R58241 DVSS.n2477 DVSS.n2454 0.5005
R58242 DVSS.n2479 DVSS.n2478 0.5005
R58243 DVSS.n2452 DVSS.n2451 0.5005
R58244 DVSS.n2484 DVSS.n2483 0.5005
R58245 DVSS.n2485 DVSS.n2450 0.5005
R58246 DVSS.n2487 DVSS.n2486 0.5005
R58247 DVSS.n2448 DVSS.n2447 0.5005
R58248 DVSS.n2492 DVSS.n2491 0.5005
R58249 DVSS.n2493 DVSS.n2446 0.5005
R58250 DVSS.n2495 DVSS.n2494 0.5005
R58251 DVSS.n2444 DVSS.n2443 0.5005
R58252 DVSS.n2500 DVSS.n2499 0.5005
R58253 DVSS.n2501 DVSS.n2442 0.5005
R58254 DVSS.n3011 DVSS.n2502 0.5005
R58255 DVSS.n3010 DVSS.n2503 0.5005
R58256 DVSS.n3009 DVSS.n2504 0.5005
R58257 DVSS.n3008 DVSS.n2505 0.5005
R58258 DVSS.n2508 DVSS.n2506 0.5005
R58259 DVSS.n3004 DVSS.n2509 0.5005
R58260 DVSS.n3003 DVSS.n2510 0.5005
R58261 DVSS.n3002 DVSS.n2511 0.5005
R58262 DVSS.n2514 DVSS.n2512 0.5005
R58263 DVSS.n2998 DVSS.n2515 0.5005
R58264 DVSS.n2997 DVSS.n2516 0.5005
R58265 DVSS.n2996 DVSS.n2517 0.5005
R58266 DVSS.n2520 DVSS.n2518 0.5005
R58267 DVSS.n2992 DVSS.n2521 0.5005
R58268 DVSS.n2991 DVSS.n2522 0.5005
R58269 DVSS.n2990 DVSS.n2523 0.5005
R58270 DVSS.n2526 DVSS.n2524 0.5005
R58271 DVSS.n2986 DVSS.n2527 0.5005
R58272 DVSS.n2985 DVSS.n2528 0.5005
R58273 DVSS.n2549 DVSS.n2529 0.5005
R58274 DVSS.n2979 DVSS.n2550 0.5005
R58275 DVSS.n2978 DVSS.n2551 0.5005
R58276 DVSS.n2977 DVSS.n2552 0.5005
R58277 DVSS.n2555 DVSS.n2553 0.5005
R58278 DVSS.n2973 DVSS.n2556 0.5005
R58279 DVSS.n2972 DVSS.n2557 0.5005
R58280 DVSS.n2971 DVSS.n2558 0.5005
R58281 DVSS.n2561 DVSS.n2559 0.5005
R58282 DVSS.n2967 DVSS.n2562 0.5005
R58283 DVSS.n2966 DVSS.n2563 0.5005
R58284 DVSS.n2965 DVSS.n2564 0.5005
R58285 DVSS.n2567 DVSS.n2565 0.5005
R58286 DVSS.n2961 DVSS.n2568 0.5005
R58287 DVSS.n2960 DVSS.n2569 0.5005
R58288 DVSS.n2959 DVSS.n2570 0.5005
R58289 DVSS.n2956 DVSS.n2571 0.5005
R58290 DVSS.n2955 DVSS.n2572 0.5005
R58291 DVSS.n2953 DVSS.n2573 0.5005
R58292 DVSS.n2576 DVSS.n2574 0.5005
R58293 DVSS.n2949 DVSS.n2577 0.5005
R58294 DVSS.n2948 DVSS.n2578 0.5005
R58295 DVSS.n2947 DVSS.n2579 0.5005
R58296 DVSS.n2582 DVSS.n2580 0.5005
R58297 DVSS.n2943 DVSS.n2583 0.5005
R58298 DVSS.n2942 DVSS.n2584 0.5005
R58299 DVSS.n2941 DVSS.n2585 0.5005
R58300 DVSS.n2588 DVSS.n2586 0.5005
R58301 DVSS.n2937 DVSS.n2589 0.5005
R58302 DVSS.n2936 DVSS.n2590 0.5005
R58303 DVSS.n2935 DVSS.n2591 0.5005
R58304 DVSS.n2594 DVSS.n2592 0.5005
R58305 DVSS.n2931 DVSS.n2595 0.5005
R58306 DVSS.n2930 DVSS.n2596 0.5005
R58307 DVSS.n2929 DVSS.n2597 0.5005
R58308 DVSS.n2908 DVSS.n2907 0.5005
R58309 DVSS.n2909 DVSS.n2899 0.5005
R58310 DVSS.n2911 DVSS.n2910 0.5005
R58311 DVSS.n2912 DVSS.n2898 0.5005
R58312 DVSS.n2914 DVSS.n2913 0.5005
R58313 DVSS.n2915 DVSS.n2893 0.5005
R58314 DVSS.n2917 DVSS.n2916 0.5005
R58315 DVSS.n2918 DVSS.n2892 0.5005
R58316 DVSS.n2920 DVSS.n2919 0.5005
R58317 DVSS.n2921 DVSS.n2887 0.5005
R58318 DVSS.n2923 DVSS.n2922 0.5005
R58319 DVSS.n2924 DVSS.n2598 0.5005
R58320 DVSS.n2463 DVSS.n2457 0.5005
R58321 DVSS.n2473 DVSS.n2456 0.5005
R58322 DVSS.n2475 DVSS.n2474 0.5005
R58323 DVSS.n2454 DVSS.n2453 0.5005
R58324 DVSS.n2480 DVSS.n2479 0.5005
R58325 DVSS.n2481 DVSS.n2452 0.5005
R58326 DVSS.n2483 DVSS.n2482 0.5005
R58327 DVSS.n2450 DVSS.n2449 0.5005
R58328 DVSS.n2488 DVSS.n2487 0.5005
R58329 DVSS.n2489 DVSS.n2448 0.5005
R58330 DVSS.n2491 DVSS.n2490 0.5005
R58331 DVSS.n2446 DVSS.n2445 0.5005
R58332 DVSS.n2496 DVSS.n2495 0.5005
R58333 DVSS.n2497 DVSS.n2444 0.5005
R58334 DVSS.n2499 DVSS.n2498 0.5005
R58335 DVSS.n2442 DVSS.n2441 0.5005
R58336 DVSS.n3012 DVSS.n3011 0.5005
R58337 DVSS.n3010 DVSS.n2435 0.5005
R58338 DVSS.n3009 DVSS.n2436 0.5005
R58339 DVSS.n3008 DVSS.n3007 0.5005
R58340 DVSS.n3006 DVSS.n2506 0.5005
R58341 DVSS.n3005 DVSS.n3004 0.5005
R58342 DVSS.n3003 DVSS.n2507 0.5005
R58343 DVSS.n3002 DVSS.n3001 0.5005
R58344 DVSS.n3000 DVSS.n2512 0.5005
R58345 DVSS.n2999 DVSS.n2998 0.5005
R58346 DVSS.n2997 DVSS.n2513 0.5005
R58347 DVSS.n2996 DVSS.n2995 0.5005
R58348 DVSS.n2994 DVSS.n2518 0.5005
R58349 DVSS.n2993 DVSS.n2992 0.5005
R58350 DVSS.n2991 DVSS.n2519 0.5005
R58351 DVSS.n2990 DVSS.n2989 0.5005
R58352 DVSS.n2988 DVSS.n2524 0.5005
R58353 DVSS.n2987 DVSS.n2986 0.5005
R58354 DVSS.n2985 DVSS.n2984 0.5005
R58355 DVSS.n2547 DVSS.n2529 0.5005
R58356 DVSS.n2980 DVSS.n2979 0.5005
R58357 DVSS.n2978 DVSS.n2548 0.5005
R58358 DVSS.n2977 DVSS.n2976 0.5005
R58359 DVSS.n2975 DVSS.n2553 0.5005
R58360 DVSS.n2974 DVSS.n2973 0.5005
R58361 DVSS.n2972 DVSS.n2554 0.5005
R58362 DVSS.n2971 DVSS.n2970 0.5005
R58363 DVSS.n2969 DVSS.n2559 0.5005
R58364 DVSS.n2968 DVSS.n2967 0.5005
R58365 DVSS.n2966 DVSS.n2560 0.5005
R58366 DVSS.n2965 DVSS.n2964 0.5005
R58367 DVSS.n2963 DVSS.n2565 0.5005
R58368 DVSS.n2962 DVSS.n2961 0.5005
R58369 DVSS.n2960 DVSS.n2566 0.5005
R58370 DVSS.n2959 DVSS.n2958 0.5005
R58371 DVSS.n2957 DVSS.n2956 0.5005
R58372 DVSS.n2955 DVSS.n2954 0.5005
R58373 DVSS.n2953 DVSS.n2952 0.5005
R58374 DVSS.n2951 DVSS.n2574 0.5005
R58375 DVSS.n2950 DVSS.n2949 0.5005
R58376 DVSS.n2948 DVSS.n2575 0.5005
R58377 DVSS.n2947 DVSS.n2946 0.5005
R58378 DVSS.n2945 DVSS.n2580 0.5005
R58379 DVSS.n2944 DVSS.n2943 0.5005
R58380 DVSS.n2942 DVSS.n2581 0.5005
R58381 DVSS.n2941 DVSS.n2940 0.5005
R58382 DVSS.n2939 DVSS.n2586 0.5005
R58383 DVSS.n2938 DVSS.n2937 0.5005
R58384 DVSS.n2936 DVSS.n2587 0.5005
R58385 DVSS.n2935 DVSS.n2934 0.5005
R58386 DVSS.n2933 DVSS.n2592 0.5005
R58387 DVSS.n2932 DVSS.n2931 0.5005
R58388 DVSS.n2930 DVSS.n2593 0.5005
R58389 DVSS.n2929 DVSS.n2928 0.5005
R58390 DVSS.n4747 DVSS.n1971 0.496843
R58391 DVSS.n3502 DVSS.n3501 0.455549
R58392 DVSS.n2248 DVSS.n2244 0.455549
R58393 DVSS.n3096 DVSS.n2365 0.455549
R58394 DVSS.n3298 DVSS.n3294 0.455549
R58395 DVSS.n2847 DVSS.n2846 0.4505
R58396 DVSS.n2849 DVSS.n2848 0.4505
R58397 DVSS.n2844 DVSS.n2843 0.4505
R58398 DVSS.n2854 DVSS.n2853 0.4505
R58399 DVSS.n2855 DVSS.n2842 0.4505
R58400 DVSS.n2857 DVSS.n2856 0.4505
R58401 DVSS.n2840 DVSS.n2839 0.4505
R58402 DVSS.n2862 DVSS.n2861 0.4505
R58403 DVSS.n2863 DVSS.n2837 0.4505
R58404 DVSS.n2865 DVSS.n2864 0.4505
R58405 DVSS.n2838 DVSS.n2835 0.4505
R58406 DVSS.n2869 DVSS.n2834 0.4505
R58407 DVSS.n2871 DVSS.n2870 0.4505
R58408 DVSS.n2681 DVSS.n2679 0.4505
R58409 DVSS.n2684 DVSS.n2683 0.4505
R58410 DVSS.n2685 DVSS.n2678 0.4505
R58411 DVSS.n2687 DVSS.n2686 0.4505
R58412 DVSS.n2676 DVSS.n2675 0.4505
R58413 DVSS.n2692 DVSS.n2691 0.4505
R58414 DVSS.n2693 DVSS.n2674 0.4505
R58415 DVSS.n2695 DVSS.n2694 0.4505
R58416 DVSS.n2672 DVSS.n2671 0.4505
R58417 DVSS.n2700 DVSS.n2699 0.4505
R58418 DVSS.n2701 DVSS.n2670 0.4505
R58419 DVSS.n2703 DVSS.n2702 0.4505
R58420 DVSS.n2668 DVSS.n2667 0.4505
R58421 DVSS.n2709 DVSS.n2708 0.4505
R58422 DVSS.n2710 DVSS.n2666 0.4505
R58423 DVSS.n2712 DVSS.n2711 0.4505
R58424 DVSS.n2713 DVSS.n2665 0.4505
R58425 DVSS.n2715 DVSS.n2714 0.4505
R58426 DVSS.n2716 DVSS.n2664 0.4505
R58427 DVSS.n2718 DVSS.n2717 0.4505
R58428 DVSS.n2662 DVSS.n2661 0.4505
R58429 DVSS.n2723 DVSS.n2722 0.4505
R58430 DVSS.n2724 DVSS.n2660 0.4505
R58431 DVSS.n2726 DVSS.n2725 0.4505
R58432 DVSS.n2658 DVSS.n2657 0.4505
R58433 DVSS.n2731 DVSS.n2730 0.4505
R58434 DVSS.n2732 DVSS.n2656 0.4505
R58435 DVSS.n2734 DVSS.n2733 0.4505
R58436 DVSS.n2654 DVSS.n2653 0.4505
R58437 DVSS.n2739 DVSS.n2738 0.4505
R58438 DVSS.n2740 DVSS.n2652 0.4505
R58439 DVSS.n2742 DVSS.n2741 0.4505
R58440 DVSS.n2650 DVSS.n2649 0.4505
R58441 DVSS.n2768 DVSS.n2767 0.4505
R58442 DVSS.n2769 DVSS.n2648 0.4505
R58443 DVSS.n2771 DVSS.n2770 0.4505
R58444 DVSS.n2646 DVSS.n2645 0.4505
R58445 DVSS.n2776 DVSS.n2775 0.4505
R58446 DVSS.n2777 DVSS.n2644 0.4505
R58447 DVSS.n2779 DVSS.n2778 0.4505
R58448 DVSS.n2642 DVSS.n2641 0.4505
R58449 DVSS.n2784 DVSS.n2783 0.4505
R58450 DVSS.n2785 DVSS.n2640 0.4505
R58451 DVSS.n2787 DVSS.n2786 0.4505
R58452 DVSS.n2638 DVSS.n2637 0.4505
R58453 DVSS.n2792 DVSS.n2791 0.4505
R58454 DVSS.n2793 DVSS.n2636 0.4505
R58455 DVSS.n2795 DVSS.n2794 0.4505
R58456 DVSS.n2634 DVSS.n2633 0.4505
R58457 DVSS.n2801 DVSS.n2800 0.4505
R58458 DVSS.n2802 DVSS.n2632 0.4505
R58459 DVSS.n2804 DVSS.n2803 0.4505
R58460 DVSS.n2805 DVSS.n2631 0.4505
R58461 DVSS.n2808 DVSS.n2807 0.4505
R58462 DVSS.n2809 DVSS.n2630 0.4505
R58463 DVSS.n2811 DVSS.n2810 0.4505
R58464 DVSS.n2628 DVSS.n2627 0.4505
R58465 DVSS.n2816 DVSS.n2815 0.4505
R58466 DVSS.n2817 DVSS.n2626 0.4505
R58467 DVSS.n2819 DVSS.n2818 0.4505
R58468 DVSS.n2624 DVSS.n2623 0.4505
R58469 DVSS.n2824 DVSS.n2823 0.4505
R58470 DVSS.n2825 DVSS.n2622 0.4505
R58471 DVSS.n2827 DVSS.n2826 0.4505
R58472 DVSS.n2620 DVSS.n2619 0.4505
R58473 DVSS.n2832 DVSS.n2831 0.4505
R58474 DVSS.n2833 DVSS.n2617 0.4505
R58475 DVSS.n2874 DVSS.n2873 0.4505
R58476 DVSS.n2872 DVSS.n2618 0.4505
R58477 DVSS.n2850 DVSS.n2849 0.4505
R58478 DVSS.n2851 DVSS.n2844 0.4505
R58479 DVSS.n2853 DVSS.n2852 0.4505
R58480 DVSS.n2842 DVSS.n2841 0.4505
R58481 DVSS.n2858 DVSS.n2857 0.4505
R58482 DVSS.n2859 DVSS.n2840 0.4505
R58483 DVSS.n2861 DVSS.n2860 0.4505
R58484 DVSS.n2837 DVSS.n2836 0.4505
R58485 DVSS.n2866 DVSS.n2865 0.4505
R58486 DVSS.n2867 DVSS.n2835 0.4505
R58487 DVSS.n2869 DVSS.n2868 0.4505
R58488 DVSS.n2870 DVSS.n2611 0.4505
R58489 DVSS.n2680 DVSS.n2098 0.4505
R58490 DVSS.n2681 DVSS.n2103 0.4505
R58491 DVSS.n2683 DVSS.n2682 0.4505
R58492 DVSS.n2678 DVSS.n2677 0.4505
R58493 DVSS.n2688 DVSS.n2687 0.4505
R58494 DVSS.n2689 DVSS.n2676 0.4505
R58495 DVSS.n2691 DVSS.n2690 0.4505
R58496 DVSS.n2674 DVSS.n2673 0.4505
R58497 DVSS.n2696 DVSS.n2695 0.4505
R58498 DVSS.n2697 DVSS.n2672 0.4505
R58499 DVSS.n2699 DVSS.n2698 0.4505
R58500 DVSS.n2670 DVSS.n2669 0.4505
R58501 DVSS.n2704 DVSS.n2703 0.4505
R58502 DVSS.n2705 DVSS.n2668 0.4505
R58503 DVSS.n2708 DVSS.n2707 0.4505
R58504 DVSS.n2706 DVSS.n2666 0.4505
R58505 DVSS.n2712 DVSS.n2433 0.4505
R58506 DVSS.n2713 DVSS.n2425 0.4505
R58507 DVSS.n2714 DVSS.n2429 0.4505
R58508 DVSS.n2664 DVSS.n2663 0.4505
R58509 DVSS.n2719 DVSS.n2718 0.4505
R58510 DVSS.n2720 DVSS.n2662 0.4505
R58511 DVSS.n2722 DVSS.n2721 0.4505
R58512 DVSS.n2660 DVSS.n2659 0.4505
R58513 DVSS.n2727 DVSS.n2726 0.4505
R58514 DVSS.n2728 DVSS.n2658 0.4505
R58515 DVSS.n2730 DVSS.n2729 0.4505
R58516 DVSS.n2656 DVSS.n2655 0.4505
R58517 DVSS.n2735 DVSS.n2734 0.4505
R58518 DVSS.n2736 DVSS.n2654 0.4505
R58519 DVSS.n2738 DVSS.n2737 0.4505
R58520 DVSS.n2652 DVSS.n2651 0.4505
R58521 DVSS.n2743 DVSS.n2742 0.4505
R58522 DVSS.n2744 DVSS.n2650 0.4505
R58523 DVSS.n2767 DVSS.n2766 0.4505
R58524 DVSS.n2761 DVSS.n2648 0.4505
R58525 DVSS.n2772 DVSS.n2771 0.4505
R58526 DVSS.n2773 DVSS.n2646 0.4505
R58527 DVSS.n2775 DVSS.n2774 0.4505
R58528 DVSS.n2644 DVSS.n2643 0.4505
R58529 DVSS.n2780 DVSS.n2779 0.4505
R58530 DVSS.n2781 DVSS.n2642 0.4505
R58531 DVSS.n2783 DVSS.n2782 0.4505
R58532 DVSS.n2640 DVSS.n2639 0.4505
R58533 DVSS.n2788 DVSS.n2787 0.4505
R58534 DVSS.n2789 DVSS.n2638 0.4505
R58535 DVSS.n2791 DVSS.n2790 0.4505
R58536 DVSS.n2636 DVSS.n2635 0.4505
R58537 DVSS.n2796 DVSS.n2795 0.4505
R58538 DVSS.n2797 DVSS.n2634 0.4505
R58539 DVSS.n2800 DVSS.n2799 0.4505
R58540 DVSS.n2798 DVSS.n2632 0.4505
R58541 DVSS.n2804 DVSS.n2402 0.4505
R58542 DVSS.n2805 DVSS.n2404 0.4505
R58543 DVSS.n2807 DVSS.n2806 0.4505
R58544 DVSS.n2630 DVSS.n2629 0.4505
R58545 DVSS.n2812 DVSS.n2811 0.4505
R58546 DVSS.n2813 DVSS.n2628 0.4505
R58547 DVSS.n2815 DVSS.n2814 0.4505
R58548 DVSS.n2626 DVSS.n2625 0.4505
R58549 DVSS.n2820 DVSS.n2819 0.4505
R58550 DVSS.n2821 DVSS.n2624 0.4505
R58551 DVSS.n2823 DVSS.n2822 0.4505
R58552 DVSS.n2622 DVSS.n2621 0.4505
R58553 DVSS.n2828 DVSS.n2827 0.4505
R58554 DVSS.n2829 DVSS.n2620 0.4505
R58555 DVSS.n2831 DVSS.n2830 0.4505
R58556 DVSS.n2617 DVSS.n2616 0.4505
R58557 DVSS.n2875 DVSS.n2874 0.4505
R58558 DVSS.n2618 DVSS.n2609 0.4505
R58559 DVSS.n5057 DVSS.n5056 0.4505
R58560 DVSS.n5059 DVSS.n5058 0.4505
R58561 DVSS.n5054 DVSS.n5053 0.4505
R58562 DVSS.n5064 DVSS.n5063 0.4505
R58563 DVSS.n5065 DVSS.n5052 0.4505
R58564 DVSS.n5067 DVSS.n5066 0.4505
R58565 DVSS.n5050 DVSS.n5049 0.4505
R58566 DVSS.n5072 DVSS.n5071 0.4505
R58567 DVSS.n5073 DVSS.n5048 0.4505
R58568 DVSS.n5075 DVSS.n5074 0.4505
R58569 DVSS.n5045 DVSS.n5044 0.4505
R58570 DVSS.n5080 DVSS.n5079 0.4505
R58571 DVSS.n5081 DVSS.n1698 0.4505
R58572 DVSS.n3690 DVSS.n3689 0.4505
R58573 DVSS.n3688 DVSS.n2092 0.4505
R58574 DVSS.n3687 DVSS.n3686 0.4505
R58575 DVSS.n3549 DVSS.n3548 0.4505
R58576 DVSS.n3682 DVSS.n3681 0.4505
R58577 DVSS.n3680 DVSS.n3551 0.4505
R58578 DVSS.n3679 DVSS.n3678 0.4505
R58579 DVSS.n3553 DVSS.n3552 0.4505
R58580 DVSS.n3674 DVSS.n3673 0.4505
R58581 DVSS.n3672 DVSS.n3555 0.4505
R58582 DVSS.n3671 DVSS.n3670 0.4505
R58583 DVSS.n3557 DVSS.n3556 0.4505
R58584 DVSS.n3666 DVSS.n3665 0.4505
R58585 DVSS.n3664 DVSS.n3559 0.4505
R58586 DVSS.n3663 DVSS.n3662 0.4505
R58587 DVSS.n3659 DVSS.n3560 0.4505
R58588 DVSS.n3658 DVSS.n3656 0.4505
R58589 DVSS.n3655 DVSS.n3561 0.4505
R58590 DVSS.n3654 DVSS.n3653 0.4505
R58591 DVSS.n3563 DVSS.n3562 0.4505
R58592 DVSS.n3649 DVSS.n3648 0.4505
R58593 DVSS.n3647 DVSS.n3566 0.4505
R58594 DVSS.n3646 DVSS.n3645 0.4505
R58595 DVSS.n3568 DVSS.n3567 0.4505
R58596 DVSS.n3641 DVSS.n3640 0.4505
R58597 DVSS.n3639 DVSS.n3570 0.4505
R58598 DVSS.n3638 DVSS.n3637 0.4505
R58599 DVSS.n3572 DVSS.n3571 0.4505
R58600 DVSS.n3633 DVSS.n3632 0.4505
R58601 DVSS.n3631 DVSS.n3574 0.4505
R58602 DVSS.n3630 DVSS.n3629 0.4505
R58603 DVSS.n3576 DVSS.n3575 0.4505
R58604 DVSS.n3625 DVSS.n3624 0.4505
R58605 DVSS.n3623 DVSS.n3578 0.4505
R58606 DVSS.n3622 DVSS.n3621 0.4505
R58607 DVSS.n3620 DVSS.n3579 0.4505
R58608 DVSS.n3583 DVSS.n3580 0.4505
R58609 DVSS.n3616 DVSS.n3615 0.4505
R58610 DVSS.n3614 DVSS.n3582 0.4505
R58611 DVSS.n3613 DVSS.n3612 0.4505
R58612 DVSS.n3585 DVSS.n3584 0.4505
R58613 DVSS.n3608 DVSS.n3607 0.4505
R58614 DVSS.n3606 DVSS.n3587 0.4505
R58615 DVSS.n3605 DVSS.n3604 0.4505
R58616 DVSS.n3589 DVSS.n3588 0.4505
R58617 DVSS.n3600 DVSS.n3599 0.4505
R58618 DVSS.n3598 DVSS.n3591 0.4505
R58619 DVSS.n3597 DVSS.n3596 0.4505
R58620 DVSS.n3593 DVSS.n3592 0.4505
R58621 DVSS.n1716 DVSS.n1715 0.4505
R58622 DVSS.n5010 DVSS.n5009 0.4505
R58623 DVSS.n5011 DVSS.n1714 0.4505
R58624 DVSS.n5013 DVSS.n5012 0.4505
R58625 DVSS.n1712 DVSS.n1711 0.4505
R58626 DVSS.n5018 DVSS.n5017 0.4505
R58627 DVSS.n5019 DVSS.n1710 0.4505
R58628 DVSS.n5021 DVSS.n5020 0.4505
R58629 DVSS.n1708 DVSS.n1707 0.4505
R58630 DVSS.n5026 DVSS.n5025 0.4505
R58631 DVSS.n5027 DVSS.n1706 0.4505
R58632 DVSS.n5029 DVSS.n5028 0.4505
R58633 DVSS.n1704 DVSS.n1703 0.4505
R58634 DVSS.n5034 DVSS.n5033 0.4505
R58635 DVSS.n5035 DVSS.n1702 0.4505
R58636 DVSS.n5037 DVSS.n5036 0.4505
R58637 DVSS.n1700 DVSS.n1699 0.4505
R58638 DVSS.n5042 DVSS.n5041 0.4505
R58639 DVSS.n5043 DVSS.n1697 0.4505
R58640 DVSS.n5083 DVSS.n5082 0.4505
R58641 DVSS.n5060 DVSS.n5059 0.4505
R58642 DVSS.n5061 DVSS.n5054 0.4505
R58643 DVSS.n5063 DVSS.n5062 0.4505
R58644 DVSS.n5052 DVSS.n5051 0.4505
R58645 DVSS.n5068 DVSS.n5067 0.4505
R58646 DVSS.n5069 DVSS.n5050 0.4505
R58647 DVSS.n5071 DVSS.n5070 0.4505
R58648 DVSS.n5048 DVSS.n5047 0.4505
R58649 DVSS.n5076 DVSS.n5075 0.4505
R58650 DVSS.n5077 DVSS.n5045 0.4505
R58651 DVSS.n5079 DVSS.n5078 0.4505
R58652 DVSS.n5046 DVSS.n1698 0.4505
R58653 DVSS.n2091 DVSS.n2084 0.4505
R58654 DVSS.n3691 DVSS.n3690 0.4505
R58655 DVSS.n2092 DVSS.n2090 0.4505
R58656 DVSS.n3686 DVSS.n3685 0.4505
R58657 DVSS.n3684 DVSS.n3549 0.4505
R58658 DVSS.n3683 DVSS.n3682 0.4505
R58659 DVSS.n3551 DVSS.n3550 0.4505
R58660 DVSS.n3678 DVSS.n3677 0.4505
R58661 DVSS.n3676 DVSS.n3553 0.4505
R58662 DVSS.n3675 DVSS.n3674 0.4505
R58663 DVSS.n3555 DVSS.n3554 0.4505
R58664 DVSS.n3670 DVSS.n3669 0.4505
R58665 DVSS.n3668 DVSS.n3557 0.4505
R58666 DVSS.n3667 DVSS.n3666 0.4505
R58667 DVSS.n3559 DVSS.n3558 0.4505
R58668 DVSS.n3662 DVSS.n3661 0.4505
R58669 DVSS.n3660 DVSS.n3659 0.4505
R58670 DVSS.n3658 DVSS.n3657 0.4505
R58671 DVSS.n3564 DVSS.n3561 0.4505
R58672 DVSS.n3653 DVSS.n3652 0.4505
R58673 DVSS.n3651 DVSS.n3563 0.4505
R58674 DVSS.n3650 DVSS.n3649 0.4505
R58675 DVSS.n3566 DVSS.n3565 0.4505
R58676 DVSS.n3645 DVSS.n3644 0.4505
R58677 DVSS.n3643 DVSS.n3568 0.4505
R58678 DVSS.n3642 DVSS.n3641 0.4505
R58679 DVSS.n3570 DVSS.n3569 0.4505
R58680 DVSS.n3637 DVSS.n3636 0.4505
R58681 DVSS.n3635 DVSS.n3572 0.4505
R58682 DVSS.n3634 DVSS.n3633 0.4505
R58683 DVSS.n3574 DVSS.n3573 0.4505
R58684 DVSS.n3629 DVSS.n3628 0.4505
R58685 DVSS.n3627 DVSS.n3576 0.4505
R58686 DVSS.n3626 DVSS.n3625 0.4505
R58687 DVSS.n3578 DVSS.n3577 0.4505
R58688 DVSS.n3621 DVSS.n1743 0.4505
R58689 DVSS.n3620 DVSS.n3619 0.4505
R58690 DVSS.n3618 DVSS.n3580 0.4505
R58691 DVSS.n3617 DVSS.n3616 0.4505
R58692 DVSS.n3582 DVSS.n3581 0.4505
R58693 DVSS.n3612 DVSS.n3611 0.4505
R58694 DVSS.n3610 DVSS.n3585 0.4505
R58695 DVSS.n3609 DVSS.n3608 0.4505
R58696 DVSS.n3587 DVSS.n3586 0.4505
R58697 DVSS.n3604 DVSS.n3603 0.4505
R58698 DVSS.n3602 DVSS.n3589 0.4505
R58699 DVSS.n3601 DVSS.n3600 0.4505
R58700 DVSS.n3591 DVSS.n3590 0.4505
R58701 DVSS.n3596 DVSS.n3595 0.4505
R58702 DVSS.n3594 DVSS.n3593 0.4505
R58703 DVSS.n1717 DVSS.n1716 0.4505
R58704 DVSS.n5009 DVSS.n5008 0.4505
R58705 DVSS.n1720 DVSS.n1714 0.4505
R58706 DVSS.n5014 DVSS.n5013 0.4505
R58707 DVSS.n5015 DVSS.n1712 0.4505
R58708 DVSS.n5017 DVSS.n5016 0.4505
R58709 DVSS.n1710 DVSS.n1709 0.4505
R58710 DVSS.n5022 DVSS.n5021 0.4505
R58711 DVSS.n5023 DVSS.n1708 0.4505
R58712 DVSS.n5025 DVSS.n5024 0.4505
R58713 DVSS.n1706 DVSS.n1705 0.4505
R58714 DVSS.n5030 DVSS.n5029 0.4505
R58715 DVSS.n5031 DVSS.n1704 0.4505
R58716 DVSS.n5033 DVSS.n5032 0.4505
R58717 DVSS.n1702 DVSS.n1701 0.4505
R58718 DVSS.n5038 DVSS.n5037 0.4505
R58719 DVSS.n5039 DVSS.n1700 0.4505
R58720 DVSS.n5041 DVSS.n5040 0.4505
R58721 DVSS.n1697 DVSS.n1686 0.4505
R58722 DVSS.n5084 DVSS.n5083 0.4505
R58723 DVSS.n5103 DVSS.n5102 0.4505
R58724 DVSS.n5105 DVSS.n5104 0.4505
R58725 DVSS.n5100 DVSS.n5099 0.4505
R58726 DVSS.n5110 DVSS.n5109 0.4505
R58727 DVSS.n5111 DVSS.n5098 0.4505
R58728 DVSS.n5113 DVSS.n5112 0.4505
R58729 DVSS.n5096 DVSS.n5095 0.4505
R58730 DVSS.n5118 DVSS.n5117 0.4505
R58731 DVSS.n5119 DVSS.n5094 0.4505
R58732 DVSS.n5121 DVSS.n5120 0.4505
R58733 DVSS.n5091 DVSS.n5090 0.4505
R58734 DVSS.n5126 DVSS.n5125 0.4505
R58735 DVSS.n5127 DVSS.n5089 0.4505
R58736 DVSS.n3881 DVSS.n3880 0.4505
R58737 DVSS.n3879 DVSS.n2078 0.4505
R58738 DVSS.n3878 DVSS.n3877 0.4505
R58739 DVSS.n3698 DVSS.n3697 0.4505
R58740 DVSS.n3873 DVSS.n3872 0.4505
R58741 DVSS.n3871 DVSS.n3700 0.4505
R58742 DVSS.n3870 DVSS.n3869 0.4505
R58743 DVSS.n3702 DVSS.n3701 0.4505
R58744 DVSS.n3865 DVSS.n3864 0.4505
R58745 DVSS.n3863 DVSS.n3704 0.4505
R58746 DVSS.n3862 DVSS.n3861 0.4505
R58747 DVSS.n3706 DVSS.n3705 0.4505
R58748 DVSS.n3857 DVSS.n3856 0.4505
R58749 DVSS.n3855 DVSS.n3708 0.4505
R58750 DVSS.n3854 DVSS.n3853 0.4505
R58751 DVSS.n3850 DVSS.n3709 0.4505
R58752 DVSS.n3849 DVSS.n3847 0.4505
R58753 DVSS.n3846 DVSS.n3710 0.4505
R58754 DVSS.n3845 DVSS.n3844 0.4505
R58755 DVSS.n3712 DVSS.n3711 0.4505
R58756 DVSS.n3840 DVSS.n3839 0.4505
R58757 DVSS.n3838 DVSS.n3715 0.4505
R58758 DVSS.n3837 DVSS.n3836 0.4505
R58759 DVSS.n3717 DVSS.n3716 0.4505
R58760 DVSS.n3832 DVSS.n3831 0.4505
R58761 DVSS.n3830 DVSS.n3719 0.4505
R58762 DVSS.n3829 DVSS.n3828 0.4505
R58763 DVSS.n3721 DVSS.n3720 0.4505
R58764 DVSS.n3824 DVSS.n3823 0.4505
R58765 DVSS.n3822 DVSS.n3723 0.4505
R58766 DVSS.n3821 DVSS.n3820 0.4505
R58767 DVSS.n3725 DVSS.n3724 0.4505
R58768 DVSS.n3816 DVSS.n3815 0.4505
R58769 DVSS.n3814 DVSS.n3727 0.4505
R58770 DVSS.n3813 DVSS.n3812 0.4505
R58771 DVSS.n3729 DVSS.n3728 0.4505
R58772 DVSS.n3786 DVSS.n3785 0.4505
R58773 DVSS.n3784 DVSS.n3737 0.4505
R58774 DVSS.n3783 DVSS.n3782 0.4505
R58775 DVSS.n3739 DVSS.n3738 0.4505
R58776 DVSS.n3778 DVSS.n3777 0.4505
R58777 DVSS.n3776 DVSS.n3741 0.4505
R58778 DVSS.n3775 DVSS.n3774 0.4505
R58779 DVSS.n3743 DVSS.n3742 0.4505
R58780 DVSS.n3770 DVSS.n3769 0.4505
R58781 DVSS.n3768 DVSS.n3745 0.4505
R58782 DVSS.n3767 DVSS.n3766 0.4505
R58783 DVSS.n3747 DVSS.n3746 0.4505
R58784 DVSS.n3762 DVSS.n3761 0.4505
R58785 DVSS.n3760 DVSS.n3749 0.4505
R58786 DVSS.n3759 DVSS.n3758 0.4505
R58787 DVSS.n1660 DVSS.n1658 0.4505
R58788 DVSS.n5162 DVSS.n5161 0.4505
R58789 DVSS.n5160 DVSS.n1659 0.4505
R58790 DVSS.n5159 DVSS.n5158 0.4505
R58791 DVSS.n1662 DVSS.n1661 0.4505
R58792 DVSS.n5154 DVSS.n5153 0.4505
R58793 DVSS.n5152 DVSS.n1664 0.4505
R58794 DVSS.n5151 DVSS.n5150 0.4505
R58795 DVSS.n1666 DVSS.n1665 0.4505
R58796 DVSS.n5146 DVSS.n5145 0.4505
R58797 DVSS.n5144 DVSS.n1668 0.4505
R58798 DVSS.n5143 DVSS.n5142 0.4505
R58799 DVSS.n1670 DVSS.n1669 0.4505
R58800 DVSS.n5138 DVSS.n5137 0.4505
R58801 DVSS.n5136 DVSS.n1672 0.4505
R58802 DVSS.n5135 DVSS.n5134 0.4505
R58803 DVSS.n1674 DVSS.n1673 0.4505
R58804 DVSS.n5129 DVSS.n5128 0.4505
R58805 DVSS.n5106 DVSS.n5105 0.4505
R58806 DVSS.n5107 DVSS.n5100 0.4505
R58807 DVSS.n5109 DVSS.n5108 0.4505
R58808 DVSS.n5098 DVSS.n5097 0.4505
R58809 DVSS.n5114 DVSS.n5113 0.4505
R58810 DVSS.n5115 DVSS.n5096 0.4505
R58811 DVSS.n5117 DVSS.n5116 0.4505
R58812 DVSS.n5094 DVSS.n5093 0.4505
R58813 DVSS.n5122 DVSS.n5121 0.4505
R58814 DVSS.n5123 DVSS.n5091 0.4505
R58815 DVSS.n5125 DVSS.n5124 0.4505
R58816 DVSS.n5092 DVSS.n5089 0.4505
R58817 DVSS.n2077 DVSS.n2070 0.4505
R58818 DVSS.n3882 DVSS.n3881 0.4505
R58819 DVSS.n2078 DVSS.n2076 0.4505
R58820 DVSS.n3877 DVSS.n3876 0.4505
R58821 DVSS.n3875 DVSS.n3698 0.4505
R58822 DVSS.n3874 DVSS.n3873 0.4505
R58823 DVSS.n3700 DVSS.n3699 0.4505
R58824 DVSS.n3869 DVSS.n3868 0.4505
R58825 DVSS.n3867 DVSS.n3702 0.4505
R58826 DVSS.n3866 DVSS.n3865 0.4505
R58827 DVSS.n3704 DVSS.n3703 0.4505
R58828 DVSS.n3861 DVSS.n3860 0.4505
R58829 DVSS.n3859 DVSS.n3706 0.4505
R58830 DVSS.n3858 DVSS.n3857 0.4505
R58831 DVSS.n3708 DVSS.n3707 0.4505
R58832 DVSS.n3853 DVSS.n3852 0.4505
R58833 DVSS.n3851 DVSS.n3850 0.4505
R58834 DVSS.n3849 DVSS.n3848 0.4505
R58835 DVSS.n3713 DVSS.n3710 0.4505
R58836 DVSS.n3844 DVSS.n3843 0.4505
R58837 DVSS.n3842 DVSS.n3712 0.4505
R58838 DVSS.n3841 DVSS.n3840 0.4505
R58839 DVSS.n3715 DVSS.n3714 0.4505
R58840 DVSS.n3836 DVSS.n3835 0.4505
R58841 DVSS.n3834 DVSS.n3717 0.4505
R58842 DVSS.n3833 DVSS.n3832 0.4505
R58843 DVSS.n3719 DVSS.n3718 0.4505
R58844 DVSS.n3828 DVSS.n3827 0.4505
R58845 DVSS.n3826 DVSS.n3721 0.4505
R58846 DVSS.n3825 DVSS.n3824 0.4505
R58847 DVSS.n3723 DVSS.n3722 0.4505
R58848 DVSS.n3820 DVSS.n3819 0.4505
R58849 DVSS.n3818 DVSS.n3725 0.4505
R58850 DVSS.n3817 DVSS.n3816 0.4505
R58851 DVSS.n3806 DVSS.n3727 0.4505
R58852 DVSS.n3812 DVSS.n3811 0.4505
R58853 DVSS.n3788 DVSS.n3729 0.4505
R58854 DVSS.n3787 DVSS.n3786 0.4505
R58855 DVSS.n3737 DVSS.n3736 0.4505
R58856 DVSS.n3782 DVSS.n3781 0.4505
R58857 DVSS.n3780 DVSS.n3739 0.4505
R58858 DVSS.n3779 DVSS.n3778 0.4505
R58859 DVSS.n3741 DVSS.n3740 0.4505
R58860 DVSS.n3774 DVSS.n3773 0.4505
R58861 DVSS.n3772 DVSS.n3743 0.4505
R58862 DVSS.n3771 DVSS.n3770 0.4505
R58863 DVSS.n3745 DVSS.n3744 0.4505
R58864 DVSS.n3766 DVSS.n3765 0.4505
R58865 DVSS.n3764 DVSS.n3747 0.4505
R58866 DVSS.n3763 DVSS.n3762 0.4505
R58867 DVSS.n3749 DVSS.n3748 0.4505
R58868 DVSS.n3758 DVSS.n3757 0.4505
R58869 DVSS.n1658 DVSS.n1651 0.4505
R58870 DVSS.n5163 DVSS.n5162 0.4505
R58871 DVSS.n1659 DVSS.n1657 0.4505
R58872 DVSS.n5158 DVSS.n5157 0.4505
R58873 DVSS.n5156 DVSS.n1662 0.4505
R58874 DVSS.n5155 DVSS.n5154 0.4505
R58875 DVSS.n1664 DVSS.n1663 0.4505
R58876 DVSS.n5150 DVSS.n5149 0.4505
R58877 DVSS.n5148 DVSS.n1666 0.4505
R58878 DVSS.n5147 DVSS.n5146 0.4505
R58879 DVSS.n1668 DVSS.n1667 0.4505
R58880 DVSS.n5142 DVSS.n5141 0.4505
R58881 DVSS.n5140 DVSS.n1670 0.4505
R58882 DVSS.n5139 DVSS.n5138 0.4505
R58883 DVSS.n1672 DVSS.n1671 0.4505
R58884 DVSS.n5134 DVSS.n5133 0.4505
R58885 DVSS.n5132 DVSS.n1674 0.4505
R58886 DVSS.n5130 DVSS.n5129 0.4505
R58887 DVSS.n5524 DVSS.n5523 0.4505
R58888 DVSS.n5526 DVSS.n5525 0.4505
R58889 DVSS.n5521 DVSS.n5520 0.4505
R58890 DVSS.n5531 DVSS.n5530 0.4505
R58891 DVSS.n5532 DVSS.n5519 0.4505
R58892 DVSS.n5534 DVSS.n5533 0.4505
R58893 DVSS.n5517 DVSS.n5516 0.4505
R58894 DVSS.n5539 DVSS.n5538 0.4505
R58895 DVSS.n5540 DVSS.n5515 0.4505
R58896 DVSS.n5542 DVSS.n5541 0.4505
R58897 DVSS.n5512 DVSS.n5511 0.4505
R58898 DVSS.n5547 DVSS.n5546 0.4505
R58899 DVSS.n5548 DVSS.n5510 0.4505
R58900 DVSS.n3939 DVSS.n3938 0.4505
R58901 DVSS.n3937 DVSS.n3899 0.4505
R58902 DVSS.n3936 DVSS.n3935 0.4505
R58903 DVSS.n3902 DVSS.n3901 0.4505
R58904 DVSS.n3931 DVSS.n3930 0.4505
R58905 DVSS.n3929 DVSS.n3904 0.4505
R58906 DVSS.n3928 DVSS.n3927 0.4505
R58907 DVSS.n3906 DVSS.n3905 0.4505
R58908 DVSS.n3923 DVSS.n3922 0.4505
R58909 DVSS.n3921 DVSS.n3908 0.4505
R58910 DVSS.n3920 DVSS.n3919 0.4505
R58911 DVSS.n3910 DVSS.n3909 0.4505
R58912 DVSS.n3915 DVSS.n3914 0.4505
R58913 DVSS.n3913 DVSS.n3912 0.4505
R58914 DVSS.n2014 DVSS.n2013 0.4505
R58915 DVSS.n4648 DVSS.n4647 0.4505
R58916 DVSS.n4649 DVSS.n2012 0.4505
R58917 DVSS.n4651 DVSS.n4650 0.4505
R58918 DVSS.n2010 DVSS.n2009 0.4505
R58919 DVSS.n4656 DVSS.n4655 0.4505
R58920 DVSS.n4657 DVSS.n2008 0.4505
R58921 DVSS.n4659 DVSS.n4658 0.4505
R58922 DVSS.n2006 DVSS.n2005 0.4505
R58923 DVSS.n4664 DVSS.n4663 0.4505
R58924 DVSS.n4665 DVSS.n2004 0.4505
R58925 DVSS.n4667 DVSS.n4666 0.4505
R58926 DVSS.n2002 DVSS.n2001 0.4505
R58927 DVSS.n4672 DVSS.n4671 0.4505
R58928 DVSS.n4673 DVSS.n2000 0.4505
R58929 DVSS.n4675 DVSS.n4674 0.4505
R58930 DVSS.n1998 DVSS.n1997 0.4505
R58931 DVSS.n4681 DVSS.n4680 0.4505
R58932 DVSS.n4682 DVSS.n1995 0.4505
R58933 DVSS.n4738 DVSS.n4737 0.4505
R58934 DVSS.n4736 DVSS.n1996 0.4505
R58935 DVSS.n4735 DVSS.n4734 0.4505
R58936 DVSS.n4733 DVSS.n4683 0.4505
R58937 DVSS.n4687 DVSS.n4684 0.4505
R58938 DVSS.n4729 DVSS.n4728 0.4505
R58939 DVSS.n4727 DVSS.n4686 0.4505
R58940 DVSS.n4726 DVSS.n4725 0.4505
R58941 DVSS.n4689 DVSS.n4688 0.4505
R58942 DVSS.n4721 DVSS.n4720 0.4505
R58943 DVSS.n4719 DVSS.n4691 0.4505
R58944 DVSS.n4718 DVSS.n4717 0.4505
R58945 DVSS.n4693 DVSS.n4692 0.4505
R58946 DVSS.n4713 DVSS.n4712 0.4505
R58947 DVSS.n4711 DVSS.n4695 0.4505
R58948 DVSS.n4710 DVSS.n4709 0.4505
R58949 DVSS.n4697 DVSS.n4696 0.4505
R58950 DVSS.n4705 DVSS.n4704 0.4505
R58951 DVSS.n1344 DVSS.n1342 0.4505
R58952 DVSS.n5583 DVSS.n5582 0.4505
R58953 DVSS.n5581 DVSS.n1343 0.4505
R58954 DVSS.n5580 DVSS.n5579 0.4505
R58955 DVSS.n1346 DVSS.n1345 0.4505
R58956 DVSS.n5575 DVSS.n5574 0.4505
R58957 DVSS.n5573 DVSS.n1348 0.4505
R58958 DVSS.n5572 DVSS.n5571 0.4505
R58959 DVSS.n1350 DVSS.n1349 0.4505
R58960 DVSS.n5567 DVSS.n5566 0.4505
R58961 DVSS.n5565 DVSS.n1352 0.4505
R58962 DVSS.n5564 DVSS.n5563 0.4505
R58963 DVSS.n1354 DVSS.n1353 0.4505
R58964 DVSS.n5559 DVSS.n5558 0.4505
R58965 DVSS.n5557 DVSS.n1356 0.4505
R58966 DVSS.n5556 DVSS.n5555 0.4505
R58967 DVSS.n1358 DVSS.n1357 0.4505
R58968 DVSS.n5550 DVSS.n5549 0.4505
R58969 DVSS.n5527 DVSS.n5526 0.4505
R58970 DVSS.n5528 DVSS.n5521 0.4505
R58971 DVSS.n5530 DVSS.n5529 0.4505
R58972 DVSS.n5519 DVSS.n5518 0.4505
R58973 DVSS.n5535 DVSS.n5534 0.4505
R58974 DVSS.n5536 DVSS.n5517 0.4505
R58975 DVSS.n5538 DVSS.n5537 0.4505
R58976 DVSS.n5515 DVSS.n5514 0.4505
R58977 DVSS.n5543 DVSS.n5542 0.4505
R58978 DVSS.n5544 DVSS.n5512 0.4505
R58979 DVSS.n5546 DVSS.n5545 0.4505
R58980 DVSS.n5513 DVSS.n5510 0.4505
R58981 DVSS.n3898 DVSS.n3896 0.4505
R58982 DVSS.n3940 DVSS.n3939 0.4505
R58983 DVSS.n3899 DVSS.n3897 0.4505
R58984 DVSS.n3935 DVSS.n3934 0.4505
R58985 DVSS.n3933 DVSS.n3902 0.4505
R58986 DVSS.n3932 DVSS.n3931 0.4505
R58987 DVSS.n3904 DVSS.n3903 0.4505
R58988 DVSS.n3927 DVSS.n3926 0.4505
R58989 DVSS.n3925 DVSS.n3906 0.4505
R58990 DVSS.n3924 DVSS.n3923 0.4505
R58991 DVSS.n3908 DVSS.n3907 0.4505
R58992 DVSS.n3919 DVSS.n3918 0.4505
R58993 DVSS.n3917 DVSS.n3910 0.4505
R58994 DVSS.n3916 DVSS.n3915 0.4505
R58995 DVSS.n3912 DVSS.n3911 0.4505
R58996 DVSS.n2015 DVSS.n2014 0.4505
R58997 DVSS.n4647 DVSS.n4646 0.4505
R58998 DVSS.n2016 DVSS.n2012 0.4505
R58999 DVSS.n4652 DVSS.n4651 0.4505
R59000 DVSS.n4653 DVSS.n2010 0.4505
R59001 DVSS.n4655 DVSS.n4654 0.4505
R59002 DVSS.n2008 DVSS.n2007 0.4505
R59003 DVSS.n4660 DVSS.n4659 0.4505
R59004 DVSS.n4661 DVSS.n2006 0.4505
R59005 DVSS.n4663 DVSS.n4662 0.4505
R59006 DVSS.n2004 DVSS.n2003 0.4505
R59007 DVSS.n4668 DVSS.n4667 0.4505
R59008 DVSS.n4669 DVSS.n2002 0.4505
R59009 DVSS.n4671 DVSS.n4670 0.4505
R59010 DVSS.n2000 DVSS.n1999 0.4505
R59011 DVSS.n4676 DVSS.n4675 0.4505
R59012 DVSS.n4677 DVSS.n1998 0.4505
R59013 DVSS.n4680 DVSS.n4679 0.4505
R59014 DVSS.n4678 DVSS.n1995 0.4505
R59015 DVSS.n4739 DVSS.n4738 0.4505
R59016 DVSS.n1996 DVSS.n1974 0.4505
R59017 DVSS.n4734 DVSS.n1980 0.4505
R59018 DVSS.n4733 DVSS.n4732 0.4505
R59019 DVSS.n4731 DVSS.n4684 0.4505
R59020 DVSS.n4730 DVSS.n4729 0.4505
R59021 DVSS.n4686 DVSS.n4685 0.4505
R59022 DVSS.n4725 DVSS.n4724 0.4505
R59023 DVSS.n4723 DVSS.n4689 0.4505
R59024 DVSS.n4722 DVSS.n4721 0.4505
R59025 DVSS.n4691 DVSS.n4690 0.4505
R59026 DVSS.n4717 DVSS.n4716 0.4505
R59027 DVSS.n4715 DVSS.n4693 0.4505
R59028 DVSS.n4714 DVSS.n4713 0.4505
R59029 DVSS.n4695 DVSS.n4694 0.4505
R59030 DVSS.n4709 DVSS.n4708 0.4505
R59031 DVSS.n4707 DVSS.n4697 0.4505
R59032 DVSS.n4706 DVSS.n4705 0.4505
R59033 DVSS.n1342 DVSS.n1335 0.4505
R59034 DVSS.n5584 DVSS.n5583 0.4505
R59035 DVSS.n1343 DVSS.n1341 0.4505
R59036 DVSS.n5579 DVSS.n5578 0.4505
R59037 DVSS.n5577 DVSS.n1346 0.4505
R59038 DVSS.n5576 DVSS.n5575 0.4505
R59039 DVSS.n1348 DVSS.n1347 0.4505
R59040 DVSS.n5571 DVSS.n5570 0.4505
R59041 DVSS.n5569 DVSS.n1350 0.4505
R59042 DVSS.n5568 DVSS.n5567 0.4505
R59043 DVSS.n1352 DVSS.n1351 0.4505
R59044 DVSS.n5563 DVSS.n5562 0.4505
R59045 DVSS.n5561 DVSS.n1354 0.4505
R59046 DVSS.n5560 DVSS.n5559 0.4505
R59047 DVSS.n1356 DVSS.n1355 0.4505
R59048 DVSS.n5555 DVSS.n5554 0.4505
R59049 DVSS.n5553 DVSS.n1358 0.4505
R59050 DVSS.n5551 DVSS.n5550 0.4505
R59051 DVSS.n5983 DVSS.n5982 0.4505
R59052 DVSS.n5985 DVSS.n5984 0.4505
R59053 DVSS.n5980 DVSS.n5979 0.4505
R59054 DVSS.n5990 DVSS.n5989 0.4505
R59055 DVSS.n5991 DVSS.n5978 0.4505
R59056 DVSS.n5993 DVSS.n5992 0.4505
R59057 DVSS.n5976 DVSS.n5975 0.4505
R59058 DVSS.n5998 DVSS.n5997 0.4505
R59059 DVSS.n5999 DVSS.n5973 0.4505
R59060 DVSS.n6001 DVSS.n6000 0.4505
R59061 DVSS.n5974 DVSS.n5971 0.4505
R59062 DVSS.n6005 DVSS.n5970 0.4505
R59063 DVSS.n6007 DVSS.n6006 0.4505
R59064 DVSS.n5857 DVSS.n5856 0.4505
R59065 DVSS.n5858 DVSS.n5854 0.4505
R59066 DVSS.n5862 DVSS.n5861 0.4505
R59067 DVSS.n5863 DVSS.n5853 0.4505
R59068 DVSS.n5865 DVSS.n5864 0.4505
R59069 DVSS.n5851 DVSS.n5850 0.4505
R59070 DVSS.n5870 DVSS.n5869 0.4505
R59071 DVSS.n5871 DVSS.n5849 0.4505
R59072 DVSS.n5873 DVSS.n5872 0.4505
R59073 DVSS.n5847 DVSS.n5846 0.4505
R59074 DVSS.n5878 DVSS.n5877 0.4505
R59075 DVSS.n5879 DVSS.n5845 0.4505
R59076 DVSS.n5882 DVSS.n5881 0.4505
R59077 DVSS.n5880 DVSS.n5842 0.4505
R59078 DVSS.n5886 DVSS.n5843 0.4505
R59079 DVSS.n5887 DVSS.n5841 0.4505
R59080 DVSS.n5889 DVSS.n5888 0.4505
R59081 DVSS.n5890 DVSS.n5840 0.4505
R59082 DVSS.n5892 DVSS.n5891 0.4505
R59083 DVSS.n5839 DVSS.n5838 0.4505
R59084 DVSS.n5897 DVSS.n5896 0.4505
R59085 DVSS.n5898 DVSS.n5837 0.4505
R59086 DVSS.n5900 DVSS.n5899 0.4505
R59087 DVSS.n5835 DVSS.n5834 0.4505
R59088 DVSS.n5905 DVSS.n5904 0.4505
R59089 DVSS.n5906 DVSS.n5833 0.4505
R59090 DVSS.n5908 DVSS.n5907 0.4505
R59091 DVSS.n5831 DVSS.n5830 0.4505
R59092 DVSS.n5913 DVSS.n5912 0.4505
R59093 DVSS.n5914 DVSS.n5829 0.4505
R59094 DVSS.n5916 DVSS.n5915 0.4505
R59095 DVSS.n5827 DVSS.n5826 0.4505
R59096 DVSS.n5921 DVSS.n5920 0.4505
R59097 DVSS.n5922 DVSS.n5825 0.4505
R59098 DVSS.n5924 DVSS.n5923 0.4505
R59099 DVSS.n5925 DVSS.n5823 0.4505
R59100 DVSS.n5928 DVSS.n5927 0.4505
R59101 DVSS.n5929 DVSS.n5822 0.4505
R59102 DVSS.n5931 DVSS.n5930 0.4505
R59103 DVSS.n5820 DVSS.n5819 0.4505
R59104 DVSS.n5936 DVSS.n5935 0.4505
R59105 DVSS.n5937 DVSS.n5818 0.4505
R59106 DVSS.n5939 DVSS.n5938 0.4505
R59107 DVSS.n5816 DVSS.n5815 0.4505
R59108 DVSS.n5944 DVSS.n5943 0.4505
R59109 DVSS.n5945 DVSS.n5814 0.4505
R59110 DVSS.n5947 DVSS.n5946 0.4505
R59111 DVSS.n5812 DVSS.n5811 0.4505
R59112 DVSS.n5952 DVSS.n5951 0.4505
R59113 DVSS.n5953 DVSS.n5809 0.4505
R59114 DVSS.n6043 DVSS.n6042 0.4505
R59115 DVSS.n6041 DVSS.n5810 0.4505
R59116 DVSS.n6040 DVSS.n6039 0.4505
R59117 DVSS.n6038 DVSS.n5954 0.4505
R59118 DVSS.n5958 DVSS.n5955 0.4505
R59119 DVSS.n6034 DVSS.n6033 0.4505
R59120 DVSS.n6032 DVSS.n5957 0.4505
R59121 DVSS.n6031 DVSS.n6030 0.4505
R59122 DVSS.n5960 DVSS.n5959 0.4505
R59123 DVSS.n6026 DVSS.n6025 0.4505
R59124 DVSS.n6024 DVSS.n5962 0.4505
R59125 DVSS.n6023 DVSS.n6022 0.4505
R59126 DVSS.n5964 DVSS.n5963 0.4505
R59127 DVSS.n6018 DVSS.n6017 0.4505
R59128 DVSS.n6016 DVSS.n5966 0.4505
R59129 DVSS.n6015 DVSS.n6014 0.4505
R59130 DVSS.n5968 DVSS.n5967 0.4505
R59131 DVSS.n6010 DVSS.n6009 0.4505
R59132 DVSS.n6008 DVSS.n5969 0.4505
R59133 DVSS.n5986 DVSS.n5985 0.4505
R59134 DVSS.n5987 DVSS.n5980 0.4505
R59135 DVSS.n5989 DVSS.n5988 0.4505
R59136 DVSS.n5978 DVSS.n5977 0.4505
R59137 DVSS.n5994 DVSS.n5993 0.4505
R59138 DVSS.n5995 DVSS.n5976 0.4505
R59139 DVSS.n5997 DVSS.n5996 0.4505
R59140 DVSS.n5973 DVSS.n5972 0.4505
R59141 DVSS.n6002 DVSS.n6001 0.4505
R59142 DVSS.n6003 DVSS.n5971 0.4505
R59143 DVSS.n6005 DVSS.n6004 0.4505
R59144 DVSS.n6006 DVSS.n1192 0.4505
R59145 DVSS.n5855 DVSS.n1159 0.4505
R59146 DVSS.n5857 DVSS.n1162 0.4505
R59147 DVSS.n5859 DVSS.n5858 0.4505
R59148 DVSS.n5861 DVSS.n5860 0.4505
R59149 DVSS.n5853 DVSS.n5852 0.4505
R59150 DVSS.n5866 DVSS.n5865 0.4505
R59151 DVSS.n5867 DVSS.n5851 0.4505
R59152 DVSS.n5869 DVSS.n5868 0.4505
R59153 DVSS.n5849 DVSS.n5848 0.4505
R59154 DVSS.n5874 DVSS.n5873 0.4505
R59155 DVSS.n5875 DVSS.n5847 0.4505
R59156 DVSS.n5877 DVSS.n5876 0.4505
R59157 DVSS.n5845 DVSS.n5844 0.4505
R59158 DVSS.n5883 DVSS.n5882 0.4505
R59159 DVSS.n5884 DVSS.n5842 0.4505
R59160 DVSS.n5886 DVSS.n5885 0.4505
R59161 DVSS.n5887 DVSS.n1152 0.4505
R59162 DVSS.n5888 DVSS.n1143 0.4505
R59163 DVSS.n5840 DVSS.n1147 0.4505
R59164 DVSS.n5893 DVSS.n5892 0.4505
R59165 DVSS.n5894 DVSS.n5839 0.4505
R59166 DVSS.n5896 DVSS.n5895 0.4505
R59167 DVSS.n5837 DVSS.n5836 0.4505
R59168 DVSS.n5901 DVSS.n5900 0.4505
R59169 DVSS.n5902 DVSS.n5835 0.4505
R59170 DVSS.n5904 DVSS.n5903 0.4505
R59171 DVSS.n5833 DVSS.n5832 0.4505
R59172 DVSS.n5909 DVSS.n5908 0.4505
R59173 DVSS.n5910 DVSS.n5831 0.4505
R59174 DVSS.n5912 DVSS.n5911 0.4505
R59175 DVSS.n5829 DVSS.n5828 0.4505
R59176 DVSS.n5917 DVSS.n5916 0.4505
R59177 DVSS.n5918 DVSS.n5827 0.4505
R59178 DVSS.n5920 DVSS.n5919 0.4505
R59179 DVSS.n5825 DVSS.n5824 0.4505
R59180 DVSS.n5924 DVSS.n5777 0.4505
R59181 DVSS.n5925 DVSS.n5781 0.4505
R59182 DVSS.n5927 DVSS.n5926 0.4505
R59183 DVSS.n5822 DVSS.n5821 0.4505
R59184 DVSS.n5932 DVSS.n5931 0.4505
R59185 DVSS.n5933 DVSS.n5820 0.4505
R59186 DVSS.n5935 DVSS.n5934 0.4505
R59187 DVSS.n5818 DVSS.n5817 0.4505
R59188 DVSS.n5940 DVSS.n5939 0.4505
R59189 DVSS.n5941 DVSS.n5816 0.4505
R59190 DVSS.n5943 DVSS.n5942 0.4505
R59191 DVSS.n5814 DVSS.n5813 0.4505
R59192 DVSS.n5948 DVSS.n5947 0.4505
R59193 DVSS.n5949 DVSS.n5812 0.4505
R59194 DVSS.n5951 DVSS.n5950 0.4505
R59195 DVSS.n5809 DVSS.n5808 0.4505
R59196 DVSS.n6044 DVSS.n6043 0.4505
R59197 DVSS.n5810 DVSS.n5802 0.4505
R59198 DVSS.n6039 DVSS.n5804 0.4505
R59199 DVSS.n6038 DVSS.n6037 0.4505
R59200 DVSS.n6036 DVSS.n5955 0.4505
R59201 DVSS.n6035 DVSS.n6034 0.4505
R59202 DVSS.n5957 DVSS.n5956 0.4505
R59203 DVSS.n6030 DVSS.n6029 0.4505
R59204 DVSS.n6028 DVSS.n5960 0.4505
R59205 DVSS.n6027 DVSS.n6026 0.4505
R59206 DVSS.n5962 DVSS.n5961 0.4505
R59207 DVSS.n6022 DVSS.n6021 0.4505
R59208 DVSS.n6020 DVSS.n5964 0.4505
R59209 DVSS.n6019 DVSS.n6018 0.4505
R59210 DVSS.n5966 DVSS.n5965 0.4505
R59211 DVSS.n6014 DVSS.n6013 0.4505
R59212 DVSS.n6012 DVSS.n5968 0.4505
R59213 DVSS.n6011 DVSS.n6010 0.4505
R59214 DVSS.n5969 DVSS.n1185 0.4505
R59215 DVSS.n2273 DVSS.n2232 0.4505
R59216 DVSS.n2272 DVSS.n2271 0.4505
R59217 DVSS.n2234 DVSS.n2233 0.4505
R59218 DVSS.n2267 DVSS.n2266 0.4505
R59219 DVSS.n2265 DVSS.n2236 0.4505
R59220 DVSS.n2264 DVSS.n2263 0.4505
R59221 DVSS.n2238 DVSS.n2237 0.4505
R59222 DVSS.n2259 DVSS.n2258 0.4505
R59223 DVSS.n2257 DVSS.n2240 0.4505
R59224 DVSS.n2256 DVSS.n2255 0.4505
R59225 DVSS.n2252 DVSS.n2241 0.4505
R59226 DVSS.n2251 DVSS.n2250 0.4505
R59227 DVSS.n2249 DVSS.n2243 0.4505
R59228 DVSS.n3500 DVSS.n3499 0.4505
R59229 DVSS.n2146 DVSS.n2145 0.4505
R59230 DVSS.n3495 DVSS.n3494 0.4505
R59231 DVSS.n3493 DVSS.n2148 0.4505
R59232 DVSS.n3492 DVSS.n3491 0.4505
R59233 DVSS.n2150 DVSS.n2149 0.4505
R59234 DVSS.n3487 DVSS.n3486 0.4505
R59235 DVSS.n3485 DVSS.n2152 0.4505
R59236 DVSS.n3484 DVSS.n3483 0.4505
R59237 DVSS.n2154 DVSS.n2153 0.4505
R59238 DVSS.n3479 DVSS.n3478 0.4505
R59239 DVSS.n3477 DVSS.n2156 0.4505
R59240 DVSS.n3476 DVSS.n3475 0.4505
R59241 DVSS.n2158 DVSS.n2157 0.4505
R59242 DVSS.n3471 DVSS.n3470 0.4505
R59243 DVSS.n3469 DVSS.n2160 0.4505
R59244 DVSS.n3468 DVSS.n3467 0.4505
R59245 DVSS.n2162 DVSS.n2161 0.4505
R59246 DVSS.n3463 DVSS.n3462 0.4505
R59247 DVSS.n3461 DVSS.n2164 0.4505
R59248 DVSS.n3460 DVSS.n3459 0.4505
R59249 DVSS.n2166 DVSS.n2165 0.4505
R59250 DVSS.n3455 DVSS.n3454 0.4505
R59251 DVSS.n3453 DVSS.n2168 0.4505
R59252 DVSS.n3452 DVSS.n3451 0.4505
R59253 DVSS.n2170 DVSS.n2169 0.4505
R59254 DVSS.n3447 DVSS.n3446 0.4505
R59255 DVSS.n3445 DVSS.n2172 0.4505
R59256 DVSS.n3444 DVSS.n3443 0.4505
R59257 DVSS.n2174 DVSS.n2173 0.4505
R59258 DVSS.n3439 DVSS.n3438 0.4505
R59259 DVSS.n3437 DVSS.n2176 0.4505
R59260 DVSS.n3436 DVSS.n3435 0.4505
R59261 DVSS.n2178 DVSS.n2177 0.4505
R59262 DVSS.n3431 DVSS.n3430 0.4505
R59263 DVSS.n3429 DVSS.n2180 0.4505
R59264 DVSS.n3428 DVSS.n3427 0.4505
R59265 DVSS.n2182 DVSS.n2181 0.4505
R59266 DVSS.n3423 DVSS.n3422 0.4505
R59267 DVSS.n3421 DVSS.n2184 0.4505
R59268 DVSS.n3420 DVSS.n3419 0.4505
R59269 DVSS.n2186 DVSS.n2185 0.4505
R59270 DVSS.n3415 DVSS.n3414 0.4505
R59271 DVSS.n3413 DVSS.n2188 0.4505
R59272 DVSS.n3412 DVSS.n3411 0.4505
R59273 DVSS.n2190 DVSS.n2189 0.4505
R59274 DVSS.n3407 DVSS.n3406 0.4505
R59275 DVSS.n3405 DVSS.n2192 0.4505
R59276 DVSS.n3404 DVSS.n3403 0.4505
R59277 DVSS.n2194 DVSS.n2193 0.4505
R59278 DVSS.n3399 DVSS.n3398 0.4505
R59279 DVSS.n3397 DVSS.n2196 0.4505
R59280 DVSS.n3396 DVSS.n3395 0.4505
R59281 DVSS.n2198 DVSS.n2197 0.4505
R59282 DVSS.n3391 DVSS.n3390 0.4505
R59283 DVSS.n3389 DVSS.n2200 0.4505
R59284 DVSS.n3388 DVSS.n3387 0.4505
R59285 DVSS.n2202 DVSS.n2201 0.4505
R59286 DVSS.n3383 DVSS.n3382 0.4505
R59287 DVSS.n3381 DVSS.n2204 0.4505
R59288 DVSS.n3380 DVSS.n3379 0.4505
R59289 DVSS.n2206 DVSS.n2205 0.4505
R59290 DVSS.n3375 DVSS.n3374 0.4505
R59291 DVSS.n3373 DVSS.n2208 0.4505
R59292 DVSS.n3372 DVSS.n3371 0.4505
R59293 DVSS.n2210 DVSS.n2209 0.4505
R59294 DVSS.n3367 DVSS.n3366 0.4505
R59295 DVSS.n3365 DVSS.n2212 0.4505
R59296 DVSS.n3364 DVSS.n3363 0.4505
R59297 DVSS.n2214 DVSS.n2213 0.4505
R59298 DVSS.n3359 DVSS.n3358 0.4505
R59299 DVSS.n3357 DVSS.n2216 0.4505
R59300 DVSS.n3356 DVSS.n3355 0.4505
R59301 DVSS.n2218 DVSS.n2217 0.4505
R59302 DVSS.n3351 DVSS.n3350 0.4505
R59303 DVSS.n3349 DVSS.n2220 0.4505
R59304 DVSS.n3348 DVSS.n3347 0.4505
R59305 DVSS.n2222 DVSS.n2221 0.4505
R59306 DVSS.n3343 DVSS.n3342 0.4505
R59307 DVSS.n3341 DVSS.n2224 0.4505
R59308 DVSS.n3340 DVSS.n3339 0.4505
R59309 DVSS.n2226 DVSS.n2225 0.4505
R59310 DVSS.n3335 DVSS.n3334 0.4505
R59311 DVSS.n3333 DVSS.n2228 0.4505
R59312 DVSS.n3332 DVSS.n3331 0.4505
R59313 DVSS.n2230 DVSS.n2229 0.4505
R59314 DVSS.n2275 DVSS.n2274 0.4505
R59315 DVSS.n3299 DVSS.n3280 0.4505
R59316 DVSS.n3301 DVSS.n3300 0.4505
R59317 DVSS.n3302 DVSS.n3278 0.4505
R59318 DVSS.n3306 DVSS.n3305 0.4505
R59319 DVSS.n3307 DVSS.n3277 0.4505
R59320 DVSS.n3309 DVSS.n3308 0.4505
R59321 DVSS.n3275 DVSS.n3274 0.4505
R59322 DVSS.n3314 DVSS.n3313 0.4505
R59323 DVSS.n3315 DVSS.n3273 0.4505
R59324 DVSS.n3317 DVSS.n3316 0.4505
R59325 DVSS.n3271 DVSS.n3270 0.4505
R59326 DVSS.n3322 DVSS.n3321 0.4505
R59327 DVSS.n3323 DVSS.n2280 0.4505
R59328 DVSS.n3100 DVSS.n3099 0.4505
R59329 DVSS.n3101 DVSS.n2364 0.4505
R59330 DVSS.n3103 DVSS.n3102 0.4505
R59331 DVSS.n2362 DVSS.n2361 0.4505
R59332 DVSS.n3108 DVSS.n3107 0.4505
R59333 DVSS.n3109 DVSS.n2360 0.4505
R59334 DVSS.n3111 DVSS.n3110 0.4505
R59335 DVSS.n2358 DVSS.n2357 0.4505
R59336 DVSS.n3116 DVSS.n3115 0.4505
R59337 DVSS.n3117 DVSS.n2356 0.4505
R59338 DVSS.n3119 DVSS.n3118 0.4505
R59339 DVSS.n2354 DVSS.n2353 0.4505
R59340 DVSS.n3124 DVSS.n3123 0.4505
R59341 DVSS.n3125 DVSS.n2352 0.4505
R59342 DVSS.n3127 DVSS.n3126 0.4505
R59343 DVSS.n2350 DVSS.n2349 0.4505
R59344 DVSS.n3132 DVSS.n3131 0.4505
R59345 DVSS.n3133 DVSS.n2348 0.4505
R59346 DVSS.n3135 DVSS.n3134 0.4505
R59347 DVSS.n2346 DVSS.n2345 0.4505
R59348 DVSS.n3140 DVSS.n3139 0.4505
R59349 DVSS.n3141 DVSS.n2344 0.4505
R59350 DVSS.n3143 DVSS.n3142 0.4505
R59351 DVSS.n2342 DVSS.n2341 0.4505
R59352 DVSS.n3148 DVSS.n3147 0.4505
R59353 DVSS.n3149 DVSS.n2340 0.4505
R59354 DVSS.n3151 DVSS.n3150 0.4505
R59355 DVSS.n2338 DVSS.n2337 0.4505
R59356 DVSS.n3156 DVSS.n3155 0.4505
R59357 DVSS.n3157 DVSS.n2336 0.4505
R59358 DVSS.n3159 DVSS.n3158 0.4505
R59359 DVSS.n2334 DVSS.n2333 0.4505
R59360 DVSS.n3164 DVSS.n3163 0.4505
R59361 DVSS.n3165 DVSS.n2332 0.4505
R59362 DVSS.n3167 DVSS.n3166 0.4505
R59363 DVSS.n2330 DVSS.n2329 0.4505
R59364 DVSS.n3172 DVSS.n3171 0.4505
R59365 DVSS.n3173 DVSS.n2328 0.4505
R59366 DVSS.n3175 DVSS.n3174 0.4505
R59367 DVSS.n2326 DVSS.n2325 0.4505
R59368 DVSS.n3180 DVSS.n3179 0.4505
R59369 DVSS.n3181 DVSS.n2324 0.4505
R59370 DVSS.n3183 DVSS.n3182 0.4505
R59371 DVSS.n2322 DVSS.n2321 0.4505
R59372 DVSS.n3188 DVSS.n3187 0.4505
R59373 DVSS.n3189 DVSS.n2320 0.4505
R59374 DVSS.n3191 DVSS.n3190 0.4505
R59375 DVSS.n2318 DVSS.n2317 0.4505
R59376 DVSS.n3196 DVSS.n3195 0.4505
R59377 DVSS.n3197 DVSS.n2316 0.4505
R59378 DVSS.n3199 DVSS.n3198 0.4505
R59379 DVSS.n2314 DVSS.n2313 0.4505
R59380 DVSS.n3204 DVSS.n3203 0.4505
R59381 DVSS.n3205 DVSS.n2312 0.4505
R59382 DVSS.n3207 DVSS.n3206 0.4505
R59383 DVSS.n2310 DVSS.n2309 0.4505
R59384 DVSS.n3212 DVSS.n3211 0.4505
R59385 DVSS.n3213 DVSS.n2308 0.4505
R59386 DVSS.n3215 DVSS.n3214 0.4505
R59387 DVSS.n2306 DVSS.n2305 0.4505
R59388 DVSS.n3220 DVSS.n3219 0.4505
R59389 DVSS.n3221 DVSS.n2304 0.4505
R59390 DVSS.n3223 DVSS.n3222 0.4505
R59391 DVSS.n2302 DVSS.n2301 0.4505
R59392 DVSS.n3228 DVSS.n3227 0.4505
R59393 DVSS.n3229 DVSS.n2300 0.4505
R59394 DVSS.n3231 DVSS.n3230 0.4505
R59395 DVSS.n2298 DVSS.n2297 0.4505
R59396 DVSS.n3236 DVSS.n3235 0.4505
R59397 DVSS.n3237 DVSS.n2296 0.4505
R59398 DVSS.n3239 DVSS.n3238 0.4505
R59399 DVSS.n2294 DVSS.n2293 0.4505
R59400 DVSS.n3244 DVSS.n3243 0.4505
R59401 DVSS.n3245 DVSS.n2292 0.4505
R59402 DVSS.n3247 DVSS.n3246 0.4505
R59403 DVSS.n2290 DVSS.n2289 0.4505
R59404 DVSS.n3252 DVSS.n3251 0.4505
R59405 DVSS.n3253 DVSS.n2288 0.4505
R59406 DVSS.n3255 DVSS.n3254 0.4505
R59407 DVSS.n2286 DVSS.n2285 0.4505
R59408 DVSS.n3260 DVSS.n3259 0.4505
R59409 DVSS.n3261 DVSS.n2284 0.4505
R59410 DVSS.n3263 DVSS.n3262 0.4505
R59411 DVSS.n2282 DVSS.n2281 0.4505
R59412 DVSS.n3268 DVSS.n3267 0.4505
R59413 DVSS.n3269 DVSS.n2279 0.4505
R59414 DVSS.n3325 DVSS.n3324 0.4505
R59415 DVSS.n2280 DVSS.n2278 0.4505
R59416 DVSS.n3321 DVSS.n3320 0.4505
R59417 DVSS.n3319 DVSS.n3271 0.4505
R59418 DVSS.n3318 DVSS.n3317 0.4505
R59419 DVSS.n3273 DVSS.n3272 0.4505
R59420 DVSS.n3313 DVSS.n3312 0.4505
R59421 DVSS.n3311 DVSS.n3275 0.4505
R59422 DVSS.n3310 DVSS.n3309 0.4505
R59423 DVSS.n3277 DVSS.n3276 0.4505
R59424 DVSS.n3305 DVSS.n3304 0.4505
R59425 DVSS.n3303 DVSS.n3302 0.4505
R59426 DVSS.n3301 DVSS.n3279 0.4505
R59427 DVSS.n3295 DVSS.n3280 0.4505
R59428 DVSS.n3297 DVSS.n3296 0.4505
R59429 DVSS.n3097 DVSS.n2366 0.4505
R59430 DVSS.n3099 DVSS.n3098 0.4505
R59431 DVSS.n2364 DVSS.n2363 0.4505
R59432 DVSS.n3104 DVSS.n3103 0.4505
R59433 DVSS.n3105 DVSS.n2362 0.4505
R59434 DVSS.n3107 DVSS.n3106 0.4505
R59435 DVSS.n2360 DVSS.n2359 0.4505
R59436 DVSS.n3112 DVSS.n3111 0.4505
R59437 DVSS.n3113 DVSS.n2358 0.4505
R59438 DVSS.n3115 DVSS.n3114 0.4505
R59439 DVSS.n2356 DVSS.n2355 0.4505
R59440 DVSS.n3120 DVSS.n3119 0.4505
R59441 DVSS.n3121 DVSS.n2354 0.4505
R59442 DVSS.n3123 DVSS.n3122 0.4505
R59443 DVSS.n2352 DVSS.n2351 0.4505
R59444 DVSS.n3128 DVSS.n3127 0.4505
R59445 DVSS.n3129 DVSS.n2350 0.4505
R59446 DVSS.n3131 DVSS.n3130 0.4505
R59447 DVSS.n2348 DVSS.n2347 0.4505
R59448 DVSS.n3136 DVSS.n3135 0.4505
R59449 DVSS.n3137 DVSS.n2346 0.4505
R59450 DVSS.n3139 DVSS.n3138 0.4505
R59451 DVSS.n2344 DVSS.n2343 0.4505
R59452 DVSS.n3144 DVSS.n3143 0.4505
R59453 DVSS.n3145 DVSS.n2342 0.4505
R59454 DVSS.n3147 DVSS.n3146 0.4505
R59455 DVSS.n2340 DVSS.n2339 0.4505
R59456 DVSS.n3152 DVSS.n3151 0.4505
R59457 DVSS.n3153 DVSS.n2338 0.4505
R59458 DVSS.n3155 DVSS.n3154 0.4505
R59459 DVSS.n2336 DVSS.n2335 0.4505
R59460 DVSS.n3160 DVSS.n3159 0.4505
R59461 DVSS.n3161 DVSS.n2334 0.4505
R59462 DVSS.n3163 DVSS.n3162 0.4505
R59463 DVSS.n2332 DVSS.n2331 0.4505
R59464 DVSS.n3168 DVSS.n3167 0.4505
R59465 DVSS.n3169 DVSS.n2330 0.4505
R59466 DVSS.n3171 DVSS.n3170 0.4505
R59467 DVSS.n2328 DVSS.n2327 0.4505
R59468 DVSS.n3176 DVSS.n3175 0.4505
R59469 DVSS.n3177 DVSS.n2326 0.4505
R59470 DVSS.n3179 DVSS.n3178 0.4505
R59471 DVSS.n2324 DVSS.n2323 0.4505
R59472 DVSS.n3184 DVSS.n3183 0.4505
R59473 DVSS.n3185 DVSS.n2322 0.4505
R59474 DVSS.n3187 DVSS.n3186 0.4505
R59475 DVSS.n2320 DVSS.n2319 0.4505
R59476 DVSS.n3192 DVSS.n3191 0.4505
R59477 DVSS.n3193 DVSS.n2318 0.4505
R59478 DVSS.n3195 DVSS.n3194 0.4505
R59479 DVSS.n2316 DVSS.n2315 0.4505
R59480 DVSS.n3200 DVSS.n3199 0.4505
R59481 DVSS.n3201 DVSS.n2314 0.4505
R59482 DVSS.n3203 DVSS.n3202 0.4505
R59483 DVSS.n2312 DVSS.n2311 0.4505
R59484 DVSS.n3208 DVSS.n3207 0.4505
R59485 DVSS.n3209 DVSS.n2310 0.4505
R59486 DVSS.n3211 DVSS.n3210 0.4505
R59487 DVSS.n2308 DVSS.n2307 0.4505
R59488 DVSS.n3216 DVSS.n3215 0.4505
R59489 DVSS.n3217 DVSS.n2306 0.4505
R59490 DVSS.n3219 DVSS.n3218 0.4505
R59491 DVSS.n2304 DVSS.n2303 0.4505
R59492 DVSS.n3224 DVSS.n3223 0.4505
R59493 DVSS.n3225 DVSS.n2302 0.4505
R59494 DVSS.n3227 DVSS.n3226 0.4505
R59495 DVSS.n2300 DVSS.n2299 0.4505
R59496 DVSS.n3232 DVSS.n3231 0.4505
R59497 DVSS.n3233 DVSS.n2298 0.4505
R59498 DVSS.n3235 DVSS.n3234 0.4505
R59499 DVSS.n2296 DVSS.n2295 0.4505
R59500 DVSS.n3240 DVSS.n3239 0.4505
R59501 DVSS.n3241 DVSS.n2294 0.4505
R59502 DVSS.n3243 DVSS.n3242 0.4505
R59503 DVSS.n2292 DVSS.n2291 0.4505
R59504 DVSS.n3248 DVSS.n3247 0.4505
R59505 DVSS.n3249 DVSS.n2290 0.4505
R59506 DVSS.n3251 DVSS.n3250 0.4505
R59507 DVSS.n2288 DVSS.n2287 0.4505
R59508 DVSS.n3256 DVSS.n3255 0.4505
R59509 DVSS.n3257 DVSS.n2286 0.4505
R59510 DVSS.n3259 DVSS.n3258 0.4505
R59511 DVSS.n2284 DVSS.n2283 0.4505
R59512 DVSS.n3264 DVSS.n3263 0.4505
R59513 DVSS.n3265 DVSS.n2282 0.4505
R59514 DVSS.n3267 DVSS.n3266 0.4505
R59515 DVSS.n2279 DVSS.n2277 0.4505
R59516 DVSS.n3326 DVSS.n3325 0.4505
R59517 DVSS.n2232 DVSS.n2231 0.4505
R59518 DVSS.n2271 DVSS.n2270 0.4505
R59519 DVSS.n2269 DVSS.n2234 0.4505
R59520 DVSS.n2268 DVSS.n2267 0.4505
R59521 DVSS.n2236 DVSS.n2235 0.4505
R59522 DVSS.n2263 DVSS.n2262 0.4505
R59523 DVSS.n2261 DVSS.n2238 0.4505
R59524 DVSS.n2260 DVSS.n2259 0.4505
R59525 DVSS.n2240 DVSS.n2239 0.4505
R59526 DVSS.n2255 DVSS.n2254 0.4505
R59527 DVSS.n2253 DVSS.n2252 0.4505
R59528 DVSS.n2251 DVSS.n2242 0.4505
R59529 DVSS.n2245 DVSS.n2243 0.4505
R59530 DVSS.n2247 DVSS.n2246 0.4505
R59531 DVSS.n2144 DVSS.n2143 0.4505
R59532 DVSS.n3499 DVSS.n3498 0.4505
R59533 DVSS.n3497 DVSS.n2146 0.4505
R59534 DVSS.n3496 DVSS.n3495 0.4505
R59535 DVSS.n2148 DVSS.n2147 0.4505
R59536 DVSS.n3491 DVSS.n3490 0.4505
R59537 DVSS.n3489 DVSS.n2150 0.4505
R59538 DVSS.n3488 DVSS.n3487 0.4505
R59539 DVSS.n2152 DVSS.n2151 0.4505
R59540 DVSS.n3483 DVSS.n3482 0.4505
R59541 DVSS.n3481 DVSS.n2154 0.4505
R59542 DVSS.n3480 DVSS.n3479 0.4505
R59543 DVSS.n2156 DVSS.n2155 0.4505
R59544 DVSS.n3475 DVSS.n3474 0.4505
R59545 DVSS.n3473 DVSS.n2158 0.4505
R59546 DVSS.n3472 DVSS.n3471 0.4505
R59547 DVSS.n2160 DVSS.n2159 0.4505
R59548 DVSS.n3467 DVSS.n3466 0.4505
R59549 DVSS.n3465 DVSS.n2162 0.4505
R59550 DVSS.n3464 DVSS.n3463 0.4505
R59551 DVSS.n2164 DVSS.n2163 0.4505
R59552 DVSS.n3459 DVSS.n3458 0.4505
R59553 DVSS.n3457 DVSS.n2166 0.4505
R59554 DVSS.n3456 DVSS.n3455 0.4505
R59555 DVSS.n2168 DVSS.n2167 0.4505
R59556 DVSS.n3451 DVSS.n3450 0.4505
R59557 DVSS.n3449 DVSS.n2170 0.4505
R59558 DVSS.n3448 DVSS.n3447 0.4505
R59559 DVSS.n2172 DVSS.n2171 0.4505
R59560 DVSS.n3443 DVSS.n3442 0.4505
R59561 DVSS.n3441 DVSS.n2174 0.4505
R59562 DVSS.n3440 DVSS.n3439 0.4505
R59563 DVSS.n2176 DVSS.n2175 0.4505
R59564 DVSS.n3435 DVSS.n3434 0.4505
R59565 DVSS.n3433 DVSS.n2178 0.4505
R59566 DVSS.n3432 DVSS.n3431 0.4505
R59567 DVSS.n2180 DVSS.n2179 0.4505
R59568 DVSS.n3427 DVSS.n3426 0.4505
R59569 DVSS.n3425 DVSS.n2182 0.4505
R59570 DVSS.n3424 DVSS.n3423 0.4505
R59571 DVSS.n2184 DVSS.n2183 0.4505
R59572 DVSS.n3419 DVSS.n3418 0.4505
R59573 DVSS.n3417 DVSS.n2186 0.4505
R59574 DVSS.n3416 DVSS.n3415 0.4505
R59575 DVSS.n2188 DVSS.n2187 0.4505
R59576 DVSS.n3411 DVSS.n3410 0.4505
R59577 DVSS.n3409 DVSS.n2190 0.4505
R59578 DVSS.n3408 DVSS.n3407 0.4505
R59579 DVSS.n2192 DVSS.n2191 0.4505
R59580 DVSS.n3403 DVSS.n3402 0.4505
R59581 DVSS.n3401 DVSS.n2194 0.4505
R59582 DVSS.n3400 DVSS.n3399 0.4505
R59583 DVSS.n2196 DVSS.n2195 0.4505
R59584 DVSS.n3395 DVSS.n3394 0.4505
R59585 DVSS.n3393 DVSS.n2198 0.4505
R59586 DVSS.n3392 DVSS.n3391 0.4505
R59587 DVSS.n2200 DVSS.n2199 0.4505
R59588 DVSS.n3387 DVSS.n3386 0.4505
R59589 DVSS.n3385 DVSS.n2202 0.4505
R59590 DVSS.n3384 DVSS.n3383 0.4505
R59591 DVSS.n2204 DVSS.n2203 0.4505
R59592 DVSS.n3379 DVSS.n3378 0.4505
R59593 DVSS.n3377 DVSS.n2206 0.4505
R59594 DVSS.n3376 DVSS.n3375 0.4505
R59595 DVSS.n2208 DVSS.n2207 0.4505
R59596 DVSS.n3371 DVSS.n3370 0.4505
R59597 DVSS.n3369 DVSS.n2210 0.4505
R59598 DVSS.n3368 DVSS.n3367 0.4505
R59599 DVSS.n2212 DVSS.n2211 0.4505
R59600 DVSS.n3363 DVSS.n3362 0.4505
R59601 DVSS.n3361 DVSS.n2214 0.4505
R59602 DVSS.n3360 DVSS.n3359 0.4505
R59603 DVSS.n2216 DVSS.n2215 0.4505
R59604 DVSS.n3355 DVSS.n3354 0.4505
R59605 DVSS.n3353 DVSS.n2218 0.4505
R59606 DVSS.n3352 DVSS.n3351 0.4505
R59607 DVSS.n2220 DVSS.n2219 0.4505
R59608 DVSS.n3347 DVSS.n3346 0.4505
R59609 DVSS.n3345 DVSS.n2222 0.4505
R59610 DVSS.n3344 DVSS.n3343 0.4505
R59611 DVSS.n2224 DVSS.n2223 0.4505
R59612 DVSS.n3339 DVSS.n3338 0.4505
R59613 DVSS.n3337 DVSS.n2226 0.4505
R59614 DVSS.n3336 DVSS.n3335 0.4505
R59615 DVSS.n2228 DVSS.n2227 0.4505
R59616 DVSS.n3331 DVSS.n3330 0.4505
R59617 DVSS.n3329 DVSS.n2230 0.4505
R59618 DVSS.n2276 DVSS.n2275 0.4505
R59619 DVSS.n3790 DVSS.n1931 0.4505
R59620 DVSS.n4748 DVSS.n4747 0.4505
R59621 DVSS.n3528 DVSS 0.435162
R59622 DVSS DVSS.n3530 0.435162
R59623 DVSS.n5659 DVSS.n5658 0.423402
R59624 DVSS.n4929 DVSS.n1791 0.400952
R59625 DVSS.n4970 DVSS.n4967 0.400952
R59626 DVSS.n4931 DVSS.n1793 0.400952
R59627 DVSS.n4983 DVSS.n4982 0.400952
R59628 DVSS.n4953 DVSS.n4952 0.400952
R59629 DVSS.n4976 DVSS.n4975 0.400952
R59630 DVSS.n3041 DVSS.n3040 0.40055
R59631 DVSS.n3028 DVSS.n3027 0.40055
R59632 DVSS.n5679 DVSS.n5678 0.400345
R59633 DVSS.n5662 DVSS.n5661 0.371929
R59634 DVSS.n5672 DVSS.n1272 0.371929
R59635 DVSS.n3534 DVSS 0.367475
R59636 DVSS.n3524 DVSS 0.367475
R59637 DVSS.n4747 DVSS.n4746 0.355295
R59638 DVSS.n3294 DVSS.n3293 0.355011
R59639 DVSS.n2244 DVSS.n2138 0.355011
R59640 DVSS.n3096 DVSS.n3095 0.354754
R59641 DVSS.n3503 DVSS.n3502 0.354754
R59642 DVSS.n3537 DVSS.n3534 0.352976
R59643 DVSS.n3524 DVSS.n3522 0.352976
R59644 DVSS.n3791 DVSS.n3790 0.349418
R59645 DVSS.n2119 DVSS 0.34295
R59646 DVSS.n5605 DVSS.n5599 0.3326
R59647 DVSS.n5588 DVSS.n1330 0.3326
R59648 DVSS.n5653 DVSS.n5652 0.3326
R59649 DVSS.n1313 DVSS.n1312 0.3326
R59650 DVSS.n2747 DVSS.n2534 0.329772
R59651 DVSS.n3809 DVSS.n3804 0.329604
R59652 DVSS.n1286 DVSS.t17 0.3281
R59653 DVSS.n1286 DVSS.t23 0.3281
R59654 DVSS.n1289 DVSS.t13 0.3281
R59655 DVSS.n1289 DVSS.t19 0.3281
R59656 DVSS.n1262 DVSS.t21 0.3281
R59657 DVSS.n1262 DVSS.t198 0.3281
R59658 DVSS.n1264 DVSS.t196 0.3281
R59659 DVSS.n1264 DVSS.t192 0.3281
R59660 DVSS.n1266 DVSS.t190 0.3281
R59661 DVSS.n1266 DVSS.t194 0.3281
R59662 DVSS.n5347 DVSS.n1379 0.321929
R59663 DVSS.n5167 DVSS.n1601 0.321929
R59664 DVSS.n4367 DVSS.n1803 0.321929
R59665 DVSS.n4431 DVSS.n4430 0.321929
R59666 DVSS.n2118 DVSS.t25 0.312926
R59667 DVSS.n2118 DVSS.t27 0.312926
R59668 DVSS.n3519 DVSS.t26 0.312926
R59669 DVSS.n3069 DVSS.t28 0.312926
R59670 DVSS.n2111 DVSS.t27 0.312926
R59671 DVSS.n2111 DVSS.t28 0.312926
R59672 DVSS.n3523 DVSS.t26 0.312926
R59673 DVSS.n3523 DVSS.t25 0.312926
R59674 DVSS.n5697 DVSS.n5696 0.3092
R59675 DVSS.n5695 DVSS.n5694 0.3092
R59676 DVSS.n4972 DVSS.n4971 0.3092
R59677 DVSS.n4968 DVSS.n1756 0.3092
R59678 DVSS.n5704 DVSS.n5703 0.3092
R59679 DVSS.n5701 DVSS.n1228 0.3092
R59680 DVSS.n4951 DVSS.n4950 0.3092
R59681 DVSS.n4947 DVSS.n4946 0.3092
R59682 DVSS.n5719 DVSS.n5718 0.3092
R59683 DVSS.n5722 DVSS.n5721 0.3092
R59684 DVSS.n5716 DVSS.n5715 0.3092
R59685 DVSS.n5724 DVSS.n1230 0.3092
R59686 DVSS.n3039 DVSS.n1771 0.30245
R59687 DVSS.n3031 DVSS.n3030 0.30245
R59688 DVSS.n3095 DVSS.n3094 0.292137
R59689 DVSS.n5713 DVSS.n218 0.273435
R59690 DVSS.n5698 DVSS.n215 0.273435
R59691 DVSS.n6427 DVSS.n217 0.273435
R59692 DVSS.n6429 DVSS.n214 0.273435
R59693 DVSS.n6426 DVSS.n219 0.273435
R59694 DVSS.n6430 DVSS.n213 0.273435
R59695 DVSS.n2383 DVSS.n1279 0.258595
R59696 DVSS.n3504 DVSS.n2142 0.252283
R59697 DVSS.n3515 DVSS.n3514 0.252283
R59698 DVSS.n3076 DVSS.n2367 0.247099
R59699 DVSS.n3501 DVSS.n3500 0.231338
R59700 DVSS.n2249 DVSS.n2248 0.231338
R59701 DVSS.n3100 DVSS.n2365 0.231338
R59702 DVSS.n3299 DVSS.n3298 0.231338
R59703 DVSS DVSS.n3527 0.222172
R59704 DVSS.n3531 DVSS 0.222172
R59705 DVSS.n5606 DVSS.n5605 0.2201
R59706 DVSS.n5606 DVSS.n1327 0.2201
R59707 DVSS.n5622 DVSS.n1327 0.2201
R59708 DVSS.n5623 DVSS.n5622 0.2201
R59709 DVSS.n5623 DVSS.n1322 0.2201
R59710 DVSS.n5639 DVSS.n1322 0.2201
R59711 DVSS.n5640 DVSS.n5639 0.2201
R59712 DVSS.n5640 DVSS.n1241 0.2201
R59713 DVSS.n5696 DVSS.n1241 0.2201
R59714 DVSS.n5694 DVSS.n1229 0.2201
R59715 DVSS.n1229 DVSS.n1227 0.2201
R59716 DVSS.n1227 DVSS.n1226 0.2201
R59717 DVSS.n1226 DVSS.n1216 0.2201
R59718 DVSS.n1216 DVSS.n1214 0.2201
R59719 DVSS.n1214 DVSS.n1213 0.2201
R59720 DVSS.n1213 DVSS.n1202 0.2201
R59721 DVSS.n1202 DVSS.n1197 0.2201
R59722 DVSS.n6068 DVSS.n1197 0.2201
R59723 DVSS.n5782 DVSS.n1138 0.2201
R59724 DVSS.n1138 DVSS.n1095 0.2201
R59725 DVSS.n6123 DVSS.n1095 0.2201
R59726 DVSS.n5611 DVSS.n1330 0.2201
R59727 DVSS.n5612 DVSS.n5611 0.2201
R59728 DVSS.n5612 DVSS.n1326 0.2201
R59729 DVSS.n5628 DVSS.n1326 0.2201
R59730 DVSS.n5629 DVSS.n5628 0.2201
R59731 DVSS.n5629 DVSS.n1323 0.2201
R59732 DVSS.n1323 DVSS.n1242 0.2201
R59733 DVSS.n5705 DVSS.n1242 0.2201
R59734 DVSS.n5705 DVSS.n5704 0.2201
R59735 DVSS.n5731 DVSS.n1228 0.2201
R59736 DVSS.n5732 DVSS.n5731 0.2201
R59737 DVSS.n5732 DVSS.n1215 0.2201
R59738 DVSS.n5748 DVSS.n1215 0.2201
R59739 DVSS.n5749 DVSS.n5748 0.2201
R59740 DVSS.n5749 DVSS.n1201 0.2201
R59741 DVSS.n5768 DVSS.n1201 0.2201
R59742 DVSS.n5769 DVSS.n5768 0.2201
R59743 DVSS.n5769 DVSS.n1198 0.2201
R59744 DVSS.n6113 DVSS.n1137 0.2201
R59745 DVSS.n6114 DVSS.n6113 0.2201
R59746 DVSS.n6114 DVSS.n1133 0.2201
R59747 DVSS.n5652 DVSS.n5651 0.2201
R59748 DVSS.n5651 DVSS.n5650 0.2201
R59749 DVSS.n5650 DVSS.n5649 0.2201
R59750 DVSS.n5649 DVSS.n5648 0.2201
R59751 DVSS.n5648 DVSS.n5647 0.2201
R59752 DVSS.n5647 DVSS.n5646 0.2201
R59753 DVSS.n5646 DVSS.n5645 0.2201
R59754 DVSS.n5645 DVSS.n1235 0.2201
R59755 DVSS.n5718 DVSS.n1235 0.2201
R59756 DVSS.n5722 DVSS.n1219 0.2201
R59757 DVSS.n5738 DVSS.n1219 0.2201
R59758 DVSS.n5739 DVSS.n5738 0.2201
R59759 DVSS.n5739 DVSS.n1206 0.2201
R59760 DVSS.n5755 DVSS.n1206 0.2201
R59761 DVSS.n5756 DVSS.n5755 0.2201
R59762 DVSS.n5756 DVSS.n1203 0.2201
R59763 DVSS.n5759 DVSS.n1203 0.2201
R59764 DVSS.n5759 DVSS.n1151 0.2201
R59765 DVSS.n6104 DVSS.n1139 0.2201
R59766 DVSS.n1139 DVSS.n426 0.2201
R59767 DVSS.n6234 DVSS.n426 0.2201
R59768 DVSS.n1314 DVSS.n1313 0.2201
R59769 DVSS.n1315 DVSS.n1314 0.2201
R59770 DVSS.n1316 DVSS.n1315 0.2201
R59771 DVSS.n1317 DVSS.n1316 0.2201
R59772 DVSS.n1318 DVSS.n1317 0.2201
R59773 DVSS.n1319 DVSS.n1318 0.2201
R59774 DVSS.n1319 DVSS.n1237 0.2201
R59775 DVSS.n5711 DVSS.n1237 0.2201
R59776 DVSS.n5716 DVSS.n5711 0.2201
R59777 DVSS.n5725 DVSS.n5724 0.2201
R59778 DVSS.n5725 DVSS.n1217 0.2201
R59779 DVSS.n5741 DVSS.n1217 0.2201
R59780 DVSS.n5742 DVSS.n5741 0.2201
R59781 DVSS.n5742 DVSS.n1204 0.2201
R59782 DVSS.n5758 DVSS.n1204 0.2201
R59783 DVSS.n5762 DVSS.n5758 0.2201
R59784 DVSS.n5762 DVSS.n5761 0.2201
R59785 DVSS.n5761 DVSS.n1166 0.2201
R59786 DVSS.n6107 DVSS.n6106 0.2201
R59787 DVSS.n6107 DVSS.n424 0.2201
R59788 DVSS.n6236 DVSS.n424 0.2201
R59789 DVSS.n5341 DVSS.n5303 0.214786
R59790 DVSS.n5323 DVSS.n5321 0.214786
R59791 DVSS.n5324 DVSS.n5320 0.214786
R59792 DVSS.n5325 DVSS.n5319 0.214786
R59793 DVSS.n5318 DVSS.n5316 0.214786
R59794 DVSS.n5329 DVSS.n5315 0.214786
R59795 DVSS.n5330 DVSS.n5314 0.214786
R59796 DVSS.n5331 DVSS.n5313 0.214786
R59797 DVSS.n5312 DVSS.n5310 0.214786
R59798 DVSS.n5335 DVSS.n5309 0.214786
R59799 DVSS.n5336 DVSS.n5308 0.214786
R59800 DVSS.n5337 DVSS.n5307 0.214786
R59801 DVSS.n5306 DVSS.n5304 0.214786
R59802 DVSS.n2055 DVSS.n2054 0.214786
R59803 DVSS.n4452 DVSS.n4451 0.214786
R59804 DVSS.n4453 DVSS.n2053 0.214786
R59805 DVSS.n4455 DVSS.n4454 0.214786
R59806 DVSS.n2051 DVSS.n2050 0.214786
R59807 DVSS.n4460 DVSS.n4459 0.214786
R59808 DVSS.n4461 DVSS.n2049 0.214786
R59809 DVSS.n4463 DVSS.n4462 0.214786
R59810 DVSS.n2047 DVSS.n2046 0.214786
R59811 DVSS.n4468 DVSS.n4467 0.214786
R59812 DVSS.n4469 DVSS.n2045 0.214786
R59813 DVSS.n4471 DVSS.n4470 0.214786
R59814 DVSS.n2043 DVSS.n2042 0.214786
R59815 DVSS.n4476 DVSS.n4475 0.214786
R59816 DVSS.n4477 DVSS.n2041 0.214786
R59817 DVSS.n4624 DVSS.n4478 0.214786
R59818 DVSS.n4623 DVSS.n4479 0.214786
R59819 DVSS.n4622 DVSS.n4480 0.214786
R59820 DVSS.n4621 DVSS.n4481 0.214786
R59821 DVSS.n4484 DVSS.n4482 0.214786
R59822 DVSS.n4617 DVSS.n4485 0.214786
R59823 DVSS.n4616 DVSS.n4486 0.214786
R59824 DVSS.n4615 DVSS.n4487 0.214786
R59825 DVSS.n4490 DVSS.n4488 0.214786
R59826 DVSS.n4611 DVSS.n4491 0.214786
R59827 DVSS.n4610 DVSS.n4492 0.214786
R59828 DVSS.n4609 DVSS.n4493 0.214786
R59829 DVSS.n4496 DVSS.n4494 0.214786
R59830 DVSS.n4605 DVSS.n4497 0.214786
R59831 DVSS.n4604 DVSS.n4498 0.214786
R59832 DVSS.n4603 DVSS.n4499 0.214786
R59833 DVSS.n4502 DVSS.n4500 0.214786
R59834 DVSS.n4599 DVSS.n4503 0.214786
R59835 DVSS.n4598 DVSS.n4504 0.214786
R59836 DVSS.n4552 DVSS.n4505 0.214786
R59837 DVSS.n4592 DVSS.n4553 0.214786
R59838 DVSS.n4591 DVSS.n4554 0.214786
R59839 DVSS.n4590 DVSS.n4555 0.214786
R59840 DVSS.n4558 DVSS.n4556 0.214786
R59841 DVSS.n4586 DVSS.n4559 0.214786
R59842 DVSS.n4585 DVSS.n4560 0.214786
R59843 DVSS.n4584 DVSS.n4561 0.214786
R59844 DVSS.n4564 DVSS.n4562 0.214786
R59845 DVSS.n4580 DVSS.n4565 0.214786
R59846 DVSS.n4579 DVSS.n4566 0.214786
R59847 DVSS.n4578 DVSS.n4567 0.214786
R59848 DVSS.n4570 DVSS.n4568 0.214786
R59849 DVSS.n4574 DVSS.n4571 0.214786
R59850 DVSS.n4573 DVSS.n4572 0.214786
R59851 DVSS.n1567 DVSS.n1566 0.214786
R59852 DVSS.n5268 DVSS.n5267 0.214786
R59853 DVSS.n5269 DVSS.n1565 0.214786
R59854 DVSS.n5271 DVSS.n5270 0.214786
R59855 DVSS.n1563 DVSS.n1562 0.214786
R59856 DVSS.n5276 DVSS.n5275 0.214786
R59857 DVSS.n5277 DVSS.n1561 0.214786
R59858 DVSS.n5279 DVSS.n5278 0.214786
R59859 DVSS.n1559 DVSS.n1558 0.214786
R59860 DVSS.n5284 DVSS.n5283 0.214786
R59861 DVSS.n5285 DVSS.n1557 0.214786
R59862 DVSS.n5287 DVSS.n5286 0.214786
R59863 DVSS.n1555 DVSS.n1554 0.214786
R59864 DVSS.n5292 DVSS.n5291 0.214786
R59865 DVSS.n5293 DVSS.n1553 0.214786
R59866 DVSS.n5295 DVSS.n5294 0.214786
R59867 DVSS.n1551 DVSS.n1550 0.214786
R59868 DVSS.n5300 DVSS.n5299 0.214786
R59869 DVSS.n5301 DVSS.n1549 0.214786
R59870 DVSS.n5342 DVSS.n5302 0.214786
R59871 DVSS.n5324 DVSS.n5317 0.214786
R59872 DVSS.n5326 DVSS.n5325 0.214786
R59873 DVSS.n5327 DVSS.n5316 0.214786
R59874 DVSS.n5329 DVSS.n5328 0.214786
R59875 DVSS.n5330 DVSS.n5311 0.214786
R59876 DVSS.n5332 DVSS.n5331 0.214786
R59877 DVSS.n5333 DVSS.n5310 0.214786
R59878 DVSS.n5335 DVSS.n5334 0.214786
R59879 DVSS.n5336 DVSS.n5305 0.214786
R59880 DVSS.n5338 DVSS.n5337 0.214786
R59881 DVSS.n5339 DVSS.n5304 0.214786
R59882 DVSS.n5341 DVSS.n5340 0.214786
R59883 DVSS.n4432 DVSS.n2056 0.214786
R59884 DVSS.n4449 DVSS.n2055 0.214786
R59885 DVSS.n4451 DVSS.n4450 0.214786
R59886 DVSS.n2053 DVSS.n2052 0.214786
R59887 DVSS.n4456 DVSS.n4455 0.214786
R59888 DVSS.n4457 DVSS.n2051 0.214786
R59889 DVSS.n4459 DVSS.n4458 0.214786
R59890 DVSS.n2049 DVSS.n2048 0.214786
R59891 DVSS.n4464 DVSS.n4463 0.214786
R59892 DVSS.n4465 DVSS.n2047 0.214786
R59893 DVSS.n4467 DVSS.n4466 0.214786
R59894 DVSS.n2045 DVSS.n2044 0.214786
R59895 DVSS.n4472 DVSS.n4471 0.214786
R59896 DVSS.n4473 DVSS.n2043 0.214786
R59897 DVSS.n4475 DVSS.n4474 0.214786
R59898 DVSS.n2041 DVSS.n2040 0.214786
R59899 DVSS.n4625 DVSS.n4624 0.214786
R59900 DVSS.n4623 DVSS.n2027 0.214786
R59901 DVSS.n4622 DVSS.n2028 0.214786
R59902 DVSS.n4621 DVSS.n4620 0.214786
R59903 DVSS.n4619 DVSS.n4482 0.214786
R59904 DVSS.n4618 DVSS.n4617 0.214786
R59905 DVSS.n4616 DVSS.n4483 0.214786
R59906 DVSS.n4615 DVSS.n4614 0.214786
R59907 DVSS.n4613 DVSS.n4488 0.214786
R59908 DVSS.n4612 DVSS.n4611 0.214786
R59909 DVSS.n4610 DVSS.n4489 0.214786
R59910 DVSS.n4609 DVSS.n4608 0.214786
R59911 DVSS.n4607 DVSS.n4494 0.214786
R59912 DVSS.n4606 DVSS.n4605 0.214786
R59913 DVSS.n4604 DVSS.n4495 0.214786
R59914 DVSS.n4603 DVSS.n4602 0.214786
R59915 DVSS.n4601 DVSS.n4500 0.214786
R59916 DVSS.n4600 DVSS.n4599 0.214786
R59917 DVSS.n4598 DVSS.n4597 0.214786
R59918 DVSS.n4550 DVSS.n4505 0.214786
R59919 DVSS.n4593 DVSS.n4592 0.214786
R59920 DVSS.n4591 DVSS.n4551 0.214786
R59921 DVSS.n4590 DVSS.n4589 0.214786
R59922 DVSS.n4588 DVSS.n4556 0.214786
R59923 DVSS.n4587 DVSS.n4586 0.214786
R59924 DVSS.n4585 DVSS.n4557 0.214786
R59925 DVSS.n4584 DVSS.n4583 0.214786
R59926 DVSS.n4582 DVSS.n4562 0.214786
R59927 DVSS.n4581 DVSS.n4580 0.214786
R59928 DVSS.n4579 DVSS.n4563 0.214786
R59929 DVSS.n4578 DVSS.n4577 0.214786
R59930 DVSS.n4576 DVSS.n4568 0.214786
R59931 DVSS.n4575 DVSS.n4574 0.214786
R59932 DVSS.n4573 DVSS.n4569 0.214786
R59933 DVSS.n1568 DVSS.n1567 0.214786
R59934 DVSS.n5267 DVSS.n5266 0.214786
R59935 DVSS.n5264 DVSS.n1565 0.214786
R59936 DVSS.n5272 DVSS.n5271 0.214786
R59937 DVSS.n5273 DVSS.n1563 0.214786
R59938 DVSS.n5275 DVSS.n5274 0.214786
R59939 DVSS.n1561 DVSS.n1560 0.214786
R59940 DVSS.n5280 DVSS.n5279 0.214786
R59941 DVSS.n5281 DVSS.n1559 0.214786
R59942 DVSS.n5283 DVSS.n5282 0.214786
R59943 DVSS.n1557 DVSS.n1556 0.214786
R59944 DVSS.n5288 DVSS.n5287 0.214786
R59945 DVSS.n5289 DVSS.n1555 0.214786
R59946 DVSS.n5291 DVSS.n5290 0.214786
R59947 DVSS.n1553 DVSS.n1552 0.214786
R59948 DVSS.n5296 DVSS.n5295 0.214786
R59949 DVSS.n5297 DVSS.n1551 0.214786
R59950 DVSS.n5299 DVSS.n5298 0.214786
R59951 DVSS.n1549 DVSS.n1527 0.214786
R59952 DVSS.n5343 DVSS.n5342 0.214786
R59953 DVSS.n1052 DVSS.n1047 0.214786
R59954 DVSS.n1053 DVSS.n1046 0.214786
R59955 DVSS.n1054 DVSS.n1045 0.214786
R59956 DVSS.n1044 DVSS.n1042 0.214786
R59957 DVSS.n1058 DVSS.n1041 0.214786
R59958 DVSS.n1059 DVSS.n1040 0.214786
R59959 DVSS.n1060 DVSS.n1039 0.214786
R59960 DVSS.n1038 DVSS.n1036 0.214786
R59961 DVSS.n1064 DVSS.n1035 0.214786
R59962 DVSS.n1065 DVSS.n1034 0.214786
R59963 DVSS.n1066 DVSS.n1033 0.214786
R59964 DVSS.n1084 DVSS.n1070 0.214786
R59965 DVSS.n753 DVSS.n397 0.214786
R59966 DVSS.n752 DVSS.n405 0.214786
R59967 DVSS.n751 DVSS.n419 0.214786
R59968 DVSS.n661 DVSS.n659 0.214786
R59969 DVSS.n747 DVSS.n662 0.214786
R59970 DVSS.n746 DVSS.n663 0.214786
R59971 DVSS.n745 DVSS.n664 0.214786
R59972 DVSS.n667 DVSS.n665 0.214786
R59973 DVSS.n741 DVSS.n668 0.214786
R59974 DVSS.n740 DVSS.n669 0.214786
R59975 DVSS.n739 DVSS.n670 0.214786
R59976 DVSS.n673 DVSS.n671 0.214786
R59977 DVSS.n735 DVSS.n674 0.214786
R59978 DVSS.n734 DVSS.n675 0.214786
R59979 DVSS.n733 DVSS.n676 0.214786
R59980 DVSS.n679 DVSS.n677 0.214786
R59981 DVSS.n729 DVSS.n680 0.214786
R59982 DVSS.n728 DVSS.n442 0.214786
R59983 DVSS.n727 DVSS.n428 0.214786
R59984 DVSS.n681 DVSS.n435 0.214786
R59985 DVSS.n723 DVSS.n683 0.214786
R59986 DVSS.n722 DVSS.n684 0.214786
R59987 DVSS.n721 DVSS.n685 0.214786
R59988 DVSS.n718 DVSS.n717 0.214786
R59989 DVSS.n715 DVSS.n714 0.214786
R59990 DVSS.n687 DVSS.n686 0.214786
R59991 DVSS.n710 DVSS.n689 0.214786
R59992 DVSS.n709 DVSS.n690 0.214786
R59993 DVSS.n708 DVSS.n691 0.214786
R59994 DVSS.n694 DVSS.n692 0.214786
R59995 DVSS.n704 DVSS.n695 0.214786
R59996 DVSS.n703 DVSS.n696 0.214786
R59997 DVSS.n702 DVSS.n697 0.214786
R59998 DVSS.n699 DVSS.n698 0.214786
R59999 DVSS.n516 DVSS.n511 0.214786
R60000 DVSS.n6188 DVSS.n6187 0.214786
R60001 DVSS.n517 DVSS.n466 0.214786
R60002 DVSS.n6183 DVSS.n475 0.214786
R60003 DVSS.n6182 DVSS.n520 0.214786
R60004 DVSS.n6181 DVSS.n521 0.214786
R60005 DVSS.n524 DVSS.n522 0.214786
R60006 DVSS.n6177 DVSS.n525 0.214786
R60007 DVSS.n6176 DVSS.n526 0.214786
R60008 DVSS.n6175 DVSS.n527 0.214786
R60009 DVSS.n530 DVSS.n528 0.214786
R60010 DVSS.n6171 DVSS.n531 0.214786
R60011 DVSS.n6170 DVSS.n532 0.214786
R60012 DVSS.n6169 DVSS.n533 0.214786
R60013 DVSS.n6165 DVSS.n998 0.214786
R60014 DVSS.n6164 DVSS.n999 0.214786
R60015 DVSS.n6163 DVSS.n1000 0.214786
R60016 DVSS.n1003 DVSS.n1001 0.214786
R60017 DVSS.n6159 DVSS.n1004 0.214786
R60018 DVSS.n6158 DVSS.n1005 0.214786
R60019 DVSS.n6157 DVSS.n1006 0.214786
R60020 DVSS.n1009 DVSS.n1007 0.214786
R60021 DVSS.n6153 DVSS.n1010 0.214786
R60022 DVSS.n6152 DVSS.n1011 0.214786
R60023 DVSS.n6151 DVSS.n1012 0.214786
R60024 DVSS.n1015 DVSS.n1013 0.214786
R60025 DVSS.n6147 DVSS.n1016 0.214786
R60026 DVSS.n6146 DVSS.n1017 0.214786
R60027 DVSS.n6145 DVSS.n1018 0.214786
R60028 DVSS.n1021 DVSS.n1019 0.214786
R60029 DVSS.n6141 DVSS.n1022 0.214786
R60030 DVSS.n6140 DVSS.n1023 0.214786
R60031 DVSS.n6139 DVSS.n1024 0.214786
R60032 DVSS.n1027 DVSS.n1025 0.214786
R60033 DVSS.n6135 DVSS.n1028 0.214786
R60034 DVSS.n6134 DVSS.n1029 0.214786
R60035 DVSS.n1050 DVSS.n1049 0.214786
R60036 DVSS.n1052 DVSS.n1051 0.214786
R60037 DVSS.n1053 DVSS.n1043 0.214786
R60038 DVSS.n1055 DVSS.n1054 0.214786
R60039 DVSS.n1056 DVSS.n1042 0.214786
R60040 DVSS.n1058 DVSS.n1057 0.214786
R60041 DVSS.n1059 DVSS.n1037 0.214786
R60042 DVSS.n1061 DVSS.n1060 0.214786
R60043 DVSS.n1062 DVSS.n1036 0.214786
R60044 DVSS.n1064 DVSS.n1063 0.214786
R60045 DVSS.n1065 DVSS.n1032 0.214786
R60046 DVSS.n1067 DVSS.n1066 0.214786
R60047 DVSS.n1070 DVSS.n1069 0.214786
R60048 DVSS.n754 DVSS.n753 0.214786
R60049 DVSS.n752 DVSS.n590 0.214786
R60050 DVSS.n751 DVSS.n750 0.214786
R60051 DVSS.n749 DVSS.n659 0.214786
R60052 DVSS.n748 DVSS.n747 0.214786
R60053 DVSS.n746 DVSS.n660 0.214786
R60054 DVSS.n745 DVSS.n744 0.214786
R60055 DVSS.n743 DVSS.n665 0.214786
R60056 DVSS.n742 DVSS.n741 0.214786
R60057 DVSS.n740 DVSS.n666 0.214786
R60058 DVSS.n739 DVSS.n738 0.214786
R60059 DVSS.n737 DVSS.n671 0.214786
R60060 DVSS.n736 DVSS.n735 0.214786
R60061 DVSS.n734 DVSS.n672 0.214786
R60062 DVSS.n733 DVSS.n732 0.214786
R60063 DVSS.n731 DVSS.n677 0.214786
R60064 DVSS.n730 DVSS.n729 0.214786
R60065 DVSS.n728 DVSS.n678 0.214786
R60066 DVSS.n727 DVSS.n726 0.214786
R60067 DVSS.n725 DVSS.n681 0.214786
R60068 DVSS.n724 DVSS.n723 0.214786
R60069 DVSS.n722 DVSS.n682 0.214786
R60070 DVSS.n721 DVSS.n720 0.214786
R60071 DVSS.n719 DVSS.n718 0.214786
R60072 DVSS.n714 DVSS.n713 0.214786
R60073 DVSS.n712 DVSS.n687 0.214786
R60074 DVSS.n711 DVSS.n710 0.214786
R60075 DVSS.n709 DVSS.n688 0.214786
R60076 DVSS.n708 DVSS.n707 0.214786
R60077 DVSS.n706 DVSS.n692 0.214786
R60078 DVSS.n705 DVSS.n704 0.214786
R60079 DVSS.n703 DVSS.n693 0.214786
R60080 DVSS.n702 DVSS.n701 0.214786
R60081 DVSS.n700 DVSS.n699 0.214786
R60082 DVSS.n518 DVSS.n516 0.214786
R60083 DVSS.n6187 DVSS.n6186 0.214786
R60084 DVSS.n6185 DVSS.n517 0.214786
R60085 DVSS.n6184 DVSS.n6183 0.214786
R60086 DVSS.n6182 DVSS.n519 0.214786
R60087 DVSS.n6181 DVSS.n6180 0.214786
R60088 DVSS.n6179 DVSS.n522 0.214786
R60089 DVSS.n6178 DVSS.n6177 0.214786
R60090 DVSS.n6176 DVSS.n523 0.214786
R60091 DVSS.n6175 DVSS.n6174 0.214786
R60092 DVSS.n6173 DVSS.n528 0.214786
R60093 DVSS.n6172 DVSS.n6171 0.214786
R60094 DVSS.n6170 DVSS.n529 0.214786
R60095 DVSS.n6169 DVSS.n6168 0.214786
R60096 DVSS.n6166 DVSS.n6165 0.214786
R60097 DVSS.n6164 DVSS.n534 0.214786
R60098 DVSS.n6163 DVSS.n6162 0.214786
R60099 DVSS.n6161 DVSS.n1001 0.214786
R60100 DVSS.n6160 DVSS.n6159 0.214786
R60101 DVSS.n6158 DVSS.n1002 0.214786
R60102 DVSS.n6157 DVSS.n6156 0.214786
R60103 DVSS.n6155 DVSS.n1007 0.214786
R60104 DVSS.n6154 DVSS.n6153 0.214786
R60105 DVSS.n6152 DVSS.n1008 0.214786
R60106 DVSS.n6151 DVSS.n6150 0.214786
R60107 DVSS.n6149 DVSS.n1013 0.214786
R60108 DVSS.n6148 DVSS.n6147 0.214786
R60109 DVSS.n6146 DVSS.n1014 0.214786
R60110 DVSS.n6145 DVSS.n6144 0.214786
R60111 DVSS.n6143 DVSS.n1019 0.214786
R60112 DVSS.n6142 DVSS.n6141 0.214786
R60113 DVSS.n6140 DVSS.n1020 0.214786
R60114 DVSS.n6139 DVSS.n6138 0.214786
R60115 DVSS.n6137 DVSS.n1025 0.214786
R60116 DVSS.n6136 DVSS.n6135 0.214786
R60117 DVSS.n6134 DVSS.n1026 0.214786
R60118 DVSS.n6133 DVSS.n1030 0.214786
R60119 DVSS.n6133 DVSS.n6132 0.214786
R60120 DVSS.n586 DVSS.n65 0.214786
R60121 DVSS.n759 DVSS.n50 0.214786
R60122 DVSS.n760 DVSS.n60 0.214786
R60123 DVSS.n762 DVSS.n761 0.214786
R60124 DVSS.n584 DVSS.n583 0.214786
R60125 DVSS.n767 DVSS.n766 0.214786
R60126 DVSS.n768 DVSS.n582 0.214786
R60127 DVSS.n770 DVSS.n769 0.214786
R60128 DVSS.n580 DVSS.n579 0.214786
R60129 DVSS.n775 DVSS.n774 0.214786
R60130 DVSS.n776 DVSS.n578 0.214786
R60131 DVSS.n778 DVSS.n777 0.214786
R60132 DVSS.n576 DVSS.n575 0.214786
R60133 DVSS.n783 DVSS.n782 0.214786
R60134 DVSS.n784 DVSS.n574 0.214786
R60135 DVSS.n787 DVSS.n786 0.214786
R60136 DVSS.n785 DVSS.n572 0.214786
R60137 DVSS.n791 DVSS.n80 0.214786
R60138 DVSS.n792 DVSS.n88 0.214786
R60139 DVSS.n793 DVSS.n102 0.214786
R60140 DVSS.n570 DVSS.n569 0.214786
R60141 DVSS.n799 DVSS.n798 0.214786
R60142 DVSS.n800 DVSS.n568 0.214786
R60143 DVSS.n802 DVSS.n801 0.214786
R60144 DVSS.n835 DVSS.n804 0.214786
R60145 DVSS.n834 DVSS.n805 0.214786
R60146 DVSS.n833 DVSS.n806 0.214786
R60147 DVSS.n809 DVSS.n807 0.214786
R60148 DVSS.n829 DVSS.n810 0.214786
R60149 DVSS.n828 DVSS.n811 0.214786
R60150 DVSS.n827 DVSS.n812 0.214786
R60151 DVSS.n815 DVSS.n813 0.214786
R60152 DVSS.n823 DVSS.n816 0.214786
R60153 DVSS.n822 DVSS.n817 0.214786
R60154 DVSS.n821 DVSS.n285 0.214786
R60155 DVSS.n818 DVSS.n299 0.214786
R60156 DVSS.n325 DVSS.n321 0.214786
R60157 DVSS.n6366 DVSS.n6365 0.214786
R60158 DVSS.n326 DVSS.n324 0.214786
R60159 DVSS.n6361 DVSS.n329 0.214786
R60160 DVSS.n6360 DVSS.n330 0.214786
R60161 DVSS.n6359 DVSS.n331 0.214786
R60162 DVSS.n334 DVSS.n332 0.214786
R60163 DVSS.n6355 DVSS.n335 0.214786
R60164 DVSS.n6354 DVSS.n336 0.214786
R60165 DVSS.n6353 DVSS.n337 0.214786
R60166 DVSS.n340 DVSS.n338 0.214786
R60167 DVSS.n6349 DVSS.n341 0.214786
R60168 DVSS.n6347 DVSS.n344 0.214786
R60169 DVSS.n347 DVSS.n345 0.214786
R60170 DVSS.n6343 DVSS.n348 0.214786
R60171 DVSS.n6342 DVSS.n349 0.214786
R60172 DVSS.n6341 DVSS.n350 0.214786
R60173 DVSS.n353 DVSS.n351 0.214786
R60174 DVSS.n6337 DVSS.n6298 0.214786
R60175 DVSS.n6336 DVSS.n6299 0.214786
R60176 DVSS.n6335 DVSS.n6300 0.214786
R60177 DVSS.n6303 DVSS.n6301 0.214786
R60178 DVSS.n6331 DVSS.n6304 0.214786
R60179 DVSS.n6330 DVSS.n6305 0.214786
R60180 DVSS.n6329 DVSS.n6306 0.214786
R60181 DVSS.n6309 DVSS.n6307 0.214786
R60182 DVSS.n6325 DVSS.n6310 0.214786
R60183 DVSS.n6324 DVSS.n6311 0.214786
R60184 DVSS.n6323 DVSS.n6312 0.214786
R60185 DVSS.n6315 DVSS.n6313 0.214786
R60186 DVSS.n6319 DVSS.n6316 0.214786
R60187 DVSS.n6318 DVSS.n6317 0.214786
R60188 DVSS.n19 DVSS.n18 0.214786
R60189 DVSS.n6502 DVSS.n6501 0.214786
R60190 DVSS.n30 DVSS.n16 0.214786
R60191 DVSS.n6507 DVSS.n6506 0.214786
R60192 DVSS.n6510 DVSS.n6509 0.214786
R60193 DVSS.n10 DVSS.n9 0.214786
R60194 DVSS.n6515 DVSS.n6514 0.214786
R60195 DVSS.n6516 DVSS.n8 0.214786
R60196 DVSS.n6518 DVSS.n6517 0.214786
R60197 DVSS.n6 DVSS.n5 0.214786
R60198 DVSS.n6523 DVSS.n6522 0.214786
R60199 DVSS.n6524 DVSS.n4 0.214786
R60200 DVSS.n6526 DVSS.n6525 0.214786
R60201 DVSS.n2 DVSS.n1 0.214786
R60202 DVSS.n6532 DVSS.n6531 0.214786
R60203 DVSS.n6533 DVSS.n0 0.214786
R60204 DVSS.n6529 DVSS.n0 0.214786
R60205 DVSS.n6531 DVSS.n6530 0.214786
R60206 DVSS.n6528 DVSS.n2 0.214786
R60207 DVSS.n6527 DVSS.n6526 0.214786
R60208 DVSS.n4 DVSS.n3 0.214786
R60209 DVSS.n6522 DVSS.n6521 0.214786
R60210 DVSS.n6520 DVSS.n6 0.214786
R60211 DVSS.n6519 DVSS.n6518 0.214786
R60212 DVSS.n8 DVSS.n7 0.214786
R60213 DVSS.n6514 DVSS.n6513 0.214786
R60214 DVSS.n6512 DVSS.n10 0.214786
R60215 DVSS.n6511 DVSS.n6510 0.214786
R60216 DVSS.n6506 DVSS.n6505 0.214786
R60217 DVSS.n6504 DVSS.n16 0.214786
R60218 DVSS.n6503 DVSS.n6502 0.214786
R60219 DVSS.n18 DVSS.n17 0.214786
R60220 DVSS.n6318 DVSS.n6314 0.214786
R60221 DVSS.n6320 DVSS.n6319 0.214786
R60222 DVSS.n6321 DVSS.n6313 0.214786
R60223 DVSS.n6323 DVSS.n6322 0.214786
R60224 DVSS.n6324 DVSS.n6308 0.214786
R60225 DVSS.n6326 DVSS.n6325 0.214786
R60226 DVSS.n6327 DVSS.n6307 0.214786
R60227 DVSS.n6329 DVSS.n6328 0.214786
R60228 DVSS.n6330 DVSS.n6302 0.214786
R60229 DVSS.n6332 DVSS.n6331 0.214786
R60230 DVSS.n6333 DVSS.n6301 0.214786
R60231 DVSS.n6335 DVSS.n6334 0.214786
R60232 DVSS.n6336 DVSS.n352 0.214786
R60233 DVSS.n6338 DVSS.n6337 0.214786
R60234 DVSS.n6339 DVSS.n351 0.214786
R60235 DVSS.n6341 DVSS.n6340 0.214786
R60236 DVSS.n6342 DVSS.n346 0.214786
R60237 DVSS.n6344 DVSS.n6343 0.214786
R60238 DVSS.n6345 DVSS.n345 0.214786
R60239 DVSS.n6347 DVSS.n6346 0.214786
R60240 DVSS.n6350 DVSS.n6349 0.214786
R60241 DVSS.n6351 DVSS.n338 0.214786
R60242 DVSS.n6353 DVSS.n6352 0.214786
R60243 DVSS.n6354 DVSS.n333 0.214786
R60244 DVSS.n6356 DVSS.n6355 0.214786
R60245 DVSS.n6357 DVSS.n332 0.214786
R60246 DVSS.n6359 DVSS.n6358 0.214786
R60247 DVSS.n6360 DVSS.n328 0.214786
R60248 DVSS.n6362 DVSS.n6361 0.214786
R60249 DVSS.n6363 DVSS.n326 0.214786
R60250 DVSS.n6365 DVSS.n6364 0.214786
R60251 DVSS.n327 DVSS.n325 0.214786
R60252 DVSS.n819 DVSS.n818 0.214786
R60253 DVSS.n821 DVSS.n820 0.214786
R60254 DVSS.n822 DVSS.n814 0.214786
R60255 DVSS.n824 DVSS.n823 0.214786
R60256 DVSS.n825 DVSS.n813 0.214786
R60257 DVSS.n827 DVSS.n826 0.214786
R60258 DVSS.n828 DVSS.n808 0.214786
R60259 DVSS.n830 DVSS.n829 0.214786
R60260 DVSS.n831 DVSS.n807 0.214786
R60261 DVSS.n833 DVSS.n832 0.214786
R60262 DVSS.n834 DVSS.n566 0.214786
R60263 DVSS.n836 DVSS.n835 0.214786
R60264 DVSS.n802 DVSS.n565 0.214786
R60265 DVSS.n796 DVSS.n568 0.214786
R60266 DVSS.n798 DVSS.n797 0.214786
R60267 DVSS.n795 DVSS.n570 0.214786
R60268 DVSS.n794 DVSS.n793 0.214786
R60269 DVSS.n792 DVSS.n571 0.214786
R60270 DVSS.n791 DVSS.n790 0.214786
R60271 DVSS.n789 DVSS.n572 0.214786
R60272 DVSS.n788 DVSS.n787 0.214786
R60273 DVSS.n574 DVSS.n573 0.214786
R60274 DVSS.n782 DVSS.n781 0.214786
R60275 DVSS.n780 DVSS.n576 0.214786
R60276 DVSS.n779 DVSS.n778 0.214786
R60277 DVSS.n578 DVSS.n577 0.214786
R60278 DVSS.n774 DVSS.n773 0.214786
R60279 DVSS.n772 DVSS.n580 0.214786
R60280 DVSS.n771 DVSS.n770 0.214786
R60281 DVSS.n582 DVSS.n581 0.214786
R60282 DVSS.n766 DVSS.n765 0.214786
R60283 DVSS.n764 DVSS.n584 0.214786
R60284 DVSS.n763 DVSS.n762 0.214786
R60285 DVSS.n760 DVSS.n585 0.214786
R60286 DVSS.n759 DVSS.n758 0.214786
R60287 DVSS.n757 DVSS.n586 0.214786
R60288 DVSS.n655 DVSS.n595 0.214786
R60289 DVSS.n596 DVSS.n224 0.214786
R60290 DVSS.n651 DVSS.n241 0.214786
R60291 DVSS.n650 DVSS.n598 0.214786
R60292 DVSS.n649 DVSS.n599 0.214786
R60293 DVSS.n602 DVSS.n600 0.214786
R60294 DVSS.n645 DVSS.n603 0.214786
R60295 DVSS.n644 DVSS.n604 0.214786
R60296 DVSS.n643 DVSS.n605 0.214786
R60297 DVSS.n608 DVSS.n606 0.214786
R60298 DVSS.n639 DVSS.n609 0.214786
R60299 DVSS.n638 DVSS.n610 0.214786
R60300 DVSS.n637 DVSS.n611 0.214786
R60301 DVSS.n614 DVSS.n612 0.214786
R60302 DVSS.n633 DVSS.n615 0.214786
R60303 DVSS.n632 DVSS.n616 0.214786
R60304 DVSS.n631 DVSS.n617 0.214786
R60305 DVSS.n618 DVSS.n109 0.214786
R60306 DVSS.n627 DVSS.n117 0.214786
R60307 DVSS.n626 DVSS.n134 0.214786
R60308 DVSS.n625 DVSS.n620 0.214786
R60309 DVSS.n622 DVSS.n621 0.214786
R60310 DVSS.n561 DVSS.n560 0.214786
R60311 DVSS.n841 DVSS.n840 0.214786
R60312 DVSS.n843 DVSS.n558 0.214786
R60313 DVSS.n845 DVSS.n844 0.214786
R60314 DVSS.n556 DVSS.n555 0.214786
R60315 DVSS.n850 DVSS.n849 0.214786
R60316 DVSS.n851 DVSS.n554 0.214786
R60317 DVSS.n853 DVSS.n852 0.214786
R60318 DVSS.n552 DVSS.n551 0.214786
R60319 DVSS.n859 DVSS.n858 0.214786
R60320 DVSS.n860 DVSS.n550 0.214786
R60321 DVSS.n862 DVSS.n861 0.214786
R60322 DVSS.n863 DVSS.n154 0.214786
R60323 DVSS.n547 DVSS.n166 0.214786
R60324 DVSS.n867 DVSS.n548 0.214786
R60325 DVSS.n869 DVSS.n868 0.214786
R60326 DVSS.n871 DVSS.n870 0.214786
R60327 DVSS.n545 DVSS.n544 0.214786
R60328 DVSS.n876 DVSS.n875 0.214786
R60329 DVSS.n877 DVSS.n543 0.214786
R60330 DVSS.n879 DVSS.n878 0.214786
R60331 DVSS.n541 DVSS.n540 0.214786
R60332 DVSS.n885 DVSS.n884 0.214786
R60333 DVSS.n886 DVSS.n539 0.214786
R60334 DVSS.n888 DVSS.n887 0.214786
R60335 DVSS.n889 DVSS.n535 0.214786
R60336 DVSS.n994 DVSS.n993 0.214786
R60337 DVSS.n537 DVSS.n536 0.214786
R60338 DVSS.n989 DVSS.n893 0.214786
R60339 DVSS.n988 DVSS.n894 0.214786
R60340 DVSS.n987 DVSS.n895 0.214786
R60341 DVSS.n896 DVSS.n183 0.214786
R60342 DVSS.n983 DVSS.n193 0.214786
R60343 DVSS.n982 DVSS.n898 0.214786
R60344 DVSS.n981 DVSS.n899 0.214786
R60345 DVSS.n902 DVSS.n900 0.214786
R60346 DVSS.n977 DVSS.n903 0.214786
R60347 DVSS.n976 DVSS.n904 0.214786
R60348 DVSS.n975 DVSS.n905 0.214786
R60349 DVSS.n908 DVSS.n906 0.214786
R60350 DVSS.n971 DVSS.n909 0.214786
R60351 DVSS.n970 DVSS.n910 0.214786
R60352 DVSS.n969 DVSS.n911 0.214786
R60353 DVSS.n914 DVSS.n912 0.214786
R60354 DVSS.n965 DVSS.n915 0.214786
R60355 DVSS.n964 DVSS.n916 0.214786
R60356 DVSS.n963 DVSS.n917 0.214786
R60357 DVSS.n918 DVSS.n273 0.214786
R60358 DVSS.n959 DVSS.n249 0.214786
R60359 DVSS.n958 DVSS.n258 0.214786
R60360 DVSS.n956 DVSS.n920 0.214786
R60361 DVSS.n924 DVSS.n921 0.214786
R60362 DVSS.n952 DVSS.n925 0.214786
R60363 DVSS.n951 DVSS.n926 0.214786
R60364 DVSS.n950 DVSS.n927 0.214786
R60365 DVSS.n930 DVSS.n928 0.214786
R60366 DVSS.n946 DVSS.n931 0.214786
R60367 DVSS.n945 DVSS.n932 0.214786
R60368 DVSS.n944 DVSS.n933 0.214786
R60369 DVSS.n936 DVSS.n934 0.214786
R60370 DVSS.n940 DVSS.n937 0.214786
R60371 DVSS.n939 DVSS.n935 0.214786
R60372 DVSS.n941 DVSS.n940 0.214786
R60373 DVSS.n942 DVSS.n934 0.214786
R60374 DVSS.n944 DVSS.n943 0.214786
R60375 DVSS.n945 DVSS.n929 0.214786
R60376 DVSS.n947 DVSS.n946 0.214786
R60377 DVSS.n948 DVSS.n928 0.214786
R60378 DVSS.n950 DVSS.n949 0.214786
R60379 DVSS.n951 DVSS.n923 0.214786
R60380 DVSS.n953 DVSS.n952 0.214786
R60381 DVSS.n954 DVSS.n921 0.214786
R60382 DVSS.n956 DVSS.n955 0.214786
R60383 DVSS.n958 DVSS.n919 0.214786
R60384 DVSS.n960 DVSS.n959 0.214786
R60385 DVSS.n961 DVSS.n918 0.214786
R60386 DVSS.n963 DVSS.n962 0.214786
R60387 DVSS.n964 DVSS.n913 0.214786
R60388 DVSS.n966 DVSS.n965 0.214786
R60389 DVSS.n967 DVSS.n912 0.214786
R60390 DVSS.n969 DVSS.n968 0.214786
R60391 DVSS.n970 DVSS.n907 0.214786
R60392 DVSS.n972 DVSS.n971 0.214786
R60393 DVSS.n973 DVSS.n906 0.214786
R60394 DVSS.n975 DVSS.n974 0.214786
R60395 DVSS.n976 DVSS.n901 0.214786
R60396 DVSS.n978 DVSS.n977 0.214786
R60397 DVSS.n979 DVSS.n900 0.214786
R60398 DVSS.n981 DVSS.n980 0.214786
R60399 DVSS.n982 DVSS.n897 0.214786
R60400 DVSS.n984 DVSS.n983 0.214786
R60401 DVSS.n985 DVSS.n896 0.214786
R60402 DVSS.n987 DVSS.n986 0.214786
R60403 DVSS.n988 DVSS.n892 0.214786
R60404 DVSS.n990 DVSS.n989 0.214786
R60405 DVSS.n991 DVSS.n537 0.214786
R60406 DVSS.n993 DVSS.n992 0.214786
R60407 DVSS.n890 DVSS.n889 0.214786
R60408 DVSS.n888 DVSS.n538 0.214786
R60409 DVSS.n882 DVSS.n539 0.214786
R60410 DVSS.n884 DVSS.n883 0.214786
R60411 DVSS.n881 DVSS.n541 0.214786
R60412 DVSS.n880 DVSS.n879 0.214786
R60413 DVSS.n543 DVSS.n542 0.214786
R60414 DVSS.n875 DVSS.n874 0.214786
R60415 DVSS.n873 DVSS.n545 0.214786
R60416 DVSS.n872 DVSS.n871 0.214786
R60417 DVSS.n868 DVSS.n546 0.214786
R60418 DVSS.n867 DVSS.n866 0.214786
R60419 DVSS.n865 DVSS.n547 0.214786
R60420 DVSS.n864 DVSS.n863 0.214786
R60421 DVSS.n862 DVSS.n549 0.214786
R60422 DVSS.n856 DVSS.n550 0.214786
R60423 DVSS.n858 DVSS.n857 0.214786
R60424 DVSS.n855 DVSS.n552 0.214786
R60425 DVSS.n854 DVSS.n853 0.214786
R60426 DVSS.n554 DVSS.n553 0.214786
R60427 DVSS.n849 DVSS.n848 0.214786
R60428 DVSS.n847 DVSS.n556 0.214786
R60429 DVSS.n846 DVSS.n845 0.214786
R60430 DVSS.n558 DVSS.n557 0.214786
R60431 DVSS.n840 DVSS.n839 0.214786
R60432 DVSS.n563 DVSS.n561 0.214786
R60433 DVSS.n623 DVSS.n622 0.214786
R60434 DVSS.n625 DVSS.n624 0.214786
R60435 DVSS.n626 DVSS.n619 0.214786
R60436 DVSS.n628 DVSS.n627 0.214786
R60437 DVSS.n629 DVSS.n618 0.214786
R60438 DVSS.n631 DVSS.n630 0.214786
R60439 DVSS.n632 DVSS.n613 0.214786
R60440 DVSS.n634 DVSS.n633 0.214786
R60441 DVSS.n635 DVSS.n612 0.214786
R60442 DVSS.n637 DVSS.n636 0.214786
R60443 DVSS.n638 DVSS.n607 0.214786
R60444 DVSS.n640 DVSS.n639 0.214786
R60445 DVSS.n641 DVSS.n606 0.214786
R60446 DVSS.n643 DVSS.n642 0.214786
R60447 DVSS.n644 DVSS.n601 0.214786
R60448 DVSS.n646 DVSS.n645 0.214786
R60449 DVSS.n647 DVSS.n600 0.214786
R60450 DVSS.n649 DVSS.n648 0.214786
R60451 DVSS.n650 DVSS.n597 0.214786
R60452 DVSS.n652 DVSS.n651 0.214786
R60453 DVSS.n653 DVSS.n596 0.214786
R60454 DVSS.n655 DVSS.n654 0.214786
R60455 DVSS.n6070 DVSS.n6068 0.2003
R60456 DVSS.n6051 DVSS.n1198 0.2003
R60457 DVSS.n6101 DVSS.n1151 0.2003
R60458 DVSS.n6092 DVSS.n1166 0.2003
R60459 DVSS DVSS.n5601 0.191946
R60460 DVSS DVSS.n5607 0.191946
R60461 DVSS DVSS.n1329 0.191946
R60462 DVSS DVSS.n5618 0.191946
R60463 DVSS DVSS.n5624 0.191946
R60464 DVSS DVSS.n1325 0.191946
R60465 DVSS DVSS.n5635 0.191946
R60466 DVSS.n5643 DVSS 0.191946
R60467 DVSS.n5709 DVSS 0.191946
R60468 DVSS DVSS.n1236 0.191946
R60469 DVSS DVSS.n1231 0.191946
R60470 DVSS DVSS.n5727 0.191946
R60471 DVSS.n5736 DVSS 0.191946
R60472 DVSS DVSS.n1218 0.191946
R60473 DVSS DVSS.n5744 0.191946
R60474 DVSS.n5753 DVSS 0.191946
R60475 DVSS DVSS.n1205 0.191946
R60476 DVSS DVSS.n5764 0.191946
R60477 DVSS DVSS.n1200 0.191946
R60478 DVSS DVSS.n6064 0.191946
R60479 DVSS DVSS.n1156 0.191946
R60480 DVSS DVSS.n1141 0.191946
R60481 DVSS DVSS.n6109 0.191946
R60482 DVSS DVSS.n1136 0.191946
R60483 DVSS DVSS.n425 0.191946
R60484 DVSS DVSS.n1103 0.191946
R60485 DVSS DVSS.n1114 0.191946
R60486 DVSS DVSS.n6205 0.191946
R60487 DVSS.n6223 DVSS 0.191946
R60488 DVSS DVSS.n6245 0.191946
R60489 DVSS DVSS.n6268 0.191946
R60490 DVSS DVSS.n6279 0.191946
R60491 DVSS DVSS.n77 0.191946
R60492 DVSS DVSS.n373 0.191946
R60493 DVSS DVSS.n6493 0.191946
R60494 DVSS DVSS.n6376 0.191946
R60495 DVSS DVSS.n6388 0.191946
R60496 DVSS DVSS.n265 0.191946
R60497 DVSS.n6407 DVSS 0.191946
R60498 DVSS DVSS.n179 0.191946
R60499 DVSS.n3064 DVSS.n2395 0.191946
R60500 DVSS.n5681 DVSS.n5680 0.189567
R60501 DVSS.n4068 DVSS.t9 0.187174
R60502 DVSS.n4123 DVSS.t3 0.187174
R60503 DVSS.n4364 DVSS.t1 0.187174
R60504 DVSS.n4364 DVSS.t9 0.187174
R60505 DVSS.n4363 DVSS.t0 0.187174
R60506 DVSS.n4363 DVSS.t3 0.187174
R60507 DVSS.n1965 DVSS.t4 0.187174
R60508 DVSS.n1965 DVSS.t1 0.187174
R60509 DVSS.n1964 DVSS.t2 0.187174
R60510 DVSS.n1964 DVSS.t0 0.187174
R60511 DVSS.n4786 DVSS.t5 0.187174
R60512 DVSS.n4786 DVSS.t4 0.187174
R60513 DVSS.n4785 DVSS.t8 0.187174
R60514 DVSS.n4785 DVSS.t2 0.187174
R60515 DVSS.n5376 DVSS.t5 0.187174
R60516 DVSS.n1412 DVSS.t8 0.187174
R60517 DVSS.n3525 DVSS.n3524 0.186867
R60518 DVSS.n3534 DVSS.n3533 0.186867
R60519 DVSS.n5659 DVSS.n1284 0.17981
R60520 DVSS.n1284 DVSS.n1282 0.17981
R60521 DVSS.n4745 DVSS.n4744 0.173833
R60522 DVSS.n4744 DVSS.n1273 0.173833
R60523 DVSS.n5595 DVSS.n1333 0.1679
R60524 DVSS.n5592 DVSS.n5586 0.1679
R60525 DVSS.n5657 DVSS.n1298 0.1679
R60526 DVSS.n3942 DVSS.n1285 0.1679
R60527 DVSS.n5593 DVSS.n1270 0.159184
R60528 DVSS.n3080 DVSS.n3079 0.159115
R60529 DVSS.n3084 DVSS.n3072 0.158395
R60530 DVSS.n3080 DVSS.n3072 0.158395
R60531 DVSS.n2390 DVSS.n2389 0.158395
R60532 DVSS.n2389 DVSS.n2376 0.158395
R60533 DVSS.n2383 DVSS.n2376 0.158395
R60534 DVSS.n2391 DVSS.n2375 0.158395
R60535 DVSS.n2391 DVSS.n2390 0.158395
R60536 DVSS.n4929 DVSS.n1780 0.155773
R60537 DVSS.n4967 DVSS.n1764 0.155773
R60538 DVSS.n2375 DVSS.n2368 0.15017
R60539 DVSS.n2752 DVSS.n2407 0.149772
R60540 DVSS.n1296 DVSS 0.149572
R60541 DVSS.n1268 DVSS 0.149572
R60542 DVSS.n1269 DVSS 0.149572
R60543 DVSS.n1287 DVSS 0.149479
R60544 DVSS.n1290 DVSS 0.149479
R60545 DVSS.n1263 DVSS 0.149479
R60546 DVSS.n1265 DVSS 0.149479
R60547 DVSS.n1267 DVSS 0.149479
R60548 DVSS.n3505 DVSS.n3504 0.146974
R60549 DVSS.n3514 DVSS.n3513 0.146974
R60550 DVSS.n3095 DVSS.n2367 0.146893
R60551 DVSS.n1291 DVSS.n1283 0.144944
R60552 DVSS.n2906 DVSS 0.144526
R60553 DVSS.n5356 DVSS.n1386 0.137755
R60554 DVSS.n2845 DVSS 0.130618
R60555 DVSS.n5055 DVSS 0.130618
R60556 DVSS.n5101 DVSS 0.130618
R60557 DVSS.n5522 DVSS 0.130618
R60558 DVSS.n5981 DVSS 0.130618
R60559 DVSS.n5782 DVSS.n1194 0.1283
R60560 DVSS.n5805 DVSS.n1137 0.1283
R60561 DVSS.n6104 DVSS.n6103 0.1283
R60562 DVSS.n6106 DVSS.n1140 0.1283
R60563 DVSS.n5347 DVSS.n5346 0.12785
R60564 DVSS.n5167 DVSS.n5166 0.12785
R60565 DVSS.n4638 DVSS.n1803 0.12785
R60566 DVSS.n4447 DVSS.n4431 0.12785
R60567 DVSS.n3066 DVSS.n2395 0.126026
R60568 DVSS.n6444 DVSS 0.126026
R60569 DVSS.n6405 DVSS 0.126026
R60570 DVSS.n267 DVSS 0.126026
R60571 DVSS.n6390 DVSS 0.126026
R60572 DVSS.n6378 DVSS 0.126026
R60573 DVSS.n6495 DVSS 0.126026
R60574 DVSS.n375 DVSS 0.126026
R60575 DVSS.n6288 DVSS 0.126026
R60576 DVSS.n6281 DVSS 0.126026
R60577 DVSS.n6270 DVSS 0.126026
R60578 DVSS.n6247 DVSS 0.126026
R60579 DVSS.n6221 DVSS 0.126026
R60580 DVSS.n6207 DVSS 0.126026
R60581 DVSS.n1116 DVSS 0.126026
R60582 DVSS.n1105 DVSS 0.126026
R60583 DVSS.n6121 DVSS 0.126026
R60584 DVSS.n6117 DVSS 0.126026
R60585 DVSS.n6111 DVSS 0.126026
R60586 DVSS.n5785 DVSS 0.126026
R60587 DVSS.n6057 DVSS 0.126026
R60588 DVSS.n6066 DVSS 0.126026
R60589 DVSS.n5772 DVSS 0.126026
R60590 DVSS.n5766 DVSS 0.126026
R60591 DVSS.n1211 DVSS 0.126026
R60592 DVSS.n5751 DVSS 0.126026
R60593 DVSS.n5746 DVSS 0.126026
R60594 DVSS.n1224 DVSS 0.126026
R60595 DVSS.n5734 DVSS 0.126026
R60596 DVSS.n5729 DVSS 0.126026
R60597 DVSS.n5692 DVSS 0.126026
R60598 DVSS.n1244 DVSS 0.126026
R60599 DVSS.n5707 DVSS 0.126026
R60600 DVSS DVSS.n5642 0.126026
R60601 DVSS.n5637 DVSS 0.126026
R60602 DVSS.n5632 DVSS 0.126026
R60603 DVSS.n5626 DVSS 0.126026
R60604 DVSS.n5620 DVSS 0.126026
R60605 DVSS.n5615 DVSS 0.126026
R60606 DVSS.n5609 DVSS 0.126026
R60607 DVSS.n5603 DVSS 0.126026
R60608 DVSS.n5600 DVSS.n1254 0.124418
R60609 DVSS.n2419 DVSS.n1774 0.115687
R60610 DVSS.n4962 DVSS.n1748 0.115687
R60611 DVSS.n5687 DVSS.n1240 0.115687
R60612 DVSS.n5690 DVSS.n5689 0.115687
R60613 DVSS.n2380 DVSS.n2378 0.115202
R60614 DVSS.n4953 DVSS.n1782 0.113608
R60615 DVSS.n4929 DVSS.n1782 0.113608
R60616 DVSS.n4932 DVSS.n4931 0.113608
R60617 DVSS.n4967 DVSS.n1759 0.113608
R60618 DVSS.n4982 DVSS.n1759 0.113608
R60619 DVSS.n4982 DVSS.n4981 0.113608
R60620 DVSS.n4930 DVSS.n4929 0.113608
R60621 DVSS.n4931 DVSS.n4930 0.113608
R60622 DVSS.n4977 DVSS.n4976 0.113608
R60623 DVSS.n4976 DVSS.n1769 0.113608
R60624 DVSS.n4967 DVSS.n1769 0.113608
R60625 DVSS.n4954 DVSS.n4953 0.113608
R60626 DVSS.n3035 DVSS.n2423 0.113168
R60627 DVSS DVSS.n2906 0.111845
R60628 DVSS.n6381 DVSS.n6380 0.1112
R60629 DVSS.n281 DVSS.n280 0.1112
R60630 DVSS.n6474 DVSS.n6473 0.1112
R60631 DVSS.n240 DVSS.n64 0.1112
R60632 DVSS.n5675 DVSS.n5674 0.108833
R60633 DVSS.n5674 DVSS.n5673 0.108833
R60634 DVSS.n2845 DVSS 0.10093
R60635 DVSS.n5055 DVSS 0.10093
R60636 DVSS.n5101 DVSS 0.10093
R60637 DVSS.n5522 DVSS 0.10093
R60638 DVSS.n5981 DVSS 0.10093
R60639 DVSS.n3512 DVSS.n3511 0.100706
R60640 DVSS.n3512 DVSS.n2138 0.100706
R60641 DVSS.n3287 DVSS.n3283 0.100706
R60642 DVSS.n3288 DVSS.n3287 0.100706
R60643 DVSS.n3288 DVSS.n3281 0.100706
R60644 DVSS.n3292 DVSS.n3281 0.100706
R60645 DVSS.n3293 DVSS.n3292 0.100706
R60646 DVSS.n3077 DVSS.n3076 0.100706
R60647 DVSS.n3507 DVSS.n2141 0.100706
R60648 DVSS.n3503 DVSS.n2141 0.100706
R60649 DVSS.n6125 DVSS.n6123 0.0932
R60650 DVSS.n1133 DVSS.n1132 0.0932
R60651 DVSS.n6234 DVSS.n6233 0.0932
R60652 DVSS.n6237 DVSS.n6236 0.0932
R60653 DVSS.n2382 DVSS.n2378 0.08969
R60654 DVSS.n2385 DVSS.n2384 0.08969
R60655 DVSS.n2386 DVSS.n2377 0.08969
R60656 DVSS.n2388 DVSS.n2387 0.08969
R60657 DVSS.n2374 DVSS.n2373 0.08969
R60658 DVSS.n3089 DVSS.n2392 0.08969
R60659 DVSS.n3090 DVSS.n2371 0.08969
R60660 DVSS.n3092 DVSS.n3091 0.08969
R60661 DVSS.n2372 DVSS.n2370 0.08969
R60662 DVSS.n3082 DVSS.n3081 0.08969
R60663 DVSS.n5600 DVSS.n1328 0.0824403
R60664 DVSS.n5616 DVSS.n1328 0.0824403
R60665 DVSS.n5617 DVSS.n5616 0.0824403
R60666 DVSS.n5617 DVSS.n1324 0.0824403
R60667 DVSS.n5633 DVSS.n1324 0.0824403
R60668 DVSS.n5634 DVSS.n5633 0.0824403
R60669 DVSS.n5634 DVSS.n1239 0.0824403
R60670 DVSS.n5708 DVSS.n1239 0.0824403
R60671 DVSS.n5708 DVSS.n1240 0.0824403
R60672 DVSS.n5690 DVSS.n1221 0.0824403
R60673 DVSS.n5735 DVSS.n1221 0.0824403
R60674 DVSS.n5735 DVSS.n1222 0.0824403
R60675 DVSS.n1222 DVSS.n1208 0.0824403
R60676 DVSS.n5752 DVSS.n1208 0.0824403
R60677 DVSS.n5752 DVSS.n1209 0.0824403
R60678 DVSS.n1209 DVSS.n1199 0.0824403
R60679 DVSS.n5773 DVSS.n1199 0.0824403
R60680 DVSS.n6062 DVSS.n5773 0.0824403
R60681 DVSS.n5786 DVSS.n1134 0.0824403
R60682 DVSS.n6118 DVSS.n1134 0.0824403
R60683 DVSS.n6119 DVSS.n6118 0.0824403
R60684 DVSS.n2470 DVSS.n2464 0.0788099
R60685 DVSS.n3508 DVSS.n2140 0.0785115
R60686 DVSS.n3510 DVSS.n2137 0.0785115
R60687 DVSS.n1072 DVSS.n29 0.0779
R60688 DVSS.n6259 DVSS.n6258 0.0779
R60689 DVSS.n498 DVSS.n87 0.0779
R60690 DVSS.n492 DVSS.n72 0.0779
R60691 DVSS.n3286 DVSS.n3285 0.0758488
R60692 DVSS.n3075 DVSS.n3074 0.0758488
R60693 DVSS.n4067 DVSS.n4066 0.0758261
R60694 DVSS.n5505 DVSS.n1371 0.0758261
R60695 DVSS.n4331 DVSS.n4329 0.0758261
R60696 DVSS.n5352 DVSS.n5350 0.0758261
R60697 DVSS.n6062 DVSS.n6061 0.0750522
R60698 DVSS.n2134 DVSS.n2123 0.0734487
R60699 DVSS.n3540 DVSS.n2106 0.0718204
R60700 DVSS.n3547 DVSS.n3546 0.0718204
R60701 DVSS.n3696 DVSS.n3695 0.0718204
R60702 DVSS.n3900 DVSS.n3895 0.0718204
R60703 DVSS.n6090 DVSS.n1167 0.0718204
R60704 DVSS.n2395 DVSS.n2134 0.0702987
R60705 DVSS.n2381 DVSS.n1279 0.0682385
R60706 DVSS.n2464 DVSS.n2455 0.0652766
R60707 DVSS.n1048 DVSS 0.0650427
R60708 DVSS.n938 DVSS 0.0646027
R60709 DVSS.n6534 DVSS 0.0645092
R60710 DVSS.n5322 DVSS 0.0638222
R60711 DVSS.n5680 DVSS.n1261 0.0629627
R60712 DVSS.n3084 DVSS.n3083 0.061538
R60713 DVSS.n6534 DVSS 0.0608995
R60714 DVSS.n3083 DVSS.n3082 0.060427
R60715 DVSS DVSS.n5602 0.059934
R60716 DVSS DVSS.n5608 0.059934
R60717 DVSS DVSS.n5614 0.059934
R60718 DVSS DVSS.n5619 0.059934
R60719 DVSS DVSS.n5625 0.059934
R60720 DVSS DVSS.n5631 0.059934
R60721 DVSS DVSS.n5636 0.059934
R60722 DVSS DVSS.n1321 0.059934
R60723 DVSS DVSS.n1238 0.059934
R60724 DVSS DVSS.n1243 0.059934
R60725 DVSS DVSS.n5691 0.059934
R60726 DVSS DVSS.n5728 0.059934
R60727 DVSS DVSS.n1220 0.059934
R60728 DVSS DVSS.n1223 0.059934
R60729 DVSS DVSS.n5745 0.059934
R60730 DVSS DVSS.n1207 0.059934
R60731 DVSS DVSS.n1210 0.059934
R60732 DVSS DVSS.n5765 0.059934
R60733 DVSS DVSS.n5771 0.059934
R60734 DVSS DVSS.n6065 0.059934
R60735 DVSS DVSS.n6056 0.059934
R60736 DVSS DVSS.n5784 0.059934
R60737 DVSS DVSS.n6110 0.059934
R60738 DVSS DVSS.n6116 0.059934
R60739 DVSS DVSS.n6120 0.059934
R60740 DVSS DVSS.n1104 0.059934
R60741 DVSS DVSS.n1115 0.059934
R60742 DVSS DVSS.n6206 0.059934
R60743 DVSS DVSS.n455 0.059934
R60744 DVSS DVSS.n6246 0.059934
R60745 DVSS DVSS.n6269 0.059934
R60746 DVSS DVSS.n6280 0.059934
R60747 DVSS DVSS.n6287 0.059934
R60748 DVSS DVSS.n374 0.059934
R60749 DVSS DVSS.n6494 0.059934
R60750 DVSS DVSS.n6377 0.059934
R60751 DVSS DVSS.n6389 0.059934
R60752 DVSS DVSS.n266 0.059934
R60753 DVSS DVSS.n246 0.059934
R60754 DVSS DVSS.n6443 0.059934
R60755 DVSS.n2679 DVSS.n2106 0.059485
R60756 DVSS.n3689 DVSS.n3547 0.059485
R60757 DVSS.n3880 DVSS.n3696 0.059485
R60758 DVSS.n3938 DVSS.n3900 0.059485
R60759 DVSS.n5856 DVSS.n1167 0.059485
R60760 DVSS.n2603 DVSS.n2602 0.0569562
R60761 DVSS.n2605 DVSS.n2604 0.0569562
R60762 DVSS.n2607 DVSS.n2606 0.0569562
R60763 DVSS.n2882 DVSS.n2881 0.0569562
R60764 DVSS.n2876 DVSS.n2615 0.0569562
R60765 DVSS.n1695 DVSS.n1688 0.0569562
R60766 DVSS.n1694 DVSS.n1689 0.0569562
R60767 DVSS.n1693 DVSS.n1690 0.0569562
R60768 DVSS.n1692 DVSS.n1691 0.0569562
R60769 DVSS.n1684 DVSS.n1676 0.0569562
R60770 DVSS.n1683 DVSS.n1677 0.0569562
R60771 DVSS.n1682 DVSS.n1678 0.0569562
R60772 DVSS.n1681 DVSS.n1679 0.0569562
R60773 DVSS.n1528 DVSS.n1526 0.0569562
R60774 DVSS.n1530 DVSS.n1529 0.0569562
R60775 DVSS.n1532 DVSS.n1531 0.0569562
R60776 DVSS.n1534 DVSS.n1533 0.0569562
R60777 DVSS.n1536 DVSS.n1535 0.0569562
R60778 DVSS.n1538 DVSS.n1537 0.0569562
R60779 DVSS.n1540 DVSS.n1539 0.0569562
R60780 DVSS.n1542 DVSS.n1541 0.0569562
R60781 DVSS.n1544 DVSS.n1543 0.0569562
R60782 DVSS.n1546 DVSS.n1545 0.0569562
R60783 DVSS.n1548 DVSS.n1547 0.0569562
R60784 DVSS.n1368 DVSS.n1360 0.0569562
R60785 DVSS.n1367 DVSS.n1361 0.0569562
R60786 DVSS.n1366 DVSS.n1362 0.0569562
R60787 DVSS.n1365 DVSS.n1363 0.0569562
R60788 DVSS.n1189 DVSS.n1188 0.0569562
R60789 DVSS.n1195 DVSS.n1190 0.0569562
R60790 DVSS.n6124 DVSS.n1076 0.0569562
R60791 DVSS.n1094 DVSS.n1093 0.0569562
R60792 DVSS.n1093 DVSS.n1077 0.0569562
R60793 DVSS.n1092 DVSS.n1091 0.0569562
R60794 DVSS.n1091 DVSS.n1079 0.0569562
R60795 DVSS.n1090 DVSS.n1089 0.0569562
R60796 DVSS.n1089 DVSS.n1081 0.0569562
R60797 DVSS.n1087 DVSS.n1086 0.0569562
R60798 DVSS.n1086 DVSS.n1083 0.0569562
R60799 DVSS.n6129 DVSS.n6127 0.0569562
R60800 DVSS.n6130 DVSS.n6128 0.0569562
R60801 DVSS.n32 DVSS.n31 0.0569562
R60802 DVSS.n34 DVSS.n33 0.0569562
R60803 DVSS.n35 DVSS.n28 0.0569562
R60804 DVSS.n37 DVSS.n25 0.0569562
R60805 DVSS.n39 DVSS.n22 0.0569562
R60806 DVSS.n42 DVSS.n41 0.0569562
R60807 DVSS.n41 DVSS.n21 0.0569562
R60808 DVSS.n6499 DVSS.n43 0.0569562
R60809 DVSS.n43 DVSS.n20 0.0569562
R60810 DVSS.n6394 DVSS.n256 0.0569562
R60811 DVSS.n278 DVSS.n256 0.0569562
R60812 DVSS.n6395 DVSS.n254 0.0569562
R60813 DVSS.n277 DVSS.n254 0.0569562
R60814 DVSS.n253 DVSS.n248 0.0569562
R60815 DVSS.n276 DVSS.n253 0.0569562
R60816 DVSS.n6396 DVSS.n251 0.0569562
R60817 DVSS.n275 DVSS.n251 0.0569562
R60818 DVSS.n274 DVSS.n250 0.0569562
R60819 DVSS.n1190 DVSS.n1189 0.0569562
R60820 DVSS.n1188 DVSS.n1187 0.0569562
R60821 DVSS.n1364 DVSS.n1363 0.0569562
R60822 DVSS.n1365 DVSS.n1362 0.0569562
R60823 DVSS.n1366 DVSS.n1361 0.0569562
R60824 DVSS.n1367 DVSS.n1360 0.0569562
R60825 DVSS.n1368 DVSS.n1359 0.0569562
R60826 DVSS.n1547 DVSS.n1546 0.0569562
R60827 DVSS.n1545 DVSS.n1544 0.0569562
R60828 DVSS.n1543 DVSS.n1542 0.0569562
R60829 DVSS.n1541 DVSS.n1540 0.0569562
R60830 DVSS.n1539 DVSS.n1538 0.0569562
R60831 DVSS.n1537 DVSS.n1536 0.0569562
R60832 DVSS.n1535 DVSS.n1534 0.0569562
R60833 DVSS.n1533 DVSS.n1532 0.0569562
R60834 DVSS.n1531 DVSS.n1530 0.0569562
R60835 DVSS.n1529 DVSS.n1528 0.0569562
R60836 DVSS.n5345 DVSS.n1526 0.0569562
R60837 DVSS.n1680 DVSS.n1679 0.0569562
R60838 DVSS.n1681 DVSS.n1678 0.0569562
R60839 DVSS.n1682 DVSS.n1677 0.0569562
R60840 DVSS.n1683 DVSS.n1676 0.0569562
R60841 DVSS.n1684 DVSS.n1675 0.0569562
R60842 DVSS.n1691 DVSS.n1685 0.0569562
R60843 DVSS.n1692 DVSS.n1690 0.0569562
R60844 DVSS.n1693 DVSS.n1689 0.0569562
R60845 DVSS.n1694 DVSS.n1688 0.0569562
R60846 DVSS.n1695 DVSS.n1687 0.0569562
R60847 DVSS.n2877 DVSS.n2612 0.0569562
R60848 DVSS.n2881 DVSS.n2615 0.0569562
R60849 DVSS.n2882 DVSS.n2608 0.0569562
R60850 DVSS.n2886 DVSS.n2607 0.0569562
R60851 DVSS.n2606 DVSS.n2605 0.0569562
R60852 DVSS.n2604 DVSS.n2603 0.0569562
R60853 DVSS.n2602 DVSS.n2601 0.0569562
R60854 DVSS.n3060 DVSS.n3059 0.0569562
R60855 DVSS.n3059 DVSS.n3058 0.0569562
R60856 DVSS.n3058 DVSS.n3057 0.0569562
R60857 DVSS.n3057 DVSS.n3056 0.0569562
R60858 DVSS.n3056 DVSS.n3055 0.0569562
R60859 DVSS.n3055 DVSS.n3054 0.0569562
R60860 DVSS.n3054 DVSS.n3053 0.0569562
R60861 DVSS.n3050 DVSS.n3049 0.0569562
R60862 DVSS.n3049 DVSS.n3048 0.0569562
R60863 DVSS.n3048 DVSS.n3047 0.0569562
R60864 DVSS.n3047 DVSS.n3046 0.0569562
R60865 DVSS.n2405 DVSS.n2403 0.0569562
R60866 DVSS.n4974 DVSS.n4973 0.0569562
R60867 DVSS.n4969 DVSS.n1772 0.0569562
R60868 DVSS.n1726 DVSS.n1725 0.0569562
R60869 DVSS.n1725 DVSS.n1724 0.0569562
R60870 DVSS.n1724 DVSS.n1723 0.0569562
R60871 DVSS.n1723 DVSS.n1722 0.0569562
R60872 DVSS.n3753 DVSS.n1652 0.0569562
R60873 DVSS.n3753 DVSS.n1653 0.0569562
R60874 DVSS.n3752 DVSS.n1653 0.0569562
R60875 DVSS.n3752 DVSS.n1654 0.0569562
R60876 DVSS.n3751 DVSS.n1654 0.0569562
R60877 DVSS.n3751 DVSS.n1655 0.0569562
R60878 DVSS.n3750 DVSS.n1655 0.0569562
R60879 DVSS.n3750 DVSS.n1656 0.0569562
R60880 DVSS.n1656 DVSS.n1650 0.0569562
R60881 DVSS.n1570 DVSS.n1569 0.0569562
R60882 DVSS.n1571 DVSS.n1570 0.0569562
R60883 DVSS.n1572 DVSS.n1571 0.0569562
R60884 DVSS.n1573 DVSS.n1572 0.0569562
R60885 DVSS.n1574 DVSS.n1573 0.0569562
R60886 DVSS.n1575 DVSS.n1574 0.0569562
R60887 DVSS.n1576 DVSS.n1575 0.0569562
R60888 DVSS.n1577 DVSS.n1576 0.0569562
R60889 DVSS.n1578 DVSS.n1577 0.0569562
R60890 DVSS.n1579 DVSS.n1578 0.0569562
R60891 DVSS.n1580 DVSS.n1579 0.0569562
R60892 DVSS.n1581 DVSS.n1580 0.0569562
R60893 DVSS.n1582 DVSS.n1581 0.0569562
R60894 DVSS.n1583 DVSS.n1582 0.0569562
R60895 DVSS.n1584 DVSS.n1583 0.0569562
R60896 DVSS.n1585 DVSS.n1584 0.0569562
R60897 DVSS.n1586 DVSS.n1585 0.0569562
R60898 DVSS.n1587 DVSS.n1586 0.0569562
R60899 DVSS.n1588 DVSS.n1587 0.0569562
R60900 DVSS.n1589 DVSS.n1588 0.0569562
R60901 DVSS.n1590 DVSS.n1589 0.0569562
R60902 DVSS.n5263 DVSS.n1590 0.0569562
R60903 DVSS.n4701 DVSS.n1336 0.0569562
R60904 DVSS.n4701 DVSS.n1337 0.0569562
R60905 DVSS.n4700 DVSS.n1337 0.0569562
R60906 DVSS.n4700 DVSS.n1338 0.0569562
R60907 DVSS.n4699 DVSS.n1338 0.0569562
R60908 DVSS.n4699 DVSS.n1339 0.0569562
R60909 DVSS.n4698 DVSS.n1339 0.0569562
R60910 DVSS.n4698 DVSS.n1340 0.0569562
R60911 DVSS.n1340 DVSS.n1334 0.0569562
R60912 DVSS.n6046 DVSS.n5807 0.0569562
R60913 DVSS.n6046 DVSS.n5806 0.0569562
R60914 DVSS.n6045 DVSS.n5806 0.0569562
R60915 DVSS.n6045 DVSS.n5803 0.0569562
R60916 DVSS.n1131 DVSS.n1130 0.0569562
R60917 DVSS.n1126 DVSS.n1125 0.0569562
R60918 DVSS.n1125 DVSS.n1124 0.0569562
R60919 DVSS.n1120 DVSS.n1119 0.0569562
R60920 DVSS.n1119 DVSS.n1118 0.0569562
R60921 DVSS.n6212 DVSS.n6211 0.0569562
R60922 DVSS.n6213 DVSS.n6212 0.0569562
R60923 DVSS.n6217 DVSS.n6216 0.0569562
R60924 DVSS.n6216 DVSS.n6215 0.0569562
R60925 DVSS.n6252 DVSS.n6251 0.0569562
R60926 DVSS.n6254 DVSS.n6253 0.0569562
R60927 DVSS.n6260 DVSS.n364 0.0569562
R60928 DVSS.n6261 DVSS.n365 0.0569562
R60929 DVSS.n385 DVSS.n362 0.0569562
R60930 DVSS.n383 DVSS.n360 0.0569562
R60931 DVSS.n381 DVSS.n358 0.0569562
R60932 DVSS.n6292 DVSS.n356 0.0569562
R60933 DVSS.n380 DVSS.n356 0.0569562
R60934 DVSS.n6293 DVSS.n354 0.0569562
R60935 DVSS.n6295 DVSS.n354 0.0569562
R60936 DVSS.n204 DVSS.n191 0.0569562
R60937 DVSS.n203 DVSS.n191 0.0569562
R60938 DVSS.n205 DVSS.n189 0.0569562
R60939 DVSS.n202 DVSS.n189 0.0569562
R60940 DVSS.n206 DVSS.n187 0.0569562
R60941 DVSS.n201 DVSS.n187 0.0569562
R60942 DVSS.n186 DVSS.n182 0.0569562
R60943 DVSS.n200 DVSS.n186 0.0569562
R60944 DVSS.n199 DVSS.n185 0.0569562
R60945 DVSS.n3014 DVSS.n2440 0.0569562
R60946 DVSS.n3014 DVSS.n2439 0.0569562
R60947 DVSS.n3015 DVSS.n2439 0.0569562
R60948 DVSS.n3015 DVSS.n2438 0.0569562
R60949 DVSS.n3016 DVSS.n2438 0.0569562
R60950 DVSS.n3016 DVSS.n2437 0.0569562
R60951 DVSS.n2437 DVSS.n2434 0.0569562
R60952 DVSS.n3022 DVSS.n2426 0.0569562
R60953 DVSS.n3022 DVSS.n2427 0.0569562
R60954 DVSS.n3024 DVSS.n2427 0.0569562
R60955 DVSS.n3025 DVSS.n3024 0.0569562
R60956 DVSS.n2428 DVSS.n2424 0.0569562
R60957 DVSS.n1789 DVSS.n1788 0.0569562
R60958 DVSS.n4948 DVSS.n1790 0.0569562
R60959 DVSS.n4942 DVSS.n4941 0.0569562
R60960 DVSS.n4941 DVSS.n4940 0.0569562
R60961 DVSS.n4940 DVSS.n4939 0.0569562
R60962 DVSS.n4939 DVSS.n4938 0.0569562
R60963 DVSS.n4924 DVSS.n4923 0.0569562
R60964 DVSS.n4923 DVSS.n4922 0.0569562
R60965 DVSS.n4922 DVSS.n4921 0.0569562
R60966 DVSS.n4921 DVSS.n4920 0.0569562
R60967 DVSS.n4920 DVSS.n4919 0.0569562
R60968 DVSS.n4919 DVSS.n4918 0.0569562
R60969 DVSS.n4918 DVSS.n4917 0.0569562
R60970 DVSS.n4917 DVSS.n4916 0.0569562
R60971 DVSS.n4916 DVSS.n4915 0.0569562
R60972 DVSS.n4637 DVSS.n2039 0.0569562
R60973 DVSS.n4626 DVSS.n2039 0.0569562
R60974 DVSS.n4626 DVSS.n2038 0.0569562
R60975 DVSS.n4627 DVSS.n2038 0.0569562
R60976 DVSS.n4627 DVSS.n2037 0.0569562
R60977 DVSS.n4628 DVSS.n2037 0.0569562
R60978 DVSS.n4628 DVSS.n2036 0.0569562
R60979 DVSS.n4629 DVSS.n2036 0.0569562
R60980 DVSS.n4629 DVSS.n2035 0.0569562
R60981 DVSS.n4630 DVSS.n2035 0.0569562
R60982 DVSS.n4630 DVSS.n2034 0.0569562
R60983 DVSS.n4631 DVSS.n2034 0.0569562
R60984 DVSS.n4631 DVSS.n2033 0.0569562
R60985 DVSS.n4632 DVSS.n2033 0.0569562
R60986 DVSS.n4632 DVSS.n2032 0.0569562
R60987 DVSS.n4633 DVSS.n2032 0.0569562
R60988 DVSS.n4633 DVSS.n2031 0.0569562
R60989 DVSS.n4634 DVSS.n2031 0.0569562
R60990 DVSS.n4634 DVSS.n2030 0.0569562
R60991 DVSS.n4635 DVSS.n2030 0.0569562
R60992 DVSS.n4635 DVSS.n2029 0.0569562
R60993 DVSS.n2029 DVSS.n2026 0.0569562
R60994 DVSS.n4643 DVSS.n2025 0.0569562
R60995 DVSS.n2025 DVSS.n2024 0.0569562
R60996 DVSS.n2024 DVSS.n2023 0.0569562
R60997 DVSS.n2023 DVSS.n2022 0.0569562
R60998 DVSS.n2022 DVSS.n2021 0.0569562
R60999 DVSS.n2021 DVSS.n2020 0.0569562
R61000 DVSS.n2020 DVSS.n2019 0.0569562
R61001 DVSS.n2019 DVSS.n2018 0.0569562
R61002 DVSS.n2018 DVSS.n2017 0.0569562
R61003 DVSS.n1154 DVSS.n1149 0.0569562
R61004 DVSS.n1154 DVSS.n1148 0.0569562
R61005 DVSS.n1153 DVSS.n1148 0.0569562
R61006 DVSS.n1153 DVSS.n1145 0.0569562
R61007 DVSS.n430 DVSS.n427 0.0569562
R61008 DVSS.n452 DVSS.n439 0.0569562
R61009 DVSS.n452 DVSS.n431 0.0569562
R61010 DVSS.n447 DVSS.n438 0.0569562
R61011 DVSS.n447 DVSS.n432 0.0569562
R61012 DVSS.n450 DVSS.n437 0.0569562
R61013 DVSS.n450 DVSS.n433 0.0569562
R61014 DVSS.n449 DVSS.n436 0.0569562
R61015 DVSS.n449 DVSS.n434 0.0569562
R61016 DVSS.n6230 DVSS.n440 0.0569562
R61017 DVSS.n6231 DVSS.n441 0.0569562
R61018 DVSS.n103 DVSS.n89 0.0569562
R61019 DVSS.n104 DVSS.n90 0.0569562
R61020 DVSS.n100 DVSS.n86 0.0569562
R61021 DVSS.n98 DVSS.n84 0.0569562
R61022 DVSS.n83 DVSS.n79 0.0569562
R61023 DVSS.n95 DVSS.n93 0.0569562
R61024 DVSS.n95 DVSS.n82 0.0569562
R61025 DVSS.n6478 DVSS.n94 0.0569562
R61026 DVSS.n94 DVSS.n81 0.0569562
R61027 DVSS.n132 DVSS.n119 0.0569562
R61028 DVSS.n132 DVSS.n116 0.0569562
R61029 DVSS.n130 DVSS.n120 0.0569562
R61030 DVSS.n130 DVSS.n115 0.0569562
R61031 DVSS.n128 DVSS.n121 0.0569562
R61032 DVSS.n128 DVSS.n114 0.0569562
R61033 DVSS.n126 DVSS.n122 0.0569562
R61034 DVSS.n126 DVSS.n113 0.0569562
R61035 DVSS.n125 DVSS.n112 0.0569562
R61036 DVSS.n2466 DVSS.n2462 0.0569562
R61037 DVSS.n2466 DVSS.n2461 0.0569562
R61038 DVSS.n2467 DVSS.n2461 0.0569562
R61039 DVSS.n2467 DVSS.n2460 0.0569562
R61040 DVSS.n2468 DVSS.n2460 0.0569562
R61041 DVSS.n2468 DVSS.n2459 0.0569562
R61042 DVSS.n2469 DVSS.n2459 0.0569562
R61043 DVSS.n2108 DVSS.n2099 0.0569562
R61044 DVSS.n2108 DVSS.n2100 0.0569562
R61045 DVSS.n3541 DVSS.n2100 0.0569562
R61046 DVSS.n3542 DVSS.n3541 0.0569562
R61047 DVSS.n2102 DVSS.n2097 0.0569562
R61048 DVSS.n2096 DVSS.n2085 0.0569562
R61049 DVSS.n2096 DVSS.n2086 0.0569562
R61050 DVSS.n2095 DVSS.n2086 0.0569562
R61051 DVSS.n2095 DVSS.n2087 0.0569562
R61052 DVSS.n2094 DVSS.n2087 0.0569562
R61053 DVSS.n2094 DVSS.n2088 0.0569562
R61054 DVSS.n2093 DVSS.n2088 0.0569562
R61055 DVSS.n2093 DVSS.n2089 0.0569562
R61056 DVSS.n2089 DVSS.n2083 0.0569562
R61057 DVSS.n2082 DVSS.n2071 0.0569562
R61058 DVSS.n2082 DVSS.n2072 0.0569562
R61059 DVSS.n2081 DVSS.n2072 0.0569562
R61060 DVSS.n2081 DVSS.n2073 0.0569562
R61061 DVSS.n2080 DVSS.n2073 0.0569562
R61062 DVSS.n2080 DVSS.n2074 0.0569562
R61063 DVSS.n2079 DVSS.n2074 0.0569562
R61064 DVSS.n2079 DVSS.n2075 0.0569562
R61065 DVSS.n2075 DVSS.n2069 0.0569562
R61066 DVSS.n4446 DVSS.n2068 0.0569562
R61067 DVSS.n4434 DVSS.n2068 0.0569562
R61068 DVSS.n4434 DVSS.n2067 0.0569562
R61069 DVSS.n4435 DVSS.n2067 0.0569562
R61070 DVSS.n4435 DVSS.n2066 0.0569562
R61071 DVSS.n4436 DVSS.n2066 0.0569562
R61072 DVSS.n4436 DVSS.n2065 0.0569562
R61073 DVSS.n4437 DVSS.n2065 0.0569562
R61074 DVSS.n4437 DVSS.n2064 0.0569562
R61075 DVSS.n4438 DVSS.n2064 0.0569562
R61076 DVSS.n4438 DVSS.n2063 0.0569562
R61077 DVSS.n4439 DVSS.n2063 0.0569562
R61078 DVSS.n4439 DVSS.n2062 0.0569562
R61079 DVSS.n4440 DVSS.n2062 0.0569562
R61080 DVSS.n4440 DVSS.n2061 0.0569562
R61081 DVSS.n4441 DVSS.n2061 0.0569562
R61082 DVSS.n4441 DVSS.n2060 0.0569562
R61083 DVSS.n4442 DVSS.n2060 0.0569562
R61084 DVSS.n4442 DVSS.n2059 0.0569562
R61085 DVSS.n4443 DVSS.n2059 0.0569562
R61086 DVSS.n4443 DVSS.n2058 0.0569562
R61087 DVSS.n4444 DVSS.n2058 0.0569562
R61088 DVSS.n3952 DVSS.n3951 0.0569562
R61089 DVSS.n3951 DVSS.n3950 0.0569562
R61090 DVSS.n3950 DVSS.n3949 0.0569562
R61091 DVSS.n3949 DVSS.n3948 0.0569562
R61092 DVSS.n3948 DVSS.n3947 0.0569562
R61093 DVSS.n3947 DVSS.n3946 0.0569562
R61094 DVSS.n3946 DVSS.n3945 0.0569562
R61095 DVSS.n3945 DVSS.n3944 0.0569562
R61096 DVSS.n3944 DVSS.n3943 0.0569562
R61097 DVSS.n1169 DVSS.n1164 0.0569562
R61098 DVSS.n1169 DVSS.n1163 0.0569562
R61099 DVSS.n1168 DVSS.n1163 0.0569562
R61100 DVSS.n1168 DVSS.n1161 0.0569562
R61101 DVSS.n414 DVSS.n400 0.0569562
R61102 DVSS.n423 DVSS.n408 0.0569562
R61103 DVSS.n415 DVSS.n408 0.0569562
R61104 DVSS.n422 DVSS.n402 0.0569562
R61105 DVSS.n416 DVSS.n402 0.0569562
R61106 DVSS.n421 DVSS.n406 0.0569562
R61107 DVSS.n417 DVSS.n406 0.0569562
R61108 DVSS.n420 DVSS.n404 0.0569562
R61109 DVSS.n418 DVSS.n404 0.0569562
R61110 DVSS.n412 DVSS.n396 0.0569562
R61111 DVSS.n6240 DVSS.n6239 0.0569562
R61112 DVSS.n73 DVSS.n61 0.0569562
R61113 DVSS.n74 DVSS.n62 0.0569562
R61114 DVSS.n71 DVSS.n58 0.0569562
R61115 DVSS.n69 DVSS.n56 0.0569562
R61116 DVSS.n67 DVSS.n54 0.0569562
R61117 DVSS.n6485 DVSS.n52 0.0569562
R61118 DVSS.n66 DVSS.n52 0.0569562
R61119 DVSS.n51 DVSS.n49 0.0569562
R61120 DVSS.n6487 DVSS.n51 0.0569562
R61121 DVSS.n238 DVSS.n237 0.0569562
R61122 DVSS.n244 DVSS.n237 0.0569562
R61123 DVSS.n235 DVSS.n234 0.0569562
R61124 DVSS.n6411 DVSS.n234 0.0569562
R61125 DVSS.n232 DVSS.n231 0.0569562
R61126 DVSS.n6416 DVSS.n231 0.0569562
R61127 DVSS.n229 DVSS.n228 0.0569562
R61128 DVSS.n228 DVSS.n227 0.0569562
R61129 DVSS.n6419 DVSS.n226 0.0569562
R61130 DVSS.n227 DVSS.n226 0.0569562
R61131 DVSS.n125 DVSS.n113 0.0569562
R61132 DVSS.n200 DVSS.n185 0.0569562
R61133 DVSS.n275 DVSS.n250 0.0569562
R61134 DVSS.n73 DVSS.n62 0.0569562
R61135 DVSS.n71 DVSS.n57 0.0569562
R61136 DVSS.n69 DVSS.n55 0.0569562
R61137 DVSS.n104 DVSS.n89 0.0569562
R61138 DVSS.n99 DVSS.n86 0.0569562
R61139 DVSS.n97 DVSS.n84 0.0569562
R61140 DVSS.n6260 DVSS.n365 0.0569562
R61141 DVSS.n385 DVSS.n361 0.0569562
R61142 DVSS.n383 DVSS.n359 0.0569562
R61143 DVSS.n33 DVSS.n32 0.0569562
R61144 DVSS.n28 DVSS.n27 0.0569562
R61145 DVSS.n25 DVSS.n24 0.0569562
R61146 DVSS.n6239 DVSS.n412 0.0569562
R61147 DVSS.n6231 DVSS.n6230 0.0569562
R61148 DVSS.n6253 DVSS.n6252 0.0569562
R61149 DVSS.n6130 DVSS.n6129 0.0569562
R61150 DVSS.n4306 DVSS.n4305 0.0568736
R61151 DVSS.n4310 DVSS.n4306 0.0568736
R61152 DVSS.n4313 DVSS.n4310 0.0568736
R61153 DVSS.n4324 DVSS.n4323 0.0568736
R61154 DVSS.n4323 DVSS.n4007 0.0568736
R61155 DVSS.n3040 DVSS.n3039 0.0563
R61156 DVSS.n4425 DVSS.n4424 0.0562609
R61157 DVSS.n4424 DVSS.n4423 0.0562609
R61158 DVSS.n4423 DVSS.n3956 0.0562609
R61159 DVSS.n4413 DVSS.n3956 0.0562609
R61160 DVSS.n4413 DVSS.n4412 0.0562609
R61161 DVSS.n4412 DVSS.n4411 0.0562609
R61162 DVSS.n4411 DVSS.n3966 0.0562609
R61163 DVSS.n4401 DVSS.n3966 0.0562609
R61164 DVSS.n4401 DVSS.n4400 0.0562609
R61165 DVSS.n4400 DVSS.n4399 0.0562609
R61166 DVSS.n4399 DVSS.n3976 0.0562609
R61167 DVSS.n4389 DVSS.n3976 0.0562609
R61168 DVSS.n4389 DVSS.n4388 0.0562609
R61169 DVSS.n4388 DVSS.n4387 0.0562609
R61170 DVSS.n4387 DVSS.n3986 0.0562609
R61171 DVSS.n4377 DVSS.n3986 0.0562609
R61172 DVSS.n4377 DVSS.n4376 0.0562609
R61173 DVSS.n4376 DVSS.n4375 0.0562609
R61174 DVSS.n4375 DVSS.n3997 0.0562609
R61175 DVSS.n3997 DVSS.n3996 0.0562609
R61176 DVSS.n4907 DVSS.n4906 0.0562609
R61177 DVSS.n4906 DVSS.n4905 0.0562609
R61178 DVSS.n4905 DVSS.n1814 0.0562609
R61179 DVSS.n4895 DVSS.n1814 0.0562609
R61180 DVSS.n4895 DVSS.n4894 0.0562609
R61181 DVSS.n4894 DVSS.n4893 0.0562609
R61182 DVSS.n4893 DVSS.n1826 0.0562609
R61183 DVSS.n4883 DVSS.n1826 0.0562609
R61184 DVSS.n4883 DVSS.n4882 0.0562609
R61185 DVSS.n4882 DVSS.n4881 0.0562609
R61186 DVSS.n4881 DVSS.n1836 0.0562609
R61187 DVSS.n4871 DVSS.n1836 0.0562609
R61188 DVSS.n4871 DVSS.n4870 0.0562609
R61189 DVSS.n4870 DVSS.n4869 0.0562609
R61190 DVSS.n4869 DVSS.n1846 0.0562609
R61191 DVSS.n4859 DVSS.n1846 0.0562609
R61192 DVSS.n4859 DVSS.n4858 0.0562609
R61193 DVSS.n4858 DVSS.n4857 0.0562609
R61194 DVSS.n4857 DVSS.n1856 0.0562609
R61195 DVSS.n1970 DVSS.n1856 0.0562609
R61196 DVSS.n4749 DVSS.n1970 0.0562609
R61197 DVSS.n4844 DVSS.n1883 0.0562609
R61198 DVSS.n4844 DVSS.n4843 0.0562609
R61199 DVSS.n4843 DVSS.n4842 0.0562609
R61200 DVSS.n4842 DVSS.n1884 0.0562609
R61201 DVSS.n4832 DVSS.n1884 0.0562609
R61202 DVSS.n4832 DVSS.n4831 0.0562609
R61203 DVSS.n4831 DVSS.n4830 0.0562609
R61204 DVSS.n4830 DVSS.n1895 0.0562609
R61205 DVSS.n4820 DVSS.n1895 0.0562609
R61206 DVSS.n4820 DVSS.n4819 0.0562609
R61207 DVSS.n4819 DVSS.n4818 0.0562609
R61208 DVSS.n4818 DVSS.n1905 0.0562609
R61209 DVSS.n4808 DVSS.n1905 0.0562609
R61210 DVSS.n4808 DVSS.n4807 0.0562609
R61211 DVSS.n4807 DVSS.n4806 0.0562609
R61212 DVSS.n4806 DVSS.n1915 0.0562609
R61213 DVSS.n4796 DVSS.n1915 0.0562609
R61214 DVSS.n4796 DVSS.n4795 0.0562609
R61215 DVSS.n4795 DVSS.n4794 0.0562609
R61216 DVSS.n4794 DVSS.n1925 0.0562609
R61217 DVSS.n1925 DVSS.n1592 0.0562609
R61218 DVSS.n5259 DVSS.n1593 0.0562609
R61219 DVSS.n5249 DVSS.n1593 0.0562609
R61220 DVSS.n5249 DVSS.n5248 0.0562609
R61221 DVSS.n5248 DVSS.n5247 0.0562609
R61222 DVSS.n5247 DVSS.n1607 0.0562609
R61223 DVSS.n5237 DVSS.n1607 0.0562609
R61224 DVSS.n5237 DVSS.n5236 0.0562609
R61225 DVSS.n5236 DVSS.n5235 0.0562609
R61226 DVSS.n5235 DVSS.n1617 0.0562609
R61227 DVSS.n5225 DVSS.n1617 0.0562609
R61228 DVSS.n5225 DVSS.n5224 0.0562609
R61229 DVSS.n5224 DVSS.n5223 0.0562609
R61230 DVSS.n5223 DVSS.n1627 0.0562609
R61231 DVSS.n5213 DVSS.n1627 0.0562609
R61232 DVSS.n5213 DVSS.n5212 0.0562609
R61233 DVSS.n5212 DVSS.n5211 0.0562609
R61234 DVSS.n5211 DVSS.n1637 0.0562609
R61235 DVSS.n5201 DVSS.n1637 0.0562609
R61236 DVSS.n5201 DVSS.n5200 0.0562609
R61237 DVSS.n5200 DVSS.n1370 0.0562609
R61238 DVSS.n4335 DVSS.n4333 0.0562609
R61239 DVSS.n4336 DVSS.n4335 0.0562609
R61240 DVSS.n4338 DVSS.n4336 0.0562609
R61241 DVSS.n4339 DVSS.n4338 0.0562609
R61242 DVSS.n4341 DVSS.n4339 0.0562609
R61243 DVSS.n4342 DVSS.n4341 0.0562609
R61244 DVSS.n4344 DVSS.n4342 0.0562609
R61245 DVSS.n4345 DVSS.n4344 0.0562609
R61246 DVSS.n4347 DVSS.n4345 0.0562609
R61247 DVSS.n4348 DVSS.n4347 0.0562609
R61248 DVSS.n4350 DVSS.n4348 0.0562609
R61249 DVSS.n4351 DVSS.n4350 0.0562609
R61250 DVSS.n4353 DVSS.n4351 0.0562609
R61251 DVSS.n4354 DVSS.n4353 0.0562609
R61252 DVSS.n4356 DVSS.n4354 0.0562609
R61253 DVSS.n4357 DVSS.n4356 0.0562609
R61254 DVSS.n4358 DVSS.n4357 0.0562609
R61255 DVSS.n4360 DVSS.n4358 0.0562609
R61256 DVSS.n4360 DVSS.n4359 0.0562609
R61257 DVSS.n4359 DVSS.n1804 0.0562609
R61258 DVSS.n4911 DVSS.n1805 0.0562609
R61259 DVSS.n1933 DVSS.n1805 0.0562609
R61260 DVSS.n1935 DVSS.n1933 0.0562609
R61261 DVSS.n1936 DVSS.n1935 0.0562609
R61262 DVSS.n1938 DVSS.n1936 0.0562609
R61263 DVSS.n1939 DVSS.n1938 0.0562609
R61264 DVSS.n1941 DVSS.n1939 0.0562609
R61265 DVSS.n1942 DVSS.n1941 0.0562609
R61266 DVSS.n1944 DVSS.n1942 0.0562609
R61267 DVSS.n1945 DVSS.n1944 0.0562609
R61268 DVSS.n1947 DVSS.n1945 0.0562609
R61269 DVSS.n1948 DVSS.n1947 0.0562609
R61270 DVSS.n1950 DVSS.n1948 0.0562609
R61271 DVSS.n1951 DVSS.n1950 0.0562609
R61272 DVSS.n1953 DVSS.n1951 0.0562609
R61273 DVSS.n1954 DVSS.n1953 0.0562609
R61274 DVSS.n1956 DVSS.n1954 0.0562609
R61275 DVSS.n1957 DVSS.n1956 0.0562609
R61276 DVSS.n1959 DVSS.n1957 0.0562609
R61277 DVSS.n1960 DVSS.n1959 0.0562609
R61278 DVSS.n1961 DVSS.n1960 0.0562609
R61279 DVSS.n4755 DVSS.n4754 0.0562609
R61280 DVSS.n4757 DVSS.n4755 0.0562609
R61281 DVSS.n4758 DVSS.n4757 0.0562609
R61282 DVSS.n4760 DVSS.n4758 0.0562609
R61283 DVSS.n4761 DVSS.n4760 0.0562609
R61284 DVSS.n4763 DVSS.n4761 0.0562609
R61285 DVSS.n4764 DVSS.n4763 0.0562609
R61286 DVSS.n4766 DVSS.n4764 0.0562609
R61287 DVSS.n4767 DVSS.n4766 0.0562609
R61288 DVSS.n4769 DVSS.n4767 0.0562609
R61289 DVSS.n4770 DVSS.n4769 0.0562609
R61290 DVSS.n4772 DVSS.n4770 0.0562609
R61291 DVSS.n4773 DVSS.n4772 0.0562609
R61292 DVSS.n4775 DVSS.n4773 0.0562609
R61293 DVSS.n4776 DVSS.n4775 0.0562609
R61294 DVSS.n4778 DVSS.n4776 0.0562609
R61295 DVSS.n4779 DVSS.n4778 0.0562609
R61296 DVSS.n4780 DVSS.n4779 0.0562609
R61297 DVSS.n4782 DVSS.n4780 0.0562609
R61298 DVSS.n4782 DVSS.n4781 0.0562609
R61299 DVSS.n4781 DVSS.n1649 0.0562609
R61300 DVSS.n5172 DVSS.n5170 0.0562609
R61301 DVSS.n5173 DVSS.n5172 0.0562609
R61302 DVSS.n5175 DVSS.n5173 0.0562609
R61303 DVSS.n5176 DVSS.n5175 0.0562609
R61304 DVSS.n5178 DVSS.n5176 0.0562609
R61305 DVSS.n5179 DVSS.n5178 0.0562609
R61306 DVSS.n5181 DVSS.n5179 0.0562609
R61307 DVSS.n5182 DVSS.n5181 0.0562609
R61308 DVSS.n5184 DVSS.n5182 0.0562609
R61309 DVSS.n5185 DVSS.n5184 0.0562609
R61310 DVSS.n5187 DVSS.n5185 0.0562609
R61311 DVSS.n5188 DVSS.n5187 0.0562609
R61312 DVSS.n5190 DVSS.n5188 0.0562609
R61313 DVSS.n5191 DVSS.n5190 0.0562609
R61314 DVSS.n5193 DVSS.n5191 0.0562609
R61315 DVSS.n5194 DVSS.n5193 0.0562609
R61316 DVSS.n5195 DVSS.n5194 0.0562609
R61317 DVSS.n5197 DVSS.n5195 0.0562609
R61318 DVSS.n5197 DVSS.n5196 0.0562609
R61319 DVSS.n5196 DVSS.n1523 0.0562609
R61320 DVSS DVSS.n2109 0.0560627
R61321 DVSS.n3520 DVSS 0.0560627
R61322 DVSS.n6126 DVSS.n392 0.0554
R61323 DVSS.n6285 DVSS.n40 0.0554
R61324 DVSS.n6250 DVSS.n6249 0.0554
R61325 DVSS.n6291 DVSS.n6290 0.0554
R61326 DVSS.n443 DVSS.n394 0.0554
R61327 DVSS.n6481 DVSS.n6480 0.0554
R61328 DVSS.n6243 DVSS.n6242 0.0554
R61329 DVSS.n6484 DVSS.n6483 0.0554
R61330 DVSS.n3515 DVSS.n2137 0.055378
R61331 DVSS.n2142 DVSS.n2140 0.055378
R61332 DVSS.n1251 DVSS.n1249 0.0540178
R61333 DVSS.n1177 DVSS.n1175 0.0540178
R61334 DVSS.n6080 DVSS.n1173 0.0540178
R61335 DVSS.n503 DVSS.n491 0.0540178
R61336 DVSS.n6073 DVSS.n1182 0.0536
R61337 DVSS.n368 DVSS.n366 0.0536
R61338 DVSS.n6393 DVSS.n6392 0.0536
R61339 DVSS.n6076 DVSS.n1179 0.0536
R61340 DVSS.n378 DVSS.n377 0.0536
R61341 DVSS.n6383 DVSS.n6382 0.0536
R61342 DVSS.n1170 DVSS.n1144 0.0536
R61343 DVSS.n370 DVSS.n105 0.0536
R61344 DVSS.n6385 DVSS.n118 0.0536
R61345 DVSS.n6085 DVSS.n1160 0.0536
R61346 DVSS.n371 DVSS.n63 0.0536
R61347 DVSS.n6386 DVSS.n243 0.0536
R61348 DVSS.n5714 DVSS.n5713 0.0533261
R61349 DVSS.n5720 DVSS.n1233 0.0533261
R61350 DVSS.n5686 DVSS.n1250 0.0533261
R61351 DVSS.n5688 DVSS.n1250 0.0533261
R61352 DVSS.n5700 DVSS.n1246 0.0533261
R61353 DVSS.n5699 DVSS.n5698 0.0533261
R61354 DVSS.n495 DVSS.n219 0.0533261
R61355 DVSS.n500 DVSS.n496 0.0533261
R61356 DVSS.n505 DVSS.n502 0.0533261
R61357 DVSS.n507 DVSS.n502 0.0533261
R61358 DVSS.n6257 DVSS.n387 0.0533261
R61359 DVSS.n388 DVSS.n213 0.0533261
R61360 DVSS.n592 DVSS.n589 0.0532401
R61361 DVSS.n1757 DVSS.n1728 0.0527
R61362 DVSS.n4984 DVSS.n1719 0.0527
R61363 DVSS.n1796 DVSS.n1794 0.0527
R61364 DVSS.n4944 DVSS.n1797 0.0527
R61365 DVSS.n2926 DVSS.n2925 0.05225
R61366 DVSS.n3062 DVSS.n2398 0.05225
R61367 DVSS.n3018 DVSS.n2394 0.05225
R61368 DVSS.n2471 DVSS.n2393 0.05225
R61369 DVSS.n3286 DVSS.n3282 0.0521279
R61370 DVSS.n3075 DVSS.n2369 0.0521279
R61371 DVSS.n3521 DVSS.n2132 0.0518
R61372 DVSS.n1085 DVSS.n458 0.0518
R61373 DVSS.n6274 DVSS.n38 0.0518
R61374 DVSS.n3526 DVSS.n2128 0.0518
R61375 DVSS.n6219 DVSS.n6218 0.0518
R61376 DVSS.n6284 DVSS.n6283 0.0518
R61377 DVSS.n3532 DVSS.n2115 0.0518
R61378 DVSS.n6226 DVSS.n448 0.0518
R61379 DVSS.n6276 DVSS.n92 0.0518
R61380 DVSS.n3539 DVSS.n3538 0.0518
R61381 DVSS.n6224 DVSS.n403 0.0518
R61382 DVSS.n6277 DVSS.n76 0.0518
R61383 DVSS.n3032 DVSS.n1786 0.0507703
R61384 DVSS.n3036 DVSS.n2406 0.0507703
R61385 DVSS.n1048 DVSS 0.0501178
R61386 DVSS.n6497 DVSS.n44 0.05
R61387 DVSS.n270 DVSS.n269 0.05
R61388 DVSS.n379 DVSS.n45 0.05
R61389 DVSS.n260 DVSS.n195 0.05
R61390 DVSS.n106 DVSS.n47 0.05
R61391 DVSS.n262 DVSS.n135 0.05
R61392 DVSS.n6491 DVSS.n48 0.05
R61393 DVSS.n263 DVSS.n245 0.05
R61394 DVSS.n5597 DVSS.n1331 0.049839
R61395 DVSS.n5590 DVSS.n5589 0.049839
R61396 DVSS.n5655 DVSS.n5654 0.049839
R61397 DVSS.n1310 DVSS.n1307 0.049839
R61398 DVSS.n938 DVSS 0.0494578
R61399 DVSS.n3291 DVSS.n1277 0.0490001
R61400 DVSS.n5322 DVSS 0.0487259
R61401 DVSS.n755 DVSS.n589 0.0485826
R61402 DVSS.n1088 DVSS.n460 0.0482
R61403 DVSS.n6263 DVSS.n36 0.0482
R61404 DVSS.n6210 DVSS.n6209 0.0482
R61405 DVSS.n6273 DVSS.n6272 0.0482
R61406 DVSS.n6202 DVSS.n451 0.0482
R61407 DVSS.n6265 DVSS.n91 0.0482
R61408 DVSS.n6203 DVSS.n407 0.0482
R61409 DVSS.n6266 DVSS.n75 0.0482
R61410 DVSS.n5787 DVSS.n5786 0.0481866
R61411 DVSS.n4069 DVSS.n4007 0.0479692
R61412 DVSS.n6072 DVSS.n1184 0.0464
R61413 DVSS.n6380 DVSS.n279 0.0464
R61414 DVSS.n6402 DVSS.n247 0.0464
R61415 DVSS.n6047 DVSS.n1180 0.0464
R61416 DVSS.n6296 DVSS.n281 0.0464
R61417 DVSS.n6403 DVSS.n196 0.0464
R61418 DVSS.n6083 DVSS.n1150 0.0464
R61419 DVSS.n6475 DVSS.n6474 0.0464
R61420 DVSS.n6408 DVSS.n136 0.0464
R61421 DVSS.n6088 DVSS.n1165 0.0464
R61422 DVSS.n6488 DVSS.n64 0.0464
R61423 DVSS.n6412 DVSS.n6410 0.0464
R61424 DVSS.n2381 DVSS.n2380 0.0459602
R61425 DVSS.n5686 DVSS.n5685 0.0457174
R61426 DVSS.n6428 DVSS.n216 0.0457174
R61427 DVSS.n505 DVSS.n504 0.0457174
R61428 DVSS.n6399 DVSS.n6398 0.0456261
R61429 DVSS.n6438 DVSS.n6437 0.0456261
R61430 DVSS.n124 DVSS.n110 0.0456261
R61431 DVSS.n6424 DVSS.n6422 0.0456261
R61432 DVSS.n2613 DVSS.n2131 0.0446
R61433 DVSS.n1109 DVSS.n1108 0.0446
R61434 DVSS.n3042 DVSS.n2127 0.0446
R61435 DVSS.n1122 DVSS.n1121 0.0446
R61436 DVSS.n2430 DVSS.n2114 0.0446
R61437 DVSS.n1111 DVSS.n446 0.0446
R61438 DVSS.n3535 DVSS.n2101 0.0446
R61439 DVSS.n1112 DVSS.n401 0.0446
R61440 DVSS.n2384 DVSS.n2383 0.04343
R61441 DVSS.n2377 DVSS.n2376 0.04343
R61442 DVSS.n2389 DVSS.n2388 0.04343
R61443 DVSS.n2390 DVSS.n2374 0.04343
R61444 DVSS.n2392 DVSS.n2391 0.04343
R61445 DVSS.n2375 DVSS.n2371 0.04343
R61446 DVSS.n3081 DVSS.n3080 0.04343
R61447 DVSS.n3073 DVSS.n3072 0.04343
R61448 DVSS.n4907 DVSS.n1813 0.0430543
R61449 DVSS.n5260 DVSS.n1592 0.0430543
R61450 DVSS.n4912 DVSS.n4911 0.0430543
R61451 DVSS.n5169 DVSS.n1649 0.0430543
R61452 DVSS.n271 DVSS.n180 0.0428
R61453 DVSS.n6441 DVSS.n181 0.0428
R61454 DVSS.n6413 DVSS.n137 0.0428
R61455 DVSS.n6417 DVSS.n6415 0.0428
R61456 DVSS.n4305 DVSS.n4301 0.0424895
R61457 DVSS.n6375 DVSS.n165 0.041806
R61458 DVSS.n1098 DVSS.n1097 0.041
R61459 DVSS.n1128 DVSS.n1127 0.041
R61460 DVSS.n1100 DVSS.n453 0.041
R61461 DVSS.n1101 DVSS.n409 0.041
R61462 DVSS.n3093 DVSS.n3092 0.04037
R61463 DVSS.n3078 DVSS.n2370 0.04037
R61464 DVSS.n6432 DVSS.n211 0.0401
R61465 DVSS.n6434 DVSS.n197 0.0401
R61466 DVSS.n6469 DVSS.n6468 0.0401
R61467 DVSS.n6420 DVSS.n6418 0.0401
R61468 DVSS DVSS.n4363 0.039875
R61469 DVSS DVSS.n4364 0.039875
R61470 DVSS DVSS.n1964 0.039875
R61471 DVSS DVSS.n1965 0.039875
R61472 DVSS DVSS.n4785 0.039875
R61473 DVSS DVSS.n4786 0.039875
R61474 DVSS DVSS.n2111 0.039875
R61475 DVSS DVSS.n3523 0.039875
R61476 DVSS DVSS.n2118 0.039875
R61477 DVSS.n4314 DVSS.n4313 0.0395659
R61478 DVSS.n4324 DVSS.n4002 0.0395659
R61479 DVSS.n3092 DVSS.n2370 0.0389615
R61480 DVSS.n2392 DVSS.n2374 0.0389615
R61481 DVSS.n3284 DVSS.n3282 0.0389615
R61482 DVSS.n2384 DVSS.n2377 0.0389615
R61483 DVSS.n2384 DVSS.n2382 0.0389615
R61484 DVSS.n2388 DVSS.n2374 0.0389615
R61485 DVSS.n2388 DVSS.n2377 0.0389615
R61486 DVSS.n3092 DVSS.n2371 0.0389615
R61487 DVSS.n2392 DVSS.n2371 0.0389615
R61488 DVSS.n3081 DVSS.n3073 0.0389615
R61489 DVSS.n3081 DVSS.n2370 0.0389615
R61490 DVSS.n4702 DVSS.n1591 0.03875
R61491 DVSS.n4644 DVSS.n4642 0.03875
R61492 DVSS.n2614 DVSS.n2129 0.0374
R61493 DVSS.n3043 DVSS.n2125 0.0374
R61494 DVSS.n2431 DVSS.n2112 0.0374
R61495 DVSS.n2110 DVSS.n2104 0.0374
R61496 DVSS.n5006 DVSS.n1729 0.03695
R61497 DVSS.n5005 DVSS.n1731 0.03695
R61498 DVSS.n4936 DVSS.n4935 0.03695
R61499 DVSS.n4934 DVSS.n4928 0.03695
R61500 DVSS.n5799 DVSS.n1191 0.0365
R61501 DVSS.n6054 DVSS.n6053 0.0365
R61502 DVSS.n6097 DVSS.n1146 0.0365
R61503 DVSS.n6095 DVSS.n6094 0.0365
R61504 DVSS.n4445 DVSS.n4433 0.0362074
R61505 DVSS.n6119 DVSS.n486 0.0350896
R61506 DVSS.n3069 DVSS 0.0338686
R61507 DVSS DVSS.n3519 0.0338686
R61508 DVSS.n3516 DVSS.n3515 0.0337188
R61509 DVSS.n3085 DVSS.n2142 0.0337188
R61510 DVSS.n593 DVSS.n588 0.033707
R61511 DVSS.n594 DVSS.n591 0.033707
R61512 DVSS.n5602 DVSS.t128 0.03326
R61513 DVSS.n5602 DVSS.t98 0.03326
R61514 DVSS.n5608 DVSS.t150 0.03326
R61515 DVSS.n5608 DVSS.t118 0.03326
R61516 DVSS.n5614 DVSS.t36 0.03326
R61517 DVSS.n5614 DVSS.t88 0.03326
R61518 DVSS.n5619 DVSS.t64 0.03326
R61519 DVSS.n5619 DVSS.t108 0.03326
R61520 DVSS.n5625 DVSS.t78 0.03326
R61521 DVSS.n5625 DVSS.t120 0.03326
R61522 DVSS.n5631 DVSS.t50 0.03326
R61523 DVSS.n5631 DVSS.t142 0.03326
R61524 DVSS.n5636 DVSS.t66 0.03326
R61525 DVSS.n5636 DVSS.t30 0.03326
R61526 DVSS.n1321 DVSS.t92 0.03326
R61527 DVSS.n1321 DVSS.t164 0.03326
R61528 DVSS.n1238 DVSS.t100 0.03326
R61529 DVSS.n1238 DVSS.t174 0.03326
R61530 DVSS.n1243 DVSS.t122 0.03326
R61531 DVSS.n1243 DVSS.t42 0.03326
R61532 DVSS.n5691 DVSS.t162 0.03326
R61533 DVSS.n5691 DVSS.t48 0.03326
R61534 DVSS.n5728 DVSS.t134 0.03326
R61535 DVSS.n5728 DVSS.t70 0.03326
R61536 DVSS.n1220 DVSS.t152 0.03326
R61537 DVSS.n1220 DVSS.t86 0.03326
R61538 DVSS.n1223 DVSS.t102 0.03326
R61539 DVSS.n1223 DVSS.t178 0.03326
R61540 DVSS.n5745 DVSS.t112 0.03326
R61541 DVSS.n5745 DVSS.t32 0.03326
R61542 DVSS.n1207 DVSS.t132 0.03326
R61543 DVSS.n1207 DVSS.t54 0.03326
R61544 DVSS.n1210 DVSS.t104 0.03326
R61545 DVSS.n1210 DVSS.t74 0.03326
R61546 DVSS.n5765 DVSS.t124 0.03326
R61547 DVSS.n5765 DVSS.t94 0.03326
R61548 DVSS.n5771 DVSS.t168 0.03326
R61549 DVSS.n5771 DVSS.t60 0.03326
R61550 DVSS.n6065 DVSS.t184 0.03326
R61551 DVSS.n6065 DVSS.t84 0.03326
R61552 DVSS.n6056 DVSS.t38 0.03326
R61553 DVSS.n6056 DVSS.t90 0.03326
R61554 DVSS.n5784 DVSS.t52 0.03326
R61555 DVSS.n5784 DVSS.t144 0.03326
R61556 DVSS.n6110 DVSS.t188 0.03326
R61557 DVSS.n6110 DVSS.t156 0.03326
R61558 DVSS.n6116 DVSS.t40 0.03326
R61559 DVSS.n6116 DVSS.t176 0.03326
R61560 DVSS.n6120 DVSS.t68 0.03326
R61561 DVSS.n6120 DVSS.t146 0.03326
R61562 DVSS.n1104 DVSS.t80 0.03326
R61563 DVSS.n1104 DVSS.t166 0.03326
R61564 DVSS.n1115 DVSS.t136 0.03326
R61565 DVSS.n1115 DVSS.t180 0.03326
R61566 DVSS.n6206 DVSS.t106 0.03326
R61567 DVSS.n6206 DVSS.t44 0.03326
R61568 DVSS.n455 DVSS.t126 0.03326
R61569 DVSS.n455 DVSS.t56 0.03326
R61570 DVSS.n6246 DVSS.t138 0.03326
R61571 DVSS.n6246 DVSS.t72 0.03326
R61572 DVSS.n6269 DVSS.t82 0.03326
R61573 DVSS.n6269 DVSS.t158 0.03326
R61574 DVSS.n6280 DVSS.t96 0.03326
R61575 DVSS.n6280 DVSS.t182 0.03326
R61576 DVSS.n6287 DVSS.t114 0.03326
R61577 DVSS.n6287 DVSS.t34 0.03326
R61578 DVSS.n374 DVSS.t116 0.03326
R61579 DVSS.n374 DVSS.t58 0.03326
R61580 DVSS.n6494 DVSS.t140 0.03326
R61581 DVSS.n6494 DVSS.t76 0.03326
R61582 DVSS.n6377 DVSS.t154 0.03326
R61583 DVSS.n6377 DVSS.t46 0.03326
R61584 DVSS.n6389 DVSS.t170 0.03326
R61585 DVSS.n6389 DVSS.t62 0.03326
R61586 DVSS.n266 DVSS.t186 0.03326
R61587 DVSS.n266 DVSS.t110 0.03326
R61588 DVSS.n246 DVSS.t160 0.03326
R61589 DVSS.n246 DVSS.t130 0.03326
R61590 DVSS.n6443 DVSS.t172 0.03326
R61591 DVSS.n6443 DVSS.t148 0.03326
R61592 DVSS.n212 DVSS.n209 0.0329
R61593 DVSS.n3506 DVSS.n3505 0.0329
R61594 DVSS.n3513 DVSS.n2139 0.0329
R61595 DVSS.n208 DVSS.n184 0.0329
R61596 DVSS.n123 DVSS.n111 0.0329
R61597 DVSS.n225 DVSS.n221 0.0329
R61598 DVSS.n4425 DVSS.n3955 0.0313152
R61599 DVSS.n5506 DVSS.n1370 0.0313152
R61600 DVSS.n4333 DVSS.n4332 0.0313152
R61601 DVSS.n5349 DVSS.n1523 0.0313152
R61602 DVSS.n1075 DVSS.n1074 0.0311
R61603 DVSS.n6256 DVSS.n6255 0.0311
R61604 DVSS.n497 DVSS.n429 0.0311
R61605 DVSS.n494 DVSS.n413 0.0311
R61606 DVSS.n756 DVSS.n588 0.0304195
R61607 DVSS.n591 DVSS.n587 0.0304195
R61608 DVSS.n4949 DVSS.n1791 0.0301809
R61609 DVSS.n4970 DVSS.n4966 0.0301809
R61610 DVSS.n4952 DVSS.n1787 0.0301809
R61611 DVSS.n4975 DVSS.n1770 0.0301809
R61612 DVSS.n4433 DVSS.n2054 0.0301532
R61613 DVSS.n1762 DVSS.n1761 0.0293889
R61614 DVSS.t24 DVSS.n1762 0.0293889
R61615 DVSS.n2409 DVSS.n1766 0.0293889
R61616 DVSS.n1766 DVSS.t24 0.0293889
R61617 DVSS.n506 DVSS.n298 0.0293806
R61618 DVSS.n2601 DVSS.n2600 0.0287281
R61619 DVSS.n2886 DVSS.n2885 0.0287281
R61620 DVSS.n2884 DVSS.n2608 0.0287281
R61621 DVSS.n2876 DVSS.n2610 0.0287281
R61622 DVSS.n2877 DVSS.n2132 0.0287281
R61623 DVSS.n2879 DVSS.n2612 0.0287281
R61624 DVSS.n2878 DVSS.n1687 0.0287281
R61625 DVSS.n5086 DVSS.n1685 0.0287281
R61626 DVSS.n5087 DVSS.n1675 0.0287281
R61627 DVSS.n1680 DVSS.n1524 0.0287281
R61628 DVSS.n5346 DVSS.n5345 0.0287281
R61629 DVSS.n5508 DVSS.n1359 0.0287281
R61630 DVSS.n1364 DVSS.n1333 0.0287281
R61631 DVSS.n6070 DVSS.n6069 0.0287281
R61632 DVSS.n1187 DVSS.n1186 0.0287281
R61633 DVSS.n1196 DVSS.n1195 0.0287281
R61634 DVSS.n1193 DVSS.n1191 0.0287281
R61635 DVSS.n27 DVSS.n26 0.0287281
R61636 DVSS.n24 DVSS.n23 0.0287281
R61637 DVSS.n6393 DVSS.n259 0.0287281
R61638 DVSS.n1194 DVSS.n1193 0.0287281
R61639 DVSS.n6069 DVSS.n1182 0.0287281
R61640 DVSS.n1548 DVSS.n1369 0.0287281
R61641 DVSS.n3053 DVSS.n3052 0.0287281
R61642 DVSS.n3041 DVSS.n2405 0.0287281
R61643 DVSS.n3754 DVSS.n1721 0.0287281
R61644 DVSS.n5165 DVSS.n1650 0.0287281
R61645 DVSS.n5263 DVSS.n5262 0.0287281
R61646 DVSS.n5586 DVSS.n1334 0.0287281
R61647 DVSS.n6050 DVSS.n1179 0.0287281
R61648 DVSS.n5805 DVSS.n5801 0.0287281
R61649 DVSS.n384 DVSS.n361 0.0287281
R61650 DVSS.n382 DVSS.n359 0.0287281
R61651 DVSS.n6382 DVSS.n194 0.0287281
R61652 DVSS.n4971 DVSS.n1772 0.0287281
R61653 DVSS.n4973 DVSS.n1771 0.0287281
R61654 DVSS.n4974 DVSS.n4972 0.0287281
R61655 DVSS.n4969 DVSS.n4968 0.0287281
R61656 DVSS.n6053 DVSS.n5801 0.0287281
R61657 DVSS.n5803 DVSS.n5800 0.0287281
R61658 DVSS.n6048 DVSS.n5807 0.0287281
R61659 DVSS.n6051 DVSS.n6050 0.0287281
R61660 DVSS.n4702 DVSS.n1336 0.0287281
R61661 DVSS.n3755 DVSS.n1652 0.0287281
R61662 DVSS.n1731 DVSS.n1721 0.0287281
R61663 DVSS.n1722 DVSS.n1718 0.0287281
R61664 DVSS.n1727 DVSS.n1726 0.0287281
R61665 DVSS.n2403 DVSS.n2128 0.0287281
R61666 DVSS.n3046 DVSS.n3045 0.0287281
R61667 DVSS.n3051 DVSS.n3050 0.0287281
R61668 DVSS.n3061 DVSS.n3060 0.0287281
R61669 DVSS.n5166 DVSS.n1569 0.0287281
R61670 DVSS.n3020 DVSS.n2434 0.0287281
R61671 DVSS.n3027 DVSS.n2424 0.0287281
R61672 DVSS.n3031 DVSS.n3029 0.0287281
R61673 DVSS.n4927 DVSS.n4926 0.0287281
R61674 DVSS.n4915 DVSS.n4914 0.0287281
R61675 DVSS.n4640 DVSS.n2026 0.0287281
R61676 DVSS.n2017 DVSS.n1298 0.0287281
R61677 DVSS.n6100 DVSS.n1144 0.0287281
R61678 DVSS.n6103 DVSS.n1142 0.0287281
R61679 DVSS.n99 DVSS.n85 0.0287281
R61680 DVSS.n97 DVSS.n78 0.0287281
R61681 DVSS.n118 DVSS.n108 0.0287281
R61682 DVSS.n3029 DVSS.n3028 0.0287281
R61683 DVSS.n4950 DVSS.n1790 0.0287281
R61684 DVSS.n3030 DVSS.n1788 0.0287281
R61685 DVSS.n4951 DVSS.n1789 0.0287281
R61686 DVSS.n4948 DVSS.n4947 0.0287281
R61687 DVSS.n1146 DVSS.n1142 0.0287281
R61688 DVSS.n6098 DVSS.n1145 0.0287281
R61689 DVSS.n1155 DVSS.n1149 0.0287281
R61690 DVSS.n6101 DVSS.n6100 0.0287281
R61691 DVSS.n4644 DVSS.n4643 0.0287281
R61692 DVSS.n4925 DVSS.n4924 0.0287281
R61693 DVSS.n4928 DVSS.n4927 0.0287281
R61694 DVSS.n4938 DVSS.n4937 0.0287281
R61695 DVSS.n4943 DVSS.n4942 0.0287281
R61696 DVSS.n2428 DVSS.n2115 0.0287281
R61697 DVSS.n3025 DVSS.n2432 0.0287281
R61698 DVSS.n3021 DVSS.n2426 0.0287281
R61699 DVSS.n3013 DVSS.n2440 0.0287281
R61700 DVSS.n4638 DVSS.n4637 0.0287281
R61701 DVSS.n2469 DVSS.n2458 0.0287281
R61702 DVSS.n3544 DVSS.n2097 0.0287281
R61703 DVSS.n3693 DVSS.n2083 0.0287281
R61704 DVSS.n3884 DVSS.n2069 0.0287281
R61705 DVSS.n4444 DVSS.n2057 0.0287281
R61706 DVSS.n3943 DVSS.n3942 0.0287281
R61707 DVSS.n6091 DVSS.n1160 0.0287281
R61708 DVSS.n1158 DVSS.n1140 0.0287281
R61709 DVSS.n70 DVSS.n57 0.0287281
R61710 DVSS.n68 DVSS.n55 0.0287281
R61711 DVSS.n243 DVSS.n242 0.0287281
R61712 DVSS.n6094 DVSS.n1158 0.0287281
R61713 DVSS.n1161 DVSS.n1157 0.0287281
R61714 DVSS.n6089 DVSS.n1164 0.0287281
R61715 DVSS.n6092 DVSS.n6091 0.0287281
R61716 DVSS.n3953 DVSS.n3952 0.0287281
R61717 DVSS.n3694 DVSS.n2071 0.0287281
R61718 DVSS.n3545 DVSS.n2085 0.0287281
R61719 DVSS.n3539 DVSS.n2102 0.0287281
R61720 DVSS.n3542 DVSS.n2105 0.0287281
R61721 DVSS.n2107 DVSS.n2099 0.0287281
R61722 DVSS.n2465 DVSS.n2462 0.0287281
R61723 DVSS.n4447 DVSS.n4446 0.0287281
R61724 DVSS.n242 DVSS.n240 0.0287281
R61725 DVSS.n239 DVSS.n238 0.0287281
R61726 DVSS.n245 DVSS.n244 0.0287281
R61727 DVSS.n236 DVSS.n235 0.0287281
R61728 DVSS.n6412 DVSS.n6411 0.0287281
R61729 DVSS.n233 DVSS.n232 0.0287281
R61730 DVSS.n6417 DVSS.n6416 0.0287281
R61731 DVSS.n230 DVSS.n229 0.0287281
R61732 DVSS.n6420 DVSS.n6419 0.0287281
R61733 DVSS.n6473 DVSS.n108 0.0287281
R61734 DVSS.n133 DVSS.n119 0.0287281
R61735 DVSS.n135 DVSS.n116 0.0287281
R61736 DVSS.n131 DVSS.n120 0.0287281
R61737 DVSS.n136 DVSS.n115 0.0287281
R61738 DVSS.n129 DVSS.n121 0.0287281
R61739 DVSS.n137 DVSS.n114 0.0287281
R61740 DVSS.n127 DVSS.n122 0.0287281
R61741 DVSS.n6469 DVSS.n112 0.0287281
R61742 DVSS.n280 DVSS.n194 0.0287281
R61743 DVSS.n204 DVSS.n192 0.0287281
R61744 DVSS.n203 DVSS.n195 0.0287281
R61745 DVSS.n205 DVSS.n190 0.0287281
R61746 DVSS.n202 DVSS.n196 0.0287281
R61747 DVSS.n206 DVSS.n188 0.0287281
R61748 DVSS.n201 DVSS.n181 0.0287281
R61749 DVSS.n6440 DVSS.n182 0.0287281
R61750 DVSS.n199 DVSS.n197 0.0287281
R61751 DVSS.n6381 DVSS.n259 0.0287281
R61752 DVSS.n6394 DVSS.n257 0.0287281
R61753 DVSS.n278 DVSS.n270 0.0287281
R61754 DVSS.n6395 DVSS.n255 0.0287281
R61755 DVSS.n277 DVSS.n247 0.0287281
R61756 DVSS.n6401 DVSS.n248 0.0287281
R61757 DVSS.n276 DVSS.n271 0.0287281
R61758 DVSS.n6396 DVSS.n252 0.0287281
R61759 DVSS.n274 DVSS.n211 0.0287281
R61760 DVSS.n72 DVSS.n61 0.0287281
R61761 DVSS.n74 DVSS.n59 0.0287281
R61762 DVSS.n75 DVSS.n58 0.0287281
R61763 DVSS.n76 DVSS.n56 0.0287281
R61764 DVSS.n6484 DVSS.n54 0.0287281
R61765 DVSS.n67 DVSS.n63 0.0287281
R61766 DVSS.n6485 DVSS.n53 0.0287281
R61767 DVSS.n66 DVSS.n48 0.0287281
R61768 DVSS.n6490 DVSS.n49 0.0287281
R61769 DVSS.n6488 DVSS.n6487 0.0287281
R61770 DVSS.n103 DVSS.n87 0.0287281
R61771 DVSS.n101 DVSS.n90 0.0287281
R61772 DVSS.n100 DVSS.n91 0.0287281
R61773 DVSS.n98 DVSS.n92 0.0287281
R61774 DVSS.n6480 DVSS.n79 0.0287281
R61775 DVSS.n105 DVSS.n83 0.0287281
R61776 DVSS.n96 DVSS.n93 0.0287281
R61777 DVSS.n106 DVSS.n82 0.0287281
R61778 DVSS.n6478 DVSS.n6477 0.0287281
R61779 DVSS.n6475 DVSS.n81 0.0287281
R61780 DVSS.n6259 DVSS.n364 0.0287281
R61781 DVSS.n6261 DVSS.n363 0.0287281
R61782 DVSS.n6273 DVSS.n362 0.0287281
R61783 DVSS.n6284 DVSS.n360 0.0287281
R61784 DVSS.n6291 DVSS.n358 0.0287281
R61785 DVSS.n381 DVSS.n378 0.0287281
R61786 DVSS.n6292 DVSS.n357 0.0287281
R61787 DVSS.n380 DVSS.n379 0.0287281
R61788 DVSS.n6293 DVSS.n355 0.0287281
R61789 DVSS.n6296 DVSS.n6295 0.0287281
R61790 DVSS.n31 DVSS.n29 0.0287281
R61791 DVSS.n6262 DVSS.n34 0.0287281
R61792 DVSS.n36 DVSS.n35 0.0287281
R61793 DVSS.n38 DVSS.n37 0.0287281
R61794 DVSS.n40 DVSS.n39 0.0287281
R61795 DVSS.n366 DVSS.n22 0.0287281
R61796 DVSS.n367 DVSS.n42 0.0287281
R61797 DVSS.n44 DVSS.n21 0.0287281
R61798 DVSS.n6499 DVSS.n6498 0.0287281
R61799 DVSS.n279 DVSS.n20 0.0287281
R61800 DVSS.n420 DVSS.n403 0.0287281
R61801 DVSS.n417 DVSS.n411 0.0287281
R61802 DVSS.n421 DVSS.n407 0.0287281
R61803 DVSS.n416 DVSS.n398 0.0287281
R61804 DVSS.n422 DVSS.n401 0.0287281
R61805 DVSS.n415 DVSS.n410 0.0287281
R61806 DVSS.n423 DVSS.n409 0.0287281
R61807 DVSS.n414 DVSS.n399 0.0287281
R61808 DVSS.n6237 DVSS.n400 0.0287281
R61809 DVSS.n6242 DVSS.n396 0.0287281
R61810 DVSS.n6240 DVSS.n413 0.0287281
R61811 DVSS.n418 DVSS.n395 0.0287281
R61812 DVSS.n448 DVSS.n436 0.0287281
R61813 DVSS.n6227 DVSS.n433 0.0287281
R61814 DVSS.n451 DVSS.n437 0.0287281
R61815 DVSS.n444 DVSS.n432 0.0287281
R61816 DVSS.n446 DVSS.n438 0.0287281
R61817 DVSS.n454 DVSS.n431 0.0287281
R61818 DVSS.n453 DVSS.n439 0.0287281
R61819 DVSS.n445 DVSS.n430 0.0287281
R61820 DVSS.n6233 DVSS.n427 0.0287281
R61821 DVSS.n443 DVSS.n440 0.0287281
R61822 DVSS.n441 DVSS.n429 0.0287281
R61823 DVSS.n6228 DVSS.n434 0.0287281
R61824 DVSS.n6218 DVSS.n6217 0.0287281
R61825 DVSS.n6214 DVSS.n6213 0.0287281
R61826 DVSS.n6211 DVSS.n6210 0.0287281
R61827 DVSS.n1118 DVSS.n459 0.0287281
R61828 DVSS.n1121 DVSS.n1120 0.0287281
R61829 DVSS.n1124 DVSS.n1123 0.0287281
R61830 DVSS.n1127 DVSS.n1126 0.0287281
R61831 DVSS.n1130 DVSS.n1129 0.0287281
R61832 DVSS.n1132 DVSS.n1131 0.0287281
R61833 DVSS.n6251 DVSS.n6250 0.0287281
R61834 DVSS.n6255 DVSS.n6254 0.0287281
R61835 DVSS.n6215 DVSS.n391 0.0287281
R61836 DVSS.n1087 DVSS.n1085 0.0287281
R61837 DVSS.n1081 DVSS.n1080 0.0287281
R61838 DVSS.n1090 DVSS.n1088 0.0287281
R61839 DVSS.n1079 DVSS.n1078 0.0287281
R61840 DVSS.n1108 DVSS.n1092 0.0287281
R61841 DVSS.n1107 DVSS.n1077 0.0287281
R61842 DVSS.n1097 DVSS.n1094 0.0287281
R61843 DVSS.n1096 DVSS.n1076 0.0287281
R61844 DVSS.n6125 DVSS.n6124 0.0287281
R61845 DVSS.n6127 DVSS.n6126 0.0287281
R61846 DVSS.n6128 DVSS.n1075 0.0287281
R61847 DVSS.n1083 DVSS.n1082 0.0287281
R61848 DVSS.n2464 DVSS.n2463 0.0287254
R61849 DVSS.n4315 DVSS.n4314 0.0283804
R61850 DVSS.n4314 DVSS.n4067 0.0283804
R61851 DVSS.n4749 DVSS.n4748 0.0283804
R61852 DVSS.n4748 DVSS.n1883 0.0283804
R61853 DVSS.n5390 DVSS.n1371 0.0283804
R61854 DVSS.n4327 DVSS.n4002 0.0283804
R61855 DVSS.n4329 DVSS.n4002 0.0283804
R61856 DVSS.n1961 DVSS.n1931 0.0283804
R61857 DVSS.n4754 DVSS.n1931 0.0283804
R61858 DVSS.n5353 DVSS.n5352 0.0283804
R61859 DVSS.n5686 DVSS.n1249 0.0272589
R61860 DVSS.n1251 DVSS.n1234 0.0272589
R61861 DVSS.n6087 DVSS.n217 0.0272589
R61862 DVSS.n6082 DVSS.n1171 0.0272589
R61863 DVSS.n6081 DVSS.n6080 0.0272589
R61864 DVSS.n1173 DVSS.n216 0.0272589
R61865 DVSS.n6078 DVSS.n1177 0.0272589
R61866 DVSS.n6077 DVSS.n1178 0.0272589
R61867 DVSS.n6074 DVSS.n1181 0.0272589
R61868 DVSS.n6075 DVSS.n1178 0.0272589
R61869 DVSS.n1181 DVSS.n214 0.0272589
R61870 DVSS.n1175 DVSS.n216 0.0272589
R61871 DVSS.n6084 DVSS.n1171 0.0272589
R61872 DVSS.n503 DVSS.n501 0.0272589
R61873 DVSS.n505 DVSS.n491 0.0272589
R61874 DVSS.n6087 DVSS.n6086 0.0272589
R61875 DVSS.n1311 DVSS.n1308 0.026913
R61876 DVSS.n1300 DVSS.n1299 0.026913
R61877 DVSS.n5684 DVSS.n1252 0.026913
R61878 DVSS.n5682 DVSS.n1259 0.026913
R61879 DVSS.n5587 DVSS.n1260 0.026913
R61880 DVSS.n5598 DVSS.n1332 0.026913
R61881 DVSS.n2680 DVSS.n2106 0.0262332
R61882 DVSS.n3547 DVSS.n2091 0.0262332
R61883 DVSS.n3696 DVSS.n2077 0.0262332
R61884 DVSS.n3900 DVSS.n3898 0.0262332
R61885 DVSS.n5855 DVSS.n1167 0.0262332
R61886 DVSS.n4933 DVSS.n1800 0.0259955
R61887 DVSS.n5000 DVSS.n4999 0.0259955
R61888 DVSS.n1736 DVSS.n1732 0.0259955
R61889 DVSS.n5004 DVSS.n5003 0.0259955
R61890 DVSS.n3034 DVSS.n3033 0.0259955
R61891 DVSS.n3038 DVSS.n1768 0.0259955
R61892 DVSS.n5003 DVSS.n1730 0.0259955
R61893 DVSS.n3038 DVSS.n3037 0.0259955
R61894 DVSS.n3033 DVSS.n2410 0.0259955
R61895 DVSS.n4999 DVSS.n1734 0.0259955
R61896 DVSS.n5002 DVSS.n1732 0.0259955
R61897 DVSS.n1800 DVSS.n1737 0.0259955
R61898 DVSS.n6398 DVSS.n272 0.0257
R61899 DVSS.n6437 DVSS.n198 0.0257
R61900 DVSS.n6471 DVSS.n124 0.0257
R61901 DVSS.n6424 DVSS.n222 0.0257
R61902 DVSS.n1761 DVSS.n1734 0.0256351
R61903 DVSS.n1761 DVSS.n1736 0.0256351
R61904 DVSS.n2410 DVSS.n2409 0.0256351
R61905 DVSS.n2409 DVSS.n2406 0.0256351
R61906 DVSS.n4066 DVSS.n3955 0.0254457
R61907 DVSS.n5506 DVSS.n5505 0.0254457
R61908 DVSS.n4332 DVSS.n4331 0.0254457
R61909 DVSS.n5350 DVSS.n5349 0.0254457
R61910 DVSS.n5599 DVSS.n1331 0.0251695
R61911 DVSS.n5695 DVSS.n1247 0.0251695
R61912 DVSS.n1073 DVSS.n1072 0.0251695
R61913 DVSS.n5589 DVSS.n5588 0.0251695
R61914 DVSS.n5702 DVSS.n5701 0.0251695
R61915 DVSS.n6258 DVSS.n386 0.0251695
R61916 DVSS.n5703 DVSS.n5702 0.0251695
R61917 DVSS.n5697 DVSS.n1247 0.0251695
R61918 DVSS.n5654 DVSS.n5653 0.0251695
R61919 DVSS.n5721 DVSS.n1232 0.0251695
R61920 DVSS.n499 DVSS.n498 0.0251695
R61921 DVSS.n5719 DVSS.n1232 0.0251695
R61922 DVSS.n499 DVSS.n497 0.0251695
R61923 DVSS.n6256 DVSS.n386 0.0251695
R61924 DVSS.n1074 DVSS.n1073 0.0251695
R61925 DVSS.n5656 DVSS.n5655 0.0251695
R61926 DVSS.n5591 DVSS.n5590 0.0251695
R61927 DVSS.n5597 DVSS.n5596 0.0251695
R61928 DVSS.n1312 DVSS.n1307 0.0251695
R61929 DVSS.n5712 DVSS.n1230 0.0251695
R61930 DVSS.n493 DVSS.n492 0.0251695
R61931 DVSS.n1310 DVSS.n1309 0.0251695
R61932 DVSS.n5715 DVSS.n5712 0.0251695
R61933 DVSS.n494 DVSS.n493 0.0251695
R61934 DVSS.n2120 DVSS.n2119 0.0248
R61935 DVSS.n2123 DVSS.n2117 0.024575
R61936 DVSS.n272 DVSS.n209 0.0239
R61937 DVSS.n208 DVSS.n198 0.0239
R61938 DVSS.n6471 DVSS.n123 0.0239
R61939 DVSS.n222 DVSS.n221 0.0239
R61940 DVSS.n658 DVSS.n589 0.0226275
R61941 DVSS.n488 DVSS.n393 0.0209851
R61942 DVSS.n6286 DVSS.n313 0.0209851
R61943 DVSS.n6079 DVSS.n1174 0.0203134
R61944 DVSS.n369 DVSS.n314 0.0203134
R61945 DVSS.n6384 DVSS.n167 0.0203134
R61946 DVSS.n5799 DVSS.n1196 0.0203
R61947 DVSS.n6054 DVSS.n5800 0.0203
R61948 DVSS.n6098 DVSS.n6097 0.0203
R61949 DVSS.n6095 DVSS.n1157 0.0203
R61950 DVSS.n1783 DVSS.n1755 0.0202719
R61951 DVSS.n1783 DVSS.t24 0.0202719
R61952 DVSS.n4961 DVSS.n4960 0.0202719
R61953 DVSS.n4960 DVSS.t24 0.0202719
R61954 DVSS.n2418 DVSS.n2417 0.0202719
R61955 DVSS.n2417 DVSS.t24 0.0202719
R61956 DVSS.n4995 DVSS.n4994 0.0199776
R61957 DVSS.n4991 DVSS.n1742 0.0199776
R61958 DVSS.n1729 DVSS.n1718 0.01985
R61959 DVSS.n5006 DVSS.n5005 0.01985
R61960 DVSS.n4937 DVSS.n4936 0.01985
R61961 DVSS.n4935 DVSS.n4934 0.01985
R61962 DVSS.n3065 DVSS.n2396 0.0198097
R61963 DVSS.n3529 DVSS.n2124 0.0196418
R61964 DVSS.n6222 DVSS.n457 0.0196418
R61965 DVSS.n6275 DVSS.n309 0.0196418
R61966 DVSS.n2610 DVSS.n2129 0.0194
R61967 DVSS.n3045 DVSS.n2125 0.0194
R61968 DVSS.n2432 DVSS.n2112 0.0194
R61969 DVSS.n2110 DVSS.n2105 0.0194
R61970 DVSS.n4190 DVSS.n4189 0.0192079
R61971 DVSS.n3082 DVSS.n2372 0.019095
R61972 DVSS.n3090 DVSS.n3089 0.019095
R61973 DVSS.n2385 DVSS.n2378 0.019095
R61974 DVSS.n2387 DVSS.n2386 0.019095
R61975 DVSS.n2386 DVSS.n2385 0.019095
R61976 DVSS.n3089 DVSS.n2373 0.019095
R61977 DVSS.n2387 DVSS.n2373 0.019095
R61978 DVSS.n3091 DVSS.n2372 0.019095
R61979 DVSS.n3091 DVSS.n3090 0.019095
R61980 DVSS.n318 DVSS.n46 0.0189701
R61981 DVSS.n261 DVSS.n171 0.0189701
R61982 DVSS.n5500 DVSS.n5499 0.0188287
R61983 DVSS.n6201 DVSS.n6200 0.0182985
R61984 DVSS.n6264 DVSS.n305 0.0182985
R61985 DVSS.n1516 DVSS.n1512 0.0180085
R61986 DVSS.n1512 DVSS.n1511 0.0180085
R61987 DVSS.n1511 DVSS.n1507 0.0180085
R61988 DVSS.n1507 DVSS.n1506 0.0180085
R61989 DVSS.n1506 DVSS.n1502 0.0180085
R61990 DVSS.n1502 DVSS.n1501 0.0180085
R61991 DVSS.n1501 DVSS.n1497 0.0180085
R61992 DVSS.n1497 DVSS.n1496 0.0180085
R61993 DVSS.n1496 DVSS.n1492 0.0180085
R61994 DVSS.n1492 DVSS.n1491 0.0180085
R61995 DVSS.n1491 DVSS.n1487 0.0180085
R61996 DVSS.n1487 DVSS.n1486 0.0180085
R61997 DVSS.n1486 DVSS.n1482 0.0180085
R61998 DVSS.n1482 DVSS.n1481 0.0180085
R61999 DVSS.n1481 DVSS.n1477 0.0180085
R62000 DVSS.n1477 DVSS.n1476 0.0180085
R62001 DVSS.n1476 DVSS.n1472 0.0180085
R62002 DVSS.n1472 DVSS.n1471 0.0180085
R62003 DVSS.n1467 DVSS.n1466 0.0180085
R62004 DVSS.n1462 DVSS.n1461 0.0180085
R62005 DVSS.n1461 DVSS.n1457 0.0180085
R62006 DVSS.n1457 DVSS.n1456 0.0180085
R62007 DVSS.n1456 DVSS.n1452 0.0180085
R62008 DVSS.n1452 DVSS.n1451 0.0180085
R62009 DVSS.n1451 DVSS.n1447 0.0180085
R62010 DVSS.n1447 DVSS.n1446 0.0180085
R62011 DVSS.n1446 DVSS.n1442 0.0180085
R62012 DVSS.n1442 DVSS.n1441 0.0180085
R62013 DVSS.n1441 DVSS.n1437 0.0180085
R62014 DVSS.n1437 DVSS.n1436 0.0180085
R62015 DVSS.n1436 DVSS.n1432 0.0180085
R62016 DVSS.n1432 DVSS.n1431 0.0180085
R62017 DVSS.n1431 DVSS.n1427 0.0180085
R62018 DVSS.n1427 DVSS.n1426 0.0180085
R62019 DVSS.n1426 DVSS.n1422 0.0180085
R62020 DVSS.n1422 DVSS.n1421 0.0180085
R62021 DVSS.n1421 DVSS.n1417 0.0180085
R62022 DVSS.n1417 DVSS.n1416 0.0180085
R62023 DVSS.n1416 DVSS.n1380 0.0180085
R62024 DVSS.n5493 DVSS.n1381 0.0180085
R62025 DVSS.n5493 DVSS.n5492 0.0180085
R62026 DVSS.n5492 DVSS.n5363 0.0180085
R62027 DVSS.n5486 DVSS.n5363 0.0180085
R62028 DVSS.n5486 DVSS.n5485 0.0180085
R62029 DVSS.n5485 DVSS.n5365 0.0180085
R62030 DVSS.n5479 DVSS.n5365 0.0180085
R62031 DVSS.n5479 DVSS.n5478 0.0180085
R62032 DVSS.n5478 DVSS.n5367 0.0180085
R62033 DVSS.n5472 DVSS.n5367 0.0180085
R62034 DVSS.n5472 DVSS.n5471 0.0180085
R62035 DVSS.n5471 DVSS.n5369 0.0180085
R62036 DVSS.n5465 DVSS.n5369 0.0180085
R62037 DVSS.n5465 DVSS.n5464 0.0180085
R62038 DVSS.n5464 DVSS.n5371 0.0180085
R62039 DVSS.n5458 DVSS.n5371 0.0180085
R62040 DVSS.n5458 DVSS.n5457 0.0180085
R62041 DVSS.n5457 DVSS.n5373 0.0180085
R62042 DVSS.n5451 DVSS.n5373 0.0180085
R62043 DVSS.n5451 DVSS.n5450 0.0180085
R62044 DVSS.n5446 DVSS.n5445 0.0180085
R62045 DVSS.n5441 DVSS.n5440 0.0180085
R62046 DVSS.n5440 DVSS.n5378 0.0180085
R62047 DVSS.n5434 DVSS.n5378 0.0180085
R62048 DVSS.n5434 DVSS.n5433 0.0180085
R62049 DVSS.n5433 DVSS.n5380 0.0180085
R62050 DVSS.n5427 DVSS.n5380 0.0180085
R62051 DVSS.n5427 DVSS.n5426 0.0180085
R62052 DVSS.n5426 DVSS.n5382 0.0180085
R62053 DVSS.n5420 DVSS.n5382 0.0180085
R62054 DVSS.n5420 DVSS.n5419 0.0180085
R62055 DVSS.n5419 DVSS.n5384 0.0180085
R62056 DVSS.n5413 DVSS.n5384 0.0180085
R62057 DVSS.n5413 DVSS.n5412 0.0180085
R62058 DVSS.n5412 DVSS.n5386 0.0180085
R62059 DVSS.n5406 DVSS.n5386 0.0180085
R62060 DVSS.n5406 DVSS.n5405 0.0180085
R62061 DVSS.n5405 DVSS.n5388 0.0180085
R62062 DVSS.n5399 DVSS.n5388 0.0180085
R62063 DVSS.n5399 DVSS.n5398 0.0180085
R62064 DVSS.n4072 DVSS.n4069 0.0178311
R62065 DVSS.n4073 DVSS.n4072 0.0178311
R62066 DVSS.n4077 DVSS.n4073 0.0178311
R62067 DVSS.n4078 DVSS.n4077 0.0178311
R62068 DVSS.n4082 DVSS.n4078 0.0178311
R62069 DVSS.n4083 DVSS.n4082 0.0178311
R62070 DVSS.n4087 DVSS.n4083 0.0178311
R62071 DVSS.n4088 DVSS.n4087 0.0178311
R62072 DVSS.n4092 DVSS.n4088 0.0178311
R62073 DVSS.n4093 DVSS.n4092 0.0178311
R62074 DVSS.n4097 DVSS.n4093 0.0178311
R62075 DVSS.n4098 DVSS.n4097 0.0178311
R62076 DVSS.n4102 DVSS.n4098 0.0178311
R62077 DVSS.n4103 DVSS.n4102 0.0178311
R62078 DVSS.n4107 DVSS.n4103 0.0178311
R62079 DVSS.n4108 DVSS.n4107 0.0178311
R62080 DVSS.n4112 DVSS.n4108 0.0178311
R62081 DVSS.n4113 DVSS.n4112 0.0178311
R62082 DVSS.n4117 DVSS.n4113 0.0178311
R62083 DVSS.n4118 DVSS.n4117 0.0178311
R62084 DVSS.n4122 DVSS.n4118 0.0178311
R62085 DVSS.n4128 DVSS.n4124 0.0178311
R62086 DVSS.n4133 DVSS.n4129 0.0178311
R62087 DVSS.n4134 DVSS.n4133 0.0178311
R62088 DVSS.n4138 DVSS.n4134 0.0178311
R62089 DVSS.n4139 DVSS.n4138 0.0178311
R62090 DVSS.n4143 DVSS.n4139 0.0178311
R62091 DVSS.n4144 DVSS.n4143 0.0178311
R62092 DVSS.n4148 DVSS.n4144 0.0178311
R62093 DVSS.n4149 DVSS.n4148 0.0178311
R62094 DVSS.n4153 DVSS.n4149 0.0178311
R62095 DVSS.n4154 DVSS.n4153 0.0178311
R62096 DVSS.n4158 DVSS.n4154 0.0178311
R62097 DVSS.n4159 DVSS.n4158 0.0178311
R62098 DVSS.n4163 DVSS.n4159 0.0178311
R62099 DVSS.n4164 DVSS.n4163 0.0178311
R62100 DVSS.n4168 DVSS.n4164 0.0178311
R62101 DVSS.n4169 DVSS.n4168 0.0178311
R62102 DVSS.n4173 DVSS.n4169 0.0178311
R62103 DVSS.n4174 DVSS.n4173 0.0178311
R62104 DVSS.n4178 DVSS.n4174 0.0178311
R62105 DVSS.n4181 DVSS.n4178 0.0178311
R62106 DVSS.n4195 DVSS.n4191 0.0178311
R62107 DVSS.n4196 DVSS.n4195 0.0178311
R62108 DVSS.n4200 DVSS.n4196 0.0178311
R62109 DVSS.n4201 DVSS.n4200 0.0178311
R62110 DVSS.n4205 DVSS.n4201 0.0178311
R62111 DVSS.n4206 DVSS.n4205 0.0178311
R62112 DVSS.n4210 DVSS.n4206 0.0178311
R62113 DVSS.n4211 DVSS.n4210 0.0178311
R62114 DVSS.n4215 DVSS.n4211 0.0178311
R62115 DVSS.n4216 DVSS.n4215 0.0178311
R62116 DVSS.n4220 DVSS.n4216 0.0178311
R62117 DVSS.n4221 DVSS.n4220 0.0178311
R62118 DVSS.n4225 DVSS.n4221 0.0178311
R62119 DVSS.n4226 DVSS.n4225 0.0178311
R62120 DVSS.n4230 DVSS.n4226 0.0178311
R62121 DVSS.n4231 DVSS.n4230 0.0178311
R62122 DVSS.n4235 DVSS.n4231 0.0178311
R62123 DVSS.n4236 DVSS.n4235 0.0178311
R62124 DVSS.n4240 DVSS.n4236 0.0178311
R62125 DVSS.n4241 DVSS.n4240 0.0178311
R62126 DVSS.n4246 DVSS.n4245 0.0178311
R62127 DVSS.n4251 DVSS.n4250 0.0178311
R62128 DVSS.n4255 DVSS.n4251 0.0178311
R62129 DVSS.n4256 DVSS.n4255 0.0178311
R62130 DVSS.n4260 DVSS.n4256 0.0178311
R62131 DVSS.n4261 DVSS.n4260 0.0178311
R62132 DVSS.n4265 DVSS.n4261 0.0178311
R62133 DVSS.n4266 DVSS.n4265 0.0178311
R62134 DVSS.n4270 DVSS.n4266 0.0178311
R62135 DVSS.n4271 DVSS.n4270 0.0178311
R62136 DVSS.n4275 DVSS.n4271 0.0178311
R62137 DVSS.n4276 DVSS.n4275 0.0178311
R62138 DVSS.n4280 DVSS.n4276 0.0178311
R62139 DVSS.n4281 DVSS.n4280 0.0178311
R62140 DVSS.n4285 DVSS.n4281 0.0178311
R62141 DVSS.n4286 DVSS.n4285 0.0178311
R62142 DVSS.n4290 DVSS.n4286 0.0178311
R62143 DVSS.n4291 DVSS.n4290 0.0178311
R62144 DVSS.n4295 DVSS.n4291 0.0178311
R62145 DVSS.n4296 DVSS.n4295 0.0178311
R62146 DVSS.n4300 DVSS.n4296 0.0178311
R62147 DVSS.n4301 DVSS.n4300 0.0178311
R62148 DVSS.n1176 DVSS.n1172 0.0176269
R62149 DVSS.n6375 DVSS.n6374 0.0176269
R62150 DVSS.n6406 DVSS.n175 0.0176269
R62151 DVSS.n3509 DVSS.n1278 0.0171667
R62152 DVSS.n3070 DVSS.n1278 0.0171667
R62153 DVSS.n5666 DVSS.n1276 0.0171667
R62154 DVSS.n5666 DVSS.n1275 0.0171667
R62155 DVSS.n5500 DVSS.n1380 0.017087
R62156 DVSS.n2122 DVSS.n2121 0.0169552
R62157 DVSS.n1110 DVSS.n471 0.0169552
R62158 DVSS.n4190 DVSS.n4181 0.0169189
R62159 DVSS.n1867 DVSS.n1861 0.0167873
R62160 DVSS.n4850 DVSS.n1873 0.0167873
R62161 DVSS.n6432 DVSS.n212 0.0167
R62162 DVSS.n6434 DVSS.n184 0.0167
R62163 DVSS.n6468 DVSS.n111 0.0167
R62164 DVSS.n6418 DVSS.n225 0.0167
R62165 DVSS.n3536 DVSS.n2109 0.0165729
R62166 DVSS.n3522 DVSS.n2130 0.0165729
R62167 DVSS.n3520 DVSS.n2130 0.0165729
R62168 DVSS.n3527 DVSS.n2126 0.0165729
R62169 DVSS.n3533 DVSS.n2113 0.0165729
R62170 DVSS.n3525 DVSS.n2126 0.0165729
R62171 DVSS.n3531 DVSS.n2113 0.0165729
R62172 DVSS.n3537 DVSS.n3536 0.0165729
R62173 DVSS.n5450 DVSS 0.0163191
R62174 DVSS.n6446 DVSS.n6445 0.0162836
R62175 DVSS.n4241 DVSS 0.0161588
R62176 DVSS.n1098 DVSS.n1096 0.0158
R62177 DVSS.n1129 DVSS.n1128 0.0158
R62178 DVSS.n1100 DVSS.n445 0.0158
R62179 DVSS.n1101 DVSS.n399 0.0158
R62180 DVSS.n1792 DVSS.n1777 0.0157916
R62181 DVSS.n4965 DVSS.n1773 0.0157916
R62182 DVSS.n1795 DVSS.n1793 0.0157916
R62183 DVSS.n4993 DVSS.n1754 0.0157916
R62184 DVSS.n4990 DVSS.n1753 0.0157916
R62185 DVSS.n4985 DVSS.n1758 0.0157916
R62186 DVSS.n2414 DVSS.n2412 0.0157916
R62187 DVSS.n2422 DVSS.n2413 0.0157916
R62188 DVSS.n4983 DVSS.n1758 0.0157916
R62189 DVSS.n4993 DVSS.n4992 0.0157916
R62190 DVSS.n4986 DVSS.n1753 0.0157916
R62191 DVSS.n4963 DVSS.n1777 0.0157916
R62192 DVSS.n2420 DVSS.n2412 0.0157916
R62193 DVSS.n2416 DVSS.n2413 0.0157916
R62194 DVSS.n1778 DVSS.n1773 0.0157916
R62195 DVSS.n4945 DVSS.n1795 0.0157916
R62196 DVSS.n5670 DVSS.n5669 0.015774
R62197 DVSS.n2379 DVSS.n1281 0.015774
R62198 DVSS.n1099 DVSS.n484 0.0156119
R62199 DVSS.n3083 DVSS.n3073 0.0155703
R62200 DVSS.n2906 DVSS.n2905 0.0154891
R62201 DVSS.n4963 DVSS.n4961 0.0153404
R62202 DVSS.n4961 DVSS.n1778 0.0153404
R62203 DVSS.n4992 DVSS.n1755 0.0153404
R62204 DVSS.n4990 DVSS.n1755 0.0153404
R62205 DVSS.n2420 DVSS.n2418 0.0153404
R62206 DVSS.n2418 DVSS.n2416 0.0153404
R62207 DVSS.n6464 DVSS.n141 0.0152761
R62208 DVSS.n4429 DVSS.n3887 0.0149101
R62209 DVSS.n4419 DVSS.n3887 0.0149101
R62210 DVSS.n4419 DVSS.n4418 0.0149101
R62211 DVSS.n4418 DVSS.n4417 0.0149101
R62212 DVSS.n4417 DVSS.n3961 0.0149101
R62213 DVSS.n4407 DVSS.n3961 0.0149101
R62214 DVSS.n4407 DVSS.n4406 0.0149101
R62215 DVSS.n4406 DVSS.n4405 0.0149101
R62216 DVSS.n4405 DVSS.n3971 0.0149101
R62217 DVSS.n4395 DVSS.n3971 0.0149101
R62218 DVSS.n4394 DVSS.n4393 0.0149101
R62219 DVSS.n4393 DVSS.n3981 0.0149101
R62220 DVSS.n4383 DVSS.n3981 0.0149101
R62221 DVSS.n4383 DVSS.n4382 0.0149101
R62222 DVSS.n4382 DVSS.n4381 0.0149101
R62223 DVSS.n4381 DVSS.n3991 0.0149101
R62224 DVSS.n4371 DVSS.n3991 0.0149101
R62225 DVSS.n4371 DVSS.n4370 0.0149101
R62226 DVSS.n4370 DVSS.n4369 0.0149101
R62227 DVSS.n4901 DVSS.n1820 0.0149101
R62228 DVSS.n4901 DVSS.n4900 0.0149101
R62229 DVSS.n4900 DVSS.n4899 0.0149101
R62230 DVSS.n4899 DVSS.n1821 0.0149101
R62231 DVSS.n4889 DVSS.n1821 0.0149101
R62232 DVSS.n4889 DVSS.n4888 0.0149101
R62233 DVSS.n4888 DVSS.n4887 0.0149101
R62234 DVSS.n4887 DVSS.n1831 0.0149101
R62235 DVSS.n4877 DVSS.n1831 0.0149101
R62236 DVSS.n4876 DVSS.n4875 0.0149101
R62237 DVSS.n4875 DVSS.n1841 0.0149101
R62238 DVSS.n4865 DVSS.n1841 0.0149101
R62239 DVSS.n4865 DVSS.n4864 0.0149101
R62240 DVSS.n4864 DVSS.n4863 0.0149101
R62241 DVSS.n4863 DVSS.n1851 0.0149101
R62242 DVSS.n4853 DVSS.n1851 0.0149101
R62243 DVSS.n4853 DVSS.n4852 0.0149101
R62244 DVSS.n4838 DVSS.n1889 0.0149101
R62245 DVSS.n4838 DVSS.n4837 0.0149101
R62246 DVSS.n4837 DVSS.n4836 0.0149101
R62247 DVSS.n4836 DVSS.n1890 0.0149101
R62248 DVSS.n4826 DVSS.n1890 0.0149101
R62249 DVSS.n4826 DVSS.n4825 0.0149101
R62250 DVSS.n4825 DVSS.n4824 0.0149101
R62251 DVSS.n4824 DVSS.n1900 0.0149101
R62252 DVSS.n4814 DVSS.n4813 0.0149101
R62253 DVSS.n4813 DVSS.n4812 0.0149101
R62254 DVSS.n4812 DVSS.n1910 0.0149101
R62255 DVSS.n4802 DVSS.n1910 0.0149101
R62256 DVSS.n4802 DVSS.n4801 0.0149101
R62257 DVSS.n4801 DVSS.n4800 0.0149101
R62258 DVSS.n4800 DVSS.n1920 0.0149101
R62259 DVSS.n4790 DVSS.n1920 0.0149101
R62260 DVSS.n4790 DVSS.n4789 0.0149101
R62261 DVSS.n5255 DVSS.n5254 0.0149101
R62262 DVSS.n5254 DVSS.n5253 0.0149101
R62263 DVSS.n5253 DVSS.n1602 0.0149101
R62264 DVSS.n5243 DVSS.n1602 0.0149101
R62265 DVSS.n5243 DVSS.n5242 0.0149101
R62266 DVSS.n5242 DVSS.n5241 0.0149101
R62267 DVSS.n5241 DVSS.n1612 0.0149101
R62268 DVSS.n5231 DVSS.n1612 0.0149101
R62269 DVSS.n5231 DVSS.n5230 0.0149101
R62270 DVSS.n5229 DVSS.n1622 0.0149101
R62271 DVSS.n5219 DVSS.n1622 0.0149101
R62272 DVSS.n5219 DVSS.n5218 0.0149101
R62273 DVSS.n5218 DVSS.n5217 0.0149101
R62274 DVSS.n5217 DVSS.n1632 0.0149101
R62275 DVSS.n5207 DVSS.n1632 0.0149101
R62276 DVSS.n5207 DVSS.n5206 0.0149101
R62277 DVSS.n5206 DVSS.n5205 0.0149101
R62278 DVSS.n5205 DVSS.n1643 0.0149101
R62279 DVSS.n1643 DVSS.n1642 0.0149101
R62280 DVSS.n4746 DVSS.n4743 0.0147724
R62281 DVSS.n5500 DVSS.n1381 0.0146297
R62282 DVSS.n4191 DVSS.n4190 0.0144865
R62283 DVSS.n2846 DVSS.n2845 0.0142903
R62284 DVSS.n5056 DVSS.n5055 0.0142903
R62285 DVSS.n5102 DVSS.n5101 0.0142903
R62286 DVSS.n5523 DVSS.n5522 0.0142903
R62287 DVSS.n5982 DVSS.n5981 0.0142903
R62288 DVSS.n1870 DVSS.n1864 0.0142781
R62289 DVSS.n4849 DVSS.n4848 0.0142781
R62290 DVSS.n2746 DVSS.n2116 0.0142687
R62291 DVSS.n1257 DVSS.n1252 0.0141679
R62292 DVSS.n1259 DVSS.n1253 0.0141679
R62293 DVSS.n1258 DVSS.n1257 0.0141679
R62294 DVSS.n5684 DVSS.n1253 0.0141679
R62295 DVSS.n6423 DVSS.n220 0.0141679
R62296 DVSS.n6466 DVSS.n138 0.0141679
R62297 DVSS.n143 DVSS.n140 0.0141679
R62298 DVSS.n145 DVSS.n143 0.0141679
R62299 DVSS.n150 DVSS.n142 0.0141679
R62300 DVSS.n147 DVSS.n142 0.0141679
R62301 DVSS.n6436 DVSS.n148 0.0141679
R62302 DVSS.n6433 DVSS.n210 0.0141679
R62303 DVSS.n6467 DVSS.n6466 0.0141679
R62304 DVSS.n6465 DVSS.n140 0.0141679
R62305 DVSS.n150 DVSS.n146 0.0141679
R62306 DVSS.n6436 DVSS.n6435 0.0141679
R62307 DVSS.n6431 DVSS.n210 0.0141679
R62308 DVSS.n146 DVSS.n145 0.0141679
R62309 DVSS.n6463 DVSS.n147 0.0141679
R62310 DVSS.n6425 DVSS.n220 0.0141679
R62311 DVSS.n4998 DVSS.n1733 0.0141007
R62312 DVSS.n5001 DVSS.n1735 0.0141007
R62313 DVSS.n252 DVSS.n180 0.014
R62314 DVSS.n6441 DVSS.n6440 0.014
R62315 DVSS.n6413 DVSS.n127 0.014
R62316 DVSS.n6415 DVSS.n230 0.014
R62317 DVSS.n6058 DVSS.n5780 0.0139328
R62318 DVSS.n1462 DVSS 0.0138618
R62319 DVSS.n4129 DVSS 0.0137264
R62320 DVSS.n3996 DVSS.n1813 0.0137065
R62321 DVSS.n5260 DVSS.n5259 0.0137065
R62322 DVSS.n4912 DVSS.n1804 0.0137065
R62323 DVSS.n5170 DVSS.n5169 0.0137065
R62324 DVSS.n4433 DVSS.n4432 0.013408
R62325 DVSS.n4789 DVSS.n4788 0.0133933
R62326 DVSS.n3290 DVSS.n3289 0.0131563
R62327 DVSS.n3291 DVSS.n3290 0.0131563
R62328 DVSS.n3285 DVSS.n3284 0.0130581
R62329 DVSS.n3079 DVSS.n3074 0.0130581
R62330 DVSS.n4852 DVSS.n4851 0.013014
R62331 DVSS.n1889 DVSS.n1872 0.013014
R62332 DVSS.n1471 DVSS.n1412 0.0127867
R62333 DVSS.n657 DVSS.n588 0.0127612
R62334 DVSS.n656 DVSS.n591 0.0127612
R62335 DVSS.n4123 DVSS.n4122 0.0126622
R62336 DVSS.n4365 DVSS.n1820 0.0126348
R62337 DVSS.n4877 DVSS 0.0126348
R62338 DVSS.n144 DVSS.n139 0.0125896
R62339 DVSS.n2614 DVSS.n2613 0.0122
R62340 DVSS.n1109 DVSS.n1107 0.0122
R62341 DVSS.n3043 DVSS.n3042 0.0122
R62342 DVSS.n1123 DVSS.n1122 0.0122
R62343 DVSS.n2431 DVSS.n2430 0.0122
R62344 DVSS.n1111 DVSS.n454 0.0122
R62345 DVSS.n3535 DVSS.n2104 0.0122
R62346 DVSS.n1112 DVSS.n410 0.0122
R62347 DVSS.n509 DVSS.n508 0.0119179
R62348 DVSS.n6462 DVSS.n6461 0.0119179
R62349 DVSS.n3517 DVSS.n3516 0.0119115
R62350 DVSS.n3086 DVSS.n3085 0.0119115
R62351 DVSS.n4814 DVSS 0.0118764
R62352 DVSS.n4367 DVSS.n4366 0.0114972
R62353 DVSS.n4787 DVSS.n1601 0.0114972
R62354 DVSS.n2982 DVSS.n2541 0.0113864
R62355 DVSS.n2542 DVSS.n2531 0.0113864
R62356 DVSS.n2540 DVSS.n2539 0.0113864
R62357 DVSS.n2543 DVSS.n2532 0.0113864
R62358 DVSS.n2538 DVSS.n2537 0.0113864
R62359 DVSS.n2544 DVSS.n2533 0.0113864
R62360 DVSS.n2536 DVSS.n2535 0.0113864
R62361 DVSS.n2545 DVSS.n2534 0.0113864
R62362 DVSS.n2757 DVSS.n2756 0.0113864
R62363 DVSS.n2759 DVSS.n2748 0.0113864
R62364 DVSS.n2755 DVSS.n2754 0.0113864
R62365 DVSS.n2760 DVSS.n2749 0.0113864
R62366 DVSS.n2764 DVSS.n2758 0.0113864
R62367 DVSS.n2751 DVSS.n2750 0.0113864
R62368 DVSS.n2762 DVSS.n2752 0.0113864
R62369 DVSS.n3035 DVSS.n2408 0.0113864
R62370 DVSS.n2421 DVSS.n2411 0.0113864
R62371 DVSS.n2419 DVSS.n2415 0.0113864
R62372 DVSS.n4964 DVSS.n1775 0.0113864
R62373 DVSS.n4962 DVSS.n1776 0.0113864
R62374 DVSS.n4988 DVSS.n4987 0.0113864
R62375 DVSS.n1749 DVSS.n1747 0.0113864
R62376 DVSS.n1751 DVSS.n1750 0.0113864
R62377 DVSS.n1746 DVSS.n1745 0.0113864
R62378 DVSS.n4997 DVSS.n1738 0.0113864
R62379 DVSS.n3804 DVSS.n1744 0.0113864
R62380 DVSS.n3805 DVSS.n3731 0.0113864
R62381 DVSS.n3803 DVSS.n3801 0.0113864
R62382 DVSS.n3802 DVSS.n3732 0.0113864
R62383 DVSS.n3800 DVSS.n3798 0.0113864
R62384 DVSS.n3799 DVSS.n3733 0.0113864
R62385 DVSS.n3797 DVSS.n3795 0.0113864
R62386 DVSS.n3796 DVSS.n3734 0.0113864
R62387 DVSS.n3794 DVSS.n3792 0.0113864
R62388 DVSS.n3793 DVSS.n3735 0.0113864
R62389 DVSS.n3791 DVSS.n3789 0.0113864
R62390 DVSS.n1868 DVSS.n1865 0.0113864
R62391 DVSS.n1871 DVSS.n1862 0.0113864
R62392 DVSS.n1869 DVSS.n1866 0.0113864
R62393 DVSS.n1875 DVSS.n1861 0.0113864
R62394 DVSS.n4595 DVSS.n4537 0.0113864
R62395 DVSS.n4538 DVSS.n4507 0.0113864
R62396 DVSS.n4536 DVSS.n4535 0.0113864
R62397 DVSS.n4539 DVSS.n4508 0.0113864
R62398 DVSS.n4534 DVSS.n4533 0.0113864
R62399 DVSS.n4540 DVSS.n4509 0.0113864
R62400 DVSS.n4532 DVSS.n4531 0.0113864
R62401 DVSS.n4541 DVSS.n4510 0.0113864
R62402 DVSS.n4530 DVSS.n4529 0.0113864
R62403 DVSS.n4542 DVSS.n4511 0.0113864
R62404 DVSS.n4528 DVSS.n4527 0.0113864
R62405 DVSS.n4543 DVSS.n4512 0.0113864
R62406 DVSS.n4526 DVSS.n4525 0.0113864
R62407 DVSS.n4544 DVSS.n4513 0.0113864
R62408 DVSS.n4524 DVSS.n4523 0.0113864
R62409 DVSS.n4545 DVSS.n4514 0.0113864
R62410 DVSS.n4522 DVSS.n4521 0.0113864
R62411 DVSS.n4546 DVSS.n4515 0.0113864
R62412 DVSS.n4520 DVSS.n4519 0.0113864
R62413 DVSS.n4547 DVSS.n4516 0.0113864
R62414 DVSS.n4518 DVSS.n4517 0.0113864
R62415 DVSS.n4548 DVSS.n1971 0.0113864
R62416 DVSS.n1975 DVSS.n1972 0.0113864
R62417 DVSS.n4741 DVSS.n1989 0.0113864
R62418 DVSS.n1990 DVSS.n1976 0.0113864
R62419 DVSS.n1987 DVSS.n1983 0.0113864
R62420 DVSS.n1991 DVSS.n1977 0.0113864
R62421 DVSS.n1986 DVSS.n1982 0.0113864
R62422 DVSS.n1992 DVSS.n1978 0.0113864
R62423 DVSS.n1985 DVSS.n1981 0.0113864
R62424 DVSS.n1993 DVSS.n1979 0.0113864
R62425 DVSS.n1984 DVSS.n1261 0.0113864
R62426 DVSS.n5774 DVSS.n1174 0.0113864
R62427 DVSS.n5791 DVSS.n5778 0.0113864
R62428 DVSS.n5797 DVSS.n5790 0.0113864
R62429 DVSS.n5789 DVSS.n5779 0.0113864
R62430 DVSS.n5796 DVSS.n5788 0.0113864
R62431 DVSS.n6059 DVSS.n5793 0.0113864
R62432 DVSS.n5795 DVSS.n5787 0.0113864
R62433 DVSS.n485 DVSS.n469 0.0113864
R62434 DVSS.n514 DVSS.n468 0.0113864
R62435 DVSS.n515 DVSS.n470 0.0113864
R62436 DVSS.n483 DVSS.n482 0.0113864
R62437 DVSS.n6191 DVSS.n487 0.0113864
R62438 DVSS.n6190 DVSS.n481 0.0113864
R62439 DVSS.n480 DVSS.n472 0.0113864
R62440 DVSS.n513 DVSS.n461 0.0113864
R62441 DVSS.n473 DVSS.n463 0.0113864
R62442 DVSS.n479 DVSS.n478 0.0113864
R62443 DVSS.n6192 DVSS.n456 0.0113864
R62444 DVSS.n6189 DVSS.n477 0.0113864
R62445 DVSS.n476 DVSS.n474 0.0113864
R62446 DVSS.n6195 DVSS.n467 0.0113864
R62447 DVSS.n6194 DVSS.n6193 0.0113864
R62448 DVSS.n512 DVSS.n489 0.0113864
R62449 DVSS.n6197 DVSS.n510 0.0113864
R62450 DVSS.n6198 DVSS.n509 0.0113864
R62451 DVSS.n301 DVSS.n300 0.0113864
R62452 DVSS.n323 DVSS.n297 0.0113864
R62453 DVSS.n303 DVSS.n302 0.0113864
R62454 DVSS.n322 DVSS.n296 0.0113864
R62455 DVSS.n304 DVSS.n294 0.0113864
R62456 DVSS.n6367 DVSS.n307 0.0113864
R62457 DVSS.n306 DVSS.n293 0.0113864
R62458 DVSS.n308 DVSS.n292 0.0113864
R62459 DVSS.n6368 DVSS.n311 0.0113864
R62460 DVSS.n310 DVSS.n291 0.0113864
R62461 DVSS.n312 DVSS.n290 0.0113864
R62462 DVSS.n6369 DVSS.n314 0.0113864
R62463 DVSS.n317 DVSS.n315 0.0113864
R62464 DVSS.n316 DVSS.n288 0.0113864
R62465 DVSS.n6370 DVSS.n318 0.0113864
R62466 DVSS.n6372 DVSS.n319 0.0113864
R62467 DVSS.n320 DVSS.n286 0.0113864
R62468 DVSS.n6374 DVSS.n282 0.0113864
R62469 DVSS.n6455 DVSS.n167 0.0113864
R62470 DVSS.n169 DVSS.n168 0.0113864
R62471 DVSS.n6453 DVSS.n163 0.0113864
R62472 DVSS.n171 DVSS.n170 0.0113864
R62473 DVSS.n173 DVSS.n172 0.0113864
R62474 DVSS.n6452 DVSS.n161 0.0113864
R62475 DVSS.n175 DVSS.n174 0.0113864
R62476 DVSS.n177 DVSS.n176 0.0113864
R62477 DVSS.n6451 DVSS.n159 0.0113864
R62478 DVSS.n6446 DVSS.n178 0.0113864
R62479 DVSS.n6448 DVSS.n6447 0.0113864
R62480 DVSS.n6450 DVSS.n157 0.0113864
R62481 DVSS.n6458 DVSS.n6449 0.0113864
R62482 DVSS.n6457 DVSS.n156 0.0113864
R62483 DVSS.n155 DVSS.n141 0.0113864
R62484 DVSS.n6459 DVSS.n151 0.0113864
R62485 DVSS.n2408 DVSS.n2407 0.0113864
R62486 DVSS.n4964 DVSS.n1776 0.0113864
R62487 DVSS.n1775 DVSS.n1774 0.0113864
R62488 DVSS.n2421 DVSS.n2415 0.0113864
R62489 DVSS.n2423 DVSS.n2411 0.0113864
R62490 DVSS.n5795 DVSS.n5780 0.0113864
R62491 DVSS.n5793 DVSS.n5788 0.0113864
R62492 DVSS.n5796 DVSS.n5779 0.0113864
R62493 DVSS.n5790 DVSS.n5789 0.0113864
R62494 DVSS.n5797 DVSS.n5778 0.0113864
R62495 DVSS.n5792 DVSS.n5791 0.0113864
R62496 DVSS.n6061 DVSS.n5774 0.0113864
R62497 DVSS.n1984 DVSS.n1979 0.0113864
R62498 DVSS.n1993 DVSS.n1981 0.0113864
R62499 DVSS.n1985 DVSS.n1978 0.0113864
R62500 DVSS.n1992 DVSS.n1982 0.0113864
R62501 DVSS.n1986 DVSS.n1977 0.0113864
R62502 DVSS.n1991 DVSS.n1983 0.0113864
R62503 DVSS.n1987 DVSS.n1976 0.0113864
R62504 DVSS.n4741 DVSS.n1990 0.0113864
R62505 DVSS.n1989 DVSS.n1975 0.0113864
R62506 DVSS.n4743 DVSS.n1972 0.0113864
R62507 DVSS.n4548 DVSS.n4518 0.0113864
R62508 DVSS.n4517 DVSS.n4516 0.0113864
R62509 DVSS.n4547 DVSS.n4520 0.0113864
R62510 DVSS.n4519 DVSS.n4515 0.0113864
R62511 DVSS.n4546 DVSS.n4522 0.0113864
R62512 DVSS.n4521 DVSS.n4514 0.0113864
R62513 DVSS.n4545 DVSS.n4524 0.0113864
R62514 DVSS.n4523 DVSS.n4513 0.0113864
R62515 DVSS.n4544 DVSS.n4526 0.0113864
R62516 DVSS.n4525 DVSS.n4512 0.0113864
R62517 DVSS.n4543 DVSS.n4528 0.0113864
R62518 DVSS.n4527 DVSS.n4511 0.0113864
R62519 DVSS.n4542 DVSS.n4530 0.0113864
R62520 DVSS.n4529 DVSS.n4510 0.0113864
R62521 DVSS.n4541 DVSS.n4532 0.0113864
R62522 DVSS.n4531 DVSS.n4509 0.0113864
R62523 DVSS.n4540 DVSS.n4534 0.0113864
R62524 DVSS.n4533 DVSS.n4508 0.0113864
R62525 DVSS.n4539 DVSS.n4536 0.0113864
R62526 DVSS.n4535 DVSS.n4507 0.0113864
R62527 DVSS.n4595 DVSS.n4538 0.0113864
R62528 DVSS.n4537 DVSS.n1873 0.0113864
R62529 DVSS.n3789 DVSS.n3735 0.0113864
R62530 DVSS.n3794 DVSS.n3793 0.0113864
R62531 DVSS.n3792 DVSS.n3734 0.0113864
R62532 DVSS.n3797 DVSS.n3796 0.0113864
R62533 DVSS.n3795 DVSS.n3733 0.0113864
R62534 DVSS.n3800 DVSS.n3799 0.0113864
R62535 DVSS.n3798 DVSS.n3732 0.0113864
R62536 DVSS.n3803 DVSS.n3802 0.0113864
R62537 DVSS.n3801 DVSS.n3731 0.0113864
R62538 DVSS.n3809 DVSS.n3805 0.0113864
R62539 DVSS.n1744 DVSS.n1735 0.0113864
R62540 DVSS.n1745 DVSS.n1738 0.0113864
R62541 DVSS.n1750 DVSS.n1746 0.0113864
R62542 DVSS.n1751 DVSS.n1749 0.0113864
R62543 DVSS.n4987 DVSS.n1747 0.0113864
R62544 DVSS.n4989 DVSS.n4988 0.0113864
R62545 DVSS.n2762 DVSS.n2751 0.0113864
R62546 DVSS.n2750 DVSS.n2124 0.0113864
R62547 DVSS.n2758 DVSS.n2749 0.0113864
R62548 DVSS.n2760 DVSS.n2755 0.0113864
R62549 DVSS.n2754 DVSS.n2748 0.0113864
R62550 DVSS.n2759 DVSS.n2757 0.0113864
R62551 DVSS.n2756 DVSS.n2747 0.0113864
R62552 DVSS.n2545 DVSS.n2536 0.0113864
R62553 DVSS.n2535 DVSS.n2533 0.0113864
R62554 DVSS.n2544 DVSS.n2538 0.0113864
R62555 DVSS.n2537 DVSS.n2532 0.0113864
R62556 DVSS.n2543 DVSS.n2540 0.0113864
R62557 DVSS.n2539 DVSS.n2531 0.0113864
R62558 DVSS.n2982 DVSS.n2542 0.0113864
R62559 DVSS.n2541 DVSS.n2397 0.0113864
R62560 DVSS.n1868 DVSS.n1863 0.0113864
R62561 DVSS.n1871 DVSS.n1865 0.0113864
R62562 DVSS.n1869 DVSS.n1862 0.0113864
R62563 DVSS.n1875 DVSS.n1866 0.0113864
R62564 DVSS.n6455 DVSS.n165 0.0113864
R62565 DVSS.n168 DVSS.n164 0.0113864
R62566 DVSS.n6453 DVSS.n169 0.0113864
R62567 DVSS.n170 DVSS.n163 0.0113864
R62568 DVSS.n172 DVSS.n162 0.0113864
R62569 DVSS.n6452 DVSS.n173 0.0113864
R62570 DVSS.n174 DVSS.n161 0.0113864
R62571 DVSS.n176 DVSS.n160 0.0113864
R62572 DVSS.n6451 DVSS.n177 0.0113864
R62573 DVSS.n178 DVSS.n159 0.0113864
R62574 DVSS.n6447 DVSS.n158 0.0113864
R62575 DVSS.n6450 DVSS.n6448 0.0113864
R62576 DVSS.n6449 DVSS.n157 0.0113864
R62577 DVSS.n6458 DVSS.n6457 0.0113864
R62578 DVSS.n156 DVSS.n155 0.0113864
R62579 DVSS.n6461 DVSS.n151 0.0113864
R62580 DVSS.n300 DVSS.n298 0.0113864
R62581 DVSS.n323 DVSS.n301 0.0113864
R62582 DVSS.n302 DVSS.n297 0.0113864
R62583 DVSS.n322 DVSS.n303 0.0113864
R62584 DVSS.n305 DVSS.n304 0.0113864
R62585 DVSS.n6367 DVSS.n294 0.0113864
R62586 DVSS.n307 DVSS.n306 0.0113864
R62587 DVSS.n309 DVSS.n308 0.0113864
R62588 DVSS.n6368 DVSS.n292 0.0113864
R62589 DVSS.n311 DVSS.n310 0.0113864
R62590 DVSS.n313 DVSS.n312 0.0113864
R62591 DVSS.n6369 DVSS.n290 0.0113864
R62592 DVSS.n315 DVSS.n289 0.0113864
R62593 DVSS.n317 DVSS.n316 0.0113864
R62594 DVSS.n6370 DVSS.n288 0.0113864
R62595 DVSS.n319 DVSS.n287 0.0113864
R62596 DVSS.n6372 DVSS.n320 0.0113864
R62597 DVSS.n286 DVSS.n282 0.0113864
R62598 DVSS.n6195 DVSS.n474 0.0113864
R62599 DVSS.n477 DVSS.n476 0.0113864
R62600 DVSS.n6189 DVSS.n457 0.0113864
R62601 DVSS.n6192 DVSS.n479 0.0113864
R62602 DVSS.n478 DVSS.n473 0.0113864
R62603 DVSS.n6200 DVSS.n463 0.0113864
R62604 DVSS.n513 DVSS.n472 0.0113864
R62605 DVSS.n481 DVSS.n480 0.0113864
R62606 DVSS.n6190 DVSS.n471 0.0113864
R62607 DVSS.n6191 DVSS.n483 0.0113864
R62608 DVSS.n482 DVSS.n470 0.0113864
R62609 DVSS.n515 DVSS.n484 0.0113864
R62610 DVSS.n514 DVSS.n469 0.0113864
R62611 DVSS.n486 DVSS.n485 0.0113864
R62612 DVSS.n6193 DVSS.n488 0.0113864
R62613 DVSS.n6194 DVSS.n489 0.0113864
R62614 DVSS.n512 DVSS.n510 0.0113864
R62615 DVSS.n6198 DVSS.n6197 0.0113864
R62616 DVSS.n3284 DVSS.n2136 0.0110469
R62617 DVSS.n6429 DVSS.n6428 0.0106562
R62618 DVSS.n6428 DVSS.n6427 0.0106562
R62619 DVSS.n2463 DVSS.n2456 0.0105
R62620 DVSS.n2475 DVSS.n2456 0.0105
R62621 DVSS.n2475 DVSS.n2454 0.0105
R62622 DVSS.n2479 DVSS.n2454 0.0105
R62623 DVSS.n2479 DVSS.n2452 0.0105
R62624 DVSS.n2483 DVSS.n2452 0.0105
R62625 DVSS.n2483 DVSS.n2450 0.0105
R62626 DVSS.n2487 DVSS.n2450 0.0105
R62627 DVSS.n2487 DVSS.n2448 0.0105
R62628 DVSS.n2491 DVSS.n2448 0.0105
R62629 DVSS.n2491 DVSS.n2446 0.0105
R62630 DVSS.n2495 DVSS.n2446 0.0105
R62631 DVSS.n2495 DVSS.n2444 0.0105
R62632 DVSS.n2499 DVSS.n2444 0.0105
R62633 DVSS.n2499 DVSS.n2442 0.0105
R62634 DVSS.n3011 DVSS.n2442 0.0105
R62635 DVSS.n3011 DVSS.n3010 0.0105
R62636 DVSS.n3010 DVSS.n3009 0.0105
R62637 DVSS.n3009 DVSS.n3008 0.0105
R62638 DVSS.n3008 DVSS.n2506 0.0105
R62639 DVSS.n3004 DVSS.n2506 0.0105
R62640 DVSS.n3004 DVSS.n3003 0.0105
R62641 DVSS.n3003 DVSS.n3002 0.0105
R62642 DVSS.n3002 DVSS.n2512 0.0105
R62643 DVSS.n2998 DVSS.n2512 0.0105
R62644 DVSS.n2998 DVSS.n2997 0.0105
R62645 DVSS.n2997 DVSS.n2996 0.0105
R62646 DVSS.n2996 DVSS.n2518 0.0105
R62647 DVSS.n2992 DVSS.n2518 0.0105
R62648 DVSS.n2992 DVSS.n2991 0.0105
R62649 DVSS.n2991 DVSS.n2990 0.0105
R62650 DVSS.n2990 DVSS.n2524 0.0105
R62651 DVSS.n2986 DVSS.n2524 0.0105
R62652 DVSS.n2986 DVSS.n2985 0.0105
R62653 DVSS.n2985 DVSS.n2529 0.0105
R62654 DVSS.n2979 DVSS.n2529 0.0105
R62655 DVSS.n2979 DVSS.n2978 0.0105
R62656 DVSS.n2978 DVSS.n2977 0.0105
R62657 DVSS.n2977 DVSS.n2553 0.0105
R62658 DVSS.n2973 DVSS.n2553 0.0105
R62659 DVSS.n2973 DVSS.n2972 0.0105
R62660 DVSS.n2972 DVSS.n2971 0.0105
R62661 DVSS.n2971 DVSS.n2559 0.0105
R62662 DVSS.n2967 DVSS.n2559 0.0105
R62663 DVSS.n2967 DVSS.n2966 0.0105
R62664 DVSS.n2966 DVSS.n2965 0.0105
R62665 DVSS.n2965 DVSS.n2565 0.0105
R62666 DVSS.n2961 DVSS.n2565 0.0105
R62667 DVSS.n2961 DVSS.n2960 0.0105
R62668 DVSS.n2960 DVSS.n2959 0.0105
R62669 DVSS.n2959 DVSS.n2956 0.0105
R62670 DVSS.n2956 DVSS.n2955 0.0105
R62671 DVSS.n2955 DVSS.n2953 0.0105
R62672 DVSS.n2953 DVSS.n2574 0.0105
R62673 DVSS.n2949 DVSS.n2574 0.0105
R62674 DVSS.n2949 DVSS.n2948 0.0105
R62675 DVSS.n2948 DVSS.n2947 0.0105
R62676 DVSS.n2947 DVSS.n2580 0.0105
R62677 DVSS.n2943 DVSS.n2580 0.0105
R62678 DVSS.n2943 DVSS.n2942 0.0105
R62679 DVSS.n2942 DVSS.n2941 0.0105
R62680 DVSS.n2941 DVSS.n2586 0.0105
R62681 DVSS.n2937 DVSS.n2586 0.0105
R62682 DVSS.n2937 DVSS.n2936 0.0105
R62683 DVSS.n2936 DVSS.n2935 0.0105
R62684 DVSS.n2935 DVSS.n2592 0.0105
R62685 DVSS.n2931 DVSS.n2592 0.0105
R62686 DVSS.n2931 DVSS.n2930 0.0105
R62687 DVSS.n2930 DVSS.n2929 0.0105
R62688 DVSS.n2929 DVSS.n2598 0.0105
R62689 DVSS.n2922 DVSS.n2598 0.0105
R62690 DVSS.n2922 DVSS.n2921 0.0105
R62691 DVSS.n2921 DVSS.n2920 0.0105
R62692 DVSS.n2920 DVSS.n2892 0.0105
R62693 DVSS.n2916 DVSS.n2892 0.0105
R62694 DVSS.n2916 DVSS.n2915 0.0105
R62695 DVSS.n2915 DVSS.n2914 0.0105
R62696 DVSS.n2914 DVSS.n2898 0.0105
R62697 DVSS.n2910 DVSS.n2898 0.0105
R62698 DVSS.n2910 DVSS.n2909 0.0105
R62699 DVSS.n2909 DVSS.n2908 0.0105
R62700 DVSS.n2474 DVSS.n2473 0.0105
R62701 DVSS.n2474 DVSS.n2453 0.0105
R62702 DVSS.n2480 DVSS.n2453 0.0105
R62703 DVSS.n2481 DVSS.n2480 0.0105
R62704 DVSS.n2482 DVSS.n2481 0.0105
R62705 DVSS.n2482 DVSS.n2449 0.0105
R62706 DVSS.n2488 DVSS.n2449 0.0105
R62707 DVSS.n2489 DVSS.n2488 0.0105
R62708 DVSS.n2490 DVSS.n2489 0.0105
R62709 DVSS.n2490 DVSS.n2445 0.0105
R62710 DVSS.n2496 DVSS.n2445 0.0105
R62711 DVSS.n2497 DVSS.n2496 0.0105
R62712 DVSS.n2498 DVSS.n2497 0.0105
R62713 DVSS.n2498 DVSS.n2441 0.0105
R62714 DVSS.n3012 DVSS.n2441 0.0105
R62715 DVSS.n3007 DVSS.n2436 0.0105
R62716 DVSS.n3007 DVSS.n3006 0.0105
R62717 DVSS.n3006 DVSS.n3005 0.0105
R62718 DVSS.n3005 DVSS.n2507 0.0105
R62719 DVSS.n3001 DVSS.n2507 0.0105
R62720 DVSS.n3001 DVSS.n3000 0.0105
R62721 DVSS.n3000 DVSS.n2999 0.0105
R62722 DVSS.n2999 DVSS.n2513 0.0105
R62723 DVSS.n2995 DVSS.n2513 0.0105
R62724 DVSS.n2995 DVSS.n2994 0.0105
R62725 DVSS.n2994 DVSS.n2993 0.0105
R62726 DVSS.n2993 DVSS.n2519 0.0105
R62727 DVSS.n2989 DVSS.n2519 0.0105
R62728 DVSS.n2989 DVSS.n2988 0.0105
R62729 DVSS.n2988 DVSS.n2987 0.0105
R62730 DVSS.n2980 DVSS.n2548 0.0105
R62731 DVSS.n2976 DVSS.n2548 0.0105
R62732 DVSS.n2976 DVSS.n2975 0.0105
R62733 DVSS.n2975 DVSS.n2974 0.0105
R62734 DVSS.n2974 DVSS.n2554 0.0105
R62735 DVSS.n2970 DVSS.n2554 0.0105
R62736 DVSS.n2970 DVSS.n2969 0.0105
R62737 DVSS.n2969 DVSS.n2968 0.0105
R62738 DVSS.n2968 DVSS.n2560 0.0105
R62739 DVSS.n2964 DVSS.n2560 0.0105
R62740 DVSS.n2964 DVSS.n2963 0.0105
R62741 DVSS.n2963 DVSS.n2962 0.0105
R62742 DVSS.n2962 DVSS.n2566 0.0105
R62743 DVSS.n2958 DVSS.n2566 0.0105
R62744 DVSS.n2958 DVSS.n2957 0.0105
R62745 DVSS.n2952 DVSS.n2951 0.0105
R62746 DVSS.n2951 DVSS.n2950 0.0105
R62747 DVSS.n2950 DVSS.n2575 0.0105
R62748 DVSS.n2946 DVSS.n2575 0.0105
R62749 DVSS.n2946 DVSS.n2945 0.0105
R62750 DVSS.n2945 DVSS.n2944 0.0105
R62751 DVSS.n2944 DVSS.n2581 0.0105
R62752 DVSS.n2940 DVSS.n2581 0.0105
R62753 DVSS.n2940 DVSS.n2939 0.0105
R62754 DVSS.n2939 DVSS.n2938 0.0105
R62755 DVSS.n2938 DVSS.n2587 0.0105
R62756 DVSS.n2934 DVSS.n2587 0.0105
R62757 DVSS.n2934 DVSS.n2933 0.0105
R62758 DVSS.n2933 DVSS.n2932 0.0105
R62759 DVSS.n2932 DVSS.n2593 0.0105
R62760 DVSS.n2924 DVSS.n2923 0.0105
R62761 DVSS.n2923 DVSS.n2887 0.0105
R62762 DVSS.n2919 DVSS.n2887 0.0105
R62763 DVSS.n2919 DVSS.n2918 0.0105
R62764 DVSS.n2918 DVSS.n2917 0.0105
R62765 DVSS.n2917 DVSS.n2893 0.0105
R62766 DVSS.n2913 DVSS.n2893 0.0105
R62767 DVSS.n2913 DVSS.n2912 0.0105
R62768 DVSS.n2912 DVSS.n2911 0.0105
R62769 DVSS.n2911 DVSS.n2899 0.0105
R62770 DVSS.n2907 DVSS.n2899 0.0105
R62771 DVSS.n1186 DVSS.n1184 0.0104
R62772 DVSS.n6402 DVSS.n6401 0.0104
R62773 DVSS.n6048 DVSS.n6047 0.0104
R62774 DVSS.n6403 DVSS.n188 0.0104
R62775 DVSS.n6083 DVSS.n1155 0.0104
R62776 DVSS.n6408 DVSS.n129 0.0104
R62777 DVSS.n6089 DVSS.n6088 0.0104
R62778 DVSS.n6410 DVSS.n233 0.0104
R62779 DVSS.n5441 DVSS.n5376 0.0103294
R62780 DVSS.n4250 DVSS.n4068 0.0102297
R62781 DVSS.n5683 DVSS.n1255 0.0100489
R62782 DVSS.n1256 DVSS.n1254 0.0100489
R62783 DVSS.n5689 DVSS.n1248 0.0100489
R62784 DVSS.n506 DVSS.n490 0.0100489
R62785 DVSS.n5687 DVSS.n1248 0.0100489
R62786 DVSS.n508 DVSS.n490 0.0100489
R62787 DVSS.n5683 DVSS.n1256 0.0100489
R62788 DVSS.n5681 DVSS.n1255 0.0100489
R62789 DVSS.n2957 DVSS.n2399 0.010007
R62790 DVSS.n6462 DVSS.n149 0.00990298
R62791 DVSS.n3019 DVSS.n2436 0.00972535
R62792 DVSS.n2681 DVSS.n2680 0.00962857
R62793 DVSS.n2683 DVSS.n2681 0.00962857
R62794 DVSS.n2683 DVSS.n2678 0.00962857
R62795 DVSS.n2687 DVSS.n2678 0.00962857
R62796 DVSS.n2687 DVSS.n2676 0.00962857
R62797 DVSS.n2691 DVSS.n2676 0.00962857
R62798 DVSS.n2691 DVSS.n2674 0.00962857
R62799 DVSS.n2695 DVSS.n2674 0.00962857
R62800 DVSS.n2695 DVSS.n2672 0.00962857
R62801 DVSS.n2699 DVSS.n2672 0.00962857
R62802 DVSS.n2699 DVSS.n2670 0.00962857
R62803 DVSS.n2703 DVSS.n2670 0.00962857
R62804 DVSS.n2703 DVSS.n2668 0.00962857
R62805 DVSS.n2708 DVSS.n2668 0.00962857
R62806 DVSS.n2708 DVSS.n2666 0.00962857
R62807 DVSS.n2712 DVSS.n2666 0.00962857
R62808 DVSS.n2713 DVSS.n2712 0.00962857
R62809 DVSS.n2714 DVSS.n2713 0.00962857
R62810 DVSS.n2714 DVSS.n2664 0.00962857
R62811 DVSS.n2718 DVSS.n2664 0.00962857
R62812 DVSS.n2718 DVSS.n2662 0.00962857
R62813 DVSS.n2722 DVSS.n2662 0.00962857
R62814 DVSS.n2722 DVSS.n2660 0.00962857
R62815 DVSS.n2726 DVSS.n2660 0.00962857
R62816 DVSS.n2726 DVSS.n2658 0.00962857
R62817 DVSS.n2730 DVSS.n2658 0.00962857
R62818 DVSS.n2730 DVSS.n2656 0.00962857
R62819 DVSS.n2734 DVSS.n2656 0.00962857
R62820 DVSS.n2734 DVSS.n2654 0.00962857
R62821 DVSS.n2738 DVSS.n2654 0.00962857
R62822 DVSS.n2738 DVSS.n2652 0.00962857
R62823 DVSS.n2742 DVSS.n2652 0.00962857
R62824 DVSS.n2742 DVSS.n2650 0.00962857
R62825 DVSS.n2767 DVSS.n2650 0.00962857
R62826 DVSS.n2767 DVSS.n2648 0.00962857
R62827 DVSS.n2771 DVSS.n2648 0.00962857
R62828 DVSS.n2771 DVSS.n2646 0.00962857
R62829 DVSS.n2775 DVSS.n2646 0.00962857
R62830 DVSS.n2775 DVSS.n2644 0.00962857
R62831 DVSS.n2779 DVSS.n2644 0.00962857
R62832 DVSS.n2779 DVSS.n2642 0.00962857
R62833 DVSS.n2783 DVSS.n2642 0.00962857
R62834 DVSS.n2783 DVSS.n2640 0.00962857
R62835 DVSS.n2787 DVSS.n2640 0.00962857
R62836 DVSS.n2787 DVSS.n2638 0.00962857
R62837 DVSS.n2791 DVSS.n2638 0.00962857
R62838 DVSS.n2791 DVSS.n2636 0.00962857
R62839 DVSS.n2795 DVSS.n2636 0.00962857
R62840 DVSS.n2795 DVSS.n2634 0.00962857
R62841 DVSS.n2800 DVSS.n2634 0.00962857
R62842 DVSS.n2800 DVSS.n2632 0.00962857
R62843 DVSS.n2804 DVSS.n2632 0.00962857
R62844 DVSS.n2805 DVSS.n2804 0.00962857
R62845 DVSS.n2807 DVSS.n2805 0.00962857
R62846 DVSS.n2807 DVSS.n2630 0.00962857
R62847 DVSS.n2811 DVSS.n2630 0.00962857
R62848 DVSS.n2811 DVSS.n2628 0.00962857
R62849 DVSS.n2815 DVSS.n2628 0.00962857
R62850 DVSS.n2815 DVSS.n2626 0.00962857
R62851 DVSS.n2819 DVSS.n2626 0.00962857
R62852 DVSS.n2819 DVSS.n2624 0.00962857
R62853 DVSS.n2823 DVSS.n2624 0.00962857
R62854 DVSS.n2823 DVSS.n2622 0.00962857
R62855 DVSS.n2827 DVSS.n2622 0.00962857
R62856 DVSS.n2827 DVSS.n2620 0.00962857
R62857 DVSS.n2831 DVSS.n2620 0.00962857
R62858 DVSS.n2831 DVSS.n2617 0.00962857
R62859 DVSS.n2874 DVSS.n2617 0.00962857
R62860 DVSS.n2874 DVSS.n2618 0.00962857
R62861 DVSS.n2870 DVSS.n2618 0.00962857
R62862 DVSS.n2870 DVSS.n2869 0.00962857
R62863 DVSS.n2869 DVSS.n2835 0.00962857
R62864 DVSS.n2865 DVSS.n2835 0.00962857
R62865 DVSS.n2865 DVSS.n2837 0.00962857
R62866 DVSS.n2861 DVSS.n2837 0.00962857
R62867 DVSS.n2861 DVSS.n2840 0.00962857
R62868 DVSS.n2857 DVSS.n2840 0.00962857
R62869 DVSS.n2857 DVSS.n2842 0.00962857
R62870 DVSS.n2853 DVSS.n2842 0.00962857
R62871 DVSS.n2853 DVSS.n2844 0.00962857
R62872 DVSS.n2849 DVSS.n2844 0.00962857
R62873 DVSS.n2682 DVSS.n2103 0.00962857
R62874 DVSS.n2682 DVSS.n2677 0.00962857
R62875 DVSS.n2688 DVSS.n2677 0.00962857
R62876 DVSS.n2689 DVSS.n2688 0.00962857
R62877 DVSS.n2690 DVSS.n2689 0.00962857
R62878 DVSS.n2690 DVSS.n2673 0.00962857
R62879 DVSS.n2696 DVSS.n2673 0.00962857
R62880 DVSS.n2697 DVSS.n2696 0.00962857
R62881 DVSS.n2698 DVSS.n2697 0.00962857
R62882 DVSS.n2698 DVSS.n2669 0.00962857
R62883 DVSS.n2704 DVSS.n2669 0.00962857
R62884 DVSS.n2705 DVSS.n2704 0.00962857
R62885 DVSS.n2707 DVSS.n2705 0.00962857
R62886 DVSS.n2707 DVSS.n2706 0.00962857
R62887 DVSS.n2706 DVSS.n2433 0.00962857
R62888 DVSS.n2663 DVSS.n2429 0.00962857
R62889 DVSS.n2719 DVSS.n2663 0.00962857
R62890 DVSS.n2720 DVSS.n2719 0.00962857
R62891 DVSS.n2721 DVSS.n2720 0.00962857
R62892 DVSS.n2721 DVSS.n2659 0.00962857
R62893 DVSS.n2727 DVSS.n2659 0.00962857
R62894 DVSS.n2728 DVSS.n2727 0.00962857
R62895 DVSS.n2729 DVSS.n2728 0.00962857
R62896 DVSS.n2729 DVSS.n2655 0.00962857
R62897 DVSS.n2735 DVSS.n2655 0.00962857
R62898 DVSS.n2736 DVSS.n2735 0.00962857
R62899 DVSS.n2737 DVSS.n2736 0.00962857
R62900 DVSS.n2737 DVSS.n2651 0.00962857
R62901 DVSS.n2743 DVSS.n2651 0.00962857
R62902 DVSS.n2744 DVSS.n2743 0.00962857
R62903 DVSS.n2773 DVSS.n2772 0.00962857
R62904 DVSS.n2774 DVSS.n2773 0.00962857
R62905 DVSS.n2774 DVSS.n2643 0.00962857
R62906 DVSS.n2780 DVSS.n2643 0.00962857
R62907 DVSS.n2781 DVSS.n2780 0.00962857
R62908 DVSS.n2782 DVSS.n2781 0.00962857
R62909 DVSS.n2782 DVSS.n2639 0.00962857
R62910 DVSS.n2788 DVSS.n2639 0.00962857
R62911 DVSS.n2789 DVSS.n2788 0.00962857
R62912 DVSS.n2790 DVSS.n2789 0.00962857
R62913 DVSS.n2790 DVSS.n2635 0.00962857
R62914 DVSS.n2796 DVSS.n2635 0.00962857
R62915 DVSS.n2797 DVSS.n2796 0.00962857
R62916 DVSS.n2799 DVSS.n2797 0.00962857
R62917 DVSS.n2799 DVSS.n2798 0.00962857
R62918 DVSS.n2806 DVSS.n2404 0.00962857
R62919 DVSS.n2806 DVSS.n2629 0.00962857
R62920 DVSS.n2812 DVSS.n2629 0.00962857
R62921 DVSS.n2813 DVSS.n2812 0.00962857
R62922 DVSS.n2814 DVSS.n2813 0.00962857
R62923 DVSS.n2814 DVSS.n2625 0.00962857
R62924 DVSS.n2820 DVSS.n2625 0.00962857
R62925 DVSS.n2821 DVSS.n2820 0.00962857
R62926 DVSS.n2822 DVSS.n2821 0.00962857
R62927 DVSS.n2822 DVSS.n2621 0.00962857
R62928 DVSS.n2828 DVSS.n2621 0.00962857
R62929 DVSS.n2829 DVSS.n2828 0.00962857
R62930 DVSS.n2830 DVSS.n2829 0.00962857
R62931 DVSS.n2830 DVSS.n2616 0.00962857
R62932 DVSS.n2875 DVSS.n2616 0.00962857
R62933 DVSS.n2868 DVSS.n2611 0.00962857
R62934 DVSS.n2868 DVSS.n2867 0.00962857
R62935 DVSS.n2867 DVSS.n2866 0.00962857
R62936 DVSS.n2866 DVSS.n2836 0.00962857
R62937 DVSS.n2860 DVSS.n2836 0.00962857
R62938 DVSS.n2860 DVSS.n2859 0.00962857
R62939 DVSS.n2859 DVSS.n2858 0.00962857
R62940 DVSS.n2858 DVSS.n2841 0.00962857
R62941 DVSS.n2852 DVSS.n2841 0.00962857
R62942 DVSS.n2852 DVSS.n2851 0.00962857
R62943 DVSS.n2851 DVSS.n2850 0.00962857
R62944 DVSS.n3690 DVSS.n2091 0.00962857
R62945 DVSS.n3690 DVSS.n2092 0.00962857
R62946 DVSS.n3686 DVSS.n2092 0.00962857
R62947 DVSS.n3686 DVSS.n3549 0.00962857
R62948 DVSS.n3682 DVSS.n3549 0.00962857
R62949 DVSS.n3682 DVSS.n3551 0.00962857
R62950 DVSS.n3678 DVSS.n3551 0.00962857
R62951 DVSS.n3678 DVSS.n3553 0.00962857
R62952 DVSS.n3674 DVSS.n3553 0.00962857
R62953 DVSS.n3674 DVSS.n3555 0.00962857
R62954 DVSS.n3670 DVSS.n3555 0.00962857
R62955 DVSS.n3670 DVSS.n3557 0.00962857
R62956 DVSS.n3666 DVSS.n3557 0.00962857
R62957 DVSS.n3666 DVSS.n3559 0.00962857
R62958 DVSS.n3662 DVSS.n3559 0.00962857
R62959 DVSS.n3662 DVSS.n3659 0.00962857
R62960 DVSS.n3659 DVSS.n3658 0.00962857
R62961 DVSS.n3658 DVSS.n3561 0.00962857
R62962 DVSS.n3653 DVSS.n3561 0.00962857
R62963 DVSS.n3653 DVSS.n3563 0.00962857
R62964 DVSS.n3649 DVSS.n3563 0.00962857
R62965 DVSS.n3649 DVSS.n3566 0.00962857
R62966 DVSS.n3645 DVSS.n3566 0.00962857
R62967 DVSS.n3645 DVSS.n3568 0.00962857
R62968 DVSS.n3641 DVSS.n3568 0.00962857
R62969 DVSS.n3641 DVSS.n3570 0.00962857
R62970 DVSS.n3637 DVSS.n3570 0.00962857
R62971 DVSS.n3637 DVSS.n3572 0.00962857
R62972 DVSS.n3633 DVSS.n3572 0.00962857
R62973 DVSS.n3633 DVSS.n3574 0.00962857
R62974 DVSS.n3629 DVSS.n3574 0.00962857
R62975 DVSS.n3629 DVSS.n3576 0.00962857
R62976 DVSS.n3625 DVSS.n3576 0.00962857
R62977 DVSS.n3625 DVSS.n3578 0.00962857
R62978 DVSS.n3621 DVSS.n3578 0.00962857
R62979 DVSS.n3621 DVSS.n3620 0.00962857
R62980 DVSS.n3620 DVSS.n3580 0.00962857
R62981 DVSS.n3616 DVSS.n3580 0.00962857
R62982 DVSS.n3616 DVSS.n3582 0.00962857
R62983 DVSS.n3612 DVSS.n3582 0.00962857
R62984 DVSS.n3612 DVSS.n3585 0.00962857
R62985 DVSS.n3608 DVSS.n3585 0.00962857
R62986 DVSS.n3608 DVSS.n3587 0.00962857
R62987 DVSS.n3604 DVSS.n3587 0.00962857
R62988 DVSS.n3604 DVSS.n3589 0.00962857
R62989 DVSS.n3600 DVSS.n3589 0.00962857
R62990 DVSS.n3600 DVSS.n3591 0.00962857
R62991 DVSS.n3596 DVSS.n3591 0.00962857
R62992 DVSS.n3596 DVSS.n3593 0.00962857
R62993 DVSS.n3593 DVSS.n1716 0.00962857
R62994 DVSS.n5009 DVSS.n1716 0.00962857
R62995 DVSS.n5009 DVSS.n1714 0.00962857
R62996 DVSS.n5013 DVSS.n1714 0.00962857
R62997 DVSS.n5013 DVSS.n1712 0.00962857
R62998 DVSS.n5017 DVSS.n1712 0.00962857
R62999 DVSS.n5017 DVSS.n1710 0.00962857
R63000 DVSS.n5021 DVSS.n1710 0.00962857
R63001 DVSS.n5021 DVSS.n1708 0.00962857
R63002 DVSS.n5025 DVSS.n1708 0.00962857
R63003 DVSS.n5025 DVSS.n1706 0.00962857
R63004 DVSS.n5029 DVSS.n1706 0.00962857
R63005 DVSS.n5029 DVSS.n1704 0.00962857
R63006 DVSS.n5033 DVSS.n1704 0.00962857
R63007 DVSS.n5033 DVSS.n1702 0.00962857
R63008 DVSS.n5037 DVSS.n1702 0.00962857
R63009 DVSS.n5037 DVSS.n1700 0.00962857
R63010 DVSS.n5041 DVSS.n1700 0.00962857
R63011 DVSS.n5041 DVSS.n1697 0.00962857
R63012 DVSS.n5083 DVSS.n1697 0.00962857
R63013 DVSS.n5083 DVSS.n1698 0.00962857
R63014 DVSS.n5079 DVSS.n1698 0.00962857
R63015 DVSS.n5079 DVSS.n5045 0.00962857
R63016 DVSS.n5075 DVSS.n5045 0.00962857
R63017 DVSS.n5075 DVSS.n5048 0.00962857
R63018 DVSS.n5071 DVSS.n5048 0.00962857
R63019 DVSS.n5071 DVSS.n5050 0.00962857
R63020 DVSS.n5067 DVSS.n5050 0.00962857
R63021 DVSS.n5067 DVSS.n5052 0.00962857
R63022 DVSS.n5063 DVSS.n5052 0.00962857
R63023 DVSS.n5063 DVSS.n5054 0.00962857
R63024 DVSS.n5059 DVSS.n5054 0.00962857
R63025 DVSS.n3691 DVSS.n2090 0.00962857
R63026 DVSS.n3685 DVSS.n2090 0.00962857
R63027 DVSS.n3685 DVSS.n3684 0.00962857
R63028 DVSS.n3684 DVSS.n3683 0.00962857
R63029 DVSS.n3683 DVSS.n3550 0.00962857
R63030 DVSS.n3677 DVSS.n3550 0.00962857
R63031 DVSS.n3677 DVSS.n3676 0.00962857
R63032 DVSS.n3676 DVSS.n3675 0.00962857
R63033 DVSS.n3675 DVSS.n3554 0.00962857
R63034 DVSS.n3669 DVSS.n3554 0.00962857
R63035 DVSS.n3669 DVSS.n3668 0.00962857
R63036 DVSS.n3668 DVSS.n3667 0.00962857
R63037 DVSS.n3667 DVSS.n3558 0.00962857
R63038 DVSS.n3661 DVSS.n3558 0.00962857
R63039 DVSS.n3661 DVSS.n3660 0.00962857
R63040 DVSS.n3652 DVSS.n3564 0.00962857
R63041 DVSS.n3652 DVSS.n3651 0.00962857
R63042 DVSS.n3651 DVSS.n3650 0.00962857
R63043 DVSS.n3650 DVSS.n3565 0.00962857
R63044 DVSS.n3644 DVSS.n3565 0.00962857
R63045 DVSS.n3644 DVSS.n3643 0.00962857
R63046 DVSS.n3643 DVSS.n3642 0.00962857
R63047 DVSS.n3642 DVSS.n3569 0.00962857
R63048 DVSS.n3636 DVSS.n3569 0.00962857
R63049 DVSS.n3636 DVSS.n3635 0.00962857
R63050 DVSS.n3635 DVSS.n3634 0.00962857
R63051 DVSS.n3634 DVSS.n3573 0.00962857
R63052 DVSS.n3628 DVSS.n3573 0.00962857
R63053 DVSS.n3628 DVSS.n3627 0.00962857
R63054 DVSS.n3627 DVSS.n3626 0.00962857
R63055 DVSS.n3619 DVSS.n3618 0.00962857
R63056 DVSS.n3618 DVSS.n3617 0.00962857
R63057 DVSS.n3617 DVSS.n3581 0.00962857
R63058 DVSS.n3611 DVSS.n3581 0.00962857
R63059 DVSS.n3611 DVSS.n3610 0.00962857
R63060 DVSS.n3610 DVSS.n3609 0.00962857
R63061 DVSS.n3609 DVSS.n3586 0.00962857
R63062 DVSS.n3603 DVSS.n3586 0.00962857
R63063 DVSS.n3603 DVSS.n3602 0.00962857
R63064 DVSS.n3602 DVSS.n3601 0.00962857
R63065 DVSS.n3601 DVSS.n3590 0.00962857
R63066 DVSS.n3595 DVSS.n3590 0.00962857
R63067 DVSS.n3595 DVSS.n3594 0.00962857
R63068 DVSS.n3594 DVSS.n1717 0.00962857
R63069 DVSS.n5008 DVSS.n1717 0.00962857
R63070 DVSS.n5015 DVSS.n5014 0.00962857
R63071 DVSS.n5016 DVSS.n5015 0.00962857
R63072 DVSS.n5016 DVSS.n1709 0.00962857
R63073 DVSS.n5022 DVSS.n1709 0.00962857
R63074 DVSS.n5023 DVSS.n5022 0.00962857
R63075 DVSS.n5024 DVSS.n5023 0.00962857
R63076 DVSS.n5024 DVSS.n1705 0.00962857
R63077 DVSS.n5030 DVSS.n1705 0.00962857
R63078 DVSS.n5031 DVSS.n5030 0.00962857
R63079 DVSS.n5032 DVSS.n5031 0.00962857
R63080 DVSS.n5032 DVSS.n1701 0.00962857
R63081 DVSS.n5038 DVSS.n1701 0.00962857
R63082 DVSS.n5039 DVSS.n5038 0.00962857
R63083 DVSS.n5040 DVSS.n5039 0.00962857
R63084 DVSS.n5040 DVSS.n1686 0.00962857
R63085 DVSS.n5078 DVSS.n5046 0.00962857
R63086 DVSS.n5078 DVSS.n5077 0.00962857
R63087 DVSS.n5077 DVSS.n5076 0.00962857
R63088 DVSS.n5076 DVSS.n5047 0.00962857
R63089 DVSS.n5070 DVSS.n5047 0.00962857
R63090 DVSS.n5070 DVSS.n5069 0.00962857
R63091 DVSS.n5069 DVSS.n5068 0.00962857
R63092 DVSS.n5068 DVSS.n5051 0.00962857
R63093 DVSS.n5062 DVSS.n5051 0.00962857
R63094 DVSS.n5062 DVSS.n5061 0.00962857
R63095 DVSS.n5061 DVSS.n5060 0.00962857
R63096 DVSS.n3881 DVSS.n2077 0.00962857
R63097 DVSS.n3881 DVSS.n2078 0.00962857
R63098 DVSS.n3877 DVSS.n2078 0.00962857
R63099 DVSS.n3877 DVSS.n3698 0.00962857
R63100 DVSS.n3873 DVSS.n3698 0.00962857
R63101 DVSS.n3873 DVSS.n3700 0.00962857
R63102 DVSS.n3869 DVSS.n3700 0.00962857
R63103 DVSS.n3869 DVSS.n3702 0.00962857
R63104 DVSS.n3865 DVSS.n3702 0.00962857
R63105 DVSS.n3865 DVSS.n3704 0.00962857
R63106 DVSS.n3861 DVSS.n3704 0.00962857
R63107 DVSS.n3861 DVSS.n3706 0.00962857
R63108 DVSS.n3857 DVSS.n3706 0.00962857
R63109 DVSS.n3857 DVSS.n3708 0.00962857
R63110 DVSS.n3853 DVSS.n3708 0.00962857
R63111 DVSS.n3853 DVSS.n3850 0.00962857
R63112 DVSS.n3850 DVSS.n3849 0.00962857
R63113 DVSS.n3849 DVSS.n3710 0.00962857
R63114 DVSS.n3844 DVSS.n3710 0.00962857
R63115 DVSS.n3844 DVSS.n3712 0.00962857
R63116 DVSS.n3840 DVSS.n3712 0.00962857
R63117 DVSS.n3840 DVSS.n3715 0.00962857
R63118 DVSS.n3836 DVSS.n3715 0.00962857
R63119 DVSS.n3836 DVSS.n3717 0.00962857
R63120 DVSS.n3832 DVSS.n3717 0.00962857
R63121 DVSS.n3832 DVSS.n3719 0.00962857
R63122 DVSS.n3828 DVSS.n3719 0.00962857
R63123 DVSS.n3828 DVSS.n3721 0.00962857
R63124 DVSS.n3824 DVSS.n3721 0.00962857
R63125 DVSS.n3824 DVSS.n3723 0.00962857
R63126 DVSS.n3820 DVSS.n3723 0.00962857
R63127 DVSS.n3820 DVSS.n3725 0.00962857
R63128 DVSS.n3816 DVSS.n3725 0.00962857
R63129 DVSS.n3816 DVSS.n3727 0.00962857
R63130 DVSS.n3812 DVSS.n3727 0.00962857
R63131 DVSS.n3812 DVSS.n3729 0.00962857
R63132 DVSS.n3786 DVSS.n3729 0.00962857
R63133 DVSS.n3786 DVSS.n3737 0.00962857
R63134 DVSS.n3782 DVSS.n3737 0.00962857
R63135 DVSS.n3782 DVSS.n3739 0.00962857
R63136 DVSS.n3778 DVSS.n3739 0.00962857
R63137 DVSS.n3778 DVSS.n3741 0.00962857
R63138 DVSS.n3774 DVSS.n3741 0.00962857
R63139 DVSS.n3774 DVSS.n3743 0.00962857
R63140 DVSS.n3770 DVSS.n3743 0.00962857
R63141 DVSS.n3770 DVSS.n3745 0.00962857
R63142 DVSS.n3766 DVSS.n3745 0.00962857
R63143 DVSS.n3766 DVSS.n3747 0.00962857
R63144 DVSS.n3762 DVSS.n3747 0.00962857
R63145 DVSS.n3762 DVSS.n3749 0.00962857
R63146 DVSS.n3758 DVSS.n3749 0.00962857
R63147 DVSS.n3758 DVSS.n1658 0.00962857
R63148 DVSS.n5162 DVSS.n1658 0.00962857
R63149 DVSS.n5162 DVSS.n1659 0.00962857
R63150 DVSS.n5158 DVSS.n1659 0.00962857
R63151 DVSS.n5158 DVSS.n1662 0.00962857
R63152 DVSS.n5154 DVSS.n1662 0.00962857
R63153 DVSS.n5154 DVSS.n1664 0.00962857
R63154 DVSS.n5150 DVSS.n1664 0.00962857
R63155 DVSS.n5150 DVSS.n1666 0.00962857
R63156 DVSS.n5146 DVSS.n1666 0.00962857
R63157 DVSS.n5146 DVSS.n1668 0.00962857
R63158 DVSS.n5142 DVSS.n1668 0.00962857
R63159 DVSS.n5142 DVSS.n1670 0.00962857
R63160 DVSS.n5138 DVSS.n1670 0.00962857
R63161 DVSS.n5138 DVSS.n1672 0.00962857
R63162 DVSS.n5134 DVSS.n1672 0.00962857
R63163 DVSS.n5134 DVSS.n1674 0.00962857
R63164 DVSS.n5129 DVSS.n1674 0.00962857
R63165 DVSS.n5129 DVSS.n5089 0.00962857
R63166 DVSS.n5125 DVSS.n5089 0.00962857
R63167 DVSS.n5125 DVSS.n5091 0.00962857
R63168 DVSS.n5121 DVSS.n5091 0.00962857
R63169 DVSS.n5121 DVSS.n5094 0.00962857
R63170 DVSS.n5117 DVSS.n5094 0.00962857
R63171 DVSS.n5117 DVSS.n5096 0.00962857
R63172 DVSS.n5113 DVSS.n5096 0.00962857
R63173 DVSS.n5113 DVSS.n5098 0.00962857
R63174 DVSS.n5109 DVSS.n5098 0.00962857
R63175 DVSS.n5109 DVSS.n5100 0.00962857
R63176 DVSS.n5105 DVSS.n5100 0.00962857
R63177 DVSS.n3882 DVSS.n2076 0.00962857
R63178 DVSS.n3876 DVSS.n2076 0.00962857
R63179 DVSS.n3876 DVSS.n3875 0.00962857
R63180 DVSS.n3875 DVSS.n3874 0.00962857
R63181 DVSS.n3874 DVSS.n3699 0.00962857
R63182 DVSS.n3868 DVSS.n3699 0.00962857
R63183 DVSS.n3868 DVSS.n3867 0.00962857
R63184 DVSS.n3867 DVSS.n3866 0.00962857
R63185 DVSS.n3866 DVSS.n3703 0.00962857
R63186 DVSS.n3860 DVSS.n3703 0.00962857
R63187 DVSS.n3860 DVSS.n3859 0.00962857
R63188 DVSS.n3859 DVSS.n3858 0.00962857
R63189 DVSS.n3858 DVSS.n3707 0.00962857
R63190 DVSS.n3852 DVSS.n3707 0.00962857
R63191 DVSS.n3852 DVSS.n3851 0.00962857
R63192 DVSS.n3843 DVSS.n3713 0.00962857
R63193 DVSS.n3843 DVSS.n3842 0.00962857
R63194 DVSS.n3842 DVSS.n3841 0.00962857
R63195 DVSS.n3841 DVSS.n3714 0.00962857
R63196 DVSS.n3835 DVSS.n3714 0.00962857
R63197 DVSS.n3835 DVSS.n3834 0.00962857
R63198 DVSS.n3834 DVSS.n3833 0.00962857
R63199 DVSS.n3833 DVSS.n3718 0.00962857
R63200 DVSS.n3827 DVSS.n3718 0.00962857
R63201 DVSS.n3827 DVSS.n3826 0.00962857
R63202 DVSS.n3826 DVSS.n3825 0.00962857
R63203 DVSS.n3825 DVSS.n3722 0.00962857
R63204 DVSS.n3819 DVSS.n3722 0.00962857
R63205 DVSS.n3819 DVSS.n3818 0.00962857
R63206 DVSS.n3818 DVSS.n3817 0.00962857
R63207 DVSS.n3788 DVSS.n3787 0.00962857
R63208 DVSS.n3787 DVSS.n3736 0.00962857
R63209 DVSS.n3781 DVSS.n3736 0.00962857
R63210 DVSS.n3781 DVSS.n3780 0.00962857
R63211 DVSS.n3780 DVSS.n3779 0.00962857
R63212 DVSS.n3779 DVSS.n3740 0.00962857
R63213 DVSS.n3773 DVSS.n3740 0.00962857
R63214 DVSS.n3773 DVSS.n3772 0.00962857
R63215 DVSS.n3772 DVSS.n3771 0.00962857
R63216 DVSS.n3771 DVSS.n3744 0.00962857
R63217 DVSS.n3765 DVSS.n3744 0.00962857
R63218 DVSS.n3765 DVSS.n3764 0.00962857
R63219 DVSS.n3764 DVSS.n3763 0.00962857
R63220 DVSS.n3763 DVSS.n3748 0.00962857
R63221 DVSS.n3757 DVSS.n3748 0.00962857
R63222 DVSS.n5163 DVSS.n1657 0.00962857
R63223 DVSS.n5157 DVSS.n1657 0.00962857
R63224 DVSS.n5157 DVSS.n5156 0.00962857
R63225 DVSS.n5156 DVSS.n5155 0.00962857
R63226 DVSS.n5155 DVSS.n1663 0.00962857
R63227 DVSS.n5149 DVSS.n1663 0.00962857
R63228 DVSS.n5149 DVSS.n5148 0.00962857
R63229 DVSS.n5148 DVSS.n5147 0.00962857
R63230 DVSS.n5147 DVSS.n1667 0.00962857
R63231 DVSS.n5141 DVSS.n1667 0.00962857
R63232 DVSS.n5141 DVSS.n5140 0.00962857
R63233 DVSS.n5140 DVSS.n5139 0.00962857
R63234 DVSS.n5139 DVSS.n1671 0.00962857
R63235 DVSS.n5133 DVSS.n1671 0.00962857
R63236 DVSS.n5133 DVSS.n5132 0.00962857
R63237 DVSS.n5124 DVSS.n5092 0.00962857
R63238 DVSS.n5124 DVSS.n5123 0.00962857
R63239 DVSS.n5123 DVSS.n5122 0.00962857
R63240 DVSS.n5122 DVSS.n5093 0.00962857
R63241 DVSS.n5116 DVSS.n5093 0.00962857
R63242 DVSS.n5116 DVSS.n5115 0.00962857
R63243 DVSS.n5115 DVSS.n5114 0.00962857
R63244 DVSS.n5114 DVSS.n5097 0.00962857
R63245 DVSS.n5108 DVSS.n5097 0.00962857
R63246 DVSS.n5108 DVSS.n5107 0.00962857
R63247 DVSS.n5107 DVSS.n5106 0.00962857
R63248 DVSS.n3939 DVSS.n3898 0.00962857
R63249 DVSS.n3939 DVSS.n3899 0.00962857
R63250 DVSS.n3935 DVSS.n3899 0.00962857
R63251 DVSS.n3935 DVSS.n3902 0.00962857
R63252 DVSS.n3931 DVSS.n3902 0.00962857
R63253 DVSS.n3931 DVSS.n3904 0.00962857
R63254 DVSS.n3927 DVSS.n3904 0.00962857
R63255 DVSS.n3927 DVSS.n3906 0.00962857
R63256 DVSS.n3923 DVSS.n3906 0.00962857
R63257 DVSS.n3923 DVSS.n3908 0.00962857
R63258 DVSS.n3919 DVSS.n3908 0.00962857
R63259 DVSS.n3919 DVSS.n3910 0.00962857
R63260 DVSS.n3915 DVSS.n3910 0.00962857
R63261 DVSS.n3915 DVSS.n3912 0.00962857
R63262 DVSS.n3912 DVSS.n2014 0.00962857
R63263 DVSS.n4647 DVSS.n2014 0.00962857
R63264 DVSS.n4647 DVSS.n2012 0.00962857
R63265 DVSS.n4651 DVSS.n2012 0.00962857
R63266 DVSS.n4651 DVSS.n2010 0.00962857
R63267 DVSS.n4655 DVSS.n2010 0.00962857
R63268 DVSS.n4655 DVSS.n2008 0.00962857
R63269 DVSS.n4659 DVSS.n2008 0.00962857
R63270 DVSS.n4659 DVSS.n2006 0.00962857
R63271 DVSS.n4663 DVSS.n2006 0.00962857
R63272 DVSS.n4663 DVSS.n2004 0.00962857
R63273 DVSS.n4667 DVSS.n2004 0.00962857
R63274 DVSS.n4667 DVSS.n2002 0.00962857
R63275 DVSS.n4671 DVSS.n2002 0.00962857
R63276 DVSS.n4671 DVSS.n2000 0.00962857
R63277 DVSS.n4675 DVSS.n2000 0.00962857
R63278 DVSS.n4675 DVSS.n1998 0.00962857
R63279 DVSS.n4680 DVSS.n1998 0.00962857
R63280 DVSS.n4680 DVSS.n1995 0.00962857
R63281 DVSS.n4738 DVSS.n1995 0.00962857
R63282 DVSS.n4738 DVSS.n1996 0.00962857
R63283 DVSS.n4734 DVSS.n1996 0.00962857
R63284 DVSS.n4734 DVSS.n4733 0.00962857
R63285 DVSS.n4733 DVSS.n4684 0.00962857
R63286 DVSS.n4729 DVSS.n4684 0.00962857
R63287 DVSS.n4729 DVSS.n4686 0.00962857
R63288 DVSS.n4725 DVSS.n4686 0.00962857
R63289 DVSS.n4725 DVSS.n4689 0.00962857
R63290 DVSS.n4721 DVSS.n4689 0.00962857
R63291 DVSS.n4721 DVSS.n4691 0.00962857
R63292 DVSS.n4717 DVSS.n4691 0.00962857
R63293 DVSS.n4717 DVSS.n4693 0.00962857
R63294 DVSS.n4713 DVSS.n4693 0.00962857
R63295 DVSS.n4713 DVSS.n4695 0.00962857
R63296 DVSS.n4709 DVSS.n4695 0.00962857
R63297 DVSS.n4709 DVSS.n4697 0.00962857
R63298 DVSS.n4705 DVSS.n4697 0.00962857
R63299 DVSS.n4705 DVSS.n1342 0.00962857
R63300 DVSS.n5583 DVSS.n1342 0.00962857
R63301 DVSS.n5583 DVSS.n1343 0.00962857
R63302 DVSS.n5579 DVSS.n1343 0.00962857
R63303 DVSS.n5579 DVSS.n1346 0.00962857
R63304 DVSS.n5575 DVSS.n1346 0.00962857
R63305 DVSS.n5575 DVSS.n1348 0.00962857
R63306 DVSS.n5571 DVSS.n1348 0.00962857
R63307 DVSS.n5571 DVSS.n1350 0.00962857
R63308 DVSS.n5567 DVSS.n1350 0.00962857
R63309 DVSS.n5567 DVSS.n1352 0.00962857
R63310 DVSS.n5563 DVSS.n1352 0.00962857
R63311 DVSS.n5563 DVSS.n1354 0.00962857
R63312 DVSS.n5559 DVSS.n1354 0.00962857
R63313 DVSS.n5559 DVSS.n1356 0.00962857
R63314 DVSS.n5555 DVSS.n1356 0.00962857
R63315 DVSS.n5555 DVSS.n1358 0.00962857
R63316 DVSS.n5550 DVSS.n1358 0.00962857
R63317 DVSS.n5550 DVSS.n5510 0.00962857
R63318 DVSS.n5546 DVSS.n5510 0.00962857
R63319 DVSS.n5546 DVSS.n5512 0.00962857
R63320 DVSS.n5542 DVSS.n5512 0.00962857
R63321 DVSS.n5542 DVSS.n5515 0.00962857
R63322 DVSS.n5538 DVSS.n5515 0.00962857
R63323 DVSS.n5538 DVSS.n5517 0.00962857
R63324 DVSS.n5534 DVSS.n5517 0.00962857
R63325 DVSS.n5534 DVSS.n5519 0.00962857
R63326 DVSS.n5530 DVSS.n5519 0.00962857
R63327 DVSS.n5530 DVSS.n5521 0.00962857
R63328 DVSS.n5526 DVSS.n5521 0.00962857
R63329 DVSS.n3940 DVSS.n3897 0.00962857
R63330 DVSS.n3934 DVSS.n3897 0.00962857
R63331 DVSS.n3934 DVSS.n3933 0.00962857
R63332 DVSS.n3933 DVSS.n3932 0.00962857
R63333 DVSS.n3932 DVSS.n3903 0.00962857
R63334 DVSS.n3926 DVSS.n3903 0.00962857
R63335 DVSS.n3926 DVSS.n3925 0.00962857
R63336 DVSS.n3925 DVSS.n3924 0.00962857
R63337 DVSS.n3924 DVSS.n3907 0.00962857
R63338 DVSS.n3918 DVSS.n3907 0.00962857
R63339 DVSS.n3918 DVSS.n3917 0.00962857
R63340 DVSS.n3917 DVSS.n3916 0.00962857
R63341 DVSS.n3916 DVSS.n3911 0.00962857
R63342 DVSS.n3911 DVSS.n2015 0.00962857
R63343 DVSS.n4646 DVSS.n2015 0.00962857
R63344 DVSS.n4653 DVSS.n4652 0.00962857
R63345 DVSS.n4654 DVSS.n4653 0.00962857
R63346 DVSS.n4654 DVSS.n2007 0.00962857
R63347 DVSS.n4660 DVSS.n2007 0.00962857
R63348 DVSS.n4661 DVSS.n4660 0.00962857
R63349 DVSS.n4662 DVSS.n4661 0.00962857
R63350 DVSS.n4662 DVSS.n2003 0.00962857
R63351 DVSS.n4668 DVSS.n2003 0.00962857
R63352 DVSS.n4669 DVSS.n4668 0.00962857
R63353 DVSS.n4670 DVSS.n4669 0.00962857
R63354 DVSS.n4670 DVSS.n1999 0.00962857
R63355 DVSS.n4676 DVSS.n1999 0.00962857
R63356 DVSS.n4677 DVSS.n4676 0.00962857
R63357 DVSS.n4679 DVSS.n4677 0.00962857
R63358 DVSS.n4679 DVSS.n4678 0.00962857
R63359 DVSS.n4732 DVSS.n1980 0.00962857
R63360 DVSS.n4732 DVSS.n4731 0.00962857
R63361 DVSS.n4731 DVSS.n4730 0.00962857
R63362 DVSS.n4730 DVSS.n4685 0.00962857
R63363 DVSS.n4724 DVSS.n4685 0.00962857
R63364 DVSS.n4724 DVSS.n4723 0.00962857
R63365 DVSS.n4723 DVSS.n4722 0.00962857
R63366 DVSS.n4722 DVSS.n4690 0.00962857
R63367 DVSS.n4716 DVSS.n4690 0.00962857
R63368 DVSS.n4716 DVSS.n4715 0.00962857
R63369 DVSS.n4715 DVSS.n4714 0.00962857
R63370 DVSS.n4714 DVSS.n4694 0.00962857
R63371 DVSS.n4708 DVSS.n4694 0.00962857
R63372 DVSS.n4708 DVSS.n4707 0.00962857
R63373 DVSS.n4707 DVSS.n4706 0.00962857
R63374 DVSS.n5584 DVSS.n1341 0.00962857
R63375 DVSS.n5578 DVSS.n1341 0.00962857
R63376 DVSS.n5578 DVSS.n5577 0.00962857
R63377 DVSS.n5577 DVSS.n5576 0.00962857
R63378 DVSS.n5576 DVSS.n1347 0.00962857
R63379 DVSS.n5570 DVSS.n1347 0.00962857
R63380 DVSS.n5570 DVSS.n5569 0.00962857
R63381 DVSS.n5569 DVSS.n5568 0.00962857
R63382 DVSS.n5568 DVSS.n1351 0.00962857
R63383 DVSS.n5562 DVSS.n1351 0.00962857
R63384 DVSS.n5562 DVSS.n5561 0.00962857
R63385 DVSS.n5561 DVSS.n5560 0.00962857
R63386 DVSS.n5560 DVSS.n1355 0.00962857
R63387 DVSS.n5554 DVSS.n1355 0.00962857
R63388 DVSS.n5554 DVSS.n5553 0.00962857
R63389 DVSS.n5545 DVSS.n5513 0.00962857
R63390 DVSS.n5545 DVSS.n5544 0.00962857
R63391 DVSS.n5544 DVSS.n5543 0.00962857
R63392 DVSS.n5543 DVSS.n5514 0.00962857
R63393 DVSS.n5537 DVSS.n5514 0.00962857
R63394 DVSS.n5537 DVSS.n5536 0.00962857
R63395 DVSS.n5536 DVSS.n5535 0.00962857
R63396 DVSS.n5535 DVSS.n5518 0.00962857
R63397 DVSS.n5529 DVSS.n5518 0.00962857
R63398 DVSS.n5529 DVSS.n5528 0.00962857
R63399 DVSS.n5528 DVSS.n5527 0.00962857
R63400 DVSS.n5857 DVSS.n5855 0.00962857
R63401 DVSS.n5858 DVSS.n5857 0.00962857
R63402 DVSS.n5861 DVSS.n5858 0.00962857
R63403 DVSS.n5861 DVSS.n5853 0.00962857
R63404 DVSS.n5865 DVSS.n5853 0.00962857
R63405 DVSS.n5865 DVSS.n5851 0.00962857
R63406 DVSS.n5869 DVSS.n5851 0.00962857
R63407 DVSS.n5869 DVSS.n5849 0.00962857
R63408 DVSS.n5873 DVSS.n5849 0.00962857
R63409 DVSS.n5873 DVSS.n5847 0.00962857
R63410 DVSS.n5877 DVSS.n5847 0.00962857
R63411 DVSS.n5877 DVSS.n5845 0.00962857
R63412 DVSS.n5882 DVSS.n5845 0.00962857
R63413 DVSS.n5882 DVSS.n5842 0.00962857
R63414 DVSS.n5886 DVSS.n5842 0.00962857
R63415 DVSS.n5887 DVSS.n5886 0.00962857
R63416 DVSS.n5888 DVSS.n5887 0.00962857
R63417 DVSS.n5888 DVSS.n5840 0.00962857
R63418 DVSS.n5892 DVSS.n5840 0.00962857
R63419 DVSS.n5892 DVSS.n5839 0.00962857
R63420 DVSS.n5896 DVSS.n5839 0.00962857
R63421 DVSS.n5896 DVSS.n5837 0.00962857
R63422 DVSS.n5900 DVSS.n5837 0.00962857
R63423 DVSS.n5900 DVSS.n5835 0.00962857
R63424 DVSS.n5904 DVSS.n5835 0.00962857
R63425 DVSS.n5904 DVSS.n5833 0.00962857
R63426 DVSS.n5908 DVSS.n5833 0.00962857
R63427 DVSS.n5908 DVSS.n5831 0.00962857
R63428 DVSS.n5912 DVSS.n5831 0.00962857
R63429 DVSS.n5912 DVSS.n5829 0.00962857
R63430 DVSS.n5916 DVSS.n5829 0.00962857
R63431 DVSS.n5916 DVSS.n5827 0.00962857
R63432 DVSS.n5920 DVSS.n5827 0.00962857
R63433 DVSS.n5920 DVSS.n5825 0.00962857
R63434 DVSS.n5924 DVSS.n5825 0.00962857
R63435 DVSS.n5925 DVSS.n5924 0.00962857
R63436 DVSS.n5927 DVSS.n5925 0.00962857
R63437 DVSS.n5927 DVSS.n5822 0.00962857
R63438 DVSS.n5931 DVSS.n5822 0.00962857
R63439 DVSS.n5931 DVSS.n5820 0.00962857
R63440 DVSS.n5935 DVSS.n5820 0.00962857
R63441 DVSS.n5935 DVSS.n5818 0.00962857
R63442 DVSS.n5939 DVSS.n5818 0.00962857
R63443 DVSS.n5939 DVSS.n5816 0.00962857
R63444 DVSS.n5943 DVSS.n5816 0.00962857
R63445 DVSS.n5943 DVSS.n5814 0.00962857
R63446 DVSS.n5947 DVSS.n5814 0.00962857
R63447 DVSS.n5947 DVSS.n5812 0.00962857
R63448 DVSS.n5951 DVSS.n5812 0.00962857
R63449 DVSS.n5951 DVSS.n5809 0.00962857
R63450 DVSS.n6043 DVSS.n5809 0.00962857
R63451 DVSS.n6043 DVSS.n5810 0.00962857
R63452 DVSS.n6039 DVSS.n5810 0.00962857
R63453 DVSS.n6039 DVSS.n6038 0.00962857
R63454 DVSS.n6038 DVSS.n5955 0.00962857
R63455 DVSS.n6034 DVSS.n5955 0.00962857
R63456 DVSS.n6034 DVSS.n5957 0.00962857
R63457 DVSS.n6030 DVSS.n5957 0.00962857
R63458 DVSS.n6030 DVSS.n5960 0.00962857
R63459 DVSS.n6026 DVSS.n5960 0.00962857
R63460 DVSS.n6026 DVSS.n5962 0.00962857
R63461 DVSS.n6022 DVSS.n5962 0.00962857
R63462 DVSS.n6022 DVSS.n5964 0.00962857
R63463 DVSS.n6018 DVSS.n5964 0.00962857
R63464 DVSS.n6018 DVSS.n5966 0.00962857
R63465 DVSS.n6014 DVSS.n5966 0.00962857
R63466 DVSS.n6014 DVSS.n5968 0.00962857
R63467 DVSS.n6010 DVSS.n5968 0.00962857
R63468 DVSS.n6010 DVSS.n5969 0.00962857
R63469 DVSS.n6006 DVSS.n5969 0.00962857
R63470 DVSS.n6006 DVSS.n6005 0.00962857
R63471 DVSS.n6005 DVSS.n5971 0.00962857
R63472 DVSS.n6001 DVSS.n5971 0.00962857
R63473 DVSS.n6001 DVSS.n5973 0.00962857
R63474 DVSS.n5997 DVSS.n5973 0.00962857
R63475 DVSS.n5997 DVSS.n5976 0.00962857
R63476 DVSS.n5993 DVSS.n5976 0.00962857
R63477 DVSS.n5993 DVSS.n5978 0.00962857
R63478 DVSS.n5989 DVSS.n5978 0.00962857
R63479 DVSS.n5989 DVSS.n5980 0.00962857
R63480 DVSS.n5985 DVSS.n5980 0.00962857
R63481 DVSS.n5859 DVSS.n1162 0.00962857
R63482 DVSS.n5860 DVSS.n5859 0.00962857
R63483 DVSS.n5860 DVSS.n5852 0.00962857
R63484 DVSS.n5866 DVSS.n5852 0.00962857
R63485 DVSS.n5867 DVSS.n5866 0.00962857
R63486 DVSS.n5868 DVSS.n5867 0.00962857
R63487 DVSS.n5868 DVSS.n5848 0.00962857
R63488 DVSS.n5874 DVSS.n5848 0.00962857
R63489 DVSS.n5875 DVSS.n5874 0.00962857
R63490 DVSS.n5876 DVSS.n5875 0.00962857
R63491 DVSS.n5876 DVSS.n5844 0.00962857
R63492 DVSS.n5883 DVSS.n5844 0.00962857
R63493 DVSS.n5884 DVSS.n5883 0.00962857
R63494 DVSS.n5885 DVSS.n5884 0.00962857
R63495 DVSS.n5885 DVSS.n1152 0.00962857
R63496 DVSS.n5893 DVSS.n1147 0.00962857
R63497 DVSS.n5894 DVSS.n5893 0.00962857
R63498 DVSS.n5895 DVSS.n5894 0.00962857
R63499 DVSS.n5895 DVSS.n5836 0.00962857
R63500 DVSS.n5901 DVSS.n5836 0.00962857
R63501 DVSS.n5902 DVSS.n5901 0.00962857
R63502 DVSS.n5903 DVSS.n5902 0.00962857
R63503 DVSS.n5903 DVSS.n5832 0.00962857
R63504 DVSS.n5909 DVSS.n5832 0.00962857
R63505 DVSS.n5910 DVSS.n5909 0.00962857
R63506 DVSS.n5911 DVSS.n5910 0.00962857
R63507 DVSS.n5911 DVSS.n5828 0.00962857
R63508 DVSS.n5917 DVSS.n5828 0.00962857
R63509 DVSS.n5918 DVSS.n5917 0.00962857
R63510 DVSS.n5919 DVSS.n5918 0.00962857
R63511 DVSS.n5926 DVSS.n5781 0.00962857
R63512 DVSS.n5926 DVSS.n5821 0.00962857
R63513 DVSS.n5932 DVSS.n5821 0.00962857
R63514 DVSS.n5933 DVSS.n5932 0.00962857
R63515 DVSS.n5934 DVSS.n5933 0.00962857
R63516 DVSS.n5934 DVSS.n5817 0.00962857
R63517 DVSS.n5940 DVSS.n5817 0.00962857
R63518 DVSS.n5941 DVSS.n5940 0.00962857
R63519 DVSS.n5942 DVSS.n5941 0.00962857
R63520 DVSS.n5942 DVSS.n5813 0.00962857
R63521 DVSS.n5948 DVSS.n5813 0.00962857
R63522 DVSS.n5949 DVSS.n5948 0.00962857
R63523 DVSS.n5950 DVSS.n5949 0.00962857
R63524 DVSS.n5950 DVSS.n5808 0.00962857
R63525 DVSS.n6044 DVSS.n5808 0.00962857
R63526 DVSS.n6037 DVSS.n5804 0.00962857
R63527 DVSS.n6037 DVSS.n6036 0.00962857
R63528 DVSS.n6036 DVSS.n6035 0.00962857
R63529 DVSS.n6035 DVSS.n5956 0.00962857
R63530 DVSS.n6029 DVSS.n5956 0.00962857
R63531 DVSS.n6029 DVSS.n6028 0.00962857
R63532 DVSS.n6028 DVSS.n6027 0.00962857
R63533 DVSS.n6027 DVSS.n5961 0.00962857
R63534 DVSS.n6021 DVSS.n5961 0.00962857
R63535 DVSS.n6021 DVSS.n6020 0.00962857
R63536 DVSS.n6020 DVSS.n6019 0.00962857
R63537 DVSS.n6019 DVSS.n5965 0.00962857
R63538 DVSS.n6013 DVSS.n5965 0.00962857
R63539 DVSS.n6013 DVSS.n6012 0.00962857
R63540 DVSS.n6012 DVSS.n6011 0.00962857
R63541 DVSS.n6004 DVSS.n1192 0.00962857
R63542 DVSS.n6004 DVSS.n6003 0.00962857
R63543 DVSS.n6003 DVSS.n6002 0.00962857
R63544 DVSS.n6002 DVSS.n5972 0.00962857
R63545 DVSS.n5996 DVSS.n5972 0.00962857
R63546 DVSS.n5996 DVSS.n5995 0.00962857
R63547 DVSS.n5995 DVSS.n5994 0.00962857
R63548 DVSS.n5994 DVSS.n5977 0.00962857
R63549 DVSS.n5988 DVSS.n5977 0.00962857
R63550 DVSS.n5988 DVSS.n5987 0.00962857
R63551 DVSS.n5987 DVSS.n5986 0.00962857
R63552 DVSS.n3499 DVSS.n2144 0.00962857
R63553 DVSS.n3499 DVSS.n2146 0.00962857
R63554 DVSS.n3495 DVSS.n2146 0.00962857
R63555 DVSS.n3495 DVSS.n2148 0.00962857
R63556 DVSS.n3491 DVSS.n2148 0.00962857
R63557 DVSS.n3491 DVSS.n2150 0.00962857
R63558 DVSS.n3487 DVSS.n2150 0.00962857
R63559 DVSS.n3487 DVSS.n2152 0.00962857
R63560 DVSS.n3483 DVSS.n2152 0.00962857
R63561 DVSS.n3483 DVSS.n2154 0.00962857
R63562 DVSS.n3479 DVSS.n2154 0.00962857
R63563 DVSS.n3479 DVSS.n2156 0.00962857
R63564 DVSS.n3475 DVSS.n2156 0.00962857
R63565 DVSS.n3475 DVSS.n2158 0.00962857
R63566 DVSS.n3471 DVSS.n2158 0.00962857
R63567 DVSS.n3471 DVSS.n2160 0.00962857
R63568 DVSS.n3467 DVSS.n2160 0.00962857
R63569 DVSS.n3467 DVSS.n2162 0.00962857
R63570 DVSS.n3463 DVSS.n2162 0.00962857
R63571 DVSS.n3463 DVSS.n2164 0.00962857
R63572 DVSS.n3459 DVSS.n2164 0.00962857
R63573 DVSS.n3459 DVSS.n2166 0.00962857
R63574 DVSS.n3455 DVSS.n2166 0.00962857
R63575 DVSS.n3455 DVSS.n2168 0.00962857
R63576 DVSS.n3451 DVSS.n2168 0.00962857
R63577 DVSS.n3451 DVSS.n2170 0.00962857
R63578 DVSS.n3447 DVSS.n2170 0.00962857
R63579 DVSS.n3447 DVSS.n2172 0.00962857
R63580 DVSS.n3443 DVSS.n2172 0.00962857
R63581 DVSS.n3443 DVSS.n2174 0.00962857
R63582 DVSS.n3439 DVSS.n2174 0.00962857
R63583 DVSS.n3439 DVSS.n2176 0.00962857
R63584 DVSS.n3435 DVSS.n2176 0.00962857
R63585 DVSS.n3435 DVSS.n2178 0.00962857
R63586 DVSS.n3431 DVSS.n2178 0.00962857
R63587 DVSS.n3431 DVSS.n2180 0.00962857
R63588 DVSS.n3427 DVSS.n2180 0.00962857
R63589 DVSS.n3427 DVSS.n2182 0.00962857
R63590 DVSS.n3423 DVSS.n2182 0.00962857
R63591 DVSS.n3423 DVSS.n2184 0.00962857
R63592 DVSS.n3419 DVSS.n2184 0.00962857
R63593 DVSS.n3419 DVSS.n2186 0.00962857
R63594 DVSS.n3415 DVSS.n2186 0.00962857
R63595 DVSS.n3415 DVSS.n2188 0.00962857
R63596 DVSS.n3411 DVSS.n2188 0.00962857
R63597 DVSS.n3411 DVSS.n2190 0.00962857
R63598 DVSS.n3407 DVSS.n2190 0.00962857
R63599 DVSS.n3407 DVSS.n2192 0.00962857
R63600 DVSS.n3403 DVSS.n2192 0.00962857
R63601 DVSS.n3403 DVSS.n2194 0.00962857
R63602 DVSS.n3399 DVSS.n2194 0.00962857
R63603 DVSS.n3399 DVSS.n2196 0.00962857
R63604 DVSS.n3395 DVSS.n2196 0.00962857
R63605 DVSS.n3395 DVSS.n2198 0.00962857
R63606 DVSS.n3391 DVSS.n2198 0.00962857
R63607 DVSS.n3391 DVSS.n2200 0.00962857
R63608 DVSS.n3387 DVSS.n2200 0.00962857
R63609 DVSS.n3387 DVSS.n2202 0.00962857
R63610 DVSS.n3383 DVSS.n2202 0.00962857
R63611 DVSS.n3383 DVSS.n2204 0.00962857
R63612 DVSS.n3379 DVSS.n2204 0.00962857
R63613 DVSS.n3379 DVSS.n2206 0.00962857
R63614 DVSS.n3375 DVSS.n2206 0.00962857
R63615 DVSS.n3375 DVSS.n2208 0.00962857
R63616 DVSS.n3371 DVSS.n2208 0.00962857
R63617 DVSS.n3371 DVSS.n2210 0.00962857
R63618 DVSS.n3367 DVSS.n2210 0.00962857
R63619 DVSS.n3367 DVSS.n2212 0.00962857
R63620 DVSS.n3363 DVSS.n2212 0.00962857
R63621 DVSS.n3363 DVSS.n2214 0.00962857
R63622 DVSS.n3359 DVSS.n2214 0.00962857
R63623 DVSS.n3359 DVSS.n2216 0.00962857
R63624 DVSS.n3355 DVSS.n2216 0.00962857
R63625 DVSS.n3355 DVSS.n2218 0.00962857
R63626 DVSS.n3351 DVSS.n2218 0.00962857
R63627 DVSS.n3351 DVSS.n2220 0.00962857
R63628 DVSS.n3347 DVSS.n2220 0.00962857
R63629 DVSS.n3347 DVSS.n2222 0.00962857
R63630 DVSS.n3343 DVSS.n2222 0.00962857
R63631 DVSS.n3343 DVSS.n2224 0.00962857
R63632 DVSS.n3339 DVSS.n2224 0.00962857
R63633 DVSS.n3339 DVSS.n2226 0.00962857
R63634 DVSS.n3335 DVSS.n2226 0.00962857
R63635 DVSS.n3335 DVSS.n2228 0.00962857
R63636 DVSS.n3331 DVSS.n2228 0.00962857
R63637 DVSS.n3331 DVSS.n2230 0.00962857
R63638 DVSS.n2275 DVSS.n2230 0.00962857
R63639 DVSS.n2275 DVSS.n2232 0.00962857
R63640 DVSS.n2271 DVSS.n2232 0.00962857
R63641 DVSS.n2271 DVSS.n2234 0.00962857
R63642 DVSS.n2267 DVSS.n2234 0.00962857
R63643 DVSS.n2267 DVSS.n2236 0.00962857
R63644 DVSS.n2263 DVSS.n2236 0.00962857
R63645 DVSS.n2263 DVSS.n2238 0.00962857
R63646 DVSS.n2259 DVSS.n2238 0.00962857
R63647 DVSS.n2259 DVSS.n2240 0.00962857
R63648 DVSS.n2255 DVSS.n2240 0.00962857
R63649 DVSS.n2252 DVSS.n2251 0.00962857
R63650 DVSS.n2251 DVSS.n2243 0.00962857
R63651 DVSS.n2247 DVSS.n2243 0.00962857
R63652 DVSS.n3099 DVSS.n2366 0.00962857
R63653 DVSS.n3099 DVSS.n2364 0.00962857
R63654 DVSS.n3103 DVSS.n2364 0.00962857
R63655 DVSS.n3103 DVSS.n2362 0.00962857
R63656 DVSS.n3107 DVSS.n2362 0.00962857
R63657 DVSS.n3107 DVSS.n2360 0.00962857
R63658 DVSS.n3111 DVSS.n2360 0.00962857
R63659 DVSS.n3111 DVSS.n2358 0.00962857
R63660 DVSS.n3115 DVSS.n2358 0.00962857
R63661 DVSS.n3115 DVSS.n2356 0.00962857
R63662 DVSS.n3119 DVSS.n2356 0.00962857
R63663 DVSS.n3119 DVSS.n2354 0.00962857
R63664 DVSS.n3123 DVSS.n2354 0.00962857
R63665 DVSS.n3123 DVSS.n2352 0.00962857
R63666 DVSS.n3127 DVSS.n2352 0.00962857
R63667 DVSS.n3127 DVSS.n2350 0.00962857
R63668 DVSS.n3131 DVSS.n2350 0.00962857
R63669 DVSS.n3131 DVSS.n2348 0.00962857
R63670 DVSS.n3135 DVSS.n2348 0.00962857
R63671 DVSS.n3135 DVSS.n2346 0.00962857
R63672 DVSS.n3139 DVSS.n2346 0.00962857
R63673 DVSS.n3139 DVSS.n2344 0.00962857
R63674 DVSS.n3143 DVSS.n2344 0.00962857
R63675 DVSS.n3143 DVSS.n2342 0.00962857
R63676 DVSS.n3147 DVSS.n2342 0.00962857
R63677 DVSS.n3147 DVSS.n2340 0.00962857
R63678 DVSS.n3151 DVSS.n2340 0.00962857
R63679 DVSS.n3151 DVSS.n2338 0.00962857
R63680 DVSS.n3155 DVSS.n2338 0.00962857
R63681 DVSS.n3155 DVSS.n2336 0.00962857
R63682 DVSS.n3159 DVSS.n2336 0.00962857
R63683 DVSS.n3159 DVSS.n2334 0.00962857
R63684 DVSS.n3163 DVSS.n2334 0.00962857
R63685 DVSS.n3163 DVSS.n2332 0.00962857
R63686 DVSS.n3167 DVSS.n2332 0.00962857
R63687 DVSS.n3167 DVSS.n2330 0.00962857
R63688 DVSS.n3171 DVSS.n2330 0.00962857
R63689 DVSS.n3171 DVSS.n2328 0.00962857
R63690 DVSS.n3175 DVSS.n2328 0.00962857
R63691 DVSS.n3175 DVSS.n2326 0.00962857
R63692 DVSS.n3179 DVSS.n2326 0.00962857
R63693 DVSS.n3179 DVSS.n2324 0.00962857
R63694 DVSS.n3183 DVSS.n2324 0.00962857
R63695 DVSS.n3183 DVSS.n2322 0.00962857
R63696 DVSS.n3187 DVSS.n2322 0.00962857
R63697 DVSS.n3187 DVSS.n2320 0.00962857
R63698 DVSS.n3191 DVSS.n2320 0.00962857
R63699 DVSS.n3191 DVSS.n2318 0.00962857
R63700 DVSS.n3195 DVSS.n2318 0.00962857
R63701 DVSS.n3195 DVSS.n2316 0.00962857
R63702 DVSS.n3199 DVSS.n2316 0.00962857
R63703 DVSS.n3199 DVSS.n2314 0.00962857
R63704 DVSS.n3203 DVSS.n2314 0.00962857
R63705 DVSS.n3203 DVSS.n2312 0.00962857
R63706 DVSS.n3207 DVSS.n2312 0.00962857
R63707 DVSS.n3207 DVSS.n2310 0.00962857
R63708 DVSS.n3211 DVSS.n2310 0.00962857
R63709 DVSS.n3211 DVSS.n2308 0.00962857
R63710 DVSS.n3215 DVSS.n2308 0.00962857
R63711 DVSS.n3215 DVSS.n2306 0.00962857
R63712 DVSS.n3219 DVSS.n2306 0.00962857
R63713 DVSS.n3219 DVSS.n2304 0.00962857
R63714 DVSS.n3223 DVSS.n2304 0.00962857
R63715 DVSS.n3223 DVSS.n2302 0.00962857
R63716 DVSS.n3227 DVSS.n2302 0.00962857
R63717 DVSS.n3227 DVSS.n2300 0.00962857
R63718 DVSS.n3231 DVSS.n2300 0.00962857
R63719 DVSS.n3231 DVSS.n2298 0.00962857
R63720 DVSS.n3235 DVSS.n2298 0.00962857
R63721 DVSS.n3235 DVSS.n2296 0.00962857
R63722 DVSS.n3239 DVSS.n2296 0.00962857
R63723 DVSS.n3239 DVSS.n2294 0.00962857
R63724 DVSS.n3243 DVSS.n2294 0.00962857
R63725 DVSS.n3243 DVSS.n2292 0.00962857
R63726 DVSS.n3247 DVSS.n2292 0.00962857
R63727 DVSS.n3247 DVSS.n2290 0.00962857
R63728 DVSS.n3251 DVSS.n2290 0.00962857
R63729 DVSS.n3251 DVSS.n2288 0.00962857
R63730 DVSS.n3255 DVSS.n2288 0.00962857
R63731 DVSS.n3255 DVSS.n2286 0.00962857
R63732 DVSS.n3259 DVSS.n2286 0.00962857
R63733 DVSS.n3259 DVSS.n2284 0.00962857
R63734 DVSS.n3263 DVSS.n2284 0.00962857
R63735 DVSS.n3263 DVSS.n2282 0.00962857
R63736 DVSS.n3267 DVSS.n2282 0.00962857
R63737 DVSS.n3267 DVSS.n2279 0.00962857
R63738 DVSS.n3325 DVSS.n2279 0.00962857
R63739 DVSS.n3325 DVSS.n2280 0.00962857
R63740 DVSS.n3321 DVSS.n2280 0.00962857
R63741 DVSS.n3321 DVSS.n3271 0.00962857
R63742 DVSS.n3317 DVSS.n3271 0.00962857
R63743 DVSS.n3317 DVSS.n3273 0.00962857
R63744 DVSS.n3313 DVSS.n3273 0.00962857
R63745 DVSS.n3313 DVSS.n3275 0.00962857
R63746 DVSS.n3309 DVSS.n3275 0.00962857
R63747 DVSS.n3309 DVSS.n3277 0.00962857
R63748 DVSS.n3305 DVSS.n3277 0.00962857
R63749 DVSS.n3302 DVSS.n3301 0.00962857
R63750 DVSS.n3301 DVSS.n3280 0.00962857
R63751 DVSS.n3297 DVSS.n3280 0.00962857
R63752 DVSS.n3097 DVSS.n3096 0.00962857
R63753 DVSS.n3098 DVSS.n3097 0.00962857
R63754 DVSS.n3098 DVSS.n2363 0.00962857
R63755 DVSS.n3104 DVSS.n2363 0.00962857
R63756 DVSS.n3105 DVSS.n3104 0.00962857
R63757 DVSS.n3106 DVSS.n3105 0.00962857
R63758 DVSS.n3106 DVSS.n2359 0.00962857
R63759 DVSS.n3112 DVSS.n2359 0.00962857
R63760 DVSS.n3113 DVSS.n3112 0.00962857
R63761 DVSS.n3114 DVSS.n3113 0.00962857
R63762 DVSS.n3114 DVSS.n2355 0.00962857
R63763 DVSS.n3120 DVSS.n2355 0.00962857
R63764 DVSS.n3121 DVSS.n3120 0.00962857
R63765 DVSS.n3122 DVSS.n3121 0.00962857
R63766 DVSS.n3122 DVSS.n2351 0.00962857
R63767 DVSS.n3128 DVSS.n2351 0.00962857
R63768 DVSS.n3129 DVSS.n3128 0.00962857
R63769 DVSS.n3130 DVSS.n3129 0.00962857
R63770 DVSS.n3130 DVSS.n2347 0.00962857
R63771 DVSS.n3136 DVSS.n2347 0.00962857
R63772 DVSS.n3137 DVSS.n3136 0.00962857
R63773 DVSS.n3138 DVSS.n3137 0.00962857
R63774 DVSS.n3138 DVSS.n2343 0.00962857
R63775 DVSS.n3144 DVSS.n2343 0.00962857
R63776 DVSS.n3145 DVSS.n3144 0.00962857
R63777 DVSS.n3146 DVSS.n3145 0.00962857
R63778 DVSS.n3146 DVSS.n2339 0.00962857
R63779 DVSS.n3152 DVSS.n2339 0.00962857
R63780 DVSS.n3153 DVSS.n3152 0.00962857
R63781 DVSS.n3154 DVSS.n3153 0.00962857
R63782 DVSS.n3154 DVSS.n2335 0.00962857
R63783 DVSS.n3160 DVSS.n2335 0.00962857
R63784 DVSS.n3161 DVSS.n3160 0.00962857
R63785 DVSS.n3162 DVSS.n3161 0.00962857
R63786 DVSS.n3162 DVSS.n2331 0.00962857
R63787 DVSS.n3168 DVSS.n2331 0.00962857
R63788 DVSS.n3169 DVSS.n3168 0.00962857
R63789 DVSS.n3170 DVSS.n3169 0.00962857
R63790 DVSS.n3170 DVSS.n2327 0.00962857
R63791 DVSS.n3176 DVSS.n2327 0.00962857
R63792 DVSS.n3177 DVSS.n3176 0.00962857
R63793 DVSS.n3178 DVSS.n3177 0.00962857
R63794 DVSS.n3178 DVSS.n2323 0.00962857
R63795 DVSS.n3184 DVSS.n2323 0.00962857
R63796 DVSS.n3185 DVSS.n3184 0.00962857
R63797 DVSS.n3186 DVSS.n3185 0.00962857
R63798 DVSS.n3186 DVSS.n2319 0.00962857
R63799 DVSS.n3192 DVSS.n2319 0.00962857
R63800 DVSS.n3193 DVSS.n3192 0.00962857
R63801 DVSS.n3194 DVSS.n3193 0.00962857
R63802 DVSS.n3194 DVSS.n2315 0.00962857
R63803 DVSS.n3200 DVSS.n2315 0.00962857
R63804 DVSS.n3201 DVSS.n3200 0.00962857
R63805 DVSS.n3202 DVSS.n3201 0.00962857
R63806 DVSS.n3202 DVSS.n2311 0.00962857
R63807 DVSS.n3208 DVSS.n2311 0.00962857
R63808 DVSS.n3209 DVSS.n3208 0.00962857
R63809 DVSS.n3210 DVSS.n3209 0.00962857
R63810 DVSS.n3210 DVSS.n2307 0.00962857
R63811 DVSS.n3216 DVSS.n2307 0.00962857
R63812 DVSS.n3217 DVSS.n3216 0.00962857
R63813 DVSS.n3218 DVSS.n3217 0.00962857
R63814 DVSS.n3218 DVSS.n2303 0.00962857
R63815 DVSS.n3224 DVSS.n2303 0.00962857
R63816 DVSS.n3225 DVSS.n3224 0.00962857
R63817 DVSS.n3226 DVSS.n3225 0.00962857
R63818 DVSS.n3226 DVSS.n2299 0.00962857
R63819 DVSS.n3232 DVSS.n2299 0.00962857
R63820 DVSS.n3233 DVSS.n3232 0.00962857
R63821 DVSS.n3234 DVSS.n3233 0.00962857
R63822 DVSS.n3234 DVSS.n2295 0.00962857
R63823 DVSS.n3240 DVSS.n2295 0.00962857
R63824 DVSS.n3241 DVSS.n3240 0.00962857
R63825 DVSS.n3242 DVSS.n3241 0.00962857
R63826 DVSS.n3242 DVSS.n2291 0.00962857
R63827 DVSS.n3248 DVSS.n2291 0.00962857
R63828 DVSS.n3249 DVSS.n3248 0.00962857
R63829 DVSS.n3250 DVSS.n3249 0.00962857
R63830 DVSS.n3250 DVSS.n2287 0.00962857
R63831 DVSS.n3256 DVSS.n2287 0.00962857
R63832 DVSS.n3257 DVSS.n3256 0.00962857
R63833 DVSS.n3258 DVSS.n3257 0.00962857
R63834 DVSS.n3258 DVSS.n2283 0.00962857
R63835 DVSS.n3264 DVSS.n2283 0.00962857
R63836 DVSS.n3265 DVSS.n3264 0.00962857
R63837 DVSS.n3266 DVSS.n3265 0.00962857
R63838 DVSS.n3266 DVSS.n2277 0.00962857
R63839 DVSS.n3326 DVSS.n2278 0.00962857
R63840 DVSS.n3320 DVSS.n2278 0.00962857
R63841 DVSS.n3320 DVSS.n3319 0.00962857
R63842 DVSS.n3319 DVSS.n3318 0.00962857
R63843 DVSS.n3318 DVSS.n3272 0.00962857
R63844 DVSS.n3312 DVSS.n3272 0.00962857
R63845 DVSS.n3312 DVSS.n3311 0.00962857
R63846 DVSS.n3311 DVSS.n3310 0.00962857
R63847 DVSS.n3310 DVSS.n3276 0.00962857
R63848 DVSS.n3304 DVSS.n3276 0.00962857
R63849 DVSS.n3303 DVSS.n3279 0.00962857
R63850 DVSS.n3295 DVSS.n3279 0.00962857
R63851 DVSS.n3296 DVSS.n3295 0.00962857
R63852 DVSS.n3296 DVSS.n3294 0.00962857
R63853 DVSS.n3502 DVSS.n2143 0.00962857
R63854 DVSS.n3498 DVSS.n2143 0.00962857
R63855 DVSS.n3498 DVSS.n3497 0.00962857
R63856 DVSS.n3497 DVSS.n3496 0.00962857
R63857 DVSS.n3496 DVSS.n2147 0.00962857
R63858 DVSS.n3490 DVSS.n2147 0.00962857
R63859 DVSS.n3490 DVSS.n3489 0.00962857
R63860 DVSS.n3489 DVSS.n3488 0.00962857
R63861 DVSS.n3488 DVSS.n2151 0.00962857
R63862 DVSS.n3482 DVSS.n2151 0.00962857
R63863 DVSS.n3482 DVSS.n3481 0.00962857
R63864 DVSS.n3481 DVSS.n3480 0.00962857
R63865 DVSS.n3480 DVSS.n2155 0.00962857
R63866 DVSS.n3474 DVSS.n2155 0.00962857
R63867 DVSS.n3474 DVSS.n3473 0.00962857
R63868 DVSS.n3473 DVSS.n3472 0.00962857
R63869 DVSS.n3472 DVSS.n2159 0.00962857
R63870 DVSS.n3466 DVSS.n2159 0.00962857
R63871 DVSS.n3466 DVSS.n3465 0.00962857
R63872 DVSS.n3465 DVSS.n3464 0.00962857
R63873 DVSS.n3464 DVSS.n2163 0.00962857
R63874 DVSS.n3458 DVSS.n2163 0.00962857
R63875 DVSS.n3458 DVSS.n3457 0.00962857
R63876 DVSS.n3457 DVSS.n3456 0.00962857
R63877 DVSS.n3456 DVSS.n2167 0.00962857
R63878 DVSS.n3450 DVSS.n2167 0.00962857
R63879 DVSS.n3450 DVSS.n3449 0.00962857
R63880 DVSS.n3449 DVSS.n3448 0.00962857
R63881 DVSS.n3448 DVSS.n2171 0.00962857
R63882 DVSS.n3442 DVSS.n2171 0.00962857
R63883 DVSS.n3442 DVSS.n3441 0.00962857
R63884 DVSS.n3441 DVSS.n3440 0.00962857
R63885 DVSS.n3440 DVSS.n2175 0.00962857
R63886 DVSS.n3434 DVSS.n2175 0.00962857
R63887 DVSS.n3434 DVSS.n3433 0.00962857
R63888 DVSS.n3433 DVSS.n3432 0.00962857
R63889 DVSS.n3432 DVSS.n2179 0.00962857
R63890 DVSS.n3426 DVSS.n2179 0.00962857
R63891 DVSS.n3426 DVSS.n3425 0.00962857
R63892 DVSS.n3425 DVSS.n3424 0.00962857
R63893 DVSS.n3424 DVSS.n2183 0.00962857
R63894 DVSS.n3418 DVSS.n2183 0.00962857
R63895 DVSS.n3418 DVSS.n3417 0.00962857
R63896 DVSS.n3417 DVSS.n3416 0.00962857
R63897 DVSS.n3416 DVSS.n2187 0.00962857
R63898 DVSS.n3410 DVSS.n2187 0.00962857
R63899 DVSS.n3410 DVSS.n3409 0.00962857
R63900 DVSS.n3409 DVSS.n3408 0.00962857
R63901 DVSS.n3408 DVSS.n2191 0.00962857
R63902 DVSS.n3402 DVSS.n2191 0.00962857
R63903 DVSS.n3402 DVSS.n3401 0.00962857
R63904 DVSS.n3401 DVSS.n3400 0.00962857
R63905 DVSS.n3400 DVSS.n2195 0.00962857
R63906 DVSS.n3394 DVSS.n2195 0.00962857
R63907 DVSS.n3394 DVSS.n3393 0.00962857
R63908 DVSS.n3393 DVSS.n3392 0.00962857
R63909 DVSS.n3392 DVSS.n2199 0.00962857
R63910 DVSS.n3386 DVSS.n2199 0.00962857
R63911 DVSS.n3386 DVSS.n3385 0.00962857
R63912 DVSS.n3385 DVSS.n3384 0.00962857
R63913 DVSS.n3384 DVSS.n2203 0.00962857
R63914 DVSS.n3378 DVSS.n2203 0.00962857
R63915 DVSS.n3378 DVSS.n3377 0.00962857
R63916 DVSS.n3377 DVSS.n3376 0.00962857
R63917 DVSS.n3376 DVSS.n2207 0.00962857
R63918 DVSS.n3370 DVSS.n2207 0.00962857
R63919 DVSS.n3370 DVSS.n3369 0.00962857
R63920 DVSS.n3369 DVSS.n3368 0.00962857
R63921 DVSS.n3368 DVSS.n2211 0.00962857
R63922 DVSS.n3362 DVSS.n2211 0.00962857
R63923 DVSS.n3362 DVSS.n3361 0.00962857
R63924 DVSS.n3361 DVSS.n3360 0.00962857
R63925 DVSS.n3360 DVSS.n2215 0.00962857
R63926 DVSS.n3354 DVSS.n2215 0.00962857
R63927 DVSS.n3354 DVSS.n3353 0.00962857
R63928 DVSS.n3353 DVSS.n3352 0.00962857
R63929 DVSS.n3352 DVSS.n2219 0.00962857
R63930 DVSS.n3346 DVSS.n2219 0.00962857
R63931 DVSS.n3346 DVSS.n3345 0.00962857
R63932 DVSS.n3345 DVSS.n3344 0.00962857
R63933 DVSS.n3344 DVSS.n2223 0.00962857
R63934 DVSS.n3338 DVSS.n2223 0.00962857
R63935 DVSS.n3338 DVSS.n3337 0.00962857
R63936 DVSS.n3337 DVSS.n3336 0.00962857
R63937 DVSS.n3336 DVSS.n2227 0.00962857
R63938 DVSS.n3330 DVSS.n2227 0.00962857
R63939 DVSS.n3330 DVSS.n3329 0.00962857
R63940 DVSS.n2276 DVSS.n2231 0.00962857
R63941 DVSS.n2270 DVSS.n2231 0.00962857
R63942 DVSS.n2270 DVSS.n2269 0.00962857
R63943 DVSS.n2269 DVSS.n2268 0.00962857
R63944 DVSS.n2268 DVSS.n2235 0.00962857
R63945 DVSS.n2262 DVSS.n2235 0.00962857
R63946 DVSS.n2262 DVSS.n2261 0.00962857
R63947 DVSS.n2261 DVSS.n2260 0.00962857
R63948 DVSS.n2260 DVSS.n2239 0.00962857
R63949 DVSS.n2254 DVSS.n2239 0.00962857
R63950 DVSS.n2253 DVSS.n2242 0.00962857
R63951 DVSS.n2245 DVSS.n2242 0.00962857
R63952 DVSS.n2246 DVSS.n2245 0.00962857
R63953 DVSS.n2246 DVSS.n2244 0.00962857
R63954 DVSS DVSS.n6534 0.00931551
R63955 DVSS.n149 DVSS.n139 0.00923134
R63956 DVSS.n2798 DVSS.n2401 0.00917857
R63957 DVSS.n5008 DVSS.n5007 0.00917857
R63958 DVSS.n3757 DVSS.n3756 0.00917857
R63959 DVSS.n4706 DVSS.n4703 0.00917857
R63960 DVSS.n6049 DVSS.n6044 0.00917857
R63961 DVSS.n5668 DVSS.n5667 0.00910927
R63962 DVSS.n5667 DVSS.n1274 0.00910927
R63963 DVSS.n5665 DVSS.n1279 0.00910927
R63964 DVSS.n5665 DVSS.n5664 0.00910927
R63965 DVSS.n3327 DVSS.n2277 0.00905
R63966 DVSS.n3329 DVSS.n3328 0.00905
R63967 DVSS.n3026 DVSS.n2429 0.00892143
R63968 DVSS.n3564 DVSS.n1799 0.00892143
R63969 DVSS.n3713 DVSS.n1802 0.00892143
R63970 DVSS.n4652 DVSS.n2011 0.00892143
R63971 DVSS.n6102 DVSS.n1147 0.00892143
R63972 DVSS.n5230 DVSS 0.0088427
R63973 DVSS.n2981 DVSS.n2547 0.00873944
R63974 DVSS.n2954 DVSS.n2400 0.00873944
R63975 DVSS.n1078 DVSS.n460 0.0086
R63976 DVSS.n6263 DVSS.n6262 0.0086
R63977 DVSS.n6209 DVSS.n459 0.0086
R63978 DVSS.n6272 DVSS.n363 0.0086
R63979 DVSS.n6202 DVSS.n444 0.0086
R63980 DVSS.n6265 DVSS.n101 0.0086
R63981 DVSS.n6203 DVSS.n398 0.0086
R63982 DVSS.n6266 DVSS.n59 0.0086
R63983 DVSS.n2908 DVSS 0.00852817
R63984 DVSS.n2907 DVSS 0.00852817
R63985 DVSS.n4430 DVSS.n4429 0.00846348
R63986 DVSS.n1642 DVSS.n1379 0.00846348
R63987 DVSS.n3017 DVSS.n2435 0.00845775
R63988 DVSS.n2984 DVSS.n2525 0.00845775
R63989 DVSS.n1049 DVSS.n1048 0.0084338
R63990 DVSS.n939 DVSS.n938 0.0084338
R63991 DVSS.n4189 DVSS.n4185 0.00819509
R63992 DVSS.n5358 DVSS.n1385 0.00819509
R63993 DVSS.n4185 DVSS.n4182 0.00819509
R63994 DVSS.n5499 DVSS.n1385 0.00819509
R63995 DVSS.n5445 DVSS.n5376 0.00817918
R63996 DVSS.n4246 DVSS.n4068 0.00810135
R63997 DVSS DVSS.n4394 0.00808427
R63998 DVSS.n2761 DVSS.n2647 0.00802143
R63999 DVSS.n3044 DVSS.n2402 0.00802143
R64000 DVSS.n1743 DVSS.n1740 0.00802143
R64001 DVSS.n1720 DVSS.n1713 0.00802143
R64002 DVSS.n3811 DVSS.n3810 0.00802143
R64003 DVSS.n5164 DVSS.n1651 0.00802143
R64004 DVSS.n4742 DVSS.n1974 0.00802143
R64005 DVSS.n5585 DVSS.n1335 0.00802143
R64006 DVSS.n6060 DVSS.n5777 0.00802143
R64007 DVSS.n6052 DVSS.n5802 0.00802143
R64008 DVSS.n1967 DVSS 0.00795787
R64009 DVSS.n6059 DVSS.n6058 0.00788806
R64010 DVSS.n2849 DVSS 0.00782857
R64011 DVSS.n2850 DVSS 0.00782857
R64012 DVSS.n5059 DVSS 0.00782857
R64013 DVSS.n5060 DVSS 0.00782857
R64014 DVSS.n5105 DVSS 0.00782857
R64015 DVSS.n5106 DVSS 0.00782857
R64016 DVSS.n5526 DVSS 0.00782857
R64017 DVSS.n5527 DVSS 0.00782857
R64018 DVSS.n5985 DVSS 0.00782857
R64019 DVSS.n5986 DVSS 0.00782857
R64020 DVSS.n2255 VSS 0.00782857
R64021 DVSS.n3305 VSS 0.00782857
R64022 DVSS.n3304 VSS 0.00782857
R64023 DVSS.n2254 VSS 0.00782857
R64024 DVSS.n3023 DVSS.n2425 0.00776429
R64025 DVSS.n2766 DVSS.n2745 0.00776429
R64026 DVSS.n3657 DVSS.n1798 0.00776429
R64027 DVSS.n3577 DVSS.n1752 0.00776429
R64028 DVSS.n3848 DVSS.n1801 0.00776429
R64029 DVSS.n3806 DVSS.n3726 0.00776429
R64030 DVSS.n4645 DVSS.n2016 0.00776429
R64031 DVSS.n4739 DVSS.n1994 0.00776429
R64032 DVSS.n6099 DVSS.n1143 0.00776429
R64033 DVSS.n5824 DVSS.n5775 0.00776429
R64034 DVSS.n5323 DVSS.n5322 0.00772462
R64035 DVSS.n4998 DVSS.n4997 0.00772015
R64036 DVSS.n5001 DVSS.n1733 0.00772015
R64037 DVSS.n2764 DVSS.n2116 0.00755224
R64038 DVSS.n4395 DVSS 0.00732584
R64039 DVSS.n1966 DVSS.n1874 0.00732584
R64040 DVSS.n2476 DVSS.n2455 0.00716667
R64041 DVSS.n2477 DVSS.n2476 0.00716667
R64042 DVSS.n2478 DVSS.n2477 0.00716667
R64043 DVSS.n2478 DVSS.n2451 0.00716667
R64044 DVSS.n2484 DVSS.n2451 0.00716667
R64045 DVSS.n2485 DVSS.n2484 0.00716667
R64046 DVSS.n2486 DVSS.n2485 0.00716667
R64047 DVSS.n2486 DVSS.n2447 0.00716667
R64048 DVSS.n2492 DVSS.n2447 0.00716667
R64049 DVSS.n2493 DVSS.n2492 0.00716667
R64050 DVSS.n2494 DVSS.n2493 0.00716667
R64051 DVSS.n2494 DVSS.n2443 0.00716667
R64052 DVSS.n2500 DVSS.n2443 0.00716667
R64053 DVSS.n2501 DVSS.n2500 0.00716667
R64054 DVSS.n2502 DVSS.n2501 0.00716667
R64055 DVSS.n2503 DVSS.n2502 0.00716667
R64056 DVSS.n2504 DVSS.n2503 0.00716667
R64057 DVSS.n2505 DVSS.n2504 0.00716667
R64058 DVSS.n2508 DVSS.n2505 0.00716667
R64059 DVSS.n2509 DVSS.n2508 0.00716667
R64060 DVSS.n2510 DVSS.n2509 0.00716667
R64061 DVSS.n2511 DVSS.n2510 0.00716667
R64062 DVSS.n2514 DVSS.n2511 0.00716667
R64063 DVSS.n2515 DVSS.n2514 0.00716667
R64064 DVSS.n2516 DVSS.n2515 0.00716667
R64065 DVSS.n2517 DVSS.n2516 0.00716667
R64066 DVSS.n2520 DVSS.n2517 0.00716667
R64067 DVSS.n2521 DVSS.n2520 0.00716667
R64068 DVSS.n2522 DVSS.n2521 0.00716667
R64069 DVSS.n2523 DVSS.n2522 0.00716667
R64070 DVSS.n2526 DVSS.n2523 0.00716667
R64071 DVSS.n2527 DVSS.n2526 0.00716667
R64072 DVSS.n2528 DVSS.n2527 0.00716667
R64073 DVSS.n2549 DVSS.n2528 0.00716667
R64074 DVSS.n2550 DVSS.n2549 0.00716667
R64075 DVSS.n2551 DVSS.n2550 0.00716667
R64076 DVSS.n2552 DVSS.n2551 0.00716667
R64077 DVSS.n2555 DVSS.n2552 0.00716667
R64078 DVSS.n2556 DVSS.n2555 0.00716667
R64079 DVSS.n2557 DVSS.n2556 0.00716667
R64080 DVSS.n2558 DVSS.n2557 0.00716667
R64081 DVSS.n2561 DVSS.n2558 0.00716667
R64082 DVSS.n2562 DVSS.n2561 0.00716667
R64083 DVSS.n2563 DVSS.n2562 0.00716667
R64084 DVSS.n2564 DVSS.n2563 0.00716667
R64085 DVSS.n2567 DVSS.n2564 0.00716667
R64086 DVSS.n2568 DVSS.n2567 0.00716667
R64087 DVSS.n2569 DVSS.n2568 0.00716667
R64088 DVSS.n2570 DVSS.n2569 0.00716667
R64089 DVSS.n2571 DVSS.n2570 0.00716667
R64090 DVSS.n2572 DVSS.n2571 0.00716667
R64091 DVSS.n2573 DVSS.n2572 0.00716667
R64092 DVSS.n2576 DVSS.n2573 0.00716667
R64093 DVSS.n2577 DVSS.n2576 0.00716667
R64094 DVSS.n2578 DVSS.n2577 0.00716667
R64095 DVSS.n2579 DVSS.n2578 0.00716667
R64096 DVSS.n2582 DVSS.n2579 0.00716667
R64097 DVSS.n2583 DVSS.n2582 0.00716667
R64098 DVSS.n2584 DVSS.n2583 0.00716667
R64099 DVSS.n2585 DVSS.n2584 0.00716667
R64100 DVSS.n2588 DVSS.n2585 0.00716667
R64101 DVSS.n2589 DVSS.n2588 0.00716667
R64102 DVSS.n2590 DVSS.n2589 0.00716667
R64103 DVSS.n2591 DVSS.n2590 0.00716667
R64104 DVSS.n2594 DVSS.n2591 0.00716667
R64105 DVSS.n2595 DVSS.n2594 0.00716667
R64106 DVSS.n2596 DVSS.n2595 0.00716667
R64107 DVSS.n2597 DVSS.n2596 0.00716667
R64108 DVSS.n2888 DVSS.n2597 0.00716667
R64109 DVSS.n2889 DVSS.n2888 0.00716667
R64110 DVSS.n2890 DVSS.n2889 0.00716667
R64111 DVSS.n2891 DVSS.n2890 0.00716667
R64112 DVSS.n2894 DVSS.n2891 0.00716667
R64113 DVSS.n2895 DVSS.n2894 0.00716667
R64114 DVSS.n2896 DVSS.n2895 0.00716667
R64115 DVSS.n2897 DVSS.n2896 0.00716667
R64116 DVSS.n2900 DVSS.n2897 0.00716667
R64117 DVSS.n2901 DVSS.n2900 0.00716667
R64118 DVSS.n2902 DVSS.n2901 0.00716667
R64119 DVSS.n2903 DVSS.n2902 0.00716667
R64120 DVSS.n2904 DVSS.n2903 0.00716667
R64121 DVSS.n4430 DVSS.n3886 0.00694663
R64122 DVSS.n5501 DVSS.n1379 0.00694663
R64123 DVSS.n2599 DVSS.n2593 0.00690845
R64124 DVSS.n3089 DVSS.n3088 0.00684146
R64125 DVSS.n6498 DVSS.n6497 0.0068
R64126 DVSS.n269 DVSS.n255 0.0068
R64127 DVSS.n355 DVSS.n45 0.0068
R64128 DVSS.n260 DVSS.n190 0.0068
R64129 DVSS.n6477 DVSS.n47 0.0068
R64130 DVSS.n262 DVSS.n131 0.0068
R64131 DVSS.n6491 DVSS.n6490 0.0068
R64132 DVSS.n263 DVSS.n236 0.0068
R64133 DVSS.n2473 DVSS.n2472 0.00662676
R64134 DVSS.n2684 DVSS.n2679 0.00658571
R64135 DVSS.n2685 DVSS.n2684 0.00658571
R64136 DVSS.n2686 DVSS.n2685 0.00658571
R64137 DVSS.n2686 DVSS.n2675 0.00658571
R64138 DVSS.n2692 DVSS.n2675 0.00658571
R64139 DVSS.n2693 DVSS.n2692 0.00658571
R64140 DVSS.n2694 DVSS.n2693 0.00658571
R64141 DVSS.n2694 DVSS.n2671 0.00658571
R64142 DVSS.n2700 DVSS.n2671 0.00658571
R64143 DVSS.n2701 DVSS.n2700 0.00658571
R64144 DVSS.n2702 DVSS.n2701 0.00658571
R64145 DVSS.n2702 DVSS.n2667 0.00658571
R64146 DVSS.n2709 DVSS.n2667 0.00658571
R64147 DVSS.n2710 DVSS.n2709 0.00658571
R64148 DVSS.n2711 DVSS.n2710 0.00658571
R64149 DVSS.n2711 DVSS.n2665 0.00658571
R64150 DVSS.n2715 DVSS.n2665 0.00658571
R64151 DVSS.n2716 DVSS.n2715 0.00658571
R64152 DVSS.n2717 DVSS.n2716 0.00658571
R64153 DVSS.n2717 DVSS.n2661 0.00658571
R64154 DVSS.n2723 DVSS.n2661 0.00658571
R64155 DVSS.n2724 DVSS.n2723 0.00658571
R64156 DVSS.n2725 DVSS.n2724 0.00658571
R64157 DVSS.n2725 DVSS.n2657 0.00658571
R64158 DVSS.n2731 DVSS.n2657 0.00658571
R64159 DVSS.n2732 DVSS.n2731 0.00658571
R64160 DVSS.n2733 DVSS.n2732 0.00658571
R64161 DVSS.n2733 DVSS.n2653 0.00658571
R64162 DVSS.n2739 DVSS.n2653 0.00658571
R64163 DVSS.n2740 DVSS.n2739 0.00658571
R64164 DVSS.n2741 DVSS.n2740 0.00658571
R64165 DVSS.n2741 DVSS.n2649 0.00658571
R64166 DVSS.n2768 DVSS.n2649 0.00658571
R64167 DVSS.n2769 DVSS.n2768 0.00658571
R64168 DVSS.n2770 DVSS.n2769 0.00658571
R64169 DVSS.n2770 DVSS.n2645 0.00658571
R64170 DVSS.n2776 DVSS.n2645 0.00658571
R64171 DVSS.n2777 DVSS.n2776 0.00658571
R64172 DVSS.n2778 DVSS.n2777 0.00658571
R64173 DVSS.n2778 DVSS.n2641 0.00658571
R64174 DVSS.n2784 DVSS.n2641 0.00658571
R64175 DVSS.n2785 DVSS.n2784 0.00658571
R64176 DVSS.n2786 DVSS.n2785 0.00658571
R64177 DVSS.n2786 DVSS.n2637 0.00658571
R64178 DVSS.n2792 DVSS.n2637 0.00658571
R64179 DVSS.n2793 DVSS.n2792 0.00658571
R64180 DVSS.n2794 DVSS.n2793 0.00658571
R64181 DVSS.n2794 DVSS.n2633 0.00658571
R64182 DVSS.n2801 DVSS.n2633 0.00658571
R64183 DVSS.n2802 DVSS.n2801 0.00658571
R64184 DVSS.n2803 DVSS.n2802 0.00658571
R64185 DVSS.n2803 DVSS.n2631 0.00658571
R64186 DVSS.n2808 DVSS.n2631 0.00658571
R64187 DVSS.n2809 DVSS.n2808 0.00658571
R64188 DVSS.n2810 DVSS.n2809 0.00658571
R64189 DVSS.n2810 DVSS.n2627 0.00658571
R64190 DVSS.n2816 DVSS.n2627 0.00658571
R64191 DVSS.n2817 DVSS.n2816 0.00658571
R64192 DVSS.n2818 DVSS.n2817 0.00658571
R64193 DVSS.n2818 DVSS.n2623 0.00658571
R64194 DVSS.n2824 DVSS.n2623 0.00658571
R64195 DVSS.n2825 DVSS.n2824 0.00658571
R64196 DVSS.n2826 DVSS.n2825 0.00658571
R64197 DVSS.n2826 DVSS.n2619 0.00658571
R64198 DVSS.n2832 DVSS.n2619 0.00658571
R64199 DVSS.n2833 DVSS.n2832 0.00658571
R64200 DVSS.n2873 DVSS.n2833 0.00658571
R64201 DVSS.n2873 DVSS.n2872 0.00658571
R64202 DVSS.n2872 DVSS.n2871 0.00658571
R64203 DVSS.n2871 DVSS.n2834 0.00658571
R64204 DVSS.n2838 DVSS.n2834 0.00658571
R64205 DVSS.n2864 DVSS.n2838 0.00658571
R64206 DVSS.n2864 DVSS.n2863 0.00658571
R64207 DVSS.n2863 DVSS.n2862 0.00658571
R64208 DVSS.n2862 DVSS.n2839 0.00658571
R64209 DVSS.n2856 DVSS.n2839 0.00658571
R64210 DVSS.n2856 DVSS.n2855 0.00658571
R64211 DVSS.n2855 DVSS.n2854 0.00658571
R64212 DVSS.n2854 DVSS.n2843 0.00658571
R64213 DVSS.n2848 DVSS.n2843 0.00658571
R64214 DVSS.n2848 DVSS.n2847 0.00658571
R64215 DVSS.n3689 DVSS.n3688 0.00658571
R64216 DVSS.n3688 DVSS.n3687 0.00658571
R64217 DVSS.n3687 DVSS.n3548 0.00658571
R64218 DVSS.n3681 DVSS.n3548 0.00658571
R64219 DVSS.n3681 DVSS.n3680 0.00658571
R64220 DVSS.n3680 DVSS.n3679 0.00658571
R64221 DVSS.n3679 DVSS.n3552 0.00658571
R64222 DVSS.n3673 DVSS.n3552 0.00658571
R64223 DVSS.n3673 DVSS.n3672 0.00658571
R64224 DVSS.n3672 DVSS.n3671 0.00658571
R64225 DVSS.n3671 DVSS.n3556 0.00658571
R64226 DVSS.n3665 DVSS.n3556 0.00658571
R64227 DVSS.n3665 DVSS.n3664 0.00658571
R64228 DVSS.n3664 DVSS.n3663 0.00658571
R64229 DVSS.n3663 DVSS.n3560 0.00658571
R64230 DVSS.n3656 DVSS.n3560 0.00658571
R64231 DVSS.n3656 DVSS.n3655 0.00658571
R64232 DVSS.n3655 DVSS.n3654 0.00658571
R64233 DVSS.n3654 DVSS.n3562 0.00658571
R64234 DVSS.n3648 DVSS.n3562 0.00658571
R64235 DVSS.n3648 DVSS.n3647 0.00658571
R64236 DVSS.n3647 DVSS.n3646 0.00658571
R64237 DVSS.n3646 DVSS.n3567 0.00658571
R64238 DVSS.n3640 DVSS.n3567 0.00658571
R64239 DVSS.n3640 DVSS.n3639 0.00658571
R64240 DVSS.n3639 DVSS.n3638 0.00658571
R64241 DVSS.n3638 DVSS.n3571 0.00658571
R64242 DVSS.n3632 DVSS.n3571 0.00658571
R64243 DVSS.n3632 DVSS.n3631 0.00658571
R64244 DVSS.n3631 DVSS.n3630 0.00658571
R64245 DVSS.n3630 DVSS.n3575 0.00658571
R64246 DVSS.n3624 DVSS.n3575 0.00658571
R64247 DVSS.n3624 DVSS.n3623 0.00658571
R64248 DVSS.n3623 DVSS.n3622 0.00658571
R64249 DVSS.n3622 DVSS.n3579 0.00658571
R64250 DVSS.n3583 DVSS.n3579 0.00658571
R64251 DVSS.n3615 DVSS.n3583 0.00658571
R64252 DVSS.n3615 DVSS.n3614 0.00658571
R64253 DVSS.n3614 DVSS.n3613 0.00658571
R64254 DVSS.n3613 DVSS.n3584 0.00658571
R64255 DVSS.n3607 DVSS.n3584 0.00658571
R64256 DVSS.n3607 DVSS.n3606 0.00658571
R64257 DVSS.n3606 DVSS.n3605 0.00658571
R64258 DVSS.n3605 DVSS.n3588 0.00658571
R64259 DVSS.n3599 DVSS.n3588 0.00658571
R64260 DVSS.n3599 DVSS.n3598 0.00658571
R64261 DVSS.n3598 DVSS.n3597 0.00658571
R64262 DVSS.n3597 DVSS.n3592 0.00658571
R64263 DVSS.n3592 DVSS.n1715 0.00658571
R64264 DVSS.n5010 DVSS.n1715 0.00658571
R64265 DVSS.n5011 DVSS.n5010 0.00658571
R64266 DVSS.n5012 DVSS.n5011 0.00658571
R64267 DVSS.n5012 DVSS.n1711 0.00658571
R64268 DVSS.n5018 DVSS.n1711 0.00658571
R64269 DVSS.n5019 DVSS.n5018 0.00658571
R64270 DVSS.n5020 DVSS.n5019 0.00658571
R64271 DVSS.n5020 DVSS.n1707 0.00658571
R64272 DVSS.n5026 DVSS.n1707 0.00658571
R64273 DVSS.n5027 DVSS.n5026 0.00658571
R64274 DVSS.n5028 DVSS.n5027 0.00658571
R64275 DVSS.n5028 DVSS.n1703 0.00658571
R64276 DVSS.n5034 DVSS.n1703 0.00658571
R64277 DVSS.n5035 DVSS.n5034 0.00658571
R64278 DVSS.n5036 DVSS.n5035 0.00658571
R64279 DVSS.n5036 DVSS.n1699 0.00658571
R64280 DVSS.n5042 DVSS.n1699 0.00658571
R64281 DVSS.n5043 DVSS.n5042 0.00658571
R64282 DVSS.n5082 DVSS.n5043 0.00658571
R64283 DVSS.n5082 DVSS.n5081 0.00658571
R64284 DVSS.n5081 DVSS.n5080 0.00658571
R64285 DVSS.n5080 DVSS.n5044 0.00658571
R64286 DVSS.n5074 DVSS.n5044 0.00658571
R64287 DVSS.n5074 DVSS.n5073 0.00658571
R64288 DVSS.n5073 DVSS.n5072 0.00658571
R64289 DVSS.n5072 DVSS.n5049 0.00658571
R64290 DVSS.n5066 DVSS.n5049 0.00658571
R64291 DVSS.n5066 DVSS.n5065 0.00658571
R64292 DVSS.n5065 DVSS.n5064 0.00658571
R64293 DVSS.n5064 DVSS.n5053 0.00658571
R64294 DVSS.n5058 DVSS.n5053 0.00658571
R64295 DVSS.n5058 DVSS.n5057 0.00658571
R64296 DVSS.n3880 DVSS.n3879 0.00658571
R64297 DVSS.n3879 DVSS.n3878 0.00658571
R64298 DVSS.n3878 DVSS.n3697 0.00658571
R64299 DVSS.n3872 DVSS.n3697 0.00658571
R64300 DVSS.n3872 DVSS.n3871 0.00658571
R64301 DVSS.n3871 DVSS.n3870 0.00658571
R64302 DVSS.n3870 DVSS.n3701 0.00658571
R64303 DVSS.n3864 DVSS.n3701 0.00658571
R64304 DVSS.n3864 DVSS.n3863 0.00658571
R64305 DVSS.n3863 DVSS.n3862 0.00658571
R64306 DVSS.n3862 DVSS.n3705 0.00658571
R64307 DVSS.n3856 DVSS.n3705 0.00658571
R64308 DVSS.n3856 DVSS.n3855 0.00658571
R64309 DVSS.n3855 DVSS.n3854 0.00658571
R64310 DVSS.n3854 DVSS.n3709 0.00658571
R64311 DVSS.n3847 DVSS.n3709 0.00658571
R64312 DVSS.n3847 DVSS.n3846 0.00658571
R64313 DVSS.n3846 DVSS.n3845 0.00658571
R64314 DVSS.n3845 DVSS.n3711 0.00658571
R64315 DVSS.n3839 DVSS.n3711 0.00658571
R64316 DVSS.n3839 DVSS.n3838 0.00658571
R64317 DVSS.n3838 DVSS.n3837 0.00658571
R64318 DVSS.n3837 DVSS.n3716 0.00658571
R64319 DVSS.n3831 DVSS.n3716 0.00658571
R64320 DVSS.n3831 DVSS.n3830 0.00658571
R64321 DVSS.n3830 DVSS.n3829 0.00658571
R64322 DVSS.n3829 DVSS.n3720 0.00658571
R64323 DVSS.n3823 DVSS.n3720 0.00658571
R64324 DVSS.n3823 DVSS.n3822 0.00658571
R64325 DVSS.n3822 DVSS.n3821 0.00658571
R64326 DVSS.n3821 DVSS.n3724 0.00658571
R64327 DVSS.n3815 DVSS.n3724 0.00658571
R64328 DVSS.n3815 DVSS.n3814 0.00658571
R64329 DVSS.n3814 DVSS.n3813 0.00658571
R64330 DVSS.n3813 DVSS.n3728 0.00658571
R64331 DVSS.n3785 DVSS.n3728 0.00658571
R64332 DVSS.n3785 DVSS.n3784 0.00658571
R64333 DVSS.n3784 DVSS.n3783 0.00658571
R64334 DVSS.n3783 DVSS.n3738 0.00658571
R64335 DVSS.n3777 DVSS.n3738 0.00658571
R64336 DVSS.n3777 DVSS.n3776 0.00658571
R64337 DVSS.n3776 DVSS.n3775 0.00658571
R64338 DVSS.n3775 DVSS.n3742 0.00658571
R64339 DVSS.n3769 DVSS.n3742 0.00658571
R64340 DVSS.n3769 DVSS.n3768 0.00658571
R64341 DVSS.n3768 DVSS.n3767 0.00658571
R64342 DVSS.n3767 DVSS.n3746 0.00658571
R64343 DVSS.n3761 DVSS.n3746 0.00658571
R64344 DVSS.n3761 DVSS.n3760 0.00658571
R64345 DVSS.n3760 DVSS.n3759 0.00658571
R64346 DVSS.n3759 DVSS.n1660 0.00658571
R64347 DVSS.n5161 DVSS.n1660 0.00658571
R64348 DVSS.n5161 DVSS.n5160 0.00658571
R64349 DVSS.n5160 DVSS.n5159 0.00658571
R64350 DVSS.n5159 DVSS.n1661 0.00658571
R64351 DVSS.n5153 DVSS.n1661 0.00658571
R64352 DVSS.n5153 DVSS.n5152 0.00658571
R64353 DVSS.n5152 DVSS.n5151 0.00658571
R64354 DVSS.n5151 DVSS.n1665 0.00658571
R64355 DVSS.n5145 DVSS.n1665 0.00658571
R64356 DVSS.n5145 DVSS.n5144 0.00658571
R64357 DVSS.n5144 DVSS.n5143 0.00658571
R64358 DVSS.n5143 DVSS.n1669 0.00658571
R64359 DVSS.n5137 DVSS.n1669 0.00658571
R64360 DVSS.n5137 DVSS.n5136 0.00658571
R64361 DVSS.n5136 DVSS.n5135 0.00658571
R64362 DVSS.n5135 DVSS.n1673 0.00658571
R64363 DVSS.n5128 DVSS.n1673 0.00658571
R64364 DVSS.n5128 DVSS.n5127 0.00658571
R64365 DVSS.n5127 DVSS.n5126 0.00658571
R64366 DVSS.n5126 DVSS.n5090 0.00658571
R64367 DVSS.n5120 DVSS.n5090 0.00658571
R64368 DVSS.n5120 DVSS.n5119 0.00658571
R64369 DVSS.n5119 DVSS.n5118 0.00658571
R64370 DVSS.n5118 DVSS.n5095 0.00658571
R64371 DVSS.n5112 DVSS.n5095 0.00658571
R64372 DVSS.n5112 DVSS.n5111 0.00658571
R64373 DVSS.n5111 DVSS.n5110 0.00658571
R64374 DVSS.n5110 DVSS.n5099 0.00658571
R64375 DVSS.n5104 DVSS.n5099 0.00658571
R64376 DVSS.n5104 DVSS.n5103 0.00658571
R64377 DVSS.n3938 DVSS.n3937 0.00658571
R64378 DVSS.n3937 DVSS.n3936 0.00658571
R64379 DVSS.n3936 DVSS.n3901 0.00658571
R64380 DVSS.n3930 DVSS.n3901 0.00658571
R64381 DVSS.n3930 DVSS.n3929 0.00658571
R64382 DVSS.n3929 DVSS.n3928 0.00658571
R64383 DVSS.n3928 DVSS.n3905 0.00658571
R64384 DVSS.n3922 DVSS.n3905 0.00658571
R64385 DVSS.n3922 DVSS.n3921 0.00658571
R64386 DVSS.n3921 DVSS.n3920 0.00658571
R64387 DVSS.n3920 DVSS.n3909 0.00658571
R64388 DVSS.n3914 DVSS.n3909 0.00658571
R64389 DVSS.n3914 DVSS.n3913 0.00658571
R64390 DVSS.n3913 DVSS.n2013 0.00658571
R64391 DVSS.n4648 DVSS.n2013 0.00658571
R64392 DVSS.n4649 DVSS.n4648 0.00658571
R64393 DVSS.n4650 DVSS.n4649 0.00658571
R64394 DVSS.n4650 DVSS.n2009 0.00658571
R64395 DVSS.n4656 DVSS.n2009 0.00658571
R64396 DVSS.n4657 DVSS.n4656 0.00658571
R64397 DVSS.n4658 DVSS.n4657 0.00658571
R64398 DVSS.n4658 DVSS.n2005 0.00658571
R64399 DVSS.n4664 DVSS.n2005 0.00658571
R64400 DVSS.n4665 DVSS.n4664 0.00658571
R64401 DVSS.n4666 DVSS.n4665 0.00658571
R64402 DVSS.n4666 DVSS.n2001 0.00658571
R64403 DVSS.n4672 DVSS.n2001 0.00658571
R64404 DVSS.n4673 DVSS.n4672 0.00658571
R64405 DVSS.n4674 DVSS.n4673 0.00658571
R64406 DVSS.n4674 DVSS.n1997 0.00658571
R64407 DVSS.n4681 DVSS.n1997 0.00658571
R64408 DVSS.n4682 DVSS.n4681 0.00658571
R64409 DVSS.n4737 DVSS.n4682 0.00658571
R64410 DVSS.n4737 DVSS.n4736 0.00658571
R64411 DVSS.n4736 DVSS.n4735 0.00658571
R64412 DVSS.n4735 DVSS.n4683 0.00658571
R64413 DVSS.n4687 DVSS.n4683 0.00658571
R64414 DVSS.n4728 DVSS.n4687 0.00658571
R64415 DVSS.n4728 DVSS.n4727 0.00658571
R64416 DVSS.n4727 DVSS.n4726 0.00658571
R64417 DVSS.n4726 DVSS.n4688 0.00658571
R64418 DVSS.n4720 DVSS.n4688 0.00658571
R64419 DVSS.n4720 DVSS.n4719 0.00658571
R64420 DVSS.n4719 DVSS.n4718 0.00658571
R64421 DVSS.n4718 DVSS.n4692 0.00658571
R64422 DVSS.n4712 DVSS.n4692 0.00658571
R64423 DVSS.n4712 DVSS.n4711 0.00658571
R64424 DVSS.n4711 DVSS.n4710 0.00658571
R64425 DVSS.n4710 DVSS.n4696 0.00658571
R64426 DVSS.n4704 DVSS.n4696 0.00658571
R64427 DVSS.n4704 DVSS.n1344 0.00658571
R64428 DVSS.n5582 DVSS.n1344 0.00658571
R64429 DVSS.n5582 DVSS.n5581 0.00658571
R64430 DVSS.n5581 DVSS.n5580 0.00658571
R64431 DVSS.n5580 DVSS.n1345 0.00658571
R64432 DVSS.n5574 DVSS.n1345 0.00658571
R64433 DVSS.n5574 DVSS.n5573 0.00658571
R64434 DVSS.n5573 DVSS.n5572 0.00658571
R64435 DVSS.n5572 DVSS.n1349 0.00658571
R64436 DVSS.n5566 DVSS.n1349 0.00658571
R64437 DVSS.n5566 DVSS.n5565 0.00658571
R64438 DVSS.n5565 DVSS.n5564 0.00658571
R64439 DVSS.n5564 DVSS.n1353 0.00658571
R64440 DVSS.n5558 DVSS.n1353 0.00658571
R64441 DVSS.n5558 DVSS.n5557 0.00658571
R64442 DVSS.n5557 DVSS.n5556 0.00658571
R64443 DVSS.n5556 DVSS.n1357 0.00658571
R64444 DVSS.n5549 DVSS.n1357 0.00658571
R64445 DVSS.n5549 DVSS.n5548 0.00658571
R64446 DVSS.n5548 DVSS.n5547 0.00658571
R64447 DVSS.n5547 DVSS.n5511 0.00658571
R64448 DVSS.n5541 DVSS.n5511 0.00658571
R64449 DVSS.n5541 DVSS.n5540 0.00658571
R64450 DVSS.n5540 DVSS.n5539 0.00658571
R64451 DVSS.n5539 DVSS.n5516 0.00658571
R64452 DVSS.n5533 DVSS.n5516 0.00658571
R64453 DVSS.n5533 DVSS.n5532 0.00658571
R64454 DVSS.n5532 DVSS.n5531 0.00658571
R64455 DVSS.n5531 DVSS.n5520 0.00658571
R64456 DVSS.n5525 DVSS.n5520 0.00658571
R64457 DVSS.n5856 DVSS.n5854 0.00658571
R64458 DVSS.n5862 DVSS.n5854 0.00658571
R64459 DVSS.n5863 DVSS.n5862 0.00658571
R64460 DVSS.n5864 DVSS.n5863 0.00658571
R64461 DVSS.n5864 DVSS.n5850 0.00658571
R64462 DVSS.n5870 DVSS.n5850 0.00658571
R64463 DVSS.n5871 DVSS.n5870 0.00658571
R64464 DVSS.n5872 DVSS.n5871 0.00658571
R64465 DVSS.n5872 DVSS.n5846 0.00658571
R64466 DVSS.n5878 DVSS.n5846 0.00658571
R64467 DVSS.n5879 DVSS.n5878 0.00658571
R64468 DVSS.n5881 DVSS.n5879 0.00658571
R64469 DVSS.n5881 DVSS.n5880 0.00658571
R64470 DVSS.n5880 DVSS.n5843 0.00658571
R64471 DVSS.n5843 DVSS.n5841 0.00658571
R64472 DVSS.n5889 DVSS.n5841 0.00658571
R64473 DVSS.n5890 DVSS.n5889 0.00658571
R64474 DVSS.n5891 DVSS.n5890 0.00658571
R64475 DVSS.n5891 DVSS.n5838 0.00658571
R64476 DVSS.n5897 DVSS.n5838 0.00658571
R64477 DVSS.n5898 DVSS.n5897 0.00658571
R64478 DVSS.n5899 DVSS.n5898 0.00658571
R64479 DVSS.n5899 DVSS.n5834 0.00658571
R64480 DVSS.n5905 DVSS.n5834 0.00658571
R64481 DVSS.n5906 DVSS.n5905 0.00658571
R64482 DVSS.n5907 DVSS.n5906 0.00658571
R64483 DVSS.n5907 DVSS.n5830 0.00658571
R64484 DVSS.n5913 DVSS.n5830 0.00658571
R64485 DVSS.n5914 DVSS.n5913 0.00658571
R64486 DVSS.n5915 DVSS.n5914 0.00658571
R64487 DVSS.n5915 DVSS.n5826 0.00658571
R64488 DVSS.n5921 DVSS.n5826 0.00658571
R64489 DVSS.n5922 DVSS.n5921 0.00658571
R64490 DVSS.n5923 DVSS.n5922 0.00658571
R64491 DVSS.n5923 DVSS.n5823 0.00658571
R64492 DVSS.n5928 DVSS.n5823 0.00658571
R64493 DVSS.n5929 DVSS.n5928 0.00658571
R64494 DVSS.n5930 DVSS.n5929 0.00658571
R64495 DVSS.n5930 DVSS.n5819 0.00658571
R64496 DVSS.n5936 DVSS.n5819 0.00658571
R64497 DVSS.n5937 DVSS.n5936 0.00658571
R64498 DVSS.n5938 DVSS.n5937 0.00658571
R64499 DVSS.n5938 DVSS.n5815 0.00658571
R64500 DVSS.n5944 DVSS.n5815 0.00658571
R64501 DVSS.n5945 DVSS.n5944 0.00658571
R64502 DVSS.n5946 DVSS.n5945 0.00658571
R64503 DVSS.n5946 DVSS.n5811 0.00658571
R64504 DVSS.n5952 DVSS.n5811 0.00658571
R64505 DVSS.n5953 DVSS.n5952 0.00658571
R64506 DVSS.n6042 DVSS.n5953 0.00658571
R64507 DVSS.n6042 DVSS.n6041 0.00658571
R64508 DVSS.n6041 DVSS.n6040 0.00658571
R64509 DVSS.n6040 DVSS.n5954 0.00658571
R64510 DVSS.n5958 DVSS.n5954 0.00658571
R64511 DVSS.n6033 DVSS.n5958 0.00658571
R64512 DVSS.n6033 DVSS.n6032 0.00658571
R64513 DVSS.n6032 DVSS.n6031 0.00658571
R64514 DVSS.n6031 DVSS.n5959 0.00658571
R64515 DVSS.n6025 DVSS.n5959 0.00658571
R64516 DVSS.n6025 DVSS.n6024 0.00658571
R64517 DVSS.n6024 DVSS.n6023 0.00658571
R64518 DVSS.n6023 DVSS.n5963 0.00658571
R64519 DVSS.n6017 DVSS.n5963 0.00658571
R64520 DVSS.n6017 DVSS.n6016 0.00658571
R64521 DVSS.n6016 DVSS.n6015 0.00658571
R64522 DVSS.n6015 DVSS.n5967 0.00658571
R64523 DVSS.n6009 DVSS.n5967 0.00658571
R64524 DVSS.n6009 DVSS.n6008 0.00658571
R64525 DVSS.n6008 DVSS.n6007 0.00658571
R64526 DVSS.n6007 DVSS.n5970 0.00658571
R64527 DVSS.n5974 DVSS.n5970 0.00658571
R64528 DVSS.n6000 DVSS.n5974 0.00658571
R64529 DVSS.n6000 DVSS.n5999 0.00658571
R64530 DVSS.n5999 DVSS.n5998 0.00658571
R64531 DVSS.n5998 DVSS.n5975 0.00658571
R64532 DVSS.n5992 DVSS.n5975 0.00658571
R64533 DVSS.n5992 DVSS.n5991 0.00658571
R64534 DVSS.n5991 DVSS.n5990 0.00658571
R64535 DVSS.n5990 DVSS.n5979 0.00658571
R64536 DVSS.n5984 DVSS.n5979 0.00658571
R64537 DVSS.n5984 DVSS.n5983 0.00658571
R64538 DVSS.n3500 DVSS.n2145 0.00658571
R64539 DVSS.n3494 DVSS.n2145 0.00658571
R64540 DVSS.n3494 DVSS.n3493 0.00658571
R64541 DVSS.n3493 DVSS.n3492 0.00658571
R64542 DVSS.n3492 DVSS.n2149 0.00658571
R64543 DVSS.n3486 DVSS.n2149 0.00658571
R64544 DVSS.n3486 DVSS.n3485 0.00658571
R64545 DVSS.n3485 DVSS.n3484 0.00658571
R64546 DVSS.n3484 DVSS.n2153 0.00658571
R64547 DVSS.n3478 DVSS.n2153 0.00658571
R64548 DVSS.n3478 DVSS.n3477 0.00658571
R64549 DVSS.n3477 DVSS.n3476 0.00658571
R64550 DVSS.n3476 DVSS.n2157 0.00658571
R64551 DVSS.n3470 DVSS.n2157 0.00658571
R64552 DVSS.n3470 DVSS.n3469 0.00658571
R64553 DVSS.n3469 DVSS.n3468 0.00658571
R64554 DVSS.n3468 DVSS.n2161 0.00658571
R64555 DVSS.n3462 DVSS.n2161 0.00658571
R64556 DVSS.n3462 DVSS.n3461 0.00658571
R64557 DVSS.n3461 DVSS.n3460 0.00658571
R64558 DVSS.n3460 DVSS.n2165 0.00658571
R64559 DVSS.n3454 DVSS.n2165 0.00658571
R64560 DVSS.n3454 DVSS.n3453 0.00658571
R64561 DVSS.n3453 DVSS.n3452 0.00658571
R64562 DVSS.n3452 DVSS.n2169 0.00658571
R64563 DVSS.n3446 DVSS.n2169 0.00658571
R64564 DVSS.n3446 DVSS.n3445 0.00658571
R64565 DVSS.n3445 DVSS.n3444 0.00658571
R64566 DVSS.n3444 DVSS.n2173 0.00658571
R64567 DVSS.n3438 DVSS.n2173 0.00658571
R64568 DVSS.n3438 DVSS.n3437 0.00658571
R64569 DVSS.n3437 DVSS.n3436 0.00658571
R64570 DVSS.n3436 DVSS.n2177 0.00658571
R64571 DVSS.n3430 DVSS.n2177 0.00658571
R64572 DVSS.n3430 DVSS.n3429 0.00658571
R64573 DVSS.n3429 DVSS.n3428 0.00658571
R64574 DVSS.n3428 DVSS.n2181 0.00658571
R64575 DVSS.n3422 DVSS.n2181 0.00658571
R64576 DVSS.n3422 DVSS.n3421 0.00658571
R64577 DVSS.n3421 DVSS.n3420 0.00658571
R64578 DVSS.n3420 DVSS.n2185 0.00658571
R64579 DVSS.n3414 DVSS.n2185 0.00658571
R64580 DVSS.n3414 DVSS.n3413 0.00658571
R64581 DVSS.n3413 DVSS.n3412 0.00658571
R64582 DVSS.n3412 DVSS.n2189 0.00658571
R64583 DVSS.n3406 DVSS.n2189 0.00658571
R64584 DVSS.n3406 DVSS.n3405 0.00658571
R64585 DVSS.n3405 DVSS.n3404 0.00658571
R64586 DVSS.n3404 DVSS.n2193 0.00658571
R64587 DVSS.n3398 DVSS.n2193 0.00658571
R64588 DVSS.n3398 DVSS.n3397 0.00658571
R64589 DVSS.n3397 DVSS.n3396 0.00658571
R64590 DVSS.n3396 DVSS.n2197 0.00658571
R64591 DVSS.n3390 DVSS.n2197 0.00658571
R64592 DVSS.n3390 DVSS.n3389 0.00658571
R64593 DVSS.n3389 DVSS.n3388 0.00658571
R64594 DVSS.n3388 DVSS.n2201 0.00658571
R64595 DVSS.n3382 DVSS.n2201 0.00658571
R64596 DVSS.n3382 DVSS.n3381 0.00658571
R64597 DVSS.n3381 DVSS.n3380 0.00658571
R64598 DVSS.n3380 DVSS.n2205 0.00658571
R64599 DVSS.n3374 DVSS.n2205 0.00658571
R64600 DVSS.n3374 DVSS.n3373 0.00658571
R64601 DVSS.n3373 DVSS.n3372 0.00658571
R64602 DVSS.n3372 DVSS.n2209 0.00658571
R64603 DVSS.n3366 DVSS.n2209 0.00658571
R64604 DVSS.n3366 DVSS.n3365 0.00658571
R64605 DVSS.n3365 DVSS.n3364 0.00658571
R64606 DVSS.n3364 DVSS.n2213 0.00658571
R64607 DVSS.n3358 DVSS.n2213 0.00658571
R64608 DVSS.n3358 DVSS.n3357 0.00658571
R64609 DVSS.n3357 DVSS.n3356 0.00658571
R64610 DVSS.n3356 DVSS.n2217 0.00658571
R64611 DVSS.n3350 DVSS.n2217 0.00658571
R64612 DVSS.n3350 DVSS.n3349 0.00658571
R64613 DVSS.n3349 DVSS.n3348 0.00658571
R64614 DVSS.n3348 DVSS.n2221 0.00658571
R64615 DVSS.n3342 DVSS.n2221 0.00658571
R64616 DVSS.n3342 DVSS.n3341 0.00658571
R64617 DVSS.n3341 DVSS.n3340 0.00658571
R64618 DVSS.n3340 DVSS.n2225 0.00658571
R64619 DVSS.n3334 DVSS.n2225 0.00658571
R64620 DVSS.n3334 DVSS.n3333 0.00658571
R64621 DVSS.n3333 DVSS.n3332 0.00658571
R64622 DVSS.n3332 DVSS.n2229 0.00658571
R64623 DVSS.n2274 DVSS.n2229 0.00658571
R64624 DVSS.n2274 DVSS.n2273 0.00658571
R64625 DVSS.n2273 DVSS.n2272 0.00658571
R64626 DVSS.n2272 DVSS.n2233 0.00658571
R64627 DVSS.n2266 DVSS.n2233 0.00658571
R64628 DVSS.n2266 DVSS.n2265 0.00658571
R64629 DVSS.n2265 DVSS.n2264 0.00658571
R64630 DVSS.n2264 DVSS.n2237 0.00658571
R64631 DVSS.n2258 DVSS.n2237 0.00658571
R64632 DVSS.n2258 DVSS.n2257 0.00658571
R64633 DVSS.n2257 DVSS.n2256 0.00658571
R64634 DVSS.n2256 DVSS.n2241 0.00658571
R64635 DVSS.n2250 DVSS.n2249 0.00658571
R64636 DVSS.n3101 DVSS.n3100 0.00658571
R64637 DVSS.n3102 DVSS.n3101 0.00658571
R64638 DVSS.n3102 DVSS.n2361 0.00658571
R64639 DVSS.n3108 DVSS.n2361 0.00658571
R64640 DVSS.n3109 DVSS.n3108 0.00658571
R64641 DVSS.n3110 DVSS.n3109 0.00658571
R64642 DVSS.n3110 DVSS.n2357 0.00658571
R64643 DVSS.n3116 DVSS.n2357 0.00658571
R64644 DVSS.n3117 DVSS.n3116 0.00658571
R64645 DVSS.n3118 DVSS.n3117 0.00658571
R64646 DVSS.n3118 DVSS.n2353 0.00658571
R64647 DVSS.n3124 DVSS.n2353 0.00658571
R64648 DVSS.n3125 DVSS.n3124 0.00658571
R64649 DVSS.n3126 DVSS.n3125 0.00658571
R64650 DVSS.n3126 DVSS.n2349 0.00658571
R64651 DVSS.n3132 DVSS.n2349 0.00658571
R64652 DVSS.n3133 DVSS.n3132 0.00658571
R64653 DVSS.n3134 DVSS.n3133 0.00658571
R64654 DVSS.n3134 DVSS.n2345 0.00658571
R64655 DVSS.n3140 DVSS.n2345 0.00658571
R64656 DVSS.n3141 DVSS.n3140 0.00658571
R64657 DVSS.n3142 DVSS.n3141 0.00658571
R64658 DVSS.n3142 DVSS.n2341 0.00658571
R64659 DVSS.n3148 DVSS.n2341 0.00658571
R64660 DVSS.n3149 DVSS.n3148 0.00658571
R64661 DVSS.n3150 DVSS.n3149 0.00658571
R64662 DVSS.n3150 DVSS.n2337 0.00658571
R64663 DVSS.n3156 DVSS.n2337 0.00658571
R64664 DVSS.n3157 DVSS.n3156 0.00658571
R64665 DVSS.n3158 DVSS.n3157 0.00658571
R64666 DVSS.n3158 DVSS.n2333 0.00658571
R64667 DVSS.n3164 DVSS.n2333 0.00658571
R64668 DVSS.n3165 DVSS.n3164 0.00658571
R64669 DVSS.n3166 DVSS.n3165 0.00658571
R64670 DVSS.n3166 DVSS.n2329 0.00658571
R64671 DVSS.n3172 DVSS.n2329 0.00658571
R64672 DVSS.n3173 DVSS.n3172 0.00658571
R64673 DVSS.n3174 DVSS.n3173 0.00658571
R64674 DVSS.n3174 DVSS.n2325 0.00658571
R64675 DVSS.n3180 DVSS.n2325 0.00658571
R64676 DVSS.n3181 DVSS.n3180 0.00658571
R64677 DVSS.n3182 DVSS.n3181 0.00658571
R64678 DVSS.n3182 DVSS.n2321 0.00658571
R64679 DVSS.n3188 DVSS.n2321 0.00658571
R64680 DVSS.n3189 DVSS.n3188 0.00658571
R64681 DVSS.n3190 DVSS.n3189 0.00658571
R64682 DVSS.n3190 DVSS.n2317 0.00658571
R64683 DVSS.n3196 DVSS.n2317 0.00658571
R64684 DVSS.n3197 DVSS.n3196 0.00658571
R64685 DVSS.n3198 DVSS.n3197 0.00658571
R64686 DVSS.n3198 DVSS.n2313 0.00658571
R64687 DVSS.n3204 DVSS.n2313 0.00658571
R64688 DVSS.n3205 DVSS.n3204 0.00658571
R64689 DVSS.n3206 DVSS.n3205 0.00658571
R64690 DVSS.n3206 DVSS.n2309 0.00658571
R64691 DVSS.n3212 DVSS.n2309 0.00658571
R64692 DVSS.n3213 DVSS.n3212 0.00658571
R64693 DVSS.n3214 DVSS.n3213 0.00658571
R64694 DVSS.n3214 DVSS.n2305 0.00658571
R64695 DVSS.n3220 DVSS.n2305 0.00658571
R64696 DVSS.n3221 DVSS.n3220 0.00658571
R64697 DVSS.n3222 DVSS.n3221 0.00658571
R64698 DVSS.n3222 DVSS.n2301 0.00658571
R64699 DVSS.n3228 DVSS.n2301 0.00658571
R64700 DVSS.n3229 DVSS.n3228 0.00658571
R64701 DVSS.n3230 DVSS.n3229 0.00658571
R64702 DVSS.n3230 DVSS.n2297 0.00658571
R64703 DVSS.n3236 DVSS.n2297 0.00658571
R64704 DVSS.n3237 DVSS.n3236 0.00658571
R64705 DVSS.n3238 DVSS.n3237 0.00658571
R64706 DVSS.n3238 DVSS.n2293 0.00658571
R64707 DVSS.n3244 DVSS.n2293 0.00658571
R64708 DVSS.n3245 DVSS.n3244 0.00658571
R64709 DVSS.n3246 DVSS.n3245 0.00658571
R64710 DVSS.n3246 DVSS.n2289 0.00658571
R64711 DVSS.n3252 DVSS.n2289 0.00658571
R64712 DVSS.n3253 DVSS.n3252 0.00658571
R64713 DVSS.n3254 DVSS.n3253 0.00658571
R64714 DVSS.n3254 DVSS.n2285 0.00658571
R64715 DVSS.n3260 DVSS.n2285 0.00658571
R64716 DVSS.n3261 DVSS.n3260 0.00658571
R64717 DVSS.n3262 DVSS.n3261 0.00658571
R64718 DVSS.n3262 DVSS.n2281 0.00658571
R64719 DVSS.n3268 DVSS.n2281 0.00658571
R64720 DVSS.n3269 DVSS.n3268 0.00658571
R64721 DVSS.n3324 DVSS.n3269 0.00658571
R64722 DVSS.n3324 DVSS.n3323 0.00658571
R64723 DVSS.n3323 DVSS.n3322 0.00658571
R64724 DVSS.n3322 DVSS.n3270 0.00658571
R64725 DVSS.n3316 DVSS.n3270 0.00658571
R64726 DVSS.n3316 DVSS.n3315 0.00658571
R64727 DVSS.n3315 DVSS.n3314 0.00658571
R64728 DVSS.n3314 DVSS.n3274 0.00658571
R64729 DVSS.n3308 DVSS.n3274 0.00658571
R64730 DVSS.n3308 DVSS.n3307 0.00658571
R64731 DVSS.n3307 DVSS.n3306 0.00658571
R64732 DVSS.n3306 DVSS.n3278 0.00658571
R64733 DVSS.n3300 DVSS.n3299 0.00658571
R64734 DVSS DVSS.n5229 0.00656742
R64735 DVSS.n6464 DVSS.n144 0.00654478
R64736 DVSS.n657 DVSS.n656 0.0065
R64737 DVSS.n803 DVSS.n562 0.0065
R64738 DVSS.n716 DVSS.n559 0.0065
R64739 DVSS.n997 DVSS.n996 0.0065
R64740 DVSS.n594 DVSS.n593 0.0065
R64741 DVSS.n842 DVSS.n559 0.0065
R64742 DVSS.n996 DVSS.n995 0.0065
R64743 DVSS.n6508 DVSS.n13 0.0065
R64744 DVSS.n6508 DVSS.n14 0.0065
R64745 DVSS.n593 DVSS.n592 0.0065
R64746 DVSS.n1031 DVSS.n12 0.0065
R64747 DVSS.n803 DVSS.n567 0.0065
R64748 DVSS.n658 DVSS.n657 0.0065
R64749 DVSS.n6348 DVSS.n342 0.0065
R64750 DVSS.n6348 DVSS.n343 0.0065
R64751 DVSS.n957 DVSS.n12 0.0065
R64752 DVSS.n2250 VSS 0.00641429
R64753 DVSS.n3300 VSS 0.00641429
R64754 DVSS.n2880 DVSS.n2875 0.00635
R64755 DVSS.n5085 DVSS.n1686 0.00635
R64756 DVSS.n5132 DVSS.n5131 0.00635
R64757 DVSS.n5553 DVSS.n5552 0.00635
R64758 DVSS.n6011 DVSS.n1183 0.00635
R64759 DVSS.n1099 DVSS.n468 0.00620896
R64760 DVSS.n3543 DVSS.n2103 0.00609286
R64761 DVSS.n3692 DVSS.n3691 0.00609286
R64762 DVSS.n3883 DVSS.n3882 0.00609286
R64763 DVSS.n3941 DVSS.n3940 0.00609286
R64764 DVSS.n6093 DVSS.n1162 0.00609286
R64765 DVSS.n1467 DVSS.n1412 0.00572184
R64766 DVSS.n4124 DVSS.n4123 0.00566892
R64767 DVSS.n2928 DVSS.n2927 0.00564085
R64768 DVSS.n6445 DVSS.n158 0.00553731
R64769 DVSS.n2248 DVSS.n2247 0.00548841
R64770 DVSS.n3501 DVSS.n2144 0.00548841
R64771 DVSS.n3298 DVSS.n3297 0.00548841
R64772 DVSS.n2366 DVSS.n2365 0.00548841
R64773 DVSS.n5525 DVSS 0.00538571
R64774 DVSS.n2546 DVSS.n2530 0.00536196
R64775 DVSS.n2983 DVSS.n2530 0.00536196
R64776 DVSS.n2470 DVSS.n2457 0.00535915
R64777 DVSS.n2927 DVSS.n2924 0.00535915
R64778 DVSS.n2883 DVSS.n2609 0.00519286
R64779 DVSS.n5084 DVSS.n1696 0.00519286
R64780 DVSS.n5130 DVSS.n5088 0.00519286
R64781 DVSS.n5551 DVSS.n5509 0.00519286
R64782 DVSS.n6071 DVSS.n1185 0.00519286
R64783 DVSS.n3528 DVSS.n2117 0.00513023
R64784 DVSS.n3530 DVSS.n2117 0.00513023
R64785 DVSS.n4850 DVSS.n1867 0.00503358
R64786 DVSS.n3521 DVSS.n2131 0.005
R64787 DVSS.n1080 DVSS.n458 0.005
R64788 DVSS.n6274 DVSS.n26 0.005
R64789 DVSS.n3526 DVSS.n2127 0.005
R64790 DVSS.n6219 DVSS.n6214 0.005
R64791 DVSS.n6283 DVSS.n384 0.005
R64792 DVSS.n3532 DVSS.n2114 0.005
R64793 DVSS.n6227 DVSS.n6226 0.005
R64794 DVSS.n6276 DVSS.n85 0.005
R64795 DVSS.n3538 DVSS.n2101 0.005
R64796 DVSS.n6224 DVSS.n411 0.005
R64797 DVSS.n6277 DVSS.n70 0.005
R64798 DVSS.n2763 DVSS.n2753 0.00498219
R64799 DVSS.n4996 DVSS.n1741 0.00498219
R64800 DVSS.n3808 DVSS.n3807 0.00498219
R64801 DVSS.n4740 DVSS.n1973 0.00498219
R64802 DVSS.n5798 DVSS.n5794 0.00498219
R64803 DVSS.n5794 DVSS.n5776 0.00498219
R64804 DVSS.n1988 DVSS.n1973 0.00498219
R64805 DVSS.n3808 DVSS.n3730 0.00498219
R64806 DVSS.n1741 DVSS.n1739 0.00498219
R64807 DVSS.n2765 DVSS.n2753 0.00498219
R64808 DVSS.n3540 DVSS.n2098 0.00493571
R64809 DVSS.n2883 DVSS.n2611 0.00493571
R64810 DVSS.n3546 DVSS.n2084 0.00493571
R64811 DVSS.n5046 DVSS.n1696 0.00493571
R64812 DVSS.n3695 DVSS.n2070 0.00493571
R64813 DVSS.n5092 DVSS.n5088 0.00493571
R64814 DVSS.n3896 DVSS.n3895 0.00493571
R64815 DVSS.n5513 DVSS.n5509 0.00493571
R64816 DVSS.n6090 DVSS.n1159 0.00493571
R64817 DVSS.n6071 DVSS.n1192 0.00493571
R64818 DVSS.n2746 DVSS.n2121 0.00486567
R64819 DVSS.n1110 DVSS.n487 0.00486567
R64820 DVSS.n4432 DVSS.n2055 0.00476
R64821 DVSS.n4451 DVSS.n2055 0.00476
R64822 DVSS.n4451 DVSS.n2053 0.00476
R64823 DVSS.n4455 DVSS.n2053 0.00476
R64824 DVSS.n4455 DVSS.n2051 0.00476
R64825 DVSS.n4459 DVSS.n2051 0.00476
R64826 DVSS.n4459 DVSS.n2049 0.00476
R64827 DVSS.n4463 DVSS.n2049 0.00476
R64828 DVSS.n4463 DVSS.n2047 0.00476
R64829 DVSS.n4467 DVSS.n2047 0.00476
R64830 DVSS.n4467 DVSS.n2045 0.00476
R64831 DVSS.n4471 DVSS.n2045 0.00476
R64832 DVSS.n4471 DVSS.n2043 0.00476
R64833 DVSS.n4475 DVSS.n2043 0.00476
R64834 DVSS.n4475 DVSS.n2041 0.00476
R64835 DVSS.n4624 DVSS.n2041 0.00476
R64836 DVSS.n4624 DVSS.n4623 0.00476
R64837 DVSS.n4623 DVSS.n4622 0.00476
R64838 DVSS.n4622 DVSS.n4621 0.00476
R64839 DVSS.n4621 DVSS.n4482 0.00476
R64840 DVSS.n4617 DVSS.n4482 0.00476
R64841 DVSS.n4617 DVSS.n4616 0.00476
R64842 DVSS.n4616 DVSS.n4615 0.00476
R64843 DVSS.n4615 DVSS.n4488 0.00476
R64844 DVSS.n4611 DVSS.n4488 0.00476
R64845 DVSS.n4611 DVSS.n4610 0.00476
R64846 DVSS.n4610 DVSS.n4609 0.00476
R64847 DVSS.n4609 DVSS.n4494 0.00476
R64848 DVSS.n4605 DVSS.n4494 0.00476
R64849 DVSS.n4605 DVSS.n4604 0.00476
R64850 DVSS.n4604 DVSS.n4603 0.00476
R64851 DVSS.n4603 DVSS.n4500 0.00476
R64852 DVSS.n4599 DVSS.n4500 0.00476
R64853 DVSS.n4599 DVSS.n4598 0.00476
R64854 DVSS.n4598 DVSS.n4505 0.00476
R64855 DVSS.n4592 DVSS.n4505 0.00476
R64856 DVSS.n4592 DVSS.n4591 0.00476
R64857 DVSS.n4591 DVSS.n4590 0.00476
R64858 DVSS.n4590 DVSS.n4556 0.00476
R64859 DVSS.n4586 DVSS.n4556 0.00476
R64860 DVSS.n4586 DVSS.n4585 0.00476
R64861 DVSS.n4585 DVSS.n4584 0.00476
R64862 DVSS.n4584 DVSS.n4562 0.00476
R64863 DVSS.n4580 DVSS.n4562 0.00476
R64864 DVSS.n4580 DVSS.n4579 0.00476
R64865 DVSS.n4579 DVSS.n4578 0.00476
R64866 DVSS.n4578 DVSS.n4568 0.00476
R64867 DVSS.n4574 DVSS.n4568 0.00476
R64868 DVSS.n4574 DVSS.n4573 0.00476
R64869 DVSS.n4573 DVSS.n1567 0.00476
R64870 DVSS.n5267 DVSS.n1567 0.00476
R64871 DVSS.n5267 DVSS.n1565 0.00476
R64872 DVSS.n5271 DVSS.n1565 0.00476
R64873 DVSS.n5271 DVSS.n1563 0.00476
R64874 DVSS.n5275 DVSS.n1563 0.00476
R64875 DVSS.n5275 DVSS.n1561 0.00476
R64876 DVSS.n5279 DVSS.n1561 0.00476
R64877 DVSS.n5279 DVSS.n1559 0.00476
R64878 DVSS.n5283 DVSS.n1559 0.00476
R64879 DVSS.n5283 DVSS.n1557 0.00476
R64880 DVSS.n5287 DVSS.n1557 0.00476
R64881 DVSS.n5287 DVSS.n1555 0.00476
R64882 DVSS.n5291 DVSS.n1555 0.00476
R64883 DVSS.n5291 DVSS.n1553 0.00476
R64884 DVSS.n5295 DVSS.n1553 0.00476
R64885 DVSS.n5295 DVSS.n1551 0.00476
R64886 DVSS.n5299 DVSS.n1551 0.00476
R64887 DVSS.n5299 DVSS.n1549 0.00476
R64888 DVSS.n5342 DVSS.n1549 0.00476
R64889 DVSS.n5342 DVSS.n5341 0.00476
R64890 DVSS.n5341 DVSS.n5304 0.00476
R64891 DVSS.n5337 DVSS.n5304 0.00476
R64892 DVSS.n5337 DVSS.n5336 0.00476
R64893 DVSS.n5336 DVSS.n5335 0.00476
R64894 DVSS.n5335 DVSS.n5310 0.00476
R64895 DVSS.n5331 DVSS.n5310 0.00476
R64896 DVSS.n5331 DVSS.n5330 0.00476
R64897 DVSS.n5330 DVSS.n5329 0.00476
R64898 DVSS.n5329 DVSS.n5316 0.00476
R64899 DVSS.n5325 DVSS.n5316 0.00476
R64900 DVSS.n5325 DVSS.n5324 0.00476
R64901 DVSS.n4450 DVSS.n4449 0.00476
R64902 DVSS.n4450 DVSS.n2052 0.00476
R64903 DVSS.n4456 DVSS.n2052 0.00476
R64904 DVSS.n4457 DVSS.n4456 0.00476
R64905 DVSS.n4458 DVSS.n4457 0.00476
R64906 DVSS.n4458 DVSS.n2048 0.00476
R64907 DVSS.n4464 DVSS.n2048 0.00476
R64908 DVSS.n4465 DVSS.n4464 0.00476
R64909 DVSS.n4466 DVSS.n4465 0.00476
R64910 DVSS.n4466 DVSS.n2044 0.00476
R64911 DVSS.n4472 DVSS.n2044 0.00476
R64912 DVSS.n4473 DVSS.n4472 0.00476
R64913 DVSS.n4474 DVSS.n4473 0.00476
R64914 DVSS.n4474 DVSS.n2040 0.00476
R64915 DVSS.n4625 DVSS.n2040 0.00476
R64916 DVSS.n4620 DVSS.n2028 0.00476
R64917 DVSS.n4620 DVSS.n4619 0.00476
R64918 DVSS.n4619 DVSS.n4618 0.00476
R64919 DVSS.n4618 DVSS.n4483 0.00476
R64920 DVSS.n4614 DVSS.n4483 0.00476
R64921 DVSS.n4614 DVSS.n4613 0.00476
R64922 DVSS.n4613 DVSS.n4612 0.00476
R64923 DVSS.n4612 DVSS.n4489 0.00476
R64924 DVSS.n4608 DVSS.n4489 0.00476
R64925 DVSS.n4608 DVSS.n4607 0.00476
R64926 DVSS.n4607 DVSS.n4606 0.00476
R64927 DVSS.n4606 DVSS.n4495 0.00476
R64928 DVSS.n4602 DVSS.n4495 0.00476
R64929 DVSS.n4602 DVSS.n4601 0.00476
R64930 DVSS.n4601 DVSS.n4600 0.00476
R64931 DVSS.n4593 DVSS.n4551 0.00476
R64932 DVSS.n4589 DVSS.n4551 0.00476
R64933 DVSS.n4589 DVSS.n4588 0.00476
R64934 DVSS.n4588 DVSS.n4587 0.00476
R64935 DVSS.n4587 DVSS.n4557 0.00476
R64936 DVSS.n4583 DVSS.n4557 0.00476
R64937 DVSS.n4583 DVSS.n4582 0.00476
R64938 DVSS.n4582 DVSS.n4581 0.00476
R64939 DVSS.n4581 DVSS.n4563 0.00476
R64940 DVSS.n4577 DVSS.n4563 0.00476
R64941 DVSS.n4577 DVSS.n4576 0.00476
R64942 DVSS.n4576 DVSS.n4575 0.00476
R64943 DVSS.n4575 DVSS.n4569 0.00476
R64944 DVSS.n4569 DVSS.n1568 0.00476
R64945 DVSS.n5266 DVSS.n1568 0.00476
R64946 DVSS.n5273 DVSS.n5272 0.00476
R64947 DVSS.n5274 DVSS.n5273 0.00476
R64948 DVSS.n5274 DVSS.n1560 0.00476
R64949 DVSS.n5280 DVSS.n1560 0.00476
R64950 DVSS.n5281 DVSS.n5280 0.00476
R64951 DVSS.n5282 DVSS.n5281 0.00476
R64952 DVSS.n5282 DVSS.n1556 0.00476
R64953 DVSS.n5288 DVSS.n1556 0.00476
R64954 DVSS.n5289 DVSS.n5288 0.00476
R64955 DVSS.n5290 DVSS.n5289 0.00476
R64956 DVSS.n5290 DVSS.n1552 0.00476
R64957 DVSS.n5296 DVSS.n1552 0.00476
R64958 DVSS.n5297 DVSS.n5296 0.00476
R64959 DVSS.n5298 DVSS.n5297 0.00476
R64960 DVSS.n5298 DVSS.n1527 0.00476
R64961 DVSS.n5340 DVSS.n5339 0.00476
R64962 DVSS.n5339 DVSS.n5338 0.00476
R64963 DVSS.n5338 DVSS.n5305 0.00476
R64964 DVSS.n5334 DVSS.n5305 0.00476
R64965 DVSS.n5334 DVSS.n5333 0.00476
R64966 DVSS.n5333 DVSS.n5332 0.00476
R64967 DVSS.n5332 DVSS.n5311 0.00476
R64968 DVSS.n5328 DVSS.n5311 0.00476
R64969 DVSS.n5328 DVSS.n5327 0.00476
R64970 DVSS.n5327 DVSS.n5326 0.00476
R64971 DVSS.n5326 DVSS.n5317 0.00476
R64972 DVSS.n598 DVSS.n241 0.00476
R64973 DVSS.n599 DVSS.n598 0.00476
R64974 DVSS.n602 DVSS.n599 0.00476
R64975 DVSS.n603 DVSS.n602 0.00476
R64976 DVSS.n604 DVSS.n603 0.00476
R64977 DVSS.n605 DVSS.n604 0.00476
R64978 DVSS.n608 DVSS.n605 0.00476
R64979 DVSS.n609 DVSS.n608 0.00476
R64980 DVSS.n610 DVSS.n609 0.00476
R64981 DVSS.n611 DVSS.n610 0.00476
R64982 DVSS.n614 DVSS.n611 0.00476
R64983 DVSS.n615 DVSS.n614 0.00476
R64984 DVSS.n616 DVSS.n615 0.00476
R64985 DVSS.n617 DVSS.n616 0.00476
R64986 DVSS.n617 DVSS.n109 0.00476
R64987 DVSS.n620 DVSS.n134 0.00476
R64988 DVSS.n621 DVSS.n620 0.00476
R64989 DVSS.n621 DVSS.n560 0.00476
R64990 DVSS.n841 DVSS.n560 0.00476
R64991 DVSS.n844 DVSS.n843 0.00476
R64992 DVSS.n844 DVSS.n555 0.00476
R64993 DVSS.n850 DVSS.n555 0.00476
R64994 DVSS.n851 DVSS.n850 0.00476
R64995 DVSS.n852 DVSS.n851 0.00476
R64996 DVSS.n852 DVSS.n551 0.00476
R64997 DVSS.n859 DVSS.n551 0.00476
R64998 DVSS.n860 DVSS.n859 0.00476
R64999 DVSS.n861 DVSS.n860 0.00476
R65000 DVSS.n861 DVSS.n154 0.00476
R65001 DVSS.n870 DVSS.n869 0.00476
R65002 DVSS.n870 DVSS.n544 0.00476
R65003 DVSS.n876 DVSS.n544 0.00476
R65004 DVSS.n877 DVSS.n876 0.00476
R65005 DVSS.n878 DVSS.n877 0.00476
R65006 DVSS.n878 DVSS.n540 0.00476
R65007 DVSS.n885 DVSS.n540 0.00476
R65008 DVSS.n886 DVSS.n885 0.00476
R65009 DVSS.n887 DVSS.n886 0.00476
R65010 DVSS.n887 DVSS.n535 0.00476
R65011 DVSS.n994 DVSS.n536 0.00476
R65012 DVSS.n893 DVSS.n536 0.00476
R65013 DVSS.n894 DVSS.n893 0.00476
R65014 DVSS.n895 DVSS.n894 0.00476
R65015 DVSS.n898 DVSS.n193 0.00476
R65016 DVSS.n899 DVSS.n898 0.00476
R65017 DVSS.n902 DVSS.n899 0.00476
R65018 DVSS.n903 DVSS.n902 0.00476
R65019 DVSS.n904 DVSS.n903 0.00476
R65020 DVSS.n905 DVSS.n904 0.00476
R65021 DVSS.n908 DVSS.n905 0.00476
R65022 DVSS.n909 DVSS.n908 0.00476
R65023 DVSS.n910 DVSS.n909 0.00476
R65024 DVSS.n911 DVSS.n910 0.00476
R65025 DVSS.n914 DVSS.n911 0.00476
R65026 DVSS.n915 DVSS.n914 0.00476
R65027 DVSS.n916 DVSS.n915 0.00476
R65028 DVSS.n917 DVSS.n916 0.00476
R65029 DVSS.n917 DVSS.n273 0.00476
R65030 DVSS.n924 DVSS.n920 0.00476
R65031 DVSS.n925 DVSS.n924 0.00476
R65032 DVSS.n926 DVSS.n925 0.00476
R65033 DVSS.n927 DVSS.n926 0.00476
R65034 DVSS.n930 DVSS.n927 0.00476
R65035 DVSS.n931 DVSS.n930 0.00476
R65036 DVSS.n932 DVSS.n931 0.00476
R65037 DVSS.n933 DVSS.n932 0.00476
R65038 DVSS.n936 DVSS.n933 0.00476
R65039 DVSS.n937 DVSS.n936 0.00476
R65040 DVSS.n761 DVSS.n60 0.00476
R65041 DVSS.n761 DVSS.n583 0.00476
R65042 DVSS.n767 DVSS.n583 0.00476
R65043 DVSS.n768 DVSS.n767 0.00476
R65044 DVSS.n769 DVSS.n768 0.00476
R65045 DVSS.n769 DVSS.n579 0.00476
R65046 DVSS.n775 DVSS.n579 0.00476
R65047 DVSS.n776 DVSS.n775 0.00476
R65048 DVSS.n777 DVSS.n776 0.00476
R65049 DVSS.n777 DVSS.n575 0.00476
R65050 DVSS.n783 DVSS.n575 0.00476
R65051 DVSS.n784 DVSS.n783 0.00476
R65052 DVSS.n786 DVSS.n784 0.00476
R65053 DVSS.n786 DVSS.n785 0.00476
R65054 DVSS.n785 DVSS.n80 0.00476
R65055 DVSS.n569 DVSS.n102 0.00476
R65056 DVSS.n799 DVSS.n569 0.00476
R65057 DVSS.n800 DVSS.n799 0.00476
R65058 DVSS.n801 DVSS.n800 0.00476
R65059 DVSS.n805 DVSS.n804 0.00476
R65060 DVSS.n806 DVSS.n805 0.00476
R65061 DVSS.n809 DVSS.n806 0.00476
R65062 DVSS.n810 DVSS.n809 0.00476
R65063 DVSS.n811 DVSS.n810 0.00476
R65064 DVSS.n812 DVSS.n811 0.00476
R65065 DVSS.n815 DVSS.n812 0.00476
R65066 DVSS.n816 DVSS.n815 0.00476
R65067 DVSS.n817 DVSS.n816 0.00476
R65068 DVSS.n817 DVSS.n285 0.00476
R65069 DVSS.n6366 DVSS.n324 0.00476
R65070 DVSS.n329 DVSS.n324 0.00476
R65071 DVSS.n330 DVSS.n329 0.00476
R65072 DVSS.n331 DVSS.n330 0.00476
R65073 DVSS.n334 DVSS.n331 0.00476
R65074 DVSS.n335 DVSS.n334 0.00476
R65075 DVSS.n336 DVSS.n335 0.00476
R65076 DVSS.n337 DVSS.n336 0.00476
R65077 DVSS.n340 DVSS.n337 0.00476
R65078 DVSS.n341 DVSS.n340 0.00476
R65079 DVSS.n347 DVSS.n344 0.00476
R65080 DVSS.n348 DVSS.n347 0.00476
R65081 DVSS.n349 DVSS.n348 0.00476
R65082 DVSS.n350 DVSS.n349 0.00476
R65083 DVSS.n6299 DVSS.n6298 0.00476
R65084 DVSS.n6300 DVSS.n6299 0.00476
R65085 DVSS.n6303 DVSS.n6300 0.00476
R65086 DVSS.n6304 DVSS.n6303 0.00476
R65087 DVSS.n6305 DVSS.n6304 0.00476
R65088 DVSS.n6306 DVSS.n6305 0.00476
R65089 DVSS.n6309 DVSS.n6306 0.00476
R65090 DVSS.n6310 DVSS.n6309 0.00476
R65091 DVSS.n6311 DVSS.n6310 0.00476
R65092 DVSS.n6312 DVSS.n6311 0.00476
R65093 DVSS.n6315 DVSS.n6312 0.00476
R65094 DVSS.n6316 DVSS.n6315 0.00476
R65095 DVSS.n6317 DVSS.n6316 0.00476
R65096 DVSS.n6317 DVSS.n19 0.00476
R65097 DVSS.n6501 DVSS.n19 0.00476
R65098 DVSS.n6509 DVSS.n9 0.00476
R65099 DVSS.n6515 DVSS.n9 0.00476
R65100 DVSS.n6516 DVSS.n6515 0.00476
R65101 DVSS.n6517 DVSS.n6516 0.00476
R65102 DVSS.n6517 DVSS.n5 0.00476
R65103 DVSS.n6523 DVSS.n5 0.00476
R65104 DVSS.n6524 DVSS.n6523 0.00476
R65105 DVSS.n6525 DVSS.n6524 0.00476
R65106 DVSS.n6525 DVSS.n1 0.00476
R65107 DVSS.n6532 DVSS.n1 0.00476
R65108 DVSS.n6533 DVSS.n6532 0.00476
R65109 DVSS.n661 DVSS.n419 0.00476
R65110 DVSS.n662 DVSS.n661 0.00476
R65111 DVSS.n663 DVSS.n662 0.00476
R65112 DVSS.n664 DVSS.n663 0.00476
R65113 DVSS.n667 DVSS.n664 0.00476
R65114 DVSS.n668 DVSS.n667 0.00476
R65115 DVSS.n669 DVSS.n668 0.00476
R65116 DVSS.n670 DVSS.n669 0.00476
R65117 DVSS.n673 DVSS.n670 0.00476
R65118 DVSS.n674 DVSS.n673 0.00476
R65119 DVSS.n675 DVSS.n674 0.00476
R65120 DVSS.n676 DVSS.n675 0.00476
R65121 DVSS.n679 DVSS.n676 0.00476
R65122 DVSS.n680 DVSS.n679 0.00476
R65123 DVSS.n680 DVSS.n442 0.00476
R65124 DVSS.n683 DVSS.n435 0.00476
R65125 DVSS.n684 DVSS.n683 0.00476
R65126 DVSS.n685 DVSS.n684 0.00476
R65127 DVSS.n717 DVSS.n685 0.00476
R65128 DVSS.n715 DVSS.n686 0.00476
R65129 DVSS.n689 DVSS.n686 0.00476
R65130 DVSS.n690 DVSS.n689 0.00476
R65131 DVSS.n691 DVSS.n690 0.00476
R65132 DVSS.n694 DVSS.n691 0.00476
R65133 DVSS.n695 DVSS.n694 0.00476
R65134 DVSS.n696 DVSS.n695 0.00476
R65135 DVSS.n697 DVSS.n696 0.00476
R65136 DVSS.n698 DVSS.n697 0.00476
R65137 DVSS.n698 DVSS.n511 0.00476
R65138 DVSS.n520 DVSS.n475 0.00476
R65139 DVSS.n521 DVSS.n520 0.00476
R65140 DVSS.n524 DVSS.n521 0.00476
R65141 DVSS.n525 DVSS.n524 0.00476
R65142 DVSS.n526 DVSS.n525 0.00476
R65143 DVSS.n527 DVSS.n526 0.00476
R65144 DVSS.n530 DVSS.n527 0.00476
R65145 DVSS.n531 DVSS.n530 0.00476
R65146 DVSS.n532 DVSS.n531 0.00476
R65147 DVSS.n533 DVSS.n532 0.00476
R65148 DVSS.n999 DVSS.n998 0.00476
R65149 DVSS.n1000 DVSS.n999 0.00476
R65150 DVSS.n1003 DVSS.n1000 0.00476
R65151 DVSS.n1004 DVSS.n1003 0.00476
R65152 DVSS.n1009 DVSS.n1006 0.00476
R65153 DVSS.n1010 DVSS.n1009 0.00476
R65154 DVSS.n1011 DVSS.n1010 0.00476
R65155 DVSS.n1012 DVSS.n1011 0.00476
R65156 DVSS.n1015 DVSS.n1012 0.00476
R65157 DVSS.n1016 DVSS.n1015 0.00476
R65158 DVSS.n1017 DVSS.n1016 0.00476
R65159 DVSS.n1018 DVSS.n1017 0.00476
R65160 DVSS.n1021 DVSS.n1018 0.00476
R65161 DVSS.n1022 DVSS.n1021 0.00476
R65162 DVSS.n1023 DVSS.n1022 0.00476
R65163 DVSS.n1024 DVSS.n1023 0.00476
R65164 DVSS.n1027 DVSS.n1024 0.00476
R65165 DVSS.n1028 DVSS.n1027 0.00476
R65166 DVSS.n1029 DVSS.n1028 0.00476
R65167 DVSS.n1034 DVSS.n1033 0.00476
R65168 DVSS.n1035 DVSS.n1034 0.00476
R65169 DVSS.n1038 DVSS.n1035 0.00476
R65170 DVSS.n1039 DVSS.n1038 0.00476
R65171 DVSS.n1040 DVSS.n1039 0.00476
R65172 DVSS.n1041 DVSS.n1040 0.00476
R65173 DVSS.n1044 DVSS.n1041 0.00476
R65174 DVSS.n1045 DVSS.n1044 0.00476
R65175 DVSS.n1046 DVSS.n1045 0.00476
R65176 DVSS.n1047 DVSS.n1046 0.00476
R65177 DVSS.n753 DVSS.n752 0.00476
R65178 DVSS.n752 DVSS.n751 0.00476
R65179 DVSS.n751 DVSS.n659 0.00476
R65180 DVSS.n747 DVSS.n659 0.00476
R65181 DVSS.n747 DVSS.n746 0.00476
R65182 DVSS.n746 DVSS.n745 0.00476
R65183 DVSS.n745 DVSS.n665 0.00476
R65184 DVSS.n741 DVSS.n665 0.00476
R65185 DVSS.n741 DVSS.n740 0.00476
R65186 DVSS.n740 DVSS.n739 0.00476
R65187 DVSS.n739 DVSS.n671 0.00476
R65188 DVSS.n735 DVSS.n671 0.00476
R65189 DVSS.n735 DVSS.n734 0.00476
R65190 DVSS.n734 DVSS.n733 0.00476
R65191 DVSS.n733 DVSS.n677 0.00476
R65192 DVSS.n729 DVSS.n677 0.00476
R65193 DVSS.n729 DVSS.n728 0.00476
R65194 DVSS.n728 DVSS.n727 0.00476
R65195 DVSS.n727 DVSS.n681 0.00476
R65196 DVSS.n723 DVSS.n681 0.00476
R65197 DVSS.n723 DVSS.n722 0.00476
R65198 DVSS.n722 DVSS.n721 0.00476
R65199 DVSS.n721 DVSS.n718 0.00476
R65200 DVSS.n714 DVSS.n687 0.00476
R65201 DVSS.n710 DVSS.n687 0.00476
R65202 DVSS.n710 DVSS.n709 0.00476
R65203 DVSS.n709 DVSS.n708 0.00476
R65204 DVSS.n708 DVSS.n692 0.00476
R65205 DVSS.n704 DVSS.n692 0.00476
R65206 DVSS.n704 DVSS.n703 0.00476
R65207 DVSS.n703 DVSS.n702 0.00476
R65208 DVSS.n702 DVSS.n699 0.00476
R65209 DVSS.n699 DVSS.n516 0.00476
R65210 DVSS.n6187 DVSS.n516 0.00476
R65211 DVSS.n6187 DVSS.n517 0.00476
R65212 DVSS.n6183 DVSS.n517 0.00476
R65213 DVSS.n6183 DVSS.n6182 0.00476
R65214 DVSS.n6182 DVSS.n6181 0.00476
R65215 DVSS.n6181 DVSS.n522 0.00476
R65216 DVSS.n6177 DVSS.n522 0.00476
R65217 DVSS.n6177 DVSS.n6176 0.00476
R65218 DVSS.n6176 DVSS.n6175 0.00476
R65219 DVSS.n6175 DVSS.n528 0.00476
R65220 DVSS.n6171 DVSS.n528 0.00476
R65221 DVSS.n6171 DVSS.n6170 0.00476
R65222 DVSS.n6170 DVSS.n6169 0.00476
R65223 DVSS.n6165 DVSS.n6164 0.00476
R65224 DVSS.n6164 DVSS.n6163 0.00476
R65225 DVSS.n6163 DVSS.n1001 0.00476
R65226 DVSS.n6159 DVSS.n1001 0.00476
R65227 DVSS.n6159 DVSS.n6158 0.00476
R65228 DVSS.n6158 DVSS.n6157 0.00476
R65229 DVSS.n6157 DVSS.n1007 0.00476
R65230 DVSS.n6153 DVSS.n1007 0.00476
R65231 DVSS.n6153 DVSS.n6152 0.00476
R65232 DVSS.n6152 DVSS.n6151 0.00476
R65233 DVSS.n6151 DVSS.n1013 0.00476
R65234 DVSS.n6147 DVSS.n1013 0.00476
R65235 DVSS.n6147 DVSS.n6146 0.00476
R65236 DVSS.n6146 DVSS.n6145 0.00476
R65237 DVSS.n6145 DVSS.n1019 0.00476
R65238 DVSS.n6141 DVSS.n1019 0.00476
R65239 DVSS.n6141 DVSS.n6140 0.00476
R65240 DVSS.n6140 DVSS.n6139 0.00476
R65241 DVSS.n6139 DVSS.n1025 0.00476
R65242 DVSS.n6135 DVSS.n1025 0.00476
R65243 DVSS.n6135 DVSS.n6134 0.00476
R65244 DVSS.n6134 DVSS.n6133 0.00476
R65245 DVSS.n6133 DVSS.n1070 0.00476
R65246 DVSS.n1066 DVSS.n1065 0.00476
R65247 DVSS.n1065 DVSS.n1064 0.00476
R65248 DVSS.n1064 DVSS.n1036 0.00476
R65249 DVSS.n1060 DVSS.n1036 0.00476
R65250 DVSS.n1060 DVSS.n1059 0.00476
R65251 DVSS.n1059 DVSS.n1058 0.00476
R65252 DVSS.n1058 DVSS.n1042 0.00476
R65253 DVSS.n1054 DVSS.n1042 0.00476
R65254 DVSS.n1054 DVSS.n1053 0.00476
R65255 DVSS.n1053 DVSS.n1052 0.00476
R65256 DVSS.n759 DVSS.n586 0.00476
R65257 DVSS.n760 DVSS.n759 0.00476
R65258 DVSS.n762 DVSS.n760 0.00476
R65259 DVSS.n762 DVSS.n584 0.00476
R65260 DVSS.n766 DVSS.n584 0.00476
R65261 DVSS.n766 DVSS.n582 0.00476
R65262 DVSS.n770 DVSS.n582 0.00476
R65263 DVSS.n770 DVSS.n580 0.00476
R65264 DVSS.n774 DVSS.n580 0.00476
R65265 DVSS.n774 DVSS.n578 0.00476
R65266 DVSS.n778 DVSS.n578 0.00476
R65267 DVSS.n778 DVSS.n576 0.00476
R65268 DVSS.n782 DVSS.n576 0.00476
R65269 DVSS.n782 DVSS.n574 0.00476
R65270 DVSS.n787 DVSS.n574 0.00476
R65271 DVSS.n787 DVSS.n572 0.00476
R65272 DVSS.n791 DVSS.n572 0.00476
R65273 DVSS.n792 DVSS.n791 0.00476
R65274 DVSS.n793 DVSS.n792 0.00476
R65275 DVSS.n793 DVSS.n570 0.00476
R65276 DVSS.n798 DVSS.n570 0.00476
R65277 DVSS.n798 DVSS.n568 0.00476
R65278 DVSS.n802 DVSS.n568 0.00476
R65279 DVSS.n835 DVSS.n834 0.00476
R65280 DVSS.n834 DVSS.n833 0.00476
R65281 DVSS.n833 DVSS.n807 0.00476
R65282 DVSS.n829 DVSS.n807 0.00476
R65283 DVSS.n829 DVSS.n828 0.00476
R65284 DVSS.n828 DVSS.n827 0.00476
R65285 DVSS.n827 DVSS.n813 0.00476
R65286 DVSS.n823 DVSS.n813 0.00476
R65287 DVSS.n823 DVSS.n822 0.00476
R65288 DVSS.n822 DVSS.n821 0.00476
R65289 DVSS.n821 DVSS.n818 0.00476
R65290 DVSS.n818 DVSS.n325 0.00476
R65291 DVSS.n6365 DVSS.n325 0.00476
R65292 DVSS.n6365 DVSS.n326 0.00476
R65293 DVSS.n6361 DVSS.n326 0.00476
R65294 DVSS.n6361 DVSS.n6360 0.00476
R65295 DVSS.n6360 DVSS.n6359 0.00476
R65296 DVSS.n6359 DVSS.n332 0.00476
R65297 DVSS.n6355 DVSS.n332 0.00476
R65298 DVSS.n6355 DVSS.n6354 0.00476
R65299 DVSS.n6354 DVSS.n6353 0.00476
R65300 DVSS.n6353 DVSS.n338 0.00476
R65301 DVSS.n6349 DVSS.n338 0.00476
R65302 DVSS.n6347 DVSS.n345 0.00476
R65303 DVSS.n6343 DVSS.n345 0.00476
R65304 DVSS.n6343 DVSS.n6342 0.00476
R65305 DVSS.n6342 DVSS.n6341 0.00476
R65306 DVSS.n6341 DVSS.n351 0.00476
R65307 DVSS.n6337 DVSS.n351 0.00476
R65308 DVSS.n6337 DVSS.n6336 0.00476
R65309 DVSS.n6336 DVSS.n6335 0.00476
R65310 DVSS.n6335 DVSS.n6301 0.00476
R65311 DVSS.n6331 DVSS.n6301 0.00476
R65312 DVSS.n6331 DVSS.n6330 0.00476
R65313 DVSS.n6330 DVSS.n6329 0.00476
R65314 DVSS.n6329 DVSS.n6307 0.00476
R65315 DVSS.n6325 DVSS.n6307 0.00476
R65316 DVSS.n6325 DVSS.n6324 0.00476
R65317 DVSS.n6324 DVSS.n6323 0.00476
R65318 DVSS.n6323 DVSS.n6313 0.00476
R65319 DVSS.n6319 DVSS.n6313 0.00476
R65320 DVSS.n6319 DVSS.n6318 0.00476
R65321 DVSS.n6318 DVSS.n18 0.00476
R65322 DVSS.n6502 DVSS.n18 0.00476
R65323 DVSS.n6502 DVSS.n16 0.00476
R65324 DVSS.n6506 DVSS.n16 0.00476
R65325 DVSS.n6510 DVSS.n10 0.00476
R65326 DVSS.n6514 DVSS.n10 0.00476
R65327 DVSS.n6514 DVSS.n8 0.00476
R65328 DVSS.n6518 DVSS.n8 0.00476
R65329 DVSS.n6518 DVSS.n6 0.00476
R65330 DVSS.n6522 DVSS.n6 0.00476
R65331 DVSS.n6522 DVSS.n4 0.00476
R65332 DVSS.n6526 DVSS.n4 0.00476
R65333 DVSS.n6526 DVSS.n2 0.00476
R65334 DVSS.n6531 DVSS.n2 0.00476
R65335 DVSS.n6531 DVSS.n0 0.00476
R65336 DVSS.n655 DVSS.n596 0.00476
R65337 DVSS.n651 DVSS.n596 0.00476
R65338 DVSS.n651 DVSS.n650 0.00476
R65339 DVSS.n650 DVSS.n649 0.00476
R65340 DVSS.n649 DVSS.n600 0.00476
R65341 DVSS.n645 DVSS.n600 0.00476
R65342 DVSS.n645 DVSS.n644 0.00476
R65343 DVSS.n644 DVSS.n643 0.00476
R65344 DVSS.n643 DVSS.n606 0.00476
R65345 DVSS.n639 DVSS.n606 0.00476
R65346 DVSS.n639 DVSS.n638 0.00476
R65347 DVSS.n638 DVSS.n637 0.00476
R65348 DVSS.n637 DVSS.n612 0.00476
R65349 DVSS.n633 DVSS.n612 0.00476
R65350 DVSS.n633 DVSS.n632 0.00476
R65351 DVSS.n632 DVSS.n631 0.00476
R65352 DVSS.n631 DVSS.n618 0.00476
R65353 DVSS.n627 DVSS.n618 0.00476
R65354 DVSS.n627 DVSS.n626 0.00476
R65355 DVSS.n626 DVSS.n625 0.00476
R65356 DVSS.n625 DVSS.n622 0.00476
R65357 DVSS.n622 DVSS.n561 0.00476
R65358 DVSS.n840 DVSS.n561 0.00476
R65359 DVSS.n845 DVSS.n558 0.00476
R65360 DVSS.n845 DVSS.n556 0.00476
R65361 DVSS.n849 DVSS.n556 0.00476
R65362 DVSS.n849 DVSS.n554 0.00476
R65363 DVSS.n853 DVSS.n554 0.00476
R65364 DVSS.n853 DVSS.n552 0.00476
R65365 DVSS.n858 DVSS.n552 0.00476
R65366 DVSS.n858 DVSS.n550 0.00476
R65367 DVSS.n862 DVSS.n550 0.00476
R65368 DVSS.n863 DVSS.n862 0.00476
R65369 DVSS.n863 DVSS.n547 0.00476
R65370 DVSS.n867 DVSS.n547 0.00476
R65371 DVSS.n868 DVSS.n867 0.00476
R65372 DVSS.n871 DVSS.n868 0.00476
R65373 DVSS.n871 DVSS.n545 0.00476
R65374 DVSS.n875 DVSS.n545 0.00476
R65375 DVSS.n875 DVSS.n543 0.00476
R65376 DVSS.n879 DVSS.n543 0.00476
R65377 DVSS.n879 DVSS.n541 0.00476
R65378 DVSS.n884 DVSS.n541 0.00476
R65379 DVSS.n884 DVSS.n539 0.00476
R65380 DVSS.n888 DVSS.n539 0.00476
R65381 DVSS.n889 DVSS.n888 0.00476
R65382 DVSS.n993 DVSS.n537 0.00476
R65383 DVSS.n989 DVSS.n537 0.00476
R65384 DVSS.n989 DVSS.n988 0.00476
R65385 DVSS.n988 DVSS.n987 0.00476
R65386 DVSS.n987 DVSS.n896 0.00476
R65387 DVSS.n983 DVSS.n896 0.00476
R65388 DVSS.n983 DVSS.n982 0.00476
R65389 DVSS.n982 DVSS.n981 0.00476
R65390 DVSS.n981 DVSS.n900 0.00476
R65391 DVSS.n977 DVSS.n900 0.00476
R65392 DVSS.n977 DVSS.n976 0.00476
R65393 DVSS.n976 DVSS.n975 0.00476
R65394 DVSS.n975 DVSS.n906 0.00476
R65395 DVSS.n971 DVSS.n906 0.00476
R65396 DVSS.n971 DVSS.n970 0.00476
R65397 DVSS.n970 DVSS.n969 0.00476
R65398 DVSS.n969 DVSS.n912 0.00476
R65399 DVSS.n965 DVSS.n912 0.00476
R65400 DVSS.n965 DVSS.n964 0.00476
R65401 DVSS.n964 DVSS.n963 0.00476
R65402 DVSS.n963 DVSS.n918 0.00476
R65403 DVSS.n959 DVSS.n918 0.00476
R65404 DVSS.n959 DVSS.n958 0.00476
R65405 DVSS.n956 DVSS.n921 0.00476
R65406 DVSS.n952 DVSS.n921 0.00476
R65407 DVSS.n952 DVSS.n951 0.00476
R65408 DVSS.n951 DVSS.n950 0.00476
R65409 DVSS.n950 DVSS.n928 0.00476
R65410 DVSS.n946 DVSS.n928 0.00476
R65411 DVSS.n946 DVSS.n945 0.00476
R65412 DVSS.n945 DVSS.n944 0.00476
R65413 DVSS.n944 DVSS.n934 0.00476
R65414 DVSS.n940 DVSS.n934 0.00476
R65415 DVSS.n2369 DVSS.n2368 0.00468605
R65416 DVSS.n1466 DVSS 0.00464676
R65417 DVSS DVSS.n4128 0.00460473
R65418 DVSS DVSS.n937 0.00458
R65419 DVSS.n940 DVSS 0.00458
R65420 DVSS.n5266 DVSS.n5265 0.00455
R65421 DVSS.n2925 DVSS.n2600 0.00455
R65422 DVSS.n3062 DVSS.n3061 0.00455
R65423 DVSS.n3013 DVSS.n2394 0.00455
R65424 DVSS.n2465 DVSS.n2393 0.00455
R65425 DVSS.n895 DVSS.n207 0.00455
R65426 DVSS.n6294 DVSS.n350 0.00455
R65427 DVSS.n1004 DVSS.n390 0.00455
R65428 DVSS.n837 DVSS.n564 0.0045
R65429 DVSS.n6167 DVSS.n339 0.0045
R65430 DVSS.n756 DVSS.n587 0.0045
R65431 DVSS.n838 DVSS.n837 0.0045
R65432 DVSS.n891 DVSS.n339 0.0045
R65433 DVSS.n1068 DVSS.n11 0.0045
R65434 DVSS.n922 DVSS.n11 0.0045
R65435 DVSS.n756 DVSS.n755 0.0045
R65436 DVSS.n3289 DVSS.n3282 0.00448437
R65437 DVSS.n4639 DVSS.n2028 0.00443
R65438 DVSS.n6470 DVSS.n134 0.00443
R65439 DVSS.n6476 DVSS.n102 0.00443
R65440 DVSS.n6232 DVSS.n435 0.00443
R65441 DVSS.n2472 DVSS.n2457 0.00437324
R65442 DVSS.n5792 DVSS.n1172 0.00419403
R65443 DVSS.n6406 DVSS.n160 0.00419403
R65444 DVSS.n1756 DVSS.n1728 0.0041
R65445 DVSS.n1757 DVSS.n1719 0.0041
R65446 DVSS.n4984 DVSS.n1727 0.0041
R65447 DVSS.n4946 DVSS.n1794 0.0041
R65448 DVSS.n1797 DVSS.n1796 0.0041
R65449 DVSS.n4944 DVSS.n4943 0.0041
R65450 DVSS.n2928 DVSS.n2599 0.00409155
R65451 DVSS.n920 DVSS.n14 0.00404
R65452 DVSS.n6509 DVSS.n6508 0.00404
R65453 DVSS.n1033 DVSS.n13 0.00404
R65454 DVSS.n1066 DVSS.n1031 0.00404
R65455 DVSS.n6510 DVSS.n12 0.00404
R65456 DVSS.n957 DVSS.n956 0.00404
R65457 DVSS.n3543 DVSS.n2098 0.00403571
R65458 DVSS.n3692 DVSS.n2084 0.00403571
R65459 DVSS.n3883 DVSS.n2070 0.00403571
R65460 DVSS.n3941 DVSS.n3896 0.00403571
R65461 DVSS.n6093 DVSS.n1159 0.00403571
R65462 DVSS.n4594 DVSS.n4550 0.00401
R65463 DVSS.n5264 DVSS.n1564 0.00401
R65464 DVSS.n548 DVSS.n152 0.00401
R65465 DVSS.n6439 DVSS.n183 0.00401
R65466 DVSS.n6371 DVSS.n321 0.00401
R65467 DVSS.n6297 DVSS.n353 0.00401
R65468 DVSS.n6199 DVSS.n466 0.00401
R65469 DVSS.n1005 DVSS.n389 0.00401
R65470 DVSS.n5324 DVSS 0.00392
R65471 DVSS DVSS.n5317 0.00392
R65472 DVSS DVSS.n1047 0.00392
R65473 DVSS.n1052 DVSS 0.00392
R65474 DVSS.n4369 DVSS.n4367 0.00391292
R65475 DVSS.n5255 DVSS.n1601 0.00391292
R65476 DVSS.n4636 DVSS.n2027 0.00389
R65477 DVSS.n4597 DVSS.n4501 0.00389
R65478 DVSS.n6472 DVSS.n117 0.00389
R65479 DVSS.n6460 DVSS.n166 0.00389
R65480 DVSS.n6479 DVSS.n88 0.00389
R65481 DVSS.n6373 DVSS.n299 0.00389
R65482 DVSS.n6229 DVSS.n428 0.00389
R65483 DVSS.n6196 DVSS.n6188 0.00389
R65484 DVSS.n995 DVSS.n994 0.0038
R65485 DVSS.n996 DVSS.n344 0.0038
R65486 DVSS.n998 DVSS.n997 0.0038
R65487 DVSS.n6165 DVSS.n342 0.0038
R65488 DVSS.n6348 DVSS.n6347 0.0038
R65489 DVSS.n993 DVSS.n343 0.0038
R65490 DVSS.n2880 DVSS.n2609 0.00377857
R65491 DVSS.n5085 DVSS.n5084 0.00377857
R65492 DVSS.n5131 DVSS.n5130 0.00377857
R65493 DVSS.n5552 DVSS.n5551 0.00377857
R65494 DVSS.n1185 DVSS.n1183 0.00377857
R65495 DVSS.n843 DVSS.n842 0.00356
R65496 DVSS.n804 DVSS.n559 0.00356
R65497 DVSS.n716 DVSS.n715 0.00356
R65498 DVSS.n714 DVSS.n567 0.00356
R65499 DVSS.n835 DVSS.n803 0.00356
R65500 DVSS.n562 DVSS.n558 0.00356
R65501 DVSS DVSS.n1900 0.00353371
R65502 DVSS.n6201 DVSS.n461 0.00352239
R65503 DVSS.n6264 DVSS.n296 0.00352239
R65504 DVSS.n2382 DVSS.n2381 0.00346697
R65505 DVSS.n654 DVSS.n653 0.00334
R65506 DVSS.n653 DVSS.n652 0.00334
R65507 DVSS.n652 DVSS.n597 0.00334
R65508 DVSS.n648 DVSS.n597 0.00334
R65509 DVSS.n648 DVSS.n647 0.00334
R65510 DVSS.n647 DVSS.n646 0.00334
R65511 DVSS.n646 DVSS.n601 0.00334
R65512 DVSS.n642 DVSS.n601 0.00334
R65513 DVSS.n642 DVSS.n641 0.00334
R65514 DVSS.n641 DVSS.n640 0.00334
R65515 DVSS.n640 DVSS.n607 0.00334
R65516 DVSS.n636 DVSS.n607 0.00334
R65517 DVSS.n636 DVSS.n635 0.00334
R65518 DVSS.n635 DVSS.n634 0.00334
R65519 DVSS.n634 DVSS.n613 0.00334
R65520 DVSS.n630 DVSS.n613 0.00334
R65521 DVSS.n630 DVSS.n629 0.00334
R65522 DVSS.n629 DVSS.n628 0.00334
R65523 DVSS.n628 DVSS.n619 0.00334
R65524 DVSS.n624 DVSS.n619 0.00334
R65525 DVSS.n624 DVSS.n623 0.00334
R65526 DVSS.n623 DVSS.n563 0.00334
R65527 DVSS.n839 DVSS.n563 0.00334
R65528 DVSS.n846 DVSS.n557 0.00334
R65529 DVSS.n847 DVSS.n846 0.00334
R65530 DVSS.n848 DVSS.n847 0.00334
R65531 DVSS.n848 DVSS.n553 0.00334
R65532 DVSS.n854 DVSS.n553 0.00334
R65533 DVSS.n855 DVSS.n854 0.00334
R65534 DVSS.n857 DVSS.n855 0.00334
R65535 DVSS.n857 DVSS.n856 0.00334
R65536 DVSS.n856 DVSS.n549 0.00334
R65537 DVSS.n864 DVSS.n549 0.00334
R65538 DVSS.n865 DVSS.n864 0.00334
R65539 DVSS.n866 DVSS.n865 0.00334
R65540 DVSS.n866 DVSS.n546 0.00334
R65541 DVSS.n872 DVSS.n546 0.00334
R65542 DVSS.n873 DVSS.n872 0.00334
R65543 DVSS.n874 DVSS.n873 0.00334
R65544 DVSS.n874 DVSS.n542 0.00334
R65545 DVSS.n880 DVSS.n542 0.00334
R65546 DVSS.n881 DVSS.n880 0.00334
R65547 DVSS.n883 DVSS.n881 0.00334
R65548 DVSS.n883 DVSS.n882 0.00334
R65549 DVSS.n882 DVSS.n538 0.00334
R65550 DVSS.n890 DVSS.n538 0.00334
R65551 DVSS.n992 DVSS.n991 0.00334
R65552 DVSS.n991 DVSS.n990 0.00334
R65553 DVSS.n990 DVSS.n892 0.00334
R65554 DVSS.n986 DVSS.n892 0.00334
R65555 DVSS.n986 DVSS.n985 0.00334
R65556 DVSS.n985 DVSS.n984 0.00334
R65557 DVSS.n984 DVSS.n897 0.00334
R65558 DVSS.n980 DVSS.n897 0.00334
R65559 DVSS.n980 DVSS.n979 0.00334
R65560 DVSS.n979 DVSS.n978 0.00334
R65561 DVSS.n978 DVSS.n901 0.00334
R65562 DVSS.n974 DVSS.n901 0.00334
R65563 DVSS.n974 DVSS.n973 0.00334
R65564 DVSS.n973 DVSS.n972 0.00334
R65565 DVSS.n972 DVSS.n907 0.00334
R65566 DVSS.n968 DVSS.n907 0.00334
R65567 DVSS.n968 DVSS.n967 0.00334
R65568 DVSS.n967 DVSS.n966 0.00334
R65569 DVSS.n966 DVSS.n913 0.00334
R65570 DVSS.n962 DVSS.n913 0.00334
R65571 DVSS.n962 DVSS.n961 0.00334
R65572 DVSS.n961 DVSS.n960 0.00334
R65573 DVSS.n960 DVSS.n919 0.00334
R65574 DVSS.n955 DVSS.n954 0.00334
R65575 DVSS.n954 DVSS.n953 0.00334
R65576 DVSS.n953 DVSS.n923 0.00334
R65577 DVSS.n949 DVSS.n923 0.00334
R65578 DVSS.n949 DVSS.n948 0.00334
R65579 DVSS.n948 DVSS.n947 0.00334
R65580 DVSS.n947 DVSS.n929 0.00334
R65581 DVSS.n943 DVSS.n929 0.00334
R65582 DVSS.n943 DVSS.n942 0.00334
R65583 DVSS.n942 DVSS.n941 0.00334
R65584 DVSS.n941 DVSS.n935 0.00334
R65585 DVSS.n758 DVSS.n757 0.00334
R65586 DVSS.n758 DVSS.n585 0.00334
R65587 DVSS.n763 DVSS.n585 0.00334
R65588 DVSS.n764 DVSS.n763 0.00334
R65589 DVSS.n765 DVSS.n764 0.00334
R65590 DVSS.n765 DVSS.n581 0.00334
R65591 DVSS.n771 DVSS.n581 0.00334
R65592 DVSS.n772 DVSS.n771 0.00334
R65593 DVSS.n773 DVSS.n772 0.00334
R65594 DVSS.n773 DVSS.n577 0.00334
R65595 DVSS.n779 DVSS.n577 0.00334
R65596 DVSS.n780 DVSS.n779 0.00334
R65597 DVSS.n781 DVSS.n780 0.00334
R65598 DVSS.n781 DVSS.n573 0.00334
R65599 DVSS.n788 DVSS.n573 0.00334
R65600 DVSS.n789 DVSS.n788 0.00334
R65601 DVSS.n790 DVSS.n789 0.00334
R65602 DVSS.n790 DVSS.n571 0.00334
R65603 DVSS.n794 DVSS.n571 0.00334
R65604 DVSS.n795 DVSS.n794 0.00334
R65605 DVSS.n797 DVSS.n795 0.00334
R65606 DVSS.n797 DVSS.n796 0.00334
R65607 DVSS.n796 DVSS.n565 0.00334
R65608 DVSS.n836 DVSS.n566 0.00334
R65609 DVSS.n832 DVSS.n566 0.00334
R65610 DVSS.n832 DVSS.n831 0.00334
R65611 DVSS.n831 DVSS.n830 0.00334
R65612 DVSS.n830 DVSS.n808 0.00334
R65613 DVSS.n826 DVSS.n808 0.00334
R65614 DVSS.n826 DVSS.n825 0.00334
R65615 DVSS.n825 DVSS.n824 0.00334
R65616 DVSS.n824 DVSS.n814 0.00334
R65617 DVSS.n820 DVSS.n814 0.00334
R65618 DVSS.n820 DVSS.n819 0.00334
R65619 DVSS.n819 DVSS.n327 0.00334
R65620 DVSS.n6364 DVSS.n327 0.00334
R65621 DVSS.n6364 DVSS.n6363 0.00334
R65622 DVSS.n6363 DVSS.n6362 0.00334
R65623 DVSS.n6362 DVSS.n328 0.00334
R65624 DVSS.n6358 DVSS.n328 0.00334
R65625 DVSS.n6358 DVSS.n6357 0.00334
R65626 DVSS.n6357 DVSS.n6356 0.00334
R65627 DVSS.n6356 DVSS.n333 0.00334
R65628 DVSS.n6352 DVSS.n333 0.00334
R65629 DVSS.n6352 DVSS.n6351 0.00334
R65630 DVSS.n6351 DVSS.n6350 0.00334
R65631 DVSS.n6346 DVSS.n6345 0.00334
R65632 DVSS.n6345 DVSS.n6344 0.00334
R65633 DVSS.n6344 DVSS.n346 0.00334
R65634 DVSS.n6340 DVSS.n346 0.00334
R65635 DVSS.n6340 DVSS.n6339 0.00334
R65636 DVSS.n6339 DVSS.n6338 0.00334
R65637 DVSS.n6338 DVSS.n352 0.00334
R65638 DVSS.n6334 DVSS.n352 0.00334
R65639 DVSS.n6334 DVSS.n6333 0.00334
R65640 DVSS.n6333 DVSS.n6332 0.00334
R65641 DVSS.n6332 DVSS.n6302 0.00334
R65642 DVSS.n6328 DVSS.n6302 0.00334
R65643 DVSS.n6328 DVSS.n6327 0.00334
R65644 DVSS.n6327 DVSS.n6326 0.00334
R65645 DVSS.n6326 DVSS.n6308 0.00334
R65646 DVSS.n6322 DVSS.n6308 0.00334
R65647 DVSS.n6322 DVSS.n6321 0.00334
R65648 DVSS.n6321 DVSS.n6320 0.00334
R65649 DVSS.n6320 DVSS.n6314 0.00334
R65650 DVSS.n6314 DVSS.n17 0.00334
R65651 DVSS.n6503 DVSS.n17 0.00334
R65652 DVSS.n6504 DVSS.n6503 0.00334
R65653 DVSS.n6505 DVSS.n6504 0.00334
R65654 DVSS.n6512 DVSS.n6511 0.00334
R65655 DVSS.n6513 DVSS.n6512 0.00334
R65656 DVSS.n6513 DVSS.n7 0.00334
R65657 DVSS.n6519 DVSS.n7 0.00334
R65658 DVSS.n6520 DVSS.n6519 0.00334
R65659 DVSS.n6521 DVSS.n6520 0.00334
R65660 DVSS.n6521 DVSS.n3 0.00334
R65661 DVSS.n6527 DVSS.n3 0.00334
R65662 DVSS.n6528 DVSS.n6527 0.00334
R65663 DVSS.n6530 DVSS.n6528 0.00334
R65664 DVSS.n6530 DVSS.n6529 0.00334
R65665 DVSS.n754 DVSS.n590 0.00334
R65666 DVSS.n750 DVSS.n590 0.00334
R65667 DVSS.n750 DVSS.n749 0.00334
R65668 DVSS.n749 DVSS.n748 0.00334
R65669 DVSS.n748 DVSS.n660 0.00334
R65670 DVSS.n744 DVSS.n660 0.00334
R65671 DVSS.n744 DVSS.n743 0.00334
R65672 DVSS.n743 DVSS.n742 0.00334
R65673 DVSS.n742 DVSS.n666 0.00334
R65674 DVSS.n738 DVSS.n666 0.00334
R65675 DVSS.n738 DVSS.n737 0.00334
R65676 DVSS.n737 DVSS.n736 0.00334
R65677 DVSS.n736 DVSS.n672 0.00334
R65678 DVSS.n732 DVSS.n672 0.00334
R65679 DVSS.n732 DVSS.n731 0.00334
R65680 DVSS.n731 DVSS.n730 0.00334
R65681 DVSS.n730 DVSS.n678 0.00334
R65682 DVSS.n726 DVSS.n678 0.00334
R65683 DVSS.n726 DVSS.n725 0.00334
R65684 DVSS.n725 DVSS.n724 0.00334
R65685 DVSS.n724 DVSS.n682 0.00334
R65686 DVSS.n720 DVSS.n682 0.00334
R65687 DVSS.n720 DVSS.n719 0.00334
R65688 DVSS.n713 DVSS.n712 0.00334
R65689 DVSS.n712 DVSS.n711 0.00334
R65690 DVSS.n711 DVSS.n688 0.00334
R65691 DVSS.n707 DVSS.n688 0.00334
R65692 DVSS.n707 DVSS.n706 0.00334
R65693 DVSS.n706 DVSS.n705 0.00334
R65694 DVSS.n705 DVSS.n693 0.00334
R65695 DVSS.n701 DVSS.n693 0.00334
R65696 DVSS.n701 DVSS.n700 0.00334
R65697 DVSS.n700 DVSS.n518 0.00334
R65698 DVSS.n6186 DVSS.n518 0.00334
R65699 DVSS.n6186 DVSS.n6185 0.00334
R65700 DVSS.n6185 DVSS.n6184 0.00334
R65701 DVSS.n6184 DVSS.n519 0.00334
R65702 DVSS.n6180 DVSS.n519 0.00334
R65703 DVSS.n6180 DVSS.n6179 0.00334
R65704 DVSS.n6179 DVSS.n6178 0.00334
R65705 DVSS.n6178 DVSS.n523 0.00334
R65706 DVSS.n6174 DVSS.n523 0.00334
R65707 DVSS.n6174 DVSS.n6173 0.00334
R65708 DVSS.n6173 DVSS.n6172 0.00334
R65709 DVSS.n6172 DVSS.n529 0.00334
R65710 DVSS.n6168 DVSS.n529 0.00334
R65711 DVSS.n6166 DVSS.n534 0.00334
R65712 DVSS.n6162 DVSS.n534 0.00334
R65713 DVSS.n6162 DVSS.n6161 0.00334
R65714 DVSS.n6161 DVSS.n6160 0.00334
R65715 DVSS.n6160 DVSS.n1002 0.00334
R65716 DVSS.n6156 DVSS.n1002 0.00334
R65717 DVSS.n6156 DVSS.n6155 0.00334
R65718 DVSS.n6155 DVSS.n6154 0.00334
R65719 DVSS.n6154 DVSS.n1008 0.00334
R65720 DVSS.n6150 DVSS.n1008 0.00334
R65721 DVSS.n6150 DVSS.n6149 0.00334
R65722 DVSS.n6149 DVSS.n6148 0.00334
R65723 DVSS.n6148 DVSS.n1014 0.00334
R65724 DVSS.n6144 DVSS.n1014 0.00334
R65725 DVSS.n6144 DVSS.n6143 0.00334
R65726 DVSS.n6143 DVSS.n6142 0.00334
R65727 DVSS.n6142 DVSS.n1020 0.00334
R65728 DVSS.n6138 DVSS.n1020 0.00334
R65729 DVSS.n6138 DVSS.n6137 0.00334
R65730 DVSS.n6137 DVSS.n6136 0.00334
R65731 DVSS.n6136 DVSS.n1026 0.00334
R65732 DVSS.n1030 DVSS.n1026 0.00334
R65733 DVSS.n1069 DVSS.n1030 0.00334
R65734 DVSS.n1067 DVSS.n1032 0.00334
R65735 DVSS.n1063 DVSS.n1032 0.00334
R65736 DVSS.n1063 DVSS.n1062 0.00334
R65737 DVSS.n1062 DVSS.n1061 0.00334
R65738 DVSS.n1061 DVSS.n1037 0.00334
R65739 DVSS.n1057 DVSS.n1037 0.00334
R65740 DVSS.n1057 DVSS.n1056 0.00334
R65741 DVSS.n1056 DVSS.n1055 0.00334
R65742 DVSS.n1055 DVSS.n1043 0.00334
R65743 DVSS.n1051 DVSS.n1043 0.00334
R65744 DVSS.n1051 DVSS.n1050 0.00334
R65745 DVSS.n4452 DVSS.n2054 0.00334
R65746 DVSS.n4453 DVSS.n4452 0.00334
R65747 DVSS.n4454 DVSS.n4453 0.00334
R65748 DVSS.n4454 DVSS.n2050 0.00334
R65749 DVSS.n4460 DVSS.n2050 0.00334
R65750 DVSS.n4461 DVSS.n4460 0.00334
R65751 DVSS.n4462 DVSS.n4461 0.00334
R65752 DVSS.n4462 DVSS.n2046 0.00334
R65753 DVSS.n4468 DVSS.n2046 0.00334
R65754 DVSS.n4469 DVSS.n4468 0.00334
R65755 DVSS.n4470 DVSS.n4469 0.00334
R65756 DVSS.n4470 DVSS.n2042 0.00334
R65757 DVSS.n4476 DVSS.n2042 0.00334
R65758 DVSS.n4477 DVSS.n4476 0.00334
R65759 DVSS.n4478 DVSS.n4477 0.00334
R65760 DVSS.n4479 DVSS.n4478 0.00334
R65761 DVSS.n4480 DVSS.n4479 0.00334
R65762 DVSS.n4481 DVSS.n4480 0.00334
R65763 DVSS.n4484 DVSS.n4481 0.00334
R65764 DVSS.n4485 DVSS.n4484 0.00334
R65765 DVSS.n4486 DVSS.n4485 0.00334
R65766 DVSS.n4487 DVSS.n4486 0.00334
R65767 DVSS.n4490 DVSS.n4487 0.00334
R65768 DVSS.n4491 DVSS.n4490 0.00334
R65769 DVSS.n4492 DVSS.n4491 0.00334
R65770 DVSS.n4493 DVSS.n4492 0.00334
R65771 DVSS.n4496 DVSS.n4493 0.00334
R65772 DVSS.n4497 DVSS.n4496 0.00334
R65773 DVSS.n4498 DVSS.n4497 0.00334
R65774 DVSS.n4499 DVSS.n4498 0.00334
R65775 DVSS.n4502 DVSS.n4499 0.00334
R65776 DVSS.n4503 DVSS.n4502 0.00334
R65777 DVSS.n4504 DVSS.n4503 0.00334
R65778 DVSS.n4552 DVSS.n4504 0.00334
R65779 DVSS.n4553 DVSS.n4552 0.00334
R65780 DVSS.n4554 DVSS.n4553 0.00334
R65781 DVSS.n4555 DVSS.n4554 0.00334
R65782 DVSS.n4558 DVSS.n4555 0.00334
R65783 DVSS.n4559 DVSS.n4558 0.00334
R65784 DVSS.n4560 DVSS.n4559 0.00334
R65785 DVSS.n4561 DVSS.n4560 0.00334
R65786 DVSS.n4564 DVSS.n4561 0.00334
R65787 DVSS.n4565 DVSS.n4564 0.00334
R65788 DVSS.n4566 DVSS.n4565 0.00334
R65789 DVSS.n4567 DVSS.n4566 0.00334
R65790 DVSS.n4570 DVSS.n4567 0.00334
R65791 DVSS.n4571 DVSS.n4570 0.00334
R65792 DVSS.n4572 DVSS.n4571 0.00334
R65793 DVSS.n4572 DVSS.n1566 0.00334
R65794 DVSS.n5268 DVSS.n1566 0.00334
R65795 DVSS.n5269 DVSS.n5268 0.00334
R65796 DVSS.n5270 DVSS.n5269 0.00334
R65797 DVSS.n5270 DVSS.n1562 0.00334
R65798 DVSS.n5276 DVSS.n1562 0.00334
R65799 DVSS.n5277 DVSS.n5276 0.00334
R65800 DVSS.n5278 DVSS.n5277 0.00334
R65801 DVSS.n5278 DVSS.n1558 0.00334
R65802 DVSS.n5284 DVSS.n1558 0.00334
R65803 DVSS.n5285 DVSS.n5284 0.00334
R65804 DVSS.n5286 DVSS.n5285 0.00334
R65805 DVSS.n5286 DVSS.n1554 0.00334
R65806 DVSS.n5292 DVSS.n1554 0.00334
R65807 DVSS.n5293 DVSS.n5292 0.00334
R65808 DVSS.n5294 DVSS.n5293 0.00334
R65809 DVSS.n5294 DVSS.n1550 0.00334
R65810 DVSS.n5300 DVSS.n1550 0.00334
R65811 DVSS.n5301 DVSS.n5300 0.00334
R65812 DVSS.n5302 DVSS.n5301 0.00334
R65813 DVSS.n5303 DVSS.n5302 0.00334
R65814 DVSS.n5306 DVSS.n5303 0.00334
R65815 DVSS.n5307 DVSS.n5306 0.00334
R65816 DVSS.n5308 DVSS.n5307 0.00334
R65817 DVSS.n5309 DVSS.n5308 0.00334
R65818 DVSS.n5312 DVSS.n5309 0.00334
R65819 DVSS.n5313 DVSS.n5312 0.00334
R65820 DVSS.n5314 DVSS.n5313 0.00334
R65821 DVSS.n5315 DVSS.n5314 0.00334
R65822 DVSS.n5318 DVSS.n5315 0.00334
R65823 DVSS.n5319 DVSS.n5318 0.00334
R65824 DVSS.n5320 DVSS.n5319 0.00334
R65825 DVSS.n5321 DVSS.n5320 0.00334
R65826 DVSS.n595 DVSS.n594 0.00332
R65827 DVSS.n593 DVSS.n65 0.00332
R65828 DVSS.n592 DVSS.n397 0.00332
R65829 DVSS.n753 DVSS.n658 0.00332
R65830 DVSS.n657 DVSS.n586 0.00332
R65831 DVSS.n656 DVSS.n655 0.00332
R65832 DVSS.n5344 DVSS.n1527 0.00323
R65833 DVSS.n6397 DVSS.n273 0.00323
R65834 DVSS.n6501 DVSS.n6500 0.00323
R65835 DVSS.n1071 DVSS.n1029 0.00323
R65836 DVSS.n6073 DVSS.n6072 0.0032
R65837 DVSS.n368 DVSS.n367 0.0032
R65838 DVSS.n6392 DVSS.n257 0.0032
R65839 DVSS.n6076 DVSS.n1180 0.0032
R65840 DVSS.n377 DVSS.n357 0.0032
R65841 DVSS.n6383 DVSS.n192 0.0032
R65842 DVSS.n1170 DVSS.n1150 0.0032
R65843 DVSS.n370 DVSS.n96 0.0032
R65844 DVSS.n6385 DVSS.n133 0.0032
R65845 DVSS.n6085 DVSS.n1165 0.0032
R65846 DVSS.n371 DVSS.n53 0.0032
R65847 DVSS.n6386 DVSS.n239 0.0032
R65848 DVSS.n4449 DVSS.n4448 0.00311
R65849 DVSS.n6421 DVSS.n241 0.00311
R65850 DVSS.n6489 DVSS.n60 0.00311
R65851 DVSS.n6238 DVSS.n419 0.00311
R65852 DVSS.n955 DVSS.n922 0.00286
R65853 DVSS.n6511 DVSS.n11 0.00286
R65854 DVSS.n1068 DVSS.n1067 0.00286
R65855 DVSS.n4549 DVSS.n4506 0.00285923
R65856 DVSS.n4596 DVSS.n4506 0.00285923
R65857 DVSS.n6456 DVSS.n6454 0.00285923
R65858 DVSS.n6454 DVSS.n153 0.00285923
R65859 DVSS.n295 DVSS.n283 0.00285923
R65860 DVSS.n295 DVSS.n284 0.00285923
R65861 DVSS.n464 DVSS.n462 0.00285923
R65862 DVSS.n465 DVSS.n464 0.00285923
R65863 DVSS.n287 DVSS.n46 0.00285075
R65864 DVSS.n261 DVSS.n162 0.00285075
R65865 DVSS.n3093 DVSS.n2369 0.00284
R65866 DVSS.n3079 DVSS.n3078 0.00284
R65867 DVSS.n4366 DVSS.n4365 0.00277528
R65868 DVSS DVSS.n4876 0.00277528
R65869 DVSS.n992 DVSS.n891 0.0027
R65870 DVSS.n6346 DVSS.n339 0.0027
R65871 DVSS.n6167 DVSS.n6166 0.0027
R65872 DVSS.n5343 DVSS.n1525 0.00269
R65873 DVSS.n595 DVSS.n223 0.00269
R65874 DVSS.n6400 DVSS.n249 0.00269
R65875 DVSS.n6486 DVSS.n65 0.00269
R65876 DVSS.n30 DVSS.n15 0.00269
R65877 DVSS.n6241 DVSS.n397 0.00269
R65878 DVSS.n6132 DVSS.n6131 0.00269
R65879 DVSS.n4445 DVSS.n2056 0.00257
R65880 DVSS.n5340 DVSS.n1525 0.00257
R65881 DVSS.n224 DVSS.n223 0.00257
R65882 DVSS.n6400 DVSS.n258 0.00257
R65883 DVSS.n6486 DVSS.n50 0.00257
R65884 DVSS.n6507 DVSS.n15 0.00257
R65885 DVSS.n6241 DVSS.n405 0.00257
R65886 DVSS.n6131 DVSS.n1084 0.00257
R65887 DVSS.n3017 DVSS.n3012 0.00254225
R65888 DVSS.n2987 DVSS.n2525 0.00254225
R65889 DVSS.n838 DVSS.n557 0.00254
R65890 DVSS.n837 DVSS.n836 0.00254
R65891 DVSS.n713 DVSS.n564 0.00254
R65892 DVSS.n2905 DVSS 0.00247183
R65893 DVSS.n4851 DVSS.n1864 0.00239607
R65894 DVSS.n4848 DVSS.n1872 0.00239607
R65895 DVSS.n654 DVSS.n587 0.00238
R65896 DVSS.n757 DVSS.n756 0.00238
R65897 DVSS.n755 DVSS.n754 0.00238
R65898 DVSS.n3023 DVSS.n2433 0.00236429
R65899 DVSS.n2745 DVSS.n2744 0.00236429
R65900 DVSS.n3660 DVSS.n1798 0.00236429
R65901 DVSS.n3626 DVSS.n1752 0.00236429
R65902 DVSS.n3851 DVSS.n1801 0.00236429
R65903 DVSS.n3817 DVSS.n3726 0.00236429
R65904 DVSS.n4646 DVSS.n4645 0.00236429
R65905 DVSS.n4678 DVSS.n1994 0.00236429
R65906 DVSS.n6099 DVSS.n1152 0.00236429
R65907 DVSS.n5919 DVSS.n5775 0.00236429
R65908 DVSS.n2846 DVSS 0.0023
R65909 DVSS.n5056 DVSS 0.0023
R65910 DVSS.n5102 DVSS 0.0023
R65911 DVSS.n5523 DVSS 0.0023
R65912 DVSS.n5982 DVSS 0.0023
R65913 DVSS.n2252 VSS 0.0023
R65914 DVSS.n3302 VSS 0.0023
R65915 VSS DVSS.n3303 0.0023
R65916 VSS DVSS.n2253 0.0023
R65917 DVSS.n3506 DVSS.n2140 0.0023
R65918 DVSS.n2139 DVSS.n2137 0.0023
R65919 DVSS.n2981 DVSS.n2980 0.00226056
R65920 DVSS.n2952 DVSS.n2400 0.00226056
R65921 DVSS.n5446 DVSS 0.00218942
R65922 DVSS.n3529 DVSS.n2122 0.0021791
R65923 DVSS.n6222 DVSS.n456 0.0021791
R65924 DVSS.n6275 DVSS.n293 0.0021791
R65925 DVSS.n4245 DVSS 0.0021723
R65926 DVSS.n4448 DVSS.n2056 0.00215
R65927 DVSS.n6421 DVSS.n224 0.00215
R65928 DVSS.n6489 DVSS.n50 0.00215
R65929 DVSS.n6238 DVSS.n405 0.00215
R65930 DVSS.n2772 DVSS.n2647 0.00210714
R65931 DVSS.n3044 DVSS.n2404 0.00210714
R65932 DVSS.n3619 DVSS.n1740 0.00210714
R65933 DVSS.n5014 DVSS.n1713 0.00210714
R65934 DVSS.n3810 DVSS.n3788 0.00210714
R65935 DVSS.n5164 DVSS.n5163 0.00210714
R65936 DVSS.n4742 DVSS.n1980 0.00210714
R65937 DVSS.n5585 DVSS.n5584 0.00210714
R65938 DVSS.n6060 DVSS.n5781 0.00210714
R65939 DVSS.n6052 DVSS.n5804 0.00210714
R65940 DVSS.n5344 DVSS.n5343 0.00203
R65941 DVSS.n6397 DVSS.n249 0.00203
R65942 DVSS.n6500 DVSS.n30 0.00203
R65943 DVSS.n6132 DVSS.n1071 0.00203
R65944 DVSS.n4788 DVSS.n4787 0.00201685
R65945 DVSS.n3065 DVSS.n2397 0.00201119
R65946 DVSS.n6529 DVSS 0.00196
R65947 DVSS.n4995 DVSS.n1748 0.00184328
R65948 DVSS.n4994 DVSS.n1742 0.00184328
R65949 DVSS.n4991 DVSS.n4989 0.00184328
R65950 DVSS DVSS.n6533 0.00173
R65951 DVSS DVSS.n0 0.00173
R65952 DVSS DVSS.n5524 0.0017
R65953 DVSS.n842 DVSS.n841 0.0017
R65954 DVSS.n801 DVSS.n559 0.0017
R65955 DVSS.n717 DVSS.n716 0.0017
R65956 DVSS.n718 DVSS.n567 0.0017
R65957 DVSS.n803 DVSS.n802 0.0017
R65958 DVSS.n840 DVSS.n562 0.0017
R65959 DVSS.n5501 DVSS.n5500 0.00163764
R65960 DVSS.n6079 DVSS.n1176 0.00150746
R65961 DVSS.n369 DVSS.n289 0.00150746
R65962 DVSS.n6384 DVSS.n164 0.00150746
R65963 DVSS.n995 DVSS.n535 0.00146
R65964 DVSS.n996 DVSS.n341 0.00146
R65965 DVSS.n997 DVSS.n533 0.00146
R65966 DVSS.n6169 DVSS.n342 0.00146
R65967 DVSS.n6349 DVSS.n6348 0.00146
R65968 DVSS.n889 DVSS.n343 0.00146
R65969 DVSS.n1082 DVSS.n392 0.0014
R65970 DVSS.n6285 DVSS.n23 0.0014
R65971 DVSS.n6249 DVSS.n391 0.0014
R65972 DVSS.n6290 DVSS.n382 0.0014
R65973 DVSS.n6228 DVSS.n394 0.0014
R65974 DVSS.n6481 DVSS.n78 0.0014
R65975 DVSS.n6243 DVSS.n395 0.0014
R65976 DVSS.n6483 DVSS.n68 0.0014
R65977 DVSS.n4636 DVSS.n4625 0.00137
R65978 DVSS.n4600 DVSS.n4501 0.00137
R65979 DVSS.n6472 DVSS.n109 0.00137
R65980 DVSS.n6460 DVSS.n154 0.00137
R65981 DVSS.n6479 DVSS.n80 0.00137
R65982 DVSS.n6373 DVSS.n285 0.00137
R65983 DVSS.n6229 DVSS.n442 0.00137
R65984 DVSS.n6196 DVSS.n511 0.00137
R65985 DVSS DVSS.n5323 0.00134
R65986 DVSS.n1049 DVSS 0.00134
R65987 DVSS.n839 DVSS.n838 0.0013
R65988 DVSS.n837 DVSS.n565 0.0013
R65989 DVSS.n719 DVSS.n564 0.0013
R65990 DVSS.n3019 DVSS.n2435 0.00127465
R65991 DVSS.n2984 DVSS.n2983 0.00127465
R65992 DVSS.n4190 DVSS.n3886 0.00125843
R65993 DVSS.n4594 DVSS.n4593 0.00125
R65994 DVSS.n5272 DVSS.n1564 0.00125
R65995 DVSS.n869 DVSS.n152 0.00125
R65996 DVSS.n6439 DVSS.n193 0.00125
R65997 DVSS.n6371 DVSS.n6366 0.00125
R65998 DVSS.n6298 DVSS.n6297 0.00125
R65999 DVSS.n6199 DVSS.n475 0.00125
R66000 DVSS.n1006 DVSS.n389 0.00125
R66001 DVSS.n258 DVSS.n14 0.00122
R66002 DVSS.n6508 DVSS.n6507 0.00122
R66003 DVSS.n1084 DVSS.n13 0.00122
R66004 DVSS.n1070 DVSS.n1031 0.00122
R66005 DVSS.n6506 DVSS.n12 0.00122
R66006 DVSS.n958 DVSS.n957 0.00122
R66007 DVSS.n3026 DVSS.n2425 0.00120714
R66008 DVSS.n2766 DVSS.n2765 0.00120714
R66009 DVSS.n3657 DVSS.n1799 0.00120714
R66010 DVSS.n3577 DVSS.n1739 0.00120714
R66011 DVSS.n3848 DVSS.n1802 0.00120714
R66012 DVSS.n3807 DVSS.n3806 0.00120714
R66013 DVSS.n2016 DVSS.n2011 0.00120714
R66014 DVSS.n4740 DVSS.n4739 0.00120714
R66015 DVSS.n6102 DVSS.n1143 0.00120714
R66016 DVSS.n5824 DVSS.n5776 0.00120714
R66017 DVSS.n891 DVSS.n890 0.00114
R66018 DVSS.n6350 DVSS.n339 0.00114
R66019 DVSS.n6168 DVSS.n6167 0.00114
R66020 DVSS.n1967 DVSS.n1870 0.00113202
R66021 DVSS.n4849 DVSS.n1874 0.00113202
R66022 DVSS.n3327 DVSS.n3326 0.00107857
R66023 DVSS.n3328 DVSS.n2276 0.00107857
R66024 DVSS DVSS.n935 0.00102
R66025 DVSS.n2547 DVSS.n2546 0.000992958
R66026 DVSS.n2954 DVSS.n2399 0.000992958
R66027 DVSS.n922 DVSS.n919 0.00098
R66028 DVSS.n6505 DVSS.n11 0.00098
R66029 DVSS.n1069 DVSS.n1068 0.00098
R66030 DVSS.n2763 DVSS.n2761 0.00095
R66031 DVSS.n2402 DVSS.n2401 0.00095
R66032 DVSS.n4996 DVSS.n1743 0.00095
R66033 DVSS.n5007 DVSS.n1720 0.00095
R66034 DVSS.n3811 DVSS.n3730 0.00095
R66035 DVSS.n3756 DVSS.n1651 0.00095
R66036 DVSS.n1988 DVSS.n1974 0.00095
R66037 DVSS.n4703 DVSS.n1335 0.00095
R66038 DVSS.n5798 DVSS.n5777 0.00095
R66039 DVSS.n6049 DVSS.n5802 0.00095
R66040 DVSS.n467 DVSS.n393 0.000835821
R66041 DVSS.n6286 DVSS.n291 0.000835821
R66042 DVSS.n4639 DVSS.n2027 0.00083
R66043 DVSS.n4597 DVSS.n4596 0.00083
R66044 DVSS.n6470 DVSS.n117 0.00083
R66045 DVSS.n6456 DVSS.n166 0.00083
R66046 DVSS.n6476 DVSS.n88 0.00083
R66047 DVSS.n299 DVSS.n283 0.00083
R66048 DVSS.n6232 DVSS.n428 0.00083
R66049 DVSS.n6188 DVSS.n465 0.00083
R66050 DVSS.n2120 DVSS.n2117 0.000725
R66051 DVSS.n4550 DVSS.n4549 0.00071
R66052 DVSS.n5265 DVSS.n5264 0.00071
R66053 DVSS.n548 DVSS.n153 0.00071
R66054 DVSS.n207 DVSS.n183 0.00071
R66055 DVSS.n321 DVSS.n284 0.00071
R66056 DVSS.n6294 DVSS.n353 0.00071
R66057 DVSS.n466 DVSS.n462 0.00071
R66058 DVSS.n1005 DVSS.n390 0.00071
R66059 DVSS.n2904 DVSS 0.000687793
R66060 DVSS DVSS.n939 0.00068
R66061 DVSS.n2847 DVSS 0.000671429
R66062 DVSS.n5057 DVSS 0.000671429
R66063 DVSS.n5103 DVSS 0.000671429
R66064 DVSS.n5524 DVSS 0.000671429
R66065 DVSS.n5983 DVSS 0.000671429
R66066 VSS DVSS.n2241 0.000671429
R66067 VSS DVSS.n3278 0.000671429
R66068 DVSS DVSS.n1966 0.000626404
R66069 DVSS.n1050 DVSS 0.00058
R66070 DVSS DVSS.n5321 0.00058
R66071 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531459_0.D.n3 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531459_0.D.t4 47.1029
R66072 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531459_0.D.n1 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531459_0.D.t9 47.1029
R66073 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531459_0.D.n6 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531459_0.D.t7 47.1029
R66074 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531459_0.D.n6 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531459_0.D.t3 47.1029
R66075 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531459_0.D.n3 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531459_0.D.t11 38.0648
R66076 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531459_0.D.n4 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531459_0.D.t8 38.0648
R66077 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531459_0.D.n1 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531459_0.D.t10 38.0648
R66078 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531459_0.D.n2 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531459_0.D.t5 38.0648
R66079 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531459_0.D.n6 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531459_0.D.t6 38.0648
R66080 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531459_0.D.n4 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531459_0.D.n3 9.0386
R66081 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531459_0.D.n2 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531459_0.D.n1 9.0386
R66082 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531459_0.D.n5 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531459_0.D.n2 4.51955
R66083 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531459_0.D.n5 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531459_0.D.n4 4.51955
R66084 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531459_0.D.n0 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531459_0.D.t2 2.8466
R66085 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531459_0.D.n0 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531459_0.D.n5 2.40746
R66086 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531459_0.D.n0 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531459_0.D.t0 1.87633
R66087 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531459_0.D.n0 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531459_0.D.n6 1.76725
R66088 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531459_0.D.n0 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531459_0.D.t1 1.65385
R66089 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/comp018green_esd_rc_v5p0_0.ppolyf_u_CDNS_406619531453_1.MINUS.t0 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/comp018green_esd_rc_v5p0_0.ppolyf_u_CDNS_406619531453_1.MINUS.t1 22.3936
R66090 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/comp018green_esd_rc_v5p0_0.ppolyf_u_CDNS_406619531453_0.PLUS.t0 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/comp018green_esd_rc_v5p0_0.ppolyf_u_CDNS_406619531453_0.PLUS 11.0117
R66091 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/comp018green_esd_rc_v5p0_0.ppolyf_u_CDNS_406619531453_0.PLUS GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/comp018green_esd_rc_v5p0_0.ppolyf_u_CDNS_406619531453_0.PLUS.t1 11.0117
R66092 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/comp018green_esd_rc_v5p0_0.VRC GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/comp018green_esd_rc_v5p0_0.VRC.t0 11.0117
R66093 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/comp018green_esd_rc_v5p0_0.VRC GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/comp018green_esd_rc_v5p0_0.VRC.n12 0.6125
R66094 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/comp018green_esd_rc_v5p0_0.VRC.n12 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/comp018green_esd_rc_v5p0_0.VRC.n18 1.2266
R66095 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/comp018green_esd_rc_v5p0_0.VRC.n19 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/comp018green_esd_rc_v5p0_0.VRC 0.225727
R66096 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/comp018green_esd_rc_v5p0_0.VRC GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/comp018green_esd_rc_v5p0_0.VRC.n18 0.00644
R66097 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/comp018green_esd_rc_v5p0_0.VRC.t9 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/comp018green_esd_rc_v5p0_0.VRC.n19 4.75334
R66098 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/comp018green_esd_rc_v5p0_0.VRC GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/comp018green_esd_rc_v5p0_0.VRC.n19 0.225727
R66099 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/comp018green_esd_rc_v5p0_0.VRC.n18 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/comp018green_esd_rc_v5p0_0.VRC.n16 0.767246
R66100 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/comp018green_esd_rc_v5p0_0.VRC.n17 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/comp018green_esd_rc_v5p0_0.VRC 0.225727
R66101 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/comp018green_esd_rc_v5p0_0.VRC GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/comp018green_esd_rc_v5p0_0.VRC.n16 0.00644
R66102 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/comp018green_esd_rc_v5p0_0.VRC.t8 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/comp018green_esd_rc_v5p0_0.VRC.n17 4.75334
R66103 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/comp018green_esd_rc_v5p0_0.VRC GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/comp018green_esd_rc_v5p0_0.VRC.n17 0.225727
R66104 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/comp018green_esd_rc_v5p0_0.VRC.n16 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/comp018green_esd_rc_v5p0_0.VRC.n14 0.767246
R66105 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/comp018green_esd_rc_v5p0_0.VRC.n15 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/comp018green_esd_rc_v5p0_0.VRC 0.225727
R66106 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/comp018green_esd_rc_v5p0_0.VRC GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/comp018green_esd_rc_v5p0_0.VRC.n14 0.00644
R66107 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/comp018green_esd_rc_v5p0_0.VRC.t11 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/comp018green_esd_rc_v5p0_0.VRC.n15 4.75334
R66108 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/comp018green_esd_rc_v5p0_0.VRC GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/comp018green_esd_rc_v5p0_0.VRC.n15 0.225727
R66109 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/comp018green_esd_rc_v5p0_0.VRC.n13 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/comp018green_esd_rc_v5p0_0.VRC 0.225727
R66110 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/comp018green_esd_rc_v5p0_0.VRC GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/comp018green_esd_rc_v5p0_0.VRC.n14 0.773185
R66111 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/comp018green_esd_rc_v5p0_0.VRC.t10 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/comp018green_esd_rc_v5p0_0.VRC.n13 4.75334
R66112 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/comp018green_esd_rc_v5p0_0.VRC GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/comp018green_esd_rc_v5p0_0.VRC.n13 0.225727
R66113 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/comp018green_esd_rc_v5p0_0.VRC.n12 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/comp018green_esd_rc_v5p0_0.VRC.n4 6.26225
R66114 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/comp018green_esd_rc_v5p0_0.VRC.n4 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/comp018green_esd_rc_v5p0_0.VRC 0.332722
R66115 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/comp018green_esd_rc_v5p0_0.VRC GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/comp018green_esd_rc_v5p0_0.VRC.n10 0.894378
R66116 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/comp018green_esd_rc_v5p0_0.VRC.n10 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/comp018green_esd_rc_v5p0_0.VRC 0.00644
R66117 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/comp018green_esd_rc_v5p0_0.VRC.n11 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/comp018green_esd_rc_v5p0_0.VRC 0.225727
R66118 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/comp018green_esd_rc_v5p0_0.VRC.t5 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/comp018green_esd_rc_v5p0_0.VRC.n11 4.75334
R66119 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/comp018green_esd_rc_v5p0_0.VRC GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/comp018green_esd_rc_v5p0_0.VRC.n11 0.225727
R66120 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/comp018green_esd_rc_v5p0_0.VRC.n10 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/comp018green_esd_rc_v5p0_0.VRC.n8 0.767246
R66121 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/comp018green_esd_rc_v5p0_0.VRC.n8 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/comp018green_esd_rc_v5p0_0.VRC 0.00644
R66122 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/comp018green_esd_rc_v5p0_0.VRC.n9 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/comp018green_esd_rc_v5p0_0.VRC 0.225727
R66123 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/comp018green_esd_rc_v5p0_0.VRC.t4 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/comp018green_esd_rc_v5p0_0.VRC.n9 4.75334
R66124 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/comp018green_esd_rc_v5p0_0.VRC GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/comp018green_esd_rc_v5p0_0.VRC.n9 0.225727
R66125 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/comp018green_esd_rc_v5p0_0.VRC.n8 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/comp018green_esd_rc_v5p0_0.VRC.n6 0.767246
R66126 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/comp018green_esd_rc_v5p0_0.VRC.n6 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/comp018green_esd_rc_v5p0_0.VRC 0.00644
R66127 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/comp018green_esd_rc_v5p0_0.VRC.n7 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/comp018green_esd_rc_v5p0_0.VRC 0.225727
R66128 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/comp018green_esd_rc_v5p0_0.VRC.t7 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/comp018green_esd_rc_v5p0_0.VRC.n7 4.75334
R66129 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/comp018green_esd_rc_v5p0_0.VRC GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/comp018green_esd_rc_v5p0_0.VRC.n7 0.225727
R66130 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/comp018green_esd_rc_v5p0_0.VRC.n6 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/comp018green_esd_rc_v5p0_0.VRC 0.773185
R66131 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/comp018green_esd_rc_v5p0_0.VRC.n5 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/comp018green_esd_rc_v5p0_0.VRC 0.225727
R66132 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/comp018green_esd_rc_v5p0_0.VRC.t6 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/comp018green_esd_rc_v5p0_0.VRC.n5 4.75334
R66133 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/comp018green_esd_rc_v5p0_0.VRC GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/comp018green_esd_rc_v5p0_0.VRC.n5 0.225727
R66134 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/comp018green_esd_rc_v5p0_0.VRC.n3 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/comp018green_esd_rc_v5p0_0.VRC.n2 1.0005
R66135 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/comp018green_esd_rc_v5p0_0.VRC.n4 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/comp018green_esd_rc_v5p0_0.VRC.n3 2.62726
R66136 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/comp018green_esd_rc_v5p0_0.VRC.n3 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/comp018green_esd_rc_v5p0_0.VRC.t3 36.8287
R66137 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/comp018green_esd_rc_v5p0_0.VRC.n2 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/comp018green_esd_rc_v5p0_0.VRC.n0 4.51955
R66138 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/comp018green_esd_rc_v5p0_0.VRC.n2 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/comp018green_esd_rc_v5p0_0.VRC.n1 4.51955
R66139 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/comp018green_esd_rc_v5p0_0.VRC.n1 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/comp018green_esd_rc_v5p0_0.VRC.t2 38.0648
R66140 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/comp018green_esd_rc_v5p0_0.VRC.n1 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/comp018green_esd_rc_v5p0_0.VRC.t1 47.1029
R66141 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/comp018green_esd_rc_v5p0_0.VRC.n0 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/comp018green_esd_rc_v5p0_0.VRC.t12 38.0648
R66142 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/comp018green_esd_rc_v5p0_0.VRC.n0 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/comp018green_esd_rc_v5p0_0.VRC.t13 47.1029
R66143 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/comp018green_esd_rc_v5p0_0.ppolyf_u_CDNS_406619531453_5.MINUS GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/comp018green_esd_rc_v5p0_0.ppolyf_u_CDNS_406619531453_5.MINUS.t0 11.0117
R66144 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/comp018green_esd_rc_v5p0_0.ppolyf_u_CDNS_406619531453_5.MINUS GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/comp018green_esd_rc_v5p0_0.ppolyf_u_CDNS_406619531453_5.MINUS.t1 11.0117
R66145 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/comp018green_esd_rc_v5p0_0.ppolyf_u_CDNS_406619531453_3.PLUS.t0 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/comp018green_esd_rc_v5p0_0.ppolyf_u_CDNS_406619531453_3.PLUS.t1 22.3936
R66146 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/comp018green_esd_rc_v5p0_0.ppolyf_u_CDNS_406619531453_2.MINUS.t0 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/comp018green_esd_rc_v5p0_0.ppolyf_u_CDNS_406619531453_2.MINUS.t1 22.3936
R66147 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/comp018green_esd_rc_v5p0_0.ppolyf_u_CDNS_406619531453_4.PLUS.t0 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/comp018green_esd_rc_v5p0_0.ppolyf_u_CDNS_406619531453_4.PLUS.t1 22.3936
R66148 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/comp018green_esd_rc_v5p0_0.ppolyf_u_CDNS_406619531453_3.MINUS.t0 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/comp018green_esd_rc_v5p0_0.ppolyf_u_CDNS_406619531453_3.MINUS.t1 22.3936
R66149 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/comp018green_esd_rc_v5p0_0.ppolyf_u_CDNS_406619531453_4.MINUS GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/comp018green_esd_rc_v5p0_0.ppolyf_u_CDNS_406619531453_4.MINUS.t0 11.0117
R66150 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/comp018green_esd_rc_v5p0_0.ppolyf_u_CDNS_406619531453_4.MINUS GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/comp018green_esd_rc_v5p0_0.ppolyf_u_CDNS_406619531453_4.MINUS.t1 11.0117
R66151 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/comp018green_esd_rc_v5p0_0.ppolyf_u_CDNS_406619531453_5.PLUS.t0 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/comp018green_esd_rc_v5p0_0.ppolyf_u_CDNS_406619531453_5.PLUS.t1 22.3936
R66152 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/comp018green_esd_rc_v5p0_0.ppolyf_u_CDNS_406619531453_2.PLUS.t0 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/comp018green_esd_rc_v5p0_0.ppolyf_u_CDNS_406619531453_2.PLUS 11.0117
R66153 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/comp018green_esd_rc_v5p0_0.ppolyf_u_CDNS_406619531453_2.PLUS GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/comp018green_esd_rc_v5p0_0.ppolyf_u_CDNS_406619531453_2.PLUS.t1 11.0117
R66154 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/comp018green_esd_rc_v5p0_0.ppolyf_u_CDNS_406619531453_1.PLUS.t0 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/comp018green_esd_rc_v5p0_0.ppolyf_u_CDNS_406619531453_1.PLUS 11.0117
R66155 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/comp018green_esd_rc_v5p0_0.ppolyf_u_CDNS_406619531453_1.PLUS GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/comp018green_esd_rc_v5p0_0.ppolyf_u_CDNS_406619531453_1.PLUS.t1 11.0117
R66156 VSS.n6455 VSS.n6454 82387.9
R66157 VSS.n6220 VSS.n6219 69392.3
R66158 VSS.n6219 VSS.n6218 69376.4
R66159 VSS.n6455 VSS.n10 20752.5
R66160 VSS.n6454 VSS.n6453 20730.8
R66161 VSS.n6221 VSS.n6220 16226.6
R66162 VSS.n6218 VSS.n6197 16226.6
R66163 VSS.n1610 VSS.n9 4180.28
R66164 VSS.n1609 VSS.n1608 4158.32
R66165 VSS.n6456 VSS.n6455 3610.1
R66166 VSS.n6454 VSS.n11 3610.1
R66167 VSS.n2912 VSS.n1127 3372.16
R66168 VSS.n2958 VSS.n1127 3372.16
R66169 VSS.n6456 VSS.n9 3351.4
R66170 VSS.n1608 VSS.n11 3351.4
R66171 VSS.n4120 VSS.n450 3055
R66172 VSS.n4119 VSS.n568 2710.64
R66173 VSS.n6223 VSS.n448 2402.48
R66174 VSS.n6223 VSS.n449 2401.2
R66175 VSS.n6201 VSS.n448 2400.01
R66176 VSS.n6201 VSS.n449 2398.73
R66177 VSS.n6196 VSS.n451 1820
R66178 VSS.n555 VSS.n476 1625.57
R66179 VSS.n5828 VSS.n478 1625.57
R66180 VSS.n6153 VSS.n476 1596.72
R66181 VSS.n6153 VSS.n478 1596.72
R66182 VSS.n6222 VSS.n6221 1409.58
R66183 VSS.n6200 VSS.n6197 1409.58
R66184 VSS.n567 VSS.n563 1373.3
R66185 VSS.n6222 VSS.n10 1327.85
R66186 VSS.n6200 VSS.n12 1327.85
R66187 VSS.n563 VSS.n451 1096.7
R66188 VSS.n4120 VSS.n4119 864.362
R66189 VSS.n568 VSS.n567 650
R66190 VSS.n1608 VSS.n1607 551.231
R66191 VSS.n1883 VSS.n9 551.231
R66192 VSS.n4118 VSS.n562 290.034
R66193 VSS.n4118 VSS.n452 266.233
R66194 VSS.n6195 VSS.n452 233.644
R66195 VSS.n4121 VSS.n562 227.811
R66196 VSS.n4121 VSS.n561 201.056
R66197 VSS.n3391 VSS.n10 177.477
R66198 VSS.n2545 VSS.n12 177.222
R66199 VSS.n6197 VSS.n6196 177.022
R66200 VSS.n6221 VSS.n450 177.022
R66201 VSS.n6195 VSS.n453 158.357
R66202 VSS.n566 VSS.n453 138.911
R66203 VSS.n2959 VSS.n1126 130.275
R66204 VSS.n2913 VSS.n1126 130.275
R66205 VSS.n2911 VSS.n2881 130.275
R66206 VSS.n2881 VSS.n1128 130.275
R66207 VSS.n2912 VSS.n2877 123.9
R66208 VSS.n2958 VSS.n1129 123.9
R66209 VSS.n2876 VSS.n2875 75.1538
R66210 VSS.n2875 VSS.n1124 75.1538
R66211 VSS.n2893 VSS.n2892 75.1538
R66212 VSS.n2893 VSS.n1132 75.1538
R66213 VSS.n2905 VSS.n2904 75.1538
R66214 VSS.n2904 VSS.n1131 75.1538
R66215 VSS.n2543 VSS.n2073 39.3263
R66216 VSS.n3397 VSS.n3101 39.3263
R66217 VSS.n566 VSS.n561 36.5561
R66218 VSS.n2681 VSS.n2073 29.1118
R66219 VSS.n2681 VSS.n2074 29.1118
R66220 VSS.n2675 VSS.n2074 29.1118
R66221 VSS.n2675 VSS.n2220 29.1118
R66222 VSS.n2669 VSS.n2220 29.1118
R66223 VSS.n2669 VSS.n2557 29.1118
R66224 VSS.n2663 VSS.n2557 29.1118
R66225 VSS.n2663 VSS.n2562 29.1118
R66226 VSS.n2657 VSS.n2562 29.1118
R66227 VSS.n2657 VSS.n2567 29.1118
R66228 VSS.n2651 VSS.n2567 29.1118
R66229 VSS.n2651 VSS.n2572 29.1118
R66230 VSS.n2645 VSS.n2572 29.1118
R66231 VSS.n2645 VSS.n2577 29.1118
R66232 VSS.n2639 VSS.n2577 29.1118
R66233 VSS.n2639 VSS.n2582 29.1118
R66234 VSS.n2633 VSS.n2582 29.1118
R66235 VSS.n2633 VSS.n2587 29.1118
R66236 VSS.n2627 VSS.n2587 29.1118
R66237 VSS.n2627 VSS.n2592 29.1118
R66238 VSS.n2592 VSS.n669 29.1118
R66239 VSS.n3927 VSS.n669 29.1118
R66240 VSS.n3927 VSS.n670 29.1118
R66241 VSS.n3920 VSS.n670 29.1118
R66242 VSS.n3920 VSS.n677 29.1118
R66243 VSS.n3914 VSS.n677 29.1118
R66244 VSS.n3914 VSS.n682 29.1118
R66245 VSS.n3908 VSS.n682 29.1118
R66246 VSS.n3908 VSS.n687 29.1118
R66247 VSS.n3902 VSS.n687 29.1118
R66248 VSS.n3902 VSS.n692 29.1118
R66249 VSS.n3896 VSS.n692 29.1118
R66250 VSS.n3896 VSS.n696 29.1118
R66251 VSS.n3890 VSS.n696 29.1118
R66252 VSS.n3890 VSS.n701 29.1118
R66253 VSS.n3884 VSS.n701 29.1118
R66254 VSS.n3884 VSS.n707 29.1118
R66255 VSS.n3878 VSS.n707 29.1118
R66256 VSS.n3878 VSS.n712 29.1118
R66257 VSS.n3872 VSS.n712 29.1118
R66258 VSS.n3872 VSS.n717 29.1118
R66259 VSS.n3866 VSS.n717 29.1118
R66260 VSS.n3866 VSS.n722 29.1118
R66261 VSS.n741 VSS.n722 29.1118
R66262 VSS.n3856 VSS.n741 29.1118
R66263 VSS.n3856 VSS.n742 29.1118
R66264 VSS.n3850 VSS.n742 29.1118
R66265 VSS.n3850 VSS.n749 29.1118
R66266 VSS.n3844 VSS.n749 29.1118
R66267 VSS.n3844 VSS.n755 29.1118
R66268 VSS.n3838 VSS.n755 29.1118
R66269 VSS.n3838 VSS.n760 29.1118
R66270 VSS.n3832 VSS.n760 29.1118
R66271 VSS.n3832 VSS.n765 29.1118
R66272 VSS.n3826 VSS.n765 29.1118
R66273 VSS.n3826 VSS.n770 29.1118
R66274 VSS.n3820 VSS.n770 29.1118
R66275 VSS.n3820 VSS.n775 29.1118
R66276 VSS.n3814 VSS.n775 29.1118
R66277 VSS.n3814 VSS.n780 29.1118
R66278 VSS.n3808 VSS.n780 29.1118
R66279 VSS.n3808 VSS.n785 29.1118
R66280 VSS.n3802 VSS.n785 29.1118
R66281 VSS.n3802 VSS.n790 29.1118
R66282 VSS.n3795 VSS.n790 29.1118
R66283 VSS.n3795 VSS.n795 29.1118
R66284 VSS.n3788 VSS.n795 29.1118
R66285 VSS.n3788 VSS.n800 29.1118
R66286 VSS.n3782 VSS.n800 29.1118
R66287 VSS.n3782 VSS.n806 29.1118
R66288 VSS.n3776 VSS.n806 29.1118
R66289 VSS.n3776 VSS.n811 29.1118
R66290 VSS.n3770 VSS.n811 29.1118
R66291 VSS.n3770 VSS.n816 29.1118
R66292 VSS.n3764 VSS.n816 29.1118
R66293 VSS.n3764 VSS.n821 29.1118
R66294 VSS.n3758 VSS.n821 29.1118
R66295 VSS.n3758 VSS.n826 29.1118
R66296 VSS.n3752 VSS.n826 29.1118
R66297 VSS.n3752 VSS.n831 29.1118
R66298 VSS.n3746 VSS.n831 29.1118
R66299 VSS.n3746 VSS.n836 29.1118
R66300 VSS.n3740 VSS.n836 29.1118
R66301 VSS.n3740 VSS.n841 29.1118
R66302 VSS.n3734 VSS.n841 29.1118
R66303 VSS.n3734 VSS.n846 29.1118
R66304 VSS.n3397 VSS.n846 29.1118
R66305 VSS.n3391 VSS.n3101 29.1118
R66306 VSS.n6453 VSS.n12 21.9617
R66307 VSS.n1610 VSS.n1609 21.96
R66308 VSS.n6271 VSS.n109 17.2463
R66309 VSS.n447 VSS.n446 7.85992
R66310 VSS.n447 VSS.n443 7.82456
R66311 VSS.n2959 VSS.n1124 7.68902
R66312 VSS.n2892 VSS.n2879 7.68902
R66313 VSS.n2879 VSS.n2876 7.68902
R66314 VSS.n2913 VSS.n2876 7.68902
R66315 VSS.n2957 VSS.n1131 7.68902
R66316 VSS.n2957 VSS.n1132 7.68902
R66317 VSS.n1132 VSS.n1130 7.68902
R66318 VSS.n1130 VSS.n1124 7.68902
R66319 VSS.n2911 VSS.n2905 7.68902
R66320 VSS.n2905 VSS.n2878 7.68902
R66321 VSS.n2892 VSS.n2878 7.68902
R66322 VSS.n1131 VSS.n1128 7.68902
R66323 VSS.n6198 VSS.n124 6.84065
R66324 VSS.n6217 VSS.n6198 6.80529
R66325 VSS.n3396 VSS.n3395 5.28481
R66326 VSS.n3268 VSS.n3102 5.28481
R66327 VSS.n3398 VSS.n3100 5.28481
R66328 VSS.n2542 VSS.n2541 5.2005
R66329 VSS.n2543 VSS.n2542 5.2005
R66330 VSS.n2542 VSS.n2444 5.2005
R66331 VSS.n2541 VSS.n2540 5.2005
R66332 VSS.n2540 VSS.n2444 5.2005
R66333 VSS.n2546 VSS.n2231 5.2005
R66334 VSS.n2546 VSS.n2545 5.2005
R66335 VSS.n2231 VSS.n2229 5.2005
R66336 VSS.n2545 VSS.n2229 5.2005
R66337 VSS.n2259 VSS.n2231 5.2005
R66338 VSS.n2545 VSS.n2259 5.2005
R66339 VSS.n2286 VSS.n2231 5.2005
R66340 VSS.n2545 VSS.n2286 5.2005
R66341 VSS.n2258 VSS.n2231 5.2005
R66342 VSS.n2545 VSS.n2258 5.2005
R66343 VSS.n2287 VSS.n2231 5.2005
R66344 VSS.n2545 VSS.n2287 5.2005
R66345 VSS.n2313 VSS.n2232 5.2005
R66346 VSS.n2545 VSS.n2232 5.2005
R66347 VSS.n2313 VSS.n2288 5.2005
R66348 VSS.n3130 VSS.n3101 5.2005
R66349 VSS.n3157 VSS.n3101 5.2005
R66350 VSS.n3158 VSS.n3101 5.2005
R66351 VSS.n3279 VSS.n3270 5.2005
R66352 VSS.n3270 VSS.n3101 5.2005
R66353 VSS.n3279 VSS.n3269 5.2005
R66354 VSS.n3269 VSS.n3101 5.2005
R66355 VSS.n3272 VSS.n3101 5.2005
R66356 VSS.n3276 VSS.n3133 5.2005
R66357 VSS.n3391 VSS.n3133 5.2005
R66358 VSS.n3279 VSS.n3268 5.2005
R66359 VSS.n3268 VSS.n3101 5.2005
R66360 VSS.n3276 VSS.n3274 5.2005
R66361 VSS.n3279 VSS.n3274 5.2005
R66362 VSS.n3274 VSS.n3101 5.2005
R66363 VSS.n3279 VSS.n3267 5.2005
R66364 VSS.n3267 VSS.n3101 5.2005
R66365 VSS.n3279 VSS.n3278 5.2005
R66366 VSS.n3278 VSS.n3101 5.2005
R66367 VSS.n3104 VSS.n3101 5.2005
R66368 VSS.n5807 VSS.n5051 5.02526
R66369 VSS.n5108 VSS.n5106 5.02526
R66370 VSS.n5097 VSS.n5095 5.02526
R66371 VSS.n5791 VSS.n5078 5.02526
R66372 VSS.n5850 VSS.n5848 5.02526
R66373 VSS.n5467 VSS.n4964 5.02526
R66374 VSS.n5638 VSS.n5255 5.02526
R66375 VSS.n5523 VSS.n5521 5.02526
R66376 VSS.n5516 VSS.n5514 5.02526
R66377 VSS.n5534 VSS.n5532 5.02526
R66378 VSS.n5989 VSS.n5987 5.02526
R66379 VSS.n4820 VSS.n4819 5.02526
R66380 VSS.n4832 VSS.n4831 5.02526
R66381 VSS.n4844 VSS.n4843 5.02526
R66382 VSS.n4856 VSS.n4855 5.02526
R66383 VSS.n4795 VSS.n4794 5.02526
R66384 VSS.n4788 VSS.n4482 5.02526
R66385 VSS.n4785 VSS.n4782 5.02526
R66386 VSS.n4781 VSS.n4780 5.02526
R66387 VSS.n4771 VSS.n4513 5.02526
R66388 VSS.n6136 VSS.n6135 5.02526
R66389 VSS.n4238 VSS.n503 5.02526
R66390 VSS.n4241 VSS.n512 5.02526
R66391 VSS.n4235 VSS.n514 5.02526
R66392 VSS.n522 VSS.n521 5.02526
R66393 VSS.n4222 VSS.n523 5.02526
R66394 VSS.n4219 VSS.n525 5.02526
R66395 VSS.n533 VSS.n532 5.02526
R66396 VSS.n4206 VSS.n534 5.02526
R66397 VSS.n4203 VSS.n4198 5.02526
R66398 VSS.n4194 VSS.n4193 5.02526
R66399 VSS.n4174 VSS.n539 5.02526
R66400 VSS.n4171 VSS.n4168 5.02526
R66401 VSS.n4167 VSS.n4166 5.02526
R66402 VSS.n4160 VSS.n544 5.02526
R66403 VSS.n4157 VSS.n4154 5.02526
R66404 VSS.n4153 VSS.n4152 5.02526
R66405 VSS.n4146 VSS.n548 5.02526
R66406 VSS.n4143 VSS.n4140 5.02526
R66407 VSS.n4139 VSS.n4138 5.02526
R66408 VSS.n6161 VSS.n459 5.02426
R66409 VSS.n6162 VSS.n460 5.02426
R66410 VSS.n6163 VSS.n461 5.02426
R66411 VSS.n6164 VSS.n462 5.02426
R66412 VSS.n6165 VSS.n463 5.02426
R66413 VSS.n6166 VSS.n464 5.02426
R66414 VSS.n6167 VSS.n465 5.02426
R66415 VSS.n6168 VSS.n466 5.02426
R66416 VSS.n6169 VSS.n467 5.02426
R66417 VSS.n6170 VSS.n468 5.02426
R66418 VSS.n4200 VSS.n4199 5.02426
R66419 VSS.n4210 VSS.n526 5.02426
R66420 VSS.n4214 VSS.n4213 5.02426
R66421 VSS.n4216 VSS.n4215 5.02426
R66422 VSS.n4226 VSS.n515 5.02426
R66423 VSS.n4230 VSS.n4229 5.02426
R66424 VSS.n4232 VSS.n4231 5.02426
R66425 VSS.n4245 VSS.n507 5.02426
R66426 VSS.n4249 VSS.n4248 5.02426
R66427 VSS.n6132 VSS.n6131 5.02426
R66428 VSS.n4511 VSS.n4510 5.02426
R66429 VSS.n6090 VSS.n4275 5.02426
R66430 VSS.n6091 VSS.n4276 5.02426
R66431 VSS.n6092 VSS.n4277 5.02426
R66432 VSS.n6093 VSS.n4278 5.02426
R66433 VSS.n4852 VSS.n4851 5.02426
R66434 VSS.n4840 VSS.n4839 5.02426
R66435 VSS.n4828 VSS.n4827 5.02426
R66436 VSS.n4816 VSS.n4815 5.02426
R66437 VSS.n6101 VSS.n6100 5.02426
R66438 VSS.n5530 VSS.n5529 5.02426
R66439 VSS.n5512 VSS.n5511 5.02426
R66440 VSS.n5626 VSS.n5625 5.02426
R66441 VSS.n5635 VSS.n5634 5.02426
R66442 VSS.n5465 VSS.n5273 5.02426
R66443 VSS.n5845 VSS.n5844 5.02426
R66444 VSS.n5788 VSS.n5787 5.02426
R66445 VSS.n5102 VSS.n5101 5.02426
R66446 VSS.n5113 VSS.n5112 5.02426
R66447 VSS.n5117 VSS.n5116 5.02426
R66448 VSS.n6448 VSS.n6447 4.83569
R66449 VSS.n6457 VSS.n8 4.72792
R66450 VSS.n6226 VSS.n8 4.60071
R66451 VSS.n136 VSS.n135 4.60071
R66452 VSS.n1886 VSS.n1229 4.5005
R66453 VSS.n1884 VSS.n1229 4.5005
R66454 VSS.n1886 VSS.n1885 4.5005
R66455 VSS.n1885 VSS.n1884 4.5005
R66456 VSS.n4859 VSS.n4808 4.5005
R66457 VSS.n4859 VSS.n4821 4.5005
R66458 VSS.n4859 VSS.n4806 4.5005
R66459 VSS.n4859 VSS.n4833 4.5005
R66460 VSS.n4859 VSS.n4804 4.5005
R66461 VSS.n4859 VSS.n4845 4.5005
R66462 VSS.n4859 VSS.n4802 4.5005
R66463 VSS.n4859 VSS.n4857 4.5005
R66464 VSS.n5985 VSS.n4796 4.5005
R66465 VSS.n6139 VSS.n500 4.5005
R66466 VSS.n6139 VSS.n497 4.5005
R66467 VSS.n6139 VSS.n502 4.5005
R66468 VSS.n6139 VSS.n492 4.5005
R66469 VSS.n6140 VSS.n489 4.5005
R66470 VSS.n6140 VSS.n6139 4.5005
R66471 VSS.n6139 VSS.n488 4.5005
R66472 VSS.n6139 VSS.n6138 4.5005
R66473 VSS.n4090 VSS.n4089 4.5005
R66474 VSS.n3728 VSS.n585 4.5005
R66475 VSS.n3727 VSS.n3726 4.5005
R66476 VSS.n3726 VSS.n3725 4.5005
R66477 VSS.n3403 VSS.n3402 4.5005
R66478 VSS.n3067 VSS.n3066 4.5005
R66479 VSS.n3065 VSS.n3064 4.5005
R66480 VSS.n1828 VSS.n1060 4.5005
R66481 VSS.n1830 VSS.n1829 4.5005
R66482 VSS.n1833 VSS.n1232 4.5005
R66483 VSS.n1833 VSS.n1231 4.5005
R66484 VSS.n1833 VSS.n1255 4.5005
R66485 VSS.n1833 VSS.n1251 4.5005
R66486 VSS.n1834 VSS.n1833 4.5005
R66487 VSS.n1836 VSS.n1835 4.5005
R66488 VSS.n1880 VSS.n1879 4.5005
R66489 VSS.n1836 VSS.n1234 4.5005
R66490 VSS.n1879 VSS.n1234 4.5005
R66491 VSS.n1830 VSS.n1255 4.5005
R66492 VSS.n1830 VSS.n1231 4.5005
R66493 VSS.n5986 VSS.n5985 4.5005
R66494 VSS.n5858 VSS.n4859 4.5005
R66495 VSS.n5856 VSS.n5855 4.5005
R66496 VSS.n5852 VSS.n4972 4.5005
R66497 VSS.n5855 VSS.n4959 4.5005
R66498 VSS.n5855 VSS.n4954 4.5005
R66499 VSS.n5855 VSS.n4960 4.5005
R66500 VSS.n5855 VSS.n4952 4.5005
R66501 VSS.n5855 VSS.n4961 4.5005
R66502 VSS.n5852 VSS.n4975 4.5005
R66503 VSS.n5852 VSS.n4966 4.5005
R66504 VSS.n5852 VSS.n4976 4.5005
R66505 VSS.n5853 VSS.n5852 4.5005
R66506 VSS.n5852 VSS.n5851 4.5005
R66507 VSS.n5849 VSS.n4943 4.5005
R66508 VSS.n5077 VSS.n4943 4.5005
R66509 VSS.n5868 VSS.n4927 4.5005
R66510 VSS.n5868 VSS.n4929 4.5005
R66511 VSS.n5868 VSS.n4925 4.5005
R66512 VSS.n5868 VSS.n4930 4.5005
R66513 VSS.n5868 VSS.n4923 4.5005
R66514 VSS.n5868 VSS.n4931 4.5005
R66515 VSS.n5868 VSS.n4921 4.5005
R66516 VSS.n5868 VSS.n4932 4.5005
R66517 VSS.n4943 VSS.n4918 4.5005
R66518 VSS.n5868 VSS.n4918 4.5005
R66519 VSS.n4943 VSS.n4933 4.5005
R66520 VSS.n5868 VSS.n4933 4.5005
R66521 VSS.n4859 VSS.n4472 4.5005
R66522 VSS.n2943 VSS.n1138 4.5005
R66523 VSS.n1140 VSS.n1138 4.5005
R66524 VSS.n2964 VSS.n1120 4.5005
R66525 VSS.n2962 VSS.n1120 4.5005
R66526 VSS.n2954 VSS.n2950 4.5005
R66527 VSS.n2946 VSS.n1137 4.5005
R66528 VSS.n2949 VSS.n2948 4.5005
R66529 VSS.n2951 VSS.n1134 4.5005
R66530 VSS.n2963 VSS.n2962 4.5005
R66531 VSS.n2964 VSS.n2963 4.5005
R66532 VSS.n2984 VSS.n1094 4.5005
R66533 VSS.n2984 VSS.n2983 4.5005
R66534 VSS.n1890 VSS.n1225 4.5005
R66535 VSS.n1888 VSS.n1225 4.5005
R66536 VSS.n1890 VSS.n1889 4.5005
R66537 VSS.n1889 VSS.n1888 4.5005
R66538 VSS.n4811 VSS.n4449 4.5005
R66539 VSS.n4823 VSS.n4449 4.5005
R66540 VSS.n4835 VSS.n4449 4.5005
R66541 VSS.n4847 VSS.n4449 4.5005
R66542 VSS.n5996 VSS.n4470 4.5005
R66543 VSS.n4768 VSS.n4519 4.5005
R66544 VSS.n4769 VSS.n4768 4.5005
R66545 VSS.n4765 VSS.n4764 4.5005
R66546 VSS.n4765 VSS.n486 4.5005
R66547 VSS.n4768 VSS.n486 4.5005
R66548 VSS.n4768 VSS.n485 4.5005
R66549 VSS.n4768 VSS.n4767 4.5005
R66550 VSS.n4104 VSS.n572 4.5005
R66551 VSS.n4115 VSS.n571 4.5005
R66552 VSS.n3640 VSS.n882 4.5005
R66553 VSS.n3640 VSS.n3639 4.5005
R66554 VSS.n3437 VSS.n3436 4.5005
R66555 VSS.n2779 VSS.n2778 4.5005
R66556 VSS.n2777 VSS.n1077 4.5005
R66557 VSS.n1095 VSS.n1077 4.5005
R66558 VSS.n2985 VSS.n1077 4.5005
R66559 VSS.n2986 VSS.n1091 4.5005
R66560 VSS.n2986 VSS.n1083 4.5005
R66561 VSS.n1083 VSS.n1077 4.5005
R66562 VSS.n2986 VSS.n1092 4.5005
R66563 VSS.n1092 VSS.n1077 4.5005
R66564 VSS.n1754 VSS.n1278 4.5005
R66565 VSS.n1751 VSS.n1228 4.5005
R66566 VSS.n1754 VSS.n1227 4.5005
R66567 VSS.n1754 VSS.n1280 4.5005
R66568 VSS.n1751 VSS.n1748 4.5005
R66569 VSS.n1747 VSS.n1746 4.5005
R66570 VSS.n1743 VSS.n1742 4.5005
R66571 VSS.n1745 VSS.n1742 4.5005
R66572 VSS.n1746 VSS.n1745 4.5005
R66573 VSS.n1751 VSS.n1281 4.5005
R66574 VSS.n1751 VSS.n1280 4.5005
R66575 VSS.n1751 VSS.n1227 4.5005
R66576 VSS.n2986 VSS.n1082 4.5005
R66577 VSS.n2986 VSS.n2985 4.5005
R66578 VSS.n4765 VSS.n4514 4.5005
R66579 VSS.n4846 VSS.n4449 4.5005
R66580 VSS.n4834 VSS.n4449 4.5005
R66581 VSS.n4822 VSS.n4449 4.5005
R66582 VSS.n4810 VSS.n4449 4.5005
R66583 VSS.n5991 VSS.n4449 4.5005
R66584 VSS.n5996 VSS.n4454 4.5005
R66585 VSS.n5646 VSS.n5185 4.5005
R66586 VSS.n5643 VSS.n5202 4.5005
R66587 VSS.n5646 VSS.n5189 4.5005
R66588 VSS.n5646 VSS.n5183 4.5005
R66589 VSS.n5646 VSS.n5190 4.5005
R66590 VSS.n5646 VSS.n5181 4.5005
R66591 VSS.n5646 VSS.n5191 4.5005
R66592 VSS.n5643 VSS.n5640 4.5005
R66593 VSS.n5643 VSS.n5196 4.5005
R66594 VSS.n5643 VSS.n5641 4.5005
R66595 VSS.n5644 VSS.n5643 4.5005
R66596 VSS.n5643 VSS.n5642 4.5005
R66597 VSS.n5797 VSS.n5076 4.5005
R66598 VSS.n5797 VSS.n5793 4.5005
R66599 VSS.n5804 VSS.n5063 4.5005
R66600 VSS.n5804 VSS.n5066 4.5005
R66601 VSS.n5804 VSS.n5061 4.5005
R66602 VSS.n5804 VSS.n5067 4.5005
R66603 VSS.n5804 VSS.n5059 4.5005
R66604 VSS.n5804 VSS.n5052 4.5005
R66605 VSS.n5805 VSS.n5804 4.5005
R66606 VSS.n5804 VSS.n5068 4.5005
R66607 VSS.n5797 VSS.n5055 4.5005
R66608 VSS.n5804 VSS.n5055 4.5005
R66609 VSS.n5797 VSS.n5069 4.5005
R66610 VSS.n5804 VSS.n5069 4.5005
R66611 VSS.n4471 VSS.n4449 4.5005
R66612 VSS.n4187 VSS.n535 4.5005
R66613 VSS.n4197 VSS.n4196 4.5005
R66614 VSS.n4187 VSS.n4186 4.5005
R66615 VSS.n4196 VSS.n4195 4.5005
R66616 VSS.n6174 VSS.n469 4.5005
R66617 VSS.n470 VSS.n469 4.5005
R66618 VSS.n2938 VSS.n1147 4.5005
R66619 VSS.n2928 VSS.n1155 4.5005
R66620 VSS.n2928 VSS.n2927 4.5005
R66621 VSS.n2932 VSS.n2931 4.5005
R66622 VSS.n2936 VSS.n2935 4.5005
R66623 VSS.n2938 VSS.n2937 4.5005
R66624 VSS.n2933 VSS.n1150 4.5005
R66625 VSS.n2929 VSS.n1153 4.5005
R66626 VSS.n2927 VSS.n2926 4.5005
R66627 VSS.n2926 VSS.n1155 4.5005
R66628 VSS.n2916 VSS.n1101 4.5005
R66629 VSS.n2916 VSS.n2915 4.5005
R66630 VSS.n1896 VSS.n1213 4.5005
R66631 VSS.n1894 VSS.n1213 4.5005
R66632 VSS.n1896 VSS.n1895 4.5005
R66633 VSS.n1895 VSS.n1894 4.5005
R66634 VSS.n6104 VSS.n4300 4.5005
R66635 VSS.n6104 VSS.n4303 4.5005
R66636 VSS.n6104 VSS.n4298 4.5005
R66637 VSS.n6104 VSS.n4305 4.5005
R66638 VSS.n6108 VSS.n6107 4.5005
R66639 VSS.n6121 VSS.n6113 4.5005
R66640 VSS.n6121 VSS.n4272 4.5005
R66641 VSS.n6116 VSS.n4268 4.5005
R66642 VSS.n6122 VSS.n4268 4.5005
R66643 VSS.n6122 VSS.n6121 4.5005
R66644 VSS.n6121 VSS.n4267 4.5005
R66645 VSS.n6121 VSS.n6120 4.5005
R66646 VSS.n3937 VSS.n456 4.5005
R66647 VSS.n3934 VSS.n3933 4.5005
R66648 VSS.n963 VSS.n664 4.5005
R66649 VSS.n3509 VSS.n963 4.5005
R66650 VSS.n2859 VSS.n968 4.5005
R66651 VSS.n2870 VSS.n1163 4.5005
R66652 VSS.n2871 VSS.n1161 4.5005
R66653 VSS.n2873 VSS.n1161 4.5005
R66654 VSS.n2917 VSS.n1161 4.5005
R66655 VSS.n2925 VSS.n1160 4.5005
R66656 VSS.n1160 VSS.n1159 4.5005
R66657 VSS.n1161 VSS.n1159 4.5005
R66658 VSS.n1160 VSS.n1156 4.5005
R66659 VSS.n1161 VSS.n1156 4.5005
R66660 VSS.n1536 VSS.n1533 4.5005
R66661 VSS.n1355 VSS.n1216 4.5005
R66662 VSS.n1536 VSS.n1215 4.5005
R66663 VSS.n1536 VSS.n1535 4.5005
R66664 VSS.n1543 VSS.n1355 4.5005
R66665 VSS.n1544 VSS.n1342 4.5005
R66666 VSS.n1617 VSS.n1347 4.5005
R66667 VSS.n1617 VSS.n1616 4.5005
R66668 VSS.n1616 VSS.n1342 4.5005
R66669 VSS.n1537 VSS.n1355 4.5005
R66670 VSS.n1535 VSS.n1355 4.5005
R66671 VSS.n1355 VSS.n1215 4.5005
R66672 VSS.n2919 VSS.n1160 4.5005
R66673 VSS.n2917 VSS.n1160 4.5005
R66674 VSS.n4507 VSS.n4268 4.5005
R66675 VSS.n6104 VSS.n4297 4.5005
R66676 VSS.n6104 VSS.n4306 4.5005
R66677 VSS.n6104 VSS.n4296 4.5005
R66678 VSS.n6104 VSS.n4307 4.5005
R66679 VSS.n6104 VSS.n4295 4.5005
R66680 VSS.n6107 VSS.n4281 4.5005
R66681 VSS.n5622 VSS.n5296 4.5005
R66682 VSS.n5619 VSS.n5311 4.5005
R66683 VSS.n5622 VSS.n5300 4.5005
R66684 VSS.n5622 VSS.n5294 4.5005
R66685 VSS.n5622 VSS.n5301 4.5005
R66686 VSS.n5622 VSS.n5287 4.5005
R66687 VSS.n5623 VSS.n5622 4.5005
R66688 VSS.n5619 VSS.n5616 4.5005
R66689 VSS.n5619 VSS.n5306 4.5005
R66690 VSS.n5619 VSS.n5617 4.5005
R66691 VSS.n5620 VSS.n5619 4.5005
R66692 VSS.n5619 VSS.n5618 4.5005
R66693 VSS.n5781 VSS.n5777 4.5005
R66694 VSS.n5781 VSS.n5080 4.5005
R66695 VSS.n5785 VSS.n5784 4.5005
R66696 VSS.n5784 VSS.n5104 4.5005
R66697 VSS.n5784 VSS.n5089 4.5005
R66698 VSS.n5784 VSS.n5115 4.5005
R66699 VSS.n5784 VSS.n5087 4.5005
R66700 VSS.n5784 VSS.n5119 4.5005
R66701 VSS.n5784 VSS.n5085 4.5005
R66702 VSS.n5784 VSS.n5014 4.5005
R66703 VSS.n5781 VSS.n5015 4.5005
R66704 VSS.n5784 VSS.n5015 4.5005
R66705 VSS.n5781 VSS.n5120 4.5005
R66706 VSS.n5784 VSS.n5120 4.5005
R66707 VSS.n6104 VSS.n6103 4.5005
R66708 VSS.n6125 VSS.n6124 4.5005
R66709 VSS.n6124 VSS.n6123 4.5005
R66710 VSS.n6146 VSS.n6145 4.5005
R66711 VSS.n6145 VSS.n6144 4.5005
R66712 VSS.n6143 VSS.n6142 4.5005
R66713 VSS.n6142 VSS.n6141 4.5005
R66714 VSS.n6127 VSS.n474 4.5005
R66715 VSS.n6127 VSS.n6126 4.5005
R66716 VSS.n6173 VSS.n472 4.5005
R66717 VSS.n6173 VSS.n6172 4.5005
R66718 VSS.n1212 VSS.n1211 4.5005
R66719 VSS.n1900 VSS.n1212 4.5005
R66720 VSS.n1901 VSS.n1211 4.5005
R66721 VSS.n1901 VSS.n1900 4.5005
R66722 VSS.n6098 VSS.n4317 4.5005
R66723 VSS.n6098 VSS.n4321 4.5005
R66724 VSS.n6098 VSS.n4315 4.5005
R66725 VSS.n6098 VSS.n4323 4.5005
R66726 VSS.n6095 VSS.n6094 4.5005
R66727 VSS.n6129 VSS.n4256 4.5005
R66728 VSS.n6129 VSS.n4254 4.5005
R66729 VSS.n4264 VSS.n4263 4.5005
R66730 VSS.n6128 VSS.n4263 4.5005
R66731 VSS.n6129 VSS.n6128 4.5005
R66732 VSS.n6129 VSS.n4252 4.5005
R66733 VSS.n6130 VSS.n6129 4.5005
R66734 VSS.n2204 VSS.n2203 4.5005
R66735 VSS.n2215 VSS.n2150 4.5005
R66736 VSS.n2149 VSS.n2148 4.5005
R66737 VSS.n2148 VSS.n2147 4.5005
R66738 VSS.n2687 VSS.n2686 4.5005
R66739 VSS.n2057 VSS.n1184 4.5005
R66740 VSS.n2056 VSS.n2055 4.5005
R66741 VSS.n1909 VSS.n1908 4.5005
R66742 VSS.n1907 VSS.n1906 4.5005
R66743 VSS.n1903 VSS.n1902 4.5005
R66744 VSS.n1906 VSS.n1203 4.5005
R66745 VSS.n1906 VSS.n1206 4.5005
R66746 VSS.n1903 VSS.n1209 4.5005
R66747 VSS.n1595 VSS.n1594 4.5005
R66748 VSS.n1604 VSS.n1548 4.5005
R66749 VSS.n1548 VSS.n1547 4.5005
R66750 VSS.n1594 VSS.n1547 4.5005
R66751 VSS.n1903 VSS.n1207 4.5005
R66752 VSS.n1903 VSS.n1206 4.5005
R66753 VSS.n1903 VSS.n1203 4.5005
R66754 VSS.n4509 VSS.n4263 4.5005
R66755 VSS.n6098 VSS.n4313 4.5005
R66756 VSS.n6098 VSS.n4324 4.5005
R66757 VSS.n6098 VSS.n4312 4.5005
R66758 VSS.n6098 VSS.n4325 4.5005
R66759 VSS.n6099 VSS.n6098 4.5005
R66760 VSS.n6095 VSS.n4327 4.5005
R66761 VSS.n5629 VSS.n5281 4.5005
R66762 VSS.n5632 VSS.n5269 4.5005
R66763 VSS.n5629 VSS.n5284 4.5005
R66764 VSS.n5629 VSS.n5279 4.5005
R66765 VSS.n5629 VSS.n5285 4.5005
R66766 VSS.n5629 VSS.n5277 4.5005
R66767 VSS.n5629 VSS.n5627 4.5005
R66768 VSS.n5632 VSS.n5258 4.5005
R66769 VSS.n5633 VSS.n5632 4.5005
R66770 VSS.n5632 VSS.n5631 4.5005
R66771 VSS.n5632 VSS.n5262 4.5005
R66772 VSS.n5632 VSS.n4980 4.5005
R66773 VSS.n5843 VSS.n5842 4.5005
R66774 VSS.n5842 VSS.n4991 4.5005
R66775 VSS.n5840 VSS.n5006 4.5005
R66776 VSS.n5840 VSS.n5008 4.5005
R66777 VSS.n5840 VSS.n5004 4.5005
R66778 VSS.n5840 VSS.n5009 4.5005
R66779 VSS.n5840 VSS.n5002 4.5005
R66780 VSS.n5840 VSS.n5010 4.5005
R66781 VSS.n5840 VSS.n5000 4.5005
R66782 VSS.n5840 VSS.n5839 4.5005
R66783 VSS.n5842 VSS.n4984 4.5005
R66784 VSS.n5840 VSS.n4984 4.5005
R66785 VSS.n5842 VSS.n5841 4.5005
R66786 VSS.n5841 VSS.n5840 4.5005
R66787 VSS.n6098 VSS.n4309 4.5005
R66788 VSS.n5492 VSS.n5490 4.5005
R66789 VSS.n5499 VSS.n5496 4.5005
R66790 VSS.n5487 VSS.n5485 4.5005
R66791 VSS.n5861 VSS.n5857 4.5005
R66792 VSS.n5491 VSS.n5490 4.5005
R66793 VSS.n5499 VSS.n5498 4.5005
R66794 VSS.n5487 VSS.n5486 4.5005
R66795 VSS.n5861 VSS.n5860 4.5005
R66796 VSS.n6160 VSS.n6159 4.5005
R66797 VSS.n6187 VSS.n458 4.5005
R66798 VSS.n4094 VSS.n4093 4.5005
R66799 VSS.n4096 VSS.n552 4.5005
R66800 VSS.n6157 VSS.n6156 4.5005
R66801 VSS.n6190 VSS.n457 4.5005
R66802 VSS.n573 VSS.n558 4.5005
R66803 VSS.n4099 VSS.n4095 4.5005
R66804 VSS.n5011 VSS.n4996 4.5005
R66805 VSS.n5837 VSS.n4996 4.5005
R66806 VSS.n5835 VSS.n5012 4.5005
R66807 VSS.n5833 VSS.n5012 4.5005
R66808 VSS.n5798 VSS.n5023 4.5005
R66809 VSS.n5800 VSS.n5798 4.5005
R66810 VSS.n4945 VSS.n4944 4.5005
R66811 VSS.n5864 VSS.n4945 4.5005
R66812 VSS.n5838 VSS.n5011 4.5005
R66813 VSS.n5838 VSS.n5837 4.5005
R66814 VSS.n5835 VSS.n5834 4.5005
R66815 VSS.n5834 VSS.n5833 4.5005
R66816 VSS.n5799 VSS.n5023 4.5005
R66817 VSS.n5800 VSS.n5799 4.5005
R66818 VSS.n5863 VSS.n4944 4.5005
R66819 VSS.n5864 VSS.n5863 4.5005
R66820 VSS.n5832 VSS.n5831 4.5005
R66821 VSS.n5831 VSS.n5020 4.5005
R66822 VSS.n5831 VSS.n5830 4.5005
R66823 VSS.n5832 VSS.n5017 4.5005
R66824 VSS.n5829 VSS.n5828 4.5005
R66825 VSS.n5829 VSS.n5025 4.5005
R66826 VSS.n5830 VSS.n5829 4.5005
R66827 VSS.n4134 VSS.n555 4.5005
R66828 VSS.n4134 VSS.n4133 4.5005
R66829 VSS.n4130 VSS.n557 4.5005
R66830 VSS.n557 VSS.n555 4.5005
R66831 VSS.n4133 VSS.n557 4.5005
R66832 VSS.n4132 VSS.n4130 4.5005
R66833 VSS.n4133 VSS.n4132 4.5005
R66834 VSS.n5503 VSS.n5482 4.5005
R66835 VSS.n5503 VSS.n5502 4.5005
R66836 VSS.n6149 VSS.n6148 4.5005
R66837 VSS.n4183 VSS.n4182 4.5005
R66838 VSS.n4188 VSS.n4183 4.5005
R66839 VSS.n4189 VSS.n4179 4.5005
R66840 VSS.n4189 VSS.n4188 4.5005
R66841 VSS.n481 VSS.n480 4.5005
R66842 VSS.n5501 VSS.n5500 4.5005
R66843 VSS.n5502 VSS.n5501 4.5005
R66844 VSS.n2942 VSS.n1142 4.5005
R66845 VSS.n1118 VSS.n1112 4.5005
R66846 VSS.n2971 VSS.n1112 4.5005
R66847 VSS.n2969 VSS.n1112 4.5005
R66848 VSS.n2965 VSS.n1112 4.5005
R66849 VSS.n2897 VSS.n2896 4.5005
R66850 VSS.n2898 VSS.n2897 4.5005
R66851 VSS.n2899 VSS.n2898 4.5005
R66852 VSS.n2885 VSS.n2883 4.5005
R66853 VSS.n2885 VSS.n1136 4.5005
R66854 VSS.n1145 VSS.n1136 4.5005
R66855 VSS.n2942 VSS.n2941 4.5005
R66856 VSS.n2941 VSS.n1144 4.5005
R66857 VSS.n2941 VSS.n2940 4.5005
R66858 VSS.n2900 VSS.n2883 4.5005
R66859 VSS.n2896 VSS.n2895 4.5005
R66860 VSS.n2970 VSS.n2965 4.5005
R66861 VSS.n2970 VSS.n2969 4.5005
R66862 VSS.n2971 VSS.n2970 4.5005
R66863 VSS.n2970 VSS.n1118 4.5005
R66864 VSS.n2981 VSS.n2980 4.5005
R66865 VSS.n2980 VSS.n1100 4.5005
R66866 VSS.n2980 VSS.n1098 4.5005
R66867 VSS.n2980 VSS.n2979 4.5005
R66868 VSS.n1893 VSS.n1221 4.5005
R66869 VSS.n1891 VSS.n1221 4.5005
R66870 VSS.n1893 VSS.n1217 4.5005
R66871 VSS.n1891 VSS.n1217 4.5005
R66872 VSS.n1893 VSS.n1892 4.5005
R66873 VSS.n1892 VSS.n1891 4.5005
R66874 VSS.n6033 VSS.n4397 4.5005
R66875 VSS.n6031 VSS.n4397 4.5005
R66876 VSS.n6033 VSS.n4398 4.5005
R66877 VSS.n6031 VSS.n4398 4.5005
R66878 VSS.n6031 VSS.n4424 4.5005
R66879 VSS.n6033 VSS.n4399 4.5005
R66880 VSS.n6031 VSS.n4399 4.5005
R66881 VSS.n6033 VSS.n4395 4.5005
R66882 VSS.n6031 VSS.n4395 4.5005
R66883 VSS.n6033 VSS.n4401 4.5005
R66884 VSS.n4420 VSS.n4401 4.5005
R66885 VSS.n6031 VSS.n4401 4.5005
R66886 VSS.n6033 VSS.n4394 4.5005
R66887 VSS.n6031 VSS.n4394 4.5005
R66888 VSS.n6033 VSS.n4403 4.5005
R66889 VSS.n6031 VSS.n4403 4.5005
R66890 VSS.n6033 VSS.n4392 4.5005
R66891 VSS.n4420 VSS.n4392 4.5005
R66892 VSS.n6031 VSS.n4392 4.5005
R66893 VSS.n6033 VSS.n4404 4.5005
R66894 VSS.n6031 VSS.n4404 4.5005
R66895 VSS.n6033 VSS.n4391 4.5005
R66896 VSS.n6031 VSS.n4391 4.5005
R66897 VSS.n6033 VSS.n4406 4.5005
R66898 VSS.n4420 VSS.n4406 4.5005
R66899 VSS.n6031 VSS.n4406 4.5005
R66900 VSS.n6033 VSS.n4390 4.5005
R66901 VSS.n6031 VSS.n4390 4.5005
R66902 VSS.n4407 VSS.n4381 4.5005
R66903 VSS.n6033 VSS.n4407 4.5005
R66904 VSS.n6031 VSS.n4407 4.5005
R66905 VSS.n4776 VSS.n4488 4.5005
R66906 VSS.n4776 VSS.n4489 4.5005
R66907 VSS.n4776 VSS.n4775 4.5005
R66908 VSS.n4495 VSS.n4488 4.5005
R66909 VSS.n4495 VSS.n4489 4.5005
R66910 VSS.n4775 VSS.n4495 4.5005
R66911 VSS.n4497 VSS.n4489 4.5005
R66912 VSS.n4775 VSS.n4497 4.5005
R66913 VSS.n4494 VSS.n4489 4.5005
R66914 VSS.n4775 VSS.n4494 4.5005
R66915 VSS.n4499 VSS.n4489 4.5005
R66916 VSS.n4775 VSS.n4499 4.5005
R66917 VSS.n4493 VSS.n4489 4.5005
R66918 VSS.n4775 VSS.n4493 4.5005
R66919 VSS.n4775 VSS.n483 4.5005
R66920 VSS.n4488 VSS.n482 4.5005
R66921 VSS.n4489 VSS.n482 4.5005
R66922 VSS.n4506 VSS.n482 4.5005
R66923 VSS.n4775 VSS.n482 4.5005
R66924 VSS.n4500 VSS.n4488 4.5005
R66925 VSS.n4500 VSS.n4489 4.5005
R66926 VSS.n4775 VSS.n4500 4.5005
R66927 VSS.n4491 VSS.n4488 4.5005
R66928 VSS.n4491 VSS.n4489 4.5005
R66929 VSS.n4775 VSS.n4491 4.5005
R66930 VSS.n3974 VSS.n559 4.5005
R66931 VSS.n3976 VSS.n559 4.5005
R66932 VSS.n3979 VSS.n559 4.5005
R66933 VSS.n3976 VSS.n628 4.5005
R66934 VSS.n3979 VSS.n628 4.5005
R66935 VSS.n3976 VSS.n630 4.5005
R66936 VSS.n3979 VSS.n630 4.5005
R66937 VSS.n3976 VSS.n626 4.5005
R66938 VSS.n3979 VSS.n626 4.5005
R66939 VSS.n3976 VSS.n632 4.5005
R66940 VSS.n3979 VSS.n632 4.5005
R66941 VSS.n3976 VSS.n625 4.5005
R66942 VSS.n3979 VSS.n625 4.5005
R66943 VSS.n3976 VSS.n634 4.5005
R66944 VSS.n3979 VSS.n634 4.5005
R66945 VSS.n3976 VSS.n624 4.5005
R66946 VSS.n3979 VSS.n624 4.5005
R66947 VSS.n3976 VSS.n636 4.5005
R66948 VSS.n3979 VSS.n636 4.5005
R66949 VSS.n3976 VSS.n623 4.5005
R66950 VSS.n3979 VSS.n623 4.5005
R66951 VSS.n3979 VSS.n3978 4.5005
R66952 VSS.n947 VSS.n924 4.5005
R66953 VSS.n3589 VSS.n924 4.5005
R66954 VSS.n3591 VSS.n924 4.5005
R66955 VSS.n3589 VSS.n925 4.5005
R66956 VSS.n3591 VSS.n925 4.5005
R66957 VSS.n3589 VSS.n921 4.5005
R66958 VSS.n3591 VSS.n921 4.5005
R66959 VSS.n3589 VSS.n926 4.5005
R66960 VSS.n3591 VSS.n926 4.5005
R66961 VSS.n3589 VSS.n920 4.5005
R66962 VSS.n3591 VSS.n920 4.5005
R66963 VSS.n3589 VSS.n927 4.5005
R66964 VSS.n3591 VSS.n927 4.5005
R66965 VSS.n3589 VSS.n919 4.5005
R66966 VSS.n3591 VSS.n919 4.5005
R66967 VSS.n3589 VSS.n928 4.5005
R66968 VSS.n3591 VSS.n928 4.5005
R66969 VSS.n3589 VSS.n918 4.5005
R66970 VSS.n3591 VSS.n918 4.5005
R66971 VSS.n3589 VSS.n929 4.5005
R66972 VSS.n3591 VSS.n929 4.5005
R66973 VSS.n3589 VSS.n917 4.5005
R66974 VSS.n3591 VSS.n917 4.5005
R66975 VSS.n3589 VSS.n930 4.5005
R66976 VSS.n3591 VSS.n930 4.5005
R66977 VSS.n3589 VSS.n916 4.5005
R66978 VSS.n3591 VSS.n916 4.5005
R66979 VSS.n3589 VSS.n931 4.5005
R66980 VSS.n3591 VSS.n931 4.5005
R66981 VSS.n3589 VSS.n915 4.5005
R66982 VSS.n3591 VSS.n915 4.5005
R66983 VSS.n3589 VSS.n932 4.5005
R66984 VSS.n3591 VSS.n932 4.5005
R66985 VSS.n3589 VSS.n914 4.5005
R66986 VSS.n3591 VSS.n914 4.5005
R66987 VSS.n3589 VSS.n933 4.5005
R66988 VSS.n3591 VSS.n933 4.5005
R66989 VSS.n3589 VSS.n913 4.5005
R66990 VSS.n3591 VSS.n913 4.5005
R66991 VSS.n3589 VSS.n934 4.5005
R66992 VSS.n3591 VSS.n934 4.5005
R66993 VSS.n3589 VSS.n912 4.5005
R66994 VSS.n3591 VSS.n912 4.5005
R66995 VSS.n3590 VSS.n3589 4.5005
R66996 VSS.n3591 VSS.n3590 4.5005
R66997 VSS.n3591 VSS.n732 4.5005
R66998 VSS.n3591 VSS.n730 4.5005
R66999 VSS.n2826 VSS.n2825 4.5005
R67000 VSS.n2825 VSS.n2746 4.5005
R67001 VSS.n2825 VSS.n2824 4.5005
R67002 VSS.n2752 VSS.n2746 4.5005
R67003 VSS.n2824 VSS.n2752 4.5005
R67004 VSS.n2812 VSS.n2746 4.5005
R67005 VSS.n2824 VSS.n2812 4.5005
R67006 VSS.n2751 VSS.n2746 4.5005
R67007 VSS.n2824 VSS.n2751 4.5005
R67008 VSS.n2813 VSS.n2746 4.5005
R67009 VSS.n2824 VSS.n2813 4.5005
R67010 VSS.n2750 VSS.n2746 4.5005
R67011 VSS.n2824 VSS.n2750 4.5005
R67012 VSS.n2814 VSS.n2746 4.5005
R67013 VSS.n2824 VSS.n2814 4.5005
R67014 VSS.n2749 VSS.n2746 4.5005
R67015 VSS.n2824 VSS.n2749 4.5005
R67016 VSS.n2815 VSS.n2746 4.5005
R67017 VSS.n2824 VSS.n2815 4.5005
R67018 VSS.n2748 VSS.n2746 4.5005
R67019 VSS.n2824 VSS.n2748 4.5005
R67020 VSS.n2824 VSS.n2823 4.5005
R67021 VSS.n2816 VSS.n1116 4.5005
R67022 VSS.n2816 VSS.n1103 4.5005
R67023 VSS.n2816 VSS.n1104 4.5005
R67024 VSS.n1116 VSS.n1099 4.5005
R67025 VSS.n1103 VSS.n1099 4.5005
R67026 VSS.n1104 VSS.n1099 4.5005
R67027 VSS.n1104 VSS.n1097 4.5005
R67028 VSS.n2976 VSS.n1104 4.5005
R67029 VSS.n1109 VSS.n1103 4.5005
R67030 VSS.n1109 VSS.n1104 4.5005
R67031 VSS.n1114 VSS.n1103 4.5005
R67032 VSS.n1114 VSS.n1104 4.5005
R67033 VSS.n1113 VSS.n1103 4.5005
R67034 VSS.n1113 VSS.n1104 4.5005
R67035 VSS.n2966 VSS.n1103 4.5005
R67036 VSS.n2966 VSS.n1104 4.5005
R67037 VSS.n2968 VSS.n1104 4.5005
R67038 VSS.n1116 VSS.n1106 4.5005
R67039 VSS.n1106 VSS.n1103 4.5005
R67040 VSS.n2975 VSS.n1106 4.5005
R67041 VSS.n1106 VSS.n1104 4.5005
R67042 VSS.n2974 VSS.n1116 4.5005
R67043 VSS.n2974 VSS.n1103 4.5005
R67044 VSS.n2975 VSS.n2974 4.5005
R67045 VSS.n2974 VSS.n1104 4.5005
R67046 VSS.n1499 VSS.n1427 4.5005
R67047 VSS.n1432 VSS.n1427 4.5005
R67048 VSS.n1496 VSS.n1427 4.5005
R67049 VSS.n1436 VSS.n1432 4.5005
R67050 VSS.n1496 VSS.n1436 4.5005
R67051 VSS.n1496 VSS.n1224 4.5005
R67052 VSS.n1497 VSS.n1432 4.5005
R67053 VSS.n1497 VSS.n1496 4.5005
R67054 VSS.n1490 VSS.n1432 4.5005
R67055 VSS.n1496 VSS.n1490 4.5005
R67056 VSS.n1435 VSS.n1432 4.5005
R67057 VSS.n1496 VSS.n1435 4.5005
R67058 VSS.n1495 VSS.n1432 4.5005
R67059 VSS.n1496 VSS.n1495 4.5005
R67060 VSS.n1434 VSS.n1432 4.5005
R67061 VSS.n1493 VSS.n1434 4.5005
R67062 VSS.n1496 VSS.n1434 4.5005
R67063 VSS.n1325 VSS.n1311 4.5005
R67064 VSS.n1661 VSS.n1311 4.5005
R67065 VSS.n1663 VSS.n1311 4.5005
R67066 VSS.n1661 VSS.n1312 4.5005
R67067 VSS.n1663 VSS.n1312 4.5005
R67068 VSS.n1661 VSS.n1310 4.5005
R67069 VSS.n1663 VSS.n1310 4.5005
R67070 VSS.n1661 VSS.n1313 4.5005
R67071 VSS.n1663 VSS.n1313 4.5005
R67072 VSS.n1661 VSS.n1309 4.5005
R67073 VSS.n1663 VSS.n1309 4.5005
R67074 VSS.n1661 VSS.n1314 4.5005
R67075 VSS.n1663 VSS.n1314 4.5005
R67076 VSS.n1661 VSS.n1308 4.5005
R67077 VSS.n1663 VSS.n1308 4.5005
R67078 VSS.n1661 VSS.n1315 4.5005
R67079 VSS.n1663 VSS.n1315 4.5005
R67080 VSS.n1663 VSS.n1307 4.5005
R67081 VSS.n1662 VSS.n1325 4.5005
R67082 VSS.n1662 VSS.n1661 4.5005
R67083 VSS.n1662 VSS.n1320 4.5005
R67084 VSS.n1663 VSS.n1662 4.5005
R67085 VSS.n1432 VSS.n1430 4.5005
R67086 VSS.n1493 VSS.n1430 4.5005
R67087 VSS.n1496 VSS.n1430 4.5005
R67088 VSS.n1499 VSS.n1424 4.5005
R67089 VSS.n1432 VSS.n1424 4.5005
R67090 VSS.n1493 VSS.n1424 4.5005
R67091 VSS.n1496 VSS.n1424 4.5005
R67092 VSS.n1499 VSS.n1222 4.5005
R67093 VSS.n1432 VSS.n1222 4.5005
R67094 VSS.n1493 VSS.n1222 4.5005
R67095 VSS.n1496 VSS.n1222 4.5005
R67096 VSS.n2976 VSS.n2975 4.5005
R67097 VSS.n2976 VSS.n1103 4.5005
R67098 VSS.n2975 VSS.n1097 4.5005
R67099 VSS.n1103 VSS.n1097 4.5005
R67100 VSS.n1116 VSS.n1097 4.5005
R67101 VSS.n3587 VSS.n730 4.5005
R67102 VSS.n3589 VSS.n730 4.5005
R67103 VSS.n947 VSS.n730 4.5005
R67104 VSS.n4774 VSS.n4489 4.5005
R67105 VSS.n4774 VSS.n4506 4.5005
R67106 VSS.n4775 VSS.n4774 4.5005
R67107 VSS.n6033 VSS.n4388 4.5005
R67108 VSS.n4420 VSS.n4388 4.5005
R67109 VSS.n6031 VSS.n4388 4.5005
R67110 VSS.n6033 VSS.n4409 4.5005
R67111 VSS.n4420 VSS.n4409 4.5005
R67112 VSS.n6031 VSS.n4409 4.5005
R67113 VSS.n6033 VSS.n4387 4.5005
R67114 VSS.n4420 VSS.n4387 4.5005
R67115 VSS.n6031 VSS.n4387 4.5005
R67116 VSS.n6033 VSS.n4411 4.5005
R67117 VSS.n4420 VSS.n4411 4.5005
R67118 VSS.n6031 VSS.n4411 4.5005
R67119 VSS.n6032 VSS.n4420 4.5005
R67120 VSS.n6032 VSS.n6031 4.5005
R67121 VSS.n6031 VSS.n6025 4.5005
R67122 VSS.n6025 VSS.n4420 4.5005
R67123 VSS.n6025 VSS.n4381 4.5005
R67124 VSS.n6027 VSS.n4420 4.5005
R67125 VSS.n6027 VSS.n4381 4.5005
R67126 VSS.n6026 VSS.n4420 4.5005
R67127 VSS.n6026 VSS.n4381 4.5005
R67128 VSS.n6029 VSS.n4420 4.5005
R67129 VSS.n6029 VSS.n4381 4.5005
R67130 VSS.n4420 VSS.n4386 4.5005
R67131 VSS.n6033 VSS.n4386 4.5005
R67132 VSS.n4386 VSS.n4381 4.5005
R67133 VSS.n5578 VSS.n5504 4.5005
R67134 VSS.n5581 VSS.n5504 4.5005
R67135 VSS.n5504 VSS.n5447 4.5005
R67136 VSS.n5581 VSS.n5506 4.5005
R67137 VSS.n5506 VSS.n5447 4.5005
R67138 VSS.n5581 VSS.n5479 4.5005
R67139 VSS.n5479 VSS.n5447 4.5005
R67140 VSS.n5581 VSS.n5507 4.5005
R67141 VSS.n5507 VSS.n5447 4.5005
R67142 VSS.n5537 VSS.n5447 4.5005
R67143 VSS.n5578 VSS.n5508 4.5005
R67144 VSS.n5581 VSS.n5508 4.5005
R67145 VSS.n5508 VSS.n5447 4.5005
R67146 VSS.n5581 VSS.n5478 4.5005
R67147 VSS.n5478 VSS.n5447 4.5005
R67148 VSS.n5581 VSS.n5509 4.5005
R67149 VSS.n5509 VSS.n5447 4.5005
R67150 VSS.n5578 VSS.n5477 4.5005
R67151 VSS.n5581 VSS.n5477 4.5005
R67152 VSS.n5477 VSS.n5447 4.5005
R67153 VSS.n5578 VSS.n5519 4.5005
R67154 VSS.n5581 VSS.n5519 4.5005
R67155 VSS.n5519 VSS.n5447 4.5005
R67156 VSS.n5581 VSS.n5476 4.5005
R67157 VSS.n5476 VSS.n5447 4.5005
R67158 VSS.n5581 VSS.n5520 4.5005
R67159 VSS.n5520 VSS.n5447 4.5005
R67160 VSS.n5578 VSS.n5475 4.5005
R67161 VSS.n5581 VSS.n5475 4.5005
R67162 VSS.n5475 VSS.n5447 4.5005
R67163 VSS.n5578 VSS.n5526 4.5005
R67164 VSS.n5581 VSS.n5526 4.5005
R67165 VSS.n5526 VSS.n5447 4.5005
R67166 VSS.n5581 VSS.n5474 4.5005
R67167 VSS.n5474 VSS.n5447 4.5005
R67168 VSS.n5581 VSS.n5464 4.5005
R67169 VSS.n5583 VSS.n5464 4.5005
R67170 VSS.n5464 VSS.n5447 4.5005
R67171 VSS.n5455 VSS.n5447 4.5005
R67172 VSS.n5583 VSS.n5455 4.5005
R67173 VSS.n5578 VSS.n5455 4.5005
R67174 VSS.n5578 VSS.n5576 4.5005
R67175 VSS.n5576 VSS.n5447 4.5005
R67176 VSS.n5581 VSS.n5473 4.5005
R67177 VSS.n5473 VSS.n5447 4.5005
R67178 VSS.n5581 VSS.n5470 4.5005
R67179 VSS.n5583 VSS.n5470 4.5005
R67180 VSS.n5470 VSS.n5447 4.5005
R67181 VSS.n5453 VSS.n5447 4.5005
R67182 VSS.n5583 VSS.n5453 4.5005
R67183 VSS.n5578 VSS.n5453 4.5005
R67184 VSS.n5579 VSS.n5578 4.5005
R67185 VSS.n5579 VSS.n5447 4.5005
R67186 VSS.n5581 VSS.n5472 4.5005
R67187 VSS.n5472 VSS.n5447 4.5005
R67188 VSS.n5582 VSS.n5581 4.5005
R67189 VSS.n5583 VSS.n5582 4.5005
R67190 VSS.n5582 VSS.n5447 4.5005
R67191 VSS.n5825 VSS.n5034 4.5005
R67192 VSS.n5034 VSS.n5026 4.5005
R67193 VSS.n5034 VSS.n5027 4.5005
R67194 VSS.n5825 VSS.n5037 4.5005
R67195 VSS.n5037 VSS.n5026 4.5005
R67196 VSS.n5037 VSS.n5027 4.5005
R67197 VSS.n5033 VSS.n5027 4.5005
R67198 VSS.n5033 VSS.n5028 4.5005
R67199 VSS.n5825 VSS.n5033 4.5005
R67200 VSS.n5825 VSS.n5039 4.5005
R67201 VSS.n5039 VSS.n5027 4.5005
R67202 VSS.n5041 VSS.n5026 4.5005
R67203 VSS.n5041 VSS.n5027 4.5005
R67204 VSS.n5094 VSS.n5027 4.5005
R67205 VSS.n5032 VSS.n5027 4.5005
R67206 VSS.n5032 VSS.n5028 4.5005
R67207 VSS.n5825 VSS.n5032 4.5005
R67208 VSS.n5825 VSS.n5044 4.5005
R67209 VSS.n5044 VSS.n5027 4.5005
R67210 VSS.n5046 VSS.n5026 4.5005
R67211 VSS.n5046 VSS.n5027 4.5005
R67212 VSS.n5105 VSS.n5026 4.5005
R67213 VSS.n5105 VSS.n5028 4.5005
R67214 VSS.n5105 VSS.n5027 4.5005
R67215 VSS.n5031 VSS.n5027 4.5005
R67216 VSS.n5031 VSS.n5028 4.5005
R67217 VSS.n5825 VSS.n5031 4.5005
R67218 VSS.n5825 VSS.n5049 4.5005
R67219 VSS.n5049 VSS.n5027 4.5005
R67220 VSS.n5812 VSS.n5026 4.5005
R67221 VSS.n5812 VSS.n5027 4.5005
R67222 VSS.n5810 VSS.n5026 4.5005
R67223 VSS.n5810 VSS.n5028 4.5005
R67224 VSS.n5810 VSS.n5027 4.5005
R67225 VSS.n5030 VSS.n5027 4.5005
R67226 VSS.n5030 VSS.n5028 4.5005
R67227 VSS.n5825 VSS.n5030 4.5005
R67228 VSS.n5825 VSS.n5815 4.5005
R67229 VSS.n5815 VSS.n5027 4.5005
R67230 VSS.n5817 VSS.n5026 4.5005
R67231 VSS.n5817 VSS.n5027 4.5005
R67232 VSS.n5819 VSS.n5026 4.5005
R67233 VSS.n5819 VSS.n5027 4.5005
R67234 VSS.n5821 VSS.n5026 4.5005
R67235 VSS.n5821 VSS.n5027 4.5005
R67236 VSS.n5026 VSS.n5024 4.5005
R67237 VSS.n5028 VSS.n5024 4.5005
R67238 VSS.n5027 VSS.n5024 4.5005
R67239 VSS.n5826 VSS.n5027 4.5005
R67240 VSS.n5826 VSS.n5028 4.5005
R67241 VSS.n5826 VSS.n5026 4.5005
R67242 VSS.n5826 VSS.n5825 4.5005
R67243 VSS.n5027 VSS.n5018 4.5005
R67244 VSS.n5028 VSS.n5018 4.5005
R67245 VSS.n5026 VSS.n5018 4.5005
R67246 VSS.n5825 VSS.n5018 4.5005
R67247 VSS.n5825 VSS.n5021 4.5005
R67248 VSS.n5026 VSS.n5021 4.5005
R67249 VSS.n5027 VSS.n5021 4.5005
R67250 VSS.n5825 VSS.n5824 4.5005
R67251 VSS.n5824 VSS.n5026 4.5005
R67252 VSS.n5824 VSS.n5027 4.5005
R67253 VSS.n6033 VSS.n6032 4.5005
R67254 VSS.n738 VSS.n731 4.5005
R67255 VSS.n3861 VSS.n738 4.5005
R67256 VSS.n738 VSS.n725 4.5005
R67257 VSS.n3861 VSS.n3860 4.5005
R67258 VSS.n3860 VSS.n725 4.5005
R67259 VSS.n3861 VSS.n737 4.5005
R67260 VSS.n737 VSS.n725 4.5005
R67261 VSS.n735 VSS.n725 4.5005
R67262 VSS.n735 VSS.n731 4.5005
R67263 VSS.n731 VSS.n726 4.5005
R67264 VSS.n3863 VSS.n726 4.5005
R67265 VSS.n726 VSS.n725 4.5005
R67266 VSS.n3862 VSS.n731 4.5005
R67267 VSS.n3862 VSS.n3861 4.5005
R67268 VSS.n3863 VSS.n3862 4.5005
R67269 VSS.n3862 VSS.n725 4.5005
R67270 VSS.n6232 VSS.n6225 4.5005
R67271 VSS.n6234 VSS.n6233 4.5005
R67272 VSS.n6235 VSS.n123 4.5005
R67273 VSS.n6227 VSS.n6226 4.5005
R67274 VSS.n6231 VSS.n6230 4.5005
R67275 VSS.n445 VSS.n444 4.5005
R67276 VSS.n6 VSS.n5 4.5005
R67277 VSS.n440 VSS.n126 4.5005
R67278 VSS.n442 VSS.n441 4.5005
R67279 VSS.n133 VSS.n132 4.5005
R67280 VSS.n135 VSS.n134 4.5005
R67281 VSS.n142 VSS.n141 4.17693
R67282 VSS.n2680 VSS.n2076 3.91226
R67283 VSS.n2680 VSS.n2077 3.91226
R67284 VSS.n2676 VSS.n2077 3.91226
R67285 VSS.n2676 VSS.n2219 3.91226
R67286 VSS.n2668 VSS.n2219 3.91226
R67287 VSS.n2668 VSS.n2559 3.91226
R67288 VSS.n2664 VSS.n2559 3.91226
R67289 VSS.n2664 VSS.n2561 3.91226
R67290 VSS.n2656 VSS.n2561 3.91226
R67291 VSS.n2656 VSS.n2569 3.91226
R67292 VSS.n2652 VSS.n2569 3.91226
R67293 VSS.n2652 VSS.n2571 3.91226
R67294 VSS.n2644 VSS.n2571 3.91226
R67295 VSS.n2644 VSS.n2579 3.91226
R67296 VSS.n2640 VSS.n2579 3.91226
R67297 VSS.n2640 VSS.n2581 3.91226
R67298 VSS.n2632 VSS.n2581 3.91226
R67299 VSS.n2632 VSS.n2589 3.91226
R67300 VSS.n2628 VSS.n2589 3.91226
R67301 VSS.n2628 VSS.n2591 3.91226
R67302 VSS.n2591 VSS.n667 3.91226
R67303 VSS.n3928 VSS.n667 3.91226
R67304 VSS.n3928 VSS.n668 3.91226
R67305 VSS.n3919 VSS.n668 3.91226
R67306 VSS.n3919 VSS.n679 3.91226
R67307 VSS.n3915 VSS.n679 3.91226
R67308 VSS.n3915 VSS.n681 3.91226
R67309 VSS.n3907 VSS.n681 3.91226
R67310 VSS.n3907 VSS.n689 3.91226
R67311 VSS.n3903 VSS.n689 3.91226
R67312 VSS.n3903 VSS.n691 3.91226
R67313 VSS.n3895 VSS.n691 3.91226
R67314 VSS.n3895 VSS.n698 3.91226
R67315 VSS.n3891 VSS.n698 3.91226
R67316 VSS.n3891 VSS.n700 3.91226
R67317 VSS.n3883 VSS.n700 3.91226
R67318 VSS.n3883 VSS.n709 3.91226
R67319 VSS.n3879 VSS.n709 3.91226
R67320 VSS.n3879 VSS.n711 3.91226
R67321 VSS.n3871 VSS.n711 3.91226
R67322 VSS.n3871 VSS.n719 3.91226
R67323 VSS.n3867 VSS.n719 3.91226
R67324 VSS.n3867 VSS.n721 3.91226
R67325 VSS.n744 VSS.n721 3.91226
R67326 VSS.n3855 VSS.n744 3.91226
R67327 VSS.n3855 VSS.n745 3.91226
R67328 VSS.n3851 VSS.n745 3.91226
R67329 VSS.n3851 VSS.n748 3.91226
R67330 VSS.n3843 VSS.n748 3.91226
R67331 VSS.n3843 VSS.n757 3.91226
R67332 VSS.n3839 VSS.n757 3.91226
R67333 VSS.n3839 VSS.n759 3.91226
R67334 VSS.n3831 VSS.n759 3.91226
R67335 VSS.n3831 VSS.n767 3.91226
R67336 VSS.n3827 VSS.n767 3.91226
R67337 VSS.n3827 VSS.n769 3.91226
R67338 VSS.n3819 VSS.n769 3.91226
R67339 VSS.n3819 VSS.n777 3.91226
R67340 VSS.n3815 VSS.n777 3.91226
R67341 VSS.n3815 VSS.n779 3.91226
R67342 VSS.n3807 VSS.n779 3.91226
R67343 VSS.n3807 VSS.n787 3.91226
R67344 VSS.n3803 VSS.n787 3.91226
R67345 VSS.n3803 VSS.n789 3.91226
R67346 VSS.n3794 VSS.n789 3.91226
R67347 VSS.n3794 VSS.n797 3.91226
R67348 VSS.n3789 VSS.n797 3.91226
R67349 VSS.n3789 VSS.n799 3.91226
R67350 VSS.n3781 VSS.n799 3.91226
R67351 VSS.n3781 VSS.n808 3.91226
R67352 VSS.n3777 VSS.n808 3.91226
R67353 VSS.n3777 VSS.n810 3.91226
R67354 VSS.n3769 VSS.n810 3.91226
R67355 VSS.n3769 VSS.n818 3.91226
R67356 VSS.n3765 VSS.n818 3.91226
R67357 VSS.n3765 VSS.n820 3.91226
R67358 VSS.n3757 VSS.n820 3.91226
R67359 VSS.n3757 VSS.n828 3.91226
R67360 VSS.n3753 VSS.n828 3.91226
R67361 VSS.n3753 VSS.n830 3.91226
R67362 VSS.n3745 VSS.n830 3.91226
R67363 VSS.n3745 VSS.n838 3.91226
R67364 VSS.n3741 VSS.n838 3.91226
R67365 VSS.n3741 VSS.n840 3.91226
R67366 VSS.n3733 VSS.n840 3.91226
R67367 VSS.n3733 VSS.n848 3.91226
R67368 VSS.n3396 VSS.n848 3.91226
R67369 VSS.n2550 VSS.n2075 3.91226
R67370 VSS.n2222 VSS.n2075 3.91226
R67371 VSS.n2674 VSS.n2222 3.91226
R67372 VSS.n2674 VSS.n2223 3.91226
R67373 VSS.n2670 VSS.n2223 3.91226
R67374 VSS.n2670 VSS.n2556 3.91226
R67375 VSS.n2662 VSS.n2556 3.91226
R67376 VSS.n2662 VSS.n2564 3.91226
R67377 VSS.n2658 VSS.n2564 3.91226
R67378 VSS.n2658 VSS.n2566 3.91226
R67379 VSS.n2650 VSS.n2566 3.91226
R67380 VSS.n2650 VSS.n2574 3.91226
R67381 VSS.n2646 VSS.n2574 3.91226
R67382 VSS.n2646 VSS.n2576 3.91226
R67383 VSS.n2638 VSS.n2576 3.91226
R67384 VSS.n2638 VSS.n2584 3.91226
R67385 VSS.n2634 VSS.n2584 3.91226
R67386 VSS.n2634 VSS.n2586 3.91226
R67387 VSS.n2626 VSS.n2586 3.91226
R67388 VSS.n2626 VSS.n2622 3.91226
R67389 VSS.n2622 VSS.n672 3.91226
R67390 VSS.n3926 VSS.n672 3.91226
R67391 VSS.n3926 VSS.n673 3.91226
R67392 VSS.n3921 VSS.n673 3.91226
R67393 VSS.n3921 VSS.n676 3.91226
R67394 VSS.n3913 VSS.n676 3.91226
R67395 VSS.n3913 VSS.n684 3.91226
R67396 VSS.n3909 VSS.n684 3.91226
R67397 VSS.n3909 VSS.n686 3.91226
R67398 VSS.n3901 VSS.n686 3.91226
R67399 VSS.n3901 VSS.n694 3.91226
R67400 VSS.n3897 VSS.n694 3.91226
R67401 VSS.n3897 VSS.n695 3.91226
R67402 VSS.n3889 VSS.n695 3.91226
R67403 VSS.n3889 VSS.n703 3.91226
R67404 VSS.n3885 VSS.n703 3.91226
R67405 VSS.n3885 VSS.n706 3.91226
R67406 VSS.n3877 VSS.n706 3.91226
R67407 VSS.n3877 VSS.n714 3.91226
R67408 VSS.n3873 VSS.n714 3.91226
R67409 VSS.n3873 VSS.n716 3.91226
R67410 VSS.n3865 VSS.n716 3.91226
R67411 VSS.n3865 VSS.n724 3.91226
R67412 VSS.n739 VSS.n724 3.91226
R67413 VSS.n3857 VSS.n739 3.91226
R67414 VSS.n3857 VSS.n740 3.91226
R67415 VSS.n3849 VSS.n740 3.91226
R67416 VSS.n3849 VSS.n751 3.91226
R67417 VSS.n3845 VSS.n751 3.91226
R67418 VSS.n3845 VSS.n754 3.91226
R67419 VSS.n3837 VSS.n754 3.91226
R67420 VSS.n3837 VSS.n762 3.91226
R67421 VSS.n3833 VSS.n762 3.91226
R67422 VSS.n3833 VSS.n764 3.91226
R67423 VSS.n3825 VSS.n764 3.91226
R67424 VSS.n3825 VSS.n772 3.91226
R67425 VSS.n3821 VSS.n772 3.91226
R67426 VSS.n3821 VSS.n774 3.91226
R67427 VSS.n3813 VSS.n774 3.91226
R67428 VSS.n3813 VSS.n782 3.91226
R67429 VSS.n3809 VSS.n782 3.91226
R67430 VSS.n3809 VSS.n784 3.91226
R67431 VSS.n3801 VSS.n784 3.91226
R67432 VSS.n3801 VSS.n792 3.91226
R67433 VSS.n3796 VSS.n792 3.91226
R67434 VSS.n3796 VSS.n794 3.91226
R67435 VSS.n3787 VSS.n794 3.91226
R67436 VSS.n3787 VSS.n802 3.91226
R67437 VSS.n3783 VSS.n802 3.91226
R67438 VSS.n3783 VSS.n805 3.91226
R67439 VSS.n3775 VSS.n805 3.91226
R67440 VSS.n3775 VSS.n813 3.91226
R67441 VSS.n3771 VSS.n813 3.91226
R67442 VSS.n3771 VSS.n815 3.91226
R67443 VSS.n3763 VSS.n815 3.91226
R67444 VSS.n3763 VSS.n823 3.91226
R67445 VSS.n3759 VSS.n823 3.91226
R67446 VSS.n3759 VSS.n825 3.91226
R67447 VSS.n3751 VSS.n825 3.91226
R67448 VSS.n3751 VSS.n833 3.91226
R67449 VSS.n3747 VSS.n833 3.91226
R67450 VSS.n3747 VSS.n835 3.91226
R67451 VSS.n3739 VSS.n835 3.91226
R67452 VSS.n3739 VSS.n843 3.91226
R67453 VSS.n3735 VSS.n843 3.91226
R67454 VSS.n3735 VSS.n845 3.91226
R67455 VSS.n3102 VSS.n845 3.91226
R67456 VSS.n2682 VSS.n2071 3.91226
R67457 VSS.n2682 VSS.n2072 3.91226
R67458 VSS.n2221 VSS.n2072 3.91226
R67459 VSS.n2597 VSS.n2221 3.91226
R67460 VSS.n2597 VSS.n2558 3.91226
R67461 VSS.n2600 VSS.n2558 3.91226
R67462 VSS.n2600 VSS.n2563 3.91226
R67463 VSS.n2603 VSS.n2563 3.91226
R67464 VSS.n2603 VSS.n2568 3.91226
R67465 VSS.n2606 VSS.n2568 3.91226
R67466 VSS.n2606 VSS.n2573 3.91226
R67467 VSS.n2609 VSS.n2573 3.91226
R67468 VSS.n2609 VSS.n2578 3.91226
R67469 VSS.n2612 VSS.n2578 3.91226
R67470 VSS.n2612 VSS.n2583 3.91226
R67471 VSS.n2615 VSS.n2583 3.91226
R67472 VSS.n2615 VSS.n2588 3.91226
R67473 VSS.n2593 VSS.n2588 3.91226
R67474 VSS.n2621 VSS.n2593 3.91226
R67475 VSS.n2621 VSS.n2595 3.91226
R67476 VSS.n2595 VSS.n2594 3.91226
R67477 VSS.n2594 VSS.n671 3.91226
R67478 VSS.n3503 VSS.n671 3.91226
R67479 VSS.n3503 VSS.n678 3.91226
R67480 VSS.n3500 VSS.n678 3.91226
R67481 VSS.n3500 VSS.n683 3.91226
R67482 VSS.n3497 VSS.n683 3.91226
R67483 VSS.n3497 VSS.n688 3.91226
R67484 VSS.n3494 VSS.n688 3.91226
R67485 VSS.n3494 VSS.n693 3.91226
R67486 VSS.n3491 VSS.n693 3.91226
R67487 VSS.n3491 VSS.n697 3.91226
R67488 VSS.n3488 VSS.n697 3.91226
R67489 VSS.n3488 VSS.n702 3.91226
R67490 VSS.n3485 VSS.n702 3.91226
R67491 VSS.n3485 VSS.n708 3.91226
R67492 VSS.n3482 VSS.n708 3.91226
R67493 VSS.n3482 VSS.n713 3.91226
R67494 VSS.n3479 VSS.n713 3.91226
R67495 VSS.n3479 VSS.n718 3.91226
R67496 VSS.n3476 VSS.n718 3.91226
R67497 VSS.n3476 VSS.n723 3.91226
R67498 VSS.n3473 VSS.n723 3.91226
R67499 VSS.n3473 VSS.n3472 3.91226
R67500 VSS.n3472 VSS.n743 3.91226
R67501 VSS.n3468 VSS.n743 3.91226
R67502 VSS.n3468 VSS.n750 3.91226
R67503 VSS.n3465 VSS.n750 3.91226
R67504 VSS.n3465 VSS.n756 3.91226
R67505 VSS.n3462 VSS.n756 3.91226
R67506 VSS.n3462 VSS.n761 3.91226
R67507 VSS.n3459 VSS.n761 3.91226
R67508 VSS.n3459 VSS.n766 3.91226
R67509 VSS.n3456 VSS.n766 3.91226
R67510 VSS.n3456 VSS.n771 3.91226
R67511 VSS.n3453 VSS.n771 3.91226
R67512 VSS.n3453 VSS.n776 3.91226
R67513 VSS.n3450 VSS.n776 3.91226
R67514 VSS.n3450 VSS.n781 3.91226
R67515 VSS.n3447 VSS.n781 3.91226
R67516 VSS.n3447 VSS.n786 3.91226
R67517 VSS.n3444 VSS.n786 3.91226
R67518 VSS.n3444 VSS.n791 3.91226
R67519 VSS.n3441 VSS.n791 3.91226
R67520 VSS.n3441 VSS.n796 3.91226
R67521 VSS.n971 VSS.n796 3.91226
R67522 VSS.n971 VSS.n801 3.91226
R67523 VSS.n3070 VSS.n801 3.91226
R67524 VSS.n3070 VSS.n807 3.91226
R67525 VSS.n3073 VSS.n807 3.91226
R67526 VSS.n3073 VSS.n812 3.91226
R67527 VSS.n3076 VSS.n812 3.91226
R67528 VSS.n3076 VSS.n817 3.91226
R67529 VSS.n3079 VSS.n817 3.91226
R67530 VSS.n3079 VSS.n822 3.91226
R67531 VSS.n3082 VSS.n822 3.91226
R67532 VSS.n3082 VSS.n827 3.91226
R67533 VSS.n3085 VSS.n827 3.91226
R67534 VSS.n3085 VSS.n832 3.91226
R67535 VSS.n3088 VSS.n832 3.91226
R67536 VSS.n3088 VSS.n837 3.91226
R67537 VSS.n3091 VSS.n837 3.91226
R67538 VSS.n3091 VSS.n842 3.91226
R67539 VSS.n3094 VSS.n842 3.91226
R67540 VSS.n3094 VSS.n847 3.91226
R67541 VSS.n3099 VSS.n847 3.91226
R67542 VSS.n3398 VSS.n3099 3.91226
R67543 VSS.n2544 VSS.n2543 3.83228
R67544 VSS.n2545 VSS.n2544 3.83228
R67545 VSS.n4117 VSS.n4116 3.81164
R67546 VSS.n1883 VSS.n1882 3.70786
R67547 VSS.n1607 VSS.n1606 3.70786
R67548 VSS.n3390 VSS.n3104 3.39586
R67549 VSS.n3390 VSS.n3389 3.39586
R67550 VSS.n1614 VSS.n1613 3.1804
R67551 VSS.n4117 VSS.n569 3.14175
R67552 VSS.n3157 VSS.n3128 3.12476
R67553 VSS.n3130 VSS.n3128 3.12476
R67554 VSS.n1611 VSS.n1233 3.11878
R67555 VSS.n1614 VSS.n1606 3.11084
R67556 VSS.n1882 VSS.n1233 3.11084
R67557 VSS.n6194 VSS.n454 3.10905
R67558 VSS.n4101 VSS.n4100 3.10905
R67559 VSS.n3932 VSS.n452 2.99652
R67560 VSS.n4138 VSS.n4137 2.87501
R67561 VSS.n4143 VSS.n4142 2.87501
R67562 VSS.n4147 VSS.n4146 2.87501
R67563 VSS.n4152 VSS.n4151 2.87501
R67564 VSS.n4157 VSS.n4156 2.87501
R67565 VSS.n4161 VSS.n4160 2.87501
R67566 VSS.n4166 VSS.n4165 2.87501
R67567 VSS.n4171 VSS.n4170 2.87501
R67568 VSS.n4175 VSS.n4174 2.87501
R67569 VSS.n4193 VSS.n4192 2.87501
R67570 VSS.n4203 VSS.n4202 2.87501
R67571 VSS.n4207 VSS.n4206 2.87501
R67572 VSS.n532 VSS.n531 2.87501
R67573 VSS.n4219 VSS.n4218 2.87501
R67574 VSS.n4223 VSS.n4222 2.87501
R67575 VSS.n521 VSS.n520 2.87501
R67576 VSS.n4235 VSS.n4234 2.87501
R67577 VSS.n4242 VSS.n4241 2.87501
R67578 VSS.n4238 VSS.n4237 2.87501
R67579 VSS.n6135 VSS.n6134 2.87501
R67580 VSS.n4772 VSS.n4771 2.87501
R67581 VSS.n4780 VSS.n4779 2.87501
R67582 VSS.n4785 VSS.n4784 2.87501
R67583 VSS.n4789 VSS.n4788 2.87501
R67584 VSS.n4794 VSS.n4793 2.87501
R67585 VSS.n4855 VSS.n4854 2.87501
R67586 VSS.n4843 VSS.n4842 2.87501
R67587 VSS.n4831 VSS.n4830 2.87501
R67588 VSS.n4819 VSS.n4818 2.87501
R67589 VSS.n5989 VSS.n5988 2.87501
R67590 VSS.n5535 VSS.n5534 2.87501
R67591 VSS.n5517 VSS.n5516 2.87501
R67592 VSS.n5524 VSS.n5523 2.87501
R67593 VSS.n5638 VSS.n5637 2.87501
R67594 VSS.n5468 VSS.n5467 2.87501
R67595 VSS.n5848 VSS.n5847 2.87501
R67596 VSS.n5791 VSS.n5790 2.87501
R67597 VSS.n5098 VSS.n5097 2.87501
R67598 VSS.n5109 VSS.n5108 2.87501
R67599 VSS.n5808 VSS.n5807 2.87501
R67600 VSS.n4136 VSS.n459 2.81339
R67601 VSS.n4141 VSS.n460 2.81339
R67602 VSS.n550 VSS.n461 2.81339
R67603 VSS.n4150 VSS.n462 2.81339
R67604 VSS.n4155 VSS.n463 2.81339
R67605 VSS.n546 VSS.n464 2.81339
R67606 VSS.n4164 VSS.n465 2.81339
R67607 VSS.n4169 VSS.n466 2.81339
R67608 VSS.n542 VSS.n467 2.81339
R67609 VSS.n4191 VSS.n468 2.81339
R67610 VSS.n4201 VSS.n4200 2.81339
R67611 VSS.n4210 VSS.n4209 2.81339
R67612 VSS.n4213 VSS.n527 2.81339
R67613 VSS.n4217 VSS.n4216 2.81339
R67614 VSS.n4226 VSS.n4225 2.81339
R67615 VSS.n4229 VSS.n516 2.81339
R67616 VSS.n4233 VSS.n4232 2.81339
R67617 VSS.n4245 VSS.n4244 2.81339
R67618 VSS.n4248 VSS.n508 2.81339
R67619 VSS.n6133 VSS.n6132 2.81339
R67620 VSS.n4512 VSS.n4511 2.81339
R67621 VSS.n4778 VSS.n4275 2.81339
R67622 VSS.n4783 VSS.n4276 2.81339
R67623 VSS.n4485 VSS.n4277 2.81339
R67624 VSS.n4792 VSS.n4278 2.81339
R67625 VSS.n4853 VSS.n4852 2.81339
R67626 VSS.n4841 VSS.n4840 2.81339
R67627 VSS.n4829 VSS.n4828 2.81339
R67628 VSS.n4817 VSS.n4816 2.81339
R67629 VSS.n6101 VSS.n4308 2.81339
R67630 VSS.n5531 VSS.n5530 2.81339
R67631 VSS.n5513 VSS.n5512 2.81339
R67632 VSS.n5625 VSS.n5286 2.81339
R67633 VSS.n5636 VSS.n5635 2.81339
R67634 VSS.n5466 VSS.n5465 2.81339
R67635 VSS.n5846 VSS.n5845 2.81339
R67636 VSS.n5789 VSS.n5788 2.81339
R67637 VSS.n5102 VSS.n5100 2.81339
R67638 VSS.n5113 VSS.n5111 2.81339
R67639 VSS.n5117 VSS.n5050 2.81339
R67640 VSS.n3401 VSS.n864 2.69735
R67641 VSS.n3438 VSS.n894 2.69735
R67642 VSS.n3508 VSS.n3507 2.69735
R67643 VSS.n2685 VSS.n2068 2.69735
R67644 VSS.n3393 VSS.n3392 2.62838
R67645 VSS.n3132 VSS.n3131 2.62838
R67646 VSS.n3131 VSS.n3130 2.62235
R67647 VSS.n3389 VSS.n3386 2.61801
R67648 VSS.n3393 VSS.n3104 2.61724
R67649 VSS.n2538 VSS.n2537 2.6005
R67650 VSS.n2536 VSS.n2535 2.6005
R67651 VSS.n2534 VSS.n2533 2.6005
R67652 VSS.n2532 VSS.n2531 2.6005
R67653 VSS.n2530 VSS.n2529 2.6005
R67654 VSS.n2528 VSS.n2527 2.6005
R67655 VSS.n2526 VSS.n2525 2.6005
R67656 VSS.n2524 VSS.n2523 2.6005
R67657 VSS.n2522 VSS.n2521 2.6005
R67658 VSS.n2520 VSS.n2519 2.6005
R67659 VSS.n2518 VSS.n2517 2.6005
R67660 VSS.n2516 VSS.n2515 2.6005
R67661 VSS.n2514 VSS.n2513 2.6005
R67662 VSS.n2512 VSS.n2511 2.6005
R67663 VSS.n2510 VSS.n2509 2.6005
R67664 VSS.n2508 VSS.n2507 2.6005
R67665 VSS.n2506 VSS.n2505 2.6005
R67666 VSS.n2504 VSS.n2503 2.6005
R67667 VSS.n2502 VSS.n2501 2.6005
R67668 VSS.n2500 VSS.n2499 2.6005
R67669 VSS.n2498 VSS.n2497 2.6005
R67670 VSS.n2496 VSS.n2495 2.6005
R67671 VSS.n2494 VSS.n2493 2.6005
R67672 VSS.n2492 VSS.n2491 2.6005
R67673 VSS.n2490 VSS.n2489 2.6005
R67674 VSS.n2488 VSS.n2487 2.6005
R67675 VSS.n2486 VSS.n2485 2.6005
R67676 VSS.n2484 VSS.n2483 2.6005
R67677 VSS.n2482 VSS.n2481 2.6005
R67678 VSS.n2480 VSS.n2479 2.6005
R67679 VSS.n2478 VSS.n2477 2.6005
R67680 VSS.n2476 VSS.n2475 2.6005
R67681 VSS.n2474 VSS.n2473 2.6005
R67682 VSS.n2472 VSS.n2471 2.6005
R67683 VSS.n2470 VSS.n2469 2.6005
R67684 VSS.n2468 VSS.n2467 2.6005
R67685 VSS.n2466 VSS.n2465 2.6005
R67686 VSS.n2464 VSS.n2463 2.6005
R67687 VSS.n2462 VSS.n2461 2.6005
R67688 VSS.n2460 VSS.n2459 2.6005
R67689 VSS.n2458 VSS.n2457 2.6005
R67690 VSS.n2456 VSS.n2455 2.6005
R67691 VSS.n2454 VSS.n2453 2.6005
R67692 VSS.n2452 VSS.n2451 2.6005
R67693 VSS.n2450 VSS.n2449 2.6005
R67694 VSS.n2448 VSS.n2447 2.6005
R67695 VSS.n2446 VSS.n2445 2.6005
R67696 VSS.n2260 VSS.n2224 2.6005
R67697 VSS.n2414 VSS.n2225 2.6005
R67698 VSS.n2413 VSS.n2412 2.6005
R67699 VSS.n2411 VSS.n2410 2.6005
R67700 VSS.n2409 VSS.n2408 2.6005
R67701 VSS.n2407 VSS.n2406 2.6005
R67702 VSS.n2405 VSS.n2404 2.6005
R67703 VSS.n2403 VSS.n2402 2.6005
R67704 VSS.n2401 VSS.n2400 2.6005
R67705 VSS.n2399 VSS.n2398 2.6005
R67706 VSS.n2397 VSS.n2396 2.6005
R67707 VSS.n2395 VSS.n2394 2.6005
R67708 VSS.n2393 VSS.n2392 2.6005
R67709 VSS.n2391 VSS.n2390 2.6005
R67710 VSS.n2389 VSS.n2388 2.6005
R67711 VSS.n2387 VSS.n2386 2.6005
R67712 VSS.n2385 VSS.n2384 2.6005
R67713 VSS.n2383 VSS.n2382 2.6005
R67714 VSS.n2381 VSS.n2380 2.6005
R67715 VSS.n2379 VSS.n2378 2.6005
R67716 VSS.n2377 VSS.n2376 2.6005
R67717 VSS.n2375 VSS.n2374 2.6005
R67718 VSS.n2373 VSS.n2372 2.6005
R67719 VSS.n2371 VSS.n2370 2.6005
R67720 VSS.n2369 VSS.n2368 2.6005
R67721 VSS.n2367 VSS.n2366 2.6005
R67722 VSS.n2365 VSS.n2364 2.6005
R67723 VSS.n2363 VSS.n2362 2.6005
R67724 VSS.n2361 VSS.n2360 2.6005
R67725 VSS.n2359 VSS.n2358 2.6005
R67726 VSS.n2357 VSS.n2356 2.6005
R67727 VSS.n2355 VSS.n2354 2.6005
R67728 VSS.n2353 VSS.n2352 2.6005
R67729 VSS.n2351 VSS.n2350 2.6005
R67730 VSS.n2349 VSS.n2348 2.6005
R67731 VSS.n2347 VSS.n2346 2.6005
R67732 VSS.n2345 VSS.n2344 2.6005
R67733 VSS.n2343 VSS.n2342 2.6005
R67734 VSS.n2341 VSS.n2340 2.6005
R67735 VSS.n2339 VSS.n2338 2.6005
R67736 VSS.n2337 VSS.n2336 2.6005
R67737 VSS.n2335 VSS.n2334 2.6005
R67738 VSS.n2333 VSS.n2332 2.6005
R67739 VSS.n2331 VSS.n2330 2.6005
R67740 VSS.n2329 VSS.n2328 2.6005
R67741 VSS.n2327 VSS.n2326 2.6005
R67742 VSS.n2325 VSS.n2324 2.6005
R67743 VSS.n2323 VSS.n2322 2.6005
R67744 VSS.n2321 VSS.n2320 2.6005
R67745 VSS.n2319 VSS.n2318 2.6005
R67746 VSS.n3391 VSS.n3132 2.6005
R67747 VSS.n3100 VSS.n3098 2.6005
R67748 VSS.n3101 VSS.n3100 2.6005
R67749 VSS.n3399 VSS.n3398 2.6005
R67750 VSS.n3398 VSS.n3397 2.6005
R67751 VSS.n3099 VSS.n3097 2.6005
R67752 VSS.n3099 VSS.n846 2.6005
R67753 VSS.n3096 VSS.n847 2.6005
R67754 VSS.n3734 VSS.n847 2.6005
R67755 VSS.n3095 VSS.n3094 2.6005
R67756 VSS.n3094 VSS.n841 2.6005
R67757 VSS.n3093 VSS.n842 2.6005
R67758 VSS.n3740 VSS.n842 2.6005
R67759 VSS.n3092 VSS.n3091 2.6005
R67760 VSS.n3091 VSS.n836 2.6005
R67761 VSS.n3090 VSS.n837 2.6005
R67762 VSS.n3746 VSS.n837 2.6005
R67763 VSS.n3089 VSS.n3088 2.6005
R67764 VSS.n3088 VSS.n831 2.6005
R67765 VSS.n3087 VSS.n832 2.6005
R67766 VSS.n3752 VSS.n832 2.6005
R67767 VSS.n3086 VSS.n3085 2.6005
R67768 VSS.n3085 VSS.n826 2.6005
R67769 VSS.n3084 VSS.n827 2.6005
R67770 VSS.n3758 VSS.n827 2.6005
R67771 VSS.n3083 VSS.n3082 2.6005
R67772 VSS.n3082 VSS.n821 2.6005
R67773 VSS.n3081 VSS.n822 2.6005
R67774 VSS.n3764 VSS.n822 2.6005
R67775 VSS.n3080 VSS.n3079 2.6005
R67776 VSS.n3079 VSS.n816 2.6005
R67777 VSS.n3078 VSS.n817 2.6005
R67778 VSS.n3770 VSS.n817 2.6005
R67779 VSS.n3077 VSS.n3076 2.6005
R67780 VSS.n3076 VSS.n811 2.6005
R67781 VSS.n3075 VSS.n812 2.6005
R67782 VSS.n3776 VSS.n812 2.6005
R67783 VSS.n3074 VSS.n3073 2.6005
R67784 VSS.n3073 VSS.n806 2.6005
R67785 VSS.n3072 VSS.n807 2.6005
R67786 VSS.n3782 VSS.n807 2.6005
R67787 VSS.n3071 VSS.n3070 2.6005
R67788 VSS.n3070 VSS.n800 2.6005
R67789 VSS.n3069 VSS.n801 2.6005
R67790 VSS.n3788 VSS.n801 2.6005
R67791 VSS.n972 VSS.n971 2.6005
R67792 VSS.n971 VSS.n795 2.6005
R67793 VSS.n3440 VSS.n796 2.6005
R67794 VSS.n3795 VSS.n796 2.6005
R67795 VSS.n3442 VSS.n3441 2.6005
R67796 VSS.n3441 VSS.n790 2.6005
R67797 VSS.n3443 VSS.n791 2.6005
R67798 VSS.n3802 VSS.n791 2.6005
R67799 VSS.n3445 VSS.n3444 2.6005
R67800 VSS.n3444 VSS.n785 2.6005
R67801 VSS.n3446 VSS.n786 2.6005
R67802 VSS.n3808 VSS.n786 2.6005
R67803 VSS.n3448 VSS.n3447 2.6005
R67804 VSS.n3447 VSS.n780 2.6005
R67805 VSS.n3449 VSS.n781 2.6005
R67806 VSS.n3814 VSS.n781 2.6005
R67807 VSS.n3451 VSS.n3450 2.6005
R67808 VSS.n3450 VSS.n775 2.6005
R67809 VSS.n3452 VSS.n776 2.6005
R67810 VSS.n3820 VSS.n776 2.6005
R67811 VSS.n3454 VSS.n3453 2.6005
R67812 VSS.n3453 VSS.n770 2.6005
R67813 VSS.n3455 VSS.n771 2.6005
R67814 VSS.n3826 VSS.n771 2.6005
R67815 VSS.n3457 VSS.n3456 2.6005
R67816 VSS.n3456 VSS.n765 2.6005
R67817 VSS.n3458 VSS.n766 2.6005
R67818 VSS.n3832 VSS.n766 2.6005
R67819 VSS.n3460 VSS.n3459 2.6005
R67820 VSS.n3459 VSS.n760 2.6005
R67821 VSS.n3461 VSS.n761 2.6005
R67822 VSS.n3838 VSS.n761 2.6005
R67823 VSS.n3463 VSS.n3462 2.6005
R67824 VSS.n3462 VSS.n755 2.6005
R67825 VSS.n3464 VSS.n756 2.6005
R67826 VSS.n3844 VSS.n756 2.6005
R67827 VSS.n3466 VSS.n3465 2.6005
R67828 VSS.n3465 VSS.n749 2.6005
R67829 VSS.n3467 VSS.n750 2.6005
R67830 VSS.n3850 VSS.n750 2.6005
R67831 VSS.n3469 VSS.n3468 2.6005
R67832 VSS.n3468 VSS.n742 2.6005
R67833 VSS.n3470 VSS.n743 2.6005
R67834 VSS.n3856 VSS.n743 2.6005
R67835 VSS.n3472 VSS.n3471 2.6005
R67836 VSS.n3472 VSS.n741 2.6005
R67837 VSS.n3474 VSS.n3473 2.6005
R67838 VSS.n3473 VSS.n722 2.6005
R67839 VSS.n3475 VSS.n723 2.6005
R67840 VSS.n3866 VSS.n723 2.6005
R67841 VSS.n3477 VSS.n3476 2.6005
R67842 VSS.n3476 VSS.n717 2.6005
R67843 VSS.n3478 VSS.n718 2.6005
R67844 VSS.n3872 VSS.n718 2.6005
R67845 VSS.n3480 VSS.n3479 2.6005
R67846 VSS.n3479 VSS.n712 2.6005
R67847 VSS.n3481 VSS.n713 2.6005
R67848 VSS.n3878 VSS.n713 2.6005
R67849 VSS.n3483 VSS.n3482 2.6005
R67850 VSS.n3482 VSS.n707 2.6005
R67851 VSS.n3484 VSS.n708 2.6005
R67852 VSS.n3884 VSS.n708 2.6005
R67853 VSS.n3486 VSS.n3485 2.6005
R67854 VSS.n3485 VSS.n701 2.6005
R67855 VSS.n3487 VSS.n702 2.6005
R67856 VSS.n3890 VSS.n702 2.6005
R67857 VSS.n3489 VSS.n3488 2.6005
R67858 VSS.n3488 VSS.n696 2.6005
R67859 VSS.n3490 VSS.n697 2.6005
R67860 VSS.n3896 VSS.n697 2.6005
R67861 VSS.n3492 VSS.n3491 2.6005
R67862 VSS.n3491 VSS.n692 2.6005
R67863 VSS.n3493 VSS.n693 2.6005
R67864 VSS.n3902 VSS.n693 2.6005
R67865 VSS.n3495 VSS.n3494 2.6005
R67866 VSS.n3494 VSS.n687 2.6005
R67867 VSS.n3496 VSS.n688 2.6005
R67868 VSS.n3908 VSS.n688 2.6005
R67869 VSS.n3498 VSS.n3497 2.6005
R67870 VSS.n3497 VSS.n682 2.6005
R67871 VSS.n3499 VSS.n683 2.6005
R67872 VSS.n3914 VSS.n683 2.6005
R67873 VSS.n3501 VSS.n3500 2.6005
R67874 VSS.n3500 VSS.n677 2.6005
R67875 VSS.n3502 VSS.n678 2.6005
R67876 VSS.n3920 VSS.n678 2.6005
R67877 VSS.n3504 VSS.n3503 2.6005
R67878 VSS.n3503 VSS.n670 2.6005
R67879 VSS.n3505 VSS.n671 2.6005
R67880 VSS.n3927 VSS.n671 2.6005
R67881 VSS.n2594 VSS.n969 2.6005
R67882 VSS.n2594 VSS.n669 2.6005
R67883 VSS.n2619 VSS.n2595 2.6005
R67884 VSS.n2595 VSS.n2592 2.6005
R67885 VSS.n2621 VSS.n2620 2.6005
R67886 VSS.n2627 VSS.n2621 2.6005
R67887 VSS.n2618 VSS.n2593 2.6005
R67888 VSS.n2593 VSS.n2587 2.6005
R67889 VSS.n2617 VSS.n2588 2.6005
R67890 VSS.n2633 VSS.n2588 2.6005
R67891 VSS.n2616 VSS.n2615 2.6005
R67892 VSS.n2615 VSS.n2582 2.6005
R67893 VSS.n2614 VSS.n2583 2.6005
R67894 VSS.n2639 VSS.n2583 2.6005
R67895 VSS.n2613 VSS.n2612 2.6005
R67896 VSS.n2612 VSS.n2577 2.6005
R67897 VSS.n2611 VSS.n2578 2.6005
R67898 VSS.n2645 VSS.n2578 2.6005
R67899 VSS.n2610 VSS.n2609 2.6005
R67900 VSS.n2609 VSS.n2572 2.6005
R67901 VSS.n2608 VSS.n2573 2.6005
R67902 VSS.n2651 VSS.n2573 2.6005
R67903 VSS.n2607 VSS.n2606 2.6005
R67904 VSS.n2606 VSS.n2567 2.6005
R67905 VSS.n2605 VSS.n2568 2.6005
R67906 VSS.n2657 VSS.n2568 2.6005
R67907 VSS.n2604 VSS.n2603 2.6005
R67908 VSS.n2603 VSS.n2562 2.6005
R67909 VSS.n2602 VSS.n2563 2.6005
R67910 VSS.n2663 VSS.n2563 2.6005
R67911 VSS.n2601 VSS.n2600 2.6005
R67912 VSS.n2600 VSS.n2557 2.6005
R67913 VSS.n2599 VSS.n2558 2.6005
R67914 VSS.n2669 VSS.n2558 2.6005
R67915 VSS.n2598 VSS.n2597 2.6005
R67916 VSS.n2597 VSS.n2220 2.6005
R67917 VSS.n2596 VSS.n2221 2.6005
R67918 VSS.n2675 VSS.n2221 2.6005
R67919 VSS.n2072 VSS.n2070 2.6005
R67920 VSS.n2074 VSS.n2072 2.6005
R67921 VSS.n2683 VSS.n2682 2.6005
R67922 VSS.n2682 VSS.n2681 2.6005
R67923 VSS.n2071 VSS.n2069 2.6005
R67924 VSS.n2073 VSS.n2071 2.6005
R67925 VSS.n3161 VSS.n3160 2.6005
R67926 VSS.n3164 VSS.n3163 2.6005
R67927 VSS.n3166 VSS.n3165 2.6005
R67928 VSS.n3169 VSS.n3168 2.6005
R67929 VSS.n3171 VSS.n3170 2.6005
R67930 VSS.n3174 VSS.n3173 2.6005
R67931 VSS.n3176 VSS.n3175 2.6005
R67932 VSS.n3179 VSS.n3178 2.6005
R67933 VSS.n3181 VSS.n3180 2.6005
R67934 VSS.n3184 VSS.n3183 2.6005
R67935 VSS.n3186 VSS.n3185 2.6005
R67936 VSS.n3189 VSS.n3188 2.6005
R67937 VSS.n3191 VSS.n3190 2.6005
R67938 VSS.n3194 VSS.n3193 2.6005
R67939 VSS.n3196 VSS.n3195 2.6005
R67940 VSS.n3199 VSS.n3198 2.6005
R67941 VSS.n3201 VSS.n3200 2.6005
R67942 VSS.n3204 VSS.n3203 2.6005
R67943 VSS.n3206 VSS.n3205 2.6005
R67944 VSS.n3209 VSS.n3208 2.6005
R67945 VSS.n3211 VSS.n3210 2.6005
R67946 VSS.n3214 VSS.n3213 2.6005
R67947 VSS.n3216 VSS.n3215 2.6005
R67948 VSS.n3219 VSS.n3218 2.6005
R67949 VSS.n3221 VSS.n3220 2.6005
R67950 VSS.n3224 VSS.n3223 2.6005
R67951 VSS.n3226 VSS.n3225 2.6005
R67952 VSS.n3229 VSS.n3228 2.6005
R67953 VSS.n3231 VSS.n3230 2.6005
R67954 VSS.n3234 VSS.n3233 2.6005
R67955 VSS.n3236 VSS.n3235 2.6005
R67956 VSS.n3239 VSS.n3238 2.6005
R67957 VSS.n3241 VSS.n3240 2.6005
R67958 VSS.n3244 VSS.n3243 2.6005
R67959 VSS.n3246 VSS.n3245 2.6005
R67960 VSS.n3249 VSS.n3248 2.6005
R67961 VSS.n3251 VSS.n3250 2.6005
R67962 VSS.n3254 VSS.n3253 2.6005
R67963 VSS.n3256 VSS.n3255 2.6005
R67964 VSS.n3259 VSS.n3258 2.6005
R67965 VSS.n3261 VSS.n3260 2.6005
R67966 VSS.n3264 VSS.n3263 2.6005
R67967 VSS.n3266 VSS.n3102 2.6005
R67968 VSS.n3397 VSS.n3102 2.6005
R67969 VSS.n845 VSS.n844 2.6005
R67970 VSS.n846 VSS.n845 2.6005
R67971 VSS.n3736 VSS.n3735 2.6005
R67972 VSS.n3735 VSS.n3734 2.6005
R67973 VSS.n3737 VSS.n843 2.6005
R67974 VSS.n843 VSS.n841 2.6005
R67975 VSS.n3739 VSS.n3738 2.6005
R67976 VSS.n3740 VSS.n3739 2.6005
R67977 VSS.n835 VSS.n834 2.6005
R67978 VSS.n836 VSS.n835 2.6005
R67979 VSS.n3748 VSS.n3747 2.6005
R67980 VSS.n3747 VSS.n3746 2.6005
R67981 VSS.n3749 VSS.n833 2.6005
R67982 VSS.n833 VSS.n831 2.6005
R67983 VSS.n3751 VSS.n3750 2.6005
R67984 VSS.n3752 VSS.n3751 2.6005
R67985 VSS.n825 VSS.n824 2.6005
R67986 VSS.n826 VSS.n825 2.6005
R67987 VSS.n3760 VSS.n3759 2.6005
R67988 VSS.n3759 VSS.n3758 2.6005
R67989 VSS.n3761 VSS.n823 2.6005
R67990 VSS.n823 VSS.n821 2.6005
R67991 VSS.n3763 VSS.n3762 2.6005
R67992 VSS.n3764 VSS.n3763 2.6005
R67993 VSS.n815 VSS.n814 2.6005
R67994 VSS.n816 VSS.n815 2.6005
R67995 VSS.n3772 VSS.n3771 2.6005
R67996 VSS.n3771 VSS.n3770 2.6005
R67997 VSS.n3773 VSS.n813 2.6005
R67998 VSS.n813 VSS.n811 2.6005
R67999 VSS.n3775 VSS.n3774 2.6005
R68000 VSS.n3776 VSS.n3775 2.6005
R68001 VSS.n805 VSS.n804 2.6005
R68002 VSS.n806 VSS.n805 2.6005
R68003 VSS.n3784 VSS.n3783 2.6005
R68004 VSS.n3783 VSS.n3782 2.6005
R68005 VSS.n3785 VSS.n802 2.6005
R68006 VSS.n802 VSS.n800 2.6005
R68007 VSS.n3787 VSS.n3786 2.6005
R68008 VSS.n3788 VSS.n3787 2.6005
R68009 VSS.n803 VSS.n794 2.6005
R68010 VSS.n795 VSS.n794 2.6005
R68011 VSS.n3797 VSS.n3796 2.6005
R68012 VSS.n3796 VSS.n3795 2.6005
R68013 VSS.n3799 VSS.n792 2.6005
R68014 VSS.n792 VSS.n790 2.6005
R68015 VSS.n3801 VSS.n3800 2.6005
R68016 VSS.n3802 VSS.n3801 2.6005
R68017 VSS.n784 VSS.n783 2.6005
R68018 VSS.n785 VSS.n784 2.6005
R68019 VSS.n3810 VSS.n3809 2.6005
R68020 VSS.n3809 VSS.n3808 2.6005
R68021 VSS.n3811 VSS.n782 2.6005
R68022 VSS.n782 VSS.n780 2.6005
R68023 VSS.n3813 VSS.n3812 2.6005
R68024 VSS.n3814 VSS.n3813 2.6005
R68025 VSS.n774 VSS.n773 2.6005
R68026 VSS.n775 VSS.n774 2.6005
R68027 VSS.n3822 VSS.n3821 2.6005
R68028 VSS.n3821 VSS.n3820 2.6005
R68029 VSS.n3823 VSS.n772 2.6005
R68030 VSS.n772 VSS.n770 2.6005
R68031 VSS.n3825 VSS.n3824 2.6005
R68032 VSS.n3826 VSS.n3825 2.6005
R68033 VSS.n764 VSS.n763 2.6005
R68034 VSS.n765 VSS.n764 2.6005
R68035 VSS.n3834 VSS.n3833 2.6005
R68036 VSS.n3833 VSS.n3832 2.6005
R68037 VSS.n3835 VSS.n762 2.6005
R68038 VSS.n762 VSS.n760 2.6005
R68039 VSS.n3837 VSS.n3836 2.6005
R68040 VSS.n3838 VSS.n3837 2.6005
R68041 VSS.n754 VSS.n753 2.6005
R68042 VSS.n755 VSS.n754 2.6005
R68043 VSS.n3846 VSS.n3845 2.6005
R68044 VSS.n3845 VSS.n3844 2.6005
R68045 VSS.n3847 VSS.n751 2.6005
R68046 VSS.n751 VSS.n749 2.6005
R68047 VSS.n3849 VSS.n3848 2.6005
R68048 VSS.n3850 VSS.n3849 2.6005
R68049 VSS.n752 VSS.n740 2.6005
R68050 VSS.n742 VSS.n740 2.6005
R68051 VSS.n3858 VSS.n3857 2.6005
R68052 VSS.n3857 VSS.n3856 2.6005
R68053 VSS.n739 VSS.n734 2.6005
R68054 VSS.n741 VSS.n739 2.6005
R68055 VSS.n727 VSS.n724 2.6005
R68056 VSS.n724 VSS.n722 2.6005
R68057 VSS.n3865 VSS.n3864 2.6005
R68058 VSS.n3866 VSS.n3865 2.6005
R68059 VSS.n716 VSS.n715 2.6005
R68060 VSS.n717 VSS.n716 2.6005
R68061 VSS.n3874 VSS.n3873 2.6005
R68062 VSS.n3873 VSS.n3872 2.6005
R68063 VSS.n3875 VSS.n714 2.6005
R68064 VSS.n714 VSS.n712 2.6005
R68065 VSS.n3877 VSS.n3876 2.6005
R68066 VSS.n3878 VSS.n3877 2.6005
R68067 VSS.n706 VSS.n705 2.6005
R68068 VSS.n707 VSS.n706 2.6005
R68069 VSS.n3886 VSS.n3885 2.6005
R68070 VSS.n3885 VSS.n3884 2.6005
R68071 VSS.n3887 VSS.n703 2.6005
R68072 VSS.n703 VSS.n701 2.6005
R68073 VSS.n3889 VSS.n3888 2.6005
R68074 VSS.n3890 VSS.n3889 2.6005
R68075 VSS.n704 VSS.n695 2.6005
R68076 VSS.n696 VSS.n695 2.6005
R68077 VSS.n3898 VSS.n3897 2.6005
R68078 VSS.n3897 VSS.n3896 2.6005
R68079 VSS.n3899 VSS.n694 2.6005
R68080 VSS.n694 VSS.n692 2.6005
R68081 VSS.n3901 VSS.n3900 2.6005
R68082 VSS.n3902 VSS.n3901 2.6005
R68083 VSS.n686 VSS.n685 2.6005
R68084 VSS.n687 VSS.n686 2.6005
R68085 VSS.n3910 VSS.n3909 2.6005
R68086 VSS.n3909 VSS.n3908 2.6005
R68087 VSS.n3911 VSS.n684 2.6005
R68088 VSS.n684 VSS.n682 2.6005
R68089 VSS.n3913 VSS.n3912 2.6005
R68090 VSS.n3914 VSS.n3913 2.6005
R68091 VSS.n676 VSS.n675 2.6005
R68092 VSS.n677 VSS.n676 2.6005
R68093 VSS.n3922 VSS.n3921 2.6005
R68094 VSS.n3921 VSS.n3920 2.6005
R68095 VSS.n3923 VSS.n673 2.6005
R68096 VSS.n673 VSS.n670 2.6005
R68097 VSS.n3926 VSS.n3925 2.6005
R68098 VSS.n3927 VSS.n3926 2.6005
R68099 VSS.n2623 VSS.n672 2.6005
R68100 VSS.n672 VSS.n669 2.6005
R68101 VSS.n2624 VSS.n2622 2.6005
R68102 VSS.n2622 VSS.n2592 2.6005
R68103 VSS.n2626 VSS.n2625 2.6005
R68104 VSS.n2627 VSS.n2626 2.6005
R68105 VSS.n2586 VSS.n2585 2.6005
R68106 VSS.n2587 VSS.n2586 2.6005
R68107 VSS.n2635 VSS.n2634 2.6005
R68108 VSS.n2634 VSS.n2633 2.6005
R68109 VSS.n2636 VSS.n2584 2.6005
R68110 VSS.n2584 VSS.n2582 2.6005
R68111 VSS.n2638 VSS.n2637 2.6005
R68112 VSS.n2639 VSS.n2638 2.6005
R68113 VSS.n2576 VSS.n2575 2.6005
R68114 VSS.n2577 VSS.n2576 2.6005
R68115 VSS.n2647 VSS.n2646 2.6005
R68116 VSS.n2646 VSS.n2645 2.6005
R68117 VSS.n2648 VSS.n2574 2.6005
R68118 VSS.n2574 VSS.n2572 2.6005
R68119 VSS.n2650 VSS.n2649 2.6005
R68120 VSS.n2651 VSS.n2650 2.6005
R68121 VSS.n2566 VSS.n2565 2.6005
R68122 VSS.n2567 VSS.n2566 2.6005
R68123 VSS.n2659 VSS.n2658 2.6005
R68124 VSS.n2658 VSS.n2657 2.6005
R68125 VSS.n2660 VSS.n2564 2.6005
R68126 VSS.n2564 VSS.n2562 2.6005
R68127 VSS.n2662 VSS.n2661 2.6005
R68128 VSS.n2663 VSS.n2662 2.6005
R68129 VSS.n2556 VSS.n2555 2.6005
R68130 VSS.n2557 VSS.n2556 2.6005
R68131 VSS.n2671 VSS.n2670 2.6005
R68132 VSS.n2670 VSS.n2669 2.6005
R68133 VSS.n2672 VSS.n2223 2.6005
R68134 VSS.n2223 VSS.n2220 2.6005
R68135 VSS.n2674 VSS.n2673 2.6005
R68136 VSS.n2675 VSS.n2674 2.6005
R68137 VSS.n2554 VSS.n2222 2.6005
R68138 VSS.n2222 VSS.n2074 2.6005
R68139 VSS.n2553 VSS.n2075 2.6005
R68140 VSS.n2681 VSS.n2075 2.6005
R68141 VSS.n2551 VSS.n2550 2.6005
R68142 VSS.n2550 VSS.n2073 2.6005
R68143 VSS.n3282 VSS.n3281 2.6005
R68144 VSS.n3285 VSS.n3284 2.6005
R68145 VSS.n3287 VSS.n3286 2.6005
R68146 VSS.n3290 VSS.n3289 2.6005
R68147 VSS.n3292 VSS.n3291 2.6005
R68148 VSS.n3295 VSS.n3294 2.6005
R68149 VSS.n3297 VSS.n3296 2.6005
R68150 VSS.n3300 VSS.n3299 2.6005
R68151 VSS.n3302 VSS.n3301 2.6005
R68152 VSS.n3305 VSS.n3304 2.6005
R68153 VSS.n3307 VSS.n3306 2.6005
R68154 VSS.n3310 VSS.n3309 2.6005
R68155 VSS.n3312 VSS.n3311 2.6005
R68156 VSS.n3315 VSS.n3314 2.6005
R68157 VSS.n3317 VSS.n3316 2.6005
R68158 VSS.n3320 VSS.n3319 2.6005
R68159 VSS.n3322 VSS.n3321 2.6005
R68160 VSS.n3325 VSS.n3324 2.6005
R68161 VSS.n3327 VSS.n3326 2.6005
R68162 VSS.n3330 VSS.n3329 2.6005
R68163 VSS.n3332 VSS.n3331 2.6005
R68164 VSS.n3335 VSS.n3334 2.6005
R68165 VSS.n3337 VSS.n3336 2.6005
R68166 VSS.n3340 VSS.n3339 2.6005
R68167 VSS.n3342 VSS.n3341 2.6005
R68168 VSS.n3345 VSS.n3344 2.6005
R68169 VSS.n3347 VSS.n3346 2.6005
R68170 VSS.n3350 VSS.n3349 2.6005
R68171 VSS.n3352 VSS.n3351 2.6005
R68172 VSS.n3355 VSS.n3354 2.6005
R68173 VSS.n3357 VSS.n3356 2.6005
R68174 VSS.n3360 VSS.n3359 2.6005
R68175 VSS.n3362 VSS.n3361 2.6005
R68176 VSS.n3365 VSS.n3364 2.6005
R68177 VSS.n3367 VSS.n3366 2.6005
R68178 VSS.n3370 VSS.n3369 2.6005
R68179 VSS.n3372 VSS.n3371 2.6005
R68180 VSS.n3375 VSS.n3374 2.6005
R68181 VSS.n3377 VSS.n3376 2.6005
R68182 VSS.n3380 VSS.n3379 2.6005
R68183 VSS.n3382 VSS.n3381 2.6005
R68184 VSS.n3385 VSS.n3384 2.6005
R68185 VSS.n3387 VSS.n3386 2.6005
R68186 VSS.n3392 VSS.n3391 2.6005
R68187 VSS.n3395 VSS.n3394 2.6005
R68188 VSS.n3395 VSS.n3101 2.6005
R68189 VSS.n3396 VSS.n849 2.6005
R68190 VSS.n3397 VSS.n3396 2.6005
R68191 VSS.n3731 VSS.n848 2.6005
R68192 VSS.n848 VSS.n846 2.6005
R68193 VSS.n3733 VSS.n3732 2.6005
R68194 VSS.n3734 VSS.n3733 2.6005
R68195 VSS.n840 VSS.n839 2.6005
R68196 VSS.n841 VSS.n840 2.6005
R68197 VSS.n3742 VSS.n3741 2.6005
R68198 VSS.n3741 VSS.n3740 2.6005
R68199 VSS.n3743 VSS.n838 2.6005
R68200 VSS.n838 VSS.n836 2.6005
R68201 VSS.n3745 VSS.n3744 2.6005
R68202 VSS.n3746 VSS.n3745 2.6005
R68203 VSS.n830 VSS.n829 2.6005
R68204 VSS.n831 VSS.n830 2.6005
R68205 VSS.n3754 VSS.n3753 2.6005
R68206 VSS.n3753 VSS.n3752 2.6005
R68207 VSS.n3755 VSS.n828 2.6005
R68208 VSS.n828 VSS.n826 2.6005
R68209 VSS.n3757 VSS.n3756 2.6005
R68210 VSS.n3758 VSS.n3757 2.6005
R68211 VSS.n820 VSS.n819 2.6005
R68212 VSS.n821 VSS.n820 2.6005
R68213 VSS.n3766 VSS.n3765 2.6005
R68214 VSS.n3765 VSS.n3764 2.6005
R68215 VSS.n3767 VSS.n818 2.6005
R68216 VSS.n818 VSS.n816 2.6005
R68217 VSS.n3769 VSS.n3768 2.6005
R68218 VSS.n3770 VSS.n3769 2.6005
R68219 VSS.n810 VSS.n809 2.6005
R68220 VSS.n811 VSS.n810 2.6005
R68221 VSS.n3778 VSS.n3777 2.6005
R68222 VSS.n3777 VSS.n3776 2.6005
R68223 VSS.n3779 VSS.n808 2.6005
R68224 VSS.n808 VSS.n806 2.6005
R68225 VSS.n3781 VSS.n3780 2.6005
R68226 VSS.n3782 VSS.n3781 2.6005
R68227 VSS.n799 VSS.n798 2.6005
R68228 VSS.n800 VSS.n799 2.6005
R68229 VSS.n3790 VSS.n3789 2.6005
R68230 VSS.n3789 VSS.n3788 2.6005
R68231 VSS.n3791 VSS.n797 2.6005
R68232 VSS.n797 VSS.n795 2.6005
R68233 VSS.n3794 VSS.n3793 2.6005
R68234 VSS.n3795 VSS.n3794 2.6005
R68235 VSS.n789 VSS.n788 2.6005
R68236 VSS.n790 VSS.n789 2.6005
R68237 VSS.n3804 VSS.n3803 2.6005
R68238 VSS.n3803 VSS.n3802 2.6005
R68239 VSS.n3805 VSS.n787 2.6005
R68240 VSS.n787 VSS.n785 2.6005
R68241 VSS.n3807 VSS.n3806 2.6005
R68242 VSS.n3808 VSS.n3807 2.6005
R68243 VSS.n779 VSS.n778 2.6005
R68244 VSS.n780 VSS.n779 2.6005
R68245 VSS.n3816 VSS.n3815 2.6005
R68246 VSS.n3815 VSS.n3814 2.6005
R68247 VSS.n3817 VSS.n777 2.6005
R68248 VSS.n777 VSS.n775 2.6005
R68249 VSS.n3819 VSS.n3818 2.6005
R68250 VSS.n3820 VSS.n3819 2.6005
R68251 VSS.n769 VSS.n768 2.6005
R68252 VSS.n770 VSS.n769 2.6005
R68253 VSS.n3828 VSS.n3827 2.6005
R68254 VSS.n3827 VSS.n3826 2.6005
R68255 VSS.n3829 VSS.n767 2.6005
R68256 VSS.n767 VSS.n765 2.6005
R68257 VSS.n3831 VSS.n3830 2.6005
R68258 VSS.n3832 VSS.n3831 2.6005
R68259 VSS.n759 VSS.n758 2.6005
R68260 VSS.n760 VSS.n759 2.6005
R68261 VSS.n3840 VSS.n3839 2.6005
R68262 VSS.n3839 VSS.n3838 2.6005
R68263 VSS.n3841 VSS.n757 2.6005
R68264 VSS.n757 VSS.n755 2.6005
R68265 VSS.n3843 VSS.n3842 2.6005
R68266 VSS.n3844 VSS.n3843 2.6005
R68267 VSS.n748 VSS.n747 2.6005
R68268 VSS.n749 VSS.n748 2.6005
R68269 VSS.n3852 VSS.n3851 2.6005
R68270 VSS.n3851 VSS.n3850 2.6005
R68271 VSS.n3853 VSS.n745 2.6005
R68272 VSS.n745 VSS.n742 2.6005
R68273 VSS.n3855 VSS.n3854 2.6005
R68274 VSS.n3856 VSS.n3855 2.6005
R68275 VSS.n746 VSS.n744 2.6005
R68276 VSS.n744 VSS.n741 2.6005
R68277 VSS.n721 VSS.n720 2.6005
R68278 VSS.n722 VSS.n721 2.6005
R68279 VSS.n3868 VSS.n3867 2.6005
R68280 VSS.n3867 VSS.n3866 2.6005
R68281 VSS.n3869 VSS.n719 2.6005
R68282 VSS.n719 VSS.n717 2.6005
R68283 VSS.n3871 VSS.n3870 2.6005
R68284 VSS.n3872 VSS.n3871 2.6005
R68285 VSS.n711 VSS.n710 2.6005
R68286 VSS.n712 VSS.n711 2.6005
R68287 VSS.n3880 VSS.n3879 2.6005
R68288 VSS.n3879 VSS.n3878 2.6005
R68289 VSS.n3881 VSS.n709 2.6005
R68290 VSS.n709 VSS.n707 2.6005
R68291 VSS.n3883 VSS.n3882 2.6005
R68292 VSS.n3884 VSS.n3883 2.6005
R68293 VSS.n700 VSS.n699 2.6005
R68294 VSS.n701 VSS.n700 2.6005
R68295 VSS.n3892 VSS.n3891 2.6005
R68296 VSS.n3891 VSS.n3890 2.6005
R68297 VSS.n3893 VSS.n698 2.6005
R68298 VSS.n698 VSS.n696 2.6005
R68299 VSS.n3895 VSS.n3894 2.6005
R68300 VSS.n3896 VSS.n3895 2.6005
R68301 VSS.n691 VSS.n690 2.6005
R68302 VSS.n692 VSS.n691 2.6005
R68303 VSS.n3904 VSS.n3903 2.6005
R68304 VSS.n3903 VSS.n3902 2.6005
R68305 VSS.n3905 VSS.n689 2.6005
R68306 VSS.n689 VSS.n687 2.6005
R68307 VSS.n3907 VSS.n3906 2.6005
R68308 VSS.n3908 VSS.n3907 2.6005
R68309 VSS.n681 VSS.n680 2.6005
R68310 VSS.n682 VSS.n681 2.6005
R68311 VSS.n3916 VSS.n3915 2.6005
R68312 VSS.n3915 VSS.n3914 2.6005
R68313 VSS.n3917 VSS.n679 2.6005
R68314 VSS.n679 VSS.n677 2.6005
R68315 VSS.n3919 VSS.n3918 2.6005
R68316 VSS.n3920 VSS.n3919 2.6005
R68317 VSS.n668 VSS.n666 2.6005
R68318 VSS.n670 VSS.n668 2.6005
R68319 VSS.n3929 VSS.n3928 2.6005
R68320 VSS.n3928 VSS.n3927 2.6005
R68321 VSS.n667 VSS.n665 2.6005
R68322 VSS.n669 VSS.n667 2.6005
R68323 VSS.n2591 VSS.n2590 2.6005
R68324 VSS.n2592 VSS.n2591 2.6005
R68325 VSS.n2629 VSS.n2628 2.6005
R68326 VSS.n2628 VSS.n2627 2.6005
R68327 VSS.n2630 VSS.n2589 2.6005
R68328 VSS.n2589 VSS.n2587 2.6005
R68329 VSS.n2632 VSS.n2631 2.6005
R68330 VSS.n2633 VSS.n2632 2.6005
R68331 VSS.n2581 VSS.n2580 2.6005
R68332 VSS.n2582 VSS.n2581 2.6005
R68333 VSS.n2641 VSS.n2640 2.6005
R68334 VSS.n2640 VSS.n2639 2.6005
R68335 VSS.n2642 VSS.n2579 2.6005
R68336 VSS.n2579 VSS.n2577 2.6005
R68337 VSS.n2644 VSS.n2643 2.6005
R68338 VSS.n2645 VSS.n2644 2.6005
R68339 VSS.n2571 VSS.n2570 2.6005
R68340 VSS.n2572 VSS.n2571 2.6005
R68341 VSS.n2653 VSS.n2652 2.6005
R68342 VSS.n2652 VSS.n2651 2.6005
R68343 VSS.n2654 VSS.n2569 2.6005
R68344 VSS.n2569 VSS.n2567 2.6005
R68345 VSS.n2656 VSS.n2655 2.6005
R68346 VSS.n2657 VSS.n2656 2.6005
R68347 VSS.n2561 VSS.n2560 2.6005
R68348 VSS.n2562 VSS.n2561 2.6005
R68349 VSS.n2665 VSS.n2664 2.6005
R68350 VSS.n2664 VSS.n2663 2.6005
R68351 VSS.n2666 VSS.n2559 2.6005
R68352 VSS.n2559 VSS.n2557 2.6005
R68353 VSS.n2668 VSS.n2667 2.6005
R68354 VSS.n2669 VSS.n2668 2.6005
R68355 VSS.n2219 VSS.n2218 2.6005
R68356 VSS.n2220 VSS.n2219 2.6005
R68357 VSS.n2677 VSS.n2676 2.6005
R68358 VSS.n2676 VSS.n2675 2.6005
R68359 VSS.n2678 VSS.n2077 2.6005
R68360 VSS.n2077 VSS.n2074 2.6005
R68361 VSS.n2680 VSS.n2679 2.6005
R68362 VSS.n2681 VSS.n2680 2.6005
R68363 VSS.n2314 VSS.n2076 2.6005
R68364 VSS.n2076 VSS.n2073 2.6005
R68365 VSS.n2416 VSS.n2226 2.5974
R68366 VSS.n3272 VSS.n3271 2.5974
R68367 VSS.n3104 VSS.n3103 2.36815
R68368 VSS.n3130 VSS.n3129 2.36815
R68369 VSS.n5868 VSS.n5867 2.25175
R68370 VSS.n5804 VSS.n5803 2.25175
R68371 VSS.n5784 VSS.n5783 2.25175
R68372 VSS.n5840 VSS.n4983 2.25175
R68373 VSS.n5867 VSS.n4943 2.251
R68374 VSS.n5803 VSS.n5797 2.251
R68375 VSS.n5783 VSS.n5781 2.251
R68376 VSS.n5842 VSS.n4983 2.251
R68377 VSS.n4103 VSS.n4102 2.2505
R68378 VSS.n6192 VSS.n6191 2.2505
R68379 VSS.n4424 VSS.n4396 2.25007
R68380 VSS.n3588 VSS.n732 2.25007
R68381 VSS.n5537 VSS.n5461 2.25007
R68382 VSS.n5094 VSS.n5093 2.25007
R68383 VSS.n3978 VSS.n3977 2.24901
R68384 VSS.n2823 VSS.n2822 2.24901
R68385 VSS.n4502 VSS.n483 2.24901
R68386 VSS.n2968 VSS.n1105 2.24901
R68387 VSS.n1491 VSS.n1224 2.24901
R68388 VSS.n1660 VSS.n1307 2.24882
R68389 VSS.n556 VSS.n553 2.24648
R68390 VSS.n4129 VSS.n4128 2.24648
R68391 VSS.n5483 VSS.n5480 2.24648
R68392 VSS.n4180 VSS.n4177 2.24648
R68393 VSS.n2891 VSS.n2887 2.24581
R68394 VSS.n2902 VSS.n2884 2.24581
R68395 VSS.n1143 VSS.n1141 2.24581
R68396 VSS.n2886 VSS.n1151 2.24581
R68397 VSS.n2890 VSS.n1154 2.24581
R68398 VSS.n4420 VSS.n4417 2.24581
R68399 VSS.n4423 VSS.n4381 2.24581
R68400 VSS.n4420 VSS.n4418 2.24581
R68401 VSS.n4400 VSS.n4381 2.24581
R68402 VSS.n4420 VSS.n4416 2.24581
R68403 VSS.n4402 VSS.n4381 2.24581
R68404 VSS.n4420 VSS.n4419 2.24581
R68405 VSS.n4405 VSS.n4381 2.24581
R68406 VSS.n4420 VSS.n4415 2.24581
R68407 VSS.n4506 VSS.n4487 2.24581
R68408 VSS.n4506 VSS.n4503 2.24581
R68409 VSS.n4498 VSS.n4488 2.24581
R68410 VSS.n4506 VSS.n4504 2.24581
R68411 VSS.n4492 VSS.n4488 2.24581
R68412 VSS.n4506 VSS.n4505 2.24581
R68413 VSS.n627 VSS.n622 2.24581
R68414 VSS.n3974 VSS.n3973 2.24581
R68415 VSS.n629 VSS.n622 2.24581
R68416 VSS.n3974 VSS.n3972 2.24581
R68417 VSS.n631 VSS.n622 2.24581
R68418 VSS.n3974 VSS.n3971 2.24581
R68419 VSS.n633 VSS.n622 2.24581
R68420 VSS.n3974 VSS.n3970 2.24581
R68421 VSS.n635 VSS.n622 2.24581
R68422 VSS.n3974 VSS.n637 2.24581
R68423 VSS.n3587 VSS.n3586 2.24581
R68424 VSS.n947 VSS.n937 2.24581
R68425 VSS.n3587 VSS.n3585 2.24581
R68426 VSS.n947 VSS.n938 2.24581
R68427 VSS.n3587 VSS.n3584 2.24581
R68428 VSS.n947 VSS.n939 2.24581
R68429 VSS.n3587 VSS.n3583 2.24581
R68430 VSS.n947 VSS.n940 2.24581
R68431 VSS.n3587 VSS.n3582 2.24581
R68432 VSS.n947 VSS.n941 2.24581
R68433 VSS.n3587 VSS.n3581 2.24581
R68434 VSS.n947 VSS.n942 2.24581
R68435 VSS.n3587 VSS.n3580 2.24581
R68436 VSS.n947 VSS.n943 2.24581
R68437 VSS.n3587 VSS.n3579 2.24581
R68438 VSS.n947 VSS.n944 2.24581
R68439 VSS.n3587 VSS.n3578 2.24581
R68440 VSS.n947 VSS.n945 2.24581
R68441 VSS.n3587 VSS.n3577 2.24581
R68442 VSS.n947 VSS.n946 2.24581
R68443 VSS.n3587 VSS.n936 2.24581
R68444 VSS.n947 VSS.n935 2.24581
R68445 VSS.n2821 VSS.n2744 2.24581
R68446 VSS.n2826 VSS.n2742 2.24581
R68447 VSS.n2821 VSS.n2817 2.24581
R68448 VSS.n2826 VSS.n2741 2.24581
R68449 VSS.n2821 VSS.n2818 2.24581
R68450 VSS.n2826 VSS.n2740 2.24581
R68451 VSS.n2821 VSS.n2819 2.24581
R68452 VSS.n2826 VSS.n2739 2.24581
R68453 VSS.n2821 VSS.n2820 2.24581
R68454 VSS.n2826 VSS.n2738 2.24581
R68455 VSS.n2975 VSS.n1108 2.24581
R68456 VSS.n2975 VSS.n1110 2.24581
R68457 VSS.n1116 VSS.n1115 2.24581
R68458 VSS.n2975 VSS.n1111 2.24581
R68459 VSS.n2967 VSS.n1116 2.24581
R68460 VSS.n1493 VSS.n1492 2.24581
R68461 VSS.n1499 VSS.n1425 2.24581
R68462 VSS.n1493 VSS.n1431 2.24581
R68463 VSS.n1499 VSS.n1428 2.24581
R68464 VSS.n1494 VSS.n1493 2.24581
R68465 VSS.n1499 VSS.n1429 2.24581
R68466 VSS.n1320 VSS.n1319 2.24581
R68467 VSS.n1325 VSS.n1321 2.24581
R68468 VSS.n1320 VSS.n1318 2.24581
R68469 VSS.n1325 VSS.n1322 2.24581
R68470 VSS.n1320 VSS.n1317 2.24581
R68471 VSS.n1325 VSS.n1323 2.24581
R68472 VSS.n1320 VSS.n1316 2.24581
R68473 VSS.n1325 VSS.n1324 2.24581
R68474 VSS.n1499 VSS.n1498 2.24581
R68475 VSS.n1116 VSS.n1102 2.24581
R68476 VSS.n4501 VSS.n4488 2.24581
R68477 VSS.n4389 VSS.n4381 2.24581
R68478 VSS.n4408 VSS.n4381 2.24581
R68479 VSS.n4393 VSS.n4381 2.24581
R68480 VSS.n4410 VSS.n4381 2.24581
R68481 VSS.n6033 VSS.n4412 2.24581
R68482 VSS.n6031 VSS.n6028 2.24581
R68483 VSS.n6033 VSS.n4413 2.24581
R68484 VSS.n6031 VSS.n6030 2.24581
R68485 VSS.n5583 VSS.n5462 2.24581
R68486 VSS.n5578 VSS.n5539 2.24581
R68487 VSS.n5583 VSS.n5463 2.24581
R68488 VSS.n5578 VSS.n5538 2.24581
R68489 VSS.n5583 VSS.n5460 2.24581
R68490 VSS.n5578 VSS.n5573 2.24581
R68491 VSS.n5583 VSS.n5459 2.24581
R68492 VSS.n5583 VSS.n5458 2.24581
R68493 VSS.n5578 VSS.n5574 2.24581
R68494 VSS.n5583 VSS.n5457 2.24581
R68495 VSS.n5583 VSS.n5456 2.24581
R68496 VSS.n5578 VSS.n5575 2.24581
R68497 VSS.n5581 VSS.n5527 2.24581
R68498 VSS.n5583 VSS.n5454 2.24581
R68499 VSS.n5578 VSS.n5577 2.24581
R68500 VSS.n5581 VSS.n5580 2.24581
R68501 VSS.n5583 VSS.n5452 2.24581
R68502 VSS.n5578 VSS.n5471 2.24581
R68503 VSS.n5036 VSS.n5028 2.24581
R68504 VSS.n5038 VSS.n5026 2.24581
R68505 VSS.n5040 VSS.n5028 2.24581
R68506 VSS.n5825 VSS.n5042 2.24581
R68507 VSS.n5043 VSS.n5026 2.24581
R68508 VSS.n5045 VSS.n5028 2.24581
R68509 VSS.n5825 VSS.n5047 2.24581
R68510 VSS.n5048 VSS.n5026 2.24581
R68511 VSS.n5811 VSS.n5028 2.24581
R68512 VSS.n5825 VSS.n5813 2.24581
R68513 VSS.n5814 VSS.n5026 2.24581
R68514 VSS.n5816 VSS.n5028 2.24581
R68515 VSS.n5825 VSS.n5818 2.24581
R68516 VSS.n5820 VSS.n5028 2.24581
R68517 VSS.n5825 VSS.n5822 2.24581
R68518 VSS.n5823 VSS.n5028 2.24581
R68519 VSS.n4414 VSS.n4381 2.24581
R68520 VSS.n3863 VSS.n728 2.24581
R68521 VSS.n3859 VSS.n731 2.24581
R68522 VSS.n3863 VSS.n729 2.24581
R68523 VSS.n3861 VSS.n736 2.24581
R68524 VSS.n5836 VSS.n4997 2.24442
R68525 VSS.n5782 VSS.n5013 2.24442
R68526 VSS.n5802 VSS.n5801 2.24442
R68527 VSS.n5866 VSS.n5865 2.24442
R68528 VSS.n5831 VSS.n5019 2.24442
R68529 VSS.n5827 VSS.n5017 2.24442
R68530 VSS.n5022 VSS.n5017 2.24442
R68531 VSS.n5829 VSS.n5016 2.24442
R68532 VSS.n4134 VSS.n554 2.24442
R68533 VSS.n4132 VSS.n4131 2.24442
R68534 VSS.n1122 VSS.n1121 2.2436
R68535 VSS.n1158 VSS.n1157 2.2436
R68536 VSS.n2973 VSS.n2972 2.2436
R68537 VSS.n2973 VSS.n1117 2.2436
R68538 VSS.n2899 VSS.n2888 2.2436
R68539 VSS.n2882 VSS.n1145 2.2436
R68540 VSS.n2901 VSS.n2900 2.2436
R68541 VSS.n2895 VSS.n2889 2.2436
R68542 VSS.n1254 VSS.n1230 2.24321
R68543 VSS.n1279 VSS.n1226 2.24321
R68544 VSS.n1534 VSS.n1214 2.24321
R68545 VSS.n1899 VSS.n1898 2.24321
R68546 VSS.n4185 VSS.n4184 2.23892
R68547 VSS.n537 VSS.n536 2.23892
R68548 VSS.n6171 VSS.n471 2.23892
R68549 VSS.n5494 VSS.n5493 2.23892
R68550 VSS.n5497 VSS.n5495 2.23892
R68551 VSS.n5488 VSS.n5484 2.23892
R68552 VSS.n5859 VSS.n4946 2.23892
R68553 VSS.n6156 VSS.n473 2.23892
R68554 VSS.n6188 VSS.n457 2.23892
R68555 VSS.n4092 VSS.n558 2.23892
R68556 VSS.n4097 VSS.n4095 2.23892
R68557 VSS.n6159 VSS.n6158 2.23892
R68558 VSS.n6189 VSS.n458 2.23892
R68559 VSS.n4094 VSS.n4091 2.23892
R68560 VSS.n4098 VSS.n4096 2.23892
R68561 VSS.n2982 VSS.n1093 2.2385
R68562 VSS.n2945 VSS.n2944 2.2385
R68563 VSS.n2918 VSS.n1162 2.2385
R68564 VSS.n2939 VSS.n1142 2.2385
R68565 VSS.n2978 VSS.n2977 2.2385
R68566 VSS.n2977 VSS.n1096 2.2385
R68567 VSS.n6176 VSS.n6175 2.23787
R68568 VSS.n4269 VSS.n4266 2.23787
R68569 VSS.n4763 VSS.n484 2.23787
R68570 VSS.n490 VSS.n487 2.23787
R68571 VSS.n4265 VSS.n4259 2.23787
R68572 VSS.n5503 VSS.n5481 2.23787
R68573 VSS.n6150 VSS.n6149 2.23787
R68574 VSS.n6149 VSS.n479 2.23787
R68575 VSS.n4183 VSS.n4181 2.23787
R68576 VSS.n4189 VSS.n4178 2.23787
R68577 VSS.n6151 VSS.n480 2.23787
R68578 VSS.n6147 VSS.n480 2.23787
R68579 VSS.n5501 VSS.n5489 2.23787
R68580 VSS.n4859 VSS.n4809 2.23714
R68581 VSS.n5985 VSS.n4800 2.23714
R68582 VSS.n4859 VSS.n4807 2.23714
R68583 VSS.n5985 VSS.n4799 2.23714
R68584 VSS.n4859 VSS.n4805 2.23714
R68585 VSS.n5985 VSS.n4798 2.23714
R68586 VSS.n4859 VSS.n4803 2.23714
R68587 VSS.n5985 VSS.n4797 2.23714
R68588 VSS.n4859 VSS.n4801 2.23714
R68589 VSS.n499 VSS.n489 2.23714
R68590 VSS.n6139 VSS.n496 2.23714
R68591 VSS.n495 VSS.n489 2.23714
R68592 VSS.n6139 VSS.n494 2.23714
R68593 VSS.n493 VSS.n489 2.23714
R68594 VSS.n6137 VSS.n489 2.23714
R68595 VSS.n585 VSS.n574 2.23714
R68596 VSS.n4089 VSS.n580 2.23714
R68597 VSS.n585 VSS.n581 2.23714
R68598 VSS.n4089 VSS.n579 2.23714
R68599 VSS.n585 VSS.n582 2.23714
R68600 VSS.n4089 VSS.n578 2.23714
R68601 VSS.n585 VSS.n583 2.23714
R68602 VSS.n4089 VSS.n577 2.23714
R68603 VSS.n585 VSS.n584 2.23714
R68604 VSS.n4089 VSS.n576 2.23714
R68605 VSS.n3723 VSS.n850 2.23714
R68606 VSS.n3726 VSS.n853 2.23714
R68607 VSS.n3723 VSS.n3722 2.23714
R68608 VSS.n3726 VSS.n854 2.23714
R68609 VSS.n3723 VSS.n3721 2.23714
R68610 VSS.n3726 VSS.n855 2.23714
R68611 VSS.n3723 VSS.n3720 2.23714
R68612 VSS.n3726 VSS.n856 2.23714
R68613 VSS.n3723 VSS.n3719 2.23714
R68614 VSS.n3726 VSS.n857 2.23714
R68615 VSS.n3723 VSS.n3718 2.23714
R68616 VSS.n3726 VSS.n858 2.23714
R68617 VSS.n3723 VSS.n3717 2.23714
R68618 VSS.n3726 VSS.n859 2.23714
R68619 VSS.n3723 VSS.n3716 2.23714
R68620 VSS.n3726 VSS.n860 2.23714
R68621 VSS.n3723 VSS.n3715 2.23714
R68622 VSS.n3726 VSS.n861 2.23714
R68623 VSS.n3723 VSS.n3714 2.23714
R68624 VSS.n3726 VSS.n862 2.23714
R68625 VSS.n3723 VSS.n3713 2.23714
R68626 VSS.n3726 VSS.n863 2.23714
R68627 VSS.n3068 VSS.n3067 2.23714
R68628 VSS.n3403 VSS.n1002 2.23714
R68629 VSS.n3067 VSS.n1045 2.23714
R68630 VSS.n3403 VSS.n1001 2.23714
R68631 VSS.n3067 VSS.n1046 2.23714
R68632 VSS.n3403 VSS.n1000 2.23714
R68633 VSS.n3067 VSS.n1047 2.23714
R68634 VSS.n3403 VSS.n999 2.23714
R68635 VSS.n3067 VSS.n1048 2.23714
R68636 VSS.n3403 VSS.n998 2.23714
R68637 VSS.n1060 VSS.n1049 2.23714
R68638 VSS.n3064 VSS.n1055 2.23714
R68639 VSS.n1060 VSS.n1056 2.23714
R68640 VSS.n3064 VSS.n1054 2.23714
R68641 VSS.n1060 VSS.n1057 2.23714
R68642 VSS.n3064 VSS.n1053 2.23714
R68643 VSS.n1060 VSS.n1058 2.23714
R68644 VSS.n3064 VSS.n1052 2.23714
R68645 VSS.n1060 VSS.n1059 2.23714
R68646 VSS.n3064 VSS.n1051 2.23714
R68647 VSS.n1833 VSS.n1253 2.23714
R68648 VSS.n1830 VSS.n1827 2.23714
R68649 VSS.n1833 VSS.n1256 2.23714
R68650 VSS.n1831 VSS.n1830 2.23714
R68651 VSS.n1833 VSS.n1832 2.23714
R68652 VSS.n1830 VSS.n1249 2.23714
R68653 VSS.n1879 VSS.n1240 2.23714
R68654 VSS.n1836 VSS.n1248 2.23714
R68655 VSS.n1879 VSS.n1239 2.23714
R68656 VSS.n1836 VSS.n1247 2.23714
R68657 VSS.n1879 VSS.n1238 2.23714
R68658 VSS.n1836 VSS.n1246 2.23714
R68659 VSS.n1879 VSS.n1237 2.23714
R68660 VSS.n1836 VSS.n1235 2.23714
R68661 VSS.n1830 VSS.n1826 2.23714
R68662 VSS.n3724 VSS.n3723 2.23714
R68663 VSS.n501 VSS.n489 2.23714
R68664 VSS.n5985 VSS.n4481 2.23714
R68665 VSS.n5985 VSS.n4480 2.23714
R68666 VSS.n5985 VSS.n4479 2.23714
R68667 VSS.n5985 VSS.n4478 2.23714
R68668 VSS.n4859 VSS.n4473 2.23714
R68669 VSS.n5985 VSS.n4477 2.23714
R68670 VSS.n4859 VSS.n4858 2.23714
R68671 VSS.n5985 VSS.n4476 2.23714
R68672 VSS.n5852 VSS.n4947 2.23714
R68673 VSS.n5855 VSS.n4957 2.23714
R68674 VSS.n5852 VSS.n4974 2.23714
R68675 VSS.n5855 VSS.n4958 2.23714
R68676 VSS.n5852 VSS.n4971 2.23714
R68677 VSS.n5855 VSS.n4955 2.23714
R68678 VSS.n5852 VSS.n4970 2.23714
R68679 VSS.n5852 VSS.n4969 2.23714
R68680 VSS.n5855 VSS.n4953 2.23714
R68681 VSS.n5852 VSS.n4968 2.23714
R68682 VSS.n5852 VSS.n4967 2.23714
R68683 VSS.n5855 VSS.n4951 2.23714
R68684 VSS.n5855 VSS.n4962 2.23714
R68685 VSS.n5852 VSS.n4965 2.23714
R68686 VSS.n5855 VSS.n4950 2.23714
R68687 VSS.n5855 VSS.n5854 2.23714
R68688 VSS.n5852 VSS.n4963 2.23714
R68689 VSS.n5855 VSS.n4949 2.23714
R68690 VSS.n5868 VSS.n4928 2.23714
R68691 VSS.n4943 VSS.n4939 2.23714
R68692 VSS.n5868 VSS.n4926 2.23714
R68693 VSS.n4943 VSS.n4938 2.23714
R68694 VSS.n4943 VSS.n4940 2.23714
R68695 VSS.n5868 VSS.n4924 2.23714
R68696 VSS.n4943 VSS.n4937 2.23714
R68697 VSS.n4943 VSS.n4941 2.23714
R68698 VSS.n5868 VSS.n4922 2.23714
R68699 VSS.n4943 VSS.n4936 2.23714
R68700 VSS.n4943 VSS.n4942 2.23714
R68701 VSS.n5868 VSS.n4920 2.23714
R68702 VSS.n4943 VSS.n4935 2.23714
R68703 VSS.n5868 VSS.n4919 2.23714
R68704 VSS.n4943 VSS.n4934 2.23714
R68705 VSS.n5985 VSS.n4475 2.23714
R68706 VSS.n2952 VSS.n1134 2.23714
R68707 VSS.n2954 VSS.n2953 2.23714
R68708 VSS.n2948 VSS.n2947 2.23714
R68709 VSS.n1137 VSS.n1135 2.23714
R68710 VSS.n4461 VSS.n4449 2.23714
R68711 VSS.n5996 VSS.n4459 2.23714
R68712 VSS.n5996 VSS.n4462 2.23714
R68713 VSS.n4463 VSS.n4449 2.23714
R68714 VSS.n5996 VSS.n4458 2.23714
R68715 VSS.n5996 VSS.n4464 2.23714
R68716 VSS.n4465 VSS.n4449 2.23714
R68717 VSS.n5996 VSS.n4457 2.23714
R68718 VSS.n5996 VSS.n4466 2.23714
R68719 VSS.n4467 VSS.n4449 2.23714
R68720 VSS.n5996 VSS.n4456 2.23714
R68721 VSS.n5996 VSS.n4468 2.23714
R68722 VSS.n4469 VSS.n4449 2.23714
R68723 VSS.n5996 VSS.n4455 2.23714
R68724 VSS.n4765 VSS.n4515 2.23714
R68725 VSS.n4765 VSS.n4761 2.23714
R68726 VSS.n4768 VSS.n4517 2.23714
R68727 VSS.n4768 VSS.n4520 2.23714
R68728 VSS.n4765 VSS.n4762 2.23714
R68729 VSS.n4768 VSS.n4521 2.23714
R68730 VSS.n4766 VSS.n4765 2.23714
R68731 VSS.n4105 VSS.n571 2.23714
R68732 VSS.n4106 VSS.n572 2.23714
R68733 VSS.n4107 VSS.n571 2.23714
R68734 VSS.n4108 VSS.n572 2.23714
R68735 VSS.n4109 VSS.n571 2.23714
R68736 VSS.n4110 VSS.n572 2.23714
R68737 VSS.n4111 VSS.n571 2.23714
R68738 VSS.n4112 VSS.n572 2.23714
R68739 VSS.n4113 VSS.n571 2.23714
R68740 VSS.n4114 VSS.n572 2.23714
R68741 VSS.n3637 VSS.n3636 2.23714
R68742 VSS.n3640 VSS.n883 2.23714
R68743 VSS.n3637 VSS.n3635 2.23714
R68744 VSS.n3640 VSS.n884 2.23714
R68745 VSS.n3637 VSS.n3634 2.23714
R68746 VSS.n3640 VSS.n885 2.23714
R68747 VSS.n3637 VSS.n3633 2.23714
R68748 VSS.n3640 VSS.n886 2.23714
R68749 VSS.n3637 VSS.n3632 2.23714
R68750 VSS.n3640 VSS.n887 2.23714
R68751 VSS.n3637 VSS.n3631 2.23714
R68752 VSS.n3640 VSS.n888 2.23714
R68753 VSS.n3637 VSS.n3630 2.23714
R68754 VSS.n3640 VSS.n889 2.23714
R68755 VSS.n3637 VSS.n3629 2.23714
R68756 VSS.n3640 VSS.n890 2.23714
R68757 VSS.n3637 VSS.n3628 2.23714
R68758 VSS.n3640 VSS.n891 2.23714
R68759 VSS.n3637 VSS.n3627 2.23714
R68760 VSS.n3640 VSS.n892 2.23714
R68761 VSS.n3637 VSS.n3626 2.23714
R68762 VSS.n3640 VSS.n893 2.23714
R68763 VSS.n3638 VSS.n3637 2.23714
R68764 VSS.n2779 VSS.n973 2.23714
R68765 VSS.n3436 VSS.n979 2.23714
R68766 VSS.n2779 VSS.n2773 2.23714
R68767 VSS.n3436 VSS.n978 2.23714
R68768 VSS.n2779 VSS.n2774 2.23714
R68769 VSS.n3436 VSS.n977 2.23714
R68770 VSS.n2779 VSS.n2775 2.23714
R68771 VSS.n3436 VSS.n976 2.23714
R68772 VSS.n2779 VSS.n2776 2.23714
R68773 VSS.n3436 VSS.n975 2.23714
R68774 VSS.n2986 VSS.n1085 2.23714
R68775 VSS.n2986 VSS.n1087 2.23714
R68776 VSS.n1086 VSS.n1077 2.23714
R68777 VSS.n1088 VSS.n1077 2.23714
R68778 VSS.n2986 VSS.n1089 2.23714
R68779 VSS.n1090 VSS.n1077 2.23714
R68780 VSS.n1751 VSS.n1750 2.23714
R68781 VSS.n1754 VSS.n1277 2.23714
R68782 VSS.n1752 VSS.n1751 2.23714
R68783 VSS.n1754 VSS.n1753 2.23714
R68784 VSS.n1754 VSS.n1276 2.23714
R68785 VSS.n1751 VSS.n1749 2.23714
R68786 VSS.n1754 VSS.n1275 2.23714
R68787 VSS.n1742 VSS.n1283 2.23714
R68788 VSS.n1746 VSS.n1286 2.23714
R68789 VSS.n1742 VSS.n1741 2.23714
R68790 VSS.n1746 VSS.n1287 2.23714
R68791 VSS.n1742 VSS.n1740 2.23714
R68792 VSS.n1746 VSS.n1288 2.23714
R68793 VSS.n1742 VSS.n1739 2.23714
R68794 VSS.n1746 VSS.n1289 2.23714
R68795 VSS.n5996 VSS.n5992 2.23714
R68796 VSS.n5994 VSS.n4449 2.23714
R68797 VSS.n5996 VSS.n5995 2.23714
R68798 VSS.n5993 VSS.n4449 2.23714
R68799 VSS.n5643 VSS.n5253 2.23714
R68800 VSS.n5646 VSS.n5187 2.23714
R68801 VSS.n5643 VSS.n5254 2.23714
R68802 VSS.n5646 VSS.n5188 2.23714
R68803 VSS.n5643 VSS.n5201 2.23714
R68804 VSS.n5646 VSS.n5184 2.23714
R68805 VSS.n5643 VSS.n5200 2.23714
R68806 VSS.n5643 VSS.n5199 2.23714
R68807 VSS.n5646 VSS.n5182 2.23714
R68808 VSS.n5643 VSS.n5198 2.23714
R68809 VSS.n5643 VSS.n5197 2.23714
R68810 VSS.n5646 VSS.n5180 2.23714
R68811 VSS.n5646 VSS.n5192 2.23714
R68812 VSS.n5643 VSS.n5195 2.23714
R68813 VSS.n5646 VSS.n5179 2.23714
R68814 VSS.n5646 VSS.n5645 2.23714
R68815 VSS.n5643 VSS.n5193 2.23714
R68816 VSS.n5646 VSS.n5178 2.23714
R68817 VSS.n5804 VSS.n5065 2.23714
R68818 VSS.n5797 VSS.n5794 2.23714
R68819 VSS.n5804 VSS.n5062 2.23714
R68820 VSS.n5797 VSS.n5075 2.23714
R68821 VSS.n5797 VSS.n5795 2.23714
R68822 VSS.n5804 VSS.n5060 2.23714
R68823 VSS.n5797 VSS.n5074 2.23714
R68824 VSS.n5797 VSS.n5796 2.23714
R68825 VSS.n5804 VSS.n5058 2.23714
R68826 VSS.n5797 VSS.n5073 2.23714
R68827 VSS.n5797 VSS.n5053 2.23714
R68828 VSS.n5804 VSS.n5057 2.23714
R68829 VSS.n5797 VSS.n5072 2.23714
R68830 VSS.n5804 VSS.n5056 2.23714
R68831 VSS.n5797 VSS.n5071 2.23714
R68832 VSS.n1153 VSS.n1152 2.23714
R68833 VSS.n2931 VSS.n2930 2.23714
R68834 VSS.n1150 VSS.n1149 2.23714
R68835 VSS.n2935 VSS.n2934 2.23714
R68836 VSS.n1148 VSS.n1146 2.23714
R68837 VSS.n6104 VSS.n4301 2.23714
R68838 VSS.n6107 VSS.n4286 2.23714
R68839 VSS.n6107 VSS.n4288 2.23714
R68840 VSS.n6104 VSS.n4302 2.23714
R68841 VSS.n6107 VSS.n4285 2.23714
R68842 VSS.n6107 VSS.n4289 2.23714
R68843 VSS.n6104 VSS.n4299 2.23714
R68844 VSS.n6107 VSS.n4284 2.23714
R68845 VSS.n6107 VSS.n4290 2.23714
R68846 VSS.n6104 VSS.n4304 2.23714
R68847 VSS.n6107 VSS.n4283 2.23714
R68848 VSS.n6107 VSS.n4291 2.23714
R68849 VSS.n6104 VSS.n4279 2.23714
R68850 VSS.n6107 VSS.n4282 2.23714
R68851 VSS.n4274 VSS.n4268 2.23714
R68852 VSS.n6114 VSS.n4268 2.23714
R68853 VSS.n6121 VSS.n4271 2.23714
R68854 VSS.n6121 VSS.n6115 2.23714
R68855 VSS.n6117 VSS.n4268 2.23714
R68856 VSS.n6121 VSS.n6118 2.23714
R68857 VSS.n6119 VSS.n4268 2.23714
R68858 VSS.n3935 VSS.n3934 2.23714
R68859 VSS.n3937 VSS.n3936 2.23714
R68860 VSS.n3934 VSS.n659 2.23714
R68861 VSS.n3937 VSS.n658 2.23714
R68862 VSS.n3934 VSS.n661 2.23714
R68863 VSS.n3937 VSS.n657 2.23714
R68864 VSS.n3934 VSS.n662 2.23714
R68865 VSS.n3937 VSS.n656 2.23714
R68866 VSS.n3934 VSS.n663 2.23714
R68867 VSS.n3937 VSS.n655 2.23714
R68868 VSS.n3534 VSS.n3532 2.23714
R68869 VSS.n3531 VSS.n963 2.23714
R68870 VSS.n3534 VSS.n3530 2.23714
R68871 VSS.n3529 VSS.n963 2.23714
R68872 VSS.n3534 VSS.n3528 2.23714
R68873 VSS.n3527 VSS.n963 2.23714
R68874 VSS.n3534 VSS.n3526 2.23714
R68875 VSS.n3525 VSS.n963 2.23714
R68876 VSS.n3534 VSS.n3524 2.23714
R68877 VSS.n3523 VSS.n963 2.23714
R68878 VSS.n3534 VSS.n3522 2.23714
R68879 VSS.n3521 VSS.n963 2.23714
R68880 VSS.n3534 VSS.n3520 2.23714
R68881 VSS.n3519 VSS.n963 2.23714
R68882 VSS.n3534 VSS.n3518 2.23714
R68883 VSS.n3517 VSS.n963 2.23714
R68884 VSS.n3534 VSS.n3516 2.23714
R68885 VSS.n3515 VSS.n963 2.23714
R68886 VSS.n3534 VSS.n3514 2.23714
R68887 VSS.n3513 VSS.n963 2.23714
R68888 VSS.n3534 VSS.n3512 2.23714
R68889 VSS.n3511 VSS.n963 2.23714
R68890 VSS.n3534 VSS.n3510 2.23714
R68891 VSS.n2860 VSS.n1163 2.23714
R68892 VSS.n2861 VSS.n2859 2.23714
R68893 VSS.n2862 VSS.n1163 2.23714
R68894 VSS.n2863 VSS.n2859 2.23714
R68895 VSS.n2864 VSS.n1163 2.23714
R68896 VSS.n2865 VSS.n2859 2.23714
R68897 VSS.n2866 VSS.n1163 2.23714
R68898 VSS.n2867 VSS.n2859 2.23714
R68899 VSS.n2868 VSS.n1163 2.23714
R68900 VSS.n2869 VSS.n2859 2.23714
R68901 VSS.n2872 VSS.n1160 2.23714
R68902 VSS.n2921 VSS.n1160 2.23714
R68903 VSS.n2920 VSS.n1161 2.23714
R68904 VSS.n2922 VSS.n1161 2.23714
R68905 VSS.n2923 VSS.n1160 2.23714
R68906 VSS.n2924 VSS.n1161 2.23714
R68907 VSS.n1532 VSS.n1355 2.23714
R68908 VSS.n1536 VSS.n1357 2.23714
R68909 VSS.n1539 VSS.n1355 2.23714
R68910 VSS.n1538 VSS.n1536 2.23714
R68911 VSS.n1540 VSS.n1536 2.23714
R68912 VSS.n1541 VSS.n1355 2.23714
R68913 VSS.n1542 VSS.n1536 2.23714
R68914 VSS.n1617 VSS.n1545 2.23714
R68915 VSS.n1354 VSS.n1342 2.23714
R68916 VSS.n1617 VSS.n1353 2.23714
R68917 VSS.n1352 VSS.n1342 2.23714
R68918 VSS.n1617 VSS.n1351 2.23714
R68919 VSS.n1350 VSS.n1342 2.23714
R68920 VSS.n1617 VSS.n1349 2.23714
R68921 VSS.n1348 VSS.n1342 2.23714
R68922 VSS.n6107 VSS.n4292 2.23714
R68923 VSS.n6105 VSS.n6104 2.23714
R68924 VSS.n6107 VSS.n6106 2.23714
R68925 VSS.n6104 VSS.n4293 2.23714
R68926 VSS.n5619 VSS.n5614 2.23714
R68927 VSS.n5622 VSS.n5298 2.23714
R68928 VSS.n5619 VSS.n5615 2.23714
R68929 VSS.n5622 VSS.n5299 2.23714
R68930 VSS.n5619 VSS.n5310 2.23714
R68931 VSS.n5622 VSS.n5295 2.23714
R68932 VSS.n5619 VSS.n5309 2.23714
R68933 VSS.n5619 VSS.n5308 2.23714
R68934 VSS.n5622 VSS.n5293 2.23714
R68935 VSS.n5619 VSS.n5307 2.23714
R68936 VSS.n5619 VSS.n5288 2.23714
R68937 VSS.n5622 VSS.n5292 2.23714
R68938 VSS.n5622 VSS.n5302 2.23714
R68939 VSS.n5619 VSS.n5305 2.23714
R68940 VSS.n5622 VSS.n5291 2.23714
R68941 VSS.n5622 VSS.n5621 2.23714
R68942 VSS.n5619 VSS.n5303 2.23714
R68943 VSS.n5622 VSS.n5290 2.23714
R68944 VSS.n5784 VSS.n5092 2.23714
R68945 VSS.n5781 VSS.n5081 2.23714
R68946 VSS.n5784 VSS.n5090 2.23714
R68947 VSS.n5781 VSS.n5776 2.23714
R68948 VSS.n5781 VSS.n5778 2.23714
R68949 VSS.n5784 VSS.n5088 2.23714
R68950 VSS.n5781 VSS.n5775 2.23714
R68951 VSS.n5781 VSS.n5779 2.23714
R68952 VSS.n5784 VSS.n5086 2.23714
R68953 VSS.n5781 VSS.n5774 2.23714
R68954 VSS.n5781 VSS.n5780 2.23714
R68955 VSS.n5784 VSS.n5084 2.23714
R68956 VSS.n5781 VSS.n5773 2.23714
R68957 VSS.n5784 VSS.n5083 2.23714
R68958 VSS.n5781 VSS.n5772 2.23714
R68959 VSS.n6098 VSS.n4318 2.23714
R68960 VSS.n6095 VSS.n4332 2.23714
R68961 VSS.n6095 VSS.n6086 2.23714
R68962 VSS.n6098 VSS.n4320 2.23714
R68963 VSS.n6095 VSS.n4331 2.23714
R68964 VSS.n6095 VSS.n6087 2.23714
R68965 VSS.n6098 VSS.n4316 2.23714
R68966 VSS.n6095 VSS.n4330 2.23714
R68967 VSS.n6095 VSS.n6088 2.23714
R68968 VSS.n6098 VSS.n4322 2.23714
R68969 VSS.n6095 VSS.n4329 2.23714
R68970 VSS.n6095 VSS.n6089 2.23714
R68971 VSS.n6098 VSS.n4314 2.23714
R68972 VSS.n6095 VSS.n4328 2.23714
R68973 VSS.n4263 VSS.n4260 2.23714
R68974 VSS.n4263 VSS.n4261 2.23714
R68975 VSS.n6129 VSS.n4253 2.23714
R68976 VSS.n6129 VSS.n4257 2.23714
R68977 VSS.n4263 VSS.n4262 2.23714
R68978 VSS.n6129 VSS.n4258 2.23714
R68979 VSS.n4263 VSS.n4250 2.23714
R68980 VSS.n2205 VSS.n2150 2.23714
R68981 VSS.n2206 VSS.n2203 2.23714
R68982 VSS.n2207 VSS.n2150 2.23714
R68983 VSS.n2208 VSS.n2203 2.23714
R68984 VSS.n2209 VSS.n2150 2.23714
R68985 VSS.n2210 VSS.n2203 2.23714
R68986 VSS.n2211 VSS.n2150 2.23714
R68987 VSS.n2212 VSS.n2203 2.23714
R68988 VSS.n2213 VSS.n2150 2.23714
R68989 VSS.n2214 VSS.n2203 2.23714
R68990 VSS.n2145 VSS.n2078 2.23714
R68991 VSS.n2148 VSS.n2081 2.23714
R68992 VSS.n2145 VSS.n2144 2.23714
R68993 VSS.n2148 VSS.n2082 2.23714
R68994 VSS.n2145 VSS.n2143 2.23714
R68995 VSS.n2148 VSS.n2083 2.23714
R68996 VSS.n2145 VSS.n2142 2.23714
R68997 VSS.n2148 VSS.n2084 2.23714
R68998 VSS.n2145 VSS.n2141 2.23714
R68999 VSS.n2148 VSS.n2085 2.23714
R69000 VSS.n2145 VSS.n2140 2.23714
R69001 VSS.n2148 VSS.n2086 2.23714
R69002 VSS.n2145 VSS.n2139 2.23714
R69003 VSS.n2148 VSS.n2087 2.23714
R69004 VSS.n2145 VSS.n2138 2.23714
R69005 VSS.n2148 VSS.n2088 2.23714
R69006 VSS.n2145 VSS.n2137 2.23714
R69007 VSS.n2148 VSS.n2089 2.23714
R69008 VSS.n2145 VSS.n2136 2.23714
R69009 VSS.n2148 VSS.n2090 2.23714
R69010 VSS.n2145 VSS.n2135 2.23714
R69011 VSS.n2148 VSS.n2091 2.23714
R69012 VSS.n2146 VSS.n2145 2.23714
R69013 VSS.n2067 VSS.n1184 2.23714
R69014 VSS.n2687 VSS.n2066 2.23714
R69015 VSS.n2065 VSS.n1184 2.23714
R69016 VSS.n2687 VSS.n2064 2.23714
R69017 VSS.n2063 VSS.n1184 2.23714
R69018 VSS.n2687 VSS.n2062 2.23714
R69019 VSS.n2061 VSS.n1184 2.23714
R69020 VSS.n2687 VSS.n2060 2.23714
R69021 VSS.n2059 VSS.n1184 2.23714
R69022 VSS.n2687 VSS.n2058 2.23714
R69023 VSS.n1909 VSS.n1185 2.23714
R69024 VSS.n2055 VSS.n1191 2.23714
R69025 VSS.n1909 VSS.n1195 2.23714
R69026 VSS.n2055 VSS.n1190 2.23714
R69027 VSS.n1909 VSS.n1196 2.23714
R69028 VSS.n2055 VSS.n1189 2.23714
R69029 VSS.n1909 VSS.n1197 2.23714
R69030 VSS.n2055 VSS.n1188 2.23714
R69031 VSS.n1909 VSS.n1198 2.23714
R69032 VSS.n2055 VSS.n1187 2.23714
R69033 VSS.n1903 VSS.n1199 2.23714
R69034 VSS.n1906 VSS.n1204 2.23714
R69035 VSS.n1904 VSS.n1903 2.23714
R69036 VSS.n1906 VSS.n1905 2.23714
R69037 VSS.n1906 VSS.n1202 2.23714
R69038 VSS.n1903 VSS.n1210 2.23714
R69039 VSS.n1906 VSS.n1201 2.23714
R69040 VSS.n1596 VSS.n1548 2.23714
R69041 VSS.n1597 VSS.n1594 2.23714
R69042 VSS.n1598 VSS.n1548 2.23714
R69043 VSS.n1599 VSS.n1594 2.23714
R69044 VSS.n1600 VSS.n1548 2.23714
R69045 VSS.n1601 VSS.n1594 2.23714
R69046 VSS.n1602 VSS.n1548 2.23714
R69047 VSS.n1603 VSS.n1594 2.23714
R69048 VSS.n6095 VSS.n4310 2.23714
R69049 VSS.n6098 VSS.n4326 2.23714
R69050 VSS.n6096 VSS.n6095 2.23714
R69051 VSS.n6098 VSS.n6097 2.23714
R69052 VSS.n5632 VSS.n5271 2.23714
R69053 VSS.n5629 VSS.n5282 2.23714
R69054 VSS.n5632 VSS.n5272 2.23714
R69055 VSS.n5629 VSS.n5283 2.23714
R69056 VSS.n5632 VSS.n5268 2.23714
R69057 VSS.n5629 VSS.n5280 2.23714
R69058 VSS.n5632 VSS.n5267 2.23714
R69059 VSS.n5632 VSS.n5266 2.23714
R69060 VSS.n5629 VSS.n5278 2.23714
R69061 VSS.n5632 VSS.n5265 2.23714
R69062 VSS.n5632 VSS.n5264 2.23714
R69063 VSS.n5629 VSS.n5276 2.23714
R69064 VSS.n5629 VSS.n5259 2.23714
R69065 VSS.n5632 VSS.n5263 2.23714
R69066 VSS.n5630 VSS.n5629 2.23714
R69067 VSS.n5629 VSS.n5628 2.23714
R69068 VSS.n5632 VSS.n5261 2.23714
R69069 VSS.n5629 VSS.n5275 2.23714
R69070 VSS.n5840 VSS.n4981 2.23714
R69071 VSS.n5842 VSS.n4992 2.23714
R69072 VSS.n5840 VSS.n5005 2.23714
R69073 VSS.n5842 VSS.n4989 2.23714
R69074 VSS.n5842 VSS.n4993 2.23714
R69075 VSS.n5840 VSS.n5003 2.23714
R69076 VSS.n5842 VSS.n4988 2.23714
R69077 VSS.n5842 VSS.n4994 2.23714
R69078 VSS.n5840 VSS.n5001 2.23714
R69079 VSS.n5842 VSS.n4987 2.23714
R69080 VSS.n5842 VSS.n4995 2.23714
R69081 VSS.n5840 VSS.n4999 2.23714
R69082 VSS.n5842 VSS.n4986 2.23714
R69083 VSS.n5840 VSS.n4998 2.23714
R69084 VSS.n5842 VSS.n4985 2.23714
R69085 VSS.n1882 VSS.n1881 2.21947
R69086 VSS.n1744 VSS.n1233 2.21947
R69087 VSS.n5807 VSS.n5806 2.21947
R69088 VSS.n5108 VSS.n5107 2.21947
R69089 VSS.n5097 VSS.n5096 2.21947
R69090 VSS.n5792 VSS.n5791 2.21947
R69091 VSS.n5848 VSS.n4977 2.21947
R69092 VSS.n5467 VSS.n5194 2.21947
R69093 VSS.n5639 VSS.n5638 2.21947
R69094 VSS.n5523 VSS.n5522 2.21947
R69095 VSS.n5516 VSS.n5515 2.21947
R69096 VSS.n5534 VSS.n5533 2.21947
R69097 VSS.n5990 VSS.n5989 2.21947
R69098 VSS.n4819 VSS.n4812 2.21947
R69099 VSS.n4831 VSS.n4824 2.21947
R69100 VSS.n4843 VSS.n4836 2.21947
R69101 VSS.n4855 VSS.n4848 2.21947
R69102 VSS.n4794 VSS.n4483 2.21947
R69103 VSS.n4788 VSS.n4787 2.21947
R69104 VSS.n4786 VSS.n4785 2.21947
R69105 VSS.n4780 VSS.n4486 2.21947
R69106 VSS.n4771 VSS.n4770 2.21947
R69107 VSS.n6135 VSS.n504 2.21947
R69108 VSS.n4239 VSS.n4238 2.21947
R69109 VSS.n4241 VSS.n4240 2.21947
R69110 VSS.n4236 VSS.n4235 2.21947
R69111 VSS.n521 VSS.n513 2.21947
R69112 VSS.n4222 VSS.n4221 2.21947
R69113 VSS.n4220 VSS.n4219 2.21947
R69114 VSS.n532 VSS.n524 2.21947
R69115 VSS.n4206 VSS.n4205 2.21947
R69116 VSS.n4204 VSS.n4203 2.21947
R69117 VSS.n4193 VSS.n540 2.21947
R69118 VSS.n4174 VSS.n4173 2.21947
R69119 VSS.n4172 VSS.n4171 2.21947
R69120 VSS.n4166 VSS.n543 2.21947
R69121 VSS.n4160 VSS.n4159 2.21947
R69122 VSS.n4158 VSS.n4157 2.21947
R69123 VSS.n4152 VSS.n547 2.21947
R69124 VSS.n4146 VSS.n4145 2.21947
R69125 VSS.n4144 VSS.n4143 2.21947
R69126 VSS.n4138 VSS.n551 2.21947
R69127 VSS.n1615 VSS.n1614 2.21947
R69128 VSS.n5118 VSS.n5117 2.21947
R69129 VSS.n5114 VSS.n5113 2.21947
R69130 VSS.n5103 VSS.n5102 2.21947
R69131 VSS.n5788 VSS.n5786 2.21947
R69132 VSS.n5845 VSS.n4979 2.21947
R69133 VSS.n5465 VSS.n5304 2.21947
R69134 VSS.n5635 VSS.n5257 2.21947
R69135 VSS.n5625 VSS.n5624 2.21947
R69136 VSS.n5512 VSS.n5510 2.21947
R69137 VSS.n5530 VSS.n5528 2.21947
R69138 VSS.n6102 VSS.n6101 2.21947
R69139 VSS.n4816 VSS.n4814 2.21947
R69140 VSS.n4828 VSS.n4826 2.21947
R69141 VSS.n4840 VSS.n4838 2.21947
R69142 VSS.n4852 VSS.n4850 2.21947
R69143 VSS.n6109 VSS.n4278 2.21947
R69144 VSS.n6110 VSS.n4277 2.21947
R69145 VSS.n6111 VSS.n4276 2.21947
R69146 VSS.n6112 VSS.n4275 2.21947
R69147 VSS.n4511 VSS.n4508 2.21947
R69148 VSS.n6132 VSS.n506 2.21947
R69149 VSS.n4248 VSS.n4247 2.21947
R69150 VSS.n4246 VSS.n4245 2.21947
R69151 VSS.n4232 VSS.n509 2.21947
R69152 VSS.n4229 VSS.n4228 2.21947
R69153 VSS.n4227 VSS.n4226 2.21947
R69154 VSS.n4216 VSS.n517 2.21947
R69155 VSS.n4213 VSS.n4212 2.21947
R69156 VSS.n4211 VSS.n4210 2.21947
R69157 VSS.n4200 VSS.n528 2.21947
R69158 VSS.n6177 VSS.n468 2.21947
R69159 VSS.n6178 VSS.n467 2.21947
R69160 VSS.n6179 VSS.n466 2.21947
R69161 VSS.n6180 VSS.n465 2.21947
R69162 VSS.n6181 VSS.n464 2.21947
R69163 VSS.n6182 VSS.n463 2.21947
R69164 VSS.n6183 VSS.n462 2.21947
R69165 VSS.n6184 VSS.n461 2.21947
R69166 VSS.n6185 VSS.n460 2.21947
R69167 VSS.n6186 VSS.n459 2.21947
R69168 VSS.n1606 VSS.n1605 2.21947
R69169 VSS.n1611 VSS.n1326 2.21947
R69170 VSS.n5809 VSS.n5050 2.21947
R69171 VSS.n5111 VSS.n5110 2.21947
R69172 VSS.n5100 VSS.n5099 2.21947
R69173 VSS.n5789 VSS.n5079 2.21947
R69174 VSS.n5846 VSS.n4978 2.21947
R69175 VSS.n5469 VSS.n5466 2.21947
R69176 VSS.n5636 VSS.n5256 2.21947
R69177 VSS.n5525 VSS.n5286 2.21947
R69178 VSS.n5518 VSS.n5513 2.21947
R69179 VSS.n5536 VSS.n5531 2.21947
R69180 VSS.n4421 VSS.n4308 2.21947
R69181 VSS.n4817 VSS.n4813 2.21947
R69182 VSS.n4829 VSS.n4825 2.21947
R69183 VSS.n4841 VSS.n4837 2.21947
R69184 VSS.n4853 VSS.n4849 2.21947
R69185 VSS.n4792 VSS.n4791 2.21947
R69186 VSS.n4790 VSS.n4485 2.21947
R69187 VSS.n4783 VSS.n4484 2.21947
R69188 VSS.n4778 VSS.n4777 2.21947
R69189 VSS.n4773 VSS.n4512 2.21947
R69190 VSS.n6133 VSS.n505 2.21947
R69191 VSS.n511 VSS.n508 2.21947
R69192 VSS.n4244 VSS.n4243 2.21947
R69193 VSS.n4233 VSS.n510 2.21947
R69194 VSS.n519 VSS.n516 2.21947
R69195 VSS.n4225 VSS.n4224 2.21947
R69196 VSS.n4217 VSS.n518 2.21947
R69197 VSS.n530 VSS.n527 2.21947
R69198 VSS.n4209 VSS.n4208 2.21947
R69199 VSS.n4201 VSS.n529 2.21947
R69200 VSS.n4191 VSS.n4190 2.21947
R69201 VSS.n4176 VSS.n542 2.21947
R69202 VSS.n4169 VSS.n541 2.21947
R69203 VSS.n4164 VSS.n4163 2.21947
R69204 VSS.n4162 VSS.n546 2.21947
R69205 VSS.n4155 VSS.n545 2.21947
R69206 VSS.n4150 VSS.n4149 2.21947
R69207 VSS.n4148 VSS.n550 2.21947
R69208 VSS.n4141 VSS.n549 2.21947
R69209 VSS.n4136 VSS.n4135 2.21947
R69210 VSS.n4102 VSS.n4101 2.16043
R69211 VSS.n3395 VSS.n3103 1.95638
R69212 VSS.n3392 VSS.n3103 1.95638
R69213 VSS.n3273 VSS.n3268 1.95638
R69214 VSS.n3273 VSS.n3133 1.95638
R69215 VSS.n3129 VSS.n3100 1.95638
R69216 VSS.n3132 VSS.n3129 1.95638
R69217 VSS.n2545 VSS.n2285 1.89035
R69218 VSS.n2543 VSS.n2443 1.89035
R69219 VSS.n2545 VSS.n2284 1.89035
R69220 VSS.n2543 VSS.n2442 1.89035
R69221 VSS.n2545 VSS.n2283 1.89035
R69222 VSS.n2543 VSS.n2441 1.89035
R69223 VSS.n2545 VSS.n2282 1.89035
R69224 VSS.n2543 VSS.n2440 1.89035
R69225 VSS.n2545 VSS.n2281 1.89035
R69226 VSS.n2543 VSS.n2439 1.89035
R69227 VSS.n2545 VSS.n2280 1.89035
R69228 VSS.n2543 VSS.n2438 1.89035
R69229 VSS.n2545 VSS.n2279 1.89035
R69230 VSS.n2543 VSS.n2437 1.89035
R69231 VSS.n2545 VSS.n2278 1.89035
R69232 VSS.n2543 VSS.n2436 1.89035
R69233 VSS.n2545 VSS.n2277 1.89035
R69234 VSS.n2543 VSS.n2435 1.89035
R69235 VSS.n2545 VSS.n2276 1.89035
R69236 VSS.n2543 VSS.n2434 1.89035
R69237 VSS.n2545 VSS.n2275 1.89035
R69238 VSS.n2543 VSS.n2433 1.89035
R69239 VSS.n2545 VSS.n2274 1.89035
R69240 VSS.n2543 VSS.n2432 1.89035
R69241 VSS.n2545 VSS.n2273 1.89035
R69242 VSS.n2543 VSS.n2431 1.89035
R69243 VSS.n2545 VSS.n2272 1.89035
R69244 VSS.n2543 VSS.n2430 1.89035
R69245 VSS.n2545 VSS.n2271 1.89035
R69246 VSS.n2543 VSS.n2429 1.89035
R69247 VSS.n2545 VSS.n2270 1.89035
R69248 VSS.n2543 VSS.n2428 1.89035
R69249 VSS.n2545 VSS.n2269 1.89035
R69250 VSS.n2543 VSS.n2427 1.89035
R69251 VSS.n2545 VSS.n2268 1.89035
R69252 VSS.n2543 VSS.n2426 1.89035
R69253 VSS.n2545 VSS.n2267 1.89035
R69254 VSS.n2543 VSS.n2425 1.89035
R69255 VSS.n2545 VSS.n2266 1.89035
R69256 VSS.n2543 VSS.n2424 1.89035
R69257 VSS.n2545 VSS.n2265 1.89035
R69258 VSS.n2543 VSS.n2423 1.89035
R69259 VSS.n2545 VSS.n2264 1.89035
R69260 VSS.n2543 VSS.n2422 1.89035
R69261 VSS.n2545 VSS.n2263 1.89035
R69262 VSS.n2543 VSS.n2421 1.89035
R69263 VSS.n2545 VSS.n2262 1.89035
R69264 VSS.n2543 VSS.n2420 1.89035
R69265 VSS.n2545 VSS.n2261 1.89035
R69266 VSS.n2543 VSS.n2230 1.89035
R69267 VSS.n2548 VSS.n2547 1.89035
R69268 VSS.n2543 VSS.n2419 1.89035
R69269 VSS.n2548 VSS.n2228 1.89035
R69270 VSS.n2543 VSS.n2418 1.89035
R69271 VSS.n2548 VSS.n2227 1.89035
R69272 VSS.n2543 VSS.n2417 1.89035
R69273 VSS.n2545 VSS.n2257 1.89035
R69274 VSS.n2543 VSS.n2415 1.89035
R69275 VSS.n2545 VSS.n2256 1.89035
R69276 VSS.n2543 VSS.n2312 1.89035
R69277 VSS.n2545 VSS.n2255 1.89035
R69278 VSS.n2543 VSS.n2311 1.89035
R69279 VSS.n2545 VSS.n2254 1.89035
R69280 VSS.n2543 VSS.n2310 1.89035
R69281 VSS.n2545 VSS.n2253 1.89035
R69282 VSS.n2543 VSS.n2309 1.89035
R69283 VSS.n2545 VSS.n2252 1.89035
R69284 VSS.n2543 VSS.n2308 1.89035
R69285 VSS.n2545 VSS.n2251 1.89035
R69286 VSS.n2543 VSS.n2307 1.89035
R69287 VSS.n2545 VSS.n2250 1.89035
R69288 VSS.n2543 VSS.n2306 1.89035
R69289 VSS.n2545 VSS.n2249 1.89035
R69290 VSS.n2543 VSS.n2305 1.89035
R69291 VSS.n2545 VSS.n2248 1.89035
R69292 VSS.n2543 VSS.n2304 1.89035
R69293 VSS.n2545 VSS.n2247 1.89035
R69294 VSS.n2543 VSS.n2303 1.89035
R69295 VSS.n2545 VSS.n2246 1.89035
R69296 VSS.n2543 VSS.n2302 1.89035
R69297 VSS.n2545 VSS.n2245 1.89035
R69298 VSS.n2543 VSS.n2301 1.89035
R69299 VSS.n2545 VSS.n2244 1.89035
R69300 VSS.n2543 VSS.n2300 1.89035
R69301 VSS.n2545 VSS.n2243 1.89035
R69302 VSS.n2543 VSS.n2299 1.89035
R69303 VSS.n2545 VSS.n2242 1.89035
R69304 VSS.n2543 VSS.n2298 1.89035
R69305 VSS.n2545 VSS.n2241 1.89035
R69306 VSS.n2543 VSS.n2297 1.89035
R69307 VSS.n2545 VSS.n2240 1.89035
R69308 VSS.n2543 VSS.n2296 1.89035
R69309 VSS.n2545 VSS.n2239 1.89035
R69310 VSS.n2543 VSS.n2295 1.89035
R69311 VSS.n2545 VSS.n2238 1.89035
R69312 VSS.n2543 VSS.n2294 1.89035
R69313 VSS.n2545 VSS.n2237 1.89035
R69314 VSS.n2543 VSS.n2293 1.89035
R69315 VSS.n2545 VSS.n2236 1.89035
R69316 VSS.n2543 VSS.n2292 1.89035
R69317 VSS.n2545 VSS.n2235 1.89035
R69318 VSS.n2543 VSS.n2291 1.89035
R69319 VSS.n2545 VSS.n2234 1.89035
R69320 VSS.n2543 VSS.n2290 1.89035
R69321 VSS.n2545 VSS.n2233 1.89035
R69322 VSS.n2543 VSS.n2289 1.89035
R69323 VSS.n2316 VSS.n2315 1.89035
R69324 VSS.n3391 VSS.n3127 1.89035
R69325 VSS.n3162 VSS.n3101 1.89035
R69326 VSS.n3391 VSS.n3126 1.89035
R69327 VSS.n3167 VSS.n3101 1.89035
R69328 VSS.n3391 VSS.n3125 1.89035
R69329 VSS.n3172 VSS.n3101 1.89035
R69330 VSS.n3391 VSS.n3124 1.89035
R69331 VSS.n3177 VSS.n3101 1.89035
R69332 VSS.n3391 VSS.n3123 1.89035
R69333 VSS.n3182 VSS.n3101 1.89035
R69334 VSS.n3391 VSS.n3122 1.89035
R69335 VSS.n3187 VSS.n3101 1.89035
R69336 VSS.n3391 VSS.n3121 1.89035
R69337 VSS.n3192 VSS.n3101 1.89035
R69338 VSS.n3391 VSS.n3120 1.89035
R69339 VSS.n3197 VSS.n3101 1.89035
R69340 VSS.n3391 VSS.n3119 1.89035
R69341 VSS.n3202 VSS.n3101 1.89035
R69342 VSS.n3391 VSS.n3118 1.89035
R69343 VSS.n3207 VSS.n3101 1.89035
R69344 VSS.n3391 VSS.n3117 1.89035
R69345 VSS.n3212 VSS.n3101 1.89035
R69346 VSS.n3391 VSS.n3116 1.89035
R69347 VSS.n3217 VSS.n3101 1.89035
R69348 VSS.n3391 VSS.n3115 1.89035
R69349 VSS.n3222 VSS.n3101 1.89035
R69350 VSS.n3391 VSS.n3114 1.89035
R69351 VSS.n3227 VSS.n3101 1.89035
R69352 VSS.n3391 VSS.n3113 1.89035
R69353 VSS.n3232 VSS.n3101 1.89035
R69354 VSS.n3391 VSS.n3112 1.89035
R69355 VSS.n3237 VSS.n3101 1.89035
R69356 VSS.n3391 VSS.n3111 1.89035
R69357 VSS.n3242 VSS.n3101 1.89035
R69358 VSS.n3391 VSS.n3110 1.89035
R69359 VSS.n3247 VSS.n3101 1.89035
R69360 VSS.n3391 VSS.n3109 1.89035
R69361 VSS.n3252 VSS.n3101 1.89035
R69362 VSS.n3391 VSS.n3108 1.89035
R69363 VSS.n3257 VSS.n3101 1.89035
R69364 VSS.n3391 VSS.n3107 1.89035
R69365 VSS.n3262 VSS.n3101 1.89035
R69366 VSS.n3391 VSS.n3106 1.89035
R69367 VSS.n3276 VSS.n3275 1.89035
R69368 VSS.n3391 VSS.n3105 1.89035
R69369 VSS.n3391 VSS.n3134 1.89035
R69370 VSS.n3277 VSS.n3276 1.89035
R69371 VSS.n3391 VSS.n3135 1.89035
R69372 VSS.n3283 VSS.n3101 1.89035
R69373 VSS.n3391 VSS.n3136 1.89035
R69374 VSS.n3288 VSS.n3101 1.89035
R69375 VSS.n3391 VSS.n3137 1.89035
R69376 VSS.n3293 VSS.n3101 1.89035
R69377 VSS.n3391 VSS.n3138 1.89035
R69378 VSS.n3298 VSS.n3101 1.89035
R69379 VSS.n3391 VSS.n3139 1.89035
R69380 VSS.n3303 VSS.n3101 1.89035
R69381 VSS.n3391 VSS.n3140 1.89035
R69382 VSS.n3308 VSS.n3101 1.89035
R69383 VSS.n3391 VSS.n3141 1.89035
R69384 VSS.n3313 VSS.n3101 1.89035
R69385 VSS.n3391 VSS.n3142 1.89035
R69386 VSS.n3318 VSS.n3101 1.89035
R69387 VSS.n3391 VSS.n3143 1.89035
R69388 VSS.n3323 VSS.n3101 1.89035
R69389 VSS.n3391 VSS.n3144 1.89035
R69390 VSS.n3328 VSS.n3101 1.89035
R69391 VSS.n3391 VSS.n3145 1.89035
R69392 VSS.n3333 VSS.n3101 1.89035
R69393 VSS.n3391 VSS.n3146 1.89035
R69394 VSS.n3338 VSS.n3101 1.89035
R69395 VSS.n3391 VSS.n3147 1.89035
R69396 VSS.n3343 VSS.n3101 1.89035
R69397 VSS.n3391 VSS.n3148 1.89035
R69398 VSS.n3348 VSS.n3101 1.89035
R69399 VSS.n3391 VSS.n3149 1.89035
R69400 VSS.n3353 VSS.n3101 1.89035
R69401 VSS.n3391 VSS.n3150 1.89035
R69402 VSS.n3358 VSS.n3101 1.89035
R69403 VSS.n3391 VSS.n3151 1.89035
R69404 VSS.n3363 VSS.n3101 1.89035
R69405 VSS.n3391 VSS.n3152 1.89035
R69406 VSS.n3368 VSS.n3101 1.89035
R69407 VSS.n3391 VSS.n3153 1.89035
R69408 VSS.n3373 VSS.n3101 1.89035
R69409 VSS.n3391 VSS.n3154 1.89035
R69410 VSS.n3378 VSS.n3101 1.89035
R69411 VSS.n3391 VSS.n3155 1.89035
R69412 VSS.n3383 VSS.n3101 1.89035
R69413 VSS.n3391 VSS.n3156 1.89035
R69414 VSS.n3388 VSS.n3101 1.89035
R69415 VSS.n6194 VSS.n6193 1.73753
R69416 VSS.n564 VSS.n561 1.73383
R69417 VSS.n568 VSS.n561 1.73383
R69418 VSS.n566 VSS.n565 1.73383
R69419 VSS.n567 VSS.n566 1.73383
R69420 VSS.n1829 VSS.n1828 1.6025
R69421 VSS.n1908 VSS.n1907 1.6025
R69422 VSS.n4096 VSS.n538 1.59898
R69423 VSS.n5864 VSS.n5862 1.59898
R69424 VSS.n6156 VSS.n6155 1.59898
R69425 VSS.n5011 VSS.n475 1.59898
R69426 VSS.n1221 VSS.n1220 1.5005
R69427 VSS.n1219 VSS.n1217 1.5005
R69428 VSS.n1892 VSS.n1223 1.5005
R69429 VSS.n20 VSS.n19 1.45763
R69430 VSS.n1613 VSS.n1326 1.44597
R69431 VSS.n5809 VSS.n5808 1.44597
R69432 VSS.n5110 VSS.n5109 1.44597
R69433 VSS.n5099 VSS.n5098 1.44597
R69434 VSS.n5790 VSS.n5079 1.44597
R69435 VSS.n5847 VSS.n4978 1.44597
R69436 VSS.n5469 VSS.n5468 1.44597
R69437 VSS.n5637 VSS.n5256 1.44597
R69438 VSS.n5525 VSS.n5524 1.44597
R69439 VSS.n5518 VSS.n5517 1.44597
R69440 VSS.n5536 VSS.n5535 1.44597
R69441 VSS.n5988 VSS.n4421 1.44597
R69442 VSS.n4818 VSS.n4813 1.44597
R69443 VSS.n4830 VSS.n4825 1.44597
R69444 VSS.n4842 VSS.n4837 1.44597
R69445 VSS.n4854 VSS.n4849 1.44597
R69446 VSS.n4793 VSS.n4791 1.44597
R69447 VSS.n4790 VSS.n4789 1.44597
R69448 VSS.n4784 VSS.n4484 1.44597
R69449 VSS.n4779 VSS.n4777 1.44597
R69450 VSS.n4773 VSS.n4772 1.44597
R69451 VSS.n6134 VSS.n505 1.44597
R69452 VSS.n4237 VSS.n511 1.44597
R69453 VSS.n4243 VSS.n4242 1.44597
R69454 VSS.n4234 VSS.n510 1.44597
R69455 VSS.n520 VSS.n519 1.44597
R69456 VSS.n4224 VSS.n4223 1.44597
R69457 VSS.n4218 VSS.n518 1.44597
R69458 VSS.n531 VSS.n530 1.44597
R69459 VSS.n4208 VSS.n4207 1.44597
R69460 VSS.n4202 VSS.n529 1.44597
R69461 VSS.n4192 VSS.n4190 1.44597
R69462 VSS.n4176 VSS.n4175 1.44597
R69463 VSS.n4170 VSS.n541 1.44597
R69464 VSS.n4165 VSS.n4163 1.44597
R69465 VSS.n4162 VSS.n4161 1.44597
R69466 VSS.n4156 VSS.n545 1.44597
R69467 VSS.n4151 VSS.n4149 1.44597
R69468 VSS.n4148 VSS.n4147 1.44597
R69469 VSS.n4142 VSS.n549 1.44597
R69470 VSS.n4137 VSS.n4135 1.44597
R69471 VSS.n538 VSS.n477 1.43659
R69472 VSS.n5862 VSS.n477 1.43659
R69473 VSS.n6155 VSS.n6154 1.43659
R69474 VSS.n6154 VSS.n475 1.43659
R69475 VSS.n3267 VSS.n3134 1.42229
R69476 VSS.n3278 VSS.n3277 1.42229
R69477 VSS.n3282 VSS.n3135 1.42229
R69478 VSS.n3283 VSS.n3282 1.42229
R69479 VSS.n3287 VSS.n3136 1.42229
R69480 VSS.n3288 VSS.n3287 1.42229
R69481 VSS.n3292 VSS.n3137 1.42229
R69482 VSS.n3293 VSS.n3292 1.42229
R69483 VSS.n3297 VSS.n3138 1.42229
R69484 VSS.n3298 VSS.n3297 1.42229
R69485 VSS.n3302 VSS.n3139 1.42229
R69486 VSS.n3303 VSS.n3302 1.42229
R69487 VSS.n3307 VSS.n3140 1.42229
R69488 VSS.n3308 VSS.n3307 1.42229
R69489 VSS.n3312 VSS.n3141 1.42229
R69490 VSS.n3313 VSS.n3312 1.42229
R69491 VSS.n3317 VSS.n3142 1.42229
R69492 VSS.n3318 VSS.n3317 1.42229
R69493 VSS.n3322 VSS.n3143 1.42229
R69494 VSS.n3323 VSS.n3322 1.42229
R69495 VSS.n3327 VSS.n3144 1.42229
R69496 VSS.n3328 VSS.n3327 1.42229
R69497 VSS.n3332 VSS.n3145 1.42229
R69498 VSS.n3333 VSS.n3332 1.42229
R69499 VSS.n3337 VSS.n3146 1.42229
R69500 VSS.n3338 VSS.n3337 1.42229
R69501 VSS.n3342 VSS.n3147 1.42229
R69502 VSS.n3343 VSS.n3342 1.42229
R69503 VSS.n3347 VSS.n3148 1.42229
R69504 VSS.n3348 VSS.n3347 1.42229
R69505 VSS.n3352 VSS.n3149 1.42229
R69506 VSS.n3353 VSS.n3352 1.42229
R69507 VSS.n3357 VSS.n3150 1.42229
R69508 VSS.n3358 VSS.n3357 1.42229
R69509 VSS.n3362 VSS.n3151 1.42229
R69510 VSS.n3363 VSS.n3362 1.42229
R69511 VSS.n3367 VSS.n3152 1.42229
R69512 VSS.n3368 VSS.n3367 1.42229
R69513 VSS.n3372 VSS.n3153 1.42229
R69514 VSS.n3373 VSS.n3372 1.42229
R69515 VSS.n3377 VSS.n3154 1.42229
R69516 VSS.n3378 VSS.n3377 1.42229
R69517 VSS.n3382 VSS.n3155 1.42229
R69518 VSS.n3383 VSS.n3382 1.42229
R69519 VSS.n3387 VSS.n3156 1.42229
R69520 VSS.n3388 VSS.n3387 1.42229
R69521 VSS.n3161 VSS.n3127 1.42229
R69522 VSS.n3162 VSS.n3161 1.42229
R69523 VSS.n3166 VSS.n3126 1.42229
R69524 VSS.n3167 VSS.n3166 1.42229
R69525 VSS.n3171 VSS.n3125 1.42229
R69526 VSS.n3172 VSS.n3171 1.42229
R69527 VSS.n3176 VSS.n3124 1.42229
R69528 VSS.n3177 VSS.n3176 1.42229
R69529 VSS.n3181 VSS.n3123 1.42229
R69530 VSS.n3182 VSS.n3181 1.42229
R69531 VSS.n3186 VSS.n3122 1.42229
R69532 VSS.n3187 VSS.n3186 1.42229
R69533 VSS.n3191 VSS.n3121 1.42229
R69534 VSS.n3192 VSS.n3191 1.42229
R69535 VSS.n3196 VSS.n3120 1.42229
R69536 VSS.n3197 VSS.n3196 1.42229
R69537 VSS.n3201 VSS.n3119 1.42229
R69538 VSS.n3202 VSS.n3201 1.42229
R69539 VSS.n3206 VSS.n3118 1.42229
R69540 VSS.n3207 VSS.n3206 1.42229
R69541 VSS.n3211 VSS.n3117 1.42229
R69542 VSS.n3212 VSS.n3211 1.42229
R69543 VSS.n3216 VSS.n3116 1.42229
R69544 VSS.n3217 VSS.n3216 1.42229
R69545 VSS.n3221 VSS.n3115 1.42229
R69546 VSS.n3222 VSS.n3221 1.42229
R69547 VSS.n3226 VSS.n3114 1.42229
R69548 VSS.n3227 VSS.n3226 1.42229
R69549 VSS.n3231 VSS.n3113 1.42229
R69550 VSS.n3232 VSS.n3231 1.42229
R69551 VSS.n3236 VSS.n3112 1.42229
R69552 VSS.n3237 VSS.n3236 1.42229
R69553 VSS.n3241 VSS.n3111 1.42229
R69554 VSS.n3242 VSS.n3241 1.42229
R69555 VSS.n3246 VSS.n3110 1.42229
R69556 VSS.n3247 VSS.n3246 1.42229
R69557 VSS.n3251 VSS.n3109 1.42229
R69558 VSS.n3252 VSS.n3251 1.42229
R69559 VSS.n3256 VSS.n3108 1.42229
R69560 VSS.n3257 VSS.n3256 1.42229
R69561 VSS.n3261 VSS.n3107 1.42229
R69562 VSS.n3262 VSS.n3261 1.42229
R69563 VSS.n3270 VSS.n3106 1.42229
R69564 VSS.n3275 VSS.n3269 1.42229
R69565 VSS.n3272 VSS.n3105 1.42229
R69566 VSS.n2540 VSS.n2285 1.42229
R69567 VSS.n2537 VSS.n2443 1.42229
R69568 VSS.n2537 VSS.n2284 1.42229
R69569 VSS.n2533 VSS.n2442 1.42229
R69570 VSS.n2533 VSS.n2283 1.42229
R69571 VSS.n2529 VSS.n2441 1.42229
R69572 VSS.n2529 VSS.n2282 1.42229
R69573 VSS.n2525 VSS.n2440 1.42229
R69574 VSS.n2525 VSS.n2281 1.42229
R69575 VSS.n2521 VSS.n2439 1.42229
R69576 VSS.n2521 VSS.n2280 1.42229
R69577 VSS.n2517 VSS.n2438 1.42229
R69578 VSS.n2517 VSS.n2279 1.42229
R69579 VSS.n2513 VSS.n2437 1.42229
R69580 VSS.n2513 VSS.n2278 1.42229
R69581 VSS.n2509 VSS.n2436 1.42229
R69582 VSS.n2509 VSS.n2277 1.42229
R69583 VSS.n2505 VSS.n2435 1.42229
R69584 VSS.n2505 VSS.n2276 1.42229
R69585 VSS.n2501 VSS.n2434 1.42229
R69586 VSS.n2501 VSS.n2275 1.42229
R69587 VSS.n2497 VSS.n2433 1.42229
R69588 VSS.n2497 VSS.n2274 1.42229
R69589 VSS.n2493 VSS.n2432 1.42229
R69590 VSS.n2493 VSS.n2273 1.42229
R69591 VSS.n2489 VSS.n2431 1.42229
R69592 VSS.n2489 VSS.n2272 1.42229
R69593 VSS.n2485 VSS.n2430 1.42229
R69594 VSS.n2485 VSS.n2271 1.42229
R69595 VSS.n2481 VSS.n2429 1.42229
R69596 VSS.n2481 VSS.n2270 1.42229
R69597 VSS.n2477 VSS.n2428 1.42229
R69598 VSS.n2477 VSS.n2269 1.42229
R69599 VSS.n2473 VSS.n2427 1.42229
R69600 VSS.n2473 VSS.n2268 1.42229
R69601 VSS.n2469 VSS.n2426 1.42229
R69602 VSS.n2469 VSS.n2267 1.42229
R69603 VSS.n2465 VSS.n2425 1.42229
R69604 VSS.n2465 VSS.n2266 1.42229
R69605 VSS.n2461 VSS.n2424 1.42229
R69606 VSS.n2461 VSS.n2265 1.42229
R69607 VSS.n2457 VSS.n2423 1.42229
R69608 VSS.n2457 VSS.n2264 1.42229
R69609 VSS.n2453 VSS.n2422 1.42229
R69610 VSS.n2453 VSS.n2263 1.42229
R69611 VSS.n2449 VSS.n2421 1.42229
R69612 VSS.n2449 VSS.n2262 1.42229
R69613 VSS.n2445 VSS.n2420 1.42229
R69614 VSS.n2445 VSS.n2261 1.42229
R69615 VSS.n2546 VSS.n2230 1.42229
R69616 VSS.n2547 VSS.n2229 1.42229
R69617 VSS.n2419 VSS.n2259 1.42229
R69618 VSS.n2286 VSS.n2228 1.42229
R69619 VSS.n2418 VSS.n2258 1.42229
R69620 VSS.n2287 VSS.n2227 1.42229
R69621 VSS.n2417 VSS.n2416 1.42229
R69622 VSS.n2416 VSS.n2257 1.42229
R69623 VSS.n2415 VSS.n2413 1.42229
R69624 VSS.n2413 VSS.n2256 1.42229
R69625 VSS.n2408 VSS.n2312 1.42229
R69626 VSS.n2408 VSS.n2255 1.42229
R69627 VSS.n2404 VSS.n2311 1.42229
R69628 VSS.n2404 VSS.n2254 1.42229
R69629 VSS.n2400 VSS.n2310 1.42229
R69630 VSS.n2400 VSS.n2253 1.42229
R69631 VSS.n2396 VSS.n2309 1.42229
R69632 VSS.n2396 VSS.n2252 1.42229
R69633 VSS.n2392 VSS.n2308 1.42229
R69634 VSS.n2392 VSS.n2251 1.42229
R69635 VSS.n2388 VSS.n2307 1.42229
R69636 VSS.n2388 VSS.n2250 1.42229
R69637 VSS.n2384 VSS.n2306 1.42229
R69638 VSS.n2384 VSS.n2249 1.42229
R69639 VSS.n2380 VSS.n2305 1.42229
R69640 VSS.n2380 VSS.n2248 1.42229
R69641 VSS.n2376 VSS.n2304 1.42229
R69642 VSS.n2376 VSS.n2247 1.42229
R69643 VSS.n2372 VSS.n2303 1.42229
R69644 VSS.n2372 VSS.n2246 1.42229
R69645 VSS.n2368 VSS.n2302 1.42229
R69646 VSS.n2368 VSS.n2245 1.42229
R69647 VSS.n2364 VSS.n2301 1.42229
R69648 VSS.n2364 VSS.n2244 1.42229
R69649 VSS.n2360 VSS.n2300 1.42229
R69650 VSS.n2360 VSS.n2243 1.42229
R69651 VSS.n2356 VSS.n2299 1.42229
R69652 VSS.n2356 VSS.n2242 1.42229
R69653 VSS.n2352 VSS.n2298 1.42229
R69654 VSS.n2352 VSS.n2241 1.42229
R69655 VSS.n2348 VSS.n2297 1.42229
R69656 VSS.n2348 VSS.n2240 1.42229
R69657 VSS.n2344 VSS.n2296 1.42229
R69658 VSS.n2344 VSS.n2239 1.42229
R69659 VSS.n2340 VSS.n2295 1.42229
R69660 VSS.n2340 VSS.n2238 1.42229
R69661 VSS.n2336 VSS.n2294 1.42229
R69662 VSS.n2336 VSS.n2237 1.42229
R69663 VSS.n2332 VSS.n2293 1.42229
R69664 VSS.n2332 VSS.n2236 1.42229
R69665 VSS.n2328 VSS.n2292 1.42229
R69666 VSS.n2328 VSS.n2235 1.42229
R69667 VSS.n2324 VSS.n2291 1.42229
R69668 VSS.n2324 VSS.n2234 1.42229
R69669 VSS.n2320 VSS.n2290 1.42229
R69670 VSS.n2320 VSS.n2233 1.42229
R69671 VSS.n2289 VSS.n2232 1.42229
R69672 VSS.n2315 VSS.n2288 1.42229
R69673 VSS.n2542 VSS.n2285 1.42229
R69674 VSS.n2540 VSS.n2443 1.42229
R69675 VSS.n2535 VSS.n2442 1.42229
R69676 VSS.n2535 VSS.n2284 1.42229
R69677 VSS.n2531 VSS.n2441 1.42229
R69678 VSS.n2531 VSS.n2283 1.42229
R69679 VSS.n2527 VSS.n2440 1.42229
R69680 VSS.n2527 VSS.n2282 1.42229
R69681 VSS.n2523 VSS.n2439 1.42229
R69682 VSS.n2523 VSS.n2281 1.42229
R69683 VSS.n2519 VSS.n2438 1.42229
R69684 VSS.n2519 VSS.n2280 1.42229
R69685 VSS.n2515 VSS.n2437 1.42229
R69686 VSS.n2515 VSS.n2279 1.42229
R69687 VSS.n2511 VSS.n2436 1.42229
R69688 VSS.n2511 VSS.n2278 1.42229
R69689 VSS.n2507 VSS.n2435 1.42229
R69690 VSS.n2507 VSS.n2277 1.42229
R69691 VSS.n2503 VSS.n2434 1.42229
R69692 VSS.n2503 VSS.n2276 1.42229
R69693 VSS.n2499 VSS.n2433 1.42229
R69694 VSS.n2499 VSS.n2275 1.42229
R69695 VSS.n2495 VSS.n2432 1.42229
R69696 VSS.n2495 VSS.n2274 1.42229
R69697 VSS.n2491 VSS.n2431 1.42229
R69698 VSS.n2491 VSS.n2273 1.42229
R69699 VSS.n2487 VSS.n2430 1.42229
R69700 VSS.n2487 VSS.n2272 1.42229
R69701 VSS.n2483 VSS.n2429 1.42229
R69702 VSS.n2483 VSS.n2271 1.42229
R69703 VSS.n2479 VSS.n2428 1.42229
R69704 VSS.n2479 VSS.n2270 1.42229
R69705 VSS.n2475 VSS.n2427 1.42229
R69706 VSS.n2475 VSS.n2269 1.42229
R69707 VSS.n2471 VSS.n2426 1.42229
R69708 VSS.n2471 VSS.n2268 1.42229
R69709 VSS.n2467 VSS.n2425 1.42229
R69710 VSS.n2467 VSS.n2267 1.42229
R69711 VSS.n2463 VSS.n2424 1.42229
R69712 VSS.n2463 VSS.n2266 1.42229
R69713 VSS.n2459 VSS.n2423 1.42229
R69714 VSS.n2459 VSS.n2265 1.42229
R69715 VSS.n2455 VSS.n2422 1.42229
R69716 VSS.n2455 VSS.n2264 1.42229
R69717 VSS.n2451 VSS.n2421 1.42229
R69718 VSS.n2451 VSS.n2263 1.42229
R69719 VSS.n2447 VSS.n2420 1.42229
R69720 VSS.n2447 VSS.n2262 1.42229
R69721 VSS.n2260 VSS.n2230 1.42229
R69722 VSS.n2261 VSS.n2260 1.42229
R69723 VSS.n2547 VSS.n2546 1.42229
R69724 VSS.n2419 VSS.n2229 1.42229
R69725 VSS.n2259 VSS.n2228 1.42229
R69726 VSS.n2418 VSS.n2286 1.42229
R69727 VSS.n2258 VSS.n2227 1.42229
R69728 VSS.n2417 VSS.n2287 1.42229
R69729 VSS.n2415 VSS.n2414 1.42229
R69730 VSS.n2414 VSS.n2257 1.42229
R69731 VSS.n2410 VSS.n2312 1.42229
R69732 VSS.n2410 VSS.n2256 1.42229
R69733 VSS.n2406 VSS.n2311 1.42229
R69734 VSS.n2406 VSS.n2255 1.42229
R69735 VSS.n2402 VSS.n2310 1.42229
R69736 VSS.n2402 VSS.n2254 1.42229
R69737 VSS.n2398 VSS.n2309 1.42229
R69738 VSS.n2398 VSS.n2253 1.42229
R69739 VSS.n2394 VSS.n2308 1.42229
R69740 VSS.n2394 VSS.n2252 1.42229
R69741 VSS.n2390 VSS.n2307 1.42229
R69742 VSS.n2390 VSS.n2251 1.42229
R69743 VSS.n2386 VSS.n2306 1.42229
R69744 VSS.n2386 VSS.n2250 1.42229
R69745 VSS.n2382 VSS.n2305 1.42229
R69746 VSS.n2382 VSS.n2249 1.42229
R69747 VSS.n2378 VSS.n2304 1.42229
R69748 VSS.n2378 VSS.n2248 1.42229
R69749 VSS.n2374 VSS.n2303 1.42229
R69750 VSS.n2374 VSS.n2247 1.42229
R69751 VSS.n2370 VSS.n2302 1.42229
R69752 VSS.n2370 VSS.n2246 1.42229
R69753 VSS.n2366 VSS.n2301 1.42229
R69754 VSS.n2366 VSS.n2245 1.42229
R69755 VSS.n2362 VSS.n2300 1.42229
R69756 VSS.n2362 VSS.n2244 1.42229
R69757 VSS.n2358 VSS.n2299 1.42229
R69758 VSS.n2358 VSS.n2243 1.42229
R69759 VSS.n2354 VSS.n2298 1.42229
R69760 VSS.n2354 VSS.n2242 1.42229
R69761 VSS.n2350 VSS.n2297 1.42229
R69762 VSS.n2350 VSS.n2241 1.42229
R69763 VSS.n2346 VSS.n2296 1.42229
R69764 VSS.n2346 VSS.n2240 1.42229
R69765 VSS.n2342 VSS.n2295 1.42229
R69766 VSS.n2342 VSS.n2239 1.42229
R69767 VSS.n2338 VSS.n2294 1.42229
R69768 VSS.n2338 VSS.n2238 1.42229
R69769 VSS.n2334 VSS.n2293 1.42229
R69770 VSS.n2334 VSS.n2237 1.42229
R69771 VSS.n2330 VSS.n2292 1.42229
R69772 VSS.n2330 VSS.n2236 1.42229
R69773 VSS.n2326 VSS.n2291 1.42229
R69774 VSS.n2326 VSS.n2235 1.42229
R69775 VSS.n2322 VSS.n2290 1.42229
R69776 VSS.n2322 VSS.n2234 1.42229
R69777 VSS.n2318 VSS.n2289 1.42229
R69778 VSS.n2318 VSS.n2233 1.42229
R69779 VSS.n2315 VSS.n2232 1.42229
R69780 VSS.n3158 VSS.n3127 1.42229
R69781 VSS.n3163 VSS.n3126 1.42229
R69782 VSS.n3163 VSS.n3162 1.42229
R69783 VSS.n3168 VSS.n3125 1.42229
R69784 VSS.n3168 VSS.n3167 1.42229
R69785 VSS.n3173 VSS.n3124 1.42229
R69786 VSS.n3173 VSS.n3172 1.42229
R69787 VSS.n3178 VSS.n3123 1.42229
R69788 VSS.n3178 VSS.n3177 1.42229
R69789 VSS.n3183 VSS.n3122 1.42229
R69790 VSS.n3183 VSS.n3182 1.42229
R69791 VSS.n3188 VSS.n3121 1.42229
R69792 VSS.n3188 VSS.n3187 1.42229
R69793 VSS.n3193 VSS.n3120 1.42229
R69794 VSS.n3193 VSS.n3192 1.42229
R69795 VSS.n3198 VSS.n3119 1.42229
R69796 VSS.n3198 VSS.n3197 1.42229
R69797 VSS.n3203 VSS.n3118 1.42229
R69798 VSS.n3203 VSS.n3202 1.42229
R69799 VSS.n3208 VSS.n3117 1.42229
R69800 VSS.n3208 VSS.n3207 1.42229
R69801 VSS.n3213 VSS.n3116 1.42229
R69802 VSS.n3213 VSS.n3212 1.42229
R69803 VSS.n3218 VSS.n3115 1.42229
R69804 VSS.n3218 VSS.n3217 1.42229
R69805 VSS.n3223 VSS.n3114 1.42229
R69806 VSS.n3223 VSS.n3222 1.42229
R69807 VSS.n3228 VSS.n3113 1.42229
R69808 VSS.n3228 VSS.n3227 1.42229
R69809 VSS.n3233 VSS.n3112 1.42229
R69810 VSS.n3233 VSS.n3232 1.42229
R69811 VSS.n3238 VSS.n3111 1.42229
R69812 VSS.n3238 VSS.n3237 1.42229
R69813 VSS.n3243 VSS.n3110 1.42229
R69814 VSS.n3243 VSS.n3242 1.42229
R69815 VSS.n3248 VSS.n3109 1.42229
R69816 VSS.n3248 VSS.n3247 1.42229
R69817 VSS.n3253 VSS.n3108 1.42229
R69818 VSS.n3253 VSS.n3252 1.42229
R69819 VSS.n3258 VSS.n3107 1.42229
R69820 VSS.n3258 VSS.n3257 1.42229
R69821 VSS.n3263 VSS.n3106 1.42229
R69822 VSS.n3263 VSS.n3262 1.42229
R69823 VSS.n3275 VSS.n3270 1.42229
R69824 VSS.n3269 VSS.n3105 1.42229
R69825 VSS.n3274 VSS.n3134 1.42229
R69826 VSS.n3277 VSS.n3267 1.42229
R69827 VSS.n3278 VSS.n3135 1.42229
R69828 VSS.n3284 VSS.n3136 1.42229
R69829 VSS.n3284 VSS.n3283 1.42229
R69830 VSS.n3289 VSS.n3137 1.42229
R69831 VSS.n3289 VSS.n3288 1.42229
R69832 VSS.n3294 VSS.n3138 1.42229
R69833 VSS.n3294 VSS.n3293 1.42229
R69834 VSS.n3299 VSS.n3139 1.42229
R69835 VSS.n3299 VSS.n3298 1.42229
R69836 VSS.n3304 VSS.n3140 1.42229
R69837 VSS.n3304 VSS.n3303 1.42229
R69838 VSS.n3309 VSS.n3141 1.42229
R69839 VSS.n3309 VSS.n3308 1.42229
R69840 VSS.n3314 VSS.n3142 1.42229
R69841 VSS.n3314 VSS.n3313 1.42229
R69842 VSS.n3319 VSS.n3143 1.42229
R69843 VSS.n3319 VSS.n3318 1.42229
R69844 VSS.n3324 VSS.n3144 1.42229
R69845 VSS.n3324 VSS.n3323 1.42229
R69846 VSS.n3329 VSS.n3145 1.42229
R69847 VSS.n3329 VSS.n3328 1.42229
R69848 VSS.n3334 VSS.n3146 1.42229
R69849 VSS.n3334 VSS.n3333 1.42229
R69850 VSS.n3339 VSS.n3147 1.42229
R69851 VSS.n3339 VSS.n3338 1.42229
R69852 VSS.n3344 VSS.n3148 1.42229
R69853 VSS.n3344 VSS.n3343 1.42229
R69854 VSS.n3349 VSS.n3149 1.42229
R69855 VSS.n3349 VSS.n3348 1.42229
R69856 VSS.n3354 VSS.n3150 1.42229
R69857 VSS.n3354 VSS.n3353 1.42229
R69858 VSS.n3359 VSS.n3151 1.42229
R69859 VSS.n3359 VSS.n3358 1.42229
R69860 VSS.n3364 VSS.n3152 1.42229
R69861 VSS.n3364 VSS.n3363 1.42229
R69862 VSS.n3369 VSS.n3153 1.42229
R69863 VSS.n3369 VSS.n3368 1.42229
R69864 VSS.n3374 VSS.n3154 1.42229
R69865 VSS.n3374 VSS.n3373 1.42229
R69866 VSS.n3379 VSS.n3155 1.42229
R69867 VSS.n3379 VSS.n3378 1.42229
R69868 VSS.n3384 VSS.n3156 1.42229
R69869 VSS.n3384 VSS.n3383 1.42229
R69870 VSS.n3389 VSS.n3388 1.42229
R69871 VSS.n2892 VSS.n2877 1.35477
R69872 VSS.n1132 VSS.n1129 1.35477
R69873 VSS.n3729 VSS.n3727 1.3307
R69874 VSS.n882 VSS.n570 1.3307
R69875 VSS.n3931 VSS.n664 1.3307
R69876 VSS.n2216 VSS.n2149 1.3307
R69877 VSS.n6195 VSS.n6194 1.32884
R69878 VSS.n4101 VSS.n562 1.32884
R69879 VSS.n443 VSS.n442 1.29118
R69880 VSS.n446 VSS.n445 1.29118
R69881 VSS.n6192 VSS.n455 1.19767
R69882 VSS.n3401 VSS.n3400 1.1255
R69883 VSS.n3730 VSS.n3729 1.1255
R69884 VSS.n3439 VSS.n3438 1.1255
R69885 VSS.n3792 VSS.n570 1.1255
R69886 VSS.n3507 VSS.n3506 1.1255
R69887 VSS.n3931 VSS.n3930 1.1255
R69888 VSS.n2685 VSS.n2684 1.1255
R69889 VSS.n2217 VSS.n2216 1.1255
R69890 VSS.n3159 VSS.n3157 1.12321
R69891 VSS.n3159 VSS.n3158 1.11525
R69892 VSS.n4179 VSS.n470 1.10985
R69893 VSS.n4188 VSS.n4187 1.10985
R69894 VSS.n6123 VSS.n481 1.10985
R69895 VSS.n6148 VSS.n6146 1.10985
R69896 VSS.n5500 VSS.n5499 1.10985
R69897 VSS.n5502 VSS.n5488 1.10985
R69898 VSS.n6174 VSS.n6173 1.10691
R69899 VSS.n4184 VSS.n537 1.10691
R69900 VSS.n6126 VSS.n6125 1.10691
R69901 VSS.n6144 VSS.n6143 1.10691
R69902 VSS.n5495 VSS.n5494 1.10691
R69903 VSS.n5487 VSS.n4946 1.10691
R69904 VSS.n3391 VSS.n3128 1.03912
R69905 VSS.n6236 VSS.n6224 1.00453
R69906 VSS.n3729 VSS.n3728 0.9896
R69907 VSS.n2216 VSS.n2215 0.9896
R69908 VSS.n4126 DVSS 0.979316
R69909 VSS.n2745 VSS.n738 0.954735
R69910 VSS.n4116 VSS.n570 0.95135
R69911 VSS.n3932 VSS.n3931 0.95135
R69912 VSS.n3402 VSS.n3401 0.9356
R69913 VSS.n3438 VSS.n3437 0.9356
R69914 VSS.n3507 VSS.n968 0.9356
R69915 VSS.n2686 VSS.n2685 0.9356
R69916 VSS.n2979 VSS.n1101 0.928878
R69917 VSS.n2983 VSS.n2981 0.928878
R69918 VSS.n2940 VSS.n2938 0.928878
R69919 VSS.n2943 VSS.n2942 0.928878
R69920 VSS.n3391 VSS.n3390 0.903572
R69921 VSS.n6224 VSS.n124 0.902201
R69922 VSS.n4127 VSS.n4126 0.9005
R69923 VSS.n455 DVSS 0.885578
R69924 VSS.n4123 DVSS 0.885578
R69925 VSS.n564 DVSS 0.884579
R69926 VSS.n565 DVSS 0.884579
R69927 VSS.n4125 DVSS 0.884579
R69928 VSS.n4124 DVSS 0.884579
R69929 VSS.n1835 VSS.n1834 0.88295
R69930 VSS.n1748 VSS.n1747 0.88295
R69931 VSS.n1544 VSS.n1543 0.88295
R69932 VSS.n1595 VSS.n1209 0.88295
R69933 VSS.n3066 VSS.n3065 0.8825
R69934 VSS.n2778 VSS.n2777 0.8825
R69935 VSS.n2871 VSS.n2870 0.8825
R69936 VSS.n2057 VSS.n2056 0.8825
R69937 VSS.n560 DVSS 0.835841
R69938 VSS.n6237 VSS.n6236 0.800919
R69939 VSS.n2915 VSS.n2914 0.791851
R69940 VSS.n2960 VSS.n1094 0.791851
R69941 VSS.n1140 VSS.n1139 0.791851
R69942 VSS.n2910 VSS.n1146 0.791851
R69943 VSS.n4123 VSS.n4122 0.786676
R69944 VSS.n3160 VSS.n3159 0.764199
R69945 VSS.n6460 VSS.n6459 0.763161
R69946 VSS.n439 VSS.n438 0.763161
R69947 VSS.n2960 VSS.n2959 0.743357
R69948 VSS.n2959 VSS.n2958 0.743357
R69949 VSS.n2906 VSS.n2879 0.743357
R69950 VSS.n2912 VSS.n2879 0.743357
R69951 VSS.n2914 VSS.n2913 0.743357
R69952 VSS.n2913 VSS.n2912 0.743357
R69953 VSS.n1130 VSS.n1123 0.743357
R69954 VSS.n2958 VSS.n1130 0.743357
R69955 VSS.n2908 VSS.n2878 0.743357
R69956 VSS.n2912 VSS.n2878 0.743357
R69957 VSS.n1139 VSS.n1128 0.743357
R69958 VSS.n2958 VSS.n1128 0.743357
R69959 VSS.n2957 VSS.n2956 0.743357
R69960 VSS.n2958 VSS.n2957 0.743357
R69961 VSS.n2911 VSS.n2910 0.743357
R69962 VSS.n2912 VSS.n2911 0.743357
R69963 VSS.n3273 VSS.n3272 0.686775
R69964 VSS.n2544 VSS.n2288 0.685361
R69965 VSS.n6217 VSS.n6216 0.670023
R69966 VSS.n6447 VSS.n19 0.661953
R69967 VSS.n4122 VSS.n560 0.564324
R69968 VSS.n3924 DVSS 0.557375
R69969 VSS.n3924 DVSS 0.557375
R69970 VSS.n733 DVSS 0.557375
R69971 VSS.n733 DVSS 0.557375
R69972 VSS.n3798 DVSS 0.557375
R69973 VSS.n3798 DVSS 0.557375
R69974 VSS.n4130 VSS.n458 0.555174
R69975 VSS.n4133 VSS.n558 0.555174
R69976 VSS.n5833 VSS.n5832 0.555174
R69977 VSS.n5830 VSS.n5023 0.555174
R69978 VSS.n6159 VSS.n457 0.553707
R69979 VSS.n4095 VSS.n4094 0.553707
R69980 VSS.n5837 VSS.n5835 0.553707
R69981 VSS.n5800 VSS.n4944 0.553707
R69982 VSS.n2931 VSS.n1154 0.548638
R69983 VSS.n2898 VSS.n1134 0.548638
R69984 VSS.n2927 VSS.n1118 0.548638
R69985 VSS.n2965 VSS.n2964 0.548638
R69986 VSS.n2935 VSS.n1151 0.548638
R69987 VSS.n2948 VSS.n1136 0.548638
R69988 VSS.n565 VSS.n564 0.545794
R69989 VSS.n565 VSS.n455 0.545794
R69990 VSS.n4125 VSS.n4124 0.545794
R69991 VSS.n4124 VSS.n4123 0.545794
R69992 VSS.n4100 VSS.n4099 0.5072
R69993 VSS.n4103 VSS.n573 0.5072
R69994 VSS.n6191 VSS.n6190 0.5072
R69995 VSS.n6157 VSS.n454 0.5072
R69996 VSS.n1859 VSS.n1858 0.5005
R69997 VSS.n1857 VSS.n1856 0.5005
R69998 VSS.n1863 VSS.n1855 0.5005
R69999 VSS.n1864 VSS.n1854 0.5005
R70000 VSS.n1865 VSS.n1853 0.5005
R70001 VSS.n1852 VSS.n1850 0.5005
R70002 VSS.n1869 VSS.n1849 0.5005
R70003 VSS.n1870 VSS.n1848 0.5005
R70004 VSS.n1871 VSS.n1847 0.5005
R70005 VSS.n1846 VSS.n1844 0.5005
R70006 VSS.n1875 VSS.n1843 0.5005
R70007 VSS.n1876 VSS.n1842 0.5005
R70008 VSS.n1877 VSS.n1841 0.5005
R70009 VSS.n1592 VSS.n1553 0.5005
R70010 VSS.n1591 VSS.n1554 0.5005
R70011 VSS.n1590 VSS.n1555 0.5005
R70012 VSS.n1558 VSS.n1556 0.5005
R70013 VSS.n1586 VSS.n1559 0.5005
R70014 VSS.n1585 VSS.n1560 0.5005
R70015 VSS.n1584 VSS.n1561 0.5005
R70016 VSS.n1564 VSS.n1562 0.5005
R70017 VSS.n1580 VSS.n1565 0.5005
R70018 VSS.n1579 VSS.n1566 0.5005
R70019 VSS.n1578 VSS.n1567 0.5005
R70020 VSS.n1570 VSS.n1568 0.5005
R70021 VSS.n1574 VSS.n1571 0.5005
R70022 VSS.n1573 VSS.n1572 0.5005
R70023 VSS.n1345 VSS.n1344 0.5005
R70024 VSS.n1620 VSS.n1619 0.5005
R70025 VSS.n1621 VSS.n1343 0.5005
R70026 VSS.n1623 VSS.n1622 0.5005
R70027 VSS.n1341 VSS.n1340 0.5005
R70028 VSS.n1628 VSS.n1627 0.5005
R70029 VSS.n1629 VSS.n1339 0.5005
R70030 VSS.n1631 VSS.n1630 0.5005
R70031 VSS.n1337 VSS.n1336 0.5005
R70032 VSS.n1636 VSS.n1635 0.5005
R70033 VSS.n1637 VSS.n1335 0.5005
R70034 VSS.n1639 VSS.n1638 0.5005
R70035 VSS.n1333 VSS.n1332 0.5005
R70036 VSS.n1644 VSS.n1643 0.5005
R70037 VSS.n1645 VSS.n1331 0.5005
R70038 VSS.n1647 VSS.n1646 0.5005
R70039 VSS.n1329 VSS.n1328 0.5005
R70040 VSS.n1653 VSS.n1652 0.5005
R70041 VSS.n1654 VSS.n1327 0.5005
R70042 VSS.n1658 VSS.n1655 0.5005
R70043 VSS.n1657 VSS.n1656 0.5005
R70044 VSS.n1305 VSS.n1304 0.5005
R70045 VSS.n1667 VSS.n1666 0.5005
R70046 VSS.n1668 VSS.n1303 0.5005
R70047 VSS.n1670 VSS.n1669 0.5005
R70048 VSS.n1301 VSS.n1300 0.5005
R70049 VSS.n1675 VSS.n1674 0.5005
R70050 VSS.n1676 VSS.n1299 0.5005
R70051 VSS.n1678 VSS.n1677 0.5005
R70052 VSS.n1297 VSS.n1296 0.5005
R70053 VSS.n1683 VSS.n1682 0.5005
R70054 VSS.n1684 VSS.n1295 0.5005
R70055 VSS.n1686 VSS.n1685 0.5005
R70056 VSS.n1293 VSS.n1292 0.5005
R70057 VSS.n1691 VSS.n1690 0.5005
R70058 VSS.n1692 VSS.n1291 0.5005
R70059 VSS.n1737 VSS.n1693 0.5005
R70060 VSS.n1736 VSS.n1694 0.5005
R70061 VSS.n1735 VSS.n1695 0.5005
R70062 VSS.n1734 VSS.n1696 0.5005
R70063 VSS.n1699 VSS.n1697 0.5005
R70064 VSS.n1730 VSS.n1700 0.5005
R70065 VSS.n1729 VSS.n1701 0.5005
R70066 VSS.n1728 VSS.n1702 0.5005
R70067 VSS.n1705 VSS.n1703 0.5005
R70068 VSS.n1724 VSS.n1706 0.5005
R70069 VSS.n1723 VSS.n1707 0.5005
R70070 VSS.n1722 VSS.n1708 0.5005
R70071 VSS.n1711 VSS.n1709 0.5005
R70072 VSS.n1718 VSS.n1712 0.5005
R70073 VSS.n1717 VSS.n1713 0.5005
R70074 VSS.n1716 VSS.n1714 0.5005
R70075 VSS.n1244 VSS.n1243 0.5005
R70076 VSS.n1839 VSS.n1838 0.5005
R70077 VSS.n1840 VSS.n1242 0.5005
R70078 VSS.n1861 VSS.n1856 0.5005
R70079 VSS.n1863 VSS.n1862 0.5005
R70080 VSS.n1864 VSS.n1851 0.5005
R70081 VSS.n1866 VSS.n1865 0.5005
R70082 VSS.n1867 VSS.n1850 0.5005
R70083 VSS.n1869 VSS.n1868 0.5005
R70084 VSS.n1870 VSS.n1845 0.5005
R70085 VSS.n1872 VSS.n1871 0.5005
R70086 VSS.n1873 VSS.n1844 0.5005
R70087 VSS.n1875 VSS.n1874 0.5005
R70088 VSS.n1876 VSS.n1241 0.5005
R70089 VSS.n1878 VSS.n1877 0.5005
R70090 VSS.n1551 VSS.n1549 0.5005
R70091 VSS.n1593 VSS.n1592 0.5005
R70092 VSS.n1591 VSS.n1550 0.5005
R70093 VSS.n1590 VSS.n1589 0.5005
R70094 VSS.n1588 VSS.n1556 0.5005
R70095 VSS.n1587 VSS.n1586 0.5005
R70096 VSS.n1585 VSS.n1557 0.5005
R70097 VSS.n1584 VSS.n1583 0.5005
R70098 VSS.n1582 VSS.n1562 0.5005
R70099 VSS.n1581 VSS.n1580 0.5005
R70100 VSS.n1579 VSS.n1563 0.5005
R70101 VSS.n1578 VSS.n1577 0.5005
R70102 VSS.n1576 VSS.n1568 0.5005
R70103 VSS.n1575 VSS.n1574 0.5005
R70104 VSS.n1573 VSS.n1569 0.5005
R70105 VSS.n1346 VSS.n1345 0.5005
R70106 VSS.n1619 VSS.n1618 0.5005
R70107 VSS.n1546 VSS.n1343 0.5005
R70108 VSS.n1624 VSS.n1623 0.5005
R70109 VSS.n1625 VSS.n1341 0.5005
R70110 VSS.n1627 VSS.n1626 0.5005
R70111 VSS.n1339 VSS.n1338 0.5005
R70112 VSS.n1632 VSS.n1631 0.5005
R70113 VSS.n1633 VSS.n1337 0.5005
R70114 VSS.n1635 VSS.n1634 0.5005
R70115 VSS.n1335 VSS.n1334 0.5005
R70116 VSS.n1640 VSS.n1639 0.5005
R70117 VSS.n1641 VSS.n1333 0.5005
R70118 VSS.n1643 VSS.n1642 0.5005
R70119 VSS.n1331 VSS.n1330 0.5005
R70120 VSS.n1648 VSS.n1647 0.5005
R70121 VSS.n1649 VSS.n1329 0.5005
R70122 VSS.n1652 VSS.n1651 0.5005
R70123 VSS.n1650 VSS.n1327 0.5005
R70124 VSS.n1659 VSS.n1658 0.5005
R70125 VSS.n1657 VSS.n1306 0.5005
R70126 VSS.n1664 VSS.n1305 0.5005
R70127 VSS.n1666 VSS.n1665 0.5005
R70128 VSS.n1303 VSS.n1302 0.5005
R70129 VSS.n1671 VSS.n1670 0.5005
R70130 VSS.n1672 VSS.n1301 0.5005
R70131 VSS.n1674 VSS.n1673 0.5005
R70132 VSS.n1299 VSS.n1298 0.5005
R70133 VSS.n1679 VSS.n1678 0.5005
R70134 VSS.n1680 VSS.n1297 0.5005
R70135 VSS.n1682 VSS.n1681 0.5005
R70136 VSS.n1295 VSS.n1294 0.5005
R70137 VSS.n1687 VSS.n1686 0.5005
R70138 VSS.n1688 VSS.n1293 0.5005
R70139 VSS.n1690 VSS.n1689 0.5005
R70140 VSS.n1291 VSS.n1290 0.5005
R70141 VSS.n1738 VSS.n1737 0.5005
R70142 VSS.n1736 VSS.n1284 0.5005
R70143 VSS.n1735 VSS.n1285 0.5005
R70144 VSS.n1734 VSS.n1733 0.5005
R70145 VSS.n1732 VSS.n1697 0.5005
R70146 VSS.n1731 VSS.n1730 0.5005
R70147 VSS.n1729 VSS.n1698 0.5005
R70148 VSS.n1728 VSS.n1727 0.5005
R70149 VSS.n1726 VSS.n1703 0.5005
R70150 VSS.n1725 VSS.n1724 0.5005
R70151 VSS.n1723 VSS.n1704 0.5005
R70152 VSS.n1722 VSS.n1721 0.5005
R70153 VSS.n1720 VSS.n1709 0.5005
R70154 VSS.n1719 VSS.n1718 0.5005
R70155 VSS.n1717 VSS.n1710 0.5005
R70156 VSS.n1716 VSS.n1715 0.5005
R70157 VSS.n1245 VSS.n1244 0.5005
R70158 VSS.n1838 VSS.n1837 0.5005
R70159 VSS.n1242 VSS.n1236 0.5005
R70160 VSS.n924 VSS.n923 0.496843
R70161 VSS.n437 VSS.n436 0.461183
R70162 VSS.n6445 VSS.n6444 0.455549
R70163 VSS.n6242 VSS.n6238 0.455549
R70164 VSS.n6461 VSS.n3 0.455549
R70165 VSS.n1797 VSS.n1796 0.4505
R70166 VSS.n1799 VSS.n1798 0.4505
R70167 VSS.n1794 VSS.n1793 0.4505
R70168 VSS.n1804 VSS.n1803 0.4505
R70169 VSS.n1805 VSS.n1792 0.4505
R70170 VSS.n1807 VSS.n1806 0.4505
R70171 VSS.n1790 VSS.n1789 0.4505
R70172 VSS.n1812 VSS.n1811 0.4505
R70173 VSS.n1813 VSS.n1787 0.4505
R70174 VSS.n1815 VSS.n1814 0.4505
R70175 VSS.n1788 VSS.n1785 0.4505
R70176 VSS.n1819 VSS.n1784 0.4505
R70177 VSS.n1821 VSS.n1820 0.4505
R70178 VSS.n1377 VSS.n1376 0.4505
R70179 VSS.n1379 VSS.n1378 0.4505
R70180 VSS.n1374 VSS.n1373 0.4505
R70181 VSS.n1384 VSS.n1383 0.4505
R70182 VSS.n1385 VSS.n1372 0.4505
R70183 VSS.n1387 VSS.n1386 0.4505
R70184 VSS.n1370 VSS.n1369 0.4505
R70185 VSS.n1392 VSS.n1391 0.4505
R70186 VSS.n1393 VSS.n1368 0.4505
R70187 VSS.n1395 VSS.n1394 0.4505
R70188 VSS.n1366 VSS.n1365 0.4505
R70189 VSS.n1400 VSS.n1399 0.4505
R70190 VSS.n1401 VSS.n1364 0.4505
R70191 VSS.n1403 VSS.n1402 0.4505
R70192 VSS.n1362 VSS.n1361 0.4505
R70193 VSS.n1408 VSS.n1407 0.4505
R70194 VSS.n1409 VSS.n1359 0.4505
R70195 VSS.n1530 VSS.n1529 0.4505
R70196 VSS.n1528 VSS.n1360 0.4505
R70197 VSS.n1527 VSS.n1526 0.4505
R70198 VSS.n1411 VSS.n1410 0.4505
R70199 VSS.n1522 VSS.n1521 0.4505
R70200 VSS.n1520 VSS.n1413 0.4505
R70201 VSS.n1519 VSS.n1518 0.4505
R70202 VSS.n1415 VSS.n1414 0.4505
R70203 VSS.n1514 VSS.n1513 0.4505
R70204 VSS.n1512 VSS.n1417 0.4505
R70205 VSS.n1511 VSS.n1510 0.4505
R70206 VSS.n1419 VSS.n1418 0.4505
R70207 VSS.n1506 VSS.n1505 0.4505
R70208 VSS.n1504 VSS.n1421 0.4505
R70209 VSS.n1503 VSS.n1502 0.4505
R70210 VSS.n1423 VSS.n1422 0.4505
R70211 VSS.n1441 VSS.n1440 0.4505
R70212 VSS.n1442 VSS.n1438 0.4505
R70213 VSS.n1488 VSS.n1487 0.4505
R70214 VSS.n1486 VSS.n1439 0.4505
R70215 VSS.n1485 VSS.n1484 0.4505
R70216 VSS.n1444 VSS.n1443 0.4505
R70217 VSS.n1480 VSS.n1479 0.4505
R70218 VSS.n1478 VSS.n1446 0.4505
R70219 VSS.n1477 VSS.n1476 0.4505
R70220 VSS.n1448 VSS.n1447 0.4505
R70221 VSS.n1472 VSS.n1471 0.4505
R70222 VSS.n1470 VSS.n1450 0.4505
R70223 VSS.n1469 VSS.n1468 0.4505
R70224 VSS.n1452 VSS.n1451 0.4505
R70225 VSS.n1464 VSS.n1463 0.4505
R70226 VSS.n1462 VSS.n1454 0.4505
R70227 VSS.n1461 VSS.n1460 0.4505
R70228 VSS.n1458 VSS.n1455 0.4505
R70229 VSS.n1457 VSS.n1456 0.4505
R70230 VSS.n1273 VSS.n1272 0.4505
R70231 VSS.n1758 VSS.n1757 0.4505
R70232 VSS.n1759 VSS.n1271 0.4505
R70233 VSS.n1761 VSS.n1760 0.4505
R70234 VSS.n1269 VSS.n1268 0.4505
R70235 VSS.n1766 VSS.n1765 0.4505
R70236 VSS.n1767 VSS.n1267 0.4505
R70237 VSS.n1769 VSS.n1768 0.4505
R70238 VSS.n1265 VSS.n1264 0.4505
R70239 VSS.n1774 VSS.n1773 0.4505
R70240 VSS.n1775 VSS.n1263 0.4505
R70241 VSS.n1777 VSS.n1776 0.4505
R70242 VSS.n1261 VSS.n1260 0.4505
R70243 VSS.n1782 VSS.n1781 0.4505
R70244 VSS.n1783 VSS.n1258 0.4505
R70245 VSS.n1824 VSS.n1823 0.4505
R70246 VSS.n1822 VSS.n1259 0.4505
R70247 VSS.n1800 VSS.n1799 0.4505
R70248 VSS.n1801 VSS.n1794 0.4505
R70249 VSS.n1803 VSS.n1802 0.4505
R70250 VSS.n1792 VSS.n1791 0.4505
R70251 VSS.n1808 VSS.n1807 0.4505
R70252 VSS.n1809 VSS.n1790 0.4505
R70253 VSS.n1811 VSS.n1810 0.4505
R70254 VSS.n1787 VSS.n1786 0.4505
R70255 VSS.n1816 VSS.n1815 0.4505
R70256 VSS.n1817 VSS.n1785 0.4505
R70257 VSS.n1819 VSS.n1818 0.4505
R70258 VSS.n1820 VSS.n1252 0.4505
R70259 VSS.n1375 VSS.n1200 0.4505
R70260 VSS.n1376 VSS.n1205 0.4505
R70261 VSS.n1380 VSS.n1379 0.4505
R70262 VSS.n1381 VSS.n1374 0.4505
R70263 VSS.n1383 VSS.n1382 0.4505
R70264 VSS.n1372 VSS.n1371 0.4505
R70265 VSS.n1388 VSS.n1387 0.4505
R70266 VSS.n1389 VSS.n1370 0.4505
R70267 VSS.n1391 VSS.n1390 0.4505
R70268 VSS.n1368 VSS.n1367 0.4505
R70269 VSS.n1396 VSS.n1395 0.4505
R70270 VSS.n1397 VSS.n1366 0.4505
R70271 VSS.n1399 VSS.n1398 0.4505
R70272 VSS.n1364 VSS.n1363 0.4505
R70273 VSS.n1404 VSS.n1403 0.4505
R70274 VSS.n1405 VSS.n1362 0.4505
R70275 VSS.n1407 VSS.n1406 0.4505
R70276 VSS.n1359 VSS.n1356 0.4505
R70277 VSS.n1531 VSS.n1530 0.4505
R70278 VSS.n1360 VSS.n1358 0.4505
R70279 VSS.n1526 VSS.n1525 0.4505
R70280 VSS.n1524 VSS.n1411 0.4505
R70281 VSS.n1523 VSS.n1522 0.4505
R70282 VSS.n1413 VSS.n1412 0.4505
R70283 VSS.n1518 VSS.n1517 0.4505
R70284 VSS.n1516 VSS.n1415 0.4505
R70285 VSS.n1515 VSS.n1514 0.4505
R70286 VSS.n1417 VSS.n1416 0.4505
R70287 VSS.n1510 VSS.n1509 0.4505
R70288 VSS.n1508 VSS.n1419 0.4505
R70289 VSS.n1507 VSS.n1506 0.4505
R70290 VSS.n1421 VSS.n1420 0.4505
R70291 VSS.n1502 VSS.n1501 0.4505
R70292 VSS.n1500 VSS.n1423 0.4505
R70293 VSS.n1440 VSS.n1426 0.4505
R70294 VSS.n1438 VSS.n1433 0.4505
R70295 VSS.n1489 VSS.n1488 0.4505
R70296 VSS.n1439 VSS.n1437 0.4505
R70297 VSS.n1484 VSS.n1483 0.4505
R70298 VSS.n1482 VSS.n1444 0.4505
R70299 VSS.n1481 VSS.n1480 0.4505
R70300 VSS.n1446 VSS.n1445 0.4505
R70301 VSS.n1476 VSS.n1475 0.4505
R70302 VSS.n1474 VSS.n1448 0.4505
R70303 VSS.n1473 VSS.n1472 0.4505
R70304 VSS.n1450 VSS.n1449 0.4505
R70305 VSS.n1468 VSS.n1467 0.4505
R70306 VSS.n1466 VSS.n1452 0.4505
R70307 VSS.n1465 VSS.n1464 0.4505
R70308 VSS.n1454 VSS.n1453 0.4505
R70309 VSS.n1460 VSS.n1459 0.4505
R70310 VSS.n1458 VSS.n1282 0.4505
R70311 VSS.n1457 VSS.n1274 0.4505
R70312 VSS.n1755 VSS.n1273 0.4505
R70313 VSS.n1757 VSS.n1756 0.4505
R70314 VSS.n1271 VSS.n1270 0.4505
R70315 VSS.n1762 VSS.n1761 0.4505
R70316 VSS.n1763 VSS.n1269 0.4505
R70317 VSS.n1765 VSS.n1764 0.4505
R70318 VSS.n1267 VSS.n1266 0.4505
R70319 VSS.n1770 VSS.n1769 0.4505
R70320 VSS.n1771 VSS.n1265 0.4505
R70321 VSS.n1773 VSS.n1772 0.4505
R70322 VSS.n1263 VSS.n1262 0.4505
R70323 VSS.n1778 VSS.n1777 0.4505
R70324 VSS.n1779 VSS.n1261 0.4505
R70325 VSS.n1781 VSS.n1780 0.4505
R70326 VSS.n1258 VSS.n1257 0.4505
R70327 VSS.n1825 VSS.n1824 0.4505
R70328 VSS.n1259 VSS.n1250 0.4505
R70329 VSS.n3036 VSS.n3035 0.4505
R70330 VSS.n3038 VSS.n3037 0.4505
R70331 VSS.n3033 VSS.n3032 0.4505
R70332 VSS.n3043 VSS.n3042 0.4505
R70333 VSS.n3044 VSS.n3031 0.4505
R70334 VSS.n3046 VSS.n3045 0.4505
R70335 VSS.n3029 VSS.n3028 0.4505
R70336 VSS.n3051 VSS.n3050 0.4505
R70337 VSS.n3052 VSS.n3027 0.4505
R70338 VSS.n3054 VSS.n3053 0.4505
R70339 VSS.n3024 VSS.n3023 0.4505
R70340 VSS.n3059 VSS.n3058 0.4505
R70341 VSS.n3060 VSS.n1062 0.4505
R70342 VSS.n2053 VSS.n2052 0.4505
R70343 VSS.n2051 VSS.n1194 0.4505
R70344 VSS.n2050 VSS.n2049 0.4505
R70345 VSS.n1912 VSS.n1911 0.4505
R70346 VSS.n2045 VSS.n2044 0.4505
R70347 VSS.n2043 VSS.n1914 0.4505
R70348 VSS.n2042 VSS.n2041 0.4505
R70349 VSS.n1916 VSS.n1915 0.4505
R70350 VSS.n2037 VSS.n2036 0.4505
R70351 VSS.n2035 VSS.n1918 0.4505
R70352 VSS.n2034 VSS.n2033 0.4505
R70353 VSS.n1920 VSS.n1919 0.4505
R70354 VSS.n2029 VSS.n2028 0.4505
R70355 VSS.n2027 VSS.n1922 0.4505
R70356 VSS.n2026 VSS.n2025 0.4505
R70357 VSS.n2022 VSS.n1923 0.4505
R70358 VSS.n2021 VSS.n2019 0.4505
R70359 VSS.n2018 VSS.n1924 0.4505
R70360 VSS.n2017 VSS.n2016 0.4505
R70361 VSS.n1926 VSS.n1925 0.4505
R70362 VSS.n2012 VSS.n2011 0.4505
R70363 VSS.n2010 VSS.n1929 0.4505
R70364 VSS.n2009 VSS.n2008 0.4505
R70365 VSS.n1931 VSS.n1930 0.4505
R70366 VSS.n2004 VSS.n2003 0.4505
R70367 VSS.n2002 VSS.n1933 0.4505
R70368 VSS.n2001 VSS.n2000 0.4505
R70369 VSS.n1935 VSS.n1934 0.4505
R70370 VSS.n1996 VSS.n1995 0.4505
R70371 VSS.n1994 VSS.n1937 0.4505
R70372 VSS.n1993 VSS.n1992 0.4505
R70373 VSS.n1939 VSS.n1938 0.4505
R70374 VSS.n1988 VSS.n1987 0.4505
R70375 VSS.n1986 VSS.n1941 0.4505
R70376 VSS.n1985 VSS.n1984 0.4505
R70377 VSS.n1983 VSS.n1942 0.4505
R70378 VSS.n1946 VSS.n1943 0.4505
R70379 VSS.n1979 VSS.n1978 0.4505
R70380 VSS.n1977 VSS.n1945 0.4505
R70381 VSS.n1976 VSS.n1975 0.4505
R70382 VSS.n1948 VSS.n1947 0.4505
R70383 VSS.n1971 VSS.n1970 0.4505
R70384 VSS.n1969 VSS.n1950 0.4505
R70385 VSS.n1968 VSS.n1967 0.4505
R70386 VSS.n1952 VSS.n1951 0.4505
R70387 VSS.n1963 VSS.n1962 0.4505
R70388 VSS.n1961 VSS.n1954 0.4505
R70389 VSS.n1960 VSS.n1959 0.4505
R70390 VSS.n1956 VSS.n1955 0.4505
R70391 VSS.n1080 VSS.n1079 0.4505
R70392 VSS.n2989 VSS.n2988 0.4505
R70393 VSS.n2990 VSS.n1078 0.4505
R70394 VSS.n2992 VSS.n2991 0.4505
R70395 VSS.n1076 VSS.n1075 0.4505
R70396 VSS.n2997 VSS.n2996 0.4505
R70397 VSS.n2998 VSS.n1074 0.4505
R70398 VSS.n3000 VSS.n2999 0.4505
R70399 VSS.n1072 VSS.n1071 0.4505
R70400 VSS.n3005 VSS.n3004 0.4505
R70401 VSS.n3006 VSS.n1070 0.4505
R70402 VSS.n3008 VSS.n3007 0.4505
R70403 VSS.n1068 VSS.n1067 0.4505
R70404 VSS.n3013 VSS.n3012 0.4505
R70405 VSS.n3014 VSS.n1066 0.4505
R70406 VSS.n3016 VSS.n3015 0.4505
R70407 VSS.n1064 VSS.n1063 0.4505
R70408 VSS.n3021 VSS.n3020 0.4505
R70409 VSS.n3022 VSS.n1061 0.4505
R70410 VSS.n3062 VSS.n3061 0.4505
R70411 VSS.n3039 VSS.n3038 0.4505
R70412 VSS.n3040 VSS.n3033 0.4505
R70413 VSS.n3042 VSS.n3041 0.4505
R70414 VSS.n3031 VSS.n3030 0.4505
R70415 VSS.n3047 VSS.n3046 0.4505
R70416 VSS.n3048 VSS.n3029 0.4505
R70417 VSS.n3050 VSS.n3049 0.4505
R70418 VSS.n3027 VSS.n3026 0.4505
R70419 VSS.n3055 VSS.n3054 0.4505
R70420 VSS.n3056 VSS.n3024 0.4505
R70421 VSS.n3058 VSS.n3057 0.4505
R70422 VSS.n3025 VSS.n1062 0.4505
R70423 VSS.n1193 VSS.n1186 0.4505
R70424 VSS.n2054 VSS.n2053 0.4505
R70425 VSS.n1194 VSS.n1192 0.4505
R70426 VSS.n2049 VSS.n2048 0.4505
R70427 VSS.n2047 VSS.n1912 0.4505
R70428 VSS.n2046 VSS.n2045 0.4505
R70429 VSS.n1914 VSS.n1913 0.4505
R70430 VSS.n2041 VSS.n2040 0.4505
R70431 VSS.n2039 VSS.n1916 0.4505
R70432 VSS.n2038 VSS.n2037 0.4505
R70433 VSS.n1918 VSS.n1917 0.4505
R70434 VSS.n2033 VSS.n2032 0.4505
R70435 VSS.n2031 VSS.n1920 0.4505
R70436 VSS.n2030 VSS.n2029 0.4505
R70437 VSS.n1922 VSS.n1921 0.4505
R70438 VSS.n2025 VSS.n2024 0.4505
R70439 VSS.n2023 VSS.n2022 0.4505
R70440 VSS.n2021 VSS.n2020 0.4505
R70441 VSS.n1927 VSS.n1924 0.4505
R70442 VSS.n2016 VSS.n2015 0.4505
R70443 VSS.n2014 VSS.n1926 0.4505
R70444 VSS.n2013 VSS.n2012 0.4505
R70445 VSS.n1929 VSS.n1928 0.4505
R70446 VSS.n2008 VSS.n2007 0.4505
R70447 VSS.n2006 VSS.n1931 0.4505
R70448 VSS.n2005 VSS.n2004 0.4505
R70449 VSS.n1933 VSS.n1932 0.4505
R70450 VSS.n2000 VSS.n1999 0.4505
R70451 VSS.n1998 VSS.n1935 0.4505
R70452 VSS.n1997 VSS.n1996 0.4505
R70453 VSS.n1937 VSS.n1936 0.4505
R70454 VSS.n1992 VSS.n1991 0.4505
R70455 VSS.n1990 VSS.n1939 0.4505
R70456 VSS.n1989 VSS.n1988 0.4505
R70457 VSS.n1941 VSS.n1940 0.4505
R70458 VSS.n1984 VSS.n1107 0.4505
R70459 VSS.n1983 VSS.n1982 0.4505
R70460 VSS.n1981 VSS.n1943 0.4505
R70461 VSS.n1980 VSS.n1979 0.4505
R70462 VSS.n1945 VSS.n1944 0.4505
R70463 VSS.n1975 VSS.n1974 0.4505
R70464 VSS.n1973 VSS.n1948 0.4505
R70465 VSS.n1972 VSS.n1971 0.4505
R70466 VSS.n1950 VSS.n1949 0.4505
R70467 VSS.n1967 VSS.n1966 0.4505
R70468 VSS.n1965 VSS.n1952 0.4505
R70469 VSS.n1964 VSS.n1963 0.4505
R70470 VSS.n1954 VSS.n1953 0.4505
R70471 VSS.n1959 VSS.n1958 0.4505
R70472 VSS.n1957 VSS.n1956 0.4505
R70473 VSS.n1081 VSS.n1080 0.4505
R70474 VSS.n2988 VSS.n2987 0.4505
R70475 VSS.n1084 VSS.n1078 0.4505
R70476 VSS.n2993 VSS.n2992 0.4505
R70477 VSS.n2994 VSS.n1076 0.4505
R70478 VSS.n2996 VSS.n2995 0.4505
R70479 VSS.n1074 VSS.n1073 0.4505
R70480 VSS.n3001 VSS.n3000 0.4505
R70481 VSS.n3002 VSS.n1072 0.4505
R70482 VSS.n3004 VSS.n3003 0.4505
R70483 VSS.n1070 VSS.n1069 0.4505
R70484 VSS.n3009 VSS.n3008 0.4505
R70485 VSS.n3010 VSS.n1068 0.4505
R70486 VSS.n3012 VSS.n3011 0.4505
R70487 VSS.n1066 VSS.n1065 0.4505
R70488 VSS.n3017 VSS.n3016 0.4505
R70489 VSS.n3018 VSS.n1064 0.4505
R70490 VSS.n3020 VSS.n3019 0.4505
R70491 VSS.n1061 VSS.n1050 0.4505
R70492 VSS.n3063 VSS.n3062 0.4505
R70493 VSS.n1019 VSS.n1018 0.4505
R70494 VSS.n1017 VSS.n1016 0.4505
R70495 VSS.n1024 VSS.n1023 0.4505
R70496 VSS.n1025 VSS.n1015 0.4505
R70497 VSS.n1027 VSS.n1026 0.4505
R70498 VSS.n1013 VSS.n1012 0.4505
R70499 VSS.n1032 VSS.n1031 0.4505
R70500 VSS.n1033 VSS.n1011 0.4505
R70501 VSS.n1035 VSS.n1034 0.4505
R70502 VSS.n1009 VSS.n1008 0.4505
R70503 VSS.n1040 VSS.n1039 0.4505
R70504 VSS.n1041 VSS.n1006 0.4505
R70505 VSS.n1043 VSS.n1042 0.4505
R70506 VSS.n2691 VSS.n1183 0.4505
R70507 VSS.n2693 VSS.n2692 0.4505
R70508 VSS.n1181 VSS.n1180 0.4505
R70509 VSS.n2698 VSS.n2697 0.4505
R70510 VSS.n2699 VSS.n1179 0.4505
R70511 VSS.n2701 VSS.n2700 0.4505
R70512 VSS.n1177 VSS.n1176 0.4505
R70513 VSS.n2706 VSS.n2705 0.4505
R70514 VSS.n2707 VSS.n1175 0.4505
R70515 VSS.n2709 VSS.n2708 0.4505
R70516 VSS.n1173 VSS.n1172 0.4505
R70517 VSS.n2714 VSS.n2713 0.4505
R70518 VSS.n2715 VSS.n1171 0.4505
R70519 VSS.n2717 VSS.n2716 0.4505
R70520 VSS.n1169 VSS.n1168 0.4505
R70521 VSS.n2722 VSS.n2721 0.4505
R70522 VSS.n2723 VSS.n1166 0.4505
R70523 VSS.n2857 VSS.n2856 0.4505
R70524 VSS.n2855 VSS.n1167 0.4505
R70525 VSS.n2854 VSS.n2853 0.4505
R70526 VSS.n2725 VSS.n2724 0.4505
R70527 VSS.n2849 VSS.n2848 0.4505
R70528 VSS.n2847 VSS.n2727 0.4505
R70529 VSS.n2846 VSS.n2845 0.4505
R70530 VSS.n2729 VSS.n2728 0.4505
R70531 VSS.n2841 VSS.n2840 0.4505
R70532 VSS.n2839 VSS.n2731 0.4505
R70533 VSS.n2838 VSS.n2837 0.4505
R70534 VSS.n2733 VSS.n2732 0.4505
R70535 VSS.n2833 VSS.n2832 0.4505
R70536 VSS.n2831 VSS.n2735 0.4505
R70537 VSS.n2830 VSS.n2829 0.4505
R70538 VSS.n2737 VSS.n2736 0.4505
R70539 VSS.n2757 VSS.n2756 0.4505
R70540 VSS.n2758 VSS.n2754 0.4505
R70541 VSS.n2810 VSS.n2809 0.4505
R70542 VSS.n2808 VSS.n2755 0.4505
R70543 VSS.n2807 VSS.n2806 0.4505
R70544 VSS.n2760 VSS.n2759 0.4505
R70545 VSS.n2802 VSS.n2801 0.4505
R70546 VSS.n2800 VSS.n2762 0.4505
R70547 VSS.n2799 VSS.n2798 0.4505
R70548 VSS.n2764 VSS.n2763 0.4505
R70549 VSS.n2794 VSS.n2793 0.4505
R70550 VSS.n2792 VSS.n2766 0.4505
R70551 VSS.n2791 VSS.n2790 0.4505
R70552 VSS.n2768 VSS.n2767 0.4505
R70553 VSS.n2786 VSS.n2785 0.4505
R70554 VSS.n2784 VSS.n2770 0.4505
R70555 VSS.n2783 VSS.n2782 0.4505
R70556 VSS.n2772 VSS.n2771 0.4505
R70557 VSS.n983 VSS.n981 0.4505
R70558 VSS.n3434 VSS.n3433 0.4505
R70559 VSS.n3432 VSS.n982 0.4505
R70560 VSS.n3431 VSS.n3430 0.4505
R70561 VSS.n985 VSS.n984 0.4505
R70562 VSS.n3426 VSS.n3425 0.4505
R70563 VSS.n3424 VSS.n987 0.4505
R70564 VSS.n3423 VSS.n3422 0.4505
R70565 VSS.n989 VSS.n988 0.4505
R70566 VSS.n3418 VSS.n3417 0.4505
R70567 VSS.n3416 VSS.n991 0.4505
R70568 VSS.n3415 VSS.n3414 0.4505
R70569 VSS.n993 VSS.n992 0.4505
R70570 VSS.n3410 VSS.n3409 0.4505
R70571 VSS.n3408 VSS.n995 0.4505
R70572 VSS.n3407 VSS.n3406 0.4505
R70573 VSS.n997 VSS.n996 0.4505
R70574 VSS.n1007 VSS.n1005 0.4505
R70575 VSS.n1021 VSS.n1017 0.4505
R70576 VSS.n1023 VSS.n1022 0.4505
R70577 VSS.n1015 VSS.n1014 0.4505
R70578 VSS.n1028 VSS.n1027 0.4505
R70579 VSS.n1029 VSS.n1013 0.4505
R70580 VSS.n1031 VSS.n1030 0.4505
R70581 VSS.n1011 VSS.n1010 0.4505
R70582 VSS.n1036 VSS.n1035 0.4505
R70583 VSS.n1037 VSS.n1009 0.4505
R70584 VSS.n1039 VSS.n1038 0.4505
R70585 VSS.n1006 VSS.n1004 0.4505
R70586 VSS.n1044 VSS.n1043 0.4505
R70587 VSS.n2689 VSS.n2688 0.4505
R70588 VSS.n1183 VSS.n1182 0.4505
R70589 VSS.n2694 VSS.n2693 0.4505
R70590 VSS.n2695 VSS.n1181 0.4505
R70591 VSS.n2697 VSS.n2696 0.4505
R70592 VSS.n1179 VSS.n1178 0.4505
R70593 VSS.n2702 VSS.n2701 0.4505
R70594 VSS.n2703 VSS.n1177 0.4505
R70595 VSS.n2705 VSS.n2704 0.4505
R70596 VSS.n1175 VSS.n1174 0.4505
R70597 VSS.n2710 VSS.n2709 0.4505
R70598 VSS.n2711 VSS.n1173 0.4505
R70599 VSS.n2713 VSS.n2712 0.4505
R70600 VSS.n1171 VSS.n1170 0.4505
R70601 VSS.n2718 VSS.n2717 0.4505
R70602 VSS.n2719 VSS.n1169 0.4505
R70603 VSS.n2721 VSS.n2720 0.4505
R70604 VSS.n1166 VSS.n1164 0.4505
R70605 VSS.n2858 VSS.n2857 0.4505
R70606 VSS.n1167 VSS.n1165 0.4505
R70607 VSS.n2853 VSS.n2852 0.4505
R70608 VSS.n2851 VSS.n2725 0.4505
R70609 VSS.n2850 VSS.n2849 0.4505
R70610 VSS.n2727 VSS.n2726 0.4505
R70611 VSS.n2845 VSS.n2844 0.4505
R70612 VSS.n2843 VSS.n2729 0.4505
R70613 VSS.n2842 VSS.n2841 0.4505
R70614 VSS.n2731 VSS.n2730 0.4505
R70615 VSS.n2837 VSS.n2836 0.4505
R70616 VSS.n2835 VSS.n2733 0.4505
R70617 VSS.n2834 VSS.n2833 0.4505
R70618 VSS.n2735 VSS.n2734 0.4505
R70619 VSS.n2829 VSS.n2828 0.4505
R70620 VSS.n2827 VSS.n2737 0.4505
R70621 VSS.n2756 VSS.n2743 0.4505
R70622 VSS.n2754 VSS.n2747 0.4505
R70623 VSS.n2811 VSS.n2810 0.4505
R70624 VSS.n2755 VSS.n2753 0.4505
R70625 VSS.n2806 VSS.n2805 0.4505
R70626 VSS.n2804 VSS.n2760 0.4505
R70627 VSS.n2803 VSS.n2802 0.4505
R70628 VSS.n2762 VSS.n2761 0.4505
R70629 VSS.n2798 VSS.n2797 0.4505
R70630 VSS.n2796 VSS.n2764 0.4505
R70631 VSS.n2795 VSS.n2794 0.4505
R70632 VSS.n2766 VSS.n2765 0.4505
R70633 VSS.n2790 VSS.n2789 0.4505
R70634 VSS.n2788 VSS.n2768 0.4505
R70635 VSS.n2787 VSS.n2786 0.4505
R70636 VSS.n2770 VSS.n2769 0.4505
R70637 VSS.n2782 VSS.n2781 0.4505
R70638 VSS.n2780 VSS.n2772 0.4505
R70639 VSS.n981 VSS.n974 0.4505
R70640 VSS.n3435 VSS.n3434 0.4505
R70641 VSS.n982 VSS.n980 0.4505
R70642 VSS.n3430 VSS.n3429 0.4505
R70643 VSS.n3428 VSS.n985 0.4505
R70644 VSS.n3427 VSS.n3426 0.4505
R70645 VSS.n987 VSS.n986 0.4505
R70646 VSS.n3422 VSS.n3421 0.4505
R70647 VSS.n3420 VSS.n989 0.4505
R70648 VSS.n3419 VSS.n3418 0.4505
R70649 VSS.n991 VSS.n990 0.4505
R70650 VSS.n3414 VSS.n3413 0.4505
R70651 VSS.n3412 VSS.n993 0.4505
R70652 VSS.n3411 VSS.n3410 0.4505
R70653 VSS.n995 VSS.n994 0.4505
R70654 VSS.n3406 VSS.n3405 0.4505
R70655 VSS.n3404 VSS.n997 0.4505
R70656 VSS.n1005 VSS.n1003 0.4505
R70657 VSS.n4061 VSS.n4060 0.4505
R70658 VSS.n4063 VSS.n4062 0.4505
R70659 VSS.n4058 VSS.n4057 0.4505
R70660 VSS.n4068 VSS.n4067 0.4505
R70661 VSS.n4069 VSS.n4056 0.4505
R70662 VSS.n4071 VSS.n4070 0.4505
R70663 VSS.n4054 VSS.n4053 0.4505
R70664 VSS.n4076 VSS.n4075 0.4505
R70665 VSS.n4077 VSS.n4052 0.4505
R70666 VSS.n4079 VSS.n4078 0.4505
R70667 VSS.n4049 VSS.n4048 0.4505
R70668 VSS.n4084 VSS.n4083 0.4505
R70669 VSS.n4085 VSS.n587 0.4505
R70670 VSS.n2201 VSS.n2200 0.4505
R70671 VSS.n2199 VSS.n2154 0.4505
R70672 VSS.n2198 VSS.n2197 0.4505
R70673 VSS.n2157 VSS.n2156 0.4505
R70674 VSS.n2193 VSS.n2192 0.4505
R70675 VSS.n2191 VSS.n2159 0.4505
R70676 VSS.n2190 VSS.n2189 0.4505
R70677 VSS.n2161 VSS.n2160 0.4505
R70678 VSS.n2185 VSS.n2184 0.4505
R70679 VSS.n2183 VSS.n2163 0.4505
R70680 VSS.n2182 VSS.n2181 0.4505
R70681 VSS.n2165 VSS.n2164 0.4505
R70682 VSS.n2177 VSS.n2176 0.4505
R70683 VSS.n2175 VSS.n2167 0.4505
R70684 VSS.n2174 VSS.n2173 0.4505
R70685 VSS.n2171 VSS.n2168 0.4505
R70686 VSS.n2170 VSS.n2169 0.4505
R70687 VSS.n653 VSS.n652 0.4505
R70688 VSS.n3941 VSS.n3940 0.4505
R70689 VSS.n3942 VSS.n651 0.4505
R70690 VSS.n3944 VSS.n3943 0.4505
R70691 VSS.n649 VSS.n648 0.4505
R70692 VSS.n3949 VSS.n3948 0.4505
R70693 VSS.n3950 VSS.n647 0.4505
R70694 VSS.n3952 VSS.n3951 0.4505
R70695 VSS.n645 VSS.n644 0.4505
R70696 VSS.n3957 VSS.n3956 0.4505
R70697 VSS.n3958 VSS.n643 0.4505
R70698 VSS.n3960 VSS.n3959 0.4505
R70699 VSS.n641 VSS.n640 0.4505
R70700 VSS.n3965 VSS.n3964 0.4505
R70701 VSS.n3966 VSS.n639 0.4505
R70702 VSS.n3968 VSS.n3967 0.4505
R70703 VSS.n621 VSS.n620 0.4505
R70704 VSS.n3982 VSS.n3981 0.4505
R70705 VSS.n3983 VSS.n619 0.4505
R70706 VSS.n3985 VSS.n3984 0.4505
R70707 VSS.n617 VSS.n616 0.4505
R70708 VSS.n3990 VSS.n3989 0.4505
R70709 VSS.n3991 VSS.n615 0.4505
R70710 VSS.n3993 VSS.n3992 0.4505
R70711 VSS.n613 VSS.n612 0.4505
R70712 VSS.n3998 VSS.n3997 0.4505
R70713 VSS.n3999 VSS.n611 0.4505
R70714 VSS.n4001 VSS.n4000 0.4505
R70715 VSS.n609 VSS.n608 0.4505
R70716 VSS.n4006 VSS.n4005 0.4505
R70717 VSS.n4007 VSS.n607 0.4505
R70718 VSS.n4009 VSS.n4008 0.4505
R70719 VSS.n605 VSS.n604 0.4505
R70720 VSS.n4014 VSS.n4013 0.4505
R70721 VSS.n4015 VSS.n603 0.4505
R70722 VSS.n4017 VSS.n4016 0.4505
R70723 VSS.n601 VSS.n600 0.4505
R70724 VSS.n4022 VSS.n4021 0.4505
R70725 VSS.n4023 VSS.n599 0.4505
R70726 VSS.n4025 VSS.n4024 0.4505
R70727 VSS.n597 VSS.n596 0.4505
R70728 VSS.n4030 VSS.n4029 0.4505
R70729 VSS.n4031 VSS.n595 0.4505
R70730 VSS.n4033 VSS.n4032 0.4505
R70731 VSS.n593 VSS.n592 0.4505
R70732 VSS.n4038 VSS.n4037 0.4505
R70733 VSS.n4039 VSS.n591 0.4505
R70734 VSS.n4041 VSS.n4040 0.4505
R70735 VSS.n589 VSS.n588 0.4505
R70736 VSS.n4046 VSS.n4045 0.4505
R70737 VSS.n4047 VSS.n586 0.4505
R70738 VSS.n4087 VSS.n4086 0.4505
R70739 VSS.n4064 VSS.n4063 0.4505
R70740 VSS.n4065 VSS.n4058 0.4505
R70741 VSS.n4067 VSS.n4066 0.4505
R70742 VSS.n4056 VSS.n4055 0.4505
R70743 VSS.n4072 VSS.n4071 0.4505
R70744 VSS.n4073 VSS.n4054 0.4505
R70745 VSS.n4075 VSS.n4074 0.4505
R70746 VSS.n4052 VSS.n4051 0.4505
R70747 VSS.n4080 VSS.n4079 0.4505
R70748 VSS.n4081 VSS.n4049 0.4505
R70749 VSS.n4083 VSS.n4082 0.4505
R70750 VSS.n4050 VSS.n587 0.4505
R70751 VSS.n2153 VSS.n2151 0.4505
R70752 VSS.n2202 VSS.n2201 0.4505
R70753 VSS.n2154 VSS.n2152 0.4505
R70754 VSS.n2197 VSS.n2196 0.4505
R70755 VSS.n2195 VSS.n2157 0.4505
R70756 VSS.n2194 VSS.n2193 0.4505
R70757 VSS.n2159 VSS.n2158 0.4505
R70758 VSS.n2189 VSS.n2188 0.4505
R70759 VSS.n2187 VSS.n2161 0.4505
R70760 VSS.n2186 VSS.n2185 0.4505
R70761 VSS.n2163 VSS.n2162 0.4505
R70762 VSS.n2181 VSS.n2180 0.4505
R70763 VSS.n2179 VSS.n2165 0.4505
R70764 VSS.n2178 VSS.n2177 0.4505
R70765 VSS.n2167 VSS.n2166 0.4505
R70766 VSS.n2173 VSS.n2172 0.4505
R70767 VSS.n2171 VSS.n660 0.4505
R70768 VSS.n2170 VSS.n654 0.4505
R70769 VSS.n3938 VSS.n653 0.4505
R70770 VSS.n3940 VSS.n3939 0.4505
R70771 VSS.n651 VSS.n650 0.4505
R70772 VSS.n3945 VSS.n3944 0.4505
R70773 VSS.n3946 VSS.n649 0.4505
R70774 VSS.n3948 VSS.n3947 0.4505
R70775 VSS.n647 VSS.n646 0.4505
R70776 VSS.n3953 VSS.n3952 0.4505
R70777 VSS.n3954 VSS.n645 0.4505
R70778 VSS.n3956 VSS.n3955 0.4505
R70779 VSS.n643 VSS.n642 0.4505
R70780 VSS.n3961 VSS.n3960 0.4505
R70781 VSS.n3962 VSS.n641 0.4505
R70782 VSS.n3964 VSS.n3963 0.4505
R70783 VSS.n639 VSS.n638 0.4505
R70784 VSS.n3969 VSS.n3968 0.4505
R70785 VSS.n3975 VSS.n621 0.4505
R70786 VSS.n3981 VSS.n3980 0.4505
R70787 VSS.n619 VSS.n618 0.4505
R70788 VSS.n3986 VSS.n3985 0.4505
R70789 VSS.n3987 VSS.n617 0.4505
R70790 VSS.n3989 VSS.n3988 0.4505
R70791 VSS.n615 VSS.n614 0.4505
R70792 VSS.n3994 VSS.n3993 0.4505
R70793 VSS.n3995 VSS.n613 0.4505
R70794 VSS.n3997 VSS.n3996 0.4505
R70795 VSS.n611 VSS.n610 0.4505
R70796 VSS.n4002 VSS.n4001 0.4505
R70797 VSS.n4003 VSS.n609 0.4505
R70798 VSS.n4005 VSS.n4004 0.4505
R70799 VSS.n607 VSS.n606 0.4505
R70800 VSS.n4010 VSS.n4009 0.4505
R70801 VSS.n4011 VSS.n605 0.4505
R70802 VSS.n4013 VSS.n4012 0.4505
R70803 VSS.n603 VSS.n602 0.4505
R70804 VSS.n4018 VSS.n4017 0.4505
R70805 VSS.n4019 VSS.n601 0.4505
R70806 VSS.n4021 VSS.n4020 0.4505
R70807 VSS.n599 VSS.n598 0.4505
R70808 VSS.n4026 VSS.n4025 0.4505
R70809 VSS.n4027 VSS.n597 0.4505
R70810 VSS.n4029 VSS.n4028 0.4505
R70811 VSS.n595 VSS.n594 0.4505
R70812 VSS.n4034 VSS.n4033 0.4505
R70813 VSS.n4035 VSS.n593 0.4505
R70814 VSS.n4037 VSS.n4036 0.4505
R70815 VSS.n591 VSS.n590 0.4505
R70816 VSS.n4042 VSS.n4041 0.4505
R70817 VSS.n4043 VSS.n589 0.4505
R70818 VSS.n4045 VSS.n4044 0.4505
R70819 VSS.n586 VSS.n575 0.4505
R70820 VSS.n4088 VSS.n4087 0.4505
R70821 VSS.n4699 VSS.n4698 0.4505
R70822 VSS.n4701 VSS.n4700 0.4505
R70823 VSS.n4696 VSS.n4695 0.4505
R70824 VSS.n4706 VSS.n4705 0.4505
R70825 VSS.n4707 VSS.n4694 0.4505
R70826 VSS.n4709 VSS.n4708 0.4505
R70827 VSS.n4692 VSS.n4691 0.4505
R70828 VSS.n4714 VSS.n4713 0.4505
R70829 VSS.n4715 VSS.n4689 0.4505
R70830 VSS.n4717 VSS.n4716 0.4505
R70831 VSS.n4690 VSS.n4687 0.4505
R70832 VSS.n4721 VSS.n4686 0.4505
R70833 VSS.n4723 VSS.n4722 0.4505
R70834 VSS.n4572 VSS.n4569 0.4505
R70835 VSS.n4574 VSS.n4573 0.4505
R70836 VSS.n4568 VSS.n4567 0.4505
R70837 VSS.n4579 VSS.n4578 0.4505
R70838 VSS.n4580 VSS.n4566 0.4505
R70839 VSS.n4582 VSS.n4581 0.4505
R70840 VSS.n4564 VSS.n4563 0.4505
R70841 VSS.n4587 VSS.n4586 0.4505
R70842 VSS.n4588 VSS.n4562 0.4505
R70843 VSS.n4590 VSS.n4589 0.4505
R70844 VSS.n4560 VSS.n4559 0.4505
R70845 VSS.n4595 VSS.n4594 0.4505
R70846 VSS.n4596 VSS.n4558 0.4505
R70847 VSS.n4599 VSS.n4598 0.4505
R70848 VSS.n4597 VSS.n4556 0.4505
R70849 VSS.n4603 VSS.n4555 0.4505
R70850 VSS.n4605 VSS.n4604 0.4505
R70851 VSS.n4606 VSS.n4554 0.4505
R70852 VSS.n4608 VSS.n4607 0.4505
R70853 VSS.n4553 VSS.n4552 0.4505
R70854 VSS.n4613 VSS.n4612 0.4505
R70855 VSS.n4614 VSS.n4551 0.4505
R70856 VSS.n4616 VSS.n4615 0.4505
R70857 VSS.n4549 VSS.n4548 0.4505
R70858 VSS.n4621 VSS.n4620 0.4505
R70859 VSS.n4622 VSS.n4547 0.4505
R70860 VSS.n4624 VSS.n4623 0.4505
R70861 VSS.n4545 VSS.n4544 0.4505
R70862 VSS.n4629 VSS.n4628 0.4505
R70863 VSS.n4630 VSS.n4543 0.4505
R70864 VSS.n4632 VSS.n4631 0.4505
R70865 VSS.n4541 VSS.n4540 0.4505
R70866 VSS.n4637 VSS.n4636 0.4505
R70867 VSS.n4638 VSS.n4539 0.4505
R70868 VSS.n4640 VSS.n4639 0.4505
R70869 VSS.n4641 VSS.n4537 0.4505
R70870 VSS.n4644 VSS.n4643 0.4505
R70871 VSS.n4645 VSS.n4536 0.4505
R70872 VSS.n4647 VSS.n4646 0.4505
R70873 VSS.n4534 VSS.n4533 0.4505
R70874 VSS.n4652 VSS.n4651 0.4505
R70875 VSS.n4653 VSS.n4532 0.4505
R70876 VSS.n4655 VSS.n4654 0.4505
R70877 VSS.n4530 VSS.n4529 0.4505
R70878 VSS.n4660 VSS.n4659 0.4505
R70879 VSS.n4661 VSS.n4528 0.4505
R70880 VSS.n4663 VSS.n4662 0.4505
R70881 VSS.n4526 VSS.n4525 0.4505
R70882 VSS.n4668 VSS.n4667 0.4505
R70883 VSS.n4669 VSS.n4523 0.4505
R70884 VSS.n4759 VSS.n4758 0.4505
R70885 VSS.n4757 VSS.n4524 0.4505
R70886 VSS.n4756 VSS.n4755 0.4505
R70887 VSS.n4754 VSS.n4670 0.4505
R70888 VSS.n4674 VSS.n4671 0.4505
R70889 VSS.n4750 VSS.n4749 0.4505
R70890 VSS.n4748 VSS.n4673 0.4505
R70891 VSS.n4747 VSS.n4746 0.4505
R70892 VSS.n4676 VSS.n4675 0.4505
R70893 VSS.n4742 VSS.n4741 0.4505
R70894 VSS.n4740 VSS.n4678 0.4505
R70895 VSS.n4739 VSS.n4738 0.4505
R70896 VSS.n4680 VSS.n4679 0.4505
R70897 VSS.n4734 VSS.n4733 0.4505
R70898 VSS.n4732 VSS.n4682 0.4505
R70899 VSS.n4731 VSS.n4730 0.4505
R70900 VSS.n4684 VSS.n4683 0.4505
R70901 VSS.n4726 VSS.n4725 0.4505
R70902 VSS.n4724 VSS.n4685 0.4505
R70903 VSS.n4702 VSS.n4701 0.4505
R70904 VSS.n4703 VSS.n4696 0.4505
R70905 VSS.n4705 VSS.n4704 0.4505
R70906 VSS.n4694 VSS.n4693 0.4505
R70907 VSS.n4710 VSS.n4709 0.4505
R70908 VSS.n4711 VSS.n4692 0.4505
R70909 VSS.n4713 VSS.n4712 0.4505
R70910 VSS.n4689 VSS.n4688 0.4505
R70911 VSS.n4718 VSS.n4717 0.4505
R70912 VSS.n4719 VSS.n4687 0.4505
R70913 VSS.n4721 VSS.n4720 0.4505
R70914 VSS.n4722 VSS.n498 0.4505
R70915 VSS.n4570 VSS.n4251 0.4505
R70916 VSS.n4569 VSS.n4255 0.4505
R70917 VSS.n4575 VSS.n4574 0.4505
R70918 VSS.n4576 VSS.n4568 0.4505
R70919 VSS.n4578 VSS.n4577 0.4505
R70920 VSS.n4566 VSS.n4565 0.4505
R70921 VSS.n4583 VSS.n4582 0.4505
R70922 VSS.n4584 VSS.n4564 0.4505
R70923 VSS.n4586 VSS.n4585 0.4505
R70924 VSS.n4562 VSS.n4561 0.4505
R70925 VSS.n4591 VSS.n4590 0.4505
R70926 VSS.n4592 VSS.n4560 0.4505
R70927 VSS.n4594 VSS.n4593 0.4505
R70928 VSS.n4558 VSS.n4557 0.4505
R70929 VSS.n4600 VSS.n4599 0.4505
R70930 VSS.n4601 VSS.n4556 0.4505
R70931 VSS.n4603 VSS.n4602 0.4505
R70932 VSS.n4604 VSS.n4270 0.4505
R70933 VSS.n4554 VSS.n4273 0.4505
R70934 VSS.n4609 VSS.n4608 0.4505
R70935 VSS.n4610 VSS.n4553 0.4505
R70936 VSS.n4612 VSS.n4611 0.4505
R70937 VSS.n4551 VSS.n4550 0.4505
R70938 VSS.n4617 VSS.n4616 0.4505
R70939 VSS.n4618 VSS.n4549 0.4505
R70940 VSS.n4620 VSS.n4619 0.4505
R70941 VSS.n4547 VSS.n4546 0.4505
R70942 VSS.n4625 VSS.n4624 0.4505
R70943 VSS.n4626 VSS.n4545 0.4505
R70944 VSS.n4628 VSS.n4627 0.4505
R70945 VSS.n4543 VSS.n4542 0.4505
R70946 VSS.n4633 VSS.n4632 0.4505
R70947 VSS.n4634 VSS.n4541 0.4505
R70948 VSS.n4636 VSS.n4635 0.4505
R70949 VSS.n4539 VSS.n4538 0.4505
R70950 VSS.n4640 VSS.n4490 0.4505
R70951 VSS.n4641 VSS.n4496 0.4505
R70952 VSS.n4643 VSS.n4642 0.4505
R70953 VSS.n4536 VSS.n4535 0.4505
R70954 VSS.n4648 VSS.n4647 0.4505
R70955 VSS.n4649 VSS.n4534 0.4505
R70956 VSS.n4651 VSS.n4650 0.4505
R70957 VSS.n4532 VSS.n4531 0.4505
R70958 VSS.n4656 VSS.n4655 0.4505
R70959 VSS.n4657 VSS.n4530 0.4505
R70960 VSS.n4659 VSS.n4658 0.4505
R70961 VSS.n4528 VSS.n4527 0.4505
R70962 VSS.n4664 VSS.n4663 0.4505
R70963 VSS.n4665 VSS.n4526 0.4505
R70964 VSS.n4667 VSS.n4666 0.4505
R70965 VSS.n4523 VSS.n4522 0.4505
R70966 VSS.n4760 VSS.n4759 0.4505
R70967 VSS.n4524 VSS.n4516 0.4505
R70968 VSS.n4755 VSS.n4518 0.4505
R70969 VSS.n4754 VSS.n4753 0.4505
R70970 VSS.n4752 VSS.n4671 0.4505
R70971 VSS.n4751 VSS.n4750 0.4505
R70972 VSS.n4673 VSS.n4672 0.4505
R70973 VSS.n4746 VSS.n4745 0.4505
R70974 VSS.n4744 VSS.n4676 0.4505
R70975 VSS.n4743 VSS.n4742 0.4505
R70976 VSS.n4678 VSS.n4677 0.4505
R70977 VSS.n4738 VSS.n4737 0.4505
R70978 VSS.n4736 VSS.n4680 0.4505
R70979 VSS.n4735 VSS.n4734 0.4505
R70980 VSS.n4682 VSS.n4681 0.4505
R70981 VSS.n4730 VSS.n4729 0.4505
R70982 VSS.n4728 VSS.n4684 0.4505
R70983 VSS.n4727 VSS.n4726 0.4505
R70984 VSS.n4685 VSS.n491 0.4505
R70985 VSS.n2745 VSS.n970 0.4505
R70986 VSS.n923 VSS.n922 0.4505
R70987 VSS.n6243 VSS.n122 0.4505
R70988 VSS.n6245 VSS.n6244 0.4505
R70989 VSS.n6246 VSS.n120 0.4505
R70990 VSS.n6250 VSS.n6249 0.4505
R70991 VSS.n6251 VSS.n119 0.4505
R70992 VSS.n6253 VSS.n6252 0.4505
R70993 VSS.n117 VSS.n116 0.4505
R70994 VSS.n6258 VSS.n6257 0.4505
R70995 VSS.n6259 VSS.n115 0.4505
R70996 VSS.n6261 VSS.n6260 0.4505
R70997 VSS.n113 VSS.n112 0.4505
R70998 VSS.n6266 VSS.n6265 0.4505
R70999 VSS.n6267 VSS.n111 0.4505
R71000 VSS.n6443 VSS.n6442 0.4505
R71001 VSS.n24 VSS.n23 0.4505
R71002 VSS.n6438 VSS.n6437 0.4505
R71003 VSS.n6436 VSS.n26 0.4505
R71004 VSS.n6435 VSS.n6434 0.4505
R71005 VSS.n28 VSS.n27 0.4505
R71006 VSS.n6430 VSS.n6429 0.4505
R71007 VSS.n6428 VSS.n30 0.4505
R71008 VSS.n6427 VSS.n6426 0.4505
R71009 VSS.n32 VSS.n31 0.4505
R71010 VSS.n6422 VSS.n6421 0.4505
R71011 VSS.n6420 VSS.n34 0.4505
R71012 VSS.n6419 VSS.n6418 0.4505
R71013 VSS.n36 VSS.n35 0.4505
R71014 VSS.n6414 VSS.n6413 0.4505
R71015 VSS.n6412 VSS.n38 0.4505
R71016 VSS.n6411 VSS.n6410 0.4505
R71017 VSS.n40 VSS.n39 0.4505
R71018 VSS.n6406 VSS.n6405 0.4505
R71019 VSS.n6404 VSS.n42 0.4505
R71020 VSS.n6403 VSS.n6402 0.4505
R71021 VSS.n44 VSS.n43 0.4505
R71022 VSS.n6398 VSS.n6397 0.4505
R71023 VSS.n6396 VSS.n46 0.4505
R71024 VSS.n6395 VSS.n6394 0.4505
R71025 VSS.n48 VSS.n47 0.4505
R71026 VSS.n6390 VSS.n6389 0.4505
R71027 VSS.n6388 VSS.n50 0.4505
R71028 VSS.n6387 VSS.n6386 0.4505
R71029 VSS.n52 VSS.n51 0.4505
R71030 VSS.n6382 VSS.n6381 0.4505
R71031 VSS.n6380 VSS.n54 0.4505
R71032 VSS.n6379 VSS.n6378 0.4505
R71033 VSS.n56 VSS.n55 0.4505
R71034 VSS.n6374 VSS.n6373 0.4505
R71035 VSS.n6372 VSS.n58 0.4505
R71036 VSS.n6371 VSS.n6370 0.4505
R71037 VSS.n60 VSS.n59 0.4505
R71038 VSS.n6366 VSS.n6365 0.4505
R71039 VSS.n6364 VSS.n62 0.4505
R71040 VSS.n6363 VSS.n6362 0.4505
R71041 VSS.n64 VSS.n63 0.4505
R71042 VSS.n6358 VSS.n6357 0.4505
R71043 VSS.n6356 VSS.n66 0.4505
R71044 VSS.n6355 VSS.n6354 0.4505
R71045 VSS.n68 VSS.n67 0.4505
R71046 VSS.n6350 VSS.n6349 0.4505
R71047 VSS.n6348 VSS.n70 0.4505
R71048 VSS.n6347 VSS.n6346 0.4505
R71049 VSS.n72 VSS.n71 0.4505
R71050 VSS.n6342 VSS.n6341 0.4505
R71051 VSS.n6340 VSS.n74 0.4505
R71052 VSS.n6339 VSS.n6338 0.4505
R71053 VSS.n76 VSS.n75 0.4505
R71054 VSS.n6334 VSS.n6333 0.4505
R71055 VSS.n6332 VSS.n78 0.4505
R71056 VSS.n6331 VSS.n6330 0.4505
R71057 VSS.n80 VSS.n79 0.4505
R71058 VSS.n6326 VSS.n6325 0.4505
R71059 VSS.n6324 VSS.n82 0.4505
R71060 VSS.n6323 VSS.n6322 0.4505
R71061 VSS.n84 VSS.n83 0.4505
R71062 VSS.n6318 VSS.n6317 0.4505
R71063 VSS.n6316 VSS.n86 0.4505
R71064 VSS.n6315 VSS.n6314 0.4505
R71065 VSS.n88 VSS.n87 0.4505
R71066 VSS.n6310 VSS.n6309 0.4505
R71067 VSS.n6308 VSS.n90 0.4505
R71068 VSS.n6307 VSS.n6306 0.4505
R71069 VSS.n92 VSS.n91 0.4505
R71070 VSS.n6302 VSS.n6301 0.4505
R71071 VSS.n6300 VSS.n94 0.4505
R71072 VSS.n6299 VSS.n6298 0.4505
R71073 VSS.n96 VSS.n95 0.4505
R71074 VSS.n6294 VSS.n6293 0.4505
R71075 VSS.n6292 VSS.n98 0.4505
R71076 VSS.n6291 VSS.n6290 0.4505
R71077 VSS.n100 VSS.n99 0.4505
R71078 VSS.n6286 VSS.n6285 0.4505
R71079 VSS.n6284 VSS.n102 0.4505
R71080 VSS.n6283 VSS.n6282 0.4505
R71081 VSS.n104 VSS.n103 0.4505
R71082 VSS.n6278 VSS.n6277 0.4505
R71083 VSS.n6276 VSS.n106 0.4505
R71084 VSS.n6275 VSS.n6274 0.4505
R71085 VSS.n108 VSS.n107 0.4505
R71086 VSS.n6269 VSS.n6268 0.4505
R71087 VSS.n111 VSS.n110 0.4505
R71088 VSS.n6265 VSS.n6264 0.4505
R71089 VSS.n6263 VSS.n113 0.4505
R71090 VSS.n6262 VSS.n6261 0.4505
R71091 VSS.n115 VSS.n114 0.4505
R71092 VSS.n6257 VSS.n6256 0.4505
R71093 VSS.n6255 VSS.n117 0.4505
R71094 VSS.n6254 VSS.n6253 0.4505
R71095 VSS.n119 VSS.n118 0.4505
R71096 VSS.n6249 VSS.n6248 0.4505
R71097 VSS.n6247 VSS.n6246 0.4505
R71098 VSS.n6245 VSS.n121 0.4505
R71099 VSS.n6239 VSS.n122 0.4505
R71100 VSS.n6241 VSS.n6240 0.4505
R71101 VSS.n22 VSS.n21 0.4505
R71102 VSS.n6442 VSS.n6441 0.4505
R71103 VSS.n6440 VSS.n24 0.4505
R71104 VSS.n6439 VSS.n6438 0.4505
R71105 VSS.n26 VSS.n25 0.4505
R71106 VSS.n6434 VSS.n6433 0.4505
R71107 VSS.n6432 VSS.n28 0.4505
R71108 VSS.n6431 VSS.n6430 0.4505
R71109 VSS.n30 VSS.n29 0.4505
R71110 VSS.n6426 VSS.n6425 0.4505
R71111 VSS.n6424 VSS.n32 0.4505
R71112 VSS.n6423 VSS.n6422 0.4505
R71113 VSS.n34 VSS.n33 0.4505
R71114 VSS.n6418 VSS.n6417 0.4505
R71115 VSS.n6416 VSS.n36 0.4505
R71116 VSS.n6415 VSS.n6414 0.4505
R71117 VSS.n38 VSS.n37 0.4505
R71118 VSS.n6410 VSS.n6409 0.4505
R71119 VSS.n6408 VSS.n40 0.4505
R71120 VSS.n6407 VSS.n6406 0.4505
R71121 VSS.n42 VSS.n41 0.4505
R71122 VSS.n6402 VSS.n6401 0.4505
R71123 VSS.n6400 VSS.n44 0.4505
R71124 VSS.n6399 VSS.n6398 0.4505
R71125 VSS.n46 VSS.n45 0.4505
R71126 VSS.n6394 VSS.n6393 0.4505
R71127 VSS.n6392 VSS.n48 0.4505
R71128 VSS.n6391 VSS.n6390 0.4505
R71129 VSS.n50 VSS.n49 0.4505
R71130 VSS.n6386 VSS.n6385 0.4505
R71131 VSS.n6384 VSS.n52 0.4505
R71132 VSS.n6383 VSS.n6382 0.4505
R71133 VSS.n54 VSS.n53 0.4505
R71134 VSS.n6378 VSS.n6377 0.4505
R71135 VSS.n6376 VSS.n56 0.4505
R71136 VSS.n6375 VSS.n6374 0.4505
R71137 VSS.n58 VSS.n57 0.4505
R71138 VSS.n6370 VSS.n6369 0.4505
R71139 VSS.n6368 VSS.n60 0.4505
R71140 VSS.n6367 VSS.n6366 0.4505
R71141 VSS.n62 VSS.n61 0.4505
R71142 VSS.n6362 VSS.n6361 0.4505
R71143 VSS.n6360 VSS.n64 0.4505
R71144 VSS.n6359 VSS.n6358 0.4505
R71145 VSS.n66 VSS.n65 0.4505
R71146 VSS.n6354 VSS.n6353 0.4505
R71147 VSS.n6352 VSS.n68 0.4505
R71148 VSS.n6351 VSS.n6350 0.4505
R71149 VSS.n70 VSS.n69 0.4505
R71150 VSS.n6346 VSS.n6345 0.4505
R71151 VSS.n6344 VSS.n72 0.4505
R71152 VSS.n6343 VSS.n6342 0.4505
R71153 VSS.n74 VSS.n73 0.4505
R71154 VSS.n6338 VSS.n6337 0.4505
R71155 VSS.n6336 VSS.n76 0.4505
R71156 VSS.n6335 VSS.n6334 0.4505
R71157 VSS.n78 VSS.n77 0.4505
R71158 VSS.n6330 VSS.n6329 0.4505
R71159 VSS.n6328 VSS.n80 0.4505
R71160 VSS.n6327 VSS.n6326 0.4505
R71161 VSS.n82 VSS.n81 0.4505
R71162 VSS.n6322 VSS.n6321 0.4505
R71163 VSS.n6320 VSS.n84 0.4505
R71164 VSS.n6319 VSS.n6318 0.4505
R71165 VSS.n86 VSS.n85 0.4505
R71166 VSS.n6314 VSS.n6313 0.4505
R71167 VSS.n6312 VSS.n88 0.4505
R71168 VSS.n6311 VSS.n6310 0.4505
R71169 VSS.n90 VSS.n89 0.4505
R71170 VSS.n6306 VSS.n6305 0.4505
R71171 VSS.n6304 VSS.n92 0.4505
R71172 VSS.n6303 VSS.n6302 0.4505
R71173 VSS.n94 VSS.n93 0.4505
R71174 VSS.n6298 VSS.n6297 0.4505
R71175 VSS.n6296 VSS.n96 0.4505
R71176 VSS.n6295 VSS.n6294 0.4505
R71177 VSS.n98 VSS.n97 0.4505
R71178 VSS.n6290 VSS.n6289 0.4505
R71179 VSS.n6288 VSS.n100 0.4505
R71180 VSS.n6287 VSS.n6286 0.4505
R71181 VSS.n102 VSS.n101 0.4505
R71182 VSS.n6282 VSS.n6281 0.4505
R71183 VSS.n6280 VSS.n104 0.4505
R71184 VSS.n6279 VSS.n6278 0.4505
R71185 VSS.n106 VSS.n105 0.4505
R71186 VSS.n6274 VSS.n6273 0.4505
R71187 VSS.n6272 VSS.n108 0.4505
R71188 VSS.n6270 VSS.n6269 0.4505
R71189 VSS.n260 VSS.n232 0.4505
R71190 VSS.n259 VSS.n258 0.4505
R71191 VSS.n234 VSS.n233 0.4505
R71192 VSS.n254 VSS.n253 0.4505
R71193 VSS.n252 VSS.n237 0.4505
R71194 VSS.n251 VSS.n250 0.4505
R71195 VSS.n239 VSS.n238 0.4505
R71196 VSS.n246 VSS.n245 0.4505
R71197 VSS.n244 VSS.n243 0.4505
R71198 VSS.n242 VSS.n0 0.4505
R71199 VSS.n6469 VSS.n6468 0.4505
R71200 VSS.n2 VSS.n1 0.4505
R71201 VSS.n6464 VSS.n6463 0.4505
R71202 VSS.n6462 VSS.n4 0.4505
R71203 VSS.n435 VSS.n144 0.4505
R71204 VSS.n434 VSS.n433 0.4505
R71205 VSS.n432 VSS.n146 0.4505
R71206 VSS.n431 VSS.n430 0.4505
R71207 VSS.n148 VSS.n147 0.4505
R71208 VSS.n426 VSS.n425 0.4505
R71209 VSS.n424 VSS.n151 0.4505
R71210 VSS.n423 VSS.n422 0.4505
R71211 VSS.n153 VSS.n152 0.4505
R71212 VSS.n418 VSS.n417 0.4505
R71213 VSS.n416 VSS.n155 0.4505
R71214 VSS.n415 VSS.n414 0.4505
R71215 VSS.n157 VSS.n156 0.4505
R71216 VSS.n410 VSS.n409 0.4505
R71217 VSS.n408 VSS.n159 0.4505
R71218 VSS.n407 VSS.n406 0.4505
R71219 VSS.n161 VSS.n160 0.4505
R71220 VSS.n402 VSS.n401 0.4505
R71221 VSS.n400 VSS.n163 0.4505
R71222 VSS.n399 VSS.n398 0.4505
R71223 VSS.n165 VSS.n164 0.4505
R71224 VSS.n394 VSS.n393 0.4505
R71225 VSS.n392 VSS.n167 0.4505
R71226 VSS.n391 VSS.n390 0.4505
R71227 VSS.n169 VSS.n168 0.4505
R71228 VSS.n386 VSS.n385 0.4505
R71229 VSS.n384 VSS.n171 0.4505
R71230 VSS.n383 VSS.n382 0.4505
R71231 VSS.n173 VSS.n172 0.4505
R71232 VSS.n378 VSS.n377 0.4505
R71233 VSS.n376 VSS.n175 0.4505
R71234 VSS.n375 VSS.n374 0.4505
R71235 VSS.n177 VSS.n176 0.4505
R71236 VSS.n370 VSS.n369 0.4505
R71237 VSS.n368 VSS.n179 0.4505
R71238 VSS.n367 VSS.n366 0.4505
R71239 VSS.n181 VSS.n180 0.4505
R71240 VSS.n362 VSS.n361 0.4505
R71241 VSS.n360 VSS.n183 0.4505
R71242 VSS.n359 VSS.n358 0.4505
R71243 VSS.n185 VSS.n184 0.4505
R71244 VSS.n354 VSS.n353 0.4505
R71245 VSS.n352 VSS.n187 0.4505
R71246 VSS.n351 VSS.n350 0.4505
R71247 VSS.n189 VSS.n188 0.4505
R71248 VSS.n346 VSS.n345 0.4505
R71249 VSS.n344 VSS.n191 0.4505
R71250 VSS.n343 VSS.n342 0.4505
R71251 VSS.n193 VSS.n192 0.4505
R71252 VSS.n338 VSS.n337 0.4505
R71253 VSS.n336 VSS.n195 0.4505
R71254 VSS.n335 VSS.n334 0.4505
R71255 VSS.n197 VSS.n196 0.4505
R71256 VSS.n330 VSS.n329 0.4505
R71257 VSS.n328 VSS.n199 0.4505
R71258 VSS.n327 VSS.n326 0.4505
R71259 VSS.n201 VSS.n200 0.4505
R71260 VSS.n322 VSS.n321 0.4505
R71261 VSS.n320 VSS.n203 0.4505
R71262 VSS.n319 VSS.n318 0.4505
R71263 VSS.n205 VSS.n204 0.4505
R71264 VSS.n314 VSS.n313 0.4505
R71265 VSS.n312 VSS.n207 0.4505
R71266 VSS.n311 VSS.n310 0.4505
R71267 VSS.n209 VSS.n208 0.4505
R71268 VSS.n306 VSS.n305 0.4505
R71269 VSS.n304 VSS.n211 0.4505
R71270 VSS.n303 VSS.n302 0.4505
R71271 VSS.n213 VSS.n212 0.4505
R71272 VSS.n298 VSS.n297 0.4505
R71273 VSS.n296 VSS.n215 0.4505
R71274 VSS.n295 VSS.n294 0.4505
R71275 VSS.n217 VSS.n216 0.4505
R71276 VSS.n290 VSS.n289 0.4505
R71277 VSS.n288 VSS.n219 0.4505
R71278 VSS.n287 VSS.n286 0.4505
R71279 VSS.n221 VSS.n220 0.4505
R71280 VSS.n282 VSS.n281 0.4505
R71281 VSS.n280 VSS.n223 0.4505
R71282 VSS.n279 VSS.n278 0.4505
R71283 VSS.n225 VSS.n224 0.4505
R71284 VSS.n274 VSS.n273 0.4505
R71285 VSS.n272 VSS.n227 0.4505
R71286 VSS.n271 VSS.n270 0.4505
R71287 VSS.n229 VSS.n228 0.4505
R71288 VSS.n266 VSS.n265 0.4505
R71289 VSS.n264 VSS.n263 0.4505
R71290 VSS.n235 VSS.n232 0.4505
R71291 VSS.n258 VSS.n257 0.4505
R71292 VSS.n256 VSS.n234 0.4505
R71293 VSS.n255 VSS.n254 0.4505
R71294 VSS.n237 VSS.n236 0.4505
R71295 VSS.n250 VSS.n249 0.4505
R71296 VSS.n248 VSS.n239 0.4505
R71297 VSS.n247 VSS.n246 0.4505
R71298 VSS.n243 VSS.n240 0.4505
R71299 VSS.n242 VSS.n241 0.4505
R71300 VSS.n6468 VSS.n6467 0.4505
R71301 VSS.n6466 VSS.n2 0.4505
R71302 VSS.n6465 VSS.n6464 0.4505
R71303 VSS.n434 VSS.n145 0.4505
R71304 VSS.n149 VSS.n146 0.4505
R71305 VSS.n430 VSS.n429 0.4505
R71306 VSS.n428 VSS.n148 0.4505
R71307 VSS.n427 VSS.n426 0.4505
R71308 VSS.n151 VSS.n150 0.4505
R71309 VSS.n422 VSS.n421 0.4505
R71310 VSS.n420 VSS.n153 0.4505
R71311 VSS.n419 VSS.n418 0.4505
R71312 VSS.n155 VSS.n154 0.4505
R71313 VSS.n414 VSS.n413 0.4505
R71314 VSS.n412 VSS.n157 0.4505
R71315 VSS.n411 VSS.n410 0.4505
R71316 VSS.n159 VSS.n158 0.4505
R71317 VSS.n406 VSS.n405 0.4505
R71318 VSS.n404 VSS.n161 0.4505
R71319 VSS.n403 VSS.n402 0.4505
R71320 VSS.n163 VSS.n162 0.4505
R71321 VSS.n398 VSS.n397 0.4505
R71322 VSS.n396 VSS.n165 0.4505
R71323 VSS.n395 VSS.n394 0.4505
R71324 VSS.n167 VSS.n166 0.4505
R71325 VSS.n390 VSS.n389 0.4505
R71326 VSS.n388 VSS.n169 0.4505
R71327 VSS.n387 VSS.n386 0.4505
R71328 VSS.n171 VSS.n170 0.4505
R71329 VSS.n382 VSS.n381 0.4505
R71330 VSS.n380 VSS.n173 0.4505
R71331 VSS.n379 VSS.n378 0.4505
R71332 VSS.n175 VSS.n174 0.4505
R71333 VSS.n374 VSS.n373 0.4505
R71334 VSS.n372 VSS.n177 0.4505
R71335 VSS.n371 VSS.n370 0.4505
R71336 VSS.n179 VSS.n178 0.4505
R71337 VSS.n366 VSS.n365 0.4505
R71338 VSS.n364 VSS.n181 0.4505
R71339 VSS.n363 VSS.n362 0.4505
R71340 VSS.n183 VSS.n182 0.4505
R71341 VSS.n358 VSS.n357 0.4505
R71342 VSS.n356 VSS.n185 0.4505
R71343 VSS.n355 VSS.n354 0.4505
R71344 VSS.n187 VSS.n186 0.4505
R71345 VSS.n350 VSS.n349 0.4505
R71346 VSS.n348 VSS.n189 0.4505
R71347 VSS.n347 VSS.n346 0.4505
R71348 VSS.n191 VSS.n190 0.4505
R71349 VSS.n342 VSS.n341 0.4505
R71350 VSS.n340 VSS.n193 0.4505
R71351 VSS.n339 VSS.n338 0.4505
R71352 VSS.n195 VSS.n194 0.4505
R71353 VSS.n334 VSS.n333 0.4505
R71354 VSS.n332 VSS.n197 0.4505
R71355 VSS.n331 VSS.n330 0.4505
R71356 VSS.n199 VSS.n198 0.4505
R71357 VSS.n326 VSS.n325 0.4505
R71358 VSS.n324 VSS.n201 0.4505
R71359 VSS.n323 VSS.n322 0.4505
R71360 VSS.n203 VSS.n202 0.4505
R71361 VSS.n318 VSS.n317 0.4505
R71362 VSS.n316 VSS.n205 0.4505
R71363 VSS.n315 VSS.n314 0.4505
R71364 VSS.n207 VSS.n206 0.4505
R71365 VSS.n310 VSS.n309 0.4505
R71366 VSS.n308 VSS.n209 0.4505
R71367 VSS.n307 VSS.n306 0.4505
R71368 VSS.n211 VSS.n210 0.4505
R71369 VSS.n302 VSS.n301 0.4505
R71370 VSS.n300 VSS.n213 0.4505
R71371 VSS.n299 VSS.n298 0.4505
R71372 VSS.n215 VSS.n214 0.4505
R71373 VSS.n294 VSS.n293 0.4505
R71374 VSS.n292 VSS.n217 0.4505
R71375 VSS.n291 VSS.n290 0.4505
R71376 VSS.n219 VSS.n218 0.4505
R71377 VSS.n286 VSS.n285 0.4505
R71378 VSS.n284 VSS.n221 0.4505
R71379 VSS.n283 VSS.n282 0.4505
R71380 VSS.n223 VSS.n222 0.4505
R71381 VSS.n278 VSS.n277 0.4505
R71382 VSS.n276 VSS.n225 0.4505
R71383 VSS.n275 VSS.n274 0.4505
R71384 VSS.n227 VSS.n226 0.4505
R71385 VSS.n270 VSS.n269 0.4505
R71386 VSS.n268 VSS.n229 0.4505
R71387 VSS.n267 VSS.n266 0.4505
R71388 VSS.n263 VSS.n230 0.4505
R71389 VSS.n262 VSS.n231 0.4505
R71390 VSS.n262 VSS.n261 0.4505
R71391 VSS.n1891 DVSS 0.435162
R71392 DVSS VSS.n1893 0.435162
R71393 VSS.n6193 VSS.n6192 0.423402
R71394 VSS.n2907 VSS.n1153 0.400952
R71395 VSS.n2955 VSS.n2954 0.400952
R71396 VSS.n2874 VSS.n1155 0.400952
R71397 VSS.n2962 VSS.n2961 0.400952
R71398 VSS.n2909 VSS.n1150 0.400952
R71399 VSS.n1137 VSS.n1133 0.400952
R71400 VSS.n1278 VSS.n1138 0.40055
R71401 VSS.n1533 VSS.n1147 0.40055
R71402 VSS.n4126 VSS.n4125 0.400345
R71403 VSS.n6196 VSS.n6195 0.371929
R71404 VSS.n562 VSS.n450 0.371929
R71405 VSS.n1887 DVSS 0.367475
R71406 VSS.n1897 DVSS 0.367475
R71407 VSS.n923 VSS.n569 0.355295
R71408 VSS.n6238 VSS.n6237 0.355011
R71409 VSS.n6461 VSS.n6460 0.355011
R71410 VSS.n6446 VSS.n6445 0.354754
R71411 VSS.n438 VSS.n437 0.354754
R71412 VSS.n1887 VSS.n1886 0.352976
R71413 VSS.n1900 VSS.n1897 0.352976
R71414 VSS.n2825 VSS.n2745 0.349418
R71415 VSS.n1219 DVSS 0.34295
R71416 VSS.n4139 VSS.n552 0.3326
R71417 VSS.n4093 VSS.n551 0.3326
R71418 VSS.n6187 VSS.n6186 0.3326
R71419 VSS.n6161 VSS.n6160 0.3326
R71420 VSS.n1434 VSS.n1311 0.329772
R71421 VSS.n2823 VSS.n2816 0.329604
R71422 VSS.n3265 VSS.n864 0.321929
R71423 VSS.n894 VSS.n793 0.321929
R71424 VSS.n3508 VSS.n674 0.321929
R71425 VSS.n2552 VSS.n2068 0.321929
R71426 VSS.n4195 VSS.n4194 0.3092
R71427 VSS.n4198 VSS.n4197 0.3092
R71428 VSS.n2950 VSS.n2949 0.3092
R71429 VSS.n2951 VSS.n1120 0.3092
R71430 VSS.n4186 VSS.n540 0.3092
R71431 VSS.n4204 VSS.n535 0.3092
R71432 VSS.n2933 VSS.n2932 0.3092
R71433 VSS.n2929 VSS.n2928 0.3092
R71434 VSS.n6177 VSS.n6176 0.3092
R71435 VSS.n528 VSS.n469 0.3092
R71436 VSS.n6172 VSS.n6170 0.3092
R71437 VSS.n4199 VSS.n472 0.3092
R71438 VSS.n2946 VSS.n2945 0.30245
R71439 VSS.n2937 VSS.n2936 0.30245
R71440 VSS.n6155 VSS.n471 0.273435
R71441 VSS.n4196 VSS.n538 0.273435
R71442 VSS.n6154 VSS.n474 0.273435
R71443 VSS.n6141 VSS.n477 0.273435
R71444 VSS.n5490 VSS.n475 0.273435
R71445 VSS.n5862 VSS.n5861 0.273435
R71446 VSS.n6204 VSS.n6202 0.258595
R71447 VSS.n6459 VSS.n6458 0.252283
R71448 VSS.n439 VSS.n143 0.252283
R71449 VSS.n6447 VSS.n6446 0.235081
R71450 VSS.n436 VSS.n145 0.233167
R71451 VSS.n6465 VSS.n3 0.231338
R71452 VSS.n6444 VSS.n6443 0.231338
R71453 VSS.n6243 VSS.n6242 0.231338
R71454 DVSS VSS.n1890 0.222172
R71455 VSS.n1894 DVSS 0.222172
R71456 VSS.n4140 VSS.n4139 0.2201
R71457 VSS.n4140 VSS.n548 0.2201
R71458 VSS.n4153 VSS.n548 0.2201
R71459 VSS.n4154 VSS.n4153 0.2201
R71460 VSS.n4154 VSS.n544 0.2201
R71461 VSS.n4167 VSS.n544 0.2201
R71462 VSS.n4168 VSS.n4167 0.2201
R71463 VSS.n4168 VSS.n539 0.2201
R71464 VSS.n4194 VSS.n539 0.2201
R71465 VSS.n4198 VSS.n534 0.2201
R71466 VSS.n534 VSS.n533 0.2201
R71467 VSS.n533 VSS.n525 0.2201
R71468 VSS.n525 VSS.n523 0.2201
R71469 VSS.n523 VSS.n522 0.2201
R71470 VSS.n522 VSS.n514 0.2201
R71471 VSS.n514 VSS.n512 0.2201
R71472 VSS.n512 VSS.n503 0.2201
R71473 VSS.n6136 VSS.n503 0.2201
R71474 VSS.n4782 VSS.n4781 0.2201
R71475 VSS.n4782 VSS.n4482 0.2201
R71476 VSS.n4795 VSS.n4482 0.2201
R71477 VSS.n4144 VSS.n551 0.2201
R71478 VSS.n4145 VSS.n4144 0.2201
R71479 VSS.n4145 VSS.n547 0.2201
R71480 VSS.n4158 VSS.n547 0.2201
R71481 VSS.n4159 VSS.n4158 0.2201
R71482 VSS.n4159 VSS.n543 0.2201
R71483 VSS.n4172 VSS.n543 0.2201
R71484 VSS.n4173 VSS.n4172 0.2201
R71485 VSS.n4173 VSS.n540 0.2201
R71486 VSS.n4205 VSS.n4204 0.2201
R71487 VSS.n4205 VSS.n524 0.2201
R71488 VSS.n4220 VSS.n524 0.2201
R71489 VSS.n4221 VSS.n4220 0.2201
R71490 VSS.n4221 VSS.n513 0.2201
R71491 VSS.n4236 VSS.n513 0.2201
R71492 VSS.n4240 VSS.n4236 0.2201
R71493 VSS.n4240 VSS.n4239 0.2201
R71494 VSS.n4239 VSS.n504 0.2201
R71495 VSS.n4786 VSS.n4486 0.2201
R71496 VSS.n4787 VSS.n4786 0.2201
R71497 VSS.n4787 VSS.n4483 0.2201
R71498 VSS.n6186 VSS.n6185 0.2201
R71499 VSS.n6185 VSS.n6184 0.2201
R71500 VSS.n6184 VSS.n6183 0.2201
R71501 VSS.n6183 VSS.n6182 0.2201
R71502 VSS.n6182 VSS.n6181 0.2201
R71503 VSS.n6181 VSS.n6180 0.2201
R71504 VSS.n6180 VSS.n6179 0.2201
R71505 VSS.n6179 VSS.n6178 0.2201
R71506 VSS.n6178 VSS.n6177 0.2201
R71507 VSS.n4211 VSS.n528 0.2201
R71508 VSS.n4212 VSS.n4211 0.2201
R71509 VSS.n4212 VSS.n517 0.2201
R71510 VSS.n4227 VSS.n517 0.2201
R71511 VSS.n4228 VSS.n4227 0.2201
R71512 VSS.n4228 VSS.n509 0.2201
R71513 VSS.n4246 VSS.n509 0.2201
R71514 VSS.n4247 VSS.n4246 0.2201
R71515 VSS.n4247 VSS.n506 0.2201
R71516 VSS.n6112 VSS.n6111 0.2201
R71517 VSS.n6111 VSS.n6110 0.2201
R71518 VSS.n6110 VSS.n6109 0.2201
R71519 VSS.n6162 VSS.n6161 0.2201
R71520 VSS.n6163 VSS.n6162 0.2201
R71521 VSS.n6164 VSS.n6163 0.2201
R71522 VSS.n6165 VSS.n6164 0.2201
R71523 VSS.n6166 VSS.n6165 0.2201
R71524 VSS.n6167 VSS.n6166 0.2201
R71525 VSS.n6168 VSS.n6167 0.2201
R71526 VSS.n6169 VSS.n6168 0.2201
R71527 VSS.n6170 VSS.n6169 0.2201
R71528 VSS.n4199 VSS.n526 0.2201
R71529 VSS.n4214 VSS.n526 0.2201
R71530 VSS.n4215 VSS.n4214 0.2201
R71531 VSS.n4215 VSS.n515 0.2201
R71532 VSS.n4230 VSS.n515 0.2201
R71533 VSS.n4231 VSS.n4230 0.2201
R71534 VSS.n4231 VSS.n507 0.2201
R71535 VSS.n4249 VSS.n507 0.2201
R71536 VSS.n6131 VSS.n4249 0.2201
R71537 VSS.n6091 VSS.n6090 0.2201
R71538 VSS.n6092 VSS.n6091 0.2201
R71539 VSS.n6093 VSS.n6092 0.2201
R71540 VSS.n3709 VSS.n3672 0.214786
R71541 VSS.n3691 VSS.n3689 0.214786
R71542 VSS.n3692 VSS.n3688 0.214786
R71543 VSS.n3687 VSS.n3686 0.214786
R71544 VSS.n3696 VSS.n3685 0.214786
R71545 VSS.n3697 VSS.n3684 0.214786
R71546 VSS.n3698 VSS.n3683 0.214786
R71547 VSS.n3682 VSS.n3680 0.214786
R71548 VSS.n3702 VSS.n3679 0.214786
R71549 VSS.n3703 VSS.n3678 0.214786
R71550 VSS.n3704 VSS.n3677 0.214786
R71551 VSS.n3676 VSS.n3674 0.214786
R71552 VSS.n3708 VSS.n3673 0.214786
R71553 VSS.n2132 VSS.n2092 0.214786
R71554 VSS.n2131 VSS.n2093 0.214786
R71555 VSS.n2096 VSS.n2094 0.214786
R71556 VSS.n2127 VSS.n2097 0.214786
R71557 VSS.n2126 VSS.n2098 0.214786
R71558 VSS.n2125 VSS.n2099 0.214786
R71559 VSS.n2102 VSS.n2100 0.214786
R71560 VSS.n2121 VSS.n2103 0.214786
R71561 VSS.n2120 VSS.n2104 0.214786
R71562 VSS.n2119 VSS.n2105 0.214786
R71563 VSS.n2108 VSS.n2106 0.214786
R71564 VSS.n2115 VSS.n2109 0.214786
R71565 VSS.n2114 VSS.n2110 0.214786
R71566 VSS.n2113 VSS.n2111 0.214786
R71567 VSS.n966 VSS.n965 0.214786
R71568 VSS.n3537 VSS.n3536 0.214786
R71569 VSS.n3538 VSS.n964 0.214786
R71570 VSS.n3540 VSS.n3539 0.214786
R71571 VSS.n962 VSS.n961 0.214786
R71572 VSS.n3545 VSS.n3544 0.214786
R71573 VSS.n3546 VSS.n960 0.214786
R71574 VSS.n3548 VSS.n3547 0.214786
R71575 VSS.n958 VSS.n957 0.214786
R71576 VSS.n3553 VSS.n3552 0.214786
R71577 VSS.n3554 VSS.n956 0.214786
R71578 VSS.n3556 VSS.n3555 0.214786
R71579 VSS.n954 VSS.n953 0.214786
R71580 VSS.n3561 VSS.n3560 0.214786
R71581 VSS.n3562 VSS.n952 0.214786
R71582 VSS.n3564 VSS.n3563 0.214786
R71583 VSS.n950 VSS.n949 0.214786
R71584 VSS.n3570 VSS.n3569 0.214786
R71585 VSS.n3571 VSS.n948 0.214786
R71586 VSS.n3575 VSS.n3572 0.214786
R71587 VSS.n3574 VSS.n3573 0.214786
R71588 VSS.n910 VSS.n909 0.214786
R71589 VSS.n3595 VSS.n3594 0.214786
R71590 VSS.n3596 VSS.n908 0.214786
R71591 VSS.n3598 VSS.n3597 0.214786
R71592 VSS.n906 VSS.n905 0.214786
R71593 VSS.n3603 VSS.n3602 0.214786
R71594 VSS.n3604 VSS.n904 0.214786
R71595 VSS.n3606 VSS.n3605 0.214786
R71596 VSS.n902 VSS.n901 0.214786
R71597 VSS.n3611 VSS.n3610 0.214786
R71598 VSS.n3612 VSS.n900 0.214786
R71599 VSS.n3614 VSS.n3613 0.214786
R71600 VSS.n898 VSS.n897 0.214786
R71601 VSS.n3619 VSS.n3618 0.214786
R71602 VSS.n3620 VSS.n896 0.214786
R71603 VSS.n3624 VSS.n3621 0.214786
R71604 VSS.n3623 VSS.n3622 0.214786
R71605 VSS.n880 VSS.n879 0.214786
R71606 VSS.n3644 VSS.n3643 0.214786
R71607 VSS.n3645 VSS.n878 0.214786
R71608 VSS.n3647 VSS.n3646 0.214786
R71609 VSS.n876 VSS.n875 0.214786
R71610 VSS.n3652 VSS.n3651 0.214786
R71611 VSS.n3653 VSS.n874 0.214786
R71612 VSS.n3655 VSS.n3654 0.214786
R71613 VSS.n872 VSS.n871 0.214786
R71614 VSS.n3660 VSS.n3659 0.214786
R71615 VSS.n3661 VSS.n870 0.214786
R71616 VSS.n3663 VSS.n3662 0.214786
R71617 VSS.n868 VSS.n867 0.214786
R71618 VSS.n3668 VSS.n3667 0.214786
R71619 VSS.n3669 VSS.n866 0.214786
R71620 VSS.n3711 VSS.n3670 0.214786
R71621 VSS.n3710 VSS.n3671 0.214786
R71622 VSS.n3693 VSS.n3692 0.214786
R71623 VSS.n3694 VSS.n3686 0.214786
R71624 VSS.n3696 VSS.n3695 0.214786
R71625 VSS.n3697 VSS.n3681 0.214786
R71626 VSS.n3699 VSS.n3698 0.214786
R71627 VSS.n3700 VSS.n3680 0.214786
R71628 VSS.n3702 VSS.n3701 0.214786
R71629 VSS.n3703 VSS.n3675 0.214786
R71630 VSS.n3705 VSS.n3704 0.214786
R71631 VSS.n3706 VSS.n3674 0.214786
R71632 VSS.n3708 VSS.n3707 0.214786
R71633 VSS.n3709 VSS.n852 0.214786
R71634 VSS.n2133 VSS.n2079 0.214786
R71635 VSS.n2132 VSS.n2080 0.214786
R71636 VSS.n2131 VSS.n2130 0.214786
R71637 VSS.n2129 VSS.n2094 0.214786
R71638 VSS.n2128 VSS.n2127 0.214786
R71639 VSS.n2126 VSS.n2095 0.214786
R71640 VSS.n2125 VSS.n2124 0.214786
R71641 VSS.n2123 VSS.n2100 0.214786
R71642 VSS.n2122 VSS.n2121 0.214786
R71643 VSS.n2120 VSS.n2101 0.214786
R71644 VSS.n2119 VSS.n2118 0.214786
R71645 VSS.n2117 VSS.n2106 0.214786
R71646 VSS.n2116 VSS.n2115 0.214786
R71647 VSS.n2114 VSS.n2107 0.214786
R71648 VSS.n2113 VSS.n2112 0.214786
R71649 VSS.n967 VSS.n966 0.214786
R71650 VSS.n3536 VSS.n3535 0.214786
R71651 VSS.n3533 VSS.n964 0.214786
R71652 VSS.n3541 VSS.n3540 0.214786
R71653 VSS.n3542 VSS.n962 0.214786
R71654 VSS.n3544 VSS.n3543 0.214786
R71655 VSS.n960 VSS.n959 0.214786
R71656 VSS.n3549 VSS.n3548 0.214786
R71657 VSS.n3550 VSS.n958 0.214786
R71658 VSS.n3552 VSS.n3551 0.214786
R71659 VSS.n956 VSS.n955 0.214786
R71660 VSS.n3557 VSS.n3556 0.214786
R71661 VSS.n3558 VSS.n954 0.214786
R71662 VSS.n3560 VSS.n3559 0.214786
R71663 VSS.n952 VSS.n951 0.214786
R71664 VSS.n3565 VSS.n3564 0.214786
R71665 VSS.n3566 VSS.n950 0.214786
R71666 VSS.n3569 VSS.n3568 0.214786
R71667 VSS.n3567 VSS.n948 0.214786
R71668 VSS.n3576 VSS.n3575 0.214786
R71669 VSS.n3574 VSS.n911 0.214786
R71670 VSS.n3592 VSS.n910 0.214786
R71671 VSS.n3594 VSS.n3593 0.214786
R71672 VSS.n908 VSS.n907 0.214786
R71673 VSS.n3599 VSS.n3598 0.214786
R71674 VSS.n3600 VSS.n906 0.214786
R71675 VSS.n3602 VSS.n3601 0.214786
R71676 VSS.n904 VSS.n903 0.214786
R71677 VSS.n3607 VSS.n3606 0.214786
R71678 VSS.n3608 VSS.n902 0.214786
R71679 VSS.n3610 VSS.n3609 0.214786
R71680 VSS.n900 VSS.n899 0.214786
R71681 VSS.n3615 VSS.n3614 0.214786
R71682 VSS.n3616 VSS.n898 0.214786
R71683 VSS.n3618 VSS.n3617 0.214786
R71684 VSS.n896 VSS.n895 0.214786
R71685 VSS.n3625 VSS.n3624 0.214786
R71686 VSS.n3623 VSS.n881 0.214786
R71687 VSS.n3641 VSS.n880 0.214786
R71688 VSS.n3643 VSS.n3642 0.214786
R71689 VSS.n878 VSS.n877 0.214786
R71690 VSS.n3648 VSS.n3647 0.214786
R71691 VSS.n3649 VSS.n876 0.214786
R71692 VSS.n3651 VSS.n3650 0.214786
R71693 VSS.n874 VSS.n873 0.214786
R71694 VSS.n3656 VSS.n3655 0.214786
R71695 VSS.n3657 VSS.n872 0.214786
R71696 VSS.n3659 VSS.n3658 0.214786
R71697 VSS.n870 VSS.n869 0.214786
R71698 VSS.n3664 VSS.n3663 0.214786
R71699 VSS.n3665 VSS.n868 0.214786
R71700 VSS.n3667 VSS.n3666 0.214786
R71701 VSS.n866 VSS.n865 0.214786
R71702 VSS.n3712 VSS.n3711 0.214786
R71703 VSS.n3710 VSS.n851 0.214786
R71704 VSS.n5961 VSS.n5960 0.214786
R71705 VSS.n5964 VSS.n5959 0.214786
R71706 VSS.n5965 VSS.n5958 0.214786
R71707 VSS.n5966 VSS.n5957 0.214786
R71708 VSS.n5956 VSS.n5954 0.214786
R71709 VSS.n5970 VSS.n5953 0.214786
R71710 VSS.n5971 VSS.n5952 0.214786
R71711 VSS.n5972 VSS.n5951 0.214786
R71712 VSS.n5950 VSS.n5948 0.214786
R71713 VSS.n5976 VSS.n5947 0.214786
R71714 VSS.n5977 VSS.n5946 0.214786
R71715 VSS.n5978 VSS.n5945 0.214786
R71716 VSS.n5982 VSS.n4906 0.214786
R71717 VSS.n5382 VSS.n5381 0.214786
R71718 VSS.n5380 VSS.n4334 0.214786
R71719 VSS.n6084 VSS.n4335 0.214786
R71720 VSS.n6083 VSS.n4336 0.214786
R71721 VSS.n6082 VSS.n4337 0.214786
R71722 VSS.n4340 VSS.n4338 0.214786
R71723 VSS.n6078 VSS.n4341 0.214786
R71724 VSS.n6077 VSS.n4342 0.214786
R71725 VSS.n6076 VSS.n4343 0.214786
R71726 VSS.n4346 VSS.n4344 0.214786
R71727 VSS.n6072 VSS.n4347 0.214786
R71728 VSS.n6071 VSS.n4348 0.214786
R71729 VSS.n6070 VSS.n4349 0.214786
R71730 VSS.n4352 VSS.n4350 0.214786
R71731 VSS.n6066 VSS.n4353 0.214786
R71732 VSS.n6065 VSS.n4354 0.214786
R71733 VSS.n6064 VSS.n4355 0.214786
R71734 VSS.n6062 VSS.n4356 0.214786
R71735 VSS.n6061 VSS.n4357 0.214786
R71736 VSS.n6060 VSS.n4358 0.214786
R71737 VSS.n6059 VSS.n4359 0.214786
R71738 VSS.n4362 VSS.n4360 0.214786
R71739 VSS.n6055 VSS.n4363 0.214786
R71740 VSS.n6054 VSS.n4364 0.214786
R71741 VSS.n6052 VSS.n4366 0.214786
R71742 VSS.n4370 VSS.n4367 0.214786
R71743 VSS.n6048 VSS.n4371 0.214786
R71744 VSS.n6047 VSS.n4372 0.214786
R71745 VSS.n6046 VSS.n4373 0.214786
R71746 VSS.n4376 VSS.n4374 0.214786
R71747 VSS.n6042 VSS.n4377 0.214786
R71748 VSS.n6041 VSS.n4378 0.214786
R71749 VSS.n6040 VSS.n4379 0.214786
R71750 VSS.n4382 VSS.n4380 0.214786
R71751 VSS.n6036 VSS.n4383 0.214786
R71752 VSS.n6035 VSS.n4384 0.214786
R71753 VSS.n4426 VSS.n4385 0.214786
R71754 VSS.n6023 VSS.n4427 0.214786
R71755 VSS.n6022 VSS.n4428 0.214786
R71756 VSS.n6021 VSS.n4429 0.214786
R71757 VSS.n4432 VSS.n4430 0.214786
R71758 VSS.n6017 VSS.n4433 0.214786
R71759 VSS.n6016 VSS.n4434 0.214786
R71760 VSS.n6015 VSS.n4435 0.214786
R71761 VSS.n4438 VSS.n4436 0.214786
R71762 VSS.n6011 VSS.n4439 0.214786
R71763 VSS.n6010 VSS.n4440 0.214786
R71764 VSS.n6009 VSS.n4441 0.214786
R71765 VSS.n6005 VSS.n4445 0.214786
R71766 VSS.n6004 VSS.n4446 0.214786
R71767 VSS.n6003 VSS.n4447 0.214786
R71768 VSS.n4450 VSS.n4448 0.214786
R71769 VSS.n5999 VSS.n4451 0.214786
R71770 VSS.n5998 VSS.n4452 0.214786
R71771 VSS.n4873 VSS.n4453 0.214786
R71772 VSS.n4875 VSS.n4874 0.214786
R71773 VSS.n4879 VSS.n4878 0.214786
R71774 VSS.n4880 VSS.n4872 0.214786
R71775 VSS.n4882 VSS.n4881 0.214786
R71776 VSS.n4870 VSS.n4869 0.214786
R71777 VSS.n4887 VSS.n4886 0.214786
R71778 VSS.n4888 VSS.n4868 0.214786
R71779 VSS.n4890 VSS.n4889 0.214786
R71780 VSS.n4866 VSS.n4865 0.214786
R71781 VSS.n4895 VSS.n4894 0.214786
R71782 VSS.n4896 VSS.n4864 0.214786
R71783 VSS.n4898 VSS.n4897 0.214786
R71784 VSS.n4862 VSS.n4861 0.214786
R71785 VSS.n4903 VSS.n4902 0.214786
R71786 VSS.n4904 VSS.n4860 0.214786
R71787 VSS.n5983 VSS.n4905 0.214786
R71788 VSS.n5924 VSS.n5922 0.214786
R71789 VSS.n5925 VSS.n5921 0.214786
R71790 VSS.n5920 VSS.n5918 0.214786
R71791 VSS.n5929 VSS.n5917 0.214786
R71792 VSS.n5930 VSS.n5916 0.214786
R71793 VSS.n5931 VSS.n5915 0.214786
R71794 VSS.n5914 VSS.n5912 0.214786
R71795 VSS.n5935 VSS.n5911 0.214786
R71796 VSS.n5936 VSS.n5910 0.214786
R71797 VSS.n5937 VSS.n5909 0.214786
R71798 VSS.n5907 VSS.n4912 0.214786
R71799 VSS.n5942 VSS.n5941 0.214786
R71800 VSS.n4913 VSS.n4911 0.214786
R71801 VSS.n5228 VSS.n5227 0.214786
R71802 VSS.n5229 VSS.n5226 0.214786
R71803 VSS.n5231 VSS.n5225 0.214786
R71804 VSS.n5232 VSS.n5224 0.214786
R71805 VSS.n5233 VSS.n5223 0.214786
R71806 VSS.n5222 VSS.n5220 0.214786
R71807 VSS.n5237 VSS.n5219 0.214786
R71808 VSS.n5238 VSS.n5218 0.214786
R71809 VSS.n5239 VSS.n5217 0.214786
R71810 VSS.n5216 VSS.n5214 0.214786
R71811 VSS.n5243 VSS.n5213 0.214786
R71812 VSS.n5244 VSS.n5212 0.214786
R71813 VSS.n5245 VSS.n5211 0.214786
R71814 VSS.n5210 VSS.n5208 0.214786
R71815 VSS.n5249 VSS.n5207 0.214786
R71816 VSS.n5250 VSS.n5206 0.214786
R71817 VSS.n5251 VSS.n5205 0.214786
R71818 VSS.n5204 VSS.n5177 0.214786
R71819 VSS.n5648 VSS.n5176 0.214786
R71820 VSS.n5649 VSS.n5175 0.214786
R71821 VSS.n5650 VSS.n5174 0.214786
R71822 VSS.n5172 VSS.n5170 0.214786
R71823 VSS.n5655 VSS.n5654 0.214786
R71824 VSS.n5557 VSS.n5169 0.214786
R71825 VSS.n5558 VSS.n5555 0.214786
R71826 VSS.n5559 VSS.n5554 0.214786
R71827 VSS.n5553 VSS.n5551 0.214786
R71828 VSS.n5563 VSS.n5550 0.214786
R71829 VSS.n5564 VSS.n5549 0.214786
R71830 VSS.n5565 VSS.n5548 0.214786
R71831 VSS.n5547 VSS.n5545 0.214786
R71832 VSS.n5569 VSS.n5544 0.214786
R71833 VSS.n5570 VSS.n5543 0.214786
R71834 VSS.n5571 VSS.n5542 0.214786
R71835 VSS.n5541 VSS.n5451 0.214786
R71836 VSS.n5585 VSS.n5450 0.214786
R71837 VSS.n5586 VSS.n5449 0.214786
R71838 VSS.n5448 VSS.n5446 0.214786
R71839 VSS.n5590 VSS.n5445 0.214786
R71840 VSS.n5591 VSS.n5444 0.214786
R71841 VSS.n5592 VSS.n5443 0.214786
R71842 VSS.n5442 VSS.n5440 0.214786
R71843 VSS.n5596 VSS.n5439 0.214786
R71844 VSS.n5597 VSS.n5438 0.214786
R71845 VSS.n5598 VSS.n5437 0.214786
R71846 VSS.n5435 VSS.n5434 0.214786
R71847 VSS.n5603 VSS.n5602 0.214786
R71848 VSS.n5606 VSS.n5605 0.214786
R71849 VSS.n5431 VSS.n5429 0.214786
R71850 VSS.n5610 VSS.n5428 0.214786
R71851 VSS.n5611 VSS.n5427 0.214786
R71852 VSS.n5612 VSS.n5426 0.214786
R71853 VSS.n5425 VSS.n5313 0.214786
R71854 VSS.n5424 VSS.n5423 0.214786
R71855 VSS.n5422 VSS.n5314 0.214786
R71856 VSS.n5416 VSS.n5315 0.214786
R71857 VSS.n5418 VSS.n5417 0.214786
R71858 VSS.n5415 VSS.n5317 0.214786
R71859 VSS.n5414 VSS.n5413 0.214786
R71860 VSS.n5319 VSS.n5318 0.214786
R71861 VSS.n5409 VSS.n5408 0.214786
R71862 VSS.n5407 VSS.n5321 0.214786
R71863 VSS.n5406 VSS.n5405 0.214786
R71864 VSS.n5323 VSS.n5322 0.214786
R71865 VSS.n5401 VSS.n5400 0.214786
R71866 VSS.n5399 VSS.n5325 0.214786
R71867 VSS.n5398 VSS.n5397 0.214786
R71868 VSS.n5394 VSS.n5326 0.214786
R71869 VSS.n5393 VSS.n5392 0.214786
R71870 VSS.n5391 VSS.n5327 0.214786
R71871 VSS.n5390 VSS.n5389 0.214786
R71872 VSS.n5887 VSS.n5885 0.214786
R71873 VSS.n5888 VSS.n5884 0.214786
R71874 VSS.n5883 VSS.n5882 0.214786
R71875 VSS.n5892 VSS.n5881 0.214786
R71876 VSS.n5893 VSS.n5880 0.214786
R71877 VSS.n5894 VSS.n5879 0.214786
R71878 VSS.n5878 VSS.n5876 0.214786
R71879 VSS.n5898 VSS.n5875 0.214786
R71880 VSS.n5899 VSS.n5874 0.214786
R71881 VSS.n5900 VSS.n5873 0.214786
R71882 VSS.n5872 VSS.n4916 0.214786
R71883 VSS.n5904 VSS.n4915 0.214786
R71884 VSS.n5688 VSS.n4914 0.214786
R71885 VSS.n5690 VSS.n5689 0.214786
R71886 VSS.n5691 VSS.n5687 0.214786
R71887 VSS.n5686 VSS.n5685 0.214786
R71888 VSS.n5695 VSS.n5684 0.214786
R71889 VSS.n5696 VSS.n5683 0.214786
R71890 VSS.n5697 VSS.n5682 0.214786
R71891 VSS.n5681 VSS.n5679 0.214786
R71892 VSS.n5701 VSS.n5678 0.214786
R71893 VSS.n5702 VSS.n5677 0.214786
R71894 VSS.n5703 VSS.n5676 0.214786
R71895 VSS.n5675 VSS.n5673 0.214786
R71896 VSS.n5707 VSS.n5672 0.214786
R71897 VSS.n5708 VSS.n5671 0.214786
R71898 VSS.n5709 VSS.n5670 0.214786
R71899 VSS.n5669 VSS.n5667 0.214786
R71900 VSS.n5713 VSS.n5666 0.214786
R71901 VSS.n5714 VSS.n5665 0.214786
R71902 VSS.n5715 VSS.n5664 0.214786
R71903 VSS.n5716 VSS.n5663 0.214786
R71904 VSS.n5717 VSS.n5662 0.214786
R71905 VSS.n5720 VSS.n5661 0.214786
R71906 VSS.n5721 VSS.n5660 0.214786
R71907 VSS.n5722 VSS.n5659 0.214786
R71908 VSS.n5657 VSS.n5165 0.214786
R71909 VSS.n5727 VSS.n5164 0.214786
R71910 VSS.n5728 VSS.n5163 0.214786
R71911 VSS.n5729 VSS.n5162 0.214786
R71912 VSS.n5161 VSS.n5159 0.214786
R71913 VSS.n5733 VSS.n5158 0.214786
R71914 VSS.n5734 VSS.n5157 0.214786
R71915 VSS.n5735 VSS.n5156 0.214786
R71916 VSS.n5155 VSS.n5153 0.214786
R71917 VSS.n5739 VSS.n5152 0.214786
R71918 VSS.n5740 VSS.n5151 0.214786
R71919 VSS.n5741 VSS.n5150 0.214786
R71920 VSS.n5743 VSS.n5149 0.214786
R71921 VSS.n5744 VSS.n5148 0.214786
R71922 VSS.n5147 VSS.n5146 0.214786
R71923 VSS.n5748 VSS.n5145 0.214786
R71924 VSS.n5749 VSS.n5144 0.214786
R71925 VSS.n5750 VSS.n5143 0.214786
R71926 VSS.n5142 VSS.n5140 0.214786
R71927 VSS.n5754 VSS.n5139 0.214786
R71928 VSS.n5755 VSS.n5138 0.214786
R71929 VSS.n5756 VSS.n5137 0.214786
R71930 VSS.n5136 VSS.n5133 0.214786
R71931 VSS.n5760 VSS.n5132 0.214786
R71932 VSS.n5762 VSS.n5131 0.214786
R71933 VSS.n5763 VSS.n5130 0.214786
R71934 VSS.n5129 VSS.n5127 0.214786
R71935 VSS.n5767 VSS.n5126 0.214786
R71936 VSS.n5768 VSS.n5125 0.214786
R71937 VSS.n5769 VSS.n5124 0.214786
R71938 VSS.n5770 VSS.n5123 0.214786
R71939 VSS.n5351 VSS.n5122 0.214786
R71940 VSS.n5354 VSS.n5352 0.214786
R71941 VSS.n5355 VSS.n5350 0.214786
R71942 VSS.n5356 VSS.n5349 0.214786
R71943 VSS.n5348 VSS.n5346 0.214786
R71944 VSS.n5360 VSS.n5345 0.214786
R71945 VSS.n5361 VSS.n5344 0.214786
R71946 VSS.n5362 VSS.n5343 0.214786
R71947 VSS.n5342 VSS.n5340 0.214786
R71948 VSS.n5366 VSS.n5339 0.214786
R71949 VSS.n5367 VSS.n5338 0.214786
R71950 VSS.n5368 VSS.n5337 0.214786
R71951 VSS.n5336 VSS.n5334 0.214786
R71952 VSS.n5372 VSS.n5333 0.214786
R71953 VSS.n5373 VSS.n5332 0.214786
R71954 VSS.n5374 VSS.n5331 0.214786
R71955 VSS.n5376 VSS.n5375 0.214786
R71956 VSS.n5375 VSS.n4982 0.214786
R71957 VSS.n5374 VSS.n4990 0.214786
R71958 VSS.n5373 VSS.n5007 0.214786
R71959 VSS.n5372 VSS.n5371 0.214786
R71960 VSS.n5370 VSS.n5334 0.214786
R71961 VSS.n5369 VSS.n5368 0.214786
R71962 VSS.n5367 VSS.n5335 0.214786
R71963 VSS.n5366 VSS.n5365 0.214786
R71964 VSS.n5364 VSS.n5340 0.214786
R71965 VSS.n5363 VSS.n5362 0.214786
R71966 VSS.n5361 VSS.n5341 0.214786
R71967 VSS.n5360 VSS.n5359 0.214786
R71968 VSS.n5358 VSS.n5346 0.214786
R71969 VSS.n5357 VSS.n5356 0.214786
R71970 VSS.n5355 VSS.n5347 0.214786
R71971 VSS.n5354 VSS.n5353 0.214786
R71972 VSS.n5122 VSS.n5121 0.214786
R71973 VSS.n5771 VSS.n5770 0.214786
R71974 VSS.n5769 VSS.n5082 0.214786
R71975 VSS.n5768 VSS.n5091 0.214786
R71976 VSS.n5767 VSS.n5766 0.214786
R71977 VSS.n5765 VSS.n5127 0.214786
R71978 VSS.n5764 VSS.n5763 0.214786
R71979 VSS.n5762 VSS.n5128 0.214786
R71980 VSS.n5760 VSS.n5759 0.214786
R71981 VSS.n5758 VSS.n5133 0.214786
R71982 VSS.n5757 VSS.n5756 0.214786
R71983 VSS.n5755 VSS.n5135 0.214786
R71984 VSS.n5754 VSS.n5753 0.214786
R71985 VSS.n5752 VSS.n5140 0.214786
R71986 VSS.n5751 VSS.n5750 0.214786
R71987 VSS.n5749 VSS.n5141 0.214786
R71988 VSS.n5748 VSS.n5747 0.214786
R71989 VSS.n5746 VSS.n5146 0.214786
R71990 VSS.n5745 VSS.n5744 0.214786
R71991 VSS.n5743 VSS.n5742 0.214786
R71992 VSS.n5741 VSS.n5029 0.214786
R71993 VSS.n5740 VSS.n5035 0.214786
R71994 VSS.n5739 VSS.n5738 0.214786
R71995 VSS.n5737 VSS.n5153 0.214786
R71996 VSS.n5736 VSS.n5735 0.214786
R71997 VSS.n5734 VSS.n5154 0.214786
R71998 VSS.n5733 VSS.n5732 0.214786
R71999 VSS.n5731 VSS.n5159 0.214786
R72000 VSS.n5730 VSS.n5729 0.214786
R72001 VSS.n5728 VSS.n5160 0.214786
R72002 VSS.n5727 VSS.n5726 0.214786
R72003 VSS.n5725 VSS.n5165 0.214786
R72004 VSS.n5723 VSS.n5722 0.214786
R72005 VSS.n5721 VSS.n5166 0.214786
R72006 VSS.n5720 VSS.n5719 0.214786
R72007 VSS.n5718 VSS.n5717 0.214786
R72008 VSS.n5716 VSS.n5070 0.214786
R72009 VSS.n5715 VSS.n5054 0.214786
R72010 VSS.n5714 VSS.n5064 0.214786
R72011 VSS.n5713 VSS.n5712 0.214786
R72012 VSS.n5711 VSS.n5667 0.214786
R72013 VSS.n5710 VSS.n5709 0.214786
R72014 VSS.n5708 VSS.n5668 0.214786
R72015 VSS.n5707 VSS.n5706 0.214786
R72016 VSS.n5705 VSS.n5673 0.214786
R72017 VSS.n5704 VSS.n5703 0.214786
R72018 VSS.n5702 VSS.n5674 0.214786
R72019 VSS.n5701 VSS.n5700 0.214786
R72020 VSS.n5699 VSS.n5679 0.214786
R72021 VSS.n5698 VSS.n5697 0.214786
R72022 VSS.n5696 VSS.n5680 0.214786
R72023 VSS.n5695 VSS.n5694 0.214786
R72024 VSS.n5693 VSS.n5685 0.214786
R72025 VSS.n5692 VSS.n5691 0.214786
R72026 VSS.n5690 VSS.n4917 0.214786
R72027 VSS.n5869 VSS.n4914 0.214786
R72028 VSS.n5904 VSS.n5903 0.214786
R72029 VSS.n5902 VSS.n4916 0.214786
R72030 VSS.n5901 VSS.n5900 0.214786
R72031 VSS.n5899 VSS.n5871 0.214786
R72032 VSS.n5898 VSS.n5897 0.214786
R72033 VSS.n5896 VSS.n5876 0.214786
R72034 VSS.n5895 VSS.n5894 0.214786
R72035 VSS.n5893 VSS.n5877 0.214786
R72036 VSS.n5892 VSS.n5891 0.214786
R72037 VSS.n5890 VSS.n5882 0.214786
R72038 VSS.n5889 VSS.n5888 0.214786
R72039 VSS.n5389 VSS.n5274 0.214786
R72040 VSS.n5327 VSS.n5260 0.214786
R72041 VSS.n5393 VSS.n5270 0.214786
R72042 VSS.n5395 VSS.n5394 0.214786
R72043 VSS.n5397 VSS.n5396 0.214786
R72044 VSS.n5325 VSS.n5324 0.214786
R72045 VSS.n5402 VSS.n5401 0.214786
R72046 VSS.n5403 VSS.n5323 0.214786
R72047 VSS.n5405 VSS.n5404 0.214786
R72048 VSS.n5321 VSS.n5320 0.214786
R72049 VSS.n5410 VSS.n5409 0.214786
R72050 VSS.n5411 VSS.n5319 0.214786
R72051 VSS.n5413 VSS.n5412 0.214786
R72052 VSS.n5317 VSS.n5316 0.214786
R72053 VSS.n5419 VSS.n5418 0.214786
R72054 VSS.n5420 VSS.n5315 0.214786
R72055 VSS.n5422 VSS.n5421 0.214786
R72056 VSS.n5423 VSS.n5289 0.214786
R72057 VSS.n5313 VSS.n5297 0.214786
R72058 VSS.n5613 VSS.n5612 0.214786
R72059 VSS.n5611 VSS.n5312 0.214786
R72060 VSS.n5610 VSS.n5609 0.214786
R72061 VSS.n5608 VSS.n5429 0.214786
R72062 VSS.n5607 VSS.n5606 0.214786
R72063 VSS.n5602 VSS.n5601 0.214786
R72064 VSS.n5600 VSS.n5435 0.214786
R72065 VSS.n5599 VSS.n5598 0.214786
R72066 VSS.n5597 VSS.n5436 0.214786
R72067 VSS.n5596 VSS.n5595 0.214786
R72068 VSS.n5594 VSS.n5440 0.214786
R72069 VSS.n5593 VSS.n5592 0.214786
R72070 VSS.n5591 VSS.n5441 0.214786
R72071 VSS.n5590 VSS.n5589 0.214786
R72072 VSS.n5588 VSS.n5446 0.214786
R72073 VSS.n5587 VSS.n5586 0.214786
R72074 VSS.n5585 VSS.n5584 0.214786
R72075 VSS.n5505 VSS.n5451 0.214786
R72076 VSS.n5572 VSS.n5571 0.214786
R72077 VSS.n5570 VSS.n5540 0.214786
R72078 VSS.n5569 VSS.n5568 0.214786
R72079 VSS.n5567 VSS.n5545 0.214786
R72080 VSS.n5566 VSS.n5565 0.214786
R72081 VSS.n5564 VSS.n5546 0.214786
R72082 VSS.n5563 VSS.n5562 0.214786
R72083 VSS.n5561 VSS.n5551 0.214786
R72084 VSS.n5560 VSS.n5559 0.214786
R72085 VSS.n5558 VSS.n5552 0.214786
R72086 VSS.n5557 VSS.n5556 0.214786
R72087 VSS.n5654 VSS.n5653 0.214786
R72088 VSS.n5652 VSS.n5172 0.214786
R72089 VSS.n5651 VSS.n5650 0.214786
R72090 VSS.n5649 VSS.n5173 0.214786
R72091 VSS.n5648 VSS.n5647 0.214786
R72092 VSS.n5186 VSS.n5177 0.214786
R72093 VSS.n5252 VSS.n5251 0.214786
R72094 VSS.n5250 VSS.n5203 0.214786
R72095 VSS.n5249 VSS.n5248 0.214786
R72096 VSS.n5247 VSS.n5208 0.214786
R72097 VSS.n5246 VSS.n5245 0.214786
R72098 VSS.n5244 VSS.n5209 0.214786
R72099 VSS.n5243 VSS.n5242 0.214786
R72100 VSS.n5241 VSS.n5214 0.214786
R72101 VSS.n5240 VSS.n5239 0.214786
R72102 VSS.n5238 VSS.n5215 0.214786
R72103 VSS.n5237 VSS.n5236 0.214786
R72104 VSS.n5235 VSS.n5220 0.214786
R72105 VSS.n5234 VSS.n5233 0.214786
R72106 VSS.n5232 VSS.n5221 0.214786
R72107 VSS.n5231 VSS.n5230 0.214786
R72108 VSS.n5229 VSS.n4948 0.214786
R72109 VSS.n5228 VSS.n4956 0.214786
R72110 VSS.n4973 VSS.n4913 0.214786
R72111 VSS.n5941 VSS.n5940 0.214786
R72112 VSS.n5939 VSS.n5907 0.214786
R72113 VSS.n5938 VSS.n5937 0.214786
R72114 VSS.n5936 VSS.n5908 0.214786
R72115 VSS.n5935 VSS.n5934 0.214786
R72116 VSS.n5933 VSS.n5912 0.214786
R72117 VSS.n5932 VSS.n5931 0.214786
R72118 VSS.n5930 VSS.n5913 0.214786
R72119 VSS.n5929 VSS.n5928 0.214786
R72120 VSS.n5927 VSS.n5918 0.214786
R72121 VSS.n5926 VSS.n5925 0.214786
R72122 VSS.n5924 VSS.n5919 0.214786
R72123 VSS.n5964 VSS.n5963 0.214786
R72124 VSS.n5965 VSS.n5955 0.214786
R72125 VSS.n5967 VSS.n5966 0.214786
R72126 VSS.n5968 VSS.n5954 0.214786
R72127 VSS.n5970 VSS.n5969 0.214786
R72128 VSS.n5971 VSS.n5949 0.214786
R72129 VSS.n5973 VSS.n5972 0.214786
R72130 VSS.n5974 VSS.n5948 0.214786
R72131 VSS.n5976 VSS.n5975 0.214786
R72132 VSS.n5977 VSS.n4909 0.214786
R72133 VSS.n5979 VSS.n5978 0.214786
R72134 VSS.n5982 VSS.n5981 0.214786
R72135 VSS.n5381 VSS.n4311 0.214786
R72136 VSS.n4334 VSS.n4319 0.214786
R72137 VSS.n6085 VSS.n6084 0.214786
R72138 VSS.n6083 VSS.n4333 0.214786
R72139 VSS.n6082 VSS.n6081 0.214786
R72140 VSS.n6080 VSS.n4338 0.214786
R72141 VSS.n6079 VSS.n6078 0.214786
R72142 VSS.n6077 VSS.n4339 0.214786
R72143 VSS.n6076 VSS.n6075 0.214786
R72144 VSS.n6074 VSS.n4344 0.214786
R72145 VSS.n6073 VSS.n6072 0.214786
R72146 VSS.n6071 VSS.n4345 0.214786
R72147 VSS.n6070 VSS.n6069 0.214786
R72148 VSS.n6068 VSS.n4350 0.214786
R72149 VSS.n6067 VSS.n6066 0.214786
R72150 VSS.n6065 VSS.n4351 0.214786
R72151 VSS.n6064 VSS.n6063 0.214786
R72152 VSS.n6062 VSS.n4294 0.214786
R72153 VSS.n6061 VSS.n4280 0.214786
R72154 VSS.n6060 VSS.n4287 0.214786
R72155 VSS.n6059 VSS.n6058 0.214786
R72156 VSS.n6057 VSS.n4360 0.214786
R72157 VSS.n6056 VSS.n6055 0.214786
R72158 VSS.n6054 VSS.n4361 0.214786
R72159 VSS.n6052 VSS.n6051 0.214786
R72160 VSS.n6050 VSS.n4367 0.214786
R72161 VSS.n6049 VSS.n6048 0.214786
R72162 VSS.n6047 VSS.n4369 0.214786
R72163 VSS.n6046 VSS.n6045 0.214786
R72164 VSS.n6044 VSS.n4374 0.214786
R72165 VSS.n6043 VSS.n6042 0.214786
R72166 VSS.n6041 VSS.n4375 0.214786
R72167 VSS.n6040 VSS.n6039 0.214786
R72168 VSS.n6038 VSS.n4380 0.214786
R72169 VSS.n6037 VSS.n6036 0.214786
R72170 VSS.n6035 VSS.n6034 0.214786
R72171 VSS.n4422 VSS.n4385 0.214786
R72172 VSS.n6024 VSS.n6023 0.214786
R72173 VSS.n6022 VSS.n4425 0.214786
R72174 VSS.n6021 VSS.n6020 0.214786
R72175 VSS.n6019 VSS.n4430 0.214786
R72176 VSS.n6018 VSS.n6017 0.214786
R72177 VSS.n6016 VSS.n4431 0.214786
R72178 VSS.n6015 VSS.n6014 0.214786
R72179 VSS.n6013 VSS.n4436 0.214786
R72180 VSS.n6012 VSS.n6011 0.214786
R72181 VSS.n6010 VSS.n4437 0.214786
R72182 VSS.n6009 VSS.n6008 0.214786
R72183 VSS.n6006 VSS.n6005 0.214786
R72184 VSS.n6004 VSS.n4444 0.214786
R72185 VSS.n6003 VSS.n6002 0.214786
R72186 VSS.n6001 VSS.n4448 0.214786
R72187 VSS.n6000 VSS.n5999 0.214786
R72188 VSS.n5998 VSS.n5997 0.214786
R72189 VSS.n4460 VSS.n4453 0.214786
R72190 VSS.n4876 VSS.n4875 0.214786
R72191 VSS.n4878 VSS.n4877 0.214786
R72192 VSS.n4872 VSS.n4871 0.214786
R72193 VSS.n4883 VSS.n4882 0.214786
R72194 VSS.n4884 VSS.n4870 0.214786
R72195 VSS.n4886 VSS.n4885 0.214786
R72196 VSS.n4868 VSS.n4867 0.214786
R72197 VSS.n4891 VSS.n4890 0.214786
R72198 VSS.n4892 VSS.n4866 0.214786
R72199 VSS.n4894 VSS.n4893 0.214786
R72200 VSS.n4864 VSS.n4863 0.214786
R72201 VSS.n4899 VSS.n4898 0.214786
R72202 VSS.n4900 VSS.n4862 0.214786
R72203 VSS.n4902 VSS.n4901 0.214786
R72204 VSS.n4860 VSS.n4474 0.214786
R72205 VSS.n5984 VSS.n5983 0.214786
R72206 VSS.n6138 VSS.n6136 0.2003
R72207 VSS.n4767 VSS.n504 0.2003
R72208 VSS.n6120 VSS.n506 0.2003
R72209 VSS.n6131 VSS.n6130 0.2003
R72210 VSS.n6446 VSS.n20 0.199895
R72211 VSS.n132 VSS.n20 0.199543
R72212 DVSS VSS.n4136 0.191946
R72213 DVSS VSS.n4141 0.191946
R72214 DVSS VSS.n550 0.191946
R72215 DVSS VSS.n4150 0.191946
R72216 DVSS VSS.n4155 0.191946
R72217 DVSS VSS.n546 0.191946
R72218 DVSS VSS.n4164 0.191946
R72219 DVSS VSS.n4169 0.191946
R72220 DVSS VSS.n542 0.191946
R72221 DVSS VSS.n4191 0.191946
R72222 DVSS VSS.n4201 0.191946
R72223 VSS.n4209 DVSS 0.191946
R72224 DVSS VSS.n527 0.191946
R72225 DVSS VSS.n4217 0.191946
R72226 VSS.n4225 DVSS 0.191946
R72227 DVSS VSS.n516 0.191946
R72228 DVSS VSS.n4233 0.191946
R72229 VSS.n4244 DVSS 0.191946
R72230 DVSS VSS.n508 0.191946
R72231 DVSS VSS.n6133 0.191946
R72232 DVSS VSS.n4512 0.191946
R72233 DVSS VSS.n4778 0.191946
R72234 DVSS VSS.n4783 0.191946
R72235 DVSS VSS.n4485 0.191946
R72236 DVSS VSS.n4792 0.191946
R72237 DVSS VSS.n4853 0.191946
R72238 DVSS VSS.n4841 0.191946
R72239 DVSS VSS.n4829 0.191946
R72240 DVSS VSS.n4817 0.191946
R72241 DVSS VSS.n4308 0.191946
R72242 DVSS VSS.n5531 0.191946
R72243 DVSS VSS.n5513 0.191946
R72244 DVSS VSS.n5286 0.191946
R72245 DVSS VSS.n5636 0.191946
R72246 DVSS VSS.n5466 0.191946
R72247 DVSS VSS.n5846 0.191946
R72248 DVSS VSS.n5789 0.191946
R72249 VSS.n5100 DVSS 0.191946
R72250 VSS.n5111 DVSS 0.191946
R72251 DVSS VSS.n5050 0.191946
R72252 VSS.n1612 VSS.n1611 0.191946
R72253 VSS.n4132 VSS.n4127 0.189567
R72254 VSS.n1888 VSS.n1887 0.186867
R72255 VSS.n1897 VSS.n1896 0.186867
R72256 VSS.n6193 VSS.n453 0.17981
R72257 VSS.n453 VSS.n451 0.17981
R72258 VSS.n4118 VSS.n4117 0.173833
R72259 VSS.n4119 VSS.n4118 0.173833
R72260 VSS.n4100 VSS.n4090 0.1679
R72261 VSS.n4104 VSS.n4103 0.1679
R72262 VSS.n6191 VSS.n456 0.1679
R72263 VSS.n2204 VSS.n454 0.1679
R72264 VSS.n4102 VSS.n560 0.159184
R72265 VSS.n131 VSS.n130 0.159115
R72266 VSS.n130 VSS.n127 0.158395
R72267 VSS.n6206 VSS.n6204 0.158395
R72268 VSS.n6208 VSS.n6206 0.158395
R72269 VSS.n6208 VSS.n6207 0.158395
R72270 VSS.n6449 VSS.n17 0.158395
R72271 VSS.n6207 VSS.n17 0.158395
R72272 VSS.n141 VSS.n127 0.158395
R72273 VSS.n2907 VSS.n2877 0.155773
R72274 VSS.n2955 VSS.n1129 0.155773
R72275 VSS.n6449 VSS.n6448 0.15017
R72276 VSS.n1427 VSS.n1142 0.149772
R72277 VSS.n6459 VSS.n6 0.146974
R72278 VSS.n440 VSS.n439 0.146974
R72279 VSS.n563 VSS.n452 0.144944
R72280 VSS.n1860 DVSS 0.144526
R72281 VSS.n3274 VSS.n3273 0.137755
R72282 VSS.n1795 DVSS 0.130618
R72283 VSS.n3034 DVSS 0.130618
R72284 VSS.n1020 DVSS 0.130618
R72285 VSS.n4059 DVSS 0.130618
R72286 VSS.n4697 DVSS 0.130618
R72287 VSS.n4781 VSS.n500 0.1283
R72288 VSS.n4519 VSS.n4486 0.1283
R72289 VSS.n6113 VSS.n6112 0.1283
R72290 VSS.n6090 VSS.n4256 0.1283
R72291 VSS.n3725 VSS.n864 0.12785
R72292 VSS.n3639 VSS.n894 0.12785
R72293 VSS.n3509 VSS.n3508 0.12785
R72294 VSS.n2147 VSS.n2068 0.12785
R72295 VSS.n1613 VSS.n1612 0.126026
R72296 VSS.n5808 DVSS 0.126026
R72297 VSS.n5109 DVSS 0.126026
R72298 VSS.n5098 DVSS 0.126026
R72299 VSS.n5790 DVSS 0.126026
R72300 VSS.n5847 DVSS 0.126026
R72301 VSS.n5468 DVSS 0.126026
R72302 VSS.n5637 DVSS 0.126026
R72303 VSS.n5524 DVSS 0.126026
R72304 VSS.n5517 DVSS 0.126026
R72305 VSS.n5535 DVSS 0.126026
R72306 VSS.n5988 DVSS 0.126026
R72307 VSS.n4818 DVSS 0.126026
R72308 VSS.n4830 DVSS 0.126026
R72309 VSS.n4842 DVSS 0.126026
R72310 VSS.n4854 DVSS 0.126026
R72311 VSS.n4793 DVSS 0.126026
R72312 VSS.n4789 DVSS 0.126026
R72313 VSS.n4784 DVSS 0.126026
R72314 VSS.n4779 DVSS 0.126026
R72315 VSS.n4772 DVSS 0.126026
R72316 VSS.n6134 DVSS 0.126026
R72317 VSS.n4237 DVSS 0.126026
R72318 VSS.n4242 DVSS 0.126026
R72319 VSS.n4234 DVSS 0.126026
R72320 VSS.n520 DVSS 0.126026
R72321 VSS.n4223 DVSS 0.126026
R72322 VSS.n4218 DVSS 0.126026
R72323 VSS.n531 DVSS 0.126026
R72324 VSS.n4207 DVSS 0.126026
R72325 VSS.n4202 DVSS 0.126026
R72326 VSS.n4192 DVSS 0.126026
R72327 VSS.n4175 DVSS 0.126026
R72328 VSS.n4170 DVSS 0.126026
R72329 VSS.n4165 DVSS 0.126026
R72330 VSS.n4161 DVSS 0.126026
R72331 VSS.n4156 DVSS 0.126026
R72332 VSS.n4151 DVSS 0.126026
R72333 VSS.n4147 DVSS 0.126026
R72334 VSS.n4142 DVSS 0.126026
R72335 VSS.n4137 DVSS 0.126026
R72336 VSS.n4135 VSS.n4134 0.124418
R72337 VSS.n2900 VSS.n2899 0.115687
R72338 VSS.n2895 VSS.n1112 0.115687
R72339 VSS.n4190 VSS.n4189 0.115687
R72340 VSS.n4183 VSS.n529 0.115687
R72341 VSS.n6216 VSS.n6199 0.115183
R72342 VSS.n2909 VSS.n2908 0.113608
R72343 VSS.n2908 VSS.n2907 0.113608
R72344 VSS.n2914 VSS.n2874 0.113608
R72345 VSS.n2955 VSS.n1123 0.113608
R72346 VSS.n2961 VSS.n1123 0.113608
R72347 VSS.n2961 VSS.n2960 0.113608
R72348 VSS.n2907 VSS.n2906 0.113608
R72349 VSS.n2906 VSS.n2874 0.113608
R72350 VSS.n1139 VSS.n1133 0.113608
R72351 VSS.n2956 VSS.n1133 0.113608
R72352 VSS.n2956 VSS.n2955 0.113608
R72353 VSS.n2910 VSS.n2909 0.113608
R72354 VSS.n2941 VSS.n1145 0.113168
R72355 DVSS VSS.n1860 0.111845
R72356 VSS.n5850 VSS.n5849 0.1112
R72357 VSS.n5076 VSS.n4977 0.1112
R72358 VSS.n5777 VSS.n4979 0.1112
R72359 VSS.n5844 VSS.n5843 0.1112
R72360 VSS.n4122 VSS.n4121 0.108833
R72361 VSS.n4121 VSS.n4120 0.108833
R72362 VSS.n1795 DVSS 0.10093
R72363 VSS.n3034 DVSS 0.10093
R72364 DVSS VSS.n1020 0.10093
R72365 VSS.n4059 DVSS 0.10093
R72366 VSS.n4697 DVSS 0.10093
R72367 VSS.n442 VSS.n126 0.100706
R72368 VSS.n438 VSS.n126 0.100706
R72369 VSS.n445 VSS.n5 0.100706
R72370 VSS.n6460 VSS.n5 0.100706
R72371 VSS.n6231 VSS.n6226 0.100706
R72372 VSS.n6232 VSS.n6231 0.100706
R72373 VSS.n6233 VSS.n6232 0.100706
R72374 VSS.n6233 VSS.n123 0.100706
R72375 VSS.n6237 VSS.n123 0.100706
R72376 VSS.n135 VSS.n132 0.100706
R72377 VSS.n4796 VSS.n4795 0.0932
R72378 VSS.n4483 VSS.n4470 0.0932
R72379 VSS.n6109 VSS.n6108 0.0932
R72380 VSS.n6094 VSS.n6093 0.0932
R72381 VSS.n6214 VSS.n6199 0.08969
R72382 VSS.n6452 VSS.n14 0.08969
R72383 VSS.n6205 VSS.n13 0.08969
R72384 VSS.n6210 VSS.n6209 0.08969
R72385 VSS.n6211 VSS.n6203 0.08969
R72386 VSS.n6213 VSS.n6212 0.08969
R72387 VSS.n139 VSS.n129 0.08969
R72388 VSS.n138 VSS.n137 0.08969
R72389 VSS.n16 VSS.n15 0.08969
R72390 VSS.n6451 VSS.n6450 0.08969
R72391 VSS.n4135 VSS.n549 0.0824403
R72392 VSS.n4148 VSS.n549 0.0824403
R72393 VSS.n4149 VSS.n4148 0.0824403
R72394 VSS.n4149 VSS.n545 0.0824403
R72395 VSS.n4162 VSS.n545 0.0824403
R72396 VSS.n4163 VSS.n4162 0.0824403
R72397 VSS.n4163 VSS.n541 0.0824403
R72398 VSS.n4176 VSS.n541 0.0824403
R72399 VSS.n4190 VSS.n4176 0.0824403
R72400 VSS.n4208 VSS.n529 0.0824403
R72401 VSS.n4208 VSS.n530 0.0824403
R72402 VSS.n530 VSS.n518 0.0824403
R72403 VSS.n4224 VSS.n518 0.0824403
R72404 VSS.n4224 VSS.n519 0.0824403
R72405 VSS.n519 VSS.n510 0.0824403
R72406 VSS.n4243 VSS.n510 0.0824403
R72407 VSS.n4243 VSS.n511 0.0824403
R72408 VSS.n511 VSS.n505 0.0824403
R72409 VSS.n4777 VSS.n4484 0.0824403
R72410 VSS.n4790 VSS.n4484 0.0824403
R72411 VSS.n4791 VSS.n4790 0.0824403
R72412 VSS.n1552 VSS.n1548 0.0788099
R72413 VSS.n446 VSS.n7 0.0785115
R72414 VSS.n443 VSS.n125 0.0785115
R72415 VSS.n5857 VSS.n5856 0.0779
R72416 VSS.n5485 VSS.n5185 0.0779
R72417 VSS.n5496 VSS.n5296 0.0779
R72418 VSS.n5492 VSS.n5281 0.0779
R72419 VSS.n6230 VSS.n6227 0.0758488
R72420 VSS.n134 VSS.n133 0.0758488
R72421 VSS.n2316 VSS.n2314 0.0758261
R72422 VSS.n3394 VSS.n849 0.0758261
R72423 VSS.n2541 VSS.n2069 0.0758261
R72424 VSS.n3399 VSS.n3098 0.0758261
R72425 VSS.n4491 VSS.n505 0.0750522
R72426 VSS.n1610 VSS.n1223 0.0734487
R72427 VSS.n1903 VSS.n1208 0.0718204
R72428 VSS.n1910 VSS.n1909 0.0718204
R72429 VSS.n2690 VSS.n1184 0.0718204
R72430 VSS.n2155 VSS.n2150 0.0718204
R72431 VSS.n4571 VSS.n4263 0.0718204
R72432 VSS.n1612 VSS.n1610 0.0702987
R72433 VSS.n6215 VSS.n6202 0.0682385
R72434 VSS.n1553 VSS.n1552 0.0652766
R72435 VSS.n3690 DVSS 0.0638222
R72436 VSS.n5962 DVSS 0.0638222
R72437 VSS.n5886 DVSS 0.0633822
R72438 VSS.n4127 VSS.n559 0.0629627
R72439 VSS.n5923 DVSS 0.0617998
R72440 VSS.n141 VSS.n140 0.061538
R72441 VSS.n140 VSS.n139 0.060427
R72442 VSS.n5923 DVSS 0.05998
R72443 VSS.n1377 VSS.n1208 0.059485
R72444 VSS.n2052 VSS.n1910 0.059485
R72445 VSS.n2691 VSS.n2690 0.059485
R72446 VSS.n2200 VSS.n2155 0.059485
R72447 VSS.n4572 VSS.n4571 0.059485
R72448 VSS.n1246 VSS.n1237 0.0569562
R72449 VSS.n1247 VSS.n1238 0.0569562
R72450 VSS.n1248 VSS.n1239 0.0569562
R72451 VSS.n1832 VSS.n1831 0.0569562
R72452 VSS.n1826 VSS.n1256 0.0569562
R72453 VSS.n1059 VSS.n1052 0.0569562
R72454 VSS.n1058 VSS.n1053 0.0569562
R72455 VSS.n1057 VSS.n1054 0.0569562
R72456 VSS.n1056 VSS.n1055 0.0569562
R72457 VSS.n1048 VSS.n999 0.0569562
R72458 VSS.n1047 VSS.n1000 0.0569562
R72459 VSS.n1046 VSS.n1001 0.0569562
R72460 VSS.n1045 VSS.n1002 0.0569562
R72461 VSS.n3713 VSS.n863 0.0569562
R72462 VSS.n3714 VSS.n862 0.0569562
R72463 VSS.n3715 VSS.n861 0.0569562
R72464 VSS.n3716 VSS.n860 0.0569562
R72465 VSS.n3717 VSS.n859 0.0569562
R72466 VSS.n3718 VSS.n858 0.0569562
R72467 VSS.n3719 VSS.n857 0.0569562
R72468 VSS.n3720 VSS.n856 0.0569562
R72469 VSS.n3721 VSS.n855 0.0569562
R72470 VSS.n3722 VSS.n854 0.0569562
R72471 VSS.n853 VSS.n850 0.0569562
R72472 VSS.n584 VSS.n577 0.0569562
R72473 VSS.n583 VSS.n578 0.0569562
R72474 VSS.n582 VSS.n579 0.0569562
R72475 VSS.n581 VSS.n580 0.0569562
R72476 VSS.n495 VSS.n494 0.0569562
R72477 VSS.n501 VSS.n496 0.0569562
R72478 VSS.n4801 VSS.n4481 0.0569562
R72479 VSS.n4803 VSS.n4480 0.0569562
R72480 VSS.n4805 VSS.n4479 0.0569562
R72481 VSS.n4807 VSS.n4478 0.0569562
R72482 VSS.n4809 VSS.n4475 0.0569562
R72483 VSS.n4477 VSS.n4473 0.0569562
R72484 VSS.n4858 VSS.n4477 0.0569562
R72485 VSS.n4858 VSS.n4476 0.0569562
R72486 VSS.n4957 VSS.n4947 0.0569562
R72487 VSS.n4974 VSS.n4958 0.0569562
R72488 VSS.n4971 VSS.n4955 0.0569562
R72489 VSS.n4969 VSS.n4953 0.0569562
R72490 VSS.n4967 VSS.n4951 0.0569562
R72491 VSS.n4965 VSS.n4962 0.0569562
R72492 VSS.n4965 VSS.n4950 0.0569562
R72493 VSS.n5854 VSS.n4963 0.0569562
R72494 VSS.n4963 VSS.n4949 0.0569562
R72495 VSS.n4939 VSS.n4926 0.0569562
R72496 VSS.n4938 VSS.n4926 0.0569562
R72497 VSS.n4940 VSS.n4924 0.0569562
R72498 VSS.n4937 VSS.n4924 0.0569562
R72499 VSS.n4941 VSS.n4922 0.0569562
R72500 VSS.n4936 VSS.n4922 0.0569562
R72501 VSS.n4942 VSS.n4920 0.0569562
R72502 VSS.n4935 VSS.n4920 0.0569562
R72503 VSS.n4934 VSS.n4919 0.0569562
R72504 VSS.n4809 VSS.n4800 0.0569562
R72505 VSS.n4807 VSS.n4799 0.0569562
R72506 VSS.n4805 VSS.n4798 0.0569562
R72507 VSS.n4803 VSS.n4797 0.0569562
R72508 VSS.n496 VSS.n495 0.0569562
R72509 VSS.n494 VSS.n493 0.0569562
R72510 VSS.n580 VSS.n574 0.0569562
R72511 VSS.n581 VSS.n579 0.0569562
R72512 VSS.n582 VSS.n578 0.0569562
R72513 VSS.n583 VSS.n577 0.0569562
R72514 VSS.n584 VSS.n576 0.0569562
R72515 VSS.n3722 VSS.n853 0.0569562
R72516 VSS.n3721 VSS.n854 0.0569562
R72517 VSS.n3720 VSS.n855 0.0569562
R72518 VSS.n3719 VSS.n856 0.0569562
R72519 VSS.n3718 VSS.n857 0.0569562
R72520 VSS.n3717 VSS.n858 0.0569562
R72521 VSS.n3716 VSS.n859 0.0569562
R72522 VSS.n3715 VSS.n860 0.0569562
R72523 VSS.n3714 VSS.n861 0.0569562
R72524 VSS.n3713 VSS.n862 0.0569562
R72525 VSS.n3724 VSS.n863 0.0569562
R72526 VSS.n3068 VSS.n1002 0.0569562
R72527 VSS.n1045 VSS.n1001 0.0569562
R72528 VSS.n1046 VSS.n1000 0.0569562
R72529 VSS.n1047 VSS.n999 0.0569562
R72530 VSS.n1048 VSS.n998 0.0569562
R72531 VSS.n1055 VSS.n1049 0.0569562
R72532 VSS.n1056 VSS.n1054 0.0569562
R72533 VSS.n1057 VSS.n1053 0.0569562
R72534 VSS.n1058 VSS.n1052 0.0569562
R72535 VSS.n1059 VSS.n1051 0.0569562
R72536 VSS.n1827 VSS.n1253 0.0569562
R72537 VSS.n1831 VSS.n1256 0.0569562
R72538 VSS.n1832 VSS.n1249 0.0569562
R72539 VSS.n1248 VSS.n1240 0.0569562
R72540 VSS.n1247 VSS.n1239 0.0569562
R72541 VSS.n1246 VSS.n1238 0.0569562
R72542 VSS.n1237 VSS.n1235 0.0569562
R72543 VSS.n4974 VSS.n4957 0.0569562
R72544 VSS.n4970 VSS.n4955 0.0569562
R72545 VSS.n4968 VSS.n4953 0.0569562
R72546 VSS.n4935 VSS.n4919 0.0569562
R72547 VSS.n1739 VSS.n1289 0.0569562
R72548 VSS.n1739 VSS.n1288 0.0569562
R72549 VSS.n1740 VSS.n1288 0.0569562
R72550 VSS.n1740 VSS.n1287 0.0569562
R72551 VSS.n1741 VSS.n1287 0.0569562
R72552 VSS.n1741 VSS.n1286 0.0569562
R72553 VSS.n1286 VSS.n1283 0.0569562
R72554 VSS.n1749 VSS.n1275 0.0569562
R72555 VSS.n1749 VSS.n1276 0.0569562
R72556 VSS.n1752 VSS.n1276 0.0569562
R72557 VSS.n1753 VSS.n1752 0.0569562
R72558 VSS.n1750 VSS.n1277 0.0569562
R72559 VSS.n2947 VSS.n1135 0.0569562
R72560 VSS.n2953 VSS.n2952 0.0569562
R72561 VSS.n1090 VSS.n1089 0.0569562
R72562 VSS.n1089 VSS.n1088 0.0569562
R72563 VSS.n1088 VSS.n1087 0.0569562
R72564 VSS.n1087 VSS.n1086 0.0569562
R72565 VSS.n2776 VSS.n975 0.0569562
R72566 VSS.n2776 VSS.n976 0.0569562
R72567 VSS.n2775 VSS.n976 0.0569562
R72568 VSS.n2775 VSS.n977 0.0569562
R72569 VSS.n2774 VSS.n977 0.0569562
R72570 VSS.n2774 VSS.n978 0.0569562
R72571 VSS.n2773 VSS.n978 0.0569562
R72572 VSS.n2773 VSS.n979 0.0569562
R72573 VSS.n979 VSS.n973 0.0569562
R72574 VSS.n3638 VSS.n893 0.0569562
R72575 VSS.n3626 VSS.n893 0.0569562
R72576 VSS.n3626 VSS.n892 0.0569562
R72577 VSS.n3627 VSS.n892 0.0569562
R72578 VSS.n3627 VSS.n891 0.0569562
R72579 VSS.n3628 VSS.n891 0.0569562
R72580 VSS.n3628 VSS.n890 0.0569562
R72581 VSS.n3629 VSS.n890 0.0569562
R72582 VSS.n3629 VSS.n889 0.0569562
R72583 VSS.n3630 VSS.n889 0.0569562
R72584 VSS.n3630 VSS.n888 0.0569562
R72585 VSS.n3631 VSS.n888 0.0569562
R72586 VSS.n3631 VSS.n887 0.0569562
R72587 VSS.n3632 VSS.n887 0.0569562
R72588 VSS.n3632 VSS.n886 0.0569562
R72589 VSS.n3633 VSS.n886 0.0569562
R72590 VSS.n3633 VSS.n885 0.0569562
R72591 VSS.n3634 VSS.n885 0.0569562
R72592 VSS.n3634 VSS.n884 0.0569562
R72593 VSS.n3635 VSS.n884 0.0569562
R72594 VSS.n3635 VSS.n883 0.0569562
R72595 VSS.n3636 VSS.n883 0.0569562
R72596 VSS.n4114 VSS.n4113 0.0569562
R72597 VSS.n4113 VSS.n4112 0.0569562
R72598 VSS.n4112 VSS.n4111 0.0569562
R72599 VSS.n4111 VSS.n4110 0.0569562
R72600 VSS.n4110 VSS.n4109 0.0569562
R72601 VSS.n4109 VSS.n4108 0.0569562
R72602 VSS.n4108 VSS.n4107 0.0569562
R72603 VSS.n4107 VSS.n4106 0.0569562
R72604 VSS.n4106 VSS.n4105 0.0569562
R72605 VSS.n4762 VSS.n4521 0.0569562
R72606 VSS.n4762 VSS.n4520 0.0569562
R72607 VSS.n4761 VSS.n4520 0.0569562
R72608 VSS.n4761 VSS.n4517 0.0569562
R72609 VSS.n4469 VSS.n4455 0.0569562
R72610 VSS.n4468 VSS.n4467 0.0569562
R72611 VSS.n4467 VSS.n4456 0.0569562
R72612 VSS.n4466 VSS.n4465 0.0569562
R72613 VSS.n4465 VSS.n4457 0.0569562
R72614 VSS.n4464 VSS.n4463 0.0569562
R72615 VSS.n4463 VSS.n4458 0.0569562
R72616 VSS.n4462 VSS.n4461 0.0569562
R72617 VSS.n4461 VSS.n4459 0.0569562
R72618 VSS.n5994 VSS.n5992 0.0569562
R72619 VSS.n5995 VSS.n5993 0.0569562
R72620 VSS.n5253 VSS.n5187 0.0569562
R72621 VSS.n5254 VSS.n5188 0.0569562
R72622 VSS.n5201 VSS.n5184 0.0569562
R72623 VSS.n5199 VSS.n5182 0.0569562
R72624 VSS.n5197 VSS.n5180 0.0569562
R72625 VSS.n5195 VSS.n5192 0.0569562
R72626 VSS.n5195 VSS.n5179 0.0569562
R72627 VSS.n5645 VSS.n5193 0.0569562
R72628 VSS.n5193 VSS.n5178 0.0569562
R72629 VSS.n5794 VSS.n5062 0.0569562
R72630 VSS.n5075 VSS.n5062 0.0569562
R72631 VSS.n5795 VSS.n5060 0.0569562
R72632 VSS.n5074 VSS.n5060 0.0569562
R72633 VSS.n5796 VSS.n5058 0.0569562
R72634 VSS.n5073 VSS.n5058 0.0569562
R72635 VSS.n5057 VSS.n5053 0.0569562
R72636 VSS.n5072 VSS.n5057 0.0569562
R72637 VSS.n5071 VSS.n5056 0.0569562
R72638 VSS.n5995 VSS.n5994 0.0569562
R72639 VSS.n5254 VSS.n5187 0.0569562
R72640 VSS.n5200 VSS.n5184 0.0569562
R72641 VSS.n5198 VSS.n5182 0.0569562
R72642 VSS.n5072 VSS.n5056 0.0569562
R72643 VSS.n1349 VSS.n1348 0.0569562
R72644 VSS.n1350 VSS.n1349 0.0569562
R72645 VSS.n1351 VSS.n1350 0.0569562
R72646 VSS.n1352 VSS.n1351 0.0569562
R72647 VSS.n1353 VSS.n1352 0.0569562
R72648 VSS.n1354 VSS.n1353 0.0569562
R72649 VSS.n1545 VSS.n1354 0.0569562
R72650 VSS.n1542 VSS.n1541 0.0569562
R72651 VSS.n1541 VSS.n1540 0.0569562
R72652 VSS.n1540 VSS.n1539 0.0569562
R72653 VSS.n1539 VSS.n1538 0.0569562
R72654 VSS.n1532 VSS.n1357 0.0569562
R72655 VSS.n2934 VSS.n1149 0.0569562
R72656 VSS.n2930 VSS.n1152 0.0569562
R72657 VSS.n2924 VSS.n2923 0.0569562
R72658 VSS.n2923 VSS.n2922 0.0569562
R72659 VSS.n2922 VSS.n2921 0.0569562
R72660 VSS.n2921 VSS.n2920 0.0569562
R72661 VSS.n2869 VSS.n2868 0.0569562
R72662 VSS.n2868 VSS.n2867 0.0569562
R72663 VSS.n2867 VSS.n2866 0.0569562
R72664 VSS.n2866 VSS.n2865 0.0569562
R72665 VSS.n2865 VSS.n2864 0.0569562
R72666 VSS.n2864 VSS.n2863 0.0569562
R72667 VSS.n2863 VSS.n2862 0.0569562
R72668 VSS.n2862 VSS.n2861 0.0569562
R72669 VSS.n2861 VSS.n2860 0.0569562
R72670 VSS.n3511 VSS.n3510 0.0569562
R72671 VSS.n3512 VSS.n3511 0.0569562
R72672 VSS.n3513 VSS.n3512 0.0569562
R72673 VSS.n3514 VSS.n3513 0.0569562
R72674 VSS.n3515 VSS.n3514 0.0569562
R72675 VSS.n3516 VSS.n3515 0.0569562
R72676 VSS.n3517 VSS.n3516 0.0569562
R72677 VSS.n3518 VSS.n3517 0.0569562
R72678 VSS.n3519 VSS.n3518 0.0569562
R72679 VSS.n3520 VSS.n3519 0.0569562
R72680 VSS.n3521 VSS.n3520 0.0569562
R72681 VSS.n3522 VSS.n3521 0.0569562
R72682 VSS.n3523 VSS.n3522 0.0569562
R72683 VSS.n3524 VSS.n3523 0.0569562
R72684 VSS.n3525 VSS.n3524 0.0569562
R72685 VSS.n3526 VSS.n3525 0.0569562
R72686 VSS.n3527 VSS.n3526 0.0569562
R72687 VSS.n3528 VSS.n3527 0.0569562
R72688 VSS.n3529 VSS.n3528 0.0569562
R72689 VSS.n3530 VSS.n3529 0.0569562
R72690 VSS.n3531 VSS.n3530 0.0569562
R72691 VSS.n3532 VSS.n3531 0.0569562
R72692 VSS.n663 VSS.n655 0.0569562
R72693 VSS.n663 VSS.n656 0.0569562
R72694 VSS.n662 VSS.n656 0.0569562
R72695 VSS.n662 VSS.n657 0.0569562
R72696 VSS.n661 VSS.n657 0.0569562
R72697 VSS.n661 VSS.n658 0.0569562
R72698 VSS.n659 VSS.n658 0.0569562
R72699 VSS.n3936 VSS.n659 0.0569562
R72700 VSS.n3936 VSS.n3935 0.0569562
R72701 VSS.n6118 VSS.n6117 0.0569562
R72702 VSS.n6117 VSS.n6115 0.0569562
R72703 VSS.n6115 VSS.n6114 0.0569562
R72704 VSS.n6114 VSS.n4271 0.0569562
R72705 VSS.n4282 VSS.n4279 0.0569562
R72706 VSS.n4304 VSS.n4291 0.0569562
R72707 VSS.n4304 VSS.n4283 0.0569562
R72708 VSS.n4299 VSS.n4290 0.0569562
R72709 VSS.n4299 VSS.n4284 0.0569562
R72710 VSS.n4302 VSS.n4289 0.0569562
R72711 VSS.n4302 VSS.n4285 0.0569562
R72712 VSS.n4301 VSS.n4288 0.0569562
R72713 VSS.n4301 VSS.n4286 0.0569562
R72714 VSS.n6105 VSS.n4292 0.0569562
R72715 VSS.n6106 VSS.n4293 0.0569562
R72716 VSS.n5614 VSS.n5298 0.0569562
R72717 VSS.n5615 VSS.n5299 0.0569562
R72718 VSS.n5310 VSS.n5295 0.0569562
R72719 VSS.n5308 VSS.n5293 0.0569562
R72720 VSS.n5292 VSS.n5288 0.0569562
R72721 VSS.n5305 VSS.n5302 0.0569562
R72722 VSS.n5305 VSS.n5291 0.0569562
R72723 VSS.n5621 VSS.n5303 0.0569562
R72724 VSS.n5303 VSS.n5290 0.0569562
R72725 VSS.n5090 VSS.n5081 0.0569562
R72726 VSS.n5776 VSS.n5090 0.0569562
R72727 VSS.n5778 VSS.n5088 0.0569562
R72728 VSS.n5775 VSS.n5088 0.0569562
R72729 VSS.n5779 VSS.n5086 0.0569562
R72730 VSS.n5774 VSS.n5086 0.0569562
R72731 VSS.n5780 VSS.n5084 0.0569562
R72732 VSS.n5773 VSS.n5084 0.0569562
R72733 VSS.n5772 VSS.n5083 0.0569562
R72734 VSS.n6106 VSS.n6105 0.0569562
R72735 VSS.n5615 VSS.n5298 0.0569562
R72736 VSS.n5309 VSS.n5295 0.0569562
R72737 VSS.n5307 VSS.n5293 0.0569562
R72738 VSS.n5773 VSS.n5083 0.0569562
R72739 VSS.n1603 VSS.n1602 0.0569562
R72740 VSS.n1602 VSS.n1601 0.0569562
R72741 VSS.n1601 VSS.n1600 0.0569562
R72742 VSS.n1600 VSS.n1599 0.0569562
R72743 VSS.n1599 VSS.n1598 0.0569562
R72744 VSS.n1598 VSS.n1597 0.0569562
R72745 VSS.n1597 VSS.n1596 0.0569562
R72746 VSS.n1210 VSS.n1201 0.0569562
R72747 VSS.n1210 VSS.n1202 0.0569562
R72748 VSS.n1904 VSS.n1202 0.0569562
R72749 VSS.n1905 VSS.n1904 0.0569562
R72750 VSS.n1204 VSS.n1199 0.0569562
R72751 VSS.n1198 VSS.n1187 0.0569562
R72752 VSS.n1198 VSS.n1188 0.0569562
R72753 VSS.n1197 VSS.n1188 0.0569562
R72754 VSS.n1197 VSS.n1189 0.0569562
R72755 VSS.n1196 VSS.n1189 0.0569562
R72756 VSS.n1196 VSS.n1190 0.0569562
R72757 VSS.n1195 VSS.n1190 0.0569562
R72758 VSS.n1195 VSS.n1191 0.0569562
R72759 VSS.n1191 VSS.n1185 0.0569562
R72760 VSS.n2059 VSS.n2058 0.0569562
R72761 VSS.n2060 VSS.n2059 0.0569562
R72762 VSS.n2061 VSS.n2060 0.0569562
R72763 VSS.n2062 VSS.n2061 0.0569562
R72764 VSS.n2063 VSS.n2062 0.0569562
R72765 VSS.n2064 VSS.n2063 0.0569562
R72766 VSS.n2065 VSS.n2064 0.0569562
R72767 VSS.n2066 VSS.n2065 0.0569562
R72768 VSS.n2067 VSS.n2066 0.0569562
R72769 VSS.n2146 VSS.n2091 0.0569562
R72770 VSS.n2135 VSS.n2091 0.0569562
R72771 VSS.n2135 VSS.n2090 0.0569562
R72772 VSS.n2136 VSS.n2090 0.0569562
R72773 VSS.n2136 VSS.n2089 0.0569562
R72774 VSS.n2137 VSS.n2089 0.0569562
R72775 VSS.n2137 VSS.n2088 0.0569562
R72776 VSS.n2138 VSS.n2088 0.0569562
R72777 VSS.n2138 VSS.n2087 0.0569562
R72778 VSS.n2139 VSS.n2087 0.0569562
R72779 VSS.n2139 VSS.n2086 0.0569562
R72780 VSS.n2140 VSS.n2086 0.0569562
R72781 VSS.n2140 VSS.n2085 0.0569562
R72782 VSS.n2141 VSS.n2085 0.0569562
R72783 VSS.n2141 VSS.n2084 0.0569562
R72784 VSS.n2142 VSS.n2084 0.0569562
R72785 VSS.n2142 VSS.n2083 0.0569562
R72786 VSS.n2143 VSS.n2083 0.0569562
R72787 VSS.n2143 VSS.n2082 0.0569562
R72788 VSS.n2144 VSS.n2082 0.0569562
R72789 VSS.n2144 VSS.n2081 0.0569562
R72790 VSS.n2081 VSS.n2078 0.0569562
R72791 VSS.n2214 VSS.n2213 0.0569562
R72792 VSS.n2213 VSS.n2212 0.0569562
R72793 VSS.n2212 VSS.n2211 0.0569562
R72794 VSS.n2211 VSS.n2210 0.0569562
R72795 VSS.n2210 VSS.n2209 0.0569562
R72796 VSS.n2209 VSS.n2208 0.0569562
R72797 VSS.n2208 VSS.n2207 0.0569562
R72798 VSS.n2207 VSS.n2206 0.0569562
R72799 VSS.n2206 VSS.n2205 0.0569562
R72800 VSS.n4262 VSS.n4258 0.0569562
R72801 VSS.n4262 VSS.n4257 0.0569562
R72802 VSS.n4261 VSS.n4257 0.0569562
R72803 VSS.n4261 VSS.n4253 0.0569562
R72804 VSS.n4328 VSS.n4314 0.0569562
R72805 VSS.n6089 VSS.n4322 0.0569562
R72806 VSS.n4329 VSS.n4322 0.0569562
R72807 VSS.n6088 VSS.n4316 0.0569562
R72808 VSS.n4330 VSS.n4316 0.0569562
R72809 VSS.n6087 VSS.n4320 0.0569562
R72810 VSS.n4331 VSS.n4320 0.0569562
R72811 VSS.n6086 VSS.n4318 0.0569562
R72812 VSS.n4332 VSS.n4318 0.0569562
R72813 VSS.n4326 VSS.n4310 0.0569562
R72814 VSS.n6097 VSS.n6096 0.0569562
R72815 VSS.n5282 VSS.n5271 0.0569562
R72816 VSS.n5283 VSS.n5272 0.0569562
R72817 VSS.n5280 VSS.n5268 0.0569562
R72818 VSS.n5278 VSS.n5266 0.0569562
R72819 VSS.n5276 VSS.n5264 0.0569562
R72820 VSS.n5263 VSS.n5259 0.0569562
R72821 VSS.n5630 VSS.n5263 0.0569562
R72822 VSS.n5628 VSS.n5261 0.0569562
R72823 VSS.n5275 VSS.n5261 0.0569562
R72824 VSS.n5005 VSS.n4992 0.0569562
R72825 VSS.n5005 VSS.n4989 0.0569562
R72826 VSS.n5003 VSS.n4993 0.0569562
R72827 VSS.n5003 VSS.n4988 0.0569562
R72828 VSS.n5001 VSS.n4994 0.0569562
R72829 VSS.n5001 VSS.n4987 0.0569562
R72830 VSS.n4999 VSS.n4995 0.0569562
R72831 VSS.n4999 VSS.n4986 0.0569562
R72832 VSS.n4998 VSS.n4985 0.0569562
R72833 VSS.n6096 VSS.n4326 0.0569562
R72834 VSS.n5282 VSS.n5272 0.0569562
R72835 VSS.n5280 VSS.n5267 0.0569562
R72836 VSS.n5278 VSS.n5265 0.0569562
R72837 VSS.n4998 VSS.n4986 0.0569562
R72838 VSS.n2325 VSS.n2323 0.0568736
R72839 VSS.n2323 VSS.n2321 0.0568736
R72840 VSS.n2321 VSS.n2319 0.0568736
R72841 VSS.n2538 VSS.n2536 0.0568736
R72842 VSS.n2536 VSS.n2534 0.0568736
R72843 VSS.n2945 VSS.n1138 0.0563
R72844 VSS.n2679 VSS.n2678 0.0562609
R72845 VSS.n2678 VSS.n2677 0.0562609
R72846 VSS.n2677 VSS.n2218 0.0562609
R72847 VSS.n2667 VSS.n2218 0.0562609
R72848 VSS.n2667 VSS.n2666 0.0562609
R72849 VSS.n2666 VSS.n2665 0.0562609
R72850 VSS.n2665 VSS.n2560 0.0562609
R72851 VSS.n2655 VSS.n2560 0.0562609
R72852 VSS.n2655 VSS.n2654 0.0562609
R72853 VSS.n2654 VSS.n2653 0.0562609
R72854 VSS.n2653 VSS.n2570 0.0562609
R72855 VSS.n2643 VSS.n2570 0.0562609
R72856 VSS.n2643 VSS.n2642 0.0562609
R72857 VSS.n2642 VSS.n2641 0.0562609
R72858 VSS.n2641 VSS.n2580 0.0562609
R72859 VSS.n2631 VSS.n2580 0.0562609
R72860 VSS.n2631 VSS.n2630 0.0562609
R72861 VSS.n2630 VSS.n2629 0.0562609
R72862 VSS.n2629 VSS.n2590 0.0562609
R72863 VSS.n2590 VSS.n665 0.0562609
R72864 VSS.n3929 VSS.n666 0.0562609
R72865 VSS.n3918 VSS.n666 0.0562609
R72866 VSS.n3918 VSS.n3917 0.0562609
R72867 VSS.n3917 VSS.n3916 0.0562609
R72868 VSS.n3916 VSS.n680 0.0562609
R72869 VSS.n3906 VSS.n680 0.0562609
R72870 VSS.n3906 VSS.n3905 0.0562609
R72871 VSS.n3905 VSS.n3904 0.0562609
R72872 VSS.n3904 VSS.n690 0.0562609
R72873 VSS.n3894 VSS.n690 0.0562609
R72874 VSS.n3894 VSS.n3893 0.0562609
R72875 VSS.n3893 VSS.n3892 0.0562609
R72876 VSS.n3892 VSS.n699 0.0562609
R72877 VSS.n3882 VSS.n699 0.0562609
R72878 VSS.n3882 VSS.n3881 0.0562609
R72879 VSS.n3881 VSS.n3880 0.0562609
R72880 VSS.n3880 VSS.n710 0.0562609
R72881 VSS.n3870 VSS.n710 0.0562609
R72882 VSS.n3870 VSS.n3869 0.0562609
R72883 VSS.n3869 VSS.n3868 0.0562609
R72884 VSS.n3868 VSS.n720 0.0562609
R72885 VSS.n3854 VSS.n746 0.0562609
R72886 VSS.n3854 VSS.n3853 0.0562609
R72887 VSS.n3853 VSS.n3852 0.0562609
R72888 VSS.n3852 VSS.n747 0.0562609
R72889 VSS.n3842 VSS.n747 0.0562609
R72890 VSS.n3842 VSS.n3841 0.0562609
R72891 VSS.n3841 VSS.n3840 0.0562609
R72892 VSS.n3840 VSS.n758 0.0562609
R72893 VSS.n3830 VSS.n758 0.0562609
R72894 VSS.n3830 VSS.n3829 0.0562609
R72895 VSS.n3829 VSS.n3828 0.0562609
R72896 VSS.n3828 VSS.n768 0.0562609
R72897 VSS.n3818 VSS.n768 0.0562609
R72898 VSS.n3818 VSS.n3817 0.0562609
R72899 VSS.n3817 VSS.n3816 0.0562609
R72900 VSS.n3816 VSS.n778 0.0562609
R72901 VSS.n3806 VSS.n778 0.0562609
R72902 VSS.n3806 VSS.n3805 0.0562609
R72903 VSS.n3805 VSS.n3804 0.0562609
R72904 VSS.n3804 VSS.n788 0.0562609
R72905 VSS.n3793 VSS.n788 0.0562609
R72906 VSS.n3791 VSS.n3790 0.0562609
R72907 VSS.n3790 VSS.n798 0.0562609
R72908 VSS.n3780 VSS.n798 0.0562609
R72909 VSS.n3780 VSS.n3779 0.0562609
R72910 VSS.n3779 VSS.n3778 0.0562609
R72911 VSS.n3778 VSS.n809 0.0562609
R72912 VSS.n3768 VSS.n809 0.0562609
R72913 VSS.n3768 VSS.n3767 0.0562609
R72914 VSS.n3767 VSS.n3766 0.0562609
R72915 VSS.n3766 VSS.n819 0.0562609
R72916 VSS.n3756 VSS.n819 0.0562609
R72917 VSS.n3756 VSS.n3755 0.0562609
R72918 VSS.n3755 VSS.n3754 0.0562609
R72919 VSS.n3754 VSS.n829 0.0562609
R72920 VSS.n3744 VSS.n829 0.0562609
R72921 VSS.n3744 VSS.n3743 0.0562609
R72922 VSS.n3743 VSS.n3742 0.0562609
R72923 VSS.n3742 VSS.n839 0.0562609
R72924 VSS.n3732 VSS.n839 0.0562609
R72925 VSS.n3732 VSS.n3731 0.0562609
R72926 VSS.n2683 VSS.n2070 0.0562609
R72927 VSS.n2596 VSS.n2070 0.0562609
R72928 VSS.n2598 VSS.n2596 0.0562609
R72929 VSS.n2599 VSS.n2598 0.0562609
R72930 VSS.n2601 VSS.n2599 0.0562609
R72931 VSS.n2602 VSS.n2601 0.0562609
R72932 VSS.n2604 VSS.n2602 0.0562609
R72933 VSS.n2605 VSS.n2604 0.0562609
R72934 VSS.n2607 VSS.n2605 0.0562609
R72935 VSS.n2608 VSS.n2607 0.0562609
R72936 VSS.n2610 VSS.n2608 0.0562609
R72937 VSS.n2611 VSS.n2610 0.0562609
R72938 VSS.n2613 VSS.n2611 0.0562609
R72939 VSS.n2614 VSS.n2613 0.0562609
R72940 VSS.n2616 VSS.n2614 0.0562609
R72941 VSS.n2617 VSS.n2616 0.0562609
R72942 VSS.n2618 VSS.n2617 0.0562609
R72943 VSS.n2620 VSS.n2618 0.0562609
R72944 VSS.n2620 VSS.n2619 0.0562609
R72945 VSS.n2619 VSS.n969 0.0562609
R72946 VSS.n3505 VSS.n3504 0.0562609
R72947 VSS.n3504 VSS.n3502 0.0562609
R72948 VSS.n3502 VSS.n3501 0.0562609
R72949 VSS.n3501 VSS.n3499 0.0562609
R72950 VSS.n3499 VSS.n3498 0.0562609
R72951 VSS.n3498 VSS.n3496 0.0562609
R72952 VSS.n3496 VSS.n3495 0.0562609
R72953 VSS.n3495 VSS.n3493 0.0562609
R72954 VSS.n3493 VSS.n3492 0.0562609
R72955 VSS.n3492 VSS.n3490 0.0562609
R72956 VSS.n3490 VSS.n3489 0.0562609
R72957 VSS.n3489 VSS.n3487 0.0562609
R72958 VSS.n3487 VSS.n3486 0.0562609
R72959 VSS.n3486 VSS.n3484 0.0562609
R72960 VSS.n3484 VSS.n3483 0.0562609
R72961 VSS.n3483 VSS.n3481 0.0562609
R72962 VSS.n3481 VSS.n3480 0.0562609
R72963 VSS.n3480 VSS.n3478 0.0562609
R72964 VSS.n3478 VSS.n3477 0.0562609
R72965 VSS.n3477 VSS.n3475 0.0562609
R72966 VSS.n3475 VSS.n3474 0.0562609
R72967 VSS.n3471 VSS.n3470 0.0562609
R72968 VSS.n3470 VSS.n3469 0.0562609
R72969 VSS.n3469 VSS.n3467 0.0562609
R72970 VSS.n3467 VSS.n3466 0.0562609
R72971 VSS.n3466 VSS.n3464 0.0562609
R72972 VSS.n3464 VSS.n3463 0.0562609
R72973 VSS.n3463 VSS.n3461 0.0562609
R72974 VSS.n3461 VSS.n3460 0.0562609
R72975 VSS.n3460 VSS.n3458 0.0562609
R72976 VSS.n3458 VSS.n3457 0.0562609
R72977 VSS.n3457 VSS.n3455 0.0562609
R72978 VSS.n3455 VSS.n3454 0.0562609
R72979 VSS.n3454 VSS.n3452 0.0562609
R72980 VSS.n3452 VSS.n3451 0.0562609
R72981 VSS.n3451 VSS.n3449 0.0562609
R72982 VSS.n3449 VSS.n3448 0.0562609
R72983 VSS.n3448 VSS.n3446 0.0562609
R72984 VSS.n3446 VSS.n3445 0.0562609
R72985 VSS.n3445 VSS.n3443 0.0562609
R72986 VSS.n3443 VSS.n3442 0.0562609
R72987 VSS.n3442 VSS.n3440 0.0562609
R72988 VSS.n3069 VSS.n972 0.0562609
R72989 VSS.n3071 VSS.n3069 0.0562609
R72990 VSS.n3072 VSS.n3071 0.0562609
R72991 VSS.n3074 VSS.n3072 0.0562609
R72992 VSS.n3075 VSS.n3074 0.0562609
R72993 VSS.n3077 VSS.n3075 0.0562609
R72994 VSS.n3078 VSS.n3077 0.0562609
R72995 VSS.n3080 VSS.n3078 0.0562609
R72996 VSS.n3081 VSS.n3080 0.0562609
R72997 VSS.n3083 VSS.n3081 0.0562609
R72998 VSS.n3084 VSS.n3083 0.0562609
R72999 VSS.n3086 VSS.n3084 0.0562609
R73000 VSS.n3087 VSS.n3086 0.0562609
R73001 VSS.n3089 VSS.n3087 0.0562609
R73002 VSS.n3090 VSS.n3089 0.0562609
R73003 VSS.n3092 VSS.n3090 0.0562609
R73004 VSS.n3093 VSS.n3092 0.0562609
R73005 VSS.n3095 VSS.n3093 0.0562609
R73006 VSS.n3096 VSS.n3095 0.0562609
R73007 VSS.n3097 VSS.n3096 0.0562609
R73008 VSS.n1884 DVSS 0.0560627
R73009 DVSS VSS.n1211 0.0560627
R73010 VSS.n5987 VSS.n5986 0.0554
R73011 VSS.n5521 VSS.n4961 0.0554
R73012 VSS.n5991 VSS.n5990 0.0554
R73013 VSS.n5522 VSS.n5191 0.0554
R73014 VSS.n6102 VSS.n4295 0.0554
R73015 VSS.n5624 VSS.n5623 0.0554
R73016 VSS.n6100 VSS.n6099 0.0554
R73017 VSS.n5627 VSS.n5626 0.0554
R73018 VSS.n143 VSS.n125 0.055378
R73019 VSS.n6458 VSS.n7 0.055378
R73020 VSS.n4181 VSS.n4178 0.0540178
R73021 VSS.n6151 VSS.n6150 0.0540178
R73022 VSS.n6147 VSS.n479 0.0540178
R73023 VSS.n5489 VSS.n5481 0.0540178
R73024 VSS.n6142 VSS.n488 0.0536
R73025 VSS.n5255 VSS.n4975 0.0536
R73026 VSS.n5078 VSS.n5077 0.0536
R73027 VSS.n6145 VSS.n485 0.0536
R73028 VSS.n5640 VSS.n5639 0.0536
R73029 VSS.n5793 VSS.n5792 0.0536
R73030 VSS.n6124 VSS.n4267 0.0536
R73031 VSS.n5616 VSS.n5257 0.0536
R73032 VSS.n5786 VSS.n5080 0.0536
R73033 VSS.n4259 VSS.n4252 0.0536
R73034 VSS.n5634 VSS.n5258 0.0536
R73035 VSS.n5787 VSS.n4991 0.0536
R73036 VSS.n6173 VSS.n471 0.0533261
R73037 VSS.n4182 VSS.n4180 0.0533261
R73038 VSS.n4188 VSS.n4180 0.0533261
R73039 VSS.n4187 VSS.n4184 0.0533261
R73040 VSS.n4196 VSS.n537 0.0533261
R73041 VSS.n5494 VSS.n5490 0.0533261
R73042 VSS.n5499 VSS.n5495 0.0533261
R73043 VSS.n5483 VSS.n5482 0.0533261
R73044 VSS.n5502 VSS.n5483 0.0533261
R73045 VSS.n5488 VSS.n5487 0.0533261
R73046 VSS.n5861 VSS.n4946 0.0533261
R73047 VSS.n1121 VSS.n1092 0.0527
R73048 VSS.n2963 VSS.n1083 0.0527
R73049 VSS.n1158 VSS.n1156 0.0527
R73050 VSS.n2926 VSS.n1159 0.0527
R73051 VSS.n1881 VSS.n1234 0.05225
R73052 VSS.n1745 VSS.n1744 0.05225
R73053 VSS.n1616 VSS.n1615 0.05225
R73054 VSS.n1605 VSS.n1547 0.05225
R73055 VSS.n6230 VSS.n6229 0.0521279
R73056 VSS.n133 VSS.n18 0.0521279
R73057 VSS.n1885 VSS.n1232 0.0518
R73058 VSS.n4820 VSS.n4808 0.0518
R73059 VSS.n5514 VSS.n4960 0.0518
R73060 VSS.n1889 VSS.n1228 0.0518
R73061 VSS.n4812 VSS.n4811 0.0518
R73062 VSS.n5515 VSS.n5190 0.0518
R73063 VSS.n1895 VSS.n1216 0.0518
R73064 VSS.n4814 VSS.n4300 0.0518
R73065 VSS.n5510 VSS.n5301 0.0518
R73066 VSS.n1902 VSS.n1901 0.0518
R73067 VSS.n4815 VSS.n4317 0.0518
R73068 VSS.n5511 VSS.n5285 0.0518
R73069 VSS.n2938 VSS.n1146 0.0507703
R73070 VSS.n2942 VSS.n1141 0.0507703
R73071 VSS.n4976 VSS.n4964 0.05
R73072 VSS.n5095 VSS.n4929 0.05
R73073 VSS.n5641 VSS.n5194 0.05
R73074 VSS.n5096 VSS.n5066 0.05
R73075 VSS.n5617 VSS.n5304 0.05
R73076 VSS.n5104 VSS.n5103 0.05
R73077 VSS.n5631 VSS.n5273 0.05
R73078 VSS.n5101 VSS.n5008 0.05
R73079 VSS.n4098 VSS.n4097 0.049839
R73080 VSS.n4092 VSS.n4091 0.049839
R73081 VSS.n6189 VSS.n6188 0.049839
R73082 VSS.n6158 VSS.n473 0.049839
R73083 VSS.n6176 VSS.n469 0.0491
R73084 VSS.n6236 VSS.n6235 0.0490001
R73085 VSS.n3690 DVSS 0.0487259
R73086 DVSS VSS.n5962 0.0487259
R73087 VSS.n4832 VSS.n4806 0.0482
R73088 VSS.n5532 VSS.n4959 0.0482
R73089 VSS.n4824 VSS.n4823 0.0482
R73090 VSS.n5533 VSS.n5189 0.0482
R73091 VSS.n4826 VSS.n4303 0.0482
R73092 VSS.n5528 VSS.n5300 0.0482
R73093 VSS.n4827 VSS.n4321 0.0482
R73094 VSS.n5529 VSS.n5284 0.0482
R73095 VSS.n4777 VSS.n4776 0.0481866
R73096 VSS.n5886 DVSS 0.0480659
R73097 VSS.n2534 VSS.n2532 0.0479692
R73098 VSS.n6140 VSS.n490 0.0464
R73099 VSS.n5851 VSS.n5850 0.0464
R73100 VSS.n5106 VSS.n4930 0.0464
R73101 VSS.n4763 VSS.n486 0.0464
R73102 VSS.n5642 VSS.n4977 0.0464
R73103 VSS.n5107 VSS.n5067 0.0464
R73104 VSS.n6122 VSS.n4269 0.0464
R73105 VSS.n5618 VSS.n4979 0.0464
R73106 VSS.n5115 VSS.n5114 0.0464
R73107 VSS.n6128 VSS.n6127 0.0464
R73108 VSS.n5844 VSS.n4980 0.0464
R73109 VSS.n5112 VSS.n5009 0.0464
R73110 VSS.n4182 VSS.n476 0.0457174
R73111 VSS.n6153 VSS.n6152 0.0457174
R73112 VSS.n5482 VSS.n478 0.0457174
R73113 VSS.n5867 VSS.n5866 0.0456261
R73114 VSS.n5803 VSS.n5802 0.0456261
R73115 VSS.n5783 VSS.n5782 0.0456261
R73116 VSS.n4997 VSS.n4983 0.0456261
R73117 VSS.n6216 VSS.n6215 0.0449833
R73118 VSS.n1254 VSS.n1231 0.0446
R73119 VSS.n4844 VSS.n4804 0.0446
R73120 VSS.n1279 VSS.n1227 0.0446
R73121 VSS.n4836 VSS.n4835 0.0446
R73122 VSS.n1534 VSS.n1215 0.0446
R73123 VSS.n4838 VSS.n4298 0.0446
R73124 VSS.n1898 VSS.n1203 0.0446
R73125 VSS.n4839 VSS.n4315 0.0446
R73126 VSS.n17 VSS.n14 0.04343
R73127 VSS.n6207 VSS.n6205 0.04343
R73128 VSS.n6209 VSS.n6208 0.04343
R73129 VSS.n6206 VSS.n6203 0.04343
R73130 VSS.n6213 VSS.n6204 0.04343
R73131 VSS.n128 VSS.n127 0.04343
R73132 VSS.n130 VSS.n129 0.04343
R73133 VSS.n6450 VSS.n6449 0.04343
R73134 VSS.n3930 VSS.n3929 0.0430543
R73135 VSS.n3793 VSS.n3792 0.0430543
R73136 VSS.n3506 VSS.n3505 0.0430543
R73137 VSS.n3440 VSS.n3439 0.0430543
R73138 VSS.n5051 VSS.n4931 0.0428
R73139 VSS.n5806 VSS.n5052 0.0428
R73140 VSS.n5119 VSS.n5118 0.0428
R73141 VSS.n5116 VSS.n5010 0.0428
R73142 VSS.n2327 VSS.n2325 0.0424895
R73143 VSS.n5034 VSS.n4978 0.041806
R73144 VSS.n4856 VSS.n4802 0.041
R73145 VSS.n4848 VSS.n4847 0.041
R73146 VSS.n4850 VSS.n4305 0.041
R73147 VSS.n4851 VSS.n4323 0.041
R73148 VSS.n137 VSS.n136 0.04037
R73149 VSS.n19 VSS.n16 0.04037
R73150 VSS.n5863 VSS.n4932 0.0401
R73151 VSS.n5799 VSS.n5068 0.0401
R73152 VSS.n5834 VSS.n5014 0.0401
R73153 VSS.n5839 VSS.n5838 0.0401
R73154 VSS.n2319 VSS.n2317 0.0395659
R73155 VSS.n2539 VSS.n2538 0.0395659
R73156 VSS.n6214 VSS.n6213 0.0389615
R73157 VSS.n6450 VSS.n14 0.0389615
R73158 VSS.n6205 VSS.n14 0.0389615
R73159 VSS.n6209 VSS.n6205 0.0389615
R73160 VSS.n6209 VSS.n6203 0.0389615
R73161 VSS.n6213 VSS.n6203 0.0389615
R73162 VSS.n6229 VSS.n6228 0.0389615
R73163 VSS.n129 VSS.n128 0.0389615
R73164 VSS.n137 VSS.n129 0.0389615
R73165 VSS.n137 VSS.n16 0.0389615
R73166 VSS.n6450 VSS.n16 0.0389615
R73167 VSS.n4116 VSS.n4115 0.03875
R73168 VSS.n3933 VSS.n3932 0.03875
R73169 VSS.n1255 VSS.n1229 0.0374
R73170 VSS.n1280 VSS.n1225 0.0374
R73171 VSS.n1535 VSS.n1213 0.0374
R73172 VSS.n1212 VSS.n1206 0.0374
R73173 VSS.n2985 VSS.n1093 0.03695
R73174 VSS.n2984 VSS.n1095 0.03695
R73175 VSS.n2918 VSS.n2917 0.03695
R73176 VSS.n2916 VSS.n2873 0.03695
R73177 VSS.n4513 VSS.n497 0.0365
R73178 VSS.n4770 VSS.n4769 0.0365
R73179 VSS.n4508 VSS.n4272 0.0365
R73180 VSS.n4510 VSS.n4254 0.0365
R73181 VSS.n2145 VSS.n2134 0.0362074
R73182 VSS.n4791 VSS.n4407 0.0350896
R73183 DVSS VSS.n1883 0.0338686
R73184 VSS.n1607 DVSS 0.0338686
R73185 VSS.n6458 VSS.n6457 0.0337188
R73186 VSS.n143 VSS.n142 0.0337188
R73187 VSS.n5379 VSS.n5378 0.0336863
R73188 VSS.n5387 VSS.n5386 0.0336863
R73189 VSS.n5385 VSS.n5384 0.0332409
R73190 VSS.n4945 VSS.n4918 0.0329
R73191 VSS.n5798 VSS.n5055 0.0329
R73192 VSS.n5015 VSS.n5012 0.0329
R73193 VSS.n4996 VSS.n4984 0.0329
R73194 VSS.n444 VSS.n6 0.0329
R73195 VSS.n441 VSS.n440 0.0329
R73196 VSS.n2679 VSS.n2217 0.0313152
R73197 VSS.n3731 VSS.n3730 0.0313152
R73198 VSS.n2684 VSS.n2683 0.0313152
R73199 VSS.n3400 VSS.n3097 0.0313152
R73200 VSS.n5860 VSS.n5858 0.0311
R73201 VSS.n5486 VSS.n4454 0.0311
R73202 VSS.n5498 VSS.n4281 0.0311
R73203 VSS.n5491 VSS.n4327 0.0311
R73204 VSS.n5384 VSS.n5383 0.0309017
R73205 VSS.n5378 VSS.n5377 0.0304416
R73206 VSS.n5387 VSS.n5328 0.0304416
R73207 VSS.n2931 VSS.n1153 0.0301809
R73208 VSS.n2954 VSS.n1134 0.0301809
R73209 VSS.n2935 VSS.n1150 0.0301809
R73210 VSS.n2948 VSS.n1137 0.0301809
R73211 VSS.n2134 VSS.n2092 0.0301532
R73212 VSS.n1126 VSS.n1125 0.0293889
R73213 VSS.n1127 VSS.n1126 0.0293889
R73214 VSS.n2881 VSS.n1127 0.0293889
R73215 VSS.n2881 VSS.n2880 0.0293889
R73216 VSS.n5504 VSS.n5503 0.0293806
R73217 VSS.n1880 VSS.n1235 0.0287281
R73218 VSS.n1835 VSS.n1240 0.0287281
R73219 VSS.n1834 VSS.n1249 0.0287281
R73220 VSS.n1826 VSS.n1251 0.0287281
R73221 VSS.n1827 VSS.n1232 0.0287281
R73222 VSS.n1829 VSS.n1253 0.0287281
R73223 VSS.n1828 VSS.n1051 0.0287281
R73224 VSS.n3065 VSS.n1049 0.0287281
R73225 VSS.n3066 VSS.n998 0.0287281
R73226 VSS.n3402 VSS.n3068 0.0287281
R73227 VSS.n3725 VSS.n3724 0.0287281
R73228 VSS.n3728 VSS.n576 0.0287281
R73229 VSS.n4090 VSS.n574 0.0287281
R73230 VSS.n6138 VSS.n6137 0.0287281
R73231 VSS.n493 VSS.n492 0.0287281
R73232 VSS.n502 VSS.n501 0.0287281
R73233 VSS.n499 VSS.n497 0.0287281
R73234 VSS.n4857 VSS.n4481 0.0287281
R73235 VSS.n4802 VSS.n4797 0.0287281
R73236 VSS.n4845 VSS.n4480 0.0287281
R73237 VSS.n4804 VSS.n4798 0.0287281
R73238 VSS.n4833 VSS.n4479 0.0287281
R73239 VSS.n4806 VSS.n4799 0.0287281
R73240 VSS.n4821 VSS.n4478 0.0287281
R73241 VSS.n4808 VSS.n4800 0.0287281
R73242 VSS.n4475 VSS.n4472 0.0287281
R73243 VSS.n5858 VSS.n4476 0.0287281
R73244 VSS.n4970 VSS.n4954 0.0287281
R73245 VSS.n4968 VSS.n4952 0.0287281
R73246 VSS.n5077 VSS.n4928 0.0287281
R73247 VSS.n4801 VSS.n4796 0.0287281
R73248 VSS.n500 VSS.n499 0.0287281
R73249 VSS.n6137 VSS.n488 0.0287281
R73250 VSS.n3727 VSS.n850 0.0287281
R73251 VSS.n5986 VSS.n4473 0.0287281
R73252 VSS.n5856 VSS.n4947 0.0287281
R73253 VSS.n4972 VSS.n4958 0.0287281
R73254 VSS.n4971 VSS.n4959 0.0287281
R73255 VSS.n4969 VSS.n4960 0.0287281
R73256 VSS.n4967 VSS.n4961 0.0287281
R73257 VSS.n4975 VSS.n4951 0.0287281
R73258 VSS.n4966 VSS.n4962 0.0287281
R73259 VSS.n4976 VSS.n4950 0.0287281
R73260 VSS.n5854 VSS.n5853 0.0287281
R73261 VSS.n5851 VSS.n4949 0.0287281
R73262 VSS.n5849 VSS.n4928 0.0287281
R73263 VSS.n4939 VSS.n4927 0.0287281
R73264 VSS.n4938 VSS.n4929 0.0287281
R73265 VSS.n4940 VSS.n4925 0.0287281
R73266 VSS.n4937 VSS.n4930 0.0287281
R73267 VSS.n4941 VSS.n4923 0.0287281
R73268 VSS.n4936 VSS.n4931 0.0287281
R73269 VSS.n4942 VSS.n4921 0.0287281
R73270 VSS.n4934 VSS.n4932 0.0287281
R73271 VSS.n1747 VSS.n1283 0.0287281
R73272 VSS.n1750 VSS.n1278 0.0287281
R73273 VSS.n2777 VSS.n1085 0.0287281
R73274 VSS.n3437 VSS.n973 0.0287281
R73275 VSS.n3636 VSS.n882 0.0287281
R73276 VSS.n4105 VSS.n4104 0.0287281
R73277 VSS.n4766 VSS.n485 0.0287281
R73278 VSS.n4519 VSS.n4515 0.0287281
R73279 VSS.n5200 VSS.n5183 0.0287281
R73280 VSS.n5198 VSS.n5181 0.0287281
R73281 VSS.n5793 VSS.n5065 0.0287281
R73282 VSS.n2952 VSS.n2950 0.0287281
R73283 VSS.n2947 VSS.n2946 0.0287281
R73284 VSS.n2949 VSS.n1135 0.0287281
R73285 VSS.n2953 VSS.n2951 0.0287281
R73286 VSS.n4811 VSS.n4462 0.0287281
R73287 VSS.n4810 VSS.n4458 0.0287281
R73288 VSS.n4823 VSS.n4464 0.0287281
R73289 VSS.n4822 VSS.n4457 0.0287281
R73290 VSS.n4835 VSS.n4466 0.0287281
R73291 VSS.n4834 VSS.n4456 0.0287281
R73292 VSS.n4847 VSS.n4468 0.0287281
R73293 VSS.n4846 VSS.n4455 0.0287281
R73294 VSS.n4470 VSS.n4469 0.0287281
R73295 VSS.n4769 VSS.n4515 0.0287281
R73296 VSS.n4517 VSS.n4514 0.0287281
R73297 VSS.n4764 VSS.n4521 0.0287281
R73298 VSS.n4767 VSS.n4766 0.0287281
R73299 VSS.n4115 VSS.n4114 0.0287281
R73300 VSS.n2778 VSS.n975 0.0287281
R73301 VSS.n1095 VSS.n1085 0.0287281
R73302 VSS.n1086 VSS.n1082 0.0287281
R73303 VSS.n1091 VSS.n1090 0.0287281
R73304 VSS.n1277 VSS.n1228 0.0287281
R73305 VSS.n1753 VSS.n1281 0.0287281
R73306 VSS.n1748 VSS.n1275 0.0287281
R73307 VSS.n1743 VSS.n1289 0.0287281
R73308 VSS.n3639 VSS.n3638 0.0287281
R73309 VSS.n5992 VSS.n5991 0.0287281
R73310 VSS.n5993 VSS.n4454 0.0287281
R73311 VSS.n5253 VSS.n5185 0.0287281
R73312 VSS.n5202 VSS.n5188 0.0287281
R73313 VSS.n5201 VSS.n5189 0.0287281
R73314 VSS.n5199 VSS.n5190 0.0287281
R73315 VSS.n5197 VSS.n5191 0.0287281
R73316 VSS.n5640 VSS.n5180 0.0287281
R73317 VSS.n5196 VSS.n5192 0.0287281
R73318 VSS.n5641 VSS.n5179 0.0287281
R73319 VSS.n5645 VSS.n5644 0.0287281
R73320 VSS.n5642 VSS.n5178 0.0287281
R73321 VSS.n5076 VSS.n5065 0.0287281
R73322 VSS.n5794 VSS.n5063 0.0287281
R73323 VSS.n5075 VSS.n5066 0.0287281
R73324 VSS.n5795 VSS.n5061 0.0287281
R73325 VSS.n5074 VSS.n5067 0.0287281
R73326 VSS.n5796 VSS.n5059 0.0287281
R73327 VSS.n5073 VSS.n5052 0.0287281
R73328 VSS.n5805 VSS.n5053 0.0287281
R73329 VSS.n5071 VSS.n5068 0.0287281
R73330 VSS.n4471 VSS.n4459 0.0287281
R73331 VSS.n1545 VSS.n1544 0.0287281
R73332 VSS.n1533 VSS.n1532 0.0287281
R73333 VSS.n2937 VSS.n1148 0.0287281
R73334 VSS.n2872 VSS.n2871 0.0287281
R73335 VSS.n2860 VSS.n968 0.0287281
R73336 VSS.n3532 VSS.n664 0.0287281
R73337 VSS.n3935 VSS.n456 0.0287281
R73338 VSS.n6119 VSS.n4267 0.0287281
R73339 VSS.n6113 VSS.n4274 0.0287281
R73340 VSS.n5309 VSS.n5294 0.0287281
R73341 VSS.n5307 VSS.n5287 0.0287281
R73342 VSS.n5092 VSS.n5080 0.0287281
R73343 VSS.n1148 VSS.n1147 0.0287281
R73344 VSS.n2932 VSS.n1152 0.0287281
R73345 VSS.n2936 VSS.n1149 0.0287281
R73346 VSS.n2934 VSS.n2933 0.0287281
R73347 VSS.n2930 VSS.n2929 0.0287281
R73348 VSS.n4300 VSS.n4288 0.0287281
R73349 VSS.n4307 VSS.n4285 0.0287281
R73350 VSS.n4303 VSS.n4289 0.0287281
R73351 VSS.n4296 VSS.n4284 0.0287281
R73352 VSS.n4298 VSS.n4290 0.0287281
R73353 VSS.n4306 VSS.n4283 0.0287281
R73354 VSS.n4305 VSS.n4291 0.0287281
R73355 VSS.n4297 VSS.n4282 0.0287281
R73356 VSS.n6108 VSS.n4279 0.0287281
R73357 VSS.n4274 VSS.n4272 0.0287281
R73358 VSS.n4507 VSS.n4271 0.0287281
R73359 VSS.n6118 VSS.n6116 0.0287281
R73360 VSS.n6120 VSS.n6119 0.0287281
R73361 VSS.n3933 VSS.n655 0.0287281
R73362 VSS.n2870 VSS.n2869 0.0287281
R73363 VSS.n2873 VSS.n2872 0.0287281
R73364 VSS.n2920 VSS.n2919 0.0287281
R73365 VSS.n2925 VSS.n2924 0.0287281
R73366 VSS.n1357 VSS.n1216 0.0287281
R73367 VSS.n1538 VSS.n1537 0.0287281
R73368 VSS.n1543 VSS.n1542 0.0287281
R73369 VSS.n1348 VSS.n1347 0.0287281
R73370 VSS.n3510 VSS.n3509 0.0287281
R73371 VSS.n4295 VSS.n4292 0.0287281
R73372 VSS.n4293 VSS.n4281 0.0287281
R73373 VSS.n5614 VSS.n5296 0.0287281
R73374 VSS.n5311 VSS.n5299 0.0287281
R73375 VSS.n5310 VSS.n5300 0.0287281
R73376 VSS.n5308 VSS.n5301 0.0287281
R73377 VSS.n5623 VSS.n5288 0.0287281
R73378 VSS.n5616 VSS.n5292 0.0287281
R73379 VSS.n5306 VSS.n5302 0.0287281
R73380 VSS.n5617 VSS.n5291 0.0287281
R73381 VSS.n5621 VSS.n5620 0.0287281
R73382 VSS.n5618 VSS.n5290 0.0287281
R73383 VSS.n5777 VSS.n5092 0.0287281
R73384 VSS.n5785 VSS.n5081 0.0287281
R73385 VSS.n5776 VSS.n5104 0.0287281
R73386 VSS.n5778 VSS.n5089 0.0287281
R73387 VSS.n5775 VSS.n5115 0.0287281
R73388 VSS.n5779 VSS.n5087 0.0287281
R73389 VSS.n5774 VSS.n5119 0.0287281
R73390 VSS.n5780 VSS.n5085 0.0287281
R73391 VSS.n5772 VSS.n5014 0.0287281
R73392 VSS.n6103 VSS.n4286 0.0287281
R73393 VSS.n1596 VSS.n1595 0.0287281
R73394 VSS.n1907 VSS.n1199 0.0287281
R73395 VSS.n2056 VSS.n1185 0.0287281
R73396 VSS.n2686 VSS.n2067 0.0287281
R73397 VSS.n2149 VSS.n2078 0.0287281
R73398 VSS.n2205 VSS.n2204 0.0287281
R73399 VSS.n4252 VSS.n4250 0.0287281
R73400 VSS.n4260 VSS.n4256 0.0287281
R73401 VSS.n5279 VSS.n5267 0.0287281
R73402 VSS.n5277 VSS.n5265 0.0287281
R73403 VSS.n4991 VSS.n4981 0.0287281
R73404 VSS.n6086 VSS.n4317 0.0287281
R73405 VSS.n4331 VSS.n4325 0.0287281
R73406 VSS.n6087 VSS.n4321 0.0287281
R73407 VSS.n4330 VSS.n4312 0.0287281
R73408 VSS.n6088 VSS.n4315 0.0287281
R73409 VSS.n4329 VSS.n4324 0.0287281
R73410 VSS.n6089 VSS.n4323 0.0287281
R73411 VSS.n4328 VSS.n4313 0.0287281
R73412 VSS.n6094 VSS.n4314 0.0287281
R73413 VSS.n4260 VSS.n4254 0.0287281
R73414 VSS.n4509 VSS.n4253 0.0287281
R73415 VSS.n4264 VSS.n4258 0.0287281
R73416 VSS.n6130 VSS.n4250 0.0287281
R73417 VSS.n2215 VSS.n2214 0.0287281
R73418 VSS.n2058 VSS.n2057 0.0287281
R73419 VSS.n1908 VSS.n1187 0.0287281
R73420 VSS.n1902 VSS.n1204 0.0287281
R73421 VSS.n1905 VSS.n1207 0.0287281
R73422 VSS.n1209 VSS.n1201 0.0287281
R73423 VSS.n1604 VSS.n1603 0.0287281
R73424 VSS.n2147 VSS.n2146 0.0287281
R73425 VSS.n6099 VSS.n4310 0.0287281
R73426 VSS.n6097 VSS.n4327 0.0287281
R73427 VSS.n5281 VSS.n5271 0.0287281
R73428 VSS.n5283 VSS.n5269 0.0287281
R73429 VSS.n5284 VSS.n5268 0.0287281
R73430 VSS.n5285 VSS.n5266 0.0287281
R73431 VSS.n5627 VSS.n5264 0.0287281
R73432 VSS.n5276 VSS.n5258 0.0287281
R73433 VSS.n5633 VSS.n5259 0.0287281
R73434 VSS.n5631 VSS.n5630 0.0287281
R73435 VSS.n5628 VSS.n5262 0.0287281
R73436 VSS.n5275 VSS.n4980 0.0287281
R73437 VSS.n5843 VSS.n4981 0.0287281
R73438 VSS.n5006 VSS.n4992 0.0287281
R73439 VSS.n5008 VSS.n4989 0.0287281
R73440 VSS.n5004 VSS.n4993 0.0287281
R73441 VSS.n5009 VSS.n4988 0.0287281
R73442 VSS.n5002 VSS.n4994 0.0287281
R73443 VSS.n5010 VSS.n4987 0.0287281
R73444 VSS.n5000 VSS.n4995 0.0287281
R73445 VSS.n5839 VSS.n4985 0.0287281
R73446 VSS.n4332 VSS.n4309 0.0287281
R73447 VSS.n1552 VSS.n1551 0.0287254
R73448 VSS.n2317 VSS.n2313 0.0283804
R73449 VSS.n2317 VSS.n2316 0.0283804
R73450 VSS.n922 VSS.n720 0.0283804
R73451 VSS.n922 VSS.n746 0.0283804
R73452 VSS.n3394 VSS.n3393 0.0283804
R73453 VSS.n2539 VSS.n2444 0.0283804
R73454 VSS.n2541 VSS.n2539 0.0283804
R73455 VSS.n3474 VSS.n970 0.0283804
R73456 VSS.n3471 VSS.n970 0.0283804
R73457 VSS.n3131 VSS.n3098 0.0283804
R73458 VSS.n6175 VSS.n470 0.0272589
R73459 VSS.n6175 VSS.n6174 0.0272589
R73460 VSS.n6126 VSS.n4265 0.0272589
R73461 VSS.n6123 VSS.n4266 0.0272589
R73462 VSS.n6146 VSS.n484 0.0272589
R73463 VSS.n6143 VSS.n487 0.0272589
R73464 VSS.n6125 VSS.n4266 0.0272589
R73465 VSS.n6144 VSS.n484 0.0272589
R73466 VSS.n6141 VSS.n487 0.0272589
R73467 VSS.n4265 VSS.n474 0.0272589
R73468 VSS.n5500 VSS.n5481 0.0272589
R73469 VSS.n6150 VSS.n481 0.0272589
R73470 VSS.n6152 VSS.n479 0.0272589
R73471 VSS.n4181 VSS.n4179 0.0272589
R73472 VSS.n4182 VSS.n4178 0.0272589
R73473 VSS.n6152 VSS.n6151 0.0272589
R73474 VSS.n6148 VSS.n6147 0.0272589
R73475 VSS.n5489 VSS.n5482 0.0272589
R73476 VSS.n6159 VSS.n6156 0.026913
R73477 VSS.n458 VSS.n457 0.026913
R73478 VSS.n4128 VSS.n555 0.026913
R73479 VSS.n4133 VSS.n556 0.026913
R73480 VSS.n4094 VSS.n558 0.026913
R73481 VSS.n4096 VSS.n4095 0.026913
R73482 VSS.n1375 VSS.n1208 0.0262332
R73483 VSS.n1910 VSS.n1193 0.0262332
R73484 VSS.n2690 VSS.n2689 0.0262332
R73485 VSS.n2155 VSS.n2153 0.0262332
R73486 VSS.n4571 VSS.n4570 0.0262332
R73487 VSS.n2915 VSS.n1162 0.0259955
R73488 VSS.n2979 VSS.n2978 0.0259955
R73489 VSS.n1100 VSS.n1096 0.0259955
R73490 VSS.n2983 VSS.n2982 0.0259955
R73491 VSS.n2940 VSS.n2939 0.0259955
R73492 VSS.n2944 VSS.n1140 0.0259955
R73493 VSS.n2982 VSS.n1094 0.0259955
R73494 VSS.n2944 VSS.n2943 0.0259955
R73495 VSS.n1162 VSS.n1101 0.0259955
R73496 VSS.n2939 VSS.n1144 0.0259955
R73497 VSS.n2978 VSS.n1098 0.0259955
R73498 VSS.n2981 VSS.n1096 0.0259955
R73499 VSS.n5866 VSS.n4933 0.0257
R73500 VSS.n5802 VSS.n5069 0.0257
R73501 VSS.n5782 VSS.n5120 0.0257
R73502 VSS.n5841 VSS.n4997 0.0257
R73503 VSS.n1125 VSS.n1098 0.0256351
R73504 VSS.n1125 VSS.n1100 0.0256351
R73505 VSS.n2880 VSS.n1144 0.0256351
R73506 VSS.n2880 VSS.n1141 0.0256351
R73507 VSS.n2314 VSS.n2217 0.0254457
R73508 VSS.n3730 VSS.n849 0.0254457
R73509 VSS.n2684 VSS.n2069 0.0254457
R73510 VSS.n3400 VSS.n3399 0.0254457
R73511 VSS.n4097 VSS.n552 0.0251695
R73512 VSS.n4197 VSS.n536 0.0251695
R73513 VSS.n5859 VSS.n5857 0.0251695
R73514 VSS.n4093 VSS.n4092 0.0251695
R73515 VSS.n4185 VSS.n535 0.0251695
R73516 VSS.n5485 VSS.n5484 0.0251695
R73517 VSS.n4186 VSS.n4185 0.0251695
R73518 VSS.n4195 VSS.n536 0.0251695
R73519 VSS.n6188 VSS.n6187 0.0251695
R73520 VSS.n5497 VSS.n5496 0.0251695
R73521 VSS.n6160 VSS.n473 0.0251695
R73522 VSS.n6171 VSS.n472 0.0251695
R73523 VSS.n5493 VSS.n5492 0.0251695
R73524 VSS.n6172 VSS.n6171 0.0251695
R73525 VSS.n5493 VSS.n5491 0.0251695
R73526 VSS.n5498 VSS.n5497 0.0251695
R73527 VSS.n5486 VSS.n5484 0.0251695
R73528 VSS.n5860 VSS.n5859 0.0251695
R73529 VSS.n6158 VSS.n6157 0.0251695
R73530 VSS.n6190 VSS.n6189 0.0251695
R73531 VSS.n4091 VSS.n573 0.0251695
R73532 VSS.n4099 VSS.n4098 0.0251695
R73533 VSS.n1220 VSS.n1219 0.0248
R73534 VSS.n1223 VSS.n1218 0.024575
R73535 VSS.n4945 VSS.n4933 0.0239
R73536 VSS.n5798 VSS.n5069 0.0239
R73537 VSS.n5120 VSS.n5012 0.0239
R73538 VSS.n5841 VSS.n4996 0.0239
R73539 VSS.n6025 VSS.n4421 0.0209851
R73540 VSS.n5526 VSS.n5525 0.0209851
R73541 VSS.n4500 VSS.n480 0.0203134
R73542 VSS.n5464 VSS.n5256 0.0203134
R73543 VSS.n5079 VSS.n5037 0.0203134
R73544 VSS.n4513 VSS.n502 0.0203
R73545 VSS.n4770 VSS.n4514 0.0203
R73546 VSS.n4508 VSS.n4507 0.0203
R73547 VSS.n4510 VSS.n4509 0.0203
R73548 VSS.n2875 VSS.n1119 0.0202719
R73549 VSS.n2894 VSS.n2893 0.0202719
R73550 VSS.n2904 VSS.n2903 0.0202719
R73551 VSS.n2875 VSS.n1127 0.0202719
R73552 VSS.n2893 VSS.n1127 0.0202719
R73553 VSS.n2904 VSS.n1127 0.0202719
R73554 VSS.n2974 VSS.n2973 0.0199776
R73555 VSS.n2970 VSS.n1106 0.0199776
R73556 VSS.n1093 VSS.n1082 0.01985
R73557 VSS.n2985 VSS.n2984 0.01985
R73558 VSS.n2919 VSS.n2918 0.01985
R73559 VSS.n2917 VSS.n2916 0.01985
R73560 VSS.n1662 VSS.n1326 0.0198097
R73561 VSS.n1892 VSS.n1224 0.0196418
R73562 VSS.n4813 VSS.n4424 0.0196418
R73563 VSS.n5519 VSS.n5518 0.0196418
R73564 VSS.n1251 VSS.n1229 0.0194
R73565 VSS.n1281 VSS.n1225 0.0194
R73566 VSS.n1537 VSS.n1213 0.0194
R73567 VSS.n1212 VSS.n1207 0.0194
R73568 VSS.n2549 VSS.n2548 0.0192079
R73569 VSS.n6452 VSS.n13 0.019095
R73570 VSS.n6210 VSS.n13 0.019095
R73571 VSS.n6211 VSS.n6210 0.019095
R73572 VSS.n6212 VSS.n6211 0.019095
R73573 VSS.n6212 VSS.n6199 0.019095
R73574 VSS.n139 VSS.n138 0.019095
R73575 VSS.n138 VSS.n15 0.019095
R73576 VSS.n6451 VSS.n15 0.019095
R73577 VSS.n6452 VSS.n6451 0.019095
R73578 VSS.n5470 VSS.n5469 0.0189701
R73579 VSS.n5099 VSS.n5094 0.0189701
R73580 VSS.n3280 VSS.n3279 0.0188287
R73581 VSS.n4825 VSS.n4401 0.0182985
R73582 VSS.n5536 VSS.n5508 0.0182985
R73583 VSS.n3209 VSS.n3205 0.0180085
R73584 VSS.n3340 VSS.n3336 0.0180085
R73585 VSS.n3164 VSS.n3160 0.0180085
R73586 VSS.n3165 VSS.n3164 0.0180085
R73587 VSS.n3169 VSS.n3165 0.0180085
R73588 VSS.n3170 VSS.n3169 0.0180085
R73589 VSS.n3174 VSS.n3170 0.0180085
R73590 VSS.n3175 VSS.n3174 0.0180085
R73591 VSS.n3179 VSS.n3175 0.0180085
R73592 VSS.n3180 VSS.n3179 0.0180085
R73593 VSS.n3184 VSS.n3180 0.0180085
R73594 VSS.n3185 VSS.n3184 0.0180085
R73595 VSS.n3189 VSS.n3185 0.0180085
R73596 VSS.n3190 VSS.n3189 0.0180085
R73597 VSS.n3194 VSS.n3190 0.0180085
R73598 VSS.n3195 VSS.n3194 0.0180085
R73599 VSS.n3199 VSS.n3195 0.0180085
R73600 VSS.n3200 VSS.n3199 0.0180085
R73601 VSS.n3204 VSS.n3200 0.0180085
R73602 VSS.n3205 VSS.n3204 0.0180085
R73603 VSS.n3210 VSS.n3209 0.0180085
R73604 VSS.n3215 VSS.n3214 0.0180085
R73605 VSS.n3219 VSS.n3215 0.0180085
R73606 VSS.n3220 VSS.n3219 0.0180085
R73607 VSS.n3224 VSS.n3220 0.0180085
R73608 VSS.n3225 VSS.n3224 0.0180085
R73609 VSS.n3229 VSS.n3225 0.0180085
R73610 VSS.n3230 VSS.n3229 0.0180085
R73611 VSS.n3234 VSS.n3230 0.0180085
R73612 VSS.n3235 VSS.n3234 0.0180085
R73613 VSS.n3239 VSS.n3235 0.0180085
R73614 VSS.n3240 VSS.n3239 0.0180085
R73615 VSS.n3244 VSS.n3240 0.0180085
R73616 VSS.n3245 VSS.n3244 0.0180085
R73617 VSS.n3249 VSS.n3245 0.0180085
R73618 VSS.n3250 VSS.n3249 0.0180085
R73619 VSS.n3254 VSS.n3250 0.0180085
R73620 VSS.n3255 VSS.n3254 0.0180085
R73621 VSS.n3259 VSS.n3255 0.0180085
R73622 VSS.n3260 VSS.n3259 0.0180085
R73623 VSS.n3264 VSS.n3260 0.0180085
R73624 VSS.n3285 VSS.n3281 0.0180085
R73625 VSS.n3286 VSS.n3285 0.0180085
R73626 VSS.n3290 VSS.n3286 0.0180085
R73627 VSS.n3291 VSS.n3290 0.0180085
R73628 VSS.n3295 VSS.n3291 0.0180085
R73629 VSS.n3296 VSS.n3295 0.0180085
R73630 VSS.n3300 VSS.n3296 0.0180085
R73631 VSS.n3301 VSS.n3300 0.0180085
R73632 VSS.n3305 VSS.n3301 0.0180085
R73633 VSS.n3306 VSS.n3305 0.0180085
R73634 VSS.n3310 VSS.n3306 0.0180085
R73635 VSS.n3311 VSS.n3310 0.0180085
R73636 VSS.n3315 VSS.n3311 0.0180085
R73637 VSS.n3316 VSS.n3315 0.0180085
R73638 VSS.n3320 VSS.n3316 0.0180085
R73639 VSS.n3321 VSS.n3320 0.0180085
R73640 VSS.n3325 VSS.n3321 0.0180085
R73641 VSS.n3326 VSS.n3325 0.0180085
R73642 VSS.n3330 VSS.n3326 0.0180085
R73643 VSS.n3331 VSS.n3330 0.0180085
R73644 VSS.n3336 VSS.n3335 0.0180085
R73645 VSS.n3341 VSS.n3340 0.0180085
R73646 VSS.n3345 VSS.n3341 0.0180085
R73647 VSS.n3346 VSS.n3345 0.0180085
R73648 VSS.n3350 VSS.n3346 0.0180085
R73649 VSS.n3351 VSS.n3350 0.0180085
R73650 VSS.n3355 VSS.n3351 0.0180085
R73651 VSS.n3356 VSS.n3355 0.0180085
R73652 VSS.n3360 VSS.n3356 0.0180085
R73653 VSS.n3361 VSS.n3360 0.0180085
R73654 VSS.n3365 VSS.n3361 0.0180085
R73655 VSS.n3366 VSS.n3365 0.0180085
R73656 VSS.n3370 VSS.n3366 0.0180085
R73657 VSS.n3371 VSS.n3370 0.0180085
R73658 VSS.n3375 VSS.n3371 0.0180085
R73659 VSS.n3376 VSS.n3375 0.0180085
R73660 VSS.n3380 VSS.n3376 0.0180085
R73661 VSS.n3381 VSS.n3380 0.0180085
R73662 VSS.n3385 VSS.n3381 0.0180085
R73663 VSS.n3386 VSS.n3385 0.0180085
R73664 VSS.n2532 VSS.n2530 0.0178311
R73665 VSS.n2530 VSS.n2528 0.0178311
R73666 VSS.n2528 VSS.n2526 0.0178311
R73667 VSS.n2526 VSS.n2524 0.0178311
R73668 VSS.n2524 VSS.n2522 0.0178311
R73669 VSS.n2522 VSS.n2520 0.0178311
R73670 VSS.n2520 VSS.n2518 0.0178311
R73671 VSS.n2518 VSS.n2516 0.0178311
R73672 VSS.n2516 VSS.n2514 0.0178311
R73673 VSS.n2514 VSS.n2512 0.0178311
R73674 VSS.n2512 VSS.n2510 0.0178311
R73675 VSS.n2510 VSS.n2508 0.0178311
R73676 VSS.n2508 VSS.n2506 0.0178311
R73677 VSS.n2506 VSS.n2504 0.0178311
R73678 VSS.n2504 VSS.n2502 0.0178311
R73679 VSS.n2502 VSS.n2500 0.0178311
R73680 VSS.n2500 VSS.n2498 0.0178311
R73681 VSS.n2498 VSS.n2496 0.0178311
R73682 VSS.n2496 VSS.n2494 0.0178311
R73683 VSS.n2494 VSS.n2492 0.0178311
R73684 VSS.n2492 VSS.n2490 0.0178311
R73685 VSS.n2490 VSS.n2488 0.0178311
R73686 VSS.n2488 VSS.n2486 0.0178311
R73687 VSS.n2484 VSS.n2482 0.0178311
R73688 VSS.n2482 VSS.n2480 0.0178311
R73689 VSS.n2480 VSS.n2478 0.0178311
R73690 VSS.n2478 VSS.n2476 0.0178311
R73691 VSS.n2476 VSS.n2474 0.0178311
R73692 VSS.n2474 VSS.n2472 0.0178311
R73693 VSS.n2472 VSS.n2470 0.0178311
R73694 VSS.n2470 VSS.n2468 0.0178311
R73695 VSS.n2468 VSS.n2466 0.0178311
R73696 VSS.n2466 VSS.n2464 0.0178311
R73697 VSS.n2464 VSS.n2462 0.0178311
R73698 VSS.n2462 VSS.n2460 0.0178311
R73699 VSS.n2460 VSS.n2458 0.0178311
R73700 VSS.n2458 VSS.n2456 0.0178311
R73701 VSS.n2456 VSS.n2454 0.0178311
R73702 VSS.n2454 VSS.n2452 0.0178311
R73703 VSS.n2452 VSS.n2450 0.0178311
R73704 VSS.n2450 VSS.n2448 0.0178311
R73705 VSS.n2448 VSS.n2446 0.0178311
R73706 VSS.n2446 VSS.n2224 0.0178311
R73707 VSS.n2412 VSS.n2225 0.0178311
R73708 VSS.n2412 VSS.n2411 0.0178311
R73709 VSS.n2411 VSS.n2409 0.0178311
R73710 VSS.n2409 VSS.n2407 0.0178311
R73711 VSS.n2407 VSS.n2405 0.0178311
R73712 VSS.n2405 VSS.n2403 0.0178311
R73713 VSS.n2403 VSS.n2401 0.0178311
R73714 VSS.n2401 VSS.n2399 0.0178311
R73715 VSS.n2399 VSS.n2397 0.0178311
R73716 VSS.n2397 VSS.n2395 0.0178311
R73717 VSS.n2395 VSS.n2393 0.0178311
R73718 VSS.n2393 VSS.n2391 0.0178311
R73719 VSS.n2391 VSS.n2389 0.0178311
R73720 VSS.n2389 VSS.n2387 0.0178311
R73721 VSS.n2387 VSS.n2385 0.0178311
R73722 VSS.n2385 VSS.n2383 0.0178311
R73723 VSS.n2383 VSS.n2381 0.0178311
R73724 VSS.n2381 VSS.n2379 0.0178311
R73725 VSS.n2379 VSS.n2377 0.0178311
R73726 VSS.n2377 VSS.n2375 0.0178311
R73727 VSS.n2373 VSS.n2371 0.0178311
R73728 VSS.n2371 VSS.n2369 0.0178311
R73729 VSS.n2369 VSS.n2367 0.0178311
R73730 VSS.n2367 VSS.n2365 0.0178311
R73731 VSS.n2365 VSS.n2363 0.0178311
R73732 VSS.n2363 VSS.n2361 0.0178311
R73733 VSS.n2361 VSS.n2359 0.0178311
R73734 VSS.n2359 VSS.n2357 0.0178311
R73735 VSS.n2357 VSS.n2355 0.0178311
R73736 VSS.n2355 VSS.n2353 0.0178311
R73737 VSS.n2353 VSS.n2351 0.0178311
R73738 VSS.n2351 VSS.n2349 0.0178311
R73739 VSS.n2349 VSS.n2347 0.0178311
R73740 VSS.n2347 VSS.n2345 0.0178311
R73741 VSS.n2345 VSS.n2343 0.0178311
R73742 VSS.n2343 VSS.n2341 0.0178311
R73743 VSS.n2341 VSS.n2339 0.0178311
R73744 VSS.n2339 VSS.n2337 0.0178311
R73745 VSS.n2337 VSS.n2335 0.0178311
R73746 VSS.n2335 VSS.n2333 0.0178311
R73747 VSS.n2333 VSS.n2331 0.0178311
R73748 VSS.n2331 VSS.n2329 0.0178311
R73749 VSS.n2329 VSS.n2327 0.0178311
R73750 VSS.n6149 VSS.n482 0.0176269
R73751 VSS.n5582 VSS.n4978 0.0176269
R73752 VSS.n5110 VSS.n5105 0.0176269
R73753 VSS.n6198 VSS.n449 0.0171667
R73754 VSS.n6219 VSS.n449 0.0171667
R73755 VSS.n448 VSS.n447 0.0171667
R73756 VSS.n1609 VSS.n448 0.0171667
R73757 VSS.n3280 VSS.n3264 0.017087
R73758 VSS.n1222 VSS.n1221 0.0169552
R73759 VSS.n4837 VSS.n4392 0.0169552
R73760 VSS.n2549 VSS.n2224 0.0169189
R73761 VSS.n730 VSS.n726 0.0167873
R73762 VSS.n3862 VSS.n732 0.0167873
R73763 VSS.n5863 VSS.n4918 0.0167
R73764 VSS.n5799 VSS.n5055 0.0167
R73765 VSS.n5834 VSS.n5015 0.0167
R73766 VSS.n5838 VSS.n4984 0.0167
R73767 VSS.n1890 VSS.n1226 0.0165729
R73768 VSS.n1886 VSS.n1230 0.0165729
R73769 VSS.n1896 VSS.n1214 0.0165729
R73770 VSS.n1899 VSS.n1211 0.0165729
R73771 VSS.n1884 VSS.n1230 0.0165729
R73772 VSS.n1888 VSS.n1226 0.0165729
R73773 VSS.n1894 VSS.n1214 0.0165729
R73774 VSS.n1900 VSS.n1899 0.0165729
R73775 VSS.n3331 DVSS 0.0163191
R73776 VSS.n5810 VSS.n5809 0.0162836
R73777 VSS.n2375 DVSS 0.0161588
R73778 VSS.n4857 VSS.n4856 0.0158
R73779 VSS.n4848 VSS.n4846 0.0158
R73780 VSS.n4850 VSS.n4297 0.0158
R73781 VSS.n4851 VSS.n4313 0.0158
R73782 VSS.n2888 VSS.n1154 0.0157916
R73783 VSS.n2898 VSS.n2889 0.0157916
R73784 VSS.n1157 VSS.n1155 0.0157916
R73785 VSS.n2972 VSS.n1118 0.0157916
R73786 VSS.n2969 VSS.n1117 0.0157916
R73787 VSS.n2964 VSS.n1122 0.0157916
R73788 VSS.n2882 VSS.n1151 0.0157916
R73789 VSS.n2901 VSS.n1136 0.0157916
R73790 VSS.n2962 VSS.n1122 0.0157916
R73791 VSS.n2927 VSS.n1157 0.0157916
R73792 VSS.n2972 VSS.n2971 0.0157916
R73793 VSS.n2965 VSS.n1117 0.0157916
R73794 VSS.n2896 VSS.n2888 0.0157916
R73795 VSS.n2883 VSS.n2882 0.0157916
R73796 VSS.n2902 VSS.n2901 0.0157916
R73797 VSS.n2891 VSS.n2889 0.0157916
R73798 VSS.n6218 VSS.n6217 0.015774
R73799 VSS.n6220 VSS.n124 0.015774
R73800 VSS.n4849 VSS.n4406 0.0156119
R73801 VSS.n140 VSS.n128 0.0155703
R73802 VSS.n1860 VSS.n1859 0.0154891
R73803 VSS.n2896 VSS.n2894 0.0153404
R73804 VSS.n2894 VSS.n2891 0.0153404
R73805 VSS.n2971 VSS.n1119 0.0153404
R73806 VSS.n2969 VSS.n1119 0.0153404
R73807 VSS.n2903 VSS.n2883 0.0153404
R73808 VSS.n2903 VSS.n2902 0.0153404
R73809 VSS.n5829 VSS.n5024 0.0152761
R73810 VSS.n2554 VSS.n2553 0.0149101
R73811 VSS.n2673 VSS.n2554 0.0149101
R73812 VSS.n2673 VSS.n2672 0.0149101
R73813 VSS.n2672 VSS.n2671 0.0149101
R73814 VSS.n2671 VSS.n2555 0.0149101
R73815 VSS.n2661 VSS.n2555 0.0149101
R73816 VSS.n2661 VSS.n2660 0.0149101
R73817 VSS.n2660 VSS.n2659 0.0149101
R73818 VSS.n2659 VSS.n2565 0.0149101
R73819 VSS.n2649 VSS.n2565 0.0149101
R73820 VSS.n2648 VSS.n2647 0.0149101
R73821 VSS.n2647 VSS.n2575 0.0149101
R73822 VSS.n2637 VSS.n2575 0.0149101
R73823 VSS.n2637 VSS.n2636 0.0149101
R73824 VSS.n2636 VSS.n2635 0.0149101
R73825 VSS.n2635 VSS.n2585 0.0149101
R73826 VSS.n2625 VSS.n2585 0.0149101
R73827 VSS.n2625 VSS.n2624 0.0149101
R73828 VSS.n2624 VSS.n2623 0.0149101
R73829 VSS.n3923 VSS.n3922 0.0149101
R73830 VSS.n3922 VSS.n675 0.0149101
R73831 VSS.n3912 VSS.n675 0.0149101
R73832 VSS.n3912 VSS.n3911 0.0149101
R73833 VSS.n3911 VSS.n3910 0.0149101
R73834 VSS.n3910 VSS.n685 0.0149101
R73835 VSS.n3900 VSS.n685 0.0149101
R73836 VSS.n3900 VSS.n3899 0.0149101
R73837 VSS.n3899 VSS.n3898 0.0149101
R73838 VSS.n3888 VSS.n704 0.0149101
R73839 VSS.n3888 VSS.n3887 0.0149101
R73840 VSS.n3887 VSS.n3886 0.0149101
R73841 VSS.n3886 VSS.n705 0.0149101
R73842 VSS.n3876 VSS.n705 0.0149101
R73843 VSS.n3876 VSS.n3875 0.0149101
R73844 VSS.n3875 VSS.n3874 0.0149101
R73845 VSS.n3874 VSS.n715 0.0149101
R73846 VSS.n3848 VSS.n752 0.0149101
R73847 VSS.n3848 VSS.n3847 0.0149101
R73848 VSS.n3847 VSS.n3846 0.0149101
R73849 VSS.n3846 VSS.n753 0.0149101
R73850 VSS.n3836 VSS.n753 0.0149101
R73851 VSS.n3836 VSS.n3835 0.0149101
R73852 VSS.n3835 VSS.n3834 0.0149101
R73853 VSS.n3834 VSS.n763 0.0149101
R73854 VSS.n3824 VSS.n3823 0.0149101
R73855 VSS.n3823 VSS.n3822 0.0149101
R73856 VSS.n3822 VSS.n773 0.0149101
R73857 VSS.n3812 VSS.n773 0.0149101
R73858 VSS.n3812 VSS.n3811 0.0149101
R73859 VSS.n3811 VSS.n3810 0.0149101
R73860 VSS.n3810 VSS.n783 0.0149101
R73861 VSS.n3800 VSS.n783 0.0149101
R73862 VSS.n3800 VSS.n3799 0.0149101
R73863 VSS.n3786 VSS.n803 0.0149101
R73864 VSS.n3786 VSS.n3785 0.0149101
R73865 VSS.n3785 VSS.n3784 0.0149101
R73866 VSS.n3784 VSS.n804 0.0149101
R73867 VSS.n3774 VSS.n804 0.0149101
R73868 VSS.n3774 VSS.n3773 0.0149101
R73869 VSS.n3773 VSS.n3772 0.0149101
R73870 VSS.n3772 VSS.n814 0.0149101
R73871 VSS.n3762 VSS.n814 0.0149101
R73872 VSS.n3761 VSS.n3760 0.0149101
R73873 VSS.n3760 VSS.n824 0.0149101
R73874 VSS.n3750 VSS.n824 0.0149101
R73875 VSS.n3750 VSS.n3749 0.0149101
R73876 VSS.n3749 VSS.n3748 0.0149101
R73877 VSS.n3748 VSS.n834 0.0149101
R73878 VSS.n3738 VSS.n834 0.0149101
R73879 VSS.n3738 VSS.n3737 0.0149101
R73880 VSS.n3737 VSS.n3736 0.0149101
R73881 VSS.n3736 VSS.n844 0.0149101
R73882 VSS.n3978 VSS.n569 0.0147724
R73883 VSS.n3281 VSS.n3280 0.0146297
R73884 VSS.n2549 VSS.n2225 0.0144865
R73885 VSS.n1796 VSS.n1795 0.0142903
R73886 VSS.n3035 VSS.n3034 0.0142903
R73887 VSS.n1020 VSS.n1019 0.0142903
R73888 VSS.n4060 VSS.n4059 0.0142903
R73889 VSS.n4698 VSS.n4697 0.0142903
R73890 VSS.n3864 VSS.n3863 0.0142781
R73891 VSS.n3861 VSS.n3858 0.0142781
R73892 VSS.n1424 VSS.n1217 0.0142687
R73893 VSS.n4128 VSS.n554 0.0141679
R73894 VSS.n4131 VSS.n555 0.0141679
R73895 VSS.n5836 VSS.n5011 0.0141679
R73896 VSS.n5835 VSS.n5013 0.0141679
R73897 VSS.n5020 VSS.n5016 0.0141679
R73898 VSS.n5827 VSS.n5020 0.0141679
R73899 VSS.n5025 VSS.n5019 0.0141679
R73900 VSS.n5025 VSS.n5022 0.0141679
R73901 VSS.n5801 VSS.n5023 0.0141679
R73902 VSS.n5865 VSS.n4944 0.0141679
R73903 VSS.n5837 VSS.n5836 0.0141679
R73904 VSS.n5833 VSS.n5013 0.0141679
R73905 VSS.n5801 VSS.n5800 0.0141679
R73906 VSS.n5865 VSS.n5864 0.0141679
R73907 VSS.n5828 VSS.n5019 0.0141679
R73908 VSS.n5828 VSS.n5827 0.0141679
R73909 VSS.n5830 VSS.n5022 0.0141679
R73910 VSS.n5832 VSS.n5016 0.0141679
R73911 VSS.n4130 VSS.n554 0.0141679
R73912 VSS.n4131 VSS.n556 0.0141679
R73913 VSS.n2977 VSS.n1097 0.0141007
R73914 VSS.n2980 VSS.n1099 0.0141007
R73915 VSS.n5051 VSS.n4921 0.014
R73916 VSS.n5806 VSS.n5805 0.014
R73917 VSS.n5118 VSS.n5085 0.014
R73918 VSS.n5116 VSS.n5000 0.014
R73919 VSS.n4773 VSS.n4495 0.0139328
R73920 VSS.n3214 DVSS 0.0138618
R73921 DVSS VSS.n2484 0.0137264
R73922 VSS.n3930 VSS.n665 0.0137065
R73923 VSS.n3792 VSS.n3791 0.0137065
R73924 VSS.n3506 VSS.n969 0.0137065
R73925 VSS.n3439 VSS.n972 0.0137065
R73926 VSS.n2134 VSS.n2133 0.013408
R73927 VSS.n3799 VSS.n3798 0.0133933
R73928 VSS.n6234 VSS.n6225 0.0131563
R73929 VSS.n6235 VSS.n6234 0.0131563
R73930 VSS.n6228 VSS.n6227 0.0130581
R73931 VSS.n134 VSS.n131 0.0130581
R73932 VSS.n725 VSS.n715 0.013014
R73933 VSS.n752 VSS.n731 0.013014
R73934 VSS.n5388 VSS.n5387 0.0127609
R73935 VSS.n5378 VSS.n5329 0.0127609
R73936 VSS.n5384 VSS.n5330 0.0127528
R73937 VSS.n3924 VSS.n3923 0.0126348
R73938 VSS.n3898 DVSS 0.0126348
R73939 VSS.n5826 VSS.n5017 0.0125896
R73940 VSS.n1255 VSS.n1254 0.0122
R73941 VSS.n4845 VSS.n4844 0.0122
R73942 VSS.n1280 VSS.n1279 0.0122
R73943 VSS.n4836 VSS.n4834 0.0122
R73944 VSS.n1535 VSS.n1534 0.0122
R73945 VSS.n4838 VSS.n4306 0.0122
R73946 VSS.n1898 VSS.n1206 0.0122
R73947 VSS.n4839 VSS.n4324 0.0122
R73948 VSS.n5501 VSS.n4386 0.0119179
R73949 VSS.n5831 VSS.n5021 0.0119179
R73950 VSS.n142 VSS.n11 0.0119115
R73951 VSS.n6457 VSS.n6456 0.0119115
R73952 VSS.n3824 DVSS 0.0118764
R73953 VSS.n3925 VSS.n674 0.0114972
R73954 VSS.n3797 VSS.n793 0.0114972
R73955 VSS.n1324 VSS.n1315 0.0113864
R73956 VSS.n1316 VSS.n1308 0.0113864
R73957 VSS.n1323 VSS.n1314 0.0113864
R73958 VSS.n1317 VSS.n1309 0.0113864
R73959 VSS.n1322 VSS.n1313 0.0113864
R73960 VSS.n1318 VSS.n1310 0.0113864
R73961 VSS.n1321 VSS.n1312 0.0113864
R73962 VSS.n1319 VSS.n1311 0.0113864
R73963 VSS.n1495 VSS.n1429 0.0113864
R73964 VSS.n1494 VSS.n1435 0.0113864
R73965 VSS.n1490 VSS.n1428 0.0113864
R73966 VSS.n1497 VSS.n1431 0.0113864
R73967 VSS.n1498 VSS.n1430 0.0113864
R73968 VSS.n1436 VSS.n1425 0.0113864
R73969 VSS.n1492 VSS.n1427 0.0113864
R73970 VSS.n2941 VSS.n1143 0.0113864
R73971 VSS.n2885 VSS.n2884 0.0113864
R73972 VSS.n2900 VSS.n2886 0.0113864
R73973 VSS.n2897 VSS.n2887 0.0113864
R73974 VSS.n2895 VSS.n2890 0.0113864
R73975 VSS.n2967 VSS.n2966 0.0113864
R73976 VSS.n1113 VSS.n1111 0.0113864
R73977 VSS.n1115 VSS.n1114 0.0113864
R73978 VSS.n1110 VSS.n1109 0.0113864
R73979 VSS.n2976 VSS.n1102 0.0113864
R73980 VSS.n2816 VSS.n1108 0.0113864
R73981 VSS.n2748 VSS.n2738 0.0113864
R73982 VSS.n2820 VSS.n2815 0.0113864
R73983 VSS.n2749 VSS.n2739 0.0113864
R73984 VSS.n2819 VSS.n2814 0.0113864
R73985 VSS.n2750 VSS.n2740 0.0113864
R73986 VSS.n2818 VSS.n2813 0.0113864
R73987 VSS.n2751 VSS.n2741 0.0113864
R73988 VSS.n2817 VSS.n2812 0.0113864
R73989 VSS.n2752 VSS.n2742 0.0113864
R73990 VSS.n2825 VSS.n2744 0.0113864
R73991 VSS.n3860 VSS.n728 0.0113864
R73992 VSS.n3859 VSS.n737 0.0113864
R73993 VSS.n735 VSS.n729 0.0113864
R73994 VSS.n736 VSS.n726 0.0113864
R73995 VSS.n3590 VSS.n935 0.0113864
R73996 VSS.n936 VSS.n912 0.0113864
R73997 VSS.n946 VSS.n934 0.0113864
R73998 VSS.n3577 VSS.n913 0.0113864
R73999 VSS.n945 VSS.n933 0.0113864
R74000 VSS.n3578 VSS.n914 0.0113864
R74001 VSS.n944 VSS.n932 0.0113864
R74002 VSS.n3579 VSS.n915 0.0113864
R74003 VSS.n943 VSS.n931 0.0113864
R74004 VSS.n3580 VSS.n916 0.0113864
R74005 VSS.n942 VSS.n930 0.0113864
R74006 VSS.n3581 VSS.n917 0.0113864
R74007 VSS.n941 VSS.n929 0.0113864
R74008 VSS.n3582 VSS.n918 0.0113864
R74009 VSS.n940 VSS.n928 0.0113864
R74010 VSS.n3583 VSS.n919 0.0113864
R74011 VSS.n939 VSS.n927 0.0113864
R74012 VSS.n3584 VSS.n920 0.0113864
R74013 VSS.n938 VSS.n926 0.0113864
R74014 VSS.n3585 VSS.n921 0.0113864
R74015 VSS.n937 VSS.n925 0.0113864
R74016 VSS.n3586 VSS.n924 0.0113864
R74017 VSS.n637 VSS.n623 0.0113864
R74018 VSS.n636 VSS.n635 0.0113864
R74019 VSS.n3970 VSS.n624 0.0113864
R74020 VSS.n634 VSS.n633 0.0113864
R74021 VSS.n3971 VSS.n625 0.0113864
R74022 VSS.n632 VSS.n631 0.0113864
R74023 VSS.n3972 VSS.n626 0.0113864
R74024 VSS.n630 VSS.n629 0.0113864
R74025 VSS.n3973 VSS.n628 0.0113864
R74026 VSS.n627 VSS.n559 0.0113864
R74027 VSS.n4505 VSS.n4500 0.0113864
R74028 VSS.n4493 VSS.n4492 0.0113864
R74029 VSS.n4504 VSS.n4499 0.0113864
R74030 VSS.n4498 VSS.n4494 0.0113864
R74031 VSS.n4503 VSS.n4497 0.0113864
R74032 VSS.n4774 VSS.n4501 0.0113864
R74033 VSS.n4776 VSS.n4487 0.0113864
R74034 VSS.n4415 VSS.n4390 0.0113864
R74035 VSS.n4389 VSS.n4388 0.0113864
R74036 VSS.n4405 VSS.n4391 0.0113864
R74037 VSS.n4419 VSS.n4404 0.0113864
R74038 VSS.n4409 VSS.n4408 0.0113864
R74039 VSS.n4403 VSS.n4402 0.0113864
R74040 VSS.n4416 VSS.n4394 0.0113864
R74041 VSS.n4393 VSS.n4387 0.0113864
R74042 VSS.n4400 VSS.n4395 0.0113864
R74043 VSS.n4418 VSS.n4399 0.0113864
R74044 VSS.n4411 VSS.n4410 0.0113864
R74045 VSS.n4423 VSS.n4398 0.0113864
R74046 VSS.n4417 VSS.n4397 0.0113864
R74047 VSS.n6032 VSS.n4414 0.0113864
R74048 VSS.n6027 VSS.n4412 0.0113864
R74049 VSS.n6028 VSS.n6026 0.0113864
R74050 VSS.n6029 VSS.n4413 0.0113864
R74051 VSS.n6030 VSS.n4386 0.0113864
R74052 VSS.n5506 VSS.n5462 0.0113864
R74053 VSS.n5539 VSS.n5479 0.0113864
R74054 VSS.n5507 VSS.n5463 0.0113864
R74055 VSS.n5538 VSS.n5537 0.0113864
R74056 VSS.n5478 VSS.n5460 0.0113864
R74057 VSS.n5573 VSS.n5509 0.0113864
R74058 VSS.n5477 VSS.n5459 0.0113864
R74059 VSS.n5476 VSS.n5458 0.0113864
R74060 VSS.n5574 VSS.n5520 0.0113864
R74061 VSS.n5475 VSS.n5457 0.0113864
R74062 VSS.n5474 VSS.n5456 0.0113864
R74063 VSS.n5575 VSS.n5464 0.0113864
R74064 VSS.n5576 VSS.n5527 0.0113864
R74065 VSS.n5473 VSS.n5454 0.0113864
R74066 VSS.n5577 VSS.n5470 0.0113864
R74067 VSS.n5580 VSS.n5579 0.0113864
R74068 VSS.n5472 VSS.n5452 0.0113864
R74069 VSS.n5582 VSS.n5471 0.0113864
R74070 VSS.n5037 VSS.n5036 0.0113864
R74071 VSS.n5039 VSS.n5038 0.0113864
R74072 VSS.n5041 VSS.n5040 0.0113864
R74073 VSS.n5094 VSS.n5042 0.0113864
R74074 VSS.n5044 VSS.n5043 0.0113864
R74075 VSS.n5046 VSS.n5045 0.0113864
R74076 VSS.n5105 VSS.n5047 0.0113864
R74077 VSS.n5049 VSS.n5048 0.0113864
R74078 VSS.n5812 VSS.n5811 0.0113864
R74079 VSS.n5813 VSS.n5810 0.0113864
R74080 VSS.n5815 VSS.n5814 0.0113864
R74081 VSS.n5817 VSS.n5816 0.0113864
R74082 VSS.n5819 VSS.n5818 0.0113864
R74083 VSS.n5821 VSS.n5820 0.0113864
R74084 VSS.n5822 VSS.n5024 0.0113864
R74085 VSS.n5824 VSS.n5823 0.0113864
R74086 VSS.n1143 VSS.n1142 0.0113864
R74087 VSS.n2897 VSS.n2890 0.0113864
R74088 VSS.n2899 VSS.n2887 0.0113864
R74089 VSS.n2886 VSS.n2885 0.0113864
R74090 VSS.n2884 VSS.n1145 0.0113864
R74091 VSS.n4414 VSS.n4397 0.0113864
R74092 VSS.n4417 VSS.n4398 0.0113864
R74093 VSS.n4424 VSS.n4423 0.0113864
R74094 VSS.n4410 VSS.n4399 0.0113864
R74095 VSS.n4418 VSS.n4395 0.0113864
R74096 VSS.n4401 VSS.n4400 0.0113864
R74097 VSS.n4394 VSS.n4393 0.0113864
R74098 VSS.n4416 VSS.n4403 0.0113864
R74099 VSS.n4402 VSS.n4392 0.0113864
R74100 VSS.n4408 VSS.n4404 0.0113864
R74101 VSS.n4419 VSS.n4391 0.0113864
R74102 VSS.n4406 VSS.n4405 0.0113864
R74103 VSS.n4390 VSS.n4389 0.0113864
R74104 VSS.n4415 VSS.n4407 0.0113864
R74105 VSS.n4495 VSS.n4487 0.0113864
R74106 VSS.n4501 VSS.n4497 0.0113864
R74107 VSS.n4503 VSS.n4494 0.0113864
R74108 VSS.n4499 VSS.n4498 0.0113864
R74109 VSS.n4504 VSS.n4493 0.0113864
R74110 VSS.n4492 VSS.n483 0.0113864
R74111 VSS.n4505 VSS.n4491 0.0113864
R74112 VSS.n628 VSS.n627 0.0113864
R74113 VSS.n3973 VSS.n630 0.0113864
R74114 VSS.n629 VSS.n626 0.0113864
R74115 VSS.n3972 VSS.n632 0.0113864
R74116 VSS.n631 VSS.n625 0.0113864
R74117 VSS.n3971 VSS.n634 0.0113864
R74118 VSS.n633 VSS.n624 0.0113864
R74119 VSS.n3970 VSS.n636 0.0113864
R74120 VSS.n635 VSS.n623 0.0113864
R74121 VSS.n3978 VSS.n637 0.0113864
R74122 VSS.n3586 VSS.n925 0.0113864
R74123 VSS.n937 VSS.n921 0.0113864
R74124 VSS.n3585 VSS.n926 0.0113864
R74125 VSS.n938 VSS.n920 0.0113864
R74126 VSS.n3584 VSS.n927 0.0113864
R74127 VSS.n939 VSS.n919 0.0113864
R74128 VSS.n3583 VSS.n928 0.0113864
R74129 VSS.n940 VSS.n918 0.0113864
R74130 VSS.n3582 VSS.n929 0.0113864
R74131 VSS.n941 VSS.n917 0.0113864
R74132 VSS.n3581 VSS.n930 0.0113864
R74133 VSS.n942 VSS.n916 0.0113864
R74134 VSS.n3580 VSS.n931 0.0113864
R74135 VSS.n943 VSS.n915 0.0113864
R74136 VSS.n3579 VSS.n932 0.0113864
R74137 VSS.n944 VSS.n914 0.0113864
R74138 VSS.n3578 VSS.n933 0.0113864
R74139 VSS.n945 VSS.n913 0.0113864
R74140 VSS.n3577 VSS.n934 0.0113864
R74141 VSS.n946 VSS.n912 0.0113864
R74142 VSS.n3590 VSS.n936 0.0113864
R74143 VSS.n935 VSS.n732 0.0113864
R74144 VSS.n2752 VSS.n2744 0.0113864
R74145 VSS.n2812 VSS.n2742 0.0113864
R74146 VSS.n2817 VSS.n2751 0.0113864
R74147 VSS.n2813 VSS.n2741 0.0113864
R74148 VSS.n2818 VSS.n2750 0.0113864
R74149 VSS.n2814 VSS.n2740 0.0113864
R74150 VSS.n2819 VSS.n2749 0.0113864
R74151 VSS.n2815 VSS.n2739 0.0113864
R74152 VSS.n2820 VSS.n2748 0.0113864
R74153 VSS.n2823 VSS.n2738 0.0113864
R74154 VSS.n1108 VSS.n1099 0.0113864
R74155 VSS.n1109 VSS.n1102 0.0113864
R74156 VSS.n1114 VSS.n1110 0.0113864
R74157 VSS.n1115 VSS.n1113 0.0113864
R74158 VSS.n2966 VSS.n1111 0.0113864
R74159 VSS.n2968 VSS.n2967 0.0113864
R74160 VSS.n1492 VSS.n1436 0.0113864
R74161 VSS.n1425 VSS.n1224 0.0113864
R74162 VSS.n1498 VSS.n1497 0.0113864
R74163 VSS.n1490 VSS.n1431 0.0113864
R74164 VSS.n1435 VSS.n1428 0.0113864
R74165 VSS.n1495 VSS.n1494 0.0113864
R74166 VSS.n1434 VSS.n1429 0.0113864
R74167 VSS.n1319 VSS.n1312 0.0113864
R74168 VSS.n1321 VSS.n1310 0.0113864
R74169 VSS.n1318 VSS.n1313 0.0113864
R74170 VSS.n1322 VSS.n1309 0.0113864
R74171 VSS.n1317 VSS.n1314 0.0113864
R74172 VSS.n1323 VSS.n1308 0.0113864
R74173 VSS.n1316 VSS.n1315 0.0113864
R74174 VSS.n1324 VSS.n1307 0.0113864
R74175 VSS.n6025 VSS.n4412 0.0113864
R74176 VSS.n6028 VSS.n6027 0.0113864
R74177 VSS.n6026 VSS.n4413 0.0113864
R74178 VSS.n6030 VSS.n6029 0.0113864
R74179 VSS.n5504 VSS.n5462 0.0113864
R74180 VSS.n5539 VSS.n5506 0.0113864
R74181 VSS.n5479 VSS.n5463 0.0113864
R74182 VSS.n5538 VSS.n5507 0.0113864
R74183 VSS.n5508 VSS.n5460 0.0113864
R74184 VSS.n5573 VSS.n5478 0.0113864
R74185 VSS.n5509 VSS.n5459 0.0113864
R74186 VSS.n5519 VSS.n5458 0.0113864
R74187 VSS.n5574 VSS.n5476 0.0113864
R74188 VSS.n5520 VSS.n5457 0.0113864
R74189 VSS.n5526 VSS.n5456 0.0113864
R74190 VSS.n5575 VSS.n5474 0.0113864
R74191 VSS.n5527 VSS.n5455 0.0113864
R74192 VSS.n5576 VSS.n5454 0.0113864
R74193 VSS.n5577 VSS.n5473 0.0113864
R74194 VSS.n5580 VSS.n5453 0.0113864
R74195 VSS.n5579 VSS.n5452 0.0113864
R74196 VSS.n5472 VSS.n5471 0.0113864
R74197 VSS.n5036 VSS.n5034 0.0113864
R74198 VSS.n5038 VSS.n5033 0.0113864
R74199 VSS.n5040 VSS.n5039 0.0113864
R74200 VSS.n5042 VSS.n5041 0.0113864
R74201 VSS.n5043 VSS.n5032 0.0113864
R74202 VSS.n5045 VSS.n5044 0.0113864
R74203 VSS.n5047 VSS.n5046 0.0113864
R74204 VSS.n5048 VSS.n5031 0.0113864
R74205 VSS.n5811 VSS.n5049 0.0113864
R74206 VSS.n5813 VSS.n5812 0.0113864
R74207 VSS.n5814 VSS.n5030 0.0113864
R74208 VSS.n5816 VSS.n5815 0.0113864
R74209 VSS.n5818 VSS.n5817 0.0113864
R74210 VSS.n5820 VSS.n5819 0.0113864
R74211 VSS.n5822 VSS.n5821 0.0113864
R74212 VSS.n5823 VSS.n5021 0.0113864
R74213 VSS.n738 VSS.n728 0.0113864
R74214 VSS.n3860 VSS.n3859 0.0113864
R74215 VSS.n737 VSS.n729 0.0113864
R74216 VSS.n736 VSS.n735 0.0113864
R74217 VSS.n6228 VSS.n8 0.0110469
R74218 VSS.n6153 VSS.n477 0.0106562
R74219 VSS.n6154 VSS.n6153 0.0106562
R74220 VSS.n1592 VSS.n1551 0.0105
R74221 VSS.n1592 VSS.n1591 0.0105
R74222 VSS.n1591 VSS.n1590 0.0105
R74223 VSS.n1590 VSS.n1556 0.0105
R74224 VSS.n1586 VSS.n1556 0.0105
R74225 VSS.n1586 VSS.n1585 0.0105
R74226 VSS.n1585 VSS.n1584 0.0105
R74227 VSS.n1584 VSS.n1562 0.0105
R74228 VSS.n1580 VSS.n1562 0.0105
R74229 VSS.n1580 VSS.n1579 0.0105
R74230 VSS.n1579 VSS.n1578 0.0105
R74231 VSS.n1578 VSS.n1568 0.0105
R74232 VSS.n1574 VSS.n1568 0.0105
R74233 VSS.n1574 VSS.n1573 0.0105
R74234 VSS.n1573 VSS.n1345 0.0105
R74235 VSS.n1619 VSS.n1345 0.0105
R74236 VSS.n1619 VSS.n1343 0.0105
R74237 VSS.n1623 VSS.n1343 0.0105
R74238 VSS.n1623 VSS.n1341 0.0105
R74239 VSS.n1627 VSS.n1341 0.0105
R74240 VSS.n1627 VSS.n1339 0.0105
R74241 VSS.n1631 VSS.n1339 0.0105
R74242 VSS.n1631 VSS.n1337 0.0105
R74243 VSS.n1635 VSS.n1337 0.0105
R74244 VSS.n1635 VSS.n1335 0.0105
R74245 VSS.n1639 VSS.n1335 0.0105
R74246 VSS.n1639 VSS.n1333 0.0105
R74247 VSS.n1643 VSS.n1333 0.0105
R74248 VSS.n1643 VSS.n1331 0.0105
R74249 VSS.n1647 VSS.n1331 0.0105
R74250 VSS.n1647 VSS.n1329 0.0105
R74251 VSS.n1652 VSS.n1329 0.0105
R74252 VSS.n1652 VSS.n1327 0.0105
R74253 VSS.n1658 VSS.n1327 0.0105
R74254 VSS.n1658 VSS.n1657 0.0105
R74255 VSS.n1657 VSS.n1305 0.0105
R74256 VSS.n1666 VSS.n1305 0.0105
R74257 VSS.n1666 VSS.n1303 0.0105
R74258 VSS.n1670 VSS.n1303 0.0105
R74259 VSS.n1670 VSS.n1301 0.0105
R74260 VSS.n1674 VSS.n1301 0.0105
R74261 VSS.n1674 VSS.n1299 0.0105
R74262 VSS.n1678 VSS.n1299 0.0105
R74263 VSS.n1678 VSS.n1297 0.0105
R74264 VSS.n1682 VSS.n1297 0.0105
R74265 VSS.n1682 VSS.n1295 0.0105
R74266 VSS.n1686 VSS.n1295 0.0105
R74267 VSS.n1686 VSS.n1293 0.0105
R74268 VSS.n1690 VSS.n1293 0.0105
R74269 VSS.n1690 VSS.n1291 0.0105
R74270 VSS.n1737 VSS.n1291 0.0105
R74271 VSS.n1737 VSS.n1736 0.0105
R74272 VSS.n1736 VSS.n1735 0.0105
R74273 VSS.n1735 VSS.n1734 0.0105
R74274 VSS.n1734 VSS.n1697 0.0105
R74275 VSS.n1730 VSS.n1697 0.0105
R74276 VSS.n1730 VSS.n1729 0.0105
R74277 VSS.n1729 VSS.n1728 0.0105
R74278 VSS.n1728 VSS.n1703 0.0105
R74279 VSS.n1724 VSS.n1703 0.0105
R74280 VSS.n1724 VSS.n1723 0.0105
R74281 VSS.n1723 VSS.n1722 0.0105
R74282 VSS.n1722 VSS.n1709 0.0105
R74283 VSS.n1718 VSS.n1709 0.0105
R74284 VSS.n1718 VSS.n1717 0.0105
R74285 VSS.n1717 VSS.n1716 0.0105
R74286 VSS.n1716 VSS.n1244 0.0105
R74287 VSS.n1838 VSS.n1244 0.0105
R74288 VSS.n1838 VSS.n1242 0.0105
R74289 VSS.n1877 VSS.n1242 0.0105
R74290 VSS.n1877 VSS.n1876 0.0105
R74291 VSS.n1876 VSS.n1875 0.0105
R74292 VSS.n1875 VSS.n1844 0.0105
R74293 VSS.n1871 VSS.n1844 0.0105
R74294 VSS.n1871 VSS.n1870 0.0105
R74295 VSS.n1870 VSS.n1869 0.0105
R74296 VSS.n1869 VSS.n1850 0.0105
R74297 VSS.n1865 VSS.n1850 0.0105
R74298 VSS.n1865 VSS.n1864 0.0105
R74299 VSS.n1864 VSS.n1863 0.0105
R74300 VSS.n1863 VSS.n1856 0.0105
R74301 VSS.n1593 VSS.n1550 0.0105
R74302 VSS.n1589 VSS.n1550 0.0105
R74303 VSS.n1589 VSS.n1588 0.0105
R74304 VSS.n1588 VSS.n1587 0.0105
R74305 VSS.n1587 VSS.n1557 0.0105
R74306 VSS.n1583 VSS.n1557 0.0105
R74307 VSS.n1583 VSS.n1582 0.0105
R74308 VSS.n1582 VSS.n1581 0.0105
R74309 VSS.n1581 VSS.n1563 0.0105
R74310 VSS.n1577 VSS.n1563 0.0105
R74311 VSS.n1577 VSS.n1576 0.0105
R74312 VSS.n1576 VSS.n1575 0.0105
R74313 VSS.n1575 VSS.n1569 0.0105
R74314 VSS.n1569 VSS.n1346 0.0105
R74315 VSS.n1618 VSS.n1346 0.0105
R74316 VSS.n1625 VSS.n1624 0.0105
R74317 VSS.n1626 VSS.n1625 0.0105
R74318 VSS.n1626 VSS.n1338 0.0105
R74319 VSS.n1632 VSS.n1338 0.0105
R74320 VSS.n1633 VSS.n1632 0.0105
R74321 VSS.n1634 VSS.n1633 0.0105
R74322 VSS.n1634 VSS.n1334 0.0105
R74323 VSS.n1640 VSS.n1334 0.0105
R74324 VSS.n1641 VSS.n1640 0.0105
R74325 VSS.n1642 VSS.n1641 0.0105
R74326 VSS.n1642 VSS.n1330 0.0105
R74327 VSS.n1648 VSS.n1330 0.0105
R74328 VSS.n1649 VSS.n1648 0.0105
R74329 VSS.n1651 VSS.n1649 0.0105
R74330 VSS.n1651 VSS.n1650 0.0105
R74331 VSS.n1665 VSS.n1664 0.0105
R74332 VSS.n1665 VSS.n1302 0.0105
R74333 VSS.n1671 VSS.n1302 0.0105
R74334 VSS.n1672 VSS.n1671 0.0105
R74335 VSS.n1673 VSS.n1672 0.0105
R74336 VSS.n1673 VSS.n1298 0.0105
R74337 VSS.n1679 VSS.n1298 0.0105
R74338 VSS.n1680 VSS.n1679 0.0105
R74339 VSS.n1681 VSS.n1680 0.0105
R74340 VSS.n1681 VSS.n1294 0.0105
R74341 VSS.n1687 VSS.n1294 0.0105
R74342 VSS.n1688 VSS.n1687 0.0105
R74343 VSS.n1689 VSS.n1688 0.0105
R74344 VSS.n1689 VSS.n1290 0.0105
R74345 VSS.n1738 VSS.n1290 0.0105
R74346 VSS.n1733 VSS.n1285 0.0105
R74347 VSS.n1733 VSS.n1732 0.0105
R74348 VSS.n1732 VSS.n1731 0.0105
R74349 VSS.n1731 VSS.n1698 0.0105
R74350 VSS.n1727 VSS.n1698 0.0105
R74351 VSS.n1727 VSS.n1726 0.0105
R74352 VSS.n1726 VSS.n1725 0.0105
R74353 VSS.n1725 VSS.n1704 0.0105
R74354 VSS.n1721 VSS.n1704 0.0105
R74355 VSS.n1721 VSS.n1720 0.0105
R74356 VSS.n1720 VSS.n1719 0.0105
R74357 VSS.n1719 VSS.n1710 0.0105
R74358 VSS.n1715 VSS.n1710 0.0105
R74359 VSS.n1715 VSS.n1245 0.0105
R74360 VSS.n1837 VSS.n1245 0.0105
R74361 VSS.n1878 VSS.n1241 0.0105
R74362 VSS.n1874 VSS.n1241 0.0105
R74363 VSS.n1874 VSS.n1873 0.0105
R74364 VSS.n1873 VSS.n1872 0.0105
R74365 VSS.n1872 VSS.n1845 0.0105
R74366 VSS.n1868 VSS.n1845 0.0105
R74367 VSS.n1868 VSS.n1867 0.0105
R74368 VSS.n1867 VSS.n1866 0.0105
R74369 VSS.n1866 VSS.n1851 0.0105
R74370 VSS.n1862 VSS.n1851 0.0105
R74371 VSS.n1862 VSS.n1861 0.0105
R74372 VSS.n492 VSS.n490 0.0104
R74373 VSS.n5106 VSS.n4923 0.0104
R74374 VSS.n4764 VSS.n4763 0.0104
R74375 VSS.n5107 VSS.n5059 0.0104
R74376 VSS.n6116 VSS.n4269 0.0104
R74377 VSS.n5114 VSS.n5087 0.0104
R74378 VSS.n6127 VSS.n4264 0.0104
R74379 VSS.n5112 VSS.n5002 0.0104
R74380 VSS.n4129 VSS.n557 0.0100489
R74381 VSS.n4134 VSS.n553 0.0100489
R74382 VSS.n4183 VSS.n4177 0.0100489
R74383 VSS.n5503 VSS.n5480 0.0100489
R74384 VSS.n557 VSS.n553 0.0100489
R74385 VSS.n4132 VSS.n4129 0.0100489
R74386 VSS.n4189 VSS.n4177 0.0100489
R74387 VSS.n5501 VSS.n5480 0.0100489
R74388 VSS.n1742 VSS.n1738 0.010007
R74389 VSS.n5831 VSS.n5018 0.00990298
R74390 VSS.n1624 VSS.n1342 0.00972535
R74391 VSS.n1376 VSS.n1375 0.00962857
R74392 VSS.n1379 VSS.n1376 0.00962857
R74393 VSS.n1379 VSS.n1374 0.00962857
R74394 VSS.n1383 VSS.n1374 0.00962857
R74395 VSS.n1383 VSS.n1372 0.00962857
R74396 VSS.n1387 VSS.n1372 0.00962857
R74397 VSS.n1387 VSS.n1370 0.00962857
R74398 VSS.n1391 VSS.n1370 0.00962857
R74399 VSS.n1391 VSS.n1368 0.00962857
R74400 VSS.n1395 VSS.n1368 0.00962857
R74401 VSS.n1395 VSS.n1366 0.00962857
R74402 VSS.n1399 VSS.n1366 0.00962857
R74403 VSS.n1399 VSS.n1364 0.00962857
R74404 VSS.n1403 VSS.n1364 0.00962857
R74405 VSS.n1403 VSS.n1362 0.00962857
R74406 VSS.n1407 VSS.n1362 0.00962857
R74407 VSS.n1407 VSS.n1359 0.00962857
R74408 VSS.n1530 VSS.n1359 0.00962857
R74409 VSS.n1530 VSS.n1360 0.00962857
R74410 VSS.n1526 VSS.n1360 0.00962857
R74411 VSS.n1526 VSS.n1411 0.00962857
R74412 VSS.n1522 VSS.n1411 0.00962857
R74413 VSS.n1522 VSS.n1413 0.00962857
R74414 VSS.n1518 VSS.n1413 0.00962857
R74415 VSS.n1518 VSS.n1415 0.00962857
R74416 VSS.n1514 VSS.n1415 0.00962857
R74417 VSS.n1514 VSS.n1417 0.00962857
R74418 VSS.n1510 VSS.n1417 0.00962857
R74419 VSS.n1510 VSS.n1419 0.00962857
R74420 VSS.n1506 VSS.n1419 0.00962857
R74421 VSS.n1506 VSS.n1421 0.00962857
R74422 VSS.n1502 VSS.n1421 0.00962857
R74423 VSS.n1502 VSS.n1423 0.00962857
R74424 VSS.n1440 VSS.n1423 0.00962857
R74425 VSS.n1440 VSS.n1438 0.00962857
R74426 VSS.n1488 VSS.n1438 0.00962857
R74427 VSS.n1488 VSS.n1439 0.00962857
R74428 VSS.n1484 VSS.n1439 0.00962857
R74429 VSS.n1484 VSS.n1444 0.00962857
R74430 VSS.n1480 VSS.n1444 0.00962857
R74431 VSS.n1480 VSS.n1446 0.00962857
R74432 VSS.n1476 VSS.n1446 0.00962857
R74433 VSS.n1476 VSS.n1448 0.00962857
R74434 VSS.n1472 VSS.n1448 0.00962857
R74435 VSS.n1472 VSS.n1450 0.00962857
R74436 VSS.n1468 VSS.n1450 0.00962857
R74437 VSS.n1468 VSS.n1452 0.00962857
R74438 VSS.n1464 VSS.n1452 0.00962857
R74439 VSS.n1464 VSS.n1454 0.00962857
R74440 VSS.n1460 VSS.n1454 0.00962857
R74441 VSS.n1460 VSS.n1458 0.00962857
R74442 VSS.n1458 VSS.n1457 0.00962857
R74443 VSS.n1457 VSS.n1273 0.00962857
R74444 VSS.n1757 VSS.n1273 0.00962857
R74445 VSS.n1757 VSS.n1271 0.00962857
R74446 VSS.n1761 VSS.n1271 0.00962857
R74447 VSS.n1761 VSS.n1269 0.00962857
R74448 VSS.n1765 VSS.n1269 0.00962857
R74449 VSS.n1765 VSS.n1267 0.00962857
R74450 VSS.n1769 VSS.n1267 0.00962857
R74451 VSS.n1769 VSS.n1265 0.00962857
R74452 VSS.n1773 VSS.n1265 0.00962857
R74453 VSS.n1773 VSS.n1263 0.00962857
R74454 VSS.n1777 VSS.n1263 0.00962857
R74455 VSS.n1777 VSS.n1261 0.00962857
R74456 VSS.n1781 VSS.n1261 0.00962857
R74457 VSS.n1781 VSS.n1258 0.00962857
R74458 VSS.n1824 VSS.n1258 0.00962857
R74459 VSS.n1824 VSS.n1259 0.00962857
R74460 VSS.n1820 VSS.n1259 0.00962857
R74461 VSS.n1820 VSS.n1819 0.00962857
R74462 VSS.n1819 VSS.n1785 0.00962857
R74463 VSS.n1815 VSS.n1785 0.00962857
R74464 VSS.n1815 VSS.n1787 0.00962857
R74465 VSS.n1811 VSS.n1787 0.00962857
R74466 VSS.n1811 VSS.n1790 0.00962857
R74467 VSS.n1807 VSS.n1790 0.00962857
R74468 VSS.n1807 VSS.n1792 0.00962857
R74469 VSS.n1803 VSS.n1792 0.00962857
R74470 VSS.n1803 VSS.n1794 0.00962857
R74471 VSS.n1799 VSS.n1794 0.00962857
R74472 VSS.n1380 VSS.n1205 0.00962857
R74473 VSS.n1381 VSS.n1380 0.00962857
R74474 VSS.n1382 VSS.n1381 0.00962857
R74475 VSS.n1382 VSS.n1371 0.00962857
R74476 VSS.n1388 VSS.n1371 0.00962857
R74477 VSS.n1389 VSS.n1388 0.00962857
R74478 VSS.n1390 VSS.n1389 0.00962857
R74479 VSS.n1390 VSS.n1367 0.00962857
R74480 VSS.n1396 VSS.n1367 0.00962857
R74481 VSS.n1397 VSS.n1396 0.00962857
R74482 VSS.n1398 VSS.n1397 0.00962857
R74483 VSS.n1398 VSS.n1363 0.00962857
R74484 VSS.n1404 VSS.n1363 0.00962857
R74485 VSS.n1405 VSS.n1404 0.00962857
R74486 VSS.n1406 VSS.n1405 0.00962857
R74487 VSS.n1531 VSS.n1358 0.00962857
R74488 VSS.n1525 VSS.n1358 0.00962857
R74489 VSS.n1525 VSS.n1524 0.00962857
R74490 VSS.n1524 VSS.n1523 0.00962857
R74491 VSS.n1523 VSS.n1412 0.00962857
R74492 VSS.n1517 VSS.n1412 0.00962857
R74493 VSS.n1517 VSS.n1516 0.00962857
R74494 VSS.n1516 VSS.n1515 0.00962857
R74495 VSS.n1515 VSS.n1416 0.00962857
R74496 VSS.n1509 VSS.n1416 0.00962857
R74497 VSS.n1509 VSS.n1508 0.00962857
R74498 VSS.n1508 VSS.n1507 0.00962857
R74499 VSS.n1507 VSS.n1420 0.00962857
R74500 VSS.n1501 VSS.n1420 0.00962857
R74501 VSS.n1501 VSS.n1500 0.00962857
R74502 VSS.n1489 VSS.n1437 0.00962857
R74503 VSS.n1483 VSS.n1437 0.00962857
R74504 VSS.n1483 VSS.n1482 0.00962857
R74505 VSS.n1482 VSS.n1481 0.00962857
R74506 VSS.n1481 VSS.n1445 0.00962857
R74507 VSS.n1475 VSS.n1445 0.00962857
R74508 VSS.n1475 VSS.n1474 0.00962857
R74509 VSS.n1474 VSS.n1473 0.00962857
R74510 VSS.n1473 VSS.n1449 0.00962857
R74511 VSS.n1467 VSS.n1449 0.00962857
R74512 VSS.n1467 VSS.n1466 0.00962857
R74513 VSS.n1466 VSS.n1465 0.00962857
R74514 VSS.n1465 VSS.n1453 0.00962857
R74515 VSS.n1459 VSS.n1453 0.00962857
R74516 VSS.n1459 VSS.n1282 0.00962857
R74517 VSS.n1756 VSS.n1755 0.00962857
R74518 VSS.n1756 VSS.n1270 0.00962857
R74519 VSS.n1762 VSS.n1270 0.00962857
R74520 VSS.n1763 VSS.n1762 0.00962857
R74521 VSS.n1764 VSS.n1763 0.00962857
R74522 VSS.n1764 VSS.n1266 0.00962857
R74523 VSS.n1770 VSS.n1266 0.00962857
R74524 VSS.n1771 VSS.n1770 0.00962857
R74525 VSS.n1772 VSS.n1771 0.00962857
R74526 VSS.n1772 VSS.n1262 0.00962857
R74527 VSS.n1778 VSS.n1262 0.00962857
R74528 VSS.n1779 VSS.n1778 0.00962857
R74529 VSS.n1780 VSS.n1779 0.00962857
R74530 VSS.n1780 VSS.n1257 0.00962857
R74531 VSS.n1825 VSS.n1257 0.00962857
R74532 VSS.n1818 VSS.n1252 0.00962857
R74533 VSS.n1818 VSS.n1817 0.00962857
R74534 VSS.n1817 VSS.n1816 0.00962857
R74535 VSS.n1816 VSS.n1786 0.00962857
R74536 VSS.n1810 VSS.n1786 0.00962857
R74537 VSS.n1810 VSS.n1809 0.00962857
R74538 VSS.n1809 VSS.n1808 0.00962857
R74539 VSS.n1808 VSS.n1791 0.00962857
R74540 VSS.n1802 VSS.n1791 0.00962857
R74541 VSS.n1802 VSS.n1801 0.00962857
R74542 VSS.n1801 VSS.n1800 0.00962857
R74543 VSS.n2053 VSS.n1193 0.00962857
R74544 VSS.n2053 VSS.n1194 0.00962857
R74545 VSS.n2049 VSS.n1194 0.00962857
R74546 VSS.n2049 VSS.n1912 0.00962857
R74547 VSS.n2045 VSS.n1912 0.00962857
R74548 VSS.n2045 VSS.n1914 0.00962857
R74549 VSS.n2041 VSS.n1914 0.00962857
R74550 VSS.n2041 VSS.n1916 0.00962857
R74551 VSS.n2037 VSS.n1916 0.00962857
R74552 VSS.n2037 VSS.n1918 0.00962857
R74553 VSS.n2033 VSS.n1918 0.00962857
R74554 VSS.n2033 VSS.n1920 0.00962857
R74555 VSS.n2029 VSS.n1920 0.00962857
R74556 VSS.n2029 VSS.n1922 0.00962857
R74557 VSS.n2025 VSS.n1922 0.00962857
R74558 VSS.n2025 VSS.n2022 0.00962857
R74559 VSS.n2022 VSS.n2021 0.00962857
R74560 VSS.n2021 VSS.n1924 0.00962857
R74561 VSS.n2016 VSS.n1924 0.00962857
R74562 VSS.n2016 VSS.n1926 0.00962857
R74563 VSS.n2012 VSS.n1926 0.00962857
R74564 VSS.n2012 VSS.n1929 0.00962857
R74565 VSS.n2008 VSS.n1929 0.00962857
R74566 VSS.n2008 VSS.n1931 0.00962857
R74567 VSS.n2004 VSS.n1931 0.00962857
R74568 VSS.n2004 VSS.n1933 0.00962857
R74569 VSS.n2000 VSS.n1933 0.00962857
R74570 VSS.n2000 VSS.n1935 0.00962857
R74571 VSS.n1996 VSS.n1935 0.00962857
R74572 VSS.n1996 VSS.n1937 0.00962857
R74573 VSS.n1992 VSS.n1937 0.00962857
R74574 VSS.n1992 VSS.n1939 0.00962857
R74575 VSS.n1988 VSS.n1939 0.00962857
R74576 VSS.n1988 VSS.n1941 0.00962857
R74577 VSS.n1984 VSS.n1941 0.00962857
R74578 VSS.n1984 VSS.n1983 0.00962857
R74579 VSS.n1983 VSS.n1943 0.00962857
R74580 VSS.n1979 VSS.n1943 0.00962857
R74581 VSS.n1979 VSS.n1945 0.00962857
R74582 VSS.n1975 VSS.n1945 0.00962857
R74583 VSS.n1975 VSS.n1948 0.00962857
R74584 VSS.n1971 VSS.n1948 0.00962857
R74585 VSS.n1971 VSS.n1950 0.00962857
R74586 VSS.n1967 VSS.n1950 0.00962857
R74587 VSS.n1967 VSS.n1952 0.00962857
R74588 VSS.n1963 VSS.n1952 0.00962857
R74589 VSS.n1963 VSS.n1954 0.00962857
R74590 VSS.n1959 VSS.n1954 0.00962857
R74591 VSS.n1959 VSS.n1956 0.00962857
R74592 VSS.n1956 VSS.n1080 0.00962857
R74593 VSS.n2988 VSS.n1080 0.00962857
R74594 VSS.n2988 VSS.n1078 0.00962857
R74595 VSS.n2992 VSS.n1078 0.00962857
R74596 VSS.n2992 VSS.n1076 0.00962857
R74597 VSS.n2996 VSS.n1076 0.00962857
R74598 VSS.n2996 VSS.n1074 0.00962857
R74599 VSS.n3000 VSS.n1074 0.00962857
R74600 VSS.n3000 VSS.n1072 0.00962857
R74601 VSS.n3004 VSS.n1072 0.00962857
R74602 VSS.n3004 VSS.n1070 0.00962857
R74603 VSS.n3008 VSS.n1070 0.00962857
R74604 VSS.n3008 VSS.n1068 0.00962857
R74605 VSS.n3012 VSS.n1068 0.00962857
R74606 VSS.n3012 VSS.n1066 0.00962857
R74607 VSS.n3016 VSS.n1066 0.00962857
R74608 VSS.n3016 VSS.n1064 0.00962857
R74609 VSS.n3020 VSS.n1064 0.00962857
R74610 VSS.n3020 VSS.n1061 0.00962857
R74611 VSS.n3062 VSS.n1061 0.00962857
R74612 VSS.n3062 VSS.n1062 0.00962857
R74613 VSS.n3058 VSS.n1062 0.00962857
R74614 VSS.n3058 VSS.n3024 0.00962857
R74615 VSS.n3054 VSS.n3024 0.00962857
R74616 VSS.n3054 VSS.n3027 0.00962857
R74617 VSS.n3050 VSS.n3027 0.00962857
R74618 VSS.n3050 VSS.n3029 0.00962857
R74619 VSS.n3046 VSS.n3029 0.00962857
R74620 VSS.n3046 VSS.n3031 0.00962857
R74621 VSS.n3042 VSS.n3031 0.00962857
R74622 VSS.n3042 VSS.n3033 0.00962857
R74623 VSS.n3038 VSS.n3033 0.00962857
R74624 VSS.n2054 VSS.n1192 0.00962857
R74625 VSS.n2048 VSS.n1192 0.00962857
R74626 VSS.n2048 VSS.n2047 0.00962857
R74627 VSS.n2047 VSS.n2046 0.00962857
R74628 VSS.n2046 VSS.n1913 0.00962857
R74629 VSS.n2040 VSS.n1913 0.00962857
R74630 VSS.n2040 VSS.n2039 0.00962857
R74631 VSS.n2039 VSS.n2038 0.00962857
R74632 VSS.n2038 VSS.n1917 0.00962857
R74633 VSS.n2032 VSS.n1917 0.00962857
R74634 VSS.n2032 VSS.n2031 0.00962857
R74635 VSS.n2031 VSS.n2030 0.00962857
R74636 VSS.n2030 VSS.n1921 0.00962857
R74637 VSS.n2024 VSS.n1921 0.00962857
R74638 VSS.n2024 VSS.n2023 0.00962857
R74639 VSS.n2015 VSS.n1927 0.00962857
R74640 VSS.n2015 VSS.n2014 0.00962857
R74641 VSS.n2014 VSS.n2013 0.00962857
R74642 VSS.n2013 VSS.n1928 0.00962857
R74643 VSS.n2007 VSS.n1928 0.00962857
R74644 VSS.n2007 VSS.n2006 0.00962857
R74645 VSS.n2006 VSS.n2005 0.00962857
R74646 VSS.n2005 VSS.n1932 0.00962857
R74647 VSS.n1999 VSS.n1932 0.00962857
R74648 VSS.n1999 VSS.n1998 0.00962857
R74649 VSS.n1998 VSS.n1997 0.00962857
R74650 VSS.n1997 VSS.n1936 0.00962857
R74651 VSS.n1991 VSS.n1936 0.00962857
R74652 VSS.n1991 VSS.n1990 0.00962857
R74653 VSS.n1990 VSS.n1989 0.00962857
R74654 VSS.n1982 VSS.n1981 0.00962857
R74655 VSS.n1981 VSS.n1980 0.00962857
R74656 VSS.n1980 VSS.n1944 0.00962857
R74657 VSS.n1974 VSS.n1944 0.00962857
R74658 VSS.n1974 VSS.n1973 0.00962857
R74659 VSS.n1973 VSS.n1972 0.00962857
R74660 VSS.n1972 VSS.n1949 0.00962857
R74661 VSS.n1966 VSS.n1949 0.00962857
R74662 VSS.n1966 VSS.n1965 0.00962857
R74663 VSS.n1965 VSS.n1964 0.00962857
R74664 VSS.n1964 VSS.n1953 0.00962857
R74665 VSS.n1958 VSS.n1953 0.00962857
R74666 VSS.n1958 VSS.n1957 0.00962857
R74667 VSS.n1957 VSS.n1081 0.00962857
R74668 VSS.n2987 VSS.n1081 0.00962857
R74669 VSS.n2994 VSS.n2993 0.00962857
R74670 VSS.n2995 VSS.n2994 0.00962857
R74671 VSS.n2995 VSS.n1073 0.00962857
R74672 VSS.n3001 VSS.n1073 0.00962857
R74673 VSS.n3002 VSS.n3001 0.00962857
R74674 VSS.n3003 VSS.n3002 0.00962857
R74675 VSS.n3003 VSS.n1069 0.00962857
R74676 VSS.n3009 VSS.n1069 0.00962857
R74677 VSS.n3010 VSS.n3009 0.00962857
R74678 VSS.n3011 VSS.n3010 0.00962857
R74679 VSS.n3011 VSS.n1065 0.00962857
R74680 VSS.n3017 VSS.n1065 0.00962857
R74681 VSS.n3018 VSS.n3017 0.00962857
R74682 VSS.n3019 VSS.n3018 0.00962857
R74683 VSS.n3019 VSS.n1050 0.00962857
R74684 VSS.n3057 VSS.n3025 0.00962857
R74685 VSS.n3057 VSS.n3056 0.00962857
R74686 VSS.n3056 VSS.n3055 0.00962857
R74687 VSS.n3055 VSS.n3026 0.00962857
R74688 VSS.n3049 VSS.n3026 0.00962857
R74689 VSS.n3049 VSS.n3048 0.00962857
R74690 VSS.n3048 VSS.n3047 0.00962857
R74691 VSS.n3047 VSS.n3030 0.00962857
R74692 VSS.n3041 VSS.n3030 0.00962857
R74693 VSS.n3041 VSS.n3040 0.00962857
R74694 VSS.n3040 VSS.n3039 0.00962857
R74695 VSS.n2689 VSS.n1183 0.00962857
R74696 VSS.n2693 VSS.n1183 0.00962857
R74697 VSS.n2693 VSS.n1181 0.00962857
R74698 VSS.n2697 VSS.n1181 0.00962857
R74699 VSS.n2697 VSS.n1179 0.00962857
R74700 VSS.n2701 VSS.n1179 0.00962857
R74701 VSS.n2701 VSS.n1177 0.00962857
R74702 VSS.n2705 VSS.n1177 0.00962857
R74703 VSS.n2705 VSS.n1175 0.00962857
R74704 VSS.n2709 VSS.n1175 0.00962857
R74705 VSS.n2709 VSS.n1173 0.00962857
R74706 VSS.n2713 VSS.n1173 0.00962857
R74707 VSS.n2713 VSS.n1171 0.00962857
R74708 VSS.n2717 VSS.n1171 0.00962857
R74709 VSS.n2717 VSS.n1169 0.00962857
R74710 VSS.n2721 VSS.n1169 0.00962857
R74711 VSS.n2721 VSS.n1166 0.00962857
R74712 VSS.n2857 VSS.n1166 0.00962857
R74713 VSS.n2857 VSS.n1167 0.00962857
R74714 VSS.n2853 VSS.n1167 0.00962857
R74715 VSS.n2853 VSS.n2725 0.00962857
R74716 VSS.n2849 VSS.n2725 0.00962857
R74717 VSS.n2849 VSS.n2727 0.00962857
R74718 VSS.n2845 VSS.n2727 0.00962857
R74719 VSS.n2845 VSS.n2729 0.00962857
R74720 VSS.n2841 VSS.n2729 0.00962857
R74721 VSS.n2841 VSS.n2731 0.00962857
R74722 VSS.n2837 VSS.n2731 0.00962857
R74723 VSS.n2837 VSS.n2733 0.00962857
R74724 VSS.n2833 VSS.n2733 0.00962857
R74725 VSS.n2833 VSS.n2735 0.00962857
R74726 VSS.n2829 VSS.n2735 0.00962857
R74727 VSS.n2829 VSS.n2737 0.00962857
R74728 VSS.n2756 VSS.n2737 0.00962857
R74729 VSS.n2756 VSS.n2754 0.00962857
R74730 VSS.n2810 VSS.n2754 0.00962857
R74731 VSS.n2810 VSS.n2755 0.00962857
R74732 VSS.n2806 VSS.n2755 0.00962857
R74733 VSS.n2806 VSS.n2760 0.00962857
R74734 VSS.n2802 VSS.n2760 0.00962857
R74735 VSS.n2802 VSS.n2762 0.00962857
R74736 VSS.n2798 VSS.n2762 0.00962857
R74737 VSS.n2798 VSS.n2764 0.00962857
R74738 VSS.n2794 VSS.n2764 0.00962857
R74739 VSS.n2794 VSS.n2766 0.00962857
R74740 VSS.n2790 VSS.n2766 0.00962857
R74741 VSS.n2790 VSS.n2768 0.00962857
R74742 VSS.n2786 VSS.n2768 0.00962857
R74743 VSS.n2786 VSS.n2770 0.00962857
R74744 VSS.n2782 VSS.n2770 0.00962857
R74745 VSS.n2782 VSS.n2772 0.00962857
R74746 VSS.n2772 VSS.n981 0.00962857
R74747 VSS.n3434 VSS.n981 0.00962857
R74748 VSS.n3434 VSS.n982 0.00962857
R74749 VSS.n3430 VSS.n982 0.00962857
R74750 VSS.n3430 VSS.n985 0.00962857
R74751 VSS.n3426 VSS.n985 0.00962857
R74752 VSS.n3426 VSS.n987 0.00962857
R74753 VSS.n3422 VSS.n987 0.00962857
R74754 VSS.n3422 VSS.n989 0.00962857
R74755 VSS.n3418 VSS.n989 0.00962857
R74756 VSS.n3418 VSS.n991 0.00962857
R74757 VSS.n3414 VSS.n991 0.00962857
R74758 VSS.n3414 VSS.n993 0.00962857
R74759 VSS.n3410 VSS.n993 0.00962857
R74760 VSS.n3410 VSS.n995 0.00962857
R74761 VSS.n3406 VSS.n995 0.00962857
R74762 VSS.n3406 VSS.n997 0.00962857
R74763 VSS.n1005 VSS.n997 0.00962857
R74764 VSS.n1043 VSS.n1005 0.00962857
R74765 VSS.n1043 VSS.n1006 0.00962857
R74766 VSS.n1039 VSS.n1006 0.00962857
R74767 VSS.n1039 VSS.n1009 0.00962857
R74768 VSS.n1035 VSS.n1009 0.00962857
R74769 VSS.n1035 VSS.n1011 0.00962857
R74770 VSS.n1031 VSS.n1011 0.00962857
R74771 VSS.n1031 VSS.n1013 0.00962857
R74772 VSS.n1027 VSS.n1013 0.00962857
R74773 VSS.n1027 VSS.n1015 0.00962857
R74774 VSS.n1023 VSS.n1015 0.00962857
R74775 VSS.n1023 VSS.n1017 0.00962857
R74776 VSS.n2694 VSS.n1182 0.00962857
R74777 VSS.n2695 VSS.n2694 0.00962857
R74778 VSS.n2696 VSS.n2695 0.00962857
R74779 VSS.n2696 VSS.n1178 0.00962857
R74780 VSS.n2702 VSS.n1178 0.00962857
R74781 VSS.n2703 VSS.n2702 0.00962857
R74782 VSS.n2704 VSS.n2703 0.00962857
R74783 VSS.n2704 VSS.n1174 0.00962857
R74784 VSS.n2710 VSS.n1174 0.00962857
R74785 VSS.n2711 VSS.n2710 0.00962857
R74786 VSS.n2712 VSS.n2711 0.00962857
R74787 VSS.n2712 VSS.n1170 0.00962857
R74788 VSS.n2718 VSS.n1170 0.00962857
R74789 VSS.n2719 VSS.n2718 0.00962857
R74790 VSS.n2720 VSS.n2719 0.00962857
R74791 VSS.n2858 VSS.n1165 0.00962857
R74792 VSS.n2852 VSS.n1165 0.00962857
R74793 VSS.n2852 VSS.n2851 0.00962857
R74794 VSS.n2851 VSS.n2850 0.00962857
R74795 VSS.n2850 VSS.n2726 0.00962857
R74796 VSS.n2844 VSS.n2726 0.00962857
R74797 VSS.n2844 VSS.n2843 0.00962857
R74798 VSS.n2843 VSS.n2842 0.00962857
R74799 VSS.n2842 VSS.n2730 0.00962857
R74800 VSS.n2836 VSS.n2730 0.00962857
R74801 VSS.n2836 VSS.n2835 0.00962857
R74802 VSS.n2835 VSS.n2834 0.00962857
R74803 VSS.n2834 VSS.n2734 0.00962857
R74804 VSS.n2828 VSS.n2734 0.00962857
R74805 VSS.n2828 VSS.n2827 0.00962857
R74806 VSS.n2811 VSS.n2753 0.00962857
R74807 VSS.n2805 VSS.n2753 0.00962857
R74808 VSS.n2805 VSS.n2804 0.00962857
R74809 VSS.n2804 VSS.n2803 0.00962857
R74810 VSS.n2803 VSS.n2761 0.00962857
R74811 VSS.n2797 VSS.n2761 0.00962857
R74812 VSS.n2797 VSS.n2796 0.00962857
R74813 VSS.n2796 VSS.n2795 0.00962857
R74814 VSS.n2795 VSS.n2765 0.00962857
R74815 VSS.n2789 VSS.n2765 0.00962857
R74816 VSS.n2789 VSS.n2788 0.00962857
R74817 VSS.n2788 VSS.n2787 0.00962857
R74818 VSS.n2787 VSS.n2769 0.00962857
R74819 VSS.n2781 VSS.n2769 0.00962857
R74820 VSS.n2781 VSS.n2780 0.00962857
R74821 VSS.n3435 VSS.n980 0.00962857
R74822 VSS.n3429 VSS.n980 0.00962857
R74823 VSS.n3429 VSS.n3428 0.00962857
R74824 VSS.n3428 VSS.n3427 0.00962857
R74825 VSS.n3427 VSS.n986 0.00962857
R74826 VSS.n3421 VSS.n986 0.00962857
R74827 VSS.n3421 VSS.n3420 0.00962857
R74828 VSS.n3420 VSS.n3419 0.00962857
R74829 VSS.n3419 VSS.n990 0.00962857
R74830 VSS.n3413 VSS.n990 0.00962857
R74831 VSS.n3413 VSS.n3412 0.00962857
R74832 VSS.n3412 VSS.n3411 0.00962857
R74833 VSS.n3411 VSS.n994 0.00962857
R74834 VSS.n3405 VSS.n994 0.00962857
R74835 VSS.n3405 VSS.n3404 0.00962857
R74836 VSS.n1044 VSS.n1004 0.00962857
R74837 VSS.n1038 VSS.n1004 0.00962857
R74838 VSS.n1038 VSS.n1037 0.00962857
R74839 VSS.n1037 VSS.n1036 0.00962857
R74840 VSS.n1036 VSS.n1010 0.00962857
R74841 VSS.n1030 VSS.n1010 0.00962857
R74842 VSS.n1030 VSS.n1029 0.00962857
R74843 VSS.n1029 VSS.n1028 0.00962857
R74844 VSS.n1028 VSS.n1014 0.00962857
R74845 VSS.n1022 VSS.n1014 0.00962857
R74846 VSS.n1022 VSS.n1021 0.00962857
R74847 VSS.n2201 VSS.n2153 0.00962857
R74848 VSS.n2201 VSS.n2154 0.00962857
R74849 VSS.n2197 VSS.n2154 0.00962857
R74850 VSS.n2197 VSS.n2157 0.00962857
R74851 VSS.n2193 VSS.n2157 0.00962857
R74852 VSS.n2193 VSS.n2159 0.00962857
R74853 VSS.n2189 VSS.n2159 0.00962857
R74854 VSS.n2189 VSS.n2161 0.00962857
R74855 VSS.n2185 VSS.n2161 0.00962857
R74856 VSS.n2185 VSS.n2163 0.00962857
R74857 VSS.n2181 VSS.n2163 0.00962857
R74858 VSS.n2181 VSS.n2165 0.00962857
R74859 VSS.n2177 VSS.n2165 0.00962857
R74860 VSS.n2177 VSS.n2167 0.00962857
R74861 VSS.n2173 VSS.n2167 0.00962857
R74862 VSS.n2173 VSS.n2171 0.00962857
R74863 VSS.n2171 VSS.n2170 0.00962857
R74864 VSS.n2170 VSS.n653 0.00962857
R74865 VSS.n3940 VSS.n653 0.00962857
R74866 VSS.n3940 VSS.n651 0.00962857
R74867 VSS.n3944 VSS.n651 0.00962857
R74868 VSS.n3944 VSS.n649 0.00962857
R74869 VSS.n3948 VSS.n649 0.00962857
R74870 VSS.n3948 VSS.n647 0.00962857
R74871 VSS.n3952 VSS.n647 0.00962857
R74872 VSS.n3952 VSS.n645 0.00962857
R74873 VSS.n3956 VSS.n645 0.00962857
R74874 VSS.n3956 VSS.n643 0.00962857
R74875 VSS.n3960 VSS.n643 0.00962857
R74876 VSS.n3960 VSS.n641 0.00962857
R74877 VSS.n3964 VSS.n641 0.00962857
R74878 VSS.n3964 VSS.n639 0.00962857
R74879 VSS.n3968 VSS.n639 0.00962857
R74880 VSS.n3968 VSS.n621 0.00962857
R74881 VSS.n3981 VSS.n621 0.00962857
R74882 VSS.n3981 VSS.n619 0.00962857
R74883 VSS.n3985 VSS.n619 0.00962857
R74884 VSS.n3985 VSS.n617 0.00962857
R74885 VSS.n3989 VSS.n617 0.00962857
R74886 VSS.n3989 VSS.n615 0.00962857
R74887 VSS.n3993 VSS.n615 0.00962857
R74888 VSS.n3993 VSS.n613 0.00962857
R74889 VSS.n3997 VSS.n613 0.00962857
R74890 VSS.n3997 VSS.n611 0.00962857
R74891 VSS.n4001 VSS.n611 0.00962857
R74892 VSS.n4001 VSS.n609 0.00962857
R74893 VSS.n4005 VSS.n609 0.00962857
R74894 VSS.n4005 VSS.n607 0.00962857
R74895 VSS.n4009 VSS.n607 0.00962857
R74896 VSS.n4009 VSS.n605 0.00962857
R74897 VSS.n4013 VSS.n605 0.00962857
R74898 VSS.n4013 VSS.n603 0.00962857
R74899 VSS.n4017 VSS.n603 0.00962857
R74900 VSS.n4017 VSS.n601 0.00962857
R74901 VSS.n4021 VSS.n601 0.00962857
R74902 VSS.n4021 VSS.n599 0.00962857
R74903 VSS.n4025 VSS.n599 0.00962857
R74904 VSS.n4025 VSS.n597 0.00962857
R74905 VSS.n4029 VSS.n597 0.00962857
R74906 VSS.n4029 VSS.n595 0.00962857
R74907 VSS.n4033 VSS.n595 0.00962857
R74908 VSS.n4033 VSS.n593 0.00962857
R74909 VSS.n4037 VSS.n593 0.00962857
R74910 VSS.n4037 VSS.n591 0.00962857
R74911 VSS.n4041 VSS.n591 0.00962857
R74912 VSS.n4041 VSS.n589 0.00962857
R74913 VSS.n4045 VSS.n589 0.00962857
R74914 VSS.n4045 VSS.n586 0.00962857
R74915 VSS.n4087 VSS.n586 0.00962857
R74916 VSS.n4087 VSS.n587 0.00962857
R74917 VSS.n4083 VSS.n587 0.00962857
R74918 VSS.n4083 VSS.n4049 0.00962857
R74919 VSS.n4079 VSS.n4049 0.00962857
R74920 VSS.n4079 VSS.n4052 0.00962857
R74921 VSS.n4075 VSS.n4052 0.00962857
R74922 VSS.n4075 VSS.n4054 0.00962857
R74923 VSS.n4071 VSS.n4054 0.00962857
R74924 VSS.n4071 VSS.n4056 0.00962857
R74925 VSS.n4067 VSS.n4056 0.00962857
R74926 VSS.n4067 VSS.n4058 0.00962857
R74927 VSS.n4063 VSS.n4058 0.00962857
R74928 VSS.n2202 VSS.n2152 0.00962857
R74929 VSS.n2196 VSS.n2152 0.00962857
R74930 VSS.n2196 VSS.n2195 0.00962857
R74931 VSS.n2195 VSS.n2194 0.00962857
R74932 VSS.n2194 VSS.n2158 0.00962857
R74933 VSS.n2188 VSS.n2158 0.00962857
R74934 VSS.n2188 VSS.n2187 0.00962857
R74935 VSS.n2187 VSS.n2186 0.00962857
R74936 VSS.n2186 VSS.n2162 0.00962857
R74937 VSS.n2180 VSS.n2162 0.00962857
R74938 VSS.n2180 VSS.n2179 0.00962857
R74939 VSS.n2179 VSS.n2178 0.00962857
R74940 VSS.n2178 VSS.n2166 0.00962857
R74941 VSS.n2172 VSS.n2166 0.00962857
R74942 VSS.n2172 VSS.n660 0.00962857
R74943 VSS.n3939 VSS.n3938 0.00962857
R74944 VSS.n3939 VSS.n650 0.00962857
R74945 VSS.n3945 VSS.n650 0.00962857
R74946 VSS.n3946 VSS.n3945 0.00962857
R74947 VSS.n3947 VSS.n3946 0.00962857
R74948 VSS.n3947 VSS.n646 0.00962857
R74949 VSS.n3953 VSS.n646 0.00962857
R74950 VSS.n3954 VSS.n3953 0.00962857
R74951 VSS.n3955 VSS.n3954 0.00962857
R74952 VSS.n3955 VSS.n642 0.00962857
R74953 VSS.n3961 VSS.n642 0.00962857
R74954 VSS.n3962 VSS.n3961 0.00962857
R74955 VSS.n3963 VSS.n3962 0.00962857
R74956 VSS.n3963 VSS.n638 0.00962857
R74957 VSS.n3969 VSS.n638 0.00962857
R74958 VSS.n3986 VSS.n618 0.00962857
R74959 VSS.n3987 VSS.n3986 0.00962857
R74960 VSS.n3988 VSS.n3987 0.00962857
R74961 VSS.n3988 VSS.n614 0.00962857
R74962 VSS.n3994 VSS.n614 0.00962857
R74963 VSS.n3995 VSS.n3994 0.00962857
R74964 VSS.n3996 VSS.n3995 0.00962857
R74965 VSS.n3996 VSS.n610 0.00962857
R74966 VSS.n4002 VSS.n610 0.00962857
R74967 VSS.n4003 VSS.n4002 0.00962857
R74968 VSS.n4004 VSS.n4003 0.00962857
R74969 VSS.n4004 VSS.n606 0.00962857
R74970 VSS.n4010 VSS.n606 0.00962857
R74971 VSS.n4011 VSS.n4010 0.00962857
R74972 VSS.n4012 VSS.n4011 0.00962857
R74973 VSS.n4019 VSS.n4018 0.00962857
R74974 VSS.n4020 VSS.n4019 0.00962857
R74975 VSS.n4020 VSS.n598 0.00962857
R74976 VSS.n4026 VSS.n598 0.00962857
R74977 VSS.n4027 VSS.n4026 0.00962857
R74978 VSS.n4028 VSS.n4027 0.00962857
R74979 VSS.n4028 VSS.n594 0.00962857
R74980 VSS.n4034 VSS.n594 0.00962857
R74981 VSS.n4035 VSS.n4034 0.00962857
R74982 VSS.n4036 VSS.n4035 0.00962857
R74983 VSS.n4036 VSS.n590 0.00962857
R74984 VSS.n4042 VSS.n590 0.00962857
R74985 VSS.n4043 VSS.n4042 0.00962857
R74986 VSS.n4044 VSS.n4043 0.00962857
R74987 VSS.n4044 VSS.n575 0.00962857
R74988 VSS.n4082 VSS.n4050 0.00962857
R74989 VSS.n4082 VSS.n4081 0.00962857
R74990 VSS.n4081 VSS.n4080 0.00962857
R74991 VSS.n4080 VSS.n4051 0.00962857
R74992 VSS.n4074 VSS.n4051 0.00962857
R74993 VSS.n4074 VSS.n4073 0.00962857
R74994 VSS.n4073 VSS.n4072 0.00962857
R74995 VSS.n4072 VSS.n4055 0.00962857
R74996 VSS.n4066 VSS.n4055 0.00962857
R74997 VSS.n4066 VSS.n4065 0.00962857
R74998 VSS.n4065 VSS.n4064 0.00962857
R74999 VSS.n4570 VSS.n4569 0.00962857
R75000 VSS.n4574 VSS.n4569 0.00962857
R75001 VSS.n4574 VSS.n4568 0.00962857
R75002 VSS.n4578 VSS.n4568 0.00962857
R75003 VSS.n4578 VSS.n4566 0.00962857
R75004 VSS.n4582 VSS.n4566 0.00962857
R75005 VSS.n4582 VSS.n4564 0.00962857
R75006 VSS.n4586 VSS.n4564 0.00962857
R75007 VSS.n4586 VSS.n4562 0.00962857
R75008 VSS.n4590 VSS.n4562 0.00962857
R75009 VSS.n4590 VSS.n4560 0.00962857
R75010 VSS.n4594 VSS.n4560 0.00962857
R75011 VSS.n4594 VSS.n4558 0.00962857
R75012 VSS.n4599 VSS.n4558 0.00962857
R75013 VSS.n4599 VSS.n4556 0.00962857
R75014 VSS.n4603 VSS.n4556 0.00962857
R75015 VSS.n4604 VSS.n4603 0.00962857
R75016 VSS.n4604 VSS.n4554 0.00962857
R75017 VSS.n4608 VSS.n4554 0.00962857
R75018 VSS.n4608 VSS.n4553 0.00962857
R75019 VSS.n4612 VSS.n4553 0.00962857
R75020 VSS.n4612 VSS.n4551 0.00962857
R75021 VSS.n4616 VSS.n4551 0.00962857
R75022 VSS.n4616 VSS.n4549 0.00962857
R75023 VSS.n4620 VSS.n4549 0.00962857
R75024 VSS.n4620 VSS.n4547 0.00962857
R75025 VSS.n4624 VSS.n4547 0.00962857
R75026 VSS.n4624 VSS.n4545 0.00962857
R75027 VSS.n4628 VSS.n4545 0.00962857
R75028 VSS.n4628 VSS.n4543 0.00962857
R75029 VSS.n4632 VSS.n4543 0.00962857
R75030 VSS.n4632 VSS.n4541 0.00962857
R75031 VSS.n4636 VSS.n4541 0.00962857
R75032 VSS.n4636 VSS.n4539 0.00962857
R75033 VSS.n4640 VSS.n4539 0.00962857
R75034 VSS.n4641 VSS.n4640 0.00962857
R75035 VSS.n4643 VSS.n4641 0.00962857
R75036 VSS.n4643 VSS.n4536 0.00962857
R75037 VSS.n4647 VSS.n4536 0.00962857
R75038 VSS.n4647 VSS.n4534 0.00962857
R75039 VSS.n4651 VSS.n4534 0.00962857
R75040 VSS.n4651 VSS.n4532 0.00962857
R75041 VSS.n4655 VSS.n4532 0.00962857
R75042 VSS.n4655 VSS.n4530 0.00962857
R75043 VSS.n4659 VSS.n4530 0.00962857
R75044 VSS.n4659 VSS.n4528 0.00962857
R75045 VSS.n4663 VSS.n4528 0.00962857
R75046 VSS.n4663 VSS.n4526 0.00962857
R75047 VSS.n4667 VSS.n4526 0.00962857
R75048 VSS.n4667 VSS.n4523 0.00962857
R75049 VSS.n4759 VSS.n4523 0.00962857
R75050 VSS.n4759 VSS.n4524 0.00962857
R75051 VSS.n4755 VSS.n4524 0.00962857
R75052 VSS.n4755 VSS.n4754 0.00962857
R75053 VSS.n4754 VSS.n4671 0.00962857
R75054 VSS.n4750 VSS.n4671 0.00962857
R75055 VSS.n4750 VSS.n4673 0.00962857
R75056 VSS.n4746 VSS.n4673 0.00962857
R75057 VSS.n4746 VSS.n4676 0.00962857
R75058 VSS.n4742 VSS.n4676 0.00962857
R75059 VSS.n4742 VSS.n4678 0.00962857
R75060 VSS.n4738 VSS.n4678 0.00962857
R75061 VSS.n4738 VSS.n4680 0.00962857
R75062 VSS.n4734 VSS.n4680 0.00962857
R75063 VSS.n4734 VSS.n4682 0.00962857
R75064 VSS.n4730 VSS.n4682 0.00962857
R75065 VSS.n4730 VSS.n4684 0.00962857
R75066 VSS.n4726 VSS.n4684 0.00962857
R75067 VSS.n4726 VSS.n4685 0.00962857
R75068 VSS.n4722 VSS.n4685 0.00962857
R75069 VSS.n4722 VSS.n4721 0.00962857
R75070 VSS.n4721 VSS.n4687 0.00962857
R75071 VSS.n4717 VSS.n4687 0.00962857
R75072 VSS.n4717 VSS.n4689 0.00962857
R75073 VSS.n4713 VSS.n4689 0.00962857
R75074 VSS.n4713 VSS.n4692 0.00962857
R75075 VSS.n4709 VSS.n4692 0.00962857
R75076 VSS.n4709 VSS.n4694 0.00962857
R75077 VSS.n4705 VSS.n4694 0.00962857
R75078 VSS.n4705 VSS.n4696 0.00962857
R75079 VSS.n4701 VSS.n4696 0.00962857
R75080 VSS.n4575 VSS.n4255 0.00962857
R75081 VSS.n4576 VSS.n4575 0.00962857
R75082 VSS.n4577 VSS.n4576 0.00962857
R75083 VSS.n4577 VSS.n4565 0.00962857
R75084 VSS.n4583 VSS.n4565 0.00962857
R75085 VSS.n4584 VSS.n4583 0.00962857
R75086 VSS.n4585 VSS.n4584 0.00962857
R75087 VSS.n4585 VSS.n4561 0.00962857
R75088 VSS.n4591 VSS.n4561 0.00962857
R75089 VSS.n4592 VSS.n4591 0.00962857
R75090 VSS.n4593 VSS.n4592 0.00962857
R75091 VSS.n4593 VSS.n4557 0.00962857
R75092 VSS.n4600 VSS.n4557 0.00962857
R75093 VSS.n4601 VSS.n4600 0.00962857
R75094 VSS.n4602 VSS.n4601 0.00962857
R75095 VSS.n4609 VSS.n4273 0.00962857
R75096 VSS.n4610 VSS.n4609 0.00962857
R75097 VSS.n4611 VSS.n4610 0.00962857
R75098 VSS.n4611 VSS.n4550 0.00962857
R75099 VSS.n4617 VSS.n4550 0.00962857
R75100 VSS.n4618 VSS.n4617 0.00962857
R75101 VSS.n4619 VSS.n4618 0.00962857
R75102 VSS.n4619 VSS.n4546 0.00962857
R75103 VSS.n4625 VSS.n4546 0.00962857
R75104 VSS.n4626 VSS.n4625 0.00962857
R75105 VSS.n4627 VSS.n4626 0.00962857
R75106 VSS.n4627 VSS.n4542 0.00962857
R75107 VSS.n4633 VSS.n4542 0.00962857
R75108 VSS.n4634 VSS.n4633 0.00962857
R75109 VSS.n4635 VSS.n4634 0.00962857
R75110 VSS.n4642 VSS.n4496 0.00962857
R75111 VSS.n4642 VSS.n4535 0.00962857
R75112 VSS.n4648 VSS.n4535 0.00962857
R75113 VSS.n4649 VSS.n4648 0.00962857
R75114 VSS.n4650 VSS.n4649 0.00962857
R75115 VSS.n4650 VSS.n4531 0.00962857
R75116 VSS.n4656 VSS.n4531 0.00962857
R75117 VSS.n4657 VSS.n4656 0.00962857
R75118 VSS.n4658 VSS.n4657 0.00962857
R75119 VSS.n4658 VSS.n4527 0.00962857
R75120 VSS.n4664 VSS.n4527 0.00962857
R75121 VSS.n4665 VSS.n4664 0.00962857
R75122 VSS.n4666 VSS.n4665 0.00962857
R75123 VSS.n4666 VSS.n4522 0.00962857
R75124 VSS.n4760 VSS.n4522 0.00962857
R75125 VSS.n4753 VSS.n4518 0.00962857
R75126 VSS.n4753 VSS.n4752 0.00962857
R75127 VSS.n4752 VSS.n4751 0.00962857
R75128 VSS.n4751 VSS.n4672 0.00962857
R75129 VSS.n4745 VSS.n4672 0.00962857
R75130 VSS.n4745 VSS.n4744 0.00962857
R75131 VSS.n4744 VSS.n4743 0.00962857
R75132 VSS.n4743 VSS.n4677 0.00962857
R75133 VSS.n4737 VSS.n4677 0.00962857
R75134 VSS.n4737 VSS.n4736 0.00962857
R75135 VSS.n4736 VSS.n4735 0.00962857
R75136 VSS.n4735 VSS.n4681 0.00962857
R75137 VSS.n4729 VSS.n4681 0.00962857
R75138 VSS.n4729 VSS.n4728 0.00962857
R75139 VSS.n4728 VSS.n4727 0.00962857
R75140 VSS.n4720 VSS.n498 0.00962857
R75141 VSS.n4720 VSS.n4719 0.00962857
R75142 VSS.n4719 VSS.n4718 0.00962857
R75143 VSS.n4718 VSS.n4688 0.00962857
R75144 VSS.n4712 VSS.n4688 0.00962857
R75145 VSS.n4712 VSS.n4711 0.00962857
R75146 VSS.n4711 VSS.n4710 0.00962857
R75147 VSS.n4710 VSS.n4693 0.00962857
R75148 VSS.n4704 VSS.n4693 0.00962857
R75149 VSS.n4704 VSS.n4703 0.00962857
R75150 VSS.n4703 VSS.n4702 0.00962857
R75151 VSS.n6442 VSS.n22 0.00962857
R75152 VSS.n6442 VSS.n24 0.00962857
R75153 VSS.n6438 VSS.n24 0.00962857
R75154 VSS.n6438 VSS.n26 0.00962857
R75155 VSS.n6434 VSS.n26 0.00962857
R75156 VSS.n6434 VSS.n28 0.00962857
R75157 VSS.n6430 VSS.n28 0.00962857
R75158 VSS.n6430 VSS.n30 0.00962857
R75159 VSS.n6426 VSS.n30 0.00962857
R75160 VSS.n6426 VSS.n32 0.00962857
R75161 VSS.n6422 VSS.n32 0.00962857
R75162 VSS.n6422 VSS.n34 0.00962857
R75163 VSS.n6418 VSS.n34 0.00962857
R75164 VSS.n6418 VSS.n36 0.00962857
R75165 VSS.n6414 VSS.n36 0.00962857
R75166 VSS.n6414 VSS.n38 0.00962857
R75167 VSS.n6410 VSS.n38 0.00962857
R75168 VSS.n6410 VSS.n40 0.00962857
R75169 VSS.n6406 VSS.n40 0.00962857
R75170 VSS.n6406 VSS.n42 0.00962857
R75171 VSS.n6402 VSS.n42 0.00962857
R75172 VSS.n6402 VSS.n44 0.00962857
R75173 VSS.n6398 VSS.n44 0.00962857
R75174 VSS.n6398 VSS.n46 0.00962857
R75175 VSS.n6394 VSS.n46 0.00962857
R75176 VSS.n6394 VSS.n48 0.00962857
R75177 VSS.n6390 VSS.n48 0.00962857
R75178 VSS.n6390 VSS.n50 0.00962857
R75179 VSS.n6386 VSS.n50 0.00962857
R75180 VSS.n6386 VSS.n52 0.00962857
R75181 VSS.n6382 VSS.n52 0.00962857
R75182 VSS.n6382 VSS.n54 0.00962857
R75183 VSS.n6378 VSS.n54 0.00962857
R75184 VSS.n6378 VSS.n56 0.00962857
R75185 VSS.n6374 VSS.n56 0.00962857
R75186 VSS.n6374 VSS.n58 0.00962857
R75187 VSS.n6370 VSS.n58 0.00962857
R75188 VSS.n6370 VSS.n60 0.00962857
R75189 VSS.n6366 VSS.n60 0.00962857
R75190 VSS.n6366 VSS.n62 0.00962857
R75191 VSS.n6362 VSS.n62 0.00962857
R75192 VSS.n6362 VSS.n64 0.00962857
R75193 VSS.n6358 VSS.n64 0.00962857
R75194 VSS.n6358 VSS.n66 0.00962857
R75195 VSS.n6354 VSS.n66 0.00962857
R75196 VSS.n6354 VSS.n68 0.00962857
R75197 VSS.n6350 VSS.n68 0.00962857
R75198 VSS.n6350 VSS.n70 0.00962857
R75199 VSS.n6346 VSS.n70 0.00962857
R75200 VSS.n6346 VSS.n72 0.00962857
R75201 VSS.n6342 VSS.n72 0.00962857
R75202 VSS.n6342 VSS.n74 0.00962857
R75203 VSS.n6338 VSS.n74 0.00962857
R75204 VSS.n6338 VSS.n76 0.00962857
R75205 VSS.n6334 VSS.n76 0.00962857
R75206 VSS.n6334 VSS.n78 0.00962857
R75207 VSS.n6330 VSS.n78 0.00962857
R75208 VSS.n6330 VSS.n80 0.00962857
R75209 VSS.n6326 VSS.n80 0.00962857
R75210 VSS.n6326 VSS.n82 0.00962857
R75211 VSS.n6322 VSS.n82 0.00962857
R75212 VSS.n6322 VSS.n84 0.00962857
R75213 VSS.n6318 VSS.n84 0.00962857
R75214 VSS.n6318 VSS.n86 0.00962857
R75215 VSS.n6314 VSS.n86 0.00962857
R75216 VSS.n6314 VSS.n88 0.00962857
R75217 VSS.n6310 VSS.n88 0.00962857
R75218 VSS.n6310 VSS.n90 0.00962857
R75219 VSS.n6306 VSS.n90 0.00962857
R75220 VSS.n6306 VSS.n92 0.00962857
R75221 VSS.n6302 VSS.n92 0.00962857
R75222 VSS.n6302 VSS.n94 0.00962857
R75223 VSS.n6298 VSS.n94 0.00962857
R75224 VSS.n6298 VSS.n96 0.00962857
R75225 VSS.n6294 VSS.n96 0.00962857
R75226 VSS.n6294 VSS.n98 0.00962857
R75227 VSS.n6290 VSS.n98 0.00962857
R75228 VSS.n6290 VSS.n100 0.00962857
R75229 VSS.n6286 VSS.n100 0.00962857
R75230 VSS.n6286 VSS.n102 0.00962857
R75231 VSS.n6282 VSS.n102 0.00962857
R75232 VSS.n6282 VSS.n104 0.00962857
R75233 VSS.n6278 VSS.n104 0.00962857
R75234 VSS.n6278 VSS.n106 0.00962857
R75235 VSS.n6274 VSS.n106 0.00962857
R75236 VSS.n6274 VSS.n108 0.00962857
R75237 VSS.n6269 VSS.n108 0.00962857
R75238 VSS.n6269 VSS.n111 0.00962857
R75239 VSS.n6265 VSS.n111 0.00962857
R75240 VSS.n6265 VSS.n113 0.00962857
R75241 VSS.n6261 VSS.n113 0.00962857
R75242 VSS.n6261 VSS.n115 0.00962857
R75243 VSS.n6257 VSS.n115 0.00962857
R75244 VSS.n6257 VSS.n117 0.00962857
R75245 VSS.n6253 VSS.n117 0.00962857
R75246 VSS.n6253 VSS.n119 0.00962857
R75247 VSS.n6249 VSS.n119 0.00962857
R75248 VSS.n6246 VSS.n6245 0.00962857
R75249 VSS.n6245 VSS.n122 0.00962857
R75250 VSS.n6241 VSS.n122 0.00962857
R75251 VSS.n6445 VSS.n21 0.00962857
R75252 VSS.n6441 VSS.n21 0.00962857
R75253 VSS.n6441 VSS.n6440 0.00962857
R75254 VSS.n6440 VSS.n6439 0.00962857
R75255 VSS.n6439 VSS.n25 0.00962857
R75256 VSS.n6433 VSS.n25 0.00962857
R75257 VSS.n6433 VSS.n6432 0.00962857
R75258 VSS.n6432 VSS.n6431 0.00962857
R75259 VSS.n6431 VSS.n29 0.00962857
R75260 VSS.n6425 VSS.n29 0.00962857
R75261 VSS.n6425 VSS.n6424 0.00962857
R75262 VSS.n6424 VSS.n6423 0.00962857
R75263 VSS.n6423 VSS.n33 0.00962857
R75264 VSS.n6417 VSS.n33 0.00962857
R75265 VSS.n6417 VSS.n6416 0.00962857
R75266 VSS.n6416 VSS.n6415 0.00962857
R75267 VSS.n6415 VSS.n37 0.00962857
R75268 VSS.n6409 VSS.n37 0.00962857
R75269 VSS.n6409 VSS.n6408 0.00962857
R75270 VSS.n6408 VSS.n6407 0.00962857
R75271 VSS.n6407 VSS.n41 0.00962857
R75272 VSS.n6401 VSS.n41 0.00962857
R75273 VSS.n6401 VSS.n6400 0.00962857
R75274 VSS.n6400 VSS.n6399 0.00962857
R75275 VSS.n6399 VSS.n45 0.00962857
R75276 VSS.n6393 VSS.n45 0.00962857
R75277 VSS.n6393 VSS.n6392 0.00962857
R75278 VSS.n6392 VSS.n6391 0.00962857
R75279 VSS.n6391 VSS.n49 0.00962857
R75280 VSS.n6385 VSS.n49 0.00962857
R75281 VSS.n6385 VSS.n6384 0.00962857
R75282 VSS.n6384 VSS.n6383 0.00962857
R75283 VSS.n6383 VSS.n53 0.00962857
R75284 VSS.n6377 VSS.n53 0.00962857
R75285 VSS.n6377 VSS.n6376 0.00962857
R75286 VSS.n6376 VSS.n6375 0.00962857
R75287 VSS.n6375 VSS.n57 0.00962857
R75288 VSS.n6369 VSS.n57 0.00962857
R75289 VSS.n6369 VSS.n6368 0.00962857
R75290 VSS.n6368 VSS.n6367 0.00962857
R75291 VSS.n6367 VSS.n61 0.00962857
R75292 VSS.n6361 VSS.n61 0.00962857
R75293 VSS.n6361 VSS.n6360 0.00962857
R75294 VSS.n6360 VSS.n6359 0.00962857
R75295 VSS.n6359 VSS.n65 0.00962857
R75296 VSS.n6353 VSS.n65 0.00962857
R75297 VSS.n6353 VSS.n6352 0.00962857
R75298 VSS.n6352 VSS.n6351 0.00962857
R75299 VSS.n6351 VSS.n69 0.00962857
R75300 VSS.n6345 VSS.n69 0.00962857
R75301 VSS.n6345 VSS.n6344 0.00962857
R75302 VSS.n6344 VSS.n6343 0.00962857
R75303 VSS.n6343 VSS.n73 0.00962857
R75304 VSS.n6337 VSS.n73 0.00962857
R75305 VSS.n6337 VSS.n6336 0.00962857
R75306 VSS.n6336 VSS.n6335 0.00962857
R75307 VSS.n6335 VSS.n77 0.00962857
R75308 VSS.n6329 VSS.n77 0.00962857
R75309 VSS.n6329 VSS.n6328 0.00962857
R75310 VSS.n6328 VSS.n6327 0.00962857
R75311 VSS.n6327 VSS.n81 0.00962857
R75312 VSS.n6321 VSS.n81 0.00962857
R75313 VSS.n6321 VSS.n6320 0.00962857
R75314 VSS.n6320 VSS.n6319 0.00962857
R75315 VSS.n6319 VSS.n85 0.00962857
R75316 VSS.n6313 VSS.n85 0.00962857
R75317 VSS.n6313 VSS.n6312 0.00962857
R75318 VSS.n6312 VSS.n6311 0.00962857
R75319 VSS.n6311 VSS.n89 0.00962857
R75320 VSS.n6305 VSS.n89 0.00962857
R75321 VSS.n6305 VSS.n6304 0.00962857
R75322 VSS.n6304 VSS.n6303 0.00962857
R75323 VSS.n6303 VSS.n93 0.00962857
R75324 VSS.n6297 VSS.n93 0.00962857
R75325 VSS.n6297 VSS.n6296 0.00962857
R75326 VSS.n6296 VSS.n6295 0.00962857
R75327 VSS.n6295 VSS.n97 0.00962857
R75328 VSS.n6289 VSS.n97 0.00962857
R75329 VSS.n6289 VSS.n6288 0.00962857
R75330 VSS.n6288 VSS.n6287 0.00962857
R75331 VSS.n6287 VSS.n101 0.00962857
R75332 VSS.n6281 VSS.n101 0.00962857
R75333 VSS.n6281 VSS.n6280 0.00962857
R75334 VSS.n6280 VSS.n6279 0.00962857
R75335 VSS.n6279 VSS.n105 0.00962857
R75336 VSS.n6273 VSS.n105 0.00962857
R75337 VSS.n6273 VSS.n6272 0.00962857
R75338 VSS.n6270 VSS.n110 0.00962857
R75339 VSS.n6264 VSS.n110 0.00962857
R75340 VSS.n6264 VSS.n6263 0.00962857
R75341 VSS.n6263 VSS.n6262 0.00962857
R75342 VSS.n6262 VSS.n114 0.00962857
R75343 VSS.n6256 VSS.n114 0.00962857
R75344 VSS.n6256 VSS.n6255 0.00962857
R75345 VSS.n6255 VSS.n6254 0.00962857
R75346 VSS.n6254 VSS.n118 0.00962857
R75347 VSS.n6248 VSS.n118 0.00962857
R75348 VSS.n6247 VSS.n121 0.00962857
R75349 VSS.n6239 VSS.n121 0.00962857
R75350 VSS.n6240 VSS.n6239 0.00962857
R75351 VSS.n6240 VSS.n6238 0.00962857
R75352 VSS.n437 VSS.n144 0.00962857
R75353 VSS.n433 VSS.n144 0.00962857
R75354 VSS.n433 VSS.n432 0.00962857
R75355 VSS.n432 VSS.n431 0.00962857
R75356 VSS.n431 VSS.n147 0.00962857
R75357 VSS.n425 VSS.n147 0.00962857
R75358 VSS.n425 VSS.n424 0.00962857
R75359 VSS.n424 VSS.n423 0.00962857
R75360 VSS.n423 VSS.n152 0.00962857
R75361 VSS.n417 VSS.n152 0.00962857
R75362 VSS.n417 VSS.n416 0.00962857
R75363 VSS.n416 VSS.n415 0.00962857
R75364 VSS.n415 VSS.n156 0.00962857
R75365 VSS.n409 VSS.n156 0.00962857
R75366 VSS.n409 VSS.n408 0.00962857
R75367 VSS.n408 VSS.n407 0.00962857
R75368 VSS.n407 VSS.n160 0.00962857
R75369 VSS.n401 VSS.n160 0.00962857
R75370 VSS.n401 VSS.n400 0.00962857
R75371 VSS.n400 VSS.n399 0.00962857
R75372 VSS.n399 VSS.n164 0.00962857
R75373 VSS.n393 VSS.n164 0.00962857
R75374 VSS.n393 VSS.n392 0.00962857
R75375 VSS.n392 VSS.n391 0.00962857
R75376 VSS.n391 VSS.n168 0.00962857
R75377 VSS.n385 VSS.n168 0.00962857
R75378 VSS.n385 VSS.n384 0.00962857
R75379 VSS.n384 VSS.n383 0.00962857
R75380 VSS.n383 VSS.n172 0.00962857
R75381 VSS.n377 VSS.n172 0.00962857
R75382 VSS.n377 VSS.n376 0.00962857
R75383 VSS.n376 VSS.n375 0.00962857
R75384 VSS.n375 VSS.n176 0.00962857
R75385 VSS.n369 VSS.n176 0.00962857
R75386 VSS.n369 VSS.n368 0.00962857
R75387 VSS.n368 VSS.n367 0.00962857
R75388 VSS.n367 VSS.n180 0.00962857
R75389 VSS.n361 VSS.n180 0.00962857
R75390 VSS.n361 VSS.n360 0.00962857
R75391 VSS.n360 VSS.n359 0.00962857
R75392 VSS.n359 VSS.n184 0.00962857
R75393 VSS.n353 VSS.n184 0.00962857
R75394 VSS.n353 VSS.n352 0.00962857
R75395 VSS.n352 VSS.n351 0.00962857
R75396 VSS.n351 VSS.n188 0.00962857
R75397 VSS.n345 VSS.n188 0.00962857
R75398 VSS.n345 VSS.n344 0.00962857
R75399 VSS.n344 VSS.n343 0.00962857
R75400 VSS.n343 VSS.n192 0.00962857
R75401 VSS.n337 VSS.n192 0.00962857
R75402 VSS.n337 VSS.n336 0.00962857
R75403 VSS.n336 VSS.n335 0.00962857
R75404 VSS.n335 VSS.n196 0.00962857
R75405 VSS.n329 VSS.n196 0.00962857
R75406 VSS.n329 VSS.n328 0.00962857
R75407 VSS.n328 VSS.n327 0.00962857
R75408 VSS.n327 VSS.n200 0.00962857
R75409 VSS.n321 VSS.n200 0.00962857
R75410 VSS.n321 VSS.n320 0.00962857
R75411 VSS.n320 VSS.n319 0.00962857
R75412 VSS.n319 VSS.n204 0.00962857
R75413 VSS.n313 VSS.n204 0.00962857
R75414 VSS.n313 VSS.n312 0.00962857
R75415 VSS.n312 VSS.n311 0.00962857
R75416 VSS.n311 VSS.n208 0.00962857
R75417 VSS.n305 VSS.n208 0.00962857
R75418 VSS.n305 VSS.n304 0.00962857
R75419 VSS.n304 VSS.n303 0.00962857
R75420 VSS.n303 VSS.n212 0.00962857
R75421 VSS.n297 VSS.n212 0.00962857
R75422 VSS.n297 VSS.n296 0.00962857
R75423 VSS.n296 VSS.n295 0.00962857
R75424 VSS.n295 VSS.n216 0.00962857
R75425 VSS.n289 VSS.n216 0.00962857
R75426 VSS.n289 VSS.n288 0.00962857
R75427 VSS.n288 VSS.n287 0.00962857
R75428 VSS.n287 VSS.n220 0.00962857
R75429 VSS.n281 VSS.n220 0.00962857
R75430 VSS.n281 VSS.n280 0.00962857
R75431 VSS.n280 VSS.n279 0.00962857
R75432 VSS.n279 VSS.n224 0.00962857
R75433 VSS.n273 VSS.n224 0.00962857
R75434 VSS.n273 VSS.n272 0.00962857
R75435 VSS.n272 VSS.n271 0.00962857
R75436 VSS.n271 VSS.n228 0.00962857
R75437 VSS.n265 VSS.n228 0.00962857
R75438 VSS.n265 VSS.n264 0.00962857
R75439 VSS.n261 VSS.n260 0.00962857
R75440 VSS.n260 VSS.n259 0.00962857
R75441 VSS.n259 VSS.n233 0.00962857
R75442 VSS.n253 VSS.n233 0.00962857
R75443 VSS.n253 VSS.n252 0.00962857
R75444 VSS.n252 VSS.n251 0.00962857
R75445 VSS.n251 VSS.n238 0.00962857
R75446 VSS.n245 VSS.n238 0.00962857
R75447 VSS.n245 VSS.n244 0.00962857
R75448 VSS.n244 VSS.n0 0.00962857
R75449 VSS.n6469 VSS.n1 0.00962857
R75450 VSS.n6463 VSS.n1 0.00962857
R75451 VSS.n6463 VSS.n6462 0.00962857
R75452 VSS.n6462 VSS.n6461 0.00962857
R75453 VSS.n435 VSS.n434 0.00962857
R75454 VSS.n434 VSS.n146 0.00962857
R75455 VSS.n430 VSS.n146 0.00962857
R75456 VSS.n430 VSS.n148 0.00962857
R75457 VSS.n426 VSS.n148 0.00962857
R75458 VSS.n426 VSS.n151 0.00962857
R75459 VSS.n422 VSS.n151 0.00962857
R75460 VSS.n422 VSS.n153 0.00962857
R75461 VSS.n418 VSS.n153 0.00962857
R75462 VSS.n418 VSS.n155 0.00962857
R75463 VSS.n414 VSS.n155 0.00962857
R75464 VSS.n414 VSS.n157 0.00962857
R75465 VSS.n410 VSS.n157 0.00962857
R75466 VSS.n410 VSS.n159 0.00962857
R75467 VSS.n406 VSS.n159 0.00962857
R75468 VSS.n406 VSS.n161 0.00962857
R75469 VSS.n402 VSS.n161 0.00962857
R75470 VSS.n402 VSS.n163 0.00962857
R75471 VSS.n398 VSS.n163 0.00962857
R75472 VSS.n398 VSS.n165 0.00962857
R75473 VSS.n394 VSS.n165 0.00962857
R75474 VSS.n394 VSS.n167 0.00962857
R75475 VSS.n390 VSS.n167 0.00962857
R75476 VSS.n390 VSS.n169 0.00962857
R75477 VSS.n386 VSS.n169 0.00962857
R75478 VSS.n386 VSS.n171 0.00962857
R75479 VSS.n382 VSS.n171 0.00962857
R75480 VSS.n382 VSS.n173 0.00962857
R75481 VSS.n378 VSS.n173 0.00962857
R75482 VSS.n378 VSS.n175 0.00962857
R75483 VSS.n374 VSS.n175 0.00962857
R75484 VSS.n374 VSS.n177 0.00962857
R75485 VSS.n370 VSS.n177 0.00962857
R75486 VSS.n370 VSS.n179 0.00962857
R75487 VSS.n366 VSS.n179 0.00962857
R75488 VSS.n366 VSS.n181 0.00962857
R75489 VSS.n362 VSS.n181 0.00962857
R75490 VSS.n362 VSS.n183 0.00962857
R75491 VSS.n358 VSS.n183 0.00962857
R75492 VSS.n358 VSS.n185 0.00962857
R75493 VSS.n354 VSS.n185 0.00962857
R75494 VSS.n354 VSS.n187 0.00962857
R75495 VSS.n350 VSS.n187 0.00962857
R75496 VSS.n350 VSS.n189 0.00962857
R75497 VSS.n346 VSS.n189 0.00962857
R75498 VSS.n346 VSS.n191 0.00962857
R75499 VSS.n342 VSS.n191 0.00962857
R75500 VSS.n342 VSS.n193 0.00962857
R75501 VSS.n338 VSS.n193 0.00962857
R75502 VSS.n338 VSS.n195 0.00962857
R75503 VSS.n334 VSS.n195 0.00962857
R75504 VSS.n334 VSS.n197 0.00962857
R75505 VSS.n330 VSS.n197 0.00962857
R75506 VSS.n330 VSS.n199 0.00962857
R75507 VSS.n326 VSS.n199 0.00962857
R75508 VSS.n326 VSS.n201 0.00962857
R75509 VSS.n322 VSS.n201 0.00962857
R75510 VSS.n322 VSS.n203 0.00962857
R75511 VSS.n318 VSS.n203 0.00962857
R75512 VSS.n318 VSS.n205 0.00962857
R75513 VSS.n314 VSS.n205 0.00962857
R75514 VSS.n314 VSS.n207 0.00962857
R75515 VSS.n310 VSS.n207 0.00962857
R75516 VSS.n310 VSS.n209 0.00962857
R75517 VSS.n306 VSS.n209 0.00962857
R75518 VSS.n306 VSS.n211 0.00962857
R75519 VSS.n302 VSS.n211 0.00962857
R75520 VSS.n302 VSS.n213 0.00962857
R75521 VSS.n298 VSS.n213 0.00962857
R75522 VSS.n298 VSS.n215 0.00962857
R75523 VSS.n294 VSS.n215 0.00962857
R75524 VSS.n294 VSS.n217 0.00962857
R75525 VSS.n290 VSS.n217 0.00962857
R75526 VSS.n290 VSS.n219 0.00962857
R75527 VSS.n286 VSS.n219 0.00962857
R75528 VSS.n286 VSS.n221 0.00962857
R75529 VSS.n282 VSS.n221 0.00962857
R75530 VSS.n282 VSS.n223 0.00962857
R75531 VSS.n278 VSS.n223 0.00962857
R75532 VSS.n278 VSS.n225 0.00962857
R75533 VSS.n274 VSS.n225 0.00962857
R75534 VSS.n274 VSS.n227 0.00962857
R75535 VSS.n270 VSS.n227 0.00962857
R75536 VSS.n270 VSS.n229 0.00962857
R75537 VSS.n266 VSS.n229 0.00962857
R75538 VSS.n266 VSS.n263 0.00962857
R75539 VSS.n263 VSS.n262 0.00962857
R75540 VSS.n262 VSS.n232 0.00962857
R75541 VSS.n258 VSS.n232 0.00962857
R75542 VSS.n258 VSS.n234 0.00962857
R75543 VSS.n254 VSS.n234 0.00962857
R75544 VSS.n254 VSS.n237 0.00962857
R75545 VSS.n250 VSS.n237 0.00962857
R75546 VSS.n250 VSS.n239 0.00962857
R75547 VSS.n246 VSS.n239 0.00962857
R75548 VSS.n246 VSS.n243 0.00962857
R75549 VSS.n243 VSS.n242 0.00962857
R75550 VSS.n6468 VSS.n2 0.00962857
R75551 VSS.n6464 VSS.n2 0.00962857
R75552 VSS.n6464 VSS.n4 0.00962857
R75553 VSS.n5018 VSS.n5017 0.00923134
R75554 VSS.n1751 VSS.n1282 0.00917857
R75555 VSS.n2987 VSS.n2986 0.00917857
R75556 VSS.n2780 VSS.n2779 0.00917857
R75557 VSS.n4012 VSS.n571 0.00917857
R75558 VSS.n4765 VSS.n4760 0.00917857
R75559 VSS.n6202 VSS.n6201 0.00910927
R75560 VSS.n6201 VSS.n6200 0.00910927
R75561 VSS.n6224 VSS.n6223 0.00910927
R75562 VSS.n6223 VSS.n6222 0.00910927
R75563 VSS.n6272 VSS.n6271 0.00905
R75564 VSS.n264 VSS.n109 0.00905
R75565 VSS.n1536 VSS.n1531 0.00892143
R75566 VSS.n1927 VSS.n1161 0.00892143
R75567 VSS.n2859 VSS.n2858 0.00892143
R75568 VSS.n3938 VSS.n3937 0.00892143
R75569 VSS.n6121 VSS.n4273 0.00892143
R75570 VSS.n3762 DVSS 0.0088427
R75571 VSS.n436 VSS.n435 0.00880017
R75572 VSS.n1663 VSS.n1306 0.00873944
R75573 VSS.n1746 VSS.n1284 0.00873944
R75574 VSS.n4833 VSS.n4832 0.0086
R75575 VSS.n5532 VSS.n4972 0.0086
R75576 VSS.n4824 VSS.n4822 0.0086
R75577 VSS.n5533 VSS.n5202 0.0086
R75578 VSS.n4826 VSS.n4296 0.0086
R75579 VSS.n5528 VSS.n5311 0.0086
R75580 VSS.n4827 VSS.n4312 0.0086
R75581 VSS.n5529 VSS.n5269 0.0086
R75582 DVSS VSS.n1856 0.00852817
R75583 VSS.n1861 DVSS 0.00852817
R75584 VSS.n2553 VSS.n2552 0.00846348
R75585 VSS.n3265 VSS.n844 0.00846348
R75586 VSS.n1617 VSS.n1546 0.00845775
R75587 VSS.n1659 VSS.n1325 0.00845775
R75588 DVSS VSS.n5923 0.00823835
R75589 VSS.n2548 VSS.n2226 0.00819509
R75590 VSS.n3276 VSS.n3271 0.00819509
R75591 VSS.n2231 VSS.n2226 0.00819509
R75592 VSS.n3279 VSS.n3271 0.00819509
R75593 DVSS VSS.n2648 0.00808427
R75594 VSS.n1496 VSS.n1433 0.00802143
R75595 VSS.n1754 VSS.n1274 0.00802143
R75596 VSS.n1107 VSS.n1104 0.00802143
R75597 VSS.n1084 VSS.n1077 0.00802143
R75598 VSS.n2824 VSS.n2747 0.00802143
R75599 VSS.n3436 VSS.n974 0.00802143
R75600 VSS.n3980 VSS.n3979 0.00802143
R75601 VSS.n602 VSS.n572 0.00802143
R75602 VSS.n4775 VSS.n4490 0.00802143
R75603 VSS.n4768 VSS.n4516 0.00802143
R75604 DVSS VSS.n727 0.00795787
R75605 VSS.n4774 VSS.n4773 0.00788806
R75606 VSS.n1799 DVSS 0.00782857
R75607 VSS.n1800 DVSS 0.00782857
R75608 VSS.n3038 DVSS 0.00782857
R75609 VSS.n3039 DVSS 0.00782857
R75610 DVSS VSS.n1017 0.00782857
R75611 VSS.n1021 DVSS 0.00782857
R75612 VSS.n4063 DVSS 0.00782857
R75613 VSS.n4064 DVSS 0.00782857
R75614 VSS.n4701 DVSS 0.00782857
R75615 VSS.n4702 DVSS 0.00782857
R75616 VSS.n6249 VSS 0.00782857
R75617 VSS.n6248 VSS 0.00782857
R75618 VSS VSS.n0 0.00782857
R75619 VSS.n242 VSS 0.00782857
R75620 VSS.n1356 VSS.n1355 0.00776429
R75621 VSS.n1499 VSS.n1426 0.00776429
R75622 VSS.n2020 VSS.n1160 0.00776429
R75623 VSS.n1940 VSS.n1116 0.00776429
R75624 VSS.n1164 VSS.n1163 0.00776429
R75625 VSS.n2826 VSS.n2743 0.00776429
R75626 VSS.n3934 VSS.n654 0.00776429
R75627 VSS.n3975 VSS.n3974 0.00776429
R75628 VSS.n4270 VSS.n4268 0.00776429
R75629 VSS.n4538 VSS.n4488 0.00776429
R75630 VSS.n3691 VSS.n3690 0.00772462
R75631 VSS.n5962 VSS.n5961 0.00772462
R75632 VSS.n5887 VSS.n5886 0.00772462
R75633 VSS.n2977 VSS.n2976 0.00772015
R75634 VSS.n2980 VSS.n1097 0.00772015
R75635 VSS.n1430 VSS.n1217 0.00755224
R75636 VSS.n2649 DVSS 0.00732584
R75637 VSS.n734 VSS.n733 0.00732584
R75638 VSS.n1554 VSS.n1553 0.00716667
R75639 VSS.n1555 VSS.n1554 0.00716667
R75640 VSS.n1558 VSS.n1555 0.00716667
R75641 VSS.n1559 VSS.n1558 0.00716667
R75642 VSS.n1560 VSS.n1559 0.00716667
R75643 VSS.n1561 VSS.n1560 0.00716667
R75644 VSS.n1564 VSS.n1561 0.00716667
R75645 VSS.n1565 VSS.n1564 0.00716667
R75646 VSS.n1566 VSS.n1565 0.00716667
R75647 VSS.n1567 VSS.n1566 0.00716667
R75648 VSS.n1570 VSS.n1567 0.00716667
R75649 VSS.n1571 VSS.n1570 0.00716667
R75650 VSS.n1572 VSS.n1571 0.00716667
R75651 VSS.n1572 VSS.n1344 0.00716667
R75652 VSS.n1620 VSS.n1344 0.00716667
R75653 VSS.n1621 VSS.n1620 0.00716667
R75654 VSS.n1622 VSS.n1621 0.00716667
R75655 VSS.n1622 VSS.n1340 0.00716667
R75656 VSS.n1628 VSS.n1340 0.00716667
R75657 VSS.n1629 VSS.n1628 0.00716667
R75658 VSS.n1630 VSS.n1629 0.00716667
R75659 VSS.n1630 VSS.n1336 0.00716667
R75660 VSS.n1636 VSS.n1336 0.00716667
R75661 VSS.n1637 VSS.n1636 0.00716667
R75662 VSS.n1638 VSS.n1637 0.00716667
R75663 VSS.n1638 VSS.n1332 0.00716667
R75664 VSS.n1644 VSS.n1332 0.00716667
R75665 VSS.n1645 VSS.n1644 0.00716667
R75666 VSS.n1646 VSS.n1645 0.00716667
R75667 VSS.n1646 VSS.n1328 0.00716667
R75668 VSS.n1653 VSS.n1328 0.00716667
R75669 VSS.n1654 VSS.n1653 0.00716667
R75670 VSS.n1655 VSS.n1654 0.00716667
R75671 VSS.n1656 VSS.n1655 0.00716667
R75672 VSS.n1656 VSS.n1304 0.00716667
R75673 VSS.n1667 VSS.n1304 0.00716667
R75674 VSS.n1668 VSS.n1667 0.00716667
R75675 VSS.n1669 VSS.n1668 0.00716667
R75676 VSS.n1669 VSS.n1300 0.00716667
R75677 VSS.n1675 VSS.n1300 0.00716667
R75678 VSS.n1676 VSS.n1675 0.00716667
R75679 VSS.n1677 VSS.n1676 0.00716667
R75680 VSS.n1677 VSS.n1296 0.00716667
R75681 VSS.n1683 VSS.n1296 0.00716667
R75682 VSS.n1684 VSS.n1683 0.00716667
R75683 VSS.n1685 VSS.n1684 0.00716667
R75684 VSS.n1685 VSS.n1292 0.00716667
R75685 VSS.n1691 VSS.n1292 0.00716667
R75686 VSS.n1692 VSS.n1691 0.00716667
R75687 VSS.n1693 VSS.n1692 0.00716667
R75688 VSS.n1694 VSS.n1693 0.00716667
R75689 VSS.n1695 VSS.n1694 0.00716667
R75690 VSS.n1696 VSS.n1695 0.00716667
R75691 VSS.n1699 VSS.n1696 0.00716667
R75692 VSS.n1700 VSS.n1699 0.00716667
R75693 VSS.n1701 VSS.n1700 0.00716667
R75694 VSS.n1702 VSS.n1701 0.00716667
R75695 VSS.n1705 VSS.n1702 0.00716667
R75696 VSS.n1706 VSS.n1705 0.00716667
R75697 VSS.n1707 VSS.n1706 0.00716667
R75698 VSS.n1708 VSS.n1707 0.00716667
R75699 VSS.n1711 VSS.n1708 0.00716667
R75700 VSS.n1712 VSS.n1711 0.00716667
R75701 VSS.n1713 VSS.n1712 0.00716667
R75702 VSS.n1714 VSS.n1713 0.00716667
R75703 VSS.n1714 VSS.n1243 0.00716667
R75704 VSS.n1839 VSS.n1243 0.00716667
R75705 VSS.n1840 VSS.n1839 0.00716667
R75706 VSS.n1841 VSS.n1840 0.00716667
R75707 VSS.n1842 VSS.n1841 0.00716667
R75708 VSS.n1843 VSS.n1842 0.00716667
R75709 VSS.n1846 VSS.n1843 0.00716667
R75710 VSS.n1847 VSS.n1846 0.00716667
R75711 VSS.n1848 VSS.n1847 0.00716667
R75712 VSS.n1849 VSS.n1848 0.00716667
R75713 VSS.n1852 VSS.n1849 0.00716667
R75714 VSS.n1853 VSS.n1852 0.00716667
R75715 VSS.n1854 VSS.n1853 0.00716667
R75716 VSS.n1855 VSS.n1854 0.00716667
R75717 VSS.n1857 VSS.n1855 0.00716667
R75718 VSS.n2552 VSS.n2551 0.00694663
R75719 VSS.n3266 VSS.n3265 0.00694663
R75720 VSS.n1837 VSS.n1836 0.00690845
R75721 VSS.n6453 VSS.n6452 0.00684146
R75722 VSS.n5853 VSS.n4964 0.0068
R75723 VSS.n5095 VSS.n4925 0.0068
R75724 VSS.n5644 VSS.n5194 0.0068
R75725 VSS.n5096 VSS.n5061 0.0068
R75726 VSS.n5620 VSS.n5304 0.0068
R75727 VSS.n5103 VSS.n5089 0.0068
R75728 VSS.n5273 VSS.n5262 0.0068
R75729 VSS.n5101 VSS.n5004 0.0068
R75730 VSS.n1594 VSS.n1593 0.00662676
R75731 VSS.n149 VSS.n145 0.00658571
R75732 VSS.n429 VSS.n149 0.00658571
R75733 VSS.n429 VSS.n428 0.00658571
R75734 VSS.n428 VSS.n427 0.00658571
R75735 VSS.n427 VSS.n150 0.00658571
R75736 VSS.n421 VSS.n150 0.00658571
R75737 VSS.n421 VSS.n420 0.00658571
R75738 VSS.n420 VSS.n419 0.00658571
R75739 VSS.n419 VSS.n154 0.00658571
R75740 VSS.n413 VSS.n154 0.00658571
R75741 VSS.n413 VSS.n412 0.00658571
R75742 VSS.n412 VSS.n411 0.00658571
R75743 VSS.n411 VSS.n158 0.00658571
R75744 VSS.n405 VSS.n158 0.00658571
R75745 VSS.n405 VSS.n404 0.00658571
R75746 VSS.n404 VSS.n403 0.00658571
R75747 VSS.n403 VSS.n162 0.00658571
R75748 VSS.n397 VSS.n162 0.00658571
R75749 VSS.n397 VSS.n396 0.00658571
R75750 VSS.n396 VSS.n395 0.00658571
R75751 VSS.n395 VSS.n166 0.00658571
R75752 VSS.n389 VSS.n166 0.00658571
R75753 VSS.n389 VSS.n388 0.00658571
R75754 VSS.n388 VSS.n387 0.00658571
R75755 VSS.n387 VSS.n170 0.00658571
R75756 VSS.n381 VSS.n170 0.00658571
R75757 VSS.n381 VSS.n380 0.00658571
R75758 VSS.n380 VSS.n379 0.00658571
R75759 VSS.n379 VSS.n174 0.00658571
R75760 VSS.n373 VSS.n174 0.00658571
R75761 VSS.n373 VSS.n372 0.00658571
R75762 VSS.n372 VSS.n371 0.00658571
R75763 VSS.n371 VSS.n178 0.00658571
R75764 VSS.n365 VSS.n178 0.00658571
R75765 VSS.n365 VSS.n364 0.00658571
R75766 VSS.n364 VSS.n363 0.00658571
R75767 VSS.n363 VSS.n182 0.00658571
R75768 VSS.n357 VSS.n182 0.00658571
R75769 VSS.n357 VSS.n356 0.00658571
R75770 VSS.n356 VSS.n355 0.00658571
R75771 VSS.n355 VSS.n186 0.00658571
R75772 VSS.n349 VSS.n186 0.00658571
R75773 VSS.n349 VSS.n348 0.00658571
R75774 VSS.n348 VSS.n347 0.00658571
R75775 VSS.n347 VSS.n190 0.00658571
R75776 VSS.n341 VSS.n190 0.00658571
R75777 VSS.n341 VSS.n340 0.00658571
R75778 VSS.n340 VSS.n339 0.00658571
R75779 VSS.n339 VSS.n194 0.00658571
R75780 VSS.n333 VSS.n194 0.00658571
R75781 VSS.n333 VSS.n332 0.00658571
R75782 VSS.n332 VSS.n331 0.00658571
R75783 VSS.n331 VSS.n198 0.00658571
R75784 VSS.n325 VSS.n198 0.00658571
R75785 VSS.n325 VSS.n324 0.00658571
R75786 VSS.n324 VSS.n323 0.00658571
R75787 VSS.n323 VSS.n202 0.00658571
R75788 VSS.n317 VSS.n202 0.00658571
R75789 VSS.n317 VSS.n316 0.00658571
R75790 VSS.n316 VSS.n315 0.00658571
R75791 VSS.n315 VSS.n206 0.00658571
R75792 VSS.n309 VSS.n206 0.00658571
R75793 VSS.n309 VSS.n308 0.00658571
R75794 VSS.n308 VSS.n307 0.00658571
R75795 VSS.n307 VSS.n210 0.00658571
R75796 VSS.n301 VSS.n210 0.00658571
R75797 VSS.n301 VSS.n300 0.00658571
R75798 VSS.n300 VSS.n299 0.00658571
R75799 VSS.n299 VSS.n214 0.00658571
R75800 VSS.n293 VSS.n214 0.00658571
R75801 VSS.n293 VSS.n292 0.00658571
R75802 VSS.n292 VSS.n291 0.00658571
R75803 VSS.n291 VSS.n218 0.00658571
R75804 VSS.n285 VSS.n218 0.00658571
R75805 VSS.n285 VSS.n284 0.00658571
R75806 VSS.n284 VSS.n283 0.00658571
R75807 VSS.n283 VSS.n222 0.00658571
R75808 VSS.n277 VSS.n222 0.00658571
R75809 VSS.n277 VSS.n276 0.00658571
R75810 VSS.n276 VSS.n275 0.00658571
R75811 VSS.n275 VSS.n226 0.00658571
R75812 VSS.n269 VSS.n226 0.00658571
R75813 VSS.n269 VSS.n268 0.00658571
R75814 VSS.n268 VSS.n267 0.00658571
R75815 VSS.n267 VSS.n230 0.00658571
R75816 VSS.n231 VSS.n230 0.00658571
R75817 VSS.n235 VSS.n231 0.00658571
R75818 VSS.n257 VSS.n235 0.00658571
R75819 VSS.n257 VSS.n256 0.00658571
R75820 VSS.n256 VSS.n255 0.00658571
R75821 VSS.n255 VSS.n236 0.00658571
R75822 VSS.n249 VSS.n236 0.00658571
R75823 VSS.n249 VSS.n248 0.00658571
R75824 VSS.n248 VSS.n247 0.00658571
R75825 VSS.n247 VSS.n240 0.00658571
R75826 VSS.n241 VSS.n240 0.00658571
R75827 VSS.n6466 VSS.n6465 0.00658571
R75828 VSS.n1378 VSS.n1377 0.00658571
R75829 VSS.n1378 VSS.n1373 0.00658571
R75830 VSS.n1384 VSS.n1373 0.00658571
R75831 VSS.n1385 VSS.n1384 0.00658571
R75832 VSS.n1386 VSS.n1385 0.00658571
R75833 VSS.n1386 VSS.n1369 0.00658571
R75834 VSS.n1392 VSS.n1369 0.00658571
R75835 VSS.n1393 VSS.n1392 0.00658571
R75836 VSS.n1394 VSS.n1393 0.00658571
R75837 VSS.n1394 VSS.n1365 0.00658571
R75838 VSS.n1400 VSS.n1365 0.00658571
R75839 VSS.n1401 VSS.n1400 0.00658571
R75840 VSS.n1402 VSS.n1401 0.00658571
R75841 VSS.n1402 VSS.n1361 0.00658571
R75842 VSS.n1408 VSS.n1361 0.00658571
R75843 VSS.n1409 VSS.n1408 0.00658571
R75844 VSS.n1529 VSS.n1409 0.00658571
R75845 VSS.n1529 VSS.n1528 0.00658571
R75846 VSS.n1528 VSS.n1527 0.00658571
R75847 VSS.n1527 VSS.n1410 0.00658571
R75848 VSS.n1521 VSS.n1410 0.00658571
R75849 VSS.n1521 VSS.n1520 0.00658571
R75850 VSS.n1520 VSS.n1519 0.00658571
R75851 VSS.n1519 VSS.n1414 0.00658571
R75852 VSS.n1513 VSS.n1414 0.00658571
R75853 VSS.n1513 VSS.n1512 0.00658571
R75854 VSS.n1512 VSS.n1511 0.00658571
R75855 VSS.n1511 VSS.n1418 0.00658571
R75856 VSS.n1505 VSS.n1418 0.00658571
R75857 VSS.n1505 VSS.n1504 0.00658571
R75858 VSS.n1504 VSS.n1503 0.00658571
R75859 VSS.n1503 VSS.n1422 0.00658571
R75860 VSS.n1441 VSS.n1422 0.00658571
R75861 VSS.n1442 VSS.n1441 0.00658571
R75862 VSS.n1487 VSS.n1442 0.00658571
R75863 VSS.n1487 VSS.n1486 0.00658571
R75864 VSS.n1486 VSS.n1485 0.00658571
R75865 VSS.n1485 VSS.n1443 0.00658571
R75866 VSS.n1479 VSS.n1443 0.00658571
R75867 VSS.n1479 VSS.n1478 0.00658571
R75868 VSS.n1478 VSS.n1477 0.00658571
R75869 VSS.n1477 VSS.n1447 0.00658571
R75870 VSS.n1471 VSS.n1447 0.00658571
R75871 VSS.n1471 VSS.n1470 0.00658571
R75872 VSS.n1470 VSS.n1469 0.00658571
R75873 VSS.n1469 VSS.n1451 0.00658571
R75874 VSS.n1463 VSS.n1451 0.00658571
R75875 VSS.n1463 VSS.n1462 0.00658571
R75876 VSS.n1462 VSS.n1461 0.00658571
R75877 VSS.n1461 VSS.n1455 0.00658571
R75878 VSS.n1456 VSS.n1455 0.00658571
R75879 VSS.n1456 VSS.n1272 0.00658571
R75880 VSS.n1758 VSS.n1272 0.00658571
R75881 VSS.n1759 VSS.n1758 0.00658571
R75882 VSS.n1760 VSS.n1759 0.00658571
R75883 VSS.n1760 VSS.n1268 0.00658571
R75884 VSS.n1766 VSS.n1268 0.00658571
R75885 VSS.n1767 VSS.n1766 0.00658571
R75886 VSS.n1768 VSS.n1767 0.00658571
R75887 VSS.n1768 VSS.n1264 0.00658571
R75888 VSS.n1774 VSS.n1264 0.00658571
R75889 VSS.n1775 VSS.n1774 0.00658571
R75890 VSS.n1776 VSS.n1775 0.00658571
R75891 VSS.n1776 VSS.n1260 0.00658571
R75892 VSS.n1782 VSS.n1260 0.00658571
R75893 VSS.n1783 VSS.n1782 0.00658571
R75894 VSS.n1823 VSS.n1783 0.00658571
R75895 VSS.n1823 VSS.n1822 0.00658571
R75896 VSS.n1822 VSS.n1821 0.00658571
R75897 VSS.n1821 VSS.n1784 0.00658571
R75898 VSS.n1788 VSS.n1784 0.00658571
R75899 VSS.n1814 VSS.n1788 0.00658571
R75900 VSS.n1814 VSS.n1813 0.00658571
R75901 VSS.n1813 VSS.n1812 0.00658571
R75902 VSS.n1812 VSS.n1789 0.00658571
R75903 VSS.n1806 VSS.n1789 0.00658571
R75904 VSS.n1806 VSS.n1805 0.00658571
R75905 VSS.n1805 VSS.n1804 0.00658571
R75906 VSS.n1804 VSS.n1793 0.00658571
R75907 VSS.n1798 VSS.n1793 0.00658571
R75908 VSS.n1798 VSS.n1797 0.00658571
R75909 VSS.n2052 VSS.n2051 0.00658571
R75910 VSS.n2051 VSS.n2050 0.00658571
R75911 VSS.n2050 VSS.n1911 0.00658571
R75912 VSS.n2044 VSS.n1911 0.00658571
R75913 VSS.n2044 VSS.n2043 0.00658571
R75914 VSS.n2043 VSS.n2042 0.00658571
R75915 VSS.n2042 VSS.n1915 0.00658571
R75916 VSS.n2036 VSS.n1915 0.00658571
R75917 VSS.n2036 VSS.n2035 0.00658571
R75918 VSS.n2035 VSS.n2034 0.00658571
R75919 VSS.n2034 VSS.n1919 0.00658571
R75920 VSS.n2028 VSS.n1919 0.00658571
R75921 VSS.n2028 VSS.n2027 0.00658571
R75922 VSS.n2027 VSS.n2026 0.00658571
R75923 VSS.n2026 VSS.n1923 0.00658571
R75924 VSS.n2019 VSS.n1923 0.00658571
R75925 VSS.n2019 VSS.n2018 0.00658571
R75926 VSS.n2018 VSS.n2017 0.00658571
R75927 VSS.n2017 VSS.n1925 0.00658571
R75928 VSS.n2011 VSS.n1925 0.00658571
R75929 VSS.n2011 VSS.n2010 0.00658571
R75930 VSS.n2010 VSS.n2009 0.00658571
R75931 VSS.n2009 VSS.n1930 0.00658571
R75932 VSS.n2003 VSS.n1930 0.00658571
R75933 VSS.n2003 VSS.n2002 0.00658571
R75934 VSS.n2002 VSS.n2001 0.00658571
R75935 VSS.n2001 VSS.n1934 0.00658571
R75936 VSS.n1995 VSS.n1934 0.00658571
R75937 VSS.n1995 VSS.n1994 0.00658571
R75938 VSS.n1994 VSS.n1993 0.00658571
R75939 VSS.n1993 VSS.n1938 0.00658571
R75940 VSS.n1987 VSS.n1938 0.00658571
R75941 VSS.n1987 VSS.n1986 0.00658571
R75942 VSS.n1986 VSS.n1985 0.00658571
R75943 VSS.n1985 VSS.n1942 0.00658571
R75944 VSS.n1946 VSS.n1942 0.00658571
R75945 VSS.n1978 VSS.n1946 0.00658571
R75946 VSS.n1978 VSS.n1977 0.00658571
R75947 VSS.n1977 VSS.n1976 0.00658571
R75948 VSS.n1976 VSS.n1947 0.00658571
R75949 VSS.n1970 VSS.n1947 0.00658571
R75950 VSS.n1970 VSS.n1969 0.00658571
R75951 VSS.n1969 VSS.n1968 0.00658571
R75952 VSS.n1968 VSS.n1951 0.00658571
R75953 VSS.n1962 VSS.n1951 0.00658571
R75954 VSS.n1962 VSS.n1961 0.00658571
R75955 VSS.n1961 VSS.n1960 0.00658571
R75956 VSS.n1960 VSS.n1955 0.00658571
R75957 VSS.n1955 VSS.n1079 0.00658571
R75958 VSS.n2989 VSS.n1079 0.00658571
R75959 VSS.n2990 VSS.n2989 0.00658571
R75960 VSS.n2991 VSS.n2990 0.00658571
R75961 VSS.n2991 VSS.n1075 0.00658571
R75962 VSS.n2997 VSS.n1075 0.00658571
R75963 VSS.n2998 VSS.n2997 0.00658571
R75964 VSS.n2999 VSS.n2998 0.00658571
R75965 VSS.n2999 VSS.n1071 0.00658571
R75966 VSS.n3005 VSS.n1071 0.00658571
R75967 VSS.n3006 VSS.n3005 0.00658571
R75968 VSS.n3007 VSS.n3006 0.00658571
R75969 VSS.n3007 VSS.n1067 0.00658571
R75970 VSS.n3013 VSS.n1067 0.00658571
R75971 VSS.n3014 VSS.n3013 0.00658571
R75972 VSS.n3015 VSS.n3014 0.00658571
R75973 VSS.n3015 VSS.n1063 0.00658571
R75974 VSS.n3021 VSS.n1063 0.00658571
R75975 VSS.n3022 VSS.n3021 0.00658571
R75976 VSS.n3061 VSS.n3022 0.00658571
R75977 VSS.n3061 VSS.n3060 0.00658571
R75978 VSS.n3060 VSS.n3059 0.00658571
R75979 VSS.n3059 VSS.n3023 0.00658571
R75980 VSS.n3053 VSS.n3023 0.00658571
R75981 VSS.n3053 VSS.n3052 0.00658571
R75982 VSS.n3052 VSS.n3051 0.00658571
R75983 VSS.n3051 VSS.n3028 0.00658571
R75984 VSS.n3045 VSS.n3028 0.00658571
R75985 VSS.n3045 VSS.n3044 0.00658571
R75986 VSS.n3044 VSS.n3043 0.00658571
R75987 VSS.n3043 VSS.n3032 0.00658571
R75988 VSS.n3037 VSS.n3032 0.00658571
R75989 VSS.n3037 VSS.n3036 0.00658571
R75990 VSS.n2692 VSS.n2691 0.00658571
R75991 VSS.n2692 VSS.n1180 0.00658571
R75992 VSS.n2698 VSS.n1180 0.00658571
R75993 VSS.n2699 VSS.n2698 0.00658571
R75994 VSS.n2700 VSS.n2699 0.00658571
R75995 VSS.n2700 VSS.n1176 0.00658571
R75996 VSS.n2706 VSS.n1176 0.00658571
R75997 VSS.n2707 VSS.n2706 0.00658571
R75998 VSS.n2708 VSS.n2707 0.00658571
R75999 VSS.n2708 VSS.n1172 0.00658571
R76000 VSS.n2714 VSS.n1172 0.00658571
R76001 VSS.n2715 VSS.n2714 0.00658571
R76002 VSS.n2716 VSS.n2715 0.00658571
R76003 VSS.n2716 VSS.n1168 0.00658571
R76004 VSS.n2722 VSS.n1168 0.00658571
R76005 VSS.n2723 VSS.n2722 0.00658571
R76006 VSS.n2856 VSS.n2723 0.00658571
R76007 VSS.n2856 VSS.n2855 0.00658571
R76008 VSS.n2855 VSS.n2854 0.00658571
R76009 VSS.n2854 VSS.n2724 0.00658571
R76010 VSS.n2848 VSS.n2724 0.00658571
R76011 VSS.n2848 VSS.n2847 0.00658571
R76012 VSS.n2847 VSS.n2846 0.00658571
R76013 VSS.n2846 VSS.n2728 0.00658571
R76014 VSS.n2840 VSS.n2728 0.00658571
R76015 VSS.n2840 VSS.n2839 0.00658571
R76016 VSS.n2839 VSS.n2838 0.00658571
R76017 VSS.n2838 VSS.n2732 0.00658571
R76018 VSS.n2832 VSS.n2732 0.00658571
R76019 VSS.n2832 VSS.n2831 0.00658571
R76020 VSS.n2831 VSS.n2830 0.00658571
R76021 VSS.n2830 VSS.n2736 0.00658571
R76022 VSS.n2757 VSS.n2736 0.00658571
R76023 VSS.n2758 VSS.n2757 0.00658571
R76024 VSS.n2809 VSS.n2758 0.00658571
R76025 VSS.n2809 VSS.n2808 0.00658571
R76026 VSS.n2808 VSS.n2807 0.00658571
R76027 VSS.n2807 VSS.n2759 0.00658571
R76028 VSS.n2801 VSS.n2759 0.00658571
R76029 VSS.n2801 VSS.n2800 0.00658571
R76030 VSS.n2800 VSS.n2799 0.00658571
R76031 VSS.n2799 VSS.n2763 0.00658571
R76032 VSS.n2793 VSS.n2763 0.00658571
R76033 VSS.n2793 VSS.n2792 0.00658571
R76034 VSS.n2792 VSS.n2791 0.00658571
R76035 VSS.n2791 VSS.n2767 0.00658571
R76036 VSS.n2785 VSS.n2767 0.00658571
R76037 VSS.n2785 VSS.n2784 0.00658571
R76038 VSS.n2784 VSS.n2783 0.00658571
R76039 VSS.n2783 VSS.n2771 0.00658571
R76040 VSS.n2771 VSS.n983 0.00658571
R76041 VSS.n3433 VSS.n983 0.00658571
R76042 VSS.n3433 VSS.n3432 0.00658571
R76043 VSS.n3432 VSS.n3431 0.00658571
R76044 VSS.n3431 VSS.n984 0.00658571
R76045 VSS.n3425 VSS.n984 0.00658571
R76046 VSS.n3425 VSS.n3424 0.00658571
R76047 VSS.n3424 VSS.n3423 0.00658571
R76048 VSS.n3423 VSS.n988 0.00658571
R76049 VSS.n3417 VSS.n988 0.00658571
R76050 VSS.n3417 VSS.n3416 0.00658571
R76051 VSS.n3416 VSS.n3415 0.00658571
R76052 VSS.n3415 VSS.n992 0.00658571
R76053 VSS.n3409 VSS.n992 0.00658571
R76054 VSS.n3409 VSS.n3408 0.00658571
R76055 VSS.n3408 VSS.n3407 0.00658571
R76056 VSS.n3407 VSS.n996 0.00658571
R76057 VSS.n1007 VSS.n996 0.00658571
R76058 VSS.n1042 VSS.n1007 0.00658571
R76059 VSS.n1042 VSS.n1041 0.00658571
R76060 VSS.n1041 VSS.n1040 0.00658571
R76061 VSS.n1040 VSS.n1008 0.00658571
R76062 VSS.n1034 VSS.n1008 0.00658571
R76063 VSS.n1034 VSS.n1033 0.00658571
R76064 VSS.n1033 VSS.n1032 0.00658571
R76065 VSS.n1032 VSS.n1012 0.00658571
R76066 VSS.n1026 VSS.n1012 0.00658571
R76067 VSS.n1026 VSS.n1025 0.00658571
R76068 VSS.n1025 VSS.n1024 0.00658571
R76069 VSS.n1024 VSS.n1016 0.00658571
R76070 VSS.n1018 VSS.n1016 0.00658571
R76071 VSS.n2200 VSS.n2199 0.00658571
R76072 VSS.n2199 VSS.n2198 0.00658571
R76073 VSS.n2198 VSS.n2156 0.00658571
R76074 VSS.n2192 VSS.n2156 0.00658571
R76075 VSS.n2192 VSS.n2191 0.00658571
R76076 VSS.n2191 VSS.n2190 0.00658571
R76077 VSS.n2190 VSS.n2160 0.00658571
R76078 VSS.n2184 VSS.n2160 0.00658571
R76079 VSS.n2184 VSS.n2183 0.00658571
R76080 VSS.n2183 VSS.n2182 0.00658571
R76081 VSS.n2182 VSS.n2164 0.00658571
R76082 VSS.n2176 VSS.n2164 0.00658571
R76083 VSS.n2176 VSS.n2175 0.00658571
R76084 VSS.n2175 VSS.n2174 0.00658571
R76085 VSS.n2174 VSS.n2168 0.00658571
R76086 VSS.n2169 VSS.n2168 0.00658571
R76087 VSS.n2169 VSS.n652 0.00658571
R76088 VSS.n3941 VSS.n652 0.00658571
R76089 VSS.n3942 VSS.n3941 0.00658571
R76090 VSS.n3943 VSS.n3942 0.00658571
R76091 VSS.n3943 VSS.n648 0.00658571
R76092 VSS.n3949 VSS.n648 0.00658571
R76093 VSS.n3950 VSS.n3949 0.00658571
R76094 VSS.n3951 VSS.n3950 0.00658571
R76095 VSS.n3951 VSS.n644 0.00658571
R76096 VSS.n3957 VSS.n644 0.00658571
R76097 VSS.n3958 VSS.n3957 0.00658571
R76098 VSS.n3959 VSS.n3958 0.00658571
R76099 VSS.n3959 VSS.n640 0.00658571
R76100 VSS.n3965 VSS.n640 0.00658571
R76101 VSS.n3966 VSS.n3965 0.00658571
R76102 VSS.n3967 VSS.n3966 0.00658571
R76103 VSS.n3967 VSS.n620 0.00658571
R76104 VSS.n3982 VSS.n620 0.00658571
R76105 VSS.n3983 VSS.n3982 0.00658571
R76106 VSS.n3984 VSS.n3983 0.00658571
R76107 VSS.n3984 VSS.n616 0.00658571
R76108 VSS.n3990 VSS.n616 0.00658571
R76109 VSS.n3991 VSS.n3990 0.00658571
R76110 VSS.n3992 VSS.n3991 0.00658571
R76111 VSS.n3992 VSS.n612 0.00658571
R76112 VSS.n3998 VSS.n612 0.00658571
R76113 VSS.n3999 VSS.n3998 0.00658571
R76114 VSS.n4000 VSS.n3999 0.00658571
R76115 VSS.n4000 VSS.n608 0.00658571
R76116 VSS.n4006 VSS.n608 0.00658571
R76117 VSS.n4007 VSS.n4006 0.00658571
R76118 VSS.n4008 VSS.n4007 0.00658571
R76119 VSS.n4008 VSS.n604 0.00658571
R76120 VSS.n4014 VSS.n604 0.00658571
R76121 VSS.n4015 VSS.n4014 0.00658571
R76122 VSS.n4016 VSS.n4015 0.00658571
R76123 VSS.n4016 VSS.n600 0.00658571
R76124 VSS.n4022 VSS.n600 0.00658571
R76125 VSS.n4023 VSS.n4022 0.00658571
R76126 VSS.n4024 VSS.n4023 0.00658571
R76127 VSS.n4024 VSS.n596 0.00658571
R76128 VSS.n4030 VSS.n596 0.00658571
R76129 VSS.n4031 VSS.n4030 0.00658571
R76130 VSS.n4032 VSS.n4031 0.00658571
R76131 VSS.n4032 VSS.n592 0.00658571
R76132 VSS.n4038 VSS.n592 0.00658571
R76133 VSS.n4039 VSS.n4038 0.00658571
R76134 VSS.n4040 VSS.n4039 0.00658571
R76135 VSS.n4040 VSS.n588 0.00658571
R76136 VSS.n4046 VSS.n588 0.00658571
R76137 VSS.n4047 VSS.n4046 0.00658571
R76138 VSS.n4086 VSS.n4047 0.00658571
R76139 VSS.n4086 VSS.n4085 0.00658571
R76140 VSS.n4085 VSS.n4084 0.00658571
R76141 VSS.n4084 VSS.n4048 0.00658571
R76142 VSS.n4078 VSS.n4048 0.00658571
R76143 VSS.n4078 VSS.n4077 0.00658571
R76144 VSS.n4077 VSS.n4076 0.00658571
R76145 VSS.n4076 VSS.n4053 0.00658571
R76146 VSS.n4070 VSS.n4053 0.00658571
R76147 VSS.n4070 VSS.n4069 0.00658571
R76148 VSS.n4069 VSS.n4068 0.00658571
R76149 VSS.n4068 VSS.n4057 0.00658571
R76150 VSS.n4062 VSS.n4057 0.00658571
R76151 VSS.n4062 VSS.n4061 0.00658571
R76152 VSS.n4573 VSS.n4572 0.00658571
R76153 VSS.n4573 VSS.n4567 0.00658571
R76154 VSS.n4579 VSS.n4567 0.00658571
R76155 VSS.n4580 VSS.n4579 0.00658571
R76156 VSS.n4581 VSS.n4580 0.00658571
R76157 VSS.n4581 VSS.n4563 0.00658571
R76158 VSS.n4587 VSS.n4563 0.00658571
R76159 VSS.n4588 VSS.n4587 0.00658571
R76160 VSS.n4589 VSS.n4588 0.00658571
R76161 VSS.n4589 VSS.n4559 0.00658571
R76162 VSS.n4595 VSS.n4559 0.00658571
R76163 VSS.n4596 VSS.n4595 0.00658571
R76164 VSS.n4598 VSS.n4596 0.00658571
R76165 VSS.n4598 VSS.n4597 0.00658571
R76166 VSS.n4597 VSS.n4555 0.00658571
R76167 VSS.n4605 VSS.n4555 0.00658571
R76168 VSS.n4606 VSS.n4605 0.00658571
R76169 VSS.n4607 VSS.n4606 0.00658571
R76170 VSS.n4607 VSS.n4552 0.00658571
R76171 VSS.n4613 VSS.n4552 0.00658571
R76172 VSS.n4614 VSS.n4613 0.00658571
R76173 VSS.n4615 VSS.n4614 0.00658571
R76174 VSS.n4615 VSS.n4548 0.00658571
R76175 VSS.n4621 VSS.n4548 0.00658571
R76176 VSS.n4622 VSS.n4621 0.00658571
R76177 VSS.n4623 VSS.n4622 0.00658571
R76178 VSS.n4623 VSS.n4544 0.00658571
R76179 VSS.n4629 VSS.n4544 0.00658571
R76180 VSS.n4630 VSS.n4629 0.00658571
R76181 VSS.n4631 VSS.n4630 0.00658571
R76182 VSS.n4631 VSS.n4540 0.00658571
R76183 VSS.n4637 VSS.n4540 0.00658571
R76184 VSS.n4638 VSS.n4637 0.00658571
R76185 VSS.n4639 VSS.n4638 0.00658571
R76186 VSS.n4639 VSS.n4537 0.00658571
R76187 VSS.n4644 VSS.n4537 0.00658571
R76188 VSS.n4645 VSS.n4644 0.00658571
R76189 VSS.n4646 VSS.n4645 0.00658571
R76190 VSS.n4646 VSS.n4533 0.00658571
R76191 VSS.n4652 VSS.n4533 0.00658571
R76192 VSS.n4653 VSS.n4652 0.00658571
R76193 VSS.n4654 VSS.n4653 0.00658571
R76194 VSS.n4654 VSS.n4529 0.00658571
R76195 VSS.n4660 VSS.n4529 0.00658571
R76196 VSS.n4661 VSS.n4660 0.00658571
R76197 VSS.n4662 VSS.n4661 0.00658571
R76198 VSS.n4662 VSS.n4525 0.00658571
R76199 VSS.n4668 VSS.n4525 0.00658571
R76200 VSS.n4669 VSS.n4668 0.00658571
R76201 VSS.n4758 VSS.n4669 0.00658571
R76202 VSS.n4758 VSS.n4757 0.00658571
R76203 VSS.n4757 VSS.n4756 0.00658571
R76204 VSS.n4756 VSS.n4670 0.00658571
R76205 VSS.n4674 VSS.n4670 0.00658571
R76206 VSS.n4749 VSS.n4674 0.00658571
R76207 VSS.n4749 VSS.n4748 0.00658571
R76208 VSS.n4748 VSS.n4747 0.00658571
R76209 VSS.n4747 VSS.n4675 0.00658571
R76210 VSS.n4741 VSS.n4675 0.00658571
R76211 VSS.n4741 VSS.n4740 0.00658571
R76212 VSS.n4740 VSS.n4739 0.00658571
R76213 VSS.n4739 VSS.n4679 0.00658571
R76214 VSS.n4733 VSS.n4679 0.00658571
R76215 VSS.n4733 VSS.n4732 0.00658571
R76216 VSS.n4732 VSS.n4731 0.00658571
R76217 VSS.n4731 VSS.n4683 0.00658571
R76218 VSS.n4725 VSS.n4683 0.00658571
R76219 VSS.n4725 VSS.n4724 0.00658571
R76220 VSS.n4724 VSS.n4723 0.00658571
R76221 VSS.n4723 VSS.n4686 0.00658571
R76222 VSS.n4690 VSS.n4686 0.00658571
R76223 VSS.n4716 VSS.n4690 0.00658571
R76224 VSS.n4716 VSS.n4715 0.00658571
R76225 VSS.n4715 VSS.n4714 0.00658571
R76226 VSS.n4714 VSS.n4691 0.00658571
R76227 VSS.n4708 VSS.n4691 0.00658571
R76228 VSS.n4708 VSS.n4707 0.00658571
R76229 VSS.n4707 VSS.n4706 0.00658571
R76230 VSS.n4706 VSS.n4695 0.00658571
R76231 VSS.n4700 VSS.n4695 0.00658571
R76232 VSS.n4700 VSS.n4699 0.00658571
R76233 VSS.n6443 VSS.n23 0.00658571
R76234 VSS.n6437 VSS.n23 0.00658571
R76235 VSS.n6437 VSS.n6436 0.00658571
R76236 VSS.n6436 VSS.n6435 0.00658571
R76237 VSS.n6435 VSS.n27 0.00658571
R76238 VSS.n6429 VSS.n27 0.00658571
R76239 VSS.n6429 VSS.n6428 0.00658571
R76240 VSS.n6428 VSS.n6427 0.00658571
R76241 VSS.n6427 VSS.n31 0.00658571
R76242 VSS.n6421 VSS.n31 0.00658571
R76243 VSS.n6421 VSS.n6420 0.00658571
R76244 VSS.n6420 VSS.n6419 0.00658571
R76245 VSS.n6419 VSS.n35 0.00658571
R76246 VSS.n6413 VSS.n35 0.00658571
R76247 VSS.n6413 VSS.n6412 0.00658571
R76248 VSS.n6412 VSS.n6411 0.00658571
R76249 VSS.n6411 VSS.n39 0.00658571
R76250 VSS.n6405 VSS.n39 0.00658571
R76251 VSS.n6405 VSS.n6404 0.00658571
R76252 VSS.n6404 VSS.n6403 0.00658571
R76253 VSS.n6403 VSS.n43 0.00658571
R76254 VSS.n6397 VSS.n43 0.00658571
R76255 VSS.n6397 VSS.n6396 0.00658571
R76256 VSS.n6396 VSS.n6395 0.00658571
R76257 VSS.n6395 VSS.n47 0.00658571
R76258 VSS.n6389 VSS.n47 0.00658571
R76259 VSS.n6389 VSS.n6388 0.00658571
R76260 VSS.n6388 VSS.n6387 0.00658571
R76261 VSS.n6387 VSS.n51 0.00658571
R76262 VSS.n6381 VSS.n51 0.00658571
R76263 VSS.n6381 VSS.n6380 0.00658571
R76264 VSS.n6380 VSS.n6379 0.00658571
R76265 VSS.n6379 VSS.n55 0.00658571
R76266 VSS.n6373 VSS.n55 0.00658571
R76267 VSS.n6373 VSS.n6372 0.00658571
R76268 VSS.n6372 VSS.n6371 0.00658571
R76269 VSS.n6371 VSS.n59 0.00658571
R76270 VSS.n6365 VSS.n59 0.00658571
R76271 VSS.n6365 VSS.n6364 0.00658571
R76272 VSS.n6364 VSS.n6363 0.00658571
R76273 VSS.n6363 VSS.n63 0.00658571
R76274 VSS.n6357 VSS.n63 0.00658571
R76275 VSS.n6357 VSS.n6356 0.00658571
R76276 VSS.n6356 VSS.n6355 0.00658571
R76277 VSS.n6355 VSS.n67 0.00658571
R76278 VSS.n6349 VSS.n67 0.00658571
R76279 VSS.n6349 VSS.n6348 0.00658571
R76280 VSS.n6348 VSS.n6347 0.00658571
R76281 VSS.n6347 VSS.n71 0.00658571
R76282 VSS.n6341 VSS.n71 0.00658571
R76283 VSS.n6341 VSS.n6340 0.00658571
R76284 VSS.n6340 VSS.n6339 0.00658571
R76285 VSS.n6339 VSS.n75 0.00658571
R76286 VSS.n6333 VSS.n75 0.00658571
R76287 VSS.n6333 VSS.n6332 0.00658571
R76288 VSS.n6332 VSS.n6331 0.00658571
R76289 VSS.n6331 VSS.n79 0.00658571
R76290 VSS.n6325 VSS.n79 0.00658571
R76291 VSS.n6325 VSS.n6324 0.00658571
R76292 VSS.n6324 VSS.n6323 0.00658571
R76293 VSS.n6323 VSS.n83 0.00658571
R76294 VSS.n6317 VSS.n83 0.00658571
R76295 VSS.n6317 VSS.n6316 0.00658571
R76296 VSS.n6316 VSS.n6315 0.00658571
R76297 VSS.n6315 VSS.n87 0.00658571
R76298 VSS.n6309 VSS.n87 0.00658571
R76299 VSS.n6309 VSS.n6308 0.00658571
R76300 VSS.n6308 VSS.n6307 0.00658571
R76301 VSS.n6307 VSS.n91 0.00658571
R76302 VSS.n6301 VSS.n91 0.00658571
R76303 VSS.n6301 VSS.n6300 0.00658571
R76304 VSS.n6300 VSS.n6299 0.00658571
R76305 VSS.n6299 VSS.n95 0.00658571
R76306 VSS.n6293 VSS.n95 0.00658571
R76307 VSS.n6293 VSS.n6292 0.00658571
R76308 VSS.n6292 VSS.n6291 0.00658571
R76309 VSS.n6291 VSS.n99 0.00658571
R76310 VSS.n6285 VSS.n99 0.00658571
R76311 VSS.n6285 VSS.n6284 0.00658571
R76312 VSS.n6284 VSS.n6283 0.00658571
R76313 VSS.n6283 VSS.n103 0.00658571
R76314 VSS.n6277 VSS.n103 0.00658571
R76315 VSS.n6277 VSS.n6276 0.00658571
R76316 VSS.n6276 VSS.n6275 0.00658571
R76317 VSS.n6275 VSS.n107 0.00658571
R76318 VSS.n6268 VSS.n107 0.00658571
R76319 VSS.n6268 VSS.n6267 0.00658571
R76320 VSS.n6267 VSS.n6266 0.00658571
R76321 VSS.n6266 VSS.n112 0.00658571
R76322 VSS.n6260 VSS.n112 0.00658571
R76323 VSS.n6260 VSS.n6259 0.00658571
R76324 VSS.n6259 VSS.n6258 0.00658571
R76325 VSS.n6258 VSS.n116 0.00658571
R76326 VSS.n6252 VSS.n116 0.00658571
R76327 VSS.n6252 VSS.n6251 0.00658571
R76328 VSS.n6251 VSS.n6250 0.00658571
R76329 VSS.n6250 VSS.n120 0.00658571
R76330 VSS.n6244 VSS.n6243 0.00658571
R76331 DVSS VSS.n3761 0.00656742
R76332 VSS.n5829 VSS.n5826 0.00654478
R76333 VSS.n5430 VSS.n4368 0.0065
R76334 VSS.n6007 VSS.n4443 0.0065
R76335 VSS.n5388 VSS.n5329 0.0065
R76336 VSS.n5761 VSS.n4365 0.0065
R76337 VSS.n5906 VSS.n4907 0.0065
R76338 VSS.n6053 VSS.n4365 0.0065
R76339 VSS.n5388 VSS.n5330 0.0065
R76340 VSS.n5171 VSS.n4442 0.0065
R76341 VSS.n5171 VSS.n5167 0.0065
R76342 VSS.n5906 VSS.n5905 0.0065
R76343 VSS.n5386 VSS.n5379 0.0065
R76344 VSS.n5430 VSS.n5134 0.0065
R76345 VSS.n5724 VSS.n4443 0.0065
R76346 VSS.n5980 VSS.n4908 0.0065
R76347 VSS.n5870 VSS.n4908 0.0065
R76348 VSS.n5386 VSS.n5385 0.0065
R76349 VSS VSS.n6466 0.00641429
R76350 VSS.n6244 VSS 0.00641429
R76351 VSS.n1830 VSS.n1825 0.00635
R76352 VSS.n3064 VSS.n1050 0.00635
R76353 VSS.n3404 VSS.n3403 0.00635
R76354 VSS.n4089 VSS.n575 0.00635
R76355 VSS.n4727 VSS.n489 0.00635
R76356 VSS.n4849 VSS.n4388 0.00620896
R76357 VSS.n1906 VSS.n1205 0.00609286
R76358 VSS.n2055 VSS.n2054 0.00609286
R76359 VSS.n2687 VSS.n1182 0.00609286
R76360 VSS.n2203 VSS.n2202 0.00609286
R76361 VSS.n6129 VSS.n4255 0.00609286
R76362 DVSS VSS.n1857 0.00585211
R76363 VSS.n1879 VSS.n1236 0.00564085
R76364 VSS.n5809 VSS.n5030 0.00553731
R76365 VSS.n6242 VSS.n6241 0.00548841
R76366 VSS.n6444 VSS.n22 0.00548841
R76367 VSS.n4 VSS.n3 0.00548841
R76368 VSS.n241 VSS 0.00538571
R76369 VSS.n1660 VSS.n1320 0.00536196
R76370 VSS.n1661 VSS.n1660 0.00536196
R76371 VSS.n1549 VSS.n1548 0.00535915
R76372 VSS.n1879 VSS.n1878 0.00535915
R76373 VSS.n1833 VSS.n1250 0.00519286
R76374 VSS.n3063 VSS.n1060 0.00519286
R76375 VSS.n3067 VSS.n1003 0.00519286
R76376 VSS.n4088 VSS.n585 0.00519286
R76377 VSS.n6139 VSS.n491 0.00519286
R76378 VSS.n1891 VSS.n1218 0.00513023
R76379 VSS.n1893 VSS.n1218 0.00513023
R76380 VSS.n3862 VSS.n730 0.00503358
R76381 VSS.n1885 VSS.n1231 0.005
R76382 VSS.n4821 VSS.n4820 0.005
R76383 VSS.n5514 VSS.n4954 0.005
R76384 VSS.n1889 VSS.n1227 0.005
R76385 VSS.n4812 VSS.n4810 0.005
R76386 VSS.n5515 VSS.n5183 0.005
R76387 VSS.n1895 VSS.n1215 0.005
R76388 VSS.n4814 VSS.n4307 0.005
R76389 VSS.n5510 VSS.n5294 0.005
R76390 VSS.n1901 VSS.n1203 0.005
R76391 VSS.n4815 VSS.n4325 0.005
R76392 VSS.n5511 VSS.n5279 0.005
R76393 VSS.n1493 VSS.n1491 0.00498219
R76394 VSS.n2975 VSS.n1105 0.00498219
R76395 VSS.n2822 VSS.n2746 0.00498219
R76396 VSS.n3977 VSS.n3976 0.00498219
R76397 VSS.n4506 VSS.n4502 0.00498219
R76398 VSS.n4502 VSS.n4489 0.00498219
R76399 VSS.n3977 VSS.n622 0.00498219
R76400 VSS.n2822 VSS.n2821 0.00498219
R76401 VSS.n1105 VSS.n1103 0.00498219
R76402 VSS.n1491 VSS.n1432 0.00498219
R76403 VSS.n1903 VSS.n1200 0.00493571
R76404 VSS.n1833 VSS.n1252 0.00493571
R76405 VSS.n1909 VSS.n1186 0.00493571
R76406 VSS.n3025 VSS.n1060 0.00493571
R76407 VSS.n2688 VSS.n1184 0.00493571
R76408 VSS.n3067 VSS.n1044 0.00493571
R76409 VSS.n2151 VSS.n2150 0.00493571
R76410 VSS.n4050 VSS.n585 0.00493571
R76411 VSS.n4263 VSS.n4251 0.00493571
R76412 VSS.n6139 VSS.n498 0.00493571
R76413 VSS.n1424 VSS.n1221 0.00486567
R76414 VSS.n4837 VSS.n4409 0.00486567
R76415 VSS.n2133 VSS.n2132 0.00476
R76416 VSS.n2132 VSS.n2131 0.00476
R76417 VSS.n2131 VSS.n2094 0.00476
R76418 VSS.n2127 VSS.n2094 0.00476
R76419 VSS.n2127 VSS.n2126 0.00476
R76420 VSS.n2126 VSS.n2125 0.00476
R76421 VSS.n2125 VSS.n2100 0.00476
R76422 VSS.n2121 VSS.n2100 0.00476
R76423 VSS.n2121 VSS.n2120 0.00476
R76424 VSS.n2120 VSS.n2119 0.00476
R76425 VSS.n2119 VSS.n2106 0.00476
R76426 VSS.n2115 VSS.n2106 0.00476
R76427 VSS.n2115 VSS.n2114 0.00476
R76428 VSS.n2114 VSS.n2113 0.00476
R76429 VSS.n2113 VSS.n966 0.00476
R76430 VSS.n3536 VSS.n966 0.00476
R76431 VSS.n3536 VSS.n964 0.00476
R76432 VSS.n3540 VSS.n964 0.00476
R76433 VSS.n3540 VSS.n962 0.00476
R76434 VSS.n3544 VSS.n962 0.00476
R76435 VSS.n3544 VSS.n960 0.00476
R76436 VSS.n3548 VSS.n960 0.00476
R76437 VSS.n3548 VSS.n958 0.00476
R76438 VSS.n3552 VSS.n958 0.00476
R76439 VSS.n3552 VSS.n956 0.00476
R76440 VSS.n3556 VSS.n956 0.00476
R76441 VSS.n3556 VSS.n954 0.00476
R76442 VSS.n3560 VSS.n954 0.00476
R76443 VSS.n3560 VSS.n952 0.00476
R76444 VSS.n3564 VSS.n952 0.00476
R76445 VSS.n3564 VSS.n950 0.00476
R76446 VSS.n3569 VSS.n950 0.00476
R76447 VSS.n3569 VSS.n948 0.00476
R76448 VSS.n3575 VSS.n948 0.00476
R76449 VSS.n3575 VSS.n3574 0.00476
R76450 VSS.n3574 VSS.n910 0.00476
R76451 VSS.n3594 VSS.n910 0.00476
R76452 VSS.n3594 VSS.n908 0.00476
R76453 VSS.n3598 VSS.n908 0.00476
R76454 VSS.n3598 VSS.n906 0.00476
R76455 VSS.n3602 VSS.n906 0.00476
R76456 VSS.n3602 VSS.n904 0.00476
R76457 VSS.n3606 VSS.n904 0.00476
R76458 VSS.n3606 VSS.n902 0.00476
R76459 VSS.n3610 VSS.n902 0.00476
R76460 VSS.n3610 VSS.n900 0.00476
R76461 VSS.n3614 VSS.n900 0.00476
R76462 VSS.n3614 VSS.n898 0.00476
R76463 VSS.n3618 VSS.n898 0.00476
R76464 VSS.n3618 VSS.n896 0.00476
R76465 VSS.n3624 VSS.n896 0.00476
R76466 VSS.n3624 VSS.n3623 0.00476
R76467 VSS.n3623 VSS.n880 0.00476
R76468 VSS.n3643 VSS.n880 0.00476
R76469 VSS.n3643 VSS.n878 0.00476
R76470 VSS.n3647 VSS.n878 0.00476
R76471 VSS.n3647 VSS.n876 0.00476
R76472 VSS.n3651 VSS.n876 0.00476
R76473 VSS.n3651 VSS.n874 0.00476
R76474 VSS.n3655 VSS.n874 0.00476
R76475 VSS.n3655 VSS.n872 0.00476
R76476 VSS.n3659 VSS.n872 0.00476
R76477 VSS.n3659 VSS.n870 0.00476
R76478 VSS.n3663 VSS.n870 0.00476
R76479 VSS.n3663 VSS.n868 0.00476
R76480 VSS.n3667 VSS.n868 0.00476
R76481 VSS.n3667 VSS.n866 0.00476
R76482 VSS.n3711 VSS.n866 0.00476
R76483 VSS.n3711 VSS.n3710 0.00476
R76484 VSS.n3710 VSS.n3709 0.00476
R76485 VSS.n3709 VSS.n3708 0.00476
R76486 VSS.n3708 VSS.n3674 0.00476
R76487 VSS.n3704 VSS.n3674 0.00476
R76488 VSS.n3704 VSS.n3703 0.00476
R76489 VSS.n3703 VSS.n3702 0.00476
R76490 VSS.n3702 VSS.n3680 0.00476
R76491 VSS.n3698 VSS.n3680 0.00476
R76492 VSS.n3698 VSS.n3697 0.00476
R76493 VSS.n3697 VSS.n3696 0.00476
R76494 VSS.n3696 VSS.n3686 0.00476
R76495 VSS.n3692 VSS.n3686 0.00476
R76496 VSS.n2130 VSS.n2080 0.00476
R76497 VSS.n2130 VSS.n2129 0.00476
R76498 VSS.n2129 VSS.n2128 0.00476
R76499 VSS.n2128 VSS.n2095 0.00476
R76500 VSS.n2124 VSS.n2095 0.00476
R76501 VSS.n2124 VSS.n2123 0.00476
R76502 VSS.n2123 VSS.n2122 0.00476
R76503 VSS.n2122 VSS.n2101 0.00476
R76504 VSS.n2118 VSS.n2101 0.00476
R76505 VSS.n2118 VSS.n2117 0.00476
R76506 VSS.n2117 VSS.n2116 0.00476
R76507 VSS.n2116 VSS.n2107 0.00476
R76508 VSS.n2112 VSS.n2107 0.00476
R76509 VSS.n2112 VSS.n967 0.00476
R76510 VSS.n3535 VSS.n967 0.00476
R76511 VSS.n3542 VSS.n3541 0.00476
R76512 VSS.n3543 VSS.n3542 0.00476
R76513 VSS.n3543 VSS.n959 0.00476
R76514 VSS.n3549 VSS.n959 0.00476
R76515 VSS.n3550 VSS.n3549 0.00476
R76516 VSS.n3551 VSS.n3550 0.00476
R76517 VSS.n3551 VSS.n955 0.00476
R76518 VSS.n3557 VSS.n955 0.00476
R76519 VSS.n3558 VSS.n3557 0.00476
R76520 VSS.n3559 VSS.n3558 0.00476
R76521 VSS.n3559 VSS.n951 0.00476
R76522 VSS.n3565 VSS.n951 0.00476
R76523 VSS.n3566 VSS.n3565 0.00476
R76524 VSS.n3568 VSS.n3566 0.00476
R76525 VSS.n3568 VSS.n3567 0.00476
R76526 VSS.n3593 VSS.n3592 0.00476
R76527 VSS.n3593 VSS.n907 0.00476
R76528 VSS.n3599 VSS.n907 0.00476
R76529 VSS.n3600 VSS.n3599 0.00476
R76530 VSS.n3601 VSS.n3600 0.00476
R76531 VSS.n3601 VSS.n903 0.00476
R76532 VSS.n3607 VSS.n903 0.00476
R76533 VSS.n3608 VSS.n3607 0.00476
R76534 VSS.n3609 VSS.n3608 0.00476
R76535 VSS.n3609 VSS.n899 0.00476
R76536 VSS.n3615 VSS.n899 0.00476
R76537 VSS.n3616 VSS.n3615 0.00476
R76538 VSS.n3617 VSS.n3616 0.00476
R76539 VSS.n3617 VSS.n895 0.00476
R76540 VSS.n3625 VSS.n895 0.00476
R76541 VSS.n3642 VSS.n3641 0.00476
R76542 VSS.n3642 VSS.n877 0.00476
R76543 VSS.n3648 VSS.n877 0.00476
R76544 VSS.n3649 VSS.n3648 0.00476
R76545 VSS.n3650 VSS.n3649 0.00476
R76546 VSS.n3650 VSS.n873 0.00476
R76547 VSS.n3656 VSS.n873 0.00476
R76548 VSS.n3657 VSS.n3656 0.00476
R76549 VSS.n3658 VSS.n3657 0.00476
R76550 VSS.n3658 VSS.n869 0.00476
R76551 VSS.n3664 VSS.n869 0.00476
R76552 VSS.n3665 VSS.n3664 0.00476
R76553 VSS.n3666 VSS.n3665 0.00476
R76554 VSS.n3666 VSS.n865 0.00476
R76555 VSS.n3712 VSS.n865 0.00476
R76556 VSS.n3707 VSS.n852 0.00476
R76557 VSS.n3707 VSS.n3706 0.00476
R76558 VSS.n3706 VSS.n3705 0.00476
R76559 VSS.n3705 VSS.n3675 0.00476
R76560 VSS.n3701 VSS.n3675 0.00476
R76561 VSS.n3701 VSS.n3700 0.00476
R76562 VSS.n3700 VSS.n3699 0.00476
R76563 VSS.n3699 VSS.n3681 0.00476
R76564 VSS.n3695 VSS.n3681 0.00476
R76565 VSS.n3695 VSS.n3694 0.00476
R76566 VSS.n3694 VSS.n3693 0.00476
R76567 VSS.n5381 VSS.n4334 0.00476
R76568 VSS.n6084 VSS.n4334 0.00476
R76569 VSS.n6084 VSS.n6083 0.00476
R76570 VSS.n6083 VSS.n6082 0.00476
R76571 VSS.n6082 VSS.n4338 0.00476
R76572 VSS.n6078 VSS.n4338 0.00476
R76573 VSS.n6078 VSS.n6077 0.00476
R76574 VSS.n6077 VSS.n6076 0.00476
R76575 VSS.n6076 VSS.n4344 0.00476
R76576 VSS.n6072 VSS.n4344 0.00476
R76577 VSS.n6072 VSS.n6071 0.00476
R76578 VSS.n6071 VSS.n6070 0.00476
R76579 VSS.n6070 VSS.n4350 0.00476
R76580 VSS.n6066 VSS.n4350 0.00476
R76581 VSS.n6066 VSS.n6065 0.00476
R76582 VSS.n6065 VSS.n6064 0.00476
R76583 VSS.n6064 VSS.n6062 0.00476
R76584 VSS.n6062 VSS.n6061 0.00476
R76585 VSS.n6061 VSS.n6060 0.00476
R76586 VSS.n6060 VSS.n6059 0.00476
R76587 VSS.n6059 VSS.n4360 0.00476
R76588 VSS.n6055 VSS.n4360 0.00476
R76589 VSS.n6055 VSS.n6054 0.00476
R76590 VSS.n6052 VSS.n4367 0.00476
R76591 VSS.n6048 VSS.n4367 0.00476
R76592 VSS.n6048 VSS.n6047 0.00476
R76593 VSS.n6047 VSS.n6046 0.00476
R76594 VSS.n6046 VSS.n4374 0.00476
R76595 VSS.n6042 VSS.n4374 0.00476
R76596 VSS.n6042 VSS.n6041 0.00476
R76597 VSS.n6041 VSS.n6040 0.00476
R76598 VSS.n6040 VSS.n4380 0.00476
R76599 VSS.n6036 VSS.n4380 0.00476
R76600 VSS.n6036 VSS.n6035 0.00476
R76601 VSS.n6035 VSS.n4385 0.00476
R76602 VSS.n6023 VSS.n4385 0.00476
R76603 VSS.n6023 VSS.n6022 0.00476
R76604 VSS.n6022 VSS.n6021 0.00476
R76605 VSS.n6021 VSS.n4430 0.00476
R76606 VSS.n6017 VSS.n4430 0.00476
R76607 VSS.n6017 VSS.n6016 0.00476
R76608 VSS.n6016 VSS.n6015 0.00476
R76609 VSS.n6015 VSS.n4436 0.00476
R76610 VSS.n6011 VSS.n4436 0.00476
R76611 VSS.n6011 VSS.n6010 0.00476
R76612 VSS.n6010 VSS.n6009 0.00476
R76613 VSS.n6005 VSS.n6004 0.00476
R76614 VSS.n6004 VSS.n6003 0.00476
R76615 VSS.n6003 VSS.n4448 0.00476
R76616 VSS.n5999 VSS.n4448 0.00476
R76617 VSS.n5999 VSS.n5998 0.00476
R76618 VSS.n5998 VSS.n4453 0.00476
R76619 VSS.n4875 VSS.n4453 0.00476
R76620 VSS.n4878 VSS.n4875 0.00476
R76621 VSS.n4878 VSS.n4872 0.00476
R76622 VSS.n4882 VSS.n4872 0.00476
R76623 VSS.n4882 VSS.n4870 0.00476
R76624 VSS.n4886 VSS.n4870 0.00476
R76625 VSS.n4886 VSS.n4868 0.00476
R76626 VSS.n4890 VSS.n4868 0.00476
R76627 VSS.n4890 VSS.n4866 0.00476
R76628 VSS.n4894 VSS.n4866 0.00476
R76629 VSS.n4894 VSS.n4864 0.00476
R76630 VSS.n4898 VSS.n4864 0.00476
R76631 VSS.n4898 VSS.n4862 0.00476
R76632 VSS.n4902 VSS.n4862 0.00476
R76633 VSS.n4902 VSS.n4860 0.00476
R76634 VSS.n5983 VSS.n4860 0.00476
R76635 VSS.n5983 VSS.n5982 0.00476
R76636 VSS.n5978 VSS.n5977 0.00476
R76637 VSS.n5977 VSS.n5976 0.00476
R76638 VSS.n5976 VSS.n5948 0.00476
R76639 VSS.n5972 VSS.n5948 0.00476
R76640 VSS.n5972 VSS.n5971 0.00476
R76641 VSS.n5971 VSS.n5970 0.00476
R76642 VSS.n5970 VSS.n5954 0.00476
R76643 VSS.n5966 VSS.n5954 0.00476
R76644 VSS.n5966 VSS.n5965 0.00476
R76645 VSS.n5965 VSS.n5964 0.00476
R76646 VSS.n5389 VSS.n5327 0.00476
R76647 VSS.n5393 VSS.n5327 0.00476
R76648 VSS.n5394 VSS.n5393 0.00476
R76649 VSS.n5397 VSS.n5394 0.00476
R76650 VSS.n5397 VSS.n5325 0.00476
R76651 VSS.n5401 VSS.n5325 0.00476
R76652 VSS.n5401 VSS.n5323 0.00476
R76653 VSS.n5405 VSS.n5323 0.00476
R76654 VSS.n5405 VSS.n5321 0.00476
R76655 VSS.n5409 VSS.n5321 0.00476
R76656 VSS.n5409 VSS.n5319 0.00476
R76657 VSS.n5413 VSS.n5319 0.00476
R76658 VSS.n5413 VSS.n5317 0.00476
R76659 VSS.n5418 VSS.n5317 0.00476
R76660 VSS.n5418 VSS.n5315 0.00476
R76661 VSS.n5422 VSS.n5315 0.00476
R76662 VSS.n5423 VSS.n5422 0.00476
R76663 VSS.n5423 VSS.n5313 0.00476
R76664 VSS.n5612 VSS.n5313 0.00476
R76665 VSS.n5612 VSS.n5611 0.00476
R76666 VSS.n5611 VSS.n5610 0.00476
R76667 VSS.n5610 VSS.n5429 0.00476
R76668 VSS.n5606 VSS.n5429 0.00476
R76669 VSS.n5602 VSS.n5435 0.00476
R76670 VSS.n5598 VSS.n5435 0.00476
R76671 VSS.n5598 VSS.n5597 0.00476
R76672 VSS.n5597 VSS.n5596 0.00476
R76673 VSS.n5596 VSS.n5440 0.00476
R76674 VSS.n5592 VSS.n5440 0.00476
R76675 VSS.n5592 VSS.n5591 0.00476
R76676 VSS.n5591 VSS.n5590 0.00476
R76677 VSS.n5590 VSS.n5446 0.00476
R76678 VSS.n5586 VSS.n5446 0.00476
R76679 VSS.n5586 VSS.n5585 0.00476
R76680 VSS.n5585 VSS.n5451 0.00476
R76681 VSS.n5571 VSS.n5451 0.00476
R76682 VSS.n5571 VSS.n5570 0.00476
R76683 VSS.n5570 VSS.n5569 0.00476
R76684 VSS.n5569 VSS.n5545 0.00476
R76685 VSS.n5565 VSS.n5545 0.00476
R76686 VSS.n5565 VSS.n5564 0.00476
R76687 VSS.n5564 VSS.n5563 0.00476
R76688 VSS.n5563 VSS.n5551 0.00476
R76689 VSS.n5559 VSS.n5551 0.00476
R76690 VSS.n5559 VSS.n5558 0.00476
R76691 VSS.n5558 VSS.n5557 0.00476
R76692 VSS.n5654 VSS.n5172 0.00476
R76693 VSS.n5650 VSS.n5172 0.00476
R76694 VSS.n5650 VSS.n5649 0.00476
R76695 VSS.n5649 VSS.n5648 0.00476
R76696 VSS.n5648 VSS.n5177 0.00476
R76697 VSS.n5251 VSS.n5177 0.00476
R76698 VSS.n5251 VSS.n5250 0.00476
R76699 VSS.n5250 VSS.n5249 0.00476
R76700 VSS.n5249 VSS.n5208 0.00476
R76701 VSS.n5245 VSS.n5208 0.00476
R76702 VSS.n5245 VSS.n5244 0.00476
R76703 VSS.n5244 VSS.n5243 0.00476
R76704 VSS.n5243 VSS.n5214 0.00476
R76705 VSS.n5239 VSS.n5214 0.00476
R76706 VSS.n5239 VSS.n5238 0.00476
R76707 VSS.n5238 VSS.n5237 0.00476
R76708 VSS.n5237 VSS.n5220 0.00476
R76709 VSS.n5233 VSS.n5220 0.00476
R76710 VSS.n5233 VSS.n5232 0.00476
R76711 VSS.n5232 VSS.n5231 0.00476
R76712 VSS.n5231 VSS.n5229 0.00476
R76713 VSS.n5229 VSS.n5228 0.00476
R76714 VSS.n5228 VSS.n4913 0.00476
R76715 VSS.n5941 VSS.n5907 0.00476
R76716 VSS.n5937 VSS.n5907 0.00476
R76717 VSS.n5937 VSS.n5936 0.00476
R76718 VSS.n5936 VSS.n5935 0.00476
R76719 VSS.n5935 VSS.n5912 0.00476
R76720 VSS.n5931 VSS.n5912 0.00476
R76721 VSS.n5931 VSS.n5930 0.00476
R76722 VSS.n5930 VSS.n5929 0.00476
R76723 VSS.n5929 VSS.n5918 0.00476
R76724 VSS.n5925 VSS.n5918 0.00476
R76725 VSS.n5925 VSS.n5924 0.00476
R76726 VSS.n5375 VSS.n5374 0.00476
R76727 VSS.n5374 VSS.n5373 0.00476
R76728 VSS.n5373 VSS.n5372 0.00476
R76729 VSS.n5372 VSS.n5334 0.00476
R76730 VSS.n5368 VSS.n5334 0.00476
R76731 VSS.n5368 VSS.n5367 0.00476
R76732 VSS.n5367 VSS.n5366 0.00476
R76733 VSS.n5366 VSS.n5340 0.00476
R76734 VSS.n5362 VSS.n5340 0.00476
R76735 VSS.n5362 VSS.n5361 0.00476
R76736 VSS.n5361 VSS.n5360 0.00476
R76737 VSS.n5360 VSS.n5346 0.00476
R76738 VSS.n5356 VSS.n5346 0.00476
R76739 VSS.n5356 VSS.n5355 0.00476
R76740 VSS.n5355 VSS.n5354 0.00476
R76741 VSS.n5354 VSS.n5122 0.00476
R76742 VSS.n5770 VSS.n5122 0.00476
R76743 VSS.n5770 VSS.n5769 0.00476
R76744 VSS.n5769 VSS.n5768 0.00476
R76745 VSS.n5768 VSS.n5767 0.00476
R76746 VSS.n5767 VSS.n5127 0.00476
R76747 VSS.n5763 VSS.n5127 0.00476
R76748 VSS.n5763 VSS.n5762 0.00476
R76749 VSS.n5760 VSS.n5133 0.00476
R76750 VSS.n5756 VSS.n5133 0.00476
R76751 VSS.n5756 VSS.n5755 0.00476
R76752 VSS.n5755 VSS.n5754 0.00476
R76753 VSS.n5754 VSS.n5140 0.00476
R76754 VSS.n5750 VSS.n5140 0.00476
R76755 VSS.n5750 VSS.n5749 0.00476
R76756 VSS.n5749 VSS.n5748 0.00476
R76757 VSS.n5748 VSS.n5146 0.00476
R76758 VSS.n5744 VSS.n5146 0.00476
R76759 VSS.n5744 VSS.n5743 0.00476
R76760 VSS.n5743 VSS.n5741 0.00476
R76761 VSS.n5741 VSS.n5740 0.00476
R76762 VSS.n5740 VSS.n5739 0.00476
R76763 VSS.n5739 VSS.n5153 0.00476
R76764 VSS.n5735 VSS.n5153 0.00476
R76765 VSS.n5735 VSS.n5734 0.00476
R76766 VSS.n5734 VSS.n5733 0.00476
R76767 VSS.n5733 VSS.n5159 0.00476
R76768 VSS.n5729 VSS.n5159 0.00476
R76769 VSS.n5729 VSS.n5728 0.00476
R76770 VSS.n5728 VSS.n5727 0.00476
R76771 VSS.n5727 VSS.n5165 0.00476
R76772 VSS.n5722 VSS.n5721 0.00476
R76773 VSS.n5721 VSS.n5720 0.00476
R76774 VSS.n5720 VSS.n5717 0.00476
R76775 VSS.n5717 VSS.n5716 0.00476
R76776 VSS.n5716 VSS.n5715 0.00476
R76777 VSS.n5715 VSS.n5714 0.00476
R76778 VSS.n5714 VSS.n5713 0.00476
R76779 VSS.n5713 VSS.n5667 0.00476
R76780 VSS.n5709 VSS.n5667 0.00476
R76781 VSS.n5709 VSS.n5708 0.00476
R76782 VSS.n5708 VSS.n5707 0.00476
R76783 VSS.n5707 VSS.n5673 0.00476
R76784 VSS.n5703 VSS.n5673 0.00476
R76785 VSS.n5703 VSS.n5702 0.00476
R76786 VSS.n5702 VSS.n5701 0.00476
R76787 VSS.n5701 VSS.n5679 0.00476
R76788 VSS.n5697 VSS.n5679 0.00476
R76789 VSS.n5697 VSS.n5696 0.00476
R76790 VSS.n5696 VSS.n5695 0.00476
R76791 VSS.n5695 VSS.n5685 0.00476
R76792 VSS.n5691 VSS.n5685 0.00476
R76793 VSS.n5691 VSS.n5690 0.00476
R76794 VSS.n5690 VSS.n4914 0.00476
R76795 VSS.n5904 VSS.n4916 0.00476
R76796 VSS.n5900 VSS.n4916 0.00476
R76797 VSS.n5900 VSS.n5899 0.00476
R76798 VSS.n5899 VSS.n5898 0.00476
R76799 VSS.n5898 VSS.n5876 0.00476
R76800 VSS.n5894 VSS.n5876 0.00476
R76801 VSS.n5894 VSS.n5893 0.00476
R76802 VSS.n5893 VSS.n5892 0.00476
R76803 VSS.n5892 VSS.n5882 0.00476
R76804 VSS.n5888 VSS.n5882 0.00476
R76805 VSS.n5371 VSS.n5007 0.00476
R76806 VSS.n5371 VSS.n5370 0.00476
R76807 VSS.n5370 VSS.n5369 0.00476
R76808 VSS.n5369 VSS.n5335 0.00476
R76809 VSS.n5365 VSS.n5335 0.00476
R76810 VSS.n5365 VSS.n5364 0.00476
R76811 VSS.n5364 VSS.n5363 0.00476
R76812 VSS.n5363 VSS.n5341 0.00476
R76813 VSS.n5359 VSS.n5341 0.00476
R76814 VSS.n5359 VSS.n5358 0.00476
R76815 VSS.n5358 VSS.n5357 0.00476
R76816 VSS.n5357 VSS.n5347 0.00476
R76817 VSS.n5353 VSS.n5347 0.00476
R76818 VSS.n5353 VSS.n5121 0.00476
R76819 VSS.n5771 VSS.n5121 0.00476
R76820 VSS.n5766 VSS.n5091 0.00476
R76821 VSS.n5766 VSS.n5765 0.00476
R76822 VSS.n5765 VSS.n5764 0.00476
R76823 VSS.n5764 VSS.n5128 0.00476
R76824 VSS.n5759 VSS.n5758 0.00476
R76825 VSS.n5758 VSS.n5757 0.00476
R76826 VSS.n5757 VSS.n5135 0.00476
R76827 VSS.n5753 VSS.n5135 0.00476
R76828 VSS.n5753 VSS.n5752 0.00476
R76829 VSS.n5752 VSS.n5751 0.00476
R76830 VSS.n5751 VSS.n5141 0.00476
R76831 VSS.n5747 VSS.n5141 0.00476
R76832 VSS.n5747 VSS.n5746 0.00476
R76833 VSS.n5746 VSS.n5745 0.00476
R76834 VSS.n5738 VSS.n5035 0.00476
R76835 VSS.n5738 VSS.n5737 0.00476
R76836 VSS.n5737 VSS.n5736 0.00476
R76837 VSS.n5736 VSS.n5154 0.00476
R76838 VSS.n5732 VSS.n5154 0.00476
R76839 VSS.n5732 VSS.n5731 0.00476
R76840 VSS.n5731 VSS.n5730 0.00476
R76841 VSS.n5730 VSS.n5160 0.00476
R76842 VSS.n5726 VSS.n5160 0.00476
R76843 VSS.n5726 VSS.n5725 0.00476
R76844 VSS.n5723 VSS.n5166 0.00476
R76845 VSS.n5719 VSS.n5166 0.00476
R76846 VSS.n5719 VSS.n5718 0.00476
R76847 VSS.n5718 VSS.n5070 0.00476
R76848 VSS.n5712 VSS.n5064 0.00476
R76849 VSS.n5712 VSS.n5711 0.00476
R76850 VSS.n5711 VSS.n5710 0.00476
R76851 VSS.n5710 VSS.n5668 0.00476
R76852 VSS.n5706 VSS.n5668 0.00476
R76853 VSS.n5706 VSS.n5705 0.00476
R76854 VSS.n5705 VSS.n5704 0.00476
R76855 VSS.n5704 VSS.n5674 0.00476
R76856 VSS.n5700 VSS.n5674 0.00476
R76857 VSS.n5700 VSS.n5699 0.00476
R76858 VSS.n5699 VSS.n5698 0.00476
R76859 VSS.n5698 VSS.n5680 0.00476
R76860 VSS.n5694 VSS.n5680 0.00476
R76861 VSS.n5694 VSS.n5693 0.00476
R76862 VSS.n5693 VSS.n5692 0.00476
R76863 VSS.n5903 VSS.n5902 0.00476
R76864 VSS.n5902 VSS.n5901 0.00476
R76865 VSS.n5901 VSS.n5871 0.00476
R76866 VSS.n5897 VSS.n5871 0.00476
R76867 VSS.n5897 VSS.n5896 0.00476
R76868 VSS.n5896 VSS.n5895 0.00476
R76869 VSS.n5895 VSS.n5877 0.00476
R76870 VSS.n5891 VSS.n5877 0.00476
R76871 VSS.n5891 VSS.n5890 0.00476
R76872 VSS.n5890 VSS.n5889 0.00476
R76873 VSS.n5395 VSS.n5270 0.00476
R76874 VSS.n5396 VSS.n5395 0.00476
R76875 VSS.n5396 VSS.n5324 0.00476
R76876 VSS.n5402 VSS.n5324 0.00476
R76877 VSS.n5403 VSS.n5402 0.00476
R76878 VSS.n5404 VSS.n5403 0.00476
R76879 VSS.n5404 VSS.n5320 0.00476
R76880 VSS.n5410 VSS.n5320 0.00476
R76881 VSS.n5411 VSS.n5410 0.00476
R76882 VSS.n5412 VSS.n5411 0.00476
R76883 VSS.n5412 VSS.n5316 0.00476
R76884 VSS.n5419 VSS.n5316 0.00476
R76885 VSS.n5420 VSS.n5419 0.00476
R76886 VSS.n5421 VSS.n5420 0.00476
R76887 VSS.n5421 VSS.n5289 0.00476
R76888 VSS.n5613 VSS.n5312 0.00476
R76889 VSS.n5609 VSS.n5312 0.00476
R76890 VSS.n5609 VSS.n5608 0.00476
R76891 VSS.n5608 VSS.n5607 0.00476
R76892 VSS.n5601 VSS.n5600 0.00476
R76893 VSS.n5600 VSS.n5599 0.00476
R76894 VSS.n5599 VSS.n5436 0.00476
R76895 VSS.n5595 VSS.n5436 0.00476
R76896 VSS.n5595 VSS.n5594 0.00476
R76897 VSS.n5594 VSS.n5593 0.00476
R76898 VSS.n5593 VSS.n5441 0.00476
R76899 VSS.n5589 VSS.n5441 0.00476
R76900 VSS.n5589 VSS.n5588 0.00476
R76901 VSS.n5588 VSS.n5587 0.00476
R76902 VSS.n5572 VSS.n5540 0.00476
R76903 VSS.n5568 VSS.n5540 0.00476
R76904 VSS.n5568 VSS.n5567 0.00476
R76905 VSS.n5567 VSS.n5566 0.00476
R76906 VSS.n5566 VSS.n5546 0.00476
R76907 VSS.n5562 VSS.n5546 0.00476
R76908 VSS.n5562 VSS.n5561 0.00476
R76909 VSS.n5561 VSS.n5560 0.00476
R76910 VSS.n5560 VSS.n5552 0.00476
R76911 VSS.n5556 VSS.n5552 0.00476
R76912 VSS.n5653 VSS.n5652 0.00476
R76913 VSS.n5652 VSS.n5651 0.00476
R76914 VSS.n5651 VSS.n5173 0.00476
R76915 VSS.n5647 VSS.n5173 0.00476
R76916 VSS.n5252 VSS.n5203 0.00476
R76917 VSS.n5248 VSS.n5203 0.00476
R76918 VSS.n5248 VSS.n5247 0.00476
R76919 VSS.n5247 VSS.n5246 0.00476
R76920 VSS.n5246 VSS.n5209 0.00476
R76921 VSS.n5242 VSS.n5209 0.00476
R76922 VSS.n5242 VSS.n5241 0.00476
R76923 VSS.n5241 VSS.n5240 0.00476
R76924 VSS.n5240 VSS.n5215 0.00476
R76925 VSS.n5236 VSS.n5215 0.00476
R76926 VSS.n5236 VSS.n5235 0.00476
R76927 VSS.n5235 VSS.n5234 0.00476
R76928 VSS.n5234 VSS.n5221 0.00476
R76929 VSS.n5230 VSS.n5221 0.00476
R76930 VSS.n5230 VSS.n4948 0.00476
R76931 VSS.n5940 VSS.n5939 0.00476
R76932 VSS.n5939 VSS.n5938 0.00476
R76933 VSS.n5938 VSS.n5908 0.00476
R76934 VSS.n5934 VSS.n5908 0.00476
R76935 VSS.n5934 VSS.n5933 0.00476
R76936 VSS.n5933 VSS.n5932 0.00476
R76937 VSS.n5932 VSS.n5913 0.00476
R76938 VSS.n5928 VSS.n5913 0.00476
R76939 VSS.n5928 VSS.n5927 0.00476
R76940 VSS.n5927 VSS.n5926 0.00476
R76941 VSS.n5926 VSS.n5919 0.00476
R76942 VSS.n6085 VSS.n4333 0.00476
R76943 VSS.n6081 VSS.n4333 0.00476
R76944 VSS.n6081 VSS.n6080 0.00476
R76945 VSS.n6080 VSS.n6079 0.00476
R76946 VSS.n6079 VSS.n4339 0.00476
R76947 VSS.n6075 VSS.n4339 0.00476
R76948 VSS.n6075 VSS.n6074 0.00476
R76949 VSS.n6074 VSS.n6073 0.00476
R76950 VSS.n6073 VSS.n4345 0.00476
R76951 VSS.n6069 VSS.n4345 0.00476
R76952 VSS.n6069 VSS.n6068 0.00476
R76953 VSS.n6068 VSS.n6067 0.00476
R76954 VSS.n6067 VSS.n4351 0.00476
R76955 VSS.n6063 VSS.n4351 0.00476
R76956 VSS.n6063 VSS.n4294 0.00476
R76957 VSS.n6058 VSS.n4287 0.00476
R76958 VSS.n6058 VSS.n6057 0.00476
R76959 VSS.n6057 VSS.n6056 0.00476
R76960 VSS.n6056 VSS.n4361 0.00476
R76961 VSS.n6051 VSS.n6050 0.00476
R76962 VSS.n6050 VSS.n6049 0.00476
R76963 VSS.n6049 VSS.n4369 0.00476
R76964 VSS.n6045 VSS.n4369 0.00476
R76965 VSS.n6045 VSS.n6044 0.00476
R76966 VSS.n6044 VSS.n6043 0.00476
R76967 VSS.n6043 VSS.n4375 0.00476
R76968 VSS.n6039 VSS.n4375 0.00476
R76969 VSS.n6039 VSS.n6038 0.00476
R76970 VSS.n6038 VSS.n6037 0.00476
R76971 VSS.n6024 VSS.n4425 0.00476
R76972 VSS.n6020 VSS.n4425 0.00476
R76973 VSS.n6020 VSS.n6019 0.00476
R76974 VSS.n6019 VSS.n6018 0.00476
R76975 VSS.n6018 VSS.n4431 0.00476
R76976 VSS.n6014 VSS.n4431 0.00476
R76977 VSS.n6014 VSS.n6013 0.00476
R76978 VSS.n6013 VSS.n6012 0.00476
R76979 VSS.n6012 VSS.n4437 0.00476
R76980 VSS.n6008 VSS.n4437 0.00476
R76981 VSS.n6006 VSS.n4444 0.00476
R76982 VSS.n6002 VSS.n4444 0.00476
R76983 VSS.n6002 VSS.n6001 0.00476
R76984 VSS.n6001 VSS.n6000 0.00476
R76985 VSS.n4876 VSS.n4460 0.00476
R76986 VSS.n4877 VSS.n4876 0.00476
R76987 VSS.n4877 VSS.n4871 0.00476
R76988 VSS.n4883 VSS.n4871 0.00476
R76989 VSS.n4884 VSS.n4883 0.00476
R76990 VSS.n4885 VSS.n4884 0.00476
R76991 VSS.n4885 VSS.n4867 0.00476
R76992 VSS.n4891 VSS.n4867 0.00476
R76993 VSS.n4892 VSS.n4891 0.00476
R76994 VSS.n4893 VSS.n4892 0.00476
R76995 VSS.n4893 VSS.n4863 0.00476
R76996 VSS.n4899 VSS.n4863 0.00476
R76997 VSS.n4900 VSS.n4899 0.00476
R76998 VSS.n4901 VSS.n4900 0.00476
R76999 VSS.n4901 VSS.n4474 0.00476
R77000 VSS.n5979 VSS.n4909 0.00476
R77001 VSS.n5975 VSS.n4909 0.00476
R77002 VSS.n5975 VSS.n5974 0.00476
R77003 VSS.n5974 VSS.n5973 0.00476
R77004 VSS.n5973 VSS.n5949 0.00476
R77005 VSS.n5969 VSS.n5949 0.00476
R77006 VSS.n5969 VSS.n5968 0.00476
R77007 VSS.n5968 VSS.n5967 0.00476
R77008 VSS.n5967 VSS.n5955 0.00476
R77009 VSS.n5963 VSS.n5955 0.00476
R77010 VSS.n6448 VSS.n18 0.00468605
R77011 VSS.n3210 DVSS 0.00464676
R77012 VSS.n2486 DVSS 0.00460473
R77013 VSS.n5888 DVSS 0.00458
R77014 VSS.n5889 DVSS 0.00458
R77015 VSS.n3637 VSS.n3625 0.00455
R77016 VSS.n5797 VSS.n5070 0.00455
R77017 VSS.n5647 VSS.n5646 0.00455
R77018 VSS.n6000 VSS.n4449 0.00455
R77019 VSS.n1881 VSS.n1880 0.00455
R77020 VSS.n1744 VSS.n1743 0.00455
R77021 VSS.n1615 VSS.n1347 0.00455
R77022 VSS.n1605 VSS.n1604 0.00455
R77023 VSS.n5604 VSS.n5432 0.0045
R77024 VSS.n5656 VSS.n5168 0.0045
R77025 VSS.n5377 VSS.n5328 0.0045
R77026 VSS.n5604 VSS.n5433 0.0045
R77027 VSS.n5658 VSS.n5656 0.0045
R77028 VSS.n5944 VSS.n5943 0.0045
R77029 VSS.n5943 VSS.n4910 0.0045
R77030 VSS.n5383 VSS.n5328 0.0045
R77031 VSS.n6229 VSS.n6225 0.00448437
R77032 VSS.n3541 VSS.n963 0.00443
R77033 VSS.n5784 VSS.n5091 0.00443
R77034 VSS.n5619 VSS.n5613 0.00443
R77035 VSS.n6107 VSS.n4287 0.00443
R77036 VSS.n1594 VSS.n1549 0.00437324
R77037 VSS.n6149 VSS.n483 0.00419403
R77038 VSS.n5110 VSS.n5031 0.00419403
R77039 VSS.n1120 VSS.n1092 0.0041
R77040 VSS.n1121 VSS.n1083 0.0041
R77041 VSS.n2963 VSS.n1091 0.0041
R77042 VSS.n2928 VSS.n1156 0.0041
R77043 VSS.n1159 VSS.n1158 0.0041
R77044 VSS.n2926 VSS.n2925 0.0041
R77045 VSS.n1836 VSS.n1236 0.00409155
R77046 VSS.n5978 VSS.n4907 0.00404
R77047 VSS.n5941 VSS.n5906 0.00404
R77048 VSS.n5905 VSS.n5904 0.00404
R77049 VSS.n5903 VSS.n5870 0.00404
R77050 VSS.n5940 VSS.n4908 0.00404
R77051 VSS.n5980 VSS.n5979 0.00404
R77052 VSS.n1906 VSS.n1200 0.00403571
R77053 VSS.n2055 VSS.n1186 0.00403571
R77054 VSS.n2688 VSS.n2687 0.00403571
R77055 VSS.n2203 VSS.n2151 0.00403571
R77056 VSS.n6129 VSS.n4251 0.00403571
R77057 VSS.n3591 VSS.n911 0.00401
R77058 VSS.n3640 VSS.n881 0.00401
R77059 VSS.n5825 VSS.n5029 0.00401
R77060 VSS.n5804 VSS.n5054 0.00401
R77061 VSS.n5578 VSS.n5505 0.00401
R77062 VSS.n5643 VSS.n5186 0.00401
R77063 VSS.n6031 VSS.n4422 0.00401
R77064 VSS.n5997 VSS.n5996 0.00401
R77065 VSS.n3692 DVSS 0.00392
R77066 VSS.n3693 DVSS 0.00392
R77067 VSS.n5964 DVSS 0.00392
R77068 VSS.n5963 DVSS 0.00392
R77069 VSS.n2623 VSS.n674 0.00391292
R77070 VSS.n803 VSS.n793 0.00391292
R77071 VSS.n3534 VSS.n3533 0.00389
R77072 VSS.n3576 VSS.n947 0.00389
R77073 VSS.n5781 VSS.n5082 0.00389
R77074 VSS.n5742 VSS.n5027 0.00389
R77075 VSS.n5622 VSS.n5297 0.00389
R77076 VSS.n5584 VSS.n5447 0.00389
R77077 VSS.n6104 VSS.n4280 0.00389
R77078 VSS.n6034 VSS.n4381 0.00389
R77079 VSS.n6005 VSS.n4442 0.0038
R77080 VSS.n5654 VSS.n5171 0.0038
R77081 VSS.n5722 VSS.n5167 0.0038
R77082 VSS.n5724 VSS.n5723 0.0038
R77083 VSS.n5653 VSS.n4443 0.0038
R77084 VSS.n6007 VSS.n6006 0.0038
R77085 VSS.n1830 VSS.n1250 0.00377857
R77086 VSS.n3064 VSS.n3063 0.00377857
R77087 VSS.n3403 VSS.n1003 0.00377857
R77088 VSS.n4089 VSS.n4088 0.00377857
R77089 VSS.n491 VSS.n489 0.00377857
R77090 VSS.n6053 VSS.n6052 0.00356
R77091 VSS.n5602 VSS.n4365 0.00356
R77092 VSS.n5761 VSS.n5760 0.00356
R77093 VSS.n5759 VSS.n5134 0.00356
R77094 VSS.n5601 VSS.n5430 0.00356
R77095 VSS.n6051 VSS.n4368 0.00356
R77096 DVSS VSS.n763 0.00353371
R77097 VSS.n4825 VSS.n4387 0.00352239
R77098 VSS.n5537 VSS.n5536 0.00352239
R77099 VSS.n6215 VSS.n6214 0.00346697
R77100 VSS.n2093 VSS.n2092 0.00334
R77101 VSS.n2096 VSS.n2093 0.00334
R77102 VSS.n2097 VSS.n2096 0.00334
R77103 VSS.n2098 VSS.n2097 0.00334
R77104 VSS.n2099 VSS.n2098 0.00334
R77105 VSS.n2102 VSS.n2099 0.00334
R77106 VSS.n2103 VSS.n2102 0.00334
R77107 VSS.n2104 VSS.n2103 0.00334
R77108 VSS.n2105 VSS.n2104 0.00334
R77109 VSS.n2108 VSS.n2105 0.00334
R77110 VSS.n2109 VSS.n2108 0.00334
R77111 VSS.n2110 VSS.n2109 0.00334
R77112 VSS.n2111 VSS.n2110 0.00334
R77113 VSS.n2111 VSS.n965 0.00334
R77114 VSS.n3537 VSS.n965 0.00334
R77115 VSS.n3538 VSS.n3537 0.00334
R77116 VSS.n3539 VSS.n3538 0.00334
R77117 VSS.n3539 VSS.n961 0.00334
R77118 VSS.n3545 VSS.n961 0.00334
R77119 VSS.n3546 VSS.n3545 0.00334
R77120 VSS.n3547 VSS.n3546 0.00334
R77121 VSS.n3547 VSS.n957 0.00334
R77122 VSS.n3553 VSS.n957 0.00334
R77123 VSS.n3554 VSS.n3553 0.00334
R77124 VSS.n3555 VSS.n3554 0.00334
R77125 VSS.n3555 VSS.n953 0.00334
R77126 VSS.n3561 VSS.n953 0.00334
R77127 VSS.n3562 VSS.n3561 0.00334
R77128 VSS.n3563 VSS.n3562 0.00334
R77129 VSS.n3563 VSS.n949 0.00334
R77130 VSS.n3570 VSS.n949 0.00334
R77131 VSS.n3571 VSS.n3570 0.00334
R77132 VSS.n3572 VSS.n3571 0.00334
R77133 VSS.n3573 VSS.n3572 0.00334
R77134 VSS.n3573 VSS.n909 0.00334
R77135 VSS.n3595 VSS.n909 0.00334
R77136 VSS.n3596 VSS.n3595 0.00334
R77137 VSS.n3597 VSS.n3596 0.00334
R77138 VSS.n3597 VSS.n905 0.00334
R77139 VSS.n3603 VSS.n905 0.00334
R77140 VSS.n3604 VSS.n3603 0.00334
R77141 VSS.n3605 VSS.n3604 0.00334
R77142 VSS.n3605 VSS.n901 0.00334
R77143 VSS.n3611 VSS.n901 0.00334
R77144 VSS.n3612 VSS.n3611 0.00334
R77145 VSS.n3613 VSS.n3612 0.00334
R77146 VSS.n3613 VSS.n897 0.00334
R77147 VSS.n3619 VSS.n897 0.00334
R77148 VSS.n3620 VSS.n3619 0.00334
R77149 VSS.n3621 VSS.n3620 0.00334
R77150 VSS.n3622 VSS.n3621 0.00334
R77151 VSS.n3622 VSS.n879 0.00334
R77152 VSS.n3644 VSS.n879 0.00334
R77153 VSS.n3645 VSS.n3644 0.00334
R77154 VSS.n3646 VSS.n3645 0.00334
R77155 VSS.n3646 VSS.n875 0.00334
R77156 VSS.n3652 VSS.n875 0.00334
R77157 VSS.n3653 VSS.n3652 0.00334
R77158 VSS.n3654 VSS.n3653 0.00334
R77159 VSS.n3654 VSS.n871 0.00334
R77160 VSS.n3660 VSS.n871 0.00334
R77161 VSS.n3661 VSS.n3660 0.00334
R77162 VSS.n3662 VSS.n3661 0.00334
R77163 VSS.n3662 VSS.n867 0.00334
R77164 VSS.n3668 VSS.n867 0.00334
R77165 VSS.n3669 VSS.n3668 0.00334
R77166 VSS.n3670 VSS.n3669 0.00334
R77167 VSS.n3671 VSS.n3670 0.00334
R77168 VSS.n3672 VSS.n3671 0.00334
R77169 VSS.n3673 VSS.n3672 0.00334
R77170 VSS.n3676 VSS.n3673 0.00334
R77171 VSS.n3677 VSS.n3676 0.00334
R77172 VSS.n3678 VSS.n3677 0.00334
R77173 VSS.n3679 VSS.n3678 0.00334
R77174 VSS.n3682 VSS.n3679 0.00334
R77175 VSS.n3683 VSS.n3682 0.00334
R77176 VSS.n3684 VSS.n3683 0.00334
R77177 VSS.n3685 VSS.n3684 0.00334
R77178 VSS.n3687 VSS.n3685 0.00334
R77179 VSS.n3688 VSS.n3687 0.00334
R77180 VSS.n3689 VSS.n3688 0.00334
R77181 VSS.n5376 VSS.n5331 0.00334
R77182 VSS.n5332 VSS.n5331 0.00334
R77183 VSS.n5333 VSS.n5332 0.00334
R77184 VSS.n5336 VSS.n5333 0.00334
R77185 VSS.n5337 VSS.n5336 0.00334
R77186 VSS.n5338 VSS.n5337 0.00334
R77187 VSS.n5339 VSS.n5338 0.00334
R77188 VSS.n5342 VSS.n5339 0.00334
R77189 VSS.n5343 VSS.n5342 0.00334
R77190 VSS.n5344 VSS.n5343 0.00334
R77191 VSS.n5345 VSS.n5344 0.00334
R77192 VSS.n5348 VSS.n5345 0.00334
R77193 VSS.n5349 VSS.n5348 0.00334
R77194 VSS.n5350 VSS.n5349 0.00334
R77195 VSS.n5352 VSS.n5350 0.00334
R77196 VSS.n5352 VSS.n5351 0.00334
R77197 VSS.n5351 VSS.n5123 0.00334
R77198 VSS.n5124 VSS.n5123 0.00334
R77199 VSS.n5125 VSS.n5124 0.00334
R77200 VSS.n5126 VSS.n5125 0.00334
R77201 VSS.n5129 VSS.n5126 0.00334
R77202 VSS.n5130 VSS.n5129 0.00334
R77203 VSS.n5131 VSS.n5130 0.00334
R77204 VSS.n5136 VSS.n5132 0.00334
R77205 VSS.n5137 VSS.n5136 0.00334
R77206 VSS.n5138 VSS.n5137 0.00334
R77207 VSS.n5139 VSS.n5138 0.00334
R77208 VSS.n5142 VSS.n5139 0.00334
R77209 VSS.n5143 VSS.n5142 0.00334
R77210 VSS.n5144 VSS.n5143 0.00334
R77211 VSS.n5145 VSS.n5144 0.00334
R77212 VSS.n5147 VSS.n5145 0.00334
R77213 VSS.n5148 VSS.n5147 0.00334
R77214 VSS.n5149 VSS.n5148 0.00334
R77215 VSS.n5150 VSS.n5149 0.00334
R77216 VSS.n5151 VSS.n5150 0.00334
R77217 VSS.n5152 VSS.n5151 0.00334
R77218 VSS.n5155 VSS.n5152 0.00334
R77219 VSS.n5156 VSS.n5155 0.00334
R77220 VSS.n5157 VSS.n5156 0.00334
R77221 VSS.n5158 VSS.n5157 0.00334
R77222 VSS.n5161 VSS.n5158 0.00334
R77223 VSS.n5162 VSS.n5161 0.00334
R77224 VSS.n5163 VSS.n5162 0.00334
R77225 VSS.n5164 VSS.n5163 0.00334
R77226 VSS.n5657 VSS.n5164 0.00334
R77227 VSS.n5660 VSS.n5659 0.00334
R77228 VSS.n5661 VSS.n5660 0.00334
R77229 VSS.n5662 VSS.n5661 0.00334
R77230 VSS.n5663 VSS.n5662 0.00334
R77231 VSS.n5664 VSS.n5663 0.00334
R77232 VSS.n5665 VSS.n5664 0.00334
R77233 VSS.n5666 VSS.n5665 0.00334
R77234 VSS.n5669 VSS.n5666 0.00334
R77235 VSS.n5670 VSS.n5669 0.00334
R77236 VSS.n5671 VSS.n5670 0.00334
R77237 VSS.n5672 VSS.n5671 0.00334
R77238 VSS.n5675 VSS.n5672 0.00334
R77239 VSS.n5676 VSS.n5675 0.00334
R77240 VSS.n5677 VSS.n5676 0.00334
R77241 VSS.n5678 VSS.n5677 0.00334
R77242 VSS.n5681 VSS.n5678 0.00334
R77243 VSS.n5682 VSS.n5681 0.00334
R77244 VSS.n5683 VSS.n5682 0.00334
R77245 VSS.n5684 VSS.n5683 0.00334
R77246 VSS.n5686 VSS.n5684 0.00334
R77247 VSS.n5687 VSS.n5686 0.00334
R77248 VSS.n5689 VSS.n5687 0.00334
R77249 VSS.n5689 VSS.n5688 0.00334
R77250 VSS.n5872 VSS.n4915 0.00334
R77251 VSS.n5873 VSS.n5872 0.00334
R77252 VSS.n5874 VSS.n5873 0.00334
R77253 VSS.n5875 VSS.n5874 0.00334
R77254 VSS.n5878 VSS.n5875 0.00334
R77255 VSS.n5879 VSS.n5878 0.00334
R77256 VSS.n5880 VSS.n5879 0.00334
R77257 VSS.n5881 VSS.n5880 0.00334
R77258 VSS.n5883 VSS.n5881 0.00334
R77259 VSS.n5884 VSS.n5883 0.00334
R77260 VSS.n5885 VSS.n5884 0.00334
R77261 VSS.n5391 VSS.n5390 0.00334
R77262 VSS.n5392 VSS.n5391 0.00334
R77263 VSS.n5392 VSS.n5326 0.00334
R77264 VSS.n5398 VSS.n5326 0.00334
R77265 VSS.n5399 VSS.n5398 0.00334
R77266 VSS.n5400 VSS.n5399 0.00334
R77267 VSS.n5400 VSS.n5322 0.00334
R77268 VSS.n5406 VSS.n5322 0.00334
R77269 VSS.n5407 VSS.n5406 0.00334
R77270 VSS.n5408 VSS.n5407 0.00334
R77271 VSS.n5408 VSS.n5318 0.00334
R77272 VSS.n5414 VSS.n5318 0.00334
R77273 VSS.n5415 VSS.n5414 0.00334
R77274 VSS.n5417 VSS.n5415 0.00334
R77275 VSS.n5417 VSS.n5416 0.00334
R77276 VSS.n5416 VSS.n5314 0.00334
R77277 VSS.n5424 VSS.n5314 0.00334
R77278 VSS.n5425 VSS.n5424 0.00334
R77279 VSS.n5426 VSS.n5425 0.00334
R77280 VSS.n5427 VSS.n5426 0.00334
R77281 VSS.n5428 VSS.n5427 0.00334
R77282 VSS.n5431 VSS.n5428 0.00334
R77283 VSS.n5605 VSS.n5431 0.00334
R77284 VSS.n5603 VSS.n5434 0.00334
R77285 VSS.n5437 VSS.n5434 0.00334
R77286 VSS.n5438 VSS.n5437 0.00334
R77287 VSS.n5439 VSS.n5438 0.00334
R77288 VSS.n5442 VSS.n5439 0.00334
R77289 VSS.n5443 VSS.n5442 0.00334
R77290 VSS.n5444 VSS.n5443 0.00334
R77291 VSS.n5445 VSS.n5444 0.00334
R77292 VSS.n5448 VSS.n5445 0.00334
R77293 VSS.n5449 VSS.n5448 0.00334
R77294 VSS.n5450 VSS.n5449 0.00334
R77295 VSS.n5541 VSS.n5450 0.00334
R77296 VSS.n5542 VSS.n5541 0.00334
R77297 VSS.n5543 VSS.n5542 0.00334
R77298 VSS.n5544 VSS.n5543 0.00334
R77299 VSS.n5547 VSS.n5544 0.00334
R77300 VSS.n5548 VSS.n5547 0.00334
R77301 VSS.n5549 VSS.n5548 0.00334
R77302 VSS.n5550 VSS.n5549 0.00334
R77303 VSS.n5553 VSS.n5550 0.00334
R77304 VSS.n5554 VSS.n5553 0.00334
R77305 VSS.n5555 VSS.n5554 0.00334
R77306 VSS.n5555 VSS.n5169 0.00334
R77307 VSS.n5655 VSS.n5170 0.00334
R77308 VSS.n5174 VSS.n5170 0.00334
R77309 VSS.n5175 VSS.n5174 0.00334
R77310 VSS.n5176 VSS.n5175 0.00334
R77311 VSS.n5204 VSS.n5176 0.00334
R77312 VSS.n5205 VSS.n5204 0.00334
R77313 VSS.n5206 VSS.n5205 0.00334
R77314 VSS.n5207 VSS.n5206 0.00334
R77315 VSS.n5210 VSS.n5207 0.00334
R77316 VSS.n5211 VSS.n5210 0.00334
R77317 VSS.n5212 VSS.n5211 0.00334
R77318 VSS.n5213 VSS.n5212 0.00334
R77319 VSS.n5216 VSS.n5213 0.00334
R77320 VSS.n5217 VSS.n5216 0.00334
R77321 VSS.n5218 VSS.n5217 0.00334
R77322 VSS.n5219 VSS.n5218 0.00334
R77323 VSS.n5222 VSS.n5219 0.00334
R77324 VSS.n5223 VSS.n5222 0.00334
R77325 VSS.n5224 VSS.n5223 0.00334
R77326 VSS.n5225 VSS.n5224 0.00334
R77327 VSS.n5226 VSS.n5225 0.00334
R77328 VSS.n5227 VSS.n5226 0.00334
R77329 VSS.n5227 VSS.n4911 0.00334
R77330 VSS.n5942 VSS.n4912 0.00334
R77331 VSS.n5909 VSS.n4912 0.00334
R77332 VSS.n5910 VSS.n5909 0.00334
R77333 VSS.n5911 VSS.n5910 0.00334
R77334 VSS.n5914 VSS.n5911 0.00334
R77335 VSS.n5915 VSS.n5914 0.00334
R77336 VSS.n5916 VSS.n5915 0.00334
R77337 VSS.n5917 VSS.n5916 0.00334
R77338 VSS.n5920 VSS.n5917 0.00334
R77339 VSS.n5921 VSS.n5920 0.00334
R77340 VSS.n5922 VSS.n5921 0.00334
R77341 VSS.n5382 VSS.n5380 0.00334
R77342 VSS.n5380 VSS.n4335 0.00334
R77343 VSS.n4336 VSS.n4335 0.00334
R77344 VSS.n4337 VSS.n4336 0.00334
R77345 VSS.n4340 VSS.n4337 0.00334
R77346 VSS.n4341 VSS.n4340 0.00334
R77347 VSS.n4342 VSS.n4341 0.00334
R77348 VSS.n4343 VSS.n4342 0.00334
R77349 VSS.n4346 VSS.n4343 0.00334
R77350 VSS.n4347 VSS.n4346 0.00334
R77351 VSS.n4348 VSS.n4347 0.00334
R77352 VSS.n4349 VSS.n4348 0.00334
R77353 VSS.n4352 VSS.n4349 0.00334
R77354 VSS.n4353 VSS.n4352 0.00334
R77355 VSS.n4354 VSS.n4353 0.00334
R77356 VSS.n4355 VSS.n4354 0.00334
R77357 VSS.n4356 VSS.n4355 0.00334
R77358 VSS.n4357 VSS.n4356 0.00334
R77359 VSS.n4358 VSS.n4357 0.00334
R77360 VSS.n4359 VSS.n4358 0.00334
R77361 VSS.n4362 VSS.n4359 0.00334
R77362 VSS.n4363 VSS.n4362 0.00334
R77363 VSS.n4364 VSS.n4363 0.00334
R77364 VSS.n4370 VSS.n4366 0.00334
R77365 VSS.n4371 VSS.n4370 0.00334
R77366 VSS.n4372 VSS.n4371 0.00334
R77367 VSS.n4373 VSS.n4372 0.00334
R77368 VSS.n4376 VSS.n4373 0.00334
R77369 VSS.n4377 VSS.n4376 0.00334
R77370 VSS.n4378 VSS.n4377 0.00334
R77371 VSS.n4379 VSS.n4378 0.00334
R77372 VSS.n4382 VSS.n4379 0.00334
R77373 VSS.n4383 VSS.n4382 0.00334
R77374 VSS.n4384 VSS.n4383 0.00334
R77375 VSS.n4426 VSS.n4384 0.00334
R77376 VSS.n4427 VSS.n4426 0.00334
R77377 VSS.n4428 VSS.n4427 0.00334
R77378 VSS.n4429 VSS.n4428 0.00334
R77379 VSS.n4432 VSS.n4429 0.00334
R77380 VSS.n4433 VSS.n4432 0.00334
R77381 VSS.n4434 VSS.n4433 0.00334
R77382 VSS.n4435 VSS.n4434 0.00334
R77383 VSS.n4438 VSS.n4435 0.00334
R77384 VSS.n4439 VSS.n4438 0.00334
R77385 VSS.n4440 VSS.n4439 0.00334
R77386 VSS.n4441 VSS.n4440 0.00334
R77387 VSS.n4446 VSS.n4445 0.00334
R77388 VSS.n4447 VSS.n4446 0.00334
R77389 VSS.n4450 VSS.n4447 0.00334
R77390 VSS.n4451 VSS.n4450 0.00334
R77391 VSS.n4452 VSS.n4451 0.00334
R77392 VSS.n4873 VSS.n4452 0.00334
R77393 VSS.n4874 VSS.n4873 0.00334
R77394 VSS.n4879 VSS.n4874 0.00334
R77395 VSS.n4880 VSS.n4879 0.00334
R77396 VSS.n4881 VSS.n4880 0.00334
R77397 VSS.n4881 VSS.n4869 0.00334
R77398 VSS.n4887 VSS.n4869 0.00334
R77399 VSS.n4888 VSS.n4887 0.00334
R77400 VSS.n4889 VSS.n4888 0.00334
R77401 VSS.n4889 VSS.n4865 0.00334
R77402 VSS.n4895 VSS.n4865 0.00334
R77403 VSS.n4896 VSS.n4895 0.00334
R77404 VSS.n4897 VSS.n4896 0.00334
R77405 VSS.n4897 VSS.n4861 0.00334
R77406 VSS.n4903 VSS.n4861 0.00334
R77407 VSS.n4904 VSS.n4903 0.00334
R77408 VSS.n4905 VSS.n4904 0.00334
R77409 VSS.n4906 VSS.n4905 0.00334
R77410 VSS.n5946 VSS.n5945 0.00334
R77411 VSS.n5947 VSS.n5946 0.00334
R77412 VSS.n5950 VSS.n5947 0.00334
R77413 VSS.n5951 VSS.n5950 0.00334
R77414 VSS.n5952 VSS.n5951 0.00334
R77415 VSS.n5953 VSS.n5952 0.00334
R77416 VSS.n5956 VSS.n5953 0.00334
R77417 VSS.n5957 VSS.n5956 0.00334
R77418 VSS.n5958 VSS.n5957 0.00334
R77419 VSS.n5959 VSS.n5958 0.00334
R77420 VSS.n5960 VSS.n5959 0.00334
R77421 VSS.n5381 VSS.n5330 0.00332
R77422 VSS.n5389 VSS.n5388 0.00332
R77423 VSS.n5375 VSS.n5329 0.00332
R77424 VSS.n5379 VSS.n4982 0.00332
R77425 VSS.n5386 VSS.n5274 0.00332
R77426 VSS.n5385 VSS.n4311 0.00332
R77427 VSS.n3723 VSS.n3712 0.00323
R77428 VSS.n5692 VSS.n4943 0.00323
R77429 VSS.n5855 VSS.n4948 0.00323
R77430 VSS.n5985 VSS.n4474 0.00323
R77431 VSS.n6142 VSS.n6140 0.0032
R77432 VSS.n5255 VSS.n4966 0.0032
R77433 VSS.n5078 VSS.n4927 0.0032
R77434 VSS.n6145 VSS.n486 0.0032
R77435 VSS.n5639 VSS.n5196 0.0032
R77436 VSS.n5792 VSS.n5063 0.0032
R77437 VSS.n6124 VSS.n6122 0.0032
R77438 VSS.n5306 VSS.n5257 0.0032
R77439 VSS.n5786 VSS.n5785 0.0032
R77440 VSS.n6128 VSS.n4259 0.0032
R77441 VSS.n5634 VSS.n5633 0.0032
R77442 VSS.n5787 VSS.n5006 0.0032
R77443 VSS.n2148 VSS.n2080 0.00311
R77444 VSS.n5840 VSS.n5007 0.00311
R77445 VSS.n5632 VSS.n5270 0.00311
R77446 VSS.n6095 VSS.n6085 0.00311
R77447 VSS.n4915 VSS.n4910 0.00286
R77448 VSS.n5943 VSS.n5942 0.00286
R77449 VSS.n5945 VSS.n5944 0.00286
R77450 VSS.n3588 VSS.n3587 0.00285923
R77451 VSS.n5093 VSS.n5028 0.00285923
R77452 VSS.n5583 VSS.n5461 0.00285923
R77453 VSS.n4420 VSS.n4396 0.00285923
R77454 VSS.n6033 VSS.n4396 0.00285923
R77455 VSS.n3589 VSS.n3588 0.00285923
R77456 VSS.n5581 VSS.n5461 0.00285923
R77457 VSS.n5093 VSS.n5026 0.00285923
R77458 VSS.n5469 VSS.n5453 0.00285075
R77459 VSS.n5099 VSS.n5032 0.00285075
R77460 VSS.n136 VSS.n131 0.00284
R77461 VSS.n19 VSS.n18 0.00284
R77462 VSS.n3925 VSS.n3924 0.00277528
R77463 VSS.n704 DVSS 0.00277528
R77464 VSS.n5659 VSS.n5658 0.0027
R77465 VSS.n5656 VSS.n5655 0.0027
R77466 VSS.n5168 VSS.n4445 0.0027
R77467 VSS.n3726 VSS.n851 0.00269
R77468 VSS.n5842 VSS.n4982 0.00269
R77469 VSS.n5868 VSS.n4917 0.00269
R77470 VSS.n5629 VSS.n5274 0.00269
R77471 VSS.n5852 VSS.n4956 0.00269
R77472 VSS.n6098 VSS.n4311 0.00269
R77473 VSS.n5984 VSS.n4859 0.00269
R77474 VSS.n2145 VSS.n2079 0.00257
R77475 VSS.n3726 VSS.n852 0.00257
R77476 VSS.n5842 VSS.n4990 0.00257
R77477 VSS.n5869 VSS.n5868 0.00257
R77478 VSS.n5629 VSS.n5260 0.00257
R77479 VSS.n5852 VSS.n4973 0.00257
R77480 VSS.n6098 VSS.n4319 0.00257
R77481 VSS.n5981 VSS.n4859 0.00257
R77482 VSS.n1618 VSS.n1617 0.00254225
R77483 VSS.n1650 VSS.n1325 0.00254225
R77484 VSS.n5433 VSS.n5132 0.00254
R77485 VSS.n5604 VSS.n5603 0.00254
R77486 VSS.n5432 VSS.n4366 0.00254
R77487 VSS.n1859 DVSS 0.00247183
R77488 VSS.n3864 VSS.n725 0.00239607
R77489 VSS.n3858 VSS.n731 0.00239607
R77490 VSS.n5377 VSS.n5376 0.00238
R77491 VSS.n5390 VSS.n5328 0.00238
R77492 VSS.n5383 VSS.n5382 0.00238
R77493 VSS.n1406 VSS.n1355 0.00236429
R77494 VSS.n1500 VSS.n1499 0.00236429
R77495 VSS.n2023 VSS.n1160 0.00236429
R77496 VSS.n1989 VSS.n1116 0.00236429
R77497 VSS.n2720 VSS.n1163 0.00236429
R77498 VSS.n2827 VSS.n2826 0.00236429
R77499 VSS.n3934 VSS.n660 0.00236429
R77500 VSS.n3974 VSS.n3969 0.00236429
R77501 VSS.n4602 VSS.n4268 0.00236429
R77502 VSS.n4635 VSS.n4488 0.00236429
R77503 VSS.n1796 DVSS 0.0023
R77504 VSS.n3035 DVSS 0.0023
R77505 VSS.n1019 DVSS 0.0023
R77506 VSS.n4060 DVSS 0.0023
R77507 VSS.n4698 DVSS 0.0023
R77508 VSS.n444 VSS.n7 0.0023
R77509 VSS.n441 VSS.n125 0.0023
R77510 VSS.n6246 VSS 0.0023
R77511 VSS VSS.n6247 0.0023
R77512 VSS VSS.n6469 0.0023
R77513 VSS.n6468 VSS 0.0023
R77514 VSS.n1664 VSS.n1663 0.00226056
R77515 VSS.n1746 VSS.n1285 0.00226056
R77516 VSS.n3335 DVSS 0.00218942
R77517 VSS.n1892 VSS.n1222 0.0021791
R77518 VSS.n4813 VSS.n4411 0.0021791
R77519 VSS.n5518 VSS.n5477 0.0021791
R77520 DVSS VSS.n2373 0.0021723
R77521 VSS.n2148 VSS.n2079 0.00215
R77522 VSS.n5840 VSS.n4990 0.00215
R77523 VSS.n5632 VSS.n5260 0.00215
R77524 VSS.n6095 VSS.n4319 0.00215
R77525 VSS.n1496 VSS.n1489 0.00210714
R77526 VSS.n1755 VSS.n1754 0.00210714
R77527 VSS.n1982 VSS.n1104 0.00210714
R77528 VSS.n2993 VSS.n1077 0.00210714
R77529 VSS.n2824 VSS.n2811 0.00210714
R77530 VSS.n3436 VSS.n3435 0.00210714
R77531 VSS.n3979 VSS.n618 0.00210714
R77532 VSS.n4018 VSS.n572 0.00210714
R77533 VSS.n4775 VSS.n4496 0.00210714
R77534 VSS.n4768 VSS.n4518 0.00210714
R77535 VSS.n3723 VSS.n851 0.00203
R77536 VSS.n4943 VSS.n4917 0.00203
R77537 VSS.n5855 VSS.n4956 0.00203
R77538 VSS.n5985 VSS.n5984 0.00203
R77539 VSS.n3798 VSS.n3797 0.00201685
R77540 VSS.n1326 VSS.n1307 0.00201119
R77541 DVSS VSS.n5922 0.00196
R77542 VSS.n2974 VSS.n1112 0.00184328
R77543 VSS.n2973 VSS.n1106 0.00184328
R77544 VSS.n2970 VSS.n2968 0.00184328
R77545 VSS.n1858 DVSS 0.00181455
R77546 VSS.n5924 DVSS 0.00173
R77547 DVSS VSS.n5919 0.00173
R77548 VSS.n6467 VSS 0.0017
R77549 VSS.n6054 VSS.n6053 0.0017
R77550 VSS.n5606 VSS.n4365 0.0017
R77551 VSS.n5762 VSS.n5761 0.0017
R77552 VSS.n5134 VSS.n5128 0.0017
R77553 VSS.n5607 VSS.n5430 0.0017
R77554 VSS.n4368 VSS.n4361 0.0017
R77555 VSS.n3280 VSS.n3266 0.00163764
R77556 VSS.n482 VSS.n480 0.00150746
R77557 VSS.n5455 VSS.n5256 0.00150746
R77558 VSS.n5079 VSS.n5033 0.00150746
R77559 VSS.n6009 VSS.n4442 0.00146
R77560 VSS.n5557 VSS.n5171 0.00146
R77561 VSS.n5167 VSS.n5165 0.00146
R77562 VSS.n5725 VSS.n5724 0.00146
R77563 VSS.n5556 VSS.n4443 0.00146
R77564 VSS.n6008 VSS.n6007 0.00146
R77565 VSS.n5987 VSS.n4472 0.0014
R77566 VSS.n5521 VSS.n4952 0.0014
R77567 VSS.n5990 VSS.n4471 0.0014
R77568 VSS.n5522 VSS.n5181 0.0014
R77569 VSS.n6103 VSS.n6102 0.0014
R77570 VSS.n5624 VSS.n5287 0.0014
R77571 VSS.n6100 VSS.n4309 0.0014
R77572 VSS.n5626 VSS.n5277 0.0014
R77573 VSS.n3535 VSS.n3534 0.00137
R77574 VSS.n3567 VSS.n947 0.00137
R77575 VSS.n5781 VSS.n5771 0.00137
R77576 VSS.n5745 VSS.n5027 0.00137
R77577 VSS.n5622 VSS.n5289 0.00137
R77578 VSS.n5587 VSS.n5447 0.00137
R77579 VSS.n6104 VSS.n4294 0.00137
R77580 VSS.n6037 VSS.n4381 0.00137
R77581 DVSS VSS.n3691 0.00134
R77582 VSS.n5961 DVSS 0.00134
R77583 VSS.n5433 VSS.n5131 0.0013
R77584 VSS.n5605 VSS.n5604 0.0013
R77585 VSS.n5432 VSS.n4364 0.0013
R77586 VSS.n1546 VSS.n1342 0.00127465
R77587 VSS.n1661 VSS.n1659 0.00127465
R77588 VSS.n2551 VSS.n2549 0.00125843
R77589 VSS.n3592 VSS.n3591 0.00125
R77590 VSS.n3641 VSS.n3640 0.00125
R77591 VSS.n5825 VSS.n5035 0.00125
R77592 VSS.n5804 VSS.n5064 0.00125
R77593 VSS.n5578 VSS.n5572 0.00125
R77594 VSS.n5643 VSS.n5252 0.00125
R77595 VSS.n6031 VSS.n6024 0.00125
R77596 VSS.n5996 VSS.n4460 0.00125
R77597 VSS.n5982 VSS.n4907 0.00122
R77598 VSS.n5906 VSS.n4913 0.00122
R77599 VSS.n5905 VSS.n4914 0.00122
R77600 VSS.n5870 VSS.n5869 0.00122
R77601 VSS.n4973 VSS.n4908 0.00122
R77602 VSS.n5981 VSS.n5980 0.00122
R77603 VSS.n1536 VSS.n1356 0.00120714
R77604 VSS.n1432 VSS.n1426 0.00120714
R77605 VSS.n2020 VSS.n1161 0.00120714
R77606 VSS.n1940 VSS.n1103 0.00120714
R77607 VSS.n2859 VSS.n1164 0.00120714
R77608 VSS.n2746 VSS.n2743 0.00120714
R77609 VSS.n3937 VSS.n654 0.00120714
R77610 VSS.n3976 VSS.n3975 0.00120714
R77611 VSS.n6121 VSS.n4270 0.00120714
R77612 VSS.n4538 VSS.n4489 0.00120714
R77613 VSS.n5658 VSS.n5657 0.00114
R77614 VSS.n5656 VSS.n5169 0.00114
R77615 VSS.n5168 VSS.n4441 0.00114
R77616 VSS.n3863 VSS.n727 0.00113202
R77617 VSS.n3861 VSS.n734 0.00113202
R77618 VSS.n6271 VSS.n6270 0.00107857
R77619 VSS.n261 VSS.n109 0.00107857
R77620 DVSS VSS.n5885 0.00102
R77621 VSS.n1320 VSS.n1306 0.000992958
R77622 VSS.n1742 VSS.n1284 0.000992958
R77623 VSS.n5688 VSS.n4910 0.00098
R77624 VSS.n5943 VSS.n4911 0.00098
R77625 VSS.n5944 VSS.n4906 0.00098
R77626 VSS.n1493 VSS.n1433 0.00095
R77627 VSS.n1751 VSS.n1274 0.00095
R77628 VSS.n2975 VSS.n1107 0.00095
R77629 VSS.n2986 VSS.n1084 0.00095
R77630 VSS.n2821 VSS.n2747 0.00095
R77631 VSS.n2779 VSS.n974 0.00095
R77632 VSS.n3980 VSS.n622 0.00095
R77633 VSS.n602 VSS.n571 0.00095
R77634 VSS.n4506 VSS.n4490 0.00095
R77635 VSS.n4765 VSS.n4516 0.00095
R77636 VSS.n6032 VSS.n4421 0.000835821
R77637 VSS.n5525 VSS.n5475 0.000835821
R77638 VSS.n3533 VSS.n963 0.00083
R77639 VSS.n3589 VSS.n3576 0.00083
R77640 VSS.n5784 VSS.n5082 0.00083
R77641 VSS.n5742 VSS.n5028 0.00083
R77642 VSS.n5619 VSS.n5297 0.00083
R77643 VSS.n5584 VSS.n5583 0.00083
R77644 VSS.n6107 VSS.n4280 0.00083
R77645 VSS.n6034 VSS.n6033 0.00083
R77646 VSS.n1220 VSS.n1218 0.000725
R77647 VSS.n3587 VSS.n911 0.00071
R77648 VSS.n3637 VSS.n881 0.00071
R77649 VSS.n5029 VSS.n5026 0.00071
R77650 VSS.n5797 VSS.n5054 0.00071
R77651 VSS.n5581 VSS.n5505 0.00071
R77652 VSS.n5646 VSS.n5186 0.00071
R77653 VSS.n4422 VSS.n4420 0.00071
R77654 VSS.n5997 VSS.n4449 0.00071
R77655 VSS.n1858 DVSS 0.000687793
R77656 DVSS VSS.n5887 0.00068
R77657 VSS.n6467 VSS 0.000671429
R77658 VSS.n1797 DVSS 0.000671429
R77659 VSS.n3036 DVSS 0.000671429
R77660 VSS.n1018 DVSS 0.000671429
R77661 VSS.n4061 DVSS 0.000671429
R77662 VSS.n4699 DVSS 0.000671429
R77663 VSS VSS.n120 0.000671429
R77664 VSS.n733 DVSS 0.000626404
R77665 DVSS VSS.n3689 0.00058
R77666 VSS.n5960 DVSS 0.00058
C0 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/comp018green_esd_rc_v5p0_0.ppolyf_u_CDNS_406619531453_4.MINUS DVDD 0.538423f
C1 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/comp018green_esd_rc_v5p0_0.ppolyf_u_CDNS_406619531453_1.PLUS DVDD 0.542321f
C2 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D DVSS 0.227121p
C3 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/comp018green_esd_rc_v5p0_0.VRC GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D 0.003635f
C4 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/comp018green_esd_rc_v5p0_0.ppolyf_u_CDNS_406619531453_2.PLUS DVDD 0.570214f
C5 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/comp018green_esd_rc_v5p0_0.ppolyf_u_CDNS_406619531453_5.MINUS DVDD 0.538226f
C6 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/comp018green_esd_rc_v5p0_0.ppolyf_u_CDNS_406619531453_0.PLUS DVDD 0.570627f
C7 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/comp018green_esd_rc_v5p0_0.VRC DVSS 61.6913f
C8 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/comp018green_esd_rc_v5p0_0.ppolyf_u_CDNS_406619531453_4.MINUS DVSS 0.003034f
C9 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/comp018green_esd_rc_v5p0_0.ppolyf_u_CDNS_406619531453_1.PLUS DVSS 6.15e-19
C10 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/comp018green_esd_rc_v5p0_0.ppolyf_u_CDNS_406619531453_2.PLUS DVSS 6.15e-19
C11 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/comp018green_esd_rc_v5p0_0.ppolyf_u_CDNS_406619531453_5.MINUS DVSS 0.003034f
C12 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/comp018green_esd_rc_v5p0_0.ppolyf_u_CDNS_406619531453_0.PLUS DVSS 0.002054f
C13 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D DVDD 0.251346p
C14 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/comp018green_esd_rc_v5p0_0.ppolyf_u_CDNS_406619531453_5.MINUS GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/comp018green_esd_rc_v5p0_0.VRC 1.19e-19
C15 DVSS DVDD 1.48144p
C16 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/comp018green_esd_rc_v5p0_0.ppolyf_u_CDNS_406619531453_4.MINUS GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/comp018green_esd_rc_v5p0_0.ppolyf_u_CDNS_406619531453_5.MINUS 0.034604f
C17 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/comp018green_esd_rc_v5p0_0.ppolyf_u_CDNS_406619531453_1.PLUS GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/comp018green_esd_rc_v5p0_0.ppolyf_u_CDNS_406619531453_0.PLUS 0.034604f
C18 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/comp018green_esd_rc_v5p0_0.VRC DVDD 0.112463p
C19 DVDD VSS 0.880631p
C20 DVSS VSS 0.211885p
C21 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D VSS 33.875786f
C22 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/comp018green_esd_rc_v5p0_0.VRC VSS 0.133911p
C23 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/comp018green_esd_rc_v5p0_0.ppolyf_u_CDNS_406619531453_0.PLUS VSS 0.157857f
C24 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/comp018green_esd_rc_v5p0_0.ppolyf_u_CDNS_406619531453_1.PLUS VSS 0.154878f
C25 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/comp018green_esd_rc_v5p0_0.ppolyf_u_CDNS_406619531453_5.MINUS VSS 0.155044f
C26 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/comp018green_esd_rc_v5p0_0.ppolyf_u_CDNS_406619531453_4.MINUS VSS 0.155044f
C27 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/comp018green_esd_rc_v5p0_0.ppolyf_u_CDNS_406619531453_2.PLUS VSS 0.159321f
C28 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/comp018green_esd_rc_v5p0_0.VRC.t0 VSS 0.017911f
C29 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/comp018green_esd_rc_v5p0_0.VRC.t13 VSS 0.170634f
C30 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/comp018green_esd_rc_v5p0_0.VRC.n0 VSS 0.152315f
C31 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/comp018green_esd_rc_v5p0_0.VRC.t12 VSS 0.154782f
C32 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/comp018green_esd_rc_v5p0_0.VRC.t1 VSS 0.170634f
C33 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/comp018green_esd_rc_v5p0_0.VRC.n1 VSS 0.152315f
C34 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/comp018green_esd_rc_v5p0_0.VRC.t2 VSS 0.154782f
C35 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/comp018green_esd_rc_v5p0_0.VRC.n2 VSS 0.005882f
C36 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/comp018green_esd_rc_v5p0_0.VRC.n3 VSS 0.999109f
C37 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/comp018green_esd_rc_v5p0_0.VRC.t3 VSS 0.153998f
C38 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/comp018green_esd_rc_v5p0_0.VRC.n4 VSS 1.87468f
C39 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/comp018green_esd_rc_v5p0_0.VRC.t6 VSS 7.174971f
C40 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/comp018green_esd_rc_v5p0_0.VRC.n6 VSS 0.519969f
C41 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/comp018green_esd_rc_v5p0_0.VRC.t7 VSS 7.174971f
C42 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/comp018green_esd_rc_v5p0_0.VRC.n8 VSS 0.518237f
C43 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/comp018green_esd_rc_v5p0_0.VRC.t4 VSS 7.174971f
C44 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/comp018green_esd_rc_v5p0_0.VRC.n10 VSS 0.561703f
C45 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/comp018green_esd_rc_v5p0_0.VRC.t5 VSS 7.174971f
C46 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/comp018green_esd_rc_v5p0_0.VRC.n12 VSS 1.57821f
C47 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/comp018green_esd_rc_v5p0_0.VRC.t10 VSS 7.174971f
C48 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/comp018green_esd_rc_v5p0_0.VRC.n14 VSS 0.519969f
C49 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/comp018green_esd_rc_v5p0_0.VRC.t11 VSS 7.174971f
C50 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/comp018green_esd_rc_v5p0_0.VRC.n16 VSS 0.518237f
C51 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/comp018green_esd_rc_v5p0_0.VRC.t8 VSS 7.174971f
C52 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/comp018green_esd_rc_v5p0_0.VRC.n18 VSS 0.628256f
C53 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/comp018green_esd_rc_v5p0_0.VRC.t9 VSS 7.174971f
C54 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531459_0.D.t2 VSS 0.62014f
C55 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531459_0.D.n0 VSS 2.84693f
C56 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531459_0.D.t0 VSS 0.813844f
C57 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531459_0.D.t1 VSS 0.632255f
C58 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531459_0.D.t9 VSS 0.752207f
C59 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531459_0.D.t10 VSS 0.682327f
C60 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531459_0.D.n1 VSS 0.684419f
C61 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531459_0.D.t5 VSS 0.682327f
C62 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531459_0.D.n2 VSS 0.37715f
C63 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531459_0.D.t4 VSS 0.752207f
C64 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531459_0.D.t11 VSS 0.682327f
C65 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531459_0.D.n3 VSS 0.684419f
C66 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531459_0.D.t8 VSS 0.682327f
C67 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531459_0.D.n4 VSS 0.37715f
C68 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531459_0.D.n5 VSS 0.514488f
C69 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531459_0.D.t3 VSS 0.752207f
C70 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531459_0.D.t7 VSS 0.752207f
C71 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531459_0.D.t6 VSS 0.682327f
C72 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531459_0.D.n6 VSS 1.02875f
C73 DVSS.n0 VSS 0.215195f
C74 DVSS.n1 VSS 0.333965f
C75 DVSS.n2 VSS 0.333965f
C76 DVSS.n3 VSS 0.333965f
C77 DVSS.n4 VSS 0.333965f
C78 DVSS.n5 VSS 0.333965f
C79 DVSS.n6 VSS 0.333965f
C80 DVSS.n7 VSS 0.333965f
C81 DVSS.n8 VSS 0.333965f
C82 DVSS.n9 VSS 0.333965f
C83 DVSS.n10 VSS 0.333965f
C84 DVSS.n11 VSS 0.637355f
C85 DVSS.n12 VSS 0.637355f
C86 DVSS.n13 VSS 0.402169f
C87 DVSS.n14 VSS 0.402169f
C88 DVSS.n15 VSS 0.166982f
C89 DVSS.n16 VSS 0.333965f
C90 DVSS.n17 VSS 0.333965f
C91 DVSS.n18 VSS 0.333965f
C92 DVSS.n19 VSS 0.333965f
C93 DVSS.n20 VSS 0.009721f
C94 DVSS.n21 VSS 0.009721f
C95 DVSS.n22 VSS 0.009721f
C96 DVSS.n23 VSS 0.009878f
C97 DVSS.n24 VSS 0.009721f
C98 DVSS.n25 VSS 0.019442f
C99 DVSS.n26 VSS 0.010505f
C100 DVSS.n27 VSS 0.009721f
C101 DVSS.n28 VSS 0.019442f
C102 DVSS.n29 VSS 0.023205f
C103 DVSS.n30 VSS 0.145816f
C104 DVSS.n31 VSS 0.009721f
C105 DVSS.n32 VSS 0.019442f
C106 DVSS.n33 VSS 0.019442f
C107 DVSS.n34 VSS 0.009721f
C108 DVSS.n35 VSS 0.009721f
C109 DVSS.n36 VSS 0.018031f
C110 DVSS.n37 VSS 0.009721f
C111 DVSS.n38 VSS 0.018658f
C112 DVSS.n39 VSS 0.009721f
C113 DVSS.n40 VSS 0.019285f
C114 DVSS.n41 VSS 0.019442f
C115 DVSS.n42 VSS 0.009721f
C116 DVSS.n43 VSS 0.019442f
C117 DVSS.n44 VSS 0.018345f
C118 DVSS.n45 VSS 0.009721f
C119 DVSS.n46 VSS 0.026052f
C120 DVSS.n47 VSS 0.009721f
C121 DVSS.n48 VSS 0.018345f
C122 DVSS.n49 VSS 0.009721f
C123 DVSS.n50 VSS 0.145816f
C124 DVSS.n51 VSS 0.019442f
C125 DVSS.n52 VSS 0.019442f
C126 DVSS.n53 VSS 0.010191f
C127 DVSS.n54 VSS 0.009721f
C128 DVSS.n55 VSS 0.009721f
C129 DVSS.n56 VSS 0.009721f
C130 DVSS.n57 VSS 0.009721f
C131 DVSS.n58 VSS 0.009721f
C132 DVSS.n59 VSS 0.011132f
C133 DVSS.n60 VSS 0.269288f
C134 DVSS.n61 VSS 0.009721f
C135 DVSS.n62 VSS 0.019442f
C136 DVSS.n63 VSS 0.018972f
C137 DVSS.n64 VSS 0.069774f
C138 DVSS.n65 VSS 0.196381f
C139 DVSS.n66 VSS 0.009721f
C140 DVSS.n67 VSS 0.009721f
C141 DVSS.n68 VSS 0.009878f
C142 DVSS.n69 VSS 0.019442f
C143 DVSS.n70 VSS 0.010505f
C144 DVSS.n71 VSS 0.019442f
C145 DVSS.n72 VSS 0.023205f
C146 DVSS.n73 VSS 0.019442f
C147 DVSS.n74 VSS 0.009721f
C148 DVSS.n75 VSS 0.018031f
C149 DVSS.n76 VSS 0.018658f
C150 DVSS.n77 VSS 0.07508f
C151 DVSS.n78 VSS 0.009878f
C152 DVSS.n79 VSS 0.009721f
C153 DVSS.n80 VSS 0.201084f
C154 DVSS.n81 VSS 0.009721f
C155 DVSS.n82 VSS 0.009721f
C156 DVSS.n83 VSS 0.009721f
C157 DVSS.n84 VSS 0.019442f
C158 DVSS.n85 VSS 0.010505f
C159 DVSS.n86 VSS 0.019442f
C160 DVSS.n87 VSS 0.023205f
C161 DVSS.n88 VSS 0.145816f
C162 DVSS.n89 VSS 0.019442f
C163 DVSS.n90 VSS 0.009721f
C164 DVSS.n91 VSS 0.018031f
C165 DVSS.n92 VSS 0.018658f
C166 DVSS.n93 VSS 0.009721f
C167 DVSS.n94 VSS 0.019442f
C168 DVSS.n95 VSS 0.019442f
C169 DVSS.n96 VSS 0.010191f
C170 DVSS.n97 VSS 0.009721f
C171 DVSS.n98 VSS 0.009721f
C172 DVSS.n99 VSS 0.009721f
C173 DVSS.n100 VSS 0.009721f
C174 DVSS.n101 VSS 0.011132f
C175 DVSS.n102 VSS 0.321029f
C176 DVSS.n103 VSS 0.009721f
C177 DVSS.n104 VSS 0.019442f
C178 DVSS.n105 VSS 0.018972f
C179 DVSS.n106 VSS 0.018345f
C180 DVSS.n107 VSS 0.174976f
C181 DVSS.n109 VSS 0.201084f
C182 DVSS.n110 VSS 0.094729f
C183 DVSS.n111 VSS 0.008467f
C184 DVSS.n112 VSS 0.009721f
C185 DVSS.n113 VSS 0.019442f
C186 DVSS.n114 VSS 0.009721f
C187 DVSS.n115 VSS 0.009721f
C188 DVSS.n116 VSS 0.009721f
C189 DVSS.n117 VSS 0.145816f
C190 DVSS.n118 VSS 0.018972f
C191 DVSS.n119 VSS 0.009721f
C192 DVSS.n120 VSS 0.009721f
C193 DVSS.n121 VSS 0.009721f
C194 DVSS.n122 VSS 0.009721f
C195 DVSS.n123 VSS 0.009721f
C196 DVSS.n124 VSS 0.014566f
C197 DVSS.n125 VSS 0.019442f
C198 DVSS.n126 VSS 0.019442f
C199 DVSS.n127 VSS 0.012073f
C200 DVSS.n128 VSS 0.019442f
C201 DVSS.n129 VSS 0.011446f
C202 DVSS.n130 VSS 0.019442f
C203 DVSS.n131 VSS 0.010819f
C204 DVSS.n132 VSS 0.019442f
C205 DVSS.n133 VSS 0.010191f
C206 DVSS.n134 VSS 0.321029f
C207 DVSS.n135 VSS 0.018345f
C208 DVSS.n136 VSS 0.017717f
C209 DVSS.n137 VSS 0.01709f
C210 DVSS.n138 VSS 0.341867f
C211 DVSS.n139 VSS 0.026052f
C212 DVSS.n141 VSS 0.044541f
C213 DVSS.n142 VSS 0.031157f
C214 DVSS.n143 VSS 0.031157f
C215 DVSS.n144 VSS 0.022691f
C216 DVSS.n146 VSS 3.11004f
C217 DVSS.n148 VSS 0.342732f
C218 DVSS.n149 VSS 0.022691f
C219 DVSS.n152 VSS 0.166982f
C220 DVSS.n153 VSS 0.154047f
C221 DVSS.n154 VSS 0.201084f
C222 DVSS.n156 VSS 0.052105f
C223 DVSS.n157 VSS 0.052105f
C224 DVSS.n158 VSS 0.032355f
C225 DVSS.n159 VSS 0.052105f
C226 DVSS.n160 VSS 0.030675f
C227 DVSS.n161 VSS 0.052105f
C228 DVSS.n162 VSS 0.028994f
C229 DVSS.n163 VSS 0.052105f
C230 DVSS.n164 VSS 0.027313f
C231 DVSS.n165 VSS 0.077737f
C232 DVSS.n166 VSS 0.145816f
C233 DVSS.n167 VSS 0.050844f
C234 DVSS.n169 VSS 0.052105f
C235 DVSS.n171 VSS 0.049163f
C236 DVSS.n173 VSS 0.052105f
C237 DVSS.n175 VSS 0.047482f
C238 DVSS.n177 VSS 0.052105f
C239 DVSS.n179 VSS 0.07508f
C240 DVSS.n180 VSS 0.052206f
C241 DVSS.n181 VSS 0.01709f
C242 DVSS.n182 VSS 0.009721f
C243 DVSS.n183 VSS 0.145816f
C244 DVSS.n184 VSS 0.008467f
C245 DVSS.n185 VSS 0.019442f
C246 DVSS.n186 VSS 0.019442f
C247 DVSS.n187 VSS 0.019442f
C248 DVSS.n188 VSS 0.011446f
C249 DVSS.n189 VSS 0.019442f
C250 DVSS.n190 VSS 0.010819f
C251 DVSS.n191 VSS 0.019442f
C252 DVSS.n192 VSS 0.010191f
C253 DVSS.n193 VSS 0.196381f
C254 DVSS.n195 VSS 0.018345f
C255 DVSS.n196 VSS 0.017717f
C256 DVSS.n197 VSS 0.01662f
C257 DVSS.n198 VSS 0.008467f
C258 DVSS.n199 VSS 0.009721f
C259 DVSS.n200 VSS 0.019442f
C260 DVSS.n201 VSS 0.009721f
C261 DVSS.n202 VSS 0.009721f
C262 DVSS.n203 VSS 0.009721f
C263 DVSS.n204 VSS 0.009721f
C264 DVSS.n205 VSS 0.009721f
C265 DVSS.n206 VSS 0.009721f
C266 DVSS.n207 VSS 0.167516f
C267 DVSS.n208 VSS 0.009721f
C268 DVSS.n209 VSS 0.009721f
C269 DVSS.n211 VSS 0.01662f
C270 DVSS.n212 VSS 0.008467f
C271 DVSS.n213 VSS 0.048035f
C272 DVSS.n214 VSS 0.048035f
C273 DVSS.n215 VSS 1.8361f
C274 DVSS.t83 VSS 4.03839f
C275 DVSS.n216 VSS -0.795461f
C276 DVSS.t37 VSS 4.03839f
C277 DVSS.n217 VSS 0.048035f
C278 DVSS.n218 VSS 1.8361f
C279 DVSS.n219 VSS 0.048035f
C280 DVSS.n221 VSS 0.009721f
C281 DVSS.n222 VSS 0.008467f
C282 DVSS.n223 VSS 0.167516f
C283 DVSS.n224 VSS 0.145816f
C284 DVSS.n225 VSS 0.008467f
C285 DVSS.n226 VSS 0.019442f
C286 DVSS.n227 VSS 0.019442f
C287 DVSS.n228 VSS 0.019442f
C288 DVSS.n229 VSS 0.009721f
C289 DVSS.n230 VSS 0.012073f
C290 DVSS.n231 VSS 0.019442f
C291 DVSS.n232 VSS 0.009721f
C292 DVSS.n233 VSS 0.011446f
C293 DVSS.n234 VSS 0.019442f
C294 DVSS.n235 VSS 0.009721f
C295 DVSS.n236 VSS 0.010819f
C296 DVSS.n237 VSS 0.019442f
C297 DVSS.n238 VSS 0.009721f
C298 DVSS.n239 VSS 0.010191f
C299 DVSS.n240 VSS 0.029006f
C300 DVSS.n241 VSS 0.269288f
C301 DVSS.n243 VSS 0.018972f
C302 DVSS.n244 VSS 0.009721f
C303 DVSS.n245 VSS 0.018345f
C304 DVSS.t160 VSS 0.203828f
C305 DVSS.t130 VSS 0.203828f
C306 DVSS.n246 VSS 0.407656f
C307 DVSS.n247 VSS 0.017717f
C308 DVSS.n248 VSS 0.009721f
C309 DVSS.n249 VSS 0.145816f
C310 DVSS.n250 VSS 0.019442f
C311 DVSS.n251 VSS 0.019442f
C312 DVSS.n252 VSS 0.012073f
C313 DVSS.n253 VSS 0.019442f
C314 DVSS.n254 VSS 0.019442f
C315 DVSS.n255 VSS 0.010819f
C316 DVSS.n256 VSS 0.019442f
C317 DVSS.n257 VSS 0.010191f
C318 DVSS.n258 VSS 0.109362f
C319 DVSS.n260 VSS 0.009721f
C320 DVSS.n261 VSS 0.026052f
C321 DVSS.n262 VSS 0.009721f
C322 DVSS.n263 VSS 0.052214f
C323 DVSS.n264 VSS 0.174976f
C324 DVSS.n265 VSS 0.07508f
C325 DVSS.t186 VSS 0.203828f
C326 DVSS.t110 VSS 0.203828f
C327 DVSS.n266 VSS 0.407656f
C328 DVSS.n267 VSS 0.073484f
C329 DVSS.n268 VSS 0.176594f
C330 DVSS.n269 VSS 0.052206f
C331 DVSS.n270 VSS 0.018345f
C332 DVSS.n271 VSS 0.01709f
C333 DVSS.n272 VSS 0.008467f
C334 DVSS.n273 VSS 0.273992f
C335 DVSS.n274 VSS 0.009721f
C336 DVSS.n275 VSS 0.019442f
C337 DVSS.n276 VSS 0.009721f
C338 DVSS.n277 VSS 0.009721f
C339 DVSS.n278 VSS 0.009721f
C340 DVSS.n279 VSS 0.017717f
C341 DVSS.n280 VSS 0.029006f
C342 DVSS.n281 VSS 0.027282f
C343 DVSS.n283 VSS 0.158751f
C344 DVSS.n284 VSS 0.154047f
C345 DVSS.n285 VSS 0.201084f
C346 DVSS.n286 VSS 0.052105f
C347 DVSS.n287 VSS 0.028994f
C348 DVSS.n288 VSS 0.052105f
C349 DVSS.n289 VSS 0.027313f
C350 DVSS.n290 VSS 0.052105f
C351 DVSS.n291 VSS 0.026473f
C352 DVSS.n292 VSS 0.052105f
C353 DVSS.n293 VSS 0.028153f
C354 DVSS.n294 VSS 0.052105f
C355 DVSS.n296 VSS 0.029834f
C356 DVSS.n297 VSS 0.052105f
C357 DVSS.n298 VSS 0.062189f
C358 DVSS.n299 VSS 0.145816f
C359 DVSS.n301 VSS 0.052105f
C360 DVSS.n303 VSS 0.052105f
C361 DVSS.n305 VSS 0.048323f
C362 DVSS.n307 VSS 0.052105f
C363 DVSS.n309 VSS 0.050004f
C364 DVSS.n311 VSS 0.052105f
C365 DVSS.n313 VSS 0.051685f
C366 DVSS.n314 VSS 0.050844f
C367 DVSS.n317 VSS 0.052105f
C368 DVSS.n318 VSS 0.049163f
C369 DVSS.n321 VSS 0.145816f
C370 DVSS.n324 VSS 0.333965f
C371 DVSS.n325 VSS 0.333965f
C372 DVSS.n326 VSS 0.333965f
C373 DVSS.n327 VSS 0.333965f
C374 DVSS.n328 VSS 0.333965f
C375 DVSS.n329 VSS 0.333965f
C376 DVSS.n330 VSS 0.333965f
C377 DVSS.n331 VSS 0.333965f
C378 DVSS.n332 VSS 0.333965f
C379 DVSS.n333 VSS 0.333965f
C380 DVSS.n334 VSS 0.333965f
C381 DVSS.n335 VSS 0.333965f
C382 DVSS.n336 VSS 0.333965f
C383 DVSS.n337 VSS 0.333965f
C384 DVSS.n338 VSS 0.333965f
C385 DVSS.n339 VSS 0.637355f
C386 DVSS.n340 VSS 0.333965f
C387 DVSS.n341 VSS 0.204612f
C388 DVSS.n342 VSS 0.402169f
C389 DVSS.n343 VSS 0.402169f
C390 DVSS.n344 VSS 0.296335f
C391 DVSS.n345 VSS 0.333965f
C392 DVSS.n346 VSS 0.333965f
C393 DVSS.n347 VSS 0.333965f
C394 DVSS.n348 VSS 0.333965f
C395 DVSS.n349 VSS 0.333965f
C396 DVSS.n350 VSS 0.325733f
C397 DVSS.n351 VSS 0.333965f
C398 DVSS.n352 VSS 0.333965f
C399 DVSS.n353 VSS 0.145816f
C400 DVSS.n354 VSS 0.019442f
C401 DVSS.n355 VSS 0.010819f
C402 DVSS.n356 VSS 0.019442f
C403 DVSS.n357 VSS 0.010191f
C404 DVSS.n358 VSS 0.009721f
C405 DVSS.n359 VSS 0.009721f
C406 DVSS.n360 VSS 0.009721f
C407 DVSS.n361 VSS 0.009721f
C408 DVSS.n362 VSS 0.009721f
C409 DVSS.n363 VSS 0.011132f
C410 DVSS.n364 VSS 0.009721f
C411 DVSS.n365 VSS 0.019442f
C412 DVSS.n366 VSS 0.018972f
C413 DVSS.n367 VSS 0.010191f
C414 DVSS.n368 VSS 0.052206f
C415 DVSS.n369 VSS 0.026052f
C416 DVSS.n370 VSS 0.009721f
C417 DVSS.n371 VSS 0.052214f
C418 DVSS.n372 VSS 0.174976f
C419 DVSS.n373 VSS 0.07508f
C420 DVSS.t116 VSS 0.203828f
C421 DVSS.t58 VSS 0.203828f
C422 DVSS.n374 VSS 0.407656f
C423 DVSS.n375 VSS 0.073484f
C424 DVSS.n376 VSS 0.176594f
C425 DVSS.n377 VSS 0.009721f
C426 DVSS.n378 VSS 0.018972f
C427 DVSS.n379 VSS 0.018345f
C428 DVSS.n380 VSS 0.009721f
C429 DVSS.n381 VSS 0.009721f
C430 DVSS.n382 VSS 0.009878f
C431 DVSS.n383 VSS 0.019442f
C432 DVSS.n384 VSS 0.010505f
C433 DVSS.n385 VSS 0.019442f
C434 DVSS.n387 VSS 0.171366f
C435 DVSS.n388 VSS 0.170933f
C436 DVSS.n389 VSS 0.166982f
C437 DVSS.n390 VSS 0.166982f
C438 DVSS.n391 VSS 0.009878f
C439 DVSS.n392 VSS 0.052206f
C440 DVSS.n393 VSS 0.026052f
C441 DVSS.n394 VSS 0.009721f
C442 DVSS.n395 VSS 0.009878f
C443 DVSS.n396 VSS 0.009721f
C444 DVSS.n397 VSS 0.196381f
C445 DVSS.n398 VSS 0.011132f
C446 DVSS.n399 VSS 0.012386f
C447 DVSS.n400 VSS 0.009721f
C448 DVSS.n401 VSS 0.017404f
C449 DVSS.n402 VSS 0.019442f
C450 DVSS.n403 VSS 0.018658f
C451 DVSS.n404 VSS 0.019442f
C452 DVSS.n405 VSS 0.145816f
C453 DVSS.n406 VSS 0.019442f
C454 DVSS.n407 VSS 0.018031f
C455 DVSS.n408 VSS 0.019442f
C456 DVSS.n409 VSS 0.016777f
C457 DVSS.n410 VSS 0.011759f
C458 DVSS.n411 VSS 0.010505f
C459 DVSS.n412 VSS 0.019442f
C460 DVSS.n413 VSS 0.015052f
C461 DVSS.n414 VSS 0.009721f
C462 DVSS.n415 VSS 0.009721f
C463 DVSS.n416 VSS 0.009721f
C464 DVSS.n417 VSS 0.009721f
C465 DVSS.n418 VSS 0.009721f
C466 DVSS.n419 VSS 0.269288f
C467 DVSS.n420 VSS 0.009721f
C468 DVSS.n421 VSS 0.009721f
C469 DVSS.n422 VSS 0.009721f
C470 DVSS.n423 VSS 0.009721f
C471 DVSS.n424 VSS 0.119007f
C472 DVSS.n425 VSS 0.07508f
C473 DVSS.n426 VSS 0.076514f
C474 DVSS.n427 VSS 0.009721f
C475 DVSS.n428 VSS 0.145816f
C476 DVSS.n429 VSS 0.015052f
C477 DVSS.n430 VSS 0.009721f
C478 DVSS.n431 VSS 0.009721f
C479 DVSS.n432 VSS 0.009721f
C480 DVSS.n433 VSS 0.009721f
C481 DVSS.n434 VSS 0.009721f
C482 DVSS.n435 VSS 0.321029f
C483 DVSS.n436 VSS 0.009721f
C484 DVSS.n437 VSS 0.009721f
C485 DVSS.n438 VSS 0.009721f
C486 DVSS.n439 VSS 0.009721f
C487 DVSS.n440 VSS 0.009721f
C488 DVSS.n441 VSS 0.009721f
C489 DVSS.n442 VSS 0.201084f
C490 DVSS.n443 VSS 0.019285f
C491 DVSS.n444 VSS 0.011132f
C492 DVSS.n445 VSS 0.012386f
C493 DVSS.n446 VSS 0.017404f
C494 DVSS.n447 VSS 0.019442f
C495 DVSS.n448 VSS 0.018658f
C496 DVSS.n449 VSS 0.019442f
C497 DVSS.n450 VSS 0.019442f
C498 DVSS.n451 VSS 0.018031f
C499 DVSS.n452 VSS 0.019442f
C500 DVSS.n453 VSS 0.016777f
C501 DVSS.n454 VSS 0.011759f
C502 DVSS.t126 VSS 0.203828f
C503 DVSS.t56 VSS 0.203828f
C504 DVSS.n455 VSS 0.407656f
C505 DVSS.n456 VSS 0.028153f
C506 DVSS.n457 VSS 0.050004f
C507 DVSS.n458 VSS 0.052206f
C508 DVSS.n459 VSS 0.011132f
C509 DVSS.n460 VSS 0.052206f
C510 DVSS.n461 VSS 0.029834f
C511 DVSS.n462 VSS 0.154047f
C512 DVSS.n465 VSS 0.158751f
C513 DVSS.n466 VSS 0.145816f
C514 DVSS.n467 VSS 0.026473f
C515 DVSS.n468 VSS 0.033196f
C516 DVSS.n469 VSS 0.052105f
C517 DVSS.n470 VSS 0.052105f
C518 DVSS.n471 VSS 0.046642f
C519 DVSS.n472 VSS 0.052105f
C520 DVSS.n473 VSS 0.052105f
C521 DVSS.n474 VSS 0.052105f
C522 DVSS.n475 VSS 0.196381f
C523 DVSS.n477 VSS 0.052105f
C524 DVSS.n479 VSS 0.052105f
C525 DVSS.n481 VSS 0.052105f
C526 DVSS.n483 VSS 0.052105f
C527 DVSS.n484 VSS 0.044961f
C528 DVSS.n486 VSS 0.069333f
C529 DVSS.n487 VSS 0.031515f
C530 DVSS.n488 VSS 0.051685f
C531 DVSS.n491 VSS 0.007789f
C532 DVSS.n492 VSS 0.021951f
C533 DVSS.n494 VSS 0.013798f
C534 DVSS.n495 VSS 0.170933f
C535 DVSS.n496 VSS 0.170933f
C536 DVSS.n497 VSS 0.013798f
C537 DVSS.n498 VSS 0.021951f
C538 DVSS.n500 VSS 0.171366f
C539 DVSS.n501 VSS 0.171366f
C540 DVSS.n502 VSS 0.015579f
C541 DVSS.n503 VSS 0.007789f
C542 DVSS.t89 VSS 2.28624f
C543 DVSS.t51 VSS 2.28624f
C544 DVSS.t143 VSS 2.28624f
C545 DVSS.t187 VSS 2.28624f
C546 DVSS.t155 VSS 2.28624f
C547 DVSS.t39 VSS 2.28624f
C548 DVSS.t175 VSS 2.28624f
C549 DVSS.t67 VSS 2.28624f
C550 DVSS.t145 VSS 2.28624f
C551 DVSS.t79 VSS 2.28624f
C552 DVSS.t165 VSS 2.28624f
C553 DVSS.t135 VSS 2.28624f
C554 DVSS.t179 VSS 2.28624f
C555 DVSS.t105 VSS 2.28624f
C556 DVSS.t43 VSS 2.28624f
C557 DVSS.t125 VSS 2.28624f
C558 DVSS.t55 VSS 2.28624f
C559 DVSS.t137 VSS 2.28624f
C560 DVSS.t71 VSS 4.03839f
C561 DVSS.t147 VSS 4.53554f
C562 DVSS.t171 VSS 2.28624f
C563 DVSS.t129 VSS 2.28624f
C564 DVSS.t159 VSS 2.28624f
C565 DVSS.t109 VSS 2.28624f
C566 DVSS.t185 VSS 2.28624f
C567 DVSS.t61 VSS 2.28624f
C568 DVSS.t169 VSS 2.28624f
C569 DVSS.t45 VSS 2.28624f
C570 DVSS.t153 VSS 2.28624f
C571 DVSS.t75 VSS 2.28624f
C572 DVSS.t139 VSS 2.28624f
C573 DVSS.t57 VSS 2.28624f
C574 DVSS.t115 VSS 2.28624f
C575 DVSS.t33 VSS 2.28624f
C576 DVSS.t113 VSS 2.28624f
C577 DVSS.t181 VSS 2.28624f
C578 DVSS.t95 VSS 2.28624f
C579 DVSS.t157 VSS 2.28624f
C580 DVSS.t81 VSS 4.03839f
C581 DVSS.n504 VSS 4.97951f
C582 DVSS.n505 VSS -0.795461f
C583 DVSS.n506 VSS 0.058828f
C584 DVSS.n507 VSS 0.171366f
C585 DVSS.n508 VSS 0.036978f
C586 DVSS.n509 VSS 0.040339f
C587 DVSS.n511 VSS 0.201084f
C588 DVSS.n512 VSS 0.052105f
C589 DVSS.n516 VSS 0.333965f
C590 DVSS.n517 VSS 0.333965f
C591 DVSS.n518 VSS 0.333965f
C592 DVSS.n519 VSS 0.333965f
C593 DVSS.n520 VSS 0.333965f
C594 DVSS.n521 VSS 0.333965f
C595 DVSS.n522 VSS 0.333965f
C596 DVSS.n523 VSS 0.333965f
C597 DVSS.n524 VSS 0.333965f
C598 DVSS.n525 VSS 0.333965f
C599 DVSS.n526 VSS 0.333965f
C600 DVSS.n527 VSS 0.333965f
C601 DVSS.n528 VSS 0.333965f
C602 DVSS.n529 VSS 0.333965f
C603 DVSS.n530 VSS 0.333965f
C604 DVSS.n531 VSS 0.333965f
C605 DVSS.n532 VSS 0.333965f
C606 DVSS.n533 VSS 0.204612f
C607 DVSS.n534 VSS 0.333965f
C608 DVSS.n535 VSS 0.204612f
C609 DVSS.n536 VSS 0.333965f
C610 DVSS.n537 VSS 0.333965f
C611 DVSS.n538 VSS 0.333965f
C612 DVSS.n539 VSS 0.333965f
C613 DVSS.n540 VSS 0.333965f
C614 DVSS.n541 VSS 0.333965f
C615 DVSS.n542 VSS 0.333965f
C616 DVSS.n543 VSS 0.333965f
C617 DVSS.n544 VSS 0.333965f
C618 DVSS.n545 VSS 0.333965f
C619 DVSS.n546 VSS 0.333965f
C620 DVSS.n547 VSS 0.333965f
C621 DVSS.n548 VSS 0.145816f
C622 DVSS.n549 VSS 0.333965f
C623 DVSS.n550 VSS 0.333965f
C624 DVSS.n551 VSS 0.333965f
C625 DVSS.n552 VSS 0.333965f
C626 DVSS.n553 VSS 0.333965f
C627 DVSS.n554 VSS 0.333965f
C628 DVSS.n555 VSS 0.333965f
C629 DVSS.n556 VSS 0.333965f
C630 DVSS.n557 VSS 0.286927f
C631 DVSS.n558 VSS 0.286927f
C632 DVSS.n559 VSS 0.637355f
C633 DVSS.n560 VSS 0.333965f
C634 DVSS.n561 VSS 0.333965f
C635 DVSS.n562 VSS 0.402169f
C636 DVSS.n563 VSS 0.333965f
C637 DVSS.n564 VSS 0.402169f
C638 DVSS.n565 VSS 0.21402f
C639 DVSS.n566 VSS 0.333965f
C640 DVSS.n567 VSS 0.402169f
C641 DVSS.n568 VSS 0.333965f
C642 DVSS.n569 VSS 0.333965f
C643 DVSS.n570 VSS 0.333965f
C644 DVSS.n571 VSS 0.333965f
C645 DVSS.n572 VSS 0.333965f
C646 DVSS.n573 VSS 0.333965f
C647 DVSS.n574 VSS 0.333965f
C648 DVSS.n575 VSS 0.333965f
C649 DVSS.n576 VSS 0.333965f
C650 DVSS.n577 VSS 0.333965f
C651 DVSS.n578 VSS 0.333965f
C652 DVSS.n579 VSS 0.333965f
C653 DVSS.n580 VSS 0.333965f
C654 DVSS.n581 VSS 0.333965f
C655 DVSS.n582 VSS 0.333965f
C656 DVSS.n583 VSS 0.333965f
C657 DVSS.n584 VSS 0.333965f
C658 DVSS.n585 VSS 0.333965f
C659 DVSS.n586 VSS 0.27752f
C660 DVSS.n587 VSS 5.70674f
C661 DVSS.n588 VSS 6.09395f
C662 DVSS.n589 VSS 3.04095f
C663 DVSS.n590 VSS 0.333965f
C664 DVSS.n591 VSS 6.09395f
C665 DVSS.n592 VSS 7.251f
C666 DVSS.n593 VSS 4.8454f
C667 DVSS.n594 VSS 4.61021f
C668 DVSS.n595 VSS 0.196381f
C669 DVSS.n596 VSS 0.333965f
C670 DVSS.n597 VSS 0.333965f
C671 DVSS.n598 VSS 0.333965f
C672 DVSS.n599 VSS 0.333965f
C673 DVSS.n600 VSS 0.333965f
C674 DVSS.n601 VSS 0.333965f
C675 DVSS.n602 VSS 0.333965f
C676 DVSS.n603 VSS 0.333965f
C677 DVSS.n604 VSS 0.333965f
C678 DVSS.n605 VSS 0.333965f
C679 DVSS.n606 VSS 0.333965f
C680 DVSS.n607 VSS 0.333965f
C681 DVSS.n608 VSS 0.333965f
C682 DVSS.n609 VSS 0.333965f
C683 DVSS.n610 VSS 0.333965f
C684 DVSS.n611 VSS 0.333965f
C685 DVSS.n612 VSS 0.333965f
C686 DVSS.n613 VSS 0.333965f
C687 DVSS.n614 VSS 0.333965f
C688 DVSS.n615 VSS 0.333965f
C689 DVSS.n616 VSS 0.333965f
C690 DVSS.n617 VSS 0.333965f
C691 DVSS.n618 VSS 0.333965f
C692 DVSS.n619 VSS 0.333965f
C693 DVSS.n620 VSS 0.333965f
C694 DVSS.n621 VSS 0.333965f
C695 DVSS.n622 VSS 0.333965f
C696 DVSS.n623 VSS 0.333965f
C697 DVSS.n624 VSS 0.333965f
C698 DVSS.n625 VSS 0.333965f
C699 DVSS.n626 VSS 0.333965f
C700 DVSS.n627 VSS 0.333965f
C701 DVSS.n628 VSS 0.333965f
C702 DVSS.n629 VSS 0.333965f
C703 DVSS.n630 VSS 0.333965f
C704 DVSS.n631 VSS 0.333965f
C705 DVSS.n632 VSS 0.333965f
C706 DVSS.n633 VSS 0.333965f
C707 DVSS.n634 VSS 0.333965f
C708 DVSS.n635 VSS 0.333965f
C709 DVSS.n636 VSS 0.333965f
C710 DVSS.n637 VSS 0.333965f
C711 DVSS.n638 VSS 0.333965f
C712 DVSS.n639 VSS 0.333965f
C713 DVSS.n640 VSS 0.333965f
C714 DVSS.n641 VSS 0.333965f
C715 DVSS.n642 VSS 0.333965f
C716 DVSS.n643 VSS 0.333965f
C717 DVSS.n644 VSS 0.333965f
C718 DVSS.n645 VSS 0.333965f
C719 DVSS.n646 VSS 0.333965f
C720 DVSS.n647 VSS 0.333965f
C721 DVSS.n648 VSS 0.333965f
C722 DVSS.n649 VSS 0.333965f
C723 DVSS.n650 VSS 0.333965f
C724 DVSS.n651 VSS 0.333965f
C725 DVSS.n652 VSS 0.333965f
C726 DVSS.n653 VSS 0.333965f
C727 DVSS.n654 VSS 0.27752f
C728 DVSS.n655 VSS 0.27752f
C729 DVSS.n656 VSS 1.29862f
C730 DVSS.n657 VSS 1.53381f
C731 DVSS.n658 VSS 1.63161f
C732 DVSS.n659 VSS 0.333965f
C733 DVSS.n660 VSS 0.333965f
C734 DVSS.n661 VSS 0.333965f
C735 DVSS.n662 VSS 0.333965f
C736 DVSS.n663 VSS 0.333965f
C737 DVSS.n664 VSS 0.333965f
C738 DVSS.n665 VSS 0.333965f
C739 DVSS.n666 VSS 0.333965f
C740 DVSS.n667 VSS 0.333965f
C741 DVSS.n668 VSS 0.333965f
C742 DVSS.n669 VSS 0.333965f
C743 DVSS.n670 VSS 0.333965f
C744 DVSS.n671 VSS 0.333965f
C745 DVSS.n672 VSS 0.333965f
C746 DVSS.n673 VSS 0.333965f
C747 DVSS.n674 VSS 0.333965f
C748 DVSS.n675 VSS 0.333965f
C749 DVSS.n676 VSS 0.333965f
C750 DVSS.n677 VSS 0.333965f
C751 DVSS.n678 VSS 0.333965f
C752 DVSS.n679 VSS 0.333965f
C753 DVSS.n680 VSS 0.333965f
C754 DVSS.n681 VSS 0.333965f
C755 DVSS.n682 VSS 0.333965f
C756 DVSS.n683 VSS 0.333965f
C757 DVSS.n684 VSS 0.333965f
C758 DVSS.n685 VSS 0.333965f
C759 DVSS.n686 VSS 0.333965f
C760 DVSS.n687 VSS 0.333965f
C761 DVSS.n688 VSS 0.333965f
C762 DVSS.n689 VSS 0.333965f
C763 DVSS.n690 VSS 0.333965f
C764 DVSS.n691 VSS 0.333965f
C765 DVSS.n692 VSS 0.333965f
C766 DVSS.n693 VSS 0.333965f
C767 DVSS.n694 VSS 0.333965f
C768 DVSS.n695 VSS 0.333965f
C769 DVSS.n696 VSS 0.333965f
C770 DVSS.n697 VSS 0.333965f
C771 DVSS.n698 VSS 0.333965f
C772 DVSS.n699 VSS 0.333965f
C773 DVSS.n700 VSS 0.333965f
C774 DVSS.n701 VSS 0.333965f
C775 DVSS.n702 VSS 0.333965f
C776 DVSS.n703 VSS 0.333965f
C777 DVSS.n704 VSS 0.333965f
C778 DVSS.n705 VSS 0.333965f
C779 DVSS.n706 VSS 0.333965f
C780 DVSS.n707 VSS 0.333965f
C781 DVSS.n708 VSS 0.333965f
C782 DVSS.n709 VSS 0.333965f
C783 DVSS.n710 VSS 0.333965f
C784 DVSS.n711 VSS 0.333965f
C785 DVSS.n712 VSS 0.333965f
C786 DVSS.n713 VSS 0.286927f
C787 DVSS.n714 VSS 0.286927f
C788 DVSS.n715 VSS 0.286927f
C789 DVSS.n716 VSS 0.402169f
C790 DVSS.n717 VSS 0.21402f
C791 DVSS.n718 VSS 0.21402f
C792 DVSS.n719 VSS 0.21402f
C793 DVSS.n720 VSS 0.333965f
C794 DVSS.n721 VSS 0.333965f
C795 DVSS.n722 VSS 0.333965f
C796 DVSS.n723 VSS 0.333965f
C797 DVSS.n724 VSS 0.333965f
C798 DVSS.n725 VSS 0.333965f
C799 DVSS.n726 VSS 0.333965f
C800 DVSS.n727 VSS 0.333965f
C801 DVSS.n728 VSS 0.333965f
C802 DVSS.n729 VSS 0.333965f
C803 DVSS.n730 VSS 0.333965f
C804 DVSS.n731 VSS 0.333965f
C805 DVSS.n732 VSS 0.333965f
C806 DVSS.n733 VSS 0.333965f
C807 DVSS.n734 VSS 0.333965f
C808 DVSS.n735 VSS 0.333965f
C809 DVSS.n736 VSS 0.333965f
C810 DVSS.n737 VSS 0.333965f
C811 DVSS.n738 VSS 0.333965f
C812 DVSS.n739 VSS 0.333965f
C813 DVSS.n740 VSS 0.333965f
C814 DVSS.n741 VSS 0.333965f
C815 DVSS.n742 VSS 0.333965f
C816 DVSS.n743 VSS 0.333965f
C817 DVSS.n744 VSS 0.333965f
C818 DVSS.n745 VSS 0.333965f
C819 DVSS.n746 VSS 0.333965f
C820 DVSS.n747 VSS 0.333965f
C821 DVSS.n748 VSS 0.333965f
C822 DVSS.n749 VSS 0.333965f
C823 DVSS.n750 VSS 0.333965f
C824 DVSS.n751 VSS 0.333965f
C825 DVSS.n752 VSS 0.333965f
C826 DVSS.n753 VSS 0.27752f
C827 DVSS.n754 VSS 0.27752f
C828 DVSS.n755 VSS 5.78597f
C829 DVSS.n756 VSS 5.94193f
C830 DVSS.n757 VSS 0.27752f
C831 DVSS.n758 VSS 0.333965f
C832 DVSS.n759 VSS 0.333965f
C833 DVSS.n760 VSS 0.333965f
C834 DVSS.n761 VSS 0.333965f
C835 DVSS.n762 VSS 0.333965f
C836 DVSS.n763 VSS 0.333965f
C837 DVSS.n764 VSS 0.333965f
C838 DVSS.n765 VSS 0.333965f
C839 DVSS.n766 VSS 0.333965f
C840 DVSS.n767 VSS 0.333965f
C841 DVSS.n768 VSS 0.333965f
C842 DVSS.n769 VSS 0.333965f
C843 DVSS.n770 VSS 0.333965f
C844 DVSS.n771 VSS 0.333965f
C845 DVSS.n772 VSS 0.333965f
C846 DVSS.n773 VSS 0.333965f
C847 DVSS.n774 VSS 0.333965f
C848 DVSS.n775 VSS 0.333965f
C849 DVSS.n776 VSS 0.333965f
C850 DVSS.n777 VSS 0.333965f
C851 DVSS.n778 VSS 0.333965f
C852 DVSS.n779 VSS 0.333965f
C853 DVSS.n780 VSS 0.333965f
C854 DVSS.n781 VSS 0.333965f
C855 DVSS.n782 VSS 0.333965f
C856 DVSS.n783 VSS 0.333965f
C857 DVSS.n784 VSS 0.333965f
C858 DVSS.n785 VSS 0.333965f
C859 DVSS.n786 VSS 0.333965f
C860 DVSS.n787 VSS 0.333965f
C861 DVSS.n788 VSS 0.333965f
C862 DVSS.n789 VSS 0.333965f
C863 DVSS.n790 VSS 0.333965f
C864 DVSS.n791 VSS 0.333965f
C865 DVSS.n792 VSS 0.333965f
C866 DVSS.n793 VSS 0.333965f
C867 DVSS.n794 VSS 0.333965f
C868 DVSS.n795 VSS 0.333965f
C869 DVSS.n796 VSS 0.333965f
C870 DVSS.n797 VSS 0.333965f
C871 DVSS.n798 VSS 0.333965f
C872 DVSS.n799 VSS 0.333965f
C873 DVSS.n800 VSS 0.333965f
C874 DVSS.n801 VSS 0.21402f
C875 DVSS.n802 VSS 0.21402f
C876 DVSS.n803 VSS 0.637355f
C877 DVSS.n804 VSS 0.286927f
C878 DVSS.n805 VSS 0.333965f
C879 DVSS.n806 VSS 0.333965f
C880 DVSS.n807 VSS 0.333965f
C881 DVSS.n808 VSS 0.333965f
C882 DVSS.n809 VSS 0.333965f
C883 DVSS.n810 VSS 0.333965f
C884 DVSS.n811 VSS 0.333965f
C885 DVSS.n812 VSS 0.333965f
C886 DVSS.n813 VSS 0.333965f
C887 DVSS.n814 VSS 0.333965f
C888 DVSS.n815 VSS 0.333965f
C889 DVSS.n816 VSS 0.333965f
C890 DVSS.n817 VSS 0.333965f
C891 DVSS.n818 VSS 0.333965f
C892 DVSS.n819 VSS 0.333965f
C893 DVSS.n820 VSS 0.333965f
C894 DVSS.n821 VSS 0.333965f
C895 DVSS.n822 VSS 0.333965f
C896 DVSS.n823 VSS 0.333965f
C897 DVSS.n824 VSS 0.333965f
C898 DVSS.n825 VSS 0.333965f
C899 DVSS.n826 VSS 0.333965f
C900 DVSS.n827 VSS 0.333965f
C901 DVSS.n828 VSS 0.333965f
C902 DVSS.n829 VSS 0.333965f
C903 DVSS.n830 VSS 0.333965f
C904 DVSS.n831 VSS 0.333965f
C905 DVSS.n832 VSS 0.333965f
C906 DVSS.n833 VSS 0.333965f
C907 DVSS.n834 VSS 0.333965f
C908 DVSS.n835 VSS 0.286927f
C909 DVSS.n836 VSS 0.286927f
C910 DVSS.n837 VSS 0.637355f
C911 DVSS.n838 VSS 0.402169f
C912 DVSS.n839 VSS 0.21402f
C913 DVSS.n840 VSS 0.21402f
C914 DVSS.n841 VSS 0.21402f
C915 DVSS.n842 VSS 0.402169f
C916 DVSS.n843 VSS 0.286927f
C917 DVSS.n844 VSS 0.333965f
C918 DVSS.n845 VSS 0.333965f
C919 DVSS.n846 VSS 0.333965f
C920 DVSS.n847 VSS 0.333965f
C921 DVSS.n848 VSS 0.333965f
C922 DVSS.n849 VSS 0.333965f
C923 DVSS.n850 VSS 0.333965f
C924 DVSS.n851 VSS 0.333965f
C925 DVSS.n852 VSS 0.333965f
C926 DVSS.n853 VSS 0.333965f
C927 DVSS.n854 VSS 0.333965f
C928 DVSS.n855 VSS 0.333965f
C929 DVSS.n856 VSS 0.333965f
C930 DVSS.n857 VSS 0.333965f
C931 DVSS.n858 VSS 0.333965f
C932 DVSS.n859 VSS 0.333965f
C933 DVSS.n860 VSS 0.333965f
C934 DVSS.n861 VSS 0.333965f
C935 DVSS.n862 VSS 0.333965f
C936 DVSS.n863 VSS 0.333965f
C937 DVSS.n864 VSS 0.333965f
C938 DVSS.n865 VSS 0.333965f
C939 DVSS.n866 VSS 0.333965f
C940 DVSS.n867 VSS 0.333965f
C941 DVSS.n868 VSS 0.333965f
C942 DVSS.n869 VSS 0.196381f
C943 DVSS.n870 VSS 0.333965f
C944 DVSS.n871 VSS 0.333965f
C945 DVSS.n872 VSS 0.333965f
C946 DVSS.n873 VSS 0.333965f
C947 DVSS.n874 VSS 0.333965f
C948 DVSS.n875 VSS 0.333965f
C949 DVSS.n876 VSS 0.333965f
C950 DVSS.n877 VSS 0.333965f
C951 DVSS.n878 VSS 0.333965f
C952 DVSS.n879 VSS 0.333965f
C953 DVSS.n880 VSS 0.333965f
C954 DVSS.n881 VSS 0.333965f
C955 DVSS.n882 VSS 0.333965f
C956 DVSS.n883 VSS 0.333965f
C957 DVSS.n884 VSS 0.333965f
C958 DVSS.n885 VSS 0.333965f
C959 DVSS.n886 VSS 0.333965f
C960 DVSS.n887 VSS 0.333965f
C961 DVSS.n888 VSS 0.333965f
C962 DVSS.n889 VSS 0.204612f
C963 DVSS.n890 VSS 0.204612f
C964 DVSS.n891 VSS 0.402169f
C965 DVSS.n892 VSS 0.333965f
C966 DVSS.n893 VSS 0.333965f
C967 DVSS.n894 VSS 0.333965f
C968 DVSS.n895 VSS 0.325733f
C969 DVSS.n896 VSS 0.333965f
C970 DVSS.n897 VSS 0.333965f
C971 DVSS.n898 VSS 0.333965f
C972 DVSS.n899 VSS 0.333965f
C973 DVSS.n900 VSS 0.333965f
C974 DVSS.n901 VSS 0.333965f
C975 DVSS.n902 VSS 0.333965f
C976 DVSS.n903 VSS 0.333965f
C977 DVSS.n904 VSS 0.333965f
C978 DVSS.n905 VSS 0.333965f
C979 DVSS.n906 VSS 0.333965f
C980 DVSS.n907 VSS 0.333965f
C981 DVSS.n908 VSS 0.333965f
C982 DVSS.n909 VSS 0.333965f
C983 DVSS.n910 VSS 0.333965f
C984 DVSS.n911 VSS 0.333965f
C985 DVSS.n912 VSS 0.333965f
C986 DVSS.n913 VSS 0.333965f
C987 DVSS.n914 VSS 0.333965f
C988 DVSS.n915 VSS 0.333965f
C989 DVSS.n916 VSS 0.333965f
C990 DVSS.n917 VSS 0.333965f
C991 DVSS.n918 VSS 0.333965f
C992 DVSS.n919 VSS 0.195205f
C993 DVSS.n920 VSS 0.305742f
C994 DVSS.n921 VSS 0.333965f
C995 DVSS.n922 VSS 0.402169f
C996 DVSS.n923 VSS 0.333965f
C997 DVSS.n924 VSS 0.333965f
C998 DVSS.n925 VSS 0.333965f
C999 DVSS.n926 VSS 0.333965f
C1000 DVSS.n927 VSS 0.333965f
C1001 DVSS.n928 VSS 0.333965f
C1002 DVSS.n929 VSS 0.333965f
C1003 DVSS.n930 VSS 0.333965f
C1004 DVSS.n931 VSS 0.333965f
C1005 DVSS.n932 VSS 0.333965f
C1006 DVSS.n933 VSS 0.333965f
C1007 DVSS.n934 VSS 0.333965f
C1008 DVSS.n935 VSS 0.197556f
C1009 DVSS.n936 VSS 0.333965f
C1010 DVSS.n937 VSS 0.326909f
C1011 DVSS.n938 VSS 1.31793f
C1012 DVSS.n939 VSS 0.553111f
C1013 DVSS.n940 VSS 0.326909f
C1014 DVSS.n941 VSS 0.333965f
C1015 DVSS.n942 VSS 0.333965f
C1016 DVSS.n943 VSS 0.333965f
C1017 DVSS.n944 VSS 0.333965f
C1018 DVSS.n945 VSS 0.333965f
C1019 DVSS.n946 VSS 0.333965f
C1020 DVSS.n947 VSS 0.333965f
C1021 DVSS.n948 VSS 0.333965f
C1022 DVSS.n949 VSS 0.333965f
C1023 DVSS.n950 VSS 0.333965f
C1024 DVSS.n951 VSS 0.333965f
C1025 DVSS.n952 VSS 0.333965f
C1026 DVSS.n953 VSS 0.333965f
C1027 DVSS.n954 VSS 0.333965f
C1028 DVSS.n955 VSS 0.305742f
C1029 DVSS.n956 VSS 0.305742f
C1030 DVSS.n957 VSS 0.402169f
C1031 DVSS.n958 VSS 0.195205f
C1032 DVSS.n959 VSS 0.333965f
C1033 DVSS.n960 VSS 0.333965f
C1034 DVSS.n961 VSS 0.333965f
C1035 DVSS.n962 VSS 0.333965f
C1036 DVSS.n963 VSS 0.333965f
C1037 DVSS.n964 VSS 0.333965f
C1038 DVSS.n965 VSS 0.333965f
C1039 DVSS.n966 VSS 0.333965f
C1040 DVSS.n967 VSS 0.333965f
C1041 DVSS.n968 VSS 0.333965f
C1042 DVSS.n969 VSS 0.333965f
C1043 DVSS.n970 VSS 0.333965f
C1044 DVSS.n971 VSS 0.333965f
C1045 DVSS.n972 VSS 0.333965f
C1046 DVSS.n973 VSS 0.333965f
C1047 DVSS.n974 VSS 0.333965f
C1048 DVSS.n975 VSS 0.333965f
C1049 DVSS.n976 VSS 0.333965f
C1050 DVSS.n977 VSS 0.333965f
C1051 DVSS.n978 VSS 0.333965f
C1052 DVSS.n979 VSS 0.333965f
C1053 DVSS.n980 VSS 0.333965f
C1054 DVSS.n981 VSS 0.333965f
C1055 DVSS.n982 VSS 0.333965f
C1056 DVSS.n983 VSS 0.333965f
C1057 DVSS.n984 VSS 0.333965f
C1058 DVSS.n985 VSS 0.333965f
C1059 DVSS.n986 VSS 0.333965f
C1060 DVSS.n987 VSS 0.333965f
C1061 DVSS.n988 VSS 0.333965f
C1062 DVSS.n989 VSS 0.333965f
C1063 DVSS.n990 VSS 0.333965f
C1064 DVSS.n991 VSS 0.333965f
C1065 DVSS.n992 VSS 0.296335f
C1066 DVSS.n993 VSS 0.296335f
C1067 DVSS.n994 VSS 0.296335f
C1068 DVSS.n995 VSS 0.402169f
C1069 DVSS.n996 VSS 0.637355f
C1070 DVSS.n997 VSS 0.402169f
C1071 DVSS.n998 VSS 0.296335f
C1072 DVSS.n999 VSS 0.333965f
C1073 DVSS.n1000 VSS 0.333965f
C1074 DVSS.n1001 VSS 0.333965f
C1075 DVSS.n1002 VSS 0.333965f
C1076 DVSS.n1003 VSS 0.333965f
C1077 DVSS.n1004 VSS 0.325733f
C1078 DVSS.n1005 VSS 0.145816f
C1079 DVSS.n1006 VSS 0.196381f
C1080 DVSS.n1007 VSS 0.333965f
C1081 DVSS.n1008 VSS 0.333965f
C1082 DVSS.n1009 VSS 0.333965f
C1083 DVSS.n1010 VSS 0.333965f
C1084 DVSS.n1011 VSS 0.333965f
C1085 DVSS.n1012 VSS 0.333965f
C1086 DVSS.n1013 VSS 0.333965f
C1087 DVSS.n1014 VSS 0.333965f
C1088 DVSS.n1015 VSS 0.333965f
C1089 DVSS.n1016 VSS 0.333965f
C1090 DVSS.n1017 VSS 0.333965f
C1091 DVSS.n1018 VSS 0.333965f
C1092 DVSS.n1019 VSS 0.333965f
C1093 DVSS.n1020 VSS 0.333965f
C1094 DVSS.n1021 VSS 0.333965f
C1095 DVSS.n1022 VSS 0.333965f
C1096 DVSS.n1023 VSS 0.333965f
C1097 DVSS.n1024 VSS 0.333965f
C1098 DVSS.n1025 VSS 0.333965f
C1099 DVSS.n1026 VSS 0.333965f
C1100 DVSS.n1027 VSS 0.333965f
C1101 DVSS.n1028 VSS 0.333965f
C1102 DVSS.n1029 VSS 0.273992f
C1103 DVSS.n1030 VSS 0.333965f
C1104 DVSS.n1031 VSS 0.402169f
C1105 DVSS.n1032 VSS 0.333965f
C1106 DVSS.n1033 VSS 0.305742f
C1107 DVSS.n1034 VSS 0.333965f
C1108 DVSS.n1035 VSS 0.333965f
C1109 DVSS.n1036 VSS 0.333965f
C1110 DVSS.n1037 VSS 0.333965f
C1111 DVSS.n1038 VSS 0.333965f
C1112 DVSS.n1039 VSS 0.333965f
C1113 DVSS.n1040 VSS 0.333965f
C1114 DVSS.n1041 VSS 0.333965f
C1115 DVSS.n1042 VSS 0.333965f
C1116 DVSS.n1043 VSS 0.333965f
C1117 DVSS.n1044 VSS 0.333965f
C1118 DVSS.n1045 VSS 0.333965f
C1119 DVSS.n1046 VSS 0.333965f
C1120 DVSS.n1047 VSS 0.301038f
C1121 DVSS.n1048 VSS 1.35288f
C1122 DVSS.n1049 VSS 0.578982f
C1123 DVSS.n1050 VSS 0.171686f
C1124 DVSS.n1051 VSS 0.333965f
C1125 DVSS.n1052 VSS 0.301038f
C1126 DVSS.n1053 VSS 0.333965f
C1127 DVSS.n1054 VSS 0.333965f
C1128 DVSS.n1055 VSS 0.333965f
C1129 DVSS.n1056 VSS 0.333965f
C1130 DVSS.n1057 VSS 0.333965f
C1131 DVSS.n1058 VSS 0.333965f
C1132 DVSS.n1059 VSS 0.333965f
C1133 DVSS.n1060 VSS 0.333965f
C1134 DVSS.n1061 VSS 0.333965f
C1135 DVSS.n1062 VSS 0.333965f
C1136 DVSS.n1063 VSS 0.333965f
C1137 DVSS.n1064 VSS 0.333965f
C1138 DVSS.n1065 VSS 0.333965f
C1139 DVSS.n1066 VSS 0.305742f
C1140 DVSS.n1067 VSS 0.305742f
C1141 DVSS.n1068 VSS 0.402169f
C1142 DVSS.n1069 VSS 0.195205f
C1143 DVSS.n1070 VSS 0.195205f
C1144 DVSS.n1071 VSS 0.166982f
C1145 DVSS.n1072 VSS 0.021951f
C1146 DVSS.n1074 VSS 0.013798f
C1147 DVSS.n1075 VSS 0.015052f
C1148 DVSS.n1076 VSS 0.009721f
C1149 DVSS.n1077 VSS 0.009721f
C1150 DVSS.n1078 VSS 0.011132f
C1151 DVSS.n1079 VSS 0.009721f
C1152 DVSS.n1080 VSS 0.010505f
C1153 DVSS.n1081 VSS 0.009721f
C1154 DVSS.n1082 VSS 0.009878f
C1155 DVSS.n1083 VSS 0.009721f
C1156 DVSS.n1084 VSS 0.109362f
C1157 DVSS.n1085 VSS 0.018658f
C1158 DVSS.n1086 VSS 0.019442f
C1159 DVSS.n1087 VSS 0.009721f
C1160 DVSS.n1088 VSS 0.018031f
C1161 DVSS.n1089 VSS 0.019442f
C1162 DVSS.n1090 VSS 0.009721f
C1163 DVSS.n1091 VSS 0.019442f
C1164 DVSS.n1092 VSS 0.009721f
C1165 DVSS.n1093 VSS 0.019442f
C1166 DVSS.n1094 VSS 0.009721f
C1167 DVSS.n1095 VSS 0.118999f
C1168 DVSS.n1096 VSS 0.012386f
C1169 DVSS.n1097 VSS 0.016777f
C1170 DVSS.n1098 VSS 0.052206f
C1171 DVSS.n1099 VSS 0.026052f
C1172 DVSS.n1100 VSS 0.009721f
C1173 DVSS.n1101 VSS 0.052214f
C1174 DVSS.n1102 VSS 0.174976f
C1175 DVSS.n1103 VSS 0.07508f
C1176 DVSS.t80 VSS 0.203828f
C1177 DVSS.t166 VSS 0.203828f
C1178 DVSS.n1104 VSS 0.407656f
C1179 DVSS.n1105 VSS 0.073484f
C1180 DVSS.n1106 VSS 0.176594f
C1181 DVSS.n1107 VSS 0.011759f
C1182 DVSS.n1108 VSS 0.017404f
C1183 DVSS.n1109 VSS 0.052206f
C1184 DVSS.n1110 VSS 0.026052f
C1185 DVSS.n1111 VSS 0.009721f
C1186 DVSS.n1112 VSS 0.052214f
C1187 DVSS.n1113 VSS 0.174976f
C1188 DVSS.n1114 VSS 0.07508f
C1189 DVSS.t136 VSS 0.203828f
C1190 DVSS.t180 VSS 0.203828f
C1191 DVSS.n1115 VSS 0.407656f
C1192 DVSS.n1116 VSS 0.073484f
C1193 DVSS.n1117 VSS 0.176594f
C1194 DVSS.n1118 VSS 0.009721f
C1195 DVSS.n1119 VSS 0.019442f
C1196 DVSS.n1120 VSS 0.009721f
C1197 DVSS.n1121 VSS 0.017404f
C1198 DVSS.n1122 VSS 0.009721f
C1199 DVSS.n1123 VSS 0.011759f
C1200 DVSS.n1124 VSS 0.009721f
C1201 DVSS.n1125 VSS 0.019442f
C1202 DVSS.n1126 VSS 0.009721f
C1203 DVSS.n1127 VSS 0.016777f
C1204 DVSS.n1128 VSS 0.009721f
C1205 DVSS.n1129 VSS 0.012386f
C1206 DVSS.n1130 VSS 0.009721f
C1207 DVSS.n1131 VSS 0.009721f
C1208 DVSS.n1132 VSS 0.025871f
C1209 DVSS.n1133 VSS 0.054406f
C1210 DVSS.n1134 VSS 0.205057f
C1211 DVSS.n1135 VSS 0.174976f
C1212 DVSS.n1136 VSS 0.07508f
C1213 DVSS.n1137 VSS 0.060521f
C1214 DVSS.n1138 VSS 0.118999f
C1215 DVSS.n1139 VSS 0.076514f
C1216 DVSS.n1140 VSS 0.031985f
C1217 DVSS.n1141 VSS 0.07508f
C1218 DVSS.n1143 VSS 0.068047f
C1219 DVSS.n1144 VSS 0.018972f
C1220 DVSS.n1145 VSS 0.009721f
C1221 DVSS.n1146 VSS 0.015993f
C1222 DVSS.n1147 VSS 0.149814f
C1223 DVSS.n1148 VSS 0.019442f
C1224 DVSS.n1149 VSS 0.009721f
C1225 DVSS.n1150 VSS 0.008467f
C1226 DVSS.n1151 VSS 0.073064f
C1227 DVSS.n1152 VSS 0.093839f
C1228 DVSS.n1153 VSS 0.019442f
C1229 DVSS.n1154 VSS 0.019442f
C1230 DVSS.n1155 VSS 0.011446f
C1231 DVSS.n1156 VSS 0.07508f
C1232 DVSS.n1157 VSS 0.01317f
C1233 DVSS.n1159 VSS 0.068047f
C1234 DVSS.n1160 VSS 0.018972f
C1235 DVSS.n1161 VSS 0.009721f
C1236 DVSS.n1162 VSS 0.125668f
C1237 DVSS.n1163 VSS 0.019442f
C1238 DVSS.n1164 VSS 0.009721f
C1239 DVSS.n1165 VSS 0.008467f
C1240 DVSS.n1166 VSS 0.115557f
C1241 DVSS.n1167 VSS 3.71965f
C1242 DVSS.n1168 VSS 0.019442f
C1243 DVSS.n1169 VSS 0.019442f
C1244 DVSS.n1170 VSS 0.009721f
C1245 DVSS.n1172 VSS 0.026052f
C1246 DVSS.n1173 VSS 0.007789f
C1247 DVSS.n1174 VSS 0.050844f
C1248 DVSS.n1175 VSS 0.007789f
C1249 DVSS.n1176 VSS 0.022691f
C1250 DVSS.n1177 VSS 0.007789f
C1251 DVSS.n1179 VSS 0.018972f
C1252 DVSS.n1180 VSS 0.008467f
C1253 DVSS.n1182 VSS 0.018972f
C1254 DVSS.n1183 VSS 0.077925f
C1255 DVSS.n1184 VSS 0.009721f
C1256 DVSS.n1185 VSS 0.068047f
C1257 DVSS.n1186 VSS 0.011446f
C1258 DVSS.n1187 VSS 0.009721f
C1259 DVSS.n1188 VSS 0.019442f
C1260 DVSS.n1189 VSS 0.019442f
C1261 DVSS.n1190 VSS 0.019442f
C1262 DVSS.n1191 VSS 0.015993f
C1263 DVSS.n1192 VSS 0.11579f
C1264 DVSS.n1194 VSS 0.031985f
C1265 DVSS.n1195 VSS 0.009721f
C1266 DVSS.n1196 VSS 0.01317f
C1267 DVSS.n1197 VSS 0.118999f
C1268 DVSS.n1198 VSS 0.073064f
C1269 DVSS.n1199 VSS 0.205057f
C1270 DVSS.n1200 VSS 0.07508f
C1271 DVSS.n1201 VSS 0.076514f
C1272 DVSS.n1202 VSS 0.118999f
C1273 DVSS.n1203 VSS 0.076514f
C1274 DVSS.n1204 VSS 0.119007f
C1275 DVSS.n1205 VSS 0.07508f
C1276 DVSS.n1206 VSS 0.076514f
C1277 DVSS.t132 VSS 0.203828f
C1278 DVSS.t54 VSS 0.203828f
C1279 DVSS.n1207 VSS 0.407656f
C1280 DVSS.n1208 VSS 0.205057f
C1281 DVSS.n1209 VSS 0.205057f
C1282 DVSS.t104 VSS 0.203828f
C1283 DVSS.t74 VSS 0.203828f
C1284 DVSS.n1210 VSS 0.407656f
C1285 DVSS.n1211 VSS 0.073484f
C1286 DVSS.n1212 VSS 0.176594f
C1287 DVSS.n1213 VSS 0.118999f
C1288 DVSS.n1214 VSS 0.118999f
C1289 DVSS.n1215 VSS 0.076514f
C1290 DVSS.n1216 VSS 0.118999f
C1291 DVSS.n1217 VSS 0.119007f
C1292 DVSS.n1218 VSS 0.07508f
C1293 DVSS.n1219 VSS 0.076514f
C1294 DVSS.t152 VSS 0.203828f
C1295 DVSS.t86 VSS 0.203828f
C1296 DVSS.n1220 VSS 0.407656f
C1297 DVSS.n1221 VSS 0.205057f
C1298 DVSS.n1222 VSS 0.205057f
C1299 DVSS.t102 VSS 0.203828f
C1300 DVSS.t178 VSS 0.203828f
C1301 DVSS.n1223 VSS 0.407656f
C1302 DVSS.n1224 VSS 0.073484f
C1303 DVSS.n1225 VSS 0.176594f
C1304 DVSS.n1226 VSS 0.118999f
C1305 DVSS.n1227 VSS 0.118999f
C1306 DVSS.n1228 VSS 0.092036f
C1307 DVSS.n1229 VSS 0.118999f
C1308 DVSS.n1230 VSS 0.062246f
C1309 DVSS.n1231 VSS 0.07508f
C1310 DVSS.n1233 VSS 0.170933f
C1311 DVSS.n1234 VSS 0.171366f
C1312 DVSS.n1235 VSS 0.076514f
C1313 DVSS.n1236 VSS 0.07508f
C1314 DVSS.n1237 VSS 0.119007f
C1315 DVSS.t100 VSS 0.203828f
C1316 DVSS.t174 VSS 0.203828f
C1317 DVSS.n1238 VSS 0.407656f
C1318 DVSS.n1239 VSS 0.205057f
C1319 DVSS.n1240 VSS 0.246657f
C1320 DVSS.n1241 VSS 0.118999f
C1321 DVSS.n1242 VSS 0.076514f
C1322 DVSS.t122 VSS 0.203828f
C1323 DVSS.t42 VSS 0.203828f
C1324 DVSS.n1243 VSS 0.407656f
C1325 DVSS.n1244 VSS 0.073484f
C1326 DVSS.n1245 VSS 0.176594f
C1327 DVSS.n1246 VSS 0.171366f
C1328 DVSS.n1249 VSS 0.007789f
C1329 DVSS.n1250 VSS 0.015579f
C1330 DVSS.n1251 VSS 0.007789f
C1331 DVSS.n1252 VSS 0.031157f
C1332 DVSS.n1254 VSS 0.177744f
C1333 DVSS.n1258 VSS 0.342732f
C1334 DVSS.n1259 VSS 0.031157f
C1335 DVSS.n1260 VSS 0.342732f
C1336 DVSS.n1261 VSS 0.104209f
C1337 DVSS.t21 VSS 0.020383f
C1338 DVSS.t198 VSS 0.020383f
C1339 DVSS.n1262 VSS 0.044773f
C1340 DVSS.n1263 VSS 0.01935f
C1341 DVSS.t196 VSS 0.020383f
C1342 DVSS.t192 VSS 0.020383f
C1343 DVSS.n1264 VSS 0.044773f
C1344 DVSS.n1265 VSS 0.01573f
C1345 DVSS.t190 VSS 0.020383f
C1346 DVSS.t194 VSS 0.020383f
C1347 DVSS.n1266 VSS 0.044773f
C1348 DVSS.n1267 VSS 0.01573f
C1349 DVSS.t11 VSS 0.054111f
C1350 DVSS.n1268 VSS 0.034585f
C1351 DVSS.t7 VSS 0.054111f
C1352 DVSS.n1269 VSS 0.03321f
C1353 DVSS.n1270 VSS 0.033619f
C1354 DVSS.n1271 VSS 0.107774f
C1355 DVSS.n1272 VSS 0.27834f
C1356 DVSS.n1273 VSS 0.694544f
C1357 DVSS.n1274 VSS 3.42532f
C1358 DVSS.n1275 VSS 0.173236p
C1359 DVSS.n1276 VSS 5.97127f
C1360 DVSS.n1277 VSS 2.41336f
C1361 DVSS.n1278 VSS 3.93009f
C1362 DVSS.n1279 VSS 0.14291f
C1363 DVSS.n1280 VSS 5.55271f
C1364 DVSS.n1281 VSS -1.89621f
C1365 DVSS.n1282 VSS 1.9427f
C1366 DVSS.n1283 VSS 0.293307f
C1367 DVSS.n1284 VSS 0.135955f
C1368 DVSS.n1285 VSS 0.125047f
C1369 DVSS.t17 VSS 0.020383f
C1370 DVSS.t23 VSS 0.020383f
C1371 DVSS.n1286 VSS 0.044773f
C1372 DVSS.n1287 VSS 0.01573f
C1373 DVSS.n1288 VSS 0.025675f
C1374 DVSS.t13 VSS 0.020383f
C1375 DVSS.t19 VSS 0.020383f
C1376 DVSS.n1289 VSS 0.044773f
C1377 DVSS.n1290 VSS 0.01573f
C1378 DVSS.n1291 VSS 1.29237f
C1379 DVSS.t14 VSS 0.786659f
C1380 DVSS.t12 VSS 0.352799f
C1381 DVSS.t10 VSS 0.343588f
C1382 DVSS.t193 VSS 0.449519f
C1383 DVSS.t189 VSS 0.449519f
C1384 DVSS.t191 VSS 0.449519f
C1385 DVSS.t195 VSS 0.449519f
C1386 DVSS.t197 VSS 0.449519f
C1387 DVSS.t20 VSS 0.449519f
C1388 DVSS.t22 VSS 0.338061f
C1389 DVSS.n1292 VSS 0.22476f
C1390 DVSS.t16 VSS 0.336218f
C1391 DVSS.t18 VSS 0.32148f
C1392 DVSS.n1293 VSS 0.22476f
C1393 DVSS.n1294 VSS 0.079587f
C1394 DVSS.n1295 VSS 0.042947f
C1395 DVSS.t15 VSS 0.054111f
C1396 DVSS.n1296 VSS 0.034585f
C1397 DVSS.n1297 VSS 0.056131f
C1398 DVSS.n1298 VSS 0.038884f
C1399 DVSS.n1299 VSS 0.341867f
C1400 DVSS.n1300 VSS 0.342732f
C1401 DVSS.n1301 VSS 0.174976f
C1402 DVSS.n1302 VSS 0.174976f
C1403 DVSS.n1303 VSS 0.174976f
C1404 DVSS.n1304 VSS 0.174976f
C1405 DVSS.n1305 VSS 0.174976f
C1406 DVSS.n1306 VSS 0.174976f
C1407 DVSS.n1307 VSS 0.008467f
C1408 DVSS.n1308 VSS 1.00544f
C1409 DVSS.n1309 VSS 0.09674f
C1410 DVSS.n1310 VSS 0.008467f
C1411 DVSS.n1311 VSS 0.341867f
C1412 DVSS.n1312 VSS 0.066322f
C1413 DVSS.n1313 VSS 0.138606f
C1414 DVSS.n1314 VSS 0.119007f
C1415 DVSS.n1315 VSS 0.119007f
C1416 DVSS.n1316 VSS 0.119007f
C1417 DVSS.n1317 VSS 0.119007f
C1418 DVSS.n1318 VSS 0.119007f
C1419 DVSS.n1319 VSS 0.119007f
C1420 DVSS.n1320 VSS 0.174976f
C1421 DVSS.t92 VSS 0.203828f
C1422 DVSS.t164 VSS 0.203828f
C1423 DVSS.n1321 VSS 0.407656f
C1424 DVSS.n1322 VSS 0.118999f
C1425 DVSS.n1323 VSS 0.076514f
C1426 DVSS.n1324 VSS 0.205057f
C1427 DVSS.n1325 VSS 0.07508f
C1428 DVSS.n1326 VSS 0.076514f
C1429 DVSS.n1327 VSS 0.118999f
C1430 DVSS.n1328 VSS 0.205057f
C1431 DVSS.n1329 VSS 0.07508f
C1432 DVSS.n1330 VSS 0.096113f
C1433 DVSS.n1331 VSS 0.008467f
C1434 DVSS.n1332 VSS 0.341867f
C1435 DVSS.n1333 VSS 0.038884f
C1436 DVSS.n1334 VSS 0.009721f
C1437 DVSS.n1335 VSS 0.068047f
C1438 DVSS.n1336 VSS 0.009721f
C1439 DVSS.n1337 VSS 0.019442f
C1440 DVSS.n1338 VSS 0.019442f
C1441 DVSS.n1339 VSS 0.019442f
C1442 DVSS.n1340 VSS 0.019442f
C1443 DVSS.n1341 VSS 0.15585f
C1444 DVSS.n1342 VSS 0.15585f
C1445 DVSS.n1343 VSS 0.15585f
C1446 DVSS.n1344 VSS 0.15585f
C1447 DVSS.n1345 VSS 0.15585f
C1448 DVSS.n1346 VSS 0.15585f
C1449 DVSS.n1347 VSS 0.15585f
C1450 DVSS.n1348 VSS 0.15585f
C1451 DVSS.n1349 VSS 0.15585f
C1452 DVSS.n1350 VSS 0.15585f
C1453 DVSS.n1351 VSS 0.15585f
C1454 DVSS.n1352 VSS 0.15585f
C1455 DVSS.n1353 VSS 0.15585f
C1456 DVSS.n1354 VSS 0.15585f
C1457 DVSS.n1355 VSS 0.15585f
C1458 DVSS.n1356 VSS 0.15585f
C1459 DVSS.n1357 VSS 0.15585f
C1460 DVSS.n1358 VSS 0.15585f
C1461 DVSS.n1359 VSS 0.009721f
C1462 DVSS.n1360 VSS 0.019442f
C1463 DVSS.n1361 VSS 0.019442f
C1464 DVSS.n1362 VSS 0.019442f
C1465 DVSS.n1363 VSS 0.019442f
C1466 DVSS.n1364 VSS 0.009721f
C1467 DVSS.n1365 VSS 0.019442f
C1468 DVSS.n1366 VSS 0.019442f
C1469 DVSS.n1367 VSS 0.019442f
C1470 DVSS.n1368 VSS 0.019442f
C1471 DVSS.n1369 VSS 0.241458f
C1472 DVSS.n1370 VSS 0.012766f
C1473 DVSS.n1371 VSS 0.015218f
C1474 DVSS.n1372 VSS 0.018232f
C1475 DVSS.n1373 VSS 0.016872f
C1476 DVSS.n1374 VSS 1.13742f
C1477 DVSS.n1375 VSS 1.33697f
C1478 DVSS.n1376 VSS 0.02143f
C1479 DVSS.n1377 VSS 0.018232f
C1480 DVSS.n1378 VSS 0.016872f
C1481 DVSS.n1379 VSS 0.031816f
C1482 DVSS.n1380 VSS 0.050993f
C1483 DVSS.n1381 VSS 0.047318f
C1484 DVSS.n1382 VSS 0.018232f
C1485 DVSS.n1383 VSS 0.018232f
C1486 DVSS.n1384 VSS 0.018232f
C1487 DVSS.n1386 VSS 0.009436f
C1488 DVSS.n1411 VSS 0.018232f
C1489 DVSS.n1412 VSS 0.111484f
C1490 DVSS.n1413 VSS 0.018232f
C1491 DVSS.n1415 VSS 0.018232f
C1492 DVSS.n1416 VSS 0.052371f
C1493 DVSS.n1417 VSS 0.052371f
C1494 DVSS.n1418 VSS 0.018232f
C1495 DVSS.n1420 VSS 0.018232f
C1496 DVSS.n1421 VSS 0.052371f
C1497 DVSS.n1422 VSS 0.052371f
C1498 DVSS.n1423 VSS 0.018232f
C1499 DVSS.n1425 VSS 0.018232f
C1500 DVSS.n1426 VSS 0.052371f
C1501 DVSS.n1427 VSS 0.052371f
C1502 DVSS.n1428 VSS 0.018232f
C1503 DVSS.n1430 VSS 0.018232f
C1504 DVSS.n1431 VSS 0.052371f
C1505 DVSS.n1432 VSS 0.052371f
C1506 DVSS.n1433 VSS 0.018232f
C1507 DVSS.n1435 VSS 0.018232f
C1508 DVSS.n1436 VSS 0.052371f
C1509 DVSS.n1437 VSS 0.052371f
C1510 DVSS.n1438 VSS 0.018232f
C1511 DVSS.n1440 VSS 0.018232f
C1512 DVSS.n1441 VSS 0.052371f
C1513 DVSS.n1442 VSS 0.052371f
C1514 DVSS.n1443 VSS 0.018232f
C1515 DVSS.n1445 VSS 0.018232f
C1516 DVSS.n1446 VSS 0.052371f
C1517 DVSS.n1447 VSS 0.052371f
C1518 DVSS.n1448 VSS 0.018232f
C1519 DVSS.n1450 VSS 0.018232f
C1520 DVSS.n1451 VSS 0.052371f
C1521 DVSS.n1452 VSS 0.052371f
C1522 DVSS.n1453 VSS 0.018232f
C1523 DVSS.n1455 VSS 0.018232f
C1524 DVSS.n1456 VSS 0.052371f
C1525 DVSS.n1457 VSS 0.052371f
C1526 DVSS.n1458 VSS 0.018232f
C1527 DVSS.n1460 VSS 0.018232f
C1528 DVSS.n1461 VSS 0.052371f
C1529 DVSS.n1462 VSS 0.046169f
C1530 DVSS.n1463 VSS 0.018232f
C1531 DVSS.n1465 VSS 0.018232f
C1532 DVSS.n1466 VSS 0.032387f
C1533 DVSS.n1467 VSS 0.033995f
C1534 DVSS.n1468 VSS 0.018232f
C1535 DVSS.n1470 VSS 0.018232f
C1536 DVSS.n1471 VSS 0.044562f
C1537 DVSS.n1472 VSS 0.052371f
C1538 DVSS.n1473 VSS 0.018232f
C1539 DVSS.n1475 VSS 0.018232f
C1540 DVSS.n1476 VSS 0.052371f
C1541 DVSS.n1477 VSS 0.052371f
C1542 DVSS.n1478 VSS 0.018232f
C1543 DVSS.n1480 VSS 0.018232f
C1544 DVSS.n1481 VSS 0.052371f
C1545 DVSS.n1482 VSS 0.052371f
C1546 DVSS.n1483 VSS 0.018232f
C1547 DVSS.n1485 VSS 0.018232f
C1548 DVSS.n1486 VSS 0.052371f
C1549 DVSS.n1487 VSS 0.052371f
C1550 DVSS.n1488 VSS 0.018232f
C1551 DVSS.n1490 VSS 0.018232f
C1552 DVSS.n1491 VSS 0.052371f
C1553 DVSS.n1492 VSS 0.052371f
C1554 DVSS.n1493 VSS 0.018232f
C1555 DVSS.n1495 VSS 0.018232f
C1556 DVSS.n1496 VSS 0.052371f
C1557 DVSS.n1497 VSS 0.052371f
C1558 DVSS.n1498 VSS 0.018232f
C1559 DVSS.n1500 VSS 0.018232f
C1560 DVSS.n1501 VSS 0.052371f
C1561 DVSS.n1502 VSS 0.052371f
C1562 DVSS.n1503 VSS 0.018232f
C1563 DVSS.n1505 VSS 0.018232f
C1564 DVSS.n1506 VSS 0.052371f
C1565 DVSS.n1507 VSS 0.052371f
C1566 DVSS.n1508 VSS 0.018232f
C1567 DVSS.n1510 VSS 0.018232f
C1568 DVSS.n1511 VSS 0.052371f
C1569 DVSS.n1512 VSS 0.052371f
C1570 DVSS.n1513 VSS 0.018232f
C1571 DVSS.n1515 VSS 0.018232f
C1572 DVSS.n1516 VSS 0.191377f
C1573 DVSS.n1517 VSS 0.003262f
C1574 DVSS.n1518 VSS 0.046185f
C1575 DVSS.n1520 VSS 22.0472f
C1576 DVSS.n1521 VSS 0.014633f
C1577 DVSS.n1522 VSS 0.042078f
C1578 DVSS.n1523 VSS 0.012766f
C1579 DVSS.n1524 VSS 0.172627f
C1580 DVSS.n1525 VSS 0.166982f
C1581 DVSS.n1526 VSS 0.019442f
C1582 DVSS.n1527 VSS 0.273992f
C1583 DVSS.n1528 VSS 0.019442f
C1584 DVSS.n1529 VSS 0.019442f
C1585 DVSS.n1530 VSS 0.019442f
C1586 DVSS.n1531 VSS 0.019442f
C1587 DVSS.n1532 VSS 0.019442f
C1588 DVSS.n1533 VSS 0.019442f
C1589 DVSS.n1534 VSS 0.019442f
C1590 DVSS.n1535 VSS 0.019442f
C1591 DVSS.n1536 VSS 0.019442f
C1592 DVSS.n1537 VSS 0.019442f
C1593 DVSS.n1538 VSS 0.019442f
C1594 DVSS.n1539 VSS 0.019442f
C1595 DVSS.n1540 VSS 0.019442f
C1596 DVSS.n1541 VSS 0.019442f
C1597 DVSS.n1542 VSS 0.019442f
C1598 DVSS.n1543 VSS 0.019442f
C1599 DVSS.n1544 VSS 0.019442f
C1600 DVSS.n1545 VSS 0.019442f
C1601 DVSS.n1546 VSS 0.019442f
C1602 DVSS.n1547 VSS 0.019442f
C1603 DVSS.n1548 VSS 0.009721f
C1604 DVSS.n1549 VSS 0.333965f
C1605 DVSS.n1550 VSS 0.333965f
C1606 DVSS.n1551 VSS 0.333965f
C1607 DVSS.n1552 VSS 0.333965f
C1608 DVSS.n1553 VSS 0.333965f
C1609 DVSS.n1554 VSS 0.333965f
C1610 DVSS.n1555 VSS 0.333965f
C1611 DVSS.n1556 VSS 0.333965f
C1612 DVSS.n1557 VSS 0.333965f
C1613 DVSS.n1558 VSS 0.333965f
C1614 DVSS.n1559 VSS 0.333965f
C1615 DVSS.n1560 VSS 0.333965f
C1616 DVSS.n1561 VSS 0.333965f
C1617 DVSS.n1562 VSS 0.333965f
C1618 DVSS.n1563 VSS 0.333965f
C1619 DVSS.n1564 VSS 0.166982f
C1620 DVSS.n1565 VSS 0.333965f
C1621 DVSS.n1566 VSS 0.333965f
C1622 DVSS.n1567 VSS 0.333965f
C1623 DVSS.n1568 VSS 0.333965f
C1624 DVSS.n1569 VSS 0.009721f
C1625 DVSS.n1570 VSS 0.019442f
C1626 DVSS.n1571 VSS 0.019442f
C1627 DVSS.n1572 VSS 0.019442f
C1628 DVSS.n1573 VSS 0.019442f
C1629 DVSS.n1574 VSS 0.019442f
C1630 DVSS.n1575 VSS 0.019442f
C1631 DVSS.n1576 VSS 0.019442f
C1632 DVSS.n1577 VSS 0.019442f
C1633 DVSS.n1578 VSS 0.019442f
C1634 DVSS.n1579 VSS 0.019442f
C1635 DVSS.n1580 VSS 0.019442f
C1636 DVSS.n1581 VSS 0.019442f
C1637 DVSS.n1582 VSS 0.019442f
C1638 DVSS.n1583 VSS 0.019442f
C1639 DVSS.n1584 VSS 0.019442f
C1640 DVSS.n1585 VSS 0.019442f
C1641 DVSS.n1586 VSS 0.019442f
C1642 DVSS.n1587 VSS 0.019442f
C1643 DVSS.n1588 VSS 0.019442f
C1644 DVSS.n1589 VSS 0.019442f
C1645 DVSS.n1590 VSS 0.019442f
C1646 DVSS.n1591 VSS 0.185235f
C1647 DVSS.n1592 VSS 0.014497f
C1648 DVSS.n1593 VSS 0.016444f
C1649 DVSS.n1594 VSS 0.018232f
C1650 DVSS.n1595 VSS 0.018232f
C1651 DVSS.n1596 VSS 1.13742f
C1652 DVSS.n1597 VSS 1.13742f
C1653 DVSS.n1598 VSS 0.018232f
C1654 DVSS.n1599 VSS 0.018232f
C1655 DVSS.n1600 VSS 0.018232f
C1656 DVSS.n1601 VSS 0.031816f
C1657 DVSS.n1602 VSS 0.063632f
C1658 DVSS.n1603 VSS 0.018232f
C1659 DVSS.n1604 VSS 1.13742f
C1660 DVSS.n1605 VSS 0.018232f
C1661 DVSS.n1606 VSS 0.018232f
C1662 DVSS.n1607 VSS 0.016444f
C1663 DVSS.n1608 VSS 0.018232f
C1664 DVSS.n1609 VSS 1.13742f
C1665 DVSS.n1610 VSS 0.018232f
C1666 DVSS.n1611 VSS 0.018232f
C1667 DVSS.n1612 VSS 0.063632f
C1668 DVSS.n1613 VSS 0.018232f
C1669 DVSS.n1614 VSS 1.13742f
C1670 DVSS.n1615 VSS 0.018232f
C1671 DVSS.n1616 VSS 0.018232f
C1672 DVSS.n1617 VSS 0.016444f
C1673 DVSS.n1618 VSS 0.018232f
C1674 DVSS.n1619 VSS 1.13742f
C1675 DVSS.n1620 VSS 0.018232f
C1676 DVSS.n1621 VSS 0.018232f
C1677 DVSS.n1622 VSS 0.063632f
C1678 DVSS.n1623 VSS 0.018232f
C1679 DVSS.n1624 VSS 1.13742f
C1680 DVSS.n1625 VSS 0.018232f
C1681 DVSS.n1626 VSS 0.018232f
C1682 DVSS.n1627 VSS 0.016444f
C1683 DVSS.n1628 VSS 0.018232f
C1684 DVSS.n1629 VSS 1.13742f
C1685 DVSS.n1630 VSS 0.018232f
C1686 DVSS.n1631 VSS 0.018232f
C1687 DVSS.n1632 VSS 0.063632f
C1688 DVSS.n1633 VSS 0.018232f
C1689 DVSS.n1634 VSS 1.13742f
C1690 DVSS.n1635 VSS 0.018232f
C1691 DVSS.n1636 VSS 0.018232f
C1692 DVSS.n1637 VSS 0.016444f
C1693 DVSS.n1638 VSS 0.018232f
C1694 DVSS.n1639 VSS 1.13742f
C1695 DVSS.n1640 VSS 0.018232f
C1696 DVSS.n1641 VSS 0.018232f
C1697 DVSS.n1642 VSS 0.049398f
C1698 DVSS.n1643 VSS 0.063632f
C1699 DVSS.n1644 VSS 0.018232f
C1700 DVSS.n1645 VSS 1.13742f
C1701 DVSS.n1646 VSS 0.018232f
C1702 DVSS.n1647 VSS 0.018232f
C1703 DVSS.n1648 VSS 0.018232f
C1704 DVSS.n1649 VSS 0.014497f
C1705 DVSS.n1650 VSS 0.009721f
C1706 DVSS.n1651 VSS 0.068047f
C1707 DVSS.n1652 VSS 0.009721f
C1708 DVSS.n1653 VSS 0.019442f
C1709 DVSS.n1654 VSS 0.019442f
C1710 DVSS.n1655 VSS 0.019442f
C1711 DVSS.n1656 VSS 0.019442f
C1712 DVSS.n1657 VSS 0.15585f
C1713 DVSS.n1658 VSS 0.15585f
C1714 DVSS.n1659 VSS 0.15585f
C1715 DVSS.n1660 VSS 0.15585f
C1716 DVSS.n1661 VSS 0.15585f
C1717 DVSS.n1662 VSS 0.15585f
C1718 DVSS.n1663 VSS 0.15585f
C1719 DVSS.n1664 VSS 0.15585f
C1720 DVSS.n1665 VSS 0.15585f
C1721 DVSS.n1666 VSS 0.15585f
C1722 DVSS.n1667 VSS 0.15585f
C1723 DVSS.n1668 VSS 0.15585f
C1724 DVSS.n1669 VSS 0.15585f
C1725 DVSS.n1670 VSS 0.15585f
C1726 DVSS.n1671 VSS 0.15585f
C1727 DVSS.n1672 VSS 0.15585f
C1728 DVSS.n1673 VSS 0.15585f
C1729 DVSS.n1674 VSS 0.15585f
C1730 DVSS.n1675 VSS 0.009721f
C1731 DVSS.n1676 VSS 0.019442f
C1732 DVSS.n1677 VSS 0.019442f
C1733 DVSS.n1678 VSS 0.019442f
C1734 DVSS.n1679 VSS 0.019442f
C1735 DVSS.n1680 VSS 0.009721f
C1736 DVSS.n1681 VSS 0.019442f
C1737 DVSS.n1682 VSS 0.019442f
C1738 DVSS.n1683 VSS 0.019442f
C1739 DVSS.n1684 VSS 0.019442f
C1740 DVSS.n1685 VSS 0.009721f
C1741 DVSS.n1686 VSS 0.127863f
C1742 DVSS.n1687 VSS 0.009721f
C1743 DVSS.n1688 VSS 0.019442f
C1744 DVSS.n1689 VSS 0.019442f
C1745 DVSS.n1690 VSS 0.019442f
C1746 DVSS.n1691 VSS 0.019442f
C1747 DVSS.n1692 VSS 0.019442f
C1748 DVSS.n1693 VSS 0.019442f
C1749 DVSS.n1694 VSS 0.019442f
C1750 DVSS.n1695 VSS 0.019442f
C1751 DVSS.n1696 VSS 0.077925f
C1752 DVSS.n1697 VSS 0.15585f
C1753 DVSS.n1698 VSS 0.15585f
C1754 DVSS.n1699 VSS 0.15585f
C1755 DVSS.n1700 VSS 0.15585f
C1756 DVSS.n1701 VSS 0.15585f
C1757 DVSS.n1702 VSS 0.15585f
C1758 DVSS.n1703 VSS 0.15585f
C1759 DVSS.n1704 VSS 0.15585f
C1760 DVSS.n1705 VSS 0.15585f
C1761 DVSS.n1706 VSS 0.15585f
C1762 DVSS.n1707 VSS 0.15585f
C1763 DVSS.n1708 VSS 0.15585f
C1764 DVSS.n1709 VSS 0.15585f
C1765 DVSS.n1710 VSS 0.15585f
C1766 DVSS.n1711 VSS 0.15585f
C1767 DVSS.n1712 VSS 0.15585f
C1768 DVSS.n1713 VSS 0.077925f
C1769 DVSS.n1714 VSS 0.15585f
C1770 DVSS.n1715 VSS 0.15585f
C1771 DVSS.n1716 VSS 0.15585f
C1772 DVSS.n1717 VSS 0.15585f
C1773 DVSS.n1718 VSS 0.013092f
C1774 DVSS.n1719 VSS 0.009721f
C1775 DVSS.n1720 VSS 0.068047f
C1776 DVSS.n1722 VSS 0.009721f
C1777 DVSS.n1723 VSS 0.019442f
C1778 DVSS.n1724 VSS 0.019442f
C1779 DVSS.n1725 VSS 0.019442f
C1780 DVSS.n1726 VSS 0.009721f
C1781 DVSS.n1727 VSS 0.010348f
C1782 DVSS.n1728 VSS 0.009721f
C1783 DVSS.n1729 VSS 0.009721f
C1784 DVSS.n1730 VSS 0.183412f
C1785 DVSS.n1731 VSS 0.016071f
C1786 DVSS.n1733 VSS 0.026052f
C1787 DVSS.n1734 VSS 0.016185f
C1788 DVSS.n1735 VSS 0.04307f
C1789 DVSS.n1736 VSS 0.016185f
C1790 DVSS.n1737 VSS 0.210064f
C1791 DVSS.n1739 VSS 0.074084f
C1792 DVSS.n1740 VSS 0.077925f
C1793 DVSS.n1742 VSS 0.026052f
C1794 DVSS.n1743 VSS 0.068047f
C1795 DVSS.n1745 VSS 0.052105f
C1796 DVSS.n1748 VSS 0.145809f
C1797 DVSS.n1749 VSS 0.052105f
C1798 DVSS.n1750 VSS 0.052105f
C1799 DVSS.n1752 VSS 0.077925f
C1800 DVSS.n1754 VSS 0.355784f
C1801 DVSS.n1755 VSS 0.018275f
C1802 DVSS.n1756 VSS 0.054406f
C1803 DVSS.n1757 VSS 0.009721f
C1804 DVSS.n1759 VSS 0.048557f
C1805 DVSS.n1760 VSS 0.755948f
C1806 DVSS.n1761 VSS 0.01079f
C1807 DVSS.n1762 VSS 0.871379f
C1808 DVSS.t24 VSS 13.3026f
C1809 DVSS.n1763 VSS 0.051264f
C1810 DVSS.n1764 VSS 0.671452f
C1811 DVSS.n1765 VSS 0.051264f
C1812 DVSS.n1766 VSS 0.871379f
C1813 DVSS.n1767 VSS 0.755948f
C1814 DVSS.n1768 VSS 0.183412f
C1815 DVSS.n1769 VSS 0.048557f
C1816 DVSS.n1770 VSS 0.355784f
C1817 DVSS.n1771 VSS 0.062324f
C1818 DVSS.n1772 VSS 0.009721f
C1819 DVSS.n1774 VSS 0.170181f
C1820 DVSS.n1778 VSS 0.027413f
C1821 DVSS.n1779 VSS 0.051264f
C1822 DVSS.n1780 VSS 0.671452f
C1823 DVSS.n1781 VSS 0.755948f
C1824 DVSS.n1782 VSS 0.048557f
C1825 DVSS.n1783 VSS 1.33324f
C1826 DVSS.n1784 VSS 0.755948f
C1827 DVSS.n1785 VSS 0.481904f
C1828 DVSS.n1786 VSS 0.183412f
C1829 DVSS.n1787 VSS 0.355784f
C1830 DVSS.n1788 VSS 0.009721f
C1831 DVSS.n1789 VSS 0.009721f
C1832 DVSS.n1790 VSS 0.009721f
C1833 DVSS.n1791 VSS 0.264848f
C1834 DVSS.n1792 VSS 0.355784f
C1835 DVSS.n1793 VSS 0.264848f
C1836 DVSS.n1794 VSS 0.009721f
C1837 DVSS.n1796 VSS 0.009721f
C1838 DVSS.n1797 VSS 0.009721f
C1839 DVSS.n1798 VSS 0.077925f
C1840 DVSS.n1799 VSS 0.077925f
C1841 DVSS.n1801 VSS 0.077925f
C1842 DVSS.n1802 VSS 0.077925f
C1843 DVSS.n1803 VSS 0.49201f
C1844 DVSS.n1804 VSS 0.01017f
C1845 DVSS.n1805 VSS 0.016444f
C1846 DVSS.n1806 VSS 0.018232f
C1847 DVSS.n1807 VSS 0.018232f
C1848 DVSS.n1808 VSS 1.13742f
C1849 DVSS.n1809 VSS 1.13742f
C1850 DVSS.n1810 VSS 0.018232f
C1851 DVSS.n1811 VSS 0.018232f
C1852 DVSS.n1812 VSS 0.018232f
C1853 DVSS.n1813 VSS 0.008222f
C1854 DVSS.n1814 VSS 0.016444f
C1855 DVSS.n1815 VSS 0.018232f
C1856 DVSS.n1816 VSS 1.13742f
C1857 DVSS.n1817 VSS 0.018232f
C1858 DVSS.n1818 VSS 0.018232f
C1859 DVSS.n1819 VSS 0.018232f
C1860 DVSS.n1820 VSS 0.058608f
C1861 DVSS.n1821 VSS 0.063632f
C1862 DVSS.n1822 VSS 0.018232f
C1863 DVSS.n1823 VSS 1.13742f
C1864 DVSS.n1824 VSS 0.018232f
C1865 DVSS.n1825 VSS 0.018232f
C1866 DVSS.n1826 VSS 0.016444f
C1867 DVSS.n1827 VSS 0.018232f
C1868 DVSS.n1828 VSS 1.13742f
C1869 DVSS.n1829 VSS 0.018232f
C1870 DVSS.n1830 VSS 0.018232f
C1871 DVSS.n1831 VSS 0.063632f
C1872 DVSS.n1832 VSS 0.018232f
C1873 DVSS.n1833 VSS 1.13742f
C1874 DVSS.n1834 VSS 0.018232f
C1875 DVSS.n1835 VSS 0.018232f
C1876 DVSS.n1836 VSS 0.016444f
C1877 DVSS.n1837 VSS 0.018232f
C1878 DVSS.n1838 VSS 1.13742f
C1879 DVSS.n1839 VSS 0.018232f
C1880 DVSS.n1840 VSS 0.018232f
C1881 DVSS.n1841 VSS 0.063632f
C1882 DVSS.n1842 VSS 0.018232f
C1883 DVSS.n1843 VSS 1.13742f
C1884 DVSS.n1844 VSS 0.018232f
C1885 DVSS.n1845 VSS 0.018232f
C1886 DVSS.n1846 VSS 0.016444f
C1887 DVSS.n1847 VSS 0.018232f
C1888 DVSS.n1848 VSS 1.13742f
C1889 DVSS.n1849 VSS 0.018232f
C1890 DVSS.n1850 VSS 0.018232f
C1891 DVSS.n1851 VSS 0.063632f
C1892 DVSS.n1852 VSS 0.018232f
C1893 DVSS.n1853 VSS 1.13742f
C1894 DVSS.n1854 VSS 0.018232f
C1895 DVSS.n1855 VSS 0.018232f
C1896 DVSS.n1856 VSS 0.016444f
C1897 DVSS.n1857 VSS 0.018232f
C1898 DVSS.n1858 VSS 1.13742f
C1899 DVSS.n1859 VSS 0.018232f
C1900 DVSS.n1860 VSS 0.018232f
C1901 DVSS.n1861 VSS 0.046432f
C1902 DVSS.n1862 VSS 0.052105f
C1903 DVSS.n1863 VSS 1.22005f
C1904 DVSS.n1864 VSS 0.034607f
C1905 DVSS.n1865 VSS 0.052105f
C1906 DVSS.n1866 VSS 0.052105f
C1907 DVSS.n1867 VSS 0.026052f
C1908 DVSS.n1870 VSS 0.031816f
C1909 DVSS.n1872 VSS 0.031816f
C1910 DVSS.n1873 VSS 0.046432f
C1911 DVSS.n1874 VSS 0.016466f
C1912 DVSS.n1876 VSS 0.018232f
C1913 DVSS.n1877 VSS 0.018232f
C1914 DVSS.n1878 VSS 1.13742f
C1915 DVSS.n1879 VSS 1.13742f
C1916 DVSS.n1880 VSS 0.018232f
C1917 DVSS.n1881 VSS 0.018232f
C1918 DVSS.n1882 VSS 0.018232f
C1919 DVSS.n1883 VSS 0.012333f
C1920 DVSS.n1884 VSS 0.016444f
C1921 DVSS.n1885 VSS 0.018232f
C1922 DVSS.n1886 VSS 1.13742f
C1923 DVSS.n1887 VSS 0.018232f
C1924 DVSS.n1888 VSS 0.018232f
C1925 DVSS.n1889 VSS 0.059446f
C1926 DVSS.n1890 VSS 0.063632f
C1927 DVSS.n1891 VSS 0.018232f
C1928 DVSS.n1892 VSS 1.13742f
C1929 DVSS.n1893 VSS 0.018232f
C1930 DVSS.n1894 VSS 0.018232f
C1931 DVSS.n1895 VSS 0.016444f
C1932 DVSS.n1896 VSS 0.018232f
C1933 DVSS.n1897 VSS 1.13742f
C1934 DVSS.n1898 VSS 0.018232f
C1935 DVSS.n1899 VSS 0.018232f
C1936 DVSS.n1900 VSS 0.038514f
C1937 DVSS.n1901 VSS 0.018232f
C1938 DVSS.n1902 VSS 1.13742f
C1939 DVSS.n1903 VSS 0.018232f
C1940 DVSS.n1904 VSS 0.018232f
C1941 DVSS.n1905 VSS 0.016444f
C1942 DVSS.n1906 VSS 0.018232f
C1943 DVSS.n1907 VSS 1.13742f
C1944 DVSS.n1908 VSS 0.018232f
C1945 DVSS.n1909 VSS 0.018232f
C1946 DVSS.n1910 VSS 0.063632f
C1947 DVSS.n1911 VSS 0.018232f
C1948 DVSS.n1912 VSS 1.13742f
C1949 DVSS.n1913 VSS 0.018232f
C1950 DVSS.n1914 VSS 0.018232f
C1951 DVSS.n1915 VSS 0.016444f
C1952 DVSS.n1916 VSS 0.018232f
C1953 DVSS.n1917 VSS 1.13742f
C1954 DVSS.n1918 VSS 0.018232f
C1955 DVSS.n1919 VSS 0.018232f
C1956 DVSS.n1920 VSS 0.063632f
C1957 DVSS.n1921 VSS 0.018232f
C1958 DVSS.n1922 VSS 1.13742f
C1959 DVSS.n1923 VSS 0.018232f
C1960 DVSS.n1924 VSS 0.018232f
C1961 DVSS.n1925 VSS 0.016444f
C1962 DVSS.n1926 VSS 0.018232f
C1963 DVSS.n1927 VSS 1.13742f
C1964 DVSS.n1928 VSS 0.018232f
C1965 DVSS.n1929 VSS 0.018232f
C1966 DVSS.n1930 VSS 0.018232f
C1967 DVSS.n1931 VSS 0.008222f
C1968 DVSS.n1932 VSS 0.018232f
C1969 DVSS.n1933 VSS 0.016444f
C1970 DVSS.n1934 VSS 0.018232f
C1971 DVSS.n1935 VSS 0.016444f
C1972 DVSS.n1936 VSS 0.016444f
C1973 DVSS.n1937 VSS 0.018232f
C1974 DVSS.n1938 VSS 0.016444f
C1975 DVSS.n1939 VSS 0.016444f
C1976 DVSS.n1940 VSS 0.018232f
C1977 DVSS.n1941 VSS 0.016444f
C1978 DVSS.n1942 VSS 0.016444f
C1979 DVSS.n1943 VSS 0.018232f
C1980 DVSS.n1944 VSS 0.016444f
C1981 DVSS.n1945 VSS 0.016444f
C1982 DVSS.n1946 VSS 0.018232f
C1983 DVSS.n1947 VSS 0.016444f
C1984 DVSS.n1948 VSS 0.016444f
C1985 DVSS.n1949 VSS 0.018232f
C1986 DVSS.n1950 VSS 0.016444f
C1987 DVSS.n1951 VSS 0.016444f
C1988 DVSS.n1952 VSS 0.018232f
C1989 DVSS.n1953 VSS 0.016444f
C1990 DVSS.n1954 VSS 0.016444f
C1991 DVSS.n1955 VSS 0.018232f
C1992 DVSS.n1956 VSS 0.016444f
C1993 DVSS.n1957 VSS 0.016444f
C1994 DVSS.n1958 VSS 0.018232f
C1995 DVSS.n1959 VSS 0.016444f
C1996 DVSS.n1960 VSS 0.016444f
C1997 DVSS.n1961 VSS 0.012333f
C1998 DVSS.n1962 VSS 1.13742f
C1999 DVSS.n1963 VSS 0.018232f
C2000 DVSS.t2 VSS 0.519282f
C2001 DVSS.n1964 VSS 0.98199f
C2002 DVSS.t4 VSS 0.519282f
C2003 DVSS.n1965 VSS 0.98199f
C2004 DVSS.n1966 VSS 0.791465f
C2005 DVSS.n1967 VSS 0.017862f
C2006 DVSS.n1968 VSS 0.018232f
C2007 DVSS.n1969 VSS 0.018232f
C2008 DVSS.n1970 VSS 0.016444f
C2009 DVSS.n1971 VSS 0.647107f
C2010 DVSS.n1974 VSS 0.068047f
C2011 DVSS.n1975 VSS 0.052105f
C2012 DVSS.n1976 VSS 0.052105f
C2013 DVSS.n1977 VSS 0.052105f
C2014 DVSS.n1978 VSS 0.052105f
C2015 DVSS.n1979 VSS 0.052105f
C2016 DVSS.n1980 VSS 0.091644f
C2017 DVSS.n1981 VSS 0.052105f
C2018 DVSS.n1982 VSS 0.052105f
C2019 DVSS.n1983 VSS 0.052105f
C2020 DVSS.n1988 VSS 0.071889f
C2021 DVSS.n1994 VSS 0.077925f
C2022 DVSS.n1995 VSS 0.15585f
C2023 DVSS.n1996 VSS 0.15585f
C2024 DVSS.n1997 VSS 0.15585f
C2025 DVSS.n1998 VSS 0.15585f
C2026 DVSS.n1999 VSS 0.15585f
C2027 DVSS.n2000 VSS 0.15585f
C2028 DVSS.n2001 VSS 0.15585f
C2029 DVSS.n2002 VSS 0.15585f
C2030 DVSS.n2003 VSS 0.15585f
C2031 DVSS.n2004 VSS 0.15585f
C2032 DVSS.n2005 VSS 0.15585f
C2033 DVSS.n2006 VSS 0.15585f
C2034 DVSS.n2007 VSS 0.15585f
C2035 DVSS.n2008 VSS 0.15585f
C2036 DVSS.n2009 VSS 0.15585f
C2037 DVSS.n2010 VSS 0.15585f
C2038 DVSS.n2011 VSS 0.077925f
C2039 DVSS.n2012 VSS 0.15585f
C2040 DVSS.n2013 VSS 0.15585f
C2041 DVSS.n2014 VSS 0.15585f
C2042 DVSS.n2015 VSS 0.15585f
C2043 DVSS.n2016 VSS 0.068047f
C2044 DVSS.n2017 VSS 0.009721f
C2045 DVSS.n2018 VSS 0.019442f
C2046 DVSS.n2019 VSS 0.019442f
C2047 DVSS.n2020 VSS 0.019442f
C2048 DVSS.n2021 VSS 0.019442f
C2049 DVSS.n2022 VSS 0.019442f
C2050 DVSS.n2023 VSS 0.019442f
C2051 DVSS.n2024 VSS 0.019442f
C2052 DVSS.n2025 VSS 0.019442f
C2053 DVSS.n2026 VSS 0.009721f
C2054 DVSS.n2027 VSS 0.145816f
C2055 DVSS.n2028 VSS 0.321029f
C2056 DVSS.n2029 VSS 0.019442f
C2057 DVSS.n2030 VSS 0.019442f
C2058 DVSS.n2031 VSS 0.019442f
C2059 DVSS.n2032 VSS 0.019442f
C2060 DVSS.n2033 VSS 0.019442f
C2061 DVSS.n2034 VSS 0.019442f
C2062 DVSS.n2035 VSS 0.019442f
C2063 DVSS.n2036 VSS 0.019442f
C2064 DVSS.n2037 VSS 0.019442f
C2065 DVSS.n2038 VSS 0.019442f
C2066 DVSS.n2039 VSS 0.019442f
C2067 DVSS.n2040 VSS 0.333965f
C2068 DVSS.n2041 VSS 0.333965f
C2069 DVSS.n2042 VSS 0.333965f
C2070 DVSS.n2043 VSS 0.333965f
C2071 DVSS.n2044 VSS 0.333965f
C2072 DVSS.n2045 VSS 0.333965f
C2073 DVSS.n2046 VSS 0.333965f
C2074 DVSS.n2047 VSS 0.333965f
C2075 DVSS.n2048 VSS 0.333965f
C2076 DVSS.n2049 VSS 0.333965f
C2077 DVSS.n2050 VSS 0.333965f
C2078 DVSS.n2051 VSS 0.333965f
C2079 DVSS.n2052 VSS 0.333965f
C2080 DVSS.n2053 VSS 0.333965f
C2081 DVSS.n2054 VSS 5.56962f
C2082 DVSS.n2055 VSS 0.333965f
C2083 DVSS.n2056 VSS 0.145816f
C2084 DVSS.n2057 VSS 0.241458f
C2085 DVSS.n2058 VSS 0.019442f
C2086 DVSS.n2059 VSS 0.019442f
C2087 DVSS.n2060 VSS 0.019442f
C2088 DVSS.n2061 VSS 0.019442f
C2089 DVSS.n2062 VSS 0.019442f
C2090 DVSS.n2063 VSS 0.019442f
C2091 DVSS.n2064 VSS 0.019442f
C2092 DVSS.n2065 VSS 0.019442f
C2093 DVSS.n2066 VSS 0.019442f
C2094 DVSS.n2067 VSS 0.019442f
C2095 DVSS.n2068 VSS 0.019442f
C2096 DVSS.n2069 VSS 0.009721f
C2097 DVSS.n2070 VSS 0.068047f
C2098 DVSS.n2071 VSS 0.009721f
C2099 DVSS.n2072 VSS 0.019442f
C2100 DVSS.n2073 VSS 0.019442f
C2101 DVSS.n2074 VSS 0.019442f
C2102 DVSS.n2075 VSS 0.019442f
C2103 DVSS.n2076 VSS 0.15585f
C2104 DVSS.n2077 VSS 0.506941f
C2105 DVSS.n2078 VSS 0.15585f
C2106 DVSS.n2079 VSS 0.019442f
C2107 DVSS.n2080 VSS 0.019442f
C2108 DVSS.n2081 VSS 0.019442f
C2109 DVSS.n2082 VSS 0.019442f
C2110 DVSS.n2083 VSS 0.009721f
C2111 DVSS.n2084 VSS 0.068047f
C2112 DVSS.n2085 VSS 0.009721f
C2113 DVSS.n2086 VSS 0.019442f
C2114 DVSS.n2087 VSS 0.019442f
C2115 DVSS.n2088 VSS 0.019442f
C2116 DVSS.n2089 VSS 0.019442f
C2117 DVSS.n2090 VSS 0.15585f
C2118 DVSS.n2091 VSS 0.506941f
C2119 DVSS.n2092 VSS 0.15585f
C2120 DVSS.n2093 VSS 0.019442f
C2121 DVSS.n2094 VSS 0.019442f
C2122 DVSS.n2095 VSS 0.019442f
C2123 DVSS.n2096 VSS 0.019442f
C2124 DVSS.n2097 VSS 0.009721f
C2125 DVSS.n2098 VSS 0.068047f
C2126 DVSS.n2099 VSS 0.009721f
C2127 DVSS.n2100 VSS 0.019442f
C2128 DVSS.n2101 VSS 0.008467f
C2129 DVSS.n2102 VSS 0.009721f
C2130 DVSS.n2103 VSS 0.125668f
C2131 DVSS.n2104 VSS 0.008467f
C2132 DVSS.n2105 VSS 0.013014f
C2133 DVSS.n2106 VSS 3.71965f
C2134 DVSS.n2107 VSS 0.163454f
C2135 DVSS.n2108 VSS 0.019442f
C2136 DVSS.n2109 VSS 0.036571f
C2137 DVSS.n2110 VSS 0.009721f
C2138 DVSS.t27 VSS 0.311996f
C2139 DVSS.n2111 VSS 0.599743f
C2140 DVSS.n2112 VSS 0.009721f
C2141 DVSS.n2114 VSS 0.008467f
C2142 DVSS.n2115 VSS 0.018658f
C2143 DVSS.n2116 VSS 0.026052f
C2144 DVSS.n2117 VSS 0.020834f
C2145 DVSS.t25 VSS 0.311996f
C2146 DVSS.n2118 VSS 0.599743f
C2147 DVSS.n2119 VSS 0.255569f
C2148 DVSS.n2120 VSS 0.01709f
C2149 DVSS.n2121 VSS 0.026052f
C2150 DVSS.n2122 VSS 0.022691f
C2151 DVSS.n2123 VSS -0.441359f
C2152 DVSS.n2124 VSS 0.050004f
C2153 DVSS.n2125 VSS 0.009721f
C2154 DVSS.n2127 VSS 0.008467f
C2155 DVSS.n2128 VSS 0.018658f
C2156 DVSS.n2129 VSS 0.009721f
C2157 DVSS.n2131 VSS 0.008467f
C2158 DVSS.n2132 VSS 0.018658f
C2159 DVSS.n2133 VSS 0.160836f
C2160 DVSS.n2134 VSS 11.080799f
C2161 DVSS.n2135 VSS 5.83802f
C2162 DVSS.n2136 VSS 2.75825f
C2163 DVSS.n2137 VSS 1.73511f
C2164 DVSS.n2138 VSS 0.048129f
C2165 DVSS.n2139 VSS 0.013406f
C2166 DVSS.n2140 VSS 1.73511f
C2167 DVSS.n2141 VSS 0.008213f
C2168 DVSS.n2142 VSS 1.76722f
C2169 DVSS.n2143 VSS 0.15585f
C2170 DVSS.n2144 VSS 0.15585f
C2171 DVSS.n2145 VSS 0.15585f
C2172 DVSS.n2146 VSS 0.15585f
C2173 DVSS.n2147 VSS 0.15585f
C2174 DVSS.n2148 VSS 0.15585f
C2175 DVSS.n2149 VSS 0.15585f
C2176 DVSS.n2150 VSS 0.15585f
C2177 DVSS.n2151 VSS 0.15585f
C2178 DVSS.n2152 VSS 0.15585f
C2179 DVSS.n2153 VSS 0.15585f
C2180 DVSS.n2154 VSS 0.15585f
C2181 DVSS.n2155 VSS 0.15585f
C2182 DVSS.n2156 VSS 0.15585f
C2183 DVSS.n2157 VSS 0.15585f
C2184 DVSS.n2158 VSS 0.15585f
C2185 DVSS.n2159 VSS 0.15585f
C2186 DVSS.n2160 VSS 0.15585f
C2187 DVSS.n2161 VSS 0.15585f
C2188 DVSS.n2162 VSS 0.15585f
C2189 DVSS.n2163 VSS 0.15585f
C2190 DVSS.n2164 VSS 0.15585f
C2191 DVSS.n2165 VSS 0.15585f
C2192 DVSS.n2166 VSS 0.15585f
C2193 DVSS.n2167 VSS 0.15585f
C2194 DVSS.n2168 VSS 0.15585f
C2195 DVSS.n2169 VSS 0.15585f
C2196 DVSS.n2170 VSS 0.15585f
C2197 DVSS.n2171 VSS 0.15585f
C2198 DVSS.n2172 VSS 0.15585f
C2199 DVSS.n2173 VSS 0.15585f
C2200 DVSS.n2174 VSS 0.15585f
C2201 DVSS.n2175 VSS 0.15585f
C2202 DVSS.n2176 VSS 0.15585f
C2203 DVSS.n2177 VSS 0.15585f
C2204 DVSS.n2178 VSS 0.15585f
C2205 DVSS.n2179 VSS 0.15585f
C2206 DVSS.n2180 VSS 0.15585f
C2207 DVSS.n2181 VSS 0.15585f
C2208 DVSS.n2182 VSS 0.15585f
C2209 DVSS.n2183 VSS 0.15585f
C2210 DVSS.n2184 VSS 0.15585f
C2211 DVSS.n2185 VSS 0.15585f
C2212 DVSS.n2186 VSS 0.15585f
C2213 DVSS.n2187 VSS 0.15585f
C2214 DVSS.n2188 VSS 0.15585f
C2215 DVSS.n2189 VSS 0.15585f
C2216 DVSS.n2190 VSS 0.15585f
C2217 DVSS.n2191 VSS 0.15585f
C2218 DVSS.n2192 VSS 0.15585f
C2219 DVSS.n2193 VSS 0.15585f
C2220 DVSS.n2194 VSS 0.15585f
C2221 DVSS.n2195 VSS 0.15585f
C2222 DVSS.n2196 VSS 0.15585f
C2223 DVSS.n2197 VSS 0.15585f
C2224 DVSS.n2198 VSS 0.15585f
C2225 DVSS.n2199 VSS 0.15585f
C2226 DVSS.n2200 VSS 0.15585f
C2227 DVSS.n2201 VSS 0.15585f
C2228 DVSS.n2202 VSS 0.15585f
C2229 DVSS.n2203 VSS 0.15585f
C2230 DVSS.n2204 VSS 0.15585f
C2231 DVSS.n2205 VSS 0.15585f
C2232 DVSS.n2206 VSS 0.15585f
C2233 DVSS.n2207 VSS 0.15585f
C2234 DVSS.n2208 VSS 0.15585f
C2235 DVSS.n2209 VSS 0.15585f
C2236 DVSS.n2210 VSS 0.15585f
C2237 DVSS.n2211 VSS 0.15585f
C2238 DVSS.n2212 VSS 0.15585f
C2239 DVSS.n2213 VSS 0.15585f
C2240 DVSS.n2214 VSS 0.15585f
C2241 DVSS.n2215 VSS 0.15585f
C2242 DVSS.n2216 VSS 0.15585f
C2243 DVSS.n2217 VSS 0.15585f
C2244 DVSS.n2218 VSS 0.15585f
C2245 DVSS.n2219 VSS 0.15585f
C2246 DVSS.n2220 VSS 0.15585f
C2247 DVSS.n2221 VSS 0.15585f
C2248 DVSS.n2222 VSS 0.15585f
C2249 DVSS.n2223 VSS 0.15585f
C2250 DVSS.n2224 VSS 0.15585f
C2251 DVSS.n2225 VSS 0.15585f
C2252 DVSS.n2226 VSS 0.15585f
C2253 DVSS.n2227 VSS 0.15585f
C2254 DVSS.n2228 VSS 0.15585f
C2255 DVSS.n2229 VSS 0.15585f
C2256 DVSS.n2230 VSS 0.15585f
C2257 DVSS.n2231 VSS 0.15585f
C2258 DVSS.n2232 VSS 0.15585f
C2259 DVSS.n2233 VSS 0.15585f
C2260 DVSS.n2234 VSS 0.15585f
C2261 DVSS.n2235 VSS 0.15585f
C2262 DVSS.n2236 VSS 0.15585f
C2263 DVSS.n2237 VSS 0.15585f
C2264 DVSS.n2238 VSS 0.15585f
C2265 DVSS.n2239 VSS 0.15585f
C2266 DVSS.n2240 VSS 0.15585f
C2267 DVSS.n2241 VSS 0.08012f
C2268 DVSS.n2242 VSS 0.15585f
C2269 DVSS.n2243 VSS 0.15585f
C2270 DVSS.n2244 VSS 0.28536f
C2271 DVSS.n2245 VSS 0.15585f
C2272 DVSS.n2246 VSS 0.15585f
C2273 DVSS.n2247 VSS 0.15585f
C2274 DVSS.n2248 VSS 0.29749f
C2275 DVSS.n2249 VSS 0.58172f
C2276 DVSS.n2250 VSS 0.153655f
C2277 DVSS.n2251 VSS 0.15585f
C2278 DVSS.n2252 VSS 0.093291f
C2279 DVSS.n2253 VSS 0.093291f
C2280 DVSS.n2254 VSS 0.140485f
C2281 DVSS.n2255 VSS 0.140485f
C2282 DVSS.n2256 VSS 0.15585f
C2283 DVSS.n2257 VSS 0.15585f
C2284 DVSS.n2258 VSS 0.15585f
C2285 DVSS.n2259 VSS 0.15585f
C2286 DVSS.n2260 VSS 0.15585f
C2287 DVSS.n2261 VSS 0.15585f
C2288 DVSS.n2262 VSS 0.15585f
C2289 DVSS.n2263 VSS 0.15585f
C2290 DVSS.n2264 VSS 0.15585f
C2291 DVSS.n2265 VSS 0.15585f
C2292 DVSS.n2266 VSS 0.15585f
C2293 DVSS.n2267 VSS 0.15585f
C2294 DVSS.n2268 VSS 0.15585f
C2295 DVSS.n2269 VSS 0.15585f
C2296 DVSS.n2270 VSS 0.15585f
C2297 DVSS.n2271 VSS 0.15585f
C2298 DVSS.n2272 VSS 0.15585f
C2299 DVSS.n2273 VSS 0.15585f
C2300 DVSS.n2274 VSS 0.15585f
C2301 DVSS.n2275 VSS 0.15585f
C2302 DVSS.n2276 VSS 0.082864f
C2303 DVSS.n2277 VSS 0.150911f
C2304 DVSS.n2278 VSS 0.15585f
C2305 DVSS.n2279 VSS 0.15585f
C2306 DVSS.n2280 VSS 0.15585f
C2307 DVSS.n2281 VSS 0.15585f
C2308 DVSS.n2282 VSS 0.15585f
C2309 DVSS.n2283 VSS 0.15585f
C2310 DVSS.n2284 VSS 0.15585f
C2311 DVSS.n2285 VSS 0.15585f
C2312 DVSS.n2286 VSS 0.15585f
C2313 DVSS.n2287 VSS 0.15585f
C2314 DVSS.n2288 VSS 0.15585f
C2315 DVSS.n2289 VSS 0.15585f
C2316 DVSS.n2290 VSS 0.15585f
C2317 DVSS.n2291 VSS 0.15585f
C2318 DVSS.n2292 VSS 0.15585f
C2319 DVSS.n2293 VSS 0.15585f
C2320 DVSS.n2294 VSS 0.15585f
C2321 DVSS.n2295 VSS 0.15585f
C2322 DVSS.n2296 VSS 0.15585f
C2323 DVSS.n2297 VSS 0.15585f
C2324 DVSS.n2298 VSS 0.15585f
C2325 DVSS.n2299 VSS 0.15585f
C2326 DVSS.n2300 VSS 0.15585f
C2327 DVSS.n2301 VSS 0.15585f
C2328 DVSS.n2302 VSS 0.15585f
C2329 DVSS.n2303 VSS 0.15585f
C2330 DVSS.n2304 VSS 0.15585f
C2331 DVSS.n2305 VSS 0.15585f
C2332 DVSS.n2306 VSS 0.15585f
C2333 DVSS.n2307 VSS 0.15585f
C2334 DVSS.n2308 VSS 0.15585f
C2335 DVSS.n2309 VSS 0.15585f
C2336 DVSS.n2310 VSS 0.15585f
C2337 DVSS.n2311 VSS 0.15585f
C2338 DVSS.n2312 VSS 0.15585f
C2339 DVSS.n2313 VSS 0.15585f
C2340 DVSS.n2314 VSS 0.15585f
C2341 DVSS.n2315 VSS 0.15585f
C2342 DVSS.n2316 VSS 0.15585f
C2343 DVSS.n2317 VSS 0.15585f
C2344 DVSS.n2318 VSS 0.15585f
C2345 DVSS.n2319 VSS 0.15585f
C2346 DVSS.n2320 VSS 0.15585f
C2347 DVSS.n2321 VSS 0.15585f
C2348 DVSS.n2322 VSS 0.15585f
C2349 DVSS.n2323 VSS 0.15585f
C2350 DVSS.n2324 VSS 0.15585f
C2351 DVSS.n2325 VSS 0.15585f
C2352 DVSS.n2326 VSS 0.15585f
C2353 DVSS.n2327 VSS 0.15585f
C2354 DVSS.n2328 VSS 0.15585f
C2355 DVSS.n2329 VSS 0.15585f
C2356 DVSS.n2330 VSS 0.15585f
C2357 DVSS.n2331 VSS 0.15585f
C2358 DVSS.n2332 VSS 0.15585f
C2359 DVSS.n2333 VSS 0.15585f
C2360 DVSS.n2334 VSS 0.15585f
C2361 DVSS.n2335 VSS 0.15585f
C2362 DVSS.n2336 VSS 0.15585f
C2363 DVSS.n2337 VSS 0.15585f
C2364 DVSS.n2338 VSS 0.15585f
C2365 DVSS.n2339 VSS 0.15585f
C2366 DVSS.n2340 VSS 0.15585f
C2367 DVSS.n2341 VSS 0.15585f
C2368 DVSS.n2342 VSS 0.15585f
C2369 DVSS.n2343 VSS 0.15585f
C2370 DVSS.n2344 VSS 0.15585f
C2371 DVSS.n2345 VSS 0.15585f
C2372 DVSS.n2346 VSS 0.15585f
C2373 DVSS.n2347 VSS 0.15585f
C2374 DVSS.n2348 VSS 0.15585f
C2375 DVSS.n2349 VSS 0.15585f
C2376 DVSS.n2350 VSS 0.15585f
C2377 DVSS.n2351 VSS 0.15585f
C2378 DVSS.n2352 VSS 0.15585f
C2379 DVSS.n2353 VSS 0.15585f
C2380 DVSS.n2354 VSS 0.15585f
C2381 DVSS.n2355 VSS 0.15585f
C2382 DVSS.n2356 VSS 0.15585f
C2383 DVSS.n2357 VSS 0.15585f
C2384 DVSS.n2358 VSS 0.15585f
C2385 DVSS.n2359 VSS 0.15585f
C2386 DVSS.n2360 VSS 0.15585f
C2387 DVSS.n2361 VSS 0.15585f
C2388 DVSS.n2362 VSS 0.15585f
C2389 DVSS.n2363 VSS 0.15585f
C2390 DVSS.n2364 VSS 0.15585f
C2391 DVSS.n2365 VSS 0.292976f
C2392 DVSS.n2366 VSS 0.15585f
C2393 DVSS.n2367 VSS 0.011149f
C2394 DVSS.n2368 VSS 0.010686f
C2395 DVSS.n2369 VSS 0.065194f
C2396 DVSS.n2370 VSS 0.635473f
C2397 DVSS.n2371 VSS 0.648801f
C2398 DVSS.n2372 VSS 0.919657f
C2399 DVSS.n2373 VSS 0.919657f
C2400 DVSS.n2374 VSS 0.648801f
C2401 DVSS.n2375 VSS 0.249142f
C2402 DVSS.n2376 VSS 0.249533f
C2403 DVSS.n2377 VSS 0.648801f
C2404 DVSS.n2378 VSS 1.62877f
C2405 DVSS.n2379 VSS 8.82012f
C2406 DVSS.n2380 VSS 2.59578f
C2407 DVSS.n2381 VSS 0.186424f
C2408 DVSS.n2382 VSS 0.559787f
C2409 DVSS.n2383 VSS 0.26825f
C2410 DVSS.n2384 VSS 0.648801f
C2411 DVSS.n2385 VSS 0.919657f
C2412 DVSS.n2386 VSS 0.919657f
C2413 DVSS.n2387 VSS 0.919657f
C2414 DVSS.n2388 VSS 0.648801f
C2415 DVSS.n2389 VSS 0.249533f
C2416 DVSS.n2390 VSS 0.249533f
C2417 DVSS.n2391 VSS 0.249533f
C2418 DVSS.n2392 VSS 0.648801f
C2419 DVSS.n2393 VSS 0.009721f
C2420 DVSS.n2394 VSS 0.009721f
C2421 DVSS.n2395 VSS -0.483269f
C2422 DVSS.n2396 VSS 0.058198f
C2423 DVSS.n2397 VSS 0.027943f
C2424 DVSS.n2398 VSS 0.021715f
C2425 DVSS.n2399 VSS 0.071134f
C2426 DVSS.n2400 VSS 0.071134f
C2427 DVSS.n2401 VSS 0.077925f
C2428 DVSS.n2402 VSS 0.068047f
C2429 DVSS.n2403 VSS 0.009721f
C2430 DVSS.n2404 VSS 0.091644f
C2431 DVSS.n2405 VSS 0.009721f
C2432 DVSS.n2406 VSS 0.016185f
C2433 DVSS.n2407 VSS 0.212831f
C2434 DVSS.n2409 VSS 0.01079f
C2435 DVSS.n2410 VSS 0.016185f
C2436 DVSS.n2414 VSS 0.355784f
C2437 DVSS.n2416 VSS 0.027413f
C2438 DVSS.n2417 VSS 1.33324f
C2439 DVSS.n2418 VSS 0.018275f
C2440 DVSS.n2419 VSS 0.170181f
C2441 DVSS.n2420 VSS 0.027413f
C2442 DVSS.n2421 VSS 0.052105f
C2443 DVSS.n2422 VSS 0.355784f
C2444 DVSS.n2423 VSS 0.167029f
C2445 DVSS.n2424 VSS 0.009721f
C2446 DVSS.n2425 VSS 0.068047f
C2447 DVSS.n2426 VSS 0.009721f
C2448 DVSS.n2427 VSS 0.019442f
C2449 DVSS.n2428 VSS 0.009721f
C2450 DVSS.n2429 VSS 0.149814f
C2451 DVSS.n2430 VSS 0.009721f
C2452 DVSS.n2431 VSS 0.008467f
C2453 DVSS.n2432 VSS 0.013014f
C2454 DVSS.n2433 VSS 0.093839f
C2455 DVSS.n2434 VSS 0.009721f
C2456 DVSS.n2435 VSS 0.062117f
C2457 DVSS.n2436 VSS 0.136758f
C2458 DVSS.n2437 VSS 0.019442f
C2459 DVSS.n2438 VSS 0.019442f
C2460 DVSS.n2439 VSS 0.019442f
C2461 DVSS.n2440 VSS 0.009721f
C2462 DVSS.n2441 VSS 0.142269f
C2463 DVSS.n2442 VSS 0.142269f
C2464 DVSS.n2443 VSS 0.142269f
C2465 DVSS.n2444 VSS 0.142269f
C2466 DVSS.n2445 VSS 0.142269f
C2467 DVSS.n2446 VSS 0.142269f
C2468 DVSS.n2447 VSS 0.142269f
C2469 DVSS.n2448 VSS 0.142269f
C2470 DVSS.n2449 VSS 0.142269f
C2471 DVSS.n2450 VSS 0.142269f
C2472 DVSS.n2451 VSS 0.142269f
C2473 DVSS.n2452 VSS 0.142269f
C2474 DVSS.n2453 VSS 0.142269f
C2475 DVSS.n2454 VSS 0.142269f
C2476 DVSS.n2455 VSS 2.21449f
C2477 DVSS.n2456 VSS 0.142269f
C2478 DVSS.n2457 VSS 0.062117f
C2479 DVSS.n2458 VSS 0.163454f
C2480 DVSS.n2459 VSS 0.019442f
C2481 DVSS.n2460 VSS 0.019442f
C2482 DVSS.n2461 VSS 0.019442f
C2483 DVSS.n2462 VSS 0.009721f
C2484 DVSS.n2463 VSS 0.462801f
C2485 DVSS.n2464 VSS 3.41655f
C2486 DVSS.n2465 VSS 0.010427f
C2487 DVSS.n2466 VSS 0.019442f
C2488 DVSS.n2467 VSS 0.019442f
C2489 DVSS.n2468 VSS 0.019442f
C2490 DVSS.n2469 VSS 0.009721f
C2491 DVSS.n2470 VSS 1.9679f
C2492 DVSS.n2471 VSS 0.021715f
C2493 DVSS.n2472 VSS 0.071134f
C2494 DVSS.n2473 VSS 0.114717f
C2495 DVSS.n2474 VSS 0.142269f
C2496 DVSS.n2475 VSS 0.142269f
C2497 DVSS.n2476 VSS 0.142269f
C2498 DVSS.n2477 VSS 0.142269f
C2499 DVSS.n2478 VSS 0.142269f
C2500 DVSS.n2479 VSS 0.142269f
C2501 DVSS.n2480 VSS 0.142269f
C2502 DVSS.n2481 VSS 0.142269f
C2503 DVSS.n2482 VSS 0.142269f
C2504 DVSS.n2483 VSS 0.142269f
C2505 DVSS.n2484 VSS 0.142269f
C2506 DVSS.n2485 VSS 0.142269f
C2507 DVSS.n2486 VSS 0.142269f
C2508 DVSS.n2487 VSS 0.142269f
C2509 DVSS.n2488 VSS 0.142269f
C2510 DVSS.n2489 VSS 0.142269f
C2511 DVSS.n2490 VSS 0.142269f
C2512 DVSS.n2491 VSS 0.142269f
C2513 DVSS.n2492 VSS 0.142269f
C2514 DVSS.n2493 VSS 0.142269f
C2515 DVSS.n2494 VSS 0.142269f
C2516 DVSS.n2495 VSS 0.142269f
C2517 DVSS.n2496 VSS 0.142269f
C2518 DVSS.n2497 VSS 0.142269f
C2519 DVSS.n2498 VSS 0.142269f
C2520 DVSS.n2499 VSS 0.142269f
C2521 DVSS.n2500 VSS 0.142269f
C2522 DVSS.n2501 VSS 0.142269f
C2523 DVSS.n2502 VSS 0.142269f
C2524 DVSS.n2503 VSS 0.142269f
C2525 DVSS.n2504 VSS 0.142269f
C2526 DVSS.n2505 VSS 0.142269f
C2527 DVSS.n2506 VSS 0.142269f
C2528 DVSS.n2507 VSS 0.142269f
C2529 DVSS.n2508 VSS 0.142269f
C2530 DVSS.n2509 VSS 0.142269f
C2531 DVSS.n2510 VSS 0.142269f
C2532 DVSS.n2511 VSS 0.142269f
C2533 DVSS.n2512 VSS 0.142269f
C2534 DVSS.n2513 VSS 0.142269f
C2535 DVSS.n2514 VSS 0.142269f
C2536 DVSS.n2515 VSS 0.142269f
C2537 DVSS.n2516 VSS 0.142269f
C2538 DVSS.n2517 VSS 0.142269f
C2539 DVSS.n2518 VSS 0.142269f
C2540 DVSS.n2519 VSS 0.142269f
C2541 DVSS.n2520 VSS 0.142269f
C2542 DVSS.n2521 VSS 0.142269f
C2543 DVSS.n2522 VSS 0.142269f
C2544 DVSS.n2523 VSS 0.142269f
C2545 DVSS.n2524 VSS 0.142269f
C2546 DVSS.n2525 VSS 0.071134f
C2547 DVSS.n2526 VSS 0.142269f
C2548 DVSS.n2527 VSS 0.142269f
C2549 DVSS.n2528 VSS 0.142269f
C2550 DVSS.n2529 VSS 0.142269f
C2551 DVSS.n2531 VSS 0.052105f
C2552 DVSS.n2532 VSS 0.052105f
C2553 DVSS.n2533 VSS 0.052105f
C2554 DVSS.n2534 VSS 0.438058f
C2555 DVSS.n2536 VSS 0.052105f
C2556 DVSS.n2538 VSS 0.052105f
C2557 DVSS.n2540 VSS 0.052105f
C2558 DVSS.n2546 VSS 0.065624f
C2559 DVSS.n2547 VSS 0.062117f
C2560 DVSS.n2548 VSS 0.142269f
C2561 DVSS.n2549 VSS 0.142269f
C2562 DVSS.n2550 VSS 0.142269f
C2563 DVSS.n2551 VSS 0.142269f
C2564 DVSS.n2552 VSS 0.142269f
C2565 DVSS.n2553 VSS 0.142269f
C2566 DVSS.n2554 VSS 0.142269f
C2567 DVSS.n2555 VSS 0.142269f
C2568 DVSS.n2556 VSS 0.142269f
C2569 DVSS.n2557 VSS 0.142269f
C2570 DVSS.n2558 VSS 0.142269f
C2571 DVSS.n2559 VSS 0.142269f
C2572 DVSS.n2560 VSS 0.142269f
C2573 DVSS.n2561 VSS 0.142269f
C2574 DVSS.n2562 VSS 0.142269f
C2575 DVSS.n2563 VSS 0.142269f
C2576 DVSS.n2564 VSS 0.142269f
C2577 DVSS.n2565 VSS 0.142269f
C2578 DVSS.n2566 VSS 0.142269f
C2579 DVSS.n2567 VSS 0.142269f
C2580 DVSS.n2568 VSS 0.142269f
C2581 DVSS.n2569 VSS 0.142269f
C2582 DVSS.n2570 VSS 0.142269f
C2583 DVSS.n2571 VSS 0.142269f
C2584 DVSS.n2572 VSS 0.142269f
C2585 DVSS.n2573 VSS 0.142269f
C2586 DVSS.n2574 VSS 0.142269f
C2587 DVSS.n2575 VSS 0.142269f
C2588 DVSS.n2576 VSS 0.142269f
C2589 DVSS.n2577 VSS 0.142269f
C2590 DVSS.n2578 VSS 0.142269f
C2591 DVSS.n2579 VSS 0.142269f
C2592 DVSS.n2580 VSS 0.142269f
C2593 DVSS.n2581 VSS 0.142269f
C2594 DVSS.n2582 VSS 0.142269f
C2595 DVSS.n2583 VSS 0.142269f
C2596 DVSS.n2584 VSS 0.142269f
C2597 DVSS.n2585 VSS 0.142269f
C2598 DVSS.n2586 VSS 0.142269f
C2599 DVSS.n2587 VSS 0.142269f
C2600 DVSS.n2588 VSS 0.142269f
C2601 DVSS.n2589 VSS 0.142269f
C2602 DVSS.n2590 VSS 0.142269f
C2603 DVSS.n2591 VSS 0.142269f
C2604 DVSS.n2592 VSS 0.142269f
C2605 DVSS.n2593 VSS 0.116721f
C2606 DVSS.n2594 VSS 0.142269f
C2607 DVSS.n2595 VSS 0.142269f
C2608 DVSS.n2596 VSS 0.142269f
C2609 DVSS.n2597 VSS 0.142269f
C2610 DVSS.n2598 VSS 0.142269f
C2611 DVSS.n2599 VSS 0.071134f
C2612 DVSS.n2600 VSS 0.010427f
C2613 DVSS.n2601 VSS 0.009721f
C2614 DVSS.n2602 VSS 0.019442f
C2615 DVSS.n2603 VSS 0.019442f
C2616 DVSS.n2604 VSS 0.019442f
C2617 DVSS.n2605 VSS 0.019442f
C2618 DVSS.n2606 VSS 0.019442f
C2619 DVSS.n2607 VSS 0.019442f
C2620 DVSS.n2608 VSS 0.009721f
C2621 DVSS.n2609 VSS 0.068047f
C2622 DVSS.n2610 VSS 0.013014f
C2623 DVSS.n2611 VSS 0.11579f
C2624 DVSS.n2612 VSS 0.009721f
C2625 DVSS.n2613 VSS 0.009721f
C2626 DVSS.n2614 VSS 0.008467f
C2627 DVSS.n2615 VSS 0.019442f
C2628 DVSS.n2616 VSS 0.15585f
C2629 DVSS.n2617 VSS 0.15585f
C2630 DVSS.n2618 VSS 0.15585f
C2631 DVSS.n2619 VSS 0.15585f
C2632 DVSS.n2620 VSS 0.15585f
C2633 DVSS.n2621 VSS 0.15585f
C2634 DVSS.n2622 VSS 0.15585f
C2635 DVSS.n2623 VSS 0.15585f
C2636 DVSS.n2624 VSS 0.15585f
C2637 DVSS.n2625 VSS 0.15585f
C2638 DVSS.n2626 VSS 0.15585f
C2639 DVSS.n2627 VSS 0.15585f
C2640 DVSS.n2628 VSS 0.15585f
C2641 DVSS.n2629 VSS 0.15585f
C2642 DVSS.n2630 VSS 0.15585f
C2643 DVSS.n2631 VSS 0.15585f
C2644 DVSS.n2632 VSS 0.15585f
C2645 DVSS.n2633 VSS 0.15585f
C2646 DVSS.n2634 VSS 0.15585f
C2647 DVSS.n2635 VSS 0.15585f
C2648 DVSS.n2636 VSS 0.15585f
C2649 DVSS.n2637 VSS 0.15585f
C2650 DVSS.n2638 VSS 0.15585f
C2651 DVSS.n2639 VSS 0.15585f
C2652 DVSS.n2640 VSS 0.15585f
C2653 DVSS.n2641 VSS 0.15585f
C2654 DVSS.n2642 VSS 0.15585f
C2655 DVSS.n2643 VSS 0.15585f
C2656 DVSS.n2644 VSS 0.15585f
C2657 DVSS.n2645 VSS 0.15585f
C2658 DVSS.n2646 VSS 0.15585f
C2659 DVSS.n2647 VSS 0.077925f
C2660 DVSS.n2648 VSS 0.15585f
C2661 DVSS.n2649 VSS 0.15585f
C2662 DVSS.n2650 VSS 0.15585f
C2663 DVSS.n2651 VSS 0.15585f
C2664 DVSS.n2652 VSS 0.15585f
C2665 DVSS.n2653 VSS 0.15585f
C2666 DVSS.n2654 VSS 0.15585f
C2667 DVSS.n2655 VSS 0.15585f
C2668 DVSS.n2656 VSS 0.15585f
C2669 DVSS.n2657 VSS 0.15585f
C2670 DVSS.n2658 VSS 0.15585f
C2671 DVSS.n2659 VSS 0.15585f
C2672 DVSS.n2660 VSS 0.15585f
C2673 DVSS.n2661 VSS 0.15585f
C2674 DVSS.n2662 VSS 0.15585f
C2675 DVSS.n2663 VSS 0.15585f
C2676 DVSS.n2664 VSS 0.15585f
C2677 DVSS.n2665 VSS 0.15585f
C2678 DVSS.n2666 VSS 0.15585f
C2679 DVSS.n2667 VSS 0.15585f
C2680 DVSS.n2668 VSS 0.15585f
C2681 DVSS.n2669 VSS 0.15585f
C2682 DVSS.n2670 VSS 0.15585f
C2683 DVSS.n2671 VSS 0.15585f
C2684 DVSS.n2672 VSS 0.15585f
C2685 DVSS.n2673 VSS 0.15585f
C2686 DVSS.n2674 VSS 0.15585f
C2687 DVSS.n2675 VSS 0.15585f
C2688 DVSS.n2676 VSS 0.15585f
C2689 DVSS.n2677 VSS 0.15585f
C2690 DVSS.n2678 VSS 0.15585f
C2691 DVSS.n2679 VSS 2.43723f
C2692 DVSS.n2680 VSS 0.506941f
C2693 DVSS.n2681 VSS 0.15585f
C2694 DVSS.n2682 VSS 0.15585f
C2695 DVSS.n2683 VSS 0.15585f
C2696 DVSS.n2684 VSS 0.15585f
C2697 DVSS.n2685 VSS 0.15585f
C2698 DVSS.n2686 VSS 0.15585f
C2699 DVSS.n2687 VSS 0.15585f
C2700 DVSS.n2688 VSS 0.15585f
C2701 DVSS.n2689 VSS 0.15585f
C2702 DVSS.n2690 VSS 0.15585f
C2703 DVSS.n2691 VSS 0.15585f
C2704 DVSS.n2692 VSS 0.15585f
C2705 DVSS.n2693 VSS 0.15585f
C2706 DVSS.n2694 VSS 0.15585f
C2707 DVSS.n2695 VSS 0.15585f
C2708 DVSS.n2696 VSS 0.15585f
C2709 DVSS.n2697 VSS 0.15585f
C2710 DVSS.n2698 VSS 0.15585f
C2711 DVSS.n2699 VSS 0.15585f
C2712 DVSS.n2700 VSS 0.15585f
C2713 DVSS.n2701 VSS 0.15585f
C2714 DVSS.n2702 VSS 0.15585f
C2715 DVSS.n2703 VSS 0.15585f
C2716 DVSS.n2704 VSS 0.15585f
C2717 DVSS.n2705 VSS 0.15585f
C2718 DVSS.n2706 VSS 0.15585f
C2719 DVSS.n2707 VSS 0.15585f
C2720 DVSS.n2708 VSS 0.15585f
C2721 DVSS.n2709 VSS 0.15585f
C2722 DVSS.n2710 VSS 0.15585f
C2723 DVSS.n2711 VSS 0.15585f
C2724 DVSS.n2712 VSS 0.15585f
C2725 DVSS.n2713 VSS 0.15585f
C2726 DVSS.n2714 VSS 0.15585f
C2727 DVSS.n2715 VSS 0.15585f
C2728 DVSS.n2716 VSS 0.15585f
C2729 DVSS.n2717 VSS 0.15585f
C2730 DVSS.n2718 VSS 0.15585f
C2731 DVSS.n2719 VSS 0.15585f
C2732 DVSS.n2720 VSS 0.15585f
C2733 DVSS.n2721 VSS 0.15585f
C2734 DVSS.n2722 VSS 0.15585f
C2735 DVSS.n2723 VSS 0.15585f
C2736 DVSS.n2724 VSS 0.15585f
C2737 DVSS.n2725 VSS 0.15585f
C2738 DVSS.n2726 VSS 0.15585f
C2739 DVSS.n2727 VSS 0.15585f
C2740 DVSS.n2728 VSS 0.15585f
C2741 DVSS.n2729 VSS 0.15585f
C2742 DVSS.n2730 VSS 0.15585f
C2743 DVSS.n2731 VSS 0.15585f
C2744 DVSS.n2732 VSS 0.15585f
C2745 DVSS.n2733 VSS 0.15585f
C2746 DVSS.n2734 VSS 0.15585f
C2747 DVSS.n2735 VSS 0.15585f
C2748 DVSS.n2736 VSS 0.15585f
C2749 DVSS.n2737 VSS 0.15585f
C2750 DVSS.n2738 VSS 0.15585f
C2751 DVSS.n2739 VSS 0.15585f
C2752 DVSS.n2740 VSS 0.15585f
C2753 DVSS.n2741 VSS 0.15585f
C2754 DVSS.n2742 VSS 0.15585f
C2755 DVSS.n2743 VSS 0.15585f
C2756 DVSS.n2744 VSS 0.093839f
C2757 DVSS.n2745 VSS 0.077925f
C2758 DVSS.n2746 VSS 0.022691f
C2759 DVSS.n2747 VSS 0.438058f
C2760 DVSS.n2748 VSS 0.052105f
C2761 DVSS.n2749 VSS 0.052105f
C2762 DVSS.n2751 VSS 0.052105f
C2763 DVSS.n2752 VSS 0.212831f
C2764 DVSS.n2755 VSS 0.052105f
C2765 DVSS.n2757 VSS 0.052105f
C2766 DVSS.n2761 VSS 0.068047f
C2767 DVSS.n2763 VSS 0.071889f
C2768 DVSS.n2764 VSS 0.034877f
C2769 DVSS.n2765 VSS 0.074084f
C2770 DVSS.n2766 VSS 0.068047f
C2771 DVSS.n2767 VSS 0.15585f
C2772 DVSS.n2768 VSS 0.15585f
C2773 DVSS.n2769 VSS 0.15585f
C2774 DVSS.n2770 VSS 0.15585f
C2775 DVSS.n2771 VSS 0.15585f
C2776 DVSS.n2772 VSS 0.091644f
C2777 DVSS.n2773 VSS 0.15585f
C2778 DVSS.n2774 VSS 0.15585f
C2779 DVSS.n2775 VSS 0.15585f
C2780 DVSS.n2776 VSS 0.15585f
C2781 DVSS.n2777 VSS 0.15585f
C2782 DVSS.n2778 VSS 0.15585f
C2783 DVSS.n2779 VSS 0.15585f
C2784 DVSS.n2780 VSS 0.15585f
C2785 DVSS.n2781 VSS 0.15585f
C2786 DVSS.n2782 VSS 0.15585f
C2787 DVSS.n2783 VSS 0.15585f
C2788 DVSS.n2784 VSS 0.15585f
C2789 DVSS.n2785 VSS 0.15585f
C2790 DVSS.n2786 VSS 0.15585f
C2791 DVSS.n2787 VSS 0.15585f
C2792 DVSS.n2788 VSS 0.15585f
C2793 DVSS.n2789 VSS 0.15585f
C2794 DVSS.n2790 VSS 0.15585f
C2795 DVSS.n2791 VSS 0.15585f
C2796 DVSS.n2792 VSS 0.15585f
C2797 DVSS.n2793 VSS 0.15585f
C2798 DVSS.n2794 VSS 0.15585f
C2799 DVSS.n2795 VSS 0.15585f
C2800 DVSS.n2796 VSS 0.15585f
C2801 DVSS.n2797 VSS 0.15585f
C2802 DVSS.n2798 VSS 0.152009f
C2803 DVSS.n2799 VSS 0.15585f
C2804 DVSS.n2800 VSS 0.15585f
C2805 DVSS.n2801 VSS 0.15585f
C2806 DVSS.n2802 VSS 0.15585f
C2807 DVSS.n2803 VSS 0.15585f
C2808 DVSS.n2804 VSS 0.15585f
C2809 DVSS.n2805 VSS 0.15585f
C2810 DVSS.n2806 VSS 0.15585f
C2811 DVSS.n2807 VSS 0.15585f
C2812 DVSS.n2808 VSS 0.15585f
C2813 DVSS.n2809 VSS 0.15585f
C2814 DVSS.n2810 VSS 0.15585f
C2815 DVSS.n2811 VSS 0.15585f
C2816 DVSS.n2812 VSS 0.15585f
C2817 DVSS.n2813 VSS 0.15585f
C2818 DVSS.n2814 VSS 0.15585f
C2819 DVSS.n2815 VSS 0.15585f
C2820 DVSS.n2816 VSS 0.15585f
C2821 DVSS.n2817 VSS 0.15585f
C2822 DVSS.n2818 VSS 0.15585f
C2823 DVSS.n2819 VSS 0.15585f
C2824 DVSS.n2820 VSS 0.15585f
C2825 DVSS.n2821 VSS 0.15585f
C2826 DVSS.n2822 VSS 0.15585f
C2827 DVSS.n2823 VSS 0.15585f
C2828 DVSS.n2824 VSS 0.15585f
C2829 DVSS.n2825 VSS 0.15585f
C2830 DVSS.n2826 VSS 0.15585f
C2831 DVSS.n2827 VSS 0.15585f
C2832 DVSS.n2828 VSS 0.15585f
C2833 DVSS.n2829 VSS 0.15585f
C2834 DVSS.n2830 VSS 0.15585f
C2835 DVSS.n2831 VSS 0.15585f
C2836 DVSS.n2832 VSS 0.15585f
C2837 DVSS.n2833 VSS 0.15585f
C2838 DVSS.n2834 VSS 0.15585f
C2839 DVSS.n2835 VSS 0.15585f
C2840 DVSS.n2836 VSS 0.15585f
C2841 DVSS.n2837 VSS 0.15585f
C2842 DVSS.n2838 VSS 0.15585f
C2843 DVSS.n2839 VSS 0.15585f
C2844 DVSS.n2840 VSS 0.15585f
C2845 DVSS.n2841 VSS 0.15585f
C2846 DVSS.n2842 VSS 0.15585f
C2847 DVSS.n2843 VSS 0.15585f
C2848 DVSS.n2844 VSS 0.15585f
C2849 DVSS.n2845 VSS 0.751144f
C2850 DVSS.n2846 VSS 0.205146f
C2851 DVSS.n2847 VSS 0.08012f
C2852 DVSS.n2848 VSS 0.15585f
C2853 DVSS.n2849 VSS 0.140485f
C2854 DVSS.n2850 VSS 0.140485f
C2855 DVSS.n2851 VSS 0.15585f
C2856 DVSS.n2852 VSS 0.15585f
C2857 DVSS.n2853 VSS 0.15585f
C2858 DVSS.n2854 VSS 0.15585f
C2859 DVSS.n2855 VSS 0.15585f
C2860 DVSS.n2856 VSS 0.15585f
C2861 DVSS.n2857 VSS 0.15585f
C2862 DVSS.n2858 VSS 0.15585f
C2863 DVSS.n2859 VSS 0.15585f
C2864 DVSS.n2860 VSS 0.15585f
C2865 DVSS.n2861 VSS 0.15585f
C2866 DVSS.n2862 VSS 0.15585f
C2867 DVSS.n2863 VSS 0.15585f
C2868 DVSS.n2864 VSS 0.15585f
C2869 DVSS.n2865 VSS 0.15585f
C2870 DVSS.n2866 VSS 0.15585f
C2871 DVSS.n2867 VSS 0.15585f
C2872 DVSS.n2868 VSS 0.15585f
C2873 DVSS.n2869 VSS 0.15585f
C2874 DVSS.n2870 VSS 0.15585f
C2875 DVSS.n2871 VSS 0.15585f
C2876 DVSS.n2872 VSS 0.15585f
C2877 DVSS.n2873 VSS 0.15585f
C2878 DVSS.n2874 VSS 0.15585f
C2879 DVSS.n2875 VSS 0.127863f
C2880 DVSS.n2876 VSS 0.009721f
C2881 DVSS.n2877 VSS 0.009721f
C2882 DVSS.n2878 VSS 0.288809f
C2883 DVSS.n2879 VSS 0.288809f
C2884 DVSS.n2880 VSS 0.077925f
C2885 DVSS.n2881 VSS 0.019442f
C2886 DVSS.n2882 VSS 0.019442f
C2887 DVSS.n2883 VSS 0.077925f
C2888 DVSS.n2884 VSS 0.163454f
C2889 DVSS.n2885 VSS 0.163454f
C2890 DVSS.n2886 VSS 0.009721f
C2891 DVSS.n2887 VSS 0.142269f
C2892 DVSS.n2888 VSS 0.142269f
C2893 DVSS.n2889 VSS 0.142269f
C2894 DVSS.n2890 VSS 0.142269f
C2895 DVSS.n2891 VSS 0.142269f
C2896 DVSS.n2892 VSS 0.142269f
C2897 DVSS.n2893 VSS 0.142269f
C2898 DVSS.n2894 VSS 0.142269f
C2899 DVSS.n2895 VSS 0.142269f
C2900 DVSS.n2896 VSS 0.142269f
C2901 DVSS.n2897 VSS 0.142269f
C2902 DVSS.n2898 VSS 0.142269f
C2903 DVSS.n2899 VSS 0.142269f
C2904 DVSS.n2900 VSS 0.142269f
C2905 DVSS.n2901 VSS 0.142269f
C2906 DVSS.n2902 VSS 0.142269f
C2907 DVSS.n2903 VSS 0.142269f
C2908 DVSS.n2904 VSS 0.073138f
C2909 DVSS.n2905 VSS 0.186193f
C2910 DVSS.n2906 VSS 0.686742f
C2911 DVSS.n2907 VSS 0.128242f
C2912 DVSS.n2908 VSS 0.128242f
C2913 DVSS.n2909 VSS 0.142269f
C2914 DVSS.n2910 VSS 0.142269f
C2915 DVSS.n2911 VSS 0.142269f
C2916 DVSS.n2912 VSS 0.142269f
C2917 DVSS.n2913 VSS 0.142269f
C2918 DVSS.n2914 VSS 0.142269f
C2919 DVSS.n2915 VSS 0.142269f
C2920 DVSS.n2916 VSS 0.142269f
C2921 DVSS.n2917 VSS 0.142269f
C2922 DVSS.n2918 VSS 0.142269f
C2923 DVSS.n2919 VSS 0.142269f
C2924 DVSS.n2920 VSS 0.142269f
C2925 DVSS.n2921 VSS 0.142269f
C2926 DVSS.n2922 VSS 0.142269f
C2927 DVSS.n2923 VSS 0.142269f
C2928 DVSS.n2924 VSS 0.1057f
C2929 DVSS.n2925 VSS 0.009721f
C2930 DVSS.n2926 VSS 0.021715f
C2931 DVSS.n2927 VSS 0.071134f
C2932 DVSS.n2928 VSS 0.062117f
C2933 DVSS.n2929 VSS 0.142269f
C2934 DVSS.n2930 VSS 0.142269f
C2935 DVSS.n2931 VSS 0.142269f
C2936 DVSS.n2932 VSS 0.142269f
C2937 DVSS.n2933 VSS 0.142269f
C2938 DVSS.n2934 VSS 0.142269f
C2939 DVSS.n2935 VSS 0.142269f
C2940 DVSS.n2936 VSS 0.142269f
C2941 DVSS.n2937 VSS 0.142269f
C2942 DVSS.n2938 VSS 0.142269f
C2943 DVSS.n2939 VSS 0.142269f
C2944 DVSS.n2940 VSS 0.142269f
C2945 DVSS.n2941 VSS 0.142269f
C2946 DVSS.n2942 VSS 0.142269f
C2947 DVSS.n2943 VSS 0.142269f
C2948 DVSS.n2944 VSS 0.142269f
C2949 DVSS.n2945 VSS 0.142269f
C2950 DVSS.n2946 VSS 0.142269f
C2951 DVSS.n2947 VSS 0.142269f
C2952 DVSS.n2948 VSS 0.142269f
C2953 DVSS.n2949 VSS 0.142269f
C2954 DVSS.n2950 VSS 0.142269f
C2955 DVSS.n2951 VSS 0.142269f
C2956 DVSS.n2952 VSS 0.083658f
C2957 DVSS.n2953 VSS 0.142269f
C2958 DVSS.n2954 VSS 0.062117f
C2959 DVSS.n2955 VSS 0.142269f
C2960 DVSS.n2956 VSS 0.142269f
C2961 DVSS.n2957 VSS 0.138762f
C2962 DVSS.n2958 VSS 0.142269f
C2963 DVSS.n2959 VSS 0.142269f
C2964 DVSS.n2960 VSS 0.142269f
C2965 DVSS.n2961 VSS 0.142269f
C2966 DVSS.n2962 VSS 0.142269f
C2967 DVSS.n2963 VSS 0.142269f
C2968 DVSS.n2964 VSS 0.142269f
C2969 DVSS.n2965 VSS 0.142269f
C2970 DVSS.n2966 VSS 0.142269f
C2971 DVSS.n2967 VSS 0.142269f
C2972 DVSS.n2968 VSS 0.142269f
C2973 DVSS.n2969 VSS 0.142269f
C2974 DVSS.n2970 VSS 0.142269f
C2975 DVSS.n2971 VSS 0.142269f
C2976 DVSS.n2972 VSS 0.142269f
C2977 DVSS.n2973 VSS 0.142269f
C2978 DVSS.n2974 VSS 0.142269f
C2979 DVSS.n2975 VSS 0.142269f
C2980 DVSS.n2976 VSS 0.142269f
C2981 DVSS.n2977 VSS 0.142269f
C2982 DVSS.n2978 VSS 0.142269f
C2983 DVSS.n2979 VSS 0.142269f
C2984 DVSS.n2980 VSS 0.083658f
C2985 DVSS.n2981 VSS 0.071134f
C2986 DVSS.n2982 VSS 0.052105f
C2987 DVSS.n2983 VSS 0.067628f
C2988 DVSS.n2984 VSS 0.062117f
C2989 DVSS.n2985 VSS 0.142269f
C2990 DVSS.n2986 VSS 0.142269f
C2991 DVSS.n2987 VSS 0.085662f
C2992 DVSS.n2988 VSS 0.142269f
C2993 DVSS.n2989 VSS 0.142269f
C2994 DVSS.n2990 VSS 0.142269f
C2995 DVSS.n2991 VSS 0.142269f
C2996 DVSS.n2992 VSS 0.142269f
C2997 DVSS.n2993 VSS 0.142269f
C2998 DVSS.n2994 VSS 0.142269f
C2999 DVSS.n2995 VSS 0.142269f
C3000 DVSS.n2996 VSS 0.142269f
C3001 DVSS.n2997 VSS 0.142269f
C3002 DVSS.n2998 VSS 0.142269f
C3003 DVSS.n2999 VSS 0.142269f
C3004 DVSS.n3000 VSS 0.142269f
C3005 DVSS.n3001 VSS 0.142269f
C3006 DVSS.n3002 VSS 0.142269f
C3007 DVSS.n3003 VSS 0.142269f
C3008 DVSS.n3004 VSS 0.142269f
C3009 DVSS.n3005 VSS 0.142269f
C3010 DVSS.n3006 VSS 0.142269f
C3011 DVSS.n3007 VSS 0.142269f
C3012 DVSS.n3008 VSS 0.142269f
C3013 DVSS.n3009 VSS 0.142269f
C3014 DVSS.n3010 VSS 0.142269f
C3015 DVSS.n3011 VSS 0.142269f
C3016 DVSS.n3012 VSS 0.085662f
C3017 DVSS.n3013 VSS 0.010427f
C3018 DVSS.n3014 VSS 0.019442f
C3019 DVSS.n3015 VSS 0.019442f
C3020 DVSS.n3016 VSS 0.019442f
C3021 DVSS.n3017 VSS 0.071134f
C3022 DVSS.n3018 VSS 0.021715f
C3023 DVSS.n3019 VSS 0.071134f
C3024 DVSS.n3020 VSS 0.163454f
C3025 DVSS.n3021 VSS 0.163454f
C3026 DVSS.n3022 VSS 0.019442f
C3027 DVSS.n3023 VSS 0.077925f
C3028 DVSS.n3024 VSS 0.019442f
C3029 DVSS.n3025 VSS 0.009721f
C3030 DVSS.n3026 VSS 0.077925f
C3031 DVSS.n3027 VSS 0.079415f
C3032 DVSS.n3028 VSS 0.079415f
C3033 DVSS.n3030 VSS 0.062324f
C3034 DVSS.n3031 VSS 0.062324f
C3035 DVSS.n3032 VSS 0.210064f
C3036 DVSS.n3034 VSS 0.210064f
C3037 DVSS.n3035 VSS 0.167029f
C3038 DVSS.n3036 VSS 0.210064f
C3039 DVSS.n3037 VSS 0.210064f
C3040 DVSS.n3039 VSS 0.062324f
C3041 DVSS.n3040 VSS 0.079415f
C3042 DVSS.n3041 VSS 0.079415f
C3043 DVSS.n3042 VSS 0.009721f
C3044 DVSS.n3043 VSS 0.008467f
C3045 DVSS.n3044 VSS 0.077925f
C3046 DVSS.n3045 VSS 0.013014f
C3047 DVSS.n3046 VSS 0.009721f
C3048 DVSS.n3047 VSS 0.019442f
C3049 DVSS.n3048 VSS 0.019442f
C3050 DVSS.n3049 VSS 0.019442f
C3051 DVSS.n3050 VSS 0.009721f
C3052 DVSS.n3051 VSS 0.163454f
C3053 DVSS.n3052 VSS 0.163454f
C3054 DVSS.n3053 VSS 0.009721f
C3055 DVSS.n3054 VSS 0.019442f
C3056 DVSS.n3055 VSS 0.019442f
C3057 DVSS.n3056 VSS 0.019442f
C3058 DVSS.n3057 VSS 0.019442f
C3059 DVSS.n3058 VSS 0.019442f
C3060 DVSS.n3059 VSS 0.019442f
C3061 DVSS.n3060 VSS 0.009721f
C3062 DVSS.n3061 VSS 0.010427f
C3063 DVSS.n3062 VSS 0.009721f
C3064 DVSS.n3063 VSS 0.127656f
C3065 DVSS.n3064 VSS 0.068207f
C3066 DVSS.n3065 VSS 0.026052f
C3067 DVSS.n3066 VSS 0.066898f
C3068 DVSS.n3067 VSS 0.128978f
C3069 DVSS.n3068 VSS 0.160836f
C3070 DVSS.t28 VSS 0.311996f
C3071 DVSS.n3069 VSS 3.60328f
C3072 DVSS.n3070 VSS 12.026401f
C3073 DVSS.n3071 VSS 16.075998f
C3074 DVSS.n3072 VSS 0.249533f
C3075 DVSS.n3073 VSS 0.648801f
C3076 DVSS.n3074 VSS 0.006371f
C3077 DVSS.n3075 VSS 0.009203f
C3078 DVSS.n3076 VSS 0.016297f
C3079 DVSS.n3077 VSS 0.016098f
C3080 DVSS.n3078 VSS 0.184013f
C3081 DVSS.n3079 VSS 0.070738f
C3082 DVSS.n3080 VSS 0.24979f
C3083 DVSS.n3081 VSS 0.648801f
C3084 DVSS.n3082 VSS 2.0355f
C3085 DVSS.n3083 VSS 1.03491f
C3086 DVSS.n3084 VSS 0.755683f
C3087 DVSS.n3085 VSS 1.70064f
C3088 DVSS.n3086 VSS 0.869181f
C3089 DVSS.n3087 VSS 5.82075f
C3090 DVSS.n3088 VSS 10.5057f
C3091 DVSS.n3089 VSS -5.09135f
C3092 DVSS.n3090 VSS 0.919657f
C3093 DVSS.n3091 VSS 0.919657f
C3094 DVSS.n3092 VSS 0.635473f
C3095 DVSS.n3093 VSS 0.183837f
C3096 DVSS.n3094 VSS 0.037283f
C3097 DVSS.n3095 VSS 0.027376f
C3098 DVSS.n3096 VSS 0.281067f
C3099 DVSS.n3097 VSS 0.15585f
C3100 DVSS.n3098 VSS 0.15585f
C3101 DVSS.n3099 VSS 0.15585f
C3102 DVSS.n3100 VSS 0.577503f
C3103 DVSS.n3101 VSS 0.15585f
C3104 DVSS.n3102 VSS 0.15585f
C3105 DVSS.n3103 VSS 0.15585f
C3106 DVSS.n3104 VSS 0.15585f
C3107 DVSS.n3105 VSS 0.15585f
C3108 DVSS.n3106 VSS 0.15585f
C3109 DVSS.n3107 VSS 0.15585f
C3110 DVSS.n3108 VSS 0.15585f
C3111 DVSS.n3109 VSS 0.15585f
C3112 DVSS.n3110 VSS 0.15585f
C3113 DVSS.n3111 VSS 0.15585f
C3114 DVSS.n3112 VSS 0.15585f
C3115 DVSS.n3113 VSS 0.15585f
C3116 DVSS.n3114 VSS 0.15585f
C3117 DVSS.n3115 VSS 0.15585f
C3118 DVSS.n3116 VSS 0.15585f
C3119 DVSS.n3117 VSS 0.15585f
C3120 DVSS.n3118 VSS 0.15585f
C3121 DVSS.n3119 VSS 0.15585f
C3122 DVSS.n3120 VSS 0.15585f
C3123 DVSS.n3121 VSS 0.15585f
C3124 DVSS.n3122 VSS 0.15585f
C3125 DVSS.n3123 VSS 0.15585f
C3126 DVSS.n3124 VSS 0.15585f
C3127 DVSS.n3125 VSS 0.15585f
C3128 DVSS.n3126 VSS 0.15585f
C3129 DVSS.n3127 VSS 0.15585f
C3130 DVSS.n3128 VSS 0.15585f
C3131 DVSS.n3129 VSS 0.15585f
C3132 DVSS.n3130 VSS 0.15585f
C3133 DVSS.n3131 VSS 0.15585f
C3134 DVSS.n3132 VSS 0.15585f
C3135 DVSS.n3133 VSS 0.15585f
C3136 DVSS.n3134 VSS 0.15585f
C3137 DVSS.n3135 VSS 0.15585f
C3138 DVSS.n3136 VSS 0.15585f
C3139 DVSS.n3137 VSS 0.15585f
C3140 DVSS.n3138 VSS 0.15585f
C3141 DVSS.n3139 VSS 0.15585f
C3142 DVSS.n3140 VSS 0.15585f
C3143 DVSS.n3141 VSS 0.15585f
C3144 DVSS.n3142 VSS 0.15585f
C3145 DVSS.n3143 VSS 0.15585f
C3146 DVSS.n3144 VSS 0.15585f
C3147 DVSS.n3145 VSS 0.15585f
C3148 DVSS.n3146 VSS 0.15585f
C3149 DVSS.n3147 VSS 0.15585f
C3150 DVSS.n3148 VSS 0.15585f
C3151 DVSS.n3149 VSS 0.15585f
C3152 DVSS.n3150 VSS 0.15585f
C3153 DVSS.n3151 VSS 0.15585f
C3154 DVSS.n3152 VSS 0.15585f
C3155 DVSS.n3153 VSS 0.15585f
C3156 DVSS.n3154 VSS 0.15585f
C3157 DVSS.n3155 VSS 0.15585f
C3158 DVSS.n3156 VSS 0.15585f
C3159 DVSS.n3157 VSS 0.15585f
C3160 DVSS.n3158 VSS 0.15585f
C3161 DVSS.n3159 VSS 0.15585f
C3162 DVSS.n3160 VSS 0.15585f
C3163 DVSS.n3161 VSS 0.15585f
C3164 DVSS.n3162 VSS 0.15585f
C3165 DVSS.n3163 VSS 0.15585f
C3166 DVSS.n3164 VSS 0.15585f
C3167 DVSS.n3165 VSS 0.15585f
C3168 DVSS.n3166 VSS 0.15585f
C3169 DVSS.n3167 VSS 0.15585f
C3170 DVSS.n3168 VSS 0.15585f
C3171 DVSS.n3169 VSS 0.15585f
C3172 DVSS.n3170 VSS 0.15585f
C3173 DVSS.n3171 VSS 0.15585f
C3174 DVSS.n3172 VSS 0.15585f
C3175 DVSS.n3173 VSS 0.15585f
C3176 DVSS.n3174 VSS 0.15585f
C3177 DVSS.n3175 VSS 0.15585f
C3178 DVSS.n3176 VSS 0.15585f
C3179 DVSS.n3177 VSS 0.15585f
C3180 DVSS.n3178 VSS 0.15585f
C3181 DVSS.n3179 VSS 0.15585f
C3182 DVSS.n3180 VSS 0.15585f
C3183 DVSS.n3181 VSS 0.15585f
C3184 DVSS.n3182 VSS 0.15585f
C3185 DVSS.n3183 VSS 0.15585f
C3186 DVSS.n3184 VSS 0.15585f
C3187 DVSS.n3185 VSS 0.15585f
C3188 DVSS.n3186 VSS 0.15585f
C3189 DVSS.n3187 VSS 0.15585f
C3190 DVSS.n3188 VSS 0.15585f
C3191 DVSS.n3189 VSS 0.15585f
C3192 DVSS.n3190 VSS 0.15585f
C3193 DVSS.n3191 VSS 0.15585f
C3194 DVSS.n3192 VSS 0.15585f
C3195 DVSS.n3193 VSS 0.15585f
C3196 DVSS.n3194 VSS 0.15585f
C3197 DVSS.n3195 VSS 0.15585f
C3198 DVSS.n3196 VSS 0.15585f
C3199 DVSS.n3197 VSS 0.15585f
C3200 DVSS.n3198 VSS 0.15585f
C3201 DVSS.n3199 VSS 0.15585f
C3202 DVSS.n3200 VSS 0.15585f
C3203 DVSS.n3201 VSS 0.15585f
C3204 DVSS.n3202 VSS 0.15585f
C3205 DVSS.n3203 VSS 0.15585f
C3206 DVSS.n3204 VSS 0.15585f
C3207 DVSS.n3205 VSS 0.15585f
C3208 DVSS.n3206 VSS 0.15585f
C3209 DVSS.n3207 VSS 0.15585f
C3210 DVSS.n3208 VSS 0.15585f
C3211 DVSS.n3209 VSS 0.15585f
C3212 DVSS.n3210 VSS 0.15585f
C3213 DVSS.n3211 VSS 0.15585f
C3214 DVSS.n3212 VSS 0.15585f
C3215 DVSS.n3213 VSS 0.15585f
C3216 DVSS.n3214 VSS 0.15585f
C3217 DVSS.n3215 VSS 0.15585f
C3218 DVSS.n3216 VSS 0.15585f
C3219 DVSS.n3217 VSS 0.15585f
C3220 DVSS.n3218 VSS 0.15585f
C3221 DVSS.n3219 VSS 0.15585f
C3222 DVSS.n3220 VSS 0.15585f
C3223 DVSS.n3221 VSS 0.15585f
C3224 DVSS.n3222 VSS 0.15585f
C3225 DVSS.n3223 VSS 0.15585f
C3226 DVSS.n3224 VSS 0.15585f
C3227 DVSS.n3225 VSS 0.15585f
C3228 DVSS.n3226 VSS 0.15585f
C3229 DVSS.n3227 VSS 0.15585f
C3230 DVSS.n3228 VSS 0.15585f
C3231 DVSS.n3229 VSS 0.15585f
C3232 DVSS.n3230 VSS 0.15585f
C3233 DVSS.n3231 VSS 0.15585f
C3234 DVSS.n3232 VSS 0.15585f
C3235 DVSS.n3233 VSS 0.15585f
C3236 DVSS.n3234 VSS 0.15585f
C3237 DVSS.n3235 VSS 0.15585f
C3238 DVSS.n3236 VSS 0.15585f
C3239 DVSS.n3237 VSS 0.15585f
C3240 DVSS.n3238 VSS 0.15585f
C3241 DVSS.n3239 VSS 0.15585f
C3242 DVSS.n3240 VSS 0.15585f
C3243 DVSS.n3241 VSS 0.15585f
C3244 DVSS.n3242 VSS 0.15585f
C3245 DVSS.n3243 VSS 0.15585f
C3246 DVSS.n3244 VSS 0.15585f
C3247 DVSS.n3245 VSS 0.15585f
C3248 DVSS.n3246 VSS 0.15585f
C3249 DVSS.n3247 VSS 0.15585f
C3250 DVSS.n3248 VSS 0.15585f
C3251 DVSS.n3249 VSS 0.15585f
C3252 DVSS.n3250 VSS 0.15585f
C3253 DVSS.n3251 VSS 0.15585f
C3254 DVSS.n3252 VSS 0.15585f
C3255 DVSS.n3253 VSS 0.15585f
C3256 DVSS.n3254 VSS 0.15585f
C3257 DVSS.n3255 VSS 0.15585f
C3258 DVSS.n3256 VSS 0.15585f
C3259 DVSS.n3257 VSS 0.15585f
C3260 DVSS.n3258 VSS 0.15585f
C3261 DVSS.n3259 VSS 0.15585f
C3262 DVSS.n3260 VSS 0.15585f
C3263 DVSS.n3261 VSS 0.15585f
C3264 DVSS.n3262 VSS 0.15585f
C3265 DVSS.n3263 VSS 0.15585f
C3266 DVSS.n3264 VSS 0.15585f
C3267 DVSS.n3265 VSS 0.15585f
C3268 DVSS.n3266 VSS 0.15585f
C3269 DVSS.n3267 VSS 0.15585f
C3270 DVSS.n3268 VSS 0.15585f
C3271 DVSS.n3269 VSS 0.15585f
C3272 DVSS.n3270 VSS 0.15585f
C3273 DVSS.n3271 VSS 0.15585f
C3274 DVSS.n3272 VSS 0.15585f
C3275 DVSS.n3273 VSS 0.15585f
C3276 DVSS.n3274 VSS 0.15585f
C3277 DVSS.n3275 VSS 0.15585f
C3278 DVSS.n3276 VSS 0.15585f
C3279 DVSS.n3277 VSS 0.15585f
C3280 DVSS.n3278 VSS 0.08012f
C3281 DVSS.n3279 VSS 0.15585f
C3282 DVSS.n3280 VSS 0.15585f
C3283 DVSS.n3281 VSS 0.008213f
C3284 DVSS.n3282 VSS 0.050666f
C3285 DVSS.n3283 VSS 0.016098f
C3286 DVSS.n3284 VSS 0.064693f
C3287 DVSS.n3285 VSS 0.006371f
C3288 DVSS.n3286 VSS 0.009203f
C3289 DVSS.n3287 VSS 0.008213f
C3290 DVSS.n3288 VSS 0.008213f
C3291 DVSS.n3289 VSS 0.042748f
C3292 DVSS.n3290 VSS 0.065024f
C3293 DVSS.n3291 VSS 0.193334f
C3294 DVSS.n3292 VSS 0.008213f
C3295 DVSS.n3293 VSS 0.048429f
C3296 DVSS.n3294 VSS 0.28536f
C3297 DVSS.n3295 VSS 0.15585f
C3298 DVSS.n3296 VSS 0.15585f
C3299 DVSS.n3297 VSS 0.15585f
C3300 DVSS.n3298 VSS 0.29749f
C3301 DVSS.n3299 VSS 0.58172f
C3302 DVSS.n3300 VSS 0.153655f
C3303 DVSS.n3301 VSS 0.15585f
C3304 DVSS.n3302 VSS 0.093291f
C3305 DVSS.n3303 VSS 0.093291f
C3306 DVSS.n3304 VSS 0.140485f
C3307 DVSS.n3305 VSS 0.140485f
C3308 DVSS.n3306 VSS 0.15585f
C3309 DVSS.n3307 VSS 0.15585f
C3310 DVSS.n3308 VSS 0.15585f
C3311 DVSS.n3309 VSS 0.15585f
C3312 DVSS.n3310 VSS 0.15585f
C3313 DVSS.n3311 VSS 0.15585f
C3314 DVSS.n3312 VSS 0.15585f
C3315 DVSS.n3313 VSS 0.15585f
C3316 DVSS.n3314 VSS 0.15585f
C3317 DVSS.n3315 VSS 0.15585f
C3318 DVSS.n3316 VSS 0.15585f
C3319 DVSS.n3317 VSS 0.15585f
C3320 DVSS.n3318 VSS 0.15585f
C3321 DVSS.n3319 VSS 0.15585f
C3322 DVSS.n3320 VSS 0.15585f
C3323 DVSS.n3321 VSS 0.15585f
C3324 DVSS.n3322 VSS 0.15585f
C3325 DVSS.n3323 VSS 0.15585f
C3326 DVSS.n3324 VSS 0.15585f
C3327 DVSS.n3325 VSS 0.15585f
C3328 DVSS.n3326 VSS 0.082864f
C3329 DVSS.n3327 VSS 0.54884f
C3330 DVSS.n3328 VSS 0.548383f
C3331 DVSS.n3329 VSS 0.150911f
C3332 DVSS.n3330 VSS 0.15585f
C3333 DVSS.n3331 VSS 0.15585f
C3334 DVSS.n3332 VSS 0.15585f
C3335 DVSS.n3333 VSS 0.15585f
C3336 DVSS.n3334 VSS 0.15585f
C3337 DVSS.n3335 VSS 0.15585f
C3338 DVSS.n3336 VSS 0.15585f
C3339 DVSS.n3337 VSS 0.15585f
C3340 DVSS.n3338 VSS 0.15585f
C3341 DVSS.n3339 VSS 0.15585f
C3342 DVSS.n3340 VSS 0.15585f
C3343 DVSS.n3341 VSS 0.15585f
C3344 DVSS.n3342 VSS 0.15585f
C3345 DVSS.n3343 VSS 0.15585f
C3346 DVSS.n3344 VSS 0.15585f
C3347 DVSS.n3345 VSS 0.15585f
C3348 DVSS.n3346 VSS 0.15585f
C3349 DVSS.n3347 VSS 0.15585f
C3350 DVSS.n3348 VSS 0.15585f
C3351 DVSS.n3349 VSS 0.15585f
C3352 DVSS.n3350 VSS 0.15585f
C3353 DVSS.n3351 VSS 0.15585f
C3354 DVSS.n3352 VSS 0.15585f
C3355 DVSS.n3353 VSS 0.15585f
C3356 DVSS.n3354 VSS 0.15585f
C3357 DVSS.n3355 VSS 0.15585f
C3358 DVSS.n3356 VSS 0.15585f
C3359 DVSS.n3357 VSS 0.15585f
C3360 DVSS.n3358 VSS 0.15585f
C3361 DVSS.n3359 VSS 0.15585f
C3362 DVSS.n3360 VSS 0.15585f
C3363 DVSS.n3361 VSS 0.15585f
C3364 DVSS.n3362 VSS 0.15585f
C3365 DVSS.n3363 VSS 0.15585f
C3366 DVSS.n3364 VSS 0.15585f
C3367 DVSS.n3365 VSS 0.15585f
C3368 DVSS.n3366 VSS 0.15585f
C3369 DVSS.n3367 VSS 0.15585f
C3370 DVSS.n3368 VSS 0.15585f
C3371 DVSS.n3369 VSS 0.15585f
C3372 DVSS.n3370 VSS 0.15585f
C3373 DVSS.n3371 VSS 0.15585f
C3374 DVSS.n3372 VSS 0.15585f
C3375 DVSS.n3373 VSS 0.15585f
C3376 DVSS.n3374 VSS 0.15585f
C3377 DVSS.n3375 VSS 0.15585f
C3378 DVSS.n3376 VSS 0.15585f
C3379 DVSS.n3377 VSS 0.15585f
C3380 DVSS.n3378 VSS 0.15585f
C3381 DVSS.n3379 VSS 0.15585f
C3382 DVSS.n3380 VSS 0.15585f
C3383 DVSS.n3381 VSS 0.15585f
C3384 DVSS.n3382 VSS 0.15585f
C3385 DVSS.n3383 VSS 0.15585f
C3386 DVSS.n3384 VSS 0.15585f
C3387 DVSS.n3385 VSS 0.15585f
C3388 DVSS.n3386 VSS 0.15585f
C3389 DVSS.n3387 VSS 0.15585f
C3390 DVSS.n3388 VSS 0.15585f
C3391 DVSS.n3389 VSS 0.15585f
C3392 DVSS.n3390 VSS 0.15585f
C3393 DVSS.n3391 VSS 0.15585f
C3394 DVSS.n3392 VSS 0.15585f
C3395 DVSS.n3393 VSS 0.15585f
C3396 DVSS.n3394 VSS 0.15585f
C3397 DVSS.n3395 VSS 0.15585f
C3398 DVSS.n3396 VSS 0.15585f
C3399 DVSS.n3397 VSS 0.15585f
C3400 DVSS.n3398 VSS 0.15585f
C3401 DVSS.n3399 VSS 0.15585f
C3402 DVSS.n3400 VSS 0.15585f
C3403 DVSS.n3401 VSS 0.15585f
C3404 DVSS.n3402 VSS 0.15585f
C3405 DVSS.n3403 VSS 0.15585f
C3406 DVSS.n3404 VSS 0.15585f
C3407 DVSS.n3405 VSS 0.15585f
C3408 DVSS.n3406 VSS 0.15585f
C3409 DVSS.n3407 VSS 0.15585f
C3410 DVSS.n3408 VSS 0.15585f
C3411 DVSS.n3409 VSS 0.15585f
C3412 DVSS.n3410 VSS 0.15585f
C3413 DVSS.n3411 VSS 0.15585f
C3414 DVSS.n3412 VSS 0.15585f
C3415 DVSS.n3413 VSS 0.15585f
C3416 DVSS.n3414 VSS 0.15585f
C3417 DVSS.n3415 VSS 0.15585f
C3418 DVSS.n3416 VSS 0.15585f
C3419 DVSS.n3417 VSS 0.15585f
C3420 DVSS.n3418 VSS 0.15585f
C3421 DVSS.n3419 VSS 0.15585f
C3422 DVSS.n3420 VSS 0.15585f
C3423 DVSS.n3421 VSS 0.15585f
C3424 DVSS.n3422 VSS 0.15585f
C3425 DVSS.n3423 VSS 0.15585f
C3426 DVSS.n3424 VSS 0.15585f
C3427 DVSS.n3425 VSS 0.15585f
C3428 DVSS.n3426 VSS 0.15585f
C3429 DVSS.n3427 VSS 0.15585f
C3430 DVSS.n3428 VSS 0.15585f
C3431 DVSS.n3429 VSS 0.15585f
C3432 DVSS.n3430 VSS 0.15585f
C3433 DVSS.n3431 VSS 0.15585f
C3434 DVSS.n3432 VSS 0.15585f
C3435 DVSS.n3433 VSS 0.15585f
C3436 DVSS.n3434 VSS 0.15585f
C3437 DVSS.n3435 VSS 0.15585f
C3438 DVSS.n3436 VSS 0.15585f
C3439 DVSS.n3437 VSS 0.15585f
C3440 DVSS.n3438 VSS 0.15585f
C3441 DVSS.n3439 VSS 0.15585f
C3442 DVSS.n3440 VSS 0.15585f
C3443 DVSS.n3441 VSS 0.15585f
C3444 DVSS.n3442 VSS 0.15585f
C3445 DVSS.n3443 VSS 0.15585f
C3446 DVSS.n3444 VSS 0.15585f
C3447 DVSS.n3445 VSS 0.15585f
C3448 DVSS.n3446 VSS 0.15585f
C3449 DVSS.n3447 VSS 0.15585f
C3450 DVSS.n3448 VSS 0.15585f
C3451 DVSS.n3449 VSS 0.15585f
C3452 DVSS.n3450 VSS 0.15585f
C3453 DVSS.n3451 VSS 0.15585f
C3454 DVSS.n3452 VSS 0.15585f
C3455 DVSS.n3453 VSS 0.15585f
C3456 DVSS.n3454 VSS 0.15585f
C3457 DVSS.n3455 VSS 0.15585f
C3458 DVSS.n3456 VSS 0.15585f
C3459 DVSS.n3457 VSS 0.15585f
C3460 DVSS.n3458 VSS 0.15585f
C3461 DVSS.n3459 VSS 0.15585f
C3462 DVSS.n3460 VSS 0.15585f
C3463 DVSS.n3461 VSS 0.15585f
C3464 DVSS.n3462 VSS 0.15585f
C3465 DVSS.n3463 VSS 0.15585f
C3466 DVSS.n3464 VSS 0.15585f
C3467 DVSS.n3465 VSS 0.15585f
C3468 DVSS.n3466 VSS 0.15585f
C3469 DVSS.n3467 VSS 0.15585f
C3470 DVSS.n3468 VSS 0.15585f
C3471 DVSS.n3469 VSS 0.15585f
C3472 DVSS.n3470 VSS 0.15585f
C3473 DVSS.n3471 VSS 0.15585f
C3474 DVSS.n3472 VSS 0.15585f
C3475 DVSS.n3473 VSS 0.15585f
C3476 DVSS.n3474 VSS 0.15585f
C3477 DVSS.n3475 VSS 0.15585f
C3478 DVSS.n3476 VSS 0.15585f
C3479 DVSS.n3477 VSS 0.15585f
C3480 DVSS.n3478 VSS 0.15585f
C3481 DVSS.n3479 VSS 0.15585f
C3482 DVSS.n3480 VSS 0.15585f
C3483 DVSS.n3481 VSS 0.15585f
C3484 DVSS.n3482 VSS 0.15585f
C3485 DVSS.n3483 VSS 0.15585f
C3486 DVSS.n3484 VSS 0.15585f
C3487 DVSS.n3485 VSS 0.15585f
C3488 DVSS.n3486 VSS 0.15585f
C3489 DVSS.n3487 VSS 0.15585f
C3490 DVSS.n3488 VSS 0.15585f
C3491 DVSS.n3489 VSS 0.15585f
C3492 DVSS.n3490 VSS 0.15585f
C3493 DVSS.n3491 VSS 0.15585f
C3494 DVSS.n3492 VSS 0.15585f
C3495 DVSS.n3493 VSS 0.15585f
C3496 DVSS.n3494 VSS 0.15585f
C3497 DVSS.n3495 VSS 0.15585f
C3498 DVSS.n3496 VSS 0.15585f
C3499 DVSS.n3497 VSS 0.15585f
C3500 DVSS.n3498 VSS 0.15585f
C3501 DVSS.n3499 VSS 0.15585f
C3502 DVSS.n3500 VSS 0.577503f
C3503 DVSS.n3501 VSS 0.292976f
C3504 DVSS.n3502 VSS 0.281067f
C3505 DVSS.n3503 VSS 0.047982f
C3506 DVSS.n3504 VSS 0.082432f
C3507 DVSS.n3505 VSS 0.077523f
C3508 DVSS.n3506 VSS 0.013406f
C3509 DVSS.n3507 VSS 0.036251f
C3510 DVSS.n3508 VSS 0.657695f
C3511 DVSS.n3509 VSS 1.68676f
C3512 DVSS.n3510 VSS 0.661498f
C3513 DVSS.n3511 VSS 0.036251f
C3514 DVSS.n3512 VSS 0.008213f
C3515 DVSS.n3513 VSS 0.077523f
C3516 DVSS.n3514 VSS 0.082432f
C3517 DVSS.n3515 VSS 1.76722f
C3518 DVSS.n3516 VSS 1.88785f
C3519 DVSS.n3517 VSS 0.869181f
C3520 DVSS.n3518 VSS 16.1392f
C3521 DVSS.n3519 VSS 3.60328f
C3522 DVSS.n3520 VSS 0.036571f
C3523 DVSS.n3521 VSS 0.009721f
C3524 DVSS.n3522 VSS 0.161646f
C3525 DVSS.t26 VSS 0.311996f
C3526 DVSS.n3523 VSS 0.599743f
C3527 DVSS.n3524 VSS 0.531318f
C3528 DVSS.n3525 VSS 0.091673f
C3529 DVSS.n3526 VSS 0.009721f
C3530 DVSS.n3527 VSS 0.106545f
C3531 DVSS.n3528 VSS 0.185052f
C3532 DVSS.n3529 VSS 0.026052f
C3533 DVSS.n3530 VSS 0.185052f
C3534 DVSS.n3531 VSS 0.106545f
C3535 DVSS.n3532 VSS 0.009721f
C3536 DVSS.n3533 VSS 0.091673f
C3537 DVSS.n3534 VSS 0.531318f
C3538 DVSS.n3535 VSS 0.009721f
C3539 DVSS.n3537 VSS 0.161646f
C3540 DVSS.n3538 VSS 0.009721f
C3541 DVSS.n3539 VSS 0.018658f
C3542 DVSS.n3540 VSS 2.1675f
C3543 DVSS.n3541 VSS 0.019442f
C3544 DVSS.n3542 VSS 0.009721f
C3545 DVSS.n3543 VSS 0.077925f
C3546 DVSS.n3544 VSS 0.288809f
C3547 DVSS.n3545 VSS 0.288809f
C3548 DVSS.n3546 VSS 2.1675f
C3549 DVSS.n3547 VSS 3.71965f
C3550 DVSS.n3548 VSS 0.15585f
C3551 DVSS.n3549 VSS 0.15585f
C3552 DVSS.n3550 VSS 0.15585f
C3553 DVSS.n3551 VSS 0.15585f
C3554 DVSS.n3552 VSS 0.15585f
C3555 DVSS.n3553 VSS 0.15585f
C3556 DVSS.n3554 VSS 0.15585f
C3557 DVSS.n3555 VSS 0.15585f
C3558 DVSS.n3556 VSS 0.15585f
C3559 DVSS.n3557 VSS 0.15585f
C3560 DVSS.n3558 VSS 0.15585f
C3561 DVSS.n3559 VSS 0.15585f
C3562 DVSS.n3560 VSS 0.15585f
C3563 DVSS.n3561 VSS 0.15585f
C3564 DVSS.n3562 VSS 0.15585f
C3565 DVSS.n3563 VSS 0.15585f
C3566 DVSS.n3564 VSS 0.149814f
C3567 DVSS.n3565 VSS 0.15585f
C3568 DVSS.n3566 VSS 0.15585f
C3569 DVSS.n3567 VSS 0.15585f
C3570 DVSS.n3568 VSS 0.15585f
C3571 DVSS.n3569 VSS 0.15585f
C3572 DVSS.n3570 VSS 0.15585f
C3573 DVSS.n3571 VSS 0.15585f
C3574 DVSS.n3572 VSS 0.15585f
C3575 DVSS.n3573 VSS 0.15585f
C3576 DVSS.n3574 VSS 0.15585f
C3577 DVSS.n3575 VSS 0.15585f
C3578 DVSS.n3576 VSS 0.15585f
C3579 DVSS.n3577 VSS 0.068047f
C3580 DVSS.n3578 VSS 0.15585f
C3581 DVSS.n3579 VSS 0.15585f
C3582 DVSS.n3580 VSS 0.15585f
C3583 DVSS.n3581 VSS 0.15585f
C3584 DVSS.n3582 VSS 0.15585f
C3585 DVSS.n3583 VSS 0.15585f
C3586 DVSS.n3584 VSS 0.15585f
C3587 DVSS.n3585 VSS 0.15585f
C3588 DVSS.n3586 VSS 0.15585f
C3589 DVSS.n3587 VSS 0.15585f
C3590 DVSS.n3588 VSS 0.15585f
C3591 DVSS.n3589 VSS 0.15585f
C3592 DVSS.n3590 VSS 0.15585f
C3593 DVSS.n3591 VSS 0.15585f
C3594 DVSS.n3592 VSS 0.15585f
C3595 DVSS.n3593 VSS 0.15585f
C3596 DVSS.n3594 VSS 0.15585f
C3597 DVSS.n3595 VSS 0.15585f
C3598 DVSS.n3596 VSS 0.15585f
C3599 DVSS.n3597 VSS 0.15585f
C3600 DVSS.n3598 VSS 0.15585f
C3601 DVSS.n3599 VSS 0.15585f
C3602 DVSS.n3600 VSS 0.15585f
C3603 DVSS.n3601 VSS 0.15585f
C3604 DVSS.n3602 VSS 0.15585f
C3605 DVSS.n3603 VSS 0.15585f
C3606 DVSS.n3604 VSS 0.15585f
C3607 DVSS.n3605 VSS 0.15585f
C3608 DVSS.n3606 VSS 0.15585f
C3609 DVSS.n3607 VSS 0.15585f
C3610 DVSS.n3608 VSS 0.15585f
C3611 DVSS.n3609 VSS 0.15585f
C3612 DVSS.n3610 VSS 0.15585f
C3613 DVSS.n3611 VSS 0.15585f
C3614 DVSS.n3612 VSS 0.15585f
C3615 DVSS.n3613 VSS 0.15585f
C3616 DVSS.n3614 VSS 0.15585f
C3617 DVSS.n3615 VSS 0.15585f
C3618 DVSS.n3616 VSS 0.15585f
C3619 DVSS.n3617 VSS 0.15585f
C3620 DVSS.n3618 VSS 0.15585f
C3621 DVSS.n3619 VSS 0.091644f
C3622 DVSS.n3620 VSS 0.15585f
C3623 DVSS.n3621 VSS 0.15585f
C3624 DVSS.n3622 VSS 0.15585f
C3625 DVSS.n3623 VSS 0.15585f
C3626 DVSS.n3624 VSS 0.15585f
C3627 DVSS.n3625 VSS 0.15585f
C3628 DVSS.n3626 VSS 0.093839f
C3629 DVSS.n3627 VSS 0.15585f
C3630 DVSS.n3628 VSS 0.15585f
C3631 DVSS.n3629 VSS 0.15585f
C3632 DVSS.n3630 VSS 0.15585f
C3633 DVSS.n3631 VSS 0.15585f
C3634 DVSS.n3632 VSS 0.15585f
C3635 DVSS.n3633 VSS 0.15585f
C3636 DVSS.n3634 VSS 0.15585f
C3637 DVSS.n3635 VSS 0.15585f
C3638 DVSS.n3636 VSS 0.15585f
C3639 DVSS.n3637 VSS 0.15585f
C3640 DVSS.n3638 VSS 0.15585f
C3641 DVSS.n3639 VSS 0.15585f
C3642 DVSS.n3640 VSS 0.15585f
C3643 DVSS.n3641 VSS 0.15585f
C3644 DVSS.n3642 VSS 0.15585f
C3645 DVSS.n3643 VSS 0.15585f
C3646 DVSS.n3644 VSS 0.15585f
C3647 DVSS.n3645 VSS 0.15585f
C3648 DVSS.n3646 VSS 0.15585f
C3649 DVSS.n3647 VSS 0.15585f
C3650 DVSS.n3648 VSS 0.15585f
C3651 DVSS.n3649 VSS 0.15585f
C3652 DVSS.n3650 VSS 0.15585f
C3653 DVSS.n3651 VSS 0.15585f
C3654 DVSS.n3652 VSS 0.15585f
C3655 DVSS.n3653 VSS 0.15585f
C3656 DVSS.n3654 VSS 0.15585f
C3657 DVSS.n3655 VSS 0.15585f
C3658 DVSS.n3656 VSS 0.15585f
C3659 DVSS.n3657 VSS 0.068047f
C3660 DVSS.n3658 VSS 0.15585f
C3661 DVSS.n3659 VSS 0.15585f
C3662 DVSS.n3660 VSS 0.093839f
C3663 DVSS.n3661 VSS 0.15585f
C3664 DVSS.n3662 VSS 0.15585f
C3665 DVSS.n3663 VSS 0.15585f
C3666 DVSS.n3664 VSS 0.15585f
C3667 DVSS.n3665 VSS 0.15585f
C3668 DVSS.n3666 VSS 0.15585f
C3669 DVSS.n3667 VSS 0.15585f
C3670 DVSS.n3668 VSS 0.15585f
C3671 DVSS.n3669 VSS 0.15585f
C3672 DVSS.n3670 VSS 0.15585f
C3673 DVSS.n3671 VSS 0.15585f
C3674 DVSS.n3672 VSS 0.15585f
C3675 DVSS.n3673 VSS 0.15585f
C3676 DVSS.n3674 VSS 0.15585f
C3677 DVSS.n3675 VSS 0.15585f
C3678 DVSS.n3676 VSS 0.15585f
C3679 DVSS.n3677 VSS 0.15585f
C3680 DVSS.n3678 VSS 0.15585f
C3681 DVSS.n3679 VSS 0.15585f
C3682 DVSS.n3680 VSS 0.15585f
C3683 DVSS.n3681 VSS 0.15585f
C3684 DVSS.n3682 VSS 0.15585f
C3685 DVSS.n3683 VSS 0.15585f
C3686 DVSS.n3684 VSS 0.15585f
C3687 DVSS.n3685 VSS 0.15585f
C3688 DVSS.n3686 VSS 0.15585f
C3689 DVSS.n3687 VSS 0.15585f
C3690 DVSS.n3688 VSS 0.15585f
C3691 DVSS.n3689 VSS 2.43723f
C3692 DVSS.n3690 VSS 0.15585f
C3693 DVSS.n3691 VSS 0.125668f
C3694 DVSS.n3692 VSS 0.077925f
C3695 DVSS.n3693 VSS 0.163376f
C3696 DVSS.n3694 VSS 0.163376f
C3697 DVSS.n3695 VSS 2.1675f
C3698 DVSS.n3696 VSS 3.71965f
C3699 DVSS.n3697 VSS 0.15585f
C3700 DVSS.n3698 VSS 0.15585f
C3701 DVSS.n3699 VSS 0.15585f
C3702 DVSS.n3700 VSS 0.15585f
C3703 DVSS.n3701 VSS 0.15585f
C3704 DVSS.n3702 VSS 0.15585f
C3705 DVSS.n3703 VSS 0.15585f
C3706 DVSS.n3704 VSS 0.15585f
C3707 DVSS.n3705 VSS 0.15585f
C3708 DVSS.n3706 VSS 0.15585f
C3709 DVSS.n3707 VSS 0.15585f
C3710 DVSS.n3708 VSS 0.15585f
C3711 DVSS.n3709 VSS 0.15585f
C3712 DVSS.n3710 VSS 0.15585f
C3713 DVSS.n3711 VSS 0.15585f
C3714 DVSS.n3712 VSS 0.15585f
C3715 DVSS.n3713 VSS 0.149814f
C3716 DVSS.n3714 VSS 0.15585f
C3717 DVSS.n3715 VSS 0.15585f
C3718 DVSS.n3716 VSS 0.15585f
C3719 DVSS.n3717 VSS 0.15585f
C3720 DVSS.n3718 VSS 0.15585f
C3721 DVSS.n3719 VSS 0.15585f
C3722 DVSS.n3720 VSS 0.15585f
C3723 DVSS.n3721 VSS 0.15585f
C3724 DVSS.n3722 VSS 0.15585f
C3725 DVSS.n3723 VSS 0.15585f
C3726 DVSS.n3724 VSS 0.15585f
C3727 DVSS.n3725 VSS 0.15585f
C3728 DVSS.n3726 VSS 0.077925f
C3729 DVSS.n3727 VSS 0.15585f
C3730 DVSS.n3728 VSS 0.15585f
C3731 DVSS.n3729 VSS 0.15585f
C3732 DVSS.n3730 VSS 0.071889f
C3733 DVSS.n3731 VSS 0.052105f
C3734 DVSS.n3732 VSS 0.052105f
C3735 DVSS.n3733 VSS 0.052105f
C3736 DVSS.n3734 VSS 0.052105f
C3737 DVSS.n3735 VSS 0.052105f
C3738 DVSS.n3736 VSS 0.15585f
C3739 DVSS.n3737 VSS 0.15585f
C3740 DVSS.n3738 VSS 0.15585f
C3741 DVSS.n3739 VSS 0.15585f
C3742 DVSS.n3740 VSS 0.15585f
C3743 DVSS.n3741 VSS 0.15585f
C3744 DVSS.n3742 VSS 0.15585f
C3745 DVSS.n3743 VSS 0.15585f
C3746 DVSS.n3744 VSS 0.15585f
C3747 DVSS.n3745 VSS 0.15585f
C3748 DVSS.n3746 VSS 0.15585f
C3749 DVSS.n3747 VSS 0.15585f
C3750 DVSS.n3748 VSS 0.15585f
C3751 DVSS.n3749 VSS 0.15585f
C3752 DVSS.n3750 VSS 0.019442f
C3753 DVSS.n3751 VSS 0.019442f
C3754 DVSS.n3752 VSS 0.019442f
C3755 DVSS.n3753 VSS 0.019442f
C3756 DVSS.n3754 VSS 0.163376f
C3757 DVSS.n3755 VSS 0.163376f
C3758 DVSS.n3756 VSS 0.077925f
C3759 DVSS.n3757 VSS 0.152009f
C3760 DVSS.n3758 VSS 0.15585f
C3761 DVSS.n3759 VSS 0.15585f
C3762 DVSS.n3760 VSS 0.15585f
C3763 DVSS.n3761 VSS 0.15585f
C3764 DVSS.n3762 VSS 0.15585f
C3765 DVSS.n3763 VSS 0.15585f
C3766 DVSS.n3764 VSS 0.15585f
C3767 DVSS.n3765 VSS 0.15585f
C3768 DVSS.n3766 VSS 0.15585f
C3769 DVSS.n3767 VSS 0.15585f
C3770 DVSS.n3768 VSS 0.15585f
C3771 DVSS.n3769 VSS 0.15585f
C3772 DVSS.n3770 VSS 0.15585f
C3773 DVSS.n3771 VSS 0.15585f
C3774 DVSS.n3772 VSS 0.15585f
C3775 DVSS.n3773 VSS 0.15585f
C3776 DVSS.n3774 VSS 0.15585f
C3777 DVSS.n3775 VSS 0.15585f
C3778 DVSS.n3776 VSS 0.15585f
C3779 DVSS.n3777 VSS 0.15585f
C3780 DVSS.n3778 VSS 0.15585f
C3781 DVSS.n3779 VSS 0.15585f
C3782 DVSS.n3780 VSS 0.15585f
C3783 DVSS.n3781 VSS 0.15585f
C3784 DVSS.n3782 VSS 0.15585f
C3785 DVSS.n3783 VSS 0.15585f
C3786 DVSS.n3784 VSS 0.15585f
C3787 DVSS.n3785 VSS 0.15585f
C3788 DVSS.n3786 VSS 0.15585f
C3789 DVSS.n3787 VSS 0.15585f
C3790 DVSS.n3788 VSS 0.091644f
C3791 DVSS.n3790 VSS 1.63058f
C3792 DVSS.n3791 VSS 0.46264f
C3793 DVSS.n3794 VSS 0.052105f
C3794 DVSS.n3797 VSS 0.052105f
C3795 DVSS.n3800 VSS 0.052105f
C3796 DVSS.n3803 VSS 0.052105f
C3797 DVSS.n3804 VSS 0.437848f
C3798 DVSS.n3806 VSS 0.068047f
C3799 DVSS.n3807 VSS 0.074084f
C3800 DVSS.n3809 VSS 0.437848f
C3801 DVSS.n3810 VSS 0.077925f
C3802 DVSS.n3811 VSS 0.068047f
C3803 DVSS.n3812 VSS 0.15585f
C3804 DVSS.n3813 VSS 0.15585f
C3805 DVSS.n3814 VSS 0.15585f
C3806 DVSS.n3815 VSS 0.15585f
C3807 DVSS.n3816 VSS 0.15585f
C3808 DVSS.n3817 VSS 0.093839f
C3809 DVSS.n3818 VSS 0.15585f
C3810 DVSS.n3819 VSS 0.15585f
C3811 DVSS.n3820 VSS 0.15585f
C3812 DVSS.n3821 VSS 0.15585f
C3813 DVSS.n3822 VSS 0.15585f
C3814 DVSS.n3823 VSS 0.15585f
C3815 DVSS.n3824 VSS 0.15585f
C3816 DVSS.n3825 VSS 0.15585f
C3817 DVSS.n3826 VSS 0.15585f
C3818 DVSS.n3827 VSS 0.15585f
C3819 DVSS.n3828 VSS 0.15585f
C3820 DVSS.n3829 VSS 0.15585f
C3821 DVSS.n3830 VSS 0.15585f
C3822 DVSS.n3831 VSS 0.15585f
C3823 DVSS.n3832 VSS 0.15585f
C3824 DVSS.n3833 VSS 0.15585f
C3825 DVSS.n3834 VSS 0.15585f
C3826 DVSS.n3835 VSS 0.15585f
C3827 DVSS.n3836 VSS 0.15585f
C3828 DVSS.n3837 VSS 0.15585f
C3829 DVSS.n3838 VSS 0.15585f
C3830 DVSS.n3839 VSS 0.15585f
C3831 DVSS.n3840 VSS 0.15585f
C3832 DVSS.n3841 VSS 0.15585f
C3833 DVSS.n3842 VSS 0.15585f
C3834 DVSS.n3843 VSS 0.15585f
C3835 DVSS.n3844 VSS 0.15585f
C3836 DVSS.n3845 VSS 0.15585f
C3837 DVSS.n3846 VSS 0.15585f
C3838 DVSS.n3847 VSS 0.15585f
C3839 DVSS.n3848 VSS 0.068047f
C3840 DVSS.n3849 VSS 0.15585f
C3841 DVSS.n3850 VSS 0.15585f
C3842 DVSS.n3851 VSS 0.093839f
C3843 DVSS.n3852 VSS 0.15585f
C3844 DVSS.n3853 VSS 0.15585f
C3845 DVSS.n3854 VSS 0.15585f
C3846 DVSS.n3855 VSS 0.15585f
C3847 DVSS.n3856 VSS 0.15585f
C3848 DVSS.n3857 VSS 0.15585f
C3849 DVSS.n3858 VSS 0.15585f
C3850 DVSS.n3859 VSS 0.15585f
C3851 DVSS.n3860 VSS 0.15585f
C3852 DVSS.n3861 VSS 0.15585f
C3853 DVSS.n3862 VSS 0.15585f
C3854 DVSS.n3863 VSS 0.15585f
C3855 DVSS.n3864 VSS 0.15585f
C3856 DVSS.n3865 VSS 0.15585f
C3857 DVSS.n3866 VSS 0.15585f
C3858 DVSS.n3867 VSS 0.15585f
C3859 DVSS.n3868 VSS 0.15585f
C3860 DVSS.n3869 VSS 0.15585f
C3861 DVSS.n3870 VSS 0.15585f
C3862 DVSS.n3871 VSS 0.15585f
C3863 DVSS.n3872 VSS 0.15585f
C3864 DVSS.n3873 VSS 0.15585f
C3865 DVSS.n3874 VSS 0.15585f
C3866 DVSS.n3875 VSS 0.15585f
C3867 DVSS.n3876 VSS 0.15585f
C3868 DVSS.n3877 VSS 0.15585f
C3869 DVSS.n3878 VSS 0.15585f
C3870 DVSS.n3879 VSS 0.15585f
C3871 DVSS.n3880 VSS 2.43723f
C3872 DVSS.n3881 VSS 0.15585f
C3873 DVSS.n3882 VSS 0.125668f
C3874 DVSS.n3883 VSS 0.077925f
C3875 DVSS.n3884 VSS 0.172627f
C3876 DVSS.n3885 VSS 0.63273f
C3877 DVSS.n3886 VSS 0.015908f
C3878 DVSS.n3887 VSS 0.063632f
C3879 DVSS.n3888 VSS 0.016313f
C3880 DVSS.n3889 VSS 0.018232f
C3881 DVSS.n3890 VSS 1.33697f
C3882 DVSS.n3891 VSS 1.13742f
C3883 DVSS.n3892 VSS 0.018232f
C3884 DVSS.n3893 VSS 0.016313f
C3885 DVSS.n3894 VSS 0.018232f
C3886 DVSS.n3895 VSS 2.1675f
C3887 DVSS.n3896 VSS 0.068047f
C3888 DVSS.n3897 VSS 0.15585f
C3889 DVSS.n3898 VSS 0.506941f
C3890 DVSS.n3899 VSS 0.15585f
C3891 DVSS.n3900 VSS 3.71965f
C3892 DVSS.n3901 VSS 0.15585f
C3893 DVSS.n3902 VSS 0.15585f
C3894 DVSS.n3903 VSS 0.15585f
C3895 DVSS.n3904 VSS 0.15585f
C3896 DVSS.n3905 VSS 0.15585f
C3897 DVSS.n3906 VSS 0.15585f
C3898 DVSS.n3907 VSS 0.15585f
C3899 DVSS.n3908 VSS 0.15585f
C3900 DVSS.n3909 VSS 0.15585f
C3901 DVSS.n3910 VSS 0.15585f
C3902 DVSS.n3911 VSS 0.15585f
C3903 DVSS.n3912 VSS 0.15585f
C3904 DVSS.n3913 VSS 0.15585f
C3905 DVSS.n3914 VSS 0.15585f
C3906 DVSS.n3915 VSS 0.15585f
C3907 DVSS.n3916 VSS 0.15585f
C3908 DVSS.n3917 VSS 0.15585f
C3909 DVSS.n3918 VSS 0.15585f
C3910 DVSS.n3919 VSS 0.15585f
C3911 DVSS.n3920 VSS 0.15585f
C3912 DVSS.n3921 VSS 0.15585f
C3913 DVSS.n3922 VSS 0.15585f
C3914 DVSS.n3923 VSS 0.15585f
C3915 DVSS.n3924 VSS 0.15585f
C3916 DVSS.n3925 VSS 0.15585f
C3917 DVSS.n3926 VSS 0.15585f
C3918 DVSS.n3927 VSS 0.15585f
C3919 DVSS.n3928 VSS 0.15585f
C3920 DVSS.n3929 VSS 0.15585f
C3921 DVSS.n3930 VSS 0.15585f
C3922 DVSS.n3931 VSS 0.15585f
C3923 DVSS.n3932 VSS 0.15585f
C3924 DVSS.n3933 VSS 0.15585f
C3925 DVSS.n3934 VSS 0.15585f
C3926 DVSS.n3935 VSS 0.15585f
C3927 DVSS.n3936 VSS 0.15585f
C3928 DVSS.n3937 VSS 0.15585f
C3929 DVSS.n3938 VSS 2.43723f
C3930 DVSS.n3939 VSS 0.15585f
C3931 DVSS.n3940 VSS 0.125668f
C3932 DVSS.n3941 VSS 0.077925f
C3933 DVSS.n3942 VSS 0.038884f
C3934 DVSS.n3943 VSS 0.009721f
C3935 DVSS.n3944 VSS 0.019442f
C3936 DVSS.n3945 VSS 0.019442f
C3937 DVSS.n3946 VSS 0.019442f
C3938 DVSS.n3947 VSS 0.019442f
C3939 DVSS.n3948 VSS 0.019442f
C3940 DVSS.n3949 VSS 0.019442f
C3941 DVSS.n3950 VSS 0.019442f
C3942 DVSS.n3951 VSS 0.019442f
C3943 DVSS.n3952 VSS 0.009721f
C3944 DVSS.n3953 VSS 0.182034f
C3945 DVSS.n3954 VSS 0.40405f
C3946 DVSS.n3955 VSS 0.008222f
C3947 DVSS.n3956 VSS 0.016444f
C3948 DVSS.n3957 VSS 0.018232f
C3949 DVSS.n3958 VSS 1.13742f
C3950 DVSS.n3959 VSS 0.018232f
C3951 DVSS.n3960 VSS 0.018232f
C3952 DVSS.n3961 VSS 0.063632f
C3953 DVSS.n3962 VSS 0.018232f
C3954 DVSS.n3963 VSS 1.13742f
C3955 DVSS.n3964 VSS 0.018232f
C3956 DVSS.n3965 VSS 0.018232f
C3957 DVSS.n3966 VSS 0.016444f
C3958 DVSS.n3967 VSS 0.018232f
C3959 DVSS.n3968 VSS 1.13742f
C3960 DVSS.n3969 VSS 0.018232f
C3961 DVSS.n3970 VSS 0.018232f
C3962 DVSS.n3971 VSS 0.063632f
C3963 DVSS.n3972 VSS 0.018232f
C3964 DVSS.n3973 VSS 1.13742f
C3965 DVSS.n3974 VSS 0.018232f
C3966 DVSS.n3975 VSS 0.018232f
C3967 DVSS.n3976 VSS 0.016444f
C3968 DVSS.n3977 VSS 0.018232f
C3969 DVSS.n3978 VSS 1.13742f
C3970 DVSS.n3979 VSS 0.018232f
C3971 DVSS.n3980 VSS 0.018232f
C3972 DVSS.n3981 VSS 0.063632f
C3973 DVSS.n3982 VSS 0.018232f
C3974 DVSS.n3983 VSS 1.13742f
C3975 DVSS.n3984 VSS 0.018232f
C3976 DVSS.n3985 VSS 0.018232f
C3977 DVSS.n3986 VSS 0.016444f
C3978 DVSS.n3987 VSS 0.018232f
C3979 DVSS.n3988 VSS 1.13742f
C3980 DVSS.n3989 VSS 0.018232f
C3981 DVSS.n3990 VSS 0.018232f
C3982 DVSS.n3991 VSS 0.063632f
C3983 DVSS.n3992 VSS 0.018232f
C3984 DVSS.n3993 VSS 1.13742f
C3985 DVSS.n3994 VSS 0.018232f
C3986 DVSS.n3995 VSS 0.018232f
C3987 DVSS.n3996 VSS 0.01017f
C3988 DVSS.n3997 VSS 0.016444f
C3989 DVSS.n3998 VSS 0.018232f
C3990 DVSS.n3999 VSS 1.13742f
C3991 DVSS.n4000 VSS 0.018232f
C3992 DVSS.n4001 VSS 0.018232f
C3993 DVSS.n4002 VSS 0.013858f
C3994 DVSS.n4003 VSS 0.016313f
C3995 DVSS.n4005 VSS 1.33697f
C3996 DVSS.n4007 VSS 0.015436f
C3997 DVSS.n4008 VSS 0.018232f
C3998 DVSS.n4009 VSS 0.018232f
C3999 DVSS.n4035 VSS 0.018232f
C4000 DVSS.n4036 VSS 0.018232f
C4001 DVSS.n4037 VSS 0.018232f
C4002 DVSS.n4061 VSS 0.018232f
C4003 DVSS.n4063 VSS 0.018232f
C4004 DVSS.n4064 VSS 0.018232f
C4005 DVSS.n4066 VSS 0.014785f
C4006 DVSS.n4067 VSS 0.015218f
C4007 DVSS.t9 VSS 0.519282f
C4008 DVSS.n4068 VSS 0.111753f
C4009 DVSS.n4069 VSS 0.043773f
C4010 DVSS.n4071 VSS 0.018232f
C4011 DVSS.n4072 VSS 0.052908f
C4012 DVSS.n4073 VSS 0.052908f
C4013 DVSS.n4074 VSS 0.018232f
C4014 DVSS.n4076 VSS 0.018232f
C4015 DVSS.n4077 VSS 0.052908f
C4016 DVSS.n4078 VSS 0.052908f
C4017 DVSS.n4079 VSS 0.018232f
C4018 DVSS.n4081 VSS 0.018232f
C4019 DVSS.n4082 VSS 0.052908f
C4020 DVSS.n4083 VSS 0.052908f
C4021 DVSS.n4084 VSS 0.018232f
C4022 DVSS.n4086 VSS 0.018232f
C4023 DVSS.n4087 VSS 0.052908f
C4024 DVSS.n4088 VSS 0.052908f
C4025 DVSS.n4089 VSS 0.018232f
C4026 DVSS.n4091 VSS 0.018232f
C4027 DVSS.n4092 VSS 0.052908f
C4028 DVSS.n4093 VSS 0.052908f
C4029 DVSS.n4094 VSS 0.018232f
C4030 DVSS.n4096 VSS 0.018232f
C4031 DVSS.n4097 VSS 0.052908f
C4032 DVSS.n4098 VSS 0.052908f
C4033 DVSS.n4099 VSS 0.018232f
C4034 DVSS.n4101 VSS 0.018232f
C4035 DVSS.n4102 VSS 0.052908f
C4036 DVSS.n4103 VSS 0.052908f
C4037 DVSS.n4104 VSS 0.018232f
C4038 DVSS.n4106 VSS 0.018232f
C4039 DVSS.n4107 VSS 0.052908f
C4040 DVSS.n4108 VSS 0.052908f
C4041 DVSS.n4109 VSS 0.018232f
C4042 DVSS.n4111 VSS 0.018232f
C4043 DVSS.n4112 VSS 0.052908f
C4044 DVSS.n4113 VSS 0.052908f
C4045 DVSS.n4114 VSS 0.018232f
C4046 DVSS.n4116 VSS 0.018232f
C4047 DVSS.n4117 VSS 0.052908f
C4048 DVSS.n4118 VSS 0.052908f
C4049 DVSS.n4119 VSS 0.018232f
C4050 DVSS.n4121 VSS 0.018232f
C4051 DVSS.n4122 VSS 0.045018f
C4052 DVSS.t3 VSS 0.519282f
C4053 DVSS.n4123 VSS 0.111753f
C4054 DVSS.n4124 VSS 0.034343f
C4055 DVSS.n4125 VSS 0.018232f
C4056 DVSS.n4127 VSS 0.018232f
C4057 DVSS.n4128 VSS 0.032719f
C4058 DVSS.n4129 VSS 0.046642f
C4059 DVSS.n4130 VSS 0.018232f
C4060 DVSS.n4132 VSS 0.018232f
C4061 DVSS.n4133 VSS 0.052908f
C4062 DVSS.n4134 VSS 0.052908f
C4063 DVSS.n4135 VSS 0.018232f
C4064 DVSS.n4137 VSS 0.018232f
C4065 DVSS.n4138 VSS 0.052908f
C4066 DVSS.n4139 VSS 0.052908f
C4067 DVSS.n4140 VSS 0.018232f
C4068 DVSS.n4142 VSS 0.018232f
C4069 DVSS.n4143 VSS 0.052908f
C4070 DVSS.n4144 VSS 0.052908f
C4071 DVSS.n4145 VSS 0.018232f
C4072 DVSS.n4147 VSS 0.018232f
C4073 DVSS.n4148 VSS 0.052908f
C4074 DVSS.n4149 VSS 0.052908f
C4075 DVSS.n4150 VSS 0.018232f
C4076 DVSS.n4152 VSS 0.018232f
C4077 DVSS.n4153 VSS 0.052908f
C4078 DVSS.n4154 VSS 0.052908f
C4079 DVSS.n4155 VSS 0.018232f
C4080 DVSS.n4157 VSS 0.018232f
C4081 DVSS.n4158 VSS 0.052908f
C4082 DVSS.n4159 VSS 0.052908f
C4083 DVSS.n4160 VSS 0.018232f
C4084 DVSS.n4162 VSS 0.018232f
C4085 DVSS.n4163 VSS 0.052908f
C4086 DVSS.n4164 VSS 0.052908f
C4087 DVSS.n4165 VSS 0.018232f
C4088 DVSS.n4167 VSS 0.018232f
C4089 DVSS.n4168 VSS 0.052908f
C4090 DVSS.n4169 VSS 0.052908f
C4091 DVSS.n4170 VSS 0.018232f
C4092 DVSS.n4172 VSS 0.018232f
C4093 DVSS.n4173 VSS 0.052908f
C4094 DVSS.n4174 VSS 0.052908f
C4095 DVSS.n4175 VSS 0.018232f
C4096 DVSS.n4177 VSS 0.018232f
C4097 DVSS.n4178 VSS 0.052908f
C4098 DVSS.n4180 VSS 0.018232f
C4099 DVSS.n4181 VSS 0.051515f
C4100 DVSS.n4182 VSS 0.050794f
C4101 DVSS.n4184 VSS 0.018232f
C4102 DVSS.n4189 VSS 0.073121f
C4103 DVSS.n4190 VSS 0.08939f
C4104 DVSS.n4191 VSS 0.047802f
C4105 DVSS.n4192 VSS 0.018232f
C4106 DVSS.n4194 VSS 0.018232f
C4107 DVSS.n4195 VSS 0.052908f
C4108 DVSS.n4196 VSS 0.052908f
C4109 DVSS.n4197 VSS 0.018232f
C4110 DVSS.n4199 VSS 0.018232f
C4111 DVSS.n4200 VSS 0.052908f
C4112 DVSS.n4201 VSS 0.052908f
C4113 DVSS.n4202 VSS 0.018232f
C4114 DVSS.n4204 VSS 0.018232f
C4115 DVSS.n4205 VSS 0.052908f
C4116 DVSS.n4206 VSS 0.052908f
C4117 DVSS.n4207 VSS 0.018232f
C4118 DVSS.n4209 VSS 0.018232f
C4119 DVSS.n4210 VSS 0.052908f
C4120 DVSS.n4211 VSS 0.052908f
C4121 DVSS.n4212 VSS 0.018232f
C4122 DVSS.n4214 VSS 0.018232f
C4123 DVSS.n4215 VSS 0.052908f
C4124 DVSS.n4216 VSS 0.052908f
C4125 DVSS.n4217 VSS 0.018232f
C4126 DVSS.n4219 VSS 0.018232f
C4127 DVSS.n4220 VSS 0.052908f
C4128 DVSS.n4221 VSS 0.052908f
C4129 DVSS.n4222 VSS 0.018232f
C4130 DVSS.n4224 VSS 0.018232f
C4131 DVSS.n4225 VSS 0.052908f
C4132 DVSS.n4226 VSS 0.052908f
C4133 DVSS.n4227 VSS 0.018232f
C4134 DVSS.n4229 VSS 0.018232f
C4135 DVSS.n4230 VSS 0.052908f
C4136 DVSS.n4231 VSS 0.052908f
C4137 DVSS.n4232 VSS 0.018232f
C4138 DVSS.n4234 VSS 0.018232f
C4139 DVSS.n4235 VSS 0.052908f
C4140 DVSS.n4236 VSS 0.052908f
C4141 DVSS.n4237 VSS 0.018232f
C4142 DVSS.n4239 VSS 0.018232f
C4143 DVSS.n4240 VSS 0.052908f
C4144 DVSS.n4241 VSS 0.050355f
C4145 DVSS.n4242 VSS 0.018232f
C4146 DVSS.n4244 VSS 0.018232f
C4147 DVSS.n4245 VSS 0.029006f
C4148 DVSS.n4246 VSS 0.038056f
C4149 DVSS.n4247 VSS 0.018232f
C4150 DVSS.n4249 VSS 0.018232f
C4151 DVSS.n4250 VSS 0.041305f
C4152 DVSS.n4251 VSS 0.052908f
C4153 DVSS.n4252 VSS 0.018232f
C4154 DVSS.n4254 VSS 0.018232f
C4155 DVSS.n4255 VSS 0.052908f
C4156 DVSS.n4256 VSS 0.052908f
C4157 DVSS.n4257 VSS 0.018232f
C4158 DVSS.n4259 VSS 0.018232f
C4159 DVSS.n4260 VSS 0.052908f
C4160 DVSS.n4261 VSS 0.052908f
C4161 DVSS.n4262 VSS 0.018232f
C4162 DVSS.n4264 VSS 0.018232f
C4163 DVSS.n4265 VSS 0.052908f
C4164 DVSS.n4266 VSS 0.052908f
C4165 DVSS.n4267 VSS 0.018232f
C4166 DVSS.n4269 VSS 0.018232f
C4167 DVSS.n4270 VSS 0.052908f
C4168 DVSS.n4271 VSS 0.052908f
C4169 DVSS.n4272 VSS 0.018232f
C4170 DVSS.n4274 VSS 0.018232f
C4171 DVSS.n4275 VSS 0.052908f
C4172 DVSS.n4276 VSS 0.052908f
C4173 DVSS.n4277 VSS 0.018232f
C4174 DVSS.n4279 VSS 0.018232f
C4175 DVSS.n4280 VSS 0.052908f
C4176 DVSS.n4281 VSS 0.052908f
C4177 DVSS.n4282 VSS 0.018232f
C4178 DVSS.n4284 VSS 0.018232f
C4179 DVSS.n4285 VSS 0.052908f
C4180 DVSS.n4286 VSS 0.052908f
C4181 DVSS.n4287 VSS 0.018232f
C4182 DVSS.n4289 VSS 0.018232f
C4183 DVSS.n4290 VSS 0.052908f
C4184 DVSS.n4291 VSS 0.052908f
C4185 DVSS.n4292 VSS 0.018232f
C4186 DVSS.n4294 VSS 0.018232f
C4187 DVSS.n4295 VSS 0.052908f
C4188 DVSS.n4296 VSS 0.052908f
C4189 DVSS.n4297 VSS 0.018232f
C4190 DVSS.n4299 VSS 0.018232f
C4191 DVSS.n4300 VSS 0.052908f
C4192 DVSS.n4301 VSS 0.048819f
C4193 DVSS.n4302 VSS 0.018232f
C4194 DVSS.n4304 VSS 0.018232f
C4195 DVSS.n4305 VSS 0.015532f
C4196 DVSS.n4306 VSS 0.016265f
C4197 DVSS.n4307 VSS 0.018232f
C4198 DVSS.n4309 VSS 0.018232f
C4199 DVSS.n4310 VSS 0.016265f
C4200 DVSS.n4312 VSS 0.018232f
C4201 DVSS.n4313 VSS 0.013769f
C4202 DVSS.n4314 VSS 0.013858f
C4203 DVSS.n4315 VSS 0.009015f
C4204 DVSS.n4316 VSS 0.016313f
C4205 DVSS.n4318 VSS 4.03086f
C4206 DVSS.n4320 VSS 0.018232f
C4207 DVSS.n4322 VSS 0.018232f
C4208 DVSS.n4323 VSS 0.016265f
C4209 DVSS.n4324 VSS 0.013769f
C4210 DVSS.n4325 VSS 0.018232f
C4211 DVSS.n4327 VSS 0.009015f
C4212 DVSS.n4328 VSS 0.018232f
C4213 DVSS.n4329 VSS 0.015218f
C4214 DVSS.n4330 VSS 0.016313f
C4215 DVSS.n4331 VSS 0.014785f
C4216 DVSS.n4332 VSS 0.008222f
C4217 DVSS.n4333 VSS 0.012766f
C4218 DVSS.n4334 VSS 0.018232f
C4219 DVSS.n4335 VSS 0.016444f
C4220 DVSS.n4336 VSS 0.016444f
C4221 DVSS.n4337 VSS 0.018232f
C4222 DVSS.n4338 VSS 0.016444f
C4223 DVSS.n4339 VSS 0.016444f
C4224 DVSS.n4340 VSS 0.018232f
C4225 DVSS.n4341 VSS 0.016444f
C4226 DVSS.n4342 VSS 0.016444f
C4227 DVSS.n4343 VSS 0.018232f
C4228 DVSS.n4344 VSS 0.016444f
C4229 DVSS.n4345 VSS 0.016444f
C4230 DVSS.n4346 VSS 0.018232f
C4231 DVSS.n4347 VSS 0.016444f
C4232 DVSS.n4348 VSS 0.016444f
C4233 DVSS.n4349 VSS 0.018232f
C4234 DVSS.n4350 VSS 0.016444f
C4235 DVSS.n4351 VSS 0.016444f
C4236 DVSS.n4352 VSS 0.018232f
C4237 DVSS.n4353 VSS 0.016444f
C4238 DVSS.n4354 VSS 0.016444f
C4239 DVSS.n4355 VSS 0.018232f
C4240 DVSS.n4356 VSS 0.016444f
C4241 DVSS.n4357 VSS 0.016444f
C4242 DVSS.n4358 VSS 0.016444f
C4243 DVSS.n4359 VSS 0.016444f
C4244 DVSS.n4360 VSS 0.016444f
C4245 DVSS.n4361 VSS 0.018232f
C4246 DVSS.n4362 VSS 0.018232f
C4247 DVSS.t0 VSS 0.519282f
C4248 DVSS.n4363 VSS 0.98199f
C4249 DVSS.t1 VSS 0.519282f
C4250 DVSS.n4364 VSS 0.98199f
C4251 DVSS.n4365 VSS 0.807931f
C4252 DVSS.n4366 VSS 0.029304f
C4253 DVSS.n4367 VSS 0.031816f
C4254 DVSS.n4368 VSS 0.018232f
C4255 DVSS.n4369 VSS 0.039351f
C4256 DVSS.n4370 VSS 0.063632f
C4257 DVSS.n4371 VSS 0.063632f
C4258 DVSS.n4372 VSS 0.018232f
C4259 DVSS.n4373 VSS 1.13742f
C4260 DVSS.n4374 VSS 0.018232f
C4261 DVSS.n4375 VSS 0.016444f
C4262 DVSS.n4376 VSS 0.016444f
C4263 DVSS.n4377 VSS 0.016444f
C4264 DVSS.n4378 VSS 0.018232f
C4265 DVSS.n4379 VSS 1.13742f
C4266 DVSS.n4380 VSS 0.018232f
C4267 DVSS.n4381 VSS 0.063632f
C4268 DVSS.n4382 VSS 0.063632f
C4269 DVSS.n4383 VSS 0.063632f
C4270 DVSS.n4384 VSS 0.018232f
C4271 DVSS.n4385 VSS 1.13742f
C4272 DVSS.n4386 VSS 0.018232f
C4273 DVSS.n4387 VSS 0.016444f
C4274 DVSS.n4388 VSS 0.016444f
C4275 DVSS.n4389 VSS 0.016444f
C4276 DVSS.n4390 VSS 0.018232f
C4277 DVSS.n4391 VSS 1.13742f
C4278 DVSS.n4392 VSS 0.018232f
C4279 DVSS.n4393 VSS 0.063632f
C4280 DVSS.n4394 VSS 0.048561f
C4281 DVSS.n4395 VSS 0.046887f
C4282 DVSS.n4396 VSS 0.018232f
C4283 DVSS.n4397 VSS 1.13742f
C4284 DVSS.n4398 VSS 0.018232f
C4285 DVSS.n4399 VSS 0.016444f
C4286 DVSS.n4400 VSS 0.016444f
C4287 DVSS.n4401 VSS 0.016444f
C4288 DVSS.n4402 VSS 0.018232f
C4289 DVSS.n4403 VSS 1.13742f
C4290 DVSS.n4404 VSS 0.018232f
C4291 DVSS.n4405 VSS 0.063632f
C4292 DVSS.n4406 VSS 0.063632f
C4293 DVSS.n4407 VSS 0.063632f
C4294 DVSS.n4408 VSS 0.018232f
C4295 DVSS.n4409 VSS 1.13742f
C4296 DVSS.n4410 VSS 0.018232f
C4297 DVSS.n4411 VSS 0.016444f
C4298 DVSS.n4412 VSS 0.016444f
C4299 DVSS.n4413 VSS 0.016444f
C4300 DVSS.n4414 VSS 0.018232f
C4301 DVSS.n4415 VSS 1.13742f
C4302 DVSS.n4416 VSS 0.018232f
C4303 DVSS.n4417 VSS 0.063632f
C4304 DVSS.n4418 VSS 0.063632f
C4305 DVSS.n4419 VSS 0.063632f
C4306 DVSS.n4420 VSS 0.018232f
C4307 DVSS.n4421 VSS 1.13742f
C4308 DVSS.n4422 VSS 0.018232f
C4309 DVSS.n4423 VSS 0.016444f
C4310 DVSS.n4424 VSS 0.016444f
C4311 DVSS.n4425 VSS 0.012766f
C4312 DVSS.n4426 VSS 0.018232f
C4313 DVSS.n4427 VSS 1.13742f
C4314 DVSS.n4428 VSS 0.018232f
C4315 DVSS.n4429 VSS 0.049398f
C4316 DVSS.n4430 VSS 0.031816f
C4317 DVSS.n4431 VSS 0.49201f
C4318 DVSS.n4432 VSS 1.15448f
C4319 DVSS.n4433 VSS 7.240029f
C4320 DVSS.n4434 VSS 0.019442f
C4321 DVSS.n4435 VSS 0.019442f
C4322 DVSS.n4436 VSS 0.019442f
C4323 DVSS.n4437 VSS 0.019442f
C4324 DVSS.n4438 VSS 0.019442f
C4325 DVSS.n4439 VSS 0.019442f
C4326 DVSS.n4440 VSS 0.019442f
C4327 DVSS.n4441 VSS 0.019442f
C4328 DVSS.n4442 VSS 0.019442f
C4329 DVSS.n4443 VSS 0.019442f
C4330 DVSS.n4444 VSS 0.009721f
C4331 DVSS.n4445 VSS 4.96014f
C4332 DVSS.n4446 VSS 0.009721f
C4333 DVSS.n4447 VSS 0.031907f
C4334 DVSS.n4448 VSS 0.166982f
C4335 DVSS.n4449 VSS 0.269288f
C4336 DVSS.n4450 VSS 0.333965f
C4337 DVSS.n4451 VSS 0.333965f
C4338 DVSS.n4452 VSS 0.333965f
C4339 DVSS.n4453 VSS 0.333965f
C4340 DVSS.n4454 VSS 0.333965f
C4341 DVSS.n4455 VSS 0.333965f
C4342 DVSS.n4456 VSS 0.333965f
C4343 DVSS.n4457 VSS 0.333965f
C4344 DVSS.n4458 VSS 0.333965f
C4345 DVSS.n4459 VSS 0.333965f
C4346 DVSS.n4460 VSS 0.333965f
C4347 DVSS.n4461 VSS 0.333965f
C4348 DVSS.n4462 VSS 0.333965f
C4349 DVSS.n4463 VSS 0.333965f
C4350 DVSS.n4464 VSS 0.333965f
C4351 DVSS.n4465 VSS 0.333965f
C4352 DVSS.n4466 VSS 0.333965f
C4353 DVSS.n4467 VSS 0.333965f
C4354 DVSS.n4468 VSS 0.333965f
C4355 DVSS.n4469 VSS 0.333965f
C4356 DVSS.n4470 VSS 0.333965f
C4357 DVSS.n4471 VSS 0.333965f
C4358 DVSS.n4472 VSS 0.333965f
C4359 DVSS.n4473 VSS 0.333965f
C4360 DVSS.n4474 VSS 0.333965f
C4361 DVSS.n4475 VSS 0.333965f
C4362 DVSS.n4476 VSS 0.333965f
C4363 DVSS.n4477 VSS 0.333965f
C4364 DVSS.n4478 VSS 0.333965f
C4365 DVSS.n4479 VSS 0.333965f
C4366 DVSS.n4480 VSS 0.333965f
C4367 DVSS.n4481 VSS 0.333965f
C4368 DVSS.n4482 VSS 0.333965f
C4369 DVSS.n4483 VSS 0.333965f
C4370 DVSS.n4484 VSS 0.333965f
C4371 DVSS.n4485 VSS 0.333965f
C4372 DVSS.n4486 VSS 0.333965f
C4373 DVSS.n4487 VSS 0.333965f
C4374 DVSS.n4488 VSS 0.333965f
C4375 DVSS.n4489 VSS 0.333965f
C4376 DVSS.n4490 VSS 0.333965f
C4377 DVSS.n4491 VSS 0.333965f
C4378 DVSS.n4492 VSS 0.333965f
C4379 DVSS.n4493 VSS 0.333965f
C4380 DVSS.n4494 VSS 0.333965f
C4381 DVSS.n4495 VSS 0.333965f
C4382 DVSS.n4496 VSS 0.333965f
C4383 DVSS.n4497 VSS 0.333965f
C4384 DVSS.n4498 VSS 0.333965f
C4385 DVSS.n4499 VSS 0.333965f
C4386 DVSS.n4500 VSS 0.333965f
C4387 DVSS.n4501 VSS 0.166982f
C4388 DVSS.n4502 VSS 0.333965f
C4389 DVSS.n4503 VSS 0.333965f
C4390 DVSS.n4504 VSS 0.333965f
C4391 DVSS.n4505 VSS 0.333965f
C4392 DVSS.n4507 VSS 0.052105f
C4393 DVSS.n4508 VSS 0.052105f
C4394 DVSS.n4509 VSS 0.052105f
C4395 DVSS.n4510 VSS 0.052105f
C4396 DVSS.n4511 VSS 0.052105f
C4397 DVSS.n4512 VSS 0.052105f
C4398 DVSS.n4513 VSS 0.052105f
C4399 DVSS.n4514 VSS 0.052105f
C4400 DVSS.n4515 VSS 0.052105f
C4401 DVSS.n4516 VSS 0.052105f
C4402 DVSS.n4518 VSS 0.052105f
C4403 DVSS.n4520 VSS 0.052105f
C4404 DVSS.n4522 VSS 0.052105f
C4405 DVSS.n4524 VSS 0.052105f
C4406 DVSS.n4526 VSS 0.052105f
C4407 DVSS.n4528 VSS 0.052105f
C4408 DVSS.n4530 VSS 0.052105f
C4409 DVSS.n4532 VSS 0.052105f
C4410 DVSS.n4534 VSS 0.052105f
C4411 DVSS.n4536 VSS 0.052105f
C4412 DVSS.n4549 VSS 0.154047f
C4413 DVSS.n4550 VSS 0.145816f
C4414 DVSS.n4551 VSS 0.333965f
C4415 DVSS.n4552 VSS 0.333965f
C4416 DVSS.n4553 VSS 0.333965f
C4417 DVSS.n4554 VSS 0.333965f
C4418 DVSS.n4555 VSS 0.333965f
C4419 DVSS.n4556 VSS 0.333965f
C4420 DVSS.n4557 VSS 0.333965f
C4421 DVSS.n4558 VSS 0.333965f
C4422 DVSS.n4559 VSS 0.333965f
C4423 DVSS.n4560 VSS 0.333965f
C4424 DVSS.n4561 VSS 0.333965f
C4425 DVSS.n4562 VSS 0.333965f
C4426 DVSS.n4563 VSS 0.333965f
C4427 DVSS.n4564 VSS 0.333965f
C4428 DVSS.n4565 VSS 0.333965f
C4429 DVSS.n4566 VSS 0.333965f
C4430 DVSS.n4567 VSS 0.333965f
C4431 DVSS.n4568 VSS 0.333965f
C4432 DVSS.n4569 VSS 0.333965f
C4433 DVSS.n4570 VSS 0.333965f
C4434 DVSS.n4571 VSS 0.333965f
C4435 DVSS.n4572 VSS 0.333965f
C4436 DVSS.n4573 VSS 0.333965f
C4437 DVSS.n4574 VSS 0.333965f
C4438 DVSS.n4575 VSS 0.333965f
C4439 DVSS.n4576 VSS 0.333965f
C4440 DVSS.n4577 VSS 0.333965f
C4441 DVSS.n4578 VSS 0.333965f
C4442 DVSS.n4579 VSS 0.333965f
C4443 DVSS.n4580 VSS 0.333965f
C4444 DVSS.n4581 VSS 0.333965f
C4445 DVSS.n4582 VSS 0.333965f
C4446 DVSS.n4583 VSS 0.333965f
C4447 DVSS.n4584 VSS 0.333965f
C4448 DVSS.n4585 VSS 0.333965f
C4449 DVSS.n4586 VSS 0.333965f
C4450 DVSS.n4587 VSS 0.333965f
C4451 DVSS.n4588 VSS 0.333965f
C4452 DVSS.n4589 VSS 0.333965f
C4453 DVSS.n4590 VSS 0.333965f
C4454 DVSS.n4591 VSS 0.333965f
C4455 DVSS.n4592 VSS 0.333965f
C4456 DVSS.n4593 VSS 0.196381f
C4457 DVSS.n4594 VSS 0.166982f
C4458 DVSS.n4595 VSS 0.052105f
C4459 DVSS.n4596 VSS 0.158751f
C4460 DVSS.n4597 VSS 0.145816f
C4461 DVSS.n4598 VSS 0.333965f
C4462 DVSS.n4599 VSS 0.333965f
C4463 DVSS.n4600 VSS 0.201084f
C4464 DVSS.n4601 VSS 0.333965f
C4465 DVSS.n4602 VSS 0.333965f
C4466 DVSS.n4603 VSS 0.333965f
C4467 DVSS.n4604 VSS 0.333965f
C4468 DVSS.n4605 VSS 0.333965f
C4469 DVSS.n4606 VSS 0.333965f
C4470 DVSS.n4607 VSS 0.333965f
C4471 DVSS.n4608 VSS 0.333965f
C4472 DVSS.n4609 VSS 0.333965f
C4473 DVSS.n4610 VSS 0.333965f
C4474 DVSS.n4611 VSS 0.333965f
C4475 DVSS.n4612 VSS 0.333965f
C4476 DVSS.n4613 VSS 0.333965f
C4477 DVSS.n4614 VSS 0.333965f
C4478 DVSS.n4615 VSS 0.333965f
C4479 DVSS.n4616 VSS 0.333965f
C4480 DVSS.n4617 VSS 0.333965f
C4481 DVSS.n4618 VSS 0.333965f
C4482 DVSS.n4619 VSS 0.333965f
C4483 DVSS.n4620 VSS 0.333965f
C4484 DVSS.n4621 VSS 0.333965f
C4485 DVSS.n4622 VSS 0.333965f
C4486 DVSS.n4623 VSS 0.333965f
C4487 DVSS.n4624 VSS 0.333965f
C4488 DVSS.n4625 VSS 0.201084f
C4489 DVSS.n4626 VSS 0.019442f
C4490 DVSS.n4627 VSS 0.019442f
C4491 DVSS.n4628 VSS 0.019442f
C4492 DVSS.n4629 VSS 0.019442f
C4493 DVSS.n4630 VSS 0.019442f
C4494 DVSS.n4631 VSS 0.019442f
C4495 DVSS.n4632 VSS 0.019442f
C4496 DVSS.n4633 VSS 0.019442f
C4497 DVSS.n4634 VSS 0.019442f
C4498 DVSS.n4635 VSS 0.019442f
C4499 DVSS.n4636 VSS 0.166982f
C4500 DVSS.n4637 VSS 0.009721f
C4501 DVSS.n4638 VSS 0.031907f
C4502 DVSS.n4639 VSS 0.166982f
C4503 DVSS.n4640 VSS 0.241458f
C4504 DVSS.n4641 VSS 0.397386f
C4505 DVSS.n4642 VSS 0.166878f
C4506 DVSS.n4643 VSS 0.009721f
C4507 DVSS.n4644 VSS 0.016385f
C4508 DVSS.n4645 VSS 0.077925f
C4509 DVSS.n4646 VSS 0.093839f
C4510 DVSS.n4647 VSS 0.15585f
C4511 DVSS.n4648 VSS 0.15585f
C4512 DVSS.n4649 VSS 0.15585f
C4513 DVSS.n4650 VSS 0.15585f
C4514 DVSS.n4651 VSS 0.15585f
C4515 DVSS.n4652 VSS 0.149814f
C4516 DVSS.n4653 VSS 0.15585f
C4517 DVSS.n4654 VSS 0.15585f
C4518 DVSS.n4655 VSS 0.15585f
C4519 DVSS.n4656 VSS 0.15585f
C4520 DVSS.n4657 VSS 0.15585f
C4521 DVSS.n4658 VSS 0.15585f
C4522 DVSS.n4659 VSS 0.15585f
C4523 DVSS.n4660 VSS 0.15585f
C4524 DVSS.n4661 VSS 0.15585f
C4525 DVSS.n4662 VSS 0.15585f
C4526 DVSS.n4663 VSS 0.15585f
C4527 DVSS.n4664 VSS 0.15585f
C4528 DVSS.n4665 VSS 0.15585f
C4529 DVSS.n4666 VSS 0.15585f
C4530 DVSS.n4667 VSS 0.15585f
C4531 DVSS.n4668 VSS 0.15585f
C4532 DVSS.n4669 VSS 0.15585f
C4533 DVSS.n4670 VSS 0.15585f
C4534 DVSS.n4671 VSS 0.15585f
C4535 DVSS.n4672 VSS 0.15585f
C4536 DVSS.n4673 VSS 0.15585f
C4537 DVSS.n4674 VSS 0.15585f
C4538 DVSS.n4675 VSS 0.15585f
C4539 DVSS.n4676 VSS 0.15585f
C4540 DVSS.n4677 VSS 0.15585f
C4541 DVSS.n4678 VSS 0.093839f
C4542 DVSS.n4679 VSS 0.15585f
C4543 DVSS.n4680 VSS 0.15585f
C4544 DVSS.n4681 VSS 0.15585f
C4545 DVSS.n4682 VSS 0.15585f
C4546 DVSS.n4683 VSS 0.15585f
C4547 DVSS.n4684 VSS 0.15585f
C4548 DVSS.n4685 VSS 0.15585f
C4549 DVSS.n4686 VSS 0.15585f
C4550 DVSS.n4687 VSS 0.15585f
C4551 DVSS.n4688 VSS 0.15585f
C4552 DVSS.n4689 VSS 0.15585f
C4553 DVSS.n4690 VSS 0.15585f
C4554 DVSS.n4691 VSS 0.15585f
C4555 DVSS.n4692 VSS 0.15585f
C4556 DVSS.n4693 VSS 0.15585f
C4557 DVSS.n4694 VSS 0.15585f
C4558 DVSS.n4695 VSS 0.15585f
C4559 DVSS.n4696 VSS 0.15585f
C4560 DVSS.n4697 VSS 0.15585f
C4561 DVSS.n4698 VSS 0.019442f
C4562 DVSS.n4699 VSS 0.019442f
C4563 DVSS.n4700 VSS 0.019442f
C4564 DVSS.n4701 VSS 0.019442f
C4565 DVSS.n4702 VSS 0.016385f
C4566 DVSS.n4703 VSS 0.077925f
C4567 DVSS.n4704 VSS 0.15585f
C4568 DVSS.n4705 VSS 0.15585f
C4569 DVSS.n4706 VSS 0.152009f
C4570 DVSS.n4707 VSS 0.15585f
C4571 DVSS.n4708 VSS 0.15585f
C4572 DVSS.n4709 VSS 0.15585f
C4573 DVSS.n4710 VSS 0.15585f
C4574 DVSS.n4711 VSS 0.15585f
C4575 DVSS.n4712 VSS 0.15585f
C4576 DVSS.n4713 VSS 0.15585f
C4577 DVSS.n4714 VSS 0.15585f
C4578 DVSS.n4715 VSS 0.15585f
C4579 DVSS.n4716 VSS 0.15585f
C4580 DVSS.n4717 VSS 0.15585f
C4581 DVSS.n4718 VSS 0.15585f
C4582 DVSS.n4719 VSS 0.15585f
C4583 DVSS.n4720 VSS 0.15585f
C4584 DVSS.n4721 VSS 0.15585f
C4585 DVSS.n4722 VSS 0.15585f
C4586 DVSS.n4723 VSS 0.15585f
C4587 DVSS.n4724 VSS 0.15585f
C4588 DVSS.n4725 VSS 0.15585f
C4589 DVSS.n4726 VSS 0.15585f
C4590 DVSS.n4727 VSS 0.15585f
C4591 DVSS.n4728 VSS 0.15585f
C4592 DVSS.n4729 VSS 0.15585f
C4593 DVSS.n4730 VSS 0.15585f
C4594 DVSS.n4731 VSS 0.15585f
C4595 DVSS.n4732 VSS 0.15585f
C4596 DVSS.n4733 VSS 0.15585f
C4597 DVSS.n4734 VSS 0.15585f
C4598 DVSS.n4735 VSS 0.15585f
C4599 DVSS.n4736 VSS 0.15585f
C4600 DVSS.n4737 VSS 0.15585f
C4601 DVSS.n4738 VSS 0.15585f
C4602 DVSS.n4739 VSS 0.068047f
C4603 DVSS.n4740 VSS 0.074084f
C4604 DVSS.n4741 VSS 0.052105f
C4605 DVSS.n4742 VSS 0.077925f
C4606 DVSS.n4743 VSS 0.043911f
C4607 DVSS.n4744 VSS 0.25307f
C4608 DVSS.n4745 VSS 0.103826f
C4609 DVSS.n4746 VSS 0.484326f
C4610 DVSS.n4747 VSS 1.065f
C4611 DVSS.n4748 VSS 0.008222f
C4612 DVSS.n4749 VSS 0.012333f
C4613 DVSS.n4750 VSS 0.018232f
C4614 DVSS.n4751 VSS 1.13742f
C4615 DVSS.n4752 VSS 0.018232f
C4616 DVSS.n4753 VSS 0.018232f
C4617 DVSS.n4754 VSS 0.012333f
C4618 DVSS.n4755 VSS 0.016444f
C4619 DVSS.n4756 VSS 0.018232f
C4620 DVSS.n4757 VSS 0.016444f
C4621 DVSS.n4758 VSS 0.016444f
C4622 DVSS.n4759 VSS 0.018232f
C4623 DVSS.n4760 VSS 0.016444f
C4624 DVSS.n4761 VSS 0.016444f
C4625 DVSS.n4762 VSS 0.018232f
C4626 DVSS.n4763 VSS 0.016444f
C4627 DVSS.n4764 VSS 0.016444f
C4628 DVSS.n4765 VSS 0.018232f
C4629 DVSS.n4766 VSS 0.016444f
C4630 DVSS.n4767 VSS 0.016444f
C4631 DVSS.n4768 VSS 0.018232f
C4632 DVSS.n4769 VSS 0.016444f
C4633 DVSS.n4770 VSS 0.016444f
C4634 DVSS.n4771 VSS 0.018232f
C4635 DVSS.n4772 VSS 0.016444f
C4636 DVSS.n4773 VSS 0.016444f
C4637 DVSS.n4774 VSS 0.018232f
C4638 DVSS.n4775 VSS 0.016444f
C4639 DVSS.n4776 VSS 0.016444f
C4640 DVSS.n4777 VSS 0.018232f
C4641 DVSS.n4778 VSS 0.016444f
C4642 DVSS.n4779 VSS 0.016444f
C4643 DVSS.n4780 VSS 0.016444f
C4644 DVSS.n4781 VSS 0.016444f
C4645 DVSS.n4782 VSS 0.016444f
C4646 DVSS.n4783 VSS 0.018232f
C4647 DVSS.n4784 VSS 0.018232f
C4648 DVSS.t8 VSS 0.519282f
C4649 DVSS.n4785 VSS 0.98199f
C4650 DVSS.t5 VSS 0.519282f
C4651 DVSS.n4786 VSS 0.98199f
C4652 DVSS.n4787 VSS 0.02763f
C4653 DVSS.n4788 VSS 0.807931f
C4654 DVSS.n4789 VSS 0.060283f
C4655 DVSS.n4790 VSS 0.063632f
C4656 DVSS.n4791 VSS 0.018232f
C4657 DVSS.n4792 VSS 1.13742f
C4658 DVSS.n4793 VSS 0.018232f
C4659 DVSS.n4794 VSS 0.016444f
C4660 DVSS.n4795 VSS 0.016444f
C4661 DVSS.n4796 VSS 0.016444f
C4662 DVSS.n4797 VSS 0.018232f
C4663 DVSS.n4798 VSS 1.13742f
C4664 DVSS.n4799 VSS 0.018232f
C4665 DVSS.n4800 VSS 0.063632f
C4666 DVSS.n4801 VSS 0.063632f
C4667 DVSS.n4802 VSS 0.063632f
C4668 DVSS.n4803 VSS 0.018232f
C4669 DVSS.n4804 VSS 1.13742f
C4670 DVSS.n4805 VSS 0.018232f
C4671 DVSS.n4806 VSS 0.016444f
C4672 DVSS.n4807 VSS 0.016444f
C4673 DVSS.n4808 VSS 0.016444f
C4674 DVSS.n4809 VSS 0.018232f
C4675 DVSS.n4810 VSS 1.13742f
C4676 DVSS.n4811 VSS 0.018232f
C4677 DVSS.n4812 VSS 0.063632f
C4678 DVSS.n4813 VSS 0.063632f
C4679 DVSS.n4814 VSS 0.056934f
C4680 DVSS.n4815 VSS 0.018232f
C4681 DVSS.n4816 VSS 1.13742f
C4682 DVSS.n4817 VSS 0.018232f
C4683 DVSS.n4818 VSS 0.016444f
C4684 DVSS.n4819 VSS 0.016444f
C4685 DVSS.n4820 VSS 0.016444f
C4686 DVSS.n4821 VSS 0.018232f
C4687 DVSS.n4822 VSS 1.13742f
C4688 DVSS.n4823 VSS 0.018232f
C4689 DVSS.n4824 VSS 0.063632f
C4690 DVSS.n4825 VSS 0.063632f
C4691 DVSS.n4826 VSS 0.063632f
C4692 DVSS.n4827 VSS 0.018232f
C4693 DVSS.n4828 VSS 1.13742f
C4694 DVSS.n4829 VSS 0.018232f
C4695 DVSS.n4830 VSS 0.016444f
C4696 DVSS.n4831 VSS 0.016444f
C4697 DVSS.n4832 VSS 0.016444f
C4698 DVSS.n4833 VSS 0.018232f
C4699 DVSS.n4834 VSS 1.13742f
C4700 DVSS.n4835 VSS 0.018232f
C4701 DVSS.n4836 VSS 0.063632f
C4702 DVSS.n4837 VSS 0.063632f
C4703 DVSS.n4838 VSS 0.063632f
C4704 DVSS.n4839 VSS 0.018232f
C4705 DVSS.n4840 VSS 1.13742f
C4706 DVSS.n4841 VSS 0.018232f
C4707 DVSS.n4842 VSS 0.016444f
C4708 DVSS.n4843 VSS 0.016444f
C4709 DVSS.n4844 VSS 0.016444f
C4710 DVSS.n4845 VSS 0.018232f
C4711 DVSS.n4846 VSS 1.13742f
C4712 DVSS.n4847 VSS 0.018232f
C4713 DVSS.n4848 VSS 0.034607f
C4714 DVSS.n4849 VSS 0.031816f
C4715 DVSS.n4850 VSS 0.026052f
C4716 DVSS.n4851 VSS 0.031816f
C4717 DVSS.n4852 VSS 0.059446f
C4718 DVSS.n4853 VSS 0.063632f
C4719 DVSS.n4854 VSS 0.018232f
C4720 DVSS.n4855 VSS 1.13742f
C4721 DVSS.n4856 VSS 0.018232f
C4722 DVSS.n4857 VSS 0.016444f
C4723 DVSS.n4858 VSS 0.016444f
C4724 DVSS.n4859 VSS 0.016444f
C4725 DVSS.n4860 VSS 0.018232f
C4726 DVSS.n4861 VSS 1.13742f
C4727 DVSS.n4862 VSS 0.018232f
C4728 DVSS.n4863 VSS 0.063632f
C4729 DVSS.n4864 VSS 0.063632f
C4730 DVSS.n4865 VSS 0.063632f
C4731 DVSS.n4866 VSS 0.018232f
C4732 DVSS.n4867 VSS 1.13742f
C4733 DVSS.n4868 VSS 0.018232f
C4734 DVSS.n4869 VSS 0.016444f
C4735 DVSS.n4870 VSS 0.016444f
C4736 DVSS.n4871 VSS 0.016444f
C4737 DVSS.n4872 VSS 0.018232f
C4738 DVSS.n4873 VSS 1.13742f
C4739 DVSS.n4874 VSS 0.018232f
C4740 DVSS.n4875 VSS 0.063632f
C4741 DVSS.n4876 VSS 0.03684f
C4742 DVSS.n4877 VSS 0.058608f
C4743 DVSS.n4878 VSS 0.018232f
C4744 DVSS.n4879 VSS 1.13742f
C4745 DVSS.n4880 VSS 0.018232f
C4746 DVSS.n4881 VSS 0.016444f
C4747 DVSS.n4882 VSS 0.016444f
C4748 DVSS.n4883 VSS 0.016444f
C4749 DVSS.n4884 VSS 0.018232f
C4750 DVSS.n4885 VSS 1.13742f
C4751 DVSS.n4886 VSS 0.018232f
C4752 DVSS.n4887 VSS 0.063632f
C4753 DVSS.n4888 VSS 0.063632f
C4754 DVSS.n4889 VSS 0.063632f
C4755 DVSS.n4890 VSS 0.018232f
C4756 DVSS.n4891 VSS 1.13742f
C4757 DVSS.n4892 VSS 0.018232f
C4758 DVSS.n4893 VSS 0.016444f
C4759 DVSS.n4894 VSS 0.016444f
C4760 DVSS.n4895 VSS 0.016444f
C4761 DVSS.n4896 VSS 0.018232f
C4762 DVSS.n4897 VSS 1.13742f
C4763 DVSS.n4898 VSS 0.018232f
C4764 DVSS.n4899 VSS 0.063632f
C4765 DVSS.n4900 VSS 0.063632f
C4766 DVSS.n4901 VSS 0.063632f
C4767 DVSS.n4902 VSS 0.018232f
C4768 DVSS.n4903 VSS 1.13742f
C4769 DVSS.n4904 VSS 0.018232f
C4770 DVSS.n4905 VSS 0.016444f
C4771 DVSS.n4906 VSS 0.016444f
C4772 DVSS.n4907 VSS 0.014497f
C4773 DVSS.n4908 VSS 0.018232f
C4774 DVSS.n4909 VSS 1.13742f
C4775 DVSS.n4910 VSS 0.018232f
C4776 DVSS.n4911 VSS 0.014497f
C4777 DVSS.n4912 VSS 0.008222f
C4778 DVSS.n4913 VSS 0.63273f
C4779 DVSS.n4914 VSS 0.172627f
C4780 DVSS.n4915 VSS 0.009721f
C4781 DVSS.n4916 VSS 0.019442f
C4782 DVSS.n4917 VSS 0.019442f
C4783 DVSS.n4918 VSS 0.019442f
C4784 DVSS.n4919 VSS 0.019442f
C4785 DVSS.n4920 VSS 0.019442f
C4786 DVSS.n4921 VSS 0.019442f
C4787 DVSS.n4922 VSS 0.019442f
C4788 DVSS.n4923 VSS 0.019442f
C4789 DVSS.n4924 VSS 0.009721f
C4790 DVSS.n4925 VSS 0.163376f
C4791 DVSS.n4926 VSS 0.163376f
C4792 DVSS.n4928 VSS 0.016071f
C4793 DVSS.n4929 VSS 0.325311f
C4794 DVSS.n4930 VSS 0.048557f
C4795 DVSS.n4931 VSS 0.327848f
C4796 DVSS.n4932 VSS 0.210696f
C4797 DVSS.n4933 VSS 0.183412f
C4798 DVSS.n4934 VSS 0.009721f
C4799 DVSS.n4935 VSS 0.009721f
C4800 DVSS.n4936 VSS 0.009721f
C4801 DVSS.n4937 VSS 0.013092f
C4802 DVSS.n4938 VSS 0.009721f
C4803 DVSS.n4939 VSS 0.019442f
C4804 DVSS.n4940 VSS 0.019442f
C4805 DVSS.n4941 VSS 0.019442f
C4806 DVSS.n4942 VSS 0.009721f
C4807 DVSS.n4943 VSS 0.010348f
C4808 DVSS.n4944 VSS 0.009721f
C4809 DVSS.n4945 VSS 0.355784f
C4810 DVSS.n4946 VSS 0.054406f
C4811 DVSS.n4947 VSS 0.0635f
C4812 DVSS.n4948 VSS 0.009721f
C4813 DVSS.n4949 VSS 0.355784f
C4814 DVSS.n4950 VSS 0.0635f
C4815 DVSS.n4951 VSS 0.0635f
C4816 DVSS.n4952 VSS 0.264848f
C4817 DVSS.n4953 VSS 0.327848f
C4818 DVSS.n4954 VSS 0.210696f
C4819 DVSS.n4955 VSS 0.481904f
C4820 DVSS.n4956 VSS 6.896141f
C4821 DVSS.n4957 VSS 0.051264f
C4822 DVSS.n4958 VSS 0.729894f
C4823 DVSS.n4959 VSS 0.729894f
C4824 DVSS.n4960 VSS 1.33324f
C4825 DVSS.n4961 VSS 0.018275f
C4826 DVSS.n4962 VSS 0.170181f
C4827 DVSS.n4963 VSS 0.027413f
C4828 DVSS.n4964 VSS 0.052105f
C4829 DVSS.n4965 VSS 0.355784f
C4830 DVSS.n4966 VSS 0.355784f
C4831 DVSS.n4967 VSS 0.325311f
C4832 DVSS.n4968 VSS 0.0635f
C4833 DVSS.n4969 VSS 0.009721f
C4834 DVSS.n4970 VSS 0.264848f
C4835 DVSS.n4971 VSS 0.0635f
C4836 DVSS.n4972 VSS 0.0635f
C4837 DVSS.n4973 VSS 0.009721f
C4838 DVSS.n4974 VSS 0.009721f
C4839 DVSS.n4975 VSS 0.264848f
C4840 DVSS.n4976 VSS 0.327848f
C4841 DVSS.n4977 VSS 0.210696f
C4842 DVSS.n4978 VSS 0.481904f
C4843 DVSS.n4979 VSS 6.896141f
C4844 DVSS.n4980 VSS 0.481904f
C4845 DVSS.n4981 VSS 0.210696f
C4846 DVSS.n4982 VSS 0.327848f
C4847 DVSS.n4983 VSS 0.264848f
C4848 DVSS.n4984 VSS 0.009721f
C4849 DVSS.n4985 VSS 0.355784f
C4850 DVSS.n4986 VSS 0.355784f
C4851 DVSS.n4987 VSS 0.052105f
C4852 DVSS.n4989 VSS 0.027733f
C4853 DVSS.n4990 VSS 0.027413f
C4854 DVSS.n4991 VSS 0.026052f
C4855 DVSS.n4992 VSS 0.027413f
C4856 DVSS.n4994 VSS 0.026052f
C4857 DVSS.n4995 VSS 0.026052f
C4858 DVSS.n4996 VSS 0.071889f
C4859 DVSS.n4997 VSS 0.035087f
C4860 DVSS.n4998 VSS 0.026052f
C4861 DVSS.n5000 VSS 0.210064f
C4862 DVSS.n5001 VSS 0.026052f
C4863 DVSS.n5002 VSS 0.210064f
C4864 DVSS.n5004 VSS 0.210064f
C4865 DVSS.n5005 VSS 0.009721f
C4866 DVSS.n5006 VSS 0.009721f
C4867 DVSS.n5007 VSS 0.077925f
C4868 DVSS.n5008 VSS 0.152009f
C4869 DVSS.n5009 VSS 0.15585f
C4870 DVSS.n5010 VSS 0.15585f
C4871 DVSS.n5011 VSS 0.15585f
C4872 DVSS.n5012 VSS 0.15585f
C4873 DVSS.n5013 VSS 0.15585f
C4874 DVSS.n5014 VSS 0.091644f
C4875 DVSS.n5015 VSS 0.15585f
C4876 DVSS.n5016 VSS 0.15585f
C4877 DVSS.n5017 VSS 0.15585f
C4878 DVSS.n5018 VSS 0.15585f
C4879 DVSS.n5019 VSS 0.15585f
C4880 DVSS.n5020 VSS 0.15585f
C4881 DVSS.n5021 VSS 0.15585f
C4882 DVSS.n5022 VSS 0.15585f
C4883 DVSS.n5023 VSS 0.15585f
C4884 DVSS.n5024 VSS 0.15585f
C4885 DVSS.n5025 VSS 0.15585f
C4886 DVSS.n5026 VSS 0.15585f
C4887 DVSS.n5027 VSS 0.15585f
C4888 DVSS.n5028 VSS 0.15585f
C4889 DVSS.n5029 VSS 0.15585f
C4890 DVSS.n5030 VSS 0.15585f
C4891 DVSS.n5031 VSS 0.15585f
C4892 DVSS.n5032 VSS 0.15585f
C4893 DVSS.n5033 VSS 0.15585f
C4894 DVSS.n5034 VSS 0.15585f
C4895 DVSS.n5035 VSS 0.15585f
C4896 DVSS.n5036 VSS 0.15585f
C4897 DVSS.n5037 VSS 0.15585f
C4898 DVSS.n5038 VSS 0.15585f
C4899 DVSS.n5039 VSS 0.15585f
C4900 DVSS.n5040 VSS 0.15585f
C4901 DVSS.n5041 VSS 0.15585f
C4902 DVSS.n5042 VSS 0.15585f
C4903 DVSS.n5043 VSS 0.15585f
C4904 DVSS.n5044 VSS 0.15585f
C4905 DVSS.n5045 VSS 0.15585f
C4906 DVSS.n5046 VSS 0.11579f
C4907 DVSS.n5047 VSS 0.15585f
C4908 DVSS.n5048 VSS 0.15585f
C4909 DVSS.n5049 VSS 0.15585f
C4910 DVSS.n5050 VSS 0.15585f
C4911 DVSS.n5051 VSS 0.15585f
C4912 DVSS.n5052 VSS 0.15585f
C4913 DVSS.n5053 VSS 0.15585f
C4914 DVSS.n5054 VSS 0.15585f
C4915 DVSS.n5055 VSS 0.751144f
C4916 DVSS.n5056 VSS 0.205146f
C4917 DVSS.n5057 VSS 0.08012f
C4918 DVSS.n5058 VSS 0.15585f
C4919 DVSS.n5059 VSS 0.140485f
C4920 DVSS.n5060 VSS 0.140485f
C4921 DVSS.n5061 VSS 0.15585f
C4922 DVSS.n5062 VSS 0.15585f
C4923 DVSS.n5063 VSS 0.15585f
C4924 DVSS.n5064 VSS 0.15585f
C4925 DVSS.n5065 VSS 0.15585f
C4926 DVSS.n5066 VSS 0.15585f
C4927 DVSS.n5067 VSS 0.15585f
C4928 DVSS.n5068 VSS 0.15585f
C4929 DVSS.n5069 VSS 0.15585f
C4930 DVSS.n5070 VSS 0.15585f
C4931 DVSS.n5071 VSS 0.15585f
C4932 DVSS.n5072 VSS 0.15585f
C4933 DVSS.n5073 VSS 0.15585f
C4934 DVSS.n5074 VSS 0.15585f
C4935 DVSS.n5075 VSS 0.15585f
C4936 DVSS.n5076 VSS 0.15585f
C4937 DVSS.n5077 VSS 0.15585f
C4938 DVSS.n5078 VSS 0.15585f
C4939 DVSS.n5079 VSS 0.15585f
C4940 DVSS.n5080 VSS 0.15585f
C4941 DVSS.n5081 VSS 0.15585f
C4942 DVSS.n5082 VSS 0.15585f
C4943 DVSS.n5083 VSS 0.15585f
C4944 DVSS.n5084 VSS 0.068047f
C4945 DVSS.n5085 VSS 0.077925f
C4946 DVSS.n5086 VSS 0.163376f
C4947 DVSS.n5087 VSS 0.163376f
C4948 DVSS.n5088 VSS 0.077925f
C4949 DVSS.n5089 VSS 0.15585f
C4950 DVSS.n5090 VSS 0.15585f
C4951 DVSS.n5091 VSS 0.15585f
C4952 DVSS.n5092 VSS 0.11579f
C4953 DVSS.n5093 VSS 0.15585f
C4954 DVSS.n5094 VSS 0.15585f
C4955 DVSS.n5095 VSS 0.15585f
C4956 DVSS.n5096 VSS 0.15585f
C4957 DVSS.n5097 VSS 0.15585f
C4958 DVSS.n5098 VSS 0.15585f
C4959 DVSS.n5099 VSS 0.15585f
C4960 DVSS.n5100 VSS 0.15585f
C4961 DVSS.n5101 VSS 0.751144f
C4962 DVSS.n5102 VSS 0.205146f
C4963 DVSS.n5103 VSS 0.08012f
C4964 DVSS.n5104 VSS 0.15585f
C4965 DVSS.n5105 VSS 0.140485f
C4966 DVSS.n5106 VSS 0.140485f
C4967 DVSS.n5107 VSS 0.15585f
C4968 DVSS.n5108 VSS 0.15585f
C4969 DVSS.n5109 VSS 0.15585f
C4970 DVSS.n5110 VSS 0.15585f
C4971 DVSS.n5111 VSS 0.15585f
C4972 DVSS.n5112 VSS 0.15585f
C4973 DVSS.n5113 VSS 0.15585f
C4974 DVSS.n5114 VSS 0.15585f
C4975 DVSS.n5115 VSS 0.15585f
C4976 DVSS.n5116 VSS 0.15585f
C4977 DVSS.n5117 VSS 0.15585f
C4978 DVSS.n5118 VSS 0.15585f
C4979 DVSS.n5119 VSS 0.15585f
C4980 DVSS.n5120 VSS 0.15585f
C4981 DVSS.n5121 VSS 0.15585f
C4982 DVSS.n5122 VSS 0.15585f
C4983 DVSS.n5123 VSS 0.15585f
C4984 DVSS.n5124 VSS 0.15585f
C4985 DVSS.n5125 VSS 0.15585f
C4986 DVSS.n5126 VSS 0.15585f
C4987 DVSS.n5127 VSS 0.15585f
C4988 DVSS.n5128 VSS 0.15585f
C4989 DVSS.n5129 VSS 0.15585f
C4990 DVSS.n5130 VSS 0.068047f
C4991 DVSS.n5131 VSS 0.077925f
C4992 DVSS.n5132 VSS 0.127863f
C4993 DVSS.n5133 VSS 0.15585f
C4994 DVSS.n5134 VSS 0.15585f
C4995 DVSS.n5135 VSS 0.15585f
C4996 DVSS.n5136 VSS 0.15585f
C4997 DVSS.n5137 VSS 0.15585f
C4998 DVSS.n5138 VSS 0.15585f
C4999 DVSS.n5139 VSS 0.15585f
C5000 DVSS.n5140 VSS 0.15585f
C5001 DVSS.n5141 VSS 0.15585f
C5002 DVSS.n5142 VSS 0.15585f
C5003 DVSS.n5143 VSS 0.15585f
C5004 DVSS.n5144 VSS 0.15585f
C5005 DVSS.n5145 VSS 0.15585f
C5006 DVSS.n5146 VSS 0.15585f
C5007 DVSS.n5147 VSS 0.15585f
C5008 DVSS.n5148 VSS 0.15585f
C5009 DVSS.n5149 VSS 0.15585f
C5010 DVSS.n5150 VSS 0.15585f
C5011 DVSS.n5151 VSS 0.15585f
C5012 DVSS.n5152 VSS 0.15585f
C5013 DVSS.n5153 VSS 0.15585f
C5014 DVSS.n5154 VSS 0.15585f
C5015 DVSS.n5155 VSS 0.15585f
C5016 DVSS.n5156 VSS 0.15585f
C5017 DVSS.n5157 VSS 0.15585f
C5018 DVSS.n5158 VSS 0.15585f
C5019 DVSS.n5159 VSS 0.15585f
C5020 DVSS.n5160 VSS 0.15585f
C5021 DVSS.n5161 VSS 0.15585f
C5022 DVSS.n5162 VSS 0.15585f
C5023 DVSS.n5163 VSS 0.091644f
C5024 DVSS.n5164 VSS 0.077925f
C5025 DVSS.n5165 VSS 0.172627f
C5026 DVSS.n5166 VSS 0.031907f
C5027 DVSS.n5167 VSS 0.49201f
C5028 DVSS.n5168 VSS 0.63273f
C5029 DVSS.n5169 VSS 0.008222f
C5030 DVSS.n5170 VSS 0.01017f
C5031 DVSS.n5171 VSS 0.018232f
C5032 DVSS.n5172 VSS 0.016444f
C5033 DVSS.n5173 VSS 0.016444f
C5034 DVSS.n5174 VSS 0.018232f
C5035 DVSS.n5175 VSS 0.016444f
C5036 DVSS.n5176 VSS 0.016444f
C5037 DVSS.n5177 VSS 0.018232f
C5038 DVSS.n5178 VSS 0.016444f
C5039 DVSS.n5179 VSS 0.016444f
C5040 DVSS.n5180 VSS 0.018232f
C5041 DVSS.n5181 VSS 0.016444f
C5042 DVSS.n5182 VSS 0.016444f
C5043 DVSS.n5183 VSS 0.018232f
C5044 DVSS.n5184 VSS 0.016444f
C5045 DVSS.n5185 VSS 0.016444f
C5046 DVSS.n5186 VSS 0.018232f
C5047 DVSS.n5187 VSS 0.016444f
C5048 DVSS.n5188 VSS 0.016444f
C5049 DVSS.n5189 VSS 0.018232f
C5050 DVSS.n5190 VSS 0.016444f
C5051 DVSS.n5191 VSS 0.016444f
C5052 DVSS.n5192 VSS 0.018232f
C5053 DVSS.n5193 VSS 0.016444f
C5054 DVSS.n5194 VSS 0.016444f
C5055 DVSS.n5195 VSS 0.016444f
C5056 DVSS.n5196 VSS 0.016444f
C5057 DVSS.n5197 VSS 0.016444f
C5058 DVSS.n5198 VSS 0.018232f
C5059 DVSS.n5199 VSS 0.018232f
C5060 DVSS.n5200 VSS 0.016444f
C5061 DVSS.n5201 VSS 0.016444f
C5062 DVSS.n5202 VSS 0.018232f
C5063 DVSS.n5203 VSS 1.13742f
C5064 DVSS.n5204 VSS 0.018232f
C5065 DVSS.n5205 VSS 0.063632f
C5066 DVSS.n5206 VSS 0.063632f
C5067 DVSS.n5207 VSS 0.063632f
C5068 DVSS.n5208 VSS 0.018232f
C5069 DVSS.n5209 VSS 1.13742f
C5070 DVSS.n5210 VSS 0.018232f
C5071 DVSS.n5211 VSS 0.016444f
C5072 DVSS.n5212 VSS 0.016444f
C5073 DVSS.n5213 VSS 0.016444f
C5074 DVSS.n5214 VSS 0.018232f
C5075 DVSS.n5215 VSS 1.13742f
C5076 DVSS.n5216 VSS 0.018232f
C5077 DVSS.n5217 VSS 0.063632f
C5078 DVSS.n5218 VSS 0.063632f
C5079 DVSS.n5219 VSS 0.063632f
C5080 DVSS.n5220 VSS 0.018232f
C5081 DVSS.n5221 VSS 1.13742f
C5082 DVSS.n5222 VSS 0.018232f
C5083 DVSS.n5223 VSS 0.016444f
C5084 DVSS.n5224 VSS 0.016444f
C5085 DVSS.n5225 VSS 0.016444f
C5086 DVSS.n5226 VSS 0.018232f
C5087 DVSS.n5227 VSS 1.13742f
C5088 DVSS.n5228 VSS 0.018232f
C5089 DVSS.n5229 VSS 0.045212f
C5090 DVSS.n5230 VSS 0.050236f
C5091 DVSS.n5231 VSS 0.063632f
C5092 DVSS.n5232 VSS 0.018232f
C5093 DVSS.n5233 VSS 1.13742f
C5094 DVSS.n5234 VSS 0.018232f
C5095 DVSS.n5235 VSS 0.016444f
C5096 DVSS.n5236 VSS 0.016444f
C5097 DVSS.n5237 VSS 0.016444f
C5098 DVSS.n5238 VSS 0.018232f
C5099 DVSS.n5239 VSS 1.13742f
C5100 DVSS.n5240 VSS 0.018232f
C5101 DVSS.n5241 VSS 0.063632f
C5102 DVSS.n5242 VSS 0.063632f
C5103 DVSS.n5243 VSS 0.063632f
C5104 DVSS.n5244 VSS 0.018232f
C5105 DVSS.n5245 VSS 1.13742f
C5106 DVSS.n5246 VSS 0.018232f
C5107 DVSS.n5247 VSS 0.016444f
C5108 DVSS.n5248 VSS 0.016444f
C5109 DVSS.n5249 VSS 0.016444f
C5110 DVSS.n5250 VSS 0.018232f
C5111 DVSS.n5251 VSS 1.13742f
C5112 DVSS.n5252 VSS 0.018232f
C5113 DVSS.n5253 VSS 0.063632f
C5114 DVSS.n5254 VSS 0.063632f
C5115 DVSS.n5255 VSS 0.039351f
C5116 DVSS.n5256 VSS 0.018232f
C5117 DVSS.n5257 VSS 1.13742f
C5118 DVSS.n5258 VSS 0.018232f
C5119 DVSS.n5259 VSS 0.01017f
C5120 DVSS.n5260 VSS 0.008222f
C5121 DVSS.n5261 VSS 0.397386f
C5122 DVSS.n5262 VSS 0.241458f
C5123 DVSS.n5263 VSS 0.009721f
C5124 DVSS.n5264 VSS 0.145816f
C5125 DVSS.n5265 VSS 0.166982f
C5126 DVSS.n5266 VSS 0.325733f
C5127 DVSS.n5267 VSS 0.333965f
C5128 DVSS.n5268 VSS 0.333965f
C5129 DVSS.n5269 VSS 0.333965f
C5130 DVSS.n5270 VSS 0.333965f
C5131 DVSS.n5271 VSS 0.333965f
C5132 DVSS.n5272 VSS 0.196381f
C5133 DVSS.n5273 VSS 0.333965f
C5134 DVSS.n5274 VSS 0.333965f
C5135 DVSS.n5275 VSS 0.333965f
C5136 DVSS.n5276 VSS 0.333965f
C5137 DVSS.n5277 VSS 0.333965f
C5138 DVSS.n5278 VSS 0.333965f
C5139 DVSS.n5279 VSS 0.333965f
C5140 DVSS.n5280 VSS 0.333965f
C5141 DVSS.n5281 VSS 0.333965f
C5142 DVSS.n5282 VSS 0.333965f
C5143 DVSS.n5283 VSS 0.333965f
C5144 DVSS.n5284 VSS 0.333965f
C5145 DVSS.n5285 VSS 0.333965f
C5146 DVSS.n5286 VSS 0.333965f
C5147 DVSS.n5287 VSS 0.333965f
C5148 DVSS.n5288 VSS 0.333965f
C5149 DVSS.n5289 VSS 0.333965f
C5150 DVSS.n5290 VSS 0.333965f
C5151 DVSS.n5291 VSS 0.333965f
C5152 DVSS.n5292 VSS 0.333965f
C5153 DVSS.n5293 VSS 0.333965f
C5154 DVSS.n5294 VSS 0.333965f
C5155 DVSS.n5295 VSS 0.333965f
C5156 DVSS.n5296 VSS 0.333965f
C5157 DVSS.n5297 VSS 0.333965f
C5158 DVSS.n5298 VSS 0.333965f
C5159 DVSS.n5299 VSS 0.333965f
C5160 DVSS.n5300 VSS 0.333965f
C5161 DVSS.n5301 VSS 0.333965f
C5162 DVSS.n5302 VSS 0.333965f
C5163 DVSS.n5303 VSS 0.333965f
C5164 DVSS.n5304 VSS 0.333965f
C5165 DVSS.n5305 VSS 0.333965f
C5166 DVSS.n5306 VSS 0.333965f
C5167 DVSS.n5307 VSS 0.333965f
C5168 DVSS.n5308 VSS 0.333965f
C5169 DVSS.n5309 VSS 0.333965f
C5170 DVSS.n5310 VSS 0.333965f
C5171 DVSS.n5311 VSS 0.333965f
C5172 DVSS.n5312 VSS 0.333965f
C5173 DVSS.n5313 VSS 0.333965f
C5174 DVSS.n5314 VSS 0.333965f
C5175 DVSS.n5315 VSS 0.333965f
C5176 DVSS.n5316 VSS 0.333965f
C5177 DVSS.n5317 VSS 0.301038f
C5178 DVSS.n5318 VSS 0.333965f
C5179 DVSS.n5319 VSS 0.333965f
C5180 DVSS.n5320 VSS 0.333965f
C5181 DVSS.n5321 VSS 0.171686f
C5182 DVSS.n5322 VSS 1.53873f
C5183 DVSS.n5323 VSS 0.474474f
C5184 DVSS.n5324 VSS 0.301038f
C5185 DVSS.n5325 VSS 0.333965f
C5186 DVSS.n5326 VSS 0.333965f
C5187 DVSS.n5327 VSS 0.333965f
C5188 DVSS.n5328 VSS 0.333965f
C5189 DVSS.n5329 VSS 0.333965f
C5190 DVSS.n5330 VSS 0.333965f
C5191 DVSS.n5331 VSS 0.333965f
C5192 DVSS.n5332 VSS 0.333965f
C5193 DVSS.n5333 VSS 0.333965f
C5194 DVSS.n5334 VSS 0.333965f
C5195 DVSS.n5335 VSS 0.333965f
C5196 DVSS.n5336 VSS 0.333965f
C5197 DVSS.n5337 VSS 0.333965f
C5198 DVSS.n5338 VSS 0.333965f
C5199 DVSS.n5339 VSS 0.333965f
C5200 DVSS.n5340 VSS 0.248122f
C5201 DVSS.n5341 VSS 0.333965f
C5202 DVSS.n5342 VSS 0.333965f
C5203 DVSS.n5343 VSS 0.145816f
C5204 DVSS.n5344 VSS 0.166982f
C5205 DVSS.n5345 VSS 0.009721f
C5206 DVSS.n5346 VSS 0.031907f
C5207 DVSS.n5347 VSS 0.49201f
C5208 DVSS.n5348 VSS 0.63273f
C5209 DVSS.n5349 VSS 0.008222f
C5210 DVSS.n5350 VSS 0.014785f
C5211 DVSS.n5351 VSS 0.016872f
C5212 DVSS.n5352 VSS 0.015218f
C5213 DVSS.n5353 VSS 0.034593f
C5214 DVSS.n5354 VSS 0.01185f
C5215 DVSS.n5355 VSS 0.010715f
C5216 DVSS.n5356 VSS 0.011035f
C5217 DVSS.n5358 VSS 0.050794f
C5218 DVSS.n5359 VSS 0.011755f
C5219 DVSS.n5361 VSS 4.03585f
C5220 DVSS.n5363 VSS 0.052371f
C5221 DVSS.n5365 VSS 0.052371f
C5222 DVSS.n5367 VSS 0.052371f
C5223 DVSS.n5369 VSS 0.052371f
C5224 DVSS.n5371 VSS 0.052371f
C5225 DVSS.n5373 VSS 0.052371f
C5226 DVSS.n5376 VSS 0.111484f
C5227 DVSS.n5378 VSS 0.052371f
C5228 DVSS.n5380 VSS 0.052371f
C5229 DVSS.n5382 VSS 0.052371f
C5230 DVSS.n5384 VSS 0.052371f
C5231 DVSS.n5386 VSS 0.052371f
C5232 DVSS.n5388 VSS 0.052371f
C5233 DVSS.n5390 VSS 0.0403f
C5234 DVSS.n5391 VSS 0.01185f
C5235 DVSS.n5392 VSS 0.014633f
C5236 DVSS.n5393 VSS 0.051194f
C5237 DVSS.n5395 VSS 0.055349f
C5238 DVSS.n5397 VSS 0.018232f
C5239 DVSS.n5398 VSS 0.149568f
C5240 DVSS.n5399 VSS 0.052371f
C5241 DVSS.n5400 VSS 0.018232f
C5242 DVSS.n5402 VSS 0.018232f
C5243 DVSS.n5404 VSS 0.018232f
C5244 DVSS.n5405 VSS 0.052371f
C5245 DVSS.n5406 VSS 0.052371f
C5246 DVSS.n5407 VSS 0.018232f
C5247 DVSS.n5409 VSS 0.018232f
C5248 DVSS.n5411 VSS 0.018232f
C5249 DVSS.n5412 VSS 0.052371f
C5250 DVSS.n5413 VSS 0.052371f
C5251 DVSS.n5414 VSS 0.018232f
C5252 DVSS.n5416 VSS 0.018232f
C5253 DVSS.n5418 VSS 0.018232f
C5254 DVSS.n5419 VSS 0.052371f
C5255 DVSS.n5420 VSS 0.052371f
C5256 DVSS.n5421 VSS 0.018232f
C5257 DVSS.n5423 VSS 0.018232f
C5258 DVSS.n5425 VSS 0.018232f
C5259 DVSS.n5426 VSS 0.052371f
C5260 DVSS.n5427 VSS 0.052371f
C5261 DVSS.n5428 VSS 0.018232f
C5262 DVSS.n5430 VSS 0.018232f
C5263 DVSS.n5432 VSS 0.018232f
C5264 DVSS.n5433 VSS 0.052371f
C5265 DVSS.n5434 VSS 0.052371f
C5266 DVSS.n5435 VSS 0.018232f
C5267 DVSS.n5437 VSS 0.018232f
C5268 DVSS.n5439 VSS 0.018232f
C5269 DVSS.n5440 VSS 0.052371f
C5270 DVSS.n5441 VSS 0.040886f
C5271 DVSS.n5442 VSS 0.018232f
C5272 DVSS.n5444 VSS 0.018232f
C5273 DVSS.n5445 VSS 0.037671f
C5274 DVSS.n5446 VSS 0.028712f
C5275 DVSS.n5447 VSS 0.018232f
C5276 DVSS.n5449 VSS 0.018232f
C5277 DVSS.n5450 VSS 0.049845f
C5278 DVSS.n5451 VSS 0.052371f
C5279 DVSS.n5452 VSS 0.018232f
C5280 DVSS.n5454 VSS 0.018232f
C5281 DVSS.n5456 VSS 0.018232f
C5282 DVSS.n5457 VSS 0.052371f
C5283 DVSS.n5458 VSS 0.052371f
C5284 DVSS.n5459 VSS 0.018232f
C5285 DVSS.n5461 VSS 0.018232f
C5286 DVSS.n5463 VSS 0.018232f
C5287 DVSS.n5464 VSS 0.052371f
C5288 DVSS.n5465 VSS 0.052371f
C5289 DVSS.n5466 VSS 0.018232f
C5290 DVSS.n5468 VSS 0.018232f
C5291 DVSS.n5470 VSS 0.018232f
C5292 DVSS.n5471 VSS 0.052371f
C5293 DVSS.n5472 VSS 0.052371f
C5294 DVSS.n5473 VSS 0.018232f
C5295 DVSS.n5475 VSS 0.018232f
C5296 DVSS.n5477 VSS 0.018232f
C5297 DVSS.n5478 VSS 0.052371f
C5298 DVSS.n5479 VSS 0.052371f
C5299 DVSS.n5480 VSS 0.018232f
C5300 DVSS.n5482 VSS 0.018232f
C5301 DVSS.n5484 VSS 0.018232f
C5302 DVSS.n5485 VSS 0.052371f
C5303 DVSS.n5486 VSS 0.052371f
C5304 DVSS.n5487 VSS 0.018232f
C5305 DVSS.n5489 VSS 0.018232f
C5306 DVSS.n5491 VSS 0.018232f
C5307 DVSS.n5492 VSS 0.052371f
C5308 DVSS.n5493 VSS 0.052371f
C5309 DVSS.n5494 VSS 0.018232f
C5310 DVSS.n5496 VSS 0.018232f
C5311 DVSS.n5498 VSS 0.018232f
C5312 DVSS.n5499 VSS 0.072284f
C5313 DVSS.n5500 VSS 0.088919f
C5314 DVSS.n5501 VSS 0.016745f
C5315 DVSS.n5502 VSS 0.02143f
C5316 DVSS.n5503 VSS 1.33697f
C5317 DVSS.n5504 VSS 0.02143f
C5318 DVSS.n5505 VSS 0.014785f
C5319 DVSS.n5506 VSS 0.008222f
C5320 DVSS.n5507 VSS 0.40405f
C5321 DVSS.n5508 VSS 0.182034f
C5322 DVSS.n5509 VSS 0.077925f
C5323 DVSS.n5510 VSS 0.15585f
C5324 DVSS.n5511 VSS 0.15585f
C5325 DVSS.n5512 VSS 0.15585f
C5326 DVSS.n5513 VSS 0.11579f
C5327 DVSS.n5514 VSS 0.15585f
C5328 DVSS.n5515 VSS 0.15585f
C5329 DVSS.n5516 VSS 0.15585f
C5330 DVSS.n5517 VSS 0.15585f
C5331 DVSS.n5518 VSS 0.15585f
C5332 DVSS.n5519 VSS 0.15585f
C5333 DVSS.n5520 VSS 0.15585f
C5334 DVSS.n5521 VSS 0.15585f
C5335 DVSS.n5522 VSS 0.751144f
C5336 DVSS.n5523 VSS 0.205146f
C5337 DVSS.n5524 VSS 0.017561f
C5338 DVSS.n5525 VSS 0.140485f
C5339 DVSS.n5526 VSS 0.140485f
C5340 DVSS.n5527 VSS 0.140485f
C5341 DVSS.n5528 VSS 0.15585f
C5342 DVSS.n5529 VSS 0.15585f
C5343 DVSS.n5530 VSS 0.15585f
C5344 DVSS.n5531 VSS 0.15585f
C5345 DVSS.n5532 VSS 0.15585f
C5346 DVSS.n5533 VSS 0.15585f
C5347 DVSS.n5534 VSS 0.15585f
C5348 DVSS.n5535 VSS 0.15585f
C5349 DVSS.n5536 VSS 0.15585f
C5350 DVSS.n5537 VSS 0.15585f
C5351 DVSS.n5538 VSS 0.15585f
C5352 DVSS.n5539 VSS 0.15585f
C5353 DVSS.n5540 VSS 0.15585f
C5354 DVSS.n5541 VSS 0.15585f
C5355 DVSS.n5542 VSS 0.15585f
C5356 DVSS.n5543 VSS 0.15585f
C5357 DVSS.n5544 VSS 0.15585f
C5358 DVSS.n5545 VSS 0.15585f
C5359 DVSS.n5546 VSS 0.15585f
C5360 DVSS.n5547 VSS 0.15585f
C5361 DVSS.n5548 VSS 0.15585f
C5362 DVSS.n5549 VSS 0.15585f
C5363 DVSS.n5550 VSS 0.15585f
C5364 DVSS.n5551 VSS 0.068047f
C5365 DVSS.n5552 VSS 0.077925f
C5366 DVSS.n5553 VSS 0.127863f
C5367 DVSS.n5554 VSS 0.15585f
C5368 DVSS.n5555 VSS 0.15585f
C5369 DVSS.n5556 VSS 0.15585f
C5370 DVSS.n5557 VSS 0.15585f
C5371 DVSS.n5558 VSS 0.15585f
C5372 DVSS.n5559 VSS 0.15585f
C5373 DVSS.n5560 VSS 0.15585f
C5374 DVSS.n5561 VSS 0.15585f
C5375 DVSS.n5562 VSS 0.15585f
C5376 DVSS.n5563 VSS 0.15585f
C5377 DVSS.n5564 VSS 0.15585f
C5378 DVSS.n5565 VSS 0.15585f
C5379 DVSS.n5566 VSS 0.15585f
C5380 DVSS.n5567 VSS 0.15585f
C5381 DVSS.n5568 VSS 0.15585f
C5382 DVSS.n5569 VSS 0.15585f
C5383 DVSS.n5570 VSS 0.15585f
C5384 DVSS.n5571 VSS 0.15585f
C5385 DVSS.n5572 VSS 0.15585f
C5386 DVSS.n5573 VSS 0.15585f
C5387 DVSS.n5574 VSS 0.15585f
C5388 DVSS.n5575 VSS 0.15585f
C5389 DVSS.n5576 VSS 0.15585f
C5390 DVSS.n5577 VSS 0.15585f
C5391 DVSS.n5578 VSS 0.15585f
C5392 DVSS.n5579 VSS 0.15585f
C5393 DVSS.n5580 VSS 0.15585f
C5394 DVSS.n5581 VSS 0.15585f
C5395 DVSS.n5582 VSS 0.15585f
C5396 DVSS.n5583 VSS 0.15585f
C5397 DVSS.n5584 VSS 0.091644f
C5398 DVSS.n5585 VSS 0.077925f
C5399 DVSS.n5586 VSS 0.038884f
C5400 DVSS.n5587 VSS 0.341867f
C5401 DVSS.n5588 VSS 0.066322f
C5402 DVSS.n5589 VSS 0.008467f
C5403 DVSS.n5590 VSS 0.008467f
C5404 DVSS.n5591 VSS 0.09674f
C5405 DVSS.n5592 VSS 0.117436f
C5406 DVSS.n5593 VSS 0.048537f
C5407 DVSS.n5594 VSS 0.119743f
C5408 DVSS.n5595 VSS 0.125047f
C5409 DVSS.n5596 VSS 0.09674f
C5410 DVSS.n5597 VSS 0.008467f
C5411 DVSS.n5598 VSS 1.00544f
C5412 DVSS.n5599 VSS 0.066322f
C5413 DVSS.n5600 VSS 0.257582f
C5414 DVSS.n5601 VSS 0.07508f
C5415 DVSS.t128 VSS 0.203828f
C5416 DVSS.t98 VSS 0.203828f
C5417 DVSS.n5602 VSS 0.407656f
C5418 DVSS.n5603 VSS 0.073484f
C5419 DVSS.n5604 VSS 0.176594f
C5420 DVSS.n5605 VSS 0.138598f
C5421 DVSS.n5606 VSS 0.118999f
C5422 DVSS.n5607 VSS 0.07508f
C5423 DVSS.t150 VSS 0.203828f
C5424 DVSS.t118 VSS 0.203828f
C5425 DVSS.n5608 VSS 0.407656f
C5426 DVSS.n5609 VSS 0.073484f
C5427 DVSS.n5610 VSS 0.176594f
C5428 DVSS.n5611 VSS 0.076514f
C5429 DVSS.n5612 VSS 0.076514f
C5430 DVSS.n5613 VSS 0.176594f
C5431 DVSS.t36 VSS 0.203828f
C5432 DVSS.t88 VSS 0.203828f
C5433 DVSS.n5614 VSS 0.407656f
C5434 DVSS.n5615 VSS 0.073484f
C5435 DVSS.n5616 VSS 0.205057f
C5436 DVSS.n5617 VSS 0.205057f
C5437 DVSS.n5618 VSS 0.07508f
C5438 DVSS.t64 VSS 0.203828f
C5439 DVSS.t108 VSS 0.203828f
C5440 DVSS.n5619 VSS 0.407656f
C5441 DVSS.n5620 VSS 0.073484f
C5442 DVSS.n5621 VSS 0.176594f
C5443 DVSS.n5622 VSS 0.118999f
C5444 DVSS.n5623 VSS 0.118999f
C5445 DVSS.n5624 VSS 0.07508f
C5446 DVSS.t78 VSS 0.203828f
C5447 DVSS.t120 VSS 0.203828f
C5448 DVSS.n5625 VSS 0.407656f
C5449 DVSS.n5626 VSS 0.073484f
C5450 DVSS.n5627 VSS 0.176594f
C5451 DVSS.n5628 VSS 0.076514f
C5452 DVSS.n5629 VSS 0.076514f
C5453 DVSS.n5630 VSS 0.176594f
C5454 DVSS.t50 VSS 0.203828f
C5455 DVSS.t142 VSS 0.203828f
C5456 DVSS.n5631 VSS 0.407656f
C5457 DVSS.n5632 VSS 0.073484f
C5458 DVSS.n5633 VSS 0.205057f
C5459 DVSS.n5634 VSS 0.205057f
C5460 DVSS.n5635 VSS 0.07508f
C5461 DVSS.t66 VSS 0.203828f
C5462 DVSS.t30 VSS 0.203828f
C5463 DVSS.n5636 VSS 0.407656f
C5464 DVSS.n5637 VSS 0.073484f
C5465 DVSS.n5638 VSS 0.176594f
C5466 DVSS.n5639 VSS 0.118999f
C5467 DVSS.n5640 VSS 0.118999f
C5468 DVSS.n5641 VSS 0.176594f
C5469 DVSS.n5642 VSS 0.073484f
C5470 DVSS.n5643 VSS 0.07508f
C5471 DVSS.n5644 VSS 0.174976f
C5472 DVSS.n5645 VSS 0.076514f
C5473 DVSS.n5646 VSS 0.076514f
C5474 DVSS.n5647 VSS 0.076514f
C5475 DVSS.n5648 VSS 0.076514f
C5476 DVSS.n5649 VSS 0.076514f
C5477 DVSS.n5650 VSS 0.076514f
C5478 DVSS.n5651 VSS 0.076514f
C5479 DVSS.n5652 VSS 0.096113f
C5480 DVSS.n5653 VSS 0.066322f
C5481 DVSS.n5654 VSS 0.008467f
C5482 DVSS.n5655 VSS 0.008467f
C5483 DVSS.n5656 VSS 0.09674f
C5484 DVSS.n5657 VSS 0.117436f
C5485 DVSS.n5658 VSS 0.034583f
C5486 DVSS.n5659 VSS 0.043638f
C5487 DVSS.n5660 VSS 0.111199f
C5488 DVSS.n5661 VSS 0.220734f
C5489 DVSS.n5662 VSS 1.33014f
C5490 DVSS.n5663 VSS 6.42185f
C5491 DVSS.n5664 VSS 3.42532f
C5492 DVSS.n5665 VSS 2.42146f
C5493 DVSS.n5666 VSS 3.9288f
C5494 DVSS.n5667 VSS 2.42546f
C5495 DVSS.n5668 VSS 4.46039f
C5496 DVSS.n5669 VSS 9.37817f
C5497 DVSS.n5670 VSS -1.87637f
C5498 DVSS.n5671 VSS 6.42185f
C5499 DVSS.n5672 VSS 1.86901f
C5500 DVSS.t6 VSS 2.03481f
C5501 DVSS.n5673 VSS 0.85943f
C5502 DVSS.n5674 VSS 0.195303f
C5503 DVSS.n5675 VSS 0.027206f
C5504 DVSS.n5676 VSS 0.047806f
C5505 DVSS.n5677 VSS 0.042947f
C5506 DVSS.n5678 VSS 0.041083f
C5507 DVSS.n5679 VSS 0.035698f
C5508 DVSS.n5680 VSS 0.314729f
C5509 DVSS.n5681 VSS 0.259263f
C5510 DVSS.n5682 VSS 0.342732f
C5511 DVSS.n5683 VSS 0.045382f
C5512 DVSS.n5684 VSS 3.11004f
C5513 DVSS.t127 VSS 4.53554f
C5514 DVSS.t97 VSS 2.28624f
C5515 DVSS.t149 VSS 2.28624f
C5516 DVSS.t117 VSS 2.28624f
C5517 DVSS.t35 VSS 2.28624f
C5518 DVSS.t87 VSS 2.28624f
C5519 DVSS.t63 VSS 2.28624f
C5520 DVSS.t107 VSS 2.28624f
C5521 DVSS.t77 VSS 2.28624f
C5522 DVSS.t119 VSS 2.28624f
C5523 DVSS.t49 VSS 2.28624f
C5524 DVSS.t141 VSS 2.28624f
C5525 DVSS.t65 VSS 2.28624f
C5526 DVSS.t29 VSS 2.28624f
C5527 DVSS.t91 VSS 2.28624f
C5528 DVSS.t163 VSS 2.28624f
C5529 DVSS.t99 VSS 2.28624f
C5530 DVSS.t173 VSS 2.28624f
C5531 DVSS.t121 VSS 2.28624f
C5532 DVSS.t41 VSS 4.03839f
C5533 DVSS.t183 VSS 2.28624f
C5534 DVSS.t59 VSS 2.28624f
C5535 DVSS.t167 VSS 2.28624f
C5536 DVSS.t93 VSS 2.28624f
C5537 DVSS.t123 VSS 2.28624f
C5538 DVSS.t73 VSS 2.28624f
C5539 DVSS.t103 VSS 2.28624f
C5540 DVSS.t53 VSS 2.28624f
C5541 DVSS.t131 VSS 2.28624f
C5542 DVSS.t31 VSS 2.28624f
C5543 DVSS.t111 VSS 2.28624f
C5544 DVSS.t177 VSS 2.28624f
C5545 DVSS.t101 VSS 2.28624f
C5546 DVSS.t85 VSS 2.28624f
C5547 DVSS.t151 VSS 2.28624f
C5548 DVSS.t69 VSS 2.28624f
C5549 DVSS.t133 VSS 2.28624f
C5550 DVSS.t47 VSS 2.28624f
C5551 DVSS.t161 VSS 4.03839f
C5552 DVSS.n5685 VSS 4.97951f
C5553 DVSS.n5686 VSS -0.795461f
C5554 DVSS.n5687 VSS 0.166819f
C5555 DVSS.n5688 VSS 0.171366f
C5556 DVSS.n5689 VSS 0.166819f
C5557 DVSS.n5690 VSS 0.246657f
C5558 DVSS.t162 VSS 0.203828f
C5559 DVSS.t48 VSS 0.203828f
C5560 DVSS.n5691 VSS 0.407656f
C5561 DVSS.n5692 VSS 0.073484f
C5562 DVSS.n5693 VSS 0.176594f
C5563 DVSS.n5694 VSS 0.134521f
C5564 DVSS.n5695 VSS 0.062246f
C5565 DVSS.n5696 VSS 0.134521f
C5566 DVSS.n5697 VSS 0.062246f
C5567 DVSS.n5698 VSS 0.048035f
C5568 DVSS.n5699 VSS 0.170933f
C5569 DVSS.n5700 VSS 0.170933f
C5570 DVSS.n5701 VSS 0.062246f
C5571 DVSS.n5703 VSS 0.062246f
C5572 DVSS.n5704 VSS 0.092036f
C5573 DVSS.n5705 VSS 0.076514f
C5574 DVSS.n5706 VSS 0.176594f
C5575 DVSS.n5707 VSS 0.073484f
C5576 DVSS.n5708 VSS 0.205057f
C5577 DVSS.n5709 VSS 0.07508f
C5578 DVSS.n5710 VSS 0.174976f
C5579 DVSS.n5711 VSS 0.119007f
C5580 DVSS.n5713 VSS 0.048035f
C5581 DVSS.n5714 VSS 0.170933f
C5582 DVSS.n5715 VSS 0.062246f
C5583 DVSS.n5716 VSS 0.134529f
C5584 DVSS.n5717 VSS 0.174976f
C5585 DVSS.n5718 VSS 0.092036f
C5586 DVSS.n5719 VSS 0.062246f
C5587 DVSS.n5720 VSS 0.171366f
C5588 DVSS.n5721 VSS 0.062246f
C5589 DVSS.n5722 VSS 0.092036f
C5590 DVSS.n5723 VSS 0.174976f
C5591 DVSS.n5724 VSS 0.134529f
C5592 DVSS.n5725 VSS 0.119007f
C5593 DVSS.n5726 VSS 0.174976f
C5594 DVSS.n5727 VSS 0.07508f
C5595 DVSS.t134 VSS 0.203828f
C5596 DVSS.t70 VSS 0.203828f
C5597 DVSS.n5728 VSS 0.407656f
C5598 DVSS.n5729 VSS 0.073484f
C5599 DVSS.n5730 VSS 0.176594f
C5600 DVSS.n5731 VSS 0.076514f
C5601 DVSS.n5732 VSS 0.076514f
C5602 DVSS.n5733 VSS 0.176594f
C5603 DVSS.n5734 VSS 0.073484f
C5604 DVSS.n5735 VSS 0.205057f
C5605 DVSS.n5736 VSS 0.07508f
C5606 DVSS.n5737 VSS 0.174976f
C5607 DVSS.n5738 VSS 0.076514f
C5608 DVSS.n5739 VSS 0.076514f
C5609 DVSS.n5740 VSS 0.174976f
C5610 DVSS.n5741 VSS 0.119007f
C5611 DVSS.n5742 VSS 0.119007f
C5612 DVSS.n5743 VSS 0.174976f
C5613 DVSS.n5744 VSS 0.07508f
C5614 DVSS.t112 VSS 0.203828f
C5615 DVSS.t32 VSS 0.203828f
C5616 DVSS.n5745 VSS 0.407656f
C5617 DVSS.n5746 VSS 0.073484f
C5618 DVSS.n5747 VSS 0.176594f
C5619 DVSS.n5748 VSS 0.076514f
C5620 DVSS.n5749 VSS 0.076514f
C5621 DVSS.n5750 VSS 0.176594f
C5622 DVSS.n5751 VSS 0.073484f
C5623 DVSS.n5752 VSS 0.205057f
C5624 DVSS.n5753 VSS 0.07508f
C5625 DVSS.n5754 VSS 0.174976f
C5626 DVSS.n5755 VSS 0.076514f
C5627 DVSS.n5756 VSS 0.076514f
C5628 DVSS.n5757 VSS 0.174976f
C5629 DVSS.n5758 VSS 0.119007f
C5630 DVSS.n5759 VSS 0.076514f
C5631 DVSS.n5760 VSS 0.174976f
C5632 DVSS.n5761 VSS 0.119007f
C5633 DVSS.n5762 VSS 0.119007f
C5634 DVSS.n5763 VSS 0.174976f
C5635 DVSS.n5764 VSS 0.07508f
C5636 DVSS.t124 VSS 0.203828f
C5637 DVSS.t94 VSS 0.203828f
C5638 DVSS.n5765 VSS 0.407656f
C5639 DVSS.n5766 VSS 0.073484f
C5640 DVSS.n5767 VSS 0.176594f
C5641 DVSS.n5768 VSS 0.076514f
C5642 DVSS.n5769 VSS 0.076514f
C5643 DVSS.n5770 VSS 0.176594f
C5644 DVSS.t168 VSS 0.203828f
C5645 DVSS.t60 VSS 0.203828f
C5646 DVSS.n5771 VSS 0.407656f
C5647 DVSS.n5772 VSS 0.073484f
C5648 DVSS.n5773 VSS 0.205057f
C5649 DVSS.n5775 VSS 0.077925f
C5650 DVSS.n5776 VSS 0.074084f
C5651 DVSS.n5777 VSS 0.068047f
C5652 DVSS.n5778 VSS 0.052105f
C5653 DVSS.n5779 VSS 0.052105f
C5654 DVSS.n5780 VSS 0.04286f
C5655 DVSS.n5781 VSS 0.091644f
C5656 DVSS.n5782 VSS 0.103006f
C5657 DVSS.n5783 VSS 0.176594f
C5658 DVSS.t52 VSS 0.203828f
C5659 DVSS.t144 VSS 0.203828f
C5660 DVSS.n5784 VSS 0.407656f
C5661 DVSS.n5785 VSS 0.073484f
C5662 DVSS.n5786 VSS 0.162197f
C5663 DVSS.n5787 VSS 0.085721f
C5664 DVSS.n5788 VSS 0.052105f
C5665 DVSS.n5790 VSS 0.052105f
C5666 DVSS.n5792 VSS 0.030675f
C5667 DVSS.n5798 VSS 0.071889f
C5668 DVSS.n5799 VSS 0.052206f
C5669 DVSS.n5800 VSS 0.01317f
C5670 DVSS.n5802 VSS 0.068047f
C5671 DVSS.n5803 VSS 0.009721f
C5672 DVSS.n5804 VSS 0.091644f
C5673 DVSS.n5805 VSS 0.031985f
C5674 DVSS.n5806 VSS 0.019442f
C5675 DVSS.n5807 VSS 0.009721f
C5676 DVSS.n5808 VSS 0.15585f
C5677 DVSS.n5809 VSS 0.15585f
C5678 DVSS.n5810 VSS 0.15585f
C5679 DVSS.n5811 VSS 0.15585f
C5680 DVSS.n5812 VSS 0.15585f
C5681 DVSS.n5813 VSS 0.15585f
C5682 DVSS.n5814 VSS 0.15585f
C5683 DVSS.n5815 VSS 0.15585f
C5684 DVSS.n5816 VSS 0.15585f
C5685 DVSS.n5817 VSS 0.15585f
C5686 DVSS.n5818 VSS 0.15585f
C5687 DVSS.n5819 VSS 0.15585f
C5688 DVSS.n5820 VSS 0.15585f
C5689 DVSS.n5821 VSS 0.15585f
C5690 DVSS.n5822 VSS 0.15585f
C5691 DVSS.n5823 VSS 0.15585f
C5692 DVSS.n5824 VSS 0.068047f
C5693 DVSS.n5825 VSS 0.15585f
C5694 DVSS.n5826 VSS 0.15585f
C5695 DVSS.n5827 VSS 0.15585f
C5696 DVSS.n5828 VSS 0.15585f
C5697 DVSS.n5829 VSS 0.15585f
C5698 DVSS.n5830 VSS 0.15585f
C5699 DVSS.n5831 VSS 0.15585f
C5700 DVSS.n5832 VSS 0.15585f
C5701 DVSS.n5833 VSS 0.15585f
C5702 DVSS.n5834 VSS 0.15585f
C5703 DVSS.n5835 VSS 0.15585f
C5704 DVSS.n5836 VSS 0.15585f
C5705 DVSS.n5837 VSS 0.15585f
C5706 DVSS.n5838 VSS 0.15585f
C5707 DVSS.n5839 VSS 0.15585f
C5708 DVSS.n5840 VSS 0.15585f
C5709 DVSS.n5841 VSS 0.15585f
C5710 DVSS.n5842 VSS 0.15585f
C5711 DVSS.n5843 VSS 0.15585f
C5712 DVSS.n5844 VSS 0.15585f
C5713 DVSS.n5845 VSS 0.15585f
C5714 DVSS.n5846 VSS 0.15585f
C5715 DVSS.n5847 VSS 0.15585f
C5716 DVSS.n5848 VSS 0.15585f
C5717 DVSS.n5849 VSS 0.15585f
C5718 DVSS.n5850 VSS 0.15585f
C5719 DVSS.n5851 VSS 0.15585f
C5720 DVSS.n5852 VSS 0.15585f
C5721 DVSS.n5853 VSS 0.15585f
C5722 DVSS.n5854 VSS 0.15585f
C5723 DVSS.n5855 VSS 0.506941f
C5724 DVSS.n5856 VSS 2.43723f
C5725 DVSS.n5857 VSS 0.15585f
C5726 DVSS.n5858 VSS 0.15585f
C5727 DVSS.n5859 VSS 0.15585f
C5728 DVSS.n5860 VSS 0.15585f
C5729 DVSS.n5861 VSS 0.15585f
C5730 DVSS.n5862 VSS 0.15585f
C5731 DVSS.n5863 VSS 0.15585f
C5732 DVSS.n5864 VSS 0.15585f
C5733 DVSS.n5865 VSS 0.15585f
C5734 DVSS.n5866 VSS 0.15585f
C5735 DVSS.n5867 VSS 0.15585f
C5736 DVSS.n5868 VSS 0.15585f
C5737 DVSS.n5869 VSS 0.15585f
C5738 DVSS.n5870 VSS 0.15585f
C5739 DVSS.n5871 VSS 0.15585f
C5740 DVSS.n5872 VSS 0.15585f
C5741 DVSS.n5873 VSS 0.15585f
C5742 DVSS.n5874 VSS 0.15585f
C5743 DVSS.n5875 VSS 0.15585f
C5744 DVSS.n5876 VSS 0.15585f
C5745 DVSS.n5877 VSS 0.15585f
C5746 DVSS.n5878 VSS 0.15585f
C5747 DVSS.n5879 VSS 0.15585f
C5748 DVSS.n5880 VSS 0.15585f
C5749 DVSS.n5881 VSS 0.15585f
C5750 DVSS.n5882 VSS 0.15585f
C5751 DVSS.n5883 VSS 0.15585f
C5752 DVSS.n5884 VSS 0.15585f
C5753 DVSS.n5885 VSS 0.15585f
C5754 DVSS.n5886 VSS 0.15585f
C5755 DVSS.n5887 VSS 0.15585f
C5756 DVSS.n5888 VSS 0.15585f
C5757 DVSS.n5889 VSS 0.15585f
C5758 DVSS.n5890 VSS 0.15585f
C5759 DVSS.n5891 VSS 0.15585f
C5760 DVSS.n5892 VSS 0.15585f
C5761 DVSS.n5893 VSS 0.15585f
C5762 DVSS.n5894 VSS 0.15585f
C5763 DVSS.n5895 VSS 0.15585f
C5764 DVSS.n5896 VSS 0.15585f
C5765 DVSS.n5897 VSS 0.15585f
C5766 DVSS.n5898 VSS 0.15585f
C5767 DVSS.n5899 VSS 0.15585f
C5768 DVSS.n5900 VSS 0.15585f
C5769 DVSS.n5901 VSS 0.15585f
C5770 DVSS.n5902 VSS 0.15585f
C5771 DVSS.n5903 VSS 0.15585f
C5772 DVSS.n5904 VSS 0.15585f
C5773 DVSS.n5905 VSS 0.15585f
C5774 DVSS.n5906 VSS 0.15585f
C5775 DVSS.n5907 VSS 0.15585f
C5776 DVSS.n5908 VSS 0.15585f
C5777 DVSS.n5909 VSS 0.15585f
C5778 DVSS.n5910 VSS 0.15585f
C5779 DVSS.n5911 VSS 0.15585f
C5780 DVSS.n5912 VSS 0.15585f
C5781 DVSS.n5913 VSS 0.15585f
C5782 DVSS.n5914 VSS 0.15585f
C5783 DVSS.n5915 VSS 0.15585f
C5784 DVSS.n5916 VSS 0.15585f
C5785 DVSS.n5917 VSS 0.15585f
C5786 DVSS.n5918 VSS 0.15585f
C5787 DVSS.n5919 VSS 0.093839f
C5788 DVSS.n5920 VSS 0.15585f
C5789 DVSS.n5921 VSS 0.15585f
C5790 DVSS.n5922 VSS 0.15585f
C5791 DVSS.n5923 VSS 0.15585f
C5792 DVSS.n5924 VSS 0.15585f
C5793 DVSS.n5925 VSS 0.15585f
C5794 DVSS.n5926 VSS 0.15585f
C5795 DVSS.n5927 VSS 0.15585f
C5796 DVSS.n5928 VSS 0.15585f
C5797 DVSS.n5929 VSS 0.15585f
C5798 DVSS.n5930 VSS 0.15585f
C5799 DVSS.n5931 VSS 0.15585f
C5800 DVSS.n5932 VSS 0.15585f
C5801 DVSS.n5933 VSS 0.15585f
C5802 DVSS.n5934 VSS 0.15585f
C5803 DVSS.n5935 VSS 0.15585f
C5804 DVSS.n5936 VSS 0.15585f
C5805 DVSS.n5937 VSS 0.15585f
C5806 DVSS.n5938 VSS 0.15585f
C5807 DVSS.n5939 VSS 0.15585f
C5808 DVSS.n5940 VSS 0.15585f
C5809 DVSS.n5941 VSS 0.15585f
C5810 DVSS.n5942 VSS 0.15585f
C5811 DVSS.n5943 VSS 0.15585f
C5812 DVSS.n5944 VSS 0.15585f
C5813 DVSS.n5945 VSS 0.15585f
C5814 DVSS.n5946 VSS 0.15585f
C5815 DVSS.n5947 VSS 0.15585f
C5816 DVSS.n5948 VSS 0.15585f
C5817 DVSS.n5949 VSS 0.15585f
C5818 DVSS.n5950 VSS 0.15585f
C5819 DVSS.n5951 VSS 0.15585f
C5820 DVSS.n5952 VSS 0.15585f
C5821 DVSS.n5953 VSS 0.15585f
C5822 DVSS.n5954 VSS 0.15585f
C5823 DVSS.n5955 VSS 0.15585f
C5824 DVSS.n5956 VSS 0.15585f
C5825 DVSS.n5957 VSS 0.15585f
C5826 DVSS.n5958 VSS 0.15585f
C5827 DVSS.n5959 VSS 0.15585f
C5828 DVSS.n5960 VSS 0.15585f
C5829 DVSS.n5961 VSS 0.15585f
C5830 DVSS.n5962 VSS 0.15585f
C5831 DVSS.n5963 VSS 0.15585f
C5832 DVSS.n5964 VSS 0.15585f
C5833 DVSS.n5965 VSS 0.15585f
C5834 DVSS.n5966 VSS 0.15585f
C5835 DVSS.n5967 VSS 0.15585f
C5836 DVSS.n5968 VSS 0.15585f
C5837 DVSS.n5969 VSS 0.15585f
C5838 DVSS.n5970 VSS 0.15585f
C5839 DVSS.n5971 VSS 0.15585f
C5840 DVSS.n5972 VSS 0.15585f
C5841 DVSS.n5973 VSS 0.15585f
C5842 DVSS.n5974 VSS 0.15585f
C5843 DVSS.n5975 VSS 0.15585f
C5844 DVSS.n5976 VSS 0.15585f
C5845 DVSS.n5977 VSS 0.15585f
C5846 DVSS.n5978 VSS 0.15585f
C5847 DVSS.n5979 VSS 0.15585f
C5848 DVSS.n5980 VSS 0.15585f
C5849 DVSS.n5981 VSS 0.751144f
C5850 DVSS.n5982 VSS 0.205146f
C5851 DVSS.n5983 VSS 0.08012f
C5852 DVSS.n5984 VSS 0.15585f
C5853 DVSS.n5985 VSS 0.140485f
C5854 DVSS.n5986 VSS 0.140485f
C5855 DVSS.n5987 VSS 0.15585f
C5856 DVSS.n5988 VSS 0.15585f
C5857 DVSS.n5989 VSS 0.15585f
C5858 DVSS.n5990 VSS 0.15585f
C5859 DVSS.n5991 VSS 0.15585f
C5860 DVSS.n5992 VSS 0.15585f
C5861 DVSS.n5993 VSS 0.15585f
C5862 DVSS.n5994 VSS 0.15585f
C5863 DVSS.n5995 VSS 0.15585f
C5864 DVSS.n5996 VSS 0.15585f
C5865 DVSS.n5997 VSS 0.15585f
C5866 DVSS.n5998 VSS 0.15585f
C5867 DVSS.n5999 VSS 0.15585f
C5868 DVSS.n6000 VSS 0.15585f
C5869 DVSS.n6001 VSS 0.15585f
C5870 DVSS.n6002 VSS 0.15585f
C5871 DVSS.n6003 VSS 0.15585f
C5872 DVSS.n6004 VSS 0.15585f
C5873 DVSS.n6005 VSS 0.15585f
C5874 DVSS.n6006 VSS 0.15585f
C5875 DVSS.n6007 VSS 0.15585f
C5876 DVSS.n6008 VSS 0.15585f
C5877 DVSS.n6009 VSS 0.15585f
C5878 DVSS.n6010 VSS 0.15585f
C5879 DVSS.n6011 VSS 0.127863f
C5880 DVSS.n6012 VSS 0.15585f
C5881 DVSS.n6013 VSS 0.15585f
C5882 DVSS.n6014 VSS 0.15585f
C5883 DVSS.n6015 VSS 0.15585f
C5884 DVSS.n6016 VSS 0.15585f
C5885 DVSS.n6017 VSS 0.15585f
C5886 DVSS.n6018 VSS 0.15585f
C5887 DVSS.n6019 VSS 0.15585f
C5888 DVSS.n6020 VSS 0.15585f
C5889 DVSS.n6021 VSS 0.15585f
C5890 DVSS.n6022 VSS 0.15585f
C5891 DVSS.n6023 VSS 0.15585f
C5892 DVSS.n6024 VSS 0.15585f
C5893 DVSS.n6025 VSS 0.15585f
C5894 DVSS.n6026 VSS 0.15585f
C5895 DVSS.n6027 VSS 0.15585f
C5896 DVSS.n6028 VSS 0.15585f
C5897 DVSS.n6029 VSS 0.15585f
C5898 DVSS.n6030 VSS 0.15585f
C5899 DVSS.n6031 VSS 0.15585f
C5900 DVSS.n6032 VSS 0.15585f
C5901 DVSS.n6033 VSS 0.15585f
C5902 DVSS.n6034 VSS 0.15585f
C5903 DVSS.n6035 VSS 0.15585f
C5904 DVSS.n6036 VSS 0.15585f
C5905 DVSS.n6037 VSS 0.15585f
C5906 DVSS.n6038 VSS 0.15585f
C5907 DVSS.n6039 VSS 0.15585f
C5908 DVSS.n6040 VSS 0.15585f
C5909 DVSS.n6041 VSS 0.15585f
C5910 DVSS.n6042 VSS 0.15585f
C5911 DVSS.n6043 VSS 0.15585f
C5912 DVSS.n6044 VSS 0.152009f
C5913 DVSS.n6045 VSS 0.019442f
C5914 DVSS.n6046 VSS 0.019442f
C5915 DVSS.n6047 VSS 0.009721f
C5916 DVSS.n6048 VSS 0.011446f
C5917 DVSS.n6049 VSS 0.077925f
C5918 DVSS.n6051 VSS 0.044529f
C5919 DVSS.n6052 VSS 0.077925f
C5920 DVSS.n6053 VSS 0.015993f
C5921 DVSS.n6054 VSS 0.009721f
C5922 DVSS.n6055 VSS 0.176594f
C5923 DVSS.t38 VSS 0.203828f
C5924 DVSS.t90 VSS 0.203828f
C5925 DVSS.n6056 VSS 0.407656f
C5926 DVSS.n6057 VSS 0.073484f
C5927 DVSS.n6058 VSS 0.026052f
C5928 DVSS.n6059 VSS 0.035297f
C5929 DVSS.n6060 VSS 0.077925f
C5930 DVSS.n6061 VSS 0.119337f
C5931 DVSS.n6062 VSS 0.195813f
C5932 DVSS.n6063 VSS 0.174976f
C5933 DVSS.n6064 VSS 0.07508f
C5934 DVSS.t184 VSS 0.203828f
C5935 DVSS.t84 VSS 0.203828f
C5936 DVSS.n6065 VSS 0.407656f
C5937 DVSS.n6066 VSS 0.073484f
C5938 DVSS.n6067 VSS 0.176594f
C5939 DVSS.n6068 VSS 0.115549f
C5940 DVSS.n6070 VSS 0.044529f
C5941 DVSS.n6071 VSS 0.077925f
C5942 DVSS.n6072 VSS 0.008467f
C5943 DVSS.n6073 VSS 0.009721f
C5944 DVSS.n6074 VSS 0.170933f
C5945 DVSS.n6075 VSS 0.170933f
C5946 DVSS.n6076 VSS 0.009721f
C5947 DVSS.n6077 VSS 0.171366f
C5948 DVSS.n6078 VSS 0.171366f
C5949 DVSS.n6079 VSS 0.026052f
C5950 DVSS.n6080 VSS 0.007789f
C5951 DVSS.n6081 VSS 0.171366f
C5952 DVSS.n6082 VSS 0.171366f
C5953 DVSS.n6083 VSS 0.009721f
C5954 DVSS.n6084 VSS 0.170933f
C5955 DVSS.n6085 VSS 0.009721f
C5956 DVSS.n6086 VSS 0.170933f
C5957 DVSS.n6088 VSS 0.009721f
C5958 DVSS.n6089 VSS 0.011446f
C5959 DVSS.n6090 VSS 2.1675f
C5960 DVSS.n6092 VSS 0.044529f
C5961 DVSS.n6093 VSS 0.077925f
C5962 DVSS.n6094 VSS 0.015993f
C5963 DVSS.n6095 VSS 0.052214f
C5964 DVSS.n6096 VSS 0.174976f
C5965 DVSS.n6097 VSS 0.009721f
C5966 DVSS.n6098 VSS 0.01317f
C5967 DVSS.n6099 VSS 0.077925f
C5968 DVSS.n6101 VSS 0.044529f
C5969 DVSS.n6102 VSS 0.077925f
C5970 DVSS.n6103 VSS 0.031985f
C5971 DVSS.n6104 VSS 0.060521f
C5972 DVSS.n6105 VSS 0.174976f
C5973 DVSS.n6106 VSS 0.103014f
C5974 DVSS.n6107 VSS 0.119007f
C5975 DVSS.n6108 VSS 0.174976f
C5976 DVSS.n6109 VSS 0.07508f
C5977 DVSS.t188 VSS 0.203828f
C5978 DVSS.t156 VSS 0.203828f
C5979 DVSS.n6110 VSS 0.407656f
C5980 DVSS.n6111 VSS 0.073484f
C5981 DVSS.n6112 VSS 0.176594f
C5982 DVSS.n6113 VSS 0.076514f
C5983 DVSS.n6114 VSS 0.076514f
C5984 DVSS.n6115 VSS 0.176594f
C5985 DVSS.t40 VSS 0.203828f
C5986 DVSS.t176 VSS 0.203828f
C5987 DVSS.n6116 VSS 0.407656f
C5988 DVSS.n6117 VSS 0.073484f
C5989 DVSS.n6118 VSS 0.205057f
C5990 DVSS.n6119 VSS 0.145809f
C5991 DVSS.t68 VSS 0.203828f
C5992 DVSS.t146 VSS 0.203828f
C5993 DVSS.n6120 VSS 0.407656f
C5994 DVSS.n6121 VSS 0.073484f
C5995 DVSS.n6122 VSS 0.176594f
C5996 DVSS.n6123 VSS 0.096891f
C5997 DVSS.n6124 VSS 0.009721f
C5998 DVSS.n6125 VSS 0.025871f
C5999 DVSS.n6126 VSS 0.019285f
C6000 DVSS.n6127 VSS 0.009721f
C6001 DVSS.n6128 VSS 0.009721f
C6002 DVSS.n6129 VSS 0.019442f
C6003 DVSS.n6130 VSS 0.019442f
C6004 DVSS.n6131 VSS 0.166982f
C6005 DVSS.n6132 VSS 0.145816f
C6006 DVSS.n6133 VSS 0.333965f
C6007 DVSS.n6134 VSS 0.333965f
C6008 DVSS.n6135 VSS 0.333965f
C6009 DVSS.n6136 VSS 0.333965f
C6010 DVSS.n6137 VSS 0.333965f
C6011 DVSS.n6138 VSS 0.333965f
C6012 DVSS.n6139 VSS 0.333965f
C6013 DVSS.n6140 VSS 0.333965f
C6014 DVSS.n6141 VSS 0.333965f
C6015 DVSS.n6142 VSS 0.333965f
C6016 DVSS.n6143 VSS 0.333965f
C6017 DVSS.n6144 VSS 0.333965f
C6018 DVSS.n6145 VSS 0.333965f
C6019 DVSS.n6146 VSS 0.333965f
C6020 DVSS.n6147 VSS 0.333965f
C6021 DVSS.n6148 VSS 0.333965f
C6022 DVSS.n6149 VSS 0.333965f
C6023 DVSS.n6150 VSS 0.333965f
C6024 DVSS.n6151 VSS 0.333965f
C6025 DVSS.n6152 VSS 0.333965f
C6026 DVSS.n6153 VSS 0.333965f
C6027 DVSS.n6154 VSS 0.333965f
C6028 DVSS.n6155 VSS 0.333965f
C6029 DVSS.n6156 VSS 0.333965f
C6030 DVSS.n6157 VSS 0.333965f
C6031 DVSS.n6158 VSS 0.333965f
C6032 DVSS.n6159 VSS 0.333965f
C6033 DVSS.n6160 VSS 0.333965f
C6034 DVSS.n6161 VSS 0.333965f
C6035 DVSS.n6162 VSS 0.333965f
C6036 DVSS.n6163 VSS 0.333965f
C6037 DVSS.n6164 VSS 0.333965f
C6038 DVSS.n6165 VSS 0.296335f
C6039 DVSS.n6166 VSS 0.296335f
C6040 DVSS.n6167 VSS 0.402169f
C6041 DVSS.n6168 VSS 0.204612f
C6042 DVSS.n6169 VSS 0.204612f
C6043 DVSS.n6170 VSS 0.333965f
C6044 DVSS.n6171 VSS 0.333965f
C6045 DVSS.n6172 VSS 0.333965f
C6046 DVSS.n6173 VSS 0.333965f
C6047 DVSS.n6174 VSS 0.333965f
C6048 DVSS.n6175 VSS 0.333965f
C6049 DVSS.n6176 VSS 0.333965f
C6050 DVSS.n6177 VSS 0.333965f
C6051 DVSS.n6178 VSS 0.333965f
C6052 DVSS.n6179 VSS 0.333965f
C6053 DVSS.n6180 VSS 0.333965f
C6054 DVSS.n6181 VSS 0.333965f
C6055 DVSS.n6182 VSS 0.333965f
C6056 DVSS.n6183 VSS 0.333965f
C6057 DVSS.n6184 VSS 0.333965f
C6058 DVSS.n6185 VSS 0.333965f
C6059 DVSS.n6186 VSS 0.333965f
C6060 DVSS.n6187 VSS 0.333965f
C6061 DVSS.n6188 VSS 0.145816f
C6062 DVSS.n6194 VSS 0.052105f
C6063 DVSS.n6196 VSS 0.166982f
C6064 DVSS.n6197 VSS 0.052105f
C6065 DVSS.n6199 VSS 0.166982f
C6066 DVSS.n6200 VSS 0.048323f
C6067 DVSS.n6201 VSS 0.026052f
C6068 DVSS.n6202 VSS 0.009721f
C6069 DVSS.n6203 VSS 0.052214f
C6070 DVSS.n6204 VSS 0.174976f
C6071 DVSS.n6205 VSS 0.07508f
C6072 DVSS.t106 VSS 0.203828f
C6073 DVSS.t44 VSS 0.203828f
C6074 DVSS.n6206 VSS 0.407656f
C6075 DVSS.n6207 VSS 0.073484f
C6076 DVSS.n6208 VSS 0.176594f
C6077 DVSS.n6209 VSS 0.009721f
C6078 DVSS.n6210 VSS 0.018031f
C6079 DVSS.n6211 VSS 0.009721f
C6080 DVSS.n6212 VSS 0.019442f
C6081 DVSS.n6213 VSS 0.009721f
C6082 DVSS.n6214 VSS 0.010505f
C6083 DVSS.n6215 VSS 0.009721f
C6084 DVSS.n6216 VSS 0.019442f
C6085 DVSS.n6217 VSS 0.009721f
C6086 DVSS.n6218 VSS 0.018658f
C6087 DVSS.n6219 VSS 0.009721f
C6088 DVSS.n6220 VSS 0.176594f
C6089 DVSS.n6221 VSS 0.073484f
C6090 DVSS.n6222 VSS 0.026052f
C6091 DVSS.n6223 VSS 0.07508f
C6092 DVSS.n6224 VSS 0.052214f
C6093 DVSS.n6225 VSS 0.174976f
C6094 DVSS.n6226 VSS 0.009721f
C6095 DVSS.n6227 VSS 0.010505f
C6096 DVSS.n6228 VSS 0.009878f
C6097 DVSS.n6229 VSS 0.166982f
C6098 DVSS.n6230 VSS 0.019442f
C6099 DVSS.n6231 VSS 0.019442f
C6100 DVSS.n6232 VSS 0.166982f
C6101 DVSS.n6233 VSS 0.025871f
C6102 DVSS.n6234 VSS 0.054406f
C6103 DVSS.n6235 VSS 0.174976f
C6104 DVSS.n6236 VSS 0.096899f
C6105 DVSS.n6237 VSS 0.025871f
C6106 DVSS.n6238 VSS 0.166982f
C6107 DVSS.n6239 VSS 0.019442f
C6108 DVSS.n6240 VSS 0.009721f
C6109 DVSS.n6241 VSS 0.166982f
C6110 DVSS.n6242 VSS 0.019285f
C6111 DVSS.n6243 VSS 0.052214f
C6112 DVSS.n6244 VSS 0.174976f
C6113 DVSS.n6245 VSS 0.07508f
C6114 DVSS.t138 VSS 0.203828f
C6115 DVSS.t72 VSS 0.203828f
C6116 DVSS.n6246 VSS 0.407656f
C6117 DVSS.n6247 VSS 0.073484f
C6118 DVSS.n6248 VSS 0.176594f
C6119 DVSS.n6249 VSS 0.009721f
C6120 DVSS.n6250 VSS 0.019285f
C6121 DVSS.n6251 VSS 0.009721f
C6122 DVSS.n6252 VSS 0.019442f
C6123 DVSS.n6253 VSS 0.019442f
C6124 DVSS.n6254 VSS 0.009721f
C6125 DVSS.n6255 VSS 0.015052f
C6126 DVSS.n6256 VSS 0.013798f
C6127 DVSS.n6257 VSS 0.170933f
C6128 DVSS.n6258 VSS 0.021951f
C6129 DVSS.n6259 VSS 0.023205f
C6130 DVSS.n6260 VSS 0.019442f
C6131 DVSS.n6261 VSS 0.009721f
C6132 DVSS.n6262 VSS 0.011132f
C6133 DVSS.n6263 VSS 0.052206f
C6134 DVSS.n6264 VSS 0.026052f
C6135 DVSS.n6265 VSS 0.009721f
C6136 DVSS.n6266 VSS 0.052214f
C6137 DVSS.n6267 VSS 0.174976f
C6138 DVSS.n6268 VSS 0.07508f
C6139 DVSS.t82 VSS 0.203828f
C6140 DVSS.t158 VSS 0.203828f
C6141 DVSS.n6269 VSS 0.407656f
C6142 DVSS.n6270 VSS 0.073484f
C6143 DVSS.n6271 VSS 0.176594f
C6144 DVSS.n6272 VSS 0.009721f
C6145 DVSS.n6273 VSS 0.018031f
C6146 DVSS.n6274 VSS 0.052206f
C6147 DVSS.n6275 VSS 0.026052f
C6148 DVSS.n6276 VSS 0.009721f
C6149 DVSS.n6277 VSS 0.052214f
C6150 DVSS.n6278 VSS 0.174976f
C6151 DVSS.n6279 VSS 0.07508f
C6152 DVSS.t96 VSS 0.203828f
C6153 DVSS.t182 VSS 0.203828f
C6154 DVSS.n6280 VSS 0.407656f
C6155 DVSS.n6281 VSS 0.073484f
C6156 DVSS.n6282 VSS 0.176594f
C6157 DVSS.n6283 VSS 0.009721f
C6158 DVSS.n6284 VSS 0.018658f
C6159 DVSS.n6285 VSS 0.052206f
C6160 DVSS.n6286 VSS 0.026052f
C6161 DVSS.t114 VSS 0.203828f
C6162 DVSS.t34 VSS 0.203828f
C6163 DVSS.n6287 VSS 0.407656f
C6164 DVSS.n6288 VSS 0.073484f
C6165 DVSS.n6289 VSS 0.176594f
C6166 DVSS.n6290 VSS 0.009721f
C6167 DVSS.n6291 VSS 0.019285f
C6168 DVSS.n6292 VSS 0.009721f
C6169 DVSS.n6293 VSS 0.009721f
C6170 DVSS.n6294 VSS 0.166982f
C6171 DVSS.n6295 VSS 0.009721f
C6172 DVSS.n6296 VSS 0.017717f
C6173 DVSS.n6297 VSS 0.166982f
C6174 DVSS.n6298 VSS 0.196381f
C6175 DVSS.n6299 VSS 0.333965f
C6176 DVSS.n6300 VSS 0.333965f
C6177 DVSS.n6301 VSS 0.333965f
C6178 DVSS.n6302 VSS 0.333965f
C6179 DVSS.n6303 VSS 0.333965f
C6180 DVSS.n6304 VSS 0.333965f
C6181 DVSS.n6305 VSS 0.333965f
C6182 DVSS.n6306 VSS 0.333965f
C6183 DVSS.n6307 VSS 0.333965f
C6184 DVSS.n6308 VSS 0.333965f
C6185 DVSS.n6309 VSS 0.333965f
C6186 DVSS.n6310 VSS 0.333965f
C6187 DVSS.n6311 VSS 0.333965f
C6188 DVSS.n6312 VSS 0.333965f
C6189 DVSS.n6313 VSS 0.333965f
C6190 DVSS.n6314 VSS 0.333965f
C6191 DVSS.n6315 VSS 0.333965f
C6192 DVSS.n6316 VSS 0.333965f
C6193 DVSS.n6317 VSS 0.333965f
C6194 DVSS.n6318 VSS 0.333965f
C6195 DVSS.n6319 VSS 0.333965f
C6196 DVSS.n6320 VSS 0.333965f
C6197 DVSS.n6321 VSS 0.333965f
C6198 DVSS.n6322 VSS 0.333965f
C6199 DVSS.n6323 VSS 0.333965f
C6200 DVSS.n6324 VSS 0.333965f
C6201 DVSS.n6325 VSS 0.333965f
C6202 DVSS.n6326 VSS 0.333965f
C6203 DVSS.n6327 VSS 0.333965f
C6204 DVSS.n6328 VSS 0.333965f
C6205 DVSS.n6329 VSS 0.333965f
C6206 DVSS.n6330 VSS 0.333965f
C6207 DVSS.n6331 VSS 0.333965f
C6208 DVSS.n6332 VSS 0.333965f
C6209 DVSS.n6333 VSS 0.333965f
C6210 DVSS.n6334 VSS 0.333965f
C6211 DVSS.n6335 VSS 0.333965f
C6212 DVSS.n6336 VSS 0.333965f
C6213 DVSS.n6337 VSS 0.333965f
C6214 DVSS.n6338 VSS 0.333965f
C6215 DVSS.n6339 VSS 0.333965f
C6216 DVSS.n6340 VSS 0.333965f
C6217 DVSS.n6341 VSS 0.333965f
C6218 DVSS.n6342 VSS 0.333965f
C6219 DVSS.n6343 VSS 0.333965f
C6220 DVSS.n6344 VSS 0.333965f
C6221 DVSS.n6345 VSS 0.333965f
C6222 DVSS.n6346 VSS 0.296335f
C6223 DVSS.n6347 VSS 0.296335f
C6224 DVSS.n6348 VSS 0.637355f
C6225 DVSS.n6349 VSS 0.204612f
C6226 DVSS.n6350 VSS 0.204612f
C6227 DVSS.n6351 VSS 0.333965f
C6228 DVSS.n6352 VSS 0.333965f
C6229 DVSS.n6353 VSS 0.333965f
C6230 DVSS.n6354 VSS 0.333965f
C6231 DVSS.n6355 VSS 0.333965f
C6232 DVSS.n6356 VSS 0.333965f
C6233 DVSS.n6357 VSS 0.333965f
C6234 DVSS.n6358 VSS 0.333965f
C6235 DVSS.n6359 VSS 0.333965f
C6236 DVSS.n6360 VSS 0.333965f
C6237 DVSS.n6361 VSS 0.333965f
C6238 DVSS.n6362 VSS 0.333965f
C6239 DVSS.n6363 VSS 0.333965f
C6240 DVSS.n6364 VSS 0.333965f
C6241 DVSS.n6365 VSS 0.333965f
C6242 DVSS.n6366 VSS 0.196381f
C6243 DVSS.n6371 VSS 0.166982f
C6244 DVSS.n6372 VSS 0.052105f
C6245 DVSS.n6373 VSS 0.166982f
C6246 DVSS.n6374 VSS 0.047482f
C6247 DVSS.n6375 VSS 0.073115f
C6248 DVSS.n6376 VSS 0.07508f
C6249 DVSS.t154 VSS 0.203828f
C6250 DVSS.t46 VSS 0.203828f
C6251 DVSS.n6377 VSS 0.407656f
C6252 DVSS.n6378 VSS 0.073484f
C6253 DVSS.n6379 VSS 0.176594f
C6254 DVSS.n6380 VSS 0.069767f
C6255 DVSS.n6381 VSS 0.029006f
C6256 DVSS.n6382 VSS 0.018972f
C6257 DVSS.n6383 VSS 0.009721f
C6258 DVSS.n6384 VSS 0.026052f
C6259 DVSS.n6385 VSS 0.009721f
C6260 DVSS.n6386 VSS 0.052214f
C6261 DVSS.n6387 VSS 0.174976f
C6262 DVSS.n6388 VSS 0.07508f
C6263 DVSS.t170 VSS 0.203828f
C6264 DVSS.t62 VSS 0.203828f
C6265 DVSS.n6389 VSS 0.407656f
C6266 DVSS.n6390 VSS 0.073484f
C6267 DVSS.n6391 VSS 0.176594f
C6268 DVSS.n6392 VSS 0.052206f
C6269 DVSS.n6393 VSS 0.018972f
C6270 DVSS.n6394 VSS 0.009721f
C6271 DVSS.n6395 VSS 0.009721f
C6272 DVSS.n6396 VSS 0.009721f
C6273 DVSS.n6397 VSS 0.167516f
C6274 DVSS.n6398 VSS 0.014566f
C6275 DVSS.n6399 VSS 0.094729f
C6276 DVSS.n6400 VSS 0.167535f
C6277 DVSS.n6401 VSS 0.011446f
C6278 DVSS.n6402 VSS 0.052206f
C6279 DVSS.n6403 VSS 0.009721f
C6280 DVSS.n6404 VSS 0.176594f
C6281 DVSS.n6405 VSS 0.073484f
C6282 DVSS.n6406 VSS 0.026052f
C6283 DVSS.n6407 VSS 0.07508f
C6284 DVSS.n6408 VSS 0.009721f
C6285 DVSS.n6409 VSS 0.174976f
C6286 DVSS.n6410 VSS 0.052214f
C6287 DVSS.n6411 VSS 0.009721f
C6288 DVSS.n6412 VSS 0.017717f
C6289 DVSS.n6413 VSS 0.009721f
C6290 DVSS.n6414 VSS 0.174976f
C6291 DVSS.n6415 VSS 0.052214f
C6292 DVSS.n6416 VSS 0.009721f
C6293 DVSS.n6417 VSS 0.01709f
C6294 DVSS.n6418 VSS 0.009721f
C6295 DVSS.n6419 VSS 0.009721f
C6296 DVSS.n6420 VSS 0.01662f
C6297 DVSS.n6421 VSS 0.167535f
C6298 DVSS.n6422 VSS 0.094729f
C6299 DVSS.n6423 VSS 0.341867f
C6300 DVSS.n6424 VSS 0.014566f
C6301 DVSS.n6425 VSS 1.00544f
C6302 DVSS.n6426 VSS 1.8361f
C6303 DVSS.n6427 VSS -1.94838f
C6304 DVSS.n6428 VSS -2.38582f
C6305 DVSS.n6429 VSS -1.94838f
C6306 DVSS.n6430 VSS 1.8346f
C6307 DVSS.n6431 VSS 1.00693f
C6308 DVSS.n6432 VSS 0.009721f
C6309 DVSS.n6433 VSS 0.341867f
C6310 DVSS.n6434 VSS 0.009721f
C6311 DVSS.n6435 VSS 0.341867f
C6312 DVSS.n6437 VSS 0.014566f
C6313 DVSS.n6438 VSS 0.094729f
C6314 DVSS.n6439 VSS 0.167535f
C6315 DVSS.n6440 VSS 0.012073f
C6316 DVSS.n6441 VSS 0.009721f
C6317 DVSS.n6442 VSS 0.176594f
C6318 DVSS.t172 VSS 0.203828f
C6319 DVSS.t148 VSS 0.203828f
C6320 DVSS.n6443 VSS 0.407656f
C6321 DVSS.n6444 VSS 0.073484f
C6322 DVSS.n6445 VSS 0.026052f
C6323 DVSS.n6446 VSS 0.045802f
C6324 DVSS.n6448 VSS 0.052105f
C6325 DVSS.n6456 VSS 0.158751f
C6326 DVSS.n6458 VSS 0.052105f
C6327 DVSS.n6459 VSS 0.229429f
C6328 DVSS.n6460 VSS 0.166982f
C6329 DVSS.n6461 VSS 0.040339f
C6330 DVSS.n6462 VSS 0.026052f
C6331 DVSS.n6463 VSS 0.342732f
C6332 DVSS.n6464 VSS 0.026052f
C6333 DVSS.n6465 VSS 0.342732f
C6334 DVSS.n6467 VSS 0.342732f
C6335 DVSS.n6468 VSS 0.009721f
C6336 DVSS.n6469 VSS 0.01662f
C6337 DVSS.n6470 VSS 0.167535f
C6338 DVSS.n6471 VSS 0.008467f
C6339 DVSS.n6472 VSS 0.167516f
C6340 DVSS.n6473 VSS 0.029006f
C6341 DVSS.n6474 VSS 0.027282f
C6342 DVSS.n6475 VSS 0.017717f
C6343 DVSS.n6476 VSS 0.166982f
C6344 DVSS.n6477 VSS 0.010819f
C6345 DVSS.n6478 VSS 0.009721f
C6346 DVSS.n6479 VSS 0.166982f
C6347 DVSS.n6480 VSS 0.019285f
C6348 DVSS.n6481 VSS 0.009721f
C6349 DVSS.n6482 VSS 0.174976f
C6350 DVSS.n6483 VSS 0.052214f
C6351 DVSS.n6484 VSS 0.019285f
C6352 DVSS.n6485 VSS 0.009721f
C6353 DVSS.n6486 VSS 0.166982f
C6354 DVSS.n6487 VSS 0.009721f
C6355 DVSS.n6488 VSS 0.017717f
C6356 DVSS.n6489 VSS 0.166982f
C6357 DVSS.n6490 VSS 0.010819f
C6358 DVSS.n6491 VSS 0.052214f
C6359 DVSS.n6492 VSS 0.174976f
C6360 DVSS.n6493 VSS 0.07508f
C6361 DVSS.t140 VSS 0.203828f
C6362 DVSS.t76 VSS 0.203828f
C6363 DVSS.n6494 VSS 0.407656f
C6364 DVSS.n6495 VSS 0.073484f
C6365 DVSS.n6496 VSS 0.176594f
C6366 DVSS.n6497 VSS 0.052206f
C6367 DVSS.n6498 VSS 0.010819f
C6368 DVSS.n6499 VSS 0.009721f
C6369 DVSS.n6500 VSS 0.166982f
C6370 DVSS.n6501 VSS 0.273992f
C6371 DVSS.n6502 VSS 0.333965f
C6372 DVSS.n6503 VSS 0.333965f
C6373 DVSS.n6504 VSS 0.333965f
C6374 DVSS.n6505 VSS 0.195205f
C6375 DVSS.n6506 VSS 0.195205f
C6376 DVSS.n6507 VSS 0.109362f
C6377 DVSS.n6508 VSS 0.637355f
C6378 DVSS.n6509 VSS 0.305742f
C6379 DVSS.n6510 VSS 0.305742f
C6380 DVSS.n6511 VSS 0.305742f
C6381 DVSS.n6512 VSS 0.333965f
C6382 DVSS.n6513 VSS 0.333965f
C6383 DVSS.n6514 VSS 0.333965f
C6384 DVSS.n6515 VSS 0.333965f
C6385 DVSS.n6516 VSS 0.333965f
C6386 DVSS.n6517 VSS 0.333965f
C6387 DVSS.n6518 VSS 0.333965f
C6388 DVSS.n6519 VSS 0.333965f
C6389 DVSS.n6520 VSS 0.333965f
C6390 DVSS.n6521 VSS 0.333965f
C6391 DVSS.n6522 VSS 0.333965f
C6392 DVSS.n6523 VSS 0.333965f
C6393 DVSS.n6524 VSS 0.333965f
C6394 DVSS.n6525 VSS 0.333965f
C6395 DVSS.n6526 VSS 0.333965f
C6396 DVSS.n6527 VSS 0.333965f
C6397 DVSS.n6528 VSS 0.333965f
C6398 DVSS.n6529 VSS 0.252825f
C6399 DVSS.n6530 VSS 0.333965f
C6400 DVSS.n6531 VSS 0.333965f
C6401 DVSS.n6532 VSS 0.333965f
C6402 DVSS.n6533 VSS 0.215195f
C6403 DVSS.n6534 VSS 1.24454f
C6404 DVDD.n0 VSS 0.05145f
C6405 DVDD.n1 VSS 0.064086f
C6406 DVDD.n2 VSS 0.128173f
C6407 DVDD.n3 VSS 0.128173f
C6408 DVDD.n4 VSS 0.376435f
C6409 DVDD.n9 VSS 0.151899f
C6410 DVDD.n11 VSS 0.882607f
C6411 DVDD.n12 VSS 0.151899f
C6412 DVDD.n13 VSS 0.075949f
C6413 DVDD.n14 VSS 0.064086f
C6414 DVDD.n15 VSS 0.064086f
C6415 DVDD.n16 VSS 0.057317f
C6416 DVDD.n17 VSS 0.064086f
C6417 DVDD.n18 VSS 0.064086f
C6418 DVDD.n20 VSS 0.055963f
C6419 DVDD.n22 VSS 0.06183f
C6420 DVDD.n23 VSS 0.064086f
C6421 DVDD.n24 VSS 0.064086f
C6422 DVDD.n25 VSS 0.062732f
C6423 DVDD.n26 VSS 0.064086f
C6424 DVDD.n27 VSS 0.103351f
C6425 DVDD.n29 VSS 0.151899f
C6426 DVDD.n30 VSS 1.27644f
C6427 DVDD.n31 VSS 0.151899f
C6428 DVDD.n32 VSS 0.151899f
C6429 DVDD.n33 VSS 0.128173f
C6430 DVDD.n34 VSS 0.055963f
C6431 DVDD.n35 VSS 0.128173f
C6432 DVDD.n36 VSS 0.128173f
C6433 DVDD.n37 VSS 0.128173f
C6434 DVDD.n38 VSS 0.11012f
C6435 DVDD.n39 VSS 0.128173f
C6436 DVDD.n40 VSS 0.128173f
C6437 DVDD.n41 VSS 0.128173f
C6438 DVDD.n42 VSS 0.064086f
C6439 DVDD.n43 VSS 0.159926f
C6440 DVDD.n44 VSS 0.163891f
C6441 DVDD.n45 VSS 0.124901f
C6442 DVDD.n46 VSS 0.163891f
C6443 DVDD.n47 VSS 0.163891f
C6444 DVDD.n49 VSS 1.37721f
C6445 DVDD.n51 VSS 0.163891f
C6446 DVDD.n52 VSS 0.120936f
C6447 DVDD.n54 VSS 0.163891f
C6448 DVDD.n56 VSS 0.163891f
C6449 DVDD.n57 VSS 0.159926f
C6450 DVDD.n58 VSS 0.059573f
C6451 DVDD.n59 VSS 0.064086f
C6452 DVDD.n60 VSS 0.064086f
C6453 DVDD.n61 VSS 0.064086f
C6454 DVDD.n62 VSS 0.058671f
C6455 DVDD.n63 VSS 0.064086f
C6456 DVDD.n64 VSS 0.055963f
C6457 DVDD.n65 VSS 0.064086f
C6458 DVDD.n66 VSS 0.081946f
C6459 DVDD.n71 VSS 0.064086f
C6460 DVDD.n73 VSS 0.061379f
C6461 DVDD.n74 VSS 0.064086f
C6462 DVDD.n75 VSS 0.064086f
C6463 DVDD.n76 VSS 0.064086f
C6464 DVDD.n78 VSS 0.060476f
C6465 DVDD.n79 VSS 0.075821f
C6466 DVDD.n80 VSS 0.128173f
C6467 DVDD.n81 VSS 0.055963f
C6468 DVDD.n82 VSS 0.128173f
C6469 DVDD.n83 VSS 0.128173f
C6470 DVDD.n84 VSS 0.128173f
C6471 DVDD.n85 VSS 0.064086f
C6472 DVDD.n86 VSS 0.128173f
C6473 DVDD.n87 VSS 0.128173f
C6474 DVDD.n88 VSS 0.128173f
C6475 DVDD.n89 VSS 0.064086f
C6476 DVDD.n90 VSS 0.159926f
C6477 DVDD.n93 VSS 0.055963f
C6478 DVDD.n96 VSS 0.120936f
C6479 DVDD.n97 VSS 0.159926f
C6480 DVDD.n98 VSS 0.064086f
C6481 DVDD.n99 VSS 0.063184f
C6482 DVDD.n100 VSS 0.064086f
C6483 DVDD.n101 VSS 0.064086f
C6484 DVDD.n102 VSS 0.064086f
C6485 DVDD.n103 VSS 0.062281f
C6486 DVDD.n104 VSS 0.081946f
C6487 DVDD.n105 VSS 0.055963f
C6488 DVDD.n106 VSS 0.057768f
C6489 DVDD.n107 VSS 0.064086f
C6490 DVDD.n108 VSS 0.064086f
C6491 DVDD.n109 VSS 0.064086f
C6492 DVDD.n110 VSS 0.056865f
C6493 DVDD.n111 VSS 0.064086f
C6494 DVDD.n112 VSS 0.095678f
C6495 DVDD.n113 VSS 0.163891f
C6496 DVDD.n114 VSS 0.124901f
C6497 DVDD.n116 VSS 0.163891f
C6498 DVDD.n117 VSS 0.163891f
C6499 DVDD.n118 VSS 0.055963f
C6500 DVDD.n121 VSS 0.163891f
C6501 DVDD.n122 VSS 0.261596f
C6502 DVDD.n123 VSS 0.11992f
C6503 DVDD.n124 VSS 0.036277f
C6504 DVDD.n125 VSS 0.163891f
C6505 DVDD.n126 VSS 0.261596f
C6506 DVDD.n127 VSS 0.11992f
C6507 DVDD.n128 VSS 1.20049f
C6508 DVDD.n129 VSS 0.151899f
C6509 DVDD.n130 VSS 0.081467f
C6510 DVDD.n131 VSS 0.038965f
C6511 DVDD.n132 VSS 0.085784f
C6512 DVDD.n133 VSS 0.037455f
C6513 DVDD.n134 VSS 0.042891f
C6514 DVDD.n135 VSS 0.165886f
C6515 DVDD.n136 VSS 0.163891f
C6516 DVDD.n137 VSS 0.151899f
C6517 DVDD.n138 VSS 0.034496f
C6518 DVDD.n139 VSS 0.11992f
C6519 DVDD.n140 VSS 0.015989f
C6520 DVDD.n141 VSS 0.015989f
C6521 DVDD.n142 VSS 0.11992f
C6522 DVDD.n143 VSS 0.034496f
C6523 DVDD.n144 VSS 0.11992f
C6524 DVDD.n145 VSS 0.163891f
C6525 DVDD.n146 VSS 0.11992f
C6526 DVDD.n147 VSS 0.165353f
C6527 DVDD.n148 VSS 0.11992f
C6528 DVDD.n149 VSS 0.11992f
C6529 DVDD.n150 VSS 0.163891f
C6530 DVDD.n151 VSS 0.11992f
C6531 DVDD.n152 VSS 0.015989f
C6532 DVDD.n153 VSS 0.015989f
C6533 DVDD.n154 VSS 0.11992f
C6534 DVDD.n155 VSS 0.037455f
C6535 DVDD.n156 VSS 0.163891f
C6536 DVDD.n157 VSS 0.151899f
C6537 DVDD.n158 VSS 0.151899f
C6538 DVDD.n159 VSS 0.042891f
C6539 DVDD.n160 VSS 0.11992f
C6540 DVDD.n161 VSS 0.01831f
C6541 DVDD.n162 VSS 0.137328f
C6542 DVDD.n163 VSS 0.01831f
C6543 DVDD.n164 VSS 0.137328f
C6544 DVDD.n165 VSS 0.163891f
C6545 DVDD.n166 VSS 0.137328f
C6546 DVDD.n167 VSS 0.274656f
C6547 DVDD.n168 VSS 0.274656f
C6548 DVDD.n169 VSS 0.274656f
C6549 DVDD.n170 VSS 0.456471f
C6550 DVDD.n171 VSS 0.333649f
C6551 DVDD.n172 VSS 0.333649f
C6552 DVDD.n173 VSS 0.11992f
C6553 DVDD.n174 VSS 0.274656f
C6554 DVDD.n175 VSS 0.202124f
C6555 DVDD.n176 VSS 0.11992f
C6556 DVDD.n177 VSS 0.11992f
C6557 DVDD.n178 VSS 0.02695f
C6558 DVDD.n179 VSS 0.039569f
C6559 DVDD.n180 VSS 0.06313f
C6560 DVDD.n181 VSS 0.209861f
C6561 DVDD.n182 VSS 0.027981f
C6562 DVDD.n183 VSS 0.058144f
C6563 DVDD.n184 VSS 0.06037f
C6564 DVDD.n185 VSS 0.202124f
C6565 DVDD.n186 VSS 0.209861f
C6566 DVDD.n187 VSS 0.163932f
C6567 DVDD.n188 VSS 0.209861f
C6568 DVDD.n189 VSS 0.202124f
C6569 DVDD.n190 VSS 0.165883f
C6570 DVDD.n191 VSS 0.02695f
C6571 DVDD.n192 VSS 0.027981f
C6572 DVDD.n193 VSS 0.202124f
C6573 DVDD.n194 VSS 0.11992f
C6574 DVDD.n195 VSS 0.274656f
C6575 DVDD.n196 VSS 1.0087f
C6576 DVDD.n197 VSS 0.274656f
C6577 DVDD.n198 VSS 0.11992f
C6578 DVDD.n199 VSS 0.11992f
C6579 DVDD.n200 VSS 0.325912f
C6580 DVDD.n201 VSS 0.440997f
C6581 DVDD.n202 VSS 0.274656f
C6582 DVDD.n203 VSS 0.11992f
C6583 DVDD.n204 VSS 0.11992f
C6584 DVDD.n205 VSS 0.11992f
C6585 DVDD.n206 VSS 0.209861f
C6586 DVDD.n207 VSS 0.06037f
C6587 DVDD.n208 VSS 0.058144f
C6588 DVDD.n209 VSS 0.027981f
C6589 DVDD.n210 VSS 0.202124f
C6590 DVDD.n211 VSS 0.209861f
C6591 DVDD.n212 VSS 0.02695f
C6592 DVDD.n213 VSS 0.06313f
C6593 DVDD.n214 VSS 0.209861f
C6594 DVDD.n215 VSS 0.202124f
C6595 DVDD.n216 VSS 0.027981f
C6596 DVDD.n217 VSS 0.165353f
C6597 DVDD.n218 VSS 0.164489f
C6598 DVDD.n219 VSS 0.202124f
C6599 DVDD.n220 VSS 0.02695f
C6600 DVDD.n221 VSS 0.209861f
C6601 DVDD.n222 VSS 0.274656f
C6602 DVDD.n223 VSS 0.744772f
C6603 DVDD.n224 VSS 0.11992f
C6604 DVDD.n225 VSS 0.11992f
C6605 DVDD.n226 VSS 0.11992f
C6606 DVDD.n227 VSS 0.274656f
C6607 DVDD.n228 VSS 0.122822f
C6608 DVDD.n229 VSS 0.296448f
C6609 DVDD.n230 VSS 0.163891f
C6610 DVDD.n231 VSS 0.319852f
C6611 DVDD.n232 VSS 0.036964f
C6612 DVDD.n233 VSS 0.122822f
C6613 DVDD.n234 VSS 0.277343f
C6614 DVDD.n235 VSS 0.163891f
C6615 DVDD.n236 VSS 0.064086f
C6616 DVDD.n238 VSS 0.064086f
C6617 DVDD.n239 VSS 0.064086f
C6618 DVDD.n240 VSS 0.064086f
C6619 DVDD.n241 VSS 0.060476f
C6620 DVDD.n242 VSS 0.064086f
C6621 DVDD.n243 VSS 0.064086f
C6622 DVDD.n244 VSS 0.064086f
C6623 DVDD.n245 VSS 0.059573f
C6624 DVDD.n246 VSS 0.064086f
C6625 DVDD.n247 VSS 0.064086f
C6626 DVDD.n248 VSS 0.064086f
C6627 DVDD.n249 VSS 0.058671f
C6628 DVDD.n250 VSS 0.064086f
C6629 DVDD.n251 VSS 0.055963f
C6630 DVDD.n252 VSS 0.163891f
C6631 DVDD.n253 VSS 0.163891f
C6632 DVDD.n254 VSS 0.163891f
C6633 DVDD.n255 VSS 0.163891f
C6634 DVDD.n256 VSS 0.163891f
C6635 DVDD.n257 VSS 0.093873f
C6636 DVDD.n260 VSS 3.48797f
C6637 DVDD.n262 VSS 0.163891f
C6638 DVDD.n264 VSS 0.163891f
C6639 DVDD.n266 VSS 0.163891f
C6640 DVDD.n272 VSS 0.055963f
C6641 DVDD.n273 VSS 0.128173f
C6642 DVDD.n274 VSS 0.055963f
C6643 DVDD.n275 VSS 0.128173f
C6644 DVDD.n276 VSS 0.128173f
C6645 DVDD.n277 VSS 0.128173f
C6646 DVDD.n278 VSS 0.128173f
C6647 DVDD.n279 VSS 0.128173f
C6648 DVDD.n280 VSS 0.128173f
C6649 DVDD.n281 VSS 0.128173f
C6650 DVDD.n282 VSS 0.128173f
C6651 DVDD.n283 VSS 0.128173f
C6652 DVDD.n284 VSS 0.128173f
C6653 DVDD.n290 VSS 0.055963f
C6654 DVDD.n293 VSS 0.064086f
C6655 DVDD.n294 VSS 0.064086f
C6656 DVDD.n295 VSS 0.064086f
C6657 DVDD.n297 VSS 0.064086f
C6658 DVDD.n298 VSS 3.48797f
C6659 DVDD.n299 VSS 0.064086f
C6660 DVDD.n300 VSS 0.064086f
C6661 DVDD.n301 VSS 0.064086f
C6662 DVDD.n302 VSS 0.064086f
C6663 DVDD.n303 VSS 0.064086f
C6664 DVDD.n304 VSS 0.055963f
C6665 DVDD.n305 VSS 0.163891f
C6666 DVDD.n306 VSS 0.163891f
C6667 DVDD.n307 VSS 0.163891f
C6668 DVDD.n308 VSS 0.163891f
C6669 DVDD.n309 VSS 0.163891f
C6670 DVDD.n310 VSS 0.090263f
C6671 DVDD.n311 VSS 0.163891f
C6672 DVDD.n312 VSS 0.163891f
C6673 DVDD.n313 VSS 0.163891f
C6674 DVDD.n314 VSS 0.163891f
C6675 DVDD.n315 VSS 0.319852f
C6676 DVDD.n320 VSS 0.064086f
C6677 DVDD.n321 VSS 0.057768f
C6678 DVDD.n322 VSS 0.056865f
C6679 DVDD.n323 VSS 0.063184f
C6680 DVDD.n324 VSS 0.055963f
C6681 DVDD.n325 VSS 0.128173f
C6682 DVDD.n326 VSS 0.055963f
C6683 DVDD.n327 VSS 0.128173f
C6684 DVDD.n328 VSS 0.128173f
C6685 DVDD.n329 VSS 0.055963f
C6686 DVDD.n330 VSS 0.128173f
C6687 DVDD.n331 VSS 0.128173f
C6688 DVDD.n332 VSS 0.128173f
C6689 DVDD.n333 VSS 0.055963f
C6690 DVDD.n334 VSS 0.128173f
C6691 DVDD.n335 VSS 0.055963f
C6692 DVDD.n336 VSS 0.128173f
C6693 DVDD.n337 VSS 0.055963f
C6694 DVDD.n338 VSS 0.128173f
C6695 DVDD.n339 VSS 0.128173f
C6696 DVDD.n340 VSS 0.128173f
C6697 DVDD.n341 VSS 0.128173f
C6698 DVDD.n342 VSS 0.055963f
C6699 DVDD.n343 VSS 0.128173f
C6700 DVDD.n344 VSS 0.055963f
C6701 DVDD.n345 VSS 0.128173f
C6702 DVDD.n346 VSS 0.055963f
C6703 DVDD.n347 VSS 0.128173f
C6704 DVDD.n348 VSS 0.128173f
C6705 DVDD.n349 VSS 0.128173f
C6706 DVDD.n350 VSS 0.128173f
C6707 DVDD.n351 VSS 0.128173f
C6708 DVDD.n352 VSS 0.128173f
C6709 DVDD.n353 VSS 0.128173f
C6710 DVDD.n354 VSS 0.128173f
C6711 DVDD.n355 VSS 0.163891f
C6712 DVDD.n356 VSS 0.163891f
C6713 DVDD.n357 VSS 0.163891f
C6714 DVDD.n358 VSS 0.163891f
C6715 DVDD.n359 VSS 0.163891f
C6716 DVDD.n360 VSS 0.055963f
C6717 DVDD.n361 VSS 3.48797f
C6718 DVDD.n362 VSS 0.163891f
C6719 DVDD.n363 VSS 0.163891f
C6720 DVDD.n364 VSS 0.163891f
C6721 DVDD.n365 VSS 0.163891f
C6722 DVDD.n366 VSS 0.319852f
C6723 DVDD.n372 VSS 0.064086f
C6724 DVDD.n374 VSS 0.061379f
C6725 DVDD.n375 VSS 0.064086f
C6726 DVDD.n376 VSS 0.064086f
C6727 DVDD.n377 VSS 0.064086f
C6728 DVDD.n378 VSS 0.060476f
C6729 DVDD.n380 VSS 0.059573f
C6730 DVDD.n381 VSS 0.064086f
C6731 DVDD.n382 VSS 0.064086f
C6732 DVDD.n383 VSS 0.064086f
C6733 DVDD.n385 VSS 0.058671f
C6734 DVDD.n386 VSS 0.064086f
C6735 DVDD.n387 VSS 0.064086f
C6736 DVDD.n388 VSS 0.055963f
C6737 DVDD.n389 VSS 0.128173f
C6738 DVDD.n390 VSS 0.128173f
C6739 DVDD.n391 VSS 0.128173f
C6740 DVDD.n392 VSS 0.128173f
C6741 DVDD.n393 VSS 0.055963f
C6742 DVDD.n394 VSS 0.128173f
C6743 DVDD.n395 VSS 0.128173f
C6744 DVDD.n396 VSS 0.055963f
C6745 DVDD.n397 VSS 0.128173f
C6746 DVDD.n398 VSS 0.128173f
C6747 DVDD.n399 VSS 0.128173f
C6748 DVDD.n400 VSS 0.128173f
C6749 DVDD.n401 VSS 0.128173f
C6750 DVDD.n402 VSS 0.055963f
C6751 DVDD.n403 VSS 0.128173f
C6752 DVDD.n404 VSS 0.055963f
C6753 DVDD.n405 VSS 0.128173f
C6754 DVDD.n406 VSS 0.055963f
C6755 DVDD.n407 VSS 0.128173f
C6756 DVDD.n408 VSS 0.128173f
C6757 DVDD.n409 VSS 0.128173f
C6758 DVDD.n410 VSS 0.128173f
C6759 DVDD.n411 VSS 0.055963f
C6760 DVDD.n412 VSS 0.128173f
C6761 DVDD.n413 VSS 0.055963f
C6762 DVDD.n414 VSS 0.128173f
C6763 DVDD.n415 VSS 0.055963f
C6764 DVDD.n416 VSS 0.128173f
C6765 DVDD.n417 VSS 0.128173f
C6766 DVDD.n418 VSS 0.128173f
C6767 DVDD.n419 VSS 0.128173f
C6768 DVDD.n420 VSS 0.128173f
C6769 DVDD.n421 VSS 0.055963f
C6770 DVDD.n426 VSS 0.064086f
C6771 DVDD.n427 VSS 0.055963f
C6772 DVDD.n428 VSS 0.128173f
C6773 DVDD.n429 VSS 0.055963f
C6774 DVDD.n430 VSS 0.128173f
C6775 DVDD.n431 VSS 0.128173f
C6776 DVDD.n432 VSS 0.128173f
C6777 DVDD.n433 VSS 0.128173f
C6778 DVDD.n434 VSS 0.128173f
C6779 DVDD.n435 VSS 0.064086f
C6780 DVDD.n436 VSS 0.128173f
C6781 DVDD.n437 VSS 0.128173f
C6782 DVDD.n438 VSS 0.128173f
C6783 DVDD.n439 VSS 0.055963f
C6784 DVDD.n440 VSS 0.064086f
C6785 DVDD.n441 VSS 0.151899f
C6786 DVDD.n442 VSS 0.151899f
C6787 DVDD.n443 VSS 0.151899f
C6788 DVDD.n444 VSS 0.151899f
C6789 DVDD.n445 VSS 0.151899f
C6790 DVDD.n446 VSS 0.055963f
C6791 DVDD.n448 VSS 0.137328f
C6792 DVDD.n449 VSS 0.137328f
C6793 DVDD.n450 VSS 0.137328f
C6794 DVDD.n451 VSS 0.122822f
C6795 DVDD.n452 VSS 0.137328f
C6796 DVDD.n453 VSS 0.137328f
C6797 DVDD.n454 VSS 0.137328f
C6798 DVDD.n455 VSS 0.137328f
C6799 DVDD.n456 VSS 0.134427f
C6800 DVDD.n457 VSS 0.137328f
C6801 DVDD.n458 VSS 0.137328f
C6802 DVDD.n459 VSS 0.110249f
C6803 DVDD.n460 VSS 0.132493f
C6804 DVDD.n461 VSS 0.11992f
C6805 DVDD.n462 VSS 0.151899f
C6806 DVDD.n463 VSS 0.151899f
C6807 DVDD.n464 VSS 0.151899f
C6808 DVDD.n465 VSS 0.151899f
C6809 DVDD.n466 VSS 0.151899f
C6810 DVDD.n467 VSS 0.151899f
C6811 DVDD.n468 VSS 0.151899f
C6812 DVDD.n469 VSS 0.151899f
C6813 DVDD.n470 VSS 0.151899f
C6814 DVDD.n471 VSS 0.151899f
C6815 DVDD.n472 VSS 0.151899f
C6816 DVDD.n474 VSS 0.292773f
C6817 DVDD.n475 VSS 1.29067f
C6818 DVDD.n476 VSS 0.057059f
C6819 DVDD.n477 VSS 0.274656f
C6820 DVDD.n478 VSS 0.11992f
C6821 DVDD.n479 VSS 0.274656f
C6822 DVDD.n480 VSS 0.11992f
C6823 DVDD.n481 VSS 0.274656f
C6824 DVDD.n482 VSS 0.11992f
C6825 DVDD.n483 VSS 0.274656f
C6826 DVDD.n484 VSS 0.11992f
C6827 DVDD.n485 VSS 0.274656f
C6828 DVDD.n486 VSS 0.251446f
C6829 DVDD.n487 VSS 0.160538f
C6830 DVDD.n488 VSS 0.085621f
C6831 DVDD.n489 VSS 0.118115f
C6832 DVDD.n490 VSS 0.21057f
C6833 DVDD.n491 VSS 0.146483f
C6834 DVDD.n492 VSS 0.251446f
C6835 DVDD.n493 VSS 0.21057f
C6836 DVDD.n494 VSS 0.146483f
C6837 DVDD.n495 VSS 0.146483f
C6838 DVDD.n496 VSS 0.073242f
C6839 DVDD.n497 VSS 0.151899f
C6840 DVDD.n498 VSS 0.151899f
C6841 DVDD.n499 VSS 0.151899f
C6842 DVDD.n500 VSS 0.151899f
C6843 DVDD.n501 VSS 0.151899f
C6844 DVDD.n502 VSS 0.063957f
C6845 DVDD.n504 VSS 0.137328f
C6846 DVDD.n505 VSS 0.137328f
C6847 DVDD.n506 VSS 0.137328f
C6848 DVDD.n507 VSS 0.122822f
C6849 DVDD.n508 VSS 0.137328f
C6850 DVDD.n509 VSS 0.137328f
C6851 DVDD.n510 VSS 0.137328f
C6852 DVDD.n511 VSS 0.137328f
C6853 DVDD.n512 VSS 0.134427f
C6854 DVDD.n513 VSS 0.137328f
C6855 DVDD.n514 VSS 0.137328f
C6856 DVDD.n515 VSS 0.110249f
C6857 DVDD.n516 VSS 0.132493f
C6858 DVDD.n517 VSS 0.11992f
C6859 DVDD.n518 VSS 0.151899f
C6860 DVDD.n519 VSS 0.151899f
C6861 DVDD.n520 VSS 0.05145f
C6862 DVDD.n521 VSS 0.06615f
C6863 DVDD.n522 VSS 0.06615f
C6864 DVDD.n523 VSS 0.06615f
C6865 DVDD.n524 VSS 0.06615f
C6866 DVDD.n525 VSS 0.06615f
C6867 DVDD.n526 VSS 0.06615f
C6868 DVDD.n527 VSS 0.132299f
C6869 DVDD.n528 VSS 0.06615f
C6870 DVDD.n529 VSS 0.06615f
C6871 DVDD.n530 VSS 0.745125f
C6872 DVDD.n532 VSS 0.06615f
C6873 DVDD.n533 VSS 0.06615f
C6874 DVDD.n534 VSS 0.06615f
C6875 DVDD.n535 VSS 0.06615f
C6876 DVDD.n536 VSS 0.06615f
C6877 DVDD.n537 VSS 0.06615f
C6878 DVDD.n538 VSS 0.06615f
C6879 DVDD.n539 VSS 0.06615f
C6880 DVDD.n540 VSS 0.0147f
C6881 DVDD.n542 VSS 0.026573f
C6882 DVDD.n543 VSS 0.06125f
C6883 DVDD.n544 VSS 0.035233f
C6884 DVDD.n546 VSS 0.0196f
C6885 DVDD.n549 VSS 0.035233f
C6886 DVDD.n550 VSS 0.098464f
C6887 DVDD.n551 VSS 0.025624f
C6888 DVDD.n552 VSS 0.06615f
C6889 DVDD.n553 VSS 0.025624f
C6890 DVDD.n554 VSS 0.137328f
C6891 DVDD.n555 VSS 0.137328f
C6892 DVDD.n556 VSS 0.122822f
C6893 DVDD.n557 VSS 0.137328f
C6894 DVDD.n558 VSS 0.124756f
C6895 DVDD.n559 VSS 0.137328f
C6896 DVDD.n560 VSS 0.137328f
C6897 DVDD.n561 VSS 0.0686f
C6898 DVDD.n562 VSS 0.137328f
C6899 DVDD.n563 VSS 0.110249f
C6900 DVDD.n564 VSS 0.132493f
C6901 DVDD.n565 VSS 0.808336f
C6902 DVDD.n566 VSS 0.137328f
C6903 DVDD.n567 VSS 0.134427f
C6904 DVDD.n568 VSS 0.137328f
C6905 DVDD.n569 VSS 0.221466f
C6906 DVDD.n570 VSS 0.06615f
C6907 DVDD.n571 VSS 0.06615f
C6908 DVDD.n572 VSS 0.06615f
C6909 DVDD.n573 VSS 0.06615f
C6910 DVDD.n574 VSS 0.06615f
C6911 DVDD.n575 VSS 0.06615f
C6912 DVDD.n576 VSS 0.06615f
C6913 DVDD.n577 VSS 0.06615f
C6914 DVDD.n578 VSS 0.06615f
C6915 DVDD.n579 VSS 0.06615f
C6916 DVDD.n582 VSS 0.06615f
C6917 DVDD.n583 VSS 0.11992f
C6918 DVDD.n584 VSS 0.06615f
C6919 DVDD.n585 VSS 0.06615f
C6920 DVDD.n586 VSS 0.06615f
C6921 DVDD.n587 VSS 0.06615f
C6922 DVDD.n588 VSS 0.132299f
C6923 DVDD.n589 VSS 0.06615f
C6924 DVDD.n590 VSS 0.06615f
C6925 DVDD.n591 VSS 0.06615f
C6926 DVDD.n592 VSS 0.06615f
C6927 DVDD.n593 VSS 0.06615f
C6928 DVDD.n594 VSS 0.075949f
C6929 DVDD.n595 VSS 0.07105f
C6930 DVDD.n596 VSS 0.0735f
C6931 DVDD.n597 VSS 0.025624f
C6932 DVDD.n598 VSS 0.075949f
C6933 DVDD.n599 VSS 0.025624f
C6934 DVDD.n600 VSS 0.075949f
C6935 DVDD.n601 VSS 0.025624f
C6936 DVDD.n602 VSS 0.075949f
C6937 DVDD.n603 VSS 0.025624f
C6938 DVDD.n604 VSS 0.075949f
C6939 DVDD.n605 VSS 0.025624f
C6940 DVDD.n606 VSS 0.075949f
C6941 DVDD.n607 VSS 0.025624f
C6942 DVDD.n608 VSS 0.075949f
C6943 DVDD.n609 VSS 0.025624f
C6944 DVDD.n610 VSS 0.025624f
C6945 DVDD.n611 VSS 0.075949f
C6946 DVDD.n612 VSS 0.025624f
C6947 DVDD.n613 VSS 0.075949f
C6948 DVDD.n614 VSS 0.025624f
C6949 DVDD.n615 VSS 0.075949f
C6950 DVDD.n616 VSS 0.025624f
C6951 DVDD.n617 VSS 0.075949f
C6952 DVDD.n618 VSS 0.025624f
C6953 DVDD.n619 VSS 0.075949f
C6954 DVDD.n620 VSS 0.025624f
C6955 DVDD.n621 VSS 0.075949f
C6956 DVDD.n622 VSS 0.025624f
C6957 DVDD.n623 VSS 0.025624f
C6958 DVDD.n624 VSS 0.0735f
C6959 DVDD.n625 VSS 0.0686f
C6960 DVDD.n626 VSS 0.025624f
C6961 DVDD.n627 VSS 0.075949f
C6962 DVDD.n628 VSS 0.025624f
C6963 DVDD.n629 VSS 0.075949f
C6964 DVDD.n630 VSS 0.025624f
C6965 DVDD.n631 VSS 0.075949f
C6966 DVDD.n632 VSS 0.025624f
C6967 DVDD.n633 VSS 0.075949f
C6968 DVDD.n634 VSS 0.025624f
C6969 DVDD.n635 VSS 0.075949f
C6970 DVDD.n636 VSS 0.025624f
C6971 DVDD.n637 VSS 0.025624f
C6972 DVDD.n638 VSS 0.025624f
C6973 DVDD.n639 VSS 0.06615f
C6974 DVDD.n640 VSS 0.025624f
C6975 DVDD.n641 VSS 0.137328f
C6976 DVDD.n642 VSS 0.137328f
C6977 DVDD.n643 VSS 0.122822f
C6978 DVDD.n644 VSS 0.137328f
C6979 DVDD.n645 VSS 0.124756f
C6980 DVDD.n646 VSS 0.137328f
C6981 DVDD.n647 VSS 0.137328f
C6982 DVDD.n648 VSS 0.075949f
C6983 DVDD.n649 VSS 0.137328f
C6984 DVDD.n650 VSS 0.110249f
C6985 DVDD.n651 VSS 0.132493f
C6986 DVDD.n652 VSS 0.808336f
C6987 DVDD.n653 VSS 0.137328f
C6988 DVDD.n654 VSS 0.134427f
C6989 DVDD.n655 VSS 0.137328f
C6990 DVDD.n656 VSS 0.221466f
C6991 DVDD.n657 VSS 0.06615f
C6992 DVDD.n658 VSS 0.06615f
C6993 DVDD.n659 VSS 0.06615f
C6994 DVDD.n660 VSS 0.06615f
C6995 DVDD.n661 VSS 0.06615f
C6996 DVDD.n662 VSS 0.06615f
C6997 DVDD.n663 VSS 0.06615f
C6998 DVDD.n664 VSS 0.06615f
C6999 DVDD.n665 VSS 0.06615f
C7000 DVDD.n666 VSS 0.06615f
C7001 DVDD.n669 VSS 0.06615f
C7002 DVDD.n670 VSS 0.11992f
C7003 DVDD.n671 VSS 0.06615f
C7004 DVDD.n672 VSS 0.06615f
C7005 DVDD.n673 VSS 0.06615f
C7006 DVDD.n674 VSS 0.06615f
C7007 DVDD.n675 VSS 0.06615f
C7008 DVDD.n676 VSS 0.06615f
C7009 DVDD.n677 VSS 0.06615f
C7010 DVDD.n678 VSS 0.06615f
C7011 DVDD.n679 VSS 0.06615f
C7012 DVDD.n680 VSS 0.06615f
C7013 DVDD.n681 VSS 0.075949f
C7014 DVDD.n682 VSS 0.132299f
C7015 DVDD.n683 VSS 0.075949f
C7016 DVDD.n684 VSS 0.025624f
C7017 DVDD.n685 VSS 0.025624f
C7018 DVDD.n686 VSS 0.0735f
C7019 DVDD.n687 VSS 0.0686f
C7020 DVDD.n688 VSS 0.025624f
C7021 DVDD.n689 VSS 0.075949f
C7022 DVDD.n690 VSS 0.025624f
C7023 DVDD.n691 VSS 0.075949f
C7024 DVDD.n692 VSS 0.025624f
C7025 DVDD.n693 VSS 0.075949f
C7026 DVDD.n694 VSS 0.025624f
C7027 DVDD.n695 VSS 0.075949f
C7028 DVDD.n696 VSS 0.025624f
C7029 DVDD.n697 VSS 0.075949f
C7030 DVDD.n698 VSS 0.025624f
C7031 DVDD.n699 VSS 0.075949f
C7032 DVDD.n700 VSS 0.025624f
C7033 DVDD.n701 VSS 0.025624f
C7034 DVDD.n702 VSS 0.07105f
C7035 DVDD.n703 VSS 0.07105f
C7036 DVDD.n704 VSS 0.025624f
C7037 DVDD.n705 VSS 0.075949f
C7038 DVDD.n706 VSS 0.025624f
C7039 DVDD.n707 VSS 0.075949f
C7040 DVDD.n708 VSS 0.025624f
C7041 DVDD.n709 VSS 0.075949f
C7042 DVDD.n710 VSS 0.025624f
C7043 DVDD.n711 VSS 0.075949f
C7044 DVDD.n712 VSS 0.025624f
C7045 DVDD.n713 VSS 0.075949f
C7046 DVDD.n714 VSS 0.025624f
C7047 DVDD.n715 VSS 0.075949f
C7048 DVDD.n716 VSS 0.025624f
C7049 DVDD.n717 VSS 0.025624f
C7050 DVDD.n718 VSS 0.0686f
C7051 DVDD.n719 VSS 0.0735f
C7052 DVDD.n720 VSS 0.025624f
C7053 DVDD.n721 VSS 0.075949f
C7054 DVDD.n722 VSS 0.025624f
C7055 DVDD.n723 VSS 0.075949f
C7056 DVDD.n724 VSS 0.025624f
C7057 DVDD.n725 VSS 0.075949f
C7058 DVDD.n726 VSS 0.025624f
C7059 DVDD.n727 VSS 0.075949f
C7060 DVDD.n728 VSS 0.025624f
C7061 DVDD.n729 VSS 0.025624f
C7062 DVDD.n730 VSS 0.025624f
C7063 DVDD.n731 VSS 0.124756f
C7064 DVDD.n732 VSS 0.137328f
C7065 DVDD.n733 VSS 0.137328f
C7066 DVDD.n734 VSS 0.137328f
C7067 DVDD.n735 VSS 0.122822f
C7068 DVDD.n736 VSS 0.137328f
C7069 DVDD.n737 VSS 0.137328f
C7070 DVDD.n738 VSS 0.075949f
C7071 DVDD.n739 VSS 0.137328f
C7072 DVDD.n740 VSS 0.137328f
C7073 DVDD.n741 VSS 0.134427f
C7074 DVDD.n742 VSS 0.137328f
C7075 DVDD.n743 VSS 0.137328f
C7076 DVDD.n744 VSS 0.110249f
C7077 DVDD.n745 VSS 0.132493f
C7078 DVDD.n746 VSS 0.11992f
C7079 DVDD.n747 VSS 0.06615f
C7080 DVDD.n748 VSS 0.06615f
C7081 DVDD.n749 VSS 0.06615f
C7082 DVDD.n750 VSS 0.06615f
C7083 DVDD.n751 VSS 0.06615f
C7084 DVDD.n752 VSS 0.06615f
C7085 DVDD.n753 VSS 0.132299f
C7086 DVDD.n754 VSS 0.06615f
C7087 DVDD.n755 VSS 0.06615f
C7088 DVDD.n756 VSS 0.06615f
C7089 DVDD.n757 VSS 0.06615f
C7090 DVDD.n760 VSS 0.06615f
C7091 DVDD.n761 VSS 0.745125f
C7092 DVDD.n762 VSS 0.06615f
C7093 DVDD.n763 VSS 0.06615f
C7094 DVDD.n764 VSS 0.06615f
C7095 DVDD.n765 VSS 0.06615f
C7096 DVDD.n766 VSS 0.06615f
C7097 DVDD.n767 VSS 0.06615f
C7098 DVDD.n768 VSS 0.06615f
C7099 DVDD.n769 VSS 0.06615f
C7100 DVDD.n770 VSS 0.06615f
C7101 DVDD.n771 VSS 0.06615f
C7102 DVDD.n772 VSS 0.075949f
C7103 DVDD.n773 VSS 0.025624f
C7104 DVDD.n774 VSS 0.025624f
C7105 DVDD.n775 VSS 0.025624f
C7106 DVDD.n776 VSS 0.132299f
C7107 DVDD.n777 VSS 0.019218f
C7108 DVDD.n778 VSS 0.132299f
C7109 DVDD.n779 VSS -3.16672f
C7110 DVDD.n780 VSS 0.025624f
C7111 DVDD.n781 VSS 0.132299f
C7112 DVDD.n782 VSS 0.025624f
C7113 DVDD.n783 VSS 0.132299f
C7114 DVDD.n784 VSS 0.025624f
C7115 DVDD.n785 VSS 0.064086f
C7116 DVDD.n786 VSS 0.064086f
C7117 DVDD.n787 VSS 0.057317f
C7118 DVDD.n788 VSS 0.064086f
C7119 DVDD.n789 VSS 0.058219f
C7120 DVDD.n790 VSS 0.064086f
C7121 DVDD.n791 VSS 0.064086f
C7122 DVDD.n792 VSS 0.075949f
C7123 DVDD.n793 VSS 0.064086f
C7124 DVDD.n794 VSS 0.05145f
C7125 DVDD.n795 VSS 0.06183f
C7126 DVDD.n796 VSS 0.37595f
C7127 DVDD.n797 VSS 0.064086f
C7128 DVDD.n798 VSS 0.062732f
C7129 DVDD.n799 VSS 0.064086f
C7130 DVDD.n800 VSS 0.103351f
C7131 DVDD.n801 VSS 0.06615f
C7132 DVDD.n802 VSS 0.06615f
C7133 DVDD.n803 VSS 0.06615f
C7134 DVDD.n804 VSS 0.06615f
C7135 DVDD.n805 VSS 0.055963f
C7136 DVDD.n808 VSS 0.06615f
C7137 DVDD.n809 VSS 0.06615f
C7138 DVDD.n810 VSS 0.06615f
C7139 DVDD.n811 VSS 0.06615f
C7140 DVDD.n812 VSS 0.06615f
C7141 DVDD.n813 VSS 0.075949f
C7142 DVDD.n814 VSS 0.069825f
C7143 DVDD.n815 VSS 0.025624f
C7144 DVDD.n816 VSS 0.075949f
C7145 DVDD.n817 VSS 0.025624f
C7146 DVDD.n818 VSS 0.025624f
C7147 DVDD.n819 VSS 0.074725f
C7148 DVDD.n820 VSS 0.067375f
C7149 DVDD.n821 VSS 0.025624f
C7150 DVDD.n822 VSS 0.075949f
C7151 DVDD.n823 VSS 0.025624f
C7152 DVDD.n824 VSS 0.075949f
C7153 DVDD.n825 VSS 0.025624f
C7154 DVDD.n826 VSS 0.075949f
C7155 DVDD.n827 VSS 0.025624f
C7156 DVDD.n828 VSS 0.075949f
C7157 DVDD.n829 VSS 0.025624f
C7158 DVDD.n830 VSS 0.075949f
C7159 DVDD.n831 VSS 0.025624f
C7160 DVDD.n832 VSS 0.025624f
C7161 DVDD.n833 VSS 0.025624f
C7162 DVDD.n834 VSS 0.132299f
C7163 DVDD.n835 VSS 0.025624f
C7164 DVDD.n836 VSS 0.132299f
C7165 DVDD.n837 VSS 0.025624f
C7166 DVDD.n838 VSS 0.132299f
C7167 DVDD.n839 VSS 0.025624f
C7168 DVDD.n840 VSS 0.132299f
C7169 DVDD.n841 VSS 0.025624f
C7170 DVDD.n842 VSS 0.132299f
C7171 DVDD.n843 VSS 0.025624f
C7172 DVDD.n844 VSS 0.132299f
C7173 DVDD.n845 VSS 0.025624f
C7174 DVDD.n846 VSS 0.132299f
C7175 DVDD.n847 VSS 0.025624f
C7176 DVDD.n848 VSS 0.132299f
C7177 DVDD.n849 VSS 0.025624f
C7178 DVDD.n850 VSS 0.132299f
C7179 DVDD.n851 VSS 0.025624f
C7180 DVDD.n852 VSS 0.132299f
C7181 DVDD.n853 VSS 0.025624f
C7182 DVDD.n854 VSS 0.132299f
C7183 DVDD.n855 VSS 0.025624f
C7184 DVDD.n856 VSS 0.132299f
C7185 DVDD.n857 VSS 0.025624f
C7186 DVDD.n858 VSS 0.132299f
C7187 DVDD.n859 VSS 0.025624f
C7188 DVDD.n860 VSS 0.132299f
C7189 DVDD.n861 VSS 0.025624f
C7190 DVDD.n862 VSS 0.132299f
C7191 DVDD.n863 VSS 0.025624f
C7192 DVDD.n864 VSS 0.132299f
C7193 DVDD.n865 VSS 0.025624f
C7194 DVDD.n866 VSS 0.132299f
C7195 DVDD.n867 VSS 0.025624f
C7196 DVDD.n868 VSS 0.132299f
C7197 DVDD.n869 VSS 0.025624f
C7198 DVDD.n870 VSS 0.132299f
C7199 DVDD.n871 VSS 0.025624f
C7200 DVDD.n872 VSS 0.132299f
C7201 DVDD.n873 VSS 0.025624f
C7202 DVDD.n874 VSS 0.132299f
C7203 DVDD.n875 VSS 0.025624f
C7204 DVDD.n876 VSS 0.132299f
C7205 DVDD.n877 VSS 0.013761f
C7206 DVDD.n878 VSS 0.025624f
C7207 DVDD.n879 VSS 0.025624f
C7208 DVDD.n880 VSS 0.06615f
C7209 DVDD.n882 VSS 0.025624f
C7210 DVDD.n884 VSS 0.06615f
C7211 DVDD.n885 VSS 0.035233f
C7212 DVDD.n886 VSS 0.06615f
C7213 DVDD.n888 VSS 0.098464f
C7214 DVDD.n890 VSS 0.031727f
C7215 DVDD.n891 VSS 0.036879f
C7216 DVDD.n892 VSS 0.106252f
C7217 DVDD.n893 VSS 0.044635f
C7218 DVDD.n894 VSS 0.059058f
C7219 DVDD.n896 VSS 0.284688f
C7220 DVDD.n897 VSS 0.088457f
C7221 DVDD.n898 VSS 0.088457f
C7222 DVDD.n900 VSS 0.048448f
C7223 DVDD.n901 VSS 0.053165f
C7224 DVDD.n902 VSS 0.05956f
C7225 DVDD.n903 VSS 0.060318f
C7226 DVDD.n904 VSS 0.05956f
C7227 DVDD.n905 VSS 0.060318f
C7228 DVDD.n906 VSS 0.522252f
C7229 DVDD.n907 VSS 0.728627f
C7230 DVDD.n908 VSS 0.041931f
C7231 DVDD.n909 VSS 0.038327f
C7232 DVDD.n910 VSS 0.041931f
C7233 DVDD.n911 VSS 0.038327f
C7234 DVDD.n912 VSS 0.028833f
C7235 DVDD.n913 VSS 0.02513f
C7236 DVDD.n914 VSS 0.02513f
C7237 DVDD.n915 VSS 0.433807f
C7238 DVDD.n916 VSS 0.033945f
C7239 DVDD.n917 VSS 0.033945f
C7240 DVDD.n918 VSS 0.028497f
C7241 DVDD.n919 VSS 0.053165f
C7242 DVDD.n920 VSS 0.05956f
C7243 DVDD.n921 VSS 0.05956f
C7244 DVDD.n963 VSS 0.019729f
C7245 DVDD.n965 VSS 0.019729f
C7246 DVDD.n966 VSS 0.031128f
C7247 DVDD.n967 VSS 0.031128f
C7248 DVDD.n968 VSS 0.031128f
C7249 DVDD.n969 VSS 0.031128f
C7250 DVDD.n970 VSS 0.031128f
C7251 DVDD.n972 VSS 0.031128f
C7252 DVDD.n973 VSS 0.031128f
C7253 DVDD.n974 VSS 0.031128f
C7254 DVDD.n975 VSS 0.031128f
C7255 DVDD.n977 VSS 0.031128f
C7256 DVDD.n978 VSS 0.031128f
C7257 DVDD.n979 VSS 0.031128f
C7258 DVDD.n980 VSS 0.031128f
C7259 DVDD.n982 VSS 0.031128f
C7260 DVDD.n983 VSS 0.031128f
C7261 DVDD.n984 VSS 0.031128f
C7262 DVDD.n985 VSS 0.031128f
C7263 DVDD.n987 VSS 0.031128f
C7264 DVDD.n988 VSS 0.031128f
C7265 DVDD.n989 VSS 0.031128f
C7266 DVDD.n990 VSS 0.031128f
C7267 DVDD.n992 VSS 0.031128f
C7268 DVDD.n993 VSS 0.031128f
C7269 DVDD.n994 VSS 0.031128f
C7270 DVDD.n995 VSS 0.031128f
C7271 DVDD.n997 VSS 0.031128f
C7272 DVDD.n998 VSS 0.031128f
C7273 DVDD.n999 VSS 0.031128f
C7274 DVDD.n1000 VSS 0.031128f
C7275 DVDD.n1002 VSS 0.031128f
C7276 DVDD.n1003 VSS 0.031128f
C7277 DVDD.n1004 VSS 0.031128f
C7278 DVDD.n1005 VSS 0.031128f
C7279 DVDD.n1007 VSS 0.031128f
C7280 DVDD.n1008 VSS 0.031128f
C7281 DVDD.n1009 VSS 0.031128f
C7282 DVDD.n1010 VSS 0.031128f
C7283 DVDD.n1012 VSS 0.031128f
C7284 DVDD.n1013 VSS 0.031128f
C7285 DVDD.n1014 VSS 0.031128f
C7286 DVDD.n1015 VSS 0.031128f
C7287 DVDD.n1017 VSS 0.031128f
C7288 DVDD.n1018 VSS 0.031128f
C7289 DVDD.n1019 VSS 0.031128f
C7290 DVDD.n1020 VSS 0.031128f
C7291 DVDD.n1022 VSS 0.031128f
C7292 DVDD.n1023 VSS 0.031128f
C7293 DVDD.n1024 VSS 0.031128f
C7294 DVDD.n1025 VSS 0.031128f
C7295 DVDD.n1027 VSS 0.031128f
C7296 DVDD.n1028 VSS 0.031128f
C7297 DVDD.n1029 VSS 0.031128f
C7298 DVDD.n1030 VSS 0.031128f
C7299 DVDD.n1032 VSS 0.031128f
C7300 DVDD.n1033 VSS 0.031128f
C7301 DVDD.n1034 VSS 0.031128f
C7302 DVDD.n1035 VSS 0.031128f
C7303 DVDD.n1037 VSS 0.031128f
C7304 DVDD.n1038 VSS 0.031128f
C7305 DVDD.n1039 VSS 0.031128f
C7306 DVDD.n1040 VSS 0.031128f
C7307 DVDD.n1042 VSS 0.031128f
C7308 DVDD.n1043 VSS 0.031128f
C7309 DVDD.n1044 VSS 0.031128f
C7310 DVDD.n1045 VSS 0.031128f
C7311 DVDD.n1047 VSS 0.031128f
C7312 DVDD.n1048 VSS 0.031128f
C7313 DVDD.n1049 VSS 0.031128f
C7314 DVDD.n1050 VSS 0.031128f
C7315 DVDD.n1052 VSS 0.031128f
C7316 DVDD.n1053 VSS 0.031128f
C7317 DVDD.n1054 VSS 0.031128f
C7318 DVDD.n1055 VSS 0.031128f
C7319 DVDD.n1057 VSS 0.031128f
C7320 DVDD.n1058 VSS 0.031128f
C7321 DVDD.n1059 VSS 0.031128f
C7322 DVDD.n1060 VSS 0.031128f
C7323 DVDD.n1062 VSS 0.031128f
C7324 DVDD.n1063 VSS 0.031128f
C7325 DVDD.n1064 VSS 0.031128f
C7326 DVDD.n1065 VSS 0.031128f
C7327 DVDD.n1067 VSS 0.031128f
C7328 DVDD.n1068 VSS 0.019729f
C7329 DVDD.n1069 VSS 0.019729f
C7330 DVDD.n1070 VSS 0.026086f
C7331 DVDD.n1071 VSS 0.031128f
C7332 DVDD.n1072 VSS 0.031128f
C7333 DVDD.n1073 VSS 0.031128f
C7334 DVDD.n1074 VSS 0.031128f
C7335 DVDD.n1075 VSS 0.031128f
C7336 DVDD.n1077 VSS 0.031128f
C7337 DVDD.n1078 VSS 0.031128f
C7338 DVDD.n1079 VSS 0.031128f
C7339 DVDD.n1080 VSS 0.031128f
C7340 DVDD.n1081 VSS 0.031128f
C7341 DVDD.n1082 VSS 0.031128f
C7342 DVDD.n1083 VSS 0.031128f
C7343 DVDD.n1084 VSS 0.031128f
C7344 DVDD.n1086 VSS 0.031128f
C7345 DVDD.n1087 VSS 0.031128f
C7346 DVDD.n1088 VSS 0.031128f
C7347 DVDD.n1089 VSS 0.031128f
C7348 DVDD.n1090 VSS 0.031128f
C7349 DVDD.n1091 VSS 0.031128f
C7350 DVDD.n1092 VSS 0.031128f
C7351 DVDD.n1093 VSS 0.031128f
C7352 DVDD.n1095 VSS 0.031128f
C7353 DVDD.n1096 VSS 0.031128f
C7354 DVDD.n1097 VSS 0.031128f
C7355 DVDD.n1098 VSS 0.031128f
C7356 DVDD.n1099 VSS 0.031128f
C7357 DVDD.n1100 VSS 0.031128f
C7358 DVDD.n1101 VSS 0.031128f
C7359 DVDD.n1102 VSS 0.031128f
C7360 DVDD.n1104 VSS 0.031128f
C7361 DVDD.n1105 VSS 0.031128f
C7362 DVDD.n1106 VSS 0.031128f
C7363 DVDD.n1107 VSS 0.031128f
C7364 DVDD.n1108 VSS 0.031128f
C7365 DVDD.n1109 VSS 0.031128f
C7366 DVDD.n1110 VSS 0.031128f
C7367 DVDD.n1111 VSS 0.031128f
C7368 DVDD.n1113 VSS 0.031128f
C7369 DVDD.n1114 VSS 0.031128f
C7370 DVDD.n1115 VSS 0.031128f
C7371 DVDD.n1116 VSS 0.031128f
C7372 DVDD.n1117 VSS 0.031128f
C7373 DVDD.n1118 VSS 0.031128f
C7374 DVDD.n1119 VSS 0.031128f
C7375 DVDD.n1120 VSS 0.031128f
C7376 DVDD.n1122 VSS 0.031128f
C7377 DVDD.n1123 VSS 0.031128f
C7378 DVDD.n1124 VSS 0.031128f
C7379 DVDD.n1125 VSS 0.031128f
C7380 DVDD.n1126 VSS 0.031128f
C7381 DVDD.n1127 VSS 0.031128f
C7382 DVDD.n1128 VSS 0.031128f
C7383 DVDD.n1129 VSS 0.031128f
C7384 DVDD.n1131 VSS 0.031128f
C7385 DVDD.n1132 VSS 0.031128f
C7386 DVDD.n1133 VSS 0.031128f
C7387 DVDD.n1134 VSS 0.031128f
C7388 DVDD.n1135 VSS 0.031128f
C7389 DVDD.n1136 VSS 0.031128f
C7390 DVDD.n1137 VSS 0.031128f
C7391 DVDD.n1138 VSS 0.031128f
C7392 DVDD.n1140 VSS 0.031128f
C7393 DVDD.n1141 VSS 0.031128f
C7394 DVDD.n1142 VSS 0.031128f
C7395 DVDD.n1143 VSS 0.031128f
C7396 DVDD.n1144 VSS 0.031128f
C7397 DVDD.n1145 VSS 0.031128f
C7398 DVDD.n1146 VSS 0.031128f
C7399 DVDD.n1147 VSS 0.031128f
C7400 DVDD.n1149 VSS 0.031128f
C7401 DVDD.n1150 VSS 0.031128f
C7402 DVDD.n1151 VSS 0.031128f
C7403 DVDD.n1152 VSS 0.031128f
C7404 DVDD.n1153 VSS 0.031128f
C7405 DVDD.n1154 VSS 0.031128f
C7406 DVDD.n1155 VSS 0.031128f
C7407 DVDD.n1156 VSS 0.031128f
C7408 DVDD.n1158 VSS 0.031128f
C7409 DVDD.n1159 VSS 0.031128f
C7410 DVDD.n1160 VSS 0.031128f
C7411 DVDD.n1161 VSS 0.031128f
C7412 DVDD.n1162 VSS 0.031128f
C7413 DVDD.n1163 VSS 0.031128f
C7414 DVDD.n1164 VSS 0.031128f
C7415 DVDD.n1165 VSS 0.031128f
C7416 DVDD.n1167 VSS 0.031128f
C7417 DVDD.n1168 VSS 0.031128f
C7418 DVDD.n1169 VSS 0.031128f
C7419 DVDD.n1170 VSS 0.031128f
C7420 DVDD.n1171 VSS 0.031128f
C7421 DVDD.n1172 VSS 0.031128f
C7422 DVDD.n1173 VSS 0.031128f
C7423 DVDD.n1174 VSS 0.031128f
C7424 DVDD.n1176 VSS 0.031128f
C7425 DVDD.n1177 VSS 0.031128f
C7426 DVDD.n1178 VSS 0.031128f
C7427 DVDD.n1179 VSS 0.031128f
C7428 DVDD.n1180 VSS 0.031128f
C7429 DVDD.n1181 VSS 0.031128f
C7430 DVDD.n1182 VSS 0.031128f
C7431 DVDD.n1183 VSS 0.031128f
C7432 DVDD.n1185 VSS 0.031128f
C7433 DVDD.n1186 VSS 0.031128f
C7434 DVDD.n1187 VSS 0.031128f
C7435 DVDD.n1188 VSS 0.031128f
C7436 DVDD.n1189 VSS 0.031128f
C7437 DVDD.n1190 VSS 0.031128f
C7438 DVDD.n1191 VSS 0.031128f
C7439 DVDD.n1192 VSS 0.031128f
C7440 DVDD.n1194 VSS 0.031128f
C7441 DVDD.n1195 VSS 0.031128f
C7442 DVDD.n1196 VSS 0.031128f
C7443 DVDD.n1197 VSS 0.031128f
C7444 DVDD.n1198 VSS 0.031128f
C7445 DVDD.n1199 VSS 0.031128f
C7446 DVDD.n1200 VSS 0.031128f
C7447 DVDD.n1201 VSS 0.031128f
C7448 DVDD.n1203 VSS 0.031128f
C7449 DVDD.n1204 VSS 0.031128f
C7450 DVDD.n1205 VSS 0.031128f
C7451 DVDD.n1206 VSS 0.031128f
C7452 DVDD.n1207 VSS 0.031128f
C7453 DVDD.n1208 VSS 0.031128f
C7454 DVDD.n1209 VSS 0.031128f
C7455 DVDD.n1210 VSS 0.031128f
C7456 DVDD.n1212 VSS 0.031128f
C7457 DVDD.n1213 VSS 0.031128f
C7458 DVDD.n1214 VSS 0.031128f
C7459 DVDD.n1215 VSS 0.031128f
C7460 DVDD.n1216 VSS 0.031128f
C7461 DVDD.n1217 VSS 0.031128f
C7462 DVDD.n1218 VSS 0.031128f
C7463 DVDD.n1219 VSS 0.031128f
C7464 DVDD.n1221 VSS 0.031128f
C7465 DVDD.n1222 VSS 0.031128f
C7466 DVDD.n1223 VSS 0.031128f
C7467 DVDD.n1224 VSS 0.031128f
C7468 DVDD.n1225 VSS 0.031128f
C7469 DVDD.n1226 VSS 0.031128f
C7470 DVDD.n1227 VSS 0.031128f
C7471 DVDD.n1228 VSS 0.031128f
C7472 DVDD.n1230 VSS 0.031128f
C7473 DVDD.n1231 VSS 0.031128f
C7474 DVDD.n1232 VSS 0.031128f
C7475 DVDD.n1233 VSS 0.031128f
C7476 DVDD.n1234 VSS 0.031128f
C7477 DVDD.n1235 VSS 0.031128f
C7478 DVDD.n1236 VSS 0.031128f
C7479 DVDD.n1237 VSS 0.031128f
C7480 DVDD.n1239 VSS 0.031128f
C7481 DVDD.n1240 VSS 0.031128f
C7482 DVDD.n1241 VSS 0.031128f
C7483 DVDD.n1242 VSS 0.031128f
C7484 DVDD.n1243 VSS 0.031128f
C7485 DVDD.n1244 VSS 0.031128f
C7486 DVDD.n1245 VSS 0.031128f
C7487 DVDD.n1246 VSS 0.031128f
C7488 DVDD.n1248 VSS 0.031128f
C7489 DVDD.n1249 VSS 0.031128f
C7490 DVDD.n1250 VSS 0.031128f
C7491 DVDD.n1251 VSS 0.031128f
C7492 DVDD.n1252 VSS 0.031128f
C7493 DVDD.n1253 VSS 0.031128f
C7494 DVDD.n1254 VSS 0.031128f
C7495 DVDD.n1256 VSS 0.509617f
C7496 DVDD.n1257 VSS 0.041931f
C7497 DVDD.n1258 VSS 0.041931f
C7498 DVDD.n1259 VSS 0.028833f
C7499 DVDD.n1260 VSS 0.02513f
C7500 DVDD.n1261 VSS 0.02513f
C7501 DVDD.n1262 VSS 0.459077f
C7502 DVDD.n1263 VSS 0.433807f
C7503 DVDD.n1264 VSS 0.534888f
C7504 DVDD.n1265 VSS 0.033945f
C7505 DVDD.n1266 VSS 0.033945f
C7506 DVDD.n1267 VSS 0.028497f
C7507 DVDD.n1268 VSS 0.053165f
C7508 DVDD.n1269 VSS 0.05956f
C7509 DVDD.n1270 VSS 0.05956f
C7510 DVDD.n1312 VSS 0.031128f
C7511 DVDD.n1314 VSS 0.031128f
C7512 DVDD.n1315 VSS 0.031128f
C7513 DVDD.n1316 VSS 0.031128f
C7514 DVDD.n1317 VSS 0.031128f
C7515 DVDD.n1318 VSS 0.031128f
C7516 DVDD.n1319 VSS 0.031128f
C7517 DVDD.n1320 VSS 0.031128f
C7518 DVDD.n1321 VSS 0.031128f
C7519 DVDD.n1322 VSS 0.031128f
C7520 DVDD.n1323 VSS 0.031128f
C7521 DVDD.n1324 VSS 0.031128f
C7522 DVDD.n1325 VSS 0.031128f
C7523 DVDD.n1326 VSS 0.031128f
C7524 DVDD.n1327 VSS 0.031128f
C7525 DVDD.n1328 VSS 0.031128f
C7526 DVDD.n1329 VSS 0.031128f
C7527 DVDD.n1330 VSS 0.031128f
C7528 DVDD.n1331 VSS 0.031128f
C7529 DVDD.n1332 VSS 0.031128f
C7530 DVDD.n1333 VSS 0.031128f
C7531 DVDD.n1334 VSS 0.031128f
C7532 DVDD.n1335 VSS 0.031128f
C7533 DVDD.n1336 VSS 0.031128f
C7534 DVDD.n1337 VSS 0.031128f
C7535 DVDD.n1338 VSS 0.031128f
C7536 DVDD.n1339 VSS 0.031128f
C7537 DVDD.n1340 VSS 0.031128f
C7538 DVDD.n1341 VSS 0.031128f
C7539 DVDD.n1342 VSS 0.031128f
C7540 DVDD.n1343 VSS 0.031128f
C7541 DVDD.n1344 VSS 0.031128f
C7542 DVDD.n1345 VSS 0.031128f
C7543 DVDD.n1346 VSS 0.031128f
C7544 DVDD.n1347 VSS 0.031128f
C7545 DVDD.n1348 VSS 0.031128f
C7546 DVDD.n1349 VSS 0.031128f
C7547 DVDD.n1350 VSS 0.031128f
C7548 DVDD.n1351 VSS 0.031128f
C7549 DVDD.n1352 VSS 0.031128f
C7550 DVDD.n1353 VSS 0.031128f
C7551 DVDD.n1354 VSS 0.031128f
C7552 DVDD.n1355 VSS 0.031128f
C7553 DVDD.n1356 VSS 0.019729f
C7554 DVDD.n1357 VSS 0.019729f
C7555 DVDD.n1358 VSS 0.026086f
C7556 DVDD.n1359 VSS 0.031128f
C7557 DVDD.n1360 VSS 0.031128f
C7558 DVDD.n1361 VSS 0.031128f
C7559 DVDD.n1363 VSS 0.031128f
C7560 DVDD.n1364 VSS 0.031128f
C7561 DVDD.n1365 VSS 0.031128f
C7562 DVDD.n1366 VSS 0.031128f
C7563 DVDD.n1368 VSS 0.031128f
C7564 DVDD.n1369 VSS 0.031128f
C7565 DVDD.n1370 VSS 0.031128f
C7566 DVDD.n1371 VSS 0.031128f
C7567 DVDD.n1372 VSS 0.031128f
C7568 DVDD.n1373 VSS 0.031128f
C7569 DVDD.n1375 VSS 0.031128f
C7570 DVDD.n1376 VSS 0.031128f
C7571 DVDD.n1377 VSS 0.031128f
C7572 DVDD.n1378 VSS 0.031128f
C7573 DVDD.n1380 VSS 0.031128f
C7574 DVDD.n1381 VSS 0.031128f
C7575 DVDD.n1382 VSS 0.031128f
C7576 DVDD.n1383 VSS 0.031128f
C7577 DVDD.n1384 VSS 0.031128f
C7578 DVDD.n1385 VSS 0.031128f
C7579 DVDD.n1387 VSS 0.031128f
C7580 DVDD.n1388 VSS 0.031128f
C7581 DVDD.n1389 VSS 0.031128f
C7582 DVDD.n1390 VSS 0.031128f
C7583 DVDD.n1392 VSS 0.031128f
C7584 DVDD.n1393 VSS 0.031128f
C7585 DVDD.n1394 VSS 0.031128f
C7586 DVDD.n1395 VSS 0.031128f
C7587 DVDD.n1396 VSS 0.031128f
C7588 DVDD.n1397 VSS 0.031128f
C7589 DVDD.n1399 VSS 0.031128f
C7590 DVDD.n1400 VSS 0.031128f
C7591 DVDD.n1401 VSS 0.031128f
C7592 DVDD.n1402 VSS 0.031128f
C7593 DVDD.n1404 VSS 0.031128f
C7594 DVDD.n1405 VSS 0.031128f
C7595 DVDD.n1406 VSS 0.031128f
C7596 DVDD.n1407 VSS 0.031128f
C7597 DVDD.n1408 VSS 0.031128f
C7598 DVDD.n1409 VSS 0.031128f
C7599 DVDD.n1411 VSS 0.031128f
C7600 DVDD.n1412 VSS 0.031128f
C7601 DVDD.n1413 VSS 0.031128f
C7602 DVDD.n1414 VSS 0.031128f
C7603 DVDD.n1416 VSS 0.031128f
C7604 DVDD.n1417 VSS 0.031128f
C7605 DVDD.n1418 VSS 0.031128f
C7606 DVDD.n1419 VSS 0.031128f
C7607 DVDD.n1420 VSS 0.031128f
C7608 DVDD.n1421 VSS 0.031128f
C7609 DVDD.n1423 VSS 0.031128f
C7610 DVDD.n1424 VSS 0.031128f
C7611 DVDD.n1425 VSS 0.031128f
C7612 DVDD.n1426 VSS 0.031128f
C7613 DVDD.n1428 VSS 0.031128f
C7614 DVDD.n1429 VSS 0.031128f
C7615 DVDD.n1430 VSS 0.031128f
C7616 DVDD.n1431 VSS 0.031128f
C7617 DVDD.n1432 VSS 0.031128f
C7618 DVDD.n1433 VSS 0.031128f
C7619 DVDD.n1435 VSS 0.031128f
C7620 DVDD.n1436 VSS 0.031128f
C7621 DVDD.n1437 VSS 0.031128f
C7622 DVDD.n1438 VSS 0.031128f
C7623 DVDD.n1440 VSS 0.031128f
C7624 DVDD.n1441 VSS 0.031128f
C7625 DVDD.n1442 VSS 0.031128f
C7626 DVDD.n1443 VSS 0.031128f
C7627 DVDD.n1444 VSS 0.031128f
C7628 DVDD.n1445 VSS 0.031128f
C7629 DVDD.n1447 VSS 0.031128f
C7630 DVDD.n1448 VSS 0.031128f
C7631 DVDD.n1449 VSS 0.031128f
C7632 DVDD.n1450 VSS 0.031128f
C7633 DVDD.n1452 VSS 0.031128f
C7634 DVDD.n1453 VSS 0.031128f
C7635 DVDD.n1454 VSS 0.031128f
C7636 DVDD.n1455 VSS 0.031128f
C7637 DVDD.n1456 VSS 0.031128f
C7638 DVDD.n1457 VSS 0.031128f
C7639 DVDD.n1459 VSS 0.031128f
C7640 DVDD.n1460 VSS 0.031128f
C7641 DVDD.n1461 VSS 0.031128f
C7642 DVDD.n1462 VSS 0.031128f
C7643 DVDD.n1464 VSS 0.031128f
C7644 DVDD.n1465 VSS 0.031128f
C7645 DVDD.n1466 VSS 0.031128f
C7646 DVDD.n1467 VSS 0.031128f
C7647 DVDD.n1468 VSS 0.031128f
C7648 DVDD.n1469 VSS 0.031128f
C7649 DVDD.n1471 VSS 0.031128f
C7650 DVDD.n1472 VSS 0.031128f
C7651 DVDD.n1473 VSS 0.031128f
C7652 DVDD.n1474 VSS 0.031128f
C7653 DVDD.n1476 VSS 0.031128f
C7654 DVDD.n1477 VSS 0.031128f
C7655 DVDD.n1478 VSS 0.031128f
C7656 DVDD.n1479 VSS 0.031128f
C7657 DVDD.n1480 VSS 0.031128f
C7658 DVDD.n1481 VSS 0.031128f
C7659 DVDD.n1483 VSS 0.031128f
C7660 DVDD.n1484 VSS 0.031128f
C7661 DVDD.n1485 VSS 0.031128f
C7662 DVDD.n1486 VSS 0.031128f
C7663 DVDD.n1488 VSS 0.031128f
C7664 DVDD.n1489 VSS 0.031128f
C7665 DVDD.n1490 VSS 0.031128f
C7666 DVDD.n1491 VSS 0.031128f
C7667 DVDD.n1492 VSS 0.031128f
C7668 DVDD.n1493 VSS 0.031128f
C7669 DVDD.n1495 VSS 0.031128f
C7670 DVDD.n1496 VSS 0.031128f
C7671 DVDD.n1497 VSS 0.031128f
C7672 DVDD.n1498 VSS 0.031128f
C7673 DVDD.n1500 VSS 0.031128f
C7674 DVDD.n1501 VSS 0.031128f
C7675 DVDD.n1502 VSS 0.031128f
C7676 DVDD.n1503 VSS 0.031128f
C7677 DVDD.n1504 VSS 0.031128f
C7678 DVDD.n1505 VSS 0.031128f
C7679 DVDD.n1507 VSS 0.031128f
C7680 DVDD.n1508 VSS 0.031128f
C7681 DVDD.n1509 VSS 0.031128f
C7682 DVDD.n1510 VSS 0.031128f
C7683 DVDD.n1512 VSS 0.031128f
C7684 DVDD.n1513 VSS 0.031128f
C7685 DVDD.n1514 VSS 0.031128f
C7686 DVDD.n1515 VSS 0.031128f
C7687 DVDD.n1516 VSS 0.031128f
C7688 DVDD.n1517 VSS 0.031128f
C7689 DVDD.n1519 VSS 0.031128f
C7690 DVDD.n1520 VSS 0.031128f
C7691 DVDD.n1521 VSS 0.031128f
C7692 DVDD.n1522 VSS 0.031128f
C7693 DVDD.n1524 VSS 0.031128f
C7694 DVDD.n1525 VSS 0.031128f
C7695 DVDD.n1526 VSS 0.031128f
C7696 DVDD.n1527 VSS 0.031128f
C7697 DVDD.n1528 VSS 0.031128f
C7698 DVDD.n1529 VSS 0.031128f
C7699 DVDD.n1531 VSS 0.031128f
C7700 DVDD.n1532 VSS 0.031128f
C7701 DVDD.n1533 VSS 0.031128f
C7702 DVDD.n1534 VSS 0.031128f
C7703 DVDD.n1536 VSS 0.031128f
C7704 DVDD.n1537 VSS 0.031128f
C7705 DVDD.n1538 VSS 0.031128f
C7706 DVDD.n1539 VSS 0.031128f
C7707 DVDD.n1540 VSS 0.031128f
C7708 DVDD.n1541 VSS 0.031128f
C7709 DVDD.n1543 VSS 0.031128f
C7710 DVDD.n1544 VSS 0.031128f
C7711 DVDD.n1545 VSS 0.031128f
C7712 DVDD.n1546 VSS 0.031128f
C7713 DVDD.n1548 VSS 0.031128f
C7714 DVDD.n1549 VSS 0.031128f
C7715 DVDD.n1550 VSS 0.031128f
C7716 DVDD.n1551 VSS 0.031128f
C7717 DVDD.n1552 VSS 0.031128f
C7718 DVDD.n1553 VSS 0.031128f
C7719 DVDD.n1555 VSS 0.031128f
C7720 DVDD.n1556 VSS 0.031128f
C7721 DVDD.n1557 VSS 0.031128f
C7722 DVDD.n1558 VSS 0.031128f
C7723 DVDD.n1560 VSS 0.031128f
C7724 DVDD.n1561 VSS 0.031128f
C7725 DVDD.n1562 VSS 0.031128f
C7726 DVDD.n1563 VSS 0.031128f
C7727 DVDD.n1564 VSS 0.031128f
C7728 DVDD.n1565 VSS 0.031128f
C7729 DVDD.n1567 VSS 0.031128f
C7730 DVDD.n1568 VSS 0.031128f
C7731 DVDD.n1569 VSS 0.031128f
C7732 DVDD.n1570 VSS 0.031128f
C7733 DVDD.n1572 VSS 0.031128f
C7734 DVDD.n1573 VSS 0.031128f
C7735 DVDD.n1574 VSS 0.031128f
C7736 DVDD.n1575 VSS 0.031128f
C7737 DVDD.n1576 VSS 0.031128f
C7738 DVDD.n1577 VSS 0.031128f
C7739 DVDD.n1579 VSS 0.031128f
C7740 DVDD.n1580 VSS 0.031128f
C7741 DVDD.n1581 VSS 0.031128f
C7742 DVDD.n1582 VSS 0.031128f
C7743 DVDD.n1584 VSS 0.031128f
C7744 DVDD.n1585 VSS 0.031128f
C7745 DVDD.n1586 VSS 0.031128f
C7746 DVDD.n1587 VSS 0.031128f
C7747 DVDD.n1588 VSS 0.031128f
C7748 DVDD.n1589 VSS 0.031128f
C7749 DVDD.n1591 VSS 0.031128f
C7750 DVDD.n1592 VSS 0.031128f
C7751 DVDD.n1593 VSS 0.031128f
C7752 DVDD.n1594 VSS 0.031128f
C7753 DVDD.n1596 VSS 0.031128f
C7754 DVDD.n1597 VSS 0.031128f
C7755 DVDD.n1598 VSS 0.031128f
C7756 DVDD.n1599 VSS 0.031128f
C7757 DVDD.n1600 VSS 0.031128f
C7758 DVDD.n1601 VSS 0.031128f
C7759 DVDD.n1602 VSS 0.019729f
C7760 DVDD.n1603 VSS 0.019729f
C7761 DVDD.n1605 VSS 0.383266f
C7762 DVDD.n1606 VSS 0.041931f
C7763 DVDD.n1607 VSS 0.041931f
C7764 DVDD.n1608 VSS 0.028833f
C7765 DVDD.n1609 VSS 0.02513f
C7766 DVDD.n1610 VSS 0.02513f
C7767 DVDD.n1611 VSS 0.560158f
C7768 DVDD.n1653 VSS 0.019729f
C7769 DVDD.n1654 VSS 0.526464f
C7770 DVDD.n1655 VSS 0.522252f
C7771 DVDD.n1656 VSS 0.560158f
C7772 DVDD.n1657 VSS 0.019729f
C7773 DVDD.n1658 VSS 0.366419f
C7774 DVDD.n1659 VSS 0.031128f
C7775 DVDD.n1660 VSS 0.031128f
C7776 DVDD.n1661 VSS 0.031128f
C7777 DVDD.n1662 VSS 0.031128f
C7778 DVDD.n1663 VSS 0.031128f
C7779 DVDD.n1664 VSS 0.031128f
C7780 DVDD.n1665 VSS 0.031128f
C7781 DVDD.n1666 VSS 0.031128f
C7782 DVDD.n1667 VSS 0.031128f
C7783 DVDD.n1668 VSS 0.031128f
C7784 DVDD.n1669 VSS 0.031128f
C7785 DVDD.n1670 VSS 0.031128f
C7786 DVDD.n1671 VSS 0.031128f
C7787 DVDD.n1672 VSS 0.031128f
C7788 DVDD.n1673 VSS 0.031128f
C7789 DVDD.n1674 VSS 0.031128f
C7790 DVDD.n1675 VSS 0.031128f
C7791 DVDD.n1676 VSS 0.031128f
C7792 DVDD.n1677 VSS 0.031128f
C7793 DVDD.n1678 VSS 0.031128f
C7794 DVDD.n1679 VSS 0.031128f
C7795 DVDD.n1680 VSS 0.031128f
C7796 DVDD.n1681 VSS 0.031128f
C7797 DVDD.n1682 VSS 0.031128f
C7798 DVDD.n1683 VSS 0.031128f
C7799 DVDD.n1684 VSS 0.031128f
C7800 DVDD.n1685 VSS 0.031128f
C7801 DVDD.n1686 VSS 0.031128f
C7802 DVDD.n1687 VSS 0.031128f
C7803 DVDD.n1688 VSS 0.031128f
C7804 DVDD.n1689 VSS 0.031128f
C7805 DVDD.n1690 VSS 0.031128f
C7806 DVDD.n1691 VSS 0.031128f
C7807 DVDD.n1692 VSS 0.031128f
C7808 DVDD.n1693 VSS 0.031128f
C7809 DVDD.n1694 VSS 0.031128f
C7810 DVDD.n1695 VSS 0.031128f
C7811 DVDD.n1696 VSS 0.031128f
C7812 DVDD.n1697 VSS 0.031128f
C7813 DVDD.n1698 VSS 0.031128f
C7814 DVDD.n1700 VSS 0.031128f
C7815 DVDD.n1701 VSS 0.031128f
C7816 DVDD.n1702 VSS 0.039516f
C7817 DVDD.n1703 VSS 0.0586f
C7818 DVDD.n1704 VSS 0.05956f
C7819 DVDD.n1705 VSS 0.05956f
C7820 DVDD.n1706 VSS 0.522252f
C7821 DVDD.n1707 VSS 0.041931f
C7822 DVDD.n1708 VSS 0.041931f
C7823 DVDD.n1709 VSS 0.028833f
C7824 DVDD.n1710 VSS 0.02513f
C7825 DVDD.n1711 VSS 0.02513f
C7826 DVDD.n1712 VSS 0.438018f
C7827 DVDD.n1754 VSS 0.019729f
C7828 DVDD.n1755 VSS 0.438018f
C7829 DVDD.n1756 VSS 0.019729f
C7830 DVDD.n1757 VSS 0.522252f
C7831 DVDD.n1758 VSS 0.031128f
C7832 DVDD.n1759 VSS 0.031128f
C7833 DVDD.n1760 VSS 0.031128f
C7834 DVDD.n1761 VSS 0.031128f
C7835 DVDD.n1762 VSS 0.031128f
C7836 DVDD.n1763 VSS 0.031128f
C7837 DVDD.n1764 VSS 0.031128f
C7838 DVDD.n1765 VSS 0.031128f
C7839 DVDD.n1766 VSS 0.031128f
C7840 DVDD.n1767 VSS 0.031128f
C7841 DVDD.n1768 VSS 0.031128f
C7842 DVDD.n1769 VSS 0.031128f
C7843 DVDD.n1770 VSS 0.031128f
C7844 DVDD.n1771 VSS 0.031128f
C7845 DVDD.n1772 VSS 0.031128f
C7846 DVDD.n1773 VSS 0.031128f
C7847 DVDD.n1774 VSS 0.031128f
C7848 DVDD.n1775 VSS 0.031128f
C7849 DVDD.n1776 VSS 0.031128f
C7850 DVDD.n1777 VSS 0.031128f
C7851 DVDD.n1778 VSS 0.031128f
C7852 DVDD.n1779 VSS 0.031128f
C7853 DVDD.n1780 VSS 0.031128f
C7854 DVDD.n1781 VSS 0.031128f
C7855 DVDD.n1782 VSS 0.031128f
C7856 DVDD.n1783 VSS 0.031128f
C7857 DVDD.n1784 VSS 0.031128f
C7858 DVDD.n1785 VSS 0.031128f
C7859 DVDD.n1786 VSS 0.031128f
C7860 DVDD.n1787 VSS 0.031128f
C7861 DVDD.n1788 VSS 0.031128f
C7862 DVDD.n1789 VSS 0.031128f
C7863 DVDD.n1790 VSS 0.031128f
C7864 DVDD.n1791 VSS 0.031128f
C7865 DVDD.n1792 VSS 0.031128f
C7866 DVDD.n1793 VSS 0.031128f
C7867 DVDD.n1794 VSS 0.031128f
C7868 DVDD.n1795 VSS 0.031128f
C7869 DVDD.n1796 VSS 0.031128f
C7870 DVDD.n1797 VSS 0.031128f
C7871 DVDD.n1799 VSS 0.031128f
C7872 DVDD.n1800 VSS 0.031128f
C7873 DVDD.n1801 VSS 0.039516f
C7874 DVDD.n1802 VSS 0.051875f
C7875 DVDD.n1803 VSS 0.05956f
C7876 DVDD.n1804 VSS 0.05956f
C7877 DVDD.n1805 VSS 0.598063f
C7878 DVDD.n1806 VSS 0.041931f
C7879 DVDD.n1807 VSS 0.041931f
C7880 DVDD.n1808 VSS 0.028833f
C7881 DVDD.n1809 VSS 0.02513f
C7882 DVDD.n1810 VSS 0.02513f
C7883 DVDD.n1811 VSS 0.315878f
C7884 DVDD.n1812 VSS 0.463288f
C7885 DVDD.n1813 VSS 0.374843f
C7886 DVDD.n1814 VSS 0.033945f
C7887 DVDD.n1815 VSS 0.033945f
C7888 DVDD.n1816 VSS 0.05956f
C7889 DVDD.n1817 VSS 0.028497f
C7890 DVDD.n1818 VSS 0.037515f
C7891 DVDD.n1819 VSS 0.05956f
C7892 DVDD.n1820 VSS 0.050915f
C7893 DVDD.n1821 VSS 0.522252f
C7894 DVDD.n1863 VSS 0.031128f
C7895 DVDD.n1865 VSS 0.031128f
C7896 DVDD.n1866 VSS 0.031128f
C7897 DVDD.n1867 VSS 0.031128f
C7898 DVDD.n1868 VSS 0.031128f
C7899 DVDD.n1869 VSS 0.031128f
C7900 DVDD.n1870 VSS 0.031128f
C7901 DVDD.n1871 VSS 0.031128f
C7902 DVDD.n1872 VSS 0.031128f
C7903 DVDD.n1873 VSS 0.031128f
C7904 DVDD.n1874 VSS 0.031128f
C7905 DVDD.n1875 VSS 0.031128f
C7906 DVDD.n1876 VSS 0.031128f
C7907 DVDD.n1877 VSS 0.031128f
C7908 DVDD.n1878 VSS 0.031128f
C7909 DVDD.n1879 VSS 0.031128f
C7910 DVDD.n1880 VSS 0.031128f
C7911 DVDD.n1881 VSS 0.031128f
C7912 DVDD.n1882 VSS 0.031128f
C7913 DVDD.n1883 VSS 0.031128f
C7914 DVDD.n1884 VSS 0.031128f
C7915 DVDD.n1885 VSS 0.031128f
C7916 DVDD.n1886 VSS 0.031128f
C7917 DVDD.n1887 VSS 0.031128f
C7918 DVDD.n1888 VSS 0.031128f
C7919 DVDD.n1889 VSS 0.031128f
C7920 DVDD.n1890 VSS 0.031128f
C7921 DVDD.n1891 VSS 0.031128f
C7922 DVDD.n1892 VSS 0.031128f
C7923 DVDD.n1893 VSS 0.031128f
C7924 DVDD.n1894 VSS 0.031128f
C7925 DVDD.n1895 VSS 0.031128f
C7926 DVDD.n1896 VSS 0.031128f
C7927 DVDD.n1897 VSS 0.031128f
C7928 DVDD.n1898 VSS 0.031128f
C7929 DVDD.n1899 VSS 0.031128f
C7930 DVDD.n1900 VSS 0.031128f
C7931 DVDD.n1901 VSS 0.031128f
C7932 DVDD.n1902 VSS 0.031128f
C7933 DVDD.n1903 VSS 0.031128f
C7934 DVDD.n1904 VSS 0.031128f
C7935 DVDD.n1905 VSS 0.031128f
C7936 DVDD.n1906 VSS 0.031128f
C7937 DVDD.n1907 VSS 0.019729f
C7938 DVDD.n1908 VSS 0.019729f
C7939 DVDD.n1909 VSS 0.026086f
C7940 DVDD.n1910 VSS 0.031128f
C7941 DVDD.n1911 VSS 0.031128f
C7942 DVDD.n1912 VSS 0.031128f
C7943 DVDD.n1914 VSS 0.031128f
C7944 DVDD.n1915 VSS 0.031128f
C7945 DVDD.n1916 VSS 0.031128f
C7946 DVDD.n1917 VSS 0.031128f
C7947 DVDD.n1919 VSS 0.031128f
C7948 DVDD.n1920 VSS 0.031128f
C7949 DVDD.n1921 VSS 0.031128f
C7950 DVDD.n1922 VSS 0.031128f
C7951 DVDD.n1923 VSS 0.031128f
C7952 DVDD.n1924 VSS 0.031128f
C7953 DVDD.n1926 VSS 0.031128f
C7954 DVDD.n1927 VSS 0.031128f
C7955 DVDD.n1928 VSS 0.031128f
C7956 DVDD.n1929 VSS 0.031128f
C7957 DVDD.n1931 VSS 0.031128f
C7958 DVDD.n1932 VSS 0.031128f
C7959 DVDD.n1933 VSS 0.031128f
C7960 DVDD.n1934 VSS 0.031128f
C7961 DVDD.n1935 VSS 0.031128f
C7962 DVDD.n1936 VSS 0.031128f
C7963 DVDD.n1938 VSS 0.031128f
C7964 DVDD.n1939 VSS 0.031128f
C7965 DVDD.n1940 VSS 0.031128f
C7966 DVDD.n1941 VSS 0.031128f
C7967 DVDD.n1943 VSS 0.031128f
C7968 DVDD.n1944 VSS 0.031128f
C7969 DVDD.n1945 VSS 0.031128f
C7970 DVDD.n1946 VSS 0.031128f
C7971 DVDD.n1947 VSS 0.031128f
C7972 DVDD.n1948 VSS 0.031128f
C7973 DVDD.n1950 VSS 0.031128f
C7974 DVDD.n1951 VSS 0.031128f
C7975 DVDD.n1952 VSS 0.031128f
C7976 DVDD.n1953 VSS 0.031128f
C7977 DVDD.n1955 VSS 0.031128f
C7978 DVDD.n1956 VSS 0.031128f
C7979 DVDD.n1957 VSS 0.031128f
C7980 DVDD.n1958 VSS 0.031128f
C7981 DVDD.n1959 VSS 0.031128f
C7982 DVDD.n1960 VSS 0.031128f
C7983 DVDD.n1962 VSS 0.031128f
C7984 DVDD.n1963 VSS 0.031128f
C7985 DVDD.n1964 VSS 0.031128f
C7986 DVDD.n1965 VSS 0.031128f
C7987 DVDD.n1967 VSS 0.031128f
C7988 DVDD.n1968 VSS 0.031128f
C7989 DVDD.n1969 VSS 0.031128f
C7990 DVDD.n1970 VSS 0.031128f
C7991 DVDD.n1971 VSS 0.031128f
C7992 DVDD.n1972 VSS 0.031128f
C7993 DVDD.n1974 VSS 0.031128f
C7994 DVDD.n1975 VSS 0.031128f
C7995 DVDD.n1976 VSS 0.031128f
C7996 DVDD.n1977 VSS 0.031128f
C7997 DVDD.n1979 VSS 0.031128f
C7998 DVDD.n1980 VSS 0.031128f
C7999 DVDD.n1981 VSS 0.031128f
C8000 DVDD.n1982 VSS 0.031128f
C8001 DVDD.n1983 VSS 0.031128f
C8002 DVDD.n1984 VSS 0.031128f
C8003 DVDD.n1986 VSS 0.031128f
C8004 DVDD.n1987 VSS 0.031128f
C8005 DVDD.n1988 VSS 0.031128f
C8006 DVDD.n1989 VSS 0.031128f
C8007 DVDD.n1991 VSS 0.031128f
C8008 DVDD.n1992 VSS 0.031128f
C8009 DVDD.n1993 VSS 0.031128f
C8010 DVDD.n1994 VSS 0.031128f
C8011 DVDD.n1995 VSS 0.031128f
C8012 DVDD.n1996 VSS 0.031128f
C8013 DVDD.n1998 VSS 0.031128f
C8014 DVDD.n1999 VSS 0.031128f
C8015 DVDD.n2000 VSS 0.031128f
C8016 DVDD.n2001 VSS 0.031128f
C8017 DVDD.n2003 VSS 0.031128f
C8018 DVDD.n2004 VSS 0.031128f
C8019 DVDD.n2005 VSS 0.031128f
C8020 DVDD.n2006 VSS 0.031128f
C8021 DVDD.n2007 VSS 0.031128f
C8022 DVDD.n2008 VSS 0.031128f
C8023 DVDD.n2010 VSS 0.031128f
C8024 DVDD.n2011 VSS 0.031128f
C8025 DVDD.n2012 VSS 0.031128f
C8026 DVDD.n2013 VSS 0.031128f
C8027 DVDD.n2015 VSS 0.031128f
C8028 DVDD.n2016 VSS 0.031128f
C8029 DVDD.n2017 VSS 0.031128f
C8030 DVDD.n2018 VSS 0.031128f
C8031 DVDD.n2019 VSS 0.031128f
C8032 DVDD.n2020 VSS 0.031128f
C8033 DVDD.n2022 VSS 0.031128f
C8034 DVDD.n2023 VSS 0.031128f
C8035 DVDD.n2024 VSS 0.031128f
C8036 DVDD.n2025 VSS 0.031128f
C8037 DVDD.n2027 VSS 0.031128f
C8038 DVDD.n2028 VSS 0.031128f
C8039 DVDD.n2029 VSS 0.031128f
C8040 DVDD.n2030 VSS 0.031128f
C8041 DVDD.n2031 VSS 0.031128f
C8042 DVDD.n2032 VSS 0.031128f
C8043 DVDD.n2034 VSS 0.031128f
C8044 DVDD.n2035 VSS 0.031128f
C8045 DVDD.n2036 VSS 0.031128f
C8046 DVDD.n2037 VSS 0.031128f
C8047 DVDD.n2039 VSS 0.031128f
C8048 DVDD.n2040 VSS 0.031128f
C8049 DVDD.n2041 VSS 0.031128f
C8050 DVDD.n2042 VSS 0.031128f
C8051 DVDD.n2043 VSS 0.031128f
C8052 DVDD.n2044 VSS 0.031128f
C8053 DVDD.n2046 VSS 0.031128f
C8054 DVDD.n2047 VSS 0.031128f
C8055 DVDD.n2048 VSS 0.031128f
C8056 DVDD.n2049 VSS 0.031128f
C8057 DVDD.n2051 VSS 0.031128f
C8058 DVDD.n2052 VSS 0.031128f
C8059 DVDD.n2053 VSS 0.031128f
C8060 DVDD.n2054 VSS 0.031128f
C8061 DVDD.n2055 VSS 0.031128f
C8062 DVDD.n2056 VSS 0.031128f
C8063 DVDD.n2058 VSS 0.031128f
C8064 DVDD.n2059 VSS 0.031128f
C8065 DVDD.n2060 VSS 0.031128f
C8066 DVDD.n2061 VSS 0.031128f
C8067 DVDD.n2063 VSS 0.031128f
C8068 DVDD.n2064 VSS 0.031128f
C8069 DVDD.n2065 VSS 0.031128f
C8070 DVDD.n2066 VSS 0.031128f
C8071 DVDD.n2067 VSS 0.031128f
C8072 DVDD.n2068 VSS 0.031128f
C8073 DVDD.n2070 VSS 0.031128f
C8074 DVDD.n2071 VSS 0.031128f
C8075 DVDD.n2072 VSS 0.031128f
C8076 DVDD.n2073 VSS 0.031128f
C8077 DVDD.n2075 VSS 0.031128f
C8078 DVDD.n2076 VSS 0.031128f
C8079 DVDD.n2077 VSS 0.031128f
C8080 DVDD.n2078 VSS 0.031128f
C8081 DVDD.n2079 VSS 0.031128f
C8082 DVDD.n2080 VSS 0.031128f
C8083 DVDD.n2082 VSS 0.031128f
C8084 DVDD.n2083 VSS 0.031128f
C8085 DVDD.n2084 VSS 0.031128f
C8086 DVDD.n2085 VSS 0.031128f
C8087 DVDD.n2087 VSS 0.031128f
C8088 DVDD.n2088 VSS 0.031128f
C8089 DVDD.n2089 VSS 0.031128f
C8090 DVDD.n2090 VSS 0.031128f
C8091 DVDD.n2091 VSS 0.031128f
C8092 DVDD.n2092 VSS 0.031128f
C8093 DVDD.n2094 VSS 0.031128f
C8094 DVDD.n2095 VSS 0.031128f
C8095 DVDD.n2096 VSS 0.031128f
C8096 DVDD.n2097 VSS 0.031128f
C8097 DVDD.n2099 VSS 0.031128f
C8098 DVDD.n2100 VSS 0.031128f
C8099 DVDD.n2101 VSS 0.031128f
C8100 DVDD.n2102 VSS 0.031128f
C8101 DVDD.n2103 VSS 0.031128f
C8102 DVDD.n2104 VSS 0.031128f
C8103 DVDD.n2106 VSS 0.031128f
C8104 DVDD.n2107 VSS 0.031128f
C8105 DVDD.n2108 VSS 0.031128f
C8106 DVDD.n2109 VSS 0.031128f
C8107 DVDD.n2111 VSS 0.031128f
C8108 DVDD.n2112 VSS 0.031128f
C8109 DVDD.n2113 VSS 0.031128f
C8110 DVDD.n2114 VSS 0.031128f
C8111 DVDD.n2115 VSS 0.031128f
C8112 DVDD.n2116 VSS 0.031128f
C8113 DVDD.n2118 VSS 0.031128f
C8114 DVDD.n2119 VSS 0.031128f
C8115 DVDD.n2120 VSS 0.031128f
C8116 DVDD.n2121 VSS 0.031128f
C8117 DVDD.n2123 VSS 0.031128f
C8118 DVDD.n2124 VSS 0.031128f
C8119 DVDD.n2125 VSS 0.031128f
C8120 DVDD.n2126 VSS 0.031128f
C8121 DVDD.n2127 VSS 0.031128f
C8122 DVDD.n2128 VSS 0.031128f
C8123 DVDD.n2130 VSS 0.031128f
C8124 DVDD.n2131 VSS 0.031128f
C8125 DVDD.n2132 VSS 0.031128f
C8126 DVDD.n2133 VSS 0.031128f
C8127 DVDD.n2135 VSS 0.031128f
C8128 DVDD.n2136 VSS 0.031128f
C8129 DVDD.n2137 VSS 0.031128f
C8130 DVDD.n2138 VSS 0.031128f
C8131 DVDD.n2139 VSS 0.031128f
C8132 DVDD.n2140 VSS 0.031128f
C8133 DVDD.n2142 VSS 0.031128f
C8134 DVDD.n2143 VSS 0.031128f
C8135 DVDD.n2144 VSS 0.031128f
C8136 DVDD.n2145 VSS 0.031128f
C8137 DVDD.n2147 VSS 0.031128f
C8138 DVDD.n2148 VSS 0.031128f
C8139 DVDD.n2149 VSS 0.031128f
C8140 DVDD.n2150 VSS 0.031128f
C8141 DVDD.n2151 VSS 0.031128f
C8142 DVDD.n2152 VSS 0.031128f
C8143 DVDD.n2153 VSS 0.019729f
C8144 DVDD.n2154 VSS 0.019729f
C8145 DVDD.n2156 VSS 0.299032f
C8146 DVDD.n2157 VSS 0.039126f
C8147 DVDD.n2158 VSS 0.039126f
C8148 DVDD.n2159 VSS 0.026086f
C8149 DVDD.n2160 VSS 0.036621f
C8150 DVDD.n2161 VSS 0.041931f
C8151 DVDD.n2162 VSS 0.02513f
C8152 DVDD.n2163 VSS 0.041931f
C8153 DVDD.n2164 VSS 0.02513f
C8154 DVDD.n2165 VSS 0.223221f
C8155 DVDD.n2207 VSS 0.019729f
C8156 DVDD.n2208 VSS 0.223221f
C8157 DVDD.n2209 VSS 0.019729f
C8158 DVDD.n2210 VSS 0.522253f
C8159 DVDD.n2211 VSS 0.031128f
C8160 DVDD.n2212 VSS 0.031128f
C8161 DVDD.n2213 VSS 0.031128f
C8162 DVDD.n2214 VSS 0.031128f
C8163 DVDD.n2215 VSS 0.031128f
C8164 DVDD.n2216 VSS 0.031128f
C8165 DVDD.n2217 VSS 0.031128f
C8166 DVDD.n2218 VSS 0.031128f
C8167 DVDD.n2219 VSS 0.031128f
C8168 DVDD.n2220 VSS 0.031128f
C8169 DVDD.n2221 VSS 0.031128f
C8170 DVDD.n2222 VSS 0.031128f
C8171 DVDD.n2223 VSS 0.031128f
C8172 DVDD.n2224 VSS 0.031128f
C8173 DVDD.n2225 VSS 0.031128f
C8174 DVDD.n2226 VSS 0.031128f
C8175 DVDD.n2227 VSS 0.031128f
C8176 DVDD.n2228 VSS 0.031128f
C8177 DVDD.n2229 VSS 0.031128f
C8178 DVDD.n2230 VSS 0.031128f
C8179 DVDD.n2231 VSS 0.031128f
C8180 DVDD.n2232 VSS 0.031128f
C8181 DVDD.n2233 VSS 0.031128f
C8182 DVDD.n2234 VSS 0.031128f
C8183 DVDD.n2235 VSS 0.031128f
C8184 DVDD.n2236 VSS 0.031128f
C8185 DVDD.n2237 VSS 0.031128f
C8186 DVDD.n2238 VSS 0.031128f
C8187 DVDD.n2239 VSS 0.031128f
C8188 DVDD.n2240 VSS 0.031128f
C8189 DVDD.n2241 VSS 0.031128f
C8190 DVDD.n2242 VSS 0.031128f
C8191 DVDD.n2243 VSS 0.031128f
C8192 DVDD.n2244 VSS 0.031128f
C8193 DVDD.n2245 VSS 0.031128f
C8194 DVDD.n2246 VSS 0.031128f
C8195 DVDD.n2247 VSS 0.031128f
C8196 DVDD.n2248 VSS 0.031128f
C8197 DVDD.n2249 VSS 0.031128f
C8198 DVDD.n2250 VSS 0.031128f
C8199 DVDD.n2252 VSS 0.031128f
C8200 DVDD.n2253 VSS 0.031128f
C8201 DVDD.n2254 VSS 0.039516f
C8202 DVDD.n2255 VSS 0.038426f
C8203 DVDD.n2265 VSS 0.025624f
C8204 DVDD.n2266 VSS 0.025624f
C8205 DVDD.n2267 VSS 0.142744f
C8206 DVDD.n2268 VSS 1.16224f
C8207 DVDD.n2269 VSS 0.025624f
C8208 DVDD.n2271 VSS 0.025624f
C8209 DVDD.n2272 VSS 0.025624f
C8210 DVDD.n2273 VSS 0.025624f
C8211 DVDD.n2274 VSS 0.025624f
C8212 DVDD.n2275 VSS 0.025624f
C8213 DVDD.n2276 VSS 0.025624f
C8214 DVDD.n2277 VSS 0.025624f
C8215 DVDD.n2278 VSS 0.025624f
C8216 DVDD.n2279 VSS 0.142744f
C8217 DVDD.n2281 VSS 0.468543f
C8218 DVDD.n2282 VSS 1.04547f
C8219 DVDD.n2284 VSS 0.025624f
C8220 DVDD.n2285 VSS 0.025624f
C8221 DVDD.n2286 VSS 0.025624f
C8222 DVDD.n2287 VSS 0.025624f
C8223 DVDD.n2288 VSS 0.025624f
C8224 DVDD.n2289 VSS 0.025624f
C8225 DVDD.n2290 VSS 0.025624f
C8226 DVDD.n2291 VSS 0.05801f
C8227 DVDD.n2292 VSS 3.49331f
C8228 DVDD.n2293 VSS 0.05801f
C8229 DVDD.n2294 VSS 0.081946f
C8230 DVDD.n2296 VSS 0.113666f
C8231 DVDD.n2297 VSS 0.025624f
C8232 DVDD.n2298 VSS 0.025624f
C8233 DVDD.n2299 VSS 0.025624f
C8234 DVDD.n2300 VSS 0.025624f
C8235 DVDD.n2301 VSS 0.025624f
C8236 DVDD.n2302 VSS 0.025624f
C8237 DVDD.n2303 VSS 0.025624f
C8238 DVDD.n2304 VSS 0.025624f
C8239 DVDD.n2305 VSS 0.025624f
C8240 DVDD.n2306 VSS 0.071372f
C8241 DVDD.n2308 VSS 0.025624f
C8242 DVDD.n2310 VSS 0.025624f
C8243 DVDD.n2312 VSS 0.025624f
C8244 DVDD.n2314 VSS 0.025624f
C8245 DVDD.n2316 VSS 0.025624f
C8246 DVDD.n2318 VSS 0.025624f
C8247 DVDD.n2320 VSS 0.025624f
C8248 DVDD.n2322 VSS 0.025624f
C8249 DVDD.n2324 VSS 0.063349f
C8250 DVDD.n2325 VSS 0.071372f
C8251 DVDD.n2335 VSS 0.123789f
C8252 DVDD.n2336 VSS 0.330748f
C8253 DVDD.n2337 VSS 0.137328f
C8254 DVDD.n2338 VSS 0.137328f
C8255 DVDD.n2339 VSS 0.121855f
C8256 DVDD.n2340 VSS 0.137328f
C8257 DVDD.n2341 VSS 0.137328f
C8258 DVDD.n2342 VSS 0.137328f
C8259 DVDD.n2343 VSS 0.135394f
C8260 DVDD.n2344 VSS 0.137328f
C8261 DVDD.n2345 VSS 0.137328f
C8262 DVDD.n2346 VSS 0.137328f
C8263 DVDD.n2347 VSS 0.13346f
C8264 DVDD.n2348 VSS 0.137328f
C8265 DVDD.n2349 VSS 0.11992f
C8266 DVDD.n2350 VSS 1.37325f
C8267 DVDD.n2351 VSS 0.163891f
C8268 DVDD.n2352 VSS 0.163891f
C8269 DVDD.n2353 VSS 0.163891f
C8270 DVDD.n2354 VSS 0.163891f
C8271 DVDD.n2355 VSS 0.085911f
C8272 DVDD.n2356 VSS 0.163891f
C8273 DVDD.n2357 VSS 0.091198f
C8274 DVDD.n2358 VSS 0.163891f
C8275 DVDD.n2361 VSS 0.244515f
C8276 DVDD.n2362 VSS 0.19342f
C8277 DVDD.n2363 VSS 0.149352f
C8278 DVDD.n2365 VSS 0.163891f
C8279 DVDD.n2366 VSS 0.154639f
C8280 DVDD.n2368 VSS 0.163891f
C8281 DVDD.n2369 VSS 0.159926f
C8282 DVDD.n2371 VSS 0.163891f
C8283 DVDD.n2373 VSS 0.163891f
C8284 DVDD.n2375 VSS 0.163891f
C8285 DVDD.n2377 VSS 0.163891f
C8286 DVDD.n2378 VSS 0.11992f
C8287 DVDD.n2379 VSS 0.274656f
C8288 DVDD.n2380 VSS 0.274656f
C8289 DVDD.n2381 VSS 0.274656f
C8290 DVDD.n2382 VSS 0.274656f
C8291 DVDD.n2383 VSS 0.274656f
C8292 DVDD.n2384 VSS 0.274656f
C8293 DVDD.n2385 VSS 0.137328f
C8294 DVDD.n2386 VSS 0.274656f
C8295 DVDD.n2387 VSS 0.274656f
C8296 DVDD.n2388 VSS 0.274656f
C8297 DVDD.n2389 VSS 0.274656f
C8298 DVDD.n2390 VSS 0.071372f
C8299 DVDD.n2391 VSS 1.37325f
C8300 DVDD.n2392 VSS 0.163891f
C8301 DVDD.n2393 VSS 0.153317f
C8302 DVDD.n2394 VSS 0.163891f
C8303 DVDD.n2395 VSS 0.163891f
C8304 DVDD.n2396 VSS 0.163891f
C8305 DVDD.n2397 VSS 0.085911f
C8306 DVDD.n2398 VSS 0.163891f
C8307 DVDD.n2399 VSS 0.091198f
C8308 DVDD.n2400 VSS 0.163891f
C8309 DVDD.n2402 VSS 0.149352f
C8310 DVDD.n2403 VSS 0.163891f
C8311 DVDD.n2404 VSS 0.154639f
C8312 DVDD.n2405 VSS 0.163891f
C8313 DVDD.n2406 VSS 0.159926f
C8314 DVDD.n2407 VSS 0.163891f
C8315 DVDD.n2408 VSS 0.163891f
C8316 DVDD.n2409 VSS 0.163891f
C8317 DVDD.n2410 VSS 0.163891f
C8318 DVDD.n2411 VSS 0.163891f
C8319 DVDD.n2412 VSS 0.113666f
C8320 DVDD.n2413 VSS 0.081946f
C8321 DVDD.n2424 VSS 0.137328f
C8322 DVDD.n2432 VSS 0.137328f
C8323 DVDD.n2433 VSS 0.131525f
C8324 DVDD.n2434 VSS 0.137328f
C8325 DVDD.n2435 VSS 0.137328f
C8326 DVDD.n2436 VSS 0.137328f
C8327 DVDD.n2437 VSS 0.129591f
C8328 DVDD.n2448 VSS 0.025624f
C8329 DVDD.n2449 VSS 0.025624f
C8330 DVDD.n2450 VSS 0.025624f
C8331 DVDD.n2451 VSS 0.025624f
C8332 DVDD.n2452 VSS 0.025624f
C8333 DVDD.n2453 VSS 0.025624f
C8334 DVDD.n2454 VSS 0.025624f
C8335 DVDD.n2455 VSS 0.025624f
C8336 DVDD.n2456 VSS 0.025624f
C8337 DVDD.n2458 VSS 0.025624f
C8338 DVDD.n2460 VSS 0.025624f
C8339 DVDD.n2462 VSS 0.025624f
C8340 DVDD.n2464 VSS 0.025624f
C8341 DVDD.n2466 VSS 0.025624f
C8342 DVDD.n2468 VSS 0.025624f
C8343 DVDD.n2470 VSS 0.025624f
C8344 DVDD.n2472 VSS 0.025624f
C8345 DVDD.n2473 VSS 0.081946f
C8346 DVDD.n2474 VSS 0.098464f
C8347 DVDD.n2475 VSS 0.081946f
C8348 DVDD.n2476 VSS 0.11992f
C8349 DVDD.n2477 VSS 0.137328f
C8350 DVDD.n2478 VSS 0.137328f
C8351 DVDD.n2479 VSS 0.137328f
C8352 DVDD.n2480 VSS 0.125723f
C8353 DVDD.n2481 VSS 0.137328f
C8354 DVDD.n2482 VSS 0.137328f
C8355 DVDD.n2483 VSS 0.11992f
C8356 DVDD.n2485 VSS 0.244515f
C8357 DVDD.n2486 VSS 0.274656f
C8358 DVDD.n2487 VSS 0.274656f
C8359 DVDD.n2488 VSS 0.274656f
C8360 DVDD.n2489 VSS 0.11992f
C8361 DVDD.n2490 VSS 0.274656f
C8362 DVDD.n2491 VSS 0.274656f
C8363 DVDD.n2492 VSS 0.11992f
C8364 DVDD.n2493 VSS 0.274656f
C8365 DVDD.n2494 VSS 0.274656f
C8366 DVDD.n2495 VSS 0.274656f
C8367 DVDD.n2496 VSS 0.11992f
C8368 DVDD.n2497 VSS 0.274656f
C8369 DVDD.n2498 VSS 0.11992f
C8370 DVDD.n2499 VSS 0.274656f
C8371 DVDD.n2500 VSS 0.274656f
C8372 DVDD.n2501 VSS 0.274656f
C8373 DVDD.n2502 VSS 0.274656f
C8374 DVDD.n2503 VSS 0.11992f
C8375 DVDD.n2504 VSS 0.274656f
C8376 DVDD.n2505 VSS 0.11992f
C8377 DVDD.n2506 VSS 0.274656f
C8378 DVDD.n2507 VSS 0.11992f
C8379 DVDD.n2508 VSS 0.274656f
C8380 DVDD.n2509 VSS 0.274656f
C8381 DVDD.n2510 VSS 0.274656f
C8382 DVDD.n2511 VSS 0.274656f
C8383 DVDD.n2512 VSS 0.11992f
C8384 DVDD.n2513 VSS 0.274656f
C8385 DVDD.n2514 VSS 0.11992f
C8386 DVDD.n2515 VSS 0.274656f
C8387 DVDD.n2516 VSS 0.11992f
C8388 DVDD.n2517 VSS 0.274656f
C8389 DVDD.n2518 VSS 0.274656f
C8390 DVDD.n2519 VSS 0.274656f
C8391 DVDD.n2520 VSS 0.274656f
C8392 DVDD.n2521 VSS 0.274656f
C8393 DVDD.n2522 VSS 0.160538f
C8394 DVDD.n2523 VSS 0.330748f
C8395 DVDD.n2524 VSS 0.251446f
C8396 DVDD.n2525 VSS 0.524168f
C8397 DVDD.n2526 VSS 0.160538f
C8398 DVDD.n2527 VSS 0.524168f
C8399 DVDD.n2528 VSS 0.274656f
C8400 DVDD.n2529 VSS 0.274656f
C8401 DVDD.n2530 VSS 0.274656f
C8402 DVDD.n2531 VSS 0.274656f
C8403 DVDD.n2532 VSS 0.274656f
C8404 DVDD.n2533 VSS 0.274656f
C8405 DVDD.n2534 VSS 0.274656f
C8406 DVDD.n2535 VSS 0.274656f
C8407 DVDD.n2536 VSS 0.274656f
C8408 DVDD.n2537 VSS 0.247577f
C8409 DVDD.n2538 VSS 0.030947f
C8410 DVDD.n2539 VSS 1.26626f
C8411 DVDD.n2540 VSS 0.355263f
C8412 DVDD.n2541 VSS 0.11992f
C8413 DVDD.n2542 VSS 0.274656f
C8414 DVDD.n2543 VSS 0.057059f
C8415 DVDD.n2544 VSS 0.164407f
C8416 DVDD.n2545 VSS 0.11992f
C8417 DVDD.n2546 VSS 0.247577f
C8418 DVDD.n2547 VSS 0.11992f
C8419 DVDD.n2548 VSS 0.274656f
C8420 DVDD.n2549 VSS 0.11992f
C8421 DVDD.n2550 VSS 0.274656f
C8422 DVDD.n2551 VSS 0.11992f
C8423 DVDD.n2552 VSS 0.274656f
C8424 DVDD.n2553 VSS 0.11992f
C8425 DVDD.n2554 VSS 0.274656f
C8426 DVDD.n2555 VSS 0.11992f
C8427 DVDD.n2556 VSS 0.274656f
C8428 DVDD.n2557 VSS 0.11992f
C8429 DVDD.n2558 VSS 0.274656f
C8430 DVDD.n2559 VSS 0.11992f
C8431 DVDD.n2560 VSS 0.274656f
C8432 DVDD.n2561 VSS 0.11992f
C8433 DVDD.n2562 VSS 0.274656f
C8434 DVDD.n2563 VSS 0.221466f
C8435 DVDD.n2564 VSS 0.274656f
C8436 DVDD.n2565 VSS 0.251446f
C8437 DVDD.n2566 VSS 0.251446f
C8438 DVDD.n2567 VSS 0.330748f
C8439 DVDD.n2568 VSS 0.524168f
C8440 DVDD.n2569 VSS 0.274656f
C8441 DVDD.n2570 VSS 0.274656f
C8442 DVDD.n2571 VSS 0.11992f
C8443 DVDD.n2572 VSS 0.085911f
C8444 DVDD.n2573 VSS 0.163891f
C8445 DVDD.n2574 VSS 0.091198f
C8446 DVDD.n2575 VSS 0.163891f
C8447 DVDD.n2576 VSS 0.096484f
C8448 DVDD.n2577 VSS 0.163891f
C8449 DVDD.n2578 VSS 0.101771f
C8450 DVDD.n2579 VSS 0.163891f
C8451 DVDD.n2580 VSS 0.107058f
C8452 DVDD.n2581 VSS 0.163891f
C8453 DVDD.n2582 VSS 0.112345f
C8454 DVDD.n2583 VSS 0.210151f
C8455 DVDD.n2584 VSS 0.163891f
C8456 DVDD.n2585 VSS 0.133492f
C8457 DVDD.n2586 VSS 0.163891f
C8458 DVDD.n2587 VSS 0.138779f
C8459 DVDD.n2588 VSS 0.163891f
C8460 DVDD.n2589 VSS 0.144066f
C8461 DVDD.n2590 VSS 0.163891f
C8462 DVDD.n2591 VSS 0.149352f
C8463 DVDD.n2592 VSS 0.163891f
C8464 DVDD.n2593 VSS 0.154639f
C8465 DVDD.n2594 VSS 0.163891f
C8466 DVDD.n2606 VSS 0.137328f
C8467 DVDD.n2613 VSS 0.137328f
C8468 DVDD.n2614 VSS 0.131525f
C8469 DVDD.n2615 VSS 0.137328f
C8470 DVDD.n2616 VSS 0.137328f
C8471 DVDD.n2617 VSS 0.137328f
C8472 DVDD.n2618 VSS 0.129591f
C8473 DVDD.n2619 VSS 0.137328f
C8474 DVDD.n2620 VSS 0.198722f
C8475 DVDD.n2622 VSS 0.127657f
C8476 DVDD.n2623 VSS 0.137328f
C8477 DVDD.n2624 VSS 0.137328f
C8478 DVDD.n2625 VSS 0.137328f
C8479 DVDD.n2627 VSS 0.125723f
C8480 DVDD.n2628 VSS 0.137328f
C8481 DVDD.n2629 VSS 0.11992f
C8482 DVDD.n2630 VSS 0.274656f
C8483 DVDD.n2631 VSS 0.274656f
C8484 DVDD.n2632 VSS 0.11992f
C8485 DVDD.n2633 VSS 0.274656f
C8486 DVDD.n2634 VSS 0.274656f
C8487 DVDD.n2635 VSS 0.11992f
C8488 DVDD.n2636 VSS 0.274656f
C8489 DVDD.n2637 VSS 0.274656f
C8490 DVDD.n2638 VSS 0.274656f
C8491 DVDD.n2639 VSS 0.274656f
C8492 DVDD.n2640 VSS 0.19342f
C8493 DVDD.n2641 VSS 0.274656f
C8494 DVDD.n2642 VSS 0.274656f
C8495 DVDD.n2643 VSS 0.274656f
C8496 DVDD.n2644 VSS 0.137328f
C8497 DVDD.n2645 VSS 0.085911f
C8498 DVDD.n2646 VSS 0.163891f
C8499 DVDD.n2647 VSS 0.091198f
C8500 DVDD.n2648 VSS 0.163891f
C8501 DVDD.n2649 VSS 0.096484f
C8502 DVDD.n2650 VSS 0.163891f
C8503 DVDD.n2651 VSS 0.101771f
C8504 DVDD.n2652 VSS 0.163891f
C8505 DVDD.n2653 VSS 0.107058f
C8506 DVDD.n2654 VSS 0.163891f
C8507 DVDD.n2655 VSS 0.112345f
C8508 DVDD.n2656 VSS 0.210151f
C8509 DVDD.n2658 VSS 0.163891f
C8510 DVDD.n2660 VSS 0.133492f
C8511 DVDD.n2662 VSS 0.163891f
C8512 DVDD.n2664 VSS 0.138779f
C8513 DVDD.n2666 VSS 0.163891f
C8514 DVDD.n2668 VSS 0.144066f
C8515 DVDD.n2670 VSS 0.163891f
C8516 DVDD.n2672 VSS 0.149352f
C8517 DVDD.n2674 VSS 0.163891f
C8518 DVDD.n2676 VSS 0.154639f
C8519 DVDD.n2678 VSS 0.163891f
C8520 DVDD.n2685 VSS 0.123789f
C8521 DVDD.n2686 VSS 0.524168f
C8522 DVDD.n2687 VSS 0.137328f
C8523 DVDD.n2688 VSS 0.137328f
C8524 DVDD.n2689 VSS 0.121855f
C8525 DVDD.n2690 VSS 0.137328f
C8526 DVDD.n2691 VSS 0.137328f
C8527 DVDD.n2692 VSS 0.081946f
C8528 DVDD.n2693 VSS 0.137328f
C8529 DVDD.n2695 VSS 0.135394f
C8530 DVDD.n2696 VSS 0.137328f
C8531 DVDD.n2697 VSS 0.137328f
C8532 DVDD.n2698 VSS 0.137328f
C8533 DVDD.n2700 VSS 0.13346f
C8534 DVDD.n2701 VSS 0.11992f
C8535 DVDD.n2702 VSS 0.243709f
C8536 DVDD.n2703 VSS 0.330748f
C8537 DVDD.n2704 VSS 0.168275f
C8538 DVDD.n2705 VSS 0.330748f
C8539 DVDD.n2706 VSS 0.168275f
C8540 DVDD.n2707 VSS 0.274656f
C8541 DVDD.n2708 VSS 0.524168f
C8542 DVDD.n2709 VSS 0.274656f
C8543 DVDD.n2710 VSS 0.524168f
C8544 DVDD.n2711 VSS 0.163891f
C8545 DVDD.n2712 VSS 0.107058f
C8546 DVDD.n2713 VSS 0.163891f
C8547 DVDD.n2714 VSS 0.163891f
C8548 DVDD.n2715 VSS 0.163891f
C8549 DVDD.n2716 VSS 0.107058f
C8550 DVDD.n2717 VSS 0.163891f
C8551 DVDD.n2718 VSS 0.112345f
C8552 DVDD.n2719 VSS 0.163891f
C8553 DVDD.n2720 VSS 0.117632f
C8554 DVDD.n2721 VSS 0.163891f
C8555 DVDD.n2723 VSS 0.122918f
C8556 DVDD.n2724 VSS 0.163891f
C8557 DVDD.n2725 VSS 0.128205f
C8558 DVDD.n2726 VSS 0.163891f
C8559 DVDD.n2727 VSS 0.133492f
C8560 DVDD.n2728 VSS 0.163891f
C8561 DVDD.n2729 VSS 0.138779f
C8562 DVDD.n2730 VSS 0.163891f
C8563 DVDD.n2731 VSS 0.163891f
C8564 DVDD.n2732 VSS 0.163891f
C8565 DVDD.n2733 VSS 0.138779f
C8566 DVDD.n2734 VSS 0.229976f
C8567 DVDD.n2746 VSS 0.137328f
C8568 DVDD.n2748 VSS 0.137328f
C8569 DVDD.n2749 VSS 0.137328f
C8570 DVDD.n2750 VSS 0.121855f
C8571 DVDD.n2751 VSS 0.137328f
C8572 DVDD.n2752 VSS 0.137328f
C8573 DVDD.n2753 VSS 0.137328f
C8574 DVDD.n2754 VSS 0.135394f
C8575 DVDD.n2755 VSS 0.137328f
C8576 DVDD.n2756 VSS 0.137328f
C8577 DVDD.n2757 VSS 0.137328f
C8578 DVDD.n2764 VSS 0.123789f
C8579 DVDD.n2765 VSS 0.11992f
C8580 DVDD.n2766 VSS 0.137328f
C8581 DVDD.n2767 VSS 0.11992f
C8582 DVDD.n2769 VSS 0.270949f
C8583 DVDD.n2770 VSS 0.274656f
C8584 DVDD.n2771 VSS 0.274656f
C8585 DVDD.n2772 VSS 0.11992f
C8586 DVDD.n2773 VSS 0.274656f
C8587 DVDD.n2774 VSS 0.274656f
C8588 DVDD.n2775 VSS 0.274656f
C8589 DVDD.n2776 VSS 0.274656f
C8590 DVDD.n2777 VSS 0.274656f
C8591 DVDD.n2778 VSS 0.274656f
C8592 DVDD.n2779 VSS 0.274656f
C8593 DVDD.n2780 VSS 0.163891f
C8594 DVDD.n2781 VSS 0.107058f
C8595 DVDD.n2782 VSS 0.163891f
C8596 DVDD.n2783 VSS 0.163891f
C8597 DVDD.n2784 VSS 0.163891f
C8598 DVDD.n2785 VSS 0.107058f
C8599 DVDD.n2786 VSS 0.163891f
C8600 DVDD.n2787 VSS 0.112345f
C8601 DVDD.n2788 VSS 0.163891f
C8602 DVDD.n2789 VSS 0.117632f
C8603 DVDD.n2790 VSS 0.163891f
C8604 DVDD.n2791 VSS 0.270949f
C8605 DVDD.n2792 VSS 0.11992f
C8606 DVDD.n2793 VSS 0.122918f
C8607 DVDD.n2794 VSS 0.163891f
C8608 DVDD.n2795 VSS 0.128205f
C8609 DVDD.n2796 VSS 0.163891f
C8610 DVDD.n2797 VSS 0.133492f
C8611 DVDD.n2798 VSS 0.163891f
C8612 DVDD.n2799 VSS 0.138779f
C8613 DVDD.n2800 VSS 0.163891f
C8614 DVDD.n2801 VSS 0.163891f
C8615 DVDD.n2802 VSS 0.163891f
C8616 DVDD.n2803 VSS 0.138779f
C8617 DVDD.n2804 VSS 0.346752f
C8618 DVDD.n2816 VSS 0.137328f
C8619 DVDD.n2818 VSS 0.131525f
C8620 DVDD.n2819 VSS 0.137328f
C8621 DVDD.n2820 VSS 0.137328f
C8622 DVDD.n2821 VSS 0.137328f
C8623 DVDD.n2822 VSS 0.129591f
C8624 DVDD.n2824 VSS 0.127657f
C8625 DVDD.n2825 VSS 0.137328f
C8626 DVDD.n2826 VSS 0.137328f
C8627 DVDD.n2827 VSS 0.137328f
C8628 DVDD.n2829 VSS 0.125723f
C8629 DVDD.n2830 VSS 0.137328f
C8630 DVDD.n2831 VSS 0.137328f
C8631 DVDD.n2832 VSS 0.11992f
C8632 DVDD.n2833 VSS 0.274656f
C8633 DVDD.n2834 VSS 0.274656f
C8634 DVDD.n2835 VSS 0.274656f
C8635 DVDD.n2836 VSS 0.11992f
C8636 DVDD.n2837 VSS 0.274656f
C8637 DVDD.n2838 VSS 0.274656f
C8638 DVDD.n2839 VSS 0.11992f
C8639 DVDD.n2840 VSS 0.274656f
C8640 DVDD.n2841 VSS 0.274656f
C8641 DVDD.n2842 VSS 0.274656f
C8642 DVDD.n2843 VSS 0.274656f
C8643 DVDD.n2844 VSS 0.274656f
C8644 DVDD.n2845 VSS 0.274656f
C8645 DVDD.n2846 VSS 0.11992f
C8646 DVDD.n2847 VSS 0.274656f
C8647 DVDD.n2848 VSS 0.11992f
C8648 DVDD.n2849 VSS 0.274656f
C8649 DVDD.n2850 VSS 0.11992f
C8650 DVDD.n2851 VSS 0.274656f
C8651 DVDD.n2852 VSS 0.274656f
C8652 DVDD.n2853 VSS 0.274656f
C8653 DVDD.n2854 VSS 0.274656f
C8654 DVDD.n2855 VSS 0.11992f
C8655 DVDD.n2856 VSS 0.274656f
C8656 DVDD.n2857 VSS 0.11992f
C8657 DVDD.n2858 VSS 0.274656f
C8658 DVDD.n2859 VSS 0.11992f
C8659 DVDD.n2860 VSS 0.274656f
C8660 DVDD.n2861 VSS 0.274656f
C8661 DVDD.n2862 VSS 0.274656f
C8662 DVDD.n2863 VSS 0.274656f
C8663 DVDD.n2864 VSS 0.274656f
C8664 DVDD.n2865 VSS 0.11992f
C8665 DVDD.n2872 VSS 0.137328f
C8666 DVDD.n2873 VSS 0.11992f
C8667 DVDD.n2874 VSS 0.274656f
C8668 DVDD.n2875 VSS 0.11992f
C8669 DVDD.n2876 VSS 0.274656f
C8670 DVDD.n2877 VSS 0.274656f
C8671 DVDD.n2878 VSS 0.274656f
C8672 DVDD.n2879 VSS 0.274656f
C8673 DVDD.n2880 VSS 0.274656f
C8674 DVDD.n2881 VSS 0.160538f
C8675 DVDD.n2882 VSS 0.160538f
C8676 DVDD.n2883 VSS 0.251446f
C8677 DVDD.n2884 VSS 0.274656f
C8678 DVDD.n2885 VSS 0.274656f
C8679 DVDD.n2886 VSS 0.274656f
C8680 DVDD.n2887 VSS 0.274656f
C8681 DVDD.n2888 VSS 0.274656f
C8682 DVDD.n2889 VSS 0.274656f
C8683 DVDD.n2890 VSS 0.274656f
C8684 DVDD.n2891 VSS 0.274656f
C8685 DVDD.n2892 VSS 0.274656f
C8686 DVDD.n2893 VSS 0.247577f
C8687 DVDD.n2894 VSS 0.030947f
C8688 DVDD.n2895 VSS 1.26626f
C8689 DVDD.n2896 VSS 0.355263f
C8690 DVDD.n2897 VSS 0.11992f
C8691 DVDD.n2898 VSS 0.274656f
C8692 DVDD.n2899 VSS 0.057059f
C8693 DVDD.n2900 VSS 0.164407f
C8694 DVDD.n2901 VSS 0.11992f
C8695 DVDD.n2902 VSS 0.247577f
C8696 DVDD.n2903 VSS 0.11992f
C8697 DVDD.n2904 VSS 0.274656f
C8698 DVDD.n2905 VSS 0.11992f
C8699 DVDD.n2906 VSS 0.274656f
C8700 DVDD.n2907 VSS 0.11992f
C8701 DVDD.n2908 VSS 0.274656f
C8702 DVDD.n2909 VSS 0.11992f
C8703 DVDD.n2910 VSS 0.274656f
C8704 DVDD.n2911 VSS 0.11992f
C8705 DVDD.n2912 VSS 0.274656f
C8706 DVDD.n2913 VSS 0.11992f
C8707 DVDD.n2914 VSS 0.274656f
C8708 DVDD.n2915 VSS 0.11992f
C8709 DVDD.n2916 VSS 0.274656f
C8710 DVDD.n2917 VSS 0.11992f
C8711 DVDD.n2918 VSS 0.274656f
C8712 DVDD.n2919 VSS 0.274656f
C8713 DVDD.n2920 VSS 0.235972f
C8714 DVDD.n2921 VSS 0.274656f
C8715 DVDD.n2922 VSS 0.274656f
C8716 DVDD.n2923 VSS 0.274656f
C8717 DVDD.n2924 VSS 0.137328f
C8718 DVDD.n2925 VSS 0.112345f
C8719 DVDD.n2926 VSS 0.281523f
C8720 DVDD.n2927 VSS 0.163891f
C8721 DVDD.n2928 VSS 0.128205f
C8722 DVDD.n2929 VSS 0.163891f
C8723 DVDD.n2930 VSS 0.122918f
C8724 DVDD.n2931 VSS 0.163891f
C8725 DVDD.n2932 VSS 0.128205f
C8726 DVDD.n2933 VSS 0.163891f
C8727 DVDD.n2934 VSS 0.163891f
C8728 DVDD.n2935 VSS 0.138779f
C8729 DVDD.n2936 VSS 0.183717f
C8730 DVDD.n2938 VSS 0.163891f
C8731 DVDD.n2940 VSS 0.163891f
C8732 DVDD.n2941 VSS 0.133492f
C8733 DVDD.n2943 VSS 0.163891f
C8734 DVDD.n2945 VSS 0.163891f
C8735 DVDD.n2946 VSS 0.122918f
C8736 DVDD.n2948 VSS 0.163891f
C8737 DVDD.n2950 VSS 0.117632f
C8738 DVDD.n2952 VSS 0.163891f
C8739 DVDD.n2954 VSS 0.112345f
C8740 DVDD.n2955 VSS 0.117632f
C8741 DVDD.n2957 VSS 0.131525f
C8742 DVDD.n2958 VSS 0.137328f
C8743 DVDD.n2959 VSS 0.137328f
C8744 DVDD.n2960 VSS 0.137328f
C8745 DVDD.n2961 VSS 0.129591f
C8746 DVDD.n2962 VSS 0.137328f
C8747 DVDD.n2963 VSS 0.198722f
C8748 DVDD.n2965 VSS 0.127657f
C8749 DVDD.n2966 VSS 0.137328f
C8750 DVDD.n2967 VSS 0.137328f
C8751 DVDD.n2968 VSS 0.137328f
C8752 DVDD.n2970 VSS 0.125723f
C8753 DVDD.n2971 VSS 0.137328f
C8754 DVDD.n2980 VSS 0.137328f
C8755 DVDD.n2981 VSS 0.11992f
C8756 DVDD.n2982 VSS 0.274656f
C8757 DVDD.n2983 VSS 0.274656f
C8758 DVDD.n2984 VSS 0.11992f
C8759 DVDD.n2985 VSS 0.274656f
C8760 DVDD.n2986 VSS 0.274656f
C8761 DVDD.n2987 VSS 0.11992f
C8762 DVDD.n2988 VSS 0.274656f
C8763 DVDD.n2989 VSS 0.274656f
C8764 DVDD.n2990 VSS 0.274656f
C8765 DVDD.n2991 VSS 0.19342f
C8766 DVDD.n2992 VSS 0.274656f
C8767 DVDD.n2993 VSS 0.274656f
C8768 DVDD.n2994 VSS 0.274656f
C8769 DVDD.n2995 VSS 0.137328f
C8770 DVDD.n2996 VSS 0.112345f
C8771 DVDD.n2997 VSS 0.281523f
C8772 DVDD.n2998 VSS 0.163891f
C8773 DVDD.n2999 VSS 0.128205f
C8774 DVDD.n3000 VSS 0.163891f
C8775 DVDD.n3001 VSS 0.122918f
C8776 DVDD.n3002 VSS 0.163891f
C8777 DVDD.n3003 VSS 0.128205f
C8778 DVDD.n3004 VSS 0.163891f
C8779 DVDD.n3005 VSS 0.163891f
C8780 DVDD.n3006 VSS 0.138779f
C8781 DVDD.n3007 VSS 0.183717f
C8782 DVDD.n3009 VSS 0.163891f
C8783 DVDD.n3011 VSS 0.163891f
C8784 DVDD.n3012 VSS 0.133492f
C8785 DVDD.n3014 VSS 0.163891f
C8786 DVDD.n3016 VSS 0.163891f
C8787 DVDD.n3017 VSS 0.122918f
C8788 DVDD.n3019 VSS 0.163891f
C8789 DVDD.n3020 VSS 0.117632f
C8790 DVDD.n3022 VSS 0.163891f
C8791 DVDD.n3023 VSS 0.112345f
C8792 DVDD.n3024 VSS 0.117632f
C8793 DVDD.n3026 VSS 0.123789f
C8794 DVDD.n3027 VSS 0.330748f
C8795 DVDD.n3028 VSS 0.137328f
C8796 DVDD.n3029 VSS 0.137328f
C8797 DVDD.n3030 VSS 0.121855f
C8798 DVDD.n3031 VSS 0.137328f
C8799 DVDD.n3032 VSS 0.081946f
C8800 DVDD.n3033 VSS 0.137328f
C8801 DVDD.n3035 VSS 0.135394f
C8802 DVDD.n3036 VSS 0.137328f
C8803 DVDD.n3037 VSS 0.137328f
C8804 DVDD.n3038 VSS 0.137328f
C8805 DVDD.n3040 VSS 0.13346f
C8806 DVDD.n3041 VSS 0.11992f
C8807 DVDD.n3042 VSS 0.274656f
C8808 DVDD.n3043 VSS 0.274656f
C8809 DVDD.n3044 VSS 0.11992f
C8810 DVDD.n3045 VSS 0.274656f
C8811 DVDD.n3046 VSS 0.274656f
C8812 DVDD.n3047 VSS 0.274656f
C8813 DVDD.n3048 VSS 0.274656f
C8814 DVDD.n3049 VSS 0.274656f
C8815 DVDD.n3050 VSS 0.274656f
C8816 DVDD.n3051 VSS 0.274656f
C8817 DVDD.n3052 VSS 0.274656f
C8818 DVDD.n3053 VSS 0.137328f
C8819 DVDD.n3054 VSS 0.274656f
C8820 DVDD.n3055 VSS 0.274656f
C8821 DVDD.n3056 VSS 0.274656f
C8822 DVDD.n3057 VSS 0.137328f
C8823 DVDD.n3058 VSS 0.112345f
C8824 DVDD.n3059 VSS 0.281523f
C8825 DVDD.n3064 VSS 0.128205f
C8826 DVDD.n3066 VSS 0.138779f
C8827 DVDD.n3068 VSS 0.11992f
C8828 DVDD.n3070 VSS 0.133492f
C8829 DVDD.n3072 VSS 0.122918f
C8830 DVDD.n3073 VSS 0.117632f
C8831 DVDD.n3075 VSS 0.137328f
C8832 DVDD.n3076 VSS 0.137328f
C8833 DVDD.n3077 VSS 0.137328f
C8834 DVDD.n3078 VSS 0.129591f
C8835 DVDD.n3079 VSS 0.137328f
C8836 DVDD.n3080 VSS 0.137328f
C8837 DVDD.n3081 VSS 0.081946f
C8838 DVDD.n3082 VSS 0.137328f
C8839 DVDD.n3083 VSS 0.127657f
C8840 DVDD.n3084 VSS 0.098644f
C8841 DVDD.n3085 VSS 0.137328f
C8842 DVDD.n3086 VSS 0.137328f
C8843 DVDD.n3087 VSS 0.11992f
C8844 DVDD.n3088 VSS 0.163891f
C8845 DVDD.n3089 VSS 0.128205f
C8846 DVDD.n3090 VSS 0.163891f
C8847 DVDD.n3091 VSS 0.122918f
C8848 DVDD.n3092 VSS 0.163891f
C8849 DVDD.n3093 VSS 0.163891f
C8850 DVDD.n3094 VSS 0.163891f
C8851 DVDD.n3096 VSS 0.163891f
C8852 DVDD.n3097 VSS 0.163891f
C8853 DVDD.n3098 VSS 0.163891f
C8854 DVDD.n3099 VSS 0.163891f
C8855 DVDD.n3100 VSS 0.163891f
C8856 DVDD.n3101 VSS 0.117632f
C8857 DVDD.n3102 VSS 0.163891f
C8858 DVDD.n3103 VSS 0.198722f
C8859 DVDD.n3104 VSS 0.081946f
C8860 DVDD.n3105 VSS 0.098809f
C8861 DVDD.t147 VSS 0.167631f
C8862 DVDD.t114 VSS 0.167631f
C8863 DVDD.n3106 VSS 0.335261f
C8864 DVDD.n3107 VSS 0.281523f
C8865 DVDD.n3109 VSS 0.137328f
C8866 DVDD.n3110 VSS 0.137328f
C8867 DVDD.n3111 VSS 0.137328f
C8868 DVDD.n3112 VSS 0.121855f
C8869 DVDD.n3113 VSS 0.137328f
C8870 DVDD.n3114 VSS 0.137328f
C8871 DVDD.n3115 VSS 0.137328f
C8872 DVDD.n3116 VSS 0.137328f
C8873 DVDD.n3117 VSS 0.137328f
C8874 DVDD.n3118 VSS 0.135394f
C8875 DVDD.n3119 VSS 0.137328f
C8876 DVDD.n3120 VSS 0.137328f
C8877 DVDD.n3121 VSS 0.137328f
C8878 DVDD.n3122 VSS 0.13346f
C8879 DVDD.n3123 VSS 0.11992f
C8880 DVDD.n3124 VSS 0.112345f
C8881 DVDD.n3125 VSS 0.163891f
C8882 DVDD.n3126 VSS 0.128205f
C8883 DVDD.n3127 VSS 0.163891f
C8884 DVDD.n3128 VSS 0.122918f
C8885 DVDD.n3129 VSS 0.163891f
C8886 DVDD.n3130 VSS 0.128205f
C8887 DVDD.n3132 VSS 0.163891f
C8888 DVDD.n3133 VSS 0.163891f
C8889 DVDD.n3134 VSS 0.138779f
C8890 DVDD.n3136 VSS 0.183717f
C8891 DVDD.n3137 VSS 0.274656f
C8892 DVDD.n3138 VSS 0.274656f
C8893 DVDD.n3139 VSS 0.274656f
C8894 DVDD.n3140 VSS 0.274656f
C8895 DVDD.n3141 VSS 0.274656f
C8896 DVDD.n3142 VSS 0.274656f
C8897 DVDD.n3143 VSS 0.274656f
C8898 DVDD.n3144 VSS 0.274656f
C8899 DVDD.n3145 VSS 0.274656f
C8900 DVDD.n3146 VSS 0.176012f
C8901 DVDD.n3147 VSS 0.330748f
C8902 DVDD.n3148 VSS 0.497089f
C8903 DVDD.n3149 VSS 0.048355f
C8904 DVDD.n3150 VSS 0.163891f
C8905 DVDD.n3151 VSS 0.107058f
C8906 DVDD.n3152 VSS 0.163891f
C8907 DVDD.n3153 VSS 0.163891f
C8908 DVDD.n3154 VSS 0.163891f
C8909 DVDD.n3155 VSS 0.107058f
C8910 DVDD.n3156 VSS 0.163891f
C8911 DVDD.n3157 VSS 0.112345f
C8912 DVDD.n3158 VSS 0.163891f
C8913 DVDD.n3159 VSS 0.117632f
C8914 DVDD.n3160 VSS 0.163891f
C8915 DVDD.n3161 VSS 0.270949f
C8916 DVDD.n3162 VSS 0.11992f
C8917 DVDD.n3163 VSS 0.122918f
C8918 DVDD.n3164 VSS 0.163891f
C8919 DVDD.n3165 VSS 0.128205f
C8920 DVDD.n3166 VSS 0.163891f
C8921 DVDD.n3167 VSS 0.133492f
C8922 DVDD.n3168 VSS 0.163891f
C8923 DVDD.n3169 VSS 0.138779f
C8924 DVDD.n3170 VSS 0.163891f
C8925 DVDD.n3171 VSS 0.163891f
C8926 DVDD.n3172 VSS 0.163891f
C8927 DVDD.n3173 VSS 0.138779f
C8928 DVDD.n3174 VSS 0.229976f
C8929 DVDD.n3186 VSS 0.137328f
C8930 DVDD.n3188 VSS 0.137328f
C8931 DVDD.n3189 VSS 0.137328f
C8932 DVDD.n3190 VSS 0.137328f
C8933 DVDD.n3191 VSS 0.129591f
C8934 DVDD.n3192 VSS 0.137328f
C8935 DVDD.n3193 VSS 0.137328f
C8936 DVDD.n3194 VSS 0.137328f
C8937 DVDD.n3196 VSS 0.127657f
C8938 DVDD.n3197 VSS 0.137328f
C8939 DVDD.n3198 VSS 0.137328f
C8940 DVDD.n3199 VSS 0.125723f
C8941 DVDD.n3200 VSS 0.137328f
C8942 DVDD.n3201 VSS 0.11992f
C8943 DVDD.n3202 VSS 0.274656f
C8944 DVDD.n3203 VSS 0.274656f
C8945 DVDD.n3204 VSS 0.274656f
C8946 DVDD.n3205 VSS 0.11992f
C8947 DVDD.n3206 VSS 0.274656f
C8948 DVDD.n3207 VSS 0.274656f
C8949 DVDD.n3208 VSS 0.235972f
C8950 DVDD.n3209 VSS 0.274656f
C8951 DVDD.n3210 VSS 0.274656f
C8952 DVDD.n3211 VSS 0.274656f
C8953 DVDD.n3212 VSS 0.274656f
C8954 DVDD.n3213 VSS 0.274656f
C8955 DVDD.n3214 VSS 0.274656f
C8956 DVDD.n3215 VSS 0.11992f
C8957 DVDD.n3216 VSS 0.274656f
C8958 DVDD.n3217 VSS 0.11992f
C8959 DVDD.n3218 VSS 0.274656f
C8960 DVDD.n3219 VSS 0.11992f
C8961 DVDD.n3220 VSS 0.274656f
C8962 DVDD.n3221 VSS 0.11992f
C8963 DVDD.n3222 VSS 0.274656f
C8964 DVDD.n3223 VSS 0.11992f
C8965 DVDD.n3224 VSS 0.235972f
C8966 DVDD.n3225 VSS 0.235972f
C8967 DVDD.n3226 VSS 0.330748f
C8968 DVDD.n3227 VSS 0.524168f
C8969 DVDD.n3228 VSS 0.274656f
C8970 DVDD.n3229 VSS 0.11992f
C8971 DVDD.n3230 VSS 0.274656f
C8972 DVDD.n3231 VSS 0.330748f
C8973 DVDD.n3232 VSS 0.176012f
C8974 DVDD.n3233 VSS 0.235972f
C8975 DVDD.n3234 VSS 0.274656f
C8976 DVDD.n3235 VSS 0.098644f
C8977 DVDD.n3236 VSS 0.085911f
C8978 DVDD.n3237 VSS 0.163891f
C8979 DVDD.n3238 VSS 0.091198f
C8980 DVDD.n3239 VSS 0.163891f
C8981 DVDD.n3240 VSS 0.096484f
C8982 DVDD.n3241 VSS 0.163891f
C8983 DVDD.n3242 VSS 0.101771f
C8984 DVDD.n3243 VSS 0.163891f
C8985 DVDD.n3244 VSS 0.107058f
C8986 DVDD.n3245 VSS 0.163891f
C8987 DVDD.n3246 VSS 0.112345f
C8988 DVDD.n3247 VSS 0.210151f
C8989 DVDD.n3248 VSS 0.11992f
C8990 DVDD.n3249 VSS 0.163891f
C8991 DVDD.n3250 VSS 0.133492f
C8992 DVDD.n3251 VSS 0.163891f
C8993 DVDD.n3252 VSS 0.138779f
C8994 DVDD.n3253 VSS 0.163891f
C8995 DVDD.n3254 VSS 0.144066f
C8996 DVDD.n3255 VSS 0.163891f
C8997 DVDD.n3256 VSS 0.149352f
C8998 DVDD.n3257 VSS 0.163891f
C8999 DVDD.n3258 VSS 0.154639f
C9000 DVDD.n3259 VSS 0.163891f
C9001 DVDD.n3260 VSS 0.244515f
C9002 DVDD.n3272 VSS 0.137328f
C9003 DVDD.n3279 VSS 0.131525f
C9004 DVDD.n3280 VSS 0.137328f
C9005 DVDD.n3281 VSS 0.137328f
C9006 DVDD.n3282 VSS 0.048355f
C9007 DVDD.n3283 VSS 0.129591f
C9008 DVDD.n3284 VSS 0.137328f
C9009 DVDD.n3285 VSS 0.137328f
C9010 DVDD.n3286 VSS 0.081946f
C9011 DVDD.n3287 VSS 0.137328f
C9012 DVDD.n3289 VSS 0.127657f
C9013 DVDD.n3290 VSS 0.137328f
C9014 DVDD.n3291 VSS 0.137328f
C9015 DVDD.n3293 VSS 0.125723f
C9016 DVDD.n3294 VSS 0.137328f
C9017 DVDD.n3295 VSS 0.11992f
C9018 DVDD.n3296 VSS 0.274656f
C9019 DVDD.n3297 VSS 0.274656f
C9020 DVDD.n3298 VSS 0.274656f
C9021 DVDD.n3299 VSS 0.11992f
C9022 DVDD.n3300 VSS 0.274656f
C9023 DVDD.n3301 VSS 0.274656f
C9024 DVDD.n3302 VSS 0.274656f
C9025 DVDD.n3303 VSS 0.11992f
C9026 DVDD.n3304 VSS 0.274656f
C9027 DVDD.n3305 VSS 0.11992f
C9028 DVDD.n3306 VSS 0.274656f
C9029 DVDD.n3307 VSS 0.274656f
C9030 DVDD.n3308 VSS 0.274656f
C9031 DVDD.n3309 VSS 0.274656f
C9032 DVDD.n3310 VSS 0.11992f
C9033 DVDD.n3311 VSS 0.274656f
C9034 DVDD.n3312 VSS 0.11992f
C9035 DVDD.n3313 VSS 0.274656f
C9036 DVDD.n3314 VSS 0.11992f
C9037 DVDD.n3315 VSS 0.274656f
C9038 DVDD.n3316 VSS 0.274656f
C9039 DVDD.n3317 VSS 0.274656f
C9040 DVDD.n3318 VSS 0.274656f
C9041 DVDD.n3319 VSS 0.274656f
C9042 DVDD.n3320 VSS 0.274656f
C9043 DVDD.n3321 VSS 0.274656f
C9044 DVDD.n3322 VSS 0.205025f
C9045 DVDD.n3323 VSS 0.274656f
C9046 DVDD.n3324 VSS 0.274656f
C9047 DVDD.n3325 VSS 0.274656f
C9048 DVDD.n3326 VSS 0.274656f
C9049 DVDD.n3327 VSS 0.274656f
C9050 DVDD.n3328 VSS 0.274656f
C9051 DVDD.n3329 VSS 0.274656f
C9052 DVDD.n3330 VSS 0.274656f
C9053 DVDD.n3331 VSS 0.274656f
C9054 DVDD.n3332 VSS 0.274656f
C9055 DVDD.n3333 VSS 0.274656f
C9056 DVDD.n3334 VSS 0.11992f
C9057 DVDD.n3335 VSS 0.274656f
C9058 DVDD.n3336 VSS 0.274656f
C9059 DVDD.n3337 VSS 0.11992f
C9060 DVDD.n3338 VSS 0.274656f
C9061 DVDD.n3339 VSS 0.274656f
C9062 DVDD.n3340 VSS 0.274656f
C9063 DVDD.n3341 VSS 0.274656f
C9064 DVDD.n3342 VSS 0.274656f
C9065 DVDD.n3343 VSS 0.274656f
C9066 DVDD.n3344 VSS 0.274656f
C9067 DVDD.n3345 VSS 0.274656f
C9068 DVDD.n3346 VSS 0.274656f
C9069 DVDD.n3347 VSS 0.11992f
C9070 DVDD.n3348 VSS 0.071372f
C9071 DVDD.n3349 VSS 1.37325f
C9072 DVDD.n3350 VSS 0.163891f
C9073 DVDD.n3351 VSS 0.153317f
C9074 DVDD.n3352 VSS 0.163891f
C9075 DVDD.n3353 VSS 0.163891f
C9076 DVDD.n3354 VSS 0.163891f
C9077 DVDD.n3355 VSS 0.085911f
C9078 DVDD.n3356 VSS 0.163891f
C9079 DVDD.n3357 VSS 0.091198f
C9080 DVDD.n3358 VSS 0.163891f
C9081 DVDD.n3359 VSS 0.149352f
C9082 DVDD.n3360 VSS 0.163891f
C9083 DVDD.n3361 VSS 0.154639f
C9084 DVDD.n3362 VSS 0.163891f
C9085 DVDD.n3363 VSS 0.159926f
C9086 DVDD.n3364 VSS 0.163891f
C9087 DVDD.n3365 VSS 0.163891f
C9088 DVDD.n3366 VSS 0.163891f
C9089 DVDD.n3367 VSS 0.163891f
C9090 DVDD.n3368 VSS 0.163891f
C9091 DVDD.n3369 VSS 0.113666f
C9092 DVDD.n3370 VSS 0.081946f
C9093 DVDD.n3381 VSS 0.137328f
C9094 DVDD.n3389 VSS 0.131525f
C9095 DVDD.n3390 VSS 0.137328f
C9096 DVDD.n3391 VSS 0.137328f
C9097 DVDD.n3392 VSS 0.137328f
C9098 DVDD.n3393 VSS 0.129591f
C9099 DVDD.n3394 VSS 0.137328f
C9100 DVDD.n3395 VSS 0.137328f
C9101 DVDD.n3396 VSS 0.081946f
C9102 DVDD.n3397 VSS 0.137328f
C9103 DVDD.n3399 VSS 0.127657f
C9104 DVDD.n3400 VSS 0.098644f
C9105 DVDD.n3401 VSS 0.137328f
C9106 DVDD.n3402 VSS 0.137328f
C9107 DVDD.n3404 VSS 0.125723f
C9108 DVDD.n3405 VSS 0.11992f
C9109 DVDD.n3406 VSS 0.274656f
C9110 DVDD.n3407 VSS 0.274656f
C9111 DVDD.n3408 VSS 0.11992f
C9112 DVDD.n3409 VSS 0.274656f
C9113 DVDD.n3410 VSS 0.274656f
C9114 DVDD.n3411 VSS 0.11992f
C9115 DVDD.n3412 VSS 0.274656f
C9116 DVDD.n3413 VSS 0.274656f
C9117 DVDD.n3414 VSS 0.274656f
C9118 DVDD.n3415 VSS 0.158604f
C9119 DVDD.n3416 VSS 0.274656f
C9120 DVDD.n3417 VSS 0.274656f
C9121 DVDD.n3418 VSS 0.274656f
C9122 DVDD.n3419 VSS 0.123789f
C9123 DVDD.n3420 VSS 0.071372f
C9124 DVDD.n3421 VSS 1.37325f
C9125 DVDD.n3422 VSS 0.163891f
C9126 DVDD.n3423 VSS 0.153317f
C9127 DVDD.n3424 VSS 0.163891f
C9128 DVDD.n3425 VSS 0.163891f
C9129 DVDD.n3426 VSS 0.163891f
C9130 DVDD.n3427 VSS 0.085911f
C9131 DVDD.n3428 VSS 0.163891f
C9132 DVDD.n3429 VSS 0.091198f
C9133 DVDD.n3430 VSS 0.163891f
C9134 DVDD.n3431 VSS 0.244515f
C9135 DVDD.n3433 VSS 0.198722f
C9136 DVDD.n3434 VSS 0.081946f
C9137 DVDD.n3435 VSS 0.098809f
C9138 DVDD.t117 VSS 0.167631f
C9139 DVDD.t76 VSS 0.167631f
C9140 DVDD.n3436 VSS 0.335261f
C9141 DVDD.n3437 VSS 0.081946f
C9142 DVDD.n3438 VSS 0.099098f
C9143 DVDD.n3439 VSS 0.198298f
C9144 DVDD.n3440 VSS 0.149352f
C9145 DVDD.n3442 VSS 0.163891f
C9146 DVDD.n3444 VSS 0.198722f
C9147 DVDD.n3445 VSS 0.081946f
C9148 DVDD.n3446 VSS 0.098809f
C9149 DVDD.t107 VSS 0.167631f
C9150 DVDD.t133 VSS 0.167631f
C9151 DVDD.n3447 VSS 0.335261f
C9152 DVDD.n3448 VSS 0.081946f
C9153 DVDD.n3449 VSS 0.099098f
C9154 DVDD.n3450 VSS 0.198298f
C9155 DVDD.n3451 VSS 0.154639f
C9156 DVDD.n3453 VSS 0.163891f
C9157 DVDD.n3455 VSS 0.198722f
C9158 DVDD.n3456 VSS 0.081946f
C9159 DVDD.n3457 VSS 0.098809f
C9160 DVDD.t122 VSS 0.425324f
C9161 DVDD.n3458 VSS 0.081946f
C9162 DVDD.n3459 VSS 0.099098f
C9163 DVDD.n3460 VSS 0.198298f
C9164 DVDD.n3461 VSS 0.159926f
C9165 DVDD.n3463 VSS 0.163891f
C9166 DVDD.n3465 VSS 0.163891f
C9167 DVDD.n3467 VSS 0.163891f
C9168 DVDD.n3469 VSS 0.163891f
C9169 DVDD.n3471 VSS 0.163891f
C9170 DVDD.n3472 VSS 0.113666f
C9171 DVDD.n3473 VSS 0.081946f
C9172 DVDD.n3481 VSS 0.137328f
C9173 DVDD.n3482 VSS 0.137328f
C9174 DVDD.n3483 VSS 0.137328f
C9175 DVDD.n3484 VSS 0.121855f
C9176 DVDD.n3485 VSS 0.137328f
C9177 DVDD.n3486 VSS 0.137328f
C9178 DVDD.n3487 VSS 0.137328f
C9179 DVDD.n3488 VSS 0.081946f
C9180 DVDD.n3489 VSS 0.137328f
C9181 DVDD.n3490 VSS 0.137328f
C9182 DVDD.n3492 VSS 0.135394f
C9183 DVDD.n3493 VSS 0.137328f
C9184 DVDD.n3494 VSS 0.137328f
C9185 DVDD.n3495 VSS 0.11992f
C9186 DVDD.n3496 VSS 0.274656f
C9187 DVDD.n3497 VSS 0.274656f
C9188 DVDD.n3498 VSS 0.11992f
C9189 DVDD.n3499 VSS 0.274656f
C9190 DVDD.n3500 VSS 0.274656f
C9191 DVDD.n3501 VSS 0.11992f
C9192 DVDD.n3502 VSS 0.274656f
C9193 DVDD.n3503 VSS 0.274656f
C9194 DVDD.n3504 VSS 0.274656f
C9195 DVDD.n3505 VSS 0.330748f
C9196 DVDD.n3506 VSS 0.330748f
C9197 DVDD.n3507 VSS 0.524168f
C9198 DVDD.n3508 VSS 0.274656f
C9199 DVDD.n3509 VSS 0.274656f
C9200 DVDD.n3510 VSS 0.11992f
C9201 DVDD.n3511 VSS 0.06615f
C9202 DVDD.n3512 VSS 0.06615f
C9203 DVDD.n3513 VSS 0.06615f
C9204 DVDD.n3514 VSS 0.06615f
C9205 DVDD.n3515 VSS 0.06615f
C9206 DVDD.n3516 VSS 0.06615f
C9207 DVDD.n3517 VSS 0.06615f
C9208 DVDD.n3518 VSS 0.06615f
C9209 DVDD.n3519 VSS 0.0147f
C9210 DVDD.n3520 VSS 0.090649f
C9211 DVDD.n3521 VSS 0.151899f
C9212 DVDD.n3523 VSS 0.073242f
C9213 DVDD.n3524 VSS 0.067568f
C9214 DVDD.n3525 VSS 0.073242f
C9215 DVDD.n3526 VSS 0.073242f
C9216 DVDD.n3527 VSS 0.073242f
C9217 DVDD.n3528 VSS 0.073242f
C9218 DVDD.n3529 VSS 0.069631f
C9219 DVDD.n3530 VSS 0.073242f
C9220 DVDD.n3531 VSS 0.073242f
C9221 DVDD.n3532 VSS 0.034496f
C9222 DVDD.n3533 VSS 0.079009f
C9223 DVDD.n3534 VSS 0.079009f
C9224 DVDD.n3535 VSS 0.079009f
C9225 DVDD.n3536 VSS 0.039504f
C9226 DVDD.n3537 VSS 0.035888f
C9227 DVDD.n3538 VSS 0.073242f
C9228 DVDD.n3540 VSS 0.056009f
C9229 DVDD.n3541 VSS 0.056009f
C9230 DVDD.n3542 VSS 0.089747f
C9231 DVDD.n3543 VSS 0.079009f
C9232 DVDD.n3544 VSS 0.079009f
C9233 DVDD.n3545 VSS 0.034496f
C9234 DVDD.n3547 VSS 0.039504f
C9235 DVDD.n3548 VSS 0.079009f
C9236 DVDD.n3549 VSS 0.034496f
C9237 DVDD.n3550 VSS 0.035331f
C9238 DVDD.n3552 VSS 0.137328f
C9239 DVDD.n3553 VSS 0.137328f
C9240 DVDD.n3554 VSS 0.137328f
C9241 DVDD.n3555 VSS 0.12669f
C9242 DVDD.n3556 VSS 0.137328f
C9243 DVDD.n3557 VSS 0.137328f
C9244 DVDD.n3558 VSS 0.137328f
C9245 DVDD.n3559 VSS 0.137328f
C9246 DVDD.n3560 VSS 0.130558f
C9247 DVDD.n3561 VSS 0.137328f
C9248 DVDD.n3562 VSS 0.137328f
C9249 DVDD.n3563 VSS 0.137328f
C9250 DVDD.n3564 VSS 0.128624f
C9251 DVDD.n3565 VSS 0.526097f
C9252 DVDD.n3566 VSS 0.151899f
C9253 DVDD.n3567 VSS 0.151899f
C9254 DVDD.n3568 VSS 0.151899f
C9255 DVDD.n3569 VSS 0.151899f
C9256 DVDD.n3570 VSS 0.151899f
C9257 DVDD.n3571 VSS 0.151899f
C9258 DVDD.n3572 VSS 0.151899f
C9259 DVDD.n3573 VSS 0.151899f
C9260 DVDD.n3574 VSS 0.151899f
C9261 DVDD.n3575 VSS 0.151899f
C9262 DVDD.n3576 VSS 0.151899f
C9263 DVDD.n3578 VSS 3.23275f
C9264 DVDD.n3579 VSS 0.11992f
C9265 DVDD.n3580 VSS 0.11992f
C9266 DVDD.n3581 VSS 0.274656f
C9267 DVDD.n3582 VSS 0.274656f
C9268 DVDD.n3583 VSS 0.11992f
C9269 DVDD.n3584 VSS 0.11992f
C9270 DVDD.n3585 VSS 0.11992f
C9271 DVDD.n3586 VSS 0.11992f
C9272 DVDD.n3587 VSS 0.274656f
C9273 DVDD.n3588 VSS 0.274656f
C9274 DVDD.n3589 VSS 0.11992f
C9275 DVDD.n3590 VSS 0.11992f
C9276 DVDD.n3591 VSS 0.11992f
C9277 DVDD.n3592 VSS 0.11992f
C9278 DVDD.n3593 VSS 0.274656f
C9279 DVDD.n3594 VSS 0.274656f
C9280 DVDD.n3595 VSS 0.11992f
C9281 DVDD.n3596 VSS 0.217597f
C9282 DVDD.n3597 VSS 0.183749f
C9283 DVDD.n3598 VSS 0.21057f
C9284 DVDD.n3599 VSS 0.228235f
C9285 DVDD.n3600 VSS 0.097999f
C9286 DVDD.n3601 VSS 0.146483f
C9287 DVDD.n3602 VSS 0.146483f
C9288 DVDD.n3603 VSS 0.116052f
C9289 DVDD.n3604 VSS 0.063957f
C9290 DVDD.n3605 VSS 0.146483f
C9291 DVDD.n3606 VSS 0.146483f
C9292 DVDD.n3607 VSS 0.063957f
C9293 DVDD.n3608 VSS 0.146483f
C9294 DVDD.n3609 VSS 0.063957f
C9295 DVDD.n3610 VSS 0.146483f
C9296 DVDD.n3611 VSS 0.057252f
C9297 DVDD.n3612 VSS 0.089747f
C9298 DVDD.n3613 VSS 0.063957f
C9299 DVDD.n3614 VSS 0.146483f
C9300 DVDD.n3615 VSS 0.146483f
C9301 DVDD.n3616 VSS 0.063957f
C9302 DVDD.n3617 VSS 0.146483f
C9303 DVDD.n3618 VSS 0.063957f
C9304 DVDD.n3619 VSS 0.146483f
C9305 DVDD.n3620 VSS 0.146483f
C9306 DVDD.n3621 VSS 0.146483f
C9307 DVDD.n3622 VSS 0.146483f
C9308 DVDD.n3623 VSS 0.146483f
C9309 DVDD.n3624 VSS 0.063957f
C9310 DVDD.n3625 VSS 0.146483f
C9311 DVDD.n3626 VSS 0.063957f
C9312 DVDD.n3627 VSS 0.146483f
C9313 DVDD.n3628 VSS 0.146483f
C9314 DVDD.n3629 VSS 0.146483f
C9315 DVDD.n3630 VSS 0.146483f
C9316 DVDD.n3631 VSS 0.146483f
C9317 DVDD.n3632 VSS 0.097999f
C9318 DVDD.n3633 VSS 0.097999f
C9319 DVDD.n3634 VSS 0.21057f
C9320 DVDD.n3635 VSS 0.073242f
C9321 DVDD.n3636 VSS 0.146483f
C9322 DVDD.n3637 VSS 0.146483f
C9323 DVDD.n3638 VSS 0.146483f
C9324 DVDD.n3639 VSS 0.063957f
C9325 DVDD.n3640 VSS 0.073242f
C9326 DVDD.n3641 VSS 0.163891f
C9327 DVDD.n3642 VSS 0.163891f
C9328 DVDD.n3643 VSS 0.130849f
C9329 DVDD.n3644 VSS 0.163891f
C9330 DVDD.n3645 VSS 0.163891f
C9331 DVDD.n3646 VSS 0.063957f
C9332 DVDD.n3647 VSS 1.37325f
C9333 DVDD.n3648 VSS 0.315887f
C9334 DVDD.n3649 VSS 0.163891f
C9335 DVDD.n3650 VSS 0.114988f
C9336 DVDD.n3651 VSS 0.163891f
C9337 DVDD.n3652 VSS 0.073242f
C9338 DVDD.n3653 VSS 0.07221f
C9339 DVDD.n3654 VSS 0.073242f
C9340 DVDD.n3655 VSS 0.017666f
C9341 DVDD.n3656 VSS 0.071178f
C9342 DVDD.n3663 VSS 0.066021f
C9343 DVDD.n3665 VSS 0.066021f
C9344 DVDD.n3667 VSS 0.064989f
C9345 DVDD.n3668 VSS 0.063957f
C9346 DVDD.n3669 VSS 0.146483f
C9347 DVDD.n3670 VSS 0.063957f
C9348 DVDD.n3671 VSS 0.146483f
C9349 DVDD.n3672 VSS 0.146483f
C9350 DVDD.n3673 VSS 0.104963f
C9351 DVDD.n3674 VSS 0.02695f
C9352 DVDD.n3675 VSS 0.027981f
C9353 DVDD.n3676 VSS 0.146483f
C9354 DVDD.n3678 VSS 0.01831f
C9355 DVDD.n3679 VSS 0.036621f
C9356 DVDD.n3680 VSS 0.036964f
C9357 DVDD.n3681 VSS 0.016376f
C9358 DVDD.n3682 VSS 0.015989f
C9359 DVDD.n3683 VSS 0.01831f
C9360 DVDD.n3684 VSS 0.015989f
C9361 DVDD.n3685 VSS 0.036621f
C9362 DVDD.n3686 VSS 0.037194f
C9363 DVDD.n3687 VSS 0.105852f
C9364 DVDD.n3688 VSS 0.02695f
C9365 DVDD.n3689 VSS 0.036621f
C9366 DVDD.n3690 VSS 0.036621f
C9367 DVDD.n3691 VSS 0.015989f
C9368 DVDD.n3692 VSS 0.01831f
C9369 DVDD.n3693 VSS 0.015989f
C9370 DVDD.n3694 VSS 0.01831f
C9371 DVDD.n3695 VSS 0.015989f
C9372 DVDD.n3696 VSS 0.036621f
C9373 DVDD.n3697 VSS 0.027981f
C9374 DVDD.n3698 VSS 0.036277f
C9375 DVDD.n3699 VSS 0.016634f
C9376 DVDD.n3700 VSS 0.015989f
C9377 DVDD.n3701 VSS 0.036621f
C9378 DVDD.n3702 VSS 0.035087f
C9379 DVDD.n3703 VSS 0.103874f
C9380 DVDD.n3704 VSS 0.036621f
C9381 DVDD.n3705 VSS 0.036621f
C9382 DVDD.n3706 VSS 0.015989f
C9383 DVDD.n3707 VSS 0.01831f
C9384 DVDD.n3708 VSS 0.015989f
C9385 DVDD.n3709 VSS 0.051321f
C9386 DVDD.n3711 VSS 0.063957f
C9387 DVDD.n3712 VSS 0.073242f
C9388 DVDD.n3713 VSS 0.037137f
C9389 DVDD.n3714 VSS 0.146483f
C9390 DVDD.n3715 VSS 0.146483f
C9391 DVDD.n3718 VSS 0.146483f
C9392 DVDD.n3719 VSS 0.146483f
C9393 DVDD.n3720 VSS 0.146483f
C9394 DVDD.n3721 VSS 0.146483f
C9395 DVDD.n3722 VSS 0.163891f
C9396 DVDD.n3723 VSS 0.163891f
C9397 DVDD.n3724 VSS 0.130849f
C9398 DVDD.n3725 VSS 0.163891f
C9399 DVDD.n3726 VSS 0.163891f
C9400 DVDD.n3727 VSS 0.063957f
C9401 DVDD.n3728 VSS 1.37325f
C9402 DVDD.n3729 VSS 0.315887f
C9403 DVDD.n3730 VSS 0.163891f
C9404 DVDD.n3731 VSS 0.114988f
C9405 DVDD.n3732 VSS 0.163891f
C9406 DVDD.n3733 VSS 0.073242f
C9407 DVDD.n3734 VSS 0.068084f
C9408 DVDD.n3735 VSS 0.05261f
C9409 DVDD.n3736 VSS 0.073242f
C9410 DVDD.n3737 VSS 0.073242f
C9411 DVDD.n3738 VSS 0.067052f
C9412 DVDD.n3739 VSS 0.073242f
C9413 DVDD.n3746 VSS 0.073242f
C9414 DVDD.n3748 VSS 0.073242f
C9415 DVDD.n3749 VSS 0.073242f
C9416 DVDD.n3750 VSS 0.073242f
C9417 DVDD.n3752 VSS 0.069115f
C9418 DVDD.n3753 VSS 0.063957f
C9419 DVDD.n3754 VSS 0.146483f
C9420 DVDD.n3755 VSS 0.093873f
C9421 DVDD.n3756 VSS 0.146483f
C9422 DVDD.n3757 VSS 0.125852f
C9423 DVDD.n3758 VSS 0.176012f
C9424 DVDD.n3759 VSS 0.274656f
C9425 DVDD.n3760 VSS 0.21057f
C9426 DVDD.n3761 VSS 0.11992f
C9427 DVDD.n3762 VSS 0.11992f
C9428 DVDD.n3763 VSS 0.11992f
C9429 DVDD.n3764 VSS 0.274656f
C9430 DVDD.n3765 VSS 0.274656f
C9431 DVDD.n3766 VSS 0.11992f
C9432 DVDD.n3767 VSS 0.11992f
C9433 DVDD.n3768 VSS 0.11992f
C9434 DVDD.n3769 VSS 0.274656f
C9435 DVDD.n3770 VSS 0.274656f
C9436 DVDD.n3771 VSS 0.11992f
C9437 DVDD.n3772 VSS 0.163891f
C9438 DVDD.n3773 VSS 0.163891f
C9439 DVDD.n3774 VSS 0.163891f
C9440 DVDD.n3775 VSS 0.163891f
C9441 DVDD.n3776 VSS 0.163891f
C9442 DVDD.n3777 VSS 0.163891f
C9443 DVDD.n3778 VSS 0.163891f
C9444 DVDD.n3779 VSS 0.163891f
C9445 DVDD.n3780 VSS 0.163891f
C9446 DVDD.n3781 VSS 0.163891f
C9447 DVDD.n3782 VSS 0.163891f
C9448 DVDD.n3783 VSS 0.315887f
C9449 DVDD.n3784 VSS 0.163891f
C9450 DVDD.n3785 VSS 0.163891f
C9451 DVDD.n3786 VSS 0.163891f
C9452 DVDD.n3787 VSS 0.163891f
C9453 DVDD.n3788 VSS 0.163891f
C9454 DVDD.n3789 VSS 0.163891f
C9455 DVDD.n3790 VSS 0.163891f
C9456 DVDD.n3791 VSS 0.163891f
C9457 DVDD.n3792 VSS 0.163891f
C9458 DVDD.n3793 VSS 0.163891f
C9459 DVDD.n3794 VSS 0.163891f
C9460 DVDD.n3807 VSS 0.131525f
C9461 DVDD.n3808 VSS 0.137328f
C9462 DVDD.n3809 VSS 0.137328f
C9463 DVDD.n3810 VSS 0.137328f
C9464 DVDD.n3811 VSS 0.129591f
C9465 DVDD.n3812 VSS 0.137328f
C9466 DVDD.n3813 VSS 0.137328f
C9467 DVDD.n3814 VSS 0.137328f
C9468 DVDD.n3816 VSS 0.127657f
C9469 DVDD.n3817 VSS 0.025789f
C9470 DVDD.n3818 VSS 0.11992f
C9471 DVDD.n3819 VSS 0.274656f
C9472 DVDD.n3820 VSS 0.11992f
C9473 DVDD.n3821 VSS 0.274656f
C9474 DVDD.n3822 VSS 0.274656f
C9475 DVDD.n3823 VSS 0.158604f
C9476 DVDD.n3824 VSS 0.274656f
C9477 DVDD.n3825 VSS 0.274656f
C9478 DVDD.n3826 VSS 0.274656f
C9479 DVDD.n3827 VSS 0.123789f
C9480 DVDD.n3828 VSS 0.163891f
C9481 DVDD.n3829 VSS 0.163891f
C9482 DVDD.n3830 VSS 0.163891f
C9483 DVDD.n3831 VSS 0.163891f
C9484 DVDD.n3832 VSS 0.163891f
C9485 DVDD.n3833 VSS 0.163891f
C9486 DVDD.n3834 VSS 0.163891f
C9487 DVDD.n3835 VSS 0.163891f
C9488 DVDD.n3836 VSS 0.163891f
C9489 DVDD.n3837 VSS 0.163891f
C9490 DVDD.n3838 VSS 0.163891f
C9491 DVDD.n3839 VSS 0.315887f
C9492 DVDD.n3841 VSS 0.163891f
C9493 DVDD.n3843 VSS 0.163891f
C9494 DVDD.n3845 VSS 0.163891f
C9495 DVDD.n3847 VSS 0.163891f
C9496 DVDD.n3849 VSS 0.163891f
C9497 DVDD.n3851 VSS 0.163891f
C9498 DVDD.n3853 VSS 0.163891f
C9499 DVDD.n3855 VSS 0.163891f
C9500 DVDD.n3857 VSS 0.163891f
C9501 DVDD.n3859 VSS 0.163891f
C9502 DVDD.n3861 VSS 0.163891f
C9503 DVDD.n3863 VSS 0.064086f
C9504 DVDD.n3864 VSS 0.064086f
C9505 DVDD.n3865 VSS 0.064086f
C9506 DVDD.n3867 VSS 0.064086f
C9507 DVDD.n3868 VSS 0.064086f
C9508 DVDD.n3869 VSS 0.064086f
C9509 DVDD.n3870 VSS 0.064086f
C9510 DVDD.n3871 VSS 0.064086f
C9511 DVDD.n3872 VSS 0.064086f
C9512 DVDD.n3873 VSS 0.064086f
C9513 DVDD.n3874 VSS 0.064086f
C9514 DVDD.n3875 VSS 0.062281f
C9515 DVDD.n3876 VSS 0.055963f
C9516 DVDD.n3878 VSS 0.163891f
C9517 DVDD.n3879 VSS 0.163891f
C9518 DVDD.n3880 VSS 0.163891f
C9519 DVDD.n3881 VSS 0.163891f
C9520 DVDD.n3882 VSS 0.163891f
C9521 DVDD.n3883 VSS 0.074015f
C9522 DVDD.n3885 VSS 0.163891f
C9523 DVDD.n3887 VSS 0.163891f
C9524 DVDD.n3889 VSS 0.163891f
C9525 DVDD.n3894 VSS 0.057768f
C9526 DVDD.n3897 VSS 0.056865f
C9527 DVDD.n3898 VSS 0.055963f
C9528 DVDD.n3899 VSS 0.128173f
C9529 DVDD.n3900 VSS 0.055963f
C9530 DVDD.n3901 VSS 0.128173f
C9531 DVDD.n3902 VSS 0.128173f
C9532 DVDD.n3903 VSS 0.128173f
C9533 DVDD.n3904 VSS 0.128173f
C9534 DVDD.n3905 VSS 0.128173f
C9535 DVDD.n3906 VSS 0.101545f
C9536 DVDD.n3907 VSS 0.128173f
C9537 DVDD.n3908 VSS 0.128173f
C9538 DVDD.n3909 VSS 0.128173f
C9539 DVDD.n3910 VSS 0.064086f
C9540 DVDD.n3911 VSS 0.151899f
C9541 DVDD.n3912 VSS 0.151899f
C9542 DVDD.n3913 VSS 0.151899f
C9543 DVDD.n3914 VSS 0.151899f
C9544 DVDD.n3915 VSS 0.151899f
C9545 DVDD.n3916 VSS 0.296448f
C9546 DVDD.n3917 VSS 0.151899f
C9547 DVDD.n3918 VSS 0.151899f
C9548 DVDD.n3919 VSS 0.151899f
C9549 DVDD.n3920 VSS 0.151899f
C9550 DVDD.n3922 VSS 0.064086f
C9551 DVDD.n3923 VSS 0.064086f
C9552 DVDD.n3924 VSS 0.059122f
C9553 DVDD.n3925 VSS 0.064086f
C9554 DVDD.n3926 VSS 0.055963f
C9555 DVDD.n3927 VSS 0.064086f
C9556 DVDD.n3929 VSS 0.060927f
C9557 DVDD.n3930 VSS 0.064086f
C9558 DVDD.n3931 VSS 0.064086f
C9559 DVDD.n3932 VSS 0.064086f
C9560 DVDD.n3934 VSS 0.353402f
C9561 DVDD.n3940 VSS 0.060025f
C9562 DVDD.n3941 VSS 0.128173f
C9563 DVDD.n3942 VSS 0.128173f
C9564 DVDD.n3943 VSS 0.055963f
C9565 DVDD.n3944 VSS 0.128173f
C9566 DVDD.n3945 VSS 0.128173f
C9567 DVDD.n3946 VSS 0.128173f
C9568 DVDD.n3947 VSS 0.055963f
C9569 DVDD.n3948 VSS 0.128173f
C9570 DVDD.n3949 VSS 0.055963f
C9571 DVDD.n3950 VSS 0.128173f
C9572 DVDD.n3951 VSS 0.055963f
C9573 DVDD.n3952 VSS 0.128173f
C9574 DVDD.n3953 VSS 0.128173f
C9575 DVDD.n3954 VSS 0.128173f
C9576 DVDD.n3955 VSS 0.128173f
C9577 DVDD.n3956 VSS 0.055963f
C9578 DVDD.n3957 VSS 0.128173f
C9579 DVDD.n3958 VSS 0.055963f
C9580 DVDD.n3959 VSS 0.128173f
C9581 DVDD.n3960 VSS 0.055963f
C9582 DVDD.n3961 VSS 0.128173f
C9583 DVDD.n3962 VSS 0.128173f
C9584 DVDD.n3963 VSS 0.128173f
C9585 DVDD.n3964 VSS 0.587849f
C9586 DVDD.n3965 VSS 0.060025f
C9587 DVDD.n3966 VSS 0.055963f
C9588 DVDD.n3971 VSS 0.064086f
C9589 DVDD.n3972 VSS 0.055963f
C9590 DVDD.n3973 VSS 0.128173f
C9591 DVDD.n3974 VSS 0.159414f
C9592 DVDD.n3975 VSS 0.055963f
C9593 DVDD.n3976 VSS 0.373774f
C9594 DVDD.n3977 VSS 3.23275f
C9595 DVDD.n3978 VSS 0.064086f
C9596 DVDD.n3979 VSS 0.055963f
C9597 DVDD.n3980 VSS 0.128173f
C9598 DVDD.n3981 VSS 0.128173f
C9599 DVDD.n3982 VSS 0.128173f
C9600 DVDD.n3983 VSS 0.128173f
C9601 DVDD.n3984 VSS 0.128173f
C9602 DVDD.n3985 VSS 0.128173f
C9603 DVDD.n3986 VSS 0.128173f
C9604 DVDD.n3987 VSS 0.111926f
C9605 DVDD.n3988 VSS 0.128173f
C9606 DVDD.n3989 VSS 0.128173f
C9607 DVDD.n3990 VSS 0.128173f
C9608 DVDD.n3991 VSS 0.128173f
C9609 DVDD.n3992 VSS 0.128173f
C9610 DVDD.n3993 VSS 0.055963f
C9611 DVDD.n3994 VSS 0.128173f
C9612 DVDD.n3995 VSS 0.055963f
C9613 DVDD.n3996 VSS 0.128173f
C9614 DVDD.n3997 VSS 0.055963f
C9615 DVDD.n3998 VSS 0.128173f
C9616 DVDD.n3999 VSS 0.128173f
C9617 DVDD.n4000 VSS 0.128173f
C9618 DVDD.n4001 VSS 0.128173f
C9619 DVDD.n4002 VSS 0.055963f
C9620 DVDD.n4003 VSS 0.128173f
C9621 DVDD.n4004 VSS 0.128173f
C9622 DVDD.n4005 VSS 0.128173f
C9623 DVDD.n4006 VSS 0.128173f
C9624 DVDD.n4007 VSS 0.128173f
C9625 DVDD.n4008 VSS 0.055963f
C9626 DVDD.n4009 VSS 0.128173f
C9627 DVDD.n4010 VSS 0.128173f
C9628 DVDD.n4011 VSS 0.055963f
C9629 DVDD.n4012 VSS 0.128173f
C9630 DVDD.n4013 VSS 0.128173f
C9631 DVDD.n4014 VSS 0.055963f
C9632 DVDD.n4015 VSS 0.128173f
C9633 DVDD.n4016 VSS 0.128173f
C9634 DVDD.n4017 VSS 0.128173f
C9635 DVDD.n4018 VSS 0.055963f
C9636 DVDD.n4019 VSS 0.128173f
C9637 DVDD.n4020 VSS 0.055963f
C9638 DVDD.n4021 VSS 0.128173f
C9639 DVDD.n4022 VSS 0.055963f
C9640 DVDD.n4023 VSS 0.128173f
C9641 DVDD.n4024 VSS 0.128173f
C9642 DVDD.n4025 VSS 0.128173f
C9643 DVDD.n4026 VSS 0.128173f
C9644 DVDD.n4027 VSS 0.055963f
C9645 DVDD.n4028 VSS 0.128173f
C9646 DVDD.n4029 VSS 0.055963f
C9647 DVDD.n4030 VSS 0.128173f
C9648 DVDD.n4031 VSS 0.055963f
C9649 DVDD.n4032 VSS 0.128173f
C9650 DVDD.n4033 VSS 0.128173f
C9651 DVDD.n4034 VSS 0.128173f
C9652 DVDD.n4035 VSS 0.128173f
C9653 DVDD.n4036 VSS 0.128173f
C9654 DVDD.n4037 VSS 0.092068f
C9655 DVDD.n4038 VSS 0.128173f
C9656 DVDD.n4039 VSS 0.128173f
C9657 DVDD.n4040 VSS 0.128173f
C9658 DVDD.n4041 VSS 0.128173f
C9659 DVDD.n4042 VSS 0.128173f
C9660 DVDD.n4043 VSS 0.128173f
C9661 DVDD.n4044 VSS 0.128173f
C9662 DVDD.n4045 VSS 0.055963f
C9663 DVDD.n4046 VSS 0.128173f
C9664 DVDD.n4047 VSS 0.055963f
C9665 DVDD.n4048 VSS 0.128173f
C9666 DVDD.n4049 VSS 0.128173f
C9667 DVDD.n4050 VSS 0.128173f
C9668 DVDD.n4051 VSS 0.128173f
C9669 DVDD.n4052 VSS 0.055963f
C9670 DVDD.n4053 VSS 0.128173f
C9671 DVDD.n4054 VSS 0.055963f
C9672 DVDD.n4055 VSS 0.128173f
C9673 DVDD.n4056 VSS 0.055963f
C9674 DVDD.n4057 VSS 0.128173f
C9675 DVDD.n4058 VSS 0.128173f
C9676 DVDD.n4059 VSS 0.128173f
C9677 DVDD.n4060 VSS 0.128173f
C9678 DVDD.n4061 VSS 0.128173f
C9679 DVDD.n4062 VSS 0.055963f
C9680 DVDD.n4063 VSS 0.063184f
C9681 DVDD.n4064 VSS 0.163891f
C9682 DVDD.n4065 VSS 0.064086f
C9683 DVDD.n4066 VSS 3.48797f
C9684 DVDD.n4079 VSS 0.137328f
C9685 DVDD.n4080 VSS 0.137328f
C9686 DVDD.n4081 VSS 0.137328f
C9687 DVDD.n4082 VSS 0.121855f
C9688 DVDD.n4083 VSS 0.137328f
C9689 DVDD.n4084 VSS 0.137328f
C9690 DVDD.n4085 VSS 0.137328f
C9691 DVDD.n4086 VSS 0.137328f
C9692 DVDD.n4087 VSS 0.137328f
C9693 DVDD.n4089 VSS 0.135394f
C9694 DVDD.n4090 VSS 0.137328f
C9695 DVDD.n4091 VSS 0.137328f
C9696 DVDD.n4092 VSS 0.11992f
C9697 DVDD.n4093 VSS 0.274656f
C9698 DVDD.n4094 VSS 0.274656f
C9699 DVDD.n4095 VSS 0.11992f
C9700 DVDD.n4096 VSS 0.274656f
C9701 DVDD.n4097 VSS 0.11992f
C9702 DVDD.n4098 VSS 0.274656f
C9703 DVDD.n4099 VSS 0.11992f
C9704 DVDD.n4100 VSS 0.274656f
C9705 DVDD.n4101 VSS 0.11992f
C9706 DVDD.n4102 VSS 0.274656f
C9707 DVDD.n4103 VSS 0.274656f
C9708 DVDD.n4104 VSS 0.274656f
C9709 DVDD.n4105 VSS 0.228235f
C9710 DVDD.n4106 VSS 0.228235f
C9711 DVDD.n4107 VSS 0.274656f
C9712 DVDD.n4108 VSS 0.239841f
C9713 DVDD.n4109 VSS 0.274656f
C9714 DVDD.n4110 VSS 0.11992f
C9715 DVDD.n4111 VSS 0.274656f
C9716 DVDD.n4112 VSS 0.274656f
C9717 DVDD.n4113 VSS 0.274656f
C9718 DVDD.n4114 VSS 0.274656f
C9719 DVDD.n4115 VSS 0.274656f
C9720 DVDD.n4116 VSS 0.11992f
C9721 DVDD.n4117 VSS 0.274656f
C9722 DVDD.n4118 VSS 0.11992f
C9723 DVDD.n4119 VSS 0.274656f
C9724 DVDD.n4120 VSS 0.274656f
C9725 DVDD.n4121 VSS 0.274656f
C9726 DVDD.n4122 VSS 0.274656f
C9727 DVDD.n4123 VSS 0.274656f
C9728 DVDD.n4124 VSS 0.11992f
C9729 DVDD.n4125 VSS 0.274656f
C9730 DVDD.n4126 VSS 0.11992f
C9731 DVDD.n4127 VSS 0.274656f
C9732 DVDD.n4128 VSS 0.274656f
C9733 DVDD.n4129 VSS 0.274656f
C9734 DVDD.n4130 VSS 0.274656f
C9735 DVDD.n4131 VSS 0.274656f
C9736 DVDD.n4132 VSS 0.11992f
C9737 DVDD.n4133 VSS 0.137328f
C9738 DVDD.n4134 VSS 0.11992f
C9739 DVDD.n4135 VSS 0.13346f
C9740 DVDD.n4136 VSS 3.48797f
C9741 DVDD.n4137 VSS 0.137328f
C9742 DVDD.n4138 VSS 0.11992f
C9743 DVDD.n4139 VSS 0.274656f
C9744 DVDD.n4140 VSS 0.274656f
C9745 DVDD.n4141 VSS 0.274656f
C9746 DVDD.n4142 VSS 0.274656f
C9747 DVDD.n4143 VSS 0.274656f
C9748 DVDD.n4144 VSS 0.274656f
C9749 DVDD.n4145 VSS 0.274656f
C9750 DVDD.n4146 VSS 0.274656f
C9751 DVDD.n4147 VSS 0.197288f
C9752 DVDD.n4148 VSS 0.274656f
C9753 DVDD.n4149 VSS 0.11992f
C9754 DVDD.n4150 VSS 0.274656f
C9755 DVDD.n4151 VSS 0.274656f
C9756 DVDD.n4152 VSS 0.274656f
C9757 DVDD.n4153 VSS 0.274656f
C9758 DVDD.n4154 VSS 0.274656f
C9759 DVDD.n4155 VSS 0.176012f
C9760 DVDD.n4156 VSS 0.048355f
C9761 DVDD.n4157 VSS 0.169049f
C9762 DVDD.n4158 VSS 0.098644f
C9763 DVDD.n4159 VSS 0.137328f
C9764 DVDD.n4160 VSS 0.11992f
C9765 DVDD.n4161 VSS 0.137328f
C9766 DVDD.n4163 VSS 0.125723f
C9767 DVDD.n4175 VSS 0.137328f
C9768 DVDD.n4176 VSS 0.11992f
C9769 DVDD.n4177 VSS 0.137328f
C9770 DVDD.n4178 VSS 3.48797f
C9771 DVDD.n4179 VSS 0.137328f
C9772 DVDD.n4180 VSS 0.201157f
C9773 DVDD.n4181 VSS 0.274656f
C9774 DVDD.n4182 VSS 0.274656f
C9775 DVDD.n4183 VSS 0.274656f
C9776 DVDD.n4184 VSS 0.274656f
C9777 DVDD.n4185 VSS 0.274656f
C9778 DVDD.n4186 VSS 0.274656f
C9779 DVDD.n4187 VSS 0.205025f
C9780 DVDD.n4188 VSS 0.274656f
C9781 DVDD.n4189 VSS 0.274656f
C9782 DVDD.n4190 VSS 0.11992f
C9783 DVDD.n4191 VSS 0.11992f
C9784 DVDD.n4192 VSS 0.11992f
C9785 DVDD.n4193 VSS 0.274656f
C9786 DVDD.n4194 VSS 0.274656f
C9787 DVDD.n4195 VSS 0.11992f
C9788 DVDD.n4196 VSS 0.11992f
C9789 DVDD.n4197 VSS 0.11992f
C9790 DVDD.n4198 VSS 0.168275f
C9791 DVDD.n4199 VSS 0.089747f
C9792 DVDD.n4200 VSS 0.129978f
C9793 DVDD.n4201 VSS 0.274656f
C9794 DVDD.n4202 VSS 0.21057f
C9795 DVDD.n4203 VSS 0.11992f
C9796 DVDD.n4204 VSS 0.11992f
C9797 DVDD.n4205 VSS 0.11992f
C9798 DVDD.n4206 VSS 0.274656f
C9799 DVDD.n4207 VSS 0.274656f
C9800 DVDD.n4208 VSS 0.19342f
C9801 DVDD.n4209 VSS 0.274656f
C9802 DVDD.n4210 VSS 0.274656f
C9803 DVDD.n4211 VSS 0.274656f
C9804 DVDD.n4212 VSS 0.274656f
C9805 DVDD.n4213 VSS 0.11992f
C9806 DVDD.n4214 VSS 0.11992f
C9807 DVDD.n4215 VSS 0.11992f
C9808 DVDD.n4216 VSS 0.274656f
C9809 DVDD.n4217 VSS 0.274656f
C9810 DVDD.n4218 VSS 0.11992f
C9811 DVDD.n4219 VSS 0.11992f
C9812 DVDD.n4220 VSS 0.11992f
C9813 DVDD.n4221 VSS 0.274656f
C9814 DVDD.n4222 VSS 0.274656f
C9815 DVDD.n4223 VSS 0.11992f
C9816 DVDD.n4224 VSS 0.11992f
C9817 DVDD.n4225 VSS 0.11992f
C9818 DVDD.n4226 VSS 0.274656f
C9819 DVDD.n4227 VSS 0.274656f
C9820 DVDD.n4228 VSS 0.11992f
C9821 DVDD.n4229 VSS 0.163891f
C9822 DVDD.n4230 VSS 0.163891f
C9823 DVDD.n4231 VSS 0.163891f
C9824 DVDD.n4232 VSS 0.163891f
C9825 DVDD.n4233 VSS 0.163891f
C9826 DVDD.n4234 VSS 0.163891f
C9827 DVDD.n4235 VSS 0.163891f
C9828 DVDD.n4236 VSS 0.163891f
C9829 DVDD.n4237 VSS 0.163891f
C9830 DVDD.n4238 VSS 0.163891f
C9831 DVDD.n4239 VSS 0.163891f
C9832 DVDD.n4240 VSS 0.070147f
C9833 DVDD.n4241 VSS 0.073242f
C9834 DVDD.n4242 VSS 0.036964f
C9835 DVDD.n4243 VSS 0.069115f
C9836 DVDD.n4244 VSS 0.073242f
C9837 DVDD.n4245 VSS 0.073242f
C9838 DVDD.n4246 VSS 0.073242f
C9839 DVDD.n4248 VSS 0.073242f
C9840 DVDD.n4249 VSS 0.068084f
C9841 DVDD.n4250 VSS 0.073242f
C9842 DVDD.n4251 VSS 0.067052f
C9843 DVDD.n4252 VSS 0.063957f
C9844 DVDD.n4253 VSS 0.163891f
C9845 DVDD.n4254 VSS 0.163891f
C9846 DVDD.n4255 VSS 0.130849f
C9847 DVDD.n4256 VSS 0.163891f
C9848 DVDD.n4257 VSS 0.163891f
C9849 DVDD.n4258 VSS 0.063957f
C9850 DVDD.n4262 VSS 1.37325f
C9851 DVDD.n4264 VSS 0.163891f
C9852 DVDD.n4265 VSS 0.104414f
C9853 DVDD.n4268 VSS 0.163891f
C9854 DVDD.n4269 VSS 0.017666f
C9855 DVDD.n4271 VSS 0.063957f
C9856 DVDD.n4274 VSS 0.146483f
C9857 DVDD.n4275 VSS 0.063957f
C9858 DVDD.n4276 VSS 0.146483f
C9859 DVDD.n4277 VSS 0.146483f
C9860 DVDD.n4278 VSS 0.063957f
C9861 DVDD.n4279 VSS 0.146483f
C9862 DVDD.n4280 VSS 0.063957f
C9863 DVDD.n4281 VSS 0.104963f
C9864 DVDD.n4282 VSS 0.104963f
C9865 DVDD.n4283 VSS 0.01831f
C9866 DVDD.n4284 VSS 0.036621f
C9867 DVDD.n4285 VSS 0.037194f
C9868 DVDD.n4286 VSS 0.036621f
C9869 DVDD.n4287 VSS 0.016376f
C9870 DVDD.n4288 VSS 0.015989f
C9871 DVDD.n4289 VSS 0.01831f
C9872 DVDD.n4290 VSS 0.015989f
C9873 DVDD.n4291 VSS 0.01831f
C9874 DVDD.n4292 VSS 0.015989f
C9875 DVDD.n4293 VSS 0.036621f
C9876 DVDD.n4294 VSS 0.105852f
C9877 DVDD.n4295 VSS 0.036621f
C9878 DVDD.n4296 VSS 0.02695f
C9879 DVDD.n4297 VSS 0.02695f
C9880 DVDD.n4298 VSS 0.015989f
C9881 DVDD.n4299 VSS 0.01831f
C9882 DVDD.n4300 VSS 0.036621f
C9883 DVDD.n4301 VSS 0.035087f
C9884 DVDD.n4302 VSS 0.015989f
C9885 DVDD.n4303 VSS 0.01831f
C9886 DVDD.n4304 VSS 0.015989f
C9887 DVDD.n4305 VSS 0.016634f
C9888 DVDD.n4306 VSS 0.036277f
C9889 DVDD.n4307 VSS 0.015989f
C9890 DVDD.n4308 VSS 0.036621f
C9891 DVDD.n4309 VSS 0.036621f
C9892 DVDD.n4310 VSS 0.103874f
C9893 DVDD.n4311 VSS 0.036621f
C9894 DVDD.n4312 VSS 0.027981f
C9895 DVDD.n4313 VSS 0.027981f
C9896 DVDD.n4314 VSS 0.015989f
C9897 DVDD.n4315 VSS 0.063957f
C9898 DVDD.n4316 VSS 0.146483f
C9899 DVDD.n4317 VSS 0.146483f
C9900 DVDD.n4318 VSS 0.146483f
C9901 DVDD.n4319 VSS 0.103157f
C9902 DVDD.n4320 VSS 0.146483f
C9903 DVDD.n4321 VSS 0.146483f
C9904 DVDD.n4322 VSS 0.146483f
C9905 DVDD.n4323 VSS 0.073242f
C9906 DVDD.n4324 VSS 0.163891f
C9907 DVDD.n4325 VSS 0.130849f
C9908 DVDD.n4326 VSS 0.163891f
C9909 DVDD.n4327 VSS 0.163891f
C9910 DVDD.n4328 VSS 0.163891f
C9911 DVDD.n4329 VSS 1.37325f
C9912 DVDD.n4331 VSS 0.163891f
C9913 DVDD.n4332 VSS 0.163891f
C9914 DVDD.t53 VSS 0.016763f
C9915 DVDD.t41 VSS 0.016763f
C9916 DVDD.n4333 VSS 0.039884f
C9917 DVDD.n4334 VSS 0.034701f
C9918 DVDD.t35 VSS 0.044262f
C9919 DVDD.n4335 VSS 0.053534f
C9920 DVDD.t23 VSS 0.016763f
C9921 DVDD.t37 VSS 0.016763f
C9922 DVDD.n4336 VSS 0.039884f
C9923 DVDD.n4337 VSS 0.034701f
C9924 DVDD.n4338 VSS 0.033491f
C9925 DVDD.n4339 VSS 0.045909f
C9926 DVDD.t9 VSS 0.016763f
C9927 DVDD.t5 VSS 0.016763f
C9928 DVDD.n4340 VSS 0.039884f
C9929 DVDD.n4341 VSS 0.034701f
C9930 DVDD.t154 VSS 0.016763f
C9931 DVDD.t11 VSS 0.016763f
C9932 DVDD.n4342 VSS 0.062036f
C9933 DVDD.n4343 VSS 0.033491f
C9934 DVDD.n4344 VSS 0.031915f
C9935 DVDD.n4345 VSS 0.050792f
C9936 DVDD.n4346 VSS 0.033491f
C9937 DVDD.n4347 VSS 0.033491f
C9938 DVDD.t3 VSS 0.016763f
C9939 DVDD.t7 VSS 0.016763f
C9940 DVDD.n4348 VSS 0.039884f
C9941 DVDD.n4349 VSS 0.034701f
C9942 DVDD.t1 VSS 0.044262f
C9943 DVDD.n4350 VSS 0.053534f
C9944 DVDD.n4351 VSS 0.078464f
C9945 DVDD.n4352 VSS 0.033043f
C9946 DVDD.n4353 VSS 0.32679f
C9947 DVDD.t0 VSS 0.338768f
C9948 DVDD.t6 VSS 0.24195f
C9949 DVDD.t2 VSS 0.24195f
C9950 DVDD.t4 VSS 0.24195f
C9951 DVDD.t8 VSS 0.24195f
C9952 DVDD.t10 VSS 0.24195f
C9953 DVDD.t153 VSS 0.327228f
C9954 DVDD.t34 VSS 0.327228f
C9955 DVDD.t36 VSS 0.24195f
C9956 DVDD.t22 VSS 0.24195f
C9957 DVDD.t40 VSS 0.24195f
C9958 DVDD.t52 VSS 0.24195f
C9959 DVDD.t18 VSS 0.24195f
C9960 DVDD.t26 VSS 0.24195f
C9961 DVDD.t56 VSS 0.199311f
C9962 DVDD.n4354 VSS -0.124359f
C9963 DVDD.t59 VSS 0.016763f
C9964 DVDD.t57 VSS 0.016763f
C9965 DVDD.n4355 VSS 0.062036f
C9966 DVDD.t47 VSS 0.016763f
C9967 DVDD.t39 VSS 0.016763f
C9968 DVDD.n4356 VSS 0.039884f
C9969 DVDD.n4357 VSS 0.034701f
C9970 DVDD.t43 VSS 0.016763f
C9971 DVDD.t15 VSS 0.016763f
C9972 DVDD.n4358 VSS 0.039884f
C9973 DVDD.n4359 VSS 0.034701f
C9974 DVDD.t21 VSS 0.016763f
C9975 DVDD.t45 VSS 0.016763f
C9976 DVDD.n4360 VSS 0.039884f
C9977 DVDD.n4361 VSS 0.034701f
C9978 DVDD.n4362 VSS 0.107265f
C9979 DVDD.t49 VSS 0.016763f
C9980 DVDD.t29 VSS 0.016763f
C9981 DVDD.n4363 VSS 0.039884f
C9982 DVDD.n4364 VSS 0.034701f
C9983 DVDD.t25 VSS 0.016763f
C9984 DVDD.t61 VSS 0.016763f
C9985 DVDD.n4365 VSS 0.062036f
C9986 DVDD.t51 VSS 0.016763f
C9987 DVDD.t33 VSS 0.016763f
C9988 DVDD.n4366 VSS 0.039884f
C9989 DVDD.n4367 VSS 0.034701f
C9990 DVDD.t31 VSS 0.016763f
C9991 DVDD.t17 VSS 0.016763f
C9992 DVDD.n4368 VSS 0.039884f
C9993 DVDD.n4369 VSS 0.034701f
C9994 DVDD.t55 VSS 0.044262f
C9995 DVDD.n4370 VSS 0.053534f
C9996 DVDD.t58 VSS 0.163614f
C9997 DVDD.t38 VSS 0.24195f
C9998 DVDD.t46 VSS 0.24195f
C9999 DVDD.t14 VSS 0.24195f
C10000 DVDD.t42 VSS 0.24195f
C10001 DVDD.t44 VSS 0.24195f
C10002 DVDD.t20 VSS 0.24195f
C10003 DVDD.t28 VSS 0.24195f
C10004 DVDD.t48 VSS 0.24195f
C10005 DVDD.t60 VSS 0.24195f
C10006 DVDD.t24 VSS 0.24195f
C10007 DVDD.t32 VSS 0.24195f
C10008 DVDD.t50 VSS 0.24195f
C10009 DVDD.t16 VSS 0.24195f
C10010 DVDD.t30 VSS 0.24195f
C10011 DVDD.t54 VSS 0.338786f
C10012 DVDD.n4371 VSS 0.100933f
C10013 DVDD.n4372 VSS 0.320853f
C10014 DVDD.n4373 VSS 0.045515f
C10015 DVDD.n4374 VSS 0.033491f
C10016 DVDD.n4375 VSS 0.033491f
C10017 DVDD.n4376 VSS 0.052371f
C10018 DVDD.n4377 VSS 0.033491f
C10019 DVDD.n4378 VSS 0.033491f
C10020 DVDD.n4379 VSS 0.033491f
C10021 DVDD.n4380 VSS 0.033491f
C10022 DVDD.n4381 VSS -0.192963f
C10023 DVDD.n4382 VSS 0.033491f
C10024 DVDD.t27 VSS 0.016763f
C10025 DVDD.t19 VSS 0.016763f
C10026 DVDD.n4383 VSS 0.039884f
C10027 DVDD.n4384 VSS 0.034701f
C10028 DVDD.n4385 VSS 0.107262f
C10029 DVDD.n4386 VSS 0.114988f
C10030 DVDD.n4387 VSS 0.163891f
C10031 DVDD.n4389 VSS 0.073242f
C10032 DVDD.n4390 VSS 0.07221f
C10033 DVDD.n4391 VSS 0.073242f
C10034 DVDD.n4392 VSS 0.073242f
C10035 DVDD.n4393 VSS 0.073242f
C10036 DVDD.n4394 VSS 0.071178f
C10037 DVDD.n4398 VSS 0.063957f
C10038 DVDD.n4399 VSS 0.073242f
C10039 DVDD.n4401 VSS 0.066021f
C10040 DVDD.n4402 VSS 0.073242f
C10041 DVDD.n4403 VSS 0.073242f
C10042 DVDD.n4405 VSS 0.064989f
C10043 DVDD.n4406 VSS 0.073242f
C10044 DVDD.n4407 VSS 0.109347f
C10045 DVDD.n4412 VSS 0.146483f
C10046 DVDD.n4413 VSS 0.063957f
C10047 DVDD.n4414 VSS 0.146483f
C10048 DVDD.n4415 VSS 0.427183f
C10049 DVDD.n4416 VSS 0.174683f
C10050 DVDD.n4419 VSS 0.073242f
C10051 DVDD.n4420 VSS 0.063957f
C10052 DVDD.n4421 VSS 0.146483f
C10053 DVDD.n4422 VSS 0.146483f
C10054 DVDD.n4423 VSS 0.063957f
C10055 DVDD.n4424 VSS 0.146483f
C10056 DVDD.n4425 VSS 0.063957f
C10057 DVDD.n4426 VSS 0.146483f
C10058 DVDD.n4427 VSS 0.063957f
C10059 DVDD.n4428 VSS 0.125852f
C10060 DVDD.n4429 VSS 0.063957f
C10061 DVDD.n4430 VSS 0.146483f
C10062 DVDD.n4431 VSS 0.146483f
C10063 DVDD.n4432 VSS 0.063957f
C10064 DVDD.n4433 VSS 0.146483f
C10065 DVDD.n4434 VSS 0.063957f
C10066 DVDD.n4435 VSS 0.146483f
C10067 DVDD.n4436 VSS 0.146483f
C10068 DVDD.n4437 VSS 0.146483f
C10069 DVDD.n4438 VSS 0.146483f
C10070 DVDD.n4439 VSS 0.146483f
C10071 DVDD.n4441 VSS 0.070147f
C10072 DVDD.n4442 VSS 0.063957f
C10073 DVDD.n4443 VSS 0.146483f
C10074 DVDD.n4444 VSS 0.063957f
C10075 DVDD.n4445 VSS 0.146483f
C10076 DVDD.n4446 VSS 0.146483f
C10077 DVDD.n4447 VSS 0.146483f
C10078 DVDD.n4448 VSS 0.135136f
C10079 DVDD.n4449 VSS 0.135136f
C10080 DVDD.n4450 VSS 0.095936f
C10081 DVDD.n4451 VSS 0.16536f
C10082 DVDD.n4452 VSS 0.165891f
C10083 DVDD.n4453 VSS 0.40999f
C10084 DVDD.n4454 VSS 0.097999f
C10085 DVDD.n4455 VSS 0.097999f
C10086 DVDD.n4456 VSS 0.097999f
C10087 DVDD.n4457 VSS 0.146483f
C10088 DVDD.n4458 VSS 0.146483f
C10089 DVDD.n4459 VSS 0.063957f
C10090 DVDD.n4460 VSS 0.146483f
C10091 DVDD.n4461 VSS 0.146483f
C10092 DVDD.n4462 VSS 0.11992f
C10093 DVDD.n4463 VSS 0.163891f
C10094 DVDD.n4464 VSS 0.163891f
C10095 DVDD.n4465 VSS 0.163891f
C10096 DVDD.n4466 VSS 0.163891f
C10097 DVDD.n4467 VSS 0.163891f
C10098 DVDD.n4468 VSS 0.163891f
C10099 DVDD.n4469 VSS 0.163891f
C10100 DVDD.n4470 VSS 0.163891f
C10101 DVDD.n4471 VSS 0.163891f
C10102 DVDD.n4472 VSS 0.163891f
C10103 DVDD.n4473 VSS 0.163891f
C10104 DVDD.n4474 VSS 0.146483f
C10105 DVDD.n4475 VSS 0.063957f
C10106 DVDD.n4476 VSS 0.146483f
C10107 DVDD.n4477 VSS 0.129978f
C10108 DVDD.n4478 VSS 0.063957f
C10109 DVDD.n4479 VSS 0.163891f
C10110 DVDD.n4480 VSS 0.163891f
C10111 DVDD.n4481 VSS 0.163891f
C10112 DVDD.n4482 VSS 0.163891f
C10113 DVDD.n4483 VSS 0.163891f
C10114 DVDD.n4484 VSS 0.163891f
C10115 DVDD.n4485 VSS 0.163891f
C10116 DVDD.n4486 VSS 0.163891f
C10117 DVDD.n4487 VSS 0.163891f
C10118 DVDD.n4488 VSS 0.163891f
C10119 DVDD.n4491 VSS 0.137328f
C10120 DVDD.n4492 VSS 0.137328f
C10121 DVDD.n4493 VSS 0.121855f
C10122 DVDD.n4494 VSS 0.137328f
C10123 DVDD.n4495 VSS 0.137328f
C10124 DVDD.n4496 VSS 0.11992f
C10125 DVDD.n4497 VSS 0.137328f
C10126 DVDD.n4498 VSS 0.135394f
C10127 DVDD.n4499 VSS 0.11992f
C10128 DVDD.n4500 VSS 0.137328f
C10129 DVDD.n4501 VSS 0.137328f
C10130 DVDD.n4502 VSS 0.137328f
C10131 DVDD.n4503 VSS 0.13346f
C10132 DVDD.n4504 VSS 0.137328f
C10133 DVDD.n4505 VSS 0.11992f
C10134 DVDD.n4516 VSS 0.137328f
C10135 DVDD.n4528 VSS 0.123789f
C10136 DVDD.n4531 VSS 0.315887f
C10137 DVDD.n4532 VSS 0.137328f
C10138 DVDD.n4533 VSS 0.163891f
C10139 DVDD.n4534 VSS 0.21057f
C10140 DVDD.n4535 VSS 0.063957f
C10141 DVDD.n4536 VSS 0.089747f
C10142 DVDD.n4537 VSS 0.063957f
C10143 DVDD.n4538 VSS 0.146483f
C10144 DVDD.n4539 VSS 0.063957f
C10145 DVDD.n4540 VSS 0.146483f
C10146 DVDD.n4541 VSS 0.146483f
C10147 DVDD.n4542 VSS 0.146483f
C10148 DVDD.n4543 VSS 0.146483f
C10149 DVDD.n4544 VSS 0.063957f
C10150 DVDD.n4545 VSS 0.146483f
C10151 DVDD.n4546 VSS 0.063957f
C10152 DVDD.n4547 VSS 0.146483f
C10153 DVDD.n4548 VSS 0.063957f
C10154 DVDD.n4549 VSS 0.146483f
C10155 DVDD.n4550 VSS 0.146483f
C10156 DVDD.n4551 VSS 0.146483f
C10157 DVDD.n4552 VSS 0.146483f
C10158 DVDD.n4553 VSS 0.146483f
C10159 DVDD.n4554 VSS 0.063957f
C10160 DVDD.n4555 VSS 0.073242f
C10161 DVDD.n4557 VSS 0.315887f
C10162 DVDD.n4558 VSS 0.073242f
C10163 DVDD.n4559 VSS 0.063957f
C10164 DVDD.n4560 VSS 0.146483f
C10165 DVDD.n4561 VSS 0.146483f
C10166 DVDD.n4562 VSS 0.146483f
C10167 DVDD.n4563 VSS 0.146483f
C10168 DVDD.n4564 VSS 0.146483f
C10169 DVDD.n4565 VSS 0.146483f
C10170 DVDD.n4566 VSS 0.146483f
C10171 DVDD.n4567 VSS 0.086652f
C10172 DVDD.n4568 VSS 0.146483f
C10173 DVDD.n4569 VSS 0.146483f
C10174 DVDD.n4570 VSS 0.146483f
C10175 DVDD.n4571 VSS 0.13101f
C10176 DVDD.n4572 VSS 0.13101f
C10177 DVDD.n4573 VSS 0.062926f
C10178 DVDD.n4574 VSS 0.104963f
C10179 DVDD.n4575 VSS 0.050547f
C10180 DVDD.n4576 VSS 0.102126f
C10181 DVDD.n4577 VSS 0.102126f
C10182 DVDD.n4578 VSS 0.146483f
C10183 DVDD.n4579 VSS 0.146483f
C10184 DVDD.n4580 VSS 0.146483f
C10185 DVDD.n4581 VSS 0.146483f
C10186 DVDD.n4582 VSS 0.146483f
C10187 DVDD.n4583 VSS 0.146483f
C10188 DVDD.n4584 VSS 0.146483f
C10189 DVDD.n4585 VSS 0.146483f
C10190 DVDD.n4586 VSS 0.085621f
C10191 DVDD.n4587 VSS 0.085621f
C10192 DVDD.n4588 VSS 0.146483f
C10193 DVDD.n4589 VSS 0.146483f
C10194 DVDD.n4590 VSS 0.125852f
C10195 DVDD.n4591 VSS 0.146483f
C10196 DVDD.n4592 VSS 0.146483f
C10197 DVDD.n4593 VSS 0.146483f
C10198 DVDD.n4594 VSS 0.146483f
C10199 DVDD.n4595 VSS 0.146483f
C10200 DVDD.n4596 VSS 0.063957f
C10201 DVDD.n4597 VSS 0.073242f
C10202 DVDD.n4599 VSS 0.163891f
C10203 DVDD.n4600 VSS 0.073242f
C10204 DVDD.n4601 VSS 0.315887f
C10205 DVDD.n4602 VSS 0.315887f
C10206 DVDD.n4603 VSS 0.163891f
C10207 DVDD.n4604 VSS 0.163891f
C10208 DVDD.n4605 VSS 0.163891f
C10209 DVDD.n4606 VSS 0.163891f
C10210 DVDD.n4607 VSS 0.163891f
C10211 DVDD.n4608 VSS 0.163891f
C10212 DVDD.n4609 VSS 0.163891f
C10213 DVDD.n4610 VSS 0.163891f
C10214 DVDD.n4611 VSS 0.163891f
C10215 DVDD.n4612 VSS 0.163891f
C10216 DVDD.n4613 VSS 0.163891f
C10217 DVDD.n4626 VSS 0.137328f
C10218 DVDD.n4627 VSS 0.131525f
C10219 DVDD.n4628 VSS 0.137328f
C10220 DVDD.n4629 VSS 0.137328f
C10221 DVDD.n4630 VSS 0.137328f
C10222 DVDD.n4631 VSS 0.129591f
C10223 DVDD.n4632 VSS 0.162473f
C10224 DVDD.n4633 VSS 0.137328f
C10225 DVDD.n4635 VSS 0.127657f
C10226 DVDD.n4636 VSS 0.137328f
C10227 DVDD.n4637 VSS 0.11992f
C10228 DVDD.n4638 VSS 0.137328f
C10229 DVDD.n4639 VSS 0.137328f
C10230 DVDD.n4640 VSS 0.11992f
C10231 DVDD.n4642 VSS 0.125723f
C10232 DVDD.n4643 VSS 0.137328f
C10233 DVDD.n4655 VSS 0.137328f
C10234 DVDD.n4656 VSS 0.11992f
C10235 DVDD.n4657 VSS 0.137328f
C10236 DVDD.n4658 VSS 3.48797f
C10237 DVDD.n4659 VSS 0.137328f
C10238 DVDD.n4660 VSS 0.235972f
C10239 DVDD.n4661 VSS 0.274656f
C10240 DVDD.n4662 VSS 0.160538f
C10241 DVDD.n4663 VSS 0.160538f
C10242 DVDD.n4664 VSS 0.274656f
C10243 DVDD.n4665 VSS 0.274656f
C10244 DVDD.n4666 VSS 0.274656f
C10245 DVDD.n4667 VSS 0.274656f
C10246 DVDD.n4668 VSS 0.274656f
C10247 DVDD.n4669 VSS 0.274656f
C10248 DVDD.n4670 VSS 0.274656f
C10249 DVDD.n4671 VSS 0.274656f
C10250 DVDD.n4672 VSS 0.274656f
C10251 DVDD.n4673 VSS 0.274656f
C10252 DVDD.n4674 VSS 0.274656f
C10253 DVDD.n4675 VSS 0.274656f
C10254 DVDD.n4676 VSS 0.274656f
C10255 DVDD.n4677 VSS 0.274656f
C10256 DVDD.n4678 VSS 0.274656f
C10257 DVDD.n4679 VSS 0.274656f
C10258 DVDD.n4680 VSS 0.274656f
C10259 DVDD.n4681 VSS 0.274656f
C10260 DVDD.n4682 VSS 0.274656f
C10261 DVDD.n4683 VSS 0.274656f
C10262 DVDD.n4684 VSS 0.274656f
C10263 DVDD.n4685 VSS 0.274656f
C10264 DVDD.n4686 VSS 0.274656f
C10265 DVDD.n4687 VSS 0.274656f
C10266 DVDD.n4688 VSS 0.274656f
C10267 DVDD.n4689 VSS 0.274656f
C10268 DVDD.n4690 VSS 0.274656f
C10269 DVDD.n4691 VSS 0.274656f
C10270 DVDD.n4692 VSS 0.274656f
C10271 DVDD.n4693 VSS 0.274656f
C10272 DVDD.n4694 VSS 0.274656f
C10273 DVDD.n4695 VSS 0.274656f
C10274 DVDD.n4696 VSS 0.274656f
C10275 DVDD.n4697 VSS 0.243709f
C10276 DVDD.n4698 VSS 0.243709f
C10277 DVDD.n4699 VSS 0.21057f
C10278 DVDD.n4700 VSS 0.168275f
C10279 DVDD.n4701 VSS 0.274656f
C10280 DVDD.n4702 VSS 0.274656f
C10281 DVDD.n4703 VSS 0.274656f
C10282 DVDD.n4704 VSS 0.274656f
C10283 DVDD.n4705 VSS 0.274656f
C10284 DVDD.n4706 VSS 0.274656f
C10285 DVDD.n4707 VSS 0.274656f
C10286 DVDD.n4708 VSS 0.274656f
C10287 DVDD.n4709 VSS 0.274656f
C10288 DVDD.n4710 VSS 0.274656f
C10289 DVDD.n4711 VSS 0.274656f
C10290 DVDD.n4712 VSS 0.274656f
C10291 DVDD.n4713 VSS 0.274656f
C10292 DVDD.n4714 VSS 0.274656f
C10293 DVDD.n4715 VSS 0.274656f
C10294 DVDD.n4716 VSS 0.274656f
C10295 DVDD.n4717 VSS 0.274656f
C10296 DVDD.n4718 VSS 0.274656f
C10297 DVDD.n4719 VSS 0.274656f
C10298 DVDD.n4720 VSS 0.274656f
C10299 DVDD.n4721 VSS 0.274656f
C10300 DVDD.n4722 VSS 0.274656f
C10301 DVDD.n4723 VSS 0.274656f
C10302 DVDD.n4724 VSS 0.274656f
C10303 DVDD.n4725 VSS 0.274656f
C10304 DVDD.n4726 VSS 0.274656f
C10305 DVDD.n4727 VSS 0.274656f
C10306 DVDD.n4728 VSS 0.274656f
C10307 DVDD.n4729 VSS 0.274656f
C10308 DVDD.n4730 VSS 0.274656f
C10309 DVDD.n4731 VSS 0.274656f
C10310 DVDD.n4732 VSS 0.274656f
C10311 DVDD.n4733 VSS 0.274656f
C10312 DVDD.n4734 VSS 0.235972f
C10313 DVDD.n4735 VSS 0.235972f
C10314 DVDD.n4736 VSS 0.21057f
C10315 DVDD.n4737 VSS 0.093873f
C10316 DVDD.n4738 VSS 0.146483f
C10317 DVDD.n4739 VSS 0.146483f
C10318 DVDD.n4740 VSS 0.063957f
C10319 DVDD.n4741 VSS 0.073242f
C10320 DVDD.n4742 VSS 0.163891f
C10321 DVDD.n4743 VSS 0.073242f
C10322 DVDD.n4744 VSS 0.10522f
C10323 DVDD.n4745 VSS 0.146483f
C10324 DVDD.n4746 VSS 0.146483f
C10325 DVDD.n4747 VSS 0.146483f
C10326 DVDD.n4748 VSS 0.146483f
C10327 DVDD.n4749 VSS 0.146483f
C10328 DVDD.n4750 VSS 0.146483f
C10329 DVDD.n4751 VSS 0.084589f
C10330 DVDD.n4752 VSS 0.073242f
C10331 DVDD.n4753 VSS 0.063957f
C10332 DVDD.n4754 VSS 0.146483f
C10333 DVDD.n4755 VSS 0.146483f
C10334 DVDD.n4756 VSS 0.146483f
C10335 DVDD.n4757 VSS 0.093873f
C10336 DVDD.n4758 VSS 0.093873f
C10337 DVDD.n4759 VSS 0.104963f
C10338 DVDD.n4760 VSS 0.063957f
C10339 DVDD.n4761 VSS 0.139262f
C10340 DVDD.n4762 VSS 0.139262f
C10341 DVDD.n4763 VSS 0.146483f
C10342 DVDD.n4764 VSS 0.146483f
C10343 DVDD.n4765 VSS 0.146483f
C10344 DVDD.n4766 VSS 0.063957f
C10345 DVDD.n4767 VSS 0.073242f
C10346 DVDD.n4768 VSS 0.163891f
C10347 DVDD.n4769 VSS 0.073242f
C10348 DVDD.n4770 VSS 0.063957f
C10349 DVDD.n4771 VSS 0.146483f
C10350 DVDD.n4772 VSS 0.146483f
C10351 DVDD.n4773 VSS 0.146483f
C10352 DVDD.n4774 VSS 0.146483f
C10353 DVDD.n4775 VSS 0.146483f
C10354 DVDD.n4776 VSS 0.127915f
C10355 DVDD.n4777 VSS 0.146483f
C10356 DVDD.n4778 VSS 0.121726f
C10357 DVDD.n4779 VSS 0.121726f
C10358 DVDD.n4780 VSS 0.121726f
C10359 DVDD.n4781 VSS 0.21057f
C10360 DVDD.n4782 VSS 0.183749f
C10361 DVDD.n4783 VSS 0.183749f
C10362 DVDD.n4784 VSS 0.274656f
C10363 DVDD.n4785 VSS 0.274656f
C10364 DVDD.n4786 VSS 0.274656f
C10365 DVDD.n4787 VSS 0.274656f
C10366 DVDD.n4788 VSS 0.274656f
C10367 DVDD.n4789 VSS 0.274656f
C10368 DVDD.n4790 VSS 0.274656f
C10369 DVDD.n4791 VSS 0.274656f
C10370 DVDD.n4792 VSS 0.274656f
C10371 DVDD.n4793 VSS 0.274656f
C10372 DVDD.n4794 VSS 0.274656f
C10373 DVDD.n4795 VSS 0.274656f
C10374 DVDD.n4796 VSS 0.274656f
C10375 DVDD.n4797 VSS 0.274656f
C10376 DVDD.n4798 VSS 0.274656f
C10377 DVDD.n4799 VSS 0.274656f
C10378 DVDD.n4800 VSS 1.26379f
C10379 DVDD.n4801 VSS 0.274656f
C10380 DVDD.n4802 VSS 0.461394f
C10381 DVDD.n4803 VSS 0.11992f
C10382 DVDD.n4805 VSS 0.151899f
C10383 DVDD.n4807 VSS 0.151899f
C10384 DVDD.n4809 VSS 0.151899f
C10385 DVDD.n4811 VSS 0.151899f
C10386 DVDD.n4813 VSS 0.151899f
C10387 DVDD.n4815 VSS 0.151899f
C10388 DVDD.n4817 VSS 0.151899f
C10389 DVDD.n4819 VSS 0.151899f
C10390 DVDD.n4821 VSS 0.151899f
C10391 DVDD.n4823 VSS 0.151899f
C10392 DVDD.n4834 VSS 0.128624f
C10393 DVDD.n4837 VSS 0.151899f
C10394 DVDD.n4838 VSS 0.908236f
C10395 DVDD.n4839 VSS 0.292773f
C10396 DVDD.n4840 VSS 0.151899f
C10397 DVDD.n4842 VSS 0.151899f
C10398 DVDD.n4845 VSS 0.292773f
C10399 DVDD.n4846 VSS 0.079661f
C10400 DVDD.n4847 VSS 0.079148f
C10401 DVDD.n4848 VSS 0.229561f
C10402 DVDD.n4849 VSS 0.079009f
C10403 DVDD.n4850 VSS 0.034496f
C10404 DVDD.n4851 VSS 0.039504f
C10405 DVDD.n4852 VSS 0.151899f
C10406 DVDD.n4854 VSS 0.151899f
C10407 DVDD.n4856 VSS 0.151899f
C10408 DVDD.n4857 VSS 0.039504f
C10409 DVDD.n4858 VSS 0.034496f
C10410 DVDD.n4859 VSS 0.058144f
C10411 DVDD.n4860 VSS 0.058144f
C10412 DVDD.n4861 VSS 0.056009f
C10413 DVDD.n4862 VSS 0.06037f
C10414 DVDD.n4863 VSS 0.06037f
C10415 DVDD.n4864 VSS 0.034496f
C10416 DVDD.n4865 VSS 0.034496f
C10417 DVDD.n4866 VSS 0.039504f
C10418 DVDD.n4867 VSS 0.151899f
C10419 DVDD.n4869 VSS 0.151899f
C10420 DVDD.n4871 VSS 0.151899f
C10421 DVDD.n4873 VSS 0.151899f
C10422 DVDD.n4874 VSS 0.038113f
C10423 DVDD.n4875 VSS 0.034496f
C10424 DVDD.n4876 VSS 0.079009f
C10425 DVDD.n4877 VSS 0.225252f
C10426 DVDD.n4878 VSS 0.074683f
C10427 DVDD.n4879 VSS 0.078141f
C10428 DVDD.n4880 VSS 1.27277f
C10429 DVDD.n4881 VSS 1.27277f
C10430 DVDD.n4882 VSS 0.151899f
C10431 DVDD.n4883 VSS 0.151899f
C10432 DVDD.n4884 VSS 0.05145f
C10433 DVDD.n4885 VSS 0.06615f
C10434 DVDD.n4886 VSS 0.06615f
C10435 DVDD.n4887 VSS 0.06615f
C10436 DVDD.n4888 VSS 0.06615f
C10437 DVDD.n4889 VSS 0.06615f
C10438 DVDD.n4890 VSS 0.06615f
C10439 DVDD.n4891 VSS 0.132299f
C10440 DVDD.n4892 VSS 0.06615f
C10441 DVDD.n4893 VSS 0.075949f
C10442 DVDD.n4896 VSS 0.128624f
C10443 DVDD.n4899 VSS 0.137328f
C10444 DVDD.n4900 VSS 0.137328f
C10445 DVDD.n4901 VSS 0.137328f
C10446 DVDD.n4902 VSS 0.12669f
C10447 DVDD.n4903 VSS 0.137328f
C10448 DVDD.n4904 VSS 0.137328f
C10449 DVDD.n4905 VSS 0.132299f
C10450 DVDD.n4906 VSS 0.026573f
C10451 DVDD.n4908 VSS 0.025624f
C10452 DVDD.n4909 VSS 0.025624f
C10453 DVDD.n4910 VSS 0.025624f
C10454 DVDD.n4911 VSS 0.025624f
C10455 DVDD.n4912 VSS 0.025624f
C10456 DVDD.n4913 VSS 0.025624f
C10457 DVDD.n4914 VSS 0.025624f
C10458 DVDD.n4915 VSS 0.025624f
C10459 DVDD.n4916 VSS 0.025624f
C10460 DVDD.n4919 VSS 0.025624f
C10461 DVDD.n4922 VSS 0.025624f
C10462 DVDD.n4925 VSS 0.025624f
C10463 DVDD.n4928 VSS 0.025624f
C10464 DVDD.n4931 VSS 0.025624f
C10465 DVDD.n4934 VSS 0.025624f
C10466 DVDD.n4937 VSS 0.025624f
C10467 DVDD.n4940 VSS 0.025624f
C10468 DVDD.n4944 VSS 0.025624f
C10469 DVDD.n4945 VSS 0.025624f
C10470 DVDD.n4946 VSS 0.025624f
C10471 DVDD.n4947 VSS 0.025624f
C10472 DVDD.n4948 VSS 0.025624f
C10473 DVDD.n4949 VSS 0.025624f
C10474 DVDD.n4950 VSS 0.025624f
C10475 DVDD.n4951 VSS 0.025624f
C10476 DVDD.n4952 VSS 0.025624f
C10477 DVDD.n4955 VSS 0.025624f
C10478 DVDD.n4958 VSS 0.025624f
C10479 DVDD.n4961 VSS 0.025624f
C10480 DVDD.n4964 VSS 0.025624f
C10481 DVDD.n4967 VSS 0.025624f
C10482 DVDD.n4970 VSS 0.025624f
C10483 DVDD.n4973 VSS 0.025624f
C10484 DVDD.n4976 VSS 0.025624f
C10485 DVDD.n4977 VSS 0.081946f
C10486 DVDD.n4978 VSS 0.063349f
C10487 DVDD.n4979 VSS 0.063349f
C10488 DVDD.n4980 VSS 0.081946f
C10489 DVDD.n4981 VSS 0.098464f
C10490 DVDD.n4982 VSS 0.098464f
C10491 DVDD.n4985 VSS 0.035233f
C10492 DVDD.n4987 VSS 0.0294f
C10493 DVDD.n4988 VSS 0.025624f
C10494 DVDD.n4989 VSS 0.025624f
C10495 DVDD.n4990 VSS 0.025624f
C10496 DVDD.n4992 VSS 0.0196f
C10497 DVDD.n4995 VSS 0.030844f
C10498 DVDD.n4996 VSS 0.05635f
C10499 DVDD.n4997 VSS 0.06615f
C10500 DVDD.n4999 VSS 0.025624f
C10501 DVDD.n5000 VSS 0.06125f
C10502 DVDD.n5001 VSS 0.035233f
C10503 DVDD.n5002 VSS 0.06125f
C10504 DVDD.n5003 VSS 0.06615f
C10505 DVDD.n5004 VSS 0.013761f
C10506 DVDD.n5005 VSS 0.075949f
C10507 DVDD.n5006 VSS 0.025624f
C10508 DVDD.n5007 VSS 0.075949f
C10509 DVDD.n5008 VSS 0.025624f
C10510 DVDD.n5009 VSS 0.075949f
C10511 DVDD.n5010 VSS 0.025624f
C10512 DVDD.n5011 VSS 0.075949f
C10513 DVDD.n5012 VSS 0.025624f
C10514 DVDD.n5013 VSS 0.075949f
C10515 DVDD.n5014 VSS 0.025624f
C10516 DVDD.n5015 VSS 0.025624f
C10517 DVDD.n5016 VSS 0.0686f
C10518 DVDD.n5017 VSS 0.0735f
C10519 DVDD.n5018 VSS 0.025624f
C10520 DVDD.n5019 VSS 0.075949f
C10521 DVDD.n5020 VSS 0.025624f
C10522 DVDD.n5021 VSS 0.075949f
C10523 DVDD.n5022 VSS 0.025624f
C10524 DVDD.n5023 VSS 0.075949f
C10525 DVDD.n5024 VSS 0.025624f
C10526 DVDD.n5025 VSS 0.075949f
C10527 DVDD.n5026 VSS 0.025624f
C10528 DVDD.n5027 VSS 0.075949f
C10529 DVDD.n5028 VSS 0.025624f
C10530 DVDD.n5029 VSS 0.075949f
C10531 DVDD.n5030 VSS 0.025624f
C10532 DVDD.n5031 VSS 0.025624f
C10533 DVDD.n5032 VSS 0.075949f
C10534 DVDD.n5033 VSS 0.025624f
C10535 DVDD.n5034 VSS 0.075949f
C10536 DVDD.n5035 VSS 0.025624f
C10537 DVDD.n5036 VSS 0.075949f
C10538 DVDD.n5037 VSS 0.025624f
C10539 DVDD.n5038 VSS 0.025624f
C10540 DVDD.n5039 VSS 0.025624f
C10541 DVDD.n5041 VSS 0.137328f
C10542 DVDD.n5042 VSS 0.137328f
C10543 DVDD.n5043 VSS 0.137328f
C10544 DVDD.n5045 VSS 0.137328f
C10545 DVDD.n5046 VSS 0.137328f
C10546 DVDD.n5047 VSS 0.075949f
C10547 DVDD.n5048 VSS 0.137328f
C10548 DVDD.n5049 VSS 0.137328f
C10549 DVDD.n5050 VSS 0.137328f
C10550 DVDD.n5051 VSS 0.137328f
C10551 DVDD.n5052 VSS 0.137328f
C10552 DVDD.n5053 VSS 0.737752f
C10553 DVDD.n5054 VSS 0.06615f
C10554 DVDD.n5055 VSS 0.06615f
C10555 DVDD.n5056 VSS 0.06615f
C10556 DVDD.n5057 VSS 0.06615f
C10557 DVDD.n5058 VSS 0.06615f
C10558 DVDD.n5059 VSS 0.06615f
C10559 DVDD.n5060 VSS 0.06615f
C10560 DVDD.n5061 VSS 0.132299f
C10561 DVDD.n5062 VSS 0.06615f
C10562 DVDD.n5063 VSS 0.06615f
C10563 DVDD.n5064 VSS 0.06615f
C10564 DVDD.n5065 VSS 0.11992f
C10565 DVDD.n5066 VSS 0.06615f
C10566 DVDD.n5067 VSS 0.06615f
C10567 DVDD.n5068 VSS 0.06615f
C10568 DVDD.n5069 VSS 0.06615f
C10569 DVDD.n5070 VSS 0.06615f
C10570 DVDD.n5071 VSS 0.06615f
C10571 DVDD.n5072 VSS 0.06615f
C10572 DVDD.n5073 VSS 0.06615f
C10573 DVDD.n5074 VSS 0.06615f
C10574 DVDD.n5075 VSS 0.06615f
C10575 DVDD.n5076 VSS 0.06615f
C10576 DVDD.n5077 VSS 0.075949f
C10577 DVDD.n5078 VSS 0.12669f
C10578 DVDD.n5079 VSS 0.128624f
C10579 DVDD.n5080 VSS 0.117599f
C10580 DVDD.n5081 VSS 0.128624f
C10581 DVDD.n5082 VSS 0.11992f
C10582 DVDD.n5083 VSS 0.274656f
C10583 DVDD.n5084 VSS 0.274656f
C10584 DVDD.n5085 VSS 0.11992f
C10585 DVDD.n5086 VSS 0.274656f
C10586 DVDD.n5087 VSS 1.26285f
C10587 DVDD.n5088 VSS 0.355263f
C10588 DVDD.n5089 VSS 0.11992f
C10589 DVDD.n5090 VSS 0.274656f
C10590 DVDD.n5091 VSS 0.11992f
C10591 DVDD.n5092 VSS 0.274656f
C10592 DVDD.n5093 VSS 0.274656f
C10593 DVDD.n5094 VSS 0.274656f
C10594 DVDD.n5095 VSS 0.274656f
C10595 DVDD.n5096 VSS 0.11992f
C10596 DVDD.n5097 VSS 0.274656f
C10597 DVDD.n5098 VSS 0.11992f
C10598 DVDD.n5099 VSS 0.274656f
C10599 DVDD.n5100 VSS 0.11992f
C10600 DVDD.n5101 VSS 0.274656f
C10601 DVDD.n5102 VSS 0.274656f
C10602 DVDD.n5103 VSS 0.274656f
C10603 DVDD.n5104 VSS 0.274656f
C10604 DVDD.n5105 VSS 0.274656f
C10605 DVDD.n5106 VSS 0.274656f
C10606 DVDD.n5107 VSS 0.274656f
C10607 DVDD.n5108 VSS 0.274656f
C10608 DVDD.n5109 VSS 0.183749f
C10609 DVDD.n5110 VSS 0.183749f
C10610 DVDD.n5111 VSS 0.524168f
C10611 DVDD.n5112 VSS 0.274656f
C10612 DVDD.n5113 VSS 0.524168f
C10613 DVDD.n5114 VSS 0.228235f
C10614 DVDD.n5115 VSS 0.274656f
C10615 DVDD.n5116 VSS 0.274656f
C10616 DVDD.n5117 VSS 0.274656f
C10617 DVDD.n5118 VSS 0.085911f
C10618 DVDD.n5119 VSS 0.163891f
C10619 DVDD.n5120 VSS 0.091198f
C10620 DVDD.n5121 VSS 0.163891f
C10621 DVDD.n5122 VSS 0.096484f
C10622 DVDD.n5123 VSS 0.163891f
C10623 DVDD.n5124 VSS 0.101771f
C10624 DVDD.n5125 VSS 0.163891f
C10625 DVDD.n5126 VSS 0.107058f
C10626 DVDD.n5127 VSS 0.163891f
C10627 DVDD.n5128 VSS 0.112345f
C10628 DVDD.n5129 VSS 0.123789f
C10629 DVDD.n5131 VSS 0.137328f
C10630 DVDD.n5132 VSS 0.137328f
C10631 DVDD.n5133 VSS 0.121855f
C10632 DVDD.n5134 VSS 0.137328f
C10633 DVDD.n5135 VSS 0.137328f
C10634 DVDD.n5136 VSS 0.137328f
C10635 DVDD.n5137 VSS 0.137328f
C10636 DVDD.n5138 VSS 0.137328f
C10637 DVDD.n5139 VSS 0.135394f
C10638 DVDD.n5140 VSS 0.137328f
C10639 DVDD.n5141 VSS 0.137328f
C10640 DVDD.n5142 VSS 0.137328f
C10641 DVDD.n5143 VSS 0.13346f
C10642 DVDD.n5144 VSS 0.11992f
C10643 DVDD.n5145 VSS 0.163891f
C10644 DVDD.n5146 VSS 0.107058f
C10645 DVDD.n5147 VSS 0.163891f
C10646 DVDD.n5148 VSS 0.163891f
C10647 DVDD.n5149 VSS 0.163891f
C10648 DVDD.n5150 VSS 0.107058f
C10649 DVDD.n5151 VSS 0.163891f
C10650 DVDD.n5152 VSS 0.112345f
C10651 DVDD.n5153 VSS 0.163891f
C10652 DVDD.n5154 VSS 0.117632f
C10653 DVDD.n5155 VSS 0.163891f
C10654 DVDD.n5158 VSS 0.270949f
C10655 DVDD.n5159 VSS 0.158604f
C10656 DVDD.n5161 VSS 0.198722f
C10657 DVDD.n5162 VSS 0.081946f
C10658 DVDD.n5163 VSS 0.098809f
C10659 DVDD.t101 VSS 0.167631f
C10660 DVDD.t109 VSS 0.167631f
C10661 DVDD.n5164 VSS 0.335261f
C10662 DVDD.n5165 VSS 0.081946f
C10663 DVDD.n5166 VSS 0.099098f
C10664 DVDD.n5167 VSS 0.198298f
C10665 DVDD.n5168 VSS 0.122918f
C10666 DVDD.n5170 VSS 0.163891f
C10667 DVDD.n5172 VSS 0.198722f
C10668 DVDD.n5173 VSS 0.081946f
C10669 DVDD.n5174 VSS 0.098809f
C10670 DVDD.t93 VSS 0.167631f
C10671 DVDD.t134 VSS 0.167631f
C10672 DVDD.n5175 VSS 0.335261f
C10673 DVDD.n5176 VSS 0.081946f
C10674 DVDD.n5177 VSS 0.099098f
C10675 DVDD.n5178 VSS 0.198298f
C10676 DVDD.n5179 VSS 0.128205f
C10677 DVDD.n5181 VSS 0.163891f
C10678 DVDD.n5183 VSS 0.198722f
C10679 DVDD.n5184 VSS 0.081946f
C10680 DVDD.n5185 VSS 0.098809f
C10681 DVDD.t82 VSS 0.167631f
C10682 DVDD.t125 VSS 0.167631f
C10683 DVDD.n5186 VSS 0.335261f
C10684 DVDD.n5187 VSS 0.081946f
C10685 DVDD.n5188 VSS 0.099098f
C10686 DVDD.n5189 VSS 0.198298f
C10687 DVDD.n5190 VSS 0.133492f
C10688 DVDD.n5192 VSS 0.163891f
C10689 DVDD.n5194 VSS 0.198722f
C10690 DVDD.n5195 VSS 0.081946f
C10691 DVDD.n5196 VSS 0.098809f
C10692 DVDD.t139 VSS 0.425324f
C10693 DVDD.n5197 VSS 0.081946f
C10694 DVDD.n5198 VSS 0.099098f
C10695 DVDD.n5199 VSS 0.198298f
C10696 DVDD.n5200 VSS 0.138779f
C10697 DVDD.n5202 VSS 0.163891f
C10698 DVDD.n5204 VSS 0.163891f
C10699 DVDD.n5206 VSS 0.163891f
C10700 DVDD.n5208 VSS 0.11992f
C10701 DVDD.n5215 VSS 0.274656f
C10702 DVDD.n5216 VSS 0.274656f
C10703 DVDD.n5217 VSS 0.11992f
C10704 DVDD.n5218 VSS 0.274656f
C10705 DVDD.n5219 VSS 0.274656f
C10706 DVDD.n5220 VSS 0.11992f
C10707 DVDD.n5221 VSS 0.274656f
C10708 DVDD.n5222 VSS 0.274656f
C10709 DVDD.n5223 VSS 0.274656f
C10710 DVDD.n5224 VSS 0.274656f
C10711 DVDD.n5225 VSS 0.524168f
C10712 DVDD.n5226 VSS 0.330748f
C10713 DVDD.n5227 VSS 0.274656f
C10714 DVDD.n5228 VSS 0.274656f
C10715 DVDD.n5229 VSS 0.11992f
C10716 DVDD.n5230 VSS 0.06615f
C10717 DVDD.n5231 VSS 0.06615f
C10718 DVDD.n5232 VSS 0.06615f
C10719 DVDD.n5233 VSS 0.06615f
C10720 DVDD.n5234 VSS 0.06615f
C10721 DVDD.n5235 VSS 0.06615f
C10722 DVDD.n5236 VSS 0.06615f
C10723 DVDD.n5237 VSS 0.06615f
C10724 DVDD.n5238 VSS 0.06615f
C10725 DVDD.n5239 VSS 0.06615f
C10726 DVDD.n5240 VSS 0.06615f
C10727 DVDD.n5241 VSS 0.06615f
C10728 DVDD.n5242 VSS 0.06615f
C10729 DVDD.n5243 VSS 0.06615f
C10730 DVDD.n5244 VSS 0.06615f
C10731 DVDD.n5245 VSS 0.06615f
C10732 DVDD.n5246 VSS 0.06615f
C10733 DVDD.n5247 VSS 0.06615f
C10734 DVDD.n5248 VSS 0.06615f
C10735 DVDD.n5249 VSS 0.06615f
C10736 DVDD.n5250 VSS 0.06615f
C10737 DVDD.n5251 VSS 0.06615f
C10738 DVDD.n5252 VSS 0.06615f
C10739 DVDD.n5253 VSS 0.075949f
C10740 DVDD.n5254 VSS 0.128624f
C10741 DVDD.n5255 VSS 0.137328f
C10742 DVDD.n5256 VSS 0.137328f
C10743 DVDD.n5257 VSS 0.137328f
C10744 DVDD.n5258 VSS 0.12669f
C10745 DVDD.n5259 VSS 0.137328f
C10746 DVDD.n5260 VSS 0.137328f
C10747 DVDD.n5261 VSS 0.132299f
C10748 DVDD.n5262 VSS 0.025624f
C10749 DVDD.n5263 VSS 0.0686f
C10750 DVDD.n5264 VSS 0.0735f
C10751 DVDD.n5265 VSS 0.025624f
C10752 DVDD.n5266 VSS 0.075949f
C10753 DVDD.n5267 VSS 0.025624f
C10754 DVDD.n5268 VSS 0.075949f
C10755 DVDD.n5269 VSS 0.025624f
C10756 DVDD.n5270 VSS 0.075949f
C10757 DVDD.n5271 VSS 0.025624f
C10758 DVDD.n5272 VSS 0.075949f
C10759 DVDD.n5273 VSS 0.025624f
C10760 DVDD.n5274 VSS 0.075949f
C10761 DVDD.n5275 VSS 0.025624f
C10762 DVDD.n5276 VSS 0.075949f
C10763 DVDD.n5277 VSS 0.025624f
C10764 DVDD.n5278 VSS 0.025624f
C10765 DVDD.n5279 VSS 0.075949f
C10766 DVDD.n5280 VSS 0.025624f
C10767 DVDD.n5281 VSS 0.075949f
C10768 DVDD.n5282 VSS 0.025624f
C10769 DVDD.n5283 VSS 0.075949f
C10770 DVDD.n5284 VSS 0.025624f
C10771 DVDD.n5285 VSS 0.075949f
C10772 DVDD.n5286 VSS 0.025624f
C10773 DVDD.n5287 VSS 0.075949f
C10774 DVDD.n5288 VSS 0.025624f
C10775 DVDD.n5289 VSS 0.075949f
C10776 DVDD.n5290 VSS 0.025624f
C10777 DVDD.n5291 VSS 0.025624f
C10778 DVDD.n5292 VSS 0.0735f
C10779 DVDD.n5293 VSS 0.0686f
C10780 DVDD.n5294 VSS 0.025624f
C10781 DVDD.n5295 VSS 0.075949f
C10782 DVDD.n5296 VSS 0.025624f
C10783 DVDD.n5297 VSS 0.075949f
C10784 DVDD.n5298 VSS 0.025624f
C10785 DVDD.n5299 VSS 0.075949f
C10786 DVDD.n5300 VSS 0.025624f
C10787 DVDD.n5301 VSS 0.075949f
C10788 DVDD.n5302 VSS 0.025624f
C10789 DVDD.n5303 VSS 0.075949f
C10790 DVDD.n5304 VSS 0.025624f
C10791 DVDD.n5305 VSS 0.075949f
C10792 DVDD.n5306 VSS 0.025624f
C10793 DVDD.n5307 VSS 0.025624f
C10794 DVDD.n5308 VSS 0.07105f
C10795 DVDD.n5309 VSS 0.07105f
C10796 DVDD.n5310 VSS 0.025624f
C10797 DVDD.n5311 VSS 0.025624f
C10798 DVDD.n5312 VSS 0.025624f
C10799 DVDD.n5313 VSS 0.025624f
C10800 DVDD.n5314 VSS 0.132299f
C10801 DVDD.n5315 VSS 0.095549f
C10802 DVDD.n5316 VSS 0.025624f
C10803 DVDD.n5317 VSS 0.075949f
C10804 DVDD.n5318 VSS 0.025624f
C10805 DVDD.n5319 VSS 0.075949f
C10806 DVDD.n5320 VSS 0.025624f
C10807 DVDD.n5321 VSS 0.075949f
C10808 DVDD.n5322 VSS 0.025624f
C10809 DVDD.n5323 VSS 0.025624f
C10810 DVDD.n5324 VSS 0.0735f
C10811 DVDD.n5325 VSS 0.0686f
C10812 DVDD.n5326 VSS 0.025624f
C10813 DVDD.n5327 VSS 0.075949f
C10814 DVDD.n5328 VSS 0.025624f
C10815 DVDD.n5329 VSS 0.075949f
C10816 DVDD.n5330 VSS 0.025624f
C10817 DVDD.n5331 VSS 0.075949f
C10818 DVDD.n5332 VSS 0.025624f
C10819 DVDD.n5333 VSS 0.075949f
C10820 DVDD.n5334 VSS 0.025624f
C10821 DVDD.n5335 VSS 0.075949f
C10822 DVDD.n5336 VSS 0.025624f
C10823 DVDD.n5337 VSS 0.075949f
C10824 DVDD.n5338 VSS 0.025624f
C10825 DVDD.n5339 VSS 0.025624f
C10826 DVDD.n5340 VSS 0.07105f
C10827 DVDD.n5341 VSS 0.07105f
C10828 DVDD.n5342 VSS 0.025624f
C10829 DVDD.n5343 VSS 0.075949f
C10830 DVDD.n5344 VSS 0.025624f
C10831 DVDD.n5345 VSS 0.075949f
C10832 DVDD.n5346 VSS 0.025624f
C10833 DVDD.n5347 VSS 0.075949f
C10834 DVDD.n5348 VSS 0.025624f
C10835 DVDD.n5349 VSS 0.075949f
C10836 DVDD.n5350 VSS 0.025624f
C10837 DVDD.n5351 VSS 0.075949f
C10838 DVDD.n5352 VSS 0.025624f
C10839 DVDD.n5353 VSS 0.075949f
C10840 DVDD.n5354 VSS 0.025624f
C10841 DVDD.n5355 VSS 0.025624f
C10842 DVDD.n5356 VSS 0.0686f
C10843 DVDD.n5357 VSS 0.0735f
C10844 DVDD.n5358 VSS 0.025624f
C10845 DVDD.n5359 VSS 0.075949f
C10846 DVDD.n5360 VSS 0.025624f
C10847 DVDD.n5361 VSS 0.075949f
C10848 DVDD.n5362 VSS 0.025624f
C10849 DVDD.n5363 VSS 0.075949f
C10850 DVDD.n5364 VSS 0.025624f
C10851 DVDD.n5365 VSS 0.075949f
C10852 DVDD.n5366 VSS 0.025624f
C10853 DVDD.n5367 VSS 0.025624f
C10854 DVDD.n5368 VSS 0.025624f
C10855 DVDD.n5369 VSS 0.137328f
C10856 DVDD.n5370 VSS 0.137328f
C10857 DVDD.n5372 VSS 0.137328f
C10858 DVDD.n5374 VSS 0.137328f
C10859 DVDD.n5375 VSS 0.137328f
C10860 DVDD.n5376 VSS 0.075949f
C10861 DVDD.n5377 VSS 0.137328f
C10862 DVDD.n5378 VSS 0.137328f
C10863 DVDD.n5379 VSS 0.803653f
C10864 DVDD.n5380 VSS 0.137328f
C10865 DVDD.n5381 VSS 0.137328f
C10866 DVDD.n5382 VSS 0.11992f
C10867 DVDD.n5383 VSS 0.06615f
C10868 DVDD.n5384 VSS 0.06615f
C10869 DVDD.n5385 VSS 0.06615f
C10870 DVDD.n5386 VSS 0.06615f
C10871 DVDD.n5387 VSS 0.06615f
C10872 DVDD.n5388 VSS 0.06615f
C10873 DVDD.n5389 VSS 0.06615f
C10874 DVDD.n5390 VSS 0.06615f
C10875 DVDD.n5391 VSS 0.06615f
C10876 DVDD.n5392 VSS 0.06615f
C10877 DVDD.n5393 VSS 0.06615f
C10878 DVDD.n5394 VSS 0.217597f
C10879 DVDD.n5395 VSS 0.06615f
C10880 DVDD.n5396 VSS 0.06615f
C10881 DVDD.n5397 VSS 0.06615f
C10882 DVDD.n5398 VSS 0.06615f
C10883 DVDD.n5399 VSS 0.06615f
C10884 DVDD.n5400 VSS 0.06615f
C10885 DVDD.n5401 VSS 0.132299f
C10886 DVDD.n5402 VSS 0.06615f
C10887 DVDD.n5403 VSS 0.06615f
C10888 DVDD.n5404 VSS 0.06615f
C10889 DVDD.n5405 VSS 0.06615f
C10890 DVDD.n5406 VSS 0.075949f
C10891 DVDD.n5407 VSS 0.12669f
C10892 DVDD.n5408 VSS 0.128624f
C10893 DVDD.n5409 VSS 0.132299f
C10894 DVDD.n5410 VSS 0.025624f
C10895 DVDD.n5411 VSS 0.075949f
C10896 DVDD.n5412 VSS 0.025624f
C10897 DVDD.n5413 VSS 0.075949f
C10898 DVDD.n5414 VSS 0.025624f
C10899 DVDD.n5415 VSS 0.075949f
C10900 DVDD.n5416 VSS 0.025624f
C10901 DVDD.n5417 VSS 0.075949f
C10902 DVDD.n5418 VSS 0.025624f
C10903 DVDD.n5419 VSS 0.075949f
C10904 DVDD.n5420 VSS 0.025624f
C10905 DVDD.n5421 VSS 0.025624f
C10906 DVDD.n5422 VSS 0.0686f
C10907 DVDD.n5423 VSS 0.0735f
C10908 DVDD.n5424 VSS 0.025624f
C10909 DVDD.n5425 VSS 0.075949f
C10910 DVDD.n5426 VSS 0.025624f
C10911 DVDD.n5427 VSS 0.075949f
C10912 DVDD.n5428 VSS 0.025624f
C10913 DVDD.n5429 VSS 0.075949f
C10914 DVDD.n5430 VSS 0.025624f
C10915 DVDD.n5431 VSS 0.075949f
C10916 DVDD.n5432 VSS 0.025624f
C10917 DVDD.n5433 VSS 0.075949f
C10918 DVDD.n5434 VSS 0.025624f
C10919 DVDD.n5435 VSS 0.075949f
C10920 DVDD.n5436 VSS 0.025624f
C10921 DVDD.n5437 VSS 0.025624f
C10922 DVDD.n5438 VSS 0.075949f
C10923 DVDD.n5439 VSS 0.025624f
C10924 DVDD.n5440 VSS 0.075949f
C10925 DVDD.n5441 VSS 0.025624f
C10926 DVDD.n5442 VSS 0.075949f
C10927 DVDD.n5443 VSS 0.025624f
C10928 DVDD.n5444 VSS 0.075949f
C10929 DVDD.n5445 VSS 0.025624f
C10930 DVDD.n5446 VSS 0.075949f
C10931 DVDD.n5447 VSS 0.025624f
C10932 DVDD.n5448 VSS 0.075949f
C10933 DVDD.n5449 VSS 0.025624f
C10934 DVDD.n5450 VSS 0.025624f
C10935 DVDD.n5451 VSS 0.0735f
C10936 DVDD.n5452 VSS 0.0686f
C10937 DVDD.n5453 VSS 0.025624f
C10938 DVDD.n5454 VSS 0.075949f
C10939 DVDD.n5455 VSS 0.025624f
C10940 DVDD.n5456 VSS 0.075949f
C10941 DVDD.n5457 VSS 0.025624f
C10942 DVDD.n5458 VSS 0.025624f
C10943 DVDD.n5459 VSS 0.025624f
C10944 DVDD.n5460 VSS 0.132299f
C10945 DVDD.n5461 VSS 0.025624f
C10946 DVDD.n5462 VSS 0.132299f
C10947 DVDD.n5463 VSS 0.025624f
C10948 DVDD.n5464 VSS 0.132299f
C10949 DVDD.n5465 VSS 0.025624f
C10950 DVDD.n5466 VSS 0.104124f
C10951 DVDD.n5467 VSS 0.025624f
C10952 DVDD.n5468 VSS 0.06615f
C10953 DVDD.n5469 VSS 0.060025f
C10954 DVDD.n5470 VSS 0.064086f
C10955 DVDD.n5471 VSS 0.064086f
C10956 DVDD.n5472 VSS 0.064086f
C10957 DVDD.n5473 VSS 0.059122f
C10958 DVDD.n5474 VSS 0.064086f
C10959 DVDD.n5475 VSS 0.064086f
C10960 DVDD.n5476 VSS 0.075949f
C10961 DVDD.n5477 VSS 0.064086f
C10962 DVDD.n5478 VSS 0.064086f
C10963 DVDD.n5480 VSS 0.060927f
C10964 DVDD.n5481 VSS 0.064086f
C10965 DVDD.n5482 VSS 0.064086f
C10966 DVDD.n5483 VSS 0.064086f
C10967 DVDD.n5485 VSS 0.060025f
C10968 DVDD.n5486 VSS 0.353402f
C10969 DVDD.n5487 VSS 0.06615f
C10970 DVDD.n5488 VSS 0.06615f
C10971 DVDD.n5489 VSS 0.06615f
C10972 DVDD.n5490 VSS 0.06615f
C10973 DVDD.n5491 VSS 0.055963f
C10974 DVDD.n5492 VSS 0.06615f
C10975 DVDD.n5493 VSS 0.06615f
C10976 DVDD.n5494 VSS 0.06615f
C10977 DVDD.n5495 VSS 0.06615f
C10978 DVDD.n5496 VSS 0.069825f
C10979 DVDD.n5497 VSS 0.132299f
C10980 DVDD.n5498 VSS 0.025624f
C10981 DVDD.n5499 VSS 0.074725f
C10982 DVDD.n5500 VSS 0.067375f
C10983 DVDD.n5501 VSS 0.025624f
C10984 DVDD.n5502 VSS 0.075949f
C10985 DVDD.n5503 VSS 0.025624f
C10986 DVDD.n5504 VSS 0.075949f
C10987 DVDD.n5505 VSS 0.025624f
C10988 DVDD.n5506 VSS 0.075949f
C10989 DVDD.n5507 VSS 0.025624f
C10990 DVDD.n5508 VSS 0.075949f
C10991 DVDD.n5509 VSS 0.025624f
C10992 DVDD.n5510 VSS 0.075949f
C10993 DVDD.n5511 VSS 0.025624f
C10994 DVDD.n5512 VSS 0.075949f
C10995 DVDD.n5513 VSS 0.025624f
C10996 DVDD.n5514 VSS 0.072275f
C10997 DVDD.n5515 VSS 0.025624f
C10998 DVDD.n5516 VSS 0.025624f
C10999 DVDD.n5517 VSS 0.025624f
C11000 DVDD.n5518 VSS 0.132299f
C11001 DVDD.n5519 VSS 0.025624f
C11002 DVDD.n5520 VSS 0.132299f
C11003 DVDD.n5521 VSS 0.025624f
C11004 DVDD.n5522 VSS 0.132299f
C11005 DVDD.n5523 VSS 0.025624f
C11006 DVDD.n5524 VSS 0.132299f
C11007 DVDD.n5525 VSS 0.025624f
C11008 DVDD.n5526 VSS 0.132299f
C11009 DVDD.n5527 VSS 0.025624f
C11010 DVDD.n5528 VSS 0.132299f
C11011 DVDD.n5529 VSS 0.025624f
C11012 DVDD.n5530 VSS 0.132299f
C11013 DVDD.n5531 VSS 0.025624f
C11014 DVDD.n5532 VSS 0.132299f
C11015 DVDD.n5533 VSS 0.025624f
C11016 DVDD.n5534 VSS 0.132299f
C11017 DVDD.n5535 VSS 0.025624f
C11018 DVDD.n5536 VSS 0.132299f
C11019 DVDD.n5537 VSS 0.025624f
C11020 DVDD.n5538 VSS 0.132299f
C11021 DVDD.n5539 VSS 0.025624f
C11022 DVDD.n5540 VSS 0.132299f
C11023 DVDD.n5541 VSS 0.025624f
C11024 DVDD.n5542 VSS 0.132299f
C11025 DVDD.n5543 VSS 0.025624f
C11026 DVDD.n5544 VSS 0.132299f
C11027 DVDD.n5545 VSS 0.025624f
C11028 DVDD.n5546 VSS 0.132299f
C11029 DVDD.n5547 VSS 0.025624f
C11030 DVDD.n5548 VSS 0.132299f
C11031 DVDD.n5549 VSS 0.025624f
C11032 DVDD.n5550 VSS 0.132299f
C11033 DVDD.n5551 VSS 0.025624f
C11034 DVDD.n5552 VSS 0.132299f
C11035 DVDD.n5553 VSS 0.025624f
C11036 DVDD.n5554 VSS 0.132299f
C11037 DVDD.n5555 VSS 0.025624f
C11038 DVDD.n5556 VSS 0.132299f
C11039 DVDD.n5557 VSS 0.025624f
C11040 DVDD.n5558 VSS 0.132299f
C11041 DVDD.n5559 VSS 0.025624f
C11042 DVDD.n5560 VSS 0.117599f
C11043 DVDD.n5563 VSS 0.06615f
C11044 DVDD.n5564 VSS 0.06615f
C11045 DVDD.n5565 VSS 0.030844f
C11046 DVDD.n5566 VSS 0.06615f
C11047 DVDD.n5568 VSS 0.098464f
C11048 DVDD.n5570 VSS 0.025624f
C11049 DVDD.n5572 VSS 0.025624f
C11050 DVDD.n5574 VSS 0.025624f
C11051 DVDD.n5575 VSS 0.025624f
C11052 DVDD.n5577 VSS 0.026154f
C11053 DVDD.n5578 VSS 0.036879f
C11054 DVDD.n5580 VSS 0.059058f
C11055 DVDD.n5582 VSS 0.053165f
C11056 DVDD.n5583 VSS 0.088457f
C11057 DVDD.n5584 VSS 0.088457f
C11058 DVDD.n5586 VSS 0.053165f
C11059 DVDD.n5587 VSS 0.106252f
C11060 DVDD.n5588 VSS 0.063957f
C11061 DVDD.n5589 VSS 0.063957f
C11062 DVDD.n5592 VSS 0.522253f
C11063 DVDD.n5593 VSS 0.522253f
C11064 DVDD.n5594 VSS 0.063957f
C11065 DVDD.n5595 VSS 0.063957f
C11066 DVDD.n5596 VSS 0.063957f
C11067 DVDD.n5597 VSS 0.063957f
C11068 DVDD.n5598 VSS 0.063957f
C11069 DVDD.n5599 VSS 0.063957f
C11070 DVDD.n5600 VSS 0.063957f
C11071 DVDD.n5601 VSS 0.063957f
C11072 DVDD.n5602 VSS 0.063957f
C11073 DVDD.n5603 VSS 0.063957f
C11074 DVDD.n5604 VSS 0.063957f
C11075 DVDD.n5605 VSS 0.063957f
C11076 DVDD.n5606 VSS 0.063957f
C11077 DVDD.n5607 VSS 0.063957f
C11078 DVDD.n5608 VSS 0.063957f
C11079 DVDD.n5609 VSS 0.063957f
C11080 DVDD.n5610 VSS 0.063957f
C11081 DVDD.n5611 VSS 0.063957f
C11082 DVDD.n5612 VSS 0.063957f
C11083 DVDD.n5613 VSS 0.063957f
C11084 DVDD.n5614 VSS 0.063957f
C11085 DVDD.n5615 VSS 0.063957f
C11086 DVDD.n5616 VSS 0.063957f
C11087 DVDD.n5617 VSS 0.063957f
C11088 DVDD.n5618 VSS 0.063957f
C11089 DVDD.n5619 VSS 0.063957f
C11090 DVDD.n5620 VSS 0.063957f
C11091 DVDD.n5621 VSS 0.063957f
C11092 DVDD.n5622 VSS 0.063957f
C11093 DVDD.n5623 VSS 0.063957f
C11094 DVDD.n5624 VSS 0.063957f
C11095 DVDD.n5625 VSS 0.063957f
C11096 DVDD.n5626 VSS 0.063957f
C11097 DVDD.n5627 VSS 0.063957f
C11098 DVDD.n5628 VSS 0.063957f
C11099 DVDD.n5629 VSS 0.063957f
C11100 DVDD.n5630 VSS 0.063957f
C11101 DVDD.n5631 VSS 0.063957f
C11102 DVDD.n5632 VSS 0.063957f
C11103 DVDD.n5633 VSS 0.063957f
C11104 DVDD.n5634 VSS 0.063957f
C11105 DVDD.n5635 VSS 0.063957f
C11106 DVDD.n5636 VSS 0.063957f
C11107 DVDD.n5637 VSS 0.063957f
C11108 DVDD.n5638 VSS 0.063957f
C11109 DVDD.n5639 VSS 0.063957f
C11110 DVDD.n5640 VSS 0.063957f
C11111 DVDD.n5641 VSS 0.063957f
C11112 DVDD.n5642 VSS 0.522253f
C11113 DVDD.n5643 VSS 0.104963f
C11114 DVDD.n5644 VSS 0.088457f
C11115 DVDD.n5645 VSS 0.063957f
C11116 DVDD.n5646 VSS 0.063957f
C11117 DVDD.n5647 VSS 0.063957f
C11118 DVDD.n5648 VSS 0.063957f
C11119 DVDD.n5649 VSS 0.063957f
C11120 DVDD.n5650 VSS 0.063957f
C11121 DVDD.n5651 VSS 0.063957f
C11122 DVDD.n5652 VSS 0.063957f
C11123 DVDD.n5653 VSS 0.063957f
C11124 DVDD.n5654 VSS 0.063957f
C11125 DVDD.n5655 VSS 0.063957f
C11126 DVDD.n5656 VSS 0.063957f
C11127 DVDD.n5657 VSS 0.063957f
C11128 DVDD.n5658 VSS 0.063957f
C11129 DVDD.n5659 VSS 0.063957f
C11130 DVDD.n5660 VSS 0.063957f
C11131 DVDD.n5661 VSS 0.063957f
C11132 DVDD.n5662 VSS 0.063957f
C11133 DVDD.n5663 VSS 0.063957f
C11134 DVDD.n5664 VSS 0.063957f
C11135 DVDD.n5665 VSS 0.063957f
C11136 DVDD.n5666 VSS 0.063957f
C11137 DVDD.n5667 VSS 0.063957f
C11138 DVDD.n5668 VSS 0.063957f
C11139 DVDD.n5669 VSS 0.063957f
C11140 DVDD.n5670 VSS 0.063957f
C11141 DVDD.n5671 VSS 0.063957f
C11142 DVDD.n5672 VSS 0.063957f
C11143 DVDD.n5673 VSS 0.063957f
C11144 DVDD.n5674 VSS 0.063957f
C11145 DVDD.n5675 VSS 0.063957f
C11146 DVDD.n5676 VSS 0.063957f
C11147 DVDD.n5677 VSS 0.063957f
C11148 DVDD.n5678 VSS 0.063957f
C11149 DVDD.n5679 VSS 0.063957f
C11150 DVDD.n5680 VSS 0.063957f
C11151 DVDD.n5681 VSS 0.063957f
C11152 DVDD.n5682 VSS 0.063957f
C11153 DVDD.n5683 VSS 0.063957f
C11154 DVDD.n5684 VSS 0.063957f
C11155 DVDD.n5685 VSS 0.063957f
C11156 DVDD.n5686 VSS 0.063957f
C11157 DVDD.n5687 VSS 0.063957f
C11158 DVDD.n5688 VSS 0.063957f
C11159 DVDD.n5689 VSS 0.063957f
C11160 DVDD.n5690 VSS 0.063957f
C11161 DVDD.n5691 VSS 0.063957f
C11162 DVDD.n5740 VSS 0.522253f
C11163 DVDD.n5741 VSS 0.03626f
C11164 DVDD.n5742 VSS 0.063957f
C11165 DVDD.n5743 VSS 0.03626f
C11166 DVDD.n5744 VSS 0.063957f
C11167 DVDD.n5745 VSS 0.063957f
C11168 DVDD.n5746 VSS 0.063957f
C11169 DVDD.n5747 VSS 0.063957f
C11170 DVDD.n5748 VSS 0.063957f
C11171 DVDD.n5749 VSS 0.063957f
C11172 DVDD.n5750 VSS 0.063957f
C11173 DVDD.n5751 VSS 0.063957f
C11174 DVDD.n5752 VSS 0.063957f
C11175 DVDD.n5753 VSS 0.063957f
C11176 DVDD.n5754 VSS 0.063957f
C11177 DVDD.n5755 VSS 0.063957f
C11178 DVDD.n5756 VSS 0.063957f
C11179 DVDD.n5757 VSS 0.063957f
C11180 DVDD.n5758 VSS 0.063957f
C11181 DVDD.n5759 VSS 0.063957f
C11182 DVDD.n5760 VSS 0.063957f
C11183 DVDD.n5761 VSS 0.063957f
C11184 DVDD.n5762 VSS 0.063957f
C11185 DVDD.n5763 VSS 0.063957f
C11186 DVDD.n5764 VSS 0.063957f
C11187 DVDD.n5765 VSS 0.063957f
C11188 DVDD.n5766 VSS 0.063957f
C11189 DVDD.n5767 VSS 0.063957f
C11190 DVDD.n5768 VSS 0.063957f
C11191 DVDD.n5769 VSS 0.063957f
C11192 DVDD.n5770 VSS 0.063957f
C11193 DVDD.n5771 VSS 0.063957f
C11194 DVDD.n5772 VSS 0.063957f
C11195 DVDD.n5773 VSS 0.063957f
C11196 DVDD.n5774 VSS 0.063957f
C11197 DVDD.n5775 VSS 0.063957f
C11198 DVDD.n5776 VSS 0.063957f
C11199 DVDD.n5777 VSS 0.063957f
C11200 DVDD.n5778 VSS 0.063957f
C11201 DVDD.n5779 VSS 0.063957f
C11202 DVDD.n5780 VSS 0.063957f
C11203 DVDD.n5781 VSS 0.063957f
C11204 DVDD.n5782 VSS 0.063957f
C11205 DVDD.n5783 VSS 0.063957f
C11206 DVDD.n5784 VSS 0.063957f
C11207 DVDD.n5785 VSS 0.063957f
C11208 DVDD.n5786 VSS 0.063957f
C11209 DVDD.n5787 VSS 0.063957f
C11210 DVDD.n5788 VSS 0.063957f
C11211 DVDD.n5789 VSS 0.063957f
C11212 DVDD.n5790 VSS 0.063957f
C11213 DVDD.n5791 VSS 0.063957f
C11214 DVDD.n5792 VSS 0.063957f
C11215 DVDD.n5793 VSS 0.063957f
C11216 DVDD.n5794 VSS 0.063957f
C11217 DVDD.n5795 VSS 0.063957f
C11218 DVDD.n5796 VSS 0.063957f
C11219 DVDD.n5797 VSS 0.063957f
C11220 DVDD.n5798 VSS 0.063957f
C11221 DVDD.n5799 VSS 0.063957f
C11222 DVDD.n5800 VSS 0.063957f
C11223 DVDD.n5801 VSS 0.063957f
C11224 DVDD.n5802 VSS 0.063957f
C11225 DVDD.n5803 VSS 0.063957f
C11226 DVDD.n5804 VSS 0.063957f
C11227 DVDD.n5805 VSS 0.063957f
C11228 DVDD.n5806 VSS 0.063957f
C11229 DVDD.n5807 VSS 0.063957f
C11230 DVDD.n5808 VSS 0.063957f
C11231 DVDD.n5809 VSS 0.063957f
C11232 DVDD.n5810 VSS 0.063957f
C11233 DVDD.n5811 VSS 0.063957f
C11234 DVDD.n5812 VSS 0.063957f
C11235 DVDD.n5813 VSS 0.063957f
C11236 DVDD.n5814 VSS 0.063957f
C11237 DVDD.n5815 VSS 0.063957f
C11238 DVDD.n5816 VSS 0.063957f
C11239 DVDD.n5817 VSS 0.063957f
C11240 DVDD.n5818 VSS 0.063957f
C11241 DVDD.n5819 VSS 0.063957f
C11242 DVDD.n5820 VSS 0.063957f
C11243 DVDD.n5821 VSS 0.063957f
C11244 DVDD.n5822 VSS 0.063957f
C11245 DVDD.n5823 VSS 0.063957f
C11246 DVDD.n5824 VSS 0.063957f
C11247 DVDD.n5825 VSS 0.063957f
C11248 DVDD.n5826 VSS 0.063957f
C11249 DVDD.n5827 VSS 0.063957f
C11250 DVDD.n5828 VSS 0.063957f
C11251 DVDD.n5829 VSS 0.063957f
C11252 DVDD.n5830 VSS 0.063957f
C11253 DVDD.n5831 VSS 0.063957f
C11254 DVDD.n5832 VSS 0.063957f
C11255 DVDD.n5833 VSS 0.063957f
C11256 DVDD.n5834 VSS 0.063957f
C11257 DVDD.n5835 VSS 0.063957f
C11258 DVDD.n5836 VSS 0.063957f
C11259 DVDD.n5837 VSS 0.063957f
C11260 DVDD.n5838 VSS 0.063957f
C11261 DVDD.n5839 VSS 0.063957f
C11262 DVDD.n5840 VSS 0.063957f
C11263 DVDD.n5841 VSS 0.063957f
C11264 DVDD.n5842 VSS 0.063957f
C11265 DVDD.n5843 VSS 0.063957f
C11266 DVDD.n5844 VSS 0.063957f
C11267 DVDD.n5845 VSS 0.063957f
C11268 DVDD.n5846 VSS 0.063957f
C11269 DVDD.n5847 VSS 0.063957f
C11270 DVDD.n5848 VSS 0.063957f
C11271 DVDD.n5849 VSS 0.063957f
C11272 DVDD.n5850 VSS 0.063957f
C11273 DVDD.n5851 VSS 0.063957f
C11274 DVDD.n5852 VSS 0.063957f
C11275 DVDD.n5853 VSS 0.063957f
C11276 DVDD.n5854 VSS 0.063957f
C11277 DVDD.n5855 VSS 0.063957f
C11278 DVDD.n5856 VSS 0.063957f
C11279 DVDD.n5857 VSS 0.063957f
C11280 DVDD.n5858 VSS 0.063957f
C11281 DVDD.n5859 VSS 0.063957f
C11282 DVDD.n5860 VSS 0.063957f
C11283 DVDD.n5861 VSS 0.063957f
C11284 DVDD.n5862 VSS 0.063957f
C11285 DVDD.n5863 VSS 0.063957f
C11286 DVDD.n5864 VSS 0.063957f
C11287 DVDD.n5865 VSS 0.063957f
C11288 DVDD.n5866 VSS 0.063957f
C11289 DVDD.n5867 VSS 0.063957f
C11290 DVDD.n5868 VSS 0.063957f
C11291 DVDD.n5869 VSS 0.063957f
C11292 DVDD.n5870 VSS 0.063957f
C11293 DVDD.n5871 VSS 0.063957f
C11294 DVDD.n5872 VSS 0.063957f
C11295 DVDD.n5873 VSS 0.063957f
C11296 DVDD.n5874 VSS 0.063957f
C11297 DVDD.n5875 VSS 0.063957f
C11298 DVDD.n5876 VSS 0.063957f
C11299 DVDD.n5877 VSS 0.063957f
C11300 DVDD.n5878 VSS 0.063957f
C11301 DVDD.n5879 VSS 0.063957f
C11302 DVDD.n5880 VSS 0.063957f
C11303 DVDD.n5881 VSS 0.063957f
C11304 DVDD.n5882 VSS 0.063957f
C11305 DVDD.n5883 VSS 0.063957f
C11306 DVDD.n5884 VSS 0.063957f
C11307 DVDD.n5885 VSS 0.063957f
C11308 DVDD.n5886 VSS 0.063957f
C11309 DVDD.n5887 VSS 0.063957f
C11310 DVDD.n5888 VSS 0.063957f
C11311 DVDD.n5889 VSS 0.063957f
C11312 DVDD.n5890 VSS 0.063957f
C11313 DVDD.n5891 VSS 0.063957f
C11314 DVDD.n5892 VSS 0.063957f
C11315 DVDD.n5893 VSS 0.063957f
C11316 DVDD.n5894 VSS 0.063957f
C11317 DVDD.n5895 VSS 0.063957f
C11318 DVDD.n5896 VSS 0.063957f
C11319 DVDD.n5897 VSS 0.063957f
C11320 DVDD.n5898 VSS 0.063957f
C11321 DVDD.n5899 VSS 0.063957f
C11322 DVDD.n5900 VSS 0.063957f
C11323 DVDD.n5901 VSS 0.063957f
C11324 DVDD.n5902 VSS 0.063957f
C11325 DVDD.n5903 VSS 0.063957f
C11326 DVDD.n5904 VSS 0.063957f
C11327 DVDD.n5905 VSS 0.063957f
C11328 DVDD.n5906 VSS 0.063957f
C11329 DVDD.n5907 VSS 0.063957f
C11330 DVDD.n5908 VSS 0.063957f
C11331 DVDD.n5909 VSS 0.063957f
C11332 DVDD.n5910 VSS 0.063957f
C11333 DVDD.n5911 VSS 0.063957f
C11334 DVDD.n5912 VSS 0.063957f
C11335 DVDD.n5913 VSS 0.063957f
C11336 DVDD.n5914 VSS 0.063957f
C11337 DVDD.n5915 VSS 0.063957f
C11338 DVDD.n5916 VSS 0.063957f
C11339 DVDD.n5917 VSS 0.063957f
C11340 DVDD.n5918 VSS 0.063957f
C11341 DVDD.n5919 VSS 0.063957f
C11342 DVDD.n5920 VSS 0.063957f
C11343 DVDD.n5921 VSS 0.063957f
C11344 DVDD.n5922 VSS 0.063957f
C11345 DVDD.n5923 VSS 0.063957f
C11346 DVDD.n5924 VSS 0.063957f
C11347 DVDD.n5925 VSS 0.063957f
C11348 DVDD.n5926 VSS 0.063957f
C11349 DVDD.n5927 VSS 0.063957f
C11350 DVDD.n5928 VSS 0.063957f
C11351 DVDD.n5929 VSS 0.063957f
C11352 DVDD.n5930 VSS 0.063957f
C11353 DVDD.n5931 VSS 0.036621f
C11354 DVDD.n5932 VSS 0.041931f
C11355 DVDD.n5933 VSS 0.041931f
C11356 DVDD.n5934 VSS 0.73705f
C11357 DVDD.n5935 VSS 0.522252f
C11358 DVDD.n5936 VSS 0.059058f
C11359 DVDD.n5938 VSS 0.522253f
C11360 DVDD.n5986 VSS 0.522253f
C11361 DVDD.n5987 VSS 0.522253f
C11362 DVDD.n5988 VSS 0.555947f
C11363 DVDD.n5990 VSS 0.106252f
C11364 DVDD.n5991 VSS 0.522253f
C11365 DVDD.n5992 VSS 0.036879f
C11366 DVDD.n5993 VSS 0.056475f
C11367 DVDD.n5994 VSS 0.05956f
C11368 DVDD.n5995 VSS 0.056475f
C11369 DVDD.n5996 VSS 0.05956f
C11370 DVDD.n5997 VSS 0.039516f
C11371 DVDD.n5998 VSS 0.033945f
C11372 DVDD.n5999 VSS 0.033945f
C11373 DVDD.n6000 VSS 0.256914f
C11374 DVDD.n6042 VSS 0.019729f
C11375 DVDD.n6043 VSS 0.181104f
C11376 DVDD.n6044 VSS 0.02513f
C11377 DVDD.n6046 VSS 0.031128f
C11378 DVDD.n6047 VSS 0.031128f
C11379 DVDD.n6048 VSS 0.031128f
C11380 DVDD.n6049 VSS 0.031128f
C11381 DVDD.n6050 VSS 0.031128f
C11382 DVDD.n6051 VSS 0.496982f
C11383 DVDD.n6091 VSS 0.019729f
C11384 DVDD.n6092 VSS 0.031128f
C11385 DVDD.n6093 VSS 0.031128f
C11386 DVDD.n6094 VSS 0.028497f
C11387 DVDD.n6095 VSS 0.031128f
C11388 DVDD.n6096 VSS 0.031128f
C11389 DVDD.n6097 VSS 0.031128f
C11390 DVDD.n6098 VSS 0.031128f
C11391 DVDD.n6099 VSS 0.031128f
C11392 DVDD.n6100 VSS 0.031128f
C11393 DVDD.n6101 VSS 0.031128f
C11394 DVDD.n6102 VSS 0.031128f
C11395 DVDD.n6103 VSS 0.031128f
C11396 DVDD.n6104 VSS 0.031128f
C11397 DVDD.n6105 VSS 0.031128f
C11398 DVDD.n6106 VSS 0.031128f
C11399 DVDD.n6107 VSS 0.031128f
C11400 DVDD.n6108 VSS 0.031128f
C11401 DVDD.n6109 VSS 0.031128f
C11402 DVDD.n6110 VSS 0.031128f
C11403 DVDD.n6111 VSS 0.031128f
C11404 DVDD.n6112 VSS 0.031128f
C11405 DVDD.n6113 VSS 0.031128f
C11406 DVDD.n6114 VSS 0.031128f
C11407 DVDD.n6115 VSS 0.031128f
C11408 DVDD.n6116 VSS 0.031128f
C11409 DVDD.n6117 VSS 0.031128f
C11410 DVDD.n6118 VSS 0.031128f
C11411 DVDD.n6119 VSS 0.031128f
C11412 DVDD.n6120 VSS 0.031128f
C11413 DVDD.n6121 VSS 0.031128f
C11414 DVDD.n6122 VSS 0.031128f
C11415 DVDD.n6123 VSS 0.031128f
C11416 DVDD.n6124 VSS 0.031128f
C11417 DVDD.n6125 VSS 0.031128f
C11418 DVDD.n6126 VSS 0.031128f
C11419 DVDD.n6127 VSS 0.031128f
C11420 DVDD.n6128 VSS 0.031128f
C11421 DVDD.n6129 VSS 0.031128f
C11422 DVDD.n6130 VSS 0.031128f
C11423 DVDD.n6131 VSS 0.031128f
C11424 DVDD.n6132 VSS 0.031128f
C11425 DVDD.n6133 VSS 0.031128f
C11426 DVDD.n6134 VSS 0.031128f
C11427 DVDD.n6135 VSS 0.031128f
C11428 DVDD.n6136 VSS 0.031128f
C11429 DVDD.n6137 VSS 0.031128f
C11430 DVDD.n6138 VSS 0.031128f
C11431 DVDD.n6139 VSS 0.031128f
C11432 DVDD.n6140 VSS 0.031128f
C11433 DVDD.n6141 VSS 0.031128f
C11434 DVDD.n6142 VSS 0.031128f
C11435 DVDD.n6143 VSS 0.031128f
C11436 DVDD.n6144 VSS 0.031128f
C11437 DVDD.n6145 VSS 0.031128f
C11438 DVDD.n6146 VSS 0.031128f
C11439 DVDD.n6147 VSS 0.031128f
C11440 DVDD.n6148 VSS 0.031128f
C11441 DVDD.n6149 VSS 0.031128f
C11442 DVDD.n6150 VSS 0.031128f
C11443 DVDD.n6151 VSS 0.031128f
C11444 DVDD.n6152 VSS 0.031128f
C11445 DVDD.n6153 VSS 0.031128f
C11446 DVDD.n6154 VSS 0.031128f
C11447 DVDD.n6155 VSS 0.031128f
C11448 DVDD.n6156 VSS 0.031128f
C11449 DVDD.n6157 VSS 0.031128f
C11450 DVDD.n6158 VSS 0.031128f
C11451 DVDD.n6159 VSS 0.031128f
C11452 DVDD.n6160 VSS 0.031128f
C11453 DVDD.n6161 VSS 0.031128f
C11454 DVDD.n6162 VSS 0.031128f
C11455 DVDD.n6163 VSS 0.031128f
C11456 DVDD.n6164 VSS 0.031128f
C11457 DVDD.n6165 VSS 0.031128f
C11458 DVDD.n6166 VSS 0.031128f
C11459 DVDD.n6167 VSS 0.031128f
C11460 DVDD.n6168 VSS 0.031128f
C11461 DVDD.n6169 VSS 0.031128f
C11462 DVDD.n6170 VSS 0.031128f
C11463 DVDD.n6171 VSS 0.031128f
C11464 DVDD.n6172 VSS 0.031128f
C11465 DVDD.n6173 VSS 0.031128f
C11466 DVDD.n6174 VSS 0.031128f
C11467 DVDD.n6175 VSS 0.031128f
C11468 DVDD.n6176 VSS 0.031128f
C11469 DVDD.n6177 VSS 0.031128f
C11470 DVDD.n6178 VSS 0.031128f
C11471 DVDD.n6179 VSS 0.031128f
C11472 DVDD.n6180 VSS 0.031128f
C11473 DVDD.n6181 VSS 0.031128f
C11474 DVDD.n6182 VSS 0.031128f
C11475 DVDD.n6183 VSS 0.031128f
C11476 DVDD.n6184 VSS 0.031128f
C11477 DVDD.n6185 VSS 0.031128f
C11478 DVDD.n6186 VSS 0.031128f
C11479 DVDD.n6187 VSS 0.031128f
C11480 DVDD.n6188 VSS 0.031128f
C11481 DVDD.n6189 VSS 0.031128f
C11482 DVDD.n6190 VSS 0.031128f
C11483 DVDD.n6191 VSS 0.031128f
C11484 DVDD.n6192 VSS 0.031128f
C11485 DVDD.n6193 VSS 0.031128f
C11486 DVDD.n6194 VSS 0.031128f
C11487 DVDD.n6195 VSS 0.031128f
C11488 DVDD.n6196 VSS 0.031128f
C11489 DVDD.n6197 VSS 0.031128f
C11490 DVDD.n6198 VSS 0.031128f
C11491 DVDD.n6199 VSS 0.031128f
C11492 DVDD.n6200 VSS 0.031128f
C11493 DVDD.n6201 VSS 0.031128f
C11494 DVDD.n6202 VSS 0.031128f
C11495 DVDD.n6203 VSS 0.031128f
C11496 DVDD.n6204 VSS 0.031128f
C11497 DVDD.n6205 VSS 0.031128f
C11498 DVDD.n6206 VSS 0.031128f
C11499 DVDD.n6207 VSS 0.031128f
C11500 DVDD.n6208 VSS 0.031128f
C11501 DVDD.n6209 VSS 0.031128f
C11502 DVDD.n6210 VSS 0.031128f
C11503 DVDD.n6211 VSS 0.031128f
C11504 DVDD.n6212 VSS 0.031128f
C11505 DVDD.n6213 VSS 0.031128f
C11506 DVDD.n6214 VSS 0.031128f
C11507 DVDD.n6215 VSS 0.031128f
C11508 DVDD.n6216 VSS 0.031128f
C11509 DVDD.n6217 VSS 0.031128f
C11510 DVDD.n6218 VSS 0.031128f
C11511 DVDD.n6219 VSS 0.031128f
C11512 DVDD.n6220 VSS 0.031128f
C11513 DVDD.n6221 VSS 0.031128f
C11514 DVDD.n6222 VSS 0.031128f
C11515 DVDD.n6223 VSS 0.031128f
C11516 DVDD.n6224 VSS 0.031128f
C11517 DVDD.n6225 VSS 0.031128f
C11518 DVDD.n6226 VSS 0.031128f
C11519 DVDD.n6227 VSS 0.031128f
C11520 DVDD.n6228 VSS 0.031128f
C11521 DVDD.n6229 VSS 0.031128f
C11522 DVDD.n6230 VSS 0.031128f
C11523 DVDD.n6231 VSS 0.031128f
C11524 DVDD.n6232 VSS 0.031128f
C11525 DVDD.n6233 VSS 0.031128f
C11526 DVDD.n6234 VSS 0.031128f
C11527 DVDD.n6235 VSS 0.031128f
C11528 DVDD.n6236 VSS 0.031128f
C11529 DVDD.n6237 VSS 0.031128f
C11530 DVDD.n6238 VSS 0.031128f
C11531 DVDD.n6239 VSS 0.031128f
C11532 DVDD.n6240 VSS 0.031128f
C11533 DVDD.n6241 VSS 0.031128f
C11534 DVDD.n6242 VSS 0.031128f
C11535 DVDD.n6243 VSS 0.031128f
C11536 DVDD.n6244 VSS 0.031128f
C11537 DVDD.n6245 VSS 0.031128f
C11538 DVDD.n6246 VSS 0.031128f
C11539 DVDD.n6247 VSS 0.031128f
C11540 DVDD.n6248 VSS 0.031128f
C11541 DVDD.n6249 VSS 0.031128f
C11542 DVDD.n6250 VSS 0.031128f
C11543 DVDD.n6251 VSS 0.031128f
C11544 DVDD.n6252 VSS 0.031128f
C11545 DVDD.n6253 VSS 0.031128f
C11546 DVDD.n6254 VSS 0.031128f
C11547 DVDD.n6255 VSS 0.031128f
C11548 DVDD.n6256 VSS 0.031128f
C11549 DVDD.n6257 VSS 0.031128f
C11550 DVDD.n6258 VSS 0.031128f
C11551 DVDD.n6259 VSS 0.031128f
C11552 DVDD.n6260 VSS 0.031128f
C11553 DVDD.n6261 VSS 0.031128f
C11554 DVDD.n6262 VSS 0.031128f
C11555 DVDD.n6263 VSS 0.031128f
C11556 DVDD.n6264 VSS 0.031128f
C11557 DVDD.n6265 VSS 0.031128f
C11558 DVDD.n6266 VSS 0.031128f
C11559 DVDD.n6267 VSS 0.031128f
C11560 DVDD.n6268 VSS 0.031128f
C11561 DVDD.n6269 VSS 0.031128f
C11562 DVDD.n6270 VSS 0.031128f
C11563 DVDD.n6271 VSS 0.031128f
C11564 DVDD.n6272 VSS 0.031128f
C11565 DVDD.n6273 VSS 0.031128f
C11566 DVDD.n6274 VSS 0.031128f
C11567 DVDD.n6275 VSS 0.031128f
C11568 DVDD.n6276 VSS 0.031128f
C11569 DVDD.n6277 VSS 0.031128f
C11570 DVDD.n6278 VSS 0.031128f
C11571 DVDD.n6279 VSS 0.031128f
C11572 DVDD.n6280 VSS 0.031128f
C11573 DVDD.n6281 VSS 0.031128f
C11574 DVDD.n6282 VSS 0.031128f
C11575 DVDD.n6283 VSS 0.031128f
C11576 DVDD.n6284 VSS 0.031128f
C11577 DVDD.n6285 VSS 0.031128f
C11578 DVDD.n6286 VSS 0.031128f
C11579 DVDD.n6287 VSS 0.031128f
C11580 DVDD.n6288 VSS 0.031128f
C11581 DVDD.n6289 VSS 0.031128f
C11582 DVDD.n6290 VSS 0.031128f
C11583 DVDD.n6291 VSS 0.031128f
C11584 DVDD.n6292 VSS 0.031128f
C11585 DVDD.n6293 VSS 0.031128f
C11586 DVDD.n6294 VSS 0.031128f
C11587 DVDD.n6295 VSS 0.031128f
C11588 DVDD.n6296 VSS 0.031128f
C11589 DVDD.n6297 VSS 0.031128f
C11590 DVDD.n6298 VSS 0.031128f
C11591 DVDD.n6299 VSS 0.031128f
C11592 DVDD.n6300 VSS 0.031128f
C11593 DVDD.n6301 VSS 0.031128f
C11594 DVDD.n6302 VSS 0.031128f
C11595 DVDD.n6303 VSS 0.031128f
C11596 DVDD.n6304 VSS 0.031128f
C11597 DVDD.n6305 VSS 0.031128f
C11598 DVDD.n6306 VSS 0.031128f
C11599 DVDD.n6307 VSS 0.031128f
C11600 DVDD.n6308 VSS 0.031128f
C11601 DVDD.n6309 VSS 0.031128f
C11602 DVDD.n6310 VSS 0.031128f
C11603 DVDD.n6311 VSS 0.031128f
C11604 DVDD.n6312 VSS 0.031128f
C11605 DVDD.n6313 VSS 0.031128f
C11606 DVDD.n6314 VSS 0.031128f
C11607 DVDD.n6315 VSS 0.031128f
C11608 DVDD.n6316 VSS 0.031128f
C11609 DVDD.n6317 VSS 0.031128f
C11610 DVDD.n6318 VSS 0.031128f
C11611 DVDD.n6319 VSS 0.031128f
C11612 DVDD.n6320 VSS 0.031128f
C11613 DVDD.n6321 VSS 0.031128f
C11614 DVDD.n6322 VSS 0.031128f
C11615 DVDD.n6323 VSS 0.031128f
C11616 DVDD.n6324 VSS 0.031128f
C11617 DVDD.n6325 VSS 0.031128f
C11618 DVDD.n6326 VSS 0.031128f
C11619 DVDD.n6327 VSS 0.031128f
C11620 DVDD.n6328 VSS 0.031128f
C11621 DVDD.n6329 VSS 0.031128f
C11622 DVDD.n6331 VSS 0.366419f
C11623 DVDD.n6333 VSS 0.031128f
C11624 DVDD.n6334 VSS 0.031128f
C11625 DVDD.n6335 VSS 0.031128f
C11626 DVDD.n6336 VSS 0.031128f
C11627 DVDD.n6337 VSS 0.026086f
C11628 DVDD.n6338 VSS 0.0282f
C11629 DVDD.n6339 VSS 0.0282f
C11630 DVDD.n6340 VSS 0.041931f
C11631 DVDD.n6341 VSS 0.034696f
C11632 DVDD.n6342 VSS 0.024629f
C11633 DVDD.n6343 VSS 0.028833f
C11634 DVDD.n6344 VSS 0.028833f
C11635 DVDD.n6345 VSS 0.02513f
C11636 DVDD.n6346 VSS 0.041931f
C11637 DVDD.n6347 VSS 0.02513f
C11638 DVDD.n6348 VSS 0.189527f
C11639 DVDD.n6391 VSS 0.522252f
C11640 DVDD.n6392 VSS 0.033945f
C11641 DVDD.n6393 VSS 0.05956f
C11642 DVDD.n6394 VSS 0.033945f
C11643 DVDD.n6395 VSS 0.05956f
C11644 DVDD.n6396 VSS 0.028497f
C11645 DVDD.n6397 VSS 0.053165f
C11646 DVDD.n6398 VSS 0.05956f
C11647 DVDD.n6399 VSS 0.050592f
C11648 DVDD.n6400 VSS 0.056679f
C11649 DVDD.n6401 VSS 0.056679f
C11650 DVDD.n6402 VSS 0.598063f
C11651 DVDD.n6403 VSS 0.522252f
C11652 DVDD.n6404 VSS 0.019729f
C11653 DVDD.n6446 VSS 0.031128f
C11654 DVDD.n6447 VSS 0.031128f
C11655 DVDD.n6448 VSS 0.031128f
C11656 DVDD.n6449 VSS 0.031128f
C11657 DVDD.n6450 VSS 0.031128f
C11658 DVDD.n6451 VSS 0.031128f
C11659 DVDD.n6452 VSS 0.031128f
C11660 DVDD.n6453 VSS 0.031128f
C11661 DVDD.n6454 VSS 0.031128f
C11662 DVDD.n6455 VSS 0.031128f
C11663 DVDD.n6456 VSS 0.031128f
C11664 DVDD.n6457 VSS 0.031128f
C11665 DVDD.n6458 VSS 0.031128f
C11666 DVDD.n6459 VSS 0.031128f
C11667 DVDD.n6460 VSS 0.031128f
C11668 DVDD.n6461 VSS 0.031128f
C11669 DVDD.n6462 VSS 0.031128f
C11670 DVDD.n6463 VSS 0.031128f
C11671 DVDD.n6464 VSS 0.031128f
C11672 DVDD.n6465 VSS 0.031128f
C11673 DVDD.n6466 VSS 0.031128f
C11674 DVDD.n6467 VSS 0.031128f
C11675 DVDD.n6468 VSS 0.031128f
C11676 DVDD.n6469 VSS 0.031128f
C11677 DVDD.n6470 VSS 0.031128f
C11678 DVDD.n6471 VSS 0.031128f
C11679 DVDD.n6472 VSS 0.031128f
C11680 DVDD.n6473 VSS 0.031128f
C11681 DVDD.n6474 VSS 0.031128f
C11682 DVDD.n6475 VSS 0.031128f
C11683 DVDD.n6476 VSS 0.031128f
C11684 DVDD.n6477 VSS 0.031128f
C11685 DVDD.n6478 VSS 0.031128f
C11686 DVDD.n6479 VSS 0.031128f
C11687 DVDD.n6480 VSS 0.031128f
C11688 DVDD.n6481 VSS 0.031128f
C11689 DVDD.n6482 VSS 0.031128f
C11690 DVDD.n6483 VSS 0.031128f
C11691 DVDD.n6484 VSS 0.031128f
C11692 DVDD.n6485 VSS 0.031128f
C11693 DVDD.n6486 VSS 0.031128f
C11694 DVDD.n6487 VSS 0.031128f
C11695 DVDD.n6488 VSS 0.031128f
C11696 DVDD.n6489 VSS 0.031128f
C11697 DVDD.n6490 VSS 0.031128f
C11698 DVDD.n6491 VSS 0.031128f
C11699 DVDD.n6492 VSS 0.031128f
C11700 DVDD.n6493 VSS 0.031128f
C11701 DVDD.n6494 VSS 0.031128f
C11702 DVDD.n6495 VSS 0.031128f
C11703 DVDD.n6496 VSS 0.031128f
C11704 DVDD.n6497 VSS 0.031128f
C11705 DVDD.n6498 VSS 0.031128f
C11706 DVDD.n6499 VSS 0.031128f
C11707 DVDD.n6500 VSS 0.031128f
C11708 DVDD.n6501 VSS 0.031128f
C11709 DVDD.n6502 VSS 0.031128f
C11710 DVDD.n6503 VSS 0.031128f
C11711 DVDD.n6504 VSS 0.031128f
C11712 DVDD.n6505 VSS 0.031128f
C11713 DVDD.n6506 VSS 0.031128f
C11714 DVDD.n6507 VSS 0.031128f
C11715 DVDD.n6508 VSS 0.019729f
C11716 DVDD.n6509 VSS 0.031128f
C11717 DVDD.n6510 VSS 0.031128f
C11718 DVDD.n6511 VSS 0.031128f
C11719 DVDD.n6512 VSS 0.031128f
C11720 DVDD.n6513 VSS 0.031128f
C11721 DVDD.n6514 VSS 0.031128f
C11722 DVDD.n6515 VSS 0.031128f
C11723 DVDD.n6516 VSS 0.031128f
C11724 DVDD.n6517 VSS 0.031128f
C11725 DVDD.n6518 VSS 0.031128f
C11726 DVDD.n6519 VSS 0.031128f
C11727 DVDD.n6520 VSS 0.031128f
C11728 DVDD.n6521 VSS 0.031128f
C11729 DVDD.n6522 VSS 0.031128f
C11730 DVDD.n6523 VSS 0.031128f
C11731 DVDD.n6524 VSS 0.031128f
C11732 DVDD.n6525 VSS 0.031128f
C11733 DVDD.n6526 VSS 0.031128f
C11734 DVDD.n6527 VSS 0.031128f
C11735 DVDD.n6528 VSS 0.031128f
C11736 DVDD.n6529 VSS 0.031128f
C11737 DVDD.n6530 VSS 0.031128f
C11738 DVDD.n6531 VSS 0.031128f
C11739 DVDD.n6532 VSS 0.031128f
C11740 DVDD.n6533 VSS 0.031128f
C11741 DVDD.n6534 VSS 0.031128f
C11742 DVDD.n6535 VSS 0.031128f
C11743 DVDD.n6536 VSS 0.031128f
C11744 DVDD.n6537 VSS 0.031128f
C11745 DVDD.n6538 VSS 0.031128f
C11746 DVDD.n6539 VSS 0.031128f
C11747 DVDD.n6540 VSS 0.031128f
C11748 DVDD.n6541 VSS 0.031128f
C11749 DVDD.n6542 VSS 0.031128f
C11750 DVDD.n6543 VSS 0.031128f
C11751 DVDD.n6544 VSS 0.031128f
C11752 DVDD.n6545 VSS 0.031128f
C11753 DVDD.n6546 VSS 0.031128f
C11754 DVDD.n6547 VSS 0.031128f
C11755 DVDD.n6548 VSS 0.031128f
C11756 DVDD.n6549 VSS 0.031128f
C11757 DVDD.n6550 VSS 0.031128f
C11758 DVDD.n6551 VSS 0.031128f
C11759 DVDD.n6552 VSS 0.031128f
C11760 DVDD.n6553 VSS 0.031128f
C11761 DVDD.n6554 VSS 0.031128f
C11762 DVDD.n6555 VSS 0.031128f
C11763 DVDD.n6556 VSS 0.031128f
C11764 DVDD.n6557 VSS 0.031128f
C11765 DVDD.n6558 VSS 0.031128f
C11766 DVDD.n6559 VSS 0.031128f
C11767 DVDD.n6560 VSS 0.031128f
C11768 DVDD.n6561 VSS 0.031128f
C11769 DVDD.n6562 VSS 0.031128f
C11770 DVDD.n6563 VSS 0.031128f
C11771 DVDD.n6564 VSS 0.031128f
C11772 DVDD.n6565 VSS 0.031128f
C11773 DVDD.n6566 VSS 0.031128f
C11774 DVDD.n6567 VSS 0.031128f
C11775 DVDD.n6568 VSS 0.031128f
C11776 DVDD.n6569 VSS 0.031128f
C11777 DVDD.n6570 VSS 0.031128f
C11778 DVDD.n6571 VSS 0.031128f
C11779 DVDD.n6572 VSS 0.031128f
C11780 DVDD.n6573 VSS 0.031128f
C11781 DVDD.n6574 VSS 0.031128f
C11782 DVDD.n6575 VSS 0.031128f
C11783 DVDD.n6576 VSS 0.031128f
C11784 DVDD.n6577 VSS 0.031128f
C11785 DVDD.n6578 VSS 0.031128f
C11786 DVDD.n6579 VSS 0.031128f
C11787 DVDD.n6580 VSS 0.031128f
C11788 DVDD.n6581 VSS 0.031128f
C11789 DVDD.n6582 VSS 0.031128f
C11790 DVDD.n6583 VSS 0.031128f
C11791 DVDD.n6584 VSS 0.031128f
C11792 DVDD.n6585 VSS 0.031128f
C11793 DVDD.n6586 VSS 0.031128f
C11794 DVDD.n6587 VSS 0.031128f
C11795 DVDD.n6588 VSS 0.031128f
C11796 DVDD.n6589 VSS 0.031128f
C11797 DVDD.n6590 VSS 0.031128f
C11798 DVDD.n6591 VSS 0.031128f
C11799 DVDD.n6592 VSS 0.031128f
C11800 DVDD.n6593 VSS 0.031128f
C11801 DVDD.n6594 VSS 0.031128f
C11802 DVDD.n6595 VSS 0.031128f
C11803 DVDD.n6596 VSS 0.031128f
C11804 DVDD.n6597 VSS 0.031128f
C11805 DVDD.n6598 VSS 0.031128f
C11806 DVDD.n6599 VSS 0.031128f
C11807 DVDD.n6600 VSS 0.031128f
C11808 DVDD.n6601 VSS 0.031128f
C11809 DVDD.n6602 VSS 0.031128f
C11810 DVDD.n6603 VSS 0.031128f
C11811 DVDD.n6604 VSS 0.031128f
C11812 DVDD.n6605 VSS 0.031128f
C11813 DVDD.n6606 VSS 0.031128f
C11814 DVDD.n6607 VSS 0.031128f
C11815 DVDD.n6608 VSS 0.031128f
C11816 DVDD.n6609 VSS 0.031128f
C11817 DVDD.n6610 VSS 0.031128f
C11818 DVDD.n6611 VSS 0.031128f
C11819 DVDD.n6612 VSS 0.031128f
C11820 DVDD.n6613 VSS 0.031128f
C11821 DVDD.n6614 VSS 0.031128f
C11822 DVDD.n6615 VSS 0.031128f
C11823 DVDD.n6616 VSS 0.031128f
C11824 DVDD.n6617 VSS 0.031128f
C11825 DVDD.n6618 VSS 0.031128f
C11826 DVDD.n6619 VSS 0.031128f
C11827 DVDD.n6620 VSS 0.031128f
C11828 DVDD.n6621 VSS 0.031128f
C11829 DVDD.n6622 VSS 0.031128f
C11830 DVDD.n6623 VSS 0.031128f
C11831 DVDD.n6624 VSS 0.031128f
C11832 DVDD.n6625 VSS 0.031128f
C11833 DVDD.n6626 VSS 0.031128f
C11834 DVDD.n6627 VSS 0.031128f
C11835 DVDD.n6628 VSS 0.031128f
C11836 DVDD.n6629 VSS 0.031128f
C11837 DVDD.n6630 VSS 0.031128f
C11838 DVDD.n6631 VSS 0.031128f
C11839 DVDD.n6632 VSS 0.031128f
C11840 DVDD.n6633 VSS 0.031128f
C11841 DVDD.n6634 VSS 0.031128f
C11842 DVDD.n6635 VSS 0.031128f
C11843 DVDD.n6636 VSS 0.031128f
C11844 DVDD.n6637 VSS 0.031128f
C11845 DVDD.n6638 VSS 0.031128f
C11846 DVDD.n6639 VSS 0.031128f
C11847 DVDD.n6640 VSS 0.031128f
C11848 DVDD.n6641 VSS 0.031128f
C11849 DVDD.n6642 VSS 0.031128f
C11850 DVDD.n6643 VSS 0.031128f
C11851 DVDD.n6644 VSS 0.031128f
C11852 DVDD.n6645 VSS 0.031128f
C11853 DVDD.n6646 VSS 0.031128f
C11854 DVDD.n6647 VSS 0.031128f
C11855 DVDD.n6648 VSS 0.031128f
C11856 DVDD.n6649 VSS 0.031128f
C11857 DVDD.n6650 VSS 0.031128f
C11858 DVDD.n6651 VSS 0.031128f
C11859 DVDD.n6652 VSS 0.031128f
C11860 DVDD.n6653 VSS 0.031128f
C11861 DVDD.n6654 VSS 0.031128f
C11862 DVDD.n6655 VSS 0.031128f
C11863 DVDD.n6656 VSS 0.031128f
C11864 DVDD.n6657 VSS 0.031128f
C11865 DVDD.n6658 VSS 0.031128f
C11866 DVDD.n6659 VSS 0.031128f
C11867 DVDD.n6660 VSS 0.031128f
C11868 DVDD.n6661 VSS 0.031128f
C11869 DVDD.n6662 VSS 0.031128f
C11870 DVDD.n6663 VSS 0.031128f
C11871 DVDD.n6664 VSS 0.031128f
C11872 DVDD.n6665 VSS 0.031128f
C11873 DVDD.n6666 VSS 0.031128f
C11874 DVDD.n6667 VSS 0.031128f
C11875 DVDD.n6668 VSS 0.031128f
C11876 DVDD.n6669 VSS 0.031128f
C11877 DVDD.n6670 VSS 0.031128f
C11878 DVDD.n6671 VSS 0.031128f
C11879 DVDD.n6672 VSS 0.031128f
C11880 DVDD.n6673 VSS 0.031128f
C11881 DVDD.n6674 VSS 0.031128f
C11882 DVDD.n6675 VSS 0.031128f
C11883 DVDD.n6676 VSS 0.031128f
C11884 DVDD.n6677 VSS 0.031128f
C11885 DVDD.n6678 VSS 0.031128f
C11886 DVDD.n6679 VSS 0.031128f
C11887 DVDD.n6680 VSS 0.031128f
C11888 DVDD.n6681 VSS 0.031128f
C11889 DVDD.n6682 VSS 0.031128f
C11890 DVDD.n6683 VSS 0.031128f
C11891 DVDD.n6684 VSS 0.031128f
C11892 DVDD.n6685 VSS 0.031128f
C11893 DVDD.n6686 VSS 0.031128f
C11894 DVDD.n6687 VSS 0.031128f
C11895 DVDD.n6688 VSS 0.031128f
C11896 DVDD.n6689 VSS 0.031128f
C11897 DVDD.n6690 VSS 0.031128f
C11898 DVDD.n6691 VSS 0.031128f
C11899 DVDD.n6692 VSS 0.031128f
C11900 DVDD.n6693 VSS 0.026086f
C11901 DVDD.n6694 VSS 0.019729f
C11902 DVDD.n6695 VSS 0.019729f
C11903 DVDD.n6696 VSS 0.522253f
C11904 DVDD.n6697 VSS 0.408536f
C11905 DVDD.n6698 VSS 0.05956f
C11906 DVDD.n6699 VSS 0.039387f
C11907 DVDD.n6700 VSS 0.039387f
C11908 DVDD.n6701 VSS 0.035157f
C11909 DVDD.n6702 VSS 0.039516f
C11910 DVDD.n6703 VSS 0.039516f
C11911 DVDD.n6704 VSS 0.033945f
C11912 DVDD.n6705 VSS 0.033945f
C11913 DVDD.n6706 VSS 0.598063f
C11914 DVDD.n6707 VSS 0.522252f
C11915 DVDD.n6749 VSS 0.522252f
C11916 DVDD.n6750 VSS 0.031128f
C11917 DVDD.n6751 VSS 0.019729f
C11918 DVDD.n6752 VSS 0.299032f
C11919 DVDD.n6794 VSS 0.446441f
C11920 DVDD.n6795 VSS 0.02513f
C11921 DVDD.n6796 VSS 0.031128f
C11922 DVDD.n6797 VSS 0.031128f
C11923 DVDD.n6798 VSS 0.031128f
C11924 DVDD.n6799 VSS 0.031128f
C11925 DVDD.n6800 VSS 0.031128f
C11926 DVDD.n6801 VSS 0.031128f
C11927 DVDD.n6802 VSS 0.031128f
C11928 DVDD.n6803 VSS 0.031128f
C11929 DVDD.n6804 VSS 0.031128f
C11930 DVDD.n6805 VSS 0.031128f
C11931 DVDD.n6806 VSS 0.031128f
C11932 DVDD.n6807 VSS 0.031128f
C11933 DVDD.n6808 VSS 0.031128f
C11934 DVDD.n6809 VSS 0.031128f
C11935 DVDD.n6810 VSS 0.031128f
C11936 DVDD.n6811 VSS 0.031128f
C11937 DVDD.n6812 VSS 0.031128f
C11938 DVDD.n6813 VSS 0.031128f
C11939 DVDD.n6814 VSS 0.031128f
C11940 DVDD.n6815 VSS 0.031128f
C11941 DVDD.n6816 VSS 0.031128f
C11942 DVDD.n6817 VSS 0.031128f
C11943 DVDD.n6818 VSS 0.031128f
C11944 DVDD.n6819 VSS 0.031128f
C11945 DVDD.n6820 VSS 0.031128f
C11946 DVDD.n6821 VSS 0.031128f
C11947 DVDD.n6822 VSS 0.031128f
C11948 DVDD.n6823 VSS 0.031128f
C11949 DVDD.n6824 VSS 0.031128f
C11950 DVDD.n6825 VSS 0.031128f
C11951 DVDD.n6826 VSS 0.031128f
C11952 DVDD.n6827 VSS 0.031128f
C11953 DVDD.n6828 VSS 0.031128f
C11954 DVDD.n6829 VSS 0.031128f
C11955 DVDD.n6830 VSS 0.031128f
C11956 DVDD.n6831 VSS 0.031128f
C11957 DVDD.n6832 VSS 0.031128f
C11958 DVDD.n6833 VSS 0.031128f
C11959 DVDD.n6834 VSS 0.031128f
C11960 DVDD.n6835 VSS 0.031128f
C11961 DVDD.n6836 VSS 0.031128f
C11962 DVDD.n6837 VSS 0.031128f
C11963 DVDD.n6838 VSS 0.031128f
C11964 DVDD.n6839 VSS 0.031128f
C11965 DVDD.n6840 VSS 0.031128f
C11966 DVDD.n6841 VSS 0.031128f
C11967 DVDD.n6842 VSS 0.031128f
C11968 DVDD.n6843 VSS 0.031128f
C11969 DVDD.n6844 VSS 0.031128f
C11970 DVDD.n6845 VSS 0.031128f
C11971 DVDD.n6846 VSS 0.031128f
C11972 DVDD.n6847 VSS 0.031128f
C11973 DVDD.n6848 VSS 0.031128f
C11974 DVDD.n6849 VSS 0.031128f
C11975 DVDD.n6850 VSS 0.031128f
C11976 DVDD.n6851 VSS 0.031128f
C11977 DVDD.n6852 VSS 0.031128f
C11978 DVDD.n6853 VSS 0.031128f
C11979 DVDD.n6854 VSS 0.031128f
C11980 DVDD.n6855 VSS 0.031128f
C11981 DVDD.n6856 VSS 0.031128f
C11982 DVDD.n6857 VSS 0.031128f
C11983 DVDD.n6858 VSS 0.028497f
C11984 DVDD.n6859 VSS 0.031128f
C11985 DVDD.n6860 VSS 0.031128f
C11986 DVDD.n6861 VSS 0.031128f
C11987 DVDD.n6862 VSS 0.031128f
C11988 DVDD.n6863 VSS 0.031128f
C11989 DVDD.n6864 VSS 0.031128f
C11990 DVDD.n6865 VSS 0.031128f
C11991 DVDD.n6866 VSS 0.031128f
C11992 DVDD.n6867 VSS 0.031128f
C11993 DVDD.n6868 VSS 0.031128f
C11994 DVDD.n6869 VSS 0.031128f
C11995 DVDD.n6870 VSS 0.031128f
C11996 DVDD.n6871 VSS 0.031128f
C11997 DVDD.n6872 VSS 0.031128f
C11998 DVDD.n6873 VSS 0.031128f
C11999 DVDD.n6874 VSS 0.031128f
C12000 DVDD.n6875 VSS 0.031128f
C12001 DVDD.n6876 VSS 0.031128f
C12002 DVDD.n6877 VSS 0.031128f
C12003 DVDD.n6878 VSS 0.031128f
C12004 DVDD.n6879 VSS 0.031128f
C12005 DVDD.n6880 VSS 0.031128f
C12006 DVDD.n6881 VSS 0.031128f
C12007 DVDD.n6882 VSS 0.031128f
C12008 DVDD.n6883 VSS 0.031128f
C12009 DVDD.n6884 VSS 0.031128f
C12010 DVDD.n6885 VSS 0.031128f
C12011 DVDD.n6886 VSS 0.031128f
C12012 DVDD.n6887 VSS 0.031128f
C12013 DVDD.n6888 VSS 0.031128f
C12014 DVDD.n6889 VSS 0.031128f
C12015 DVDD.n6890 VSS 0.031128f
C12016 DVDD.n6891 VSS 0.031128f
C12017 DVDD.n6892 VSS 0.031128f
C12018 DVDD.n6893 VSS 0.031128f
C12019 DVDD.n6894 VSS 0.031128f
C12020 DVDD.n6895 VSS 0.031128f
C12021 DVDD.n6896 VSS 0.031128f
C12022 DVDD.n6897 VSS 0.031128f
C12023 DVDD.n6898 VSS 0.031128f
C12024 DVDD.n6899 VSS 0.031128f
C12025 DVDD.n6900 VSS 0.031128f
C12026 DVDD.n6901 VSS 0.031128f
C12027 DVDD.n6902 VSS 0.031128f
C12028 DVDD.n6903 VSS 0.031128f
C12029 DVDD.n6904 VSS 0.031128f
C12030 DVDD.n6905 VSS 0.031128f
C12031 DVDD.n6906 VSS 0.031128f
C12032 DVDD.n6907 VSS 0.031128f
C12033 DVDD.n6908 VSS 0.031128f
C12034 DVDD.n6909 VSS 0.031128f
C12035 DVDD.n6910 VSS 0.031128f
C12036 DVDD.n6911 VSS 0.031128f
C12037 DVDD.n6912 VSS 0.031128f
C12038 DVDD.n6913 VSS 0.031128f
C12039 DVDD.n6914 VSS 0.031128f
C12040 DVDD.n6915 VSS 0.031128f
C12041 DVDD.n6916 VSS 0.031128f
C12042 DVDD.n6917 VSS 0.031128f
C12043 DVDD.n6918 VSS 0.031128f
C12044 DVDD.n6919 VSS 0.031128f
C12045 DVDD.n6920 VSS 0.031128f
C12046 DVDD.n6921 VSS 0.031128f
C12047 DVDD.n6922 VSS 0.031128f
C12048 DVDD.n6923 VSS 0.031128f
C12049 DVDD.n6924 VSS 0.031128f
C12050 DVDD.n6925 VSS 0.031128f
C12051 DVDD.n6926 VSS 0.031128f
C12052 DVDD.n6927 VSS 0.031128f
C12053 DVDD.n6928 VSS 0.031128f
C12054 DVDD.n6929 VSS 0.031128f
C12055 DVDD.n6930 VSS 0.031128f
C12056 DVDD.n6931 VSS 0.031128f
C12057 DVDD.n6932 VSS 0.031128f
C12058 DVDD.n6933 VSS 0.031128f
C12059 DVDD.n6934 VSS 0.031128f
C12060 DVDD.n6935 VSS 0.031128f
C12061 DVDD.n6936 VSS 0.031128f
C12062 DVDD.n6937 VSS 0.031128f
C12063 DVDD.n6938 VSS 0.031128f
C12064 DVDD.n6939 VSS 0.031128f
C12065 DVDD.n6940 VSS 0.031128f
C12066 DVDD.n6941 VSS 0.031128f
C12067 DVDD.n6942 VSS 0.031128f
C12068 DVDD.n6943 VSS 0.031128f
C12069 DVDD.n6944 VSS 0.031128f
C12070 DVDD.n6945 VSS 0.031128f
C12071 DVDD.n6946 VSS 0.031128f
C12072 DVDD.n6947 VSS 0.031128f
C12073 DVDD.n6948 VSS 0.031128f
C12074 DVDD.n6949 VSS 0.031128f
C12075 DVDD.n6950 VSS 0.031128f
C12076 DVDD.n6951 VSS 0.031128f
C12077 DVDD.n6952 VSS 0.031128f
C12078 DVDD.n6953 VSS 0.031128f
C12079 DVDD.n6954 VSS 0.031128f
C12080 DVDD.n6955 VSS 0.031128f
C12081 DVDD.n6956 VSS 0.031128f
C12082 DVDD.n6957 VSS 0.031128f
C12083 DVDD.n6958 VSS 0.031128f
C12084 DVDD.n6959 VSS 0.031128f
C12085 DVDD.n6960 VSS 0.031128f
C12086 DVDD.n6961 VSS 0.031128f
C12087 DVDD.n6962 VSS 0.031128f
C12088 DVDD.n6963 VSS 0.031128f
C12089 DVDD.n6964 VSS 0.031128f
C12090 DVDD.n6965 VSS 0.031128f
C12091 DVDD.n6966 VSS 0.031128f
C12092 DVDD.n6967 VSS 0.031128f
C12093 DVDD.n6968 VSS 0.031128f
C12094 DVDD.n6969 VSS 0.031128f
C12095 DVDD.n6970 VSS 0.031128f
C12096 DVDD.n6971 VSS 0.031128f
C12097 DVDD.n6972 VSS 0.031128f
C12098 DVDD.n6973 VSS 0.031128f
C12099 DVDD.n6974 VSS 0.031128f
C12100 DVDD.n6975 VSS 0.031128f
C12101 DVDD.n6976 VSS 0.031128f
C12102 DVDD.n6977 VSS 0.031128f
C12103 DVDD.n6978 VSS 0.031128f
C12104 DVDD.n6979 VSS 0.031128f
C12105 DVDD.n6980 VSS 0.031128f
C12106 DVDD.n6981 VSS 0.031128f
C12107 DVDD.n6982 VSS 0.031128f
C12108 DVDD.n6983 VSS 0.031128f
C12109 DVDD.n6984 VSS 0.031128f
C12110 DVDD.n6985 VSS 0.031128f
C12111 DVDD.n6986 VSS 0.031128f
C12112 DVDD.n6987 VSS 0.031128f
C12113 DVDD.n6988 VSS 0.031128f
C12114 DVDD.n6989 VSS 0.031128f
C12115 DVDD.n6990 VSS 0.031128f
C12116 DVDD.n6991 VSS 0.031128f
C12117 DVDD.n6992 VSS 0.031128f
C12118 DVDD.n6993 VSS 0.031128f
C12119 DVDD.n6994 VSS 0.031128f
C12120 DVDD.n6995 VSS 0.031128f
C12121 DVDD.n6996 VSS 0.031128f
C12122 DVDD.n6997 VSS 0.031128f
C12123 DVDD.n6998 VSS 0.031128f
C12124 DVDD.n6999 VSS 0.031128f
C12125 DVDD.n7000 VSS 0.031128f
C12126 DVDD.n7001 VSS 0.031128f
C12127 DVDD.n7002 VSS 0.031128f
C12128 DVDD.n7003 VSS 0.031128f
C12129 DVDD.n7004 VSS 0.031128f
C12130 DVDD.n7005 VSS 0.031128f
C12131 DVDD.n7006 VSS 0.031128f
C12132 DVDD.n7007 VSS 0.031128f
C12133 DVDD.n7008 VSS 0.031128f
C12134 DVDD.n7009 VSS 0.031128f
C12135 DVDD.n7010 VSS 0.031128f
C12136 DVDD.n7011 VSS 0.031128f
C12137 DVDD.n7012 VSS 0.031128f
C12138 DVDD.n7013 VSS 0.031128f
C12139 DVDD.n7014 VSS 0.031128f
C12140 DVDD.n7015 VSS 0.031128f
C12141 DVDD.n7016 VSS 0.031128f
C12142 DVDD.n7017 VSS 0.031128f
C12143 DVDD.n7018 VSS 0.031128f
C12144 DVDD.n7019 VSS 0.031128f
C12145 DVDD.n7020 VSS 0.031128f
C12146 DVDD.n7021 VSS 0.031128f
C12147 DVDD.n7022 VSS 0.031128f
C12148 DVDD.n7023 VSS 0.031128f
C12149 DVDD.n7024 VSS 0.031128f
C12150 DVDD.n7025 VSS 0.031128f
C12151 DVDD.n7026 VSS 0.031128f
C12152 DVDD.n7027 VSS 0.031128f
C12153 DVDD.n7028 VSS 0.031128f
C12154 DVDD.n7029 VSS 0.031128f
C12155 DVDD.n7030 VSS 0.031128f
C12156 DVDD.n7031 VSS 0.031128f
C12157 DVDD.n7032 VSS 0.031128f
C12158 DVDD.n7033 VSS 0.031128f
C12159 DVDD.n7034 VSS 0.031128f
C12160 DVDD.n7035 VSS 0.031128f
C12161 DVDD.n7036 VSS 0.031128f
C12162 DVDD.n7037 VSS 0.031128f
C12163 DVDD.n7038 VSS 0.031128f
C12164 DVDD.n7039 VSS 0.031128f
C12165 DVDD.n7040 VSS 0.031128f
C12166 DVDD.n7041 VSS 0.031128f
C12167 DVDD.n7042 VSS 0.026086f
C12168 DVDD.n7043 VSS 0.041488f
C12169 DVDD.n7044 VSS 0.041931f
C12170 DVDD.n7045 VSS 0.021408f
C12171 DVDD.n7046 VSS 0.041488f
C12172 DVDD.n7047 VSS 0.038535f
C12173 DVDD.n7048 VSS 0.038535f
C12174 DVDD.n7049 VSS 0.033655f
C12175 DVDD.n7050 VSS 0.036234f
C12176 DVDD.n7051 VSS 0.028833f
C12177 DVDD.n7052 VSS 0.028833f
C12178 DVDD.n7053 VSS 0.02513f
C12179 DVDD.n7054 VSS 0.041931f
C12180 DVDD.n7055 VSS 0.02513f
C12181 DVDD.n7056 VSS 0.598063f
C12182 DVDD.n7057 VSS 0.522252f
C12183 DVDD.n7058 VSS 0.05956f
C12184 DVDD.n7059 VSS 0.033945f
C12185 DVDD.n7060 VSS 0.05956f
C12186 DVDD.n7061 VSS 0.033945f
C12187 DVDD.n7062 VSS 0.043229f
C12188 DVDD.n7063 VSS 0.043229f
C12189 DVDD.n7064 VSS 0.038587f
C12190 DVDD.n7065 VSS 0.053165f
C12191 DVDD.n7066 VSS 0.028497f
C12192 DVDD.n7067 VSS 0.053165f
C12193 DVDD.n7068 VSS 0.05956f
C12194 DVDD.n7069 VSS 0.05956f
C12195 DVDD.n7111 VSS 0.019729f
C12196 DVDD.n7112 VSS 0.019729f
C12197 DVDD.n7113 VSS 0.031128f
C12198 DVDD.n7114 VSS 0.031128f
C12199 DVDD.n7115 VSS 0.031128f
C12200 DVDD.n7116 VSS 0.031128f
C12201 DVDD.n7117 VSS 0.031128f
C12202 DVDD.n7118 VSS 0.031128f
C12203 DVDD.n7119 VSS 0.031128f
C12204 DVDD.n7120 VSS 0.031128f
C12205 DVDD.n7121 VSS 0.031128f
C12206 DVDD.n7122 VSS 0.031128f
C12207 DVDD.n7123 VSS 0.031128f
C12208 DVDD.n7124 VSS 0.031128f
C12209 DVDD.n7125 VSS 0.031128f
C12210 DVDD.n7126 VSS 0.031128f
C12211 DVDD.n7127 VSS 0.031128f
C12212 DVDD.n7128 VSS 0.031128f
C12213 DVDD.n7129 VSS 0.031128f
C12214 DVDD.n7130 VSS 0.031128f
C12215 DVDD.n7131 VSS 0.031128f
C12216 DVDD.n7132 VSS 0.031128f
C12217 DVDD.n7133 VSS 0.031128f
C12218 DVDD.n7134 VSS 0.031128f
C12219 DVDD.n7135 VSS 0.031128f
C12220 DVDD.n7136 VSS 0.031128f
C12221 DVDD.n7137 VSS 0.031128f
C12222 DVDD.n7138 VSS 0.031128f
C12223 DVDD.n7139 VSS 0.031128f
C12224 DVDD.n7140 VSS 0.031128f
C12225 DVDD.n7141 VSS 0.031128f
C12226 DVDD.n7142 VSS 0.031128f
C12227 DVDD.n7143 VSS 0.031128f
C12228 DVDD.n7144 VSS 0.031128f
C12229 DVDD.n7145 VSS 0.031128f
C12230 DVDD.n7146 VSS 0.031128f
C12231 DVDD.n7147 VSS 0.031128f
C12232 DVDD.n7148 VSS 0.031128f
C12233 DVDD.n7149 VSS 0.031128f
C12234 DVDD.n7150 VSS 0.031128f
C12235 DVDD.n7151 VSS 0.031128f
C12236 DVDD.n7152 VSS 0.031128f
C12237 DVDD.n7153 VSS 0.019729f
C12238 DVDD.n7155 VSS 0.031128f
C12239 DVDD.n7156 VSS 0.031128f
C12240 DVDD.n7157 VSS 0.031128f
C12241 DVDD.n7158 VSS 0.031128f
C12242 DVDD.n7159 VSS 0.031128f
C12243 DVDD.n7160 VSS 0.031128f
C12244 DVDD.n7162 VSS 0.031128f
C12245 DVDD.n7163 VSS 0.031128f
C12246 DVDD.n7164 VSS 0.031128f
C12247 DVDD.n7166 VSS 0.031128f
C12248 DVDD.n7167 VSS 0.031128f
C12249 DVDD.n7168 VSS 0.031128f
C12250 DVDD.n7169 VSS 0.031128f
C12251 DVDD.n7170 VSS 0.031128f
C12252 DVDD.n7171 VSS 0.031128f
C12253 DVDD.n7172 VSS 0.031128f
C12254 DVDD.n7174 VSS 0.031128f
C12255 DVDD.n7175 VSS 0.031128f
C12256 DVDD.n7176 VSS 0.031128f
C12257 DVDD.n7178 VSS 0.031128f
C12258 DVDD.n7179 VSS 0.031128f
C12259 DVDD.n7180 VSS 0.031128f
C12260 DVDD.n7181 VSS 0.031128f
C12261 DVDD.n7182 VSS 0.031128f
C12262 DVDD.n7183 VSS 0.031128f
C12263 DVDD.n7184 VSS 0.031128f
C12264 DVDD.n7186 VSS 0.031128f
C12265 DVDD.n7187 VSS 0.031128f
C12266 DVDD.n7188 VSS 0.031128f
C12267 DVDD.n7190 VSS 0.031128f
C12268 DVDD.n7191 VSS 0.031128f
C12269 DVDD.n7192 VSS 0.031128f
C12270 DVDD.n7193 VSS 0.031128f
C12271 DVDD.n7194 VSS 0.031128f
C12272 DVDD.n7195 VSS 0.031128f
C12273 DVDD.n7196 VSS 0.031128f
C12274 DVDD.n7198 VSS 0.031128f
C12275 DVDD.n7199 VSS 0.031128f
C12276 DVDD.n7200 VSS 0.031128f
C12277 DVDD.n7202 VSS 0.031128f
C12278 DVDD.n7203 VSS 0.031128f
C12279 DVDD.n7204 VSS 0.031128f
C12280 DVDD.n7205 VSS 0.031128f
C12281 DVDD.n7206 VSS 0.031128f
C12282 DVDD.n7207 VSS 0.031128f
C12283 DVDD.n7208 VSS 0.031128f
C12284 DVDD.n7210 VSS 0.031128f
C12285 DVDD.n7211 VSS 0.031128f
C12286 DVDD.n7212 VSS 0.031128f
C12287 DVDD.n7214 VSS 0.031128f
C12288 DVDD.n7215 VSS 0.031128f
C12289 DVDD.n7216 VSS 0.031128f
C12290 DVDD.n7217 VSS 0.031128f
C12291 DVDD.n7218 VSS 0.031128f
C12292 DVDD.n7219 VSS 0.031128f
C12293 DVDD.n7220 VSS 0.031128f
C12294 DVDD.n7222 VSS 0.031128f
C12295 DVDD.n7223 VSS 0.031128f
C12296 DVDD.n7224 VSS 0.031128f
C12297 DVDD.n7226 VSS 0.031128f
C12298 DVDD.n7227 VSS 0.031128f
C12299 DVDD.n7228 VSS 0.031128f
C12300 DVDD.n7229 VSS 0.031128f
C12301 DVDD.n7230 VSS 0.031128f
C12302 DVDD.n7231 VSS 0.031128f
C12303 DVDD.n7232 VSS 0.031128f
C12304 DVDD.n7234 VSS 0.031128f
C12305 DVDD.n7235 VSS 0.031128f
C12306 DVDD.n7236 VSS 0.031128f
C12307 DVDD.n7238 VSS 0.031128f
C12308 DVDD.n7239 VSS 0.031128f
C12309 DVDD.n7240 VSS 0.031128f
C12310 DVDD.n7241 VSS 0.031128f
C12311 DVDD.n7242 VSS 0.031128f
C12312 DVDD.n7243 VSS 0.031128f
C12313 DVDD.n7244 VSS 0.031128f
C12314 DVDD.n7246 VSS 0.031128f
C12315 DVDD.n7247 VSS 0.031128f
C12316 DVDD.n7248 VSS 0.031128f
C12317 DVDD.n7250 VSS 0.031128f
C12318 DVDD.n7251 VSS 0.031128f
C12319 DVDD.n7252 VSS 0.031128f
C12320 DVDD.n7253 VSS 0.031128f
C12321 DVDD.n7254 VSS 0.031128f
C12322 DVDD.n7255 VSS 0.031128f
C12323 DVDD.n7256 VSS 0.031128f
C12324 DVDD.n7258 VSS 0.031128f
C12325 DVDD.n7259 VSS 0.031128f
C12326 DVDD.n7260 VSS 0.031128f
C12327 DVDD.n7262 VSS 0.031128f
C12328 DVDD.n7263 VSS 0.031128f
C12329 DVDD.n7264 VSS 0.031128f
C12330 DVDD.n7265 VSS 0.031128f
C12331 DVDD.n7266 VSS 0.031128f
C12332 DVDD.n7267 VSS 0.031128f
C12333 DVDD.n7268 VSS 0.031128f
C12334 DVDD.n7270 VSS 0.031128f
C12335 DVDD.n7271 VSS 0.031128f
C12336 DVDD.n7272 VSS 0.031128f
C12337 DVDD.n7274 VSS 0.031128f
C12338 DVDD.n7275 VSS 0.031128f
C12339 DVDD.n7276 VSS 0.031128f
C12340 DVDD.n7277 VSS 0.031128f
C12341 DVDD.n7278 VSS 0.031128f
C12342 DVDD.n7279 VSS 0.031128f
C12343 DVDD.n7280 VSS 0.031128f
C12344 DVDD.n7282 VSS 0.031128f
C12345 DVDD.n7283 VSS 0.031128f
C12346 DVDD.n7284 VSS 0.031128f
C12347 DVDD.n7286 VSS 0.031128f
C12348 DVDD.n7287 VSS 0.031128f
C12349 DVDD.n7288 VSS 0.031128f
C12350 DVDD.n7289 VSS 0.031128f
C12351 DVDD.n7290 VSS 0.031128f
C12352 DVDD.n7291 VSS 0.031128f
C12353 DVDD.n7292 VSS 0.031128f
C12354 DVDD.n7294 VSS 0.031128f
C12355 DVDD.n7295 VSS 0.031128f
C12356 DVDD.n7296 VSS 0.031128f
C12357 DVDD.n7298 VSS 0.031128f
C12358 DVDD.n7299 VSS 0.031128f
C12359 DVDD.n7300 VSS 0.031128f
C12360 DVDD.n7301 VSS 0.031128f
C12361 DVDD.n7302 VSS 0.031128f
C12362 DVDD.n7303 VSS 0.031128f
C12363 DVDD.n7304 VSS 0.031128f
C12364 DVDD.n7306 VSS 0.031128f
C12365 DVDD.n7307 VSS 0.031128f
C12366 DVDD.n7308 VSS 0.031128f
C12367 DVDD.n7310 VSS 0.031128f
C12368 DVDD.n7311 VSS 0.031128f
C12369 DVDD.n7312 VSS 0.031128f
C12370 DVDD.n7313 VSS 0.031128f
C12371 DVDD.n7314 VSS 0.031128f
C12372 DVDD.n7315 VSS 0.031128f
C12373 DVDD.n7316 VSS 0.031128f
C12374 DVDD.n7318 VSS 0.031128f
C12375 DVDD.n7319 VSS 0.031128f
C12376 DVDD.n7320 VSS 0.031128f
C12377 DVDD.n7322 VSS 0.031128f
C12378 DVDD.n7323 VSS 0.031128f
C12379 DVDD.n7324 VSS 0.031128f
C12380 DVDD.n7325 VSS 0.031128f
C12381 DVDD.n7326 VSS 0.031128f
C12382 DVDD.n7327 VSS 0.031128f
C12383 DVDD.n7328 VSS 0.031128f
C12384 DVDD.n7330 VSS 0.031128f
C12385 DVDD.n7331 VSS 0.031128f
C12386 DVDD.n7332 VSS 0.031128f
C12387 DVDD.n7334 VSS 0.031128f
C12388 DVDD.n7335 VSS 0.031128f
C12389 DVDD.n7336 VSS 0.031128f
C12390 DVDD.n7337 VSS 0.031128f
C12391 DVDD.n7338 VSS 0.031128f
C12392 DVDD.n7339 VSS 0.031128f
C12393 DVDD.n7340 VSS 0.031128f
C12394 DVDD.n7342 VSS 0.031128f
C12395 DVDD.n7343 VSS 0.031128f
C12396 DVDD.n7344 VSS 0.031128f
C12397 DVDD.n7346 VSS 0.031128f
C12398 DVDD.n7347 VSS 0.031128f
C12399 DVDD.n7348 VSS 0.031128f
C12400 DVDD.n7349 VSS 0.031128f
C12401 DVDD.n7350 VSS 0.031128f
C12402 DVDD.n7351 VSS 0.031128f
C12403 DVDD.n7352 VSS 0.031128f
C12404 DVDD.n7354 VSS 0.031128f
C12405 DVDD.n7355 VSS 0.031128f
C12406 DVDD.n7356 VSS 0.031128f
C12407 DVDD.n7358 VSS 0.031128f
C12408 DVDD.n7359 VSS 0.031128f
C12409 DVDD.n7360 VSS 0.031128f
C12410 DVDD.n7361 VSS 0.031128f
C12411 DVDD.n7362 VSS 0.031128f
C12412 DVDD.n7363 VSS 0.031128f
C12413 DVDD.n7364 VSS 0.031128f
C12414 DVDD.n7366 VSS 0.031128f
C12415 DVDD.n7367 VSS 0.031128f
C12416 DVDD.n7368 VSS 0.031128f
C12417 DVDD.n7370 VSS 0.031128f
C12418 DVDD.n7371 VSS 0.031128f
C12419 DVDD.n7372 VSS 0.031128f
C12420 DVDD.n7373 VSS 0.031128f
C12421 DVDD.n7374 VSS 0.031128f
C12422 DVDD.n7375 VSS 0.031128f
C12423 DVDD.n7376 VSS 0.031128f
C12424 DVDD.n7378 VSS 0.031128f
C12425 DVDD.n7379 VSS 0.031128f
C12426 DVDD.n7380 VSS 0.031128f
C12427 DVDD.n7382 VSS 0.031128f
C12428 DVDD.n7383 VSS 0.031128f
C12429 DVDD.n7384 VSS 0.031128f
C12430 DVDD.n7385 VSS 0.031128f
C12431 DVDD.n7386 VSS 0.031128f
C12432 DVDD.n7387 VSS 0.031128f
C12433 DVDD.n7388 VSS 0.031128f
C12434 DVDD.n7390 VSS 0.031128f
C12435 DVDD.n7391 VSS 0.031128f
C12436 DVDD.n7392 VSS 0.031128f
C12437 DVDD.n7394 VSS 0.031128f
C12438 DVDD.n7395 VSS 0.031128f
C12439 DVDD.n7396 VSS 0.031128f
C12440 DVDD.n7397 VSS 0.031128f
C12441 DVDD.n7398 VSS 0.026086f
C12442 DVDD.n7399 VSS 0.031128f
C12443 DVDD.n7400 VSS 0.031128f
C12444 DVDD.n7401 VSS 0.031128f
C12445 DVDD.n7403 VSS 0.019729f
C12446 DVDD.n7404 VSS 0.518041f
C12447 DVDD.n7405 VSS 0.041931f
C12448 DVDD.n7406 VSS 0.041931f
C12449 DVDD.n7407 VSS 0.028833f
C12450 DVDD.n7408 VSS 0.02513f
C12451 DVDD.n7409 VSS 0.02513f
C12452 DVDD.n7410 VSS 0.387477f
C12453 DVDD.n7411 VSS 0.522252f
C12454 DVDD.n7412 VSS 0.598063f
C12455 DVDD.n7454 VSS 0.509617f
C12456 DVDD.n7455 VSS 0.031128f
C12457 DVDD.n7456 VSS 0.063725f
C12458 DVDD.n7457 VSS 0.019729f
C12459 DVDD.n7458 VSS 0.32009f
C12460 DVDD.n7500 VSS 0.509617f
C12461 DVDD.n7501 VSS 0.031128f
C12462 DVDD.n7502 VSS 0.031128f
C12463 DVDD.n7503 VSS 0.031128f
C12464 DVDD.n7504 VSS 0.031128f
C12465 DVDD.n7505 VSS 0.031128f
C12466 DVDD.n7506 VSS 0.031128f
C12467 DVDD.n7507 VSS 0.031128f
C12468 DVDD.n7508 VSS 0.031128f
C12469 DVDD.n7509 VSS 0.031128f
C12470 DVDD.n7510 VSS 0.031128f
C12471 DVDD.n7511 VSS 0.031128f
C12472 DVDD.n7512 VSS 0.031128f
C12473 DVDD.n7513 VSS 0.031128f
C12474 DVDD.n7514 VSS 0.031128f
C12475 DVDD.n7515 VSS 0.031128f
C12476 DVDD.n7516 VSS 0.031128f
C12477 DVDD.n7517 VSS 0.031128f
C12478 DVDD.n7518 VSS 0.031128f
C12479 DVDD.n7519 VSS 0.031128f
C12480 DVDD.n7520 VSS 0.031128f
C12481 DVDD.n7521 VSS 0.031128f
C12482 DVDD.n7522 VSS 0.031128f
C12483 DVDD.n7523 VSS 0.031128f
C12484 DVDD.n7524 VSS 0.031128f
C12485 DVDD.n7525 VSS 0.031128f
C12486 DVDD.n7526 VSS 0.031128f
C12487 DVDD.n7527 VSS 0.031128f
C12488 DVDD.n7528 VSS 0.031128f
C12489 DVDD.n7529 VSS 0.031128f
C12490 DVDD.n7530 VSS 0.031128f
C12491 DVDD.n7531 VSS 0.031128f
C12492 DVDD.n7532 VSS 0.031128f
C12493 DVDD.n7533 VSS 0.031128f
C12494 DVDD.n7534 VSS 0.031128f
C12495 DVDD.n7535 VSS 0.031128f
C12496 DVDD.n7536 VSS 0.031128f
C12497 DVDD.n7537 VSS 0.031128f
C12498 DVDD.n7538 VSS 0.031128f
C12499 DVDD.n7539 VSS 0.031128f
C12500 DVDD.n7540 VSS 0.031128f
C12501 DVDD.n7541 VSS 0.031128f
C12502 DVDD.n7542 VSS 0.031128f
C12503 DVDD.n7543 VSS 0.031128f
C12504 DVDD.n7544 VSS 0.031128f
C12505 DVDD.n7545 VSS 0.031128f
C12506 DVDD.n7546 VSS 0.031128f
C12507 DVDD.n7547 VSS 0.031128f
C12508 DVDD.n7548 VSS 0.031128f
C12509 DVDD.n7549 VSS 0.031128f
C12510 DVDD.n7550 VSS 0.031128f
C12511 DVDD.n7551 VSS 0.031128f
C12512 DVDD.n7552 VSS 0.031128f
C12513 DVDD.n7553 VSS 0.031128f
C12514 DVDD.n7554 VSS 0.031128f
C12515 DVDD.n7555 VSS 0.031128f
C12516 DVDD.n7556 VSS 0.031128f
C12517 DVDD.n7557 VSS 0.031128f
C12518 DVDD.n7558 VSS 0.031128f
C12519 DVDD.n7559 VSS 0.031128f
C12520 DVDD.n7560 VSS 0.031128f
C12521 DVDD.n7561 VSS 0.031128f
C12522 DVDD.n7562 VSS 0.031128f
C12523 DVDD.n7563 VSS 0.053165f
C12524 DVDD.n7564 VSS 0.053165f
C12525 DVDD.n7565 VSS 0.05956f
C12526 DVDD.n7566 VSS 0.05956f
C12527 DVDD.n7567 VSS 0.05956f
C12528 DVDD.n7568 VSS 0.036505f
C12529 DVDD.n7569 VSS 0.522252f
C12530 DVDD.n7611 VSS 0.160045f
C12531 DVDD.n7612 VSS 0.031128f
C12532 DVDD.n7613 VSS 0.033945f
C12533 DVDD.n7614 VSS 0.019729f
C12534 DVDD.n7615 VSS 0.577005f
C12535 DVDD.n7657 VSS 0.084234f
C12536 DVDD.n7658 VSS 0.02513f
C12537 DVDD.n7659 VSS 0.031128f
C12538 DVDD.n7660 VSS 0.031128f
C12539 DVDD.n7661 VSS 0.026086f
C12540 DVDD.n7662 VSS 0.029972f
C12541 DVDD.n7663 VSS 0.041931f
C12542 DVDD.n7664 VSS 0.032925f
C12543 DVDD.n7665 VSS 0.025402f
C12544 DVDD.n7666 VSS 0.029086f
C12545 DVDD.n7667 VSS 0.029086f
C12546 DVDD.n7668 VSS 0.029972f
C12547 DVDD.n7669 VSS 0.041931f
C12548 DVDD.n7670 VSS 0.041931f
C12549 DVDD.n7671 VSS 0.036621f
C12550 DVDD.n7672 VSS 0.026176f
C12551 DVDD.n7673 VSS 0.028833f
C12552 DVDD.n7674 VSS 0.028833f
C12553 DVDD.n7675 VSS 0.02513f
C12554 DVDD.n7676 VSS 0.041931f
C12555 DVDD.n7677 VSS 0.02513f
C12556 DVDD.n7678 VSS 0.14741f
C12557 DVDD.n7679 VSS 0.164257f
C12558 DVDD.n7680 VSS 0.033945f
C12559 DVDD.n7681 VSS 0.05956f
C12560 DVDD.n7682 VSS 0.033945f
C12561 DVDD.n7683 VSS 0.05956f
C12562 DVDD.n7684 VSS 0.039516f
C12563 DVDD.n7685 VSS 0.039516f
C12564 DVDD.n7686 VSS 0.033945f
C12565 DVDD.n7687 VSS 0.033945f
C12566 DVDD.n7688 VSS 0.522252f
C12567 DVDD.n7730 VSS 0.446441f
C12568 DVDD.n7731 VSS 0.031128f
C12569 DVDD.n7732 VSS 0.019729f
C12570 DVDD.n7733 VSS 0.357996f
C12571 DVDD.n7775 VSS 0.37063f
C12572 DVDD.n7776 VSS 0.02513f
C12573 DVDD.n7777 VSS 0.031128f
C12574 DVDD.n7778 VSS 0.031128f
C12575 DVDD.n7779 VSS 0.031128f
C12576 DVDD.n7780 VSS 0.031128f
C12577 DVDD.n7781 VSS 0.031128f
C12578 DVDD.n7782 VSS 0.031128f
C12579 DVDD.n7783 VSS 0.031128f
C12580 DVDD.n7784 VSS 0.031128f
C12581 DVDD.n7785 VSS 0.031128f
C12582 DVDD.n7786 VSS 0.031128f
C12583 DVDD.n7787 VSS 0.031128f
C12584 DVDD.n7788 VSS 0.031128f
C12585 DVDD.n7789 VSS 0.031128f
C12586 DVDD.n7790 VSS 0.031128f
C12587 DVDD.n7791 VSS 0.031128f
C12588 DVDD.n7792 VSS 0.031128f
C12589 DVDD.n7793 VSS 0.031128f
C12590 DVDD.n7794 VSS 0.031128f
C12591 DVDD.n7795 VSS 0.031128f
C12592 DVDD.n7796 VSS 0.031128f
C12593 DVDD.n7797 VSS 0.031128f
C12594 DVDD.n7798 VSS 0.031128f
C12595 DVDD.n7799 VSS 0.031128f
C12596 DVDD.n7800 VSS 0.031128f
C12597 DVDD.n7801 VSS 0.031128f
C12598 DVDD.n7802 VSS 0.031128f
C12599 DVDD.n7803 VSS 0.031128f
C12600 DVDD.n7804 VSS 0.031128f
C12601 DVDD.n7805 VSS 0.031128f
C12602 DVDD.n7806 VSS 0.031128f
C12603 DVDD.n7807 VSS 0.031128f
C12604 DVDD.n7808 VSS 0.031128f
C12605 DVDD.n7809 VSS 0.031128f
C12606 DVDD.n7810 VSS 0.031128f
C12607 DVDD.n7811 VSS 0.031128f
C12608 DVDD.n7812 VSS 0.031128f
C12609 DVDD.n7813 VSS 0.031128f
C12610 DVDD.n7814 VSS 0.031128f
C12611 DVDD.n7815 VSS 0.031128f
C12612 DVDD.n7816 VSS 0.031128f
C12613 DVDD.n7817 VSS 0.031128f
C12614 DVDD.n7818 VSS 0.031128f
C12615 DVDD.n7819 VSS 0.031128f
C12616 DVDD.n7820 VSS 0.031128f
C12617 DVDD.n7821 VSS 0.031128f
C12618 DVDD.n7822 VSS 0.031128f
C12619 DVDD.n7823 VSS 0.031128f
C12620 DVDD.n7824 VSS 0.031128f
C12621 DVDD.n7825 VSS 0.031128f
C12622 DVDD.n7826 VSS 0.031128f
C12623 DVDD.n7827 VSS 0.031128f
C12624 DVDD.n7828 VSS 0.031128f
C12625 DVDD.n7829 VSS 0.031128f
C12626 DVDD.n7830 VSS 0.031128f
C12627 DVDD.n7831 VSS 0.031128f
C12628 DVDD.n7832 VSS 0.031128f
C12629 DVDD.n7833 VSS 0.031128f
C12630 DVDD.n7834 VSS 0.031128f
C12631 DVDD.n7835 VSS 0.031128f
C12632 DVDD.n7836 VSS 0.031128f
C12633 DVDD.n7837 VSS 0.031128f
C12634 DVDD.n7838 VSS 0.031128f
C12635 DVDD.n7839 VSS 0.028497f
C12636 DVDD.n7840 VSS 0.031128f
C12637 DVDD.n7841 VSS 0.031128f
C12638 DVDD.n7842 VSS 0.031128f
C12639 DVDD.n7843 VSS 0.031128f
C12640 DVDD.n7844 VSS 0.031128f
C12641 DVDD.n7845 VSS 0.031128f
C12642 DVDD.n7846 VSS 0.031128f
C12643 DVDD.n7847 VSS 0.031128f
C12644 DVDD.n7848 VSS 0.031128f
C12645 DVDD.n7849 VSS 0.031128f
C12646 DVDD.n7850 VSS 0.031128f
C12647 DVDD.n7851 VSS 0.031128f
C12648 DVDD.n7852 VSS 0.031128f
C12649 DVDD.n7853 VSS 0.031128f
C12650 DVDD.n7854 VSS 0.031128f
C12651 DVDD.n7855 VSS 0.031128f
C12652 DVDD.n7856 VSS 0.031128f
C12653 DVDD.n7857 VSS 0.031128f
C12654 DVDD.n7858 VSS 0.031128f
C12655 DVDD.n7859 VSS 0.031128f
C12656 DVDD.n7860 VSS 0.031128f
C12657 DVDD.n7861 VSS 0.031128f
C12658 DVDD.n7862 VSS 0.031128f
C12659 DVDD.n7863 VSS 0.031128f
C12660 DVDD.n7864 VSS 0.031128f
C12661 DVDD.n7865 VSS 0.031128f
C12662 DVDD.n7866 VSS 0.031128f
C12663 DVDD.n7867 VSS 0.031128f
C12664 DVDD.n7868 VSS 0.031128f
C12665 DVDD.n7869 VSS 0.031128f
C12666 DVDD.n7870 VSS 0.031128f
C12667 DVDD.n7871 VSS 0.031128f
C12668 DVDD.n7872 VSS 0.031128f
C12669 DVDD.n7873 VSS 0.031128f
C12670 DVDD.n7874 VSS 0.031128f
C12671 DVDD.n7875 VSS 0.031128f
C12672 DVDD.n7876 VSS 0.031128f
C12673 DVDD.n7877 VSS 0.031128f
C12674 DVDD.n7878 VSS 0.031128f
C12675 DVDD.n7879 VSS 0.031128f
C12676 DVDD.n7880 VSS 0.031128f
C12677 DVDD.n7881 VSS 0.031128f
C12678 DVDD.n7882 VSS 0.031128f
C12679 DVDD.n7883 VSS 0.031128f
C12680 DVDD.n7884 VSS 0.031128f
C12681 DVDD.n7885 VSS 0.031128f
C12682 DVDD.n7886 VSS 0.031128f
C12683 DVDD.n7887 VSS 0.031128f
C12684 DVDD.n7888 VSS 0.031128f
C12685 DVDD.n7889 VSS 0.031128f
C12686 DVDD.n7890 VSS 0.031128f
C12687 DVDD.n7891 VSS 0.031128f
C12688 DVDD.n7892 VSS 0.031128f
C12689 DVDD.n7893 VSS 0.031128f
C12690 DVDD.n7894 VSS 0.031128f
C12691 DVDD.n7895 VSS 0.031128f
C12692 DVDD.n7896 VSS 0.031128f
C12693 DVDD.n7897 VSS 0.031128f
C12694 DVDD.n7898 VSS 0.031128f
C12695 DVDD.n7899 VSS 0.031128f
C12696 DVDD.n7900 VSS 0.031128f
C12697 DVDD.n7901 VSS 0.031128f
C12698 DVDD.n7902 VSS 0.031128f
C12699 DVDD.n7903 VSS 0.031128f
C12700 DVDD.n7904 VSS 0.031128f
C12701 DVDD.n7905 VSS 0.031128f
C12702 DVDD.n7906 VSS 0.031128f
C12703 DVDD.n7907 VSS 0.031128f
C12704 DVDD.n7908 VSS 0.031128f
C12705 DVDD.n7909 VSS 0.031128f
C12706 DVDD.n7910 VSS 0.031128f
C12707 DVDD.n7911 VSS 0.031128f
C12708 DVDD.n7912 VSS 0.031128f
C12709 DVDD.n7913 VSS 0.031128f
C12710 DVDD.n7914 VSS 0.031128f
C12711 DVDD.n7915 VSS 0.031128f
C12712 DVDD.n7916 VSS 0.031128f
C12713 DVDD.n7917 VSS 0.031128f
C12714 DVDD.n7918 VSS 0.031128f
C12715 DVDD.n7919 VSS 0.031128f
C12716 DVDD.n7920 VSS 0.031128f
C12717 DVDD.n7921 VSS 0.031128f
C12718 DVDD.n7922 VSS 0.031128f
C12719 DVDD.n7923 VSS 0.031128f
C12720 DVDD.n7924 VSS 0.031128f
C12721 DVDD.n7925 VSS 0.031128f
C12722 DVDD.n7926 VSS 0.031128f
C12723 DVDD.n7927 VSS 0.031128f
C12724 DVDD.n7928 VSS 0.031128f
C12725 DVDD.n7929 VSS 0.031128f
C12726 DVDD.n7930 VSS 0.031128f
C12727 DVDD.n7931 VSS 0.031128f
C12728 DVDD.n7932 VSS 0.031128f
C12729 DVDD.n7933 VSS 0.031128f
C12730 DVDD.n7934 VSS 0.031128f
C12731 DVDD.n7935 VSS 0.031128f
C12732 DVDD.n7936 VSS 0.031128f
C12733 DVDD.n7937 VSS 0.031128f
C12734 DVDD.n7938 VSS 0.031128f
C12735 DVDD.n7939 VSS 0.031128f
C12736 DVDD.n7940 VSS 0.031128f
C12737 DVDD.n7941 VSS 0.031128f
C12738 DVDD.n7942 VSS 0.031128f
C12739 DVDD.n7943 VSS 0.031128f
C12740 DVDD.n7944 VSS 0.031128f
C12741 DVDD.n7945 VSS 0.031128f
C12742 DVDD.n7946 VSS 0.031128f
C12743 DVDD.n7947 VSS 0.031128f
C12744 DVDD.n7948 VSS 0.031128f
C12745 DVDD.n7949 VSS 0.031128f
C12746 DVDD.n7950 VSS 0.031128f
C12747 DVDD.n7951 VSS 0.031128f
C12748 DVDD.n7952 VSS 0.031128f
C12749 DVDD.n7953 VSS 0.031128f
C12750 DVDD.n7954 VSS 0.031128f
C12751 DVDD.n7955 VSS 0.031128f
C12752 DVDD.n7956 VSS 0.031128f
C12753 DVDD.n7957 VSS 0.031128f
C12754 DVDD.n7958 VSS 0.031128f
C12755 DVDD.n7959 VSS 0.031128f
C12756 DVDD.n7960 VSS 0.031128f
C12757 DVDD.n7961 VSS 0.031128f
C12758 DVDD.n7962 VSS 0.031128f
C12759 DVDD.n7963 VSS 0.031128f
C12760 DVDD.n7964 VSS 0.031128f
C12761 DVDD.n7965 VSS 0.031128f
C12762 DVDD.n7966 VSS 0.031128f
C12763 DVDD.n7967 VSS 0.031128f
C12764 DVDD.n7968 VSS 0.031128f
C12765 DVDD.n7969 VSS 0.031128f
C12766 DVDD.n7970 VSS 0.031128f
C12767 DVDD.n7971 VSS 0.031128f
C12768 DVDD.n7972 VSS 0.031128f
C12769 DVDD.n7973 VSS 0.031128f
C12770 DVDD.n7974 VSS 0.031128f
C12771 DVDD.n7975 VSS 0.031128f
C12772 DVDD.n7976 VSS 0.031128f
C12773 DVDD.n7977 VSS 0.031128f
C12774 DVDD.n7978 VSS 0.031128f
C12775 DVDD.n7979 VSS 0.031128f
C12776 DVDD.n7980 VSS 0.031128f
C12777 DVDD.n7981 VSS 0.031128f
C12778 DVDD.n7982 VSS 0.031128f
C12779 DVDD.n7983 VSS 0.031128f
C12780 DVDD.n7984 VSS 0.031128f
C12781 DVDD.n7985 VSS 0.031128f
C12782 DVDD.n7986 VSS 0.031128f
C12783 DVDD.n7987 VSS 0.031128f
C12784 DVDD.n7988 VSS 0.031128f
C12785 DVDD.n7989 VSS 0.031128f
C12786 DVDD.n7990 VSS 0.031128f
C12787 DVDD.n7991 VSS 0.031128f
C12788 DVDD.n7992 VSS 0.031128f
C12789 DVDD.n7993 VSS 0.031128f
C12790 DVDD.n7994 VSS 0.031128f
C12791 DVDD.n7995 VSS 0.031128f
C12792 DVDD.n7996 VSS 0.031128f
C12793 DVDD.n7997 VSS 0.031128f
C12794 DVDD.n7998 VSS 0.031128f
C12795 DVDD.n7999 VSS 0.031128f
C12796 DVDD.n8000 VSS 0.031128f
C12797 DVDD.n8001 VSS 0.031128f
C12798 DVDD.n8002 VSS 0.031128f
C12799 DVDD.n8003 VSS 0.031128f
C12800 DVDD.n8004 VSS 0.031128f
C12801 DVDD.n8005 VSS 0.031128f
C12802 DVDD.n8006 VSS 0.031128f
C12803 DVDD.n8007 VSS 0.031128f
C12804 DVDD.n8008 VSS 0.031128f
C12805 DVDD.n8009 VSS 0.031128f
C12806 DVDD.n8010 VSS 0.031128f
C12807 DVDD.n8011 VSS 0.031128f
C12808 DVDD.n8012 VSS 0.031128f
C12809 DVDD.n8013 VSS 0.031128f
C12810 DVDD.n8014 VSS 0.031128f
C12811 DVDD.n8015 VSS 0.031128f
C12812 DVDD.n8016 VSS 0.031128f
C12813 DVDD.n8017 VSS 0.031128f
C12814 DVDD.n8018 VSS 0.031128f
C12815 DVDD.n8019 VSS 0.031128f
C12816 DVDD.n8020 VSS 0.031128f
C12817 DVDD.n8021 VSS 0.031128f
C12818 DVDD.n8022 VSS 0.031128f
C12819 DVDD.n8023 VSS 0.026086f
C12820 DVDD.n8024 VSS 0.022294f
C12821 DVDD.n8025 VSS 0.039421f
C12822 DVDD.n8026 VSS 0.040602f
C12823 DVDD.n8027 VSS 0.032108f
C12824 DVDD.n8028 VSS 0.036763f
C12825 DVDD.n8029 VSS 0.598063f
C12826 DVDD.n8030 VSS 0.505405f
C12827 DVDD.n8031 VSS 0.036763f
C12828 DVDD.n8032 VSS 0.022294f
C12829 DVDD.n8033 VSS 0.041931f
C12830 DVDD.n8034 VSS 0.041931f
C12831 DVDD.n8035 VSS 0.036621f
C12832 DVDD.n8036 VSS 0.019471f
C12833 DVDD.n8037 VSS 0.028833f
C12834 DVDD.n8038 VSS 0.026086f
C12835 DVDD.n8039 VSS 0.036621f
C12836 DVDD.n8040 VSS 0.02513f
C12837 DVDD.n8041 VSS 0.041931f
C12838 DVDD.n8042 VSS 0.02513f
C12839 DVDD.n8043 VSS 0.041931f
C12840 DVDD.n8044 VSS 0.362207f
C12841 DVDD.n8086 VSS 0.019729f
C12842 DVDD.n8087 VSS 0.362207f
C12843 DVDD.n8088 VSS 0.019729f
C12844 DVDD.n8089 VSS 0.522252f
C12845 DVDD.n8090 VSS 0.031128f
C12846 DVDD.n8091 VSS 0.031128f
C12847 DVDD.n8092 VSS 0.031128f
C12848 DVDD.n8093 VSS 0.031128f
C12849 DVDD.n8094 VSS 0.031128f
C12850 DVDD.n8095 VSS 0.031128f
C12851 DVDD.n8096 VSS 0.031128f
C12852 DVDD.n8097 VSS 0.031128f
C12853 DVDD.n8098 VSS 0.031128f
C12854 DVDD.n8099 VSS 0.031128f
C12855 DVDD.n8100 VSS 0.031128f
C12856 DVDD.n8101 VSS 0.031128f
C12857 DVDD.n8102 VSS 0.031128f
C12858 DVDD.n8103 VSS 0.031128f
C12859 DVDD.n8104 VSS 0.031128f
C12860 DVDD.n8105 VSS 0.031128f
C12861 DVDD.n8106 VSS 0.031128f
C12862 DVDD.n8107 VSS 0.031128f
C12863 DVDD.n8108 VSS 0.031128f
C12864 DVDD.n8109 VSS 0.031128f
C12865 DVDD.n8110 VSS 0.031128f
C12866 DVDD.n8111 VSS 0.031128f
C12867 DVDD.n8112 VSS 0.031128f
C12868 DVDD.n8113 VSS 0.031128f
C12869 DVDD.n8114 VSS 0.031128f
C12870 DVDD.n8115 VSS 0.031128f
C12871 DVDD.n8116 VSS 0.031128f
C12872 DVDD.n8117 VSS 0.031128f
C12873 DVDD.n8118 VSS 0.031128f
C12874 DVDD.n8119 VSS 0.031128f
C12875 DVDD.n8120 VSS 0.031128f
C12876 DVDD.n8121 VSS 0.031128f
C12877 DVDD.n8122 VSS 0.031128f
C12878 DVDD.n8123 VSS 0.031128f
C12879 DVDD.n8124 VSS 0.031128f
C12880 DVDD.n8125 VSS 0.031128f
C12881 DVDD.n8126 VSS 0.031128f
C12882 DVDD.n8127 VSS 0.031128f
C12883 DVDD.n8128 VSS 0.031128f
C12884 DVDD.n8129 VSS 0.031128f
C12885 DVDD.n8131 VSS 0.031128f
C12886 DVDD.n8132 VSS 0.031128f
C12887 DVDD.n8133 VSS 0.039516f
C12888 DVDD.n8134 VSS 0.056679f
C12889 DVDD.n8135 VSS 0.05956f
C12890 DVDD.n8136 VSS 0.039387f
C12891 DVDD.n8137 VSS 0.039387f
C12892 DVDD.n8138 VSS 0.035157f
C12893 DVDD.n8139 VSS 0.050592f
C12894 DVDD.n8140 VSS 0.053165f
C12895 DVDD.n8141 VSS 0.05956f
C12896 DVDD.n8142 VSS 0.05956f
C12897 DVDD.n8143 VSS 0.598063f
C12898 DVDD.n8144 VSS 0.039421f
C12899 DVDD.n8145 VSS 0.522252f
C12900 DVDD.n8146 VSS 0.235856f
C12901 DVDD.n8147 VSS 0.056679f
C12902 DVDD.n8148 VSS 0.033945f
C12903 DVDD.n8149 VSS 0.032662f
C12904 DVDD.n8150 VSS 0.030012f
C12905 DVDD.n8151 VSS 0.033623f
C12906 DVDD.n8152 VSS 0.05956f
C12907 DVDD.n8153 VSS 0.033623f
C12908 DVDD.n8154 VSS 0.522252f
C12909 DVDD.n8155 VSS 0.349572f
C12910 DVDD.n8156 VSS 0.02513f
C12911 DVDD.n8157 VSS 0.02513f
C12912 DVDD.n8158 VSS 0.026086f
C12913 DVDD.n8159 VSS 0.036621f
C12914 DVDD.n8160 VSS 0.041931f
C12915 DVDD.n8161 VSS 0.041931f
C12916 DVDD.n8162 VSS 0.484347f
C12917 DVDD.n8204 VSS 0.019729f
C12918 DVDD.n8205 VSS 0.484347f
C12919 DVDD.n8206 VSS 0.019729f
C12920 DVDD.n8207 VSS 0.031128f
C12921 DVDD.n8208 VSS 0.031128f
C12922 DVDD.n8209 VSS 0.031128f
C12923 DVDD.n8210 VSS 0.031128f
C12924 DVDD.n8211 VSS 0.031128f
C12925 DVDD.n8212 VSS 0.031128f
C12926 DVDD.n8213 VSS 0.031128f
C12927 DVDD.n8214 VSS 0.031128f
C12928 DVDD.n8215 VSS 0.031128f
C12929 DVDD.n8216 VSS 0.031128f
C12930 DVDD.n8217 VSS 0.031128f
C12931 DVDD.n8218 VSS 0.031128f
C12932 DVDD.n8219 VSS 0.031128f
C12933 DVDD.n8220 VSS 0.031128f
C12934 DVDD.n8221 VSS 0.031128f
C12935 DVDD.n8222 VSS 0.031128f
C12936 DVDD.n8223 VSS 0.031128f
C12937 DVDD.n8224 VSS 0.031128f
C12938 DVDD.n8225 VSS 0.031128f
C12939 DVDD.n8226 VSS 0.031128f
C12940 DVDD.n8227 VSS 0.031128f
C12941 DVDD.n8228 VSS 0.031128f
C12942 DVDD.n8229 VSS 0.031128f
C12943 DVDD.n8230 VSS 0.031128f
C12944 DVDD.n8231 VSS 0.031128f
C12945 DVDD.n8232 VSS 0.031128f
C12946 DVDD.n8233 VSS 0.031128f
C12947 DVDD.n8234 VSS 0.031128f
C12948 DVDD.n8235 VSS 0.031128f
C12949 DVDD.n8236 VSS 0.031128f
C12950 DVDD.n8237 VSS 0.031128f
C12951 DVDD.n8238 VSS 0.031128f
C12952 DVDD.n8239 VSS 0.031128f
C12953 DVDD.n8240 VSS 0.031128f
C12954 DVDD.n8241 VSS 0.031128f
C12955 DVDD.n8242 VSS 0.031128f
C12956 DVDD.n8243 VSS 0.031128f
C12957 DVDD.n8244 VSS 0.031128f
C12958 DVDD.n8245 VSS 0.031128f
C12959 DVDD.n8246 VSS 0.031128f
C12960 DVDD.n8248 VSS 0.031128f
C12961 DVDD.n8249 VSS 0.031128f
C12962 DVDD.n8250 VSS 0.039516f
C12963 DVDD.n8251 VSS 0.05956f
C12964 DVDD.n8252 VSS 0.033945f
C12965 DVDD.n8253 VSS 0.055718f
C12966 DVDD.n8254 VSS 0.039516f
C12967 DVDD.n8255 VSS 0.033945f
C12968 DVDD.n8256 VSS 0.05956f
C12969 DVDD.n8257 VSS 0.033945f
C12970 DVDD.n8258 VSS 0.122139f
C12971 DVDD.n8259 VSS 0.046329f
C12972 DVDD.n8260 VSS 0.02513f
C12973 DVDD.n8261 VSS 0.041931f
C12974 DVDD.n8262 VSS 0.02513f
C12975 DVDD.n8263 VSS 0.041931f
C12976 DVDD.n8264 VSS 0.031128f
C12977 DVDD.n8265 VSS 0.031128f
C12978 DVDD.n8266 VSS 0.031128f
C12979 DVDD.n8268 VSS 0.031128f
C12980 DVDD.n8269 VSS 0.031128f
C12981 DVDD.n8270 VSS 0.031128f
C12982 DVDD.n8272 VSS 0.031128f
C12983 DVDD.n8273 VSS 0.031128f
C12984 DVDD.n8274 VSS 0.031128f
C12985 DVDD.n8276 VSS 0.031128f
C12986 DVDD.n8277 VSS 0.031128f
C12987 DVDD.n8278 VSS 0.031128f
C12988 DVDD.n8280 VSS 0.031128f
C12989 DVDD.n8281 VSS 0.031128f
C12990 DVDD.n8282 VSS 0.031128f
C12991 DVDD.n8284 VSS 0.031128f
C12992 DVDD.n8285 VSS 0.031128f
C12993 DVDD.n8286 VSS 0.031128f
C12994 DVDD.n8288 VSS 0.031128f
C12995 DVDD.n8289 VSS 0.031128f
C12996 DVDD.n8290 VSS 0.031128f
C12997 DVDD.n8292 VSS 0.031128f
C12998 DVDD.n8293 VSS 0.031128f
C12999 DVDD.n8294 VSS 0.031128f
C13000 DVDD.n8296 VSS 0.031128f
C13001 DVDD.n8297 VSS 0.031128f
C13002 DVDD.n8298 VSS 0.031128f
C13003 DVDD.n8300 VSS 0.031128f
C13004 DVDD.n8301 VSS 0.031128f
C13005 DVDD.n8302 VSS 0.031128f
C13006 DVDD.n8304 VSS 0.031128f
C13007 DVDD.n8305 VSS 0.031128f
C13008 DVDD.n8306 VSS 0.031128f
C13009 DVDD.n8308 VSS 0.031128f
C13010 DVDD.n8309 VSS 0.031128f
C13011 DVDD.n8310 VSS 0.031128f
C13012 DVDD.n8312 VSS 0.031128f
C13013 DVDD.n8313 VSS 0.031128f
C13014 DVDD.n8314 VSS 0.031128f
C13015 DVDD.n8316 VSS 0.031128f
C13016 DVDD.n8317 VSS 0.031128f
C13017 DVDD.n8318 VSS 0.031128f
C13018 DVDD.n8320 VSS 0.031128f
C13019 DVDD.n8321 VSS 0.031128f
C13020 DVDD.n8322 VSS 0.031128f
C13021 DVDD.n8324 VSS 0.031128f
C13022 DVDD.n8325 VSS 0.031128f
C13023 DVDD.n8326 VSS 0.031128f
C13024 DVDD.n8328 VSS 0.031128f
C13025 DVDD.n8329 VSS 0.031128f
C13026 DVDD.n8330 VSS 0.031128f
C13027 DVDD.n8332 VSS 0.031128f
C13028 DVDD.n8333 VSS 0.031128f
C13029 DVDD.n8334 VSS 0.031128f
C13030 DVDD.n8336 VSS 0.031128f
C13031 DVDD.n8337 VSS 0.031128f
C13032 DVDD.n8338 VSS 0.031128f
C13033 DVDD.n8340 VSS 0.031128f
C13034 DVDD.n8341 VSS 0.031128f
C13035 DVDD.n8342 VSS 0.031128f
C13036 DVDD.n8344 VSS 0.031128f
C13037 DVDD.n8345 VSS 0.031128f
C13038 DVDD.n8346 VSS 0.031128f
C13039 DVDD.n8347 VSS 0.028497f
C13040 DVDD.n8348 VSS 0.019729f
C13041 DVDD.n8349 VSS 0.019729f
C13042 DVDD.n8351 VSS 0.031128f
C13043 DVDD.n8353 VSS 0.031128f
C13044 DVDD.n8355 VSS 0.031128f
C13045 DVDD.n8356 VSS 0.031128f
C13046 DVDD.n8357 VSS 0.031128f
C13047 DVDD.n8358 VSS 0.031128f
C13048 DVDD.n8359 VSS 0.031128f
C13049 DVDD.n8360 VSS 0.031128f
C13050 DVDD.n8361 VSS 0.031128f
C13051 DVDD.n8363 VSS 0.031128f
C13052 DVDD.n8365 VSS 0.031128f
C13053 DVDD.n8367 VSS 0.031128f
C13054 DVDD.n8368 VSS 0.031128f
C13055 DVDD.n8369 VSS 0.031128f
C13056 DVDD.n8370 VSS 0.031128f
C13057 DVDD.n8371 VSS 0.031128f
C13058 DVDD.n8372 VSS 0.031128f
C13059 DVDD.n8373 VSS 0.031128f
C13060 DVDD.n8375 VSS 0.031128f
C13061 DVDD.n8377 VSS 0.031128f
C13062 DVDD.n8379 VSS 0.031128f
C13063 DVDD.n8380 VSS 0.031128f
C13064 DVDD.n8381 VSS 0.031128f
C13065 DVDD.n8382 VSS 0.031128f
C13066 DVDD.n8383 VSS 0.031128f
C13067 DVDD.n8384 VSS 0.031128f
C13068 DVDD.n8385 VSS 0.031128f
C13069 DVDD.n8387 VSS 0.031128f
C13070 DVDD.n8389 VSS 0.031128f
C13071 DVDD.n8391 VSS 0.031128f
C13072 DVDD.n8392 VSS 0.031128f
C13073 DVDD.n8393 VSS 0.031128f
C13074 DVDD.n8394 VSS 0.031128f
C13075 DVDD.n8395 VSS 0.031128f
C13076 DVDD.n8396 VSS 0.031128f
C13077 DVDD.n8397 VSS 0.031128f
C13078 DVDD.n8399 VSS 0.031128f
C13079 DVDD.n8401 VSS 0.031128f
C13080 DVDD.n8403 VSS 0.031128f
C13081 DVDD.n8404 VSS 0.031128f
C13082 DVDD.n8405 VSS 0.031128f
C13083 DVDD.n8406 VSS 0.031128f
C13084 DVDD.n8407 VSS 0.031128f
C13085 DVDD.n8408 VSS 0.031128f
C13086 DVDD.n8409 VSS 0.031128f
C13087 DVDD.n8411 VSS 0.031128f
C13088 DVDD.n8413 VSS 0.031128f
C13089 DVDD.n8415 VSS 0.031128f
C13090 DVDD.n8416 VSS 0.031128f
C13091 DVDD.n8417 VSS 0.031128f
C13092 DVDD.n8418 VSS 0.031128f
C13093 DVDD.n8419 VSS 0.031128f
C13094 DVDD.n8420 VSS 0.031128f
C13095 DVDD.n8421 VSS 0.031128f
C13096 DVDD.n8423 VSS 0.031128f
C13097 DVDD.n8425 VSS 0.031128f
C13098 DVDD.n8427 VSS 0.031128f
C13099 DVDD.n8428 VSS 0.031128f
C13100 DVDD.n8429 VSS 0.031128f
C13101 DVDD.n8430 VSS 0.031128f
C13102 DVDD.n8431 VSS 0.031128f
C13103 DVDD.n8432 VSS 0.031128f
C13104 DVDD.n8433 VSS 0.031128f
C13105 DVDD.n8435 VSS 0.031128f
C13106 DVDD.n8437 VSS 0.031128f
C13107 DVDD.n8439 VSS 0.031128f
C13108 DVDD.n8440 VSS 0.031128f
C13109 DVDD.n8441 VSS 0.031128f
C13110 DVDD.n8442 VSS 0.031128f
C13111 DVDD.n8443 VSS 0.031128f
C13112 DVDD.n8444 VSS 0.031128f
C13113 DVDD.n8445 VSS 0.031128f
C13114 DVDD.n8447 VSS 0.031128f
C13115 DVDD.n8449 VSS 0.031128f
C13116 DVDD.n8451 VSS 0.031128f
C13117 DVDD.n8452 VSS 0.031128f
C13118 DVDD.n8453 VSS 0.031128f
C13119 DVDD.n8454 VSS 0.031128f
C13120 DVDD.n8455 VSS 0.031128f
C13121 DVDD.n8456 VSS 0.031128f
C13122 DVDD.n8457 VSS 0.031128f
C13123 DVDD.n8459 VSS 0.031128f
C13124 DVDD.n8461 VSS 0.031128f
C13125 DVDD.n8463 VSS 0.031128f
C13126 DVDD.n8464 VSS 0.031128f
C13127 DVDD.n8465 VSS 0.031128f
C13128 DVDD.n8466 VSS 0.031128f
C13129 DVDD.n8467 VSS 0.031128f
C13130 DVDD.n8468 VSS 0.031128f
C13131 DVDD.n8469 VSS 0.031128f
C13132 DVDD.n8471 VSS 0.031128f
C13133 DVDD.n8473 VSS 0.031128f
C13134 DVDD.n8475 VSS 0.031128f
C13135 DVDD.n8476 VSS 0.031128f
C13136 DVDD.n8477 VSS 0.031128f
C13137 DVDD.n8478 VSS 0.031128f
C13138 DVDD.n8479 VSS 0.031128f
C13139 DVDD.n8480 VSS 0.031128f
C13140 DVDD.n8481 VSS 0.031128f
C13141 DVDD.n8483 VSS 0.031128f
C13142 DVDD.n8485 VSS 0.031128f
C13143 DVDD.n8487 VSS 0.031128f
C13144 DVDD.n8488 VSS 0.031128f
C13145 DVDD.n8489 VSS 0.031128f
C13146 DVDD.n8490 VSS 0.031128f
C13147 DVDD.n8491 VSS 0.031128f
C13148 DVDD.n8492 VSS 0.031128f
C13149 DVDD.n8493 VSS 0.031128f
C13150 DVDD.n8495 VSS 0.031128f
C13151 DVDD.n8497 VSS 0.031128f
C13152 DVDD.n8499 VSS 0.031128f
C13153 DVDD.n8500 VSS 0.031128f
C13154 DVDD.n8501 VSS 0.031128f
C13155 DVDD.n8502 VSS 0.031128f
C13156 DVDD.n8503 VSS 0.031128f
C13157 DVDD.n8504 VSS 0.031128f
C13158 DVDD.n8505 VSS 0.031128f
C13159 DVDD.n8507 VSS 0.031128f
C13160 DVDD.n8509 VSS 0.031128f
C13161 DVDD.n8511 VSS 0.031128f
C13162 DVDD.n8512 VSS 0.031128f
C13163 DVDD.n8513 VSS 0.031128f
C13164 DVDD.n8514 VSS 0.031128f
C13165 DVDD.n8515 VSS 0.031128f
C13166 DVDD.n8516 VSS 0.031128f
C13167 DVDD.n8517 VSS 0.031128f
C13168 DVDD.n8519 VSS 0.031128f
C13169 DVDD.n8521 VSS 0.031128f
C13170 DVDD.n8523 VSS 0.031128f
C13171 DVDD.n8524 VSS 0.031128f
C13172 DVDD.n8525 VSS 0.031128f
C13173 DVDD.n8526 VSS 0.031128f
C13174 DVDD.n8527 VSS 0.031128f
C13175 DVDD.n8528 VSS 0.031128f
C13176 DVDD.n8529 VSS 0.031128f
C13177 DVDD.n8531 VSS 0.031128f
C13178 DVDD.n8533 VSS 0.031128f
C13179 DVDD.n8535 VSS 0.031128f
C13180 DVDD.n8536 VSS 0.031128f
C13181 DVDD.n8537 VSS 0.031128f
C13182 DVDD.n8538 VSS 0.031128f
C13183 DVDD.n8539 VSS 0.031128f
C13184 DVDD.n8540 VSS 0.031128f
C13185 DVDD.n8541 VSS 0.031128f
C13186 DVDD.n8543 VSS 0.031128f
C13187 DVDD.n8545 VSS 0.031128f
C13188 DVDD.n8547 VSS 0.031128f
C13189 DVDD.n8548 VSS 0.031128f
C13190 DVDD.n8549 VSS 0.031128f
C13191 DVDD.n8550 VSS 0.031128f
C13192 DVDD.n8551 VSS 0.031128f
C13193 DVDD.n8552 VSS 0.031128f
C13194 DVDD.n8553 VSS 0.031128f
C13195 DVDD.n8555 VSS 0.031128f
C13196 DVDD.n8557 VSS 0.031128f
C13197 DVDD.n8559 VSS 0.031128f
C13198 DVDD.n8560 VSS 0.031128f
C13199 DVDD.n8561 VSS 0.031128f
C13200 DVDD.n8562 VSS 0.031128f
C13201 DVDD.n8563 VSS 0.031128f
C13202 DVDD.n8564 VSS 0.031128f
C13203 DVDD.n8565 VSS 0.031128f
C13204 DVDD.n8567 VSS 0.031128f
C13205 DVDD.n8569 VSS 0.031128f
C13206 DVDD.n8571 VSS 0.031128f
C13207 DVDD.n8572 VSS 0.031128f
C13208 DVDD.n8573 VSS 0.031128f
C13209 DVDD.n8574 VSS 0.031128f
C13210 DVDD.n8575 VSS 0.031128f
C13211 DVDD.n8576 VSS 0.031128f
C13212 DVDD.n8577 VSS 0.031128f
C13213 DVDD.n8579 VSS 0.031128f
C13214 DVDD.n8581 VSS 0.031128f
C13215 DVDD.n8583 VSS 0.031128f
C13216 DVDD.n8584 VSS 0.031128f
C13217 DVDD.n8585 VSS 0.031128f
C13218 DVDD.n8586 VSS 0.031128f
C13219 DVDD.n8587 VSS 0.031128f
C13220 DVDD.n8588 VSS 0.031128f
C13221 DVDD.n8589 VSS 0.031128f
C13222 DVDD.n8590 VSS 0.031128f
C13223 DVDD.n8592 VSS 0.031128f
C13224 DVDD.n8594 VSS 0.031128f
C13225 DVDD.n8596 VSS 0.019729f
C13226 DVDD.n8597 VSS 0.019729f
C13227 DVDD.n8598 VSS 0.026086f
C13228 DVDD.n8599 VSS 0.522252f
C13229 DVDD.n8600 VSS 0.598063f
C13230 DVDD.n8601 VSS 0.404324f
C13231 DVDD.n8602 VSS 0.031743f
C13232 DVDD.n8603 VSS 0.031743f
C13233 DVDD.n8604 VSS 0.027723f
C13234 DVDD.n8605 VSS 0.028833f
C13235 DVDD.n8606 VSS 0.028833f
C13236 DVDD.n8607 VSS 0.02513f
C13237 DVDD.n8608 VSS 0.02513f
C13238 DVDD.n8609 VSS 0.105293f
C13239 DVDD.n8610 VSS 0.181104f
C13240 DVDD.n8611 VSS 0.033945f
C13241 DVDD.n8612 VSS 0.05956f
C13242 DVDD.n8613 VSS 0.033945f
C13243 DVDD.n8614 VSS 0.05956f
C13244 DVDD.n8615 VSS 0.031128f
C13245 DVDD.n8616 VSS 0.031128f
C13246 DVDD.n8618 VSS 0.031128f
C13247 DVDD.n8619 VSS 0.031128f
C13248 DVDD.n8620 VSS 0.031128f
C13249 DVDD.n8621 VSS 0.031128f
C13250 DVDD.n8624 VSS 0.031128f
C13251 DVDD.n8625 VSS 0.031128f
C13252 DVDD.n8626 VSS 0.031128f
C13253 DVDD.n8627 VSS 0.031128f
C13254 DVDD.n8630 VSS 0.031128f
C13255 DVDD.n8631 VSS 0.031128f
C13256 DVDD.n8632 VSS 0.031128f
C13257 DVDD.n8633 VSS 0.031128f
C13258 DVDD.n8636 VSS 0.031128f
C13259 DVDD.n8637 VSS 0.031128f
C13260 DVDD.n8638 VSS 0.031128f
C13261 DVDD.n8639 VSS 0.031128f
C13262 DVDD.n8642 VSS 0.031128f
C13263 DVDD.n8643 VSS 0.031128f
C13264 DVDD.n8644 VSS 0.031128f
C13265 DVDD.n8645 VSS 0.031128f
C13266 DVDD.n8648 VSS 0.031128f
C13267 DVDD.n8649 VSS 0.031128f
C13268 DVDD.n8650 VSS 0.031128f
C13269 DVDD.n8651 VSS 0.031128f
C13270 DVDD.n8654 VSS 0.031128f
C13271 DVDD.n8655 VSS 0.031128f
C13272 DVDD.n8656 VSS 0.031128f
C13273 DVDD.n8657 VSS 0.031128f
C13274 DVDD.n8660 VSS 0.031128f
C13275 DVDD.n8661 VSS 0.031128f
C13276 DVDD.n8662 VSS 0.031128f
C13277 DVDD.n8663 VSS 0.031128f
C13278 DVDD.n8666 VSS 0.031128f
C13279 DVDD.n8667 VSS 0.031128f
C13280 DVDD.n8668 VSS 0.031128f
C13281 DVDD.n8669 VSS 0.031128f
C13282 DVDD.n8672 VSS 0.031128f
C13283 DVDD.n8673 VSS 0.031128f
C13284 DVDD.n8674 VSS 0.031128f
C13285 DVDD.n8675 VSS 0.031128f
C13286 DVDD.n8678 VSS 0.031128f
C13287 DVDD.n8679 VSS 0.031128f
C13288 DVDD.n8680 VSS 0.031128f
C13289 DVDD.n8681 VSS 0.031128f
C13290 DVDD.n8684 VSS 0.031128f
C13291 DVDD.n8685 VSS 0.031128f
C13292 DVDD.n8686 VSS 0.031128f
C13293 DVDD.n8687 VSS 0.031128f
C13294 DVDD.n8690 VSS 0.031128f
C13295 DVDD.n8691 VSS 0.031128f
C13296 DVDD.n8692 VSS 0.031128f
C13297 DVDD.n8693 VSS 0.031128f
C13298 DVDD.n8696 VSS 0.031128f
C13299 DVDD.n8697 VSS 0.031128f
C13300 DVDD.n8698 VSS 0.031128f
C13301 DVDD.n8699 VSS 0.031128f
C13302 DVDD.n8702 VSS 0.031128f
C13303 DVDD.n8703 VSS 0.031128f
C13304 DVDD.n8704 VSS 0.031128f
C13305 DVDD.n8705 VSS 0.031128f
C13306 DVDD.n8708 VSS 0.031128f
C13307 DVDD.n8709 VSS 0.031128f
C13308 DVDD.n8710 VSS 0.031128f
C13309 DVDD.n8711 VSS 0.031128f
C13310 DVDD.n8714 VSS 0.031128f
C13311 DVDD.n8715 VSS 0.031128f
C13312 DVDD.n8716 VSS 0.031128f
C13313 DVDD.n8717 VSS 0.031128f
C13314 DVDD.n8720 VSS 0.031128f
C13315 DVDD.n8721 VSS 0.031128f
C13316 DVDD.n8722 VSS 0.031128f
C13317 DVDD.n8723 VSS 0.031128f
C13318 DVDD.n8726 VSS 0.031128f
C13319 DVDD.n8727 VSS 0.031128f
C13320 DVDD.n8728 VSS 0.031128f
C13321 DVDD.n8729 VSS 0.031128f
C13322 DVDD.n8732 VSS 0.031128f
C13323 DVDD.n8733 VSS 0.031128f
C13324 DVDD.n8734 VSS 0.031128f
C13325 DVDD.n8735 VSS 0.031128f
C13326 DVDD.n8738 VSS 0.019729f
C13327 DVDD.n8739 VSS 0.019729f
C13328 DVDD.n8740 VSS 0.026086f
C13329 DVDD.n8741 VSS 0.031128f
C13330 DVDD.n8742 VSS 0.031128f
C13331 DVDD.n8743 VSS 0.031128f
C13332 DVDD.n8745 VSS 0.031128f
C13333 DVDD.n8747 VSS 0.031128f
C13334 DVDD.n8748 VSS 0.031128f
C13335 DVDD.n8749 VSS 0.031128f
C13336 DVDD.n8750 VSS 0.031128f
C13337 DVDD.n8751 VSS 0.031128f
C13338 DVDD.n8752 VSS 0.031128f
C13339 DVDD.n8753 VSS 0.031128f
C13340 DVDD.n8755 VSS 0.031128f
C13341 DVDD.n8757 VSS 0.031128f
C13342 DVDD.n8758 VSS 0.031128f
C13343 DVDD.n8759 VSS 0.031128f
C13344 DVDD.n8760 VSS 0.031128f
C13345 DVDD.n8761 VSS 0.031128f
C13346 DVDD.n8762 VSS 0.031128f
C13347 DVDD.n8763 VSS 0.031128f
C13348 DVDD.n8765 VSS 0.031128f
C13349 DVDD.n8767 VSS 0.031128f
C13350 DVDD.n8768 VSS 0.031128f
C13351 DVDD.n8769 VSS 0.031128f
C13352 DVDD.n8770 VSS 0.031128f
C13353 DVDD.n8771 VSS 0.031128f
C13354 DVDD.n8772 VSS 0.031128f
C13355 DVDD.n8773 VSS 0.031128f
C13356 DVDD.n8775 VSS 0.031128f
C13357 DVDD.n8777 VSS 0.031128f
C13358 DVDD.n8778 VSS 0.031128f
C13359 DVDD.n8779 VSS 0.031128f
C13360 DVDD.n8780 VSS 0.031128f
C13361 DVDD.n8781 VSS 0.031128f
C13362 DVDD.n8782 VSS 0.031128f
C13363 DVDD.n8783 VSS 0.031128f
C13364 DVDD.n8785 VSS 0.031128f
C13365 DVDD.n8787 VSS 0.031128f
C13366 DVDD.n8788 VSS 0.031128f
C13367 DVDD.n8789 VSS 0.031128f
C13368 DVDD.n8790 VSS 0.031128f
C13369 DVDD.n8791 VSS 0.031128f
C13370 DVDD.n8792 VSS 0.031128f
C13371 DVDD.n8793 VSS 0.031128f
C13372 DVDD.n8795 VSS 0.031128f
C13373 DVDD.n8797 VSS 0.031128f
C13374 DVDD.n8798 VSS 0.031128f
C13375 DVDD.n8799 VSS 0.031128f
C13376 DVDD.n8800 VSS 0.031128f
C13377 DVDD.n8801 VSS 0.031128f
C13378 DVDD.n8802 VSS 0.031128f
C13379 DVDD.n8803 VSS 0.031128f
C13380 DVDD.n8805 VSS 0.031128f
C13381 DVDD.n8807 VSS 0.031128f
C13382 DVDD.n8808 VSS 0.031128f
C13383 DVDD.n8809 VSS 0.031128f
C13384 DVDD.n8810 VSS 0.031128f
C13385 DVDD.n8811 VSS 0.031128f
C13386 DVDD.n8812 VSS 0.031128f
C13387 DVDD.n8813 VSS 0.031128f
C13388 DVDD.n8815 VSS 0.031128f
C13389 DVDD.n8817 VSS 0.031128f
C13390 DVDD.n8818 VSS 0.031128f
C13391 DVDD.n8819 VSS 0.031128f
C13392 DVDD.n8820 VSS 0.031128f
C13393 DVDD.n8821 VSS 0.031128f
C13394 DVDD.n8822 VSS 0.031128f
C13395 DVDD.n8823 VSS 0.031128f
C13396 DVDD.n8825 VSS 0.031128f
C13397 DVDD.n8827 VSS 0.031128f
C13398 DVDD.n8828 VSS 0.031128f
C13399 DVDD.n8829 VSS 0.031128f
C13400 DVDD.n8830 VSS 0.031128f
C13401 DVDD.n8831 VSS 0.031128f
C13402 DVDD.n8832 VSS 0.031128f
C13403 DVDD.n8833 VSS 0.031128f
C13404 DVDD.n8835 VSS 0.031128f
C13405 DVDD.n8837 VSS 0.031128f
C13406 DVDD.n8838 VSS 0.031128f
C13407 DVDD.n8839 VSS 0.031128f
C13408 DVDD.n8840 VSS 0.031128f
C13409 DVDD.n8841 VSS 0.031128f
C13410 DVDD.n8842 VSS 0.031128f
C13411 DVDD.n8843 VSS 0.031128f
C13412 DVDD.n8845 VSS 0.031128f
C13413 DVDD.n8847 VSS 0.031128f
C13414 DVDD.n8848 VSS 0.031128f
C13415 DVDD.n8849 VSS 0.031128f
C13416 DVDD.n8850 VSS 0.031128f
C13417 DVDD.n8851 VSS 0.031128f
C13418 DVDD.n8852 VSS 0.031128f
C13419 DVDD.n8853 VSS 0.031128f
C13420 DVDD.n8855 VSS 0.031128f
C13421 DVDD.n8857 VSS 0.031128f
C13422 DVDD.n8858 VSS 0.031128f
C13423 DVDD.n8859 VSS 0.031128f
C13424 DVDD.n8860 VSS 0.031128f
C13425 DVDD.n8861 VSS 0.031128f
C13426 DVDD.n8862 VSS 0.031128f
C13427 DVDD.n8863 VSS 0.031128f
C13428 DVDD.n8865 VSS 0.031128f
C13429 DVDD.n8867 VSS 0.031128f
C13430 DVDD.n8868 VSS 0.031128f
C13431 DVDD.n8869 VSS 0.031128f
C13432 DVDD.n8870 VSS 0.031128f
C13433 DVDD.n8871 VSS 0.031128f
C13434 DVDD.n8872 VSS 0.031128f
C13435 DVDD.n8873 VSS 0.031128f
C13436 DVDD.n8875 VSS 0.031128f
C13437 DVDD.n8877 VSS 0.031128f
C13438 DVDD.n8878 VSS 0.031128f
C13439 DVDD.n8879 VSS 0.031128f
C13440 DVDD.n8880 VSS 0.031128f
C13441 DVDD.n8881 VSS 0.031128f
C13442 DVDD.n8882 VSS 0.031128f
C13443 DVDD.n8883 VSS 0.031128f
C13444 DVDD.n8885 VSS 0.031128f
C13445 DVDD.n8887 VSS 0.031128f
C13446 DVDD.n8888 VSS 0.031128f
C13447 DVDD.n8889 VSS 0.031128f
C13448 DVDD.n8890 VSS 0.031128f
C13449 DVDD.n8891 VSS 0.031128f
C13450 DVDD.n8892 VSS 0.031128f
C13451 DVDD.n8893 VSS 0.031128f
C13452 DVDD.n8895 VSS 0.031128f
C13453 DVDD.n8897 VSS 0.031128f
C13454 DVDD.n8898 VSS 0.031128f
C13455 DVDD.n8899 VSS 0.031128f
C13456 DVDD.n8900 VSS 0.031128f
C13457 DVDD.n8901 VSS 0.031128f
C13458 DVDD.n8902 VSS 0.031128f
C13459 DVDD.n8903 VSS 0.031128f
C13460 DVDD.n8905 VSS 0.031128f
C13461 DVDD.n8907 VSS 0.031128f
C13462 DVDD.n8908 VSS 0.031128f
C13463 DVDD.n8909 VSS 0.031128f
C13464 DVDD.n8910 VSS 0.031128f
C13465 DVDD.n8911 VSS 0.031128f
C13466 DVDD.n8912 VSS 0.031128f
C13467 DVDD.n8913 VSS 0.031128f
C13468 DVDD.n8915 VSS 0.031128f
C13469 DVDD.n8917 VSS 0.031128f
C13470 DVDD.n8918 VSS 0.031128f
C13471 DVDD.n8919 VSS 0.031128f
C13472 DVDD.n8920 VSS 0.031128f
C13473 DVDD.n8921 VSS 0.031128f
C13474 DVDD.n8922 VSS 0.031128f
C13475 DVDD.n8923 VSS 0.031128f
C13476 DVDD.n8925 VSS 0.031128f
C13477 DVDD.n8927 VSS 0.031128f
C13478 DVDD.n8928 VSS 0.031128f
C13479 DVDD.n8929 VSS 0.031128f
C13480 DVDD.n8930 VSS 0.031128f
C13481 DVDD.n8931 VSS 0.031128f
C13482 DVDD.n8932 VSS 0.031128f
C13483 DVDD.n8933 VSS 0.031128f
C13484 DVDD.n8935 VSS 0.031128f
C13485 DVDD.n8937 VSS 0.031128f
C13486 DVDD.n8938 VSS 0.031128f
C13487 DVDD.n8939 VSS 0.031128f
C13488 DVDD.n8940 VSS 0.031128f
C13489 DVDD.n8941 VSS 0.031128f
C13490 DVDD.n8942 VSS 0.031128f
C13491 DVDD.n8943 VSS 0.031128f
C13492 DVDD.n8945 VSS 0.031128f
C13493 DVDD.n8947 VSS 0.019729f
C13494 DVDD.n8948 VSS 0.019729f
C13495 DVDD.n8949 VSS 0.028497f
C13496 DVDD.n8959 VSS 0.025624f
C13497 DVDD.n8960 VSS 0.142744f
C13498 DVDD.n8961 VSS 0.025624f
C13499 DVDD.n8962 VSS 1.04547f
C13500 DVDD.n8964 VSS 0.025624f
C13501 DVDD.n8965 VSS 0.025624f
C13502 DVDD.n8966 VSS 0.025624f
C13503 DVDD.n8967 VSS 0.025624f
C13504 DVDD.n8968 VSS 0.025624f
C13505 DVDD.n8969 VSS 0.025624f
C13506 DVDD.n8970 VSS 0.025624f
C13507 DVDD.n8971 VSS 0.025624f
C13508 DVDD.n8972 VSS 0.142744f
C13509 DVDD.n8974 VSS 0.040945f
C13510 DVDD.n8975 VSS 0.031128f
C13511 DVDD.n8976 VSS 0.031128f
C13512 DVDD.n8977 VSS 0.031128f
C13513 DVDD.n8978 VSS 0.031128f
C13514 DVDD.n8979 VSS 0.031128f
C13515 DVDD.n8980 VSS 0.031128f
C13516 DVDD.n8981 VSS 0.031128f
C13517 DVDD.n8982 VSS 0.031128f
C13518 DVDD.n8983 VSS 0.031128f
C13519 DVDD.n8984 VSS 0.031128f
C13520 DVDD.n8985 VSS 0.031128f
C13521 DVDD.n8986 VSS 0.031128f
C13522 DVDD.n8987 VSS 0.031128f
C13523 DVDD.n8988 VSS 0.031128f
C13524 DVDD.n8989 VSS 0.031128f
C13525 DVDD.n8990 VSS 0.031128f
C13526 DVDD.n8991 VSS 0.031128f
C13527 DVDD.n8992 VSS 0.031128f
C13528 DVDD.n8993 VSS 0.031128f
C13529 DVDD.n8994 VSS 0.031128f
C13530 DVDD.n8995 VSS 0.031128f
C13531 DVDD.n8996 VSS 0.031128f
C13532 DVDD.n8997 VSS 0.031128f
C13533 DVDD.n8998 VSS 0.031128f
C13534 DVDD.n8999 VSS 0.031128f
C13535 DVDD.n9000 VSS 0.031128f
C13536 DVDD.n9001 VSS 0.031128f
C13537 DVDD.n9002 VSS 0.031128f
C13538 DVDD.n9003 VSS 0.031128f
C13539 DVDD.n9004 VSS 0.031128f
C13540 DVDD.n9005 VSS 0.031128f
C13541 DVDD.n9006 VSS 0.031128f
C13542 DVDD.n9007 VSS 0.031128f
C13543 DVDD.n9008 VSS 0.031128f
C13544 DVDD.n9009 VSS 0.031128f
C13545 DVDD.n9010 VSS 0.031128f
C13546 DVDD.n9011 VSS 0.031128f
C13547 DVDD.n9012 VSS 0.031128f
C13548 DVDD.n9013 VSS 0.031128f
C13549 DVDD.n9014 VSS 0.031128f
C13550 DVDD.n9015 VSS 0.031128f
C13551 DVDD.n9016 VSS 0.031128f
C13552 DVDD.n9017 VSS 0.031128f
C13553 DVDD.n9018 VSS 0.031128f
C13554 DVDD.n9019 VSS 0.031128f
C13555 DVDD.n9020 VSS 0.031128f
C13556 DVDD.n9021 VSS 0.031128f
C13557 DVDD.n9022 VSS 0.031128f
C13558 DVDD.n9023 VSS 0.031128f
C13559 DVDD.n9024 VSS 0.031128f
C13560 DVDD.n9025 VSS 0.031128f
C13561 DVDD.n9026 VSS 0.031128f
C13562 DVDD.n9027 VSS 0.031128f
C13563 DVDD.n9028 VSS 0.031128f
C13564 DVDD.n9029 VSS 0.031128f
C13565 DVDD.n9030 VSS 0.031128f
C13566 DVDD.n9031 VSS 0.031128f
C13567 DVDD.n9032 VSS 0.031128f
C13568 DVDD.n9033 VSS 0.031128f
C13569 DVDD.n9034 VSS 0.031128f
C13570 DVDD.n9035 VSS 0.031128f
C13571 DVDD.n9036 VSS 0.031128f
C13572 DVDD.n9037 VSS 0.031128f
C13573 DVDD.n9038 VSS 0.031128f
C13574 DVDD.n9039 VSS 0.031128f
C13575 DVDD.n9040 VSS 0.031128f
C13576 DVDD.n9041 VSS 0.031128f
C13577 DVDD.n9042 VSS 0.031128f
C13578 DVDD.n9043 VSS 0.031128f
C13579 DVDD.n9044 VSS 0.031128f
C13580 DVDD.n9045 VSS 0.031128f
C13581 DVDD.n9046 VSS 0.031128f
C13582 DVDD.n9047 VSS 0.031128f
C13583 DVDD.n9048 VSS 0.031128f
C13584 DVDD.n9049 VSS 0.031128f
C13585 DVDD.n9050 VSS 0.031128f
C13586 DVDD.n9051 VSS 0.031128f
C13587 DVDD.n9052 VSS 0.031128f
C13588 DVDD.n9053 VSS 0.031128f
C13589 DVDD.n9054 VSS 0.031128f
C13590 DVDD.n9055 VSS 0.031128f
C13591 DVDD.n9056 VSS 0.031128f
C13592 DVDD.n9057 VSS 0.031128f
C13593 DVDD.n9058 VSS 0.031128f
C13594 DVDD.n9059 VSS 0.031128f
C13595 DVDD.n9060 VSS 0.031128f
C13596 DVDD.n9061 VSS 0.031128f
C13597 DVDD.n9062 VSS 0.031128f
C13598 DVDD.n9063 VSS 0.031128f
C13599 DVDD.n9064 VSS 0.031128f
C13600 DVDD.n9065 VSS 0.031128f
C13601 DVDD.n9066 VSS 0.031128f
C13602 DVDD.n9067 VSS 0.031128f
C13603 DVDD.n9068 VSS 0.031128f
C13604 DVDD.n9069 VSS 0.031128f
C13605 DVDD.n9070 VSS 0.031128f
C13606 DVDD.n9071 VSS 0.031128f
C13607 DVDD.n9072 VSS 0.031128f
C13608 DVDD.n9073 VSS 0.031128f
C13609 DVDD.n9074 VSS 0.031128f
C13610 DVDD.n9075 VSS 0.031128f
C13611 DVDD.n9076 VSS 0.031128f
C13612 DVDD.n9077 VSS 0.031128f
C13613 DVDD.n9078 VSS 0.031128f
C13614 DVDD.n9079 VSS 0.031128f
C13615 DVDD.n9080 VSS 0.031128f
C13616 DVDD.n9081 VSS 0.031128f
C13617 DVDD.n9082 VSS 0.031128f
C13618 DVDD.n9083 VSS 0.031128f
C13619 DVDD.n9084 VSS 0.031128f
C13620 DVDD.n9085 VSS 0.031128f
C13621 DVDD.n9086 VSS 0.031128f
C13622 DVDD.n9087 VSS 0.031128f
C13623 DVDD.n9088 VSS 0.031128f
C13624 DVDD.n9089 VSS 0.031128f
C13625 DVDD.n9090 VSS 0.031128f
C13626 DVDD.n9091 VSS 0.031128f
C13627 DVDD.n9092 VSS 0.031128f
C13628 DVDD.n9093 VSS 0.031128f
C13629 DVDD.n9094 VSS 0.031128f
C13630 DVDD.n9095 VSS 0.031128f
C13631 DVDD.n9096 VSS 0.031128f
C13632 DVDD.n9097 VSS 0.031128f
C13633 DVDD.n9098 VSS 0.031128f
C13634 DVDD.n9099 VSS 0.031128f
C13635 DVDD.n9100 VSS 0.031128f
C13636 DVDD.n9101 VSS 0.031128f
C13637 DVDD.n9102 VSS 0.031128f
C13638 DVDD.n9103 VSS 0.031128f
C13639 DVDD.n9104 VSS 0.031128f
C13640 DVDD.n9105 VSS 0.031128f
C13641 DVDD.n9106 VSS 0.031128f
C13642 DVDD.n9107 VSS 0.031128f
C13643 DVDD.n9108 VSS 0.031128f
C13644 DVDD.n9109 VSS 0.031128f
C13645 DVDD.n9110 VSS 0.031128f
C13646 DVDD.n9111 VSS 0.031128f
C13647 DVDD.n9112 VSS 0.031128f
C13648 DVDD.n9113 VSS 0.031128f
C13649 DVDD.n9114 VSS 0.031128f
C13650 DVDD.n9115 VSS 0.031128f
C13651 DVDD.n9116 VSS 0.031128f
C13652 DVDD.n9117 VSS 0.031128f
C13653 DVDD.n9118 VSS 0.031128f
C13654 DVDD.n9119 VSS 0.031128f
C13655 DVDD.n9120 VSS 0.031128f
C13656 DVDD.n9121 VSS 0.031128f
C13657 DVDD.n9122 VSS 0.031128f
C13658 DVDD.n9123 VSS 0.031128f
C13659 DVDD.n9124 VSS 0.031128f
C13660 DVDD.n9125 VSS 0.031128f
C13661 DVDD.n9126 VSS 0.031128f
C13662 DVDD.n9127 VSS 0.031128f
C13663 DVDD.n9128 VSS 0.031128f
C13664 DVDD.n9129 VSS 0.031128f
C13665 DVDD.n9130 VSS 0.031128f
C13666 DVDD.n9131 VSS 0.031128f
C13667 DVDD.n9132 VSS 0.031128f
C13668 DVDD.n9133 VSS 0.031128f
C13669 DVDD.n9134 VSS 0.031128f
C13670 DVDD.n9135 VSS 0.031128f
C13671 DVDD.n9136 VSS 0.031128f
C13672 DVDD.n9137 VSS 0.031128f
C13673 DVDD.n9138 VSS 0.031128f
C13674 DVDD.n9139 VSS 0.031128f
C13675 DVDD.n9140 VSS 0.031128f
C13676 DVDD.n9141 VSS 0.031128f
C13677 DVDD.n9142 VSS 0.031128f
C13678 DVDD.n9143 VSS 0.031128f
C13679 DVDD.n9144 VSS 0.031128f
C13680 DVDD.n9145 VSS 0.031128f
C13681 DVDD.n9146 VSS 0.031128f
C13682 DVDD.n9147 VSS 0.031128f
C13683 DVDD.n9148 VSS 0.031128f
C13684 DVDD.n9149 VSS 0.031128f
C13685 DVDD.n9150 VSS 0.031128f
C13686 DVDD.n9151 VSS 0.031128f
C13687 DVDD.n9152 VSS 0.031128f
C13688 DVDD.n9153 VSS 0.031128f
C13689 DVDD.n9154 VSS 0.031128f
C13690 DVDD.n9155 VSS 0.031128f
C13691 DVDD.n9156 VSS 0.031128f
C13692 DVDD.n9157 VSS 0.031128f
C13693 DVDD.n9158 VSS 0.031128f
C13694 DVDD.n9159 VSS 0.031128f
C13695 DVDD.n9160 VSS 0.031128f
C13696 DVDD.n9161 VSS 0.031128f
C13697 DVDD.n9162 VSS 0.031128f
C13698 DVDD.n9163 VSS 0.031128f
C13699 DVDD.n9164 VSS 0.031128f
C13700 DVDD.n9165 VSS 0.031128f
C13701 DVDD.n9166 VSS 0.031128f
C13702 DVDD.n9167 VSS 0.031128f
C13703 DVDD.n9168 VSS 0.031128f
C13704 DVDD.n9169 VSS 0.031128f
C13705 DVDD.n9170 VSS 0.031128f
C13706 DVDD.n9171 VSS 0.031128f
C13707 DVDD.n9172 VSS 0.031128f
C13708 DVDD.n9173 VSS 0.031128f
C13709 DVDD.n9174 VSS 0.031128f
C13710 DVDD.n9175 VSS 0.031128f
C13711 DVDD.n9176 VSS 0.031128f
C13712 DVDD.n9177 VSS 0.031128f
C13713 DVDD.n9178 VSS 0.031128f
C13714 DVDD.n9179 VSS 0.031128f
C13715 DVDD.n9180 VSS 0.031128f
C13716 DVDD.n9181 VSS 0.031128f
C13717 DVDD.n9182 VSS 0.031128f
C13718 DVDD.n9183 VSS 0.031128f
C13719 DVDD.n9184 VSS 0.031128f
C13720 DVDD.n9185 VSS 0.031128f
C13721 DVDD.n9186 VSS 0.031128f
C13722 DVDD.n9187 VSS 0.031128f
C13723 DVDD.n9188 VSS 0.031128f
C13724 DVDD.n9189 VSS 0.031128f
C13725 DVDD.n9190 VSS 0.031128f
C13726 DVDD.n9191 VSS 0.031128f
C13727 DVDD.n9192 VSS 0.031128f
C13728 DVDD.n9193 VSS 0.031128f
C13729 DVDD.n9194 VSS 0.031128f
C13730 DVDD.n9195 VSS 0.031128f
C13731 DVDD.n9196 VSS 0.031128f
C13732 DVDD.n9197 VSS 0.031128f
C13733 DVDD.n9198 VSS 0.031128f
C13734 DVDD.n9199 VSS 0.031128f
C13735 DVDD.n9200 VSS 0.031128f
C13736 DVDD.n9201 VSS 0.031128f
C13737 DVDD.n9202 VSS 0.031128f
C13738 DVDD.n9203 VSS 0.031128f
C13739 DVDD.n9204 VSS 0.031128f
C13740 DVDD.n9205 VSS 0.031128f
C13741 DVDD.n9206 VSS 0.031128f
C13742 DVDD.n9207 VSS 0.031128f
C13743 DVDD.n9208 VSS 0.031128f
C13744 DVDD.n9209 VSS 0.031128f
C13745 DVDD.n9210 VSS 0.031128f
C13746 DVDD.n9211 VSS 0.031128f
C13747 DVDD.n9212 VSS 0.031128f
C13748 DVDD.n9213 VSS 0.031128f
C13749 DVDD.n9214 VSS 0.031128f
C13750 DVDD.n9215 VSS 0.031128f
C13751 DVDD.n9216 VSS 0.031128f
C13752 DVDD.n9217 VSS 0.031128f
C13753 DVDD.n9218 VSS 0.028497f
C13754 DVDD.n9219 VSS 0.039516f
C13755 DVDD.n9220 VSS 0.05956f
C13756 DVDD.n9221 VSS 0.052836f
C13757 DVDD.n9222 VSS 0.585428f
C13758 DVDD.n9264 VSS 0.031128f
C13759 DVDD.n9265 VSS 0.028497f
C13760 DVDD.n9267 VSS 0.031128f
C13761 DVDD.n9268 VSS 0.031128f
C13762 DVDD.n9269 VSS 0.031128f
C13763 DVDD.n9270 VSS 0.031128f
C13764 DVDD.n9271 VSS 0.031128f
C13765 DVDD.n9272 VSS 0.031128f
C13766 DVDD.n9273 VSS 0.031128f
C13767 DVDD.n9274 VSS 0.031128f
C13768 DVDD.n9275 VSS 0.031128f
C13769 DVDD.n9276 VSS 0.031128f
C13770 DVDD.n9277 VSS 0.031128f
C13771 DVDD.n9278 VSS 0.031128f
C13772 DVDD.n9279 VSS 0.031128f
C13773 DVDD.n9280 VSS 0.031128f
C13774 DVDD.n9281 VSS 0.031128f
C13775 DVDD.n9282 VSS 0.031128f
C13776 DVDD.n9283 VSS 0.031128f
C13777 DVDD.n9284 VSS 0.031128f
C13778 DVDD.n9285 VSS 0.031128f
C13779 DVDD.n9286 VSS 0.031128f
C13780 DVDD.n9287 VSS 0.031128f
C13781 DVDD.n9288 VSS 0.031128f
C13782 DVDD.n9289 VSS 0.031128f
C13783 DVDD.n9290 VSS 0.031128f
C13784 DVDD.n9291 VSS 0.031128f
C13785 DVDD.n9292 VSS 0.031128f
C13786 DVDD.n9293 VSS 0.031128f
C13787 DVDD.n9294 VSS 0.031128f
C13788 DVDD.n9295 VSS 0.031128f
C13789 DVDD.n9296 VSS 0.031128f
C13790 DVDD.n9297 VSS 0.031128f
C13791 DVDD.n9298 VSS 0.031128f
C13792 DVDD.n9299 VSS 0.031128f
C13793 DVDD.n9300 VSS 0.031128f
C13794 DVDD.n9301 VSS 0.031128f
C13795 DVDD.n9302 VSS 0.031128f
C13796 DVDD.n9303 VSS 0.031128f
C13797 DVDD.n9304 VSS 0.031128f
C13798 DVDD.n9305 VSS 0.031128f
C13799 DVDD.n9306 VSS 0.031128f
C13800 DVDD.n9307 VSS 0.031128f
C13801 DVDD.n9308 VSS 0.031128f
C13802 DVDD.n9309 VSS 0.019729f
C13803 DVDD.n9310 VSS 0.019729f
C13804 DVDD.n9311 VSS 0.026086f
C13805 DVDD.n9312 VSS 0.031128f
C13806 DVDD.n9313 VSS 0.031128f
C13807 DVDD.n9314 VSS 0.031128f
C13808 DVDD.n9316 VSS 0.031128f
C13809 DVDD.n9317 VSS 0.031128f
C13810 DVDD.n9318 VSS 0.031128f
C13811 DVDD.n9319 VSS 0.031128f
C13812 DVDD.n9321 VSS 0.031128f
C13813 DVDD.n9322 VSS 0.031128f
C13814 DVDD.n9323 VSS 0.031128f
C13815 DVDD.n9324 VSS 0.031128f
C13816 DVDD.n9325 VSS 0.031128f
C13817 DVDD.n9326 VSS 0.031128f
C13818 DVDD.n9328 VSS 0.031128f
C13819 DVDD.n9329 VSS 0.031128f
C13820 DVDD.n9330 VSS 0.031128f
C13821 DVDD.n9331 VSS 0.031128f
C13822 DVDD.n9333 VSS 0.031128f
C13823 DVDD.n9334 VSS 0.031128f
C13824 DVDD.n9335 VSS 0.031128f
C13825 DVDD.n9336 VSS 0.031128f
C13826 DVDD.n9337 VSS 0.031128f
C13827 DVDD.n9338 VSS 0.031128f
C13828 DVDD.n9340 VSS 0.031128f
C13829 DVDD.n9341 VSS 0.031128f
C13830 DVDD.n9342 VSS 0.031128f
C13831 DVDD.n9343 VSS 0.031128f
C13832 DVDD.n9345 VSS 0.031128f
C13833 DVDD.n9346 VSS 0.031128f
C13834 DVDD.n9347 VSS 0.031128f
C13835 DVDD.n9348 VSS 0.031128f
C13836 DVDD.n9349 VSS 0.031128f
C13837 DVDD.n9350 VSS 0.031128f
C13838 DVDD.n9352 VSS 0.031128f
C13839 DVDD.n9353 VSS 0.031128f
C13840 DVDD.n9354 VSS 0.031128f
C13841 DVDD.n9355 VSS 0.031128f
C13842 DVDD.n9357 VSS 0.031128f
C13843 DVDD.n9358 VSS 0.031128f
C13844 DVDD.n9359 VSS 0.031128f
C13845 DVDD.n9360 VSS 0.031128f
C13846 DVDD.n9361 VSS 0.031128f
C13847 DVDD.n9362 VSS 0.031128f
C13848 DVDD.n9364 VSS 0.031128f
C13849 DVDD.n9365 VSS 0.031128f
C13850 DVDD.n9366 VSS 0.031128f
C13851 DVDD.n9367 VSS 0.031128f
C13852 DVDD.n9369 VSS 0.031128f
C13853 DVDD.n9370 VSS 0.031128f
C13854 DVDD.n9371 VSS 0.031128f
C13855 DVDD.n9372 VSS 0.031128f
C13856 DVDD.n9373 VSS 0.031128f
C13857 DVDD.n9374 VSS 0.031128f
C13858 DVDD.n9376 VSS 0.031128f
C13859 DVDD.n9377 VSS 0.031128f
C13860 DVDD.n9378 VSS 0.031128f
C13861 DVDD.n9379 VSS 0.031128f
C13862 DVDD.n9381 VSS 0.031128f
C13863 DVDD.n9382 VSS 0.031128f
C13864 DVDD.n9383 VSS 0.031128f
C13865 DVDD.n9384 VSS 0.031128f
C13866 DVDD.n9385 VSS 0.031128f
C13867 DVDD.n9386 VSS 0.031128f
C13868 DVDD.n9388 VSS 0.031128f
C13869 DVDD.n9389 VSS 0.031128f
C13870 DVDD.n9390 VSS 0.031128f
C13871 DVDD.n9391 VSS 0.031128f
C13872 DVDD.n9393 VSS 0.031128f
C13873 DVDD.n9394 VSS 0.031128f
C13874 DVDD.n9395 VSS 0.031128f
C13875 DVDD.n9396 VSS 0.031128f
C13876 DVDD.n9397 VSS 0.031128f
C13877 DVDD.n9398 VSS 0.031128f
C13878 DVDD.n9400 VSS 0.031128f
C13879 DVDD.n9401 VSS 0.031128f
C13880 DVDD.n9402 VSS 0.031128f
C13881 DVDD.n9403 VSS 0.031128f
C13882 DVDD.n9405 VSS 0.031128f
C13883 DVDD.n9406 VSS 0.031128f
C13884 DVDD.n9407 VSS 0.031128f
C13885 DVDD.n9408 VSS 0.031128f
C13886 DVDD.n9409 VSS 0.031128f
C13887 DVDD.n9410 VSS 0.031128f
C13888 DVDD.n9412 VSS 0.031128f
C13889 DVDD.n9413 VSS 0.031128f
C13890 DVDD.n9414 VSS 0.031128f
C13891 DVDD.n9415 VSS 0.031128f
C13892 DVDD.n9417 VSS 0.031128f
C13893 DVDD.n9418 VSS 0.031128f
C13894 DVDD.n9419 VSS 0.031128f
C13895 DVDD.n9420 VSS 0.031128f
C13896 DVDD.n9421 VSS 0.031128f
C13897 DVDD.n9422 VSS 0.031128f
C13898 DVDD.n9424 VSS 0.031128f
C13899 DVDD.n9425 VSS 0.031128f
C13900 DVDD.n9426 VSS 0.031128f
C13901 DVDD.n9427 VSS 0.031128f
C13902 DVDD.n9429 VSS 0.031128f
C13903 DVDD.n9430 VSS 0.031128f
C13904 DVDD.n9431 VSS 0.031128f
C13905 DVDD.n9432 VSS 0.031128f
C13906 DVDD.n9433 VSS 0.031128f
C13907 DVDD.n9434 VSS 0.031128f
C13908 DVDD.n9436 VSS 0.031128f
C13909 DVDD.n9437 VSS 0.031128f
C13910 DVDD.n9438 VSS 0.031128f
C13911 DVDD.n9439 VSS 0.031128f
C13912 DVDD.n9441 VSS 0.031128f
C13913 DVDD.n9442 VSS 0.031128f
C13914 DVDD.n9443 VSS 0.031128f
C13915 DVDD.n9444 VSS 0.031128f
C13916 DVDD.n9445 VSS 0.031128f
C13917 DVDD.n9446 VSS 0.031128f
C13918 DVDD.n9448 VSS 0.031128f
C13919 DVDD.n9449 VSS 0.031128f
C13920 DVDD.n9450 VSS 0.031128f
C13921 DVDD.n9451 VSS 0.031128f
C13922 DVDD.n9453 VSS 0.031128f
C13923 DVDD.n9454 VSS 0.031128f
C13924 DVDD.n9455 VSS 0.031128f
C13925 DVDD.n9456 VSS 0.031128f
C13926 DVDD.n9457 VSS 0.031128f
C13927 DVDD.n9458 VSS 0.031128f
C13928 DVDD.n9460 VSS 0.031128f
C13929 DVDD.n9461 VSS 0.031128f
C13930 DVDD.n9462 VSS 0.031128f
C13931 DVDD.n9463 VSS 0.031128f
C13932 DVDD.n9465 VSS 0.031128f
C13933 DVDD.n9466 VSS 0.031128f
C13934 DVDD.n9467 VSS 0.031128f
C13935 DVDD.n9468 VSS 0.031128f
C13936 DVDD.n9469 VSS 0.031128f
C13937 DVDD.n9470 VSS 0.031128f
C13938 DVDD.n9472 VSS 0.031128f
C13939 DVDD.n9473 VSS 0.031128f
C13940 DVDD.n9474 VSS 0.031128f
C13941 DVDD.n9475 VSS 0.031128f
C13942 DVDD.n9477 VSS 0.031128f
C13943 DVDD.n9478 VSS 0.031128f
C13944 DVDD.n9479 VSS 0.031128f
C13945 DVDD.n9480 VSS 0.031128f
C13946 DVDD.n9481 VSS 0.031128f
C13947 DVDD.n9482 VSS 0.031128f
C13948 DVDD.n9484 VSS 0.031128f
C13949 DVDD.n9485 VSS 0.031128f
C13950 DVDD.n9486 VSS 0.031128f
C13951 DVDD.n9487 VSS 0.031128f
C13952 DVDD.n9489 VSS 0.031128f
C13953 DVDD.n9490 VSS 0.031128f
C13954 DVDD.n9491 VSS 0.031128f
C13955 DVDD.n9492 VSS 0.031128f
C13956 DVDD.n9493 VSS 0.031128f
C13957 DVDD.n9494 VSS 0.031128f
C13958 DVDD.n9496 VSS 0.031128f
C13959 DVDD.n9497 VSS 0.031128f
C13960 DVDD.n9498 VSS 0.031128f
C13961 DVDD.n9499 VSS 0.031128f
C13962 DVDD.n9501 VSS 0.031128f
C13963 DVDD.n9502 VSS 0.031128f
C13964 DVDD.n9503 VSS 0.031128f
C13965 DVDD.n9504 VSS 0.031128f
C13966 DVDD.n9505 VSS 0.031128f
C13967 DVDD.n9506 VSS 0.031128f
C13968 DVDD.n9508 VSS 0.031128f
C13969 DVDD.n9509 VSS 0.031128f
C13970 DVDD.n9510 VSS 0.031128f
C13971 DVDD.n9511 VSS 0.031128f
C13972 DVDD.n9513 VSS 0.031128f
C13973 DVDD.n9514 VSS 0.031128f
C13974 DVDD.n9515 VSS 0.031128f
C13975 DVDD.n9516 VSS 0.031128f
C13976 DVDD.n9517 VSS 0.031128f
C13977 DVDD.n9518 VSS 0.031128f
C13978 DVDD.n9520 VSS 0.031128f
C13979 DVDD.n9521 VSS 0.031128f
C13980 DVDD.n9522 VSS 0.031128f
C13981 DVDD.n9523 VSS 0.031128f
C13982 DVDD.n9525 VSS 0.031128f
C13983 DVDD.n9526 VSS 0.031128f
C13984 DVDD.n9527 VSS 0.031128f
C13985 DVDD.n9528 VSS 0.031128f
C13986 DVDD.n9529 VSS 0.031128f
C13987 DVDD.n9530 VSS 0.031128f
C13988 DVDD.n9532 VSS 0.031128f
C13989 DVDD.n9533 VSS 0.031128f
C13990 DVDD.n9534 VSS 0.031128f
C13991 DVDD.n9535 VSS 0.031128f
C13992 DVDD.n9537 VSS 0.031128f
C13993 DVDD.n9538 VSS 0.031128f
C13994 DVDD.n9539 VSS 0.031128f
C13995 DVDD.n9540 VSS 0.031128f
C13996 DVDD.n9541 VSS 0.031128f
C13997 DVDD.n9542 VSS 0.031128f
C13998 DVDD.n9544 VSS 0.031128f
C13999 DVDD.n9545 VSS 0.031128f
C14000 DVDD.n9546 VSS 0.031128f
C14001 DVDD.n9547 VSS 0.031128f
C14002 DVDD.n9549 VSS 0.031128f
C14003 DVDD.n9550 VSS 0.031128f
C14004 DVDD.n9551 VSS 0.031128f
C14005 DVDD.n9552 VSS 0.031128f
C14006 DVDD.n9553 VSS 0.031128f
C14007 DVDD.n9554 VSS 0.031128f
C14008 DVDD.n9555 VSS 0.019729f
C14009 DVDD.n9556 VSS 0.019729f
C14010 DVDD.n9558 VSS 0.509617f
C14011 DVDD.n9559 VSS 0.463288f
C14012 DVDD.n9560 VSS 0.534888f
C14013 DVDD.n9561 VSS 0.05956f
C14014 DVDD.n9562 VSS 0.043229f
C14015 DVDD.n9563 VSS 0.043229f
C14016 DVDD.n9564 VSS 0.038587f
C14017 DVDD.n9565 VSS 0.053165f
C14018 DVDD.n9566 VSS 0.047162f
C14019 DVDD.n9567 VSS 0.052836f
C14020 DVDD.n9568 VSS 0.033945f
C14021 DVDD.n9569 VSS 0.036505f
C14022 DVDD.n9570 VSS 0.018221f
C14023 DVDD.n9571 VSS 0.423753f
C14024 DVDD.n9572 VSS 0.468543f
C14025 DVDD.n9573 VSS 0.761343f
C14026 DVDD.t123 VSS 0.167631f
C14027 DVDD.t144 VSS 0.167631f
C14028 DVDD.n9574 VSS 0.335261f
C14029 DVDD.n9575 VSS 0.644991f
C14030 DVDD.n9576 VSS 0.761767f
C14031 DVDD.n9577 VSS 0.644991f
C14032 DVDD.n9578 VSS 0.761767f
C14033 DVDD.n9579 VSS 0.761343f
C14034 DVDD.t81 VSS 0.167631f
C14035 DVDD.t143 VSS 0.167631f
C14036 DVDD.n9580 VSS 0.335261f
C14037 DVDD.n9581 VSS 0.644991f
C14038 DVDD.n9582 VSS 0.098809f
C14039 DVDD.n9583 VSS 0.761767f
C14040 DVDD.n9584 VSS 0.761767f
C14041 DVDD.n9585 VSS 0.644991f
C14042 DVDD.n9586 VSS 0.761767f
C14043 DVDD.n9587 VSS 0.761343f
C14044 DVDD.t75 VSS 0.167631f
C14045 DVDD.t116 VSS 0.167631f
C14046 DVDD.n9588 VSS 0.335261f
C14047 DVDD.n9589 VSS 0.644991f
C14048 DVDD.n9590 VSS 0.098809f
C14049 DVDD.n9591 VSS 0.761767f
C14050 DVDD.n9592 VSS 0.761767f
C14051 DVDD.n9593 VSS 0.97806f
C14052 DVDD.n9594 VSS 0.761767f
C14053 DVDD.n9595 VSS 1.09441f
C14054 DVDD.t99 VSS 0.425324f
C14055 DVDD.n9596 VSS 0.644991f
C14056 DVDD.n9597 VSS 0.098809f
C14057 DVDD.n9598 VSS 1.09484f
C14058 DVDD.n9599 VSS 1.09484f
C14059 DVDD.n9600 VSS 0.644991f
C14060 DVDD.n9601 VSS 0.761767f
C14061 DVDD.n9602 VSS 0.761343f
C14062 DVDD.t80 VSS 0.167631f
C14063 DVDD.t121 VSS 0.167631f
C14064 DVDD.n9603 VSS 0.335261f
C14065 DVDD.n9604 VSS 0.644991f
C14066 DVDD.n9605 VSS 0.098809f
C14067 DVDD.n9606 VSS 0.761767f
C14068 DVDD.n9607 VSS 0.761767f
C14069 DVDD.n9608 VSS 0.581549f
C14070 DVDD.n9609 VSS 0.761767f
C14071 DVDD.n9610 VSS 0.322495f
C14072 DVDD.t131 VSS 0.167631f
C14073 DVDD.t98 VSS 0.167631f
C14074 DVDD.n9611 VSS 0.335261f
C14075 DVDD.n9612 VSS 0.081946f
C14076 DVDD.n9613 VSS 0.064086f
C14077 DVDD.n9615 VSS 0.064086f
C14078 DVDD.n9616 VSS 0.064086f
C14079 DVDD.n9617 VSS 0.064086f
C14080 DVDD.n9619 VSS 0.064086f
C14081 DVDD.n9620 VSS 0.064086f
C14082 DVDD.n9621 VSS 0.064086f
C14083 DVDD.n9622 VSS 0.064086f
C14084 DVDD.n9623 VSS 0.064086f
C14085 DVDD.n9624 VSS 0.064086f
C14086 DVDD.n9625 VSS 0.064086f
C14087 DVDD.n9626 VSS 0.055963f
C14088 DVDD.n9627 VSS 0.105736f
C14089 DVDD.n9628 VSS 0.293418f
C14090 DVDD.n9629 VSS 0.163891f
C14091 DVDD.n9630 VSS 0.1401f
C14092 DVDD.n9631 VSS 0.163891f
C14093 DVDD.n9632 VSS 0.093873f
C14094 DVDD.n9634 VSS 0.163891f
C14095 DVDD.n9636 VSS 0.163891f
C14096 DVDD.n9637 VSS 0.134814f
C14097 DVDD.n9639 VSS 0.111023f
C14098 DVDD.n9641 VSS 0.060476f
C14099 DVDD.n9642 VSS 0.059573f
C14100 DVDD.n9643 VSS 0.055963f
C14101 DVDD.n9644 VSS 0.128173f
C14102 DVDD.n9648 VSS 0.061379f
C14103 DVDD.n9649 VSS 0.055963f
C14104 DVDD.n9650 VSS 0.128173f
C14105 DVDD.n9651 VSS 0.128173f
C14106 DVDD.n9652 VSS 0.128173f
C14107 DVDD.n9653 VSS 0.128173f
C14108 DVDD.n9654 VSS 0.128173f
C14109 DVDD.n9655 VSS 0.128173f
C14110 DVDD.n9656 VSS 0.128173f
C14111 DVDD.n9657 VSS 0.095678f
C14112 DVDD.n9658 VSS 0.128173f
C14113 DVDD.n9659 VSS 0.128173f
C14114 DVDD.n9660 VSS 0.128173f
C14115 DVDD.n9661 VSS 0.064086f
C14116 DVDD.n9662 VSS 0.105736f
C14117 DVDD.n9663 VSS 0.293418f
C14118 DVDD.n9664 VSS 0.163891f
C14119 DVDD.n9665 VSS 0.1401f
C14120 DVDD.n9666 VSS 0.163891f
C14121 DVDD.n9667 VSS 0.055963f
C14122 DVDD.n9668 VSS 0.322495f
C14123 DVDD.n9670 VSS 0.163891f
C14124 DVDD.n9672 VSS 0.163891f
C14125 DVDD.n9674 VSS 0.134814f
C14126 DVDD.n9676 VSS 0.111023f
C14127 DVDD.n9680 VSS 0.064086f
C14128 DVDD.n9681 VSS 0.057768f
C14129 DVDD.n9682 VSS 0.064086f
C14130 DVDD.n9683 VSS 0.064086f
C14131 DVDD.n9684 VSS 0.064086f
C14132 DVDD.n9685 VSS 0.056865f
C14133 DVDD.n9686 VSS 0.064086f
C14134 DVDD.n9687 VSS 0.081946f
C14135 DVDD.n9689 VSS 0.063184f
C14136 DVDD.n9690 VSS 0.064086f
C14137 DVDD.n9691 VSS 0.064086f
C14138 DVDD.n9692 VSS 0.064086f
C14139 DVDD.n9694 VSS 0.062281f
C14140 DVDD.n9695 VSS 0.064086f
C14141 DVDD.n9696 VSS 0.055963f
C14142 DVDD.n9697 VSS 0.128173f
C14143 DVDD.n9698 VSS 0.128173f
C14144 DVDD.n9699 VSS 0.128173f
C14145 DVDD.n9700 VSS 0.128173f
C14146 DVDD.n9701 VSS 0.055963f
C14147 DVDD.n9702 VSS 0.128173f
C14148 DVDD.n9703 VSS 0.128173f
C14149 DVDD.n9704 VSS 0.055963f
C14150 DVDD.n9705 VSS 0.128173f
C14151 DVDD.n9706 VSS 0.128173f
C14152 DVDD.n9707 VSS 0.055963f
C14153 DVDD.n9708 VSS 0.128173f
C14154 DVDD.n9709 VSS 0.055963f
C14155 DVDD.n9710 VSS 0.128173f
C14156 DVDD.n9711 VSS 0.128173f
C14157 DVDD.n9712 VSS 0.128173f
C14158 DVDD.n9713 VSS 0.128173f
C14159 DVDD.n9714 VSS 0.055963f
C14160 DVDD.n9715 VSS 0.128173f
C14161 DVDD.n9716 VSS 0.055963f
C14162 DVDD.n9717 VSS 0.128173f
C14163 DVDD.n9718 VSS 0.055963f
C14164 DVDD.n9719 VSS 0.128173f
C14165 DVDD.n9720 VSS 0.128173f
C14166 DVDD.n9721 VSS 0.128173f
C14167 DVDD.n9722 VSS 0.128173f
C14168 DVDD.n9723 VSS 0.055963f
C14169 DVDD.n9724 VSS 0.128173f
C14170 DVDD.n9725 VSS 0.055963f
C14171 DVDD.n9726 VSS 0.128173f
C14172 DVDD.n9727 VSS 0.055963f
C14173 DVDD.n9728 VSS 0.128173f
C14174 DVDD.n9729 VSS 0.128173f
C14175 DVDD.n9730 VSS 0.128173f
C14176 DVDD.n9731 VSS 0.128173f
C14177 DVDD.n9732 VSS 0.128173f
C14178 DVDD.n9733 VSS 0.105736f
C14179 DVDD.n9734 VSS 0.293418f
C14180 DVDD.n9735 VSS 0.163891f
C14181 DVDD.n9736 VSS 0.1401f
C14182 DVDD.n9737 VSS 0.163891f
C14183 DVDD.n9738 VSS 0.055963f
C14184 DVDD.n9739 VSS 0.098809f
C14185 DVDD.n9740 VSS 0.698325f
C14186 DVDD.n9741 VSS 0.322495f
C14187 DVDD.n9742 VSS 0.163891f
C14188 DVDD.n9743 VSS 0.163891f
C14189 DVDD.n9744 VSS 0.134814f
C14190 DVDD.n9745 VSS 0.111023f
C14191 DVDD.n9750 VSS 0.064086f
C14192 DVDD.n9751 VSS 0.061379f
C14193 DVDD.n9752 VSS 0.064086f
C14194 DVDD.n9753 VSS 0.064086f
C14195 DVDD.n9754 VSS 0.064086f
C14196 DVDD.n9755 VSS 0.060476f
C14197 DVDD.n9757 VSS 0.057768f
C14198 DVDD.n9758 VSS 0.064086f
C14199 DVDD.n9759 VSS 0.064086f
C14200 DVDD.n9760 VSS 0.056865f
C14201 DVDD.n9761 VSS 0.064086f
C14202 DVDD.n9762 VSS 0.064086f
C14203 DVDD.n9763 VSS 0.064086f
C14204 DVDD.n9764 VSS 0.064086f
C14205 DVDD.n9765 VSS 0.064086f
C14206 DVDD.n9767 VSS 0.063184f
C14207 DVDD.n9768 VSS 0.064086f
C14208 DVDD.n9769 VSS 0.064086f
C14209 DVDD.n9770 VSS 0.064086f
C14210 DVDD.n9772 VSS 0.062281f
C14211 DVDD.n9773 VSS 0.055963f
C14212 DVDD.n9774 VSS 0.105736f
C14213 DVDD.n9775 VSS 1.09441f
C14214 DVDD.t103 VSS 0.167631f
C14215 DVDD.t84 VSS 0.167631f
C14216 DVDD.n9776 VSS 0.335261f
C14217 DVDD.n9778 VSS 0.183717f
C14218 DVDD.n9779 VSS 0.757335f
C14219 DVDD.n9780 VSS 1.09484f
C14220 DVDD.n9781 VSS 0.874112f
C14221 DVDD.n9782 VSS 0.873688f
C14222 DVDD.n9783 VSS 0.099098f
C14223 DVDD.t100 VSS 0.425324f
C14224 DVDD.n9784 VSS 0.098809f
C14225 DVDD.n9785 VSS 0.757335f
C14226 DVDD.n9786 VSS 0.650744f
C14227 DVDD.n9787 VSS 0.098809f
C14228 DVDD.n9788 VSS 0.533968f
C14229 DVDD.n9789 VSS 0.97806f
C14230 DVDD.n9790 VSS 0.098809f
C14231 DVDD.t77 VSS 0.425324f
C14232 DVDD.n9791 VSS 0.099098f
C14233 DVDD.n9792 VSS 0.97806f
C14234 DVDD.n9793 VSS 0.533968f
C14235 DVDD.n9794 VSS 0.099098f
C14236 DVDD.n9795 VSS 0.65032f
C14237 DVDD.n9796 VSS 0.293418f
C14238 DVDD.n9797 VSS 0.163891f
C14239 DVDD.n9798 VSS 0.198722f
C14240 DVDD.n9799 VSS 0.081946f
C14241 DVDD.n9800 VSS 0.098809f
C14242 DVDD.t136 VSS 0.167631f
C14243 DVDD.t78 VSS 0.167631f
C14244 DVDD.n9801 VSS 0.335261f
C14245 DVDD.n9802 VSS 0.081946f
C14246 DVDD.n9803 VSS 0.099098f
C14247 DVDD.n9804 VSS 0.198298f
C14248 DVDD.n9805 VSS 0.1401f
C14249 DVDD.n9806 VSS 0.163891f
C14250 DVDD.n9807 VSS 0.074015f
C14251 DVDD.n9809 VSS 0.163891f
C14252 DVDD.n9811 VSS 0.163891f
C14253 DVDD.n9812 VSS 0.134814f
C14254 DVDD.n9814 VSS 0.055963f
C14255 DVDD.n9817 VSS 0.128173f
C14256 DVDD.n9818 VSS 0.128173f
C14257 DVDD.n9819 VSS 0.128173f
C14258 DVDD.n9820 VSS 0.055963f
C14259 DVDD.n9821 VSS 0.128173f
C14260 DVDD.n9822 VSS 0.128173f
C14261 DVDD.n9823 VSS 0.055963f
C14262 DVDD.n9824 VSS 0.128173f
C14263 DVDD.n9825 VSS 0.128173f
C14264 DVDD.n9826 VSS 0.128173f
C14265 DVDD.n9827 VSS 0.128173f
C14266 DVDD.n9828 VSS 0.128173f
C14267 DVDD.n9829 VSS 0.128173f
C14268 DVDD.n9830 VSS 0.128173f
C14269 DVDD.n9831 VSS 0.055963f
C14270 DVDD.n9832 VSS 0.128173f
C14271 DVDD.n9833 VSS 0.128173f
C14272 DVDD.n9834 VSS 0.055963f
C14273 DVDD.n9835 VSS 0.128173f
C14274 DVDD.n9836 VSS 0.128173f
C14275 DVDD.n9837 VSS 0.159414f
C14276 DVDD.n9838 VSS 0.055963f
C14277 DVDD.n9839 VSS 0.128173f
C14278 DVDD.n9840 VSS 0.587849f
C14279 DVDD.n9841 VSS 0.128173f
C14280 DVDD.n9842 VSS 0.055963f
C14281 DVDD.n9843 VSS 0.128173f
C14282 DVDD.n9844 VSS 0.055963f
C14283 DVDD.n9845 VSS 0.128173f
C14284 DVDD.n9846 VSS 0.055963f
C14285 DVDD.n9847 VSS 0.128173f
C14286 DVDD.n9848 VSS 0.128173f
C14287 DVDD.n9849 VSS 0.128173f
C14288 DVDD.n9850 VSS 0.128173f
C14289 DVDD.n9851 VSS 0.055963f
C14290 DVDD.n9852 VSS 0.128173f
C14291 DVDD.n9853 VSS 0.055963f
C14292 DVDD.n9854 VSS 0.128173f
C14293 DVDD.n9855 VSS 0.055963f
C14294 DVDD.n9856 VSS 0.128173f
C14295 DVDD.n9857 VSS 0.128173f
C14296 DVDD.n9858 VSS 0.128173f
C14297 DVDD.n9859 VSS 0.128173f
C14298 DVDD.n9860 VSS 0.055963f
C14299 DVDD.n9861 VSS 0.128173f
C14300 DVDD.n9862 VSS 0.055963f
C14301 DVDD.n9863 VSS 0.128173f
C14302 DVDD.n9864 VSS 0.101545f
C14303 DVDD.n9865 VSS 0.128173f
C14304 DVDD.n9866 VSS 0.128173f
C14305 DVDD.n9867 VSS 0.128173f
C14306 DVDD.n9868 VSS 0.128173f
C14307 DVDD.n9869 VSS 0.128173f
C14308 DVDD.n9870 VSS 0.128173f
C14309 DVDD.n9871 VSS 0.128173f
C14310 DVDD.n9872 VSS 0.128173f
C14311 DVDD.n9873 VSS 0.111926f
C14312 DVDD.n9874 VSS 0.128173f
C14313 DVDD.n9875 VSS 0.055963f
C14314 DVDD.n9876 VSS 0.128173f
C14315 DVDD.n9877 VSS 0.055963f
C14316 DVDD.n9878 VSS 0.128173f
C14317 DVDD.n9879 VSS 0.128173f
C14318 DVDD.n9880 VSS 0.128173f
C14319 DVDD.n9881 VSS 0.128173f
C14320 DVDD.n9882 VSS 0.055963f
C14321 DVDD.n9883 VSS 0.128173f
C14322 DVDD.n9884 VSS 0.055963f
C14323 DVDD.n9885 VSS 0.128173f
C14324 DVDD.n9886 VSS 0.055963f
C14325 DVDD.n9887 VSS 0.128173f
C14326 DVDD.n9888 VSS 0.128173f
C14327 DVDD.n9889 VSS 0.128173f
C14328 DVDD.n9890 VSS 0.128173f
C14329 DVDD.n9891 VSS 0.055963f
C14330 DVDD.n9892 VSS 0.128173f
C14331 DVDD.n9893 VSS 0.055963f
C14332 DVDD.n9894 VSS 0.128173f
C14333 DVDD.n9895 VSS 0.055963f
C14334 DVDD.n9896 VSS 0.128173f
C14335 DVDD.n9897 VSS 0.128173f
C14336 DVDD.n9898 VSS 0.128173f
C14337 DVDD.n9899 VSS 0.128173f
C14338 DVDD.n9900 VSS 0.128173f
C14339 DVDD.n9901 VSS 0.055963f
C14340 DVDD.n9902 VSS 0.128173f
C14341 DVDD.n9903 VSS 0.128173f
C14342 DVDD.n9904 VSS 0.128173f
C14343 DVDD.n9905 VSS 0.055963f
C14344 DVDD.n9906 VSS 0.128173f
C14345 DVDD.n9907 VSS 0.128173f
C14346 DVDD.n9908 VSS 0.128173f
C14347 DVDD.n9909 VSS 0.055963f
C14348 DVDD.n9910 VSS 0.128173f
C14349 DVDD.n9911 VSS 0.055963f
C14350 DVDD.n9912 VSS 0.128173f
C14351 DVDD.n9913 VSS 0.055963f
C14352 DVDD.n9914 VSS 0.128173f
C14353 DVDD.n9915 VSS 0.128173f
C14354 DVDD.n9916 VSS 0.128173f
C14355 DVDD.n9917 VSS 0.128173f
C14356 DVDD.n9918 VSS 0.055963f
C14357 DVDD.n9919 VSS 0.128173f
C14358 DVDD.n9920 VSS 0.055963f
C14359 DVDD.n9921 VSS 0.128173f
C14360 DVDD.n9922 VSS 0.055963f
C14361 DVDD.n9923 VSS 0.128173f
C14362 DVDD.n9924 VSS 0.128173f
C14363 DVDD.n9925 VSS 0.128173f
C14364 DVDD.n9926 VSS 0.128173f
C14365 DVDD.n9927 VSS 0.128173f
C14366 DVDD.n9928 VSS 0.092068f
C14367 DVDD.n9929 VSS 0.128173f
C14368 DVDD.n9930 VSS 0.128173f
C14369 DVDD.n9931 VSS 0.128173f
C14370 DVDD.n9932 VSS 0.128173f
C14371 DVDD.n9933 VSS 0.128173f
C14372 DVDD.n9934 VSS 0.128173f
C14373 DVDD.n9935 VSS 0.128173f
C14374 DVDD.n9936 VSS 0.128173f
C14375 DVDD.n9937 VSS 0.055963f
C14376 DVDD.n9939 VSS 0.064086f
C14377 DVDD.n9940 VSS 0.198722f
C14378 DVDD.n9941 VSS 0.081946f
C14379 DVDD.n9942 VSS 0.098809f
C14380 DVDD.t130 VSS 0.167631f
C14381 DVDD.t152 VSS 0.167631f
C14382 DVDD.n9943 VSS 0.335261f
C14383 DVDD.n9944 VSS 0.081946f
C14384 DVDD.n9945 VSS 0.099098f
C14385 DVDD.n9946 VSS 0.198298f
C14386 DVDD.n9947 VSS 0.111023f
C14387 DVDD.n9948 VSS 0.064086f
C14388 DVDD.n9949 VSS 0.100449f
C14389 DVDD.n9950 VSS 0.198298f
C14390 DVDD.n9951 VSS 0.099098f
C14391 DVDD.t146 VSS 0.167631f
C14392 DVDD.t92 VSS 0.167631f
C14393 DVDD.n9952 VSS 0.335261f
C14394 DVDD.n9953 VSS 0.098809f
C14395 DVDD.n9954 VSS 0.198722f
C14396 DVDD.n9956 VSS 0.059573f
C14397 DVDD.n9957 VSS 0.064086f
C14398 DVDD.n9958 VSS 0.064086f
C14399 DVDD.n9959 VSS 0.064086f
C14400 DVDD.n9961 VSS 0.058671f
C14401 DVDD.n9962 VSS 0.064086f
C14402 DVDD.n9963 VSS 0.064086f
C14403 DVDD.n9964 VSS 0.055963f
C14404 DVDD.n9965 VSS 0.128173f
C14405 DVDD.n9966 VSS 0.128173f
C14406 DVDD.n9967 VSS 0.128173f
C14407 DVDD.n9968 VSS 0.128173f
C14408 DVDD.n9969 VSS 0.055963f
C14409 DVDD.n9970 VSS 0.128173f
C14410 DVDD.n9971 VSS 0.128173f
C14411 DVDD.n9972 VSS 0.055963f
C14412 DVDD.n9973 VSS 0.128173f
C14413 DVDD.n9974 VSS 0.128173f
C14414 DVDD.n9975 VSS 0.128173f
C14415 DVDD.n9976 VSS 0.128173f
C14416 DVDD.n9977 VSS 0.128173f
C14417 DVDD.n9978 VSS 0.055963f
C14418 DVDD.n9979 VSS 0.128173f
C14419 DVDD.n9980 VSS 0.055963f
C14420 DVDD.n9981 VSS 0.128173f
C14421 DVDD.n9982 VSS 0.055963f
C14422 DVDD.n9983 VSS 0.128173f
C14423 DVDD.n9984 VSS 0.128173f
C14424 DVDD.n9985 VSS 0.128173f
C14425 DVDD.n9986 VSS 0.128173f
C14426 DVDD.n9987 VSS 0.055963f
C14427 DVDD.n9988 VSS 0.128173f
C14428 DVDD.n9989 VSS 0.055963f
C14429 DVDD.n9990 VSS 0.128173f
C14430 DVDD.n9991 VSS 0.055963f
C14431 DVDD.n9992 VSS 0.128173f
C14432 DVDD.n9993 VSS 0.128173f
C14433 DVDD.n9994 VSS 0.128173f
C14434 DVDD.n9995 VSS 0.128173f
C14435 DVDD.n9996 VSS 0.128173f
C14436 DVDD.n9997 VSS 0.055963f
C14437 DVDD.n10001 VSS 0.064086f
C14438 DVDD.n10002 VSS 0.055963f
C14439 DVDD.n10003 VSS 0.128173f
C14440 DVDD.n10004 VSS 0.055963f
C14441 DVDD.n10005 VSS 0.128173f
C14442 DVDD.n10006 VSS 0.128173f
C14443 DVDD.n10007 VSS 0.128173f
C14444 DVDD.n10008 VSS 0.128173f
C14445 DVDD.n10009 VSS 0.128173f
C14446 DVDD.n10010 VSS 0.128173f
C14447 DVDD.n10011 VSS 0.055963f
C14448 DVDD.n10012 VSS 0.128173f
C14449 DVDD.n10013 VSS 0.128173f
C14450 DVDD.n10014 VSS 0.055963f
C14451 DVDD.n10015 VSS 0.115536f
C14452 DVDD.n10016 VSS 0.055963f
C14453 DVDD.n10017 VSS 0.159414f
C14454 DVDD.n10018 VSS 0.35687f
C14455 DVDD.n10019 VSS 0.589426f
C14456 DVDD.n10020 VSS 0.055963f
C14457 DVDD.n10021 VSS 0.128173f
C14458 DVDD.n10022 VSS 0.026627f
C14459 DVDD.n10023 VSS 0.076723f
C14460 DVDD.n10024 VSS 0.065892f
C14461 DVDD.n10025 VSS 0.128173f
C14462 DVDD.n10026 VSS 0.128173f
C14463 DVDD.n10027 VSS 0.055963f
C14464 DVDD.n10028 VSS 0.128173f
C14465 DVDD.n10029 VSS 0.055963f
C14466 DVDD.n10030 VSS 0.128173f
C14467 DVDD.n10031 VSS 0.055963f
C14468 DVDD.n10032 VSS 0.128173f
C14469 DVDD.n10033 VSS 0.128173f
C14470 DVDD.n10034 VSS 0.128173f
C14471 DVDD.n10035 VSS 0.128173f
C14472 DVDD.n10036 VSS 0.055963f
C14473 DVDD.n10037 VSS 0.128173f
C14474 DVDD.n10038 VSS 0.055963f
C14475 DVDD.n10039 VSS 0.128173f
C14476 DVDD.n10040 VSS 0.055963f
C14477 DVDD.n10041 VSS 0.128173f
C14478 DVDD.n10042 VSS 0.128173f
C14479 DVDD.n10043 VSS 0.128173f
C14480 DVDD.n10044 VSS 0.128173f
C14481 DVDD.n10045 VSS 0.128173f
C14482 DVDD.n10046 VSS 0.128173f
C14483 DVDD.n10047 VSS 0.128173f
C14484 DVDD.n10048 VSS 0.128173f
C14485 DVDD.n10049 VSS 0.128173f
C14486 DVDD.n10050 VSS 0.128173f
C14487 DVDD.n10051 VSS 0.128173f
C14488 DVDD.n10052 VSS 0.128173f
C14489 DVDD.n10053 VSS 0.128173f
C14490 DVDD.n10054 VSS 0.11012f
C14491 DVDD.n10055 VSS 0.064086f
C14492 DVDD.n10056 VSS 0.100449f
C14493 DVDD.n10057 VSS 0.064086f
C14494 DVDD.n10058 VSS 0.075821f
C14495 DVDD.n10059 VSS 0.128173f
C14496 DVDD.n10060 VSS 0.128173f
C14497 DVDD.n10061 VSS 0.128173f
C14498 DVDD.n10062 VSS 0.128173f
C14499 DVDD.n10063 VSS 0.128173f
C14500 DVDD.n10064 VSS 0.128173f
C14501 DVDD.n10065 VSS 0.090263f
C14502 DVDD.n10066 VSS 0.064086f
C14503 DVDD.n10067 VSS 0.100449f
C14504 DVDD.n10068 VSS 0.064086f
C14505 DVDD.n10069 VSS 0.055963f
C14506 DVDD.n10070 VSS 0.128173f
C14507 DVDD.n10071 VSS 0.128173f
C14508 DVDD.n10072 VSS 0.128173f
C14509 DVDD.n10073 VSS 0.128173f
C14510 DVDD.n10074 VSS 0.128173f
C14511 DVDD.n10075 VSS 0.128173f
C14512 DVDD.n10076 VSS 0.128173f
C14513 DVDD.n10077 VSS 0.128173f
C14514 DVDD.n10078 VSS 0.128173f
C14515 DVDD.n10079 VSS 0.128173f
C14516 DVDD.n10080 VSS 0.128173f
C14517 DVDD.n10081 VSS 0.128173f
C14518 DVDD.n10082 VSS 0.128173f
C14519 DVDD.n10083 VSS 0.128173f
C14520 DVDD.n10084 VSS 0.055963f
C14521 DVDD.n10085 VSS 0.128173f
C14522 DVDD.n10086 VSS 0.128173f
C14523 DVDD.n10087 VSS 0.128173f
C14524 DVDD.n10088 VSS 0.128173f
C14525 DVDD.n10089 VSS 0.128173f
C14526 DVDD.n10090 VSS 0.055963f
C14527 DVDD.n10091 VSS 0.058671f
C14528 DVDD.n10092 VSS 0.100449f
C14529 DVDD.n10093 VSS 0.064086f
C14530 DVDD.n10094 VSS 0.322495f
C14531 DVDD.n10095 VSS 0.581549f
C14532 DVDD.n10096 VSS 0.099098f
C14533 DVDD.n10097 VSS 0.697901f
C14534 DVDD.n10098 VSS 0.761343f
C14535 DVDD.n10099 VSS 0.099098f
C14536 DVDD.t141 VSS 0.167631f
C14537 DVDD.t126 VSS 0.167631f
C14538 DVDD.n10100 VSS 0.335261f
C14539 DVDD.n10101 VSS 0.098809f
C14540 DVDD.n10102 VSS 0.644991f
C14541 DVDD.n10103 VSS 0.644991f
C14542 DVDD.n10104 VSS 0.098809f
C14543 DVDD.t148 VSS 0.167631f
C14544 DVDD.t111 VSS 0.167631f
C14545 DVDD.n10105 VSS 0.335261f
C14546 DVDD.n10106 VSS 0.099098f
C14547 DVDD.n10107 VSS 0.644991f
C14548 DVDD.n10108 VSS 0.644991f
C14549 DVDD.n10109 VSS 0.099098f
C14550 DVDD.n10110 VSS 0.761343f
C14551 DVDD.n10111 VSS 0.761343f
C14552 DVDD.n10112 VSS 0.099098f
C14553 DVDD.t86 VSS 0.167631f
C14554 DVDD.t127 VSS 0.167631f
C14555 DVDD.n10113 VSS 0.335261f
C14556 DVDD.n10114 VSS 0.098809f
C14557 DVDD.n10115 VSS 0.644991f
C14558 DVDD.n10116 VSS 0.97806f
C14559 DVDD.n10117 VSS 0.098809f
C14560 DVDD.t94 VSS 0.425324f
C14561 DVDD.n10118 VSS 0.099098f
C14562 DVDD.n10119 VSS 0.97806f
C14563 DVDD.n10120 VSS 0.97806f
C14564 DVDD.n10121 VSS 0.099098f
C14565 DVDD.n10122 VSS 1.09441f
C14566 DVDD.n10123 VSS 0.761343f
C14567 DVDD.n10124 VSS 0.099098f
C14568 DVDD.t137 VSS 0.167631f
C14569 DVDD.t106 VSS 0.167631f
C14570 DVDD.n10125 VSS 0.335261f
C14571 DVDD.n10126 VSS 0.098809f
C14572 DVDD.n10127 VSS 0.644991f
C14573 DVDD.n10128 VSS 0.644991f
C14574 DVDD.n10129 VSS 0.098809f
C14575 DVDD.t149 VSS 0.167631f
C14576 DVDD.t115 VSS 0.167631f
C14577 DVDD.n10130 VSS 0.335261f
C14578 DVDD.n10131 VSS 0.099098f
C14579 DVDD.n10132 VSS 0.644991f
C14580 DVDD.n10133 VSS 0.644991f
C14581 DVDD.n10134 VSS 0.099098f
C14582 DVDD.n10135 VSS 0.761343f
C14583 DVDD.n10136 VSS 0.761343f
C14584 DVDD.n10137 VSS 0.099098f
C14585 DVDD.t87 VSS 0.167631f
C14586 DVDD.t128 VSS 0.167631f
C14587 DVDD.n10138 VSS 0.335261f
C14588 DVDD.n10139 VSS 0.098809f
C14589 DVDD.n10140 VSS 0.644991f
C14590 DVDD.n10141 VSS 0.644991f
C14591 DVDD.n10142 VSS 0.098809f
C14592 DVDD.t96 VSS 0.167631f
C14593 DVDD.t135 VSS 0.167631f
C14594 DVDD.n10143 VSS 0.335261f
C14595 DVDD.n10144 VSS 0.099098f
C14596 DVDD.n10145 VSS 0.644991f
C14597 DVDD.n10146 VSS 0.644991f
C14598 DVDD.n10147 VSS 0.099098f
C14599 DVDD.n10148 VSS 0.761343f
C14600 DVDD.n10149 VSS 0.761343f
C14601 DVDD.n10150 VSS 0.099098f
C14602 DVDD.t89 VSS 0.167631f
C14603 DVDD.t151 VSS 0.167631f
C14604 DVDD.n10151 VSS 0.335261f
C14605 DVDD.n10152 VSS 0.098809f
C14606 DVDD.n10153 VSS 0.644991f
C14607 DVDD.n10154 VSS 0.761754f
C14608 DVDD.n10155 VSS 0.098828f
C14609 DVDD.n10156 VSS 0.644991f
C14610 DVDD.n10157 VSS 0.644991f
C14611 DVDD.n10158 VSS 0.098809f
C14612 DVDD.t113 VSS 0.167631f
C14613 DVDD.t138 VSS 0.167631f
C14614 DVDD.n10159 VSS 0.335261f
C14615 DVDD.n10160 VSS 0.099098f
C14616 DVDD.n10161 VSS 0.644991f
C14617 DVDD.n10162 VSS 0.644991f
C14618 DVDD.n10163 VSS 0.099098f
C14619 DVDD.n10164 VSS 0.761343f
C14620 DVDD.n10165 VSS 0.098815f
C14621 DVDD.t132 VSS 0.425324f
C14622 DVDD.n10166 VSS 0.099098f
C14623 DVDD.n10167 VSS 1.16182f
C14624 DVDD.n10169 VSS 0.025624f
C14625 DVDD.n10170 VSS 0.025624f
C14626 DVDD.n10171 VSS 0.025624f
C14627 DVDD.n10172 VSS 0.025624f
C14628 DVDD.n10173 VSS 0.025624f
C14629 DVDD.n10174 VSS 0.025624f
C14630 DVDD.n10175 VSS 0.025624f
C14631 DVDD.n10177 VSS 0.098464f
C14632 DVDD.n10180 VSS 0.025624f
C14633 DVDD.n10183 VSS 0.025624f
C14634 DVDD.n10186 VSS 0.025624f
C14635 DVDD.n10189 VSS 0.025624f
C14636 DVDD.n10192 VSS 0.025624f
C14637 DVDD.n10195 VSS 0.025624f
C14638 DVDD.n10197 VSS 0.025624f
C14639 DVDD.n10199 VSS 0.025624f
C14640 DVDD.n10200 VSS 0.025624f
C14641 DVDD.n10202 VSS 0.794343f
C14642 DVDD.n10203 VSS 0.063349f
C14643 DVDD.n10204 VSS 0.063349f
C14644 DVDD.n10206 VSS 0.025624f
C14645 DVDD.n10208 VSS 0.025624f
C14646 DVDD.n10210 VSS 0.025624f
C14647 DVDD.n10212 VSS 0.025624f
C14648 DVDD.n10214 VSS 0.025624f
C14649 DVDD.n10216 VSS 0.025624f
C14650 DVDD.n10218 VSS 0.025624f
C14651 DVDD.n10219 VSS 0.794343f
C14652 DVDD.n10221 VSS 0.025624f
C14653 DVDD.n10222 VSS 0.468543f
C14654 DVDD.n10223 VSS 0.423753f
C14655 DVDD.n10224 VSS 0.05956f
C14656 DVDD.n10225 VSS 0.05956f
C14657 DVDD.n10226 VSS 0.043946f
C14658 DVDD.n10227 VSS 0.043732f
C14659 DVDD.n10228 VSS 0.048993f
C14660 DVDD.n10229 VSS 0.048993f
C14661 DVDD.n10230 VSS 0.56437f
C14662 DVDD.n10231 VSS 0.551735f
C14663 DVDD.n10232 VSS 0.522252f
C14664 DVDD.n10233 VSS 0.496982f
C14665 DVDD.n10234 VSS 0.047072f
C14666 DVDD.n10235 VSS 0.047072f
C14667 DVDD.n10236 VSS 0.024653f
C14668 DVDD.n10237 VSS 0.039516f
C14669 DVDD.n10238 VSS 0.039516f
C14670 DVDD.n10239 VSS 0.033945f
C14671 DVDD.n10240 VSS 0.033945f
C14672 DVDD.n10241 VSS 0.522252f
C14673 DVDD.n10283 VSS 0.425383f
C14674 DVDD.n10284 VSS 0.031128f
C14675 DVDD.n10285 VSS 0.019729f
C14676 DVDD.n10286 VSS 0.362207f
C14677 DVDD.n10328 VSS 0.349572f
C14678 DVDD.n10329 VSS 0.02513f
C14679 DVDD.n10330 VSS 0.031128f
C14680 DVDD.n10331 VSS 0.031128f
C14681 DVDD.n10332 VSS 0.031128f
C14682 DVDD.n10333 VSS 0.031128f
C14683 DVDD.n10334 VSS 0.031128f
C14684 DVDD.n10335 VSS 0.031128f
C14685 DVDD.n10336 VSS 0.031128f
C14686 DVDD.n10337 VSS 0.031128f
C14687 DVDD.n10338 VSS 0.031128f
C14688 DVDD.n10339 VSS 0.031128f
C14689 DVDD.n10340 VSS 0.031128f
C14690 DVDD.n10341 VSS 0.031128f
C14691 DVDD.n10342 VSS 0.031128f
C14692 DVDD.n10343 VSS 0.031128f
C14693 DVDD.n10344 VSS 0.031128f
C14694 DVDD.n10345 VSS 0.031128f
C14695 DVDD.n10346 VSS 0.031128f
C14696 DVDD.n10347 VSS 0.031128f
C14697 DVDD.n10348 VSS 0.031128f
C14698 DVDD.n10349 VSS 0.031128f
C14699 DVDD.n10350 VSS 0.031128f
C14700 DVDD.n10351 VSS 0.031128f
C14701 DVDD.n10352 VSS 0.031128f
C14702 DVDD.n10353 VSS 0.031128f
C14703 DVDD.n10354 VSS 0.031128f
C14704 DVDD.n10355 VSS 0.031128f
C14705 DVDD.n10356 VSS 0.031128f
C14706 DVDD.n10357 VSS 0.031128f
C14707 DVDD.n10358 VSS 0.031128f
C14708 DVDD.n10359 VSS 0.031128f
C14709 DVDD.n10360 VSS 0.031128f
C14710 DVDD.n10361 VSS 0.031128f
C14711 DVDD.n10362 VSS 0.031128f
C14712 DVDD.n10363 VSS 0.031128f
C14713 DVDD.n10364 VSS 0.031128f
C14714 DVDD.n10365 VSS 0.031128f
C14715 DVDD.n10366 VSS 0.031128f
C14716 DVDD.n10367 VSS 0.031128f
C14717 DVDD.n10368 VSS 0.031128f
C14718 DVDD.n10369 VSS 0.031128f
C14719 DVDD.n10370 VSS 0.031128f
C14720 DVDD.n10371 VSS 0.031128f
C14721 DVDD.n10372 VSS 0.031128f
C14722 DVDD.n10373 VSS 0.031128f
C14723 DVDD.n10374 VSS 0.031128f
C14724 DVDD.n10375 VSS 0.031128f
C14725 DVDD.n10376 VSS 0.031128f
C14726 DVDD.n10377 VSS 0.031128f
C14727 DVDD.n10378 VSS 0.031128f
C14728 DVDD.n10379 VSS 0.031128f
C14729 DVDD.n10380 VSS 0.031128f
C14730 DVDD.n10381 VSS 0.031128f
C14731 DVDD.n10382 VSS 0.031128f
C14732 DVDD.n10383 VSS 0.031128f
C14733 DVDD.n10384 VSS 0.031128f
C14734 DVDD.n10385 VSS 0.031128f
C14735 DVDD.n10386 VSS 0.031128f
C14736 DVDD.n10387 VSS 0.031128f
C14737 DVDD.n10388 VSS 0.031128f
C14738 DVDD.n10389 VSS 0.031128f
C14739 DVDD.n10390 VSS 0.031128f
C14740 DVDD.n10391 VSS 0.031128f
C14741 DVDD.n10392 VSS 0.028497f
C14742 DVDD.n10393 VSS 0.031128f
C14743 DVDD.n10394 VSS 0.031128f
C14744 DVDD.n10395 VSS 0.031128f
C14745 DVDD.n10396 VSS 0.031128f
C14746 DVDD.n10397 VSS 0.031128f
C14747 DVDD.n10398 VSS 0.031128f
C14748 DVDD.n10399 VSS 0.031128f
C14749 DVDD.n10400 VSS 0.031128f
C14750 DVDD.n10401 VSS 0.031128f
C14751 DVDD.n10402 VSS 0.031128f
C14752 DVDD.n10403 VSS 0.031128f
C14753 DVDD.n10404 VSS 0.031128f
C14754 DVDD.n10405 VSS 0.031128f
C14755 DVDD.n10406 VSS 0.031128f
C14756 DVDD.n10407 VSS 0.031128f
C14757 DVDD.n10408 VSS 0.031128f
C14758 DVDD.n10409 VSS 0.031128f
C14759 DVDD.n10410 VSS 0.031128f
C14760 DVDD.n10411 VSS 0.031128f
C14761 DVDD.n10412 VSS 0.031128f
C14762 DVDD.n10413 VSS 0.031128f
C14763 DVDD.n10414 VSS 0.031128f
C14764 DVDD.n10415 VSS 0.031128f
C14765 DVDD.n10416 VSS 0.031128f
C14766 DVDD.n10417 VSS 0.031128f
C14767 DVDD.n10418 VSS 0.031128f
C14768 DVDD.n10419 VSS 0.031128f
C14769 DVDD.n10420 VSS 0.031128f
C14770 DVDD.n10421 VSS 0.031128f
C14771 DVDD.n10422 VSS 0.031128f
C14772 DVDD.n10423 VSS 0.031128f
C14773 DVDD.n10424 VSS 0.031128f
C14774 DVDD.n10425 VSS 0.031128f
C14775 DVDD.n10426 VSS 0.031128f
C14776 DVDD.n10427 VSS 0.031128f
C14777 DVDD.n10428 VSS 0.031128f
C14778 DVDD.n10429 VSS 0.031128f
C14779 DVDD.n10430 VSS 0.031128f
C14780 DVDD.n10431 VSS 0.031128f
C14781 DVDD.n10432 VSS 0.031128f
C14782 DVDD.n10433 VSS 0.031128f
C14783 DVDD.n10434 VSS 0.031128f
C14784 DVDD.n10435 VSS 0.031128f
C14785 DVDD.n10436 VSS 0.031128f
C14786 DVDD.n10437 VSS 0.031128f
C14787 DVDD.n10438 VSS 0.031128f
C14788 DVDD.n10439 VSS 0.031128f
C14789 DVDD.n10440 VSS 0.031128f
C14790 DVDD.n10441 VSS 0.031128f
C14791 DVDD.n10442 VSS 0.031128f
C14792 DVDD.n10443 VSS 0.031128f
C14793 DVDD.n10444 VSS 0.031128f
C14794 DVDD.n10445 VSS 0.031128f
C14795 DVDD.n10446 VSS 0.031128f
C14796 DVDD.n10447 VSS 0.031128f
C14797 DVDD.n10448 VSS 0.031128f
C14798 DVDD.n10449 VSS 0.031128f
C14799 DVDD.n10450 VSS 0.031128f
C14800 DVDD.n10451 VSS 0.031128f
C14801 DVDD.n10452 VSS 0.031128f
C14802 DVDD.n10453 VSS 0.031128f
C14803 DVDD.n10454 VSS 0.031128f
C14804 DVDD.n10455 VSS 0.031128f
C14805 DVDD.n10456 VSS 0.031128f
C14806 DVDD.n10457 VSS 0.031128f
C14807 DVDD.n10458 VSS 0.031128f
C14808 DVDD.n10459 VSS 0.031128f
C14809 DVDD.n10460 VSS 0.031128f
C14810 DVDD.n10461 VSS 0.031128f
C14811 DVDD.n10462 VSS 0.031128f
C14812 DVDD.n10463 VSS 0.031128f
C14813 DVDD.n10464 VSS 0.031128f
C14814 DVDD.n10465 VSS 0.031128f
C14815 DVDD.n10466 VSS 0.031128f
C14816 DVDD.n10467 VSS 0.031128f
C14817 DVDD.n10468 VSS 0.031128f
C14818 DVDD.n10469 VSS 0.031128f
C14819 DVDD.n10470 VSS 0.031128f
C14820 DVDD.n10471 VSS 0.031128f
C14821 DVDD.n10472 VSS 0.031128f
C14822 DVDD.n10473 VSS 0.031128f
C14823 DVDD.n10474 VSS 0.031128f
C14824 DVDD.n10475 VSS 0.031128f
C14825 DVDD.n10476 VSS 0.031128f
C14826 DVDD.n10477 VSS 0.031128f
C14827 DVDD.n10478 VSS 0.031128f
C14828 DVDD.n10479 VSS 0.031128f
C14829 DVDD.n10480 VSS 0.031128f
C14830 DVDD.n10481 VSS 0.031128f
C14831 DVDD.n10482 VSS 0.031128f
C14832 DVDD.n10483 VSS 0.031128f
C14833 DVDD.n10484 VSS 0.031128f
C14834 DVDD.n10485 VSS 0.031128f
C14835 DVDD.n10486 VSS 0.031128f
C14836 DVDD.n10487 VSS 0.031128f
C14837 DVDD.n10488 VSS 0.031128f
C14838 DVDD.n10489 VSS 0.031128f
C14839 DVDD.n10490 VSS 0.031128f
C14840 DVDD.n10491 VSS 0.031128f
C14841 DVDD.n10492 VSS 0.031128f
C14842 DVDD.n10493 VSS 0.031128f
C14843 DVDD.n10494 VSS 0.031128f
C14844 DVDD.n10495 VSS 0.031128f
C14845 DVDD.n10496 VSS 0.031128f
C14846 DVDD.n10497 VSS 0.031128f
C14847 DVDD.n10498 VSS 0.031128f
C14848 DVDD.n10499 VSS 0.031128f
C14849 DVDD.n10500 VSS 0.031128f
C14850 DVDD.n10501 VSS 0.031128f
C14851 DVDD.n10502 VSS 0.031128f
C14852 DVDD.n10503 VSS 0.031128f
C14853 DVDD.n10504 VSS 0.031128f
C14854 DVDD.n10505 VSS 0.031128f
C14855 DVDD.n10506 VSS 0.031128f
C14856 DVDD.n10507 VSS 0.031128f
C14857 DVDD.n10508 VSS 0.031128f
C14858 DVDD.n10509 VSS 0.031128f
C14859 DVDD.n10510 VSS 0.031128f
C14860 DVDD.n10511 VSS 0.031128f
C14861 DVDD.n10512 VSS 0.031128f
C14862 DVDD.n10513 VSS 0.031128f
C14863 DVDD.n10514 VSS 0.031128f
C14864 DVDD.n10515 VSS 0.031128f
C14865 DVDD.n10516 VSS 0.031128f
C14866 DVDD.n10517 VSS 0.031128f
C14867 DVDD.n10518 VSS 0.031128f
C14868 DVDD.n10519 VSS 0.031128f
C14869 DVDD.n10520 VSS 0.031128f
C14870 DVDD.n10521 VSS 0.031128f
C14871 DVDD.n10522 VSS 0.031128f
C14872 DVDD.n10523 VSS 0.031128f
C14873 DVDD.n10524 VSS 0.031128f
C14874 DVDD.n10525 VSS 0.031128f
C14875 DVDD.n10526 VSS 0.031128f
C14876 DVDD.n10527 VSS 0.031128f
C14877 DVDD.n10528 VSS 0.031128f
C14878 DVDD.n10529 VSS 0.031128f
C14879 DVDD.n10530 VSS 0.031128f
C14880 DVDD.n10531 VSS 0.031128f
C14881 DVDD.n10532 VSS 0.031128f
C14882 DVDD.n10533 VSS 0.031128f
C14883 DVDD.n10534 VSS 0.031128f
C14884 DVDD.n10535 VSS 0.031128f
C14885 DVDD.n10536 VSS 0.031128f
C14886 DVDD.n10537 VSS 0.031128f
C14887 DVDD.n10538 VSS 0.031128f
C14888 DVDD.n10539 VSS 0.031128f
C14889 DVDD.n10540 VSS 0.031128f
C14890 DVDD.n10541 VSS 0.031128f
C14891 DVDD.n10542 VSS 0.031128f
C14892 DVDD.n10543 VSS 0.031128f
C14893 DVDD.n10544 VSS 0.031128f
C14894 DVDD.n10545 VSS 0.031128f
C14895 DVDD.n10546 VSS 0.031128f
C14896 DVDD.n10547 VSS 0.031128f
C14897 DVDD.n10548 VSS 0.031128f
C14898 DVDD.n10549 VSS 0.031128f
C14899 DVDD.n10550 VSS 0.031128f
C14900 DVDD.n10551 VSS 0.031128f
C14901 DVDD.n10552 VSS 0.031128f
C14902 DVDD.n10553 VSS 0.031128f
C14903 DVDD.n10554 VSS 0.031128f
C14904 DVDD.n10555 VSS 0.031128f
C14905 DVDD.n10556 VSS 0.031128f
C14906 DVDD.n10557 VSS 0.031128f
C14907 DVDD.n10558 VSS 0.031128f
C14908 DVDD.n10559 VSS 0.031128f
C14909 DVDD.n10560 VSS 0.031128f
C14910 DVDD.n10561 VSS 0.031128f
C14911 DVDD.n10562 VSS 0.031128f
C14912 DVDD.n10563 VSS 0.031128f
C14913 DVDD.n10564 VSS 0.031128f
C14914 DVDD.n10565 VSS 0.031128f
C14915 DVDD.n10566 VSS 0.031128f
C14916 DVDD.n10567 VSS 0.031128f
C14917 DVDD.n10568 VSS 0.031128f
C14918 DVDD.n10569 VSS 0.031128f
C14919 DVDD.n10570 VSS 0.031128f
C14920 DVDD.n10571 VSS 0.031128f
C14921 DVDD.n10572 VSS 0.031128f
C14922 DVDD.n10573 VSS 0.031128f
C14923 DVDD.n10574 VSS 0.031128f
C14924 DVDD.n10575 VSS 0.031128f
C14925 DVDD.n10576 VSS 0.026086f
C14926 DVDD.n10577 VSS 0.024066f
C14927 DVDD.n10578 VSS 0.041193f
C14928 DVDD.n10579 VSS 0.03883f
C14929 DVDD.n10580 VSS 0.03056f
C14930 DVDD.n10581 VSS 0.034992f
C14931 DVDD.n10582 VSS 0.598063f
C14932 DVDD.n10583 VSS 0.44223f
C14933 DVDD.n10584 VSS 0.034992f
C14934 DVDD.n10585 VSS 0.024066f
C14935 DVDD.n10586 VSS 0.041931f
C14936 DVDD.n10587 VSS 0.041931f
C14937 DVDD.n10588 VSS 0.036621f
C14938 DVDD.n10589 VSS 0.021018f
C14939 DVDD.n10590 VSS 0.028833f
C14940 DVDD.n10591 VSS 0.026086f
C14941 DVDD.n10592 VSS 0.036621f
C14942 DVDD.n10593 VSS 0.02513f
C14943 DVDD.n10594 VSS 0.041931f
C14944 DVDD.n10595 VSS 0.02513f
C14945 DVDD.n10596 VSS 0.041931f
C14946 DVDD.n10597 VSS 0.332725f
C14947 DVDD.n10639 VSS 0.019729f
C14948 DVDD.n10640 VSS 0.332725f
C14949 DVDD.n10641 VSS 0.019729f
C14950 DVDD.n10642 VSS 0.522253f
C14951 DVDD.n10643 VSS 0.031128f
C14952 DVDD.n10644 VSS 0.031128f
C14953 DVDD.n10645 VSS 0.031128f
C14954 DVDD.n10646 VSS 0.031128f
C14955 DVDD.n10647 VSS 0.031128f
C14956 DVDD.n10648 VSS 0.031128f
C14957 DVDD.n10649 VSS 0.031128f
C14958 DVDD.n10650 VSS 0.031128f
C14959 DVDD.n10651 VSS 0.031128f
C14960 DVDD.n10652 VSS 0.031128f
C14961 DVDD.n10653 VSS 0.031128f
C14962 DVDD.n10654 VSS 0.031128f
C14963 DVDD.n10655 VSS 0.031128f
C14964 DVDD.n10656 VSS 0.031128f
C14965 DVDD.n10657 VSS 0.031128f
C14966 DVDD.n10658 VSS 0.031128f
C14967 DVDD.n10659 VSS 0.031128f
C14968 DVDD.n10660 VSS 0.031128f
C14969 DVDD.n10661 VSS 0.031128f
C14970 DVDD.n10662 VSS 0.031128f
C14971 DVDD.n10663 VSS 0.031128f
C14972 DVDD.n10664 VSS 0.031128f
C14973 DVDD.n10665 VSS 0.031128f
C14974 DVDD.n10666 VSS 0.031128f
C14975 DVDD.n10667 VSS 0.031128f
C14976 DVDD.n10668 VSS 0.031128f
C14977 DVDD.n10669 VSS 0.031128f
C14978 DVDD.n10670 VSS 0.031128f
C14979 DVDD.n10671 VSS 0.031128f
C14980 DVDD.n10672 VSS 0.031128f
C14981 DVDD.n10673 VSS 0.031128f
C14982 DVDD.n10674 VSS 0.031128f
C14983 DVDD.n10675 VSS 0.031128f
C14984 DVDD.n10676 VSS 0.031128f
C14985 DVDD.n10677 VSS 0.031128f
C14986 DVDD.n10678 VSS 0.031128f
C14987 DVDD.n10679 VSS 0.031128f
C14988 DVDD.n10680 VSS 0.031128f
C14989 DVDD.n10681 VSS 0.031128f
C14990 DVDD.n10682 VSS 0.031128f
C14991 DVDD.n10684 VSS 0.031128f
C14992 DVDD.n10685 VSS 0.031128f
C14993 DVDD.n10686 VSS 0.039516f
C14994 DVDD.n10687 VSS 0.030741f
C14995 DVDD.n10688 VSS 0.05956f
C14996 DVDD.n10689 VSS 0.05956f
C14997 DVDD.n10690 VSS 0.598063f
C14998 DVDD.n10691 VSS 0.041193f
C14999 DVDD.n10692 VSS 0.522252f
C15000 DVDD.n10693 VSS 0.265338f
C15001 DVDD.n10694 VSS 0.05956f
C15002 DVDD.n10695 VSS 0.035544f
C15003 DVDD.n10696 VSS 0.035544f
C15004 DVDD.n10697 VSS 0.031727f
C15005 DVDD.n10698 VSS 0.053165f
C15006 DVDD.n10699 VSS 0.02744f
C15007 DVDD.n10700 VSS 0.053165f
C15008 DVDD.n10701 VSS 0.05956f
C15009 DVDD.n10702 VSS 0.05956f
C15010 DVDD.n10703 VSS 0.030741f
C15011 DVDD.n10704 VSS 0.033945f
C15012 DVDD.n10705 VSS 0.0586f
C15013 DVDD.n10706 VSS 0.039516f
C15014 DVDD.n10707 VSS 0.033945f
C15015 DVDD.n10708 VSS 0.05956f
C15016 DVDD.n10709 VSS 0.033945f
C15017 DVDD.n10710 VSS 0.332725f
C15018 DVDD.n10711 VSS 0.256914f
C15019 DVDD.n10712 VSS 0.02513f
C15020 DVDD.n10713 VSS 0.041931f
C15021 DVDD.n10714 VSS 0.02513f
C15022 DVDD.n10715 VSS 0.041931f
C15023 DVDD.n10716 VSS 0.031128f
C15024 DVDD.n10717 VSS 0.031128f
C15025 DVDD.n10718 VSS 0.031128f
C15026 DVDD.n10720 VSS 0.031128f
C15027 DVDD.n10721 VSS 0.031128f
C15028 DVDD.n10722 VSS 0.031128f
C15029 DVDD.n10724 VSS 0.031128f
C15030 DVDD.n10725 VSS 0.031128f
C15031 DVDD.n10726 VSS 0.031128f
C15032 DVDD.n10728 VSS 0.031128f
C15033 DVDD.n10729 VSS 0.031128f
C15034 DVDD.n10730 VSS 0.031128f
C15035 DVDD.n10732 VSS 0.031128f
C15036 DVDD.n10733 VSS 0.031128f
C15037 DVDD.n10734 VSS 0.031128f
C15038 DVDD.n10736 VSS 0.031128f
C15039 DVDD.n10737 VSS 0.031128f
C15040 DVDD.n10738 VSS 0.031128f
C15041 DVDD.n10740 VSS 0.031128f
C15042 DVDD.n10741 VSS 0.031128f
C15043 DVDD.n10742 VSS 0.031128f
C15044 DVDD.n10744 VSS 0.031128f
C15045 DVDD.n10745 VSS 0.031128f
C15046 DVDD.n10746 VSS 0.031128f
C15047 DVDD.n10748 VSS 0.031128f
C15048 DVDD.n10749 VSS 0.031128f
C15049 DVDD.n10750 VSS 0.031128f
C15050 DVDD.n10752 VSS 0.031128f
C15051 DVDD.n10753 VSS 0.031128f
C15052 DVDD.n10754 VSS 0.031128f
C15053 DVDD.n10756 VSS 0.031128f
C15054 DVDD.n10757 VSS 0.031128f
C15055 DVDD.n10758 VSS 0.031128f
C15056 DVDD.n10760 VSS 0.031128f
C15057 DVDD.n10761 VSS 0.031128f
C15058 DVDD.n10762 VSS 0.031128f
C15059 DVDD.n10764 VSS 0.031128f
C15060 DVDD.n10765 VSS 0.031128f
C15061 DVDD.n10766 VSS 0.031128f
C15062 DVDD.n10768 VSS 0.031128f
C15063 DVDD.n10769 VSS 0.031128f
C15064 DVDD.n10770 VSS 0.031128f
C15065 DVDD.n10772 VSS 0.031128f
C15066 DVDD.n10773 VSS 0.031128f
C15067 DVDD.n10774 VSS 0.031128f
C15068 DVDD.n10776 VSS 0.031128f
C15069 DVDD.n10777 VSS 0.031128f
C15070 DVDD.n10778 VSS 0.031128f
C15071 DVDD.n10780 VSS 0.031128f
C15072 DVDD.n10781 VSS 0.031128f
C15073 DVDD.n10782 VSS 0.031128f
C15074 DVDD.n10784 VSS 0.031128f
C15075 DVDD.n10785 VSS 0.031128f
C15076 DVDD.n10786 VSS 0.031128f
C15077 DVDD.n10788 VSS 0.031128f
C15078 DVDD.n10789 VSS 0.031128f
C15079 DVDD.n10790 VSS 0.031128f
C15080 DVDD.n10792 VSS 0.031128f
C15081 DVDD.n10793 VSS 0.031128f
C15082 DVDD.n10794 VSS 0.031128f
C15083 DVDD.n10796 VSS 0.031128f
C15084 DVDD.n10797 VSS 0.031128f
C15085 DVDD.n10798 VSS 0.031128f
C15086 DVDD.n10799 VSS 0.028497f
C15087 DVDD.n10800 VSS 0.019729f
C15088 DVDD.n10801 VSS 0.019729f
C15089 DVDD.n10803 VSS 0.031128f
C15090 DVDD.n10805 VSS 0.031128f
C15091 DVDD.n10807 VSS 0.031128f
C15092 DVDD.n10808 VSS 0.031128f
C15093 DVDD.n10809 VSS 0.031128f
C15094 DVDD.n10810 VSS 0.031128f
C15095 DVDD.n10811 VSS 0.031128f
C15096 DVDD.n10812 VSS 0.031128f
C15097 DVDD.n10813 VSS 0.031128f
C15098 DVDD.n10815 VSS 0.031128f
C15099 DVDD.n10817 VSS 0.031128f
C15100 DVDD.n10819 VSS 0.031128f
C15101 DVDD.n10820 VSS 0.031128f
C15102 DVDD.n10821 VSS 0.031128f
C15103 DVDD.n10822 VSS 0.031128f
C15104 DVDD.n10823 VSS 0.031128f
C15105 DVDD.n10824 VSS 0.031128f
C15106 DVDD.n10825 VSS 0.031128f
C15107 DVDD.n10827 VSS 0.031128f
C15108 DVDD.n10829 VSS 0.031128f
C15109 DVDD.n10831 VSS 0.031128f
C15110 DVDD.n10832 VSS 0.031128f
C15111 DVDD.n10833 VSS 0.031128f
C15112 DVDD.n10834 VSS 0.031128f
C15113 DVDD.n10835 VSS 0.031128f
C15114 DVDD.n10836 VSS 0.031128f
C15115 DVDD.n10837 VSS 0.031128f
C15116 DVDD.n10839 VSS 0.031128f
C15117 DVDD.n10841 VSS 0.031128f
C15118 DVDD.n10843 VSS 0.031128f
C15119 DVDD.n10844 VSS 0.031128f
C15120 DVDD.n10845 VSS 0.031128f
C15121 DVDD.n10846 VSS 0.031128f
C15122 DVDD.n10847 VSS 0.031128f
C15123 DVDD.n10848 VSS 0.031128f
C15124 DVDD.n10849 VSS 0.031128f
C15125 DVDD.n10851 VSS 0.031128f
C15126 DVDD.n10853 VSS 0.031128f
C15127 DVDD.n10855 VSS 0.031128f
C15128 DVDD.n10856 VSS 0.031128f
C15129 DVDD.n10857 VSS 0.031128f
C15130 DVDD.n10858 VSS 0.031128f
C15131 DVDD.n10859 VSS 0.031128f
C15132 DVDD.n10860 VSS 0.031128f
C15133 DVDD.n10861 VSS 0.031128f
C15134 DVDD.n10863 VSS 0.031128f
C15135 DVDD.n10865 VSS 0.031128f
C15136 DVDD.n10867 VSS 0.031128f
C15137 DVDD.n10868 VSS 0.031128f
C15138 DVDD.n10869 VSS 0.031128f
C15139 DVDD.n10870 VSS 0.031128f
C15140 DVDD.n10871 VSS 0.031128f
C15141 DVDD.n10872 VSS 0.031128f
C15142 DVDD.n10873 VSS 0.031128f
C15143 DVDD.n10875 VSS 0.031128f
C15144 DVDD.n10877 VSS 0.031128f
C15145 DVDD.n10879 VSS 0.031128f
C15146 DVDD.n10880 VSS 0.031128f
C15147 DVDD.n10881 VSS 0.031128f
C15148 DVDD.n10882 VSS 0.031128f
C15149 DVDD.n10883 VSS 0.031128f
C15150 DVDD.n10884 VSS 0.031128f
C15151 DVDD.n10885 VSS 0.031128f
C15152 DVDD.n10887 VSS 0.031128f
C15153 DVDD.n10889 VSS 0.031128f
C15154 DVDD.n10891 VSS 0.031128f
C15155 DVDD.n10892 VSS 0.031128f
C15156 DVDD.n10893 VSS 0.031128f
C15157 DVDD.n10894 VSS 0.031128f
C15158 DVDD.n10895 VSS 0.031128f
C15159 DVDD.n10896 VSS 0.031128f
C15160 DVDD.n10897 VSS 0.031128f
C15161 DVDD.n10899 VSS 0.031128f
C15162 DVDD.n10901 VSS 0.031128f
C15163 DVDD.n10903 VSS 0.031128f
C15164 DVDD.n10904 VSS 0.031128f
C15165 DVDD.n10905 VSS 0.031128f
C15166 DVDD.n10906 VSS 0.031128f
C15167 DVDD.n10907 VSS 0.031128f
C15168 DVDD.n10908 VSS 0.031128f
C15169 DVDD.n10909 VSS 0.031128f
C15170 DVDD.n10911 VSS 0.031128f
C15171 DVDD.n10913 VSS 0.031128f
C15172 DVDD.n10915 VSS 0.031128f
C15173 DVDD.n10916 VSS 0.031128f
C15174 DVDD.n10917 VSS 0.031128f
C15175 DVDD.n10918 VSS 0.031128f
C15176 DVDD.n10919 VSS 0.031128f
C15177 DVDD.n10920 VSS 0.031128f
C15178 DVDD.n10921 VSS 0.031128f
C15179 DVDD.n10923 VSS 0.031128f
C15180 DVDD.n10925 VSS 0.031128f
C15181 DVDD.n10927 VSS 0.031128f
C15182 DVDD.n10928 VSS 0.031128f
C15183 DVDD.n10929 VSS 0.031128f
C15184 DVDD.n10930 VSS 0.031128f
C15185 DVDD.n10931 VSS 0.031128f
C15186 DVDD.n10932 VSS 0.031128f
C15187 DVDD.n10933 VSS 0.031128f
C15188 DVDD.n10935 VSS 0.031128f
C15189 DVDD.n10937 VSS 0.031128f
C15190 DVDD.n10939 VSS 0.031128f
C15191 DVDD.n10940 VSS 0.031128f
C15192 DVDD.n10941 VSS 0.031128f
C15193 DVDD.n10942 VSS 0.031128f
C15194 DVDD.n10943 VSS 0.031128f
C15195 DVDD.n10944 VSS 0.031128f
C15196 DVDD.n10945 VSS 0.031128f
C15197 DVDD.n10947 VSS 0.031128f
C15198 DVDD.n10949 VSS 0.031128f
C15199 DVDD.n10951 VSS 0.031128f
C15200 DVDD.n10952 VSS 0.031128f
C15201 DVDD.n10953 VSS 0.031128f
C15202 DVDD.n10954 VSS 0.031128f
C15203 DVDD.n10955 VSS 0.031128f
C15204 DVDD.n10956 VSS 0.031128f
C15205 DVDD.n10957 VSS 0.031128f
C15206 DVDD.n10959 VSS 0.031128f
C15207 DVDD.n10961 VSS 0.031128f
C15208 DVDD.n10963 VSS 0.031128f
C15209 DVDD.n10964 VSS 0.031128f
C15210 DVDD.n10965 VSS 0.031128f
C15211 DVDD.n10966 VSS 0.031128f
C15212 DVDD.n10967 VSS 0.031128f
C15213 DVDD.n10968 VSS 0.031128f
C15214 DVDD.n10969 VSS 0.031128f
C15215 DVDD.n10971 VSS 0.031128f
C15216 DVDD.n10973 VSS 0.031128f
C15217 DVDD.n10975 VSS 0.031128f
C15218 DVDD.n10976 VSS 0.031128f
C15219 DVDD.n10977 VSS 0.031128f
C15220 DVDD.n10978 VSS 0.031128f
C15221 DVDD.n10979 VSS 0.031128f
C15222 DVDD.n10980 VSS 0.031128f
C15223 DVDD.n10981 VSS 0.031128f
C15224 DVDD.n10983 VSS 0.031128f
C15225 DVDD.n10985 VSS 0.031128f
C15226 DVDD.n10987 VSS 0.031128f
C15227 DVDD.n10988 VSS 0.031128f
C15228 DVDD.n10989 VSS 0.031128f
C15229 DVDD.n10990 VSS 0.031128f
C15230 DVDD.n10991 VSS 0.031128f
C15231 DVDD.n10992 VSS 0.031128f
C15232 DVDD.n10993 VSS 0.031128f
C15233 DVDD.n10995 VSS 0.031128f
C15234 DVDD.n10997 VSS 0.031128f
C15235 DVDD.n10999 VSS 0.031128f
C15236 DVDD.n11000 VSS 0.031128f
C15237 DVDD.n11001 VSS 0.031128f
C15238 DVDD.n11002 VSS 0.031128f
C15239 DVDD.n11003 VSS 0.031128f
C15240 DVDD.n11004 VSS 0.031128f
C15241 DVDD.n11005 VSS 0.031128f
C15242 DVDD.n11007 VSS 0.031128f
C15243 DVDD.n11009 VSS 0.031128f
C15244 DVDD.n11011 VSS 0.031128f
C15245 DVDD.n11012 VSS 0.031128f
C15246 DVDD.n11013 VSS 0.031128f
C15247 DVDD.n11014 VSS 0.031128f
C15248 DVDD.n11015 VSS 0.031128f
C15249 DVDD.n11016 VSS 0.031128f
C15250 DVDD.n11017 VSS 0.031128f
C15251 DVDD.n11019 VSS 0.031128f
C15252 DVDD.n11021 VSS 0.031128f
C15253 DVDD.n11023 VSS 0.031128f
C15254 DVDD.n11024 VSS 0.031128f
C15255 DVDD.n11025 VSS 0.031128f
C15256 DVDD.n11026 VSS 0.031128f
C15257 DVDD.n11027 VSS 0.031128f
C15258 DVDD.n11028 VSS 0.031128f
C15259 DVDD.n11029 VSS 0.031128f
C15260 DVDD.n11031 VSS 0.031128f
C15261 DVDD.n11033 VSS 0.031128f
C15262 DVDD.n11035 VSS 0.031128f
C15263 DVDD.n11036 VSS 0.031128f
C15264 DVDD.n11037 VSS 0.031128f
C15265 DVDD.n11038 VSS 0.031128f
C15266 DVDD.n11039 VSS 0.031128f
C15267 DVDD.n11040 VSS 0.031128f
C15268 DVDD.n11041 VSS 0.031128f
C15269 DVDD.n11042 VSS 0.031128f
C15270 DVDD.n11044 VSS 0.031128f
C15271 DVDD.n11046 VSS 0.031128f
C15272 DVDD.n11048 VSS 0.019729f
C15273 DVDD.n11049 VSS 0.019729f
C15274 DVDD.n11050 VSS 0.026086f
C15275 DVDD.n11051 VSS 0.160045f
C15276 DVDD.n11052 VSS 0.551735f
C15277 DVDD.n11053 VSS 0.353784f
C15278 DVDD.n11054 VSS 0.037354f
C15279 DVDD.n11055 VSS 0.037354f
C15280 DVDD.n11056 VSS 0.032623f
C15281 DVDD.n11057 VSS 0.028833f
C15282 DVDD.n11058 VSS 0.028833f
C15283 DVDD.n11059 VSS 0.02513f
C15284 DVDD.n11060 VSS 0.02513f
C15285 DVDD.n11061 VSS 0.598063f
C15286 DVDD.n11103 VSS 0.530676f
C15287 DVDD.n11104 VSS 0.031128f
C15288 DVDD.n11105 VSS 0.033945f
C15289 DVDD.n11106 VSS 0.019729f
C15290 DVDD.n11107 VSS 0.067387f
C15291 DVDD.n11149 VSS 0.530676f
C15292 DVDD.n11150 VSS 0.031128f
C15293 DVDD.n11151 VSS 0.031128f
C15294 DVDD.n11152 VSS 0.031128f
C15295 DVDD.n11153 VSS 0.031128f
C15296 DVDD.n11154 VSS 0.031128f
C15297 DVDD.n11155 VSS 0.031128f
C15298 DVDD.n11156 VSS 0.031128f
C15299 DVDD.n11157 VSS 0.031128f
C15300 DVDD.n11158 VSS 0.031128f
C15301 DVDD.n11159 VSS 0.031128f
C15302 DVDD.n11160 VSS 0.031128f
C15303 DVDD.n11161 VSS 0.031128f
C15304 DVDD.n11162 VSS 0.031128f
C15305 DVDD.n11163 VSS 0.031128f
C15306 DVDD.n11164 VSS 0.031128f
C15307 DVDD.n11165 VSS 0.031128f
C15308 DVDD.n11166 VSS 0.031128f
C15309 DVDD.n11167 VSS 0.031128f
C15310 DVDD.n11168 VSS 0.031128f
C15311 DVDD.n11169 VSS 0.031128f
C15312 DVDD.n11170 VSS 0.031128f
C15313 DVDD.n11171 VSS 0.031128f
C15314 DVDD.n11172 VSS 0.031128f
C15315 DVDD.n11173 VSS 0.031128f
C15316 DVDD.n11174 VSS 0.031128f
C15317 DVDD.n11175 VSS 0.031128f
C15318 DVDD.n11176 VSS 0.031128f
C15319 DVDD.n11177 VSS 0.031128f
C15320 DVDD.n11178 VSS 0.031128f
C15321 DVDD.n11179 VSS 0.031128f
C15322 DVDD.n11180 VSS 0.031128f
C15323 DVDD.n11181 VSS 0.031128f
C15324 DVDD.n11182 VSS 0.031128f
C15325 DVDD.n11183 VSS 0.031128f
C15326 DVDD.n11184 VSS 0.031128f
C15327 DVDD.n11185 VSS 0.031128f
C15328 DVDD.n11186 VSS 0.031128f
C15329 DVDD.n11187 VSS 0.031128f
C15330 DVDD.n11188 VSS 0.031128f
C15331 DVDD.n11189 VSS 0.031128f
C15332 DVDD.n11190 VSS 0.031128f
C15333 DVDD.n11191 VSS 0.031128f
C15334 DVDD.n11192 VSS 0.031128f
C15335 DVDD.n11193 VSS 0.031128f
C15336 DVDD.n11194 VSS 0.031128f
C15337 DVDD.n11195 VSS 0.031128f
C15338 DVDD.n11196 VSS 0.031128f
C15339 DVDD.n11197 VSS 0.031128f
C15340 DVDD.n11198 VSS 0.031128f
C15341 DVDD.n11199 VSS 0.031128f
C15342 DVDD.n11200 VSS 0.031128f
C15343 DVDD.n11201 VSS 0.031128f
C15344 DVDD.n11202 VSS 0.031128f
C15345 DVDD.n11203 VSS 0.031128f
C15346 DVDD.n11204 VSS 0.031128f
C15347 DVDD.n11205 VSS 0.031128f
C15348 DVDD.n11206 VSS 0.031128f
C15349 DVDD.n11207 VSS 0.031128f
C15350 DVDD.n11208 VSS 0.031128f
C15351 DVDD.n11209 VSS 0.031128f
C15352 DVDD.n11210 VSS 0.031128f
C15353 DVDD.n11211 VSS 0.031128f
C15354 DVDD.n11212 VSS 0.039445f
C15355 DVDD.n11213 VSS 0.053165f
C15356 DVDD.n11214 VSS 0.05956f
C15357 DVDD.n11215 VSS 0.522252f
C15358 DVDD.n11216 VSS 0.433807f
C15359 DVDD.n11217 VSS 0.053165f
C15360 DVDD.n11218 VSS 0.046305f
C15361 DVDD.n11219 VSS 0.051875f
C15362 DVDD.n11220 VSS 0.051875f
C15363 DVDD.n11221 VSS 0.05956f
C15364 DVDD.n11222 VSS 0.04419f
C15365 DVDD.n11223 VSS 0.04419f
C15366 DVDD.n11224 VSS 0.033945f
C15367 DVDD.n11225 VSS 0.05956f
C15368 DVDD.n11226 VSS 0.033945f
C15369 DVDD.n11227 VSS 0.543311f
C15370 DVDD.n11228 VSS 0.033945f
C15371 DVDD.n11229 VSS 0.028497f
C15372 DVDD.n11230 VSS 0.053165f
C15373 DVDD.n11231 VSS 0.05956f
C15374 DVDD.n11232 VSS 0.05956f
C15375 DVDD.n11233 VSS 0.454865f
C15376 DVDD.n11275 VSS 0.019729f
C15377 DVDD.n11276 VSS 0.379054f
C15378 DVDD.n11277 VSS 0.02513f
C15379 DVDD.n11278 VSS 0.019729f
C15380 DVDD.n11279 VSS 0.122139f
C15381 DVDD.n11280 VSS 0.031128f
C15382 DVDD.n11281 VSS 0.031128f
C15383 DVDD.n11282 VSS 0.031128f
C15384 DVDD.n11283 VSS 0.031128f
C15385 DVDD.n11284 VSS 0.031128f
C15386 DVDD.n11285 VSS 0.031128f
C15387 DVDD.n11286 VSS 0.031128f
C15388 DVDD.n11287 VSS 0.031128f
C15389 DVDD.n11288 VSS 0.031128f
C15390 DVDD.n11289 VSS 0.031128f
C15391 DVDD.n11290 VSS 0.031128f
C15392 DVDD.n11291 VSS 0.031128f
C15393 DVDD.n11292 VSS 0.031128f
C15394 DVDD.n11293 VSS 0.031128f
C15395 DVDD.n11294 VSS 0.031128f
C15396 DVDD.n11295 VSS 0.031128f
C15397 DVDD.n11296 VSS 0.031128f
C15398 DVDD.n11297 VSS 0.031128f
C15399 DVDD.n11298 VSS 0.031128f
C15400 DVDD.n11299 VSS 0.031128f
C15401 DVDD.n11300 VSS 0.031128f
C15402 DVDD.n11301 VSS 0.031128f
C15403 DVDD.n11302 VSS 0.031128f
C15404 DVDD.n11303 VSS 0.031128f
C15405 DVDD.n11304 VSS 0.031128f
C15406 DVDD.n11305 VSS 0.031128f
C15407 DVDD.n11306 VSS 0.031128f
C15408 DVDD.n11307 VSS 0.031128f
C15409 DVDD.n11308 VSS 0.031128f
C15410 DVDD.n11309 VSS 0.031128f
C15411 DVDD.n11310 VSS 0.031128f
C15412 DVDD.n11311 VSS 0.031128f
C15413 DVDD.n11312 VSS 0.031128f
C15414 DVDD.n11313 VSS 0.031128f
C15415 DVDD.n11314 VSS 0.031128f
C15416 DVDD.n11315 VSS 0.031128f
C15417 DVDD.n11316 VSS 0.031128f
C15418 DVDD.n11317 VSS 0.031128f
C15419 DVDD.n11318 VSS 0.031128f
C15420 DVDD.n11319 VSS 0.031128f
C15421 DVDD.n11320 VSS 0.019729f
C15422 DVDD.n11322 VSS 0.031128f
C15423 DVDD.n11323 VSS 0.031128f
C15424 DVDD.n11324 VSS 0.031128f
C15425 DVDD.n11325 VSS 0.031128f
C15426 DVDD.n11326 VSS 0.031128f
C15427 DVDD.n11327 VSS 0.031128f
C15428 DVDD.n11329 VSS 0.031128f
C15429 DVDD.n11330 VSS 0.031128f
C15430 DVDD.n11331 VSS 0.031128f
C15431 DVDD.n11333 VSS 0.031128f
C15432 DVDD.n11334 VSS 0.031128f
C15433 DVDD.n11335 VSS 0.031128f
C15434 DVDD.n11336 VSS 0.031128f
C15435 DVDD.n11337 VSS 0.031128f
C15436 DVDD.n11338 VSS 0.031128f
C15437 DVDD.n11339 VSS 0.031128f
C15438 DVDD.n11341 VSS 0.031128f
C15439 DVDD.n11342 VSS 0.031128f
C15440 DVDD.n11343 VSS 0.031128f
C15441 DVDD.n11345 VSS 0.031128f
C15442 DVDD.n11346 VSS 0.031128f
C15443 DVDD.n11347 VSS 0.031128f
C15444 DVDD.n11348 VSS 0.031128f
C15445 DVDD.n11349 VSS 0.031128f
C15446 DVDD.n11350 VSS 0.031128f
C15447 DVDD.n11351 VSS 0.031128f
C15448 DVDD.n11353 VSS 0.031128f
C15449 DVDD.n11354 VSS 0.031128f
C15450 DVDD.n11355 VSS 0.031128f
C15451 DVDD.n11357 VSS 0.031128f
C15452 DVDD.n11358 VSS 0.031128f
C15453 DVDD.n11359 VSS 0.031128f
C15454 DVDD.n11360 VSS 0.031128f
C15455 DVDD.n11361 VSS 0.031128f
C15456 DVDD.n11362 VSS 0.031128f
C15457 DVDD.n11363 VSS 0.031128f
C15458 DVDD.n11365 VSS 0.031128f
C15459 DVDD.n11366 VSS 0.031128f
C15460 DVDD.n11367 VSS 0.031128f
C15461 DVDD.n11369 VSS 0.031128f
C15462 DVDD.n11370 VSS 0.031128f
C15463 DVDD.n11371 VSS 0.031128f
C15464 DVDD.n11372 VSS 0.031128f
C15465 DVDD.n11373 VSS 0.031128f
C15466 DVDD.n11374 VSS 0.031128f
C15467 DVDD.n11375 VSS 0.031128f
C15468 DVDD.n11377 VSS 0.031128f
C15469 DVDD.n11378 VSS 0.031128f
C15470 DVDD.n11379 VSS 0.031128f
C15471 DVDD.n11381 VSS 0.031128f
C15472 DVDD.n11382 VSS 0.031128f
C15473 DVDD.n11383 VSS 0.031128f
C15474 DVDD.n11384 VSS 0.031128f
C15475 DVDD.n11385 VSS 0.031128f
C15476 DVDD.n11386 VSS 0.031128f
C15477 DVDD.n11387 VSS 0.031128f
C15478 DVDD.n11389 VSS 0.031128f
C15479 DVDD.n11390 VSS 0.031128f
C15480 DVDD.n11391 VSS 0.031128f
C15481 DVDD.n11393 VSS 0.031128f
C15482 DVDD.n11394 VSS 0.031128f
C15483 DVDD.n11395 VSS 0.031128f
C15484 DVDD.n11396 VSS 0.031128f
C15485 DVDD.n11397 VSS 0.031128f
C15486 DVDD.n11398 VSS 0.031128f
C15487 DVDD.n11399 VSS 0.031128f
C15488 DVDD.n11401 VSS 0.031128f
C15489 DVDD.n11402 VSS 0.031128f
C15490 DVDD.n11403 VSS 0.031128f
C15491 DVDD.n11405 VSS 0.031128f
C15492 DVDD.n11406 VSS 0.031128f
C15493 DVDD.n11407 VSS 0.031128f
C15494 DVDD.n11408 VSS 0.031128f
C15495 DVDD.n11409 VSS 0.031128f
C15496 DVDD.n11410 VSS 0.031128f
C15497 DVDD.n11411 VSS 0.031128f
C15498 DVDD.n11413 VSS 0.031128f
C15499 DVDD.n11414 VSS 0.031128f
C15500 DVDD.n11415 VSS 0.031128f
C15501 DVDD.n11417 VSS 0.031128f
C15502 DVDD.n11418 VSS 0.031128f
C15503 DVDD.n11419 VSS 0.031128f
C15504 DVDD.n11420 VSS 0.031128f
C15505 DVDD.n11421 VSS 0.031128f
C15506 DVDD.n11422 VSS 0.031128f
C15507 DVDD.n11423 VSS 0.031128f
C15508 DVDD.n11425 VSS 0.031128f
C15509 DVDD.n11426 VSS 0.031128f
C15510 DVDD.n11427 VSS 0.031128f
C15511 DVDD.n11429 VSS 0.031128f
C15512 DVDD.n11430 VSS 0.031128f
C15513 DVDD.n11431 VSS 0.031128f
C15514 DVDD.n11432 VSS 0.031128f
C15515 DVDD.n11433 VSS 0.031128f
C15516 DVDD.n11434 VSS 0.031128f
C15517 DVDD.n11435 VSS 0.031128f
C15518 DVDD.n11437 VSS 0.031128f
C15519 DVDD.n11438 VSS 0.031128f
C15520 DVDD.n11439 VSS 0.031128f
C15521 DVDD.n11441 VSS 0.031128f
C15522 DVDD.n11442 VSS 0.031128f
C15523 DVDD.n11443 VSS 0.031128f
C15524 DVDD.n11444 VSS 0.031128f
C15525 DVDD.n11445 VSS 0.031128f
C15526 DVDD.n11446 VSS 0.031128f
C15527 DVDD.n11447 VSS 0.031128f
C15528 DVDD.n11449 VSS 0.031128f
C15529 DVDD.n11450 VSS 0.031128f
C15530 DVDD.n11451 VSS 0.031128f
C15531 DVDD.n11453 VSS 0.031128f
C15532 DVDD.n11454 VSS 0.031128f
C15533 DVDD.n11455 VSS 0.031128f
C15534 DVDD.n11456 VSS 0.031128f
C15535 DVDD.n11457 VSS 0.031128f
C15536 DVDD.n11458 VSS 0.031128f
C15537 DVDD.n11459 VSS 0.031128f
C15538 DVDD.n11461 VSS 0.031128f
C15539 DVDD.n11462 VSS 0.031128f
C15540 DVDD.n11463 VSS 0.031128f
C15541 DVDD.n11465 VSS 0.031128f
C15542 DVDD.n11466 VSS 0.031128f
C15543 DVDD.n11467 VSS 0.031128f
C15544 DVDD.n11468 VSS 0.031128f
C15545 DVDD.n11469 VSS 0.031128f
C15546 DVDD.n11470 VSS 0.031128f
C15547 DVDD.n11471 VSS 0.031128f
C15548 DVDD.n11473 VSS 0.031128f
C15549 DVDD.n11474 VSS 0.031128f
C15550 DVDD.n11475 VSS 0.031128f
C15551 DVDD.n11477 VSS 0.031128f
C15552 DVDD.n11478 VSS 0.031128f
C15553 DVDD.n11479 VSS 0.031128f
C15554 DVDD.n11480 VSS 0.031128f
C15555 DVDD.n11481 VSS 0.031128f
C15556 DVDD.n11482 VSS 0.031128f
C15557 DVDD.n11483 VSS 0.031128f
C15558 DVDD.n11485 VSS 0.031128f
C15559 DVDD.n11486 VSS 0.031128f
C15560 DVDD.n11487 VSS 0.031128f
C15561 DVDD.n11489 VSS 0.031128f
C15562 DVDD.n11490 VSS 0.031128f
C15563 DVDD.n11491 VSS 0.031128f
C15564 DVDD.n11492 VSS 0.031128f
C15565 DVDD.n11493 VSS 0.031128f
C15566 DVDD.n11494 VSS 0.031128f
C15567 DVDD.n11495 VSS 0.031128f
C15568 DVDD.n11497 VSS 0.031128f
C15569 DVDD.n11498 VSS 0.031128f
C15570 DVDD.n11499 VSS 0.031128f
C15571 DVDD.n11501 VSS 0.031128f
C15572 DVDD.n11502 VSS 0.031128f
C15573 DVDD.n11503 VSS 0.031128f
C15574 DVDD.n11504 VSS 0.031128f
C15575 DVDD.n11505 VSS 0.031128f
C15576 DVDD.n11506 VSS 0.031128f
C15577 DVDD.n11507 VSS 0.031128f
C15578 DVDD.n11509 VSS 0.031128f
C15579 DVDD.n11510 VSS 0.031128f
C15580 DVDD.n11511 VSS 0.031128f
C15581 DVDD.n11513 VSS 0.031128f
C15582 DVDD.n11514 VSS 0.031128f
C15583 DVDD.n11515 VSS 0.031128f
C15584 DVDD.n11516 VSS 0.031128f
C15585 DVDD.n11517 VSS 0.031128f
C15586 DVDD.n11518 VSS 0.031128f
C15587 DVDD.n11519 VSS 0.031128f
C15588 DVDD.n11521 VSS 0.031128f
C15589 DVDD.n11522 VSS 0.031128f
C15590 DVDD.n11523 VSS 0.031128f
C15591 DVDD.n11525 VSS 0.031128f
C15592 DVDD.n11526 VSS 0.031128f
C15593 DVDD.n11527 VSS 0.031128f
C15594 DVDD.n11528 VSS 0.031128f
C15595 DVDD.n11529 VSS 0.031128f
C15596 DVDD.n11530 VSS 0.031128f
C15597 DVDD.n11531 VSS 0.031128f
C15598 DVDD.n11533 VSS 0.031128f
C15599 DVDD.n11534 VSS 0.031128f
C15600 DVDD.n11535 VSS 0.031128f
C15601 DVDD.n11537 VSS 0.031128f
C15602 DVDD.n11538 VSS 0.031128f
C15603 DVDD.n11539 VSS 0.031128f
C15604 DVDD.n11540 VSS 0.031128f
C15605 DVDD.n11541 VSS 0.031128f
C15606 DVDD.n11542 VSS 0.031128f
C15607 DVDD.n11543 VSS 0.031128f
C15608 DVDD.n11545 VSS 0.031128f
C15609 DVDD.n11546 VSS 0.031128f
C15610 DVDD.n11547 VSS 0.031128f
C15611 DVDD.n11549 VSS 0.031128f
C15612 DVDD.n11550 VSS 0.031128f
C15613 DVDD.n11551 VSS 0.031128f
C15614 DVDD.n11552 VSS 0.031128f
C15615 DVDD.n11553 VSS 0.031128f
C15616 DVDD.n11554 VSS 0.031128f
C15617 DVDD.n11555 VSS 0.031128f
C15618 DVDD.n11557 VSS 0.031128f
C15619 DVDD.n11558 VSS 0.031128f
C15620 DVDD.n11559 VSS 0.031128f
C15621 DVDD.n11561 VSS 0.031128f
C15622 DVDD.n11562 VSS 0.031128f
C15623 DVDD.n11563 VSS 0.031128f
C15624 DVDD.n11564 VSS 0.031128f
C15625 DVDD.n11565 VSS 0.025918f
C15626 DVDD.n11566 VSS 0.036621f
C15627 DVDD.n11567 VSS 0.041931f
C15628 DVDD.n11568 VSS 0.522252f
C15629 DVDD.n11569 VSS 0.036621f
C15630 DVDD.n11570 VSS 0.02566f
C15631 DVDD.n11571 VSS 0.029381f
C15632 DVDD.n11572 VSS 0.029381f
C15633 DVDD.n11573 VSS 0.522252f
C15634 DVDD.n11574 VSS 0.041931f
C15635 DVDD.n11575 VSS 0.029676f
C15636 DVDD.n11576 VSS 0.029676f
C15637 DVDD.n11577 VSS 0.02513f
C15638 DVDD.n11578 VSS 0.041931f
C15639 DVDD.n11579 VSS 0.025838f
C15640 DVDD.n11580 VSS 0.598063f
C15641 DVDD.n11581 VSS 0.349572f
C15642 DVDD.n11582 VSS 0.033945f
C15643 DVDD.n11583 VSS 0.033945f
C15644 DVDD.n11584 VSS 0.028497f
C15645 DVDD.n11585 VSS 0.03923f
C15646 DVDD.n11586 VSS 0.05956f
C15647 DVDD.n11587 VSS 0.05956f
C15648 DVDD.n11588 VSS 0.349572f
C15649 DVDD.n11630 VSS 0.019729f
C15650 DVDD.n11631 VSS 0.273761f
C15651 DVDD.n11632 VSS 0.02513f
C15652 DVDD.n11633 VSS 0.019729f
C15653 DVDD.n11634 VSS 0.031128f
C15654 DVDD.n11635 VSS 0.031128f
C15655 DVDD.n11636 VSS 0.031128f
C15656 DVDD.n11637 VSS 0.031128f
C15657 DVDD.n11638 VSS 0.031128f
C15658 DVDD.n11639 VSS 0.031128f
C15659 DVDD.n11640 VSS 0.031128f
C15660 DVDD.n11641 VSS 0.031128f
C15661 DVDD.n11642 VSS 0.031128f
C15662 DVDD.n11643 VSS 0.031128f
C15663 DVDD.n11644 VSS 0.031128f
C15664 DVDD.n11645 VSS 0.031128f
C15665 DVDD.n11646 VSS 0.031128f
C15666 DVDD.n11647 VSS 0.031128f
C15667 DVDD.n11648 VSS 0.031128f
C15668 DVDD.n11649 VSS 0.031128f
C15669 DVDD.n11650 VSS 0.031128f
C15670 DVDD.n11651 VSS 0.031128f
C15671 DVDD.n11652 VSS 0.031128f
C15672 DVDD.n11653 VSS 0.031128f
C15673 DVDD.n11654 VSS 0.031128f
C15674 DVDD.n11655 VSS 0.031128f
C15675 DVDD.n11656 VSS 0.031128f
C15676 DVDD.n11657 VSS 0.031128f
C15677 DVDD.n11658 VSS 0.031128f
C15678 DVDD.n11659 VSS 0.031128f
C15679 DVDD.n11660 VSS 0.031128f
C15680 DVDD.n11661 VSS 0.031128f
C15681 DVDD.n11662 VSS 0.031128f
C15682 DVDD.n11663 VSS 0.031128f
C15683 DVDD.n11664 VSS 0.031128f
C15684 DVDD.n11665 VSS 0.031128f
C15685 DVDD.n11666 VSS 0.031128f
C15686 DVDD.n11667 VSS 0.031128f
C15687 DVDD.n11668 VSS 0.031128f
C15688 DVDD.n11669 VSS 0.031128f
C15689 DVDD.n11670 VSS 0.031128f
C15690 DVDD.n11671 VSS 0.031128f
C15691 DVDD.n11672 VSS 0.031128f
C15692 DVDD.n11673 VSS 0.031128f
C15693 DVDD.n11674 VSS 0.019729f
C15694 DVDD.n11676 VSS 0.031128f
C15695 DVDD.n11677 VSS 0.031128f
C15696 DVDD.n11678 VSS 0.031128f
C15697 DVDD.n11679 VSS 0.031128f
C15698 DVDD.n11680 VSS 0.031128f
C15699 DVDD.n11681 VSS 0.031128f
C15700 DVDD.n11683 VSS 0.031128f
C15701 DVDD.n11684 VSS 0.031128f
C15702 DVDD.n11685 VSS 0.031128f
C15703 DVDD.n11687 VSS 0.031128f
C15704 DVDD.n11688 VSS 0.031128f
C15705 DVDD.n11689 VSS 0.031128f
C15706 DVDD.n11690 VSS 0.031128f
C15707 DVDD.n11691 VSS 0.031128f
C15708 DVDD.n11692 VSS 0.031128f
C15709 DVDD.n11693 VSS 0.031128f
C15710 DVDD.n11695 VSS 0.031128f
C15711 DVDD.n11696 VSS 0.031128f
C15712 DVDD.n11697 VSS 0.031128f
C15713 DVDD.n11699 VSS 0.031128f
C15714 DVDD.n11700 VSS 0.031128f
C15715 DVDD.n11701 VSS 0.031128f
C15716 DVDD.n11702 VSS 0.031128f
C15717 DVDD.n11703 VSS 0.031128f
C15718 DVDD.n11704 VSS 0.031128f
C15719 DVDD.n11705 VSS 0.031128f
C15720 DVDD.n11707 VSS 0.031128f
C15721 DVDD.n11708 VSS 0.031128f
C15722 DVDD.n11709 VSS 0.031128f
C15723 DVDD.n11711 VSS 0.031128f
C15724 DVDD.n11712 VSS 0.031128f
C15725 DVDD.n11713 VSS 0.031128f
C15726 DVDD.n11714 VSS 0.031128f
C15727 DVDD.n11715 VSS 0.031128f
C15728 DVDD.n11716 VSS 0.031128f
C15729 DVDD.n11717 VSS 0.031128f
C15730 DVDD.n11719 VSS 0.031128f
C15731 DVDD.n11720 VSS 0.031128f
C15732 DVDD.n11721 VSS 0.031128f
C15733 DVDD.n11723 VSS 0.031128f
C15734 DVDD.n11724 VSS 0.031128f
C15735 DVDD.n11725 VSS 0.031128f
C15736 DVDD.n11726 VSS 0.031128f
C15737 DVDD.n11727 VSS 0.031128f
C15738 DVDD.n11728 VSS 0.031128f
C15739 DVDD.n11729 VSS 0.031128f
C15740 DVDD.n11731 VSS 0.031128f
C15741 DVDD.n11732 VSS 0.031128f
C15742 DVDD.n11733 VSS 0.031128f
C15743 DVDD.n11735 VSS 0.031128f
C15744 DVDD.n11736 VSS 0.031128f
C15745 DVDD.n11737 VSS 0.031128f
C15746 DVDD.n11738 VSS 0.031128f
C15747 DVDD.n11739 VSS 0.031128f
C15748 DVDD.n11740 VSS 0.031128f
C15749 DVDD.n11741 VSS 0.031128f
C15750 DVDD.n11743 VSS 0.031128f
C15751 DVDD.n11744 VSS 0.031128f
C15752 DVDD.n11745 VSS 0.031128f
C15753 DVDD.n11747 VSS 0.031128f
C15754 DVDD.n11748 VSS 0.031128f
C15755 DVDD.n11749 VSS 0.031128f
C15756 DVDD.n11750 VSS 0.031128f
C15757 DVDD.n11751 VSS 0.031128f
C15758 DVDD.n11752 VSS 0.031128f
C15759 DVDD.n11753 VSS 0.031128f
C15760 DVDD.n11755 VSS 0.031128f
C15761 DVDD.n11756 VSS 0.031128f
C15762 DVDD.n11757 VSS 0.031128f
C15763 DVDD.n11759 VSS 0.031128f
C15764 DVDD.n11760 VSS 0.031128f
C15765 DVDD.n11761 VSS 0.031128f
C15766 DVDD.n11762 VSS 0.031128f
C15767 DVDD.n11763 VSS 0.031128f
C15768 DVDD.n11764 VSS 0.031128f
C15769 DVDD.n11765 VSS 0.031128f
C15770 DVDD.n11767 VSS 0.031128f
C15771 DVDD.n11768 VSS 0.031128f
C15772 DVDD.n11769 VSS 0.031128f
C15773 DVDD.n11771 VSS 0.031128f
C15774 DVDD.n11772 VSS 0.031128f
C15775 DVDD.n11773 VSS 0.031128f
C15776 DVDD.n11774 VSS 0.031128f
C15777 DVDD.n11775 VSS 0.031128f
C15778 DVDD.n11776 VSS 0.031128f
C15779 DVDD.n11777 VSS 0.031128f
C15780 DVDD.n11779 VSS 0.031128f
C15781 DVDD.n11780 VSS 0.031128f
C15782 DVDD.n11781 VSS 0.031128f
C15783 DVDD.n11783 VSS 0.031128f
C15784 DVDD.n11784 VSS 0.031128f
C15785 DVDD.n11785 VSS 0.031128f
C15786 DVDD.n11786 VSS 0.031128f
C15787 DVDD.n11787 VSS 0.031128f
C15788 DVDD.n11788 VSS 0.031128f
C15789 DVDD.n11789 VSS 0.031128f
C15790 DVDD.n11791 VSS 0.031128f
C15791 DVDD.n11792 VSS 0.031128f
C15792 DVDD.n11793 VSS 0.031128f
C15793 DVDD.n11795 VSS 0.031128f
C15794 DVDD.n11796 VSS 0.031128f
C15795 DVDD.n11797 VSS 0.031128f
C15796 DVDD.n11798 VSS 0.031128f
C15797 DVDD.n11799 VSS 0.031128f
C15798 DVDD.n11800 VSS 0.031128f
C15799 DVDD.n11801 VSS 0.031128f
C15800 DVDD.n11803 VSS 0.031128f
C15801 DVDD.n11804 VSS 0.031128f
C15802 DVDD.n11805 VSS 0.031128f
C15803 DVDD.n11807 VSS 0.031128f
C15804 DVDD.n11808 VSS 0.031128f
C15805 DVDD.n11809 VSS 0.031128f
C15806 DVDD.n11810 VSS 0.031128f
C15807 DVDD.n11811 VSS 0.031128f
C15808 DVDD.n11812 VSS 0.031128f
C15809 DVDD.n11813 VSS 0.031128f
C15810 DVDD.n11815 VSS 0.031128f
C15811 DVDD.n11816 VSS 0.031128f
C15812 DVDD.n11817 VSS 0.031128f
C15813 DVDD.n11819 VSS 0.031128f
C15814 DVDD.n11820 VSS 0.031128f
C15815 DVDD.n11821 VSS 0.031128f
C15816 DVDD.n11822 VSS 0.031128f
C15817 DVDD.n11823 VSS 0.031128f
C15818 DVDD.n11824 VSS 0.031128f
C15819 DVDD.n11825 VSS 0.031128f
C15820 DVDD.n11827 VSS 0.031128f
C15821 DVDD.n11828 VSS 0.031128f
C15822 DVDD.n11829 VSS 0.031128f
C15823 DVDD.n11831 VSS 0.031128f
C15824 DVDD.n11832 VSS 0.031128f
C15825 DVDD.n11833 VSS 0.031128f
C15826 DVDD.n11834 VSS 0.031128f
C15827 DVDD.n11835 VSS 0.031128f
C15828 DVDD.n11836 VSS 0.031128f
C15829 DVDD.n11837 VSS 0.031128f
C15830 DVDD.n11839 VSS 0.031128f
C15831 DVDD.n11840 VSS 0.031128f
C15832 DVDD.n11841 VSS 0.031128f
C15833 DVDD.n11843 VSS 0.031128f
C15834 DVDD.n11844 VSS 0.031128f
C15835 DVDD.n11845 VSS 0.031128f
C15836 DVDD.n11846 VSS 0.031128f
C15837 DVDD.n11847 VSS 0.031128f
C15838 DVDD.n11848 VSS 0.031128f
C15839 DVDD.n11849 VSS 0.031128f
C15840 DVDD.n11851 VSS 0.031128f
C15841 DVDD.n11852 VSS 0.031128f
C15842 DVDD.n11853 VSS 0.031128f
C15843 DVDD.n11855 VSS 0.031128f
C15844 DVDD.n11856 VSS 0.031128f
C15845 DVDD.n11857 VSS 0.031128f
C15846 DVDD.n11858 VSS 0.031128f
C15847 DVDD.n11859 VSS 0.031128f
C15848 DVDD.n11860 VSS 0.031128f
C15849 DVDD.n11861 VSS 0.031128f
C15850 DVDD.n11863 VSS 0.031128f
C15851 DVDD.n11864 VSS 0.031128f
C15852 DVDD.n11865 VSS 0.031128f
C15853 DVDD.n11867 VSS 0.031128f
C15854 DVDD.n11868 VSS 0.031128f
C15855 DVDD.n11869 VSS 0.031128f
C15856 DVDD.n11870 VSS 0.031128f
C15857 DVDD.n11871 VSS 0.031128f
C15858 DVDD.n11872 VSS 0.031128f
C15859 DVDD.n11873 VSS 0.031128f
C15860 DVDD.n11875 VSS 0.031128f
C15861 DVDD.n11876 VSS 0.031128f
C15862 DVDD.n11877 VSS 0.031128f
C15863 DVDD.n11879 VSS 0.031128f
C15864 DVDD.n11880 VSS 0.031128f
C15865 DVDD.n11881 VSS 0.031128f
C15866 DVDD.n11882 VSS 0.031128f
C15867 DVDD.n11883 VSS 0.031128f
C15868 DVDD.n11884 VSS 0.031128f
C15869 DVDD.n11885 VSS 0.031128f
C15870 DVDD.n11887 VSS 0.031128f
C15871 DVDD.n11888 VSS 0.031128f
C15872 DVDD.n11889 VSS 0.031128f
C15873 DVDD.n11891 VSS 0.031128f
C15874 DVDD.n11892 VSS 0.031128f
C15875 DVDD.n11893 VSS 0.031128f
C15876 DVDD.n11894 VSS 0.031128f
C15877 DVDD.n11895 VSS 0.031128f
C15878 DVDD.n11896 VSS 0.031128f
C15879 DVDD.n11897 VSS 0.031128f
C15880 DVDD.n11899 VSS 0.031128f
C15881 DVDD.n11900 VSS 0.031128f
C15882 DVDD.n11901 VSS 0.031128f
C15883 DVDD.n11903 VSS 0.031128f
C15884 DVDD.n11904 VSS 0.031128f
C15885 DVDD.n11905 VSS 0.031128f
C15886 DVDD.n11906 VSS 0.031128f
C15887 DVDD.n11907 VSS 0.031128f
C15888 DVDD.n11908 VSS 0.031128f
C15889 DVDD.n11909 VSS 0.031128f
C15890 DVDD.n11911 VSS 0.031128f
C15891 DVDD.n11912 VSS 0.031128f
C15892 DVDD.n11913 VSS 0.031128f
C15893 DVDD.n11915 VSS 0.031128f
C15894 DVDD.n11916 VSS 0.031128f
C15895 DVDD.n11917 VSS 0.031128f
C15896 DVDD.n11918 VSS 0.031128f
C15897 DVDD.n11919 VSS 0.022566f
C15898 DVDD.n11920 VSS 0.036621f
C15899 DVDD.n11921 VSS 0.025838f
C15900 DVDD.n11922 VSS 0.02513f
C15901 DVDD.n11923 VSS 0.041931f
C15902 DVDD.n11924 VSS 0.021999f
C15903 DVDD.n11925 VSS 0.598063f
C15904 DVDD.n11926 VSS 0.522253f
C15905 DVDD.n11927 VSS 0.034583f
C15906 DVDD.n11928 VSS 0.034583f
C15907 DVDD.n11929 VSS 0.423753f
C15908 DVDD.n11930 VSS 0.028497f
C15909 DVDD.n11931 VSS 0.053165f
C15910 DVDD.n11932 VSS 0.033945f
C15911 DVDD.n11933 VSS 0.05956f
C15912 DVDD.n11934 VSS 0.033945f
C15913 DVDD.n11935 VSS 0.05956f
C15914 DVDD.n11936 VSS 0.265338f
C15915 DVDD.n11937 VSS 0.387477f
C15916 DVDD.n11938 VSS 0.4675f
C15917 DVDD.n11939 VSS 0.598063f
C15918 DVDD.n11940 VSS 0.02513f
C15919 DVDD.n11941 VSS 0.039126f
C15920 DVDD.n11942 VSS 0.02513f
C15921 DVDD.n11943 VSS 0.039126f
C15922 DVDD.n11944 VSS 0.031128f
C15923 DVDD.n11945 VSS 0.031128f
C15924 DVDD.n11946 VSS 0.031128f
C15925 DVDD.n11948 VSS 0.031128f
C15926 DVDD.n11949 VSS 0.031128f
C15927 DVDD.n11950 VSS 0.031128f
C15928 DVDD.n11952 VSS 0.031128f
C15929 DVDD.n11953 VSS 0.031128f
C15930 DVDD.n11954 VSS 0.031128f
C15931 DVDD.n11956 VSS 0.031128f
C15932 DVDD.n11957 VSS 0.031128f
C15933 DVDD.n11958 VSS 0.031128f
C15934 DVDD.n11960 VSS 0.031128f
C15935 DVDD.n11961 VSS 0.031128f
C15936 DVDD.n11962 VSS 0.031128f
C15937 DVDD.n11964 VSS 0.031128f
C15938 DVDD.n11965 VSS 0.031128f
C15939 DVDD.n11966 VSS 0.031128f
C15940 DVDD.n11968 VSS 0.031128f
C15941 DVDD.n11969 VSS 0.031128f
C15942 DVDD.n11970 VSS 0.031128f
C15943 DVDD.n11972 VSS 0.031128f
C15944 DVDD.n11973 VSS 0.031128f
C15945 DVDD.n11974 VSS 0.031128f
C15946 DVDD.n11976 VSS 0.031128f
C15947 DVDD.n11977 VSS 0.031128f
C15948 DVDD.n11978 VSS 0.031128f
C15949 DVDD.n11980 VSS 0.031128f
C15950 DVDD.n11981 VSS 0.031128f
C15951 DVDD.n11982 VSS 0.031128f
C15952 DVDD.n11984 VSS 0.031128f
C15953 DVDD.n11985 VSS 0.031128f
C15954 DVDD.n11986 VSS 0.031128f
C15955 DVDD.n11988 VSS 0.031128f
C15956 DVDD.n11989 VSS 0.031128f
C15957 DVDD.n11990 VSS 0.031128f
C15958 DVDD.n11992 VSS 0.031128f
C15959 DVDD.n11993 VSS 0.031128f
C15960 DVDD.n11994 VSS 0.031128f
C15961 DVDD.n11996 VSS 0.031128f
C15962 DVDD.n11997 VSS 0.031128f
C15963 DVDD.n11998 VSS 0.031128f
C15964 DVDD.n12000 VSS 0.031128f
C15965 DVDD.n12001 VSS 0.031128f
C15966 DVDD.n12002 VSS 0.031128f
C15967 DVDD.n12004 VSS 0.031128f
C15968 DVDD.n12005 VSS 0.031128f
C15969 DVDD.n12006 VSS 0.031128f
C15970 DVDD.n12008 VSS 0.031128f
C15971 DVDD.n12009 VSS 0.031128f
C15972 DVDD.n12010 VSS 0.031128f
C15973 DVDD.n12012 VSS 0.031128f
C15974 DVDD.n12013 VSS 0.031128f
C15975 DVDD.n12014 VSS 0.031128f
C15976 DVDD.n12016 VSS 0.031128f
C15977 DVDD.n12017 VSS 0.031128f
C15978 DVDD.n12018 VSS 0.031128f
C15979 DVDD.n12020 VSS 0.031128f
C15980 DVDD.n12021 VSS 0.031128f
C15981 DVDD.n12022 VSS 0.031128f
C15982 DVDD.n12024 VSS 0.031128f
C15983 DVDD.n12025 VSS 0.031128f
C15984 DVDD.n12026 VSS 0.031128f
C15985 DVDD.n12027 VSS 0.019729f
C15986 DVDD.n12028 VSS 0.019729f
C15987 DVDD.n12030 VSS 0.031128f
C15988 DVDD.n12032 VSS 0.031128f
C15989 DVDD.n12034 VSS 0.031128f
C15990 DVDD.n12035 VSS 0.031128f
C15991 DVDD.n12036 VSS 0.031128f
C15992 DVDD.n12037 VSS 0.031128f
C15993 DVDD.n12038 VSS 0.031128f
C15994 DVDD.n12039 VSS 0.031128f
C15995 DVDD.n12040 VSS 0.031128f
C15996 DVDD.n12042 VSS 0.031128f
C15997 DVDD.n12044 VSS 0.031128f
C15998 DVDD.n12046 VSS 0.031128f
C15999 DVDD.n12047 VSS 0.031128f
C16000 DVDD.n12048 VSS 0.031128f
C16001 DVDD.n12049 VSS 0.031128f
C16002 DVDD.n12050 VSS 0.031128f
C16003 DVDD.n12051 VSS 0.031128f
C16004 DVDD.n12052 VSS 0.031128f
C16005 DVDD.n12054 VSS 0.031128f
C16006 DVDD.n12056 VSS 0.031128f
C16007 DVDD.n12058 VSS 0.031128f
C16008 DVDD.n12059 VSS 0.031128f
C16009 DVDD.n12060 VSS 0.031128f
C16010 DVDD.n12061 VSS 0.031128f
C16011 DVDD.n12062 VSS 0.031128f
C16012 DVDD.n12063 VSS 0.031128f
C16013 DVDD.n12064 VSS 0.031128f
C16014 DVDD.n12066 VSS 0.031128f
C16015 DVDD.n12068 VSS 0.031128f
C16016 DVDD.n12070 VSS 0.031128f
C16017 DVDD.n12071 VSS 0.031128f
C16018 DVDD.n12072 VSS 0.031128f
C16019 DVDD.n12073 VSS 0.031128f
C16020 DVDD.n12074 VSS 0.031128f
C16021 DVDD.n12075 VSS 0.031128f
C16022 DVDD.n12076 VSS 0.031128f
C16023 DVDD.n12078 VSS 0.031128f
C16024 DVDD.n12080 VSS 0.031128f
C16025 DVDD.n12082 VSS 0.031128f
C16026 DVDD.n12083 VSS 0.031128f
C16027 DVDD.n12084 VSS 0.031128f
C16028 DVDD.n12085 VSS 0.031128f
C16029 DVDD.n12086 VSS 0.031128f
C16030 DVDD.n12087 VSS 0.031128f
C16031 DVDD.n12088 VSS 0.031128f
C16032 DVDD.n12090 VSS 0.031128f
C16033 DVDD.n12092 VSS 0.031128f
C16034 DVDD.n12094 VSS 0.031128f
C16035 DVDD.n12095 VSS 0.031128f
C16036 DVDD.n12096 VSS 0.031128f
C16037 DVDD.n12097 VSS 0.031128f
C16038 DVDD.n12098 VSS 0.031128f
C16039 DVDD.n12099 VSS 0.031128f
C16040 DVDD.n12100 VSS 0.031128f
C16041 DVDD.n12102 VSS 0.031128f
C16042 DVDD.n12104 VSS 0.031128f
C16043 DVDD.n12106 VSS 0.031128f
C16044 DVDD.n12107 VSS 0.031128f
C16045 DVDD.n12108 VSS 0.031128f
C16046 DVDD.n12109 VSS 0.031128f
C16047 DVDD.n12110 VSS 0.031128f
C16048 DVDD.n12111 VSS 0.031128f
C16049 DVDD.n12112 VSS 0.031128f
C16050 DVDD.n12114 VSS 0.031128f
C16051 DVDD.n12116 VSS 0.031128f
C16052 DVDD.n12118 VSS 0.031128f
C16053 DVDD.n12119 VSS 0.031128f
C16054 DVDD.n12120 VSS 0.031128f
C16055 DVDD.n12121 VSS 0.031128f
C16056 DVDD.n12122 VSS 0.031128f
C16057 DVDD.n12123 VSS 0.031128f
C16058 DVDD.n12124 VSS 0.031128f
C16059 DVDD.n12126 VSS 0.031128f
C16060 DVDD.n12128 VSS 0.031128f
C16061 DVDD.n12130 VSS 0.031128f
C16062 DVDD.n12131 VSS 0.031128f
C16063 DVDD.n12132 VSS 0.031128f
C16064 DVDD.n12133 VSS 0.031128f
C16065 DVDD.n12134 VSS 0.031128f
C16066 DVDD.n12135 VSS 0.031128f
C16067 DVDD.n12136 VSS 0.031128f
C16068 DVDD.n12138 VSS 0.031128f
C16069 DVDD.n12140 VSS 0.031128f
C16070 DVDD.n12142 VSS 0.031128f
C16071 DVDD.n12143 VSS 0.031128f
C16072 DVDD.n12144 VSS 0.031128f
C16073 DVDD.n12145 VSS 0.031128f
C16074 DVDD.n12146 VSS 0.031128f
C16075 DVDD.n12147 VSS 0.031128f
C16076 DVDD.n12148 VSS 0.031128f
C16077 DVDD.n12150 VSS 0.031128f
C16078 DVDD.n12152 VSS 0.031128f
C16079 DVDD.n12154 VSS 0.031128f
C16080 DVDD.n12155 VSS 0.031128f
C16081 DVDD.n12156 VSS 0.031128f
C16082 DVDD.n12157 VSS 0.031128f
C16083 DVDD.n12158 VSS 0.031128f
C16084 DVDD.n12159 VSS 0.031128f
C16085 DVDD.n12160 VSS 0.031128f
C16086 DVDD.n12162 VSS 0.031128f
C16087 DVDD.n12164 VSS 0.031128f
C16088 DVDD.n12166 VSS 0.031128f
C16089 DVDD.n12167 VSS 0.031128f
C16090 DVDD.n12168 VSS 0.031128f
C16091 DVDD.n12169 VSS 0.031128f
C16092 DVDD.n12170 VSS 0.031128f
C16093 DVDD.n12171 VSS 0.031128f
C16094 DVDD.n12172 VSS 0.031128f
C16095 DVDD.n12174 VSS 0.031128f
C16096 DVDD.n12176 VSS 0.031128f
C16097 DVDD.n12178 VSS 0.031128f
C16098 DVDD.n12179 VSS 0.031128f
C16099 DVDD.n12180 VSS 0.031128f
C16100 DVDD.n12181 VSS 0.031128f
C16101 DVDD.n12182 VSS 0.031128f
C16102 DVDD.n12183 VSS 0.031128f
C16103 DVDD.n12184 VSS 0.031128f
C16104 DVDD.n12186 VSS 0.031128f
C16105 DVDD.n12188 VSS 0.031128f
C16106 DVDD.n12190 VSS 0.031128f
C16107 DVDD.n12191 VSS 0.031128f
C16108 DVDD.n12192 VSS 0.031128f
C16109 DVDD.n12193 VSS 0.031128f
C16110 DVDD.n12194 VSS 0.031128f
C16111 DVDD.n12195 VSS 0.031128f
C16112 DVDD.n12196 VSS 0.031128f
C16113 DVDD.n12198 VSS 0.031128f
C16114 DVDD.n12200 VSS 0.031128f
C16115 DVDD.n12202 VSS 0.031128f
C16116 DVDD.n12203 VSS 0.031128f
C16117 DVDD.n12204 VSS 0.031128f
C16118 DVDD.n12205 VSS 0.031128f
C16119 DVDD.n12206 VSS 0.031128f
C16120 DVDD.n12207 VSS 0.031128f
C16121 DVDD.n12208 VSS 0.031128f
C16122 DVDD.n12210 VSS 0.031128f
C16123 DVDD.n12212 VSS 0.031128f
C16124 DVDD.n12214 VSS 0.031128f
C16125 DVDD.n12215 VSS 0.031128f
C16126 DVDD.n12216 VSS 0.031128f
C16127 DVDD.n12217 VSS 0.031128f
C16128 DVDD.n12218 VSS 0.031128f
C16129 DVDD.n12219 VSS 0.031128f
C16130 DVDD.n12220 VSS 0.031128f
C16131 DVDD.n12222 VSS 0.031128f
C16132 DVDD.n12224 VSS 0.031128f
C16133 DVDD.n12226 VSS 0.031128f
C16134 DVDD.n12227 VSS 0.031128f
C16135 DVDD.n12228 VSS 0.031128f
C16136 DVDD.n12229 VSS 0.031128f
C16137 DVDD.n12230 VSS 0.031128f
C16138 DVDD.n12231 VSS 0.031128f
C16139 DVDD.n12232 VSS 0.031128f
C16140 DVDD.n12234 VSS 0.031128f
C16141 DVDD.n12236 VSS 0.031128f
C16142 DVDD.n12238 VSS 0.031128f
C16143 DVDD.n12239 VSS 0.031128f
C16144 DVDD.n12240 VSS 0.031128f
C16145 DVDD.n12241 VSS 0.031128f
C16146 DVDD.n12242 VSS 0.031128f
C16147 DVDD.n12243 VSS 0.031128f
C16148 DVDD.n12244 VSS 0.031128f
C16149 DVDD.n12246 VSS 0.031128f
C16150 DVDD.n12248 VSS 0.031128f
C16151 DVDD.n12250 VSS 0.031128f
C16152 DVDD.n12251 VSS 0.031128f
C16153 DVDD.n12252 VSS 0.031128f
C16154 DVDD.n12253 VSS 0.031128f
C16155 DVDD.n12254 VSS 0.031128f
C16156 DVDD.n12255 VSS 0.031128f
C16157 DVDD.n12256 VSS 0.031128f
C16158 DVDD.n12258 VSS 0.031128f
C16159 DVDD.n12260 VSS 0.031128f
C16160 DVDD.n12262 VSS 0.031128f
C16161 DVDD.n12263 VSS 0.031128f
C16162 DVDD.n12264 VSS 0.031128f
C16163 DVDD.n12265 VSS 0.031128f
C16164 DVDD.n12266 VSS 0.031128f
C16165 DVDD.n12267 VSS 0.031128f
C16166 DVDD.n12268 VSS 0.031128f
C16167 DVDD.n12269 VSS 0.031128f
C16168 DVDD.n12271 VSS 0.031128f
C16169 DVDD.n12273 VSS 0.031128f
C16170 DVDD.n12275 VSS 0.019729f
C16171 DVDD.n12276 VSS 0.019729f
C16172 DVDD.n12277 VSS 0.026086f
C16173 DVDD.n12278 VSS 0.021999f
C16174 DVDD.n12279 VSS 0.019213f
C16175 DVDD.n12280 VSS 0.028833f
C16176 DVDD.n12281 VSS 0.026086f
C16177 DVDD.n12282 VSS 0.036621f
C16178 DVDD.n12283 VSS 0.02513f
C16179 DVDD.n12284 VSS 0.041931f
C16180 DVDD.n12285 VSS 0.02513f
C16181 DVDD.n12286 VSS 0.041931f
C16182 DVDD.n12287 VSS 0.374843f
C16183 DVDD.n12329 VSS 0.019729f
C16184 DVDD.n12330 VSS 0.374843f
C16185 DVDD.n12331 VSS 0.019729f
C16186 DVDD.n12332 VSS 0.429595f
C16187 DVDD.n12333 VSS 0.315878f
C16188 DVDD.n12334 VSS 0.031128f
C16189 DVDD.n12335 VSS 0.031128f
C16190 DVDD.n12336 VSS 0.031128f
C16191 DVDD.n12337 VSS 0.031128f
C16192 DVDD.n12338 VSS 0.031128f
C16193 DVDD.n12339 VSS 0.031128f
C16194 DVDD.n12340 VSS 0.031128f
C16195 DVDD.n12341 VSS 0.031128f
C16196 DVDD.n12342 VSS 0.031128f
C16197 DVDD.n12343 VSS 0.031128f
C16198 DVDD.n12344 VSS 0.031128f
C16199 DVDD.n12345 VSS 0.031128f
C16200 DVDD.n12346 VSS 0.031128f
C16201 DVDD.n12347 VSS 0.031128f
C16202 DVDD.n12348 VSS 0.031128f
C16203 DVDD.n12349 VSS 0.031128f
C16204 DVDD.n12350 VSS 0.031128f
C16205 DVDD.n12351 VSS 0.031128f
C16206 DVDD.n12352 VSS 0.031128f
C16207 DVDD.n12353 VSS 0.031128f
C16208 DVDD.n12354 VSS 0.031128f
C16209 DVDD.n12355 VSS 0.031128f
C16210 DVDD.n12356 VSS 0.031128f
C16211 DVDD.n12357 VSS 0.031128f
C16212 DVDD.n12358 VSS 0.031128f
C16213 DVDD.n12359 VSS 0.031128f
C16214 DVDD.n12360 VSS 0.031128f
C16215 DVDD.n12361 VSS 0.031128f
C16216 DVDD.n12362 VSS 0.031128f
C16217 DVDD.n12363 VSS 0.031128f
C16218 DVDD.n12364 VSS 0.031128f
C16219 DVDD.n12365 VSS 0.031128f
C16220 DVDD.n12366 VSS 0.031128f
C16221 DVDD.n12367 VSS 0.031128f
C16222 DVDD.n12368 VSS 0.031128f
C16223 DVDD.n12369 VSS 0.031128f
C16224 DVDD.n12370 VSS 0.031128f
C16225 DVDD.n12371 VSS 0.031128f
C16226 DVDD.n12372 VSS 0.031128f
C16227 DVDD.n12373 VSS 0.031128f
C16228 DVDD.n12375 VSS 0.031128f
C16229 DVDD.n12376 VSS 0.031128f
C16230 DVDD.n12377 VSS 0.039516f
C16231 DVDD.n12378 VSS 0.036872f
C16232 DVDD.n12379 VSS 0.041308f
C16233 DVDD.n12380 VSS 0.05956f
C16234 DVDD.n12381 VSS 0.041308f
C16235 DVDD.n12382 VSS 0.033945f
C16236 DVDD.n12383 VSS 0.048033f
C16237 DVDD.n12384 VSS 0.039516f
C16238 DVDD.n12385 VSS 0.033945f
C16239 DVDD.n12386 VSS 0.05956f
C16240 DVDD.n12387 VSS 0.033945f
C16241 DVDD.n12388 VSS 0.522252f
C16242 DVDD.n12389 VSS 0.598063f
C16243 DVDD.n12390 VSS 0.522252f
C16244 DVDD.n12432 VSS 0.475924f
C16245 DVDD.n12433 VSS 0.031128f
C16246 DVDD.n12434 VSS 0.019729f
C16247 DVDD.n12435 VSS 0.134774f
C16248 DVDD.n12477 VSS 0.463288f
C16249 DVDD.n12478 VSS 0.02513f
C16250 DVDD.n12479 VSS 0.031128f
C16251 DVDD.n12480 VSS 0.031128f
C16252 DVDD.n12481 VSS 0.031128f
C16253 DVDD.n12482 VSS 0.031128f
C16254 DVDD.n12483 VSS 0.031128f
C16255 DVDD.n12484 VSS 0.031128f
C16256 DVDD.n12485 VSS 0.031128f
C16257 DVDD.n12486 VSS 0.031128f
C16258 DVDD.n12487 VSS 0.031128f
C16259 DVDD.n12488 VSS 0.031128f
C16260 DVDD.n12489 VSS 0.031128f
C16261 DVDD.n12490 VSS 0.031128f
C16262 DVDD.n12491 VSS 0.031128f
C16263 DVDD.n12492 VSS 0.031128f
C16264 DVDD.n12493 VSS 0.031128f
C16265 DVDD.n12494 VSS 0.031128f
C16266 DVDD.n12495 VSS 0.031128f
C16267 DVDD.n12496 VSS 0.031128f
C16268 DVDD.n12497 VSS 0.031128f
C16269 DVDD.n12498 VSS 0.031128f
C16270 DVDD.n12499 VSS 0.031128f
C16271 DVDD.n12500 VSS 0.031128f
C16272 DVDD.n12501 VSS 0.031128f
C16273 DVDD.n12502 VSS 0.031128f
C16274 DVDD.n12503 VSS 0.031128f
C16275 DVDD.n12504 VSS 0.031128f
C16276 DVDD.n12505 VSS 0.031128f
C16277 DVDD.n12506 VSS 0.031128f
C16278 DVDD.n12507 VSS 0.031128f
C16279 DVDD.n12508 VSS 0.031128f
C16280 DVDD.n12509 VSS 0.031128f
C16281 DVDD.n12510 VSS 0.031128f
C16282 DVDD.n12511 VSS 0.031128f
C16283 DVDD.n12512 VSS 0.031128f
C16284 DVDD.n12513 VSS 0.031128f
C16285 DVDD.n12514 VSS 0.031128f
C16286 DVDD.n12515 VSS 0.031128f
C16287 DVDD.n12516 VSS 0.031128f
C16288 DVDD.n12517 VSS 0.031128f
C16289 DVDD.n12518 VSS 0.031128f
C16290 DVDD.n12519 VSS 0.031128f
C16291 DVDD.n12520 VSS 0.031128f
C16292 DVDD.n12521 VSS 0.031128f
C16293 DVDD.n12522 VSS 0.031128f
C16294 DVDD.n12523 VSS 0.031128f
C16295 DVDD.n12524 VSS 0.031128f
C16296 DVDD.n12525 VSS 0.031128f
C16297 DVDD.n12526 VSS 0.031128f
C16298 DVDD.n12527 VSS 0.031128f
C16299 DVDD.n12528 VSS 0.031128f
C16300 DVDD.n12529 VSS 0.031128f
C16301 DVDD.n12530 VSS 0.031128f
C16302 DVDD.n12531 VSS 0.031128f
C16303 DVDD.n12532 VSS 0.031128f
C16304 DVDD.n12533 VSS 0.031128f
C16305 DVDD.n12534 VSS 0.031128f
C16306 DVDD.n12535 VSS 0.031128f
C16307 DVDD.n12536 VSS 0.031128f
C16308 DVDD.n12537 VSS 0.031128f
C16309 DVDD.n12538 VSS 0.031128f
C16310 DVDD.n12539 VSS 0.031128f
C16311 DVDD.n12540 VSS 0.031128f
C16312 DVDD.n12541 VSS 0.028497f
C16313 DVDD.n12542 VSS 0.031128f
C16314 DVDD.n12543 VSS 0.031128f
C16315 DVDD.n12544 VSS 0.031128f
C16316 DVDD.n12545 VSS 0.031128f
C16317 DVDD.n12546 VSS 0.031128f
C16318 DVDD.n12547 VSS 0.031128f
C16319 DVDD.n12548 VSS 0.031128f
C16320 DVDD.n12549 VSS 0.031128f
C16321 DVDD.n12550 VSS 0.031128f
C16322 DVDD.n12551 VSS 0.031128f
C16323 DVDD.n12552 VSS 0.031128f
C16324 DVDD.n12553 VSS 0.031128f
C16325 DVDD.n12554 VSS 0.031128f
C16326 DVDD.n12555 VSS 0.031128f
C16327 DVDD.n12556 VSS 0.031128f
C16328 DVDD.n12557 VSS 0.031128f
C16329 DVDD.n12558 VSS 0.031128f
C16330 DVDD.n12559 VSS 0.031128f
C16331 DVDD.n12560 VSS 0.031128f
C16332 DVDD.n12561 VSS 0.031128f
C16333 DVDD.n12562 VSS 0.031128f
C16334 DVDD.n12563 VSS 0.031128f
C16335 DVDD.n12564 VSS 0.031128f
C16336 DVDD.n12565 VSS 0.031128f
C16337 DVDD.n12566 VSS 0.031128f
C16338 DVDD.n12567 VSS 0.031128f
C16339 DVDD.n12568 VSS 0.031128f
C16340 DVDD.n12569 VSS 0.031128f
C16341 DVDD.n12570 VSS 0.031128f
C16342 DVDD.n12571 VSS 0.031128f
C16343 DVDD.n12572 VSS 0.031128f
C16344 DVDD.n12573 VSS 0.031128f
C16345 DVDD.n12574 VSS 0.031128f
C16346 DVDD.n12575 VSS 0.031128f
C16347 DVDD.n12576 VSS 0.031128f
C16348 DVDD.n12577 VSS 0.031128f
C16349 DVDD.n12578 VSS 0.031128f
C16350 DVDD.n12579 VSS 0.031128f
C16351 DVDD.n12580 VSS 0.031128f
C16352 DVDD.n12581 VSS 0.031128f
C16353 DVDD.n12582 VSS 0.031128f
C16354 DVDD.n12583 VSS 0.031128f
C16355 DVDD.n12584 VSS 0.031128f
C16356 DVDD.n12585 VSS 0.031128f
C16357 DVDD.n12586 VSS 0.031128f
C16358 DVDD.n12587 VSS 0.031128f
C16359 DVDD.n12588 VSS 0.031128f
C16360 DVDD.n12589 VSS 0.031128f
C16361 DVDD.n12590 VSS 0.031128f
C16362 DVDD.n12591 VSS 0.031128f
C16363 DVDD.n12592 VSS 0.031128f
C16364 DVDD.n12593 VSS 0.031128f
C16365 DVDD.n12594 VSS 0.031128f
C16366 DVDD.n12595 VSS 0.031128f
C16367 DVDD.n12596 VSS 0.031128f
C16368 DVDD.n12597 VSS 0.031128f
C16369 DVDD.n12598 VSS 0.031128f
C16370 DVDD.n12599 VSS 0.031128f
C16371 DVDD.n12600 VSS 0.031128f
C16372 DVDD.n12601 VSS 0.031128f
C16373 DVDD.n12602 VSS 0.031128f
C16374 DVDD.n12603 VSS 0.031128f
C16375 DVDD.n12604 VSS 0.031128f
C16376 DVDD.n12605 VSS 0.031128f
C16377 DVDD.n12606 VSS 0.031128f
C16378 DVDD.n12607 VSS 0.031128f
C16379 DVDD.n12608 VSS 0.031128f
C16380 DVDD.n12609 VSS 0.031128f
C16381 DVDD.n12610 VSS 0.031128f
C16382 DVDD.n12611 VSS 0.031128f
C16383 DVDD.n12612 VSS 0.031128f
C16384 DVDD.n12613 VSS 0.031128f
C16385 DVDD.n12614 VSS 0.031128f
C16386 DVDD.n12615 VSS 0.031128f
C16387 DVDD.n12616 VSS 0.031128f
C16388 DVDD.n12617 VSS 0.031128f
C16389 DVDD.n12618 VSS 0.031128f
C16390 DVDD.n12619 VSS 0.031128f
C16391 DVDD.n12620 VSS 0.031128f
C16392 DVDD.n12621 VSS 0.031128f
C16393 DVDD.n12622 VSS 0.031128f
C16394 DVDD.n12623 VSS 0.031128f
C16395 DVDD.n12624 VSS 0.031128f
C16396 DVDD.n12625 VSS 0.031128f
C16397 DVDD.n12626 VSS 0.031128f
C16398 DVDD.n12627 VSS 0.031128f
C16399 DVDD.n12628 VSS 0.031128f
C16400 DVDD.n12629 VSS 0.031128f
C16401 DVDD.n12630 VSS 0.031128f
C16402 DVDD.n12631 VSS 0.031128f
C16403 DVDD.n12632 VSS 0.031128f
C16404 DVDD.n12633 VSS 0.031128f
C16405 DVDD.n12634 VSS 0.031128f
C16406 DVDD.n12635 VSS 0.031128f
C16407 DVDD.n12636 VSS 0.031128f
C16408 DVDD.n12637 VSS 0.031128f
C16409 DVDD.n12638 VSS 0.031128f
C16410 DVDD.n12639 VSS 0.031128f
C16411 DVDD.n12640 VSS 0.031128f
C16412 DVDD.n12641 VSS 0.031128f
C16413 DVDD.n12642 VSS 0.031128f
C16414 DVDD.n12643 VSS 0.031128f
C16415 DVDD.n12644 VSS 0.031128f
C16416 DVDD.n12645 VSS 0.031128f
C16417 DVDD.n12646 VSS 0.031128f
C16418 DVDD.n12647 VSS 0.031128f
C16419 DVDD.n12648 VSS 0.031128f
C16420 DVDD.n12649 VSS 0.031128f
C16421 DVDD.n12650 VSS 0.031128f
C16422 DVDD.n12651 VSS 0.031128f
C16423 DVDD.n12652 VSS 0.031128f
C16424 DVDD.n12653 VSS 0.031128f
C16425 DVDD.n12654 VSS 0.031128f
C16426 DVDD.n12655 VSS 0.031128f
C16427 DVDD.n12656 VSS 0.031128f
C16428 DVDD.n12657 VSS 0.031128f
C16429 DVDD.n12658 VSS 0.031128f
C16430 DVDD.n12659 VSS 0.031128f
C16431 DVDD.n12660 VSS 0.031128f
C16432 DVDD.n12661 VSS 0.031128f
C16433 DVDD.n12662 VSS 0.031128f
C16434 DVDD.n12663 VSS 0.031128f
C16435 DVDD.n12664 VSS 0.031128f
C16436 DVDD.n12665 VSS 0.031128f
C16437 DVDD.n12666 VSS 0.031128f
C16438 DVDD.n12667 VSS 0.031128f
C16439 DVDD.n12668 VSS 0.031128f
C16440 DVDD.n12669 VSS 0.031128f
C16441 DVDD.n12670 VSS 0.031128f
C16442 DVDD.n12671 VSS 0.031128f
C16443 DVDD.n12672 VSS 0.031128f
C16444 DVDD.n12673 VSS 0.031128f
C16445 DVDD.n12674 VSS 0.031128f
C16446 DVDD.n12675 VSS 0.031128f
C16447 DVDD.n12676 VSS 0.031128f
C16448 DVDD.n12677 VSS 0.031128f
C16449 DVDD.n12678 VSS 0.031128f
C16450 DVDD.n12679 VSS 0.031128f
C16451 DVDD.n12680 VSS 0.031128f
C16452 DVDD.n12681 VSS 0.031128f
C16453 DVDD.n12682 VSS 0.031128f
C16454 DVDD.n12683 VSS 0.031128f
C16455 DVDD.n12684 VSS 0.031128f
C16456 DVDD.n12685 VSS 0.031128f
C16457 DVDD.n12686 VSS 0.031128f
C16458 DVDD.n12687 VSS 0.031128f
C16459 DVDD.n12688 VSS 0.031128f
C16460 DVDD.n12689 VSS 0.031128f
C16461 DVDD.n12690 VSS 0.031128f
C16462 DVDD.n12691 VSS 0.031128f
C16463 DVDD.n12692 VSS 0.031128f
C16464 DVDD.n12693 VSS 0.031128f
C16465 DVDD.n12694 VSS 0.031128f
C16466 DVDD.n12695 VSS 0.031128f
C16467 DVDD.n12696 VSS 0.031128f
C16468 DVDD.n12697 VSS 0.031128f
C16469 DVDD.n12698 VSS 0.031128f
C16470 DVDD.n12699 VSS 0.031128f
C16471 DVDD.n12700 VSS 0.031128f
C16472 DVDD.n12701 VSS 0.031128f
C16473 DVDD.n12702 VSS 0.031128f
C16474 DVDD.n12703 VSS 0.031128f
C16475 DVDD.n12704 VSS 0.031128f
C16476 DVDD.n12705 VSS 0.031128f
C16477 DVDD.n12706 VSS 0.031128f
C16478 DVDD.n12707 VSS 0.031128f
C16479 DVDD.n12708 VSS 0.031128f
C16480 DVDD.n12709 VSS 0.031128f
C16481 DVDD.n12710 VSS 0.031128f
C16482 DVDD.n12711 VSS 0.031128f
C16483 DVDD.n12712 VSS 0.031128f
C16484 DVDD.n12713 VSS 0.031128f
C16485 DVDD.n12714 VSS 0.031128f
C16486 DVDD.n12715 VSS 0.031128f
C16487 DVDD.n12716 VSS 0.031128f
C16488 DVDD.n12717 VSS 0.031128f
C16489 DVDD.n12718 VSS 0.031128f
C16490 DVDD.n12719 VSS 0.031128f
C16491 DVDD.n12720 VSS 0.031128f
C16492 DVDD.n12721 VSS 0.031128f
C16493 DVDD.n12722 VSS 0.031128f
C16494 DVDD.n12723 VSS 0.031128f
C16495 DVDD.n12724 VSS 0.031128f
C16496 DVDD.n12725 VSS 0.026086f
C16497 DVDD.n12726 VSS 0.035287f
C16498 DVDD.n12727 VSS 0.035287f
C16499 DVDD.n12728 VSS 0.041931f
C16500 DVDD.n12729 VSS 0.027609f
C16501 DVDD.n12730 VSS 0.030818f
C16502 DVDD.n12731 VSS 0.028833f
C16503 DVDD.n12732 VSS 0.028833f
C16504 DVDD.n12733 VSS 0.02513f
C16505 DVDD.n12734 VSS 0.041931f
C16506 DVDD.n12735 VSS 0.02513f
C16507 DVDD.n12736 VSS 0.522252f
C16508 DVDD.n12737 VSS 0.598063f
C16509 DVDD.n12779 VSS 0.585428f
C16510 DVDD.n12780 VSS 0.031128f
C16511 DVDD.n12781 VSS 0.033945f
C16512 DVDD.n12782 VSS 0.019729f
C16513 DVDD.n12783 VSS 0.227432f
C16514 DVDD.n12825 VSS 0.585428f
C16515 DVDD.n12826 VSS 0.031128f
C16516 DVDD.n12827 VSS 0.031128f
C16517 DVDD.n12828 VSS 0.031128f
C16518 DVDD.n12829 VSS 0.031128f
C16519 DVDD.n12830 VSS 0.031128f
C16520 DVDD.n12831 VSS 0.031128f
C16521 DVDD.n12832 VSS 0.031128f
C16522 DVDD.n12833 VSS 0.031128f
C16523 DVDD.n12834 VSS 0.031128f
C16524 DVDD.n12835 VSS 0.031128f
C16525 DVDD.n12836 VSS 0.031128f
C16526 DVDD.n12837 VSS 0.031128f
C16527 DVDD.n12838 VSS 0.031128f
C16528 DVDD.n12839 VSS 0.031128f
C16529 DVDD.n12840 VSS 0.031128f
C16530 DVDD.n12841 VSS 0.031128f
C16531 DVDD.n12842 VSS 0.031128f
C16532 DVDD.n12843 VSS 0.031128f
C16533 DVDD.n12844 VSS 0.031128f
C16534 DVDD.n12845 VSS 0.031128f
C16535 DVDD.n12846 VSS 0.031128f
C16536 DVDD.n12847 VSS 0.031128f
C16537 DVDD.n12848 VSS 0.031128f
C16538 DVDD.n12849 VSS 0.031128f
C16539 DVDD.n12850 VSS 0.031128f
C16540 DVDD.n12851 VSS 0.031128f
C16541 DVDD.n12852 VSS 0.031128f
C16542 DVDD.n12853 VSS 0.031128f
C16543 DVDD.n12854 VSS 0.031128f
C16544 DVDD.n12855 VSS 0.031128f
C16545 DVDD.n12856 VSS 0.031128f
C16546 DVDD.n12857 VSS 0.031128f
C16547 DVDD.n12858 VSS 0.031128f
C16548 DVDD.n12859 VSS 0.031128f
C16549 DVDD.n12860 VSS 0.031128f
C16550 DVDD.n12861 VSS 0.031128f
C16551 DVDD.n12862 VSS 0.031128f
C16552 DVDD.n12863 VSS 0.031128f
C16553 DVDD.n12864 VSS 0.031128f
C16554 DVDD.n12865 VSS 0.031128f
C16555 DVDD.n12866 VSS 0.031128f
C16556 DVDD.n12867 VSS 0.031128f
C16557 DVDD.n12868 VSS 0.031128f
C16558 DVDD.n12869 VSS 0.031128f
C16559 DVDD.n12870 VSS 0.031128f
C16560 DVDD.n12871 VSS 0.031128f
C16561 DVDD.n12872 VSS 0.031128f
C16562 DVDD.n12873 VSS 0.031128f
C16563 DVDD.n12874 VSS 0.031128f
C16564 DVDD.n12875 VSS 0.031128f
C16565 DVDD.n12876 VSS 0.031128f
C16566 DVDD.n12877 VSS 0.031128f
C16567 DVDD.n12878 VSS 0.031128f
C16568 DVDD.n12879 VSS 0.031128f
C16569 DVDD.n12880 VSS 0.031128f
C16570 DVDD.n12881 VSS 0.031128f
C16571 DVDD.n12882 VSS 0.031128f
C16572 DVDD.n12883 VSS 0.031128f
C16573 DVDD.n12884 VSS 0.031128f
C16574 DVDD.n12885 VSS 0.031128f
C16575 DVDD.n12886 VSS 0.031128f
C16576 DVDD.n12887 VSS 0.031128f
C16577 DVDD.n12888 VSS 0.048877f
C16578 DVDD.n12889 VSS 0.053165f
C16579 DVDD.n12890 VSS 0.05956f
C16580 DVDD.n12891 VSS 0.053165f
C16581 DVDD.n12892 VSS 0.036872f
C16582 DVDD.n12893 VSS 0.041308f
C16583 DVDD.n12894 VSS 0.041308f
C16584 DVDD.n12895 VSS 0.05956f
C16585 DVDD.n12896 VSS 0.054757f
C16586 DVDD.n12897 VSS 0.054757f
C16587 DVDD.n12898 VSS 0.033945f
C16588 DVDD.n12899 VSS 0.05956f
C16589 DVDD.n12900 VSS 0.031701f
C16590 DVDD.n12901 VSS 0.501194f
C16591 DVDD.n12902 VSS 0.031701f
C16592 DVDD.n12903 VSS 0.028497f
C16593 DVDD.n12904 VSS 0.0343f
C16594 DVDD.n12905 VSS 0.053165f
C16595 DVDD.n12906 VSS 0.033945f
C16596 DVDD.n12907 VSS 0.05956f
C16597 DVDD.n12908 VSS 0.033945f
C16598 DVDD.n12909 VSS 0.033945f
C16599 DVDD.n12910 VSS 0.038426f
C16600 DVDD.n12911 VSS 0.05956f
C16601 DVDD.n12912 VSS 0.44223f
C16602 DVDD.n12913 VSS 0.02513f
C16603 DVDD.n12914 VSS 0.02513f
C16604 DVDD.n12915 VSS 0.026086f
C16605 DVDD.n12916 VSS 0.036621f
C16606 DVDD.n12917 VSS 0.041931f
C16607 DVDD.n12918 VSS 0.027466f
C16608 DVDD.n12919 VSS 0.031448f
C16609 DVDD.n12920 VSS 0.031448f
C16610 DVDD.n12921 VSS 0.522252f
C16611 DVDD.n12922 VSS 0.041931f
C16612 DVDD.n12964 VSS 0.031128f
C16613 DVDD.n12966 VSS 0.031128f
C16614 DVDD.n12967 VSS 0.031128f
C16615 DVDD.n12968 VSS 0.031128f
C16616 DVDD.n12969 VSS 0.031128f
C16617 DVDD.n12970 VSS 0.031128f
C16618 DVDD.n12971 VSS 0.031128f
C16619 DVDD.n12972 VSS 0.031128f
C16620 DVDD.n12973 VSS 0.031128f
C16621 DVDD.n12974 VSS 0.031128f
C16622 DVDD.n12975 VSS 0.031128f
C16623 DVDD.n12976 VSS 0.031128f
C16624 DVDD.n12977 VSS 0.031128f
C16625 DVDD.n12978 VSS 0.031128f
C16626 DVDD.n12979 VSS 0.031128f
C16627 DVDD.n12980 VSS 0.031128f
C16628 DVDD.n12981 VSS 0.031128f
C16629 DVDD.n12982 VSS 0.031128f
C16630 DVDD.n12983 VSS 0.031128f
C16631 DVDD.n12984 VSS 0.031128f
C16632 DVDD.n12985 VSS 0.031128f
C16633 DVDD.n12986 VSS 0.031128f
C16634 DVDD.n12987 VSS 0.031128f
C16635 DVDD.n12988 VSS 0.031128f
C16636 DVDD.n12989 VSS 0.031128f
C16637 DVDD.n12990 VSS 0.031128f
C16638 DVDD.n12991 VSS 0.031128f
C16639 DVDD.n12992 VSS 0.031128f
C16640 DVDD.n12993 VSS 0.031128f
C16641 DVDD.n12994 VSS 0.031128f
C16642 DVDD.n12995 VSS 0.031128f
C16643 DVDD.n12996 VSS 0.031128f
C16644 DVDD.n12997 VSS 0.031128f
C16645 DVDD.n12998 VSS 0.031128f
C16646 DVDD.n12999 VSS 0.031128f
C16647 DVDD.n13000 VSS 0.031128f
C16648 DVDD.n13001 VSS 0.031128f
C16649 DVDD.n13002 VSS 0.031128f
C16650 DVDD.n13003 VSS 0.031128f
C16651 DVDD.n13004 VSS 0.031128f
C16652 DVDD.n13005 VSS 0.031128f
C16653 DVDD.n13006 VSS 0.031128f
C16654 DVDD.n13007 VSS 0.019729f
C16655 DVDD.n13008 VSS 0.019729f
C16656 DVDD.n13009 VSS 0.031128f
C16657 DVDD.n13010 VSS 0.031128f
C16658 DVDD.n13011 VSS 0.031128f
C16659 DVDD.n13012 VSS 0.031128f
C16660 DVDD.n13014 VSS 0.031128f
C16661 DVDD.n13015 VSS 0.031128f
C16662 DVDD.n13016 VSS 0.031128f
C16663 DVDD.n13017 VSS 0.031128f
C16664 DVDD.n13019 VSS 0.031128f
C16665 DVDD.n13020 VSS 0.031128f
C16666 DVDD.n13021 VSS 0.031128f
C16667 DVDD.n13022 VSS 0.031128f
C16668 DVDD.n13023 VSS 0.031128f
C16669 DVDD.n13024 VSS 0.031128f
C16670 DVDD.n13026 VSS 0.031128f
C16671 DVDD.n13027 VSS 0.031128f
C16672 DVDD.n13028 VSS 0.031128f
C16673 DVDD.n13029 VSS 0.031128f
C16674 DVDD.n13031 VSS 0.031128f
C16675 DVDD.n13032 VSS 0.031128f
C16676 DVDD.n13033 VSS 0.031128f
C16677 DVDD.n13034 VSS 0.031128f
C16678 DVDD.n13035 VSS 0.031128f
C16679 DVDD.n13036 VSS 0.031128f
C16680 DVDD.n13038 VSS 0.031128f
C16681 DVDD.n13039 VSS 0.031128f
C16682 DVDD.n13040 VSS 0.031128f
C16683 DVDD.n13041 VSS 0.031128f
C16684 DVDD.n13043 VSS 0.031128f
C16685 DVDD.n13044 VSS 0.031128f
C16686 DVDD.n13045 VSS 0.031128f
C16687 DVDD.n13046 VSS 0.031128f
C16688 DVDD.n13047 VSS 0.031128f
C16689 DVDD.n13048 VSS 0.031128f
C16690 DVDD.n13050 VSS 0.031128f
C16691 DVDD.n13051 VSS 0.031128f
C16692 DVDD.n13052 VSS 0.031128f
C16693 DVDD.n13053 VSS 0.031128f
C16694 DVDD.n13055 VSS 0.031128f
C16695 DVDD.n13056 VSS 0.031128f
C16696 DVDD.n13057 VSS 0.031128f
C16697 DVDD.n13058 VSS 0.031128f
C16698 DVDD.n13059 VSS 0.031128f
C16699 DVDD.n13060 VSS 0.031128f
C16700 DVDD.n13062 VSS 0.031128f
C16701 DVDD.n13063 VSS 0.031128f
C16702 DVDD.n13064 VSS 0.031128f
C16703 DVDD.n13065 VSS 0.031128f
C16704 DVDD.n13067 VSS 0.031128f
C16705 DVDD.n13068 VSS 0.031128f
C16706 DVDD.n13069 VSS 0.031128f
C16707 DVDD.n13070 VSS 0.031128f
C16708 DVDD.n13071 VSS 0.031128f
C16709 DVDD.n13072 VSS 0.031128f
C16710 DVDD.n13074 VSS 0.031128f
C16711 DVDD.n13075 VSS 0.031128f
C16712 DVDD.n13076 VSS 0.031128f
C16713 DVDD.n13077 VSS 0.031128f
C16714 DVDD.n13079 VSS 0.031128f
C16715 DVDD.n13080 VSS 0.031128f
C16716 DVDD.n13081 VSS 0.031128f
C16717 DVDD.n13082 VSS 0.031128f
C16718 DVDD.n13083 VSS 0.031128f
C16719 DVDD.n13084 VSS 0.031128f
C16720 DVDD.n13086 VSS 0.031128f
C16721 DVDD.n13087 VSS 0.031128f
C16722 DVDD.n13088 VSS 0.031128f
C16723 DVDD.n13089 VSS 0.031128f
C16724 DVDD.n13091 VSS 0.031128f
C16725 DVDD.n13092 VSS 0.031128f
C16726 DVDD.n13093 VSS 0.031128f
C16727 DVDD.n13094 VSS 0.031128f
C16728 DVDD.n13095 VSS 0.031128f
C16729 DVDD.n13096 VSS 0.031128f
C16730 DVDD.n13098 VSS 0.031128f
C16731 DVDD.n13099 VSS 0.031128f
C16732 DVDD.n13100 VSS 0.031128f
C16733 DVDD.n13101 VSS 0.031128f
C16734 DVDD.n13103 VSS 0.031128f
C16735 DVDD.n13104 VSS 0.031128f
C16736 DVDD.n13105 VSS 0.031128f
C16737 DVDD.n13106 VSS 0.031128f
C16738 DVDD.n13107 VSS 0.031128f
C16739 DVDD.n13108 VSS 0.031128f
C16740 DVDD.n13110 VSS 0.031128f
C16741 DVDD.n13111 VSS 0.031128f
C16742 DVDD.n13112 VSS 0.031128f
C16743 DVDD.n13113 VSS 0.031128f
C16744 DVDD.n13115 VSS 0.031128f
C16745 DVDD.n13116 VSS 0.031128f
C16746 DVDD.n13117 VSS 0.031128f
C16747 DVDD.n13118 VSS 0.031128f
C16748 DVDD.n13119 VSS 0.031128f
C16749 DVDD.n13120 VSS 0.031128f
C16750 DVDD.n13122 VSS 0.031128f
C16751 DVDD.n13123 VSS 0.031128f
C16752 DVDD.n13124 VSS 0.031128f
C16753 DVDD.n13125 VSS 0.031128f
C16754 DVDD.n13127 VSS 0.031128f
C16755 DVDD.n13128 VSS 0.031128f
C16756 DVDD.n13129 VSS 0.031128f
C16757 DVDD.n13130 VSS 0.031128f
C16758 DVDD.n13131 VSS 0.031128f
C16759 DVDD.n13132 VSS 0.031128f
C16760 DVDD.n13134 VSS 0.031128f
C16761 DVDD.n13135 VSS 0.031128f
C16762 DVDD.n13136 VSS 0.031128f
C16763 DVDD.n13137 VSS 0.031128f
C16764 DVDD.n13139 VSS 0.031128f
C16765 DVDD.n13140 VSS 0.031128f
C16766 DVDD.n13141 VSS 0.031128f
C16767 DVDD.n13142 VSS 0.031128f
C16768 DVDD.n13143 VSS 0.031128f
C16769 DVDD.n13144 VSS 0.031128f
C16770 DVDD.n13146 VSS 0.031128f
C16771 DVDD.n13147 VSS 0.031128f
C16772 DVDD.n13148 VSS 0.031128f
C16773 DVDD.n13149 VSS 0.031128f
C16774 DVDD.n13151 VSS 0.031128f
C16775 DVDD.n13152 VSS 0.031128f
C16776 DVDD.n13153 VSS 0.031128f
C16777 DVDD.n13154 VSS 0.031128f
C16778 DVDD.n13155 VSS 0.031128f
C16779 DVDD.n13156 VSS 0.031128f
C16780 DVDD.n13158 VSS 0.031128f
C16781 DVDD.n13159 VSS 0.031128f
C16782 DVDD.n13160 VSS 0.031128f
C16783 DVDD.n13161 VSS 0.031128f
C16784 DVDD.n13163 VSS 0.031128f
C16785 DVDD.n13164 VSS 0.031128f
C16786 DVDD.n13165 VSS 0.031128f
C16787 DVDD.n13166 VSS 0.031128f
C16788 DVDD.n13167 VSS 0.031128f
C16789 DVDD.n13168 VSS 0.031128f
C16790 DVDD.n13170 VSS 0.031128f
C16791 DVDD.n13171 VSS 0.031128f
C16792 DVDD.n13172 VSS 0.031128f
C16793 DVDD.n13173 VSS 0.031128f
C16794 DVDD.n13175 VSS 0.031128f
C16795 DVDD.n13176 VSS 0.031128f
C16796 DVDD.n13177 VSS 0.031128f
C16797 DVDD.n13178 VSS 0.031128f
C16798 DVDD.n13179 VSS 0.031128f
C16799 DVDD.n13180 VSS 0.031128f
C16800 DVDD.n13182 VSS 0.031128f
C16801 DVDD.n13183 VSS 0.031128f
C16802 DVDD.n13184 VSS 0.031128f
C16803 DVDD.n13185 VSS 0.031128f
C16804 DVDD.n13187 VSS 0.031128f
C16805 DVDD.n13188 VSS 0.031128f
C16806 DVDD.n13189 VSS 0.031128f
C16807 DVDD.n13190 VSS 0.031128f
C16808 DVDD.n13191 VSS 0.031128f
C16809 DVDD.n13192 VSS 0.031128f
C16810 DVDD.n13194 VSS 0.031128f
C16811 DVDD.n13195 VSS 0.031128f
C16812 DVDD.n13196 VSS 0.031128f
C16813 DVDD.n13197 VSS 0.031128f
C16814 DVDD.n13199 VSS 0.031128f
C16815 DVDD.n13200 VSS 0.031128f
C16816 DVDD.n13201 VSS 0.031128f
C16817 DVDD.n13202 VSS 0.031128f
C16818 DVDD.n13203 VSS 0.031128f
C16819 DVDD.n13204 VSS 0.031128f
C16820 DVDD.n13206 VSS 0.031128f
C16821 DVDD.n13207 VSS 0.031128f
C16822 DVDD.n13208 VSS 0.031128f
C16823 DVDD.n13209 VSS 0.031128f
C16824 DVDD.n13211 VSS 0.031128f
C16825 DVDD.n13212 VSS 0.031128f
C16826 DVDD.n13213 VSS 0.031128f
C16827 DVDD.n13214 VSS 0.031128f
C16828 DVDD.n13215 VSS 0.031128f
C16829 DVDD.n13216 VSS 0.031128f
C16830 DVDD.n13218 VSS 0.031128f
C16831 DVDD.n13219 VSS 0.031128f
C16832 DVDD.n13220 VSS 0.031128f
C16833 DVDD.n13221 VSS 0.031128f
C16834 DVDD.n13223 VSS 0.031128f
C16835 DVDD.n13224 VSS 0.031128f
C16836 DVDD.n13225 VSS 0.031128f
C16837 DVDD.n13226 VSS 0.031128f
C16838 DVDD.n13227 VSS 0.031128f
C16839 DVDD.n13228 VSS 0.031128f
C16840 DVDD.n13230 VSS 0.031128f
C16841 DVDD.n13231 VSS 0.031128f
C16842 DVDD.n13232 VSS 0.031128f
C16843 DVDD.n13233 VSS 0.031128f
C16844 DVDD.n13235 VSS 0.031128f
C16845 DVDD.n13236 VSS 0.031128f
C16846 DVDD.n13237 VSS 0.031128f
C16847 DVDD.n13238 VSS 0.031128f
C16848 DVDD.n13239 VSS 0.031128f
C16849 DVDD.n13240 VSS 0.031128f
C16850 DVDD.n13242 VSS 0.031128f
C16851 DVDD.n13243 VSS 0.031128f
C16852 DVDD.n13244 VSS 0.031128f
C16853 DVDD.n13245 VSS 0.031128f
C16854 DVDD.n13247 VSS 0.031128f
C16855 DVDD.n13248 VSS 0.031128f
C16856 DVDD.n13249 VSS 0.031128f
C16857 DVDD.n13250 VSS 0.031128f
C16858 DVDD.n13251 VSS 0.031128f
C16859 DVDD.n13252 VSS 0.031128f
C16860 DVDD.n13253 VSS 0.019729f
C16861 DVDD.n13254 VSS 0.019729f
C16862 DVDD.n13256 VSS 0.366419f
C16863 DVDD.n13257 VSS 0.501194f
C16864 DVDD.n13258 VSS 0.252702f
C16865 DVDD.n13259 VSS 0.027609f
C16866 DVDD.n13260 VSS 0.027609f
C16867 DVDD.n13261 VSS 0.024113f
C16868 DVDD.n13262 VSS 0.028833f
C16869 DVDD.n13263 VSS 0.030818f
C16870 DVDD.n13264 VSS 0.035287f
C16871 DVDD.n13265 VSS 0.035287f
C16872 DVDD.n13266 VSS 0.176891f
C16873 DVDD.n13267 VSS 0.374843f
C16874 DVDD.n13268 VSS 0.522252f
C16875 DVDD.n13269 VSS 0.598063f
C16876 DVDD.n13270 VSS 0.057639f
C16877 DVDD.n13271 VSS 0.057639f
C16878 DVDD.n13272 VSS 0.05145f
C16879 DVDD.n13273 VSS 0.039516f
C16880 DVDD.n13274 VSS 0.028297f
C16881 DVDD.n13275 VSS 0.053165f
C16882 DVDD.n13276 VSS 0.05956f
C16883 DVDD.n13277 VSS 0.05956f
C16884 DVDD.n13278 VSS 0.05956f
C16885 DVDD.n13279 VSS 0.034583f
C16886 DVDD.n13280 VSS 0.034583f
C16887 DVDD.n13281 VSS 0.03087f
C16888 DVDD.n13282 VSS 0.039516f
C16889 DVDD.n13283 VSS 0.028497f
C16890 DVDD.n13284 VSS 0.031128f
C16891 DVDD.n13285 VSS 0.031128f
C16892 DVDD.n13286 VSS 0.031128f
C16893 DVDD.n13287 VSS 0.031128f
C16894 DVDD.n13288 VSS 0.031128f
C16895 DVDD.n13289 VSS 0.031128f
C16896 DVDD.n13290 VSS 0.031128f
C16897 DVDD.n13291 VSS 0.031128f
C16898 DVDD.n13292 VSS 0.031128f
C16899 DVDD.n13293 VSS 0.031128f
C16900 DVDD.n13294 VSS 0.031128f
C16901 DVDD.n13295 VSS 0.031128f
C16902 DVDD.n13296 VSS 0.031128f
C16903 DVDD.n13297 VSS 0.031128f
C16904 DVDD.n13298 VSS 0.031128f
C16905 DVDD.n13299 VSS 0.031128f
C16906 DVDD.n13300 VSS 0.031128f
C16907 DVDD.n13301 VSS 0.031128f
C16908 DVDD.n13302 VSS 0.031128f
C16909 DVDD.n13303 VSS 0.031128f
C16910 DVDD.n13304 VSS 0.031128f
C16911 DVDD.n13305 VSS 0.031128f
C16912 DVDD.n13306 VSS 0.031128f
C16913 DVDD.n13307 VSS 0.031128f
C16914 DVDD.n13308 VSS 0.031128f
C16915 DVDD.n13309 VSS 0.031128f
C16916 DVDD.n13310 VSS 0.031128f
C16917 DVDD.n13311 VSS 0.031128f
C16918 DVDD.n13312 VSS 0.031128f
C16919 DVDD.n13313 VSS 0.031128f
C16920 DVDD.n13314 VSS 0.031128f
C16921 DVDD.n13315 VSS 0.031128f
C16922 DVDD.n13316 VSS 0.031128f
C16923 DVDD.n13317 VSS 0.031128f
C16924 DVDD.n13318 VSS 0.031128f
C16925 DVDD.n13319 VSS 0.031128f
C16926 DVDD.n13320 VSS 0.031128f
C16927 DVDD.n13321 VSS 0.031128f
C16928 DVDD.n13322 VSS 0.031128f
C16929 DVDD.n13323 VSS 0.031128f
C16930 DVDD.n13324 VSS 0.031128f
C16931 DVDD.n13325 VSS 0.031128f
C16932 DVDD.n13326 VSS 0.031128f
C16933 DVDD.n13327 VSS 0.031128f
C16934 DVDD.n13328 VSS 0.031128f
C16935 DVDD.n13329 VSS 0.031128f
C16936 DVDD.n13330 VSS 0.031128f
C16937 DVDD.n13331 VSS 0.031128f
C16938 DVDD.n13332 VSS 0.031128f
C16939 DVDD.n13333 VSS 0.031128f
C16940 DVDD.n13334 VSS 0.031128f
C16941 DVDD.n13335 VSS 0.031128f
C16942 DVDD.n13336 VSS 0.031128f
C16943 DVDD.n13337 VSS 0.031128f
C16944 DVDD.n13338 VSS 0.031128f
C16945 DVDD.n13339 VSS 0.031128f
C16946 DVDD.n13340 VSS 0.031128f
C16947 DVDD.n13341 VSS 0.031128f
C16948 DVDD.n13342 VSS 0.031128f
C16949 DVDD.n13343 VSS 0.031128f
C16950 DVDD.n13344 VSS 0.031128f
C16951 DVDD.n13345 VSS 0.031128f
C16952 DVDD.n13346 VSS 0.031128f
C16953 DVDD.n13347 VSS 0.031128f
C16954 DVDD.n13348 VSS 0.031128f
C16955 DVDD.n13349 VSS 0.031128f
C16956 DVDD.n13350 VSS 0.031128f
C16957 DVDD.n13351 VSS 0.031128f
C16958 DVDD.n13352 VSS 0.031128f
C16959 DVDD.n13353 VSS 0.031128f
C16960 DVDD.n13354 VSS 0.031128f
C16961 DVDD.n13355 VSS 0.031128f
C16962 DVDD.n13356 VSS 0.031128f
C16963 DVDD.n13357 VSS 0.031128f
C16964 DVDD.n13358 VSS 0.031128f
C16965 DVDD.n13359 VSS 0.031128f
C16966 DVDD.n13360 VSS 0.031128f
C16967 DVDD.n13361 VSS 0.031128f
C16968 DVDD.n13362 VSS 0.031128f
C16969 DVDD.n13363 VSS 0.031128f
C16970 DVDD.n13364 VSS 0.031128f
C16971 DVDD.n13365 VSS 0.031128f
C16972 DVDD.n13366 VSS 0.031128f
C16973 DVDD.n13367 VSS 0.031128f
C16974 DVDD.n13368 VSS 0.031128f
C16975 DVDD.n13369 VSS 0.031128f
C16976 DVDD.n13370 VSS 0.031128f
C16977 DVDD.n13371 VSS 0.031128f
C16978 DVDD.n13372 VSS 0.031128f
C16979 DVDD.n13373 VSS 0.031128f
C16980 DVDD.n13374 VSS 0.031128f
C16981 DVDD.n13375 VSS 0.031128f
C16982 DVDD.n13376 VSS 0.031128f
C16983 DVDD.n13377 VSS 0.031128f
C16984 DVDD.n13378 VSS 0.031128f
C16985 DVDD.n13379 VSS 0.031128f
C16986 DVDD.n13380 VSS 0.031128f
C16987 DVDD.n13381 VSS 0.031128f
C16988 DVDD.n13382 VSS 0.031128f
C16989 DVDD.n13383 VSS 0.031128f
C16990 DVDD.n13384 VSS 0.031128f
C16991 DVDD.n13385 VSS 0.031128f
C16992 DVDD.n13386 VSS 0.031128f
C16993 DVDD.n13387 VSS 0.031128f
C16994 DVDD.n13388 VSS 0.031128f
C16995 DVDD.n13389 VSS 0.031128f
C16996 DVDD.n13390 VSS 0.031128f
C16997 DVDD.n13391 VSS 0.031128f
C16998 DVDD.n13392 VSS 0.031128f
C16999 DVDD.n13393 VSS 0.031128f
C17000 DVDD.n13394 VSS 0.031128f
C17001 DVDD.n13395 VSS 0.031128f
C17002 DVDD.n13396 VSS 0.031128f
C17003 DVDD.n13397 VSS 0.031128f
C17004 DVDD.n13398 VSS 0.031128f
C17005 DVDD.n13399 VSS 0.031128f
C17006 DVDD.n13400 VSS 0.031128f
C17007 DVDD.n13401 VSS 0.031128f
C17008 DVDD.n13402 VSS 0.031128f
C17009 DVDD.n13403 VSS 0.031128f
C17010 DVDD.n13404 VSS 0.031128f
C17011 DVDD.n13405 VSS 0.031128f
C17012 DVDD.n13406 VSS 0.031128f
C17013 DVDD.n13407 VSS 0.031128f
C17014 DVDD.n13408 VSS 0.031128f
C17015 DVDD.n13409 VSS 0.031128f
C17016 DVDD.n13410 VSS 0.031128f
C17017 DVDD.n13411 VSS 0.031128f
C17018 DVDD.n13412 VSS 0.031128f
C17019 DVDD.n13413 VSS 0.031128f
C17020 DVDD.n13414 VSS 0.031128f
C17021 DVDD.n13415 VSS 0.031128f
C17022 DVDD.n13416 VSS 0.031128f
C17023 DVDD.n13417 VSS 0.031128f
C17024 DVDD.n13418 VSS 0.031128f
C17025 DVDD.n13419 VSS 0.031128f
C17026 DVDD.n13420 VSS 0.031128f
C17027 DVDD.n13421 VSS 0.031128f
C17028 DVDD.n13422 VSS 0.031128f
C17029 DVDD.n13423 VSS 0.031128f
C17030 DVDD.n13424 VSS 0.031128f
C17031 DVDD.n13425 VSS 0.031128f
C17032 DVDD.n13426 VSS 0.031128f
C17033 DVDD.n13427 VSS 0.031128f
C17034 DVDD.n13428 VSS 0.031128f
C17035 DVDD.n13429 VSS 0.031128f
C17036 DVDD.n13430 VSS 0.031128f
C17037 DVDD.n13431 VSS 0.031128f
C17038 DVDD.n13432 VSS 0.031128f
C17039 DVDD.n13433 VSS 0.031128f
C17040 DVDD.n13434 VSS 0.031128f
C17041 DVDD.n13435 VSS 0.031128f
C17042 DVDD.n13436 VSS 0.031128f
C17043 DVDD.n13437 VSS 0.031128f
C17044 DVDD.n13438 VSS 0.031128f
C17045 DVDD.n13439 VSS 0.031128f
C17046 DVDD.n13440 VSS 0.031128f
C17047 DVDD.n13441 VSS 0.031128f
C17048 DVDD.n13442 VSS 0.031128f
C17049 DVDD.n13443 VSS 0.031128f
C17050 DVDD.n13444 VSS 0.031128f
C17051 DVDD.n13445 VSS 0.031128f
C17052 DVDD.n13446 VSS 0.031128f
C17053 DVDD.n13447 VSS 0.031128f
C17054 DVDD.n13448 VSS 0.031128f
C17055 DVDD.n13449 VSS 0.031128f
C17056 DVDD.n13450 VSS 0.031128f
C17057 DVDD.n13451 VSS 0.031128f
C17058 DVDD.n13452 VSS 0.031128f
C17059 DVDD.n13453 VSS 0.031128f
C17060 DVDD.n13454 VSS 0.031128f
C17061 DVDD.n13455 VSS 0.031128f
C17062 DVDD.n13456 VSS 0.031128f
C17063 DVDD.n13457 VSS 0.031128f
C17064 DVDD.n13458 VSS 0.031128f
C17065 DVDD.n13459 VSS 0.031128f
C17066 DVDD.n13460 VSS 0.031128f
C17067 DVDD.n13461 VSS 0.031128f
C17068 DVDD.n13462 VSS 0.031128f
C17069 DVDD.n13463 VSS 0.031128f
C17070 DVDD.n13464 VSS 0.031128f
C17071 DVDD.n13465 VSS 0.031128f
C17072 DVDD.n13466 VSS 0.031128f
C17073 DVDD.n13467 VSS 0.026086f
C17074 DVDD.n13468 VSS 0.019729f
C17075 DVDD.n13469 VSS 0.019729f
C17076 DVDD.n13470 VSS 0.307455f
C17077 DVDD.n13471 VSS 0.019729f
C17078 DVDD.n13473 VSS 0.383266f
C17079 DVDD.n13474 VSS 0.151621f
C17080 DVDD.n13475 VSS 0.031448f
C17081 DVDD.n13476 VSS 0.031448f
C17082 DVDD.n13477 VSS 0.027466f
C17083 DVDD.n13478 VSS 0.036621f
C17084 DVDD.n13479 VSS 0.024113f
C17085 DVDD.n13480 VSS 0.027609f
C17086 DVDD.n13481 VSS 0.02513f
C17087 DVDD.n13482 VSS 0.019729f
C17088 DVDD.n13483 VSS 0.019729f
C17089 DVDD.n13484 VSS 0.522252f
C17090 DVDD.n13485 VSS 0.019729f
C17091 DVDD.n13487 VSS 0.509617f
C17092 DVDD.n13488 VSS 0.134774f
C17093 DVDD.n13489 VSS 0.048033f
C17094 DVDD.n13490 VSS 0.048033f
C17095 DVDD.n13491 VSS 0.042875f
C17096 DVDD.n13492 VSS 0.053165f
C17097 DVDD.n13493 VSS 0.042875f
C17098 DVDD.n13494 VSS 0.048033f
C17099 DVDD.n13495 VSS 0.033945f
C17100 DVDD.n13496 VSS 0.019729f
C17101 DVDD.n13497 VSS 0.028497f
C17102 DVDD.n13498 VSS 0.031128f
C17103 DVDD.n13499 VSS 0.031128f
C17104 DVDD.n13500 VSS 0.031128f
C17105 DVDD.n13501 VSS 0.031128f
C17106 DVDD.n13503 VSS 0.031128f
C17107 DVDD.n13504 VSS 0.031128f
C17108 DVDD.n13505 VSS 0.031128f
C17109 DVDD.n13507 VSS 0.031128f
C17110 DVDD.n13508 VSS 0.031128f
C17111 DVDD.n13509 VSS 0.031128f
C17112 DVDD.n13510 VSS 0.031128f
C17113 DVDD.n13511 VSS 0.031128f
C17114 DVDD.n13512 VSS 0.031128f
C17115 DVDD.n13513 VSS 0.031128f
C17116 DVDD.n13515 VSS 0.031128f
C17117 DVDD.n13516 VSS 0.031128f
C17118 DVDD.n13517 VSS 0.031128f
C17119 DVDD.n13519 VSS 0.031128f
C17120 DVDD.n13520 VSS 0.031128f
C17121 DVDD.n13521 VSS 0.031128f
C17122 DVDD.n13522 VSS 0.031128f
C17123 DVDD.n13523 VSS 0.031128f
C17124 DVDD.n13524 VSS 0.031128f
C17125 DVDD.n13525 VSS 0.031128f
C17126 DVDD.n13527 VSS 0.031128f
C17127 DVDD.n13528 VSS 0.031128f
C17128 DVDD.n13529 VSS 0.031128f
C17129 DVDD.n13531 VSS 0.031128f
C17130 DVDD.n13532 VSS 0.031128f
C17131 DVDD.n13533 VSS 0.031128f
C17132 DVDD.n13534 VSS 0.031128f
C17133 DVDD.n13535 VSS 0.031128f
C17134 DVDD.n13536 VSS 0.031128f
C17135 DVDD.n13537 VSS 0.031128f
C17136 DVDD.n13539 VSS 0.031128f
C17137 DVDD.n13540 VSS 0.031128f
C17138 DVDD.n13541 VSS 0.031128f
C17139 DVDD.n13543 VSS 0.031128f
C17140 DVDD.n13544 VSS 0.031128f
C17141 DVDD.n13545 VSS 0.031128f
C17142 DVDD.n13546 VSS 0.031128f
C17143 DVDD.n13547 VSS 0.031128f
C17144 DVDD.n13548 VSS 0.031128f
C17145 DVDD.n13549 VSS 0.031128f
C17146 DVDD.n13551 VSS 0.031128f
C17147 DVDD.n13552 VSS 0.031128f
C17148 DVDD.n13553 VSS 0.031128f
C17149 DVDD.n13555 VSS 0.031128f
C17150 DVDD.n13556 VSS 0.031128f
C17151 DVDD.n13557 VSS 0.031128f
C17152 DVDD.n13558 VSS 0.031128f
C17153 DVDD.n13559 VSS 0.031128f
C17154 DVDD.n13560 VSS 0.031128f
C17155 DVDD.n13561 VSS 0.031128f
C17156 DVDD.n13563 VSS 0.031128f
C17157 DVDD.n13564 VSS 0.031128f
C17158 DVDD.n13565 VSS 0.031128f
C17159 DVDD.n13567 VSS 0.031128f
C17160 DVDD.n13568 VSS 0.031128f
C17161 DVDD.n13569 VSS 0.031128f
C17162 DVDD.n13570 VSS 0.031128f
C17163 DVDD.n13571 VSS 0.031128f
C17164 DVDD.n13572 VSS 0.031128f
C17165 DVDD.n13573 VSS 0.031128f
C17166 DVDD.n13575 VSS 0.031128f
C17167 DVDD.n13576 VSS 0.031128f
C17168 DVDD.n13577 VSS 0.031128f
C17169 DVDD.n13579 VSS 0.031128f
C17170 DVDD.n13580 VSS 0.031128f
C17171 DVDD.n13581 VSS 0.031128f
C17172 DVDD.n13582 VSS 0.031128f
C17173 DVDD.n13583 VSS 0.031128f
C17174 DVDD.n13584 VSS 0.031128f
C17175 DVDD.n13585 VSS 0.031128f
C17176 DVDD.n13587 VSS 0.031128f
C17177 DVDD.n13588 VSS 0.031128f
C17178 DVDD.n13589 VSS 0.031128f
C17179 DVDD.n13591 VSS 0.031128f
C17180 DVDD.n13592 VSS 0.031128f
C17181 DVDD.n13593 VSS 0.031128f
C17182 DVDD.n13594 VSS 0.031128f
C17183 DVDD.n13595 VSS 0.031128f
C17184 DVDD.n13596 VSS 0.031128f
C17185 DVDD.n13597 VSS 0.031128f
C17186 DVDD.n13599 VSS 0.031128f
C17187 DVDD.n13600 VSS 0.031128f
C17188 DVDD.n13601 VSS 0.031128f
C17189 DVDD.n13603 VSS 0.031128f
C17190 DVDD.n13604 VSS 0.031128f
C17191 DVDD.n13605 VSS 0.031128f
C17192 DVDD.n13606 VSS 0.031128f
C17193 DVDD.n13607 VSS 0.031128f
C17194 DVDD.n13608 VSS 0.031128f
C17195 DVDD.n13609 VSS 0.031128f
C17196 DVDD.n13611 VSS 0.031128f
C17197 DVDD.n13612 VSS 0.031128f
C17198 DVDD.n13613 VSS 0.031128f
C17199 DVDD.n13615 VSS 0.031128f
C17200 DVDD.n13616 VSS 0.031128f
C17201 DVDD.n13617 VSS 0.031128f
C17202 DVDD.n13618 VSS 0.031128f
C17203 DVDD.n13619 VSS 0.031128f
C17204 DVDD.n13620 VSS 0.031128f
C17205 DVDD.n13621 VSS 0.031128f
C17206 DVDD.n13623 VSS 0.031128f
C17207 DVDD.n13624 VSS 0.031128f
C17208 DVDD.n13625 VSS 0.031128f
C17209 DVDD.n13627 VSS 0.031128f
C17210 DVDD.n13628 VSS 0.031128f
C17211 DVDD.n13629 VSS 0.031128f
C17212 DVDD.n13630 VSS 0.031128f
C17213 DVDD.n13631 VSS 0.031128f
C17214 DVDD.n13632 VSS 0.031128f
C17215 DVDD.n13633 VSS 0.031128f
C17216 DVDD.n13635 VSS 0.031128f
C17217 DVDD.n13636 VSS 0.031128f
C17218 DVDD.n13637 VSS 0.031128f
C17219 DVDD.n13639 VSS 0.031128f
C17220 DVDD.n13640 VSS 0.031128f
C17221 DVDD.n13641 VSS 0.031128f
C17222 DVDD.n13642 VSS 0.031128f
C17223 DVDD.n13643 VSS 0.031128f
C17224 DVDD.n13644 VSS 0.031128f
C17225 DVDD.n13645 VSS 0.031128f
C17226 DVDD.n13647 VSS 0.031128f
C17227 DVDD.n13648 VSS 0.031128f
C17228 DVDD.n13649 VSS 0.031128f
C17229 DVDD.n13651 VSS 0.031128f
C17230 DVDD.n13652 VSS 0.031128f
C17231 DVDD.n13653 VSS 0.031128f
C17232 DVDD.n13654 VSS 0.031128f
C17233 DVDD.n13655 VSS 0.031128f
C17234 DVDD.n13656 VSS 0.031128f
C17235 DVDD.n13657 VSS 0.031128f
C17236 DVDD.n13659 VSS 0.031128f
C17237 DVDD.n13660 VSS 0.031128f
C17238 DVDD.n13661 VSS 0.031128f
C17239 DVDD.n13663 VSS 0.031128f
C17240 DVDD.n13664 VSS 0.031128f
C17241 DVDD.n13665 VSS 0.031128f
C17242 DVDD.n13666 VSS 0.031128f
C17243 DVDD.n13667 VSS 0.031128f
C17244 DVDD.n13668 VSS 0.031128f
C17245 DVDD.n13669 VSS 0.031128f
C17246 DVDD.n13671 VSS 0.031128f
C17247 DVDD.n13672 VSS 0.031128f
C17248 DVDD.n13673 VSS 0.031128f
C17249 DVDD.n13675 VSS 0.031128f
C17250 DVDD.n13676 VSS 0.031128f
C17251 DVDD.n13677 VSS 0.031128f
C17252 DVDD.n13678 VSS 0.031128f
C17253 DVDD.n13679 VSS 0.031128f
C17254 DVDD.n13680 VSS 0.031128f
C17255 DVDD.n13681 VSS 0.031128f
C17256 DVDD.n13683 VSS 0.031128f
C17257 DVDD.n13684 VSS 0.031128f
C17258 DVDD.n13685 VSS 0.031128f
C17259 DVDD.n13687 VSS 0.031128f
C17260 DVDD.n13688 VSS 0.031128f
C17261 DVDD.n13689 VSS 0.031128f
C17262 DVDD.n13690 VSS 0.031128f
C17263 DVDD.n13691 VSS 0.031128f
C17264 DVDD.n13692 VSS 0.031128f
C17265 DVDD.n13693 VSS 0.031128f
C17266 DVDD.n13695 VSS 0.031128f
C17267 DVDD.n13696 VSS 0.031128f
C17268 DVDD.n13697 VSS 0.031128f
C17269 DVDD.n13699 VSS 0.031128f
C17270 DVDD.n13700 VSS 0.031128f
C17271 DVDD.n13701 VSS 0.031128f
C17272 DVDD.n13702 VSS 0.031128f
C17273 DVDD.n13703 VSS 0.031128f
C17274 DVDD.n13704 VSS 0.031128f
C17275 DVDD.n13705 VSS 0.031128f
C17276 DVDD.n13707 VSS 0.031128f
C17277 DVDD.n13708 VSS 0.031128f
C17278 DVDD.n13709 VSS 0.031128f
C17279 DVDD.n13711 VSS 0.031128f
C17280 DVDD.n13712 VSS 0.031128f
C17281 DVDD.n13713 VSS 0.031128f
C17282 DVDD.n13714 VSS 0.031128f
C17283 DVDD.n13715 VSS 0.031128f
C17284 DVDD.n13716 VSS 0.031128f
C17285 DVDD.n13717 VSS 0.031128f
C17286 DVDD.n13719 VSS 0.031128f
C17287 DVDD.n13720 VSS 0.031128f
C17288 DVDD.n13721 VSS 0.031128f
C17289 DVDD.n13723 VSS 0.031128f
C17290 DVDD.n13724 VSS 0.031128f
C17291 DVDD.n13725 VSS 0.031128f
C17292 DVDD.n13726 VSS 0.031128f
C17293 DVDD.n13727 VSS 0.031128f
C17294 DVDD.n13728 VSS 0.031128f
C17295 DVDD.n13729 VSS 0.031128f
C17296 DVDD.n13731 VSS 0.031128f
C17297 DVDD.n13732 VSS 0.031128f
C17298 DVDD.n13733 VSS 0.031128f
C17299 DVDD.n13735 VSS 0.031128f
C17300 DVDD.n13736 VSS 0.031128f
C17301 DVDD.n13737 VSS 0.031128f
C17302 DVDD.n13738 VSS 0.031128f
C17303 DVDD.n13739 VSS 0.031128f
C17304 DVDD.n13740 VSS 0.031128f
C17305 DVDD.n13741 VSS 0.031128f
C17306 DVDD.n13743 VSS 0.019729f
C17307 DVDD.n13744 VSS 0.240068f
C17308 DVDD.n13745 VSS 0.505405f
C17309 DVDD.n13746 VSS 0.023771f
C17310 DVDD.n13747 VSS 0.023771f
C17311 DVDD.n13748 VSS 0.02076f
C17312 DVDD.n13749 VSS 0.028833f
C17313 DVDD.n13750 VSS 0.034171f
C17314 DVDD.n13751 VSS 0.035718f
C17315 DVDD.n13752 VSS 0.040897f
C17316 DVDD.n13753 VSS 0.040897f
C17317 DVDD.n13754 VSS 0.522252f
C17318 DVDD.n13755 VSS 0.265338f
C17319 DVDD.n13756 VSS 0.054757f
C17320 DVDD.n13757 VSS 0.054757f
C17321 DVDD.n13758 VSS 0.048877f
C17322 DVDD.n13759 VSS 0.039516f
C17323 DVDD.n13760 VSS 0.03087f
C17324 DVDD.n13761 VSS 0.040516f
C17325 DVDD.n13762 VSS 0.05956f
C17326 DVDD.n13763 VSS 0.05956f
C17327 DVDD.n13764 VSS 0.332725f
C17328 DVDD.n13765 VSS 0.522252f
C17329 DVDD.n13766 VSS 0.041931f
C17330 DVDD.n13767 VSS 0.037059f
C17331 DVDD.n13768 VSS 0.037059f
C17332 DVDD.n13769 VSS 0.032366f
C17333 DVDD.n13770 VSS 0.028833f
C17334 DVDD.n13771 VSS 0.026086f
C17335 DVDD.n13772 VSS 0.031128f
C17336 DVDD.n13773 VSS 0.031128f
C17337 DVDD.n13774 VSS 0.031128f
C17338 DVDD.n13776 VSS 0.019729f
C17339 DVDD.n13777 VSS 0.425383f
C17340 DVDD.n13778 VSS 0.421171f
C17341 DVDD.n13779 VSS 0.031701f
C17342 DVDD.n13780 VSS 0.031701f
C17343 DVDD.n13781 VSS 0.028297f
C17344 DVDD.n13782 VSS 0.039516f
C17345 DVDD.n13783 VSS 0.05145f
C17346 DVDD.n13784 VSS 0.057639f
C17347 DVDD.n13785 VSS 0.057639f
C17348 DVDD.n13786 VSS 0.421171f
C17349 DVDD.n13787 VSS 0.522252f
C17350 DVDD.n13788 VSS 0.041931f
C17351 DVDD.n13789 VSS 0.03322f
C17352 DVDD.n13790 VSS 0.03322f
C17353 DVDD.n13791 VSS 0.029013f
C17354 DVDD.n13792 VSS 0.028833f
C17355 DVDD.n13793 VSS 0.026086f
C17356 DVDD.n13794 VSS 0.031128f
C17357 DVDD.n13795 VSS 0.031128f
C17358 DVDD.n13796 VSS 0.031128f
C17359 DVDD.n13798 VSS 0.019729f
C17360 DVDD.n13799 VSS 0.19795f
C17361 DVDD.n13800 VSS 0.543311f
C17362 DVDD.n13801 VSS 0.038426f
C17363 DVDD.n13802 VSS 0.038426f
C17364 DVDD.n13803 VSS 0.0343f
C17365 DVDD.n13804 VSS 0.039516f
C17366 DVDD.n13805 VSS 0.045447f
C17367 DVDD.n13806 VSS 0.050915f
C17368 DVDD.n13807 VSS 0.050915f
C17369 DVDD.n13808 VSS 0.05956f
C17370 DVDD.n13809 VSS 0.045151f
C17371 DVDD.n13810 VSS 0.045151f
C17372 DVDD.n13811 VSS 0.040302f
C17373 DVDD.n13812 VSS 0.039516f
C17374 DVDD.n13813 VSS 0.028497f
C17375 DVDD.n13814 VSS 0.031128f
C17376 DVDD.n13815 VSS 0.031128f
C17377 DVDD.n13816 VSS 0.031128f
C17378 DVDD.n13817 VSS 0.031128f
C17379 DVDD.n13818 VSS 0.031128f
C17380 DVDD.n13819 VSS 0.031128f
C17381 DVDD.n13820 VSS 0.031128f
C17382 DVDD.n13821 VSS 0.031128f
C17383 DVDD.n13822 VSS 0.031128f
C17384 DVDD.n13823 VSS 0.031128f
C17385 DVDD.n13824 VSS 0.031128f
C17386 DVDD.n13825 VSS 0.031128f
C17387 DVDD.n13826 VSS 0.031128f
C17388 DVDD.n13827 VSS 0.031128f
C17389 DVDD.n13828 VSS 0.031128f
C17390 DVDD.n13829 VSS 0.031128f
C17391 DVDD.n13830 VSS 0.031128f
C17392 DVDD.n13831 VSS 0.031128f
C17393 DVDD.n13832 VSS 0.031128f
C17394 DVDD.n13833 VSS 0.031128f
C17395 DVDD.n13834 VSS 0.031128f
C17396 DVDD.n13835 VSS 0.031128f
C17397 DVDD.n13836 VSS 0.031128f
C17398 DVDD.n13837 VSS 0.031128f
C17399 DVDD.n13838 VSS 0.031128f
C17400 DVDD.n13839 VSS 0.031128f
C17401 DVDD.n13840 VSS 0.031128f
C17402 DVDD.n13841 VSS 0.031128f
C17403 DVDD.n13842 VSS 0.031128f
C17404 DVDD.n13843 VSS 0.031128f
C17405 DVDD.n13844 VSS 0.031128f
C17406 DVDD.n13845 VSS 0.031128f
C17407 DVDD.n13846 VSS 0.031128f
C17408 DVDD.n13847 VSS 0.031128f
C17409 DVDD.n13848 VSS 0.031128f
C17410 DVDD.n13849 VSS 0.031128f
C17411 DVDD.n13850 VSS 0.031128f
C17412 DVDD.n13851 VSS 0.031128f
C17413 DVDD.n13852 VSS 0.031128f
C17414 DVDD.n13853 VSS 0.031128f
C17415 DVDD.n13854 VSS 0.031128f
C17416 DVDD.n13855 VSS 0.031128f
C17417 DVDD.n13856 VSS 0.031128f
C17418 DVDD.n13857 VSS 0.031128f
C17419 DVDD.n13858 VSS 0.031128f
C17420 DVDD.n13859 VSS 0.031128f
C17421 DVDD.n13860 VSS 0.031128f
C17422 DVDD.n13861 VSS 0.031128f
C17423 DVDD.n13862 VSS 0.031128f
C17424 DVDD.n13863 VSS 0.031128f
C17425 DVDD.n13864 VSS 0.031128f
C17426 DVDD.n13865 VSS 0.031128f
C17427 DVDD.n13866 VSS 0.031128f
C17428 DVDD.n13867 VSS 0.031128f
C17429 DVDD.n13868 VSS 0.031128f
C17430 DVDD.n13869 VSS 0.031128f
C17431 DVDD.n13870 VSS 0.031128f
C17432 DVDD.n13871 VSS 0.031128f
C17433 DVDD.n13872 VSS 0.031128f
C17434 DVDD.n13873 VSS 0.031128f
C17435 DVDD.n13874 VSS 0.031128f
C17436 DVDD.n13875 VSS 0.031128f
C17437 DVDD.n13876 VSS 0.031128f
C17438 DVDD.n13877 VSS 0.031128f
C17439 DVDD.n13878 VSS 0.031128f
C17440 DVDD.n13879 VSS 0.031128f
C17441 DVDD.n13880 VSS 0.031128f
C17442 DVDD.n13881 VSS 0.031128f
C17443 DVDD.n13882 VSS 0.031128f
C17444 DVDD.n13883 VSS 0.031128f
C17445 DVDD.n13884 VSS 0.031128f
C17446 DVDD.n13885 VSS 0.031128f
C17447 DVDD.n13886 VSS 0.031128f
C17448 DVDD.n13887 VSS 0.031128f
C17449 DVDD.n13888 VSS 0.031128f
C17450 DVDD.n13889 VSS 0.031128f
C17451 DVDD.n13890 VSS 0.031128f
C17452 DVDD.n13891 VSS 0.031128f
C17453 DVDD.n13892 VSS 0.031128f
C17454 DVDD.n13893 VSS 0.031128f
C17455 DVDD.n13894 VSS 0.031128f
C17456 DVDD.n13895 VSS 0.031128f
C17457 DVDD.n13896 VSS 0.031128f
C17458 DVDD.n13897 VSS 0.031128f
C17459 DVDD.n13898 VSS 0.031128f
C17460 DVDD.n13899 VSS 0.031128f
C17461 DVDD.n13900 VSS 0.031128f
C17462 DVDD.n13901 VSS 0.031128f
C17463 DVDD.n13902 VSS 0.031128f
C17464 DVDD.n13903 VSS 0.031128f
C17465 DVDD.n13904 VSS 0.031128f
C17466 DVDD.n13905 VSS 0.031128f
C17467 DVDD.n13906 VSS 0.031128f
C17468 DVDD.n13907 VSS 0.031128f
C17469 DVDD.n13908 VSS 0.031128f
C17470 DVDD.n13909 VSS 0.031128f
C17471 DVDD.n13910 VSS 0.031128f
C17472 DVDD.n13911 VSS 0.031128f
C17473 DVDD.n13912 VSS 0.031128f
C17474 DVDD.n13913 VSS 0.031128f
C17475 DVDD.n13914 VSS 0.031128f
C17476 DVDD.n13915 VSS 0.031128f
C17477 DVDD.n13916 VSS 0.031128f
C17478 DVDD.n13917 VSS 0.031128f
C17479 DVDD.n13918 VSS 0.031128f
C17480 DVDD.n13919 VSS 0.031128f
C17481 DVDD.n13920 VSS 0.031128f
C17482 DVDD.n13921 VSS 0.031128f
C17483 DVDD.n13922 VSS 0.031128f
C17484 DVDD.n13923 VSS 0.031128f
C17485 DVDD.n13924 VSS 0.031128f
C17486 DVDD.n13925 VSS 0.031128f
C17487 DVDD.n13926 VSS 0.031128f
C17488 DVDD.n13927 VSS 0.031128f
C17489 DVDD.n13928 VSS 0.031128f
C17490 DVDD.n13929 VSS 0.031128f
C17491 DVDD.n13930 VSS 0.031128f
C17492 DVDD.n13931 VSS 0.031128f
C17493 DVDD.n13932 VSS 0.031128f
C17494 DVDD.n13933 VSS 0.031128f
C17495 DVDD.n13934 VSS 0.031128f
C17496 DVDD.n13935 VSS 0.031128f
C17497 DVDD.n13936 VSS 0.031128f
C17498 DVDD.n13937 VSS 0.031128f
C17499 DVDD.n13938 VSS 0.031128f
C17500 DVDD.n13939 VSS 0.031128f
C17501 DVDD.n13940 VSS 0.031128f
C17502 DVDD.n13941 VSS 0.031128f
C17503 DVDD.n13942 VSS 0.031128f
C17504 DVDD.n13943 VSS 0.031128f
C17505 DVDD.n13944 VSS 0.031128f
C17506 DVDD.n13945 VSS 0.031128f
C17507 DVDD.n13946 VSS 0.031128f
C17508 DVDD.n13947 VSS 0.031128f
C17509 DVDD.n13948 VSS 0.031128f
C17510 DVDD.n13949 VSS 0.031128f
C17511 DVDD.n13950 VSS 0.031128f
C17512 DVDD.n13951 VSS 0.031128f
C17513 DVDD.n13952 VSS 0.031128f
C17514 DVDD.n13953 VSS 0.031128f
C17515 DVDD.n13954 VSS 0.031128f
C17516 DVDD.n13955 VSS 0.031128f
C17517 DVDD.n13956 VSS 0.031128f
C17518 DVDD.n13957 VSS 0.031128f
C17519 DVDD.n13958 VSS 0.031128f
C17520 DVDD.n13959 VSS 0.031128f
C17521 DVDD.n13960 VSS 0.031128f
C17522 DVDD.n13961 VSS 0.031128f
C17523 DVDD.n13962 VSS 0.031128f
C17524 DVDD.n13963 VSS 0.031128f
C17525 DVDD.n13964 VSS 0.031128f
C17526 DVDD.n13965 VSS 0.031128f
C17527 DVDD.n13966 VSS 0.031128f
C17528 DVDD.n13967 VSS 0.031128f
C17529 DVDD.n13968 VSS 0.031128f
C17530 DVDD.n13969 VSS 0.031128f
C17531 DVDD.n13970 VSS 0.031128f
C17532 DVDD.n13971 VSS 0.031128f
C17533 DVDD.n13972 VSS 0.031128f
C17534 DVDD.n13973 VSS 0.031128f
C17535 DVDD.n13974 VSS 0.031128f
C17536 DVDD.n13975 VSS 0.031128f
C17537 DVDD.n13976 VSS 0.031128f
C17538 DVDD.n13977 VSS 0.031128f
C17539 DVDD.n13978 VSS 0.031128f
C17540 DVDD.n13979 VSS 0.031128f
C17541 DVDD.n13980 VSS 0.031128f
C17542 DVDD.n13981 VSS 0.031128f
C17543 DVDD.n13982 VSS 0.031128f
C17544 DVDD.n13983 VSS 0.031128f
C17545 DVDD.n13984 VSS 0.031128f
C17546 DVDD.n13985 VSS 0.031128f
C17547 DVDD.n13986 VSS 0.031128f
C17548 DVDD.n13987 VSS 0.031128f
C17549 DVDD.n13988 VSS 0.031128f
C17550 DVDD.n13989 VSS 0.031128f
C17551 DVDD.n13990 VSS 0.031128f
C17552 DVDD.n13991 VSS 0.031128f
C17553 DVDD.n13992 VSS 0.031128f
C17554 DVDD.n13993 VSS 0.031128f
C17555 DVDD.n13994 VSS 0.031128f
C17556 DVDD.n13995 VSS 0.031128f
C17557 DVDD.n13996 VSS 0.031128f
C17558 DVDD.n13997 VSS 0.026086f
C17559 DVDD.n13998 VSS 0.019729f
C17560 DVDD.n13999 VSS 0.019729f
C17561 DVDD.n14000 VSS 0.522252f
C17562 DVDD.n14001 VSS 0.019729f
C17563 DVDD.n14003 VSS 0.105293f
C17564 DVDD.n14004 VSS 0.484347f
C17565 DVDD.n14005 VSS 0.033515f
C17566 DVDD.n14006 VSS 0.033515f
C17567 DVDD.n14007 VSS 0.029271f
C17568 DVDD.n14008 VSS 0.036621f
C17569 DVDD.n14009 VSS 0.022308f
C17570 DVDD.n14010 VSS 0.025542f
C17571 DVDD.n14011 VSS 0.025542f
C17572 DVDD.n14012 VSS 0.429595f
C17573 DVDD.n14013 VSS 0.433807f
C17574 DVDD.n14014 VSS 0.037465f
C17575 DVDD.n14015 VSS 0.037465f
C17576 DVDD.n14016 VSS 0.033442f
C17577 DVDD.n14017 VSS 0.053165f
C17578 DVDD.n14018 VSS 0.052307f
C17579 DVDD.n14019 VSS 0.0586f
C17580 DVDD.n14020 VSS 0.033945f
C17581 DVDD.n14021 VSS 0.019729f
C17582 DVDD.n14022 VSS 0.028497f
C17583 DVDD.n14023 VSS 0.031128f
C17584 DVDD.n14024 VSS 0.031128f
C17585 DVDD.n14025 VSS 0.031128f
C17586 DVDD.n14026 VSS 0.031128f
C17587 DVDD.n14028 VSS 0.031128f
C17588 DVDD.n14029 VSS 0.031128f
C17589 DVDD.n14030 VSS 0.031128f
C17590 DVDD.n14032 VSS 0.031128f
C17591 DVDD.n14033 VSS 0.031128f
C17592 DVDD.n14034 VSS 0.031128f
C17593 DVDD.n14035 VSS 0.031128f
C17594 DVDD.n14036 VSS 0.031128f
C17595 DVDD.n14037 VSS 0.031128f
C17596 DVDD.n14038 VSS 0.031128f
C17597 DVDD.n14040 VSS 0.031128f
C17598 DVDD.n14041 VSS 0.031128f
C17599 DVDD.n14042 VSS 0.031128f
C17600 DVDD.n14044 VSS 0.031128f
C17601 DVDD.n14045 VSS 0.031128f
C17602 DVDD.n14046 VSS 0.031128f
C17603 DVDD.n14047 VSS 0.031128f
C17604 DVDD.n14048 VSS 0.031128f
C17605 DVDD.n14049 VSS 0.031128f
C17606 DVDD.n14050 VSS 0.031128f
C17607 DVDD.n14052 VSS 0.031128f
C17608 DVDD.n14053 VSS 0.031128f
C17609 DVDD.n14054 VSS 0.031128f
C17610 DVDD.n14056 VSS 0.031128f
C17611 DVDD.n14057 VSS 0.031128f
C17612 DVDD.n14058 VSS 0.031128f
C17613 DVDD.n14059 VSS 0.031128f
C17614 DVDD.n14060 VSS 0.031128f
C17615 DVDD.n14061 VSS 0.031128f
C17616 DVDD.n14062 VSS 0.031128f
C17617 DVDD.n14064 VSS 0.031128f
C17618 DVDD.n14065 VSS 0.031128f
C17619 DVDD.n14066 VSS 0.031128f
C17620 DVDD.n14068 VSS 0.031128f
C17621 DVDD.n14069 VSS 0.031128f
C17622 DVDD.n14070 VSS 0.031128f
C17623 DVDD.n14071 VSS 0.031128f
C17624 DVDD.n14072 VSS 0.031128f
C17625 DVDD.n14073 VSS 0.031128f
C17626 DVDD.n14074 VSS 0.031128f
C17627 DVDD.n14076 VSS 0.031128f
C17628 DVDD.n14077 VSS 0.031128f
C17629 DVDD.n14078 VSS 0.031128f
C17630 DVDD.n14080 VSS 0.031128f
C17631 DVDD.n14081 VSS 0.031128f
C17632 DVDD.n14082 VSS 0.031128f
C17633 DVDD.n14083 VSS 0.031128f
C17634 DVDD.n14084 VSS 0.031128f
C17635 DVDD.n14085 VSS 0.031128f
C17636 DVDD.n14086 VSS 0.031128f
C17637 DVDD.n14088 VSS 0.031128f
C17638 DVDD.n14089 VSS 0.031128f
C17639 DVDD.n14090 VSS 0.031128f
C17640 DVDD.n14092 VSS 0.031128f
C17641 DVDD.n14093 VSS 0.031128f
C17642 DVDD.n14094 VSS 0.031128f
C17643 DVDD.n14095 VSS 0.031128f
C17644 DVDD.n14096 VSS 0.031128f
C17645 DVDD.n14097 VSS 0.031128f
C17646 DVDD.n14098 VSS 0.031128f
C17647 DVDD.n14100 VSS 0.031128f
C17648 DVDD.n14101 VSS 0.031128f
C17649 DVDD.n14102 VSS 0.031128f
C17650 DVDD.n14104 VSS 0.031128f
C17651 DVDD.n14105 VSS 0.031128f
C17652 DVDD.n14106 VSS 0.031128f
C17653 DVDD.n14107 VSS 0.031128f
C17654 DVDD.n14108 VSS 0.031128f
C17655 DVDD.n14109 VSS 0.031128f
C17656 DVDD.n14110 VSS 0.031128f
C17657 DVDD.n14112 VSS 0.031128f
C17658 DVDD.n14113 VSS 0.031128f
C17659 DVDD.n14114 VSS 0.031128f
C17660 DVDD.n14116 VSS 0.031128f
C17661 DVDD.n14117 VSS 0.031128f
C17662 DVDD.n14118 VSS 0.031128f
C17663 DVDD.n14119 VSS 0.031128f
C17664 DVDD.n14120 VSS 0.031128f
C17665 DVDD.n14121 VSS 0.031128f
C17666 DVDD.n14122 VSS 0.031128f
C17667 DVDD.n14124 VSS 0.031128f
C17668 DVDD.n14125 VSS 0.031128f
C17669 DVDD.n14126 VSS 0.031128f
C17670 DVDD.n14128 VSS 0.031128f
C17671 DVDD.n14129 VSS 0.031128f
C17672 DVDD.n14130 VSS 0.031128f
C17673 DVDD.n14131 VSS 0.031128f
C17674 DVDD.n14132 VSS 0.031128f
C17675 DVDD.n14133 VSS 0.031128f
C17676 DVDD.n14134 VSS 0.031128f
C17677 DVDD.n14136 VSS 0.031128f
C17678 DVDD.n14137 VSS 0.031128f
C17679 DVDD.n14138 VSS 0.031128f
C17680 DVDD.n14140 VSS 0.031128f
C17681 DVDD.n14141 VSS 0.031128f
C17682 DVDD.n14142 VSS 0.031128f
C17683 DVDD.n14143 VSS 0.031128f
C17684 DVDD.n14144 VSS 0.031128f
C17685 DVDD.n14145 VSS 0.031128f
C17686 DVDD.n14146 VSS 0.031128f
C17687 DVDD.n14148 VSS 0.031128f
C17688 DVDD.n14149 VSS 0.031128f
C17689 DVDD.n14150 VSS 0.031128f
C17690 DVDD.n14152 VSS 0.031128f
C17691 DVDD.n14153 VSS 0.031128f
C17692 DVDD.n14154 VSS 0.031128f
C17693 DVDD.n14155 VSS 0.031128f
C17694 DVDD.n14156 VSS 0.031128f
C17695 DVDD.n14157 VSS 0.031128f
C17696 DVDD.n14158 VSS 0.031128f
C17697 DVDD.n14160 VSS 0.031128f
C17698 DVDD.n14161 VSS 0.031128f
C17699 DVDD.n14162 VSS 0.031128f
C17700 DVDD.n14164 VSS 0.031128f
C17701 DVDD.n14165 VSS 0.031128f
C17702 DVDD.n14166 VSS 0.031128f
C17703 DVDD.n14167 VSS 0.031128f
C17704 DVDD.n14168 VSS 0.031128f
C17705 DVDD.n14169 VSS 0.031128f
C17706 DVDD.n14170 VSS 0.031128f
C17707 DVDD.n14172 VSS 0.031128f
C17708 DVDD.n14173 VSS 0.031128f
C17709 DVDD.n14174 VSS 0.031128f
C17710 DVDD.n14176 VSS 0.031128f
C17711 DVDD.n14177 VSS 0.031128f
C17712 DVDD.n14178 VSS 0.031128f
C17713 DVDD.n14179 VSS 0.031128f
C17714 DVDD.n14180 VSS 0.031128f
C17715 DVDD.n14181 VSS 0.031128f
C17716 DVDD.n14182 VSS 0.031128f
C17717 DVDD.n14184 VSS 0.031128f
C17718 DVDD.n14185 VSS 0.031128f
C17719 DVDD.n14186 VSS 0.031128f
C17720 DVDD.n14188 VSS 0.031128f
C17721 DVDD.n14189 VSS 0.031128f
C17722 DVDD.n14190 VSS 0.031128f
C17723 DVDD.n14191 VSS 0.031128f
C17724 DVDD.n14192 VSS 0.031128f
C17725 DVDD.n14193 VSS 0.031128f
C17726 DVDD.n14194 VSS 0.031128f
C17727 DVDD.n14196 VSS 0.031128f
C17728 DVDD.n14197 VSS 0.031128f
C17729 DVDD.n14198 VSS 0.031128f
C17730 DVDD.n14200 VSS 0.031128f
C17731 DVDD.n14201 VSS 0.031128f
C17732 DVDD.n14202 VSS 0.031128f
C17733 DVDD.n14203 VSS 0.031128f
C17734 DVDD.n14204 VSS 0.031128f
C17735 DVDD.n14205 VSS 0.031128f
C17736 DVDD.n14206 VSS 0.031128f
C17737 DVDD.n14208 VSS 0.031128f
C17738 DVDD.n14209 VSS 0.031128f
C17739 DVDD.n14210 VSS 0.031128f
C17740 DVDD.n14212 VSS 0.031128f
C17741 DVDD.n14213 VSS 0.031128f
C17742 DVDD.n14214 VSS 0.031128f
C17743 DVDD.n14215 VSS 0.031128f
C17744 DVDD.n14216 VSS 0.031128f
C17745 DVDD.n14217 VSS 0.031128f
C17746 DVDD.n14218 VSS 0.031128f
C17747 DVDD.n14220 VSS 0.031128f
C17748 DVDD.n14221 VSS 0.031128f
C17749 DVDD.n14222 VSS 0.031128f
C17750 DVDD.n14224 VSS 0.031128f
C17751 DVDD.n14225 VSS 0.031128f
C17752 DVDD.n14226 VSS 0.031128f
C17753 DVDD.n14227 VSS 0.031128f
C17754 DVDD.n14228 VSS 0.031128f
C17755 DVDD.n14229 VSS 0.031128f
C17756 DVDD.n14230 VSS 0.031128f
C17757 DVDD.n14232 VSS 0.031128f
C17758 DVDD.n14233 VSS 0.031128f
C17759 DVDD.n14234 VSS 0.031128f
C17760 DVDD.n14236 VSS 0.031128f
C17761 DVDD.n14237 VSS 0.031128f
C17762 DVDD.n14238 VSS 0.031128f
C17763 DVDD.n14239 VSS 0.031128f
C17764 DVDD.n14240 VSS 0.031128f
C17765 DVDD.n14241 VSS 0.031128f
C17766 DVDD.n14242 VSS 0.031128f
C17767 DVDD.n14244 VSS 0.031128f
C17768 DVDD.n14245 VSS 0.031128f
C17769 DVDD.n14246 VSS 0.031128f
C17770 DVDD.n14248 VSS 0.031128f
C17771 DVDD.n14249 VSS 0.031128f
C17772 DVDD.n14250 VSS 0.031128f
C17773 DVDD.n14251 VSS 0.031128f
C17774 DVDD.n14252 VSS 0.031128f
C17775 DVDD.n14253 VSS 0.031128f
C17776 DVDD.n14254 VSS 0.031128f
C17777 DVDD.n14256 VSS 0.031128f
C17778 DVDD.n14257 VSS 0.031128f
C17779 DVDD.n14258 VSS 0.031128f
C17780 DVDD.n14260 VSS 0.031128f
C17781 DVDD.n14261 VSS 0.031128f
C17782 DVDD.n14262 VSS 0.031128f
C17783 DVDD.n14263 VSS 0.031128f
C17784 DVDD.n14264 VSS 0.031128f
C17785 DVDD.n14265 VSS 0.031128f
C17786 DVDD.n14266 VSS 0.031128f
C17787 DVDD.n14268 VSS 0.019729f
C17788 DVDD.n14269 VSS 0.484347f
C17789 DVDD.n14270 VSS 0.303243f
C17790 DVDD.n14271 VSS 0.021704f
C17791 DVDD.n14272 VSS 0.021704f
C17792 DVDD.n14273 VSS 0.018955f
C17793 DVDD.n14274 VSS 0.028833f
C17794 DVDD.n14275 VSS 0.035976f
C17795 DVDD.n14276 VSS 0.033913f
C17796 DVDD.n14277 VSS 0.03883f
C17797 DVDD.n14278 VSS 0.02513f
C17798 DVDD.n14279 VSS 0.019729f
C17799 DVDD.n14280 VSS 0.019729f
C17800 DVDD.n14281 VSS 0.408536f
C17801 DVDD.n14282 VSS 0.019729f
C17802 DVDD.n14284 VSS 0.332725f
C17803 DVDD.n14285 VSS 0.362207f
C17804 DVDD.n14286 VSS 0.053796f
C17805 DVDD.n14287 VSS 0.053796f
C17806 DVDD.n14288 VSS 0.04802f
C17807 DVDD.n14289 VSS 0.053165f
C17808 DVDD.n14290 VSS 0.03773f
C17809 DVDD.n14291 VSS 0.042269f
C17810 DVDD.n14292 VSS 0.042269f
C17811 DVDD.n14293 VSS 0.496982f
C17812 DVDD.n14294 VSS 0.518041f
C17813 DVDD.n14295 VSS 0.027905f
C17814 DVDD.n14296 VSS 0.027905f
C17815 DVDD.n14297 VSS 0.024371f
C17816 DVDD.n14298 VSS 0.036621f
C17817 DVDD.n14299 VSS 0.027208f
C17818 DVDD.n14300 VSS 0.031153f
C17819 DVDD.n14301 VSS 0.031153f
C17820 DVDD.n14302 VSS 0.480135f
C17821 DVDD.n14303 VSS 0.593852f
C17822 DVDD.n14304 VSS 0.040347f
C17823 DVDD.n14305 VSS 0.040347f
C17824 DVDD.n14306 VSS 0.036015f
C17825 DVDD.n14307 VSS 0.053165f
C17826 DVDD.n14308 VSS 0.049735f
C17827 DVDD.n14309 VSS 0.055718f
C17828 DVDD.n14310 VSS 0.033945f
C17829 DVDD.n14311 VSS 0.019729f
C17830 DVDD.n14312 VSS 0.028497f
C17831 DVDD.n14313 VSS 0.031128f
C17832 DVDD.n14314 VSS 0.031128f
C17833 DVDD.n14315 VSS 0.031128f
C17834 DVDD.n14316 VSS 0.031128f
C17835 DVDD.n14318 VSS 0.031128f
C17836 DVDD.n14319 VSS 0.031128f
C17837 DVDD.n14320 VSS 0.031128f
C17838 DVDD.n14322 VSS 0.031128f
C17839 DVDD.n14323 VSS 0.031128f
C17840 DVDD.n14324 VSS 0.031128f
C17841 DVDD.n14325 VSS 0.031128f
C17842 DVDD.n14326 VSS 0.031128f
C17843 DVDD.n14327 VSS 0.031128f
C17844 DVDD.n14328 VSS 0.031128f
C17845 DVDD.n14330 VSS 0.031128f
C17846 DVDD.n14331 VSS 0.031128f
C17847 DVDD.n14332 VSS 0.031128f
C17848 DVDD.n14334 VSS 0.031128f
C17849 DVDD.n14335 VSS 0.031128f
C17850 DVDD.n14336 VSS 0.031128f
C17851 DVDD.n14337 VSS 0.031128f
C17852 DVDD.n14338 VSS 0.031128f
C17853 DVDD.n14339 VSS 0.031128f
C17854 DVDD.n14340 VSS 0.031128f
C17855 DVDD.n14342 VSS 0.031128f
C17856 DVDD.n14343 VSS 0.031128f
C17857 DVDD.n14344 VSS 0.031128f
C17858 DVDD.n14346 VSS 0.031128f
C17859 DVDD.n14347 VSS 0.031128f
C17860 DVDD.n14348 VSS 0.031128f
C17861 DVDD.n14349 VSS 0.031128f
C17862 DVDD.n14350 VSS 0.031128f
C17863 DVDD.n14351 VSS 0.031128f
C17864 DVDD.n14352 VSS 0.031128f
C17865 DVDD.n14354 VSS 0.031128f
C17866 DVDD.n14355 VSS 0.031128f
C17867 DVDD.n14356 VSS 0.031128f
C17868 DVDD.n14358 VSS 0.031128f
C17869 DVDD.n14359 VSS 0.031128f
C17870 DVDD.n14360 VSS 0.031128f
C17871 DVDD.n14361 VSS 0.031128f
C17872 DVDD.n14362 VSS 0.031128f
C17873 DVDD.n14363 VSS 0.031128f
C17874 DVDD.n14364 VSS 0.031128f
C17875 DVDD.n14366 VSS 0.031128f
C17876 DVDD.n14367 VSS 0.031128f
C17877 DVDD.n14368 VSS 0.031128f
C17878 DVDD.n14370 VSS 0.031128f
C17879 DVDD.n14371 VSS 0.031128f
C17880 DVDD.n14372 VSS 0.031128f
C17881 DVDD.n14373 VSS 0.031128f
C17882 DVDD.n14374 VSS 0.031128f
C17883 DVDD.n14375 VSS 0.031128f
C17884 DVDD.n14376 VSS 0.031128f
C17885 DVDD.n14378 VSS 0.031128f
C17886 DVDD.n14379 VSS 0.031128f
C17887 DVDD.n14380 VSS 0.031128f
C17888 DVDD.n14382 VSS 0.031128f
C17889 DVDD.n14383 VSS 0.031128f
C17890 DVDD.n14384 VSS 0.031128f
C17891 DVDD.n14385 VSS 0.031128f
C17892 DVDD.n14386 VSS 0.031128f
C17893 DVDD.n14387 VSS 0.031128f
C17894 DVDD.n14388 VSS 0.031128f
C17895 DVDD.n14390 VSS 0.031128f
C17896 DVDD.n14391 VSS 0.031128f
C17897 DVDD.n14392 VSS 0.031128f
C17898 DVDD.n14394 VSS 0.031128f
C17899 DVDD.n14395 VSS 0.031128f
C17900 DVDD.n14396 VSS 0.031128f
C17901 DVDD.n14397 VSS 0.031128f
C17902 DVDD.n14398 VSS 0.031128f
C17903 DVDD.n14399 VSS 0.031128f
C17904 DVDD.n14400 VSS 0.031128f
C17905 DVDD.n14402 VSS 0.031128f
C17906 DVDD.n14403 VSS 0.031128f
C17907 DVDD.n14404 VSS 0.031128f
C17908 DVDD.n14406 VSS 0.031128f
C17909 DVDD.n14407 VSS 0.031128f
C17910 DVDD.n14408 VSS 0.031128f
C17911 DVDD.n14409 VSS 0.031128f
C17912 DVDD.n14410 VSS 0.031128f
C17913 DVDD.n14411 VSS 0.031128f
C17914 DVDD.n14412 VSS 0.031128f
C17915 DVDD.n14414 VSS 0.031128f
C17916 DVDD.n14415 VSS 0.031128f
C17917 DVDD.n14416 VSS 0.031128f
C17918 DVDD.n14418 VSS 0.031128f
C17919 DVDD.n14419 VSS 0.031128f
C17920 DVDD.n14420 VSS 0.031128f
C17921 DVDD.n14421 VSS 0.031128f
C17922 DVDD.n14422 VSS 0.031128f
C17923 DVDD.n14423 VSS 0.031128f
C17924 DVDD.n14424 VSS 0.031128f
C17925 DVDD.n14426 VSS 0.031128f
C17926 DVDD.n14427 VSS 0.031128f
C17927 DVDD.n14428 VSS 0.031128f
C17928 DVDD.n14430 VSS 0.031128f
C17929 DVDD.n14431 VSS 0.031128f
C17930 DVDD.n14432 VSS 0.031128f
C17931 DVDD.n14433 VSS 0.031128f
C17932 DVDD.n14434 VSS 0.031128f
C17933 DVDD.n14435 VSS 0.031128f
C17934 DVDD.n14436 VSS 0.031128f
C17935 DVDD.n14438 VSS 0.031128f
C17936 DVDD.n14439 VSS 0.031128f
C17937 DVDD.n14440 VSS 0.031128f
C17938 DVDD.n14442 VSS 0.031128f
C17939 DVDD.n14443 VSS 0.031128f
C17940 DVDD.n14444 VSS 0.031128f
C17941 DVDD.n14445 VSS 0.031128f
C17942 DVDD.n14446 VSS 0.031128f
C17943 DVDD.n14447 VSS 0.031128f
C17944 DVDD.n14448 VSS 0.031128f
C17945 DVDD.n14450 VSS 0.031128f
C17946 DVDD.n14451 VSS 0.031128f
C17947 DVDD.n14452 VSS 0.031128f
C17948 DVDD.n14454 VSS 0.031128f
C17949 DVDD.n14455 VSS 0.031128f
C17950 DVDD.n14456 VSS 0.031128f
C17951 DVDD.n14457 VSS 0.031128f
C17952 DVDD.n14458 VSS 0.031128f
C17953 DVDD.n14459 VSS 0.031128f
C17954 DVDD.n14460 VSS 0.031128f
C17955 DVDD.n14462 VSS 0.031128f
C17956 DVDD.n14463 VSS 0.031128f
C17957 DVDD.n14464 VSS 0.031128f
C17958 DVDD.n14466 VSS 0.031128f
C17959 DVDD.n14467 VSS 0.031128f
C17960 DVDD.n14468 VSS 0.031128f
C17961 DVDD.n14469 VSS 0.031128f
C17962 DVDD.n14470 VSS 0.031128f
C17963 DVDD.n14471 VSS 0.031128f
C17964 DVDD.n14472 VSS 0.031128f
C17965 DVDD.n14474 VSS 0.031128f
C17966 DVDD.n14475 VSS 0.031128f
C17967 DVDD.n14476 VSS 0.031128f
C17968 DVDD.n14478 VSS 0.031128f
C17969 DVDD.n14479 VSS 0.031128f
C17970 DVDD.n14480 VSS 0.031128f
C17971 DVDD.n14481 VSS 0.031128f
C17972 DVDD.n14482 VSS 0.031128f
C17973 DVDD.n14483 VSS 0.031128f
C17974 DVDD.n14484 VSS 0.031128f
C17975 DVDD.n14486 VSS 0.031128f
C17976 DVDD.n14487 VSS 0.031128f
C17977 DVDD.n14488 VSS 0.031128f
C17978 DVDD.n14490 VSS 0.031128f
C17979 DVDD.n14491 VSS 0.031128f
C17980 DVDD.n14492 VSS 0.031128f
C17981 DVDD.n14493 VSS 0.031128f
C17982 DVDD.n14494 VSS 0.031128f
C17983 DVDD.n14495 VSS 0.031128f
C17984 DVDD.n14496 VSS 0.031128f
C17985 DVDD.n14498 VSS 0.031128f
C17986 DVDD.n14499 VSS 0.031128f
C17987 DVDD.n14500 VSS 0.031128f
C17988 DVDD.n14502 VSS 0.031128f
C17989 DVDD.n14503 VSS 0.031128f
C17990 DVDD.n14504 VSS 0.031128f
C17991 DVDD.n14505 VSS 0.031128f
C17992 DVDD.n14506 VSS 0.031128f
C17993 DVDD.n14507 VSS 0.031128f
C17994 DVDD.n14508 VSS 0.031128f
C17995 DVDD.n14510 VSS 0.031128f
C17996 DVDD.n14511 VSS 0.031128f
C17997 DVDD.n14512 VSS 0.031128f
C17998 DVDD.n14514 VSS 0.031128f
C17999 DVDD.n14515 VSS 0.031128f
C18000 DVDD.n14516 VSS 0.031128f
C18001 DVDD.n14517 VSS 0.031128f
C18002 DVDD.n14518 VSS 0.031128f
C18003 DVDD.n14519 VSS 0.031128f
C18004 DVDD.n14520 VSS 0.031128f
C18005 DVDD.n14522 VSS 0.031128f
C18006 DVDD.n14523 VSS 0.031128f
C18007 DVDD.n14524 VSS 0.031128f
C18008 DVDD.n14526 VSS 0.031128f
C18009 DVDD.n14527 VSS 0.031128f
C18010 DVDD.n14528 VSS 0.031128f
C18011 DVDD.n14529 VSS 0.031128f
C18012 DVDD.n14530 VSS 0.031128f
C18013 DVDD.n14531 VSS 0.031128f
C18014 DVDD.n14532 VSS 0.031128f
C18015 DVDD.n14534 VSS 0.031128f
C18016 DVDD.n14535 VSS 0.031128f
C18017 DVDD.n14536 VSS 0.031128f
C18018 DVDD.n14538 VSS 0.031128f
C18019 DVDD.n14539 VSS 0.031128f
C18020 DVDD.n14540 VSS 0.031128f
C18021 DVDD.n14541 VSS 0.031128f
C18022 DVDD.n14542 VSS 0.031128f
C18023 DVDD.n14543 VSS 0.031128f
C18024 DVDD.n14544 VSS 0.031128f
C18025 DVDD.n14546 VSS 0.031128f
C18026 DVDD.n14547 VSS 0.031128f
C18027 DVDD.n14548 VSS 0.031128f
C18028 DVDD.n14550 VSS 0.031128f
C18029 DVDD.n14551 VSS 0.031128f
C18030 DVDD.n14552 VSS 0.031128f
C18031 DVDD.n14553 VSS 0.031128f
C18032 DVDD.n14554 VSS 0.031128f
C18033 DVDD.n14555 VSS 0.031128f
C18034 DVDD.n14556 VSS 0.031128f
C18035 DVDD.n14558 VSS 0.019729f
C18036 DVDD.n14559 VSS 0.273761f
C18037 DVDD.n14560 VSS 0.362207f
C18038 DVDD.n14561 VSS 0.027314f
C18039 DVDD.n14562 VSS 0.027314f
C18040 DVDD.n14563 VSS 0.023855f
C18041 DVDD.n14564 VSS 0.028833f
C18042 DVDD.n14565 VSS 0.031076f
C18043 DVDD.n14566 VSS 0.035582f
C18044 DVDD.n14567 VSS 0.035582f
C18045 DVDD.n14568 VSS 0.286396f
C18046 DVDD.n14569 VSS 0.598063f
C18047 DVDD.n14570 VSS 0.05956f
C18048 DVDD.n14571 VSS 0.05956f
C18049 DVDD.n14572 VSS 0.053165f
C18050 DVDD.n14573 VSS 0.053165f
C18051 DVDD.n14574 VSS 0.029155f
C18052 DVDD.n14575 VSS 0.032662f
C18053 DVDD.n14576 VSS 0.033945f
C18054 DVDD.n14577 VSS 0.019729f
C18055 DVDD.n14578 VSS 0.028497f
C18056 DVDD.n14579 VSS 0.031128f
C18057 DVDD.n14580 VSS 0.031128f
C18058 DVDD.n14581 VSS 0.031128f
C18059 DVDD.n14582 VSS 0.031128f
C18060 DVDD.n14584 VSS 0.031128f
C18061 DVDD.n14585 VSS 0.031128f
C18062 DVDD.n14586 VSS 0.031128f
C18063 DVDD.n14588 VSS 0.031128f
C18064 DVDD.n14589 VSS 0.031128f
C18065 DVDD.n14590 VSS 0.031128f
C18066 DVDD.n14591 VSS 0.031128f
C18067 DVDD.n14592 VSS 0.031128f
C18068 DVDD.n14593 VSS 0.031128f
C18069 DVDD.n14594 VSS 0.031128f
C18070 DVDD.n14596 VSS 0.031128f
C18071 DVDD.n14597 VSS 0.031128f
C18072 DVDD.n14598 VSS 0.031128f
C18073 DVDD.n14600 VSS 0.031128f
C18074 DVDD.n14601 VSS 0.031128f
C18075 DVDD.n14602 VSS 0.031128f
C18076 DVDD.n14603 VSS 0.031128f
C18077 DVDD.n14604 VSS 0.031128f
C18078 DVDD.n14605 VSS 0.031128f
C18079 DVDD.n14606 VSS 0.031128f
C18080 DVDD.n14608 VSS 0.031128f
C18081 DVDD.n14609 VSS 0.031128f
C18082 DVDD.n14610 VSS 0.031128f
C18083 DVDD.n14612 VSS 0.031128f
C18084 DVDD.n14613 VSS 0.031128f
C18085 DVDD.n14614 VSS 0.031128f
C18086 DVDD.n14615 VSS 0.031128f
C18087 DVDD.n14616 VSS 0.031128f
C18088 DVDD.n14617 VSS 0.031128f
C18089 DVDD.n14618 VSS 0.031128f
C18090 DVDD.n14620 VSS 0.031128f
C18091 DVDD.n14621 VSS 0.031128f
C18092 DVDD.n14622 VSS 0.031128f
C18093 DVDD.n14624 VSS 0.031128f
C18094 DVDD.n14625 VSS 0.031128f
C18095 DVDD.n14626 VSS 0.031128f
C18096 DVDD.n14627 VSS 0.031128f
C18097 DVDD.n14628 VSS 0.031128f
C18098 DVDD.n14629 VSS 0.031128f
C18099 DVDD.n14630 VSS 0.031128f
C18100 DVDD.n14632 VSS 0.031128f
C18101 DVDD.n14633 VSS 0.031128f
C18102 DVDD.n14634 VSS 0.031128f
C18103 DVDD.n14636 VSS 0.031128f
C18104 DVDD.n14637 VSS 0.031128f
C18105 DVDD.n14638 VSS 0.031128f
C18106 DVDD.n14639 VSS 0.031128f
C18107 DVDD.n14640 VSS 0.031128f
C18108 DVDD.n14641 VSS 0.031128f
C18109 DVDD.n14642 VSS 0.031128f
C18110 DVDD.n14644 VSS 0.031128f
C18111 DVDD.n14645 VSS 0.031128f
C18112 DVDD.n14646 VSS 0.031128f
C18113 DVDD.n14648 VSS 0.031128f
C18114 DVDD.n14649 VSS 0.031128f
C18115 DVDD.n14650 VSS 0.031128f
C18116 DVDD.n14651 VSS 0.031128f
C18117 DVDD.n14652 VSS 0.031128f
C18118 DVDD.n14653 VSS 0.031128f
C18119 DVDD.n14654 VSS 0.031128f
C18120 DVDD.n14656 VSS 0.031128f
C18121 DVDD.n14657 VSS 0.031128f
C18122 DVDD.n14658 VSS 0.031128f
C18123 DVDD.n14660 VSS 0.031128f
C18124 DVDD.n14661 VSS 0.031128f
C18125 DVDD.n14662 VSS 0.031128f
C18126 DVDD.n14663 VSS 0.031128f
C18127 DVDD.n14664 VSS 0.031128f
C18128 DVDD.n14665 VSS 0.031128f
C18129 DVDD.n14666 VSS 0.031128f
C18130 DVDD.n14668 VSS 0.031128f
C18131 DVDD.n14669 VSS 0.031128f
C18132 DVDD.n14670 VSS 0.031128f
C18133 DVDD.n14672 VSS 0.031128f
C18134 DVDD.n14673 VSS 0.031128f
C18135 DVDD.n14674 VSS 0.031128f
C18136 DVDD.n14675 VSS 0.031128f
C18137 DVDD.n14676 VSS 0.031128f
C18138 DVDD.n14677 VSS 0.031128f
C18139 DVDD.n14678 VSS 0.031128f
C18140 DVDD.n14680 VSS 0.031128f
C18141 DVDD.n14681 VSS 0.031128f
C18142 DVDD.n14682 VSS 0.031128f
C18143 DVDD.n14684 VSS 0.031128f
C18144 DVDD.n14685 VSS 0.031128f
C18145 DVDD.n14686 VSS 0.031128f
C18146 DVDD.n14687 VSS 0.031128f
C18147 DVDD.n14688 VSS 0.031128f
C18148 DVDD.n14689 VSS 0.031128f
C18149 DVDD.n14690 VSS 0.031128f
C18150 DVDD.n14692 VSS 0.031128f
C18151 DVDD.n14693 VSS 0.031128f
C18152 DVDD.n14694 VSS 0.031128f
C18153 DVDD.n14696 VSS 0.031128f
C18154 DVDD.n14697 VSS 0.031128f
C18155 DVDD.n14698 VSS 0.031128f
C18156 DVDD.n14699 VSS 0.031128f
C18157 DVDD.n14700 VSS 0.031128f
C18158 DVDD.n14701 VSS 0.031128f
C18159 DVDD.n14702 VSS 0.031128f
C18160 DVDD.n14704 VSS 0.031128f
C18161 DVDD.n14705 VSS 0.031128f
C18162 DVDD.n14706 VSS 0.031128f
C18163 DVDD.n14708 VSS 0.031128f
C18164 DVDD.n14709 VSS 0.031128f
C18165 DVDD.n14710 VSS 0.031128f
C18166 DVDD.n14711 VSS 0.031128f
C18167 DVDD.n14712 VSS 0.031128f
C18168 DVDD.n14713 VSS 0.031128f
C18169 DVDD.n14714 VSS 0.031128f
C18170 DVDD.n14716 VSS 0.031128f
C18171 DVDD.n14717 VSS 0.031128f
C18172 DVDD.n14718 VSS 0.031128f
C18173 DVDD.n14720 VSS 0.031128f
C18174 DVDD.n14721 VSS 0.031128f
C18175 DVDD.n14722 VSS 0.031128f
C18176 DVDD.n14723 VSS 0.031128f
C18177 DVDD.n14724 VSS 0.031128f
C18178 DVDD.n14725 VSS 0.031128f
C18179 DVDD.n14726 VSS 0.031128f
C18180 DVDD.n14728 VSS 0.031128f
C18181 DVDD.n14729 VSS 0.031128f
C18182 DVDD.n14730 VSS 0.031128f
C18183 DVDD.n14732 VSS 0.031128f
C18184 DVDD.n14733 VSS 0.031128f
C18185 DVDD.n14734 VSS 0.031128f
C18186 DVDD.n14735 VSS 0.031128f
C18187 DVDD.n14736 VSS 0.031128f
C18188 DVDD.n14737 VSS 0.031128f
C18189 DVDD.n14738 VSS 0.031128f
C18190 DVDD.n14740 VSS 0.031128f
C18191 DVDD.n14741 VSS 0.031128f
C18192 DVDD.n14742 VSS 0.031128f
C18193 DVDD.n14744 VSS 0.031128f
C18194 DVDD.n14745 VSS 0.031128f
C18195 DVDD.n14746 VSS 0.031128f
C18196 DVDD.n14747 VSS 0.031128f
C18197 DVDD.n14748 VSS 0.031128f
C18198 DVDD.n14749 VSS 0.031128f
C18199 DVDD.n14750 VSS 0.031128f
C18200 DVDD.n14752 VSS 0.031128f
C18201 DVDD.n14753 VSS 0.031128f
C18202 DVDD.n14754 VSS 0.031128f
C18203 DVDD.n14756 VSS 0.031128f
C18204 DVDD.n14757 VSS 0.031128f
C18205 DVDD.n14758 VSS 0.031128f
C18206 DVDD.n14759 VSS 0.031128f
C18207 DVDD.n14760 VSS 0.031128f
C18208 DVDD.n14761 VSS 0.031128f
C18209 DVDD.n14762 VSS 0.031128f
C18210 DVDD.n14764 VSS 0.031128f
C18211 DVDD.n14765 VSS 0.031128f
C18212 DVDD.n14766 VSS 0.031128f
C18213 DVDD.n14768 VSS 0.031128f
C18214 DVDD.n14769 VSS 0.031128f
C18215 DVDD.n14770 VSS 0.031128f
C18216 DVDD.n14771 VSS 0.031128f
C18217 DVDD.n14772 VSS 0.031128f
C18218 DVDD.n14773 VSS 0.031128f
C18219 DVDD.n14774 VSS 0.031128f
C18220 DVDD.n14776 VSS 0.031128f
C18221 DVDD.n14777 VSS 0.031128f
C18222 DVDD.n14778 VSS 0.031128f
C18223 DVDD.n14780 VSS 0.031128f
C18224 DVDD.n14781 VSS 0.031128f
C18225 DVDD.n14782 VSS 0.031128f
C18226 DVDD.n14783 VSS 0.031128f
C18227 DVDD.n14784 VSS 0.031128f
C18228 DVDD.n14785 VSS 0.031128f
C18229 DVDD.n14786 VSS 0.031128f
C18230 DVDD.n14788 VSS 0.031128f
C18231 DVDD.n14789 VSS 0.031128f
C18232 DVDD.n14790 VSS 0.031128f
C18233 DVDD.n14792 VSS 0.031128f
C18234 DVDD.n14793 VSS 0.031128f
C18235 DVDD.n14794 VSS 0.031128f
C18236 DVDD.n14795 VSS 0.031128f
C18237 DVDD.n14796 VSS 0.031128f
C18238 DVDD.n14797 VSS 0.031128f
C18239 DVDD.n14798 VSS 0.031128f
C18240 DVDD.n14800 VSS 0.031128f
C18241 DVDD.n14801 VSS 0.031128f
C18242 DVDD.n14802 VSS 0.031128f
C18243 DVDD.n14804 VSS 0.031128f
C18244 DVDD.n14805 VSS 0.031128f
C18245 DVDD.n14806 VSS 0.031128f
C18246 DVDD.n14807 VSS 0.031128f
C18247 DVDD.n14808 VSS 0.031128f
C18248 DVDD.n14809 VSS 0.031128f
C18249 DVDD.n14810 VSS 0.031128f
C18250 DVDD.n14812 VSS 0.031128f
C18251 DVDD.n14813 VSS 0.031128f
C18252 DVDD.n14814 VSS 0.031128f
C18253 DVDD.n14816 VSS 0.031128f
C18254 DVDD.n14817 VSS 0.031128f
C18255 DVDD.n14818 VSS 0.031128f
C18256 DVDD.n14819 VSS 0.031128f
C18257 DVDD.n14820 VSS 0.031128f
C18258 DVDD.n14821 VSS 0.031128f
C18259 DVDD.n14822 VSS 0.031128f
C18260 DVDD.n14824 VSS 0.019729f
C18261 DVDD.n14825 VSS 0.501194f
C18262 DVDD.n14826 VSS 0.256914f
C18263 DVDD.n14827 VSS 0.023475f
C18264 DVDD.n14828 VSS 0.023475f
C18265 DVDD.n14829 VSS 0.020503f
C18266 DVDD.n14830 VSS 0.028833f
C18267 DVDD.n14831 VSS 0.034429f
C18268 DVDD.n14832 VSS 0.03546f
C18269 DVDD.n14833 VSS 0.040602f
C18270 DVDD.n14834 VSS 0.02513f
C18271 DVDD.n14835 VSS 0.019729f
C18272 DVDD.n14836 VSS 0.019729f
C18273 DVDD.n14837 VSS 0.391689f
C18274 DVDD.n14838 VSS 0.019729f
C18275 DVDD.n14840 VSS 0.315878f
C18276 DVDD.n14841 VSS 0.357996f
C18277 DVDD.n14842 VSS 0.049954f
C18278 DVDD.n14843 VSS 0.049954f
C18279 DVDD.n14844 VSS 0.04459f
C18280 DVDD.n14845 VSS 0.053165f
C18281 DVDD.n14846 VSS 0.04116f
C18282 DVDD.n14847 VSS 0.046111f
C18283 DVDD.n14848 VSS 0.046111f
C18284 DVDD.n14849 VSS 0.450653f
C18285 DVDD.n14850 VSS 0.522252f
C18286 DVDD.n14851 VSS 0.026133f
C18287 DVDD.n14852 VSS 0.026133f
C18288 DVDD.n14853 VSS 0.022823f
C18289 DVDD.n14854 VSS 0.036621f
C18290 DVDD.n14855 VSS 0.028755f
C18291 DVDD.n14856 VSS 0.032925f
C18292 DVDD.n14857 VSS 0.02513f
C18293 DVDD.n14858 VSS 0.019729f
C18294 DVDD.n14859 VSS 0.019729f
C18295 DVDD.n14860 VSS 0.459077f
C18296 DVDD.n14861 VSS 0.019729f
C18297 DVDD.n14863 VSS 0.383266f
C18298 DVDD.n14864 VSS 0.577005f
C18299 DVDD.n14865 VSS 0.05956f
C18300 DVDD.n14866 VSS 0.05956f
C18301 DVDD.n14867 VSS 0.05956f
C18302 DVDD.n14868 VSS 0.063725f
C18303 DVDD.n14869 VSS 0.066098f
C18304 DVDD.n14870 VSS 0.028497f
C18305 DVDD.n14871 VSS 0.031128f
C18306 DVDD.n14872 VSS 0.031128f
C18307 DVDD.n14873 VSS 0.031128f
C18308 DVDD.n14874 VSS 0.031128f
C18309 DVDD.n14875 VSS 0.031128f
C18310 DVDD.n14876 VSS 0.031128f
C18311 DVDD.n14877 VSS 0.031128f
C18312 DVDD.n14878 VSS 0.031128f
C18313 DVDD.n14879 VSS 0.031128f
C18314 DVDD.n14880 VSS 0.031128f
C18315 DVDD.n14881 VSS 0.031128f
C18316 DVDD.n14882 VSS 0.031128f
C18317 DVDD.n14883 VSS 0.031128f
C18318 DVDD.n14884 VSS 0.031128f
C18319 DVDD.n14885 VSS 0.031128f
C18320 DVDD.n14886 VSS 0.031128f
C18321 DVDD.n14887 VSS 0.031128f
C18322 DVDD.n14888 VSS 0.031128f
C18323 DVDD.n14889 VSS 0.031128f
C18324 DVDD.n14890 VSS 0.031128f
C18325 DVDD.n14891 VSS 0.031128f
C18326 DVDD.n14892 VSS 0.031128f
C18327 DVDD.n14893 VSS 0.031128f
C18328 DVDD.n14894 VSS 0.031128f
C18329 DVDD.n14895 VSS 0.031128f
C18330 DVDD.n14896 VSS 0.031128f
C18331 DVDD.n14897 VSS 0.031128f
C18332 DVDD.n14898 VSS 0.031128f
C18333 DVDD.n14899 VSS 0.031128f
C18334 DVDD.n14900 VSS 0.031128f
C18335 DVDD.n14901 VSS 0.031128f
C18336 DVDD.n14902 VSS 0.031128f
C18337 DVDD.n14903 VSS 0.031128f
C18338 DVDD.n14904 VSS 0.031128f
C18339 DVDD.n14905 VSS 0.031128f
C18340 DVDD.n14906 VSS 0.031128f
C18341 DVDD.n14907 VSS 0.031128f
C18342 DVDD.n14908 VSS 0.031128f
C18343 DVDD.n14909 VSS 0.031128f
C18344 DVDD.n14910 VSS 0.031128f
C18345 DVDD.n14911 VSS 0.031128f
C18346 DVDD.n14912 VSS 0.031128f
C18347 DVDD.n14913 VSS 0.031128f
C18348 DVDD.n14914 VSS 0.031128f
C18349 DVDD.n14915 VSS 0.031128f
C18350 DVDD.n14916 VSS 0.031128f
C18351 DVDD.n14917 VSS 0.031128f
C18352 DVDD.n14918 VSS 0.031128f
C18353 DVDD.n14919 VSS 0.031128f
C18354 DVDD.n14920 VSS 0.031128f
C18355 DVDD.n14921 VSS 0.031128f
C18356 DVDD.n14922 VSS 0.031128f
C18357 DVDD.n14923 VSS 0.031128f
C18358 DVDD.n14924 VSS 0.031128f
C18359 DVDD.n14925 VSS 0.031128f
C18360 DVDD.n14926 VSS 0.031128f
C18361 DVDD.n14927 VSS 0.031128f
C18362 DVDD.n14928 VSS 0.031128f
C18363 DVDD.n14929 VSS 0.031128f
C18364 DVDD.n14930 VSS 0.031128f
C18365 DVDD.n14931 VSS 0.031128f
C18366 DVDD.n14932 VSS 0.031128f
C18367 DVDD.n14933 VSS 0.031128f
C18368 DVDD.n14934 VSS 0.031128f
C18369 DVDD.n14935 VSS 0.031128f
C18370 DVDD.n14936 VSS 0.031128f
C18371 DVDD.n14937 VSS 0.031128f
C18372 DVDD.n14938 VSS 0.031128f
C18373 DVDD.n14939 VSS 0.031128f
C18374 DVDD.n14940 VSS 0.031128f
C18375 DVDD.n14941 VSS 0.031128f
C18376 DVDD.n14942 VSS 0.031128f
C18377 DVDD.n14943 VSS 0.031128f
C18378 DVDD.n14944 VSS 0.031128f
C18379 DVDD.n14945 VSS 0.031128f
C18380 DVDD.n14946 VSS 0.031128f
C18381 DVDD.n14947 VSS 0.031128f
C18382 DVDD.n14948 VSS 0.031128f
C18383 DVDD.n14949 VSS 0.031128f
C18384 DVDD.n14950 VSS 0.031128f
C18385 DVDD.n14951 VSS 0.031128f
C18386 DVDD.n14952 VSS 0.031128f
C18387 DVDD.n14953 VSS 0.031128f
C18388 DVDD.n14954 VSS 0.031128f
C18389 DVDD.n14955 VSS 0.031128f
C18390 DVDD.n14956 VSS 0.031128f
C18391 DVDD.n14957 VSS 0.031128f
C18392 DVDD.n14958 VSS 0.031128f
C18393 DVDD.n14959 VSS 0.031128f
C18394 DVDD.n14960 VSS 0.031128f
C18395 DVDD.n14961 VSS 0.031128f
C18396 DVDD.n14962 VSS 0.031128f
C18397 DVDD.n14963 VSS 0.031128f
C18398 DVDD.n14964 VSS 0.031128f
C18399 DVDD.n14965 VSS 0.031128f
C18400 DVDD.n14966 VSS 0.031128f
C18401 DVDD.n14967 VSS 0.031128f
C18402 DVDD.n14968 VSS 0.031128f
C18403 DVDD.n14969 VSS 0.031128f
C18404 DVDD.n14970 VSS 0.031128f
C18405 DVDD.n14971 VSS 0.031128f
C18406 DVDD.n14972 VSS 0.031128f
C18407 DVDD.n14973 VSS 0.031128f
C18408 DVDD.n14974 VSS 0.031128f
C18409 DVDD.n14975 VSS 0.031128f
C18410 DVDD.n14976 VSS 0.031128f
C18411 DVDD.n14977 VSS 0.031128f
C18412 DVDD.n14978 VSS 0.031128f
C18413 DVDD.n14979 VSS 0.031128f
C18414 DVDD.n14980 VSS 0.031128f
C18415 DVDD.n14981 VSS 0.031128f
C18416 DVDD.n14982 VSS 0.031128f
C18417 DVDD.n14983 VSS 0.031128f
C18418 DVDD.n14984 VSS 0.031128f
C18419 DVDD.n14985 VSS 0.031128f
C18420 DVDD.n14986 VSS 0.031128f
C18421 DVDD.n14987 VSS 0.031128f
C18422 DVDD.n14988 VSS 0.031128f
C18423 DVDD.n14989 VSS 0.031128f
C18424 DVDD.n14990 VSS 0.031128f
C18425 DVDD.n14991 VSS 0.031128f
C18426 DVDD.n14992 VSS 0.031128f
C18427 DVDD.n14993 VSS 0.031128f
C18428 DVDD.n14994 VSS 0.031128f
C18429 DVDD.n14995 VSS 0.031128f
C18430 DVDD.n14996 VSS 0.031128f
C18431 DVDD.n14997 VSS 0.031128f
C18432 DVDD.n14998 VSS 0.031128f
C18433 DVDD.n14999 VSS 0.031128f
C18434 DVDD.n15000 VSS 0.031128f
C18435 DVDD.n15001 VSS 0.031128f
C18436 DVDD.n15002 VSS 0.031128f
C18437 DVDD.n15003 VSS 0.031128f
C18438 DVDD.n15004 VSS 0.031128f
C18439 DVDD.n15005 VSS 0.031128f
C18440 DVDD.n15006 VSS 0.031128f
C18441 DVDD.n15007 VSS 0.031128f
C18442 DVDD.n15008 VSS 0.031128f
C18443 DVDD.n15009 VSS 0.031128f
C18444 DVDD.n15010 VSS 0.031128f
C18445 DVDD.n15011 VSS 0.031128f
C18446 DVDD.n15012 VSS 0.031128f
C18447 DVDD.n15013 VSS 0.031128f
C18448 DVDD.n15014 VSS 0.031128f
C18449 DVDD.n15015 VSS 0.031128f
C18450 DVDD.n15016 VSS 0.031128f
C18451 DVDD.n15017 VSS 0.031128f
C18452 DVDD.n15018 VSS 0.031128f
C18453 DVDD.n15019 VSS 0.031128f
C18454 DVDD.n15020 VSS 0.031128f
C18455 DVDD.n15021 VSS 0.031128f
C18456 DVDD.n15022 VSS 0.031128f
C18457 DVDD.n15023 VSS 0.031128f
C18458 DVDD.n15024 VSS 0.031128f
C18459 DVDD.n15025 VSS 0.031128f
C18460 DVDD.n15026 VSS 0.031128f
C18461 DVDD.n15027 VSS 0.031128f
C18462 DVDD.n15028 VSS 0.031128f
C18463 DVDD.n15029 VSS 0.031128f
C18464 DVDD.n15030 VSS 0.031128f
C18465 DVDD.n15031 VSS 0.031128f
C18466 DVDD.n15032 VSS 0.031128f
C18467 DVDD.n15033 VSS 0.031128f
C18468 DVDD.n15034 VSS 0.031128f
C18469 DVDD.n15035 VSS 0.031128f
C18470 DVDD.n15036 VSS 0.031128f
C18471 DVDD.n15037 VSS 0.031128f
C18472 DVDD.n15038 VSS 0.031128f
C18473 DVDD.n15039 VSS 0.031128f
C18474 DVDD.n15040 VSS 0.031128f
C18475 DVDD.n15041 VSS 0.031128f
C18476 DVDD.n15042 VSS 0.031128f
C18477 DVDD.n15043 VSS 0.031128f
C18478 DVDD.n15044 VSS 0.031128f
C18479 DVDD.n15045 VSS 0.031128f
C18480 DVDD.n15046 VSS 0.031128f
C18481 DVDD.n15047 VSS 0.031128f
C18482 DVDD.n15048 VSS 0.031128f
C18483 DVDD.n15049 VSS 0.031128f
C18484 DVDD.n15050 VSS 0.031128f
C18485 DVDD.n15051 VSS 0.031128f
C18486 DVDD.n15052 VSS 0.031128f
C18487 DVDD.n15053 VSS 0.031128f
C18488 DVDD.n15054 VSS 0.026086f
C18489 DVDD.n15055 VSS 0.019729f
C18490 DVDD.n15056 VSS 0.019729f
C18491 DVDD.n15057 VSS 0.290608f
C18492 DVDD.n15058 VSS 0.019729f
C18493 DVDD.n15060 VSS 0.366419f
C18494 DVDD.n15061 VSS 0.244279f
C18495 DVDD.n15062 VSS 0.03381f
C18496 DVDD.n15063 VSS 0.03381f
C18497 DVDD.n15064 VSS 0.029529f
C18498 DVDD.n15065 VSS 0.036621f
C18499 DVDD.n15066 VSS 0.02205f
C18500 DVDD.n15067 VSS 0.025247f
C18501 DVDD.n15068 VSS 0.025247f
C18502 DVDD.n15069 VSS 0.214797f
C18503 DVDD.n15070 VSS 0.387477f
C18504 DVDD.n15071 VSS 0.036505f
C18505 DVDD.n15072 VSS 0.036505f
C18506 DVDD.n15073 VSS 0.032585f
C18507 DVDD.n15074 VSS 0.039516f
C18508 DVDD.n15075 VSS 0.047162f
C18509 DVDD.n15076 VSS 0.052836f
C18510 DVDD.n15077 VSS 0.052836f
C18511 DVDD.n15078 VSS 0.210585f
C18512 DVDD.n15079 VSS 0.522252f
C18513 DVDD.n15080 VSS 0.037649f
C18514 DVDD.n15081 VSS 0.037649f
C18515 DVDD.n15082 VSS 0.032881f
C18516 DVDD.n15083 VSS 0.036621f
C18517 DVDD.n15084 VSS 0.018697f
C18518 DVDD.n15085 VSS 0.021408f
C18519 DVDD.n15086 VSS 0.02513f
C18520 DVDD.n15087 VSS 0.019729f
C18521 DVDD.n15088 VSS 0.019729f
C18522 DVDD.n15089 VSS 0.374843f
C18523 DVDD.n15090 VSS 0.019729f
C18524 DVDD.n15092 VSS 0.598063f
C18525 DVDD.n15093 VSS 0.046111f
C18526 DVDD.n15094 VSS 0.046111f
C18527 DVDD.n15095 VSS 0.04116f
C18528 DVDD.n15096 VSS 0.053165f
C18529 DVDD.n15097 VSS 0.04459f
C18530 DVDD.n15098 VSS 0.049954f
C18531 DVDD.n15099 VSS 0.049954f
C18532 DVDD.n15100 VSS 0.189527f
C18533 DVDD.n15101 VSS 0.450653f
C18534 DVDD.n15102 VSS 0.480135f
C18535 DVDD.n15103 VSS 0.024361f
C18536 DVDD.n15104 VSS 0.024361f
C18537 DVDD.n15105 VSS 0.021276f
C18538 DVDD.n15106 VSS 0.036621f
C18539 DVDD.n15107 VSS 0.030302f
C18540 DVDD.n15108 VSS 0.034696f
C18541 DVDD.n15109 VSS 0.02513f
C18542 DVDD.n15110 VSS 0.019729f
C18543 DVDD.n15111 VSS 0.019729f
C18544 DVDD.n15112 VSS 0.44223f
C18545 DVDD.n15113 VSS 0.496982f
C18546 DVDD.n15114 VSS 0.032662f
C18547 DVDD.n15115 VSS 0.032662f
C18548 DVDD.n15116 VSS 0.029155f
C18549 DVDD.n15117 VSS 0.053165f
C18550 DVDD.n15118 VSS 0.053165f
C18551 DVDD.n15119 VSS 0.054277f
C18552 DVDD.n15120 VSS 0.054277f
C18553 DVDD.n15121 VSS 0.598063f
C18554 DVDD.n15122 VSS 0.522252f
C18555 DVDD.n15123 VSS 0.025247f
C18556 DVDD.n15124 VSS 0.025247f
C18557 DVDD.n15125 VSS 0.02205f
C18558 DVDD.n15126 VSS 0.10523f
C18559 DVDD.n15127 VSS 0.132934f
C18560 DVDD.n15128 VSS 0.058284f
C18561 DVDD.n15129 VSS 0.050805f
C18562 DVDD.n15130 VSS 0.050805f
C18563 DVDD.n15131 VSS 1.29721f
C18564 DVDD.n15132 VSS 0.063957f
C18565 DVDD.n15133 VSS 0.063957f
C18566 DVDD.n15134 VSS 0.063957f
C18567 DVDD.n15135 VSS 0.050031f
C18568 DVDD.n15136 VSS 0.044635f
C18569 DVDD.n15138 VSS 0.051878f
C18570 DVDD.n15139 VSS 0.277828f
C18571 DVDD.n15140 VSS 0.088457f
C18572 DVDD.n15141 VSS 0.028297f
C18573 DVDD.n15142 VSS 0.379993f
C18574 DVDD.n15143 VSS 0.36811f
C18575 DVDD.n15144 VSS 0.06615f
C18576 DVDD.n15145 VSS 0.035233f
C18577 DVDD.n15146 VSS 0.035233f
C18578 DVDD.n15147 VSS 0.06615f
C18579 DVDD.n15148 VSS 0.026573f
C18580 DVDD.n15149 VSS 0.013761f
C18581 DVDD.n15150 VSS 0.025624f
C18582 DVDD.n15151 VSS 0.132299f
C18583 DVDD.n15152 VSS 0.132299f
C18584 DVDD.n15153 VSS 0.132299f
C18585 DVDD.n15154 VSS 0.025624f
C18586 DVDD.n15155 VSS 0.025624f
C18587 DVDD.n15156 VSS 0.025624f
C18588 DVDD.n15157 VSS 0.132299f
C18589 DVDD.n15158 VSS 0.132299f
C18590 DVDD.n15159 VSS 0.132299f
C18591 DVDD.n15160 VSS 0.025624f
C18592 DVDD.n15161 VSS 0.025624f
C18593 DVDD.n15162 VSS 0.025624f
C18594 DVDD.n15163 VSS 0.132299f
C18595 DVDD.n15164 VSS 0.132299f
C18596 DVDD.n15165 VSS 0.132299f
C18597 DVDD.n15166 VSS 0.025624f
C18598 DVDD.n15167 VSS 0.025624f
C18599 DVDD.n15168 VSS 0.025624f
C18600 DVDD.n15169 VSS 0.132299f
C18601 DVDD.n15170 VSS 0.132299f
C18602 DVDD.n15171 VSS 0.132299f
C18603 DVDD.n15172 VSS 0.025624f
C18604 DVDD.n15173 VSS 0.025624f
C18605 DVDD.n15174 VSS 0.025624f
C18606 DVDD.n15175 VSS 0.132299f
C18607 DVDD.n15176 VSS 0.132299f
C18608 DVDD.n15177 VSS 0.132299f
C18609 DVDD.n15178 VSS 0.025624f
C18610 DVDD.n15179 VSS 0.025624f
C18611 DVDD.n15180 VSS 0.025624f
C18612 DVDD.n15181 VSS 0.132299f
C18613 DVDD.n15182 VSS 0.132299f
C18614 DVDD.n15183 VSS 0.132299f
C18615 DVDD.n15184 VSS 0.025624f
C18616 DVDD.n15185 VSS 0.025624f
C18617 DVDD.n15186 VSS 0.025624f
C18618 DVDD.n15187 VSS 0.132299f
C18619 DVDD.n15188 VSS 0.132299f
C18620 DVDD.n15189 VSS 0.132299f
C18621 DVDD.n15190 VSS 0.025624f
C18622 DVDD.n15191 VSS 0.025624f
C18623 DVDD.n15192 VSS 0.025624f
C18624 DVDD.n15193 VSS 0.132299f
C18625 DVDD.n15194 VSS 0.132299f
C18626 DVDD.n15195 VSS 0.132299f
C18627 DVDD.n15196 VSS 0.025624f
C18628 DVDD.n15197 VSS 0.025624f
C18629 DVDD.n15198 VSS 0.025624f
C18630 DVDD.n15199 VSS 0.132299f
C18631 DVDD.n15200 VSS 0.132299f
C18632 DVDD.n15201 VSS 0.132299f
C18633 DVDD.n15202 VSS 0.025624f
C18634 DVDD.n15203 VSS 0.025624f
C18635 DVDD.n15204 VSS 0.025624f
C18636 DVDD.n15205 VSS 0.132299f
C18637 DVDD.n15206 VSS 0.132299f
C18638 DVDD.n15207 VSS 0.132299f
C18639 DVDD.n15208 VSS 0.025624f
C18640 DVDD.n15209 VSS 0.025624f
C18641 DVDD.n15210 VSS 0.025624f
C18642 DVDD.n15211 VSS 0.132299f
C18643 DVDD.n15212 VSS 0.132299f
C18644 DVDD.n15213 VSS 0.132299f
C18645 DVDD.n15214 VSS 0.025624f
C18646 DVDD.n15215 VSS 0.025624f
C18647 DVDD.n15216 VSS 0.025624f
C18648 DVDD.n15217 VSS 0.132299f
C18649 DVDD.n15218 VSS 0.132299f
C18650 DVDD.n15219 VSS 0.132299f
C18651 DVDD.n15220 VSS 0.025624f
C18652 DVDD.n15221 VSS 0.025624f
C18653 DVDD.n15222 VSS 0.025624f
C18654 DVDD.n15223 VSS 0.132299f
C18655 DVDD.n15224 VSS 0.132299f
C18656 DVDD.n15225 VSS 0.132299f
C18657 DVDD.n15226 VSS 0.025624f
C18658 DVDD.n15227 VSS 0.025624f
C18659 DVDD.n15228 VSS 0.025624f
C18660 DVDD.n15229 VSS 0.132299f
C18661 DVDD.n15230 VSS 0.132299f
C18662 DVDD.n15231 VSS 0.132299f
C18663 DVDD.n15232 VSS 0.025624f
C18664 DVDD.n15233 VSS 0.025624f
C18665 DVDD.n15234 VSS 0.025624f
C18666 DVDD.n15235 VSS 0.132299f
C18667 DVDD.n15236 VSS 0.132299f
C18668 DVDD.n15237 VSS 0.132299f
C18669 DVDD.n15238 VSS 0.025624f
C18670 DVDD.n15239 VSS 0.025624f
C18671 DVDD.n15240 VSS 0.025624f
C18672 DVDD.n15241 VSS 0.132299f
C18673 DVDD.n15242 VSS 0.132299f
C18674 DVDD.n15243 VSS 0.132299f
C18675 DVDD.n15244 VSS 0.025624f
C18676 DVDD.n15245 VSS 0.025624f
C18677 DVDD.n15246 VSS 0.025624f
C18678 DVDD.n15247 VSS 0.132299f
C18679 DVDD.n15248 VSS 0.132299f
C18680 DVDD.n15249 VSS 0.132299f
C18681 DVDD.n15250 VSS 0.025624f
C18682 DVDD.n15251 VSS 0.025624f
C18683 DVDD.n15252 VSS 0.025624f
C18684 DVDD.n15253 VSS 0.132299f
C18685 DVDD.n15254 VSS 0.132299f
C18686 DVDD.n15255 VSS 0.132299f
C18687 DVDD.n15256 VSS 0.025624f
C18688 DVDD.n15257 VSS 0.025624f
C18689 DVDD.n15258 VSS 0.025624f
C18690 DVDD.n15259 VSS 0.132299f
C18691 DVDD.n15260 VSS 0.132299f
C18692 DVDD.n15261 VSS 0.132299f
C18693 DVDD.n15262 VSS 0.025624f
C18694 DVDD.n15263 VSS 0.025624f
C18695 DVDD.n15264 VSS 0.025624f
C18696 DVDD.n15265 VSS 0.132299f
C18697 DVDD.n15266 VSS 0.132299f
C18698 DVDD.n15267 VSS 0.132299f
C18699 DVDD.n15268 VSS 0.025624f
C18700 DVDD.n15269 VSS 0.025624f
C18701 DVDD.n15270 VSS 0.025624f
C18702 DVDD.n15271 VSS 0.132299f
C18703 DVDD.n15272 VSS 0.132299f
C18704 DVDD.n15273 VSS 0.132299f
C18705 DVDD.n15274 VSS 0.025624f
C18706 DVDD.n15275 VSS 0.025624f
C18707 DVDD.n15276 VSS 0.025624f
C18708 DVDD.n15277 VSS 0.132299f
C18709 DVDD.n15278 VSS 0.132299f
C18710 DVDD.n15279 VSS 0.132299f
C18711 DVDD.n15280 VSS 0.025624f
C18712 DVDD.n15281 VSS 0.025624f
C18713 DVDD.n15282 VSS 0.025624f
C18714 DVDD.n15283 VSS 0.128624f
C18715 DVDD.n15284 VSS 0.06615f
C18716 DVDD.n15285 VSS 0.373774f
C18717 DVDD.n15286 VSS 0.06615f
C18718 DVDD.n15287 VSS 0.075949f
C18719 DVDD.n15288 VSS 0.025624f
C18720 DVDD.n15289 VSS 0.025624f
C18721 DVDD.n15290 VSS 0.025624f
C18722 DVDD.n15291 VSS 0.132299f
C18723 DVDD.n15292 VSS 0.132299f
C18724 DVDD.n15293 VSS 0.132299f
C18725 DVDD.n15294 VSS 0.025624f
C18726 DVDD.n15295 VSS 0.025624f
C18727 DVDD.n15296 VSS 0.025624f
C18728 DVDD.n15297 VSS 0.132299f
C18729 DVDD.n15298 VSS 0.132299f
C18730 DVDD.n15299 VSS 0.132299f
C18731 DVDD.n15300 VSS 0.025624f
C18732 DVDD.n15301 VSS 0.025624f
C18733 DVDD.n15302 VSS 0.025624f
C18734 DVDD.n15303 VSS 0.132299f
C18735 DVDD.n15304 VSS 0.132299f
C18736 DVDD.n15305 VSS 0.132299f
C18737 DVDD.n15306 VSS 0.019218f
C18738 DVDD.n15307 VSS -3.16672f
C18739 DVDD.n15308 VSS 0.019218f
C18740 DVDD.n15309 VSS 0.025624f
C18741 DVDD.n15310 VSS 0.132299f
C18742 DVDD.n15311 VSS 0.132299f
C18743 DVDD.n15312 VSS 0.132299f
C18744 DVDD.n15313 VSS 0.025624f
C18745 DVDD.n15314 VSS 0.025624f
C18746 DVDD.n15315 VSS 0.025624f
C18747 DVDD.n15316 VSS 0.100449f
C18748 DVDD.n15317 VSS 0.128624f
C18749 DVDD.n15318 VSS 0.11992f
C18750 DVDD.n15319 VSS 0.274656f
C18751 DVDD.n15320 VSS 0.274656f
C18752 DVDD.n15321 VSS 0.11992f
C18753 DVDD.n15322 VSS 0.274656f
C18754 DVDD.n15323 VSS 1.26285f
C18755 DVDD.n15324 VSS 0.737752f
C18756 DVDD.n15325 VSS 0.11992f
C18757 DVDD.n15326 VSS 0.355263f
C18758 DVDD.n15327 VSS 0.11992f
C18759 DVDD.n15328 VSS 0.274656f
C18760 DVDD.n15329 VSS 0.11992f
C18761 DVDD.n15330 VSS 0.274656f
C18762 DVDD.n15331 VSS 0.274656f
C18763 DVDD.n15332 VSS 0.274656f
C18764 DVDD.n15333 VSS 0.274656f
C18765 DVDD.n15334 VSS 0.11992f
C18766 DVDD.n15335 VSS 0.274656f
C18767 DVDD.n15336 VSS 0.11992f
C18768 DVDD.n15337 VSS 0.274656f
C18769 DVDD.n15338 VSS 0.11992f
C18770 DVDD.n15339 VSS 0.274656f
C18771 DVDD.n15340 VSS 0.274656f
C18772 DVDD.n15341 VSS 0.274656f
C18773 DVDD.n15342 VSS 0.274656f
C18774 DVDD.n15343 VSS 0.274656f
C18775 DVDD.n15344 VSS 0.274656f
C18776 DVDD.n15345 VSS 0.274656f
C18777 DVDD.n15346 VSS 0.274656f
C18778 DVDD.n15347 VSS 0.183749f
C18779 DVDD.n15348 VSS 0.330748f
C18780 DVDD.n15349 VSS 0.274656f
C18781 DVDD.n15350 VSS 0.228235f
C18782 DVDD.n15351 VSS 0.274656f
C18783 DVDD.n15352 VSS 0.274656f
C18784 DVDD.n15353 VSS 0.274656f
C18785 DVDD.n15354 VSS 0.274656f
C18786 DVDD.n15355 VSS 0.274656f
C18787 DVDD.n15356 VSS 0.274656f
C18788 DVDD.n15357 VSS 0.274656f
C18789 DVDD.n15358 VSS 0.274656f
C18790 DVDD.n15359 VSS 0.274656f
C18791 DVDD.n15360 VSS 0.274656f
C18792 DVDD.n15361 VSS 0.274656f
C18793 DVDD.n15362 VSS 0.274656f
C18794 DVDD.n15363 VSS 0.274656f
C18795 DVDD.n15364 VSS 0.274656f
C18796 DVDD.n15365 VSS 0.274656f
C18797 DVDD.n15366 VSS 0.11992f
C18798 DVDD.n15367 VSS 0.274656f
C18799 DVDD.n15368 VSS 0.11992f
C18800 DVDD.n15369 VSS 0.274656f
C18801 DVDD.n15370 VSS 0.11992f
C18802 DVDD.n15371 VSS 0.274656f
C18803 DVDD.n15372 VSS 0.11992f
C18804 DVDD.n15373 VSS 0.274656f
C18805 DVDD.n15374 VSS 0.11992f
C18806 DVDD.n15375 VSS 0.274656f
C18807 DVDD.n15376 VSS 0.11992f
C18808 DVDD.n15377 VSS 0.274656f
C18809 DVDD.n15378 VSS 0.11992f
C18810 DVDD.n15379 VSS 0.274656f
C18811 DVDD.n15380 VSS 0.11992f
C18812 DVDD.n15381 VSS 0.274656f
C18813 DVDD.n15382 VSS 0.11992f
C18814 DVDD.n15383 VSS 0.274656f
C18815 DVDD.n15384 VSS 0.11992f
C18816 DVDD.n15385 VSS 0.274656f
C18817 DVDD.n15386 VSS 0.11992f
C18818 DVDD.n15387 VSS 0.274656f
C18819 DVDD.n15388 VSS 0.11992f
C18820 DVDD.n15389 VSS 0.274656f
C18821 DVDD.n15390 VSS 0.239841f
C18822 DVDD.n15391 VSS 0.274656f
C18823 DVDD.n15392 VSS 0.274656f
C18824 DVDD.n15393 VSS 0.228235f
C18825 DVDD.n15394 VSS 0.228235f
C18826 DVDD.n15395 VSS 0.330748f
C18827 DVDD.n15396 VSS 0.183749f
C18828 DVDD.n15397 VSS 0.183749f
C18829 DVDD.n15398 VSS 0.274656f
C18830 DVDD.n15399 VSS 0.274656f
C18831 DVDD.n15400 VSS 0.11992f
C18832 DVDD.n15401 VSS 0.274656f
C18833 DVDD.n15402 VSS 0.11992f
C18834 DVDD.n15403 VSS 0.274656f
C18835 DVDD.n15404 VSS 0.274656f
C18836 DVDD.n15405 VSS 0.11992f
C18837 DVDD.n15406 VSS 0.130558f
C18838 DVDD.n15407 VSS 0.06615f
C18839 DVDD.n15408 VSS 0.137328f
C18840 DVDD.n15409 VSS 0.06615f
C18841 DVDD.n15410 VSS 0.07105f
C18842 DVDD.n15411 VSS 0.132299f
C18843 DVDD.n15412 VSS 0.025624f
C18844 DVDD.n15413 VSS 0.025624f
C18845 DVDD.n15414 VSS 0.025624f
C18846 DVDD.n15415 VSS 0.075949f
C18847 DVDD.n15416 VSS 0.137328f
C18848 DVDD.n15418 VSS 0.130558f
C18849 DVDD.n15419 VSS 0.137328f
C18850 DVDD.n15420 VSS 0.137328f
C18851 DVDD.n15421 VSS 0.137328f
C18852 DVDD.n15423 VSS 0.128624f
C18853 DVDD.n15424 VSS 0.737752f
C18854 DVDD.n15425 VSS 1.26285f
C18855 DVDD.n15426 VSS 0.274656f
C18856 DVDD.n15427 VSS 0.274656f
C18857 DVDD.n15428 VSS 0.274656f
C18858 DVDD.n15429 VSS 0.274656f
C18859 DVDD.n15430 VSS 0.274656f
C18860 DVDD.n15431 VSS 0.274656f
C18861 DVDD.n15432 VSS 0.274656f
C18862 DVDD.n15433 VSS 0.274656f
C18863 DVDD.n15434 VSS 0.274656f
C18864 DVDD.n15435 VSS 0.274656f
C18865 DVDD.n15436 VSS 0.274656f
C18866 DVDD.n15437 VSS 0.11992f
C18867 DVDD.n15438 VSS 0.274656f
C18868 DVDD.n15439 VSS 0.11992f
C18869 DVDD.n15440 VSS 0.274656f
C18870 DVDD.n15441 VSS 0.11992f
C18871 DVDD.n15442 VSS 0.274656f
C18872 DVDD.n15443 VSS 0.11992f
C18873 DVDD.n15444 VSS 0.274656f
C18874 DVDD.n15445 VSS 0.11992f
C18875 DVDD.n15446 VSS 0.274656f
C18876 DVDD.n15447 VSS 0.11992f
C18877 DVDD.n15448 VSS 0.274656f
C18878 DVDD.n15449 VSS 0.11992f
C18879 DVDD.n15450 VSS 0.274656f
C18880 DVDD.n15451 VSS 0.11992f
C18881 DVDD.n15452 VSS 0.274656f
C18882 DVDD.n15453 VSS 0.11992f
C18883 DVDD.n15454 VSS 0.274656f
C18884 DVDD.n15455 VSS 0.11992f
C18885 DVDD.n15456 VSS 0.274656f
C18886 DVDD.n15457 VSS 0.355263f
C18887 DVDD.n15458 VSS 0.11992f
C18888 DVDD.n15459 VSS 0.803653f
C18889 DVDD.n15460 VSS 0.06615f
C18890 DVDD.n15461 VSS 0.137328f
C18891 DVDD.n15462 VSS 0.217597f
C18892 DVDD.n15463 VSS 0.183749f
C18893 DVDD.n15464 VSS 0.183749f
C18894 DVDD.n15465 VSS 0.183749f
C18895 DVDD.n15466 VSS 0.524168f
C18896 DVDD.n15467 VSS 0.274656f
C18897 DVDD.n15468 VSS 0.228235f
C18898 DVDD.n15469 VSS 0.228235f
C18899 DVDD.n15470 VSS 0.228235f
C18900 DVDD.n15471 VSS 0.274656f
C18901 DVDD.n15472 VSS 0.239841f
C18902 DVDD.n15473 VSS 0.274656f
C18903 DVDD.n15474 VSS 0.11992f
C18904 DVDD.n15475 VSS 0.274656f
C18905 DVDD.n15476 VSS 0.11992f
C18906 DVDD.n15477 VSS 0.274656f
C18907 DVDD.n15478 VSS 0.274656f
C18908 DVDD.n15479 VSS 0.274656f
C18909 DVDD.n15480 VSS 0.274656f
C18910 DVDD.n15481 VSS 0.11992f
C18911 DVDD.n15482 VSS 0.274656f
C18912 DVDD.n15483 VSS 0.11992f
C18913 DVDD.n15484 VSS 0.274656f
C18914 DVDD.n15485 VSS 0.11992f
C18915 DVDD.n15486 VSS 0.274656f
C18916 DVDD.n15487 VSS 0.274656f
C18917 DVDD.n15488 VSS 0.274656f
C18918 DVDD.n15489 VSS 0.274656f
C18919 DVDD.n15490 VSS 0.11992f
C18920 DVDD.n15491 VSS 0.274656f
C18921 DVDD.n15492 VSS 0.11992f
C18922 DVDD.n15493 VSS 0.274656f
C18923 DVDD.n15494 VSS 0.11992f
C18924 DVDD.n15495 VSS 0.274656f
C18925 DVDD.n15496 VSS 0.274656f
C18926 DVDD.n15497 VSS 0.274656f
C18927 DVDD.n15498 VSS 0.274656f
C18928 DVDD.n15499 VSS 0.274656f
C18929 DVDD.n15500 VSS 0.274656f
C18930 DVDD.n15501 VSS 0.274656f
C18931 DVDD.n15502 VSS 0.274656f
C18932 DVDD.n15503 VSS 0.274656f
C18933 DVDD.n15504 VSS 0.274656f
C18934 DVDD.n15505 VSS 0.274656f
C18935 DVDD.n15506 VSS 0.274656f
C18936 DVDD.n15507 VSS 0.11992f
C18937 DVDD.n15508 VSS 0.274656f
C18938 DVDD.n15509 VSS 0.11992f
C18939 DVDD.n15510 VSS 0.274656f
C18940 DVDD.n15511 VSS 0.274656f
C18941 DVDD.n15512 VSS 0.197288f
C18942 DVDD.n15513 VSS 0.274656f
C18943 DVDD.n15514 VSS 0.274656f
C18944 DVDD.n15515 VSS 0.274656f
C18945 DVDD.n15516 VSS 0.274656f
C18946 DVDD.n15517 VSS 0.274656f
C18947 DVDD.n15518 VSS 0.274656f
C18948 DVDD.n15519 VSS 0.11992f
C18949 DVDD.n15520 VSS 0.137328f
C18950 DVDD.n15521 VSS 0.198722f
C18951 DVDD.n15522 VSS 0.081946f
C18952 DVDD.n15523 VSS 0.098809f
C18953 DVDD.t79 VSS 0.425324f
C18954 DVDD.n15524 VSS 0.081946f
C18955 DVDD.n15525 VSS 0.099098f
C18956 DVDD.n15526 VSS 0.198298f
C18957 DVDD.n15527 VSS 0.138779f
C18958 DVDD.n15528 VSS 0.137328f
C18959 DVDD.n15529 VSS 0.183717f
C18960 DVDD.n15530 VSS 0.098809f
C18961 DVDD.t145 VSS 0.167631f
C18962 DVDD.t119 VSS 0.167631f
C18963 DVDD.n15531 VSS 0.335261f
C18964 DVDD.n15532 VSS 0.099098f
C18965 DVDD.n15533 VSS 0.346328f
C18966 DVDD.n15534 VSS 0.210151f
C18967 DVDD.n15535 VSS 0.11992f
C18968 DVDD.n15536 VSS 0.163891f
C18969 DVDD.n15537 VSS 0.198722f
C18970 DVDD.n15538 VSS 0.081946f
C18971 DVDD.n15539 VSS 0.098809f
C18972 DVDD.t140 VSS 0.167631f
C18973 DVDD.t108 VSS 0.167631f
C18974 DVDD.n15540 VSS 0.335261f
C18975 DVDD.n15541 VSS 0.081946f
C18976 DVDD.n15542 VSS 0.099098f
C18977 DVDD.n15543 VSS 0.198298f
C18978 DVDD.n15544 VSS 0.133492f
C18979 DVDD.n15545 VSS 0.163891f
C18980 DVDD.n15546 VSS 0.198722f
C18981 DVDD.n15547 VSS 0.081946f
C18982 DVDD.n15548 VSS 0.098809f
C18983 DVDD.t73 VSS 0.167631f
C18984 DVDD.t104 VSS 0.167631f
C18985 DVDD.n15549 VSS 0.335261f
C18986 DVDD.n15550 VSS 0.081946f
C18987 DVDD.n15551 VSS 0.099098f
C18988 DVDD.n15552 VSS 0.198298f
C18989 DVDD.n15553 VSS 0.138779f
C18990 DVDD.n15554 VSS 0.163891f
C18991 DVDD.n15555 VSS 0.198722f
C18992 DVDD.n15556 VSS 0.081946f
C18993 DVDD.n15557 VSS 0.098809f
C18994 DVDD.t129 VSS 0.167631f
C18995 DVDD.t91 VSS 0.167631f
C18996 DVDD.n15558 VSS 0.335261f
C18997 DVDD.n15559 VSS 0.081946f
C18998 DVDD.n15560 VSS 0.099098f
C18999 DVDD.n15561 VSS 0.198298f
C19000 DVDD.n15562 VSS 0.144066f
C19001 DVDD.n15563 VSS 0.163891f
C19002 DVDD.n15564 VSS 0.198722f
C19003 DVDD.n15565 VSS 0.081946f
C19004 DVDD.n15566 VSS 0.098809f
C19005 DVDD.t118 VSS 0.167631f
C19006 DVDD.t83 VSS 0.167631f
C19007 DVDD.n15567 VSS 0.335261f
C19008 DVDD.n15568 VSS 0.081946f
C19009 DVDD.n15569 VSS 0.099098f
C19010 DVDD.n15570 VSS 0.198298f
C19011 DVDD.n15571 VSS 0.149352f
C19012 DVDD.n15572 VSS 0.163891f
C19013 DVDD.n15573 VSS 0.198722f
C19014 DVDD.n15574 VSS 0.081946f
C19015 DVDD.n15575 VSS 0.098809f
C19016 DVDD.t112 VSS 0.167631f
C19017 DVDD.t97 VSS 0.167631f
C19018 DVDD.n15576 VSS 0.335261f
C19019 DVDD.n15577 VSS 0.081946f
C19020 DVDD.n15578 VSS 0.099098f
C19021 DVDD.n15579 VSS 0.198298f
C19022 DVDD.n15580 VSS 0.154639f
C19023 DVDD.n15581 VSS 0.163891f
C19024 DVDD.n15593 VSS 0.123789f
C19025 DVDD.n15600 VSS 0.137328f
C19026 DVDD.n15601 VSS 0.137328f
C19027 DVDD.n15602 VSS 0.137328f
C19028 DVDD.n15603 VSS 0.121855f
C19029 DVDD.n15604 VSS 0.137328f
C19030 DVDD.n15605 VSS 0.137328f
C19031 DVDD.n15606 VSS 0.098809f
C19032 DVDD.t102 VSS 0.167631f
C19033 DVDD.t90 VSS 0.167631f
C19034 DVDD.n15607 VSS 0.335261f
C19035 DVDD.n15608 VSS 0.099098f
C19036 DVDD.n15609 VSS 0.198298f
C19037 DVDD.n15610 VSS 0.137328f
C19038 DVDD.n15611 VSS 0.137328f
C19039 DVDD.n15613 VSS 0.135394f
C19040 DVDD.n15614 VSS 0.137328f
C19041 DVDD.n15615 VSS 0.137328f
C19042 DVDD.n15616 VSS 0.137328f
C19043 DVDD.n15618 VSS 0.13346f
C19044 DVDD.n15619 VSS 0.11992f
C19045 DVDD.n15620 VSS 0.274656f
C19046 DVDD.n15621 VSS 0.274656f
C19047 DVDD.n15622 VSS 0.274656f
C19048 DVDD.n15623 VSS 0.11992f
C19049 DVDD.n15624 VSS 0.274656f
C19050 DVDD.n15625 VSS 0.274656f
C19051 DVDD.n15626 VSS 0.11992f
C19052 DVDD.n15627 VSS 0.274656f
C19053 DVDD.n15628 VSS 0.274656f
C19054 DVDD.n15629 VSS 0.274656f
C19055 DVDD.n15630 VSS 0.274656f
C19056 DVDD.n15631 VSS 0.11992f
C19057 DVDD.n15632 VSS 0.274656f
C19058 DVDD.n15633 VSS 0.11992f
C19059 DVDD.n15634 VSS 0.274656f
C19060 DVDD.n15635 VSS 0.11992f
C19061 DVDD.n15636 VSS 0.274656f
C19062 DVDD.n15637 VSS 0.274656f
C19063 DVDD.n15638 VSS 0.274656f
C19064 DVDD.n15639 VSS 0.274656f
C19065 DVDD.n15640 VSS 0.11992f
C19066 DVDD.n15641 VSS 0.274656f
C19067 DVDD.n15642 VSS 0.11992f
C19068 DVDD.n15643 VSS 0.274656f
C19069 DVDD.n15644 VSS 0.11992f
C19070 DVDD.n15645 VSS 0.274656f
C19071 DVDD.n15646 VSS 0.274656f
C19072 DVDD.n15647 VSS 0.274656f
C19073 DVDD.n15648 VSS 0.274656f
C19074 DVDD.n15649 VSS 0.11992f
C19075 DVDD.n15650 VSS 0.274656f
C19076 DVDD.n15651 VSS 0.11992f
C19077 DVDD.n15652 VSS 0.274656f
C19078 DVDD.n15653 VSS 0.11992f
C19079 DVDD.n15654 VSS 0.274656f
C19080 DVDD.n15655 VSS 0.274656f
C19081 DVDD.n15656 VSS 0.274656f
C19082 DVDD.n15657 VSS 0.274656f
C19083 DVDD.n15658 VSS 0.274656f
C19084 DVDD.n15659 VSS 0.274656f
C19085 DVDD.n15660 VSS 0.274656f
C19086 DVDD.n15661 VSS 0.274656f
C19087 DVDD.n15662 VSS 0.274656f
C19088 DVDD.n15663 VSS 0.176012f
C19089 DVDD.n15664 VSS 0.274656f
C19090 DVDD.n15665 VSS 0.11992f
C19091 DVDD.n15666 VSS 0.274656f
C19092 DVDD.n15667 VSS 0.11992f
C19093 DVDD.n15668 VSS 0.274656f
C19094 DVDD.n15669 VSS 0.11992f
C19095 DVDD.n15670 VSS 0.274656f
C19096 DVDD.n15671 VSS 0.274656f
C19097 DVDD.n15672 VSS 0.197288f
C19098 DVDD.n15673 VSS 0.274656f
C19099 DVDD.n15674 VSS 0.274656f
C19100 DVDD.n15675 VSS 0.274656f
C19101 DVDD.n15676 VSS 0.274656f
C19102 DVDD.n15677 VSS 0.158604f
C19103 DVDD.n15678 VSS 0.137328f
C19104 DVDD.n15679 VSS 0.307957f
C19105 DVDD.n15680 VSS 0.137328f
C19106 DVDD.n15681 VSS 0.239841f
C19107 DVDD.n15682 VSS 0.274656f
C19108 DVDD.n15683 VSS 0.274656f
C19109 DVDD.n15684 VSS 0.228235f
C19110 DVDD.n15685 VSS 0.228235f
C19111 DVDD.n15686 VSS 0.524168f
C19112 DVDD.n15687 VSS 0.183749f
C19113 DVDD.n15688 VSS 0.217597f
C19114 DVDD.n15689 VSS 0.274656f
C19115 DVDD.n15690 VSS 0.11992f
C19116 DVDD.n15691 VSS 0.274656f
C19117 DVDD.n15692 VSS 0.11992f
C19118 DVDD.n15693 VSS 0.274656f
C19119 DVDD.n15694 VSS 0.11992f
C19120 DVDD.n15695 VSS 0.274656f
C19121 DVDD.n15696 VSS 0.274656f
C19122 DVDD.n15697 VSS 0.11992f
C19123 DVDD.n15698 VSS 0.130558f
C19124 DVDD.n15699 VSS 0.06615f
C19125 DVDD.n15700 VSS 0.803653f
C19126 DVDD.n15701 VSS 0.06615f
C19127 DVDD.n15702 VSS 0.120049f
C19128 DVDD.n15703 VSS 0.025624f
C19129 DVDD.n15704 VSS 0.025624f
C19130 DVDD.n15705 VSS 0.025624f
C19131 DVDD.n15706 VSS 0.093099f
C19132 DVDD.n15707 VSS 0.137328f
C19133 DVDD.n15709 VSS 0.130558f
C19134 DVDD.n15710 VSS 0.137328f
C19135 DVDD.n15711 VSS 0.137328f
C19136 DVDD.n15712 VSS 0.137328f
C19137 DVDD.n15714 VSS 0.128624f
C19138 DVDD.n15715 VSS 0.737752f
C19139 DVDD.n15716 VSS 1.26285f
C19140 DVDD.n15717 VSS 0.274656f
C19141 DVDD.n15718 VSS 0.274656f
C19142 DVDD.n15719 VSS 0.274656f
C19143 DVDD.n15720 VSS 0.274656f
C19144 DVDD.n15721 VSS 0.274656f
C19145 DVDD.n15722 VSS 0.274656f
C19146 DVDD.n15723 VSS 0.274656f
C19147 DVDD.n15724 VSS 0.274656f
C19148 DVDD.n15725 VSS 0.274656f
C19149 DVDD.n15726 VSS 0.274656f
C19150 DVDD.n15727 VSS 0.274656f
C19151 DVDD.n15728 VSS 0.11992f
C19152 DVDD.n15729 VSS 0.274656f
C19153 DVDD.n15730 VSS 0.11992f
C19154 DVDD.n15731 VSS 0.274656f
C19155 DVDD.n15732 VSS 0.11992f
C19156 DVDD.n15733 VSS 0.274656f
C19157 DVDD.n15734 VSS 0.11992f
C19158 DVDD.n15735 VSS 0.274656f
C19159 DVDD.n15736 VSS 0.11992f
C19160 DVDD.n15737 VSS 0.274656f
C19161 DVDD.n15738 VSS 0.11992f
C19162 DVDD.n15739 VSS 0.274656f
C19163 DVDD.n15740 VSS 0.11992f
C19164 DVDD.n15741 VSS 0.274656f
C19165 DVDD.n15742 VSS 0.11992f
C19166 DVDD.n15743 VSS 0.274656f
C19167 DVDD.n15744 VSS 0.11992f
C19168 DVDD.n15745 VSS 0.274656f
C19169 DVDD.n15746 VSS 0.11992f
C19170 DVDD.n15747 VSS 0.274656f
C19171 DVDD.n15748 VSS 0.355263f
C19172 DVDD.n15749 VSS 0.11992f
C19173 DVDD.n15750 VSS 0.803653f
C19174 DVDD.n15751 VSS 0.06615f
C19175 DVDD.n15752 VSS 0.137328f
C19176 DVDD.n15753 VSS 0.217597f
C19177 DVDD.n15754 VSS 0.183749f
C19178 DVDD.n15755 VSS 0.183749f
C19179 DVDD.n15756 VSS 0.183749f
C19180 DVDD.n15757 VSS 0.330748f
C19181 DVDD.n15758 VSS 0.274656f
C19182 DVDD.n15759 VSS 0.228235f
C19183 DVDD.n15760 VSS 0.228235f
C19184 DVDD.n15761 VSS 0.228235f
C19185 DVDD.n15762 VSS 0.274656f
C19186 DVDD.n15763 VSS 0.239841f
C19187 DVDD.n15764 VSS 0.274656f
C19188 DVDD.n15765 VSS 0.11992f
C19189 DVDD.n15766 VSS 0.274656f
C19190 DVDD.n15767 VSS 0.274656f
C19191 DVDD.n15768 VSS 0.274656f
C19192 DVDD.n15769 VSS 0.274656f
C19193 DVDD.n15770 VSS 0.11992f
C19194 DVDD.n15771 VSS 0.274656f
C19195 DVDD.n15772 VSS 0.11992f
C19196 DVDD.n15773 VSS 0.274656f
C19197 DVDD.n15774 VSS 0.11992f
C19198 DVDD.n15775 VSS 0.274656f
C19199 DVDD.n15776 VSS 0.274656f
C19200 DVDD.n15777 VSS 0.274656f
C19201 DVDD.n15778 VSS 0.274656f
C19202 DVDD.n15779 VSS 0.11992f
C19203 DVDD.n15780 VSS 0.274656f
C19204 DVDD.n15781 VSS 0.11992f
C19205 DVDD.n15782 VSS 0.274656f
C19206 DVDD.n15783 VSS 0.11992f
C19207 DVDD.n15784 VSS 0.274656f
C19208 DVDD.n15785 VSS 0.274656f
C19209 DVDD.n15786 VSS 0.274656f
C19210 DVDD.n15787 VSS 0.274656f
C19211 DVDD.n15788 VSS 0.274656f
C19212 DVDD.n15789 VSS 0.11992f
C19213 DVDD.n15790 VSS 0.137328f
C19214 DVDD.n15791 VSS 0.11992f
C19215 DVDD.n15793 VSS 0.13346f
C19216 DVDD.n15794 VSS 0.071372f
C19217 DVDD.n15795 VSS 0.137328f
C19218 DVDD.n15796 VSS 0.11992f
C19219 DVDD.n15797 VSS 0.274656f
C19220 DVDD.n15798 VSS 0.274656f
C19221 DVDD.n15799 VSS 0.274656f
C19222 DVDD.n15800 VSS 0.274656f
C19223 DVDD.n15801 VSS 0.274656f
C19224 DVDD.n15802 VSS 0.274656f
C19225 DVDD.n15803 VSS 0.274656f
C19226 DVDD.n15804 VSS 0.197288f
C19227 DVDD.n15805 VSS 0.274656f
C19228 DVDD.n15806 VSS 0.274656f
C19229 DVDD.n15807 VSS 0.274656f
C19230 DVDD.n15808 VSS 0.274656f
C19231 DVDD.n15809 VSS 0.11992f
C19232 DVDD.n15810 VSS 0.274656f
C19233 DVDD.n15811 VSS 0.11992f
C19234 DVDD.n15812 VSS 0.274656f
C19235 DVDD.n15813 VSS 0.303669f
C19236 DVDD.n15814 VSS 0.048355f
C19237 DVDD.n15815 VSS 0.176012f
C19238 DVDD.n15816 VSS 0.176012f
C19239 DVDD.n15817 VSS 0.330748f
C19240 DVDD.n15818 VSS 0.235972f
C19241 DVDD.n15819 VSS 0.11992f
C19242 DVDD.n15820 VSS 0.235972f
C19243 DVDD.n15821 VSS 0.11992f
C19244 DVDD.n15822 VSS 0.274656f
C19245 DVDD.n15823 VSS 0.274656f
C19246 DVDD.n15824 VSS 0.274656f
C19247 DVDD.n15825 VSS 0.274656f
C19248 DVDD.n15826 VSS 0.11992f
C19249 DVDD.n15827 VSS 0.274656f
C19250 DVDD.n15828 VSS 0.11992f
C19251 DVDD.n15829 VSS 0.274656f
C19252 DVDD.n15830 VSS 0.11992f
C19253 DVDD.n15831 VSS 0.274656f
C19254 DVDD.n15832 VSS 0.274656f
C19255 DVDD.n15833 VSS 0.274656f
C19256 DVDD.n15834 VSS 0.274656f
C19257 DVDD.n15835 VSS 0.274656f
C19258 DVDD.n15836 VSS 0.11992f
C19259 DVDD.n15837 VSS 0.137328f
C19260 DVDD.n15838 VSS 0.071372f
C19261 DVDD.n15839 VSS 0.137328f
C19262 DVDD.n15840 VSS 0.201157f
C19263 DVDD.n15841 VSS 0.274656f
C19264 DVDD.n15842 VSS 0.274656f
C19265 DVDD.n15843 VSS 0.274656f
C19266 DVDD.n15844 VSS 0.274656f
C19267 DVDD.n15845 VSS 0.274656f
C19268 DVDD.n15846 VSS 0.274656f
C19269 DVDD.n15847 VSS 0.274656f
C19270 DVDD.n15848 VSS 0.205025f
C19271 DVDD.n15849 VSS 0.274656f
C19272 DVDD.n15850 VSS 0.274656f
C19273 DVDD.n15851 VSS 0.274656f
C19274 DVDD.n15852 VSS 0.274656f
C19275 DVDD.n15853 VSS 0.274656f
C19276 DVDD.n15854 VSS 0.11992f
C19277 DVDD.n15855 VSS 0.274656f
C19278 DVDD.n15856 VSS 0.11992f
C19279 DVDD.n15857 VSS 0.274656f
C19280 DVDD.n15858 VSS 0.11992f
C19281 DVDD.n15859 VSS 0.274656f
C19282 DVDD.n15860 VSS 0.274656f
C19283 DVDD.n15861 VSS 0.274656f
C19284 DVDD.n15862 VSS 0.274656f
C19285 DVDD.n15863 VSS 0.11992f
C19286 DVDD.n15864 VSS 0.274656f
C19287 DVDD.n15865 VSS 0.11992f
C19288 DVDD.n15866 VSS 0.274656f
C19289 DVDD.n15867 VSS 0.11992f
C19290 DVDD.n15868 VSS 0.274656f
C19291 DVDD.n15869 VSS 0.274656f
C19292 DVDD.n15870 VSS 0.274656f
C19293 DVDD.n15871 VSS 0.168275f
C19294 DVDD.n15872 VSS 0.11992f
C19295 DVDD.n15873 VSS 0.168275f
C19296 DVDD.n15874 VSS 0.274656f
C19297 DVDD.n15875 VSS 0.243709f
C19298 DVDD.n15876 VSS 0.11992f
C19299 DVDD.n15877 VSS 0.243709f
C19300 DVDD.n15878 VSS 0.330748f
C19301 DVDD.n15879 VSS 0.524168f
C19302 DVDD.n15880 VSS 0.11992f
C19303 DVDD.n15881 VSS 0.168275f
C19304 DVDD.n15882 VSS 0.11992f
C19305 DVDD.n15883 VSS 0.274656f
C19306 DVDD.n15884 VSS 0.11992f
C19307 DVDD.n15885 VSS 0.274656f
C19308 DVDD.n15886 VSS 0.11992f
C19309 DVDD.n15887 VSS 0.274656f
C19310 DVDD.n15888 VSS 0.11992f
C19311 DVDD.n15889 VSS 0.274656f
C19312 DVDD.n15890 VSS 0.11992f
C19313 DVDD.n15891 VSS 0.274656f
C19314 DVDD.n15892 VSS 0.11992f
C19315 DVDD.n15893 VSS 0.274656f
C19316 DVDD.n15894 VSS 0.11992f
C19317 DVDD.n15895 VSS 0.274656f
C19318 DVDD.n15896 VSS 0.11992f
C19319 DVDD.n15897 VSS 0.274656f
C19320 DVDD.n15898 VSS 0.274656f
C19321 DVDD.n15899 VSS 0.274656f
C19322 DVDD.n15900 VSS 0.274656f
C19323 DVDD.n15901 VSS 0.274656f
C19324 DVDD.n15902 VSS 0.274656f
C19325 DVDD.n15903 VSS 0.274656f
C19326 DVDD.n15904 VSS 0.274656f
C19327 DVDD.n15905 VSS 0.274656f
C19328 DVDD.n15906 VSS 0.201157f
C19329 DVDD.n15907 VSS 0.137328f
C19330 DVDD.n15908 VSS 0.307957f
C19331 DVDD.n15909 VSS 0.137328f
C19332 DVDD.n15910 VSS 0.11992f
C19333 DVDD.n15911 VSS 0.235972f
C19334 DVDD.n15912 VSS 0.524168f
C19335 DVDD.n15913 VSS 0.524168f
C19336 DVDD.n15914 VSS 0.176012f
C19337 DVDD.n15915 VSS 0.176012f
C19338 DVDD.n15916 VSS 0.524168f
C19339 DVDD.n15917 VSS 0.235972f
C19340 DVDD.n15918 VSS 0.274656f
C19341 DVDD.n15919 VSS 0.11992f
C19342 DVDD.n15920 VSS 0.274656f
C19343 DVDD.n15921 VSS 0.11992f
C19344 DVDD.n15922 VSS 0.274656f
C19345 DVDD.n15923 VSS 0.11992f
C19346 DVDD.n15924 VSS 0.274656f
C19347 DVDD.n15925 VSS 0.274656f
C19348 DVDD.n15926 VSS 0.274656f
C19349 DVDD.n15927 VSS 0.274656f
C19350 DVDD.n15928 VSS 0.11992f
C19351 DVDD.n15929 VSS 0.274656f
C19352 DVDD.n15937 VSS 0.131525f
C19353 DVDD.n15938 VSS 0.11992f
C19354 DVDD.n15939 VSS 0.274656f
C19355 DVDD.n15940 VSS 0.11992f
C19356 DVDD.n15941 VSS 0.274656f
C19357 DVDD.n15942 VSS 0.274656f
C19358 DVDD.n15943 VSS 0.274656f
C19359 DVDD.n15944 VSS 0.274656f
C19360 DVDD.n15945 VSS 0.274656f
C19361 DVDD.n15946 VSS 0.274656f
C19362 DVDD.n15947 VSS 0.274656f
C19363 DVDD.n15948 VSS 0.205025f
C19364 DVDD.n15949 VSS 0.274656f
C19365 DVDD.n15950 VSS 0.274656f
C19366 DVDD.n15951 VSS 0.274656f
C19367 DVDD.n15952 VSS 0.274656f
C19368 DVDD.n15953 VSS 0.274656f
C19369 DVDD.n15954 VSS 0.274656f
C19370 DVDD.n15955 VSS 0.274656f
C19371 DVDD.n15956 VSS 0.274656f
C19372 DVDD.n15957 VSS 0.274656f
C19373 DVDD.n15958 VSS 0.274656f
C19374 DVDD.n15959 VSS 0.274656f
C19375 DVDD.n15960 VSS 0.11992f
C19376 DVDD.n15961 VSS 0.168275f
C19377 DVDD.n15962 VSS 0.11992f
C19378 DVDD.n15963 VSS 0.274656f
C19379 DVDD.n15964 VSS 0.11992f
C19380 DVDD.n15965 VSS 0.274656f
C19381 DVDD.n15966 VSS 0.11992f
C19382 DVDD.n15967 VSS 0.274656f
C19383 DVDD.n15968 VSS 0.11992f
C19384 DVDD.n15969 VSS 0.274656f
C19385 DVDD.n15970 VSS 0.11992f
C19386 DVDD.n15971 VSS 0.274656f
C19387 DVDD.n15972 VSS 0.11992f
C19388 DVDD.n15973 VSS 0.274656f
C19389 DVDD.n15974 VSS 0.11992f
C19390 DVDD.n15975 VSS 0.274656f
C19391 DVDD.n15976 VSS 0.11992f
C19392 DVDD.n15977 VSS 0.274656f
C19393 DVDD.n15978 VSS 0.274656f
C19394 DVDD.n15979 VSS 0.274656f
C19395 DVDD.n15980 VSS 0.274656f
C19396 DVDD.n15981 VSS 0.274656f
C19397 DVDD.n15982 VSS 0.274656f
C19398 DVDD.n15983 VSS 0.274656f
C19399 DVDD.n15984 VSS 0.274656f
C19400 DVDD.n15985 VSS 0.274656f
C19401 DVDD.n15986 VSS 0.201157f
C19402 DVDD.n15987 VSS 0.137328f
C19403 DVDD.n15988 VSS 0.183717f
C19404 DVDD.n15989 VSS 0.098644f
C19405 DVDD.n15990 VSS 0.497089f
C19406 DVDD.n15991 VSS 0.303669f
C19407 DVDD.n15992 VSS 0.048355f
C19408 DVDD.n15993 VSS 0.176012f
C19409 DVDD.n15994 VSS 0.11992f
C19410 DVDD.n15995 VSS 0.274656f
C19411 DVDD.n15996 VSS 0.11992f
C19412 DVDD.n15997 VSS 0.274656f
C19413 DVDD.n15998 VSS 0.11992f
C19414 DVDD.n15999 VSS 0.274656f
C19415 DVDD.n16000 VSS 0.274656f
C19416 DVDD.n16001 VSS 0.197288f
C19417 DVDD.n16002 VSS 0.274656f
C19418 DVDD.n16003 VSS 0.274656f
C19419 DVDD.n16004 VSS 0.274656f
C19420 DVDD.n16005 VSS 0.274656f
C19421 DVDD.n16006 VSS 0.158604f
C19422 DVDD.n16008 VSS 0.163891f
C19423 DVDD.n16009 VSS 0.163891f
C19424 DVDD.n16010 VSS 0.198722f
C19425 DVDD.n16011 VSS 0.081946f
C19426 DVDD.n16012 VSS 0.098809f
C19427 DVDD.t105 VSS 0.167631f
C19428 DVDD.t142 VSS 0.167631f
C19429 DVDD.n16013 VSS 0.335261f
C19430 DVDD.n16014 VSS 0.081946f
C19431 DVDD.n16015 VSS 0.099098f
C19432 DVDD.n16016 VSS 0.198298f
C19433 DVDD.n16018 VSS 0.133492f
C19434 DVDD.n16020 VSS 0.163891f
C19435 DVDD.n16021 VSS 0.163891f
C19436 DVDD.n16022 VSS 0.198722f
C19437 DVDD.n16023 VSS 0.081946f
C19438 DVDD.n16024 VSS 0.098809f
C19439 DVDD.t85 VSS 0.167631f
C19440 DVDD.t110 VSS 0.167631f
C19441 DVDD.n16025 VSS 0.335261f
C19442 DVDD.n16026 VSS 0.081946f
C19443 DVDD.n16027 VSS 0.099098f
C19444 DVDD.n16028 VSS 0.198298f
C19445 DVDD.n16030 VSS 0.122918f
C19446 DVDD.n16032 VSS 0.163891f
C19447 DVDD.n16033 VSS 0.198722f
C19448 DVDD.n16034 VSS 0.081946f
C19449 DVDD.n16035 VSS 0.098809f
C19450 DVDD.t74 VSS 0.167631f
C19451 DVDD.t124 VSS 0.167631f
C19452 DVDD.n16036 VSS 0.335261f
C19453 DVDD.n16037 VSS 0.081946f
C19454 DVDD.n16038 VSS 0.099098f
C19455 DVDD.n16039 VSS 0.198298f
C19456 DVDD.n16040 VSS 0.117632f
C19457 DVDD.n16042 VSS 0.163891f
C19458 DVDD.n16044 VSS 0.198722f
C19459 DVDD.n16045 VSS 0.081946f
C19460 DVDD.n16046 VSS 0.098809f
C19461 DVDD.t95 VSS 0.167631f
C19462 DVDD.t120 VSS 0.167631f
C19463 DVDD.n16047 VSS 0.335261f
C19464 DVDD.n16048 VSS 0.081946f
C19465 DVDD.n16049 VSS 0.099098f
C19466 DVDD.n16050 VSS 0.198298f
C19467 DVDD.n16051 VSS 0.117632f
C19468 DVDD.n16061 VSS 0.123789f
C19469 DVDD.n16062 VSS 0.098809f
C19470 DVDD.t88 VSS 0.167631f
C19471 DVDD.t150 VSS 0.167631f
C19472 DVDD.n16063 VSS 0.335261f
C19473 DVDD.n16064 VSS 0.099098f
C19474 DVDD.n16065 VSS 0.198298f
C19475 DVDD.n16066 VSS 0.107058f
C19476 DVDD.n16067 VSS 0.137328f
C19477 DVDD.n16068 VSS 0.112345f
C19478 DVDD.n16069 VSS 0.198298f
C19479 DVDD.n16070 VSS 0.099098f
C19480 DVDD.n16071 VSS 0.081946f
C19481 DVDD.n16075 VSS 0.11992f
C19482 DVDD.n16081 VSS 0.131525f
C19483 DVDD.n16082 VSS 0.112345f
C19484 DVDD.n16083 VSS 0.125723f
C19485 DVDD.n16084 VSS 0.107058f
C19486 DVDD.n16085 VSS 0.137328f
C19487 DVDD.n16086 VSS 0.11992f
C19488 DVDD.n16087 VSS 0.274656f
C19489 DVDD.n16088 VSS 0.274656f
C19490 DVDD.n16089 VSS 0.274656f
C19491 DVDD.n16090 VSS 0.274656f
C19492 DVDD.n16091 VSS 0.274656f
C19493 DVDD.n16092 VSS 0.201157f
C19494 DVDD.n16093 VSS 0.274656f
C19495 DVDD.n16094 VSS 0.274656f
C19496 DVDD.n16095 VSS 0.274656f
C19497 DVDD.n16096 VSS 0.274656f
C19498 DVDD.n16097 VSS 0.274656f
C19499 DVDD.n16098 VSS 0.274656f
C19500 DVDD.n16099 VSS 0.274656f
C19501 DVDD.n16100 VSS 0.274656f
C19502 DVDD.n16101 VSS 0.274656f
C19503 DVDD.n16102 VSS 0.205025f
C19504 DVDD.n16113 VSS 0.137328f
C19505 DVDD.n16114 VSS 0.11992f
C19506 DVDD.n16115 VSS 0.274656f
C19507 DVDD.n16116 VSS 0.11992f
C19508 DVDD.n16117 VSS 0.274656f
C19509 DVDD.n16118 VSS 0.11992f
C19510 DVDD.n16119 VSS 0.274656f
C19511 DVDD.n16120 VSS 0.274656f
C19512 DVDD.n16121 VSS 0.274656f
C19513 DVDD.n16122 VSS 0.274656f
C19514 DVDD.n16123 VSS 0.11992f
C19515 DVDD.n16124 VSS 0.274656f
C19516 DVDD.n16125 VSS 0.11992f
C19517 DVDD.n16126 VSS 0.274656f
C19518 DVDD.n16127 VSS 0.11992f
C19519 DVDD.n16128 VSS 0.274656f
C19520 DVDD.n16129 VSS 0.274656f
C19521 DVDD.n16130 VSS 0.274656f
C19522 DVDD.n16131 VSS 0.168275f
C19523 DVDD.n16132 VSS 0.11992f
C19524 DVDD.n16133 VSS 0.168275f
C19525 DVDD.n16134 VSS 0.330748f
C19526 DVDD.n16135 VSS 0.11992f
C19527 DVDD.n16136 VSS 0.243709f
C19528 DVDD.n16137 VSS 0.243709f
C19529 DVDD.n16138 VSS 0.274656f
C19530 DVDD.n16139 VSS 0.274656f
C19531 DVDD.n16140 VSS 0.11992f
C19532 DVDD.n16141 VSS 0.11992f
C19533 DVDD.n16142 VSS 0.137328f
C19534 DVDD.n16143 VSS 0.107058f
C19535 DVDD.n16144 VSS 0.137328f
C19536 DVDD.n16145 VSS 0.11992f
C19537 DVDD.n16146 VSS 0.274656f
C19538 DVDD.n16147 VSS 0.274656f
C19539 DVDD.n16148 VSS 0.274656f
C19540 DVDD.n16149 VSS 0.274656f
C19541 DVDD.n16150 VSS 0.274656f
C19542 DVDD.n16151 VSS 0.274656f
C19543 DVDD.n16152 VSS 0.274656f
C19544 DVDD.n16153 VSS 0.274656f
C19545 DVDD.n16154 VSS 0.162473f
C19546 DVDD.n16155 VSS 0.274656f
C19547 DVDD.n16156 VSS 0.11992f
C19548 DVDD.n16157 VSS 0.274656f
C19549 DVDD.n16158 VSS 0.274656f
C19550 DVDD.n16159 VSS 0.274656f
C19551 DVDD.n16160 VSS 0.274656f
C19552 DVDD.n16161 VSS 0.11992f
C19553 DVDD.n16162 VSS 0.274656f
C19554 DVDD.n16163 VSS 0.11992f
C19555 DVDD.n16164 VSS 0.274656f
C19556 DVDD.n16165 VSS 0.11992f
C19557 DVDD.n16166 VSS 0.274656f
C19558 DVDD.n16167 VSS 0.274656f
C19559 DVDD.n16168 VSS 0.274656f
C19560 DVDD.n16169 VSS 0.274656f
C19561 DVDD.n16170 VSS 0.11992f
C19562 DVDD.n16171 VSS 0.274656f
C19563 DVDD.n16172 VSS 0.11992f
C19564 DVDD.n16173 VSS 0.274656f
C19565 DVDD.n16174 VSS 0.11992f
C19566 DVDD.n16175 VSS 0.274656f
C19567 DVDD.n16176 VSS 0.274656f
C19568 DVDD.n16177 VSS 0.274656f
C19569 DVDD.n16178 VSS 0.274656f
C19570 DVDD.n16179 VSS 0.274656f
C19571 DVDD.n16180 VSS 0.11992f
C19572 DVDD.n16181 VSS 0.11992f
C19573 DVDD.n16182 VSS 0.137328f
C19574 DVDD.n16183 VSS 0.107058f
C19575 DVDD.n16184 VSS 0.137328f
C19576 DVDD.n16185 VSS 0.11992f
C19577 DVDD.n16186 VSS 0.274656f
C19578 DVDD.n16187 VSS 0.274656f
C19579 DVDD.n16188 VSS 0.274656f
C19580 DVDD.n16189 VSS 0.330748f
C19581 DVDD.n16190 VSS 0.160538f
C19582 DVDD.n16191 VSS 0.274656f
C19583 DVDD.n16192 VSS 0.274656f
C19584 DVDD.n16193 VSS 0.274656f
C19585 DVDD.n16194 VSS 0.160538f
C19586 DVDD.n16195 VSS 0.330748f
C19587 DVDD.n16196 VSS 0.221466f
C19588 DVDD.n16197 VSS 0.251446f
C19589 DVDD.n16198 VSS 0.251446f
C19590 DVDD.n16199 VSS 0.330748f
C19591 DVDD.n16200 VSS 0.251446f
C19592 DVDD.n16201 VSS 0.274656f
C19593 DVDD.n16202 VSS 0.274656f
C19594 DVDD.n16203 VSS 0.274656f
C19595 DVDD.n16204 VSS 0.274656f
C19596 DVDD.n16205 VSS 0.274656f
C19597 DVDD.n16206 VSS 0.274656f
C19598 DVDD.n16207 VSS 0.274656f
C19599 DVDD.n16208 VSS 0.274656f
C19600 DVDD.n16209 VSS 0.274656f
C19601 DVDD.n16210 VSS 0.247577f
C19602 DVDD.n16211 VSS 0.030947f
C19603 DVDD.n16212 VSS 1.26626f
C19604 DVDD.n16213 VSS 0.745125f
C19605 DVDD.n16214 VSS 0.11992f
C19606 DVDD.n16215 VSS 0.355263f
C19607 DVDD.n16216 VSS 0.11992f
C19608 DVDD.n16217 VSS 0.274656f
C19609 DVDD.n16218 VSS 0.057059f
C19610 DVDD.n16219 VSS 0.164407f
C19611 DVDD.n16220 VSS 0.11992f
C19612 DVDD.n16221 VSS 0.247577f
C19613 DVDD.n16222 VSS 0.11992f
C19614 DVDD.n16223 VSS 0.274656f
C19615 DVDD.n16224 VSS 0.11992f
C19616 DVDD.n16225 VSS 0.274656f
C19617 DVDD.n16226 VSS 0.11992f
C19618 DVDD.n16227 VSS 0.274656f
C19619 DVDD.n16228 VSS 0.11992f
C19620 DVDD.n16229 VSS 0.274656f
C19621 DVDD.n16230 VSS 0.11992f
C19622 DVDD.n16231 VSS 0.274656f
C19623 DVDD.n16232 VSS 0.11992f
C19624 DVDD.n16233 VSS 0.274656f
C19625 DVDD.n16234 VSS 0.11992f
C19626 DVDD.n16235 VSS 0.274656f
C19627 DVDD.n16236 VSS 0.274656f
C19628 DVDD.n16237 VSS 0.274656f
C19629 DVDD.n16238 VSS 0.251446f
C19630 DVDD.n16239 VSS 0.251446f
C19631 DVDD.n16240 VSS 0.524168f
C19632 DVDD.n16241 VSS 0.160538f
C19633 DVDD.n16242 VSS 0.160538f
C19634 DVDD.n16243 VSS 0.274656f
C19635 DVDD.n16244 VSS 0.274656f
C19636 DVDD.n16245 VSS 0.235972f
C19637 DVDD.n16246 VSS 0.137328f
C19638 DVDD.n16247 VSS 0.183717f
C19639 DVDD.n16248 VSS 0.137328f
C19640 DVDD.n16249 VSS 0.162473f
C19641 DVDD.n16250 VSS 0.274656f
C19642 DVDD.n16251 VSS 0.274656f
C19643 DVDD.n16252 VSS 0.274656f
C19644 DVDD.n16253 VSS 0.274656f
C19645 DVDD.n16254 VSS 0.19342f
C19646 DVDD.n16255 VSS 0.137328f
C19647 DVDD.n16256 VSS 0.183717f
C19648 DVDD.n16257 VSS 0.13346f
C19649 DVDD.n16258 VSS 0.11992f
C19650 DVDD.n16259 VSS 0.243709f
C19651 DVDD.n16260 VSS 0.243709f
C19652 DVDD.n16261 VSS 0.524168f
C19653 DVDD.n16262 VSS 0.524168f
C19654 DVDD.n16263 VSS 0.243709f
C19655 DVDD.n16264 VSS 0.274656f
C19656 DVDD.n16265 VSS 0.274656f
C19657 DVDD.n16266 VSS 0.11992f
C19658 DVDD.n16267 VSS 0.11992f
C19659 DVDD.n16268 VSS 0.137328f
C19660 DVDD.n16269 VSS 0.307957f
C19661 DVDD.n16270 VSS 0.137328f
C19662 DVDD.n16271 VSS 0.11992f
C19663 DVDD.n16272 VSS 0.274656f
C19664 DVDD.n16273 VSS 0.274656f
C19665 DVDD.n16274 VSS 0.274656f
C19666 DVDD.n16275 VSS 0.274656f
C19667 DVDD.n16276 VSS 0.274656f
C19668 DVDD.n16277 VSS 0.274656f
C19669 DVDD.n16278 VSS 0.274656f
C19670 DVDD.n16279 VSS 0.274656f
C19671 DVDD.n16280 VSS 0.162473f
C19672 DVDD.n16281 VSS 0.274656f
C19673 DVDD.n16282 VSS 0.11992f
C19674 DVDD.n16283 VSS 0.274656f
C19675 DVDD.n16284 VSS 0.11992f
C19676 DVDD.n16285 VSS 0.274656f
C19677 DVDD.n16286 VSS 0.274656f
C19678 DVDD.n16287 VSS 0.274656f
C19679 DVDD.n16288 VSS 0.274656f
C19680 DVDD.n16289 VSS 0.11992f
C19681 DVDD.n16290 VSS 0.274656f
C19682 DVDD.n16291 VSS 0.11992f
C19683 DVDD.n16292 VSS 0.274656f
C19684 DVDD.n16293 VSS 0.11992f
C19685 DVDD.n16294 VSS 0.274656f
C19686 DVDD.n16295 VSS 0.274656f
C19687 DVDD.n16296 VSS 0.274656f
C19688 DVDD.n16297 VSS 0.274656f
C19689 DVDD.n16298 VSS 0.11992f
C19690 DVDD.n16299 VSS 0.274656f
C19691 DVDD.n16300 VSS 0.11992f
C19692 DVDD.n16301 VSS 0.274656f
C19693 DVDD.n16302 VSS 0.11992f
C19694 DVDD.n16303 VSS 0.274656f
C19695 DVDD.n16304 VSS 0.274656f
C19696 DVDD.n16305 VSS 0.274656f
C19697 DVDD.n16306 VSS 0.274656f
C19698 DVDD.n16307 VSS 0.274656f
C19699 DVDD.n16308 VSS 0.274656f
C19700 DVDD.n16309 VSS 0.274656f
C19701 DVDD.n16310 VSS 0.274656f
C19702 DVDD.n16311 VSS 0.11992f
C19703 DVDD.n16312 VSS 0.137328f
C19704 DVDD.n16313 VSS 0.307957f
C19705 DVDD.n16314 VSS 0.137328f
C19706 DVDD.n16315 VSS 0.235972f
C19707 DVDD.n16316 VSS 0.274656f
C19708 DVDD.n16317 VSS 0.274656f
C19709 DVDD.n16318 VSS 0.160538f
C19710 DVDD.n16319 VSS 0.160538f
C19711 DVDD.n16320 VSS 0.524168f
C19712 DVDD.n16321 VSS 0.251446f
C19713 DVDD.n16322 VSS 0.274656f
C19714 DVDD.n16323 VSS 0.274656f
C19715 DVDD.n16324 VSS 0.274656f
C19716 DVDD.n16325 VSS 0.274656f
C19717 DVDD.n16326 VSS 0.274656f
C19718 DVDD.n16327 VSS 0.274656f
C19719 DVDD.n16328 VSS 0.274656f
C19720 DVDD.n16329 VSS 0.274656f
C19721 DVDD.n16330 VSS 0.274656f
C19722 DVDD.n16331 VSS 0.274656f
C19723 DVDD.n16332 VSS 0.141196f
C19724 DVDD.n16333 VSS 1.26626f
C19725 DVDD.n16334 VSS 0.745125f
C19726 DVDD.n16335 VSS 0.11992f
C19727 DVDD.n16336 VSS 0.355263f
C19728 DVDD.n16337 VSS 0.11992f
C19729 DVDD.n16338 VSS 0.274656f
C19730 DVDD.n16339 VSS 0.057059f
C19731 DVDD.n16340 VSS 0.164407f
C19732 DVDD.n16341 VSS 0.11992f
C19733 DVDD.n16342 VSS 0.247577f
C19734 DVDD.n16343 VSS 0.11992f
C19735 DVDD.n16344 VSS 0.274656f
C19736 DVDD.n16345 VSS 0.11992f
C19737 DVDD.n16346 VSS 0.274656f
C19738 DVDD.n16347 VSS 0.11992f
C19739 DVDD.n16348 VSS 0.274656f
C19740 DVDD.n16349 VSS 0.11992f
C19741 DVDD.n16350 VSS 0.274656f
C19742 DVDD.n16351 VSS 0.11992f
C19743 DVDD.n16352 VSS 0.274656f
C19744 DVDD.n16353 VSS 0.11992f
C19745 DVDD.n16354 VSS 0.274656f
C19746 DVDD.n16355 VSS 0.11992f
C19747 DVDD.n16356 VSS 0.274656f
C19748 DVDD.n16357 VSS 0.274656f
C19749 DVDD.n16358 VSS 0.274656f
C19750 DVDD.n16359 VSS 0.251446f
C19751 DVDD.n16360 VSS 0.251446f
C19752 DVDD.n16361 VSS 0.524168f
C19753 DVDD.n16362 VSS 0.330748f
C19754 DVDD.n16363 VSS 0.160538f
C19755 DVDD.n16364 VSS 0.160538f
C19756 DVDD.n16365 VSS 0.274656f
C19757 DVDD.n16366 VSS 0.274656f
C19758 DVDD.n16367 VSS 0.235972f
C19759 DVDD.n16368 VSS 0.137328f
C19760 DVDD.n16369 VSS 0.071372f
C19761 DVDD.n16370 VSS 0.127657f
C19762 DVDD.n16371 VSS 0.11992f
C19763 DVDD.n16372 VSS 0.274656f
C19764 DVDD.n16373 VSS 0.274656f
C19765 DVDD.n16374 VSS 0.162473f
C19766 DVDD.n16375 VSS 0.274656f
C19767 DVDD.n16376 VSS 0.274656f
C19768 DVDD.n16377 VSS 0.274656f
C19769 DVDD.n16378 VSS 0.274656f
C19770 DVDD.n16379 VSS 0.274656f
C19771 DVDD.n16380 VSS 0.274656f
C19772 DVDD.n16381 VSS 0.11992f
C19773 DVDD.n16390 VSS 0.137328f
C19774 DVDD.n16393 VSS 0.163891f
C19775 DVDD.n16394 VSS 0.137328f
C19776 DVDD.n16395 VSS 0.153317f
C19777 DVDD.n16396 VSS 0.081946f
C19778 DVDD.n16397 VSS 0.063349f
C19779 DVDD.n16398 VSS 0.081946f
C19780 DVDD.n16399 VSS 0.05801f
C19781 DVDD.n16400 VSS -1.41702f
C19782 DVDD.n16401 VSS 5.22944f
C19783 DVDD.n16402 VSS 3.49331f
C19784 DVDD.n16403 VSS 5.22944f
C19785 DVDD.n16404 VSS -1.41702f
C19786 DVDD.n16406 VSS 0.05801f
C19787 DVDD.n16409 VSS 0.025624f
C19788 DVDD.n16412 VSS 0.025624f
C19789 DVDD.n16415 VSS 0.025624f
C19790 DVDD.n16418 VSS 0.025624f
C19791 DVDD.n16421 VSS 0.025624f
C19792 DVDD.n16424 VSS 0.025624f
C19793 DVDD.n16426 VSS 0.025624f
C19794 DVDD.n16428 VSS 0.025624f
C19795 DVDD.n16429 VSS 0.025624f
C19796 DVDD.n16431 VSS 0.794343f
C19797 DVDD.n16432 VSS 0.063349f
C19798 DVDD.n16433 VSS 0.063349f
C19799 DVDD.n16435 VSS 0.025624f
C19800 DVDD.n16437 VSS 0.025624f
C19801 DVDD.n16439 VSS 0.025624f
C19802 DVDD.n16441 VSS 0.025624f
C19803 DVDD.n16443 VSS 0.025624f
C19804 DVDD.n16445 VSS 0.025624f
C19805 DVDD.n16447 VSS 0.025624f
C19806 DVDD.n16449 VSS 0.794343f
C19807 DVDD.n16450 VSS 0.098464f
C19808 DVDD.n16451 VSS 0.468543f
C19809 DVDD.n16452 VSS 0.423753f
C19810 DVDD.n16453 VSS 0.034514f
C19811 DVDD.n16454 VSS 0.050915f
C19812 DVDD.n16455 VSS 0.033945f
C19813 DVDD.n16456 VSS 0.019729f
C19814 DVDD.n16457 VSS 0.028497f
C19815 DVDD.n16458 VSS 0.031128f
C19816 DVDD.n16459 VSS 0.031128f
C19817 DVDD.n16460 VSS 0.031128f
C19818 DVDD.n16461 VSS 0.031128f
C19819 DVDD.n16463 VSS 0.031128f
C19820 DVDD.n16464 VSS 0.031128f
C19821 DVDD.n16465 VSS 0.031128f
C19822 DVDD.n16467 VSS 0.031128f
C19823 DVDD.n16468 VSS 0.031128f
C19824 DVDD.n16469 VSS 0.031128f
C19825 DVDD.n16470 VSS 0.031128f
C19826 DVDD.n16471 VSS 0.031128f
C19827 DVDD.n16472 VSS 0.031128f
C19828 DVDD.n16473 VSS 0.031128f
C19829 DVDD.n16475 VSS 0.031128f
C19830 DVDD.n16476 VSS 0.031128f
C19831 DVDD.n16477 VSS 0.031128f
C19832 DVDD.n16479 VSS 0.031128f
C19833 DVDD.n16480 VSS 0.031128f
C19834 DVDD.n16481 VSS 0.031128f
C19835 DVDD.n16482 VSS 0.031128f
C19836 DVDD.n16483 VSS 0.031128f
C19837 DVDD.n16484 VSS 0.031128f
C19838 DVDD.n16485 VSS 0.031128f
C19839 DVDD.n16487 VSS 0.031128f
C19840 DVDD.n16488 VSS 0.031128f
C19841 DVDD.n16489 VSS 0.031128f
C19842 DVDD.n16491 VSS 0.031128f
C19843 DVDD.n16492 VSS 0.031128f
C19844 DVDD.n16493 VSS 0.031128f
C19845 DVDD.n16494 VSS 0.031128f
C19846 DVDD.n16495 VSS 0.031128f
C19847 DVDD.n16496 VSS 0.031128f
C19848 DVDD.n16497 VSS 0.031128f
C19849 DVDD.n16499 VSS 0.031128f
C19850 DVDD.n16500 VSS 0.031128f
C19851 DVDD.n16501 VSS 0.031128f
C19852 DVDD.n16503 VSS 0.031128f
C19853 DVDD.n16504 VSS 0.031128f
C19854 DVDD.n16505 VSS 0.031128f
C19855 DVDD.n16506 VSS 0.031128f
C19856 DVDD.n16507 VSS 0.031128f
C19857 DVDD.n16508 VSS 0.031128f
C19858 DVDD.n16509 VSS 0.031128f
C19859 DVDD.n16511 VSS 0.031128f
C19860 DVDD.n16512 VSS 0.031128f
C19861 DVDD.n16513 VSS 0.031128f
C19862 DVDD.n16515 VSS 0.031128f
C19863 DVDD.n16516 VSS 0.031128f
C19864 DVDD.n16517 VSS 0.031128f
C19865 DVDD.n16518 VSS 0.031128f
C19866 DVDD.n16519 VSS 0.031128f
C19867 DVDD.n16520 VSS 0.031128f
C19868 DVDD.n16521 VSS 0.031128f
C19869 DVDD.n16523 VSS 0.031128f
C19870 DVDD.n16524 VSS 0.031128f
C19871 DVDD.n16525 VSS 0.031128f
C19872 DVDD.n16527 VSS 0.031128f
C19873 DVDD.n16528 VSS 0.031128f
C19874 DVDD.n16529 VSS 0.031128f
C19875 DVDD.n16530 VSS 0.031128f
C19876 DVDD.n16531 VSS 0.031128f
C19877 DVDD.n16532 VSS 0.031128f
C19878 DVDD.n16533 VSS 0.031128f
C19879 DVDD.n16535 VSS 0.031128f
C19880 DVDD.n16536 VSS 0.031128f
C19881 DVDD.n16537 VSS 0.031128f
C19882 DVDD.n16539 VSS 0.031128f
C19883 DVDD.n16540 VSS 0.031128f
C19884 DVDD.n16541 VSS 0.031128f
C19885 DVDD.n16542 VSS 0.031128f
C19886 DVDD.n16543 VSS 0.031128f
C19887 DVDD.n16544 VSS 0.031128f
C19888 DVDD.n16545 VSS 0.031128f
C19889 DVDD.n16547 VSS 0.031128f
C19890 DVDD.n16548 VSS 0.031128f
C19891 DVDD.n16549 VSS 0.031128f
C19892 DVDD.n16551 VSS 0.031128f
C19893 DVDD.n16552 VSS 0.031128f
C19894 DVDD.n16553 VSS 0.031128f
C19895 DVDD.n16554 VSS 0.031128f
C19896 DVDD.n16555 VSS 0.031128f
C19897 DVDD.n16556 VSS 0.031128f
C19898 DVDD.n16557 VSS 0.031128f
C19899 DVDD.n16559 VSS 0.031128f
C19900 DVDD.n16560 VSS 0.031128f
C19901 DVDD.n16561 VSS 0.031128f
C19902 DVDD.n16563 VSS 0.031128f
C19903 DVDD.n16564 VSS 0.031128f
C19904 DVDD.n16565 VSS 0.031128f
C19905 DVDD.n16566 VSS 0.031128f
C19906 DVDD.n16567 VSS 0.031128f
C19907 DVDD.n16568 VSS 0.031128f
C19908 DVDD.n16569 VSS 0.031128f
C19909 DVDD.n16571 VSS 0.031128f
C19910 DVDD.n16572 VSS 0.031128f
C19911 DVDD.n16573 VSS 0.031128f
C19912 DVDD.n16575 VSS 0.031128f
C19913 DVDD.n16576 VSS 0.031128f
C19914 DVDD.n16577 VSS 0.031128f
C19915 DVDD.n16578 VSS 0.031128f
C19916 DVDD.n16579 VSS 0.031128f
C19917 DVDD.n16580 VSS 0.031128f
C19918 DVDD.n16581 VSS 0.031128f
C19919 DVDD.n16583 VSS 0.031128f
C19920 DVDD.n16584 VSS 0.031128f
C19921 DVDD.n16585 VSS 0.031128f
C19922 DVDD.n16587 VSS 0.031128f
C19923 DVDD.n16588 VSS 0.031128f
C19924 DVDD.n16589 VSS 0.031128f
C19925 DVDD.n16590 VSS 0.031128f
C19926 DVDD.n16591 VSS 0.031128f
C19927 DVDD.n16592 VSS 0.031128f
C19928 DVDD.n16593 VSS 0.031128f
C19929 DVDD.n16595 VSS 0.031128f
C19930 DVDD.n16596 VSS 0.031128f
C19931 DVDD.n16597 VSS 0.031128f
C19932 DVDD.n16599 VSS 0.031128f
C19933 DVDD.n16600 VSS 0.031128f
C19934 DVDD.n16601 VSS 0.031128f
C19935 DVDD.n16602 VSS 0.031128f
C19936 DVDD.n16603 VSS 0.031128f
C19937 DVDD.n16604 VSS 0.031128f
C19938 DVDD.n16605 VSS 0.031128f
C19939 DVDD.n16607 VSS 0.031128f
C19940 DVDD.n16608 VSS 0.031128f
C19941 DVDD.n16609 VSS 0.031128f
C19942 DVDD.n16611 VSS 0.031128f
C19943 DVDD.n16612 VSS 0.031128f
C19944 DVDD.n16613 VSS 0.031128f
C19945 DVDD.n16614 VSS 0.031128f
C19946 DVDD.n16615 VSS 0.031128f
C19947 DVDD.n16616 VSS 0.031128f
C19948 DVDD.n16617 VSS 0.031128f
C19949 DVDD.n16619 VSS 0.031128f
C19950 DVDD.n16620 VSS 0.031128f
C19951 DVDD.n16621 VSS 0.031128f
C19952 DVDD.n16623 VSS 0.031128f
C19953 DVDD.n16624 VSS 0.031128f
C19954 DVDD.n16625 VSS 0.031128f
C19955 DVDD.n16626 VSS 0.031128f
C19956 DVDD.n16627 VSS 0.031128f
C19957 DVDD.n16628 VSS 0.031128f
C19958 DVDD.n16629 VSS 0.031128f
C19959 DVDD.n16631 VSS 0.031128f
C19960 DVDD.n16632 VSS 0.031128f
C19961 DVDD.n16633 VSS 0.031128f
C19962 DVDD.n16635 VSS 0.031128f
C19963 DVDD.n16636 VSS 0.031128f
C19964 DVDD.n16637 VSS 0.031128f
C19965 DVDD.n16638 VSS 0.031128f
C19966 DVDD.n16639 VSS 0.031128f
C19967 DVDD.n16640 VSS 0.031128f
C19968 DVDD.n16641 VSS 0.031128f
C19969 DVDD.n16643 VSS 0.031128f
C19970 DVDD.n16644 VSS 0.031128f
C19971 DVDD.n16645 VSS 0.031128f
C19972 DVDD.n16647 VSS 0.031128f
C19973 DVDD.n16648 VSS 0.031128f
C19974 DVDD.n16649 VSS 0.031128f
C19975 DVDD.n16650 VSS 0.031128f
C19976 DVDD.n16651 VSS 0.031128f
C19977 DVDD.n16652 VSS 0.031128f
C19978 DVDD.n16653 VSS 0.031128f
C19979 DVDD.n16655 VSS 0.031128f
C19980 DVDD.n16656 VSS 0.031128f
C19981 DVDD.n16657 VSS 0.031128f
C19982 DVDD.n16659 VSS 0.031128f
C19983 DVDD.n16660 VSS 0.031128f
C19984 DVDD.n16661 VSS 0.031128f
C19985 DVDD.n16662 VSS 0.031128f
C19986 DVDD.n16663 VSS 0.031128f
C19987 DVDD.n16664 VSS 0.031128f
C19988 DVDD.n16665 VSS 0.031128f
C19989 DVDD.n16667 VSS 0.031128f
C19990 DVDD.n16668 VSS 0.031128f
C19991 DVDD.n16669 VSS 0.031128f
C19992 DVDD.n16671 VSS 0.031128f
C19993 DVDD.n16672 VSS 0.031128f
C19994 DVDD.n16673 VSS 0.031128f
C19995 DVDD.n16674 VSS 0.031128f
C19996 DVDD.n16675 VSS 0.031128f
C19997 DVDD.n16676 VSS 0.031128f
C19998 DVDD.n16677 VSS 0.031128f
C19999 DVDD.n16679 VSS 0.031128f
C20000 DVDD.n16680 VSS 0.031128f
C20001 DVDD.n16681 VSS 0.031128f
C20002 DVDD.n16683 VSS 0.031128f
C20003 DVDD.n16684 VSS 0.031128f
C20004 DVDD.n16685 VSS 0.031128f
C20005 DVDD.n16686 VSS 0.031128f
C20006 DVDD.n16687 VSS 0.031128f
C20007 DVDD.n16688 VSS 0.031128f
C20008 DVDD.n16689 VSS 0.031128f
C20009 DVDD.n16691 VSS 0.031128f
C20010 DVDD.n16692 VSS 0.031128f
C20011 DVDD.n16693 VSS 0.031128f
C20012 DVDD.n16695 VSS 0.031128f
C20013 DVDD.n16696 VSS 0.031128f
C20014 DVDD.n16697 VSS 0.031128f
C20015 DVDD.n16698 VSS 0.031128f
C20016 DVDD.n16699 VSS 0.031128f
C20017 DVDD.n16700 VSS 0.031128f
C20018 DVDD.n16701 VSS 0.031128f
C20019 DVDD.n16703 VSS 0.019729f
C20020 DVDD.n16704 VSS 0.450653f
C20021 DVDD.n16705 VSS 0.446441f
C20022 DVDD.n16706 VSS 0.023771f
C20023 DVDD.n16707 VSS 0.023771f
C20024 DVDD.n16708 VSS 0.02076f
C20025 DVDD.n16709 VSS 0.028833f
C20026 DVDD.n16710 VSS 0.034171f
C20027 DVDD.n16711 VSS 0.035718f
C20028 DVDD.n16712 VSS 0.040897f
C20029 DVDD.n16713 VSS 0.040897f
C20030 DVDD.n16714 VSS 0.505405f
C20031 DVDD.n16715 VSS 0.598063f
C20032 DVDD.n16716 VSS 0.05956f
C20033 DVDD.n16717 VSS 0.045151f
C20034 DVDD.n16718 VSS 0.045151f
C20035 DVDD.n16719 VSS 0.040302f
C20036 DVDD.n16720 VSS 0.039516f
C20037 DVDD.n16721 VSS 0.046305f
C20038 DVDD.n16722 VSS 0.053165f
C20039 DVDD.n16723 VSS 0.039445f
C20040 DVDD.n16724 VSS 0.04419f
C20041 DVDD.n16725 VSS 0.04419f
C20042 DVDD.n16726 VSS 0.282185f
C20043 DVDD.n16727 VSS 0.522252f
C20044 DVDD.n16728 VSS 0.021999f
C20045 DVDD.n16729 VSS 0.021999f
C20046 DVDD.n16730 VSS 0.019213f
C20047 DVDD.n16731 VSS 0.036621f
C20048 DVDD.n16732 VSS 0.032366f
C20049 DVDD.n16733 VSS 0.037059f
C20050 DVDD.n16734 VSS 0.037059f
C20051 DVDD.n16735 VSS 0.522252f
C20052 DVDD.n16736 VSS 0.160045f
C20053 DVDD.n16737 VSS 0.051875f
C20054 DVDD.n16738 VSS 0.033945f
C20055 DVDD.n16739 VSS 0.037465f
C20056 DVDD.n16740 VSS 0.052307f
C20057 DVDD.n16741 VSS 0.053165f
C20058 DVDD.n16742 VSS 0.033442f
C20059 DVDD.n16743 VSS 0.037465f
C20060 DVDD.n16744 VSS 0.033945f
C20061 DVDD.n16745 VSS 0.019729f
C20062 DVDD.n16746 VSS 0.028497f
C20063 DVDD.n16747 VSS 0.031128f
C20064 DVDD.n16748 VSS 0.031128f
C20065 DVDD.n16749 VSS 0.031128f
C20066 DVDD.n16750 VSS 0.031128f
C20067 DVDD.n16752 VSS 0.031128f
C20068 DVDD.n16753 VSS 0.031128f
C20069 DVDD.n16754 VSS 0.031128f
C20070 DVDD.n16756 VSS 0.031128f
C20071 DVDD.n16757 VSS 0.031128f
C20072 DVDD.n16758 VSS 0.031128f
C20073 DVDD.n16759 VSS 0.031128f
C20074 DVDD.n16760 VSS 0.031128f
C20075 DVDD.n16761 VSS 0.031128f
C20076 DVDD.n16762 VSS 0.031128f
C20077 DVDD.n16764 VSS 0.031128f
C20078 DVDD.n16765 VSS 0.031128f
C20079 DVDD.n16766 VSS 0.031128f
C20080 DVDD.n16768 VSS 0.031128f
C20081 DVDD.n16769 VSS 0.031128f
C20082 DVDD.n16770 VSS 0.031128f
C20083 DVDD.n16771 VSS 0.031128f
C20084 DVDD.n16772 VSS 0.031128f
C20085 DVDD.n16773 VSS 0.031128f
C20086 DVDD.n16774 VSS 0.031128f
C20087 DVDD.n16776 VSS 0.031128f
C20088 DVDD.n16777 VSS 0.031128f
C20089 DVDD.n16778 VSS 0.031128f
C20090 DVDD.n16780 VSS 0.031128f
C20091 DVDD.n16781 VSS 0.031128f
C20092 DVDD.n16782 VSS 0.031128f
C20093 DVDD.n16783 VSS 0.031128f
C20094 DVDD.n16784 VSS 0.031128f
C20095 DVDD.n16785 VSS 0.031128f
C20096 DVDD.n16786 VSS 0.031128f
C20097 DVDD.n16788 VSS 0.031128f
C20098 DVDD.n16789 VSS 0.031128f
C20099 DVDD.n16790 VSS 0.031128f
C20100 DVDD.n16792 VSS 0.031128f
C20101 DVDD.n16793 VSS 0.031128f
C20102 DVDD.n16794 VSS 0.031128f
C20103 DVDD.n16795 VSS 0.031128f
C20104 DVDD.n16796 VSS 0.031128f
C20105 DVDD.n16797 VSS 0.031128f
C20106 DVDD.n16798 VSS 0.031128f
C20107 DVDD.n16800 VSS 0.031128f
C20108 DVDD.n16801 VSS 0.031128f
C20109 DVDD.n16802 VSS 0.031128f
C20110 DVDD.n16804 VSS 0.031128f
C20111 DVDD.n16805 VSS 0.031128f
C20112 DVDD.n16806 VSS 0.031128f
C20113 DVDD.n16807 VSS 0.031128f
C20114 DVDD.n16808 VSS 0.031128f
C20115 DVDD.n16809 VSS 0.031128f
C20116 DVDD.n16810 VSS 0.031128f
C20117 DVDD.n16812 VSS 0.031128f
C20118 DVDD.n16813 VSS 0.031128f
C20119 DVDD.n16814 VSS 0.031128f
C20120 DVDD.n16816 VSS 0.031128f
C20121 DVDD.n16817 VSS 0.031128f
C20122 DVDD.n16818 VSS 0.031128f
C20123 DVDD.n16819 VSS 0.031128f
C20124 DVDD.n16820 VSS 0.031128f
C20125 DVDD.n16821 VSS 0.031128f
C20126 DVDD.n16822 VSS 0.031128f
C20127 DVDD.n16824 VSS 0.031128f
C20128 DVDD.n16825 VSS 0.031128f
C20129 DVDD.n16826 VSS 0.031128f
C20130 DVDD.n16828 VSS 0.031128f
C20131 DVDD.n16829 VSS 0.031128f
C20132 DVDD.n16830 VSS 0.031128f
C20133 DVDD.n16831 VSS 0.031128f
C20134 DVDD.n16832 VSS 0.031128f
C20135 DVDD.n16833 VSS 0.031128f
C20136 DVDD.n16834 VSS 0.031128f
C20137 DVDD.n16836 VSS 0.031128f
C20138 DVDD.n16837 VSS 0.031128f
C20139 DVDD.n16838 VSS 0.031128f
C20140 DVDD.n16840 VSS 0.031128f
C20141 DVDD.n16841 VSS 0.031128f
C20142 DVDD.n16842 VSS 0.031128f
C20143 DVDD.n16843 VSS 0.031128f
C20144 DVDD.n16844 VSS 0.031128f
C20145 DVDD.n16845 VSS 0.031128f
C20146 DVDD.n16846 VSS 0.031128f
C20147 DVDD.n16848 VSS 0.031128f
C20148 DVDD.n16849 VSS 0.031128f
C20149 DVDD.n16850 VSS 0.031128f
C20150 DVDD.n16852 VSS 0.031128f
C20151 DVDD.n16853 VSS 0.031128f
C20152 DVDD.n16854 VSS 0.031128f
C20153 DVDD.n16855 VSS 0.031128f
C20154 DVDD.n16856 VSS 0.031128f
C20155 DVDD.n16857 VSS 0.031128f
C20156 DVDD.n16858 VSS 0.031128f
C20157 DVDD.n16860 VSS 0.031128f
C20158 DVDD.n16861 VSS 0.031128f
C20159 DVDD.n16862 VSS 0.031128f
C20160 DVDD.n16864 VSS 0.031128f
C20161 DVDD.n16865 VSS 0.031128f
C20162 DVDD.n16866 VSS 0.031128f
C20163 DVDD.n16867 VSS 0.031128f
C20164 DVDD.n16868 VSS 0.031128f
C20165 DVDD.n16869 VSS 0.031128f
C20166 DVDD.n16870 VSS 0.031128f
C20167 DVDD.n16872 VSS 0.031128f
C20168 DVDD.n16873 VSS 0.031128f
C20169 DVDD.n16874 VSS 0.031128f
C20170 DVDD.n16876 VSS 0.031128f
C20171 DVDD.n16877 VSS 0.031128f
C20172 DVDD.n16878 VSS 0.031128f
C20173 DVDD.n16879 VSS 0.031128f
C20174 DVDD.n16880 VSS 0.031128f
C20175 DVDD.n16881 VSS 0.031128f
C20176 DVDD.n16882 VSS 0.031128f
C20177 DVDD.n16884 VSS 0.031128f
C20178 DVDD.n16885 VSS 0.031128f
C20179 DVDD.n16886 VSS 0.031128f
C20180 DVDD.n16888 VSS 0.031128f
C20181 DVDD.n16889 VSS 0.031128f
C20182 DVDD.n16890 VSS 0.031128f
C20183 DVDD.n16891 VSS 0.031128f
C20184 DVDD.n16892 VSS 0.031128f
C20185 DVDD.n16893 VSS 0.031128f
C20186 DVDD.n16894 VSS 0.031128f
C20187 DVDD.n16896 VSS 0.031128f
C20188 DVDD.n16897 VSS 0.031128f
C20189 DVDD.n16898 VSS 0.031128f
C20190 DVDD.n16900 VSS 0.031128f
C20191 DVDD.n16901 VSS 0.031128f
C20192 DVDD.n16902 VSS 0.031128f
C20193 DVDD.n16903 VSS 0.031128f
C20194 DVDD.n16904 VSS 0.031128f
C20195 DVDD.n16905 VSS 0.031128f
C20196 DVDD.n16906 VSS 0.031128f
C20197 DVDD.n16908 VSS 0.031128f
C20198 DVDD.n16909 VSS 0.031128f
C20199 DVDD.n16910 VSS 0.031128f
C20200 DVDD.n16912 VSS 0.031128f
C20201 DVDD.n16913 VSS 0.031128f
C20202 DVDD.n16914 VSS 0.031128f
C20203 DVDD.n16915 VSS 0.031128f
C20204 DVDD.n16916 VSS 0.031128f
C20205 DVDD.n16917 VSS 0.031128f
C20206 DVDD.n16918 VSS 0.031128f
C20207 DVDD.n16920 VSS 0.031128f
C20208 DVDD.n16921 VSS 0.031128f
C20209 DVDD.n16922 VSS 0.031128f
C20210 DVDD.n16924 VSS 0.031128f
C20211 DVDD.n16925 VSS 0.031128f
C20212 DVDD.n16926 VSS 0.031128f
C20213 DVDD.n16927 VSS 0.031128f
C20214 DVDD.n16928 VSS 0.031128f
C20215 DVDD.n16929 VSS 0.031128f
C20216 DVDD.n16930 VSS 0.031128f
C20217 DVDD.n16932 VSS 0.031128f
C20218 DVDD.n16933 VSS 0.031128f
C20219 DVDD.n16934 VSS 0.031128f
C20220 DVDD.n16936 VSS 0.031128f
C20221 DVDD.n16937 VSS 0.031128f
C20222 DVDD.n16938 VSS 0.031128f
C20223 DVDD.n16939 VSS 0.031128f
C20224 DVDD.n16940 VSS 0.031128f
C20225 DVDD.n16941 VSS 0.031128f
C20226 DVDD.n16942 VSS 0.031128f
C20227 DVDD.n16944 VSS 0.031128f
C20228 DVDD.n16945 VSS 0.031128f
C20229 DVDD.n16946 VSS 0.031128f
C20230 DVDD.n16948 VSS 0.031128f
C20231 DVDD.n16949 VSS 0.031128f
C20232 DVDD.n16950 VSS 0.031128f
C20233 DVDD.n16951 VSS 0.031128f
C20234 DVDD.n16952 VSS 0.031128f
C20235 DVDD.n16953 VSS 0.031128f
C20236 DVDD.n16954 VSS 0.031128f
C20237 DVDD.n16956 VSS 0.031128f
C20238 DVDD.n16957 VSS 0.031128f
C20239 DVDD.n16958 VSS 0.031128f
C20240 DVDD.n16960 VSS 0.031128f
C20241 DVDD.n16961 VSS 0.031128f
C20242 DVDD.n16962 VSS 0.031128f
C20243 DVDD.n16963 VSS 0.031128f
C20244 DVDD.n16964 VSS 0.031128f
C20245 DVDD.n16965 VSS 0.031128f
C20246 DVDD.n16966 VSS 0.031128f
C20247 DVDD.n16968 VSS 0.031128f
C20248 DVDD.n16969 VSS 0.031128f
C20249 DVDD.n16970 VSS 0.031128f
C20250 DVDD.n16972 VSS 0.031128f
C20251 DVDD.n16973 VSS 0.031128f
C20252 DVDD.n16974 VSS 0.031128f
C20253 DVDD.n16975 VSS 0.031128f
C20254 DVDD.n16976 VSS 0.031128f
C20255 DVDD.n16977 VSS 0.031128f
C20256 DVDD.n16978 VSS 0.031128f
C20257 DVDD.n16980 VSS 0.031128f
C20258 DVDD.n16981 VSS 0.031128f
C20259 DVDD.n16982 VSS 0.031128f
C20260 DVDD.n16984 VSS 0.031128f
C20261 DVDD.n16985 VSS 0.031128f
C20262 DVDD.n16986 VSS 0.031128f
C20263 DVDD.n16987 VSS 0.031128f
C20264 DVDD.n16988 VSS 0.026086f
C20265 DVDD.n16989 VSS 0.031128f
C20266 DVDD.n16990 VSS 0.031128f
C20267 DVDD.n16991 VSS 0.031128f
C20268 DVDD.n16993 VSS 0.019729f
C20269 DVDD.n16994 VSS 0.518041f
C20270 DVDD.n16995 VSS 0.164257f
C20271 DVDD.n16996 VSS 0.025838f
C20272 DVDD.n16997 VSS 0.025838f
C20273 DVDD.n16998 VSS 0.022566f
C20274 DVDD.n16999 VSS 0.036621f
C20275 DVDD.n17000 VSS 0.029013f
C20276 DVDD.n17001 VSS 0.03322f
C20277 DVDD.n17002 VSS 0.03322f
C20278 DVDD.n17003 VSS 0.193738f
C20279 DVDD.n17004 VSS 0.598063f
C20280 DVDD.n17005 VSS 0.0586f
C20281 DVDD.n17006 VSS 0.033945f
C20282 DVDD.n17007 VSS 0.05956f
C20283 DVDD.n17008 VSS 0.030741f
C20284 DVDD.n17009 VSS 0.053165f
C20285 DVDD.n17010 VSS 0.02744f
C20286 DVDD.n17011 VSS 0.030741f
C20287 DVDD.n17012 VSS 0.033945f
C20288 DVDD.n17013 VSS 0.019729f
C20289 DVDD.n17014 VSS 0.028497f
C20290 DVDD.n17015 VSS 0.031128f
C20291 DVDD.n17016 VSS 0.031128f
C20292 DVDD.n17017 VSS 0.031128f
C20293 DVDD.n17018 VSS 0.031128f
C20294 DVDD.n17020 VSS 0.031128f
C20295 DVDD.n17021 VSS 0.031128f
C20296 DVDD.n17022 VSS 0.031128f
C20297 DVDD.n17024 VSS 0.031128f
C20298 DVDD.n17025 VSS 0.031128f
C20299 DVDD.n17026 VSS 0.031128f
C20300 DVDD.n17027 VSS 0.031128f
C20301 DVDD.n17028 VSS 0.031128f
C20302 DVDD.n17029 VSS 0.031128f
C20303 DVDD.n17030 VSS 0.031128f
C20304 DVDD.n17032 VSS 0.031128f
C20305 DVDD.n17033 VSS 0.031128f
C20306 DVDD.n17034 VSS 0.031128f
C20307 DVDD.n17036 VSS 0.031128f
C20308 DVDD.n17037 VSS 0.031128f
C20309 DVDD.n17038 VSS 0.031128f
C20310 DVDD.n17039 VSS 0.031128f
C20311 DVDD.n17040 VSS 0.031128f
C20312 DVDD.n17041 VSS 0.031128f
C20313 DVDD.n17042 VSS 0.031128f
C20314 DVDD.n17044 VSS 0.031128f
C20315 DVDD.n17045 VSS 0.031128f
C20316 DVDD.n17046 VSS 0.031128f
C20317 DVDD.n17048 VSS 0.031128f
C20318 DVDD.n17049 VSS 0.031128f
C20319 DVDD.n17050 VSS 0.031128f
C20320 DVDD.n17051 VSS 0.031128f
C20321 DVDD.n17052 VSS 0.031128f
C20322 DVDD.n17053 VSS 0.031128f
C20323 DVDD.n17054 VSS 0.031128f
C20324 DVDD.n17056 VSS 0.031128f
C20325 DVDD.n17057 VSS 0.031128f
C20326 DVDD.n17058 VSS 0.031128f
C20327 DVDD.n17060 VSS 0.031128f
C20328 DVDD.n17061 VSS 0.031128f
C20329 DVDD.n17062 VSS 0.031128f
C20330 DVDD.n17063 VSS 0.031128f
C20331 DVDD.n17064 VSS 0.031128f
C20332 DVDD.n17065 VSS 0.031128f
C20333 DVDD.n17066 VSS 0.031128f
C20334 DVDD.n17068 VSS 0.031128f
C20335 DVDD.n17069 VSS 0.031128f
C20336 DVDD.n17070 VSS 0.031128f
C20337 DVDD.n17072 VSS 0.031128f
C20338 DVDD.n17073 VSS 0.031128f
C20339 DVDD.n17074 VSS 0.031128f
C20340 DVDD.n17075 VSS 0.031128f
C20341 DVDD.n17076 VSS 0.031128f
C20342 DVDD.n17077 VSS 0.031128f
C20343 DVDD.n17078 VSS 0.031128f
C20344 DVDD.n17080 VSS 0.031128f
C20345 DVDD.n17081 VSS 0.031128f
C20346 DVDD.n17082 VSS 0.031128f
C20347 DVDD.n17084 VSS 0.031128f
C20348 DVDD.n17085 VSS 0.031128f
C20349 DVDD.n17086 VSS 0.031128f
C20350 DVDD.n17087 VSS 0.031128f
C20351 DVDD.n17088 VSS 0.031128f
C20352 DVDD.n17089 VSS 0.031128f
C20353 DVDD.n17090 VSS 0.031128f
C20354 DVDD.n17092 VSS 0.031128f
C20355 DVDD.n17093 VSS 0.031128f
C20356 DVDD.n17094 VSS 0.031128f
C20357 DVDD.n17096 VSS 0.031128f
C20358 DVDD.n17097 VSS 0.031128f
C20359 DVDD.n17098 VSS 0.031128f
C20360 DVDD.n17099 VSS 0.031128f
C20361 DVDD.n17100 VSS 0.031128f
C20362 DVDD.n17101 VSS 0.031128f
C20363 DVDD.n17102 VSS 0.031128f
C20364 DVDD.n17104 VSS 0.031128f
C20365 DVDD.n17105 VSS 0.031128f
C20366 DVDD.n17106 VSS 0.031128f
C20367 DVDD.n17108 VSS 0.031128f
C20368 DVDD.n17109 VSS 0.031128f
C20369 DVDD.n17110 VSS 0.031128f
C20370 DVDD.n17111 VSS 0.031128f
C20371 DVDD.n17112 VSS 0.031128f
C20372 DVDD.n17113 VSS 0.031128f
C20373 DVDD.n17114 VSS 0.031128f
C20374 DVDD.n17116 VSS 0.031128f
C20375 DVDD.n17117 VSS 0.031128f
C20376 DVDD.n17118 VSS 0.031128f
C20377 DVDD.n17120 VSS 0.031128f
C20378 DVDD.n17121 VSS 0.031128f
C20379 DVDD.n17122 VSS 0.031128f
C20380 DVDD.n17123 VSS 0.031128f
C20381 DVDD.n17124 VSS 0.031128f
C20382 DVDD.n17125 VSS 0.031128f
C20383 DVDD.n17126 VSS 0.031128f
C20384 DVDD.n17128 VSS 0.031128f
C20385 DVDD.n17129 VSS 0.031128f
C20386 DVDD.n17130 VSS 0.031128f
C20387 DVDD.n17132 VSS 0.031128f
C20388 DVDD.n17133 VSS 0.031128f
C20389 DVDD.n17134 VSS 0.031128f
C20390 DVDD.n17135 VSS 0.031128f
C20391 DVDD.n17136 VSS 0.031128f
C20392 DVDD.n17137 VSS 0.031128f
C20393 DVDD.n17138 VSS 0.031128f
C20394 DVDD.n17140 VSS 0.031128f
C20395 DVDD.n17141 VSS 0.031128f
C20396 DVDD.n17142 VSS 0.031128f
C20397 DVDD.n17144 VSS 0.031128f
C20398 DVDD.n17145 VSS 0.031128f
C20399 DVDD.n17146 VSS 0.031128f
C20400 DVDD.n17147 VSS 0.031128f
C20401 DVDD.n17148 VSS 0.031128f
C20402 DVDD.n17149 VSS 0.031128f
C20403 DVDD.n17150 VSS 0.031128f
C20404 DVDD.n17152 VSS 0.031128f
C20405 DVDD.n17153 VSS 0.031128f
C20406 DVDD.n17154 VSS 0.031128f
C20407 DVDD.n17156 VSS 0.031128f
C20408 DVDD.n17157 VSS 0.031128f
C20409 DVDD.n17158 VSS 0.031128f
C20410 DVDD.n17159 VSS 0.031128f
C20411 DVDD.n17160 VSS 0.031128f
C20412 DVDD.n17161 VSS 0.031128f
C20413 DVDD.n17162 VSS 0.031128f
C20414 DVDD.n17164 VSS 0.031128f
C20415 DVDD.n17165 VSS 0.031128f
C20416 DVDD.n17166 VSS 0.031128f
C20417 DVDD.n17168 VSS 0.031128f
C20418 DVDD.n17169 VSS 0.031128f
C20419 DVDD.n17170 VSS 0.031128f
C20420 DVDD.n17171 VSS 0.031128f
C20421 DVDD.n17172 VSS 0.031128f
C20422 DVDD.n17173 VSS 0.031128f
C20423 DVDD.n17174 VSS 0.031128f
C20424 DVDD.n17176 VSS 0.031128f
C20425 DVDD.n17177 VSS 0.031128f
C20426 DVDD.n17178 VSS 0.031128f
C20427 DVDD.n17180 VSS 0.031128f
C20428 DVDD.n17181 VSS 0.031128f
C20429 DVDD.n17182 VSS 0.031128f
C20430 DVDD.n17183 VSS 0.031128f
C20431 DVDD.n17184 VSS 0.031128f
C20432 DVDD.n17185 VSS 0.031128f
C20433 DVDD.n17186 VSS 0.031128f
C20434 DVDD.n17188 VSS 0.031128f
C20435 DVDD.n17189 VSS 0.031128f
C20436 DVDD.n17190 VSS 0.031128f
C20437 DVDD.n17192 VSS 0.031128f
C20438 DVDD.n17193 VSS 0.031128f
C20439 DVDD.n17194 VSS 0.031128f
C20440 DVDD.n17195 VSS 0.031128f
C20441 DVDD.n17196 VSS 0.031128f
C20442 DVDD.n17197 VSS 0.031128f
C20443 DVDD.n17198 VSS 0.031128f
C20444 DVDD.n17200 VSS 0.031128f
C20445 DVDD.n17201 VSS 0.031128f
C20446 DVDD.n17202 VSS 0.031128f
C20447 DVDD.n17204 VSS 0.031128f
C20448 DVDD.n17205 VSS 0.031128f
C20449 DVDD.n17206 VSS 0.031128f
C20450 DVDD.n17207 VSS 0.031128f
C20451 DVDD.n17208 VSS 0.031128f
C20452 DVDD.n17209 VSS 0.031128f
C20453 DVDD.n17210 VSS 0.031128f
C20454 DVDD.n17212 VSS 0.031128f
C20455 DVDD.n17213 VSS 0.031128f
C20456 DVDD.n17214 VSS 0.031128f
C20457 DVDD.n17216 VSS 0.031128f
C20458 DVDD.n17217 VSS 0.031128f
C20459 DVDD.n17218 VSS 0.031128f
C20460 DVDD.n17219 VSS 0.031128f
C20461 DVDD.n17220 VSS 0.031128f
C20462 DVDD.n17221 VSS 0.031128f
C20463 DVDD.n17222 VSS 0.031128f
C20464 DVDD.n17224 VSS 0.031128f
C20465 DVDD.n17225 VSS 0.031128f
C20466 DVDD.n17226 VSS 0.031128f
C20467 DVDD.n17228 VSS 0.031128f
C20468 DVDD.n17229 VSS 0.031128f
C20469 DVDD.n17230 VSS 0.031128f
C20470 DVDD.n17231 VSS 0.031128f
C20471 DVDD.n17232 VSS 0.031128f
C20472 DVDD.n17233 VSS 0.031128f
C20473 DVDD.n17234 VSS 0.031128f
C20474 DVDD.n17236 VSS 0.031128f
C20475 DVDD.n17237 VSS 0.031128f
C20476 DVDD.n17238 VSS 0.031128f
C20477 DVDD.n17240 VSS 0.031128f
C20478 DVDD.n17241 VSS 0.031128f
C20479 DVDD.n17242 VSS 0.031128f
C20480 DVDD.n17243 VSS 0.031128f
C20481 DVDD.n17244 VSS 0.031128f
C20482 DVDD.n17245 VSS 0.031128f
C20483 DVDD.n17246 VSS 0.031128f
C20484 DVDD.n17248 VSS 0.031128f
C20485 DVDD.n17249 VSS 0.031128f
C20486 DVDD.n17250 VSS 0.031128f
C20487 DVDD.n17252 VSS 0.031128f
C20488 DVDD.n17253 VSS 0.031128f
C20489 DVDD.n17254 VSS 0.031128f
C20490 DVDD.n17255 VSS 0.031128f
C20491 DVDD.n17256 VSS 0.026086f
C20492 DVDD.n17257 VSS 0.031128f
C20493 DVDD.n17258 VSS 0.031128f
C20494 DVDD.n17259 VSS 0.031128f
C20495 DVDD.n17261 VSS 0.019729f
C20496 DVDD.n17262 VSS 0.290608f
C20497 DVDD.n17263 VSS 0.269549f
C20498 DVDD.n17264 VSS 0.029676f
C20499 DVDD.n17265 VSS 0.029676f
C20500 DVDD.n17266 VSS 0.025918f
C20501 DVDD.n17267 VSS 0.036621f
C20502 DVDD.n17268 VSS 0.02566f
C20503 DVDD.n17269 VSS 0.029381f
C20504 DVDD.n17270 VSS 0.029381f
C20505 DVDD.n17271 VSS 0.210585f
C20506 DVDD.n17272 VSS 0.526464f
C20507 DVDD.n17273 VSS 0.035544f
C20508 DVDD.n17274 VSS 0.035544f
C20509 DVDD.n17275 VSS 0.031727f
C20510 DVDD.n17276 VSS 0.039516f
C20511 DVDD.n17277 VSS 0.04802f
C20512 DVDD.n17278 VSS 0.053796f
C20513 DVDD.n17279 VSS 0.053796f
C20514 DVDD.n17280 VSS 0.585428f
C20515 DVDD.n17281 VSS 0.134774f
C20516 DVDD.n17282 VSS 0.033515f
C20517 DVDD.n17283 VSS 0.033515f
C20518 DVDD.n17284 VSS 0.029271f
C20519 DVDD.n17285 VSS 0.036621f
C20520 DVDD.n17286 VSS 0.022308f
C20521 DVDD.n17287 VSS 0.025542f
C20522 DVDD.n17288 VSS 0.025542f
C20523 DVDD.n17289 VSS 0.509617f
C20524 DVDD.n17290 VSS 0.176891f
C20525 DVDD.n17291 VSS 0.042269f
C20526 DVDD.n17292 VSS 0.042269f
C20527 DVDD.n17293 VSS 0.03773f
C20528 DVDD.n17294 VSS 0.039516f
C20529 DVDD.n17295 VSS 0.042017f
C20530 DVDD.n17296 VSS 0.047072f
C20531 DVDD.n17297 VSS 0.047072f
C20532 DVDD.n17298 VSS 0.176891f
C20533 DVDD.n17299 VSS 0.598063f
C20534 DVDD.n17300 VSS 0.522252f
C20535 DVDD.n17301 VSS 0.037354f
C20536 DVDD.n17302 VSS 0.037354f
C20537 DVDD.n17303 VSS 0.032623f
C20538 DVDD.n17304 VSS 0.036621f
C20539 DVDD.n17305 VSS 0.058284f
C20540 DVDD.n17306 VSS 0.522253f
C20541 DVDD.n17307 VSS 0.522253f
C20542 DVDD.n17308 VSS 1.3309f
C20543 DVDD.n17309 VSS 0.522253f
C20544 DVDD.n17311 VSS 0.657028f
C20545 DVDD.n17312 VSS 0.088457f
C20546 DVDD.n17313 VSS 0.063957f
C20547 DVDD.n17314 VSS 0.063957f
C20548 DVDD.n17315 VSS 0.063957f
C20549 DVDD.n17316 VSS 0.063957f
C20550 DVDD.n17317 VSS 0.063957f
C20551 DVDD.n17318 VSS 0.063957f
C20552 DVDD.n17319 VSS 0.063957f
C20553 DVDD.n17320 VSS 0.063957f
C20554 DVDD.n17321 VSS 0.063957f
C20555 DVDD.n17322 VSS 0.063957f
C20556 DVDD.n17323 VSS 0.063957f
C20557 DVDD.n17324 VSS 0.063957f
C20558 DVDD.n17325 VSS 0.063957f
C20559 DVDD.n17326 VSS 0.063957f
C20560 DVDD.n17327 VSS 0.063957f
C20561 DVDD.n17328 VSS 0.063957f
C20562 DVDD.n17329 VSS 0.063957f
C20563 DVDD.n17330 VSS 0.063957f
C20564 DVDD.n17331 VSS 0.063957f
C20565 DVDD.n17332 VSS 0.063957f
C20566 DVDD.n17333 VSS 0.063957f
C20567 DVDD.n17334 VSS 0.063957f
C20568 DVDD.n17335 VSS 0.063957f
C20569 DVDD.n17336 VSS 0.063957f
C20570 DVDD.n17337 VSS 0.063957f
C20571 DVDD.n17338 VSS 0.063957f
C20572 DVDD.n17339 VSS 0.063957f
C20573 DVDD.n17340 VSS 0.063957f
C20574 DVDD.n17341 VSS 0.063957f
C20575 DVDD.n17342 VSS 0.063957f
C20576 DVDD.n17343 VSS 0.063957f
C20577 DVDD.n17344 VSS 0.063957f
C20578 DVDD.n17345 VSS 0.063957f
C20579 DVDD.n17346 VSS 0.063957f
C20580 DVDD.n17347 VSS 0.063957f
C20581 DVDD.n17348 VSS 0.063957f
C20582 DVDD.n17349 VSS 0.063957f
C20583 DVDD.n17350 VSS 0.063957f
C20584 DVDD.n17351 VSS 0.063957f
C20585 DVDD.n17352 VSS 0.063957f
C20586 DVDD.n17353 VSS 0.063957f
C20587 DVDD.n17354 VSS 0.063957f
C20588 DVDD.n17355 VSS 0.063957f
C20589 DVDD.n17356 VSS 0.063957f
C20590 DVDD.n17357 VSS 0.063957f
C20591 DVDD.n17358 VSS 0.063957f
C20592 DVDD.n17359 VSS 0.063957f
C20593 DVDD.n17360 VSS 0.063957f
C20594 DVDD.n17361 VSS 0.059058f
C20595 DVDD.n17362 VSS 0.036879f
C20596 DVDD.n17364 VSS 0.522253f
C20597 DVDD.n17366 VSS 0.522253f
C20598 DVDD.n17367 VSS 0.522253f
C20599 DVDD.n17368 VSS 0.106252f
C20600 DVDD.n17369 VSS 0.522253f
C20601 DVDD.n17371 VSS 0.050805f
C20602 DVDD.n17374 VSS 0.063957f
C20603 DVDD.n17377 VSS 0.063957f
C20604 DVDD.n17380 VSS 0.063957f
C20605 DVDD.n17383 VSS 0.063957f
C20606 DVDD.n17386 VSS 0.063957f
C20607 DVDD.n17389 VSS 0.063957f
C20608 DVDD.n17392 VSS 0.063957f
C20609 DVDD.n17395 VSS 0.063957f
C20610 DVDD.n17398 VSS 0.063957f
C20611 DVDD.n17401 VSS 0.063957f
C20612 DVDD.n17404 VSS 0.063957f
C20613 DVDD.n17407 VSS 0.063957f
C20614 DVDD.n17410 VSS 0.063957f
C20615 DVDD.n17413 VSS 0.063957f
C20616 DVDD.n17416 VSS 0.063957f
C20617 DVDD.n17419 VSS 0.063957f
C20618 DVDD.n17422 VSS 0.063957f
C20619 DVDD.n17425 VSS 0.063957f
C20620 DVDD.n17428 VSS 0.063957f
C20621 DVDD.n17431 VSS 0.063957f
C20622 DVDD.n17434 VSS 0.063957f
C20623 DVDD.n17437 VSS 0.063957f
C20624 DVDD.n17440 VSS 0.063957f
C20625 DVDD.n17443 VSS 0.063957f
C20626 DVDD.n17446 VSS 0.063957f
C20627 DVDD.n17449 VSS 0.063957f
C20628 DVDD.n17452 VSS 0.063957f
C20629 DVDD.n17455 VSS 0.063957f
C20630 DVDD.n17458 VSS 0.063957f
C20631 DVDD.n17461 VSS 0.063957f
C20632 DVDD.n17464 VSS 0.063957f
C20633 DVDD.n17467 VSS 0.063957f
C20634 DVDD.n17470 VSS 0.063957f
C20635 DVDD.n17473 VSS 0.063957f
C20636 DVDD.n17476 VSS 0.063957f
C20637 DVDD.n17479 VSS 0.063957f
C20638 DVDD.n17482 VSS 0.063957f
C20639 DVDD.n17485 VSS 0.063957f
C20640 DVDD.n17488 VSS 0.063957f
C20641 DVDD.n17491 VSS 0.063957f
C20642 DVDD.n17494 VSS 0.063957f
C20643 DVDD.n17497 VSS 0.063957f
C20644 DVDD.n17500 VSS 0.063957f
C20645 DVDD.n17503 VSS 0.063957f
C20646 DVDD.n17506 VSS 0.063957f
C20647 DVDD.n17509 VSS 0.063957f
C20648 DVDD.n17512 VSS 0.063957f
C20649 DVDD.n17515 VSS 0.050031f
C20650 DVDD.n17516 VSS 0.063957f
C20651 DVDD.n17517 VSS 0.063957f
C20652 DVDD.n17518 VSS 0.063957f
C20653 DVDD.n17519 VSS 0.063957f
C20654 DVDD.n17520 VSS 0.063957f
C20655 DVDD.n17521 VSS 0.063957f
C20656 DVDD.n17522 VSS 0.063957f
C20657 DVDD.n17523 VSS 0.063957f
C20658 DVDD.n17524 VSS 0.063957f
C20659 DVDD.n17525 VSS 0.063957f
C20660 DVDD.n17526 VSS 0.063957f
C20661 DVDD.n17527 VSS 0.063957f
C20662 DVDD.n17528 VSS 0.063957f
C20663 DVDD.n17529 VSS 0.063957f
C20664 DVDD.n17530 VSS 0.063957f
C20665 DVDD.n17531 VSS 0.063957f
C20666 DVDD.n17532 VSS 0.063957f
C20667 DVDD.n17533 VSS 0.063957f
C20668 DVDD.n17534 VSS 0.063957f
C20669 DVDD.n17535 VSS 0.063957f
C20670 DVDD.n17536 VSS 0.063957f
C20671 DVDD.n17537 VSS 0.063957f
C20672 DVDD.n17538 VSS 0.063957f
C20673 DVDD.n17539 VSS 0.063957f
C20674 DVDD.n17540 VSS 0.063957f
C20675 DVDD.n17541 VSS 0.063957f
C20676 DVDD.n17542 VSS 0.063957f
C20677 DVDD.n17543 VSS 0.063957f
C20678 DVDD.n17544 VSS 0.063957f
C20679 DVDD.n17545 VSS 0.063957f
C20680 DVDD.n17546 VSS 0.063957f
C20681 DVDD.n17547 VSS 0.063957f
C20682 DVDD.n17548 VSS 0.063957f
C20683 DVDD.n17549 VSS 0.063957f
C20684 DVDD.n17550 VSS 0.063957f
C20685 DVDD.n17551 VSS 0.063957f
C20686 DVDD.n17552 VSS 0.063957f
C20687 DVDD.n17553 VSS 0.063957f
C20688 DVDD.n17554 VSS 0.063957f
C20689 DVDD.n17555 VSS 0.063957f
C20690 DVDD.n17556 VSS 0.063957f
C20691 DVDD.n17557 VSS 0.063957f
C20692 DVDD.n17558 VSS 0.063957f
C20693 DVDD.n17559 VSS 0.063957f
C20694 DVDD.n17560 VSS 0.063957f
C20695 DVDD.n17561 VSS 0.063957f
C20696 DVDD.n17562 VSS 0.063957f
C20697 DVDD.n17563 VSS 0.063957f
C20698 DVDD.n17564 VSS 0.063957f
C20699 DVDD.n17565 VSS 0.063957f
C20700 DVDD.n17566 VSS 0.063957f
C20701 DVDD.n17567 VSS 0.063957f
C20702 DVDD.n17568 VSS 0.063957f
C20703 DVDD.n17569 VSS 0.063957f
C20704 DVDD.n17570 VSS 0.063957f
C20705 DVDD.n17571 VSS 0.063957f
C20706 DVDD.n17572 VSS 0.063957f
C20707 DVDD.n17573 VSS 0.063957f
C20708 DVDD.n17574 VSS 0.063957f
C20709 DVDD.n17575 VSS 0.063957f
C20710 DVDD.n17576 VSS 0.063957f
C20711 DVDD.n17577 VSS 0.063957f
C20712 DVDD.n17578 VSS 0.063957f
C20713 DVDD.n17579 VSS 0.063957f
C20714 DVDD.n17580 VSS 0.063957f
C20715 DVDD.n17581 VSS 0.063957f
C20716 DVDD.n17582 VSS 0.063957f
C20717 DVDD.n17583 VSS 0.063957f
C20718 DVDD.n17584 VSS 0.063957f
C20719 DVDD.n17585 VSS 0.063957f
C20720 DVDD.n17586 VSS 0.063957f
C20721 DVDD.n17587 VSS 0.063957f
C20722 DVDD.n17588 VSS 0.063957f
C20723 DVDD.n17589 VSS 0.063957f
C20724 DVDD.n17590 VSS 0.063957f
C20725 DVDD.n17591 VSS 0.063957f
C20726 DVDD.n17592 VSS 0.063957f
C20727 DVDD.n17593 VSS 0.063957f
C20728 DVDD.n17594 VSS 0.063957f
C20729 DVDD.n17595 VSS 0.063957f
C20730 DVDD.n17596 VSS 0.063957f
C20731 DVDD.n17597 VSS 0.063957f
C20732 DVDD.n17598 VSS 0.063957f
C20733 DVDD.n17599 VSS 0.063957f
C20734 DVDD.n17600 VSS 0.063957f
C20735 DVDD.n17601 VSS 0.063957f
C20736 DVDD.n17602 VSS 0.063957f
C20737 DVDD.n17603 VSS 0.063957f
C20738 DVDD.n17604 VSS 0.063957f
C20739 DVDD.n17605 VSS 0.063957f
C20740 DVDD.n17606 VSS 0.063957f
C20741 DVDD.n17607 VSS 0.063957f
C20742 DVDD.n17608 VSS 0.063957f
C20743 DVDD.n17609 VSS 0.063957f
C20744 DVDD.n17610 VSS 0.063957f
C20745 DVDD.n17611 VSS 0.063957f
C20746 DVDD.n17612 VSS 0.050805f
C20747 DVDD.n17613 VSS 0.063957f
C20748 DVDD.n17614 VSS 0.063957f
C20749 DVDD.n17615 VSS 0.063957f
C20750 DVDD.n17616 VSS 0.063957f
C20751 DVDD.n17617 VSS 0.063957f
C20752 DVDD.n17618 VSS 0.063957f
C20753 DVDD.n17619 VSS 0.063957f
C20754 DVDD.n17620 VSS 0.063957f
C20755 DVDD.n17621 VSS 0.063957f
C20756 DVDD.n17622 VSS 0.063957f
C20757 DVDD.n17623 VSS 0.063957f
C20758 DVDD.n17624 VSS 0.063957f
C20759 DVDD.n17625 VSS 0.063957f
C20760 DVDD.n17626 VSS 0.063957f
C20761 DVDD.n17627 VSS 0.063957f
C20762 DVDD.n17628 VSS 0.063957f
C20763 DVDD.n17629 VSS 0.063957f
C20764 DVDD.n17630 VSS 0.063957f
C20765 DVDD.n17631 VSS 0.063957f
C20766 DVDD.n17632 VSS 0.063957f
C20767 DVDD.n17633 VSS 0.063957f
C20768 DVDD.n17634 VSS 0.063957f
C20769 DVDD.n17635 VSS 0.063957f
C20770 DVDD.n17636 VSS 0.063957f
C20771 DVDD.n17637 VSS 0.063957f
C20772 DVDD.n17638 VSS 0.063957f
C20773 DVDD.n17639 VSS 0.063957f
C20774 DVDD.n17640 VSS 0.063957f
C20775 DVDD.n17641 VSS 0.063957f
C20776 DVDD.n17642 VSS 0.063957f
C20777 DVDD.n17643 VSS 0.063957f
C20778 DVDD.n17644 VSS 0.063957f
C20779 DVDD.n17645 VSS 0.063957f
C20780 DVDD.n17646 VSS 0.063957f
C20781 DVDD.n17647 VSS 0.063957f
C20782 DVDD.n17648 VSS 0.063957f
C20783 DVDD.n17649 VSS 0.063957f
C20784 DVDD.n17650 VSS 0.063957f
C20785 DVDD.n17651 VSS 0.063957f
C20786 DVDD.n17652 VSS 0.063957f
C20787 DVDD.n17653 VSS 0.063957f
C20788 DVDD.n17654 VSS 0.063957f
C20789 DVDD.n17655 VSS 0.063957f
C20790 DVDD.n17656 VSS 0.063957f
C20791 DVDD.n17657 VSS 0.063957f
C20792 DVDD.n17658 VSS 0.063957f
C20793 DVDD.n17659 VSS 0.063957f
C20794 DVDD.n17660 VSS 0.063957f
C20795 DVDD.n17661 VSS 0.063957f
C20796 DVDD.n17662 VSS 0.063957f
C20797 DVDD.n17663 VSS 0.063957f
C20798 DVDD.n17664 VSS 0.063957f
C20799 DVDD.n17665 VSS 0.063957f
C20800 DVDD.n17666 VSS 0.063957f
C20801 DVDD.n17667 VSS 0.063957f
C20802 DVDD.n17668 VSS 0.063957f
C20803 DVDD.n17669 VSS 0.063957f
C20804 DVDD.n17670 VSS 0.063957f
C20805 DVDD.n17671 VSS 0.063957f
C20806 DVDD.n17672 VSS 0.063957f
C20807 DVDD.n17673 VSS 0.063957f
C20808 DVDD.n17674 VSS 0.063957f
C20809 DVDD.n17675 VSS 0.063957f
C20810 DVDD.n17676 VSS 0.063957f
C20811 DVDD.n17677 VSS 0.063957f
C20812 DVDD.n17678 VSS 0.063957f
C20813 DVDD.n17679 VSS 0.063957f
C20814 DVDD.n17680 VSS 0.063957f
C20815 DVDD.n17681 VSS 0.063957f
C20816 DVDD.n17682 VSS 0.063957f
C20817 DVDD.n17683 VSS 0.063957f
C20818 DVDD.n17684 VSS 0.063957f
C20819 DVDD.n17685 VSS 0.063957f
C20820 DVDD.n17686 VSS 0.063957f
C20821 DVDD.n17687 VSS 0.063957f
C20822 DVDD.n17688 VSS 0.063957f
C20823 DVDD.n17689 VSS 0.063957f
C20824 DVDD.n17690 VSS 0.063957f
C20825 DVDD.n17691 VSS 0.063957f
C20826 DVDD.n17692 VSS 0.063957f
C20827 DVDD.n17693 VSS 0.063957f
C20828 DVDD.n17694 VSS 0.063957f
C20829 DVDD.n17695 VSS 0.063957f
C20830 DVDD.n17696 VSS 0.063957f
C20831 DVDD.n17697 VSS 0.063957f
C20832 DVDD.n17698 VSS 0.063957f
C20833 DVDD.n17699 VSS 0.063957f
C20834 DVDD.n17700 VSS 0.063957f
C20835 DVDD.n17701 VSS 0.063957f
C20836 DVDD.n17702 VSS 0.063957f
C20837 DVDD.n17703 VSS 0.063957f
C20838 DVDD.n17704 VSS 0.063957f
C20839 DVDD.n17705 VSS 0.063957f
C20840 DVDD.n17706 VSS 0.063957f
C20841 DVDD.n17707 VSS 0.063957f
C20842 DVDD.n17708 VSS 0.063957f
C20843 DVDD.n17709 VSS 0.063957f
C20844 DVDD.n17710 VSS 0.522253f
C20845 DVDD.n17711 VSS 0.104963f
C20846 DVDD.n17712 VSS 0.10523f
C20847 DVDD.n17713 VSS 0.13474f
C20848 DVDD.n17714 VSS 0.023855f
C20849 DVDD.n17715 VSS 0.027314f
C20850 DVDD.n17716 VSS 0.027314f
C20851 DVDD.n17717 VSS 0.522252f
C20852 DVDD.n17718 VSS 0.598063f
C20853 DVDD.n17719 VSS 0.058119f
C20854 DVDD.n17720 VSS 0.058119f
C20855 DVDD.n17721 VSS 0.053165f
C20856 DVDD.n17723 VSS 0.053165f
C20857 DVDD.n17724 VSS 0.053165f
C20858 DVDD.n17725 VSS 0.088457f
C20859 DVDD.n17726 VSS 0.026154f
C20860 DVDD.n17727 VSS 0.379993f
C20861 DVDD.n17728 VSS 0.026573f
C20862 DVDD.n17730 VSS 0.030844f
C20863 DVDD.n17731 VSS 0.36811f
C20864 DVDD.n17733 VSS 0.025624f
C20865 DVDD.n17734 VSS 0.06615f
C20866 DVDD.n17736 VSS 0.035233f
C20867 DVDD.n17737 VSS 0.06615f
C20868 DVDD.n17738 VSS 0.117599f
C20869 DVDD.n17739 VSS 0.132299f
C20870 DVDD.n17740 VSS 0.025624f
C20871 DVDD.n17741 VSS 0.025624f
C20872 DVDD.n17742 VSS 0.025624f
C20873 DVDD.n17743 VSS 0.132299f
C20874 DVDD.n17744 VSS 0.132299f
C20875 DVDD.n17745 VSS 0.132299f
C20876 DVDD.n17746 VSS 0.025624f
C20877 DVDD.n17747 VSS 0.025624f
C20878 DVDD.n17748 VSS 0.025624f
C20879 DVDD.n17749 VSS 0.132299f
C20880 DVDD.n17750 VSS 0.132299f
C20881 DVDD.n17751 VSS 0.132299f
C20882 DVDD.n17752 VSS 0.025624f
C20883 DVDD.n17753 VSS 0.025624f
C20884 DVDD.n17754 VSS 0.025624f
C20885 DVDD.n17755 VSS 0.132299f
C20886 DVDD.n17756 VSS 0.132299f
C20887 DVDD.n17757 VSS 0.132299f
C20888 DVDD.n17758 VSS 0.025624f
C20889 DVDD.n17759 VSS 0.025624f
C20890 DVDD.n17760 VSS 0.025624f
C20891 DVDD.n17761 VSS 0.132299f
C20892 DVDD.n17762 VSS 0.132299f
C20893 DVDD.n17763 VSS 0.132299f
C20894 DVDD.n17764 VSS 0.025624f
C20895 DVDD.n17765 VSS 0.025624f
C20896 DVDD.n17766 VSS 0.025624f
C20897 DVDD.n17767 VSS 0.132299f
C20898 DVDD.n17768 VSS 0.132299f
C20899 DVDD.n17769 VSS 0.132299f
C20900 DVDD.n17770 VSS 0.025624f
C20901 DVDD.n17771 VSS 0.025624f
C20902 DVDD.n17772 VSS 0.025624f
C20903 DVDD.n17773 VSS 0.132299f
C20904 DVDD.n17774 VSS 0.132299f
C20905 DVDD.n17775 VSS 0.132299f
C20906 DVDD.n17776 VSS 0.025624f
C20907 DVDD.n17777 VSS 0.025624f
C20908 DVDD.n17778 VSS 0.025624f
C20909 DVDD.n17779 VSS 0.132299f
C20910 DVDD.n17780 VSS 0.132299f
C20911 DVDD.n17781 VSS 0.132299f
C20912 DVDD.n17782 VSS 0.025624f
C20913 DVDD.n17783 VSS 0.025624f
C20914 DVDD.n17784 VSS 0.025624f
C20915 DVDD.n17785 VSS 0.132299f
C20916 DVDD.n17786 VSS 0.132299f
C20917 DVDD.n17787 VSS 0.132299f
C20918 DVDD.n17788 VSS 0.025624f
C20919 DVDD.n17789 VSS 0.025624f
C20920 DVDD.n17790 VSS 0.025624f
C20921 DVDD.n17791 VSS 0.132299f
C20922 DVDD.n17792 VSS 0.132299f
C20923 DVDD.n17793 VSS 0.132299f
C20924 DVDD.n17794 VSS 0.025624f
C20925 DVDD.n17795 VSS 0.025624f
C20926 DVDD.n17796 VSS 0.025624f
C20927 DVDD.n17797 VSS 0.132299f
C20928 DVDD.n17798 VSS 0.132299f
C20929 DVDD.n17799 VSS 0.132299f
C20930 DVDD.n17800 VSS 0.025624f
C20931 DVDD.n17801 VSS 0.025624f
C20932 DVDD.n17802 VSS 0.025624f
C20933 DVDD.n17803 VSS 0.132299f
C20934 DVDD.n17804 VSS 0.132299f
C20935 DVDD.n17805 VSS 0.132299f
C20936 DVDD.n17806 VSS 0.025624f
C20937 DVDD.n17807 VSS 0.025624f
C20938 DVDD.n17808 VSS 0.025624f
C20939 DVDD.n17809 VSS 0.132299f
C20940 DVDD.n17810 VSS 0.132299f
C20941 DVDD.n17811 VSS 0.132299f
C20942 DVDD.n17812 VSS 0.025624f
C20943 DVDD.n17813 VSS 0.025624f
C20944 DVDD.n17814 VSS 0.025624f
C20945 DVDD.n17815 VSS 0.132299f
C20946 DVDD.n17816 VSS 0.132299f
C20947 DVDD.n17817 VSS 0.132299f
C20948 DVDD.n17818 VSS 0.025624f
C20949 DVDD.n17819 VSS 0.025624f
C20950 DVDD.n17820 VSS 0.025624f
C20951 DVDD.n17821 VSS 0.132299f
C20952 DVDD.n17822 VSS 0.132299f
C20953 DVDD.n17823 VSS 0.132299f
C20954 DVDD.n17824 VSS 0.025624f
C20955 DVDD.n17825 VSS 0.025624f
C20956 DVDD.n17826 VSS 0.025624f
C20957 DVDD.n17827 VSS 0.132299f
C20958 DVDD.n17828 VSS 0.132299f
C20959 DVDD.n17829 VSS 0.132299f
C20960 DVDD.n17830 VSS 0.025624f
C20961 DVDD.n17831 VSS 0.025624f
C20962 DVDD.n17832 VSS 0.025624f
C20963 DVDD.n17833 VSS 0.132299f
C20964 DVDD.n17834 VSS 0.132299f
C20965 DVDD.n17835 VSS 0.132299f
C20966 DVDD.n17836 VSS 0.025624f
C20967 DVDD.n17837 VSS 0.025624f
C20968 DVDD.n17838 VSS 0.025624f
C20969 DVDD.n17839 VSS 0.132299f
C20970 DVDD.n17840 VSS 0.132299f
C20971 DVDD.n17841 VSS 0.132299f
C20972 DVDD.n17842 VSS 0.025624f
C20973 DVDD.n17843 VSS 0.025624f
C20974 DVDD.n17844 VSS 0.025624f
C20975 DVDD.n17845 VSS 0.132299f
C20976 DVDD.n17846 VSS 0.132299f
C20977 DVDD.n17847 VSS 0.132299f
C20978 DVDD.n17848 VSS 0.025624f
C20979 DVDD.n17849 VSS 0.025624f
C20980 DVDD.n17850 VSS 0.025624f
C20981 DVDD.n17851 VSS 0.132299f
C20982 DVDD.n17852 VSS 0.132299f
C20983 DVDD.n17853 VSS 0.132299f
C20984 DVDD.n17854 VSS 0.025624f
C20985 DVDD.n17855 VSS 0.025624f
C20986 DVDD.n17856 VSS 0.025624f
C20987 DVDD.n17857 VSS 0.132299f
C20988 DVDD.n17858 VSS 0.132299f
C20989 DVDD.n17859 VSS 0.132299f
C20990 DVDD.n17860 VSS 0.025624f
C20991 DVDD.n17861 VSS 0.025624f
C20992 DVDD.n17862 VSS 0.025624f
C20993 DVDD.n17863 VSS 0.132299f
C20994 DVDD.n17864 VSS 0.132299f
C20995 DVDD.n17865 VSS 0.132299f
C20996 DVDD.n17866 VSS 0.025624f
C20997 DVDD.n17867 VSS 0.025624f
C20998 DVDD.n17868 VSS 0.025624f
C20999 DVDD.n17869 VSS 0.132299f
C21000 DVDD.n17870 VSS 0.132299f
C21001 DVDD.n17871 VSS 0.128624f
C21002 DVDD.n17872 VSS 0.025624f
C21003 DVDD.n17873 VSS 0.025624f
C21004 DVDD.n17874 VSS 0.025624f
C21005 DVDD.n17875 VSS 0.072275f
C21006 DVDD.n17876 VSS 0.06615f
C21007 DVDD.n17877 VSS 0.064086f
C21008 DVDD.n17878 VSS 0.06615f
C21009 DVDD.n17879 VSS 0.104124f
C21010 DVDD.n17880 VSS 0.132299f
C21011 DVDD.n17881 VSS 0.025624f
C21012 DVDD.n17882 VSS 0.025624f
C21013 DVDD.n17883 VSS 0.025624f
C21014 DVDD.n17884 VSS 0.132299f
C21015 DVDD.n17885 VSS 0.132299f
C21016 DVDD.n17886 VSS 0.132299f
C21017 DVDD.n17887 VSS 0.025624f
C21018 DVDD.n17888 VSS 0.025624f
C21019 DVDD.n17889 VSS 0.025624f
C21020 DVDD.n17890 VSS 0.132299f
C21021 DVDD.n17891 VSS 0.132299f
C21022 DVDD.n17892 VSS 0.132299f
C21023 DVDD.n17893 VSS 0.025624f
C21024 DVDD.n17894 VSS 0.025624f
C21025 DVDD.n17895 VSS 0.019218f
C21026 DVDD.n17896 VSS 0.132299f
C21027 DVDD.n17897 VSS 0.132299f
C21028 DVDD.n17898 VSS 0.132299f
C21029 DVDD.n17899 VSS 0.025624f
C21030 DVDD.n17900 VSS 0.025624f
C21031 DVDD.n17901 VSS 0.025624f
C21032 DVDD.n17902 VSS 0.132299f
C21033 DVDD.n17903 VSS 0.132299f
C21034 DVDD.n17904 VSS 0.100449f
C21035 DVDD.n17905 VSS 0.025624f
C21036 DVDD.n17906 VSS 0.075949f
C21037 DVDD.n17907 VSS 0.025624f
C21038 DVDD.n17908 VSS 0.075949f
C21039 DVDD.n17909 VSS 0.025624f
C21040 DVDD.n17910 VSS 0.075949f
C21041 DVDD.n17911 VSS 0.025624f
C21042 DVDD.n17912 VSS 0.025624f
C21043 DVDD.n17913 VSS 0.0686f
C21044 DVDD.n17914 VSS 0.0735f
C21045 DVDD.n17915 VSS 0.025624f
C21046 DVDD.n17916 VSS 0.075949f
C21047 DVDD.n17917 VSS 0.025624f
C21048 DVDD.n17918 VSS 0.075949f
C21049 DVDD.n17919 VSS 0.025624f
C21050 DVDD.n17920 VSS 0.075949f
C21051 DVDD.n17921 VSS 0.025624f
C21052 DVDD.n17922 VSS 0.075949f
C21053 DVDD.n17923 VSS 0.025624f
C21054 DVDD.n17924 VSS 0.075949f
C21055 DVDD.n17925 VSS 0.025624f
C21056 DVDD.n17926 VSS 0.075949f
C21057 DVDD.n17927 VSS 0.025624f
C21058 DVDD.n17928 VSS 0.025624f
C21059 DVDD.n17929 VSS 0.075949f
C21060 DVDD.n17930 VSS 0.025624f
C21061 DVDD.n17931 VSS 0.075949f
C21062 DVDD.n17932 VSS 0.025624f
C21063 DVDD.n17933 VSS 0.075949f
C21064 DVDD.n17934 VSS 0.025624f
C21065 DVDD.n17935 VSS 0.075949f
C21066 DVDD.n17936 VSS 0.025624f
C21067 DVDD.n17937 VSS 0.075949f
C21068 DVDD.n17938 VSS 0.025624f
C21069 DVDD.n17939 VSS 0.075949f
C21070 DVDD.n17940 VSS 0.025624f
C21071 DVDD.n17941 VSS 0.025624f
C21072 DVDD.n17942 VSS 0.0735f
C21073 DVDD.n17943 VSS 0.0686f
C21074 DVDD.n17944 VSS 0.025624f
C21075 DVDD.n17945 VSS 0.075949f
C21076 DVDD.n17946 VSS 0.025624f
C21077 DVDD.n17947 VSS 0.075949f
C21078 DVDD.n17948 VSS 0.025624f
C21079 DVDD.n17949 VSS 0.075949f
C21080 DVDD.n17950 VSS 0.025624f
C21081 DVDD.n17951 VSS 0.025624f
C21082 DVDD.n17952 VSS 0.075949f
C21083 DVDD.n17953 VSS 0.06615f
C21084 DVDD.n17954 VSS 0.808336f
C21085 DVDD.n17955 VSS 0.06615f
C21086 DVDD.n17956 VSS 0.07105f
C21087 DVDD.n17957 VSS 0.132299f
C21088 DVDD.n17958 VSS 0.025624f
C21089 DVDD.n17959 VSS 0.025624f
C21090 DVDD.n17960 VSS 0.025624f
C21091 DVDD.n17961 VSS 0.075949f
C21092 DVDD.n17962 VSS 0.06615f
C21093 DVDD.n17963 VSS 0.137328f
C21094 DVDD.n17964 VSS 0.06615f
C21095 DVDD.n17965 VSS 0.075949f
C21096 DVDD.n17966 VSS 0.025624f
C21097 DVDD.n17967 VSS 0.025624f
C21098 DVDD.n17968 VSS 0.095549f
C21099 DVDD.n17969 VSS 0.132299f
C21100 DVDD.n17970 VSS 0.117599f
C21101 DVDD.n17971 VSS 0.025624f
C21102 DVDD.n17972 VSS 0.075949f
C21103 DVDD.n17973 VSS 0.025624f
C21104 DVDD.n17974 VSS 0.025624f
C21105 DVDD.n17975 VSS 0.025624f
C21106 DVDD.n17976 VSS 0.07105f
C21107 DVDD.n17977 VSS 0.06615f
C21108 DVDD.n17978 VSS 0.137328f
C21109 DVDD.n17979 VSS 0.06615f
C21110 DVDD.n17980 VSS 0.075949f
C21111 DVDD.n17981 VSS 0.025624f
C21112 DVDD.n17982 VSS 0.025624f
C21113 DVDD.n17983 VSS 0.120049f
C21114 DVDD.n17984 VSS 0.132299f
C21115 DVDD.n17985 VSS 0.093099f
C21116 DVDD.n17986 VSS 0.025624f
C21117 DVDD.n17987 VSS 0.075949f
C21118 DVDD.n17988 VSS 0.025624f
C21119 DVDD.n17989 VSS 0.075949f
C21120 DVDD.n17990 VSS 0.025624f
C21121 DVDD.n17991 VSS 0.075949f
C21122 DVDD.n17992 VSS 0.025624f
C21123 DVDD.n17993 VSS 0.075949f
C21124 DVDD.n17994 VSS 0.025624f
C21125 DVDD.n17995 VSS 0.025624f
C21126 DVDD.n17996 VSS 0.075949f
C21127 DVDD.n17997 VSS 0.025624f
C21128 DVDD.n17998 VSS 0.075949f
C21129 DVDD.n17999 VSS 0.025624f
C21130 DVDD.n18000 VSS 0.075949f
C21131 DVDD.n18001 VSS 0.025624f
C21132 DVDD.n18002 VSS 0.075949f
C21133 DVDD.n18003 VSS 0.025624f
C21134 DVDD.n18004 VSS 0.075949f
C21135 DVDD.n18005 VSS 0.025624f
C21136 DVDD.n18006 VSS 0.075949f
C21137 DVDD.n18007 VSS 0.025624f
C21138 DVDD.n18008 VSS 0.025624f
C21139 DVDD.n18009 VSS 0.0735f
C21140 DVDD.n18010 VSS 0.0686f
C21141 DVDD.n18011 VSS 0.025624f
C21142 DVDD.n18012 VSS 0.075949f
C21143 DVDD.n18013 VSS 0.025624f
C21144 DVDD.n18014 VSS 0.075949f
C21145 DVDD.n18015 VSS 0.025624f
C21146 DVDD.n18016 VSS 0.075949f
C21147 DVDD.n18017 VSS 0.025624f
C21148 DVDD.n18018 VSS 0.075949f
C21149 DVDD.n18019 VSS 0.025624f
C21150 DVDD.n18020 VSS 0.075949f
C21151 DVDD.n18021 VSS 0.025624f
C21152 DVDD.n18022 VSS 0.013761f
C21153 DVDD.n18023 VSS 0.06615f
C21154 DVDD.n18024 VSS 0.025624f
C21155 DVDD.n18025 VSS 0.025624f
C21156 DVDD.n18027 VSS 0.06125f
C21157 DVDD.n18028 VSS 0.025624f
C21158 DVDD.n18030 VSS 0.025624f
C21159 DVDD.n18032 VSS 0.06615f
C21160 DVDD.n18034 VSS 0.05635f
C21161 DVDD.n18035 VSS 0.030844f
C21162 DVDD.n18036 VSS 0.0294f
C21163 DVDD.n18037 VSS 0.090649f
C21164 DVDD.n18040 VSS 0.124756f
C21165 DVDD.n18042 VSS 0.151899f
C21166 DVDD.n18043 VSS 0.808336f
C21167 DVDD.n18044 VSS 1.27277f
C21168 DVDD.n18045 VSS 1.27277f
C21169 DVDD.n18046 VSS 0.151899f
C21170 DVDD.n18047 VSS 0.151899f
C21171 DVDD.n18048 VSS 0.151899f
C21172 DVDD.n18049 VSS 0.151899f
C21173 DVDD.n18054 VSS 0.053642f
C21174 DVDD.n18057 VSS 0.065505f
C21175 DVDD.n18058 VSS 0.073242f
C21176 DVDD.n18059 VSS 0.073242f
C21177 DVDD.n18061 VSS 0.071694f
C21178 DVDD.n18062 VSS 0.073242f
C21179 DVDD.n18063 VSS 0.073242f
C21180 DVDD.n18064 VSS 0.086309f
C21181 DVDD.n18065 VSS 0.042891f
C21182 DVDD.n18066 VSS 0.085784f
C21183 DVDD.n18067 VSS 0.037455f
C21184 DVDD.n18068 VSS 0.077504f
C21185 DVDD.n18069 VSS 0.146483f
C21186 DVDD.n18070 VSS 0.063957f
C21187 DVDD.n18071 VSS 0.146483f
C21188 DVDD.n18072 VSS 0.063957f
C21189 DVDD.n18073 VSS 0.146483f
C21190 DVDD.n18074 VSS 0.063957f
C21191 DVDD.n18075 VSS 0.146483f
C21192 DVDD.n18076 VSS 0.146483f
C21193 DVDD.n18077 VSS 0.146483f
C21194 DVDD.n18078 VSS 0.063957f
C21195 DVDD.n18079 VSS 0.146483f
C21196 DVDD.n18084 VSS 0.063957f
C21197 DVDD.n18085 VSS 0.073242f
C21198 DVDD.n18086 VSS 0.063957f
C21199 DVDD.n18087 VSS 0.146483f
C21200 DVDD.n18088 VSS 0.146483f
C21201 DVDD.n18089 VSS 0.146483f
C21202 DVDD.n18090 VSS 0.126883f
C21203 DVDD.n18091 VSS 0.126883f
C21204 DVDD.n18092 VSS 0.077504f
C21205 DVDD.n18093 VSS 0.042891f
C21206 DVDD.n18094 VSS 0.037455f
C21207 DVDD.n18095 VSS 0.042891f
C21208 DVDD.n18097 VSS 0.042891f
C21209 DVDD.n18098 VSS 0.085784f
C21210 DVDD.n18099 VSS 0.081467f
C21211 DVDD.n18100 VSS 0.085784f
C21212 DVDD.n18101 VSS 0.037455f
C21213 DVDD.n18102 VSS 0.042891f
C21214 DVDD.n18103 VSS 0.084905f
C21215 DVDD.n18104 VSS 0.037455f
C21216 DVDD.n18105 VSS 0.038965f
C21217 DVDD.n18106 VSS 0.041382f
C21218 DVDD.n18107 VSS 0.037455f
C21219 DVDD.n18108 VSS 0.085784f
C21220 DVDD.n18109 VSS 0.244123f
C21221 DVDD.n18110 VSS 0.085784f
C21222 DVDD.n18111 VSS 0.061921f
C21223 DVDD.n18112 VSS 0.061921f
C21224 DVDD.n18113 VSS 0.03383f
C21225 DVDD.n18114 VSS 0.042946f
C21226 DVDD.n18115 VSS 0.037455f
C21227 DVDD.n18116 VSS 0.06313f
C21228 DVDD.n18117 VSS 0.06313f
C21229 DVDD.n18118 VSS 0.085784f
C21230 DVDD.n18119 VSS 0.248786f
C21231 DVDD.n18120 VSS 0.085784f
C21232 DVDD.n18121 VSS 0.085784f
C21233 DVDD.n18122 VSS 0.037455f
C21234 DVDD.n18123 VSS 0.038361f
C21235 DVDD.n18124 VSS 0.086577f
C21236 DVDD.n18125 VSS 0.292773f
C21237 DVDD.n18126 VSS 0.073242f
C21238 DVDD.n18127 VSS 0.063957f
C21239 DVDD.n18128 VSS 0.146483f
C21240 DVDD.n18129 VSS 0.146483f
C21241 DVDD.n18130 VSS 0.146483f
C21242 DVDD.n18131 VSS 0.134104f
C21243 DVDD.n18132 VSS 0.134104f
C21244 DVDD.n18133 VSS 0.134104f
C21245 DVDD.n18134 VSS 0.21057f
C21246 DVDD.n18135 VSS 0.251446f
C21247 DVDD.n18136 VSS 0.221466f
C21248 DVDD.n18137 VSS 0.274656f
C21249 DVDD.n18138 VSS 0.11992f
C21250 DVDD.n18139 VSS 0.274656f
C21251 DVDD.n18140 VSS 0.274656f
C21252 DVDD.n18141 VSS 0.274656f
C21253 DVDD.n18142 VSS 0.274656f
C21254 DVDD.n18143 VSS 0.274656f
C21255 DVDD.n18144 VSS 0.11992f
C21256 DVDD.n18145 VSS 0.274656f
C21257 DVDD.n18146 VSS 0.11992f
C21258 DVDD.n18147 VSS 0.274656f
C21259 DVDD.n18148 VSS 0.274656f
C21260 DVDD.n18149 VSS 0.274656f
C21261 DVDD.n18150 VSS 0.274656f
C21262 DVDD.n18151 VSS 0.274656f
C21263 DVDD.n18152 VSS 0.11992f
C21264 DVDD.n18153 VSS 0.274656f
C21265 DVDD.n18154 VSS 0.11992f
C21266 DVDD.n18155 VSS 0.247577f
C21267 DVDD.n18156 VSS 0.247577f
C21268 DVDD.n18157 VSS 0.030947f
C21269 DVDD.n18158 VSS 0.164407f
C21270 DVDD.n18159 VSS 0.11992f
C21271 DVDD.n18160 VSS 0.274656f
C21272 DVDD.n18161 VSS 0.478216f
C21273 DVDD.n18162 VSS 0.529582f
C21274 DVDD.n18164 VSS 0.151899f
C21275 DVDD.n18166 VSS 0.151899f
C21276 DVDD.n18168 VSS 0.151899f
C21277 DVDD.n18170 VSS 0.151899f
C21278 DVDD.n18172 VSS 0.151899f
C21279 DVDD.n18174 VSS 0.151899f
C21280 DVDD.n18176 VSS 0.151899f
C21281 DVDD.n18178 VSS 0.151899f
C21282 DVDD.n18180 VSS 0.151899f
C21283 DVDD.n18182 VSS 0.151899f
C21284 DVDD.n18194 VSS 0.124756f
C21285 DVDD.n18196 VSS 0.151899f
C21286 DVDD.n18197 VSS 0.876514f
C21287 DVDD.n18198 VSS 3.23275f
C21288 DVDD.n18199 VSS 3.23275f
C21289 DVDD.n18200 VSS 0.151899f
C21290 DVDD.n18201 VSS 0.151899f
C21291 DVDD.n18202 VSS 0.151899f
C21292 DVDD.n18203 VSS 0.151899f
C21293 DVDD.n18204 VSS 0.151899f
C21294 DVDD.n18205 VSS 0.277582f
C21295 DVDD.n18206 VSS 0.038361f
C21296 DVDD.n18207 VSS 0.085784f
C21297 DVDD.n18208 VSS 0.085784f
C21298 DVDD.n18209 VSS 0.085784f
C21299 DVDD.n18210 VSS 0.042891f
C21300 DVDD.n18211 VSS 0.037455f
C21301 DVDD.n18212 VSS 0.151899f
C21302 DVDD.n18213 VSS 0.11992f
C21303 DVDD.n18214 VSS 0.11992f
C21304 DVDD.n18215 VSS 0.163891f
C21305 DVDD.n18216 VSS 0.01831f
C21306 DVDD.n18217 VSS 0.137328f
C21307 DVDD.n18218 VSS 0.016376f
C21308 DVDD.n18219 VSS 0.11992f
C21309 DVDD.n18220 VSS 0.163891f
C21310 DVDD.n18221 VSS 0.274656f
C21311 DVDD.n18222 VSS 0.274656f
C21312 DVDD.n18223 VSS 0.274656f
C21313 DVDD.n18224 VSS 0.11992f
C21314 DVDD.n18225 VSS 0.163891f
C21315 DVDD.n18226 VSS 0.202124f
C21316 DVDD.n18227 VSS 0.11992f
C21317 DVDD.n18228 VSS 0.163891f
C21318 DVDD.n18229 VSS 0.01831f
C21319 DVDD.n18230 VSS 0.11992f
C21320 DVDD.n18231 VSS 0.137328f
C21321 DVDD.n18232 VSS 0.202124f
C21322 DVDD.n18233 VSS 0.274656f
C21323 DVDD.n18234 VSS 0.274656f
C21324 DVDD.n18235 VSS 0.277343f
C21325 DVDD.n18236 VSS 0.795146f
C21326 DVDD.n18237 VSS 0.274656f
C21327 DVDD.n18238 VSS 0.274656f
C21328 DVDD.n18239 VSS 0.11992f
C21329 DVDD.n18240 VSS 0.151899f
C21330 DVDD.n18241 VSS 0.11992f
C21331 DVDD.n18242 VSS 0.11992f
C21332 DVDD.n18243 VSS 0.151899f
C21333 DVDD.n18244 VSS 0.034496f
C21334 DVDD.n18245 VSS 0.034496f
C21335 DVDD.n18246 VSS 0.015989f
C21336 DVDD.n18247 VSS 0.015989f
C21337 DVDD.n18248 VSS 0.11992f
C21338 DVDD.n18249 VSS 0.11992f
C21339 DVDD.n18250 VSS 0.015989f
C21340 DVDD.n18251 VSS 0.015989f
C21341 DVDD.n18252 VSS 0.01831f
C21342 DVDD.n18253 VSS 0.015989f
C21343 DVDD.n18254 VSS 0.036621f
C21344 DVDD.n18255 VSS 0.036964f
C21345 DVDD.n18256 VSS 0.015989f
C21346 DVDD.n18257 VSS 0.036621f
C21347 DVDD.n18258 VSS 0.037194f
C21348 DVDD.n18259 VSS 0.105852f
C21349 DVDD.n18260 VSS 0.036621f
C21350 DVDD.n18261 VSS 0.036621f
C21351 DVDD.n18262 VSS 0.02695f
C21352 DVDD.n18263 VSS 0.015989f
C21353 DVDD.n18264 VSS 0.11992f
C21354 DVDD.n18265 VSS 0.163891f
C21355 DVDD.n18266 VSS 0.163891f
C21356 DVDD.n18267 VSS 0.137328f
C21357 DVDD.n18268 VSS 0.01831f
C21358 DVDD.n18269 VSS 0.163891f
C21359 DVDD.n18270 VSS 0.124756f
C21360 DVDD.n18271 VSS 0.163891f
C21361 DVDD.n18272 VSS 0.132493f
C21362 DVDD.n18273 VSS 0.016634f
C21363 DVDD.n18274 VSS 0.01831f
C21364 DVDD.n18275 VSS 0.036621f
C21365 DVDD.n18276 VSS 0.015989f
C21366 DVDD.n18277 VSS 0.027981f
C21367 DVDD.n18278 VSS 0.036621f
C21368 DVDD.n18279 VSS 0.015989f
C21369 DVDD.n18280 VSS 0.319852f
C21370 DVDD.n18281 VSS 0.137328f
C21371 DVDD.n18282 VSS 0.325912f
C21372 DVDD.n18283 VSS 0.163891f
C21373 DVDD.n18284 VSS 0.132493f
C21374 DVDD.n18285 VSS 0.163891f
C21375 DVDD.n18286 VSS 0.124756f
C21376 DVDD.n18287 VSS 0.017666f
C21377 DVDD.n18288 VSS 0.036277f
C21378 DVDD.n18289 VSS 0.036621f
C21379 DVDD.n18290 VSS 0.027981f
C21380 DVDD.n18291 VSS 0.01831f
C21381 DVDD.n18292 VSS 0.015989f
C21382 DVDD.n18293 VSS 0.163891f
C21383 DVDD.n18294 VSS 0.137328f
C21384 DVDD.n18295 VSS 0.11992f
C21385 DVDD.n18296 VSS 0.163891f
C21386 DVDD.n18297 VSS 0.037455f
C21387 DVDD.n18298 VSS 0.163891f
C21388 DVDD.n18299 VSS 0.11992f
C21389 DVDD.n18300 VSS 0.11992f
C21390 DVDD.n18301 VSS 0.151899f
C21391 DVDD.n18302 VSS 0.034496f
C21392 DVDD.n18303 VSS 0.11992f
C21393 DVDD.n18304 VSS 0.015989f
C21394 DVDD.n18305 VSS 0.015989f
C21395 DVDD.n18306 VSS 0.11992f
C21396 DVDD.n18307 VSS 0.151899f
C21397 DVDD.n18308 VSS 0.039504f
C21398 DVDD.n18309 VSS 0.079009f
C21399 DVDD.n18310 VSS 0.06037f
C21400 DVDD.n18311 VSS 0.078141f
C21401 DVDD.n18312 VSS 0.034496f
C21402 DVDD.n18313 VSS 0.038113f
C21403 DVDD.n18314 VSS 0.151899f
C21404 DVDD.n18315 VSS 0.296448f
C21405 DVDD.n18316 VSS 0.11992f
C21406 DVDD.n18317 VSS 0.325912f
C21407 DVDD.n18318 VSS 0.274656f
C21408 DVDD.n18319 VSS 0.440997f
C21409 DVDD.n18320 VSS 0.209861f
C21410 DVDD.n18321 VSS 0.274656f
C21411 DVDD.n18322 VSS 0.274656f
C21412 DVDD.n18323 VSS 0.132493f
C21413 DVDD.n18324 VSS 0.11992f
C21414 DVDD.n18325 VSS 0.274656f
C21415 DVDD.n18326 VSS 0.274656f
C21416 DVDD.n18327 VSS 0.274656f
C21417 DVDD.n18328 VSS 0.274656f
C21418 DVDD.n18329 VSS 0.11992f
C21419 DVDD.n18330 VSS 0.11992f
C21420 DVDD.n18331 VSS 0.151899f
C21421 DVDD.n18332 VSS 0.151899f
C21422 DVDD.n18333 VSS 0.034496f
C21423 DVDD.n18334 VSS 0.039504f
C21424 DVDD.n18335 VSS 0.079009f
C21425 DVDD.n18336 VSS 0.06037f
C21426 DVDD.n18337 VSS 0.078195f
C21427 DVDD.n18338 VSS 0.038113f
C21428 DVDD.n18339 VSS 0.124756f
C21429 DVDD.n18340 VSS 0.151899f
C21430 DVDD.n18341 VSS 0.035888f
C21431 DVDD.n18342 VSS 0.034496f
C21432 DVDD.n18343 VSS 0.079009f
C21433 DVDD.n18344 VSS 0.074628f
C21434 DVDD.n18345 VSS 0.225253f
C21435 DVDD.n18346 VSS 0.079009f
C21436 DVDD.n18347 VSS 0.079009f
C21437 DVDD.n18348 VSS 0.034496f
C21438 DVDD.n18349 VSS 0.039504f
C21439 DVDD.n18350 VSS 0.151899f
C21440 DVDD.n18351 VSS 0.137328f
C21441 DVDD.n18352 VSS 0.11992f
C21442 DVDD.n18353 VSS 0.209861f
C21443 DVDD.n18354 VSS 0.274656f
C21444 DVDD.n18355 VSS 0.274656f
C21445 DVDD.n18356 VSS 0.274656f
C21446 DVDD.n18357 VSS 0.274656f
C21447 DVDD.n18358 VSS 0.274656f
C21448 DVDD.n18359 VSS 0.440997f
C21449 DVDD.n18360 VSS 0.440997f
C21450 DVDD.n18361 VSS 0.440997f
C21451 DVDD.n18362 VSS 0.325912f
C21452 DVDD.n18363 VSS 0.137328f
C21453 DVDD.n18364 VSS 0.296448f
C21454 DVDD.n18365 VSS 0.151899f
C21455 DVDD.n18366 VSS 0.035888f
C21456 DVDD.n18367 VSS 0.034496f
C21457 DVDD.n18368 VSS 0.079009f
C21458 DVDD.n18369 VSS 0.074683f
C21459 DVDD.n18370 VSS 0.225252f
C21460 DVDD.n18371 VSS 0.079009f
C21461 DVDD.n18372 VSS 0.079009f
C21462 DVDD.n18373 VSS 0.034496f
C21463 DVDD.n18374 VSS 0.039504f
C21464 DVDD.n18375 VSS 0.151899f
C21465 DVDD.n18376 VSS 0.137328f
C21466 DVDD.n18377 VSS 0.11992f
C21467 DVDD.n18378 VSS 0.034496f
C21468 DVDD.n18379 VSS 0.015989f
C21469 DVDD.n18380 VSS 0.015989f
C21470 DVDD.n18381 VSS 0.11992f
C21471 DVDD.n18382 VSS 0.163891f
C21472 DVDD.n18383 VSS 0.11992f
C21473 DVDD.n18384 VSS 0.163891f
C21474 DVDD.n18385 VSS 0.037455f
C21475 DVDD.n18386 VSS 0.151899f
C21476 DVDD.n18387 VSS 0.137328f
C21477 DVDD.n18388 VSS 0.042891f
C21478 DVDD.n18389 VSS 0.085784f
C21479 DVDD.n18390 VSS 0.085784f
C21480 DVDD.n18391 VSS 0.038361f
C21481 DVDD.n18392 VSS 0.229686f
C21482 DVDD.n18393 VSS 0.134427f
C21483 DVDD.n18394 VSS 0.122822f
C21484 DVDD.n18395 VSS 0.11992f
C21485 DVDD.n18396 VSS 0.163891f
C21486 DVDD.n18397 VSS 0.01831f
C21487 DVDD.n18398 VSS 0.137328f
C21488 DVDD.n18399 VSS 0.01831f
C21489 DVDD.n18400 VSS 0.137328f
C21490 DVDD.n18401 VSS 0.01831f
C21491 DVDD.n18402 VSS 0.11992f
C21492 DVDD.n18403 VSS 0.319852f
C21493 DVDD.n18404 VSS 0.134427f
C21494 DVDD.n18405 VSS 0.456471f
C21495 DVDD.n18406 VSS 0.274656f
C21496 DVDD.n18407 VSS 0.274656f
C21497 DVDD.n18408 VSS 0.122822f
C21498 DVDD.n18409 VSS 0.247819f
C21499 DVDD.n18410 VSS 0.081946f
C21500 DVDD.n18411 VSS 0.036964f
C21501 DVDD.n18412 VSS 0.037178f
C21502 DVDD.n18413 VSS 0.015989f
C21503 DVDD.n18414 VSS 0.015989f
C21504 DVDD.n18415 VSS 0.036621f
C21505 DVDD.n18416 VSS 0.02695f
C21506 DVDD.n18417 VSS 0.036621f
C21507 DVDD.n18418 VSS 0.105853f
C21508 DVDD.n18419 VSS 0.036621f
C21509 DVDD.n18420 VSS 0.036621f
C21510 DVDD.n18421 VSS 0.015989f
C21511 DVDD.n18422 VSS 0.016376f
C21512 DVDD.n18423 VSS 0.036979f
C21513 DVDD.n18424 VSS 0.319852f
C21514 DVDD.n18425 VSS 0.11992f
C21515 DVDD.n18426 VSS 0.153978f
C21516 DVDD.n18427 VSS 0.151899f
C21517 DVDD.n18428 VSS 0.075949f
C21518 DVDD.n18429 VSS 0.037455f
C21519 DVDD.n18430 VSS 0.085784f
C21520 DVDD.n18431 VSS 0.085784f
C21521 DVDD.n18432 VSS 0.743981f
C21522 DVDD.n18433 VSS 0.06037f
C21523 DVDD.n18434 VSS 0.058144f
C21524 DVDD.n18435 VSS 0.036621f
C21525 DVDD.n18436 VSS 0.015989f
C21526 DVDD.n18437 VSS 0.015989f
C21527 DVDD.n18438 VSS 0.01831f
C21528 DVDD.n18439 VSS 0.016376f
C21529 DVDD.n18440 VSS 0.015989f
C21530 DVDD.n18441 VSS 0.036621f
C21531 DVDD.n18442 VSS 0.037194f
C21532 DVDD.n18443 VSS 0.105852f
C21533 DVDD.n18444 VSS 0.036621f
C21534 DVDD.n18445 VSS 0.036621f
C21535 DVDD.n18446 VSS 0.02695f
C21536 DVDD.n18447 VSS 0.02695f
C21537 DVDD.n18448 VSS 0.027981f
C21538 DVDD.n18449 VSS 0.202124f
C21539 DVDD.n18450 VSS 0.209861f
C21540 DVDD.n18451 VSS 0.202124f
C21541 DVDD.n18452 VSS 0.202124f
C21542 DVDD.n18453 VSS 0.274656f
C21543 DVDD.n18454 VSS 0.274656f
C21544 DVDD.n18455 VSS 0.780268f
C21545 DVDD.n18456 VSS 0.274656f
C21546 DVDD.n18457 VSS 0.137328f
C21547 DVDD.n18458 VSS 0.163891f
C21548 DVDD.n18459 VSS 0.01831f
C21549 DVDD.n18460 VSS 0.11992f
C21550 DVDD.n18461 VSS 0.163891f
C21551 DVDD.n18462 VSS 0.124756f
C21552 DVDD.n18463 VSS 0.016634f
C21553 DVDD.n18464 VSS 0.01831f
C21554 DVDD.n18465 VSS 0.015989f
C21555 DVDD.n18466 VSS 0.036621f
C21556 DVDD.n18467 VSS 0.015989f
C21557 DVDD.n18468 VSS 0.027981f
C21558 DVDD.n18469 VSS 0.036621f
C21559 DVDD.n18470 VSS 0.035087f
C21560 DVDD.n18471 VSS 0.036621f
C21561 DVDD.n18472 VSS 0.103874f
C21562 DVDD.n18473 VSS 0.036621f
C21563 DVDD.n18474 VSS 0.015989f
C21564 DVDD.n18475 VSS 0.017666f
C21565 DVDD.n18476 VSS 0.124756f
C21566 DVDD.n18477 VSS 0.11992f
C21567 DVDD.n18478 VSS 0.037455f
C21568 DVDD.n18479 VSS 0.042891f
C21569 DVDD.n18480 VSS 0.151899f
C21570 DVDD.n18481 VSS 0.041382f
C21571 DVDD.n18482 VSS 0.151899f
C21572 DVDD.n18483 VSS 0.132493f
C21573 DVDD.n18484 VSS 0.163891f
C21574 DVDD.n18485 VSS 0.132493f
C21575 DVDD.n18486 VSS 0.274656f
C21576 DVDD.n18487 VSS 0.780268f
C21577 DVDD.n18488 VSS 0.274656f
C21578 DVDD.n18489 VSS 0.209861f
C21579 DVDD.n18490 VSS 0.274656f
C21580 DVDD.n18491 VSS 0.274656f
C21581 DVDD.n18492 VSS 0.11992f
C21582 DVDD.n18493 VSS 0.137328f
C21583 DVDD.n18494 VSS 0.163891f
C21584 DVDD.n18495 VSS 0.163891f
C21585 DVDD.n18496 VSS 0.137328f
C21586 DVDD.n18497 VSS 0.163891f
C21587 DVDD.n18498 VSS 0.137328f
C21588 DVDD.n18499 VSS 0.11992f
C21589 DVDD.n18500 VSS 0.274656f
C21590 DVDD.n18501 VSS 0.209861f
C21591 DVDD.n18502 VSS 0.209861f
C21592 DVDD.n18503 VSS 0.027981f
C21593 DVDD.n18504 VSS 0.202124f
C21594 DVDD.n18505 VSS 0.209861f
C21595 DVDD.n18506 VSS 0.02695f
C21596 DVDD.n18507 VSS 0.209861f
C21597 DVDD.n18508 VSS 0.274656f
C21598 DVDD.n18509 VSS 0.11992f
C21599 DVDD.n18510 VSS 0.11992f
C21600 DVDD.n18511 VSS 0.274656f
C21601 DVDD.n18512 VSS 0.456471f
C21602 DVDD.n18513 VSS 0.333649f
C21603 DVDD.n18514 VSS 0.333649f
C21604 DVDD.n18515 VSS 0.11992f
C21605 DVDD.n18516 VSS 0.274656f
C21606 DVDD.n18517 VSS 0.202124f
C21607 DVDD.n18518 VSS 0.137328f
C21608 DVDD.n18519 VSS 0.163891f
C21609 DVDD.n18520 VSS 0.137328f
C21610 DVDD.n18521 VSS 0.01831f
C21611 DVDD.n18522 VSS 0.036621f
C21612 DVDD.n18523 VSS 0.036979f
C21613 DVDD.n18524 VSS 0.016376f
C21614 DVDD.n18525 VSS 0.015989f
C21615 DVDD.n18526 VSS 0.163891f
C21616 DVDD.n18527 VSS 0.137328f
C21617 DVDD.n18528 VSS 0.11992f
C21618 DVDD.n18529 VSS 0.319852f
C21619 DVDD.n18530 VSS 0.247819f
C21620 DVDD.n18531 VSS 0.333649f
C21621 DVDD.n18532 VSS 0.122822f
C21622 DVDD.n18533 VSS 0.229686f
C21623 DVDD.n18534 VSS 0.151899f
C21624 DVDD.n18535 VSS 0.079206f
C21625 DVDD.n18536 VSS 0.039504f
C21626 DVDD.n18537 VSS 0.034496f
C21627 DVDD.n18538 VSS 0.039504f
C21628 DVDD.n18539 VSS 0.151899f
C21629 DVDD.n18540 VSS 0.11992f
C21630 DVDD.n18541 VSS 0.274656f
C21631 DVDD.n18542 VSS 0.456471f
C21632 DVDD.n18543 VSS 0.274656f
C21633 DVDD.n18544 VSS 0.333649f
C21634 DVDD.n18545 VSS 0.274656f
C21635 DVDD.n18546 VSS 0.202124f
C21636 DVDD.n18547 VSS 0.274656f
C21637 DVDD.n18548 VSS 0.137328f
C21638 DVDD.n18549 VSS 0.151899f
C21639 DVDD.n18550 VSS 0.11992f
C21640 DVDD.n18551 VSS 0.163891f
C21641 DVDD.n18552 VSS 0.153978f
C21642 DVDD.n18553 VSS 0.01831f
C21643 DVDD.n18554 VSS 0.11992f
C21644 DVDD.n18555 VSS 0.137328f
C21645 DVDD.n18556 VSS 0.163891f
C21646 DVDD.n18557 VSS 0.005071f
C21647 DVDD.n18558 VSS 0.005096f
C21648 DVDD.n18560 VSS 1.82078f
C21649 DVDD.n18561 VSS 0.006035f
C21650 DVDD.n18562 VSS 0.005096f
C21651 DVDD.n18564 VSS 0.006035f
C21652 DVDD.n18565 VSS 0.005096f
C21653 DVDD.n18567 VSS 0.006035f
C21654 DVDD.n18568 VSS 0.005096f
C21655 DVDD.n18570 VSS 0.006035f
C21656 DVDD.n18571 VSS 0.005096f
C21657 DVDD.n18573 VSS 0.006035f
C21658 DVDD.n18574 VSS 0.005096f
C21659 DVDD.n18576 VSS 0.006035f
C21660 DVDD.n18577 VSS 0.005096f
C21661 DVDD.n18579 VSS 0.006035f
C21662 DVDD.n18580 VSS 0.005096f
C21663 DVDD.n18582 VSS 0.006035f
C21664 DVDD.n18583 VSS 0.005096f
C21665 DVDD.n18585 VSS 0.006035f
C21666 DVDD.n18586 VSS 0.005096f
C21667 DVDD.n18588 VSS 0.006035f
C21668 DVDD.n18589 VSS 0.005096f
C21669 DVDD.n18591 VSS 0.006035f
C21670 DVDD.n18592 VSS 0.005096f
C21671 DVDD.n18594 VSS 0.006035f
C21672 DVDD.n18595 VSS 0.002548f
C21673 DVDD.n18597 VSS 0.003062f
C21674 DVDD.n18598 VSS 0.006035f
C21675 DVDD.n18599 VSS 0.005096f
C21676 DVDD.n18601 VSS 0.006035f
C21677 DVDD.n18602 VSS 0.005096f
C21678 DVDD.n18604 VSS 0.006035f
C21679 DVDD.n18605 VSS 0.005096f
C21680 DVDD.n18607 VSS 0.006035f
C21681 DVDD.n18608 VSS 0.005096f
C21682 DVDD.n18610 VSS 0.006035f
C21683 DVDD.n18611 VSS 0.002842f
C21684 DVDD.n18613 VSS 0.006035f
C21685 DVDD.n18614 VSS 0.002548f
C21686 DVDD.n18615 VSS 0.003008f
C21687 DVDD.n18616 VSS 0.011124f
C21688 DVDD.n18617 VSS 0.006035f
C21689 DVDD.n18618 VSS 0.006321f
C21690 DVDD.n18619 VSS 0.781602f
C21691 DVDD.n18620 VSS 0.006035f
C21692 DVDD.n18621 VSS 0.008791f
C21693 DVDD.n18622 VSS 0.005096f
C21694 DVDD.n18623 VSS 0.006035f
C21695 DVDD.n18624 VSS 0.923711f
C21696 DVDD.n18625 VSS 0.006035f
C21697 DVDD.n18626 VSS 0.005096f
C21698 DVDD.n18627 VSS 0.006035f
C21699 DVDD.t69 VSS 0.461856f
C21700 DVDD.n18628 VSS 0.006035f
C21701 DVDD.n18629 VSS 0.005096f
C21702 DVDD.n18630 VSS 0.006035f
C21703 DVDD.n18631 VSS 0.497383f
C21704 DVDD.n18632 VSS 0.006035f
C21705 DVDD.n18633 VSS 0.005096f
C21706 DVDD.n18634 VSS 0.006035f
C21707 DVDD.n18635 VSS 0.817129f
C21708 DVDD.t12 VSS 0.461856f
C21709 DVDD.n18636 VSS 0.006035f
C21710 DVDD.n18637 VSS 0.005096f
C21711 DVDD.n18638 VSS 0.006035f
C21712 DVDD.n18639 VSS 0.923711f
C21713 DVDD.n18640 VSS 0.006035f
C21714 DVDD.n18641 VSS 0.005096f
C21715 DVDD.n18642 VSS 0.006035f
C21716 DVDD.t66 VSS 0.461856f
C21717 DVDD.n18643 VSS 0.006035f
C21718 DVDD.n18644 VSS 0.005096f
C21719 DVDD.n18645 VSS 0.006035f
C21720 DVDD.n18646 VSS 0.53291f
C21721 DVDD.n18647 VSS 0.006035f
C21722 DVDD.n18648 VSS 0.002548f
C21723 DVDD.n18649 VSS 0.006035f
C21724 DVDD.n18650 VSS 0.852657f
C21725 DVDD.t13 VSS 0.461856f
C21726 DVDD.n18651 VSS 0.006035f
C21727 DVDD.n18652 VSS 0.003871f
C21728 DVDD.n18653 VSS 0.882607f
C21729 DVDD.n18654 VSS 0.151899f
C21730 DVDD.n18655 VSS 0.272424f
C21731 DVDD.n18656 VSS 0.074683f
C21732 DVDD.n18657 VSS 0.035888f
C21733 DVDD.n18658 VSS 0.034496f
C21734 DVDD.n18659 VSS 0.039504f
C21735 DVDD.n18660 VSS 0.151899f
C21736 DVDD.n18661 VSS 0.11992f
C21737 DVDD.n18662 VSS 0.163891f
C21738 DVDD.n18663 VSS 0.01831f
C21739 DVDD.n18664 VSS 0.11992f
C21740 DVDD.n18665 VSS 0.163891f
C21741 DVDD.n18666 VSS 0.132493f
C21742 DVDD.n18667 VSS 0.274656f
C21743 DVDD.n18668 VSS 0.209861f
C21744 DVDD.n18669 VSS 0.274656f
C21745 DVDD.n18670 VSS 0.11992f
C21746 DVDD.n18671 VSS 1.37721f
C21747 DVDD.n18674 VSS 0.064086f
C21748 DVDD.n18675 VSS 0.064086f
C21749 DVDD.n18676 VSS 0.064086f
C21750 DVDD.n18677 VSS 0.064086f
C21751 DVDD.n18678 VSS 0.064086f
C21752 DVDD.n18679 VSS 0.064086f
C21753 DVDD.n18681 VSS 0.064086f
C21754 DVDD.n18682 VSS 0.064086f
C21755 DVDD.n18683 VSS 0.064086f
C21756 DVDD.n18684 VSS 0.064086f
C21757 DVDD.n18685 VSS 0.111926f
C21758 DVDD.n18686 VSS 0.159926f
C21759 DVDD.n18687 VSS 0.163891f
C21760 DVDD.n18688 VSS 0.124901f
C21761 DVDD.n18689 VSS 0.163891f
C21762 DVDD.n18690 VSS 0.163891f
C21763 DVDD.n18691 VSS 0.055963f
C21764 DVDD.n18693 VSS 0.163891f
C21765 DVDD.n18694 VSS 0.120936f
C21766 DVDD.n18696 VSS 0.163891f
C21767 DVDD.n18698 VSS 0.163891f
C21768 DVDD.n18699 VSS 0.159926f
C21769 DVDD.n18700 VSS 0.063184f
C21770 DVDD.n18701 VSS 0.062281f
C21771 DVDD.n18702 VSS 0.064086f
C21772 DVDD.n18703 VSS 0.081946f
C21773 DVDD.n18708 VSS 0.057768f
C21774 DVDD.n18709 VSS 0.055963f
C21775 DVDD.n18710 VSS 0.128173f
C21776 DVDD.n18711 VSS 0.055963f
C21777 DVDD.n18712 VSS 0.128173f
C21778 DVDD.n18713 VSS 0.128173f
C21779 DVDD.n18714 VSS 0.128173f
C21780 DVDD.n18715 VSS 0.055963f
C21781 DVDD.n18716 VSS 0.128173f
C21782 DVDD.n18717 VSS 0.055963f
C21783 DVDD.n18718 VSS 0.128173f
C21784 DVDD.n18719 VSS 0.128173f
C21785 DVDD.n18720 VSS 0.074015f
C21786 DVDD.n18721 VSS 0.128173f
C21787 DVDD.n18722 VSS 0.128173f
C21788 DVDD.n18723 VSS 0.128173f
C21789 DVDD.n18724 VSS 0.159926f
C21790 DVDD.n18725 VSS 0.163891f
C21791 DVDD.n18726 VSS 0.124901f
C21792 DVDD.n18727 VSS 0.163891f
C21793 DVDD.n18728 VSS 0.163891f
C21794 DVDD.n18729 VSS 0.055963f
C21795 DVDD.n18730 VSS 1.37721f
C21796 DVDD.n18731 VSS 0.163891f
C21797 DVDD.n18732 VSS 0.120936f
C21798 DVDD.n18733 VSS 0.163891f
C21799 DVDD.n18734 VSS 0.163891f
C21800 DVDD.n18735 VSS 0.159926f
C21801 DVDD.n18736 VSS 0.064086f
C21802 DVDD.n18737 VSS 0.059573f
C21803 DVDD.n18738 VSS 0.064086f
C21804 DVDD.n18739 VSS 0.064086f
C21805 DVDD.n18740 VSS 0.064086f
C21806 DVDD.n18741 VSS 0.058671f
C21807 DVDD.n18742 VSS 0.064086f
C21808 DVDD.n18743 VSS 0.064086f
C21809 DVDD.n18751 VSS 0.075212f
C21810 DVDD.n18752 VSS 0.02942f
C21811 DVDD.n18753 VSS -1.02989f
C21812 DVDD.n18755 VSS 0.007995f
C21813 DVDD.n18756 VSS 0.015989f
C21814 DVDD.n18757 VSS 0.015989f
C21815 DVDD.n18758 VSS 0.015989f
C21816 DVDD.n18759 VSS 0.015989f
C21817 DVDD.n18760 VSS 0.015989f
C21818 DVDD.n18761 VSS 0.007995f
C21819 DVDD.n18762 VSS 0.040554f
C21820 DVDD.n18763 VSS 0.58221f
C21821 DVDD.n18764 VSS 0.015989f
C21822 DVDD.n18765 VSS 0.015989f
C21823 DVDD.n18766 VSS 0.015989f
C21824 DVDD.n18767 VSS 0.015989f
C21825 DVDD.n18768 VSS 0.015989f
C21826 DVDD.n18769 VSS 0.015989f
C21827 DVDD.n18770 VSS 0.617235f
C21828 DVDD.n18771 VSS 0.015989f
C21829 DVDD.n18773 VSS 0.015989f
C21830 DVDD.n18774 VSS 0.007995f
C21831 DVDD.n18775 VSS 0.015989f
C21832 DVDD.n18776 VSS 0.015989f
C21833 DVDD.n18777 VSS 0.015989f
C21834 DVDD.n18778 VSS 0.015989f
C21835 DVDD.n18779 VSS 0.015989f
C21836 DVDD.n18780 VSS 0.015989f
C21837 DVDD.n18781 VSS 0.015989f
C21838 DVDD.n18782 VSS 0.015989f
C21839 DVDD.n18783 VSS 0.015989f
C21840 DVDD.n18784 VSS 0.015989f
C21841 DVDD.n18785 VSS 0.015989f
C21842 DVDD.n18786 VSS 0.007995f
C21843 DVDD.n18787 VSS 0.02942f
C21844 DVDD.n18788 VSS 0.02942f
C21845 DVDD.n18789 VSS 0.02942f
C21846 DVDD.n18790 VSS 0.02942f
C21847 DVDD.n18791 VSS 0.02942f
C21848 DVDD.n18792 VSS 0.02942f
C21849 DVDD.n18794 VSS 0.02942f
C21850 DVDD.n18797 VSS 0.02942f
C21851 DVDD.n18799 VSS 0.064891f
C21852 DVDD.n18801 VSS 0.02942f
C21853 DVDD.n18804 VSS 0.02942f
C21854 DVDD.n18807 VSS 0.02942f
C21855 DVDD.n18810 VSS 0.02942f
C21856 DVDD.n18813 VSS 0.02942f
C21857 DVDD.n18816 VSS 0.02942f
C21858 DVDD.n18819 VSS 0.561072f
C21859 DVDD.n18820 VSS 0.319382f
C21860 DVDD.n18821 VSS 1.35823f
C21861 DVDD.n18822 VSS 0.319382f
C21862 DVDD.n18825 VSS 0.007995f
C21863 DVDD.n18826 VSS 0.015989f
C21864 DVDD.n18827 VSS 0.015989f
C21865 DVDD.n18828 VSS 0.007995f
C21866 DVDD.n18829 VSS 0.081946f
C21867 DVDD.n18830 VSS 0.066473f
C21868 DVDD.n18832 VSS 0.064086f
C21869 DVDD.n18833 VSS 0.064086f
C21870 DVDD.n18834 VSS 0.064086f
C21871 DVDD.n18835 VSS 0.056865f
C21872 DVDD.n18836 VSS 0.064086f
C21873 DVDD.n18837 VSS 0.064086f
C21874 DVDD.n18838 VSS 0.064086f
C21875 DVDD.n18839 VSS 0.064086f
C21876 DVDD.n18840 VSS 0.064086f
C21877 DVDD.n18842 VSS 0.063184f
C21878 DVDD.n18843 VSS 0.064086f
C21879 DVDD.n18844 VSS 0.064086f
C21880 DVDD.n18845 VSS 0.064086f
C21881 DVDD.n18846 VSS 0.062281f
C21882 DVDD.n18847 VSS 0.055963f
C21883 DVDD.n18848 VSS 0.08525f
C21884 DVDD.n18850 VSS 0.163891f
C21885 DVDD.n18851 VSS 0.163891f
C21886 DVDD.n18852 VSS 0.163891f
C21887 DVDD.n18853 VSS 0.074015f
C21888 DVDD.n18855 VSS 0.163891f
C21889 DVDD.n18857 VSS 0.163891f
C21890 DVDD.n18858 VSS 0.160587f
C21891 DVDD.n18859 VSS 0.45004f
C21892 DVDD.n18860 VSS 0.096137f
C21893 DVDD.n18865 VSS 0.057768f
C21894 DVDD.n18866 VSS 0.081946f
C21895 DVDD.n18867 VSS 0.081946f
C21896 DVDD.n18868 VSS 0.081946f
C21897 DVDD.n18869 VSS 0.081946f
C21898 DVDD.n18870 VSS 0.096197f
C21899 DVDD.n18871 VSS 0.08525f
C21900 DVDD.n18872 VSS 0.059573f
C21901 DVDD.n18873 VSS 0.064086f
C21902 DVDD.n18874 VSS 0.064086f
C21903 DVDD.n18875 VSS 0.064086f
C21904 DVDD.n18876 VSS 0.064086f
C21905 DVDD.n18877 VSS 0.064086f
C21906 DVDD.n18878 VSS 0.064086f
C21907 DVDD.n18879 VSS 0.058671f
C21908 DVDD.n18880 VSS 0.061379f
C21909 DVDD.n18881 VSS 0.064086f
C21910 DVDD.n18882 VSS 0.064086f
C21911 DVDD.n18883 VSS 0.064086f
C21912 DVDD.n18884 VSS 0.064086f
C21913 DVDD.n18885 VSS 0.064086f
C21914 DVDD.n18886 VSS 0.060476f
C21915 DVDD.n18887 VSS 0.075821f
C21916 DVDD.n18889 VSS 0.163891f
C21917 DVDD.n18890 VSS 0.163891f
C21918 DVDD.n18891 VSS 0.163891f
C21919 DVDD.n18892 VSS 0.128866f
C21920 DVDD.n18893 VSS 0.055963f
C21921 DVDD.n18896 VSS 0.081946f
C21922 DVDD.n18899 VSS 0.163891f
C21923 DVDD.n18902 VSS 0.163891f
C21924 DVDD.n18904 VSS 0.160587f
C21925 DVDD.n18906 VSS 0.091557f
C21926 DVDD.n18907 VSS 0.040554f
C21927 DVDD.n18908 VSS 0.163891f
C21928 DVDD.n18909 VSS 0.075212f
C21929 DVDD.n18917 VSS 0.02942f
C21930 DVDD.n18919 VSS 0.163891f
C21931 DVDD.n18920 VSS 0.115237f
C21932 DVDD.n18921 VSS 0.079947f
C21933 DVDD.n18922 VSS 0.115237f
C21934 DVDD.n18923 VSS 0.115237f
C21935 DVDD.n18924 VSS 0.079947f
C21936 DVDD.n18925 VSS 0.151899f
C21937 DVDD.n18926 VSS 0.079947f
C21938 DVDD.n18927 VSS 0.109637f
C21939 DVDD.n18928 VSS 0.079947f
C21940 DVDD.n18929 VSS 0.075949f
C21941 DVDD.n18930 VSS 0.058219f
C21942 DVDD.n18931 VSS 0.064086f
C21943 DVDD.n18932 VSS 0.064086f
C21944 DVDD.n18933 VSS 0.064086f
C21945 DVDD.n18934 VSS 0.057317f
C21946 DVDD.n18935 VSS 0.064086f
C21947 DVDD.n18936 VSS 0.064086f
C21948 DVDD.n18937 VSS 0.075949f
C21949 DVDD.n18938 VSS 0.064086f
C21950 DVDD.n18939 VSS 0.064086f
C21951 DVDD.n18940 VSS 0.062732f
C21952 DVDD.n18941 VSS 0.064086f
C21953 DVDD.n18942 VSS 0.064086f
C21954 DVDD.n18943 VSS 0.05145f
C21955 DVDD.n18944 VSS 0.06183f
C21956 DVDD.n18945 VSS 0.055963f
C21957 DVDD.n18946 VSS 0.075949f
C21958 DVDD.n18947 VSS 0.075949f
C21959 DVDD.n18948 VSS 0.075949f
C21960 DVDD.n18949 VSS 0.075949f
C21961 DVDD.n18950 VSS 0.35687f
C21962 DVDD.n18953 VSS 0.075949f
C21963 DVDD.n18954 VSS 0.075949f
C21964 DVDD.n18955 VSS 0.075949f
C21965 DVDD.n18956 VSS 0.075949f
C21966 DVDD.n18957 VSS 0.079947f
C21967 DVDD.n18958 VSS 0.151899f
C21968 DVDD.n18959 VSS 0.079947f
C21969 DVDD.n18961 VSS 0.064086f
C21970 DVDD.n18962 VSS 0.064086f
C21971 DVDD.n18963 VSS 0.057317f
C21972 DVDD.n18964 VSS 0.064086f
C21973 DVDD.n18965 VSS 0.064086f
C21974 DVDD.n18966 VSS 0.064086f
C21975 DVDD.n18967 VSS 0.064086f
C21976 DVDD.n18968 VSS 0.062732f
C21977 DVDD.n18969 VSS 0.064086f
C21978 DVDD.n18970 VSS 0.064086f
C21979 DVDD.n18971 VSS 0.05145f
C21980 DVDD.n18973 VSS 0.055963f
C21981 DVDD.n18974 VSS 0.151899f
C21982 DVDD.n18975 VSS 0.151899f
C21983 DVDD.n18976 VSS 0.151899f
C21984 DVDD.n18977 VSS 0.151899f
C21985 DVDD.n18978 VSS 0.151899f
C21986 DVDD.n18979 VSS 0.35687f
C21987 DVDD.n18981 VSS 1.27644f
C21988 DVDD.n18982 VSS 0.151899f
C21989 DVDD.n18983 VSS 0.151899f
C21990 DVDD.n18984 VSS 0.151899f
C21991 DVDD.n18989 VSS 0.058219f
C21992 DVDD.n18995 VSS 0.064086f
C21993 DVDD.n18996 VSS 0.026627f
C21994 DVDD.n18997 VSS 0.076723f
C21995 DVDD.n18998 VSS 0.159414f
C21996 DVDD.n18999 VSS 0.128173f
C21997 DVDD.n19000 VSS 0.055963f
C21998 DVDD.n19001 VSS 0.128173f
C21999 DVDD.n19002 VSS 0.128173f
C22000 DVDD.n19003 VSS 0.055963f
C22001 DVDD.n19004 VSS 0.128173f
C22002 DVDD.n19005 VSS 0.128173f
C22003 DVDD.n19006 VSS 0.128173f
C22004 DVDD.n19007 VSS 0.128173f
C22005 DVDD.n19008 VSS 0.128173f
C22006 DVDD.n19009 VSS 0.128173f
C22007 DVDD.n19010 VSS 0.055963f
C22008 DVDD.n19011 VSS 0.128173f
C22009 DVDD.n19012 VSS 0.128173f
C22010 DVDD.n19013 VSS 0.055963f
C22011 DVDD.n19014 VSS 0.128173f
C22012 DVDD.n19015 VSS 0.128173f
C22013 DVDD.n19016 VSS 0.055963f
C22014 DVDD.n19017 VSS 0.128173f
C22015 DVDD.n19018 VSS 0.128173f
C22016 DVDD.n19019 VSS 0.128173f
C22017 DVDD.n19020 VSS 0.128173f
C22018 DVDD.n19021 VSS 0.128173f
C22019 DVDD.n19022 VSS 0.055963f
C22020 DVDD.n19023 VSS 0.163891f
C22021 DVDD.n19024 VSS 0.081946f
C22022 DVDD.n19025 VSS 0.163891f
C22023 DVDD.n19026 VSS 0.163891f
C22024 DVDD.n19027 VSS 0.128866f
C22025 DVDD.n19028 VSS 0.081946f
C22026 DVDD.n19029 VSS 0.163891f
C22027 DVDD.n19030 VSS 0.163891f
C22028 DVDD.n19031 VSS 0.160587f
C22029 DVDD.n19032 VSS 0.08525f
C22030 DVDD.n19033 VSS 0.45004f
C22031 DVDD.n19035 VSS 0.057768f
C22032 DVDD.n19036 VSS 0.064086f
C22033 DVDD.n19037 VSS 0.064086f
C22034 DVDD.n19038 VSS 0.064086f
C22035 DVDD.n19039 VSS 0.056865f
C22036 DVDD.n19040 VSS 0.064086f
C22037 DVDD.n19045 VSS 0.064086f
C22038 DVDD.n19046 VSS 0.064086f
C22039 DVDD.n19048 VSS 0.063184f
C22040 DVDD.n19049 VSS 0.064086f
C22041 DVDD.n19050 VSS 0.064086f
C22042 DVDD.n19051 VSS 0.064086f
C22043 DVDD.n19053 VSS 0.062281f
C22044 DVDD.n19054 VSS 0.055963f
C22045 DVDD.n19057 VSS 0.064086f
C22046 DVDD.n19058 VSS 0.128173f
C22047 DVDD.n19059 VSS 0.128173f
C22048 DVDD.n19060 VSS 0.128173f
C22049 DVDD.n19061 VSS 0.055963f
C22050 DVDD.n19062 VSS 0.128173f
C22051 DVDD.n19063 VSS 0.128173f
C22052 DVDD.n19064 VSS 0.055963f
C22053 DVDD.n19065 VSS 0.128173f
C22054 DVDD.n19066 VSS 0.128173f
C22055 DVDD.n19067 VSS 0.128173f
C22056 DVDD.n19068 VSS 0.128173f
C22057 DVDD.n19069 VSS 0.128173f
C22058 DVDD.n19070 VSS 0.128173f
C22059 DVDD.n19071 VSS 0.128173f
C22060 DVDD.n19072 VSS 0.128173f
C22061 DVDD.n19073 VSS 0.055963f
C22062 DVDD.n19074 VSS 0.163891f
C22063 DVDD.n19075 VSS 0.081946f
C22064 DVDD.n19076 VSS 0.163891f
C22065 DVDD.n19077 VSS 0.163891f
C22066 DVDD.n19078 VSS 0.128866f
C22067 DVDD.n19079 VSS 0.007995f
C22068 DVDD.n19080 VSS 0.015989f
C22069 DVDD.n19081 VSS 0.015989f
C22070 DVDD.n19082 VSS 0.015989f
C22071 DVDD.n19083 VSS 0.015989f
C22072 DVDD.n19084 VSS 0.015989f
C22073 DVDD.n19085 VSS 0.015989f
C22074 DVDD.n19086 VSS 0.015989f
C22075 DVDD.n19087 VSS 0.015989f
C22076 DVDD.n19088 VSS 0.015989f
C22077 DVDD.n19089 VSS 0.015989f
C22078 DVDD.n19090 VSS 0.015989f
C22079 DVDD.n19091 VSS 0.015989f
C22080 DVDD.n19092 VSS 0.015989f
C22081 DVDD.n19093 VSS 0.007995f
C22082 DVDD.n19094 VSS 0.081946f
C22083 DVDD.n19095 VSS 0.58221f
C22084 DVDD.n19097 VSS 0.091557f
C22085 DVDD.n19098 VSS 0.040554f
C22086 DVDD.n19099 VSS 0.040896f
C22087 DVDD.n19100 VSS 0.040554f
C22088 DVDD.n19101 VSS 0.625132f
C22089 DVDD.n19102 VSS 0.596461f
C22090 DVDD.n19103 VSS 0.096137f
C22091 DVDD.n19104 VSS 0.13448f
C22092 DVDD.n19105 VSS 0.066473f
C22093 DVDD.n19106 VSS 0.007995f
C22094 DVDD.n19107 VSS 0.015989f
C22095 DVDD.n19108 VSS 0.015989f
C22096 DVDD.n19109 VSS 0.015989f
C22097 DVDD.n19110 VSS 0.015989f
C22098 DVDD.n19111 VSS 0.015989f
C22099 DVDD.n19112 VSS 0.015989f
C22100 DVDD.n19113 VSS 0.015989f
C22101 DVDD.n19114 VSS 0.015989f
C22102 DVDD.n19115 VSS 0.015989f
C22103 DVDD.n19116 VSS 0.015989f
C22104 DVDD.n19117 VSS 0.015989f
C22105 DVDD.n19118 VSS 0.015989f
C22106 DVDD.n19119 VSS 0.015989f
C22107 DVDD.n19120 VSS 0.007995f
C22108 DVDD.n19121 VSS 0.035267f
C22109 DVDD.t159 VSS 1.03157f
C22110 DVDD.n19122 VSS 0.035267f
C22111 DVDD.n19123 VSS 0.081946f
C22112 DVDD.n19124 VSS 0.081946f
C22113 DVDD.n19125 VSS 0.163891f
C22114 DVDD.n19126 VSS 0.163891f
C22115 DVDD.n19127 VSS 0.160587f
C22116 DVDD.n19128 VSS 0.08525f
C22117 DVDD.n19129 VSS 0.45004f
C22118 DVDD.n19134 VSS 0.061379f
C22119 DVDD.n19135 VSS 0.064086f
C22120 DVDD.n19136 VSS 0.064086f
C22121 DVDD.n19137 VSS 0.064086f
C22122 DVDD.n19138 VSS 0.060476f
C22123 DVDD.n19139 VSS 0.064086f
C22124 DVDD.n19140 VSS 0.064086f
C22125 DVDD.n19141 VSS 0.064086f
C22126 DVDD.n19143 VSS 0.059573f
C22127 DVDD.n19144 VSS 0.064086f
C22128 DVDD.n19145 VSS 0.064086f
C22129 DVDD.n19146 VSS 0.064086f
C22130 DVDD.n19148 VSS 0.058671f
C22131 DVDD.n19149 VSS 0.055963f
C22132 DVDD.n19153 VSS 0.064086f
C22133 DVDD.n19154 VSS 0.128173f
C22134 DVDD.n19155 VSS 0.128173f
C22135 DVDD.n19156 VSS 0.128173f
C22136 DVDD.n19157 VSS 0.055963f
C22137 DVDD.n19158 VSS 0.128173f
C22138 DVDD.n19159 VSS 0.128173f
C22139 DVDD.n19160 VSS 0.055963f
C22140 DVDD.n19161 VSS 0.128173f
C22141 DVDD.n19162 VSS 0.128173f
C22142 DVDD.n19163 VSS 0.128173f
C22143 DVDD.n19164 VSS 0.128173f
C22144 DVDD.n19165 VSS 0.128173f
C22145 DVDD.n19166 VSS 0.128173f
C22146 DVDD.n19167 VSS 0.055963f
C22147 DVDD.n19168 VSS 0.128173f
C22148 DVDD.n19169 VSS 0.128173f
C22149 DVDD.n19170 VSS 0.055963f
C22150 DVDD.n19171 VSS 0.128173f
C22151 DVDD.n19172 VSS 0.128173f
C22152 DVDD.n19173 VSS 0.055963f
C22153 DVDD.n19174 VSS 0.128173f
C22154 DVDD.n19175 VSS 0.128173f
C22155 DVDD.n19176 VSS 0.128173f
C22156 DVDD.n19177 VSS 0.128173f
C22157 DVDD.n19178 VSS 0.128173f
C22158 DVDD.n19179 VSS 0.128173f
C22159 DVDD.n19180 VSS 0.128173f
C22160 DVDD.n19181 VSS 0.055963f
C22161 DVDD.n19182 VSS 0.151899f
C22162 DVDD.n19183 VSS 0.151899f
C22163 DVDD.n19184 VSS 0.151899f
C22164 DVDD.n19185 VSS 0.151899f
C22165 DVDD.n19186 VSS 0.151899f
C22166 DVDD.n19188 VSS 0.064086f
C22167 DVDD.n19189 VSS 0.059122f
C22168 DVDD.n19190 VSS 0.064086f
C22169 DVDD.n19191 VSS 0.064086f
C22170 DVDD.n19192 VSS 0.064086f
C22171 DVDD.n19193 VSS 0.060025f
C22172 DVDD.n19194 VSS 0.374251f
C22173 DVDD.n19195 VSS 0.060025f
C22174 DVDD.n19196 VSS 0.064086f
C22175 DVDD.n19197 VSS 0.064086f
C22176 DVDD.n19198 VSS 0.064086f
C22177 DVDD.n19199 VSS 0.060927f
C22178 DVDD.n19200 VSS 0.064086f
C22179 DVDD.n19201 VSS 0.055963f
C22180 DVDD.n19203 VSS 0.151899f
C22181 DVDD.n19204 VSS 0.151899f
C22182 DVDD.n19205 VSS 0.151899f
C22183 DVDD.n19206 VSS 0.151899f
C22184 DVDD.n19207 VSS 0.101545f
C22185 DVDD.n19210 VSS 0.115762f
C22186 DVDD.n19212 VSS 0.151899f
C22187 DVDD.n19214 VSS 0.151899f
C22188 DVDD.n19215 VSS 0.003332f
C22189 DVDD.n19216 VSS 0.005096f
C22190 DVDD.n19218 VSS 1.82078f
C22191 DVDD.n19219 VSS 0.006035f
C22192 DVDD.n19220 VSS 0.005096f
C22193 DVDD.n19222 VSS 0.006035f
C22194 DVDD.n19223 VSS 0.005096f
C22195 DVDD.n19225 VSS 0.006035f
C22196 DVDD.n19226 VSS 0.005096f
C22197 DVDD.n19228 VSS 0.006035f
C22198 DVDD.n19229 VSS 0.005096f
C22199 DVDD.n19231 VSS 0.006035f
C22200 DVDD.n19232 VSS 0.003062f
C22201 DVDD.n19234 VSS 0.006035f
C22202 DVDD.n19235 VSS 0.081946f
C22203 DVDD.n19236 VSS 0.002548f
C22204 DVDD.n19237 VSS 0.005096f
C22205 DVDD.n19239 VSS 0.006035f
C22206 DVDD.n19240 VSS 0.005096f
C22207 DVDD.n19242 VSS 0.006035f
C22208 DVDD.n19243 VSS 0.005096f
C22209 DVDD.n19245 VSS 0.006035f
C22210 DVDD.n19246 VSS 0.005096f
C22211 DVDD.n19248 VSS 0.006035f
C22212 DVDD.n19249 VSS 0.005096f
C22213 DVDD.n19251 VSS 0.006035f
C22214 DVDD.n19252 VSS 0.005096f
C22215 DVDD.n19254 VSS 0.006035f
C22216 DVDD.n19255 VSS 0.005096f
C22217 DVDD.n19257 VSS 0.006035f
C22218 DVDD.n19258 VSS 0.005096f
C22219 DVDD.n19260 VSS 0.006035f
C22220 DVDD.n19261 VSS 0.005096f
C22221 DVDD.n19263 VSS 0.006035f
C22222 DVDD.n19264 VSS 0.005096f
C22223 DVDD.n19266 VSS 0.006035f
C22224 DVDD.n19267 VSS 0.005096f
C22225 DVDD.n19269 VSS 0.006035f
C22226 DVDD.n19270 VSS 0.005096f
C22227 DVDD.n19272 VSS 0.006035f
C22228 DVDD.n19273 VSS 0.005096f
C22229 DVDD.n19275 VSS 0.006035f
C22230 DVDD.n19276 VSS 0.005096f
C22231 DVDD.n19278 VSS 0.006035f
C22232 DVDD.n19279 VSS 0.005096f
C22233 DVDD.n19281 VSS 0.006035f
C22234 DVDD.n19282 VSS 0.005096f
C22235 DVDD.n19284 VSS 0.006035f
C22236 DVDD.n19285 VSS 0.005096f
C22237 DVDD.n19287 VSS 0.006035f
C22238 DVDD.n19288 VSS 0.081946f
C22239 DVDD.n19289 VSS 0.002548f
C22240 DVDD.n19291 VSS 0.003062f
C22241 DVDD.n19292 VSS 0.006035f
C22242 DVDD.n19293 VSS 0.005096f
C22243 DVDD.n19295 VSS 0.006035f
C22244 DVDD.n19296 VSS 0.005096f
C22245 DVDD.n19298 VSS 0.006035f
C22246 DVDD.n19299 VSS 0.005096f
C22247 DVDD.n19301 VSS 0.006035f
C22248 DVDD.n19302 VSS 0.005096f
C22249 DVDD.n19304 VSS 0.006035f
C22250 DVDD.n19305 VSS 0.005096f
C22251 DVDD.n19307 VSS 0.006035f
C22252 DVDD.n19308 VSS 0.005096f
C22253 DVDD.n19310 VSS 0.006035f
C22254 DVDD.t64 VSS 0.008576f
C22255 DVDD.n19311 VSS 0.005096f
C22256 DVDD.n19313 VSS 0.005096f
C22257 DVDD.n19314 VSS 0.006035f
C22258 DVDD.n19315 VSS 0.005629f
C22259 DVDD.t63 VSS 0.461856f
C22260 DVDD.n19316 VSS 0.006035f
C22261 DVDD.n19317 VSS 0.005096f
C22262 DVDD.n19318 VSS 0.006035f
C22263 DVDD.n19319 VSS 0.005096f
C22264 DVDD.n19321 VSS 0.006035f
C22265 DVDD.n19322 VSS 0.005096f
C22266 DVDD.n19323 VSS 0.006035f
C22267 DVDD.n19325 VSS 0.006035f
C22268 DVDD.n19326 VSS 0.006035f
C22269 DVDD.n19327 VSS 0.005096f
C22270 DVDD.n19328 VSS 0.005096f
C22271 DVDD.n19329 VSS 0.005096f
C22272 DVDD.n19330 VSS 0.006035f
C22273 DVDD.n19332 VSS 0.006035f
C22274 DVDD.n19333 VSS 0.005629f
C22275 DVDD.n19334 VSS 0.007288f
C22276 DVDD.n19335 VSS 0.00555f
C22277 DVDD.n19336 VSS 0.005096f
C22278 DVDD.n19337 VSS 0.006035f
C22279 DVDD.n19338 VSS 0.603965f
C22280 DVDD.n19339 VSS 0.006035f
C22281 DVDD.n19340 VSS 0.006035f
C22282 DVDD.n19341 VSS 0.006035f
C22283 DVDD.n19342 VSS 0.923711f
C22284 DVDD.n19343 VSS 0.006035f
C22285 DVDD.n19344 VSS 0.005096f
C22286 DVDD.n19345 VSS 0.006035f
C22287 DVDD.n19346 VSS 0.006035f
C22288 DVDD.n19347 VSS 0.006035f
C22289 DVDD.n19348 VSS 0.006035f
C22290 DVDD.t70 VSS 0.461856f
C22291 DVDD.n19349 VSS 0.006035f
C22292 DVDD.n19350 VSS 0.005096f
C22293 DVDD.n19351 VSS 0.006035f
C22294 DVDD.n19352 VSS 0.568438f
C22295 DVDD.n19353 VSS 0.006035f
C22296 DVDD.n19354 VSS 0.006035f
C22297 DVDD.n19355 VSS 0.006035f
C22298 DVDD.n19356 VSS 0.923711f
C22299 DVDD.n19357 VSS 0.006035f
C22300 DVDD.n19358 VSS 0.006035f
C22301 DVDD.n19359 VSS 0.006035f
C22302 DVDD.n19360 VSS 0.005096f
C22303 DVDD.n19361 VSS 0.005096f
C22304 DVDD.n19362 VSS 0.005096f
C22305 DVDD.n19363 VSS 0.005096f
C22306 DVDD.n19364 VSS 0.006035f
C22307 DVDD.n19365 VSS 0.005096f
C22308 DVDD.n19366 VSS 0.005096f
C22309 DVDD.n19367 VSS 0.005096f
C22310 DVDD.n19368 VSS 0.005096f
C22311 DVDD.n19369 VSS 0.006035f
C22312 DVDD.n19370 VSS 0.005096f
C22313 DVDD.n19371 VSS 0.005096f
C22314 DVDD.n19372 VSS 0.005096f
C22315 DVDD.n19373 VSS 0.005096f
C22316 DVDD.n19374 VSS 0.005096f
C22317 DVDD.n19375 VSS 0.003871f
C22318 DVDD.n19376 VSS 0.005096f
C22319 DVDD.n19377 VSS 0.006035f
C22320 DVDD.t72 VSS 0.461856f
C22321 DVDD.n19378 VSS 0.53291f
C22322 DVDD.n19379 VSS 0.006035f
C22323 DVDD.n19380 VSS 0.005096f
C22324 DVDD.n19381 VSS 0.005096f
C22325 DVDD.n19382 VSS 0.005096f
C22326 DVDD.n19383 VSS 0.006035f
C22327 DVDD.n19384 VSS 0.710547f
C22328 DVDD.t67 VSS 0.461856f
C22329 DVDD.n19385 VSS 0.67502f
C22330 DVDD.n19386 VSS 0.923711f
C22331 DVDD.n19387 VSS 0.006035f
C22332 DVDD.n19388 VSS 0.005096f
C22333 DVDD.n19389 VSS 0.005096f
C22334 DVDD.n19390 VSS 0.005096f
C22335 DVDD.n19391 VSS 0.006035f
C22336 DVDD.n19392 VSS 0.817129f
C22337 DVDD.n19393 VSS 0.888184f
C22338 DVDD.t68 VSS 0.461856f
C22339 DVDD.n19394 VSS 0.497383f
C22340 DVDD.n19395 VSS 0.006035f
C22341 DVDD.n19396 VSS 0.005096f
C22342 DVDD.n19397 VSS 0.005096f
C22343 DVDD.n19398 VSS 0.005096f
C22344 DVDD.n19399 VSS 0.006035f
C22345 DVDD.n19400 VSS 0.746075f
C22346 DVDD.t62 VSS 0.461856f
C22347 DVDD.n19401 VSS 0.639492f
C22348 DVDD.n19402 VSS 0.923711f
C22349 DVDD.n19403 VSS 0.006035f
C22350 DVDD.n19404 VSS 0.005096f
C22351 DVDD.n19405 VSS 0.005096f
C22352 DVDD.n19406 VSS 0.005096f
C22353 DVDD.n19407 VSS 0.006035f
C22354 DVDD.n19408 VSS 0.781602f
C22355 DVDD.n19409 VSS 1.14576f
C22356 DVDD.n19410 VSS 0.005629f
C22357 DVDD.n19411 VSS 0.00555f
C22358 DVDD.n19412 VSS 0.008797f
C22359 DVDD.n19413 VSS 0.00412f
C22360 DVDD.n19414 VSS 0.006035f
C22361 DVDD.n19415 VSS 0.006035f
C22362 DVDD.n19416 VSS 0.005096f
C22363 DVDD.n19417 VSS 0.011056f
C22364 DVDD.n19418 VSS 0.002989f
C22365 DVDD.n19419 VSS 0.006035f
C22366 DVDD.n19421 VSS 0.006035f
C22367 DVDD.n19422 VSS 0.006035f
C22368 DVDD.n19423 VSS 0.005096f
C22369 DVDD.n19424 VSS 0.00365f
C22370 DVDD.n19425 VSS 0.002548f
C22371 DVDD.n19426 VSS 0.003993f
C22372 DVDD.n19427 VSS 0.006035f
C22373 DVDD.n19429 VSS 0.006035f
C22374 DVDD.n19430 VSS 0.006035f
C22375 DVDD.n19431 VSS 0.005096f
C22376 DVDD.n19432 VSS 0.005096f
C22377 DVDD.n19433 VSS 0.005096f
C22378 DVDD.n19434 VSS 0.006035f
C22379 DVDD.n19436 VSS 0.006035f
C22380 DVDD.n19437 VSS 0.006035f
C22381 DVDD.n19438 VSS 0.005096f
C22382 DVDD.n19439 VSS 0.005096f
C22383 DVDD.n19440 VSS 0.005096f
C22384 DVDD.n19441 VSS 0.006035f
C22385 DVDD.n19443 VSS 0.006035f
C22386 DVDD.n19444 VSS 0.006035f
C22387 DVDD.n19445 VSS 0.005096f
C22388 DVDD.n19446 VSS 0.005096f
C22389 DVDD.n19447 VSS 0.005096f
C22390 DVDD.n19448 VSS 0.006035f
C22391 DVDD.n19450 VSS 0.006035f
C22392 DVDD.n19451 VSS 0.006035f
C22393 DVDD.n19452 VSS 0.005096f
C22394 DVDD.n19453 VSS 0.005096f
C22395 DVDD.n19454 VSS 0.005096f
C22396 DVDD.n19455 VSS 0.006035f
C22397 DVDD.n19457 VSS 0.006035f
C22398 DVDD.n19458 VSS 0.006035f
C22399 DVDD.n19459 VSS 0.005096f
C22400 DVDD.n19460 VSS 0.005096f
C22401 DVDD.n19461 VSS 0.005096f
C22402 DVDD.n19462 VSS 0.006035f
C22403 DVDD.n19464 VSS 0.006035f
C22404 DVDD.n19465 VSS 0.006035f
C22405 DVDD.n19466 VSS 0.004581f
C22406 DVDD.n19467 VSS 0.005096f
C22407 DVDD.n19468 VSS 0.005096f
C22408 DVDD.n19469 VSS 0.006035f
C22409 DVDD.n19471 VSS 0.006035f
C22410 DVDD.n19472 VSS 0.006035f
C22411 DVDD.n19473 VSS 0.005096f
C22412 DVDD.n19474 VSS 0.005096f
C22413 DVDD.n19475 VSS 0.005096f
C22414 DVDD.n19476 VSS 0.006035f
C22415 DVDD.n19478 VSS 0.006035f
C22416 DVDD.n19479 VSS 0.006035f
C22417 DVDD.n19480 VSS 0.005096f
C22418 DVDD.n19481 VSS 0.005096f
C22419 DVDD.n19482 VSS 0.005096f
C22420 DVDD.n19483 VSS 0.006035f
C22421 DVDD.n19485 VSS 0.006035f
C22422 DVDD.n19486 VSS 0.006035f
C22423 DVDD.n19487 VSS 0.005096f
C22424 DVDD.n19488 VSS 0.005096f
C22425 DVDD.n19489 VSS 0.005096f
C22426 DVDD.n19490 VSS 0.006035f
C22427 DVDD.n19492 VSS 0.006035f
C22428 DVDD.n19493 VSS 0.006035f
C22429 DVDD.n19494 VSS 0.005096f
C22430 DVDD.n19495 VSS 0.005096f
C22431 DVDD.n19496 VSS 0.005096f
C22432 DVDD.n19497 VSS 0.006035f
C22433 DVDD.n19499 VSS 0.006035f
C22434 DVDD.n19500 VSS 0.006035f
C22435 DVDD.n19501 VSS 0.005096f
C22436 DVDD.n19502 VSS 0.005071f
C22437 DVDD.n19503 VSS 0.081946f
C22438 DVDD.n19504 VSS 0.002548f
C22439 DVDD.n19505 VSS 0.002572f
C22440 DVDD.n19506 VSS 0.006035f
C22441 DVDD.n19508 VSS 0.006035f
C22442 DVDD.n19509 VSS 0.006035f
C22443 DVDD.n19510 VSS 0.005096f
C22444 DVDD.n19511 VSS 0.005096f
C22445 DVDD.n19512 VSS 0.005096f
C22446 DVDD.n19513 VSS 0.006035f
C22447 DVDD.n19515 VSS 0.006035f
C22448 DVDD.n19516 VSS 0.006035f
C22449 DVDD.n19517 VSS 0.005096f
C22450 DVDD.n19518 VSS 0.005096f
C22451 DVDD.n19519 VSS 0.005096f
C22452 DVDD.n19520 VSS 0.006035f
C22453 DVDD.n19522 VSS 0.006035f
C22454 DVDD.n19523 VSS 0.006035f
C22455 DVDD.n19524 VSS 0.005096f
C22456 DVDD.n19525 VSS 0.005096f
C22457 DVDD.n19526 VSS 0.005096f
C22458 DVDD.n19527 VSS 0.006035f
C22459 DVDD.n19529 VSS 0.006035f
C22460 DVDD.n19530 VSS 0.006035f
C22461 DVDD.n19531 VSS 0.005096f
C22462 DVDD.n19532 VSS 0.005096f
C22463 DVDD.n19533 VSS 0.005096f
C22464 DVDD.n19534 VSS 0.006035f
C22465 DVDD.n19536 VSS 0.006035f
C22466 DVDD.n19537 VSS 0.006035f
C22467 DVDD.n19538 VSS 0.005096f
C22468 DVDD.n19539 VSS 0.005096f
C22469 DVDD.n19540 VSS 0.005096f
C22470 DVDD.n19541 VSS 0.006035f
C22471 DVDD.n19543 VSS 0.006035f
C22472 DVDD.n19544 VSS 0.006035f
C22473 DVDD.n19545 VSS 0.005096f
C22474 DVDD.n19546 VSS 0.005096f
C22475 DVDD.n19547 VSS 0.005096f
C22476 DVDD.n19548 VSS 0.006035f
C22477 DVDD.n19550 VSS 0.006035f
C22478 DVDD.n19551 VSS 0.006035f
C22479 DVDD.n19552 VSS 0.002572f
C22480 DVDD.n19553 VSS 0.081946f
C22481 DVDD.n19554 VSS 0.002548f
C22482 DVDD.n19555 VSS 0.005071f
C22483 DVDD.n19556 VSS 0.005096f
C22484 DVDD.n19557 VSS 0.006035f
C22485 DVDD.n19559 VSS 0.006035f
C22486 DVDD.n19560 VSS 0.006035f
C22487 DVDD.n19561 VSS 0.005096f
C22488 DVDD.n19562 VSS 0.005096f
C22489 DVDD.n19563 VSS 0.005096f
C22490 DVDD.n19564 VSS 0.006035f
C22491 DVDD.n19566 VSS 0.006035f
C22492 DVDD.n19567 VSS 0.006035f
C22493 DVDD.n19568 VSS 0.005096f
C22494 DVDD.n19569 VSS 0.005096f
C22495 DVDD.n19570 VSS 0.005096f
C22496 DVDD.n19571 VSS 0.006035f
C22497 DVDD.n19573 VSS 0.006035f
C22498 DVDD.n19574 VSS 0.006035f
C22499 DVDD.n19575 VSS 0.005096f
C22500 DVDD.n19576 VSS 0.005096f
C22501 DVDD.n19577 VSS 0.005096f
C22502 DVDD.n19578 VSS 0.006035f
C22503 DVDD.n19580 VSS 0.006035f
C22504 DVDD.n19581 VSS 0.006035f
C22505 DVDD.n19582 VSS 0.005096f
C22506 DVDD.n19583 VSS 0.005096f
C22507 DVDD.n19584 VSS 0.005096f
C22508 DVDD.n19585 VSS 0.006035f
C22509 DVDD.n19587 VSS 0.006035f
C22510 DVDD.n19588 VSS 0.006035f
C22511 DVDD.n19589 VSS 0.005096f
C22512 DVDD.n19590 VSS 0.005096f
C22513 DVDD.n19591 VSS 0.004581f
C22514 DVDD.n19592 VSS 0.006035f
C22515 DVDD.n19594 VSS 0.006035f
C22516 DVDD.n19595 VSS 0.006035f
C22517 DVDD.n19596 VSS 0.005096f
C22518 DVDD.n19597 VSS 0.005096f
C22519 DVDD.n19598 VSS 0.005096f
C22520 DVDD.n19599 VSS 0.006035f
C22521 DVDD.n19601 VSS 0.006035f
C22522 DVDD.n19602 VSS 0.006035f
C22523 DVDD.n19603 VSS 0.005096f
C22524 DVDD.n19604 VSS 0.005096f
C22525 DVDD.n19605 VSS 0.005096f
C22526 DVDD.n19606 VSS 0.006035f
C22527 DVDD.n19608 VSS 0.006035f
C22528 DVDD.n19609 VSS 0.006035f
C22529 DVDD.n19610 VSS 0.005096f
C22530 DVDD.n19611 VSS 0.005096f
C22531 DVDD.n19612 VSS 0.005096f
C22532 DVDD.n19613 VSS 0.006035f
C22533 DVDD.n19615 VSS 0.006035f
C22534 DVDD.n19616 VSS 0.006035f
C22535 DVDD.n19617 VSS 0.005096f
C22536 DVDD.n19618 VSS 0.005096f
C22537 DVDD.n19619 VSS 0.005096f
C22538 DVDD.n19620 VSS 0.006035f
C22539 DVDD.n19622 VSS 0.006035f
C22540 DVDD.n19623 VSS 0.006035f
C22541 DVDD.n19624 VSS 0.005096f
C22542 DVDD.n19625 VSS 0.005096f
C22543 DVDD.n19626 VSS 0.005096f
C22544 DVDD.n19627 VSS 0.006035f
C22545 DVDD.n19629 VSS 0.006035f
C22546 DVDD.n19630 VSS 0.006035f
C22547 DVDD.n19631 VSS 0.004312f
C22548 DVDD.n19632 VSS 0.002548f
C22549 DVDD.n19633 VSS 0.075949f
C22550 DVDD.n19635 VSS 0.112087f
C22551 DVDD.n19638 VSS 0.055963f
C22552 DVDD.n19639 VSS 0.128173f
C22553 DVDD.n19640 VSS 0.128173f
C22554 DVDD.n19641 VSS 0.128173f
C22555 DVDD.n19642 VSS 0.055963f
C22556 DVDD.n19643 VSS 0.128173f
C22557 DVDD.n19644 VSS 0.055963f
C22558 DVDD.n19645 VSS 0.128173f
C22559 DVDD.n19646 VSS 0.055963f
C22560 DVDD.n19647 VSS 0.128173f
C22561 DVDD.n19648 VSS 0.055963f
C22562 DVDD.n19649 VSS 0.159421f
C22563 DVDD.n19650 VSS 0.353461f
C22564 DVDD.n19651 VSS 0.587306f
C22565 DVDD.n19652 VSS 0.128173f
C22566 DVDD.n19653 VSS 0.055963f
C22567 DVDD.n19654 VSS 0.128173f
C22568 DVDD.n19655 VSS 0.055963f
C22569 DVDD.n19656 VSS 0.128173f
C22570 DVDD.n19657 VSS 0.055963f
C22571 DVDD.n19658 VSS 0.128173f
C22572 DVDD.n19659 VSS 0.128173f
C22573 DVDD.n19660 VSS 0.128173f
C22574 DVDD.n19661 VSS 0.128173f
C22575 DVDD.n19662 VSS 0.128173f
C22576 DVDD.n19663 VSS 0.055963f
C22577 DVDD.n19664 VSS 0.128173f
C22578 DVDD.n19665 VSS 0.055963f
C22579 DVDD.n19666 VSS 0.128173f
C22580 DVDD.n19667 VSS 0.128173f
C22581 DVDD.n19668 VSS 0.128173f
C22582 DVDD.n19669 VSS 0.128173f
C22583 DVDD.n19670 VSS 0.128173f
C22584 DVDD.n19671 VSS 0.128173f
C22585 DVDD.n19672 VSS 0.128173f
C22586 DVDD.n19673 VSS 0.128173f
C22587 DVDD.n19674 VSS 0.055963f
C22588 DVDD.n19675 VSS 0.128173f
C22589 DVDD.n19676 VSS 0.055963f
C22590 DVDD.n19677 VSS 0.128173f
C22591 DVDD.n19678 VSS 0.128173f
C22592 DVDD.n19679 VSS 0.128173f
C22593 DVDD.n19680 VSS 0.055963f
C22594 DVDD.n19681 VSS 0.128173f
C22595 DVDD.n19682 VSS 0.128173f
C22596 DVDD.n19683 VSS 0.128173f
C22597 DVDD.n19684 VSS 0.128173f
C22598 DVDD.n19685 VSS 0.128173f
C22599 DVDD.n19686 VSS 0.128173f
C22600 DVDD.n19687 VSS 0.128173f
C22601 DVDD.n19688 VSS 0.128173f
C22602 DVDD.n19689 VSS 0.128173f
C22603 DVDD.n19690 VSS 0.128173f
C22604 DVDD.n19691 VSS 0.128173f
C22605 DVDD.n19692 VSS 0.128173f
C22606 DVDD.n19693 VSS 0.128173f
C22607 DVDD.n19694 VSS 0.128173f
C22608 DVDD.n19695 VSS 0.128173f
C22609 DVDD.n19696 VSS 0.055963f
C22610 DVDD.n19699 VSS 0.064086f
C22611 DVDD.n19700 VSS 0.151899f
C22612 DVDD.n19701 VSS 0.064086f
C22613 DVDD.n19702 VSS 1.27644f
C22614 DVDD.n19703 VSS 1.27644f
C22615 DVDD.n19704 VSS 0.151899f
C22616 DVDD.n19705 VSS 0.151899f
C22617 DVDD.n19706 VSS 0.151899f
C22618 DVDD.n19707 VSS 0.151899f
C22619 DVDD.n19708 VSS 0.151899f
C22620 DVDD.n19709 VSS 0.079947f
C22621 DVDD.n19710 VSS 0.115237f
C22622 DVDD.n19711 VSS 0.115237f
C22623 DVDD.n19712 VSS 0.079947f
C22624 DVDD.n19713 VSS 0.163891f
C22625 DVDD.n19714 VSS 0.079947f
C22626 DVDD.n19715 VSS 0.163891f
C22627 DVDD.n19716 VSS 0.079947f
C22628 DVDD.n19717 VSS 0.163891f
C22629 DVDD.n19718 VSS 0.079947f
C22630 DVDD.n19719 VSS 0.118292f
C22631 DVDD.n19720 VSS 0.079947f
C22632 DVDD.n19721 VSS 0.081946f
C22633 DVDD.n19722 VSS 0.081946f
C22634 DVDD.n19723 VSS 0.079947f
C22635 DVDD.n19724 VSS 0.057768f
C22636 DVDD.n19725 VSS 0.064086f
C22637 DVDD.n19726 VSS 0.064086f
C22638 DVDD.n19727 VSS 0.064086f
C22639 DVDD.n19728 VSS 0.056865f
C22640 DVDD.n19729 VSS 0.064086f
C22641 DVDD.n19730 VSS 0.064086f
C22642 DVDD.n19731 VSS 0.064086f
C22643 DVDD.n19732 VSS 0.081946f
C22644 DVDD.n19733 VSS 0.064086f
C22645 DVDD.n19734 VSS 0.064086f
C22646 DVDD.n19735 VSS 0.063184f
C22647 DVDD.n19736 VSS 0.064086f
C22648 DVDD.n19737 VSS 0.064086f
C22649 DVDD.n19738 VSS 0.064086f
C22650 DVDD.n19739 VSS 0.062281f
C22651 DVDD.n19740 VSS 0.055963f
C22652 DVDD.n19741 VSS 0.081946f
C22653 DVDD.n19742 VSS 0.081946f
C22654 DVDD.n19743 VSS 0.081946f
C22655 DVDD.n19744 VSS 0.081946f
C22656 DVDD.n19745 VSS 0.074015f
C22657 DVDD.n19748 VSS 0.081946f
C22658 DVDD.n19749 VSS 0.081946f
C22659 DVDD.n19750 VSS 0.081946f
C22660 DVDD.n19751 VSS 0.081946f
C22661 DVDD.n19752 VSS 0.079947f
C22662 DVDD.n19753 VSS 0.079947f
C22663 DVDD.n19754 VSS 0.079947f
C22664 DVDD.n19755 VSS 0.079947f
C22665 DVDD.n19756 VSS 0.079947f
C22666 DVDD.n19757 VSS 0.079947f
C22667 DVDD.n19758 VSS 0.079947f
C22668 DVDD.n19759 VSS 0.079947f
C22669 DVDD.n19760 VSS 0.163891f
C22670 DVDD.n19761 VSS 0.079947f
C22671 DVDD.n19762 VSS 0.163891f
C22672 DVDD.n19763 VSS 0.079947f
C22673 DVDD.n19764 VSS 0.812186f
C22674 DVDD.n19765 VSS 0.079947f
C22675 DVDD.n19766 VSS 0.163891f
C22676 DVDD.n19768 VSS 0.02942f
C22677 DVDD.n19769 VSS 0.02942f
C22678 DVDD.n19770 VSS 0.02942f
C22679 DVDD.n19771 VSS 0.02942f
C22680 DVDD.n19772 VSS 0.02942f
C22681 DVDD.n19773 VSS 0.075212f
C22682 DVDD.n19774 VSS 0.02942f
C22683 DVDD.n19775 VSS 0.02942f
C22684 DVDD.n19776 VSS 0.02942f
C22685 DVDD.n19777 VSS 0.02942f
C22686 DVDD.n19778 VSS 0.02942f
C22687 DVDD.n19779 VSS 0.02942f
C22688 DVDD.n19781 VSS 0.02942f
C22689 DVDD.n19788 VSS 0.163891f
C22690 DVDD.n19789 VSS -1.02989f
C22691 DVDD.n19798 VSS 0.015989f
C22692 DVDD.n19799 VSS 0.015989f
C22693 DVDD.n19800 VSS 0.015989f
C22694 DVDD.n19801 VSS 0.015989f
C22695 DVDD.n19802 VSS 0.015989f
C22696 DVDD.n19803 VSS 0.015989f
C22697 DVDD.n19804 VSS 0.015989f
C22698 DVDD.n19805 VSS 0.015989f
C22699 DVDD.n19806 VSS 0.015989f
C22700 DVDD.n19807 VSS 0.015989f
C22701 DVDD.n19808 VSS 0.015989f
C22702 DVDD.n19809 VSS 0.007995f
C22703 DVDD.n19817 VSS 0.064891f
C22704 DVDD.n19818 VSS 0.02942f
C22705 DVDD.n19819 VSS 0.02942f
C22706 DVDD.n19820 VSS 0.163891f
C22707 DVDD.n19821 VSS 0.163891f
C22708 DVDD.n19822 VSS 0.079947f
C22709 DVDD.n19823 VSS 0.115237f
C22710 DVDD.n19824 VSS 0.079947f
C22711 DVDD.n19825 VSS 0.163891f
C22712 DVDD.n19826 VSS 0.079947f
C22713 DVDD.n19827 VSS 0.163891f
C22714 DVDD.n19828 VSS 0.079947f
C22715 DVDD.n19829 VSS 0.079947f
C22716 DVDD.n19830 VSS 0.163891f
C22717 DVDD.n19831 VSS 0.079947f
C22718 DVDD.n19832 VSS 0.081946f
C22719 DVDD.n19833 VSS 0.079947f
C22720 DVDD.n19834 VSS 0.064086f
C22721 DVDD.n19835 VSS 0.064086f
C22722 DVDD.n19836 VSS 0.061379f
C22723 DVDD.n19837 VSS 0.064086f
C22724 DVDD.n19838 VSS 0.064086f
C22725 DVDD.n19839 VSS 0.064086f
C22726 DVDD.n19840 VSS 0.060476f
C22727 DVDD.n19841 VSS 0.064086f
C22728 DVDD.n19842 VSS 0.081946f
C22729 DVDD.n19843 VSS 0.059573f
C22730 DVDD.n19844 VSS 0.064086f
C22731 DVDD.n19845 VSS 0.064086f
C22732 DVDD.n19846 VSS 0.064086f
C22733 DVDD.n19847 VSS 0.058671f
C22734 DVDD.n19848 VSS 0.064086f
C22735 DVDD.n19849 VSS 0.064086f
C22736 DVDD.n19850 VSS 0.055963f
C22737 DVDD.n19851 VSS 0.081946f
C22738 DVDD.n19852 VSS 0.081946f
C22739 DVDD.n19853 VSS 0.081946f
C22740 DVDD.n19854 VSS 0.081946f
C22741 DVDD.n19855 VSS 0.128173f
C22742 DVDD.n19856 VSS 0.128173f
C22743 DVDD.n19857 VSS 0.128173f
C22744 DVDD.n19858 VSS 0.128173f
C22745 DVDD.n19859 VSS 0.055963f
C22746 DVDD.n19860 VSS 0.128173f
C22747 DVDD.n19861 VSS 0.128173f
C22748 DVDD.n19862 VSS 0.055963f
C22749 DVDD.n19863 VSS 0.128173f
C22750 DVDD.n19864 VSS 0.128173f
C22751 DVDD.n19865 VSS 0.055963f
C22752 DVDD.n19866 VSS 0.128173f
C22753 DVDD.n19867 VSS 0.128173f
C22754 DVDD.n19868 VSS 0.128173f
C22755 DVDD.n19869 VSS 0.090263f
C22756 DVDD.n19870 VSS 0.128173f
C22757 DVDD.n19871 VSS 0.128173f
C22758 DVDD.n19872 VSS 0.128173f
C22759 DVDD.n19873 VSS 0.064086f
C22760 DVDD.n19874 VSS 0.081946f
C22761 DVDD.n19875 VSS 0.081946f
C22762 DVDD.n19876 VSS 0.081946f
C22763 DVDD.n19877 VSS 0.081946f
C22764 DVDD.n19878 VSS 0.081946f
C22765 DVDD.n19879 VSS 0.081946f
C22766 DVDD.n19880 VSS 0.081946f
C22767 DVDD.n19881 VSS 0.081946f
C22768 DVDD.n19882 VSS 0.081946f
C22769 DVDD.n19883 VSS 0.081946f
C22770 DVDD.n19884 VSS 0.118292f
C22771 DVDD.n19885 VSS 0.057768f
C22772 DVDD.n19886 VSS 0.064086f
C22773 DVDD.n19887 VSS 0.064086f
C22774 DVDD.n19888 VSS 0.064086f
C22775 DVDD.n19889 VSS 0.056865f
C22776 DVDD.n19890 VSS 0.064086f
C22777 DVDD.n19891 VSS 0.064086f
C22778 DVDD.n19892 VSS 0.079947f
C22779 DVDD.n19893 VSS 0.163891f
C22780 DVDD.n19894 VSS 0.079947f
C22781 DVDD.n19895 VSS 0.648295f
C22782 DVDD.n19896 VSS 0.163891f
C22783 DVDD.n19897 VSS 0.163891f
C22784 DVDD.n19898 VSS 0.079947f
C22785 DVDD.n19899 VSS 0.079947f
C22786 DVDD.n19900 VSS 0.079947f
C22787 DVDD.n19901 VSS 0.163891f
C22788 DVDD.n19902 VSS 0.163891f
C22789 DVDD.n19903 VSS 0.163891f
C22790 DVDD.n19904 VSS 0.079947f
C22791 DVDD.n19905 VSS 0.079947f
C22792 DVDD.n19906 VSS 0.079947f
C22793 DVDD.n19907 VSS 0.163891f
C22794 DVDD.n19908 VSS 0.163891f
C22795 DVDD.n19909 VSS 0.079947f
C22796 DVDD.n19910 VSS 0.079947f
C22797 DVDD.n19911 VSS 0.079947f
C22798 DVDD.n19912 VSS 0.163891f
C22799 DVDD.n19913 VSS 0.163891f
C22800 DVDD.n19914 VSS 0.127544f
C22801 DVDD.n19915 VSS 0.079947f
C22802 DVDD.n19916 VSS 0.081946f
C22803 DVDD.n19917 VSS 0.079947f
C22804 DVDD.n19918 VSS 0.081946f
C22805 DVDD.n19919 VSS 0.079947f
C22806 DVDD.n19920 VSS 0.081946f
C22807 DVDD.n19921 VSS 0.079947f
C22808 DVDD.n19922 VSS 0.081946f
C22809 DVDD.n19923 VSS 0.079947f
C22810 DVDD.n19924 VSS 0.081946f
C22811 DVDD.n19925 VSS 0.079947f
C22812 DVDD.n19926 VSS 0.081946f
C22813 DVDD.n19927 VSS 0.079947f
C22814 DVDD.n19928 VSS 0.081946f
C22815 DVDD.n19929 VSS 0.079947f
C22816 DVDD.n19930 VSS 0.081946f
C22817 DVDD.n19931 VSS 0.079947f
C22818 DVDD.n19932 VSS 0.081946f
C22819 DVDD.n19933 VSS 0.079947f
C22820 DVDD.n19934 VSS 0.079947f
C22821 DVDD.n19935 VSS 0.081946f
C22822 DVDD.n19936 VSS 0.064086f
C22823 DVDD.n19938 VSS 0.063184f
C22824 DVDD.n19939 VSS 0.064086f
C22825 DVDD.n19940 VSS 0.064086f
C22826 DVDD.n19941 VSS 0.064086f
C22827 DVDD.n19943 VSS 0.062281f
C22828 DVDD.n19944 VSS 0.055963f
C22829 DVDD.n19945 VSS 0.128173f
C22830 DVDD.n19946 VSS 0.128173f
C22831 DVDD.n19947 VSS 0.055963f
C22832 DVDD.n19948 VSS 0.128173f
C22833 DVDD.n19949 VSS 0.128173f
C22834 DVDD.n19950 VSS 0.055963f
C22835 DVDD.n19951 VSS 0.128173f
C22836 DVDD.n19952 VSS 0.128173f
C22837 DVDD.n19953 VSS 0.128173f
C22838 DVDD.n19954 VSS 0.128173f
C22839 DVDD.n19955 VSS 0.128173f
C22840 DVDD.n19956 VSS 0.128173f
C22841 DVDD.n19957 VSS 0.128173f
C22842 DVDD.n19958 VSS 0.055963f
C22843 DVDD.n19959 VSS 0.081946f
C22844 DVDD.n19960 VSS 0.081946f
C22845 DVDD.n19961 VSS 0.081946f
C22846 DVDD.n19962 VSS 0.081946f
C22847 DVDD.n19963 VSS 0.081946f
C22848 DVDD.n19964 VSS 0.081946f
C22849 DVDD.n19965 VSS 0.081946f
C22850 DVDD.n19966 VSS 0.081946f
C22851 DVDD.n19967 VSS 0.081946f
C22852 DVDD.n19968 VSS 0.081946f
C22853 DVDD.n19969 VSS 0.118292f
C22854 DVDD.n19970 VSS 0.064086f
C22855 DVDD.n19971 VSS 0.061379f
C22856 DVDD.n19972 VSS 0.064086f
C22857 DVDD.n19973 VSS 0.064086f
C22858 DVDD.n19974 VSS 0.064086f
C22859 DVDD.n19975 VSS 0.060476f
C22860 DVDD.n19976 VSS 0.064086f
C22861 DVDD.n19977 VSS 0.064086f
C22862 DVDD.n19978 VSS 0.079947f
C22863 DVDD.n19979 VSS 0.163891f
C22864 DVDD.n19980 VSS 0.079947f
C22865 DVDD.n19981 VSS 0.115237f
C22866 DVDD.n19982 VSS 0.648295f
C22867 DVDD.n19983 VSS 0.163891f
C22868 DVDD.n19984 VSS 0.163891f
C22869 DVDD.n19985 VSS 0.079947f
C22870 DVDD.n19986 VSS 0.079947f
C22871 DVDD.n19987 VSS 0.079947f
C22872 DVDD.n19988 VSS 0.163891f
C22873 DVDD.n19989 VSS 0.163891f
C22874 DVDD.n19990 VSS 0.163891f
C22875 DVDD.n19991 VSS 0.079947f
C22876 DVDD.n19992 VSS 0.079947f
C22877 DVDD.n19993 VSS 0.079947f
C22878 DVDD.n19994 VSS 0.163891f
C22879 DVDD.n19995 VSS 0.163891f
C22880 DVDD.n19996 VSS 0.079947f
C22881 DVDD.n19997 VSS 0.079947f
C22882 DVDD.n19998 VSS 0.079947f
C22883 DVDD.n19999 VSS 0.163891f
C22884 DVDD.n20000 VSS 0.163891f
C22885 DVDD.n20001 VSS 0.127544f
C22886 DVDD.n20002 VSS 0.079947f
C22887 DVDD.n20003 VSS 0.081946f
C22888 DVDD.n20004 VSS 0.079947f
C22889 DVDD.n20005 VSS 0.081946f
C22890 DVDD.n20006 VSS 0.079947f
C22891 DVDD.n20007 VSS 0.081946f
C22892 DVDD.n20008 VSS 0.079947f
C22893 DVDD.n20009 VSS 0.081946f
C22894 DVDD.n20010 VSS 0.079947f
C22895 DVDD.n20011 VSS 0.081946f
C22896 DVDD.n20012 VSS 0.079947f
C22897 DVDD.n20013 VSS 0.081946f
C22898 DVDD.n20014 VSS 0.079947f
C22899 DVDD.n20015 VSS 0.081946f
C22900 DVDD.n20016 VSS 0.079947f
C22901 DVDD.n20017 VSS 0.081946f
C22902 DVDD.n20018 VSS 0.079947f
C22903 DVDD.n20019 VSS 0.081946f
C22904 DVDD.n20020 VSS 0.079947f
C22905 DVDD.n20021 VSS 0.079947f
C22906 DVDD.n20022 VSS 0.081946f
C22907 DVDD.n20023 VSS 0.064086f
C22908 DVDD.n20025 VSS 0.059573f
C22909 DVDD.n20026 VSS 0.064086f
C22910 DVDD.n20027 VSS 0.064086f
C22911 DVDD.n20028 VSS 0.064086f
C22912 DVDD.n20030 VSS 0.058671f
C22913 DVDD.n20031 VSS 0.055963f
C22914 DVDD.n20032 VSS 0.128173f
C22915 DVDD.n20033 VSS 0.128173f
C22916 DVDD.n20034 VSS 0.128173f
C22917 DVDD.n20035 VSS 0.055963f
C22918 DVDD.n20036 VSS 0.128173f
C22919 DVDD.n20037 VSS 0.128173f
C22920 DVDD.n20038 VSS 0.055963f
C22921 DVDD.n20039 VSS 0.128173f
C22922 DVDD.n20040 VSS 0.128173f
C22923 DVDD.n20041 VSS 0.128173f
C22924 DVDD.n20042 VSS 0.128173f
C22925 DVDD.n20043 VSS 0.128173f
C22926 DVDD.n20044 VSS 0.128173f
C22927 DVDD.n20045 VSS 0.055963f
C22928 DVDD.n20046 VSS 0.128173f
C22929 DVDD.n20047 VSS 0.128173f
C22930 DVDD.n20048 VSS 0.055963f
C22931 DVDD.n20049 VSS 0.128173f
C22932 DVDD.n20050 VSS 0.128173f
C22933 DVDD.n20051 VSS 0.055963f
C22934 DVDD.n20052 VSS 0.128173f
C22935 DVDD.n20053 VSS 0.128173f
C22936 DVDD.n20054 VSS 0.128173f
C22937 DVDD.n20055 VSS 0.128173f
C22938 DVDD.n20056 VSS 0.128173f
C22939 DVDD.n20057 VSS 0.128173f
C22940 DVDD.n20058 VSS 0.128173f
C22941 DVDD.n20059 VSS 0.055963f
C22942 DVDD.n20060 VSS 0.075949f
C22943 DVDD.n20061 VSS 0.075949f
C22944 DVDD.n20062 VSS 0.075949f
C22945 DVDD.n20063 VSS 0.075949f
C22946 DVDD.n20064 VSS 0.075949f
C22947 DVDD.n20065 VSS 0.075949f
C22948 DVDD.n20066 VSS 0.075949f
C22949 DVDD.n20067 VSS 0.075949f
C22950 DVDD.n20068 VSS 0.075949f
C22951 DVDD.n20069 VSS 0.075949f
C22952 DVDD.n20070 VSS 0.109637f
C22953 DVDD.n20071 VSS 0.064086f
C22954 DVDD.n20072 VSS 0.064086f
C22955 DVDD.n20073 VSS 0.059122f
C22956 DVDD.n20074 VSS 0.064086f
C22957 DVDD.n20075 VSS 0.064086f
C22958 DVDD.n20076 VSS 0.064086f
C22959 DVDD.n20077 VSS 0.060025f
C22960 DVDD.n20078 VSS 0.079947f
C22961 DVDD.n20079 VSS 0.151899f
C22962 DVDD.n20080 VSS 0.079947f
C22963 DVDD.n20081 VSS 0.600859f
C22964 DVDD.n20082 VSS 0.151899f
C22965 DVDD.n20083 VSS 0.151899f
C22966 DVDD.n20084 VSS 0.079947f
C22967 DVDD.n20085 VSS 0.079947f
C22968 DVDD.n20086 VSS 0.079947f
C22969 DVDD.n20087 VSS 0.151899f
C22970 DVDD.n20088 VSS 0.151899f
C22971 DVDD.n20089 VSS 0.151899f
C22972 DVDD.n20090 VSS 0.079947f
C22973 DVDD.n20091 VSS 0.079947f
C22974 DVDD.n20092 VSS 0.079947f
C22975 DVDD.n20093 VSS 0.151899f
C22976 DVDD.n20094 VSS 0.151899f
C22977 DVDD.n20095 VSS 0.079947f
C22978 DVDD.n20096 VSS 0.079947f
C22979 DVDD.n20097 VSS 0.079947f
C22980 DVDD.n20098 VSS 0.151899f
C22981 DVDD.n20099 VSS 0.151899f
C22982 DVDD.n20100 VSS 0.118212f
C22983 DVDD.n20101 VSS 0.079947f
C22984 DVDD.n20102 VSS 0.075949f
C22985 DVDD.n20103 VSS 0.079947f
C22986 DVDD.n20104 VSS 0.075949f
C22987 DVDD.n20105 VSS 0.079947f
C22988 DVDD.n20106 VSS 0.075949f
C22989 DVDD.n20107 VSS 0.079947f
C22990 DVDD.n20108 VSS 0.075949f
C22991 DVDD.n20109 VSS 0.079947f
C22992 DVDD.n20110 VSS 0.075949f
C22993 DVDD.n20111 VSS 0.079947f
C22994 DVDD.n20112 VSS 0.075949f
C22995 DVDD.n20113 VSS 0.079947f
C22996 DVDD.n20114 VSS 0.075949f
C22997 DVDD.n20115 VSS 0.079947f
C22998 DVDD.n20116 VSS 0.075949f
C22999 DVDD.n20117 VSS 0.079947f
C23000 DVDD.n20118 VSS 0.075949f
C23001 DVDD.n20119 VSS 0.079947f
C23002 DVDD.n20120 VSS 0.079947f
C23003 DVDD.n20121 VSS 0.075949f
C23004 DVDD.n20122 VSS 0.373774f
C23005 DVDD.n20124 VSS 0.060025f
C23006 DVDD.n20125 VSS 0.064086f
C23007 DVDD.n20126 VSS 0.064086f
C23008 DVDD.n20127 VSS 0.064086f
C23009 DVDD.n20129 VSS 0.060927f
C23010 DVDD.n20130 VSS 0.055963f
C23011 DVDD.n20131 VSS 0.128173f
C23012 DVDD.n20132 VSS 0.128173f
C23013 DVDD.n20133 VSS 0.055963f
C23014 DVDD.n20134 VSS 0.128173f
C23015 DVDD.n20135 VSS 0.128173f
C23016 DVDD.n20136 VSS 0.055963f
C23017 DVDD.n20137 VSS 0.128173f
C23018 DVDD.n20138 VSS 0.055963f
C23019 DVDD.n20139 VSS 0.159414f
C23020 DVDD.n20140 VSS 0.353402f
C23021 DVDD.n20141 VSS 0.587849f
C23022 DVDD.n20142 VSS 0.128173f
C23023 DVDD.n20143 VSS 0.055963f
C23024 DVDD.n20144 VSS 0.128173f
C23025 DVDD.n20145 VSS 0.055963f
C23026 DVDD.n20146 VSS 0.128173f
C23027 DVDD.n20147 VSS 0.055963f
C23028 DVDD.n20148 VSS 0.128173f
C23029 DVDD.n20149 VSS 0.128173f
C23030 DVDD.n20150 VSS 0.128173f
C23031 DVDD.n20151 VSS 0.128173f
C23032 DVDD.n20152 VSS 0.055963f
C23033 DVDD.n20153 VSS 0.128173f
C23034 DVDD.n20154 VSS 0.055963f
C23035 DVDD.n20155 VSS 0.128173f
C23036 DVDD.n20156 VSS 0.055963f
C23037 DVDD.n20157 VSS 0.128173f
C23038 DVDD.n20158 VSS 0.128173f
C23039 DVDD.n20159 VSS 0.128173f
C23040 DVDD.n20160 VSS 0.128173f
C23041 DVDD.n20161 VSS 0.128173f
C23042 DVDD.n20162 VSS 0.055963f
C23043 DVDD.n20163 VSS 0.064086f
C23044 DVDD.n20164 VSS 0.075949f
C23045 DVDD.n20165 VSS 0.064086f
C23046 DVDD.n20166 VSS 0.101545f
C23047 DVDD.n20167 VSS 0.128173f
C23048 DVDD.n20168 VSS 0.128173f
C23049 DVDD.n20169 VSS 0.128173f
C23050 DVDD.n20170 VSS 0.128173f
C23051 DVDD.n20171 VSS 0.128173f
C23052 DVDD.n20172 VSS 0.128173f
C23053 DVDD.n20173 VSS 0.128173f
C23054 DVDD.n20174 VSS 0.128173f
C23055 DVDD.n20175 VSS 0.111926f
C23056 DVDD.n20176 VSS 0.128173f
C23057 DVDD.n20177 VSS 0.055963f
C23058 DVDD.n20178 VSS 0.128173f
C23059 DVDD.n20179 VSS 0.128173f
C23060 DVDD.n20180 VSS 0.128173f
C23061 DVDD.n20181 VSS 0.128173f
C23062 DVDD.n20182 VSS 0.055963f
C23063 DVDD.n20183 VSS 0.128173f
C23064 DVDD.n20184 VSS 0.055963f
C23065 DVDD.n20185 VSS 0.128173f
C23066 DVDD.n20186 VSS 0.055963f
C23067 DVDD.n20187 VSS 0.128173f
C23068 DVDD.n20188 VSS 0.128173f
C23069 DVDD.n20189 VSS 0.128173f
C23070 DVDD.n20190 VSS 0.128173f
C23071 DVDD.n20191 VSS 0.055963f
C23072 DVDD.n20192 VSS 0.128173f
C23073 DVDD.n20193 VSS 0.055963f
C23074 DVDD.n20194 VSS 0.128173f
C23075 DVDD.n20195 VSS 0.055963f
C23076 DVDD.n20196 VSS 0.128173f
C23077 DVDD.n20197 VSS 0.128173f
C23078 DVDD.n20198 VSS 0.128173f
C23079 DVDD.n20199 VSS 0.128173f
C23080 DVDD.n20200 VSS 0.055963f
C23081 DVDD.n20201 VSS 0.128173f
C23082 DVDD.n20202 VSS 0.055963f
C23083 DVDD.n20203 VSS 0.128173f
C23084 DVDD.n20204 VSS 0.128173f
C23085 DVDD.n20205 VSS 0.128173f
C23086 DVDD.n20206 VSS 0.128173f
C23087 DVDD.n20207 VSS 0.128173f
C23088 DVDD.n20208 VSS 0.128173f
C23089 DVDD.n20209 VSS 0.128173f
C23090 DVDD.n20210 VSS 0.128173f
C23091 DVDD.n20211 VSS 0.128173f
C23092 DVDD.n20212 VSS 0.092068f
C23093 DVDD.n20213 VSS 0.128173f
C23094 DVDD.n20214 VSS 0.055963f
C23095 DVDD.n20215 VSS 0.128173f
C23096 DVDD.n20216 VSS 0.055963f
C23097 DVDD.n20217 VSS 0.128173f
C23098 DVDD.n20218 VSS 0.128173f
C23099 DVDD.n20219 VSS 0.128173f
C23100 DVDD.n20220 VSS 0.128173f
C23101 DVDD.n20221 VSS 0.055963f
C23102 DVDD.n20222 VSS 0.128173f
C23103 DVDD.n20223 VSS 0.055963f
C23104 DVDD.n20224 VSS 0.128173f
C23105 DVDD.n20225 VSS 0.055963f
C23106 DVDD.n20226 VSS 0.128173f
C23107 DVDD.n20227 VSS 0.128173f
C23108 DVDD.n20228 VSS 0.128173f
C23109 DVDD.n20229 VSS 0.128173f
C23110 DVDD.n20230 VSS 0.055963f
C23111 DVDD.n20231 VSS 0.128173f
C23112 DVDD.n20232 VSS 0.055963f
C23113 DVDD.n20233 VSS 0.128173f
C23114 DVDD.n20234 VSS 0.055963f
C23115 DVDD.n20235 VSS 0.128173f
C23116 DVDD.n20236 VSS 0.128173f
C23117 DVDD.n20237 VSS 0.128173f
C23118 DVDD.n20238 VSS 0.128173f
C23119 DVDD.n20239 VSS 0.128173f
C23120 DVDD.n20240 VSS 0.128173f
C23121 DVDD.n20241 VSS 0.055963f
C23122 DVDD.n20242 VSS 0.064086f
C23123 DVDD.n20243 VSS 0.081946f
C23124 DVDD.n20244 VSS 0.064086f
C23125 DVDD.n20245 VSS 0.093873f
C23126 DVDD.n20246 VSS 0.128173f
C23127 DVDD.n20247 VSS 0.128173f
C23128 DVDD.n20248 VSS 0.128173f
C23129 DVDD.n20249 VSS 0.128173f
C23130 DVDD.n20250 VSS 0.128173f
C23131 DVDD.n20251 VSS 0.128173f
C23132 DVDD.n20252 VSS 0.128173f
C23133 DVDD.n20253 VSS 0.128173f
C23134 DVDD.n20254 VSS 0.128173f
C23135 DVDD.n20255 VSS 0.095678f
C23136 DVDD.n20256 VSS 0.128173f
C23137 DVDD.n20257 VSS 0.055963f
C23138 DVDD.n20258 VSS 0.128173f
C23139 DVDD.n20259 VSS 0.128173f
C23140 DVDD.n20260 VSS 0.128173f
C23141 DVDD.n20261 VSS 0.128173f
C23142 DVDD.n20262 VSS 0.055963f
C23143 DVDD.n20263 VSS 0.128173f
C23144 DVDD.n20264 VSS 0.055963f
C23145 DVDD.n20265 VSS 0.128173f
C23146 DVDD.n20266 VSS 0.055963f
C23147 DVDD.n20267 VSS 0.128173f
C23148 DVDD.n20268 VSS 0.128173f
C23149 DVDD.n20269 VSS 0.128173f
C23150 DVDD.n20270 VSS 0.128173f
C23151 DVDD.n20271 VSS 0.055963f
C23152 DVDD.n20272 VSS 0.128173f
C23153 DVDD.n20273 VSS 0.055963f
C23154 DVDD.n20274 VSS 0.128173f
C23155 DVDD.n20275 VSS 0.055963f
C23156 DVDD.n20276 VSS 0.128173f
C23157 DVDD.n20277 VSS 0.128173f
C23158 DVDD.n20278 VSS 0.128173f
C23159 DVDD.n20279 VSS 0.128173f
C23160 DVDD.n20280 VSS 0.128173f
C23161 DVDD.n20281 VSS 0.055963f
C23162 DVDD.n20282 VSS 0.055963f
C23163 DVDD.n20283 VSS 0.064086f
C23164 DVDD.n20284 VSS 0.081946f
C23165 DVDD.n20285 VSS 0.064086f
C23166 DVDD.n20286 VSS 0.055963f
C23167 DVDD.n20287 VSS 0.128173f
C23168 DVDD.n20288 VSS 0.128173f
C23169 DVDD.n20289 VSS 0.128173f
C23170 DVDD.n20290 VSS 0.128173f
C23171 DVDD.n20291 VSS 0.128173f
C23172 DVDD.n20292 VSS 0.128173f
C23173 DVDD.n20293 VSS 0.128173f
C23174 DVDD.n20294 VSS 0.075821f
C23175 DVDD.n20295 VSS 0.128173f
C23176 DVDD.n20296 VSS 0.128173f
C23177 DVDD.n20297 VSS 0.128173f
C23178 DVDD.n20298 VSS 0.128173f
C23179 DVDD.n20299 VSS 0.055963f
C23180 DVDD.n20300 VSS 0.128173f
C23181 DVDD.n20301 VSS 0.055963f
C23182 DVDD.n20302 VSS 0.128173f
C23183 DVDD.n20303 VSS 0.055963f
C23184 DVDD.n20304 VSS 0.128173f
C23185 DVDD.n20305 VSS 0.128173f
C23186 DVDD.n20306 VSS 0.128173f
C23187 DVDD.n20307 VSS 0.128173f
C23188 DVDD.n20308 VSS 0.055963f
C23189 DVDD.n20309 VSS 0.128173f
C23190 DVDD.n20310 VSS 0.055963f
C23191 DVDD.n20311 VSS 0.128173f
C23192 DVDD.n20312 VSS 0.055963f
C23193 DVDD.n20313 VSS 0.128173f
C23194 DVDD.n20314 VSS 0.128173f
C23195 DVDD.n20315 VSS 0.128173f
C23196 DVDD.n20316 VSS 0.128173f
C23197 DVDD.n20317 VSS 0.055963f
C23198 DVDD.n20318 VSS 0.128173f
C23199 DVDD.n20319 VSS 0.055963f
C23200 DVDD.n20320 VSS 0.128173f
C23201 DVDD.n20321 VSS 0.055963f
C23202 DVDD.n20322 VSS 0.128173f
C23203 DVDD.n20323 VSS 0.128173f
C23204 DVDD.n20324 VSS 0.128173f
C23205 DVDD.n20325 VSS 0.128173f
C23206 DVDD.n20326 VSS 0.128173f
C23207 DVDD.n20327 VSS 0.055963f
C23208 DVDD.n20328 VSS 0.128173f
C23209 DVDD.n20329 VSS 0.128173f
C23210 DVDD.n20330 VSS 0.055963f
C23211 DVDD.n20331 VSS 0.128173f
C23212 DVDD.n20332 VSS 0.128173f
C23213 DVDD.n20333 VSS 0.055963f
C23214 DVDD.n20334 VSS 0.115536f
C23215 DVDD.n20335 VSS 0.159414f
C23216 DVDD.n20336 VSS 0.589426f
C23217 DVDD.n20337 VSS 0.055963f
C23218 DVDD.n20338 VSS 0.128173f
C23219 DVDD.n20339 VSS 0.026627f
C23220 DVDD.n20340 VSS 0.076723f
C23221 DVDD.n20341 VSS 0.065892f
C23222 DVDD.n20342 VSS 0.128173f
C23223 DVDD.n20343 VSS 0.128173f
C23224 DVDD.n20344 VSS 0.055963f
C23225 DVDD.n20345 VSS 0.128173f
C23226 DVDD.n20346 VSS 0.055963f
C23227 DVDD.n20347 VSS 0.128173f
C23228 DVDD.n20348 VSS 0.055963f
C23229 DVDD.n20349 VSS 0.128173f
C23230 DVDD.n20350 VSS 0.128173f
C23231 DVDD.n20351 VSS 0.128173f
C23232 DVDD.n20352 VSS 0.128173f
C23233 DVDD.n20353 VSS 0.055963f
C23234 DVDD.n20354 VSS 0.128173f
C23235 DVDD.n20355 VSS 0.055963f
C23236 DVDD.n20356 VSS 0.128173f
C23237 DVDD.n20357 VSS 0.055963f
C23238 DVDD.n20358 VSS 0.128173f
C23239 DVDD.n20359 VSS 0.128173f
C23240 DVDD.n20360 VSS 0.128173f
C23241 DVDD.n20361 VSS 0.128173f
C23242 DVDD.n20362 VSS 0.128173f
C23243 DVDD.n20363 VSS 0.103351f
C23244 DVDD.n20364 VSS 0.128173f
C23245 DVDD.n20365 VSS 0.128173f
C23246 DVDD.n20366 VSS 0.128173f
C23247 DVDD.n20367 VSS 0.128173f
C23248 DVDD.n20368 VSS 0.128173f
C23249 DVDD.n20369 VSS 0.128173f
C23250 DVDD.n20370 VSS 0.128173f
C23251 DVDD.n20371 VSS 0.11012f
C23252 DVDD.n20374 VSS 0.081946f
C23253 DVDD.n20375 VSS 0.081946f
C23254 DVDD.n20376 VSS 0.081946f
C23255 DVDD.n20377 VSS 0.081946f
C23256 DVDD.n20378 VSS 0.079947f
C23257 DVDD.n20379 VSS 0.079947f
C23258 DVDD.n20380 VSS 0.079947f
C23259 DVDD.n20381 VSS 0.079947f
C23260 DVDD.n20382 VSS 0.079947f
C23261 DVDD.n20383 VSS 0.079947f
C23262 DVDD.n20384 VSS 0.079947f
C23263 DVDD.n20385 VSS 0.163891f
C23264 DVDD.n20386 VSS 0.079947f
C23265 DVDD.n20387 VSS 0.079947f
C23266 DVDD.n20388 VSS 0.163891f
C23267 DVDD.n20389 VSS 0.079947f
C23268 DVDD.n20390 VSS 0.079947f
C23269 DVDD.n20391 VSS 0.079947f
C23270 DVDD.n20392 VSS 0.163891f
C23271 DVDD.n20393 VSS 0.079947f
C23272 DVDD.n20394 VSS 0.079947f
C23273 DVDD.n20395 VSS 0.079947f
C23274 DVDD.n20396 VSS 0.163891f
C23275 DVDD.n20397 VSS 0.127544f
C23276 DVDD.n20398 VSS 0.079947f
C23277 DVDD.n20399 VSS 0.079947f
C23278 DVDD.n20400 VSS 0.081946f
C23279 DVDD.n20401 VSS 0.079947f
C23280 DVDD.n20402 VSS 0.081946f
C23281 DVDD.n20403 VSS 0.079947f
C23282 DVDD.n20404 VSS 0.079947f
C23283 DVDD.n20405 VSS 0.081946f
C23284 DVDD.n20406 VSS 0.079947f
C23285 DVDD.n20407 VSS 0.081946f
C23286 DVDD.n20408 VSS 0.079947f
C23287 DVDD.n20409 VSS 0.079947f
C23288 DVDD.n20410 VSS 0.081946f
C23289 DVDD.n20411 VSS 0.079947f
C23290 DVDD.n20412 VSS 0.081946f
C23291 DVDD.n20413 VSS 0.079947f
C23292 DVDD.n20414 VSS 0.079947f
C23293 DVDD.n20415 VSS 0.081946f
C23294 DVDD.n20416 VSS 0.079947f
C23295 DVDD.n20417 VSS 0.079947f
C23296 DVDD.n20418 VSS 0.081946f
C23297 DVDD.n20419 VSS 0.081946f
C23298 DVDD.n20420 VSS 0.064086f
C23299 DVDD.n20421 VSS 0.081946f
C23300 DVDD.n20422 VSS 0.081946f
C23301 DVDD.n20423 VSS 0.079947f
C23302 DVDD.n20424 VSS 0.079947f
C23303 DVDD.n20425 VSS 0.118292f
C23304 DVDD.n20426 VSS 0.079947f
C23305 DVDD.n20427 VSS 0.079947f
C23306 DVDD.n20428 VSS 0.079947f
C23307 DVDD.n20429 VSS 0.163891f
C23308 DVDD.n20430 VSS 0.079947f
C23309 DVDD.n20431 VSS 0.079947f
C23310 DVDD.n20432 VSS 0.079947f
C23311 DVDD.n20433 VSS 0.163891f
C23312 DVDD.n20434 VSS 0.079947f
C23313 DVDD.n20435 VSS 0.079947f
C23314 DVDD.n20436 VSS 0.079947f
C23315 DVDD.n20437 VSS 0.163891f
C23316 DVDD.n20438 VSS 0.648295f
C23317 DVDD.n20439 VSS 0.115237f
C23318 DVDD.t161 VSS 3.21054f
C23319 DVDD.n20440 VSS 0.115237f
C23320 DVDD.n20441 VSS 0.812186f
C23321 DVDD.n20442 VSS 0.02942f
C23322 DVDD.n20444 VSS 0.02942f
C23323 DVDD.n20445 VSS 0.02942f
C23324 DVDD.n20446 VSS 0.02942f
C23325 DVDD.n20447 VSS 0.02942f
C23326 DVDD.n20448 VSS 0.02942f
C23327 DVDD.n20450 VSS 0.02942f
C23328 DVDD.n20452 VSS 0.02942f
C23329 DVDD.n20454 VSS 0.02942f
C23330 DVDD.n20456 VSS 0.02942f
C23331 DVDD.n20458 VSS 0.02942f
C23332 DVDD.n20460 VSS 0.02942f
C23333 DVDD.n20462 VSS 0.812186f
C23334 DVDD.n20463 VSS 0.075212f
C23335 DVDD.n20464 VSS 0.553132f
C23336 DVDD.n20465 VSS 0.553132f
C23337 DVDD.n20466 VSS 0.007995f
C23338 DVDD.n20467 VSS 0.015989f
C23339 DVDD.n20468 VSS 0.015989f
C23340 DVDD.n20469 VSS 0.015989f
C23341 DVDD.n20470 VSS 0.015989f
C23342 DVDD.n20471 VSS 0.015989f
C23343 DVDD.n20472 VSS 0.015989f
C23344 DVDD.n20473 VSS 0.015989f
C23345 DVDD.n20474 VSS 0.015989f
C23346 DVDD.n20475 VSS 0.015989f
C23347 DVDD.n20476 VSS 0.015989f
C23348 DVDD.n20477 VSS 0.015989f
C23349 DVDD.n20478 VSS 0.007995f
C23350 DVDD.n20479 VSS 0.015989f
C23351 DVDD.n20481 VSS 0.015989f
C23352 DVDD.n20482 VSS 0.035267f
C23353 DVDD.t162 VSS 1.03157f
C23354 DVDD.n20483 VSS 0.035267f
C23355 DVDD.n20484 VSS 0.007995f
C23356 DVDD.n20485 VSS 0.015989f
C23357 DVDD.n20486 VSS 0.007995f
C23358 DVDD.n20487 VSS 0.163891f
C23359 DVDD.n20488 VSS 0.075212f
C23360 DVDD.n20496 VSS 0.02942f
C23361 DVDD.n20498 VSS 0.02942f
C23362 DVDD.n20499 VSS 0.02942f
C23363 DVDD.n20500 VSS 0.02942f
C23364 DVDD.n20501 VSS 0.02942f
C23365 DVDD.n20502 VSS 0.02942f
C23366 DVDD.n20503 VSS 0.02942f
C23367 DVDD.n20505 VSS 0.02942f
C23368 DVDD.n20507 VSS 0.02942f
C23369 DVDD.n20509 VSS 0.02942f
C23370 DVDD.n20511 VSS 0.02942f
C23371 DVDD.n20513 VSS 0.02942f
C23372 DVDD.n20515 VSS 0.02942f
C23373 DVDD.n20516 VSS 0.812186f
C23374 DVDD.n20517 VSS 0.02942f
C23375 DVDD.n20519 VSS 0.553132f
C23376 DVDD.n20521 VSS 0.015989f
C23377 DVDD.n20522 VSS 0.015989f
C23378 DVDD.n20523 VSS 0.015989f
C23379 DVDD.n20524 VSS 0.015989f
C23380 DVDD.n20525 VSS 0.015989f
C23381 DVDD.n20526 VSS 0.007995f
C23382 DVDD.n20527 VSS 0.015989f
C23383 DVDD.n20528 VSS 0.015989f
C23384 DVDD.n20529 VSS 0.45004f
C23385 DVDD.n20530 VSS 0.020374f
C23386 DVDD.n20531 VSS 0.553132f
C23387 DVDD.n20532 VSS 0.040554f
C23388 DVDD.n20533 VSS 0.015989f
C23389 DVDD.n20534 VSS 0.040554f
C23390 DVDD.n20535 VSS 0.553132f
C23391 DVDD.n20536 VSS 0.02942f
C23392 DVDD.n20537 VSS 0.02942f
C23393 DVDD.n20538 VSS 0.553132f
C23394 DVDD.n20539 VSS 0.064891f
C23395 DVDD.n20540 VSS 0.812186f
C23396 DVDD.n20541 VSS 0.812186f
C23397 DVDD.n20542 VSS 0.115237f
C23398 DVDD.t157 VSS 3.21054f
C23399 DVDD.n20543 VSS 0.115237f
C23400 DVDD.n20544 VSS 0.079947f
C23401 DVDD.n20545 VSS 0.163891f
C23402 DVDD.n20546 VSS 0.079947f
C23403 DVDD.n20547 VSS 0.079947f
C23404 DVDD.n20548 VSS 0.079947f
C23405 DVDD.n20549 VSS 0.163891f
C23406 DVDD.n20550 VSS 0.079947f
C23407 DVDD.n20551 VSS 0.079947f
C23408 DVDD.n20552 VSS 0.079947f
C23409 DVDD.n20553 VSS 0.163891f
C23410 DVDD.n20554 VSS 0.127544f
C23411 DVDD.n20555 VSS 0.079947f
C23412 DVDD.n20556 VSS 0.079947f
C23413 DVDD.n20557 VSS 0.081946f
C23414 DVDD.n20558 VSS 0.079947f
C23415 DVDD.n20559 VSS 0.081946f
C23416 DVDD.n20560 VSS 0.079947f
C23417 DVDD.n20561 VSS 0.079947f
C23418 DVDD.n20562 VSS 0.081946f
C23419 DVDD.n20563 VSS 0.079947f
C23420 DVDD.n20564 VSS 0.081946f
C23421 DVDD.n20565 VSS 0.079947f
C23422 DVDD.n20566 VSS 0.079947f
C23423 DVDD.n20567 VSS 0.081946f
C23424 DVDD.n20568 VSS 0.079947f
C23425 DVDD.n20569 VSS 0.079947f
C23426 DVDD.n20570 VSS 0.081946f
C23427 DVDD.n20571 VSS 0.081946f
C23428 DVDD.n20572 VSS 0.064086f
C23429 DVDD.n20573 VSS 0.081946f
C23430 DVDD.n20574 VSS 0.081946f
C23431 DVDD.n20575 VSS 0.079947f
C23432 DVDD.n20576 VSS 0.079947f
C23433 DVDD.n20577 VSS 0.081946f
C23434 DVDD.n20578 VSS 0.079947f
C23435 DVDD.n20579 VSS 0.079947f
C23436 DVDD.n20580 VSS 0.079947f
C23437 DVDD.n20581 VSS 0.163891f
C23438 DVDD.n20582 VSS 0.079947f
C23439 DVDD.n20583 VSS 0.079947f
C23440 DVDD.n20584 VSS 0.079947f
C23441 DVDD.n20585 VSS 0.163891f
C23442 DVDD.n20586 VSS 0.079947f
C23443 DVDD.n20587 VSS 0.079947f
C23444 DVDD.n20588 VSS 0.079947f
C23445 DVDD.n20589 VSS 0.163891f
C23446 DVDD.n20590 VSS 0.079947f
C23447 DVDD.n20591 VSS 0.079947f
C23448 DVDD.n20592 VSS 0.115237f
C23449 DVDD.n20593 VSS 0.648295f
C23450 DVDD.n20594 VSS 0.115237f
C23451 DVDD.t155 VSS 3.21054f
C23452 DVDD.n20595 VSS 0.115237f
C23453 DVDD.n20596 VSS 1.75848f
C23454 DVDD.n20602 VSS 0.064086f
C23455 DVDD.n20604 VSS 0.059122f
C23456 DVDD.n20605 VSS 0.064086f
C23457 DVDD.n20606 VSS 0.064086f
C23458 DVDD.n20607 VSS 0.064086f
C23459 DVDD.n20608 VSS 0.060025f
C23460 DVDD.n20609 VSS 0.373774f
C23461 DVDD.n20611 VSS 0.060025f
C23462 DVDD.n20612 VSS 0.064086f
C23463 DVDD.n20613 VSS 0.064086f
C23464 DVDD.n20614 VSS 0.064086f
C23465 DVDD.n20616 VSS 0.060927f
C23466 DVDD.n20617 VSS 0.055963f
C23467 DVDD.n20618 VSS 0.128173f
C23468 DVDD.n20619 VSS 0.128173f
C23469 DVDD.n20620 VSS 0.055963f
C23470 DVDD.n20621 VSS 0.128173f
C23471 DVDD.n20622 VSS 0.128173f
C23472 DVDD.n20623 VSS 0.055963f
C23473 DVDD.n20624 VSS 0.128173f
C23474 DVDD.n20625 VSS 0.055963f
C23475 DVDD.n20626 VSS 0.159414f
C23476 DVDD.n20627 VSS 0.353402f
C23477 DVDD.n20628 VSS 0.587849f
C23478 DVDD.n20629 VSS 0.128173f
C23479 DVDD.n20630 VSS 0.055963f
C23480 DVDD.n20631 VSS 0.128173f
C23481 DVDD.n20632 VSS 0.055963f
C23482 DVDD.n20633 VSS 0.128173f
C23483 DVDD.n20634 VSS 0.055963f
C23484 DVDD.n20635 VSS 0.128173f
C23485 DVDD.n20636 VSS 0.128173f
C23486 DVDD.n20637 VSS 0.128173f
C23487 DVDD.n20638 VSS 0.128173f
C23488 DVDD.n20639 VSS 0.055963f
C23489 DVDD.n20640 VSS 0.128173f
C23490 DVDD.n20641 VSS 0.055963f
C23491 DVDD.n20642 VSS 0.128173f
C23492 DVDD.n20647 VSS 0.064086f
C23493 DVDD.n20648 VSS 0.055963f
C23494 DVDD.n20649 VSS 0.128173f
C23495 DVDD.n20650 VSS 0.128173f
C23496 DVDD.n20651 VSS 0.128173f
C23497 DVDD.n20652 VSS 0.128173f
C23498 DVDD.n20653 VSS 0.128173f
C23499 DVDD.n20654 VSS 0.055963f
C23500 DVDD.n20655 VSS 0.064086f
C23501 DVDD.n20656 VSS 1.75848f
C23502 DVDD.n20657 VSS 0.064086f
C23503 DVDD.n20658 VSS 0.101545f
C23504 DVDD.n20659 VSS 0.128173f
C23505 DVDD.n20660 VSS 0.128173f
C23506 DVDD.n20661 VSS 0.128173f
C23507 DVDD.n20662 VSS 0.128173f
C23508 DVDD.n20663 VSS 0.128173f
C23509 DVDD.n20664 VSS 0.128173f
C23510 DVDD.n20665 VSS 0.128173f
C23511 DVDD.n20666 VSS 0.128173f
C23512 DVDD.n20667 VSS 0.111926f
C23513 DVDD.n20668 VSS 0.128173f
C23514 DVDD.n20669 VSS 0.055963f
C23515 DVDD.n20670 VSS 0.128173f
C23516 DVDD.n20671 VSS 0.128173f
C23517 DVDD.n20672 VSS 0.128173f
C23518 DVDD.n20673 VSS 0.128173f
C23519 DVDD.n20674 VSS 0.055963f
C23520 DVDD.n20675 VSS 0.128173f
C23521 DVDD.n20676 VSS 0.055963f
C23522 DVDD.n20677 VSS 0.128173f
C23523 DVDD.n20678 VSS 0.055963f
C23524 DVDD.n20679 VSS 0.128173f
C23525 DVDD.n20680 VSS 0.128173f
C23526 DVDD.n20681 VSS 0.128173f
C23527 DVDD.n20682 VSS 0.128173f
C23528 DVDD.n20683 VSS 0.055963f
C23529 DVDD.n20684 VSS 0.128173f
C23530 DVDD.n20685 VSS 0.055963f
C23531 DVDD.n20686 VSS 0.128173f
C23532 DVDD.n20687 VSS 0.055963f
C23533 DVDD.n20688 VSS 0.128173f
C23534 DVDD.n20689 VSS 0.128173f
C23535 DVDD.n20690 VSS 0.128173f
C23536 DVDD.n20691 VSS 0.128173f
C23537 DVDD.n20692 VSS 0.055963f
C23538 DVDD.n20693 VSS 0.128173f
C23539 DVDD.n20694 VSS 0.055963f
C23540 DVDD.n20695 VSS 0.128173f
C23541 DVDD.n20696 VSS 0.128173f
C23542 DVDD.n20697 VSS 0.128173f
C23543 DVDD.n20698 VSS 0.128173f
C23544 DVDD.n20699 VSS 0.128173f
C23545 DVDD.n20700 VSS 0.128173f
C23546 DVDD.n20701 VSS 0.128173f
C23547 DVDD.n20702 VSS 0.128173f
C23548 DVDD.n20703 VSS 0.128173f
C23549 DVDD.n20704 VSS 0.092068f
C23550 DVDD.n20705 VSS 0.128173f
C23551 DVDD.n20706 VSS 0.055963f
C23552 DVDD.n20707 VSS 0.128173f
C23553 DVDD.n20708 VSS 0.055963f
C23554 DVDD.n20709 VSS 0.128173f
C23555 DVDD.n20710 VSS 0.128173f
C23556 DVDD.n20711 VSS 0.128173f
C23557 DVDD.n20712 VSS 0.128173f
C23558 DVDD.n20713 VSS 0.055963f
C23559 DVDD.n20714 VSS 0.128173f
C23560 DVDD.n20715 VSS 0.055963f
C23561 DVDD.n20716 VSS 0.128173f
C23562 DVDD.n20717 VSS 0.055963f
C23563 DVDD.n20718 VSS 0.128173f
C23564 DVDD.n20719 VSS 0.128173f
C23565 DVDD.n20720 VSS 0.128173f
C23566 DVDD.n20721 VSS 0.128173f
C23567 DVDD.n20722 VSS 0.055963f
C23568 DVDD.n20723 VSS 0.128173f
C23569 DVDD.n20724 VSS 0.055963f
C23570 DVDD.n20725 VSS 0.128173f
C23571 DVDD.n20726 VSS 0.055963f
C23572 DVDD.n20727 VSS 0.128173f
C23573 DVDD.n20728 VSS 0.128173f
C23574 DVDD.n20729 VSS 0.128173f
C23575 DVDD.n20730 VSS 0.128173f
C23576 DVDD.n20731 VSS 0.128173f
C23577 DVDD.n20732 VSS 0.128173f
C23578 DVDD.n20733 VSS 0.055963f
C23579 DVDD.n20734 VSS 0.064086f
C23580 DVDD.n20735 VSS 0.45004f
C23581 DVDD.n20736 VSS 0.064086f
C23582 DVDD.n20737 VSS 0.093873f
C23583 DVDD.n20738 VSS 0.128173f
C23584 DVDD.n20739 VSS 0.128173f
C23585 DVDD.n20740 VSS 0.128173f
C23586 DVDD.n20741 VSS 0.128173f
C23587 DVDD.n20742 VSS 0.128173f
C23588 DVDD.n20743 VSS 0.128173f
C23589 DVDD.n20744 VSS 0.128173f
C23590 DVDD.n20745 VSS 0.128173f
C23591 DVDD.n20746 VSS 0.128173f
C23592 DVDD.n20747 VSS 0.095678f
C23593 DVDD.n20748 VSS 0.128173f
C23594 DVDD.n20749 VSS 0.055963f
C23595 DVDD.n20750 VSS 0.128173f
C23596 DVDD.n20751 VSS 0.055963f
C23597 DVDD.n20752 VSS 0.128173f
C23598 DVDD.n20753 VSS 0.128173f
C23599 DVDD.n20754 VSS 0.128173f
C23600 DVDD.n20755 VSS 0.128173f
C23601 DVDD.n20756 VSS 0.055963f
C23602 DVDD.n20757 VSS 0.128173f
C23603 DVDD.n20758 VSS 0.055963f
C23604 DVDD.n20759 VSS 0.128173f
C23605 DVDD.n20760 VSS 0.055963f
C23606 DVDD.n20761 VSS 0.128173f
C23607 DVDD.n20762 VSS 0.128173f
C23608 DVDD.n20763 VSS 0.128173f
C23609 DVDD.n20764 VSS 0.128173f
C23610 DVDD.n20765 VSS 0.055963f
C23611 DVDD.n20766 VSS 0.128173f
C23612 DVDD.n20767 VSS 0.055963f
C23613 DVDD.n20768 VSS 0.128173f
C23614 DVDD.n20769 VSS 0.055963f
C23615 DVDD.n20770 VSS 0.128173f
C23616 DVDD.n20771 VSS 0.128173f
C23617 DVDD.n20772 VSS 0.128173f
C23618 DVDD.n20773 VSS 0.128173f
C23619 DVDD.n20774 VSS 0.128173f
C23620 DVDD.n20775 VSS 0.128173f
C23621 DVDD.n20776 VSS 0.055963f
C23622 DVDD.n20777 VSS 0.064086f
C23623 DVDD.n20778 VSS 0.45004f
C23624 DVDD.n20779 VSS 0.064086f
C23625 DVDD.n20780 VSS 0.090263f
C23626 DVDD.n20781 VSS 0.128173f
C23627 DVDD.n20782 VSS 0.128173f
C23628 DVDD.n20783 VSS 0.128173f
C23629 DVDD.n20784 VSS 0.128173f
C23630 DVDD.n20785 VSS 0.128173f
C23631 DVDD.n20786 VSS 0.128173f
C23632 DVDD.n20787 VSS 0.128173f
C23633 DVDD.n20788 VSS 0.128173f
C23634 DVDD.n20789 VSS 0.055963f
C23635 DVDD.n20790 VSS 0.128173f
C23636 DVDD.n20791 VSS 0.128173f
C23637 DVDD.n20792 VSS 0.128173f
C23638 DVDD.n20793 VSS 0.128173f
C23639 DVDD.n20794 VSS 0.055963f
C23640 DVDD.n20795 VSS 0.128173f
C23641 DVDD.n20796 VSS 0.055963f
C23642 DVDD.n20797 VSS 0.128173f
C23643 DVDD.n20798 VSS 0.055963f
C23644 DVDD.n20799 VSS 0.128173f
C23645 DVDD.n20800 VSS 0.128173f
C23646 DVDD.n20801 VSS 0.128173f
C23647 DVDD.n20802 VSS 0.128173f
C23648 DVDD.n20803 VSS 0.055963f
C23649 DVDD.n20804 VSS 0.128173f
C23650 DVDD.n20805 VSS 0.055963f
C23651 DVDD.n20806 VSS 0.128173f
C23652 DVDD.n20807 VSS 0.055963f
C23653 DVDD.n20808 VSS 0.128173f
C23654 DVDD.n20809 VSS 0.128173f
C23655 DVDD.n20810 VSS 0.128173f
C23656 DVDD.n20811 VSS 0.128173f
C23657 DVDD.n20812 VSS 0.055963f
C23658 DVDD.n20813 VSS 0.128173f
C23659 DVDD.n20814 VSS 0.055963f
C23660 DVDD.n20815 VSS 0.128173f
C23661 DVDD.n20816 VSS 0.11012f
C23662 DVDD.n20817 VSS 0.128173f
C23663 DVDD.n20818 VSS 0.128173f
C23664 DVDD.n20819 VSS 0.128173f
C23665 DVDD.n20820 VSS 0.128173f
C23666 DVDD.n20821 VSS 0.128173f
C23667 DVDD.n20822 VSS 0.128173f
C23668 DVDD.n20823 VSS 0.128173f
C23669 DVDD.n20824 VSS 0.128173f
C23670 DVDD.n20825 VSS 0.103351f
C23671 DVDD.n20826 VSS 0.128173f
C23672 DVDD.n20827 VSS 0.055963f
C23673 DVDD.n20828 VSS 0.128173f
C23674 DVDD.n20829 VSS 0.128173f
C23675 DVDD.n20830 VSS 0.128173f
C23676 DVDD.n20831 VSS 0.128173f
C23677 DVDD.n20832 VSS 0.055963f
C23678 DVDD.n20833 VSS 0.128173f
C23679 DVDD.n20834 VSS 0.055963f
C23680 DVDD.n20835 VSS 0.128173f
C23681 DVDD.n20836 VSS 0.055963f
C23682 DVDD.n20837 VSS 0.128173f
C23683 DVDD.n20838 VSS 0.128173f
C23684 DVDD.n20839 VSS 0.128173f
C23685 DVDD.n20840 VSS 0.128173f
C23686 DVDD.n20841 VSS 0.055963f
C23687 DVDD.n20842 VSS 0.128173f
C23688 DVDD.n20843 VSS 0.055963f
C23689 DVDD.n20844 VSS 0.128173f
C23690 DVDD.n20845 VSS 0.055963f
C23691 DVDD.n20846 VSS 0.115536f
C23692 DVDD.n20847 VSS 0.128173f
C23693 DVDD.n20848 VSS 0.065892f
C23694 DVDD.n20849 VSS 0.589426f
C23695 DVDD.n20850 VSS 0.128173f
C23696 DVDD.n20851 VSS 0.055963f
C23697 DVDD.n20852 VSS 0.06183f
C23698 DVDD.n20853 VSS 0.151899f
C23699 DVDD.n20854 VSS 0.37595f
C23700 DVDD.n20855 VSS 1.75848f
C23701 DVDD.n20856 VSS 1.75848f
C23702 DVDD.n20857 VSS 0.151899f
C23703 DVDD.n20858 VSS 0.151899f
C23704 DVDD.n20859 VSS 0.079947f
C23705 DVDD.n20860 VSS 0.079947f
C23706 DVDD.n20861 VSS 0.079947f
C23707 DVDD.n20862 VSS 0.151899f
C23708 DVDD.n20863 VSS 0.151899f
C23709 DVDD.n20864 VSS 0.118212f
C23710 DVDD.n20865 VSS 0.079947f
C23711 DVDD.n20866 VSS 0.075949f
C23712 DVDD.n20867 VSS 0.079947f
C23713 DVDD.n20868 VSS 0.075949f
C23714 DVDD.n20869 VSS 0.079947f
C23715 DVDD.n20870 VSS 0.075949f
C23716 DVDD.n20871 VSS 0.079947f
C23717 DVDD.n20872 VSS 0.075949f
C23718 DVDD.n20873 VSS 0.079947f
C23719 DVDD.n20874 VSS 0.075949f
C23720 DVDD.n20875 VSS 0.079947f
C23721 DVDD.n20876 VSS 0.075949f
C23722 DVDD.n20877 VSS 0.079947f
C23723 DVDD.n20878 VSS 0.075949f
C23724 DVDD.n20879 VSS 0.079947f
C23725 DVDD.n20880 VSS 0.079947f
C23726 DVDD.n20881 VSS 0.075949f
C23727 DVDD.n20882 VSS 0.075949f
C23728 DVDD.n20883 VSS 0.37595f
C23729 DVDD.n20884 VSS 0.075949f
C23730 DVDD.n20885 VSS 0.075949f
C23731 DVDD.n20886 VSS 0.079947f
C23732 DVDD.n20887 VSS 0.079947f
C23733 DVDD.n20888 VSS 0.079947f
C23734 DVDD.n20889 VSS 0.151899f
C23735 DVDD.n20890 VSS 0.151899f
C23736 DVDD.n20891 VSS 0.151899f
C23737 DVDD.n20892 VSS 0.079947f
C23738 DVDD.n20893 VSS 0.079947f
C23739 DVDD.n20894 VSS 0.079947f
C23740 DVDD.n20895 VSS 0.151899f
C23741 DVDD.n20896 VSS 0.151899f
C23742 DVDD.n20897 VSS 0.600859f
C23743 DVDD.n20898 VSS 0.115237f
C23744 DVDD.t158 VSS 3.21054f
C23745 DVDD.n20899 VSS 0.115237f
C23746 DVDD.n20900 VSS 0.812186f
C23747 DVDD.n20901 VSS 0.02942f
C23748 DVDD.n20902 VSS 0.02942f
C23749 DVDD.n20903 VSS 0.02942f
C23750 DVDD.n20904 VSS 0.02942f
C23751 DVDD.n20905 VSS 0.02942f
C23752 DVDD.n20906 VSS 0.02942f
C23753 DVDD.n20908 VSS 0.02942f
C23754 DVDD.n20910 VSS 0.02942f
C23755 DVDD.n20912 VSS 0.02942f
C23756 DVDD.n20914 VSS 0.02942f
C23757 DVDD.n20916 VSS 0.02942f
C23758 DVDD.n20918 VSS 0.02942f
C23759 DVDD.n20919 VSS 0.812186f
C23760 DVDD.n20920 VSS 0.02942f
C23761 DVDD.n20922 VSS 0.553132f
C23762 DVDD.n20923 VSS 0.561029f
C23763 DVDD.n20924 VSS 0.040896f
C23764 DVDD.n20925 VSS 0.040554f
C23765 DVDD.n20926 VSS 0.457979f
C23766 DVDD.n20928 VSS 0.45004f
C23767 DVDD.n20929 VSS 0.064086f
C23768 DVDD.n20930 VSS 0.081946f
C23769 DVDD.n20931 VSS 0.096137f
C23770 DVDD.n20932 VSS 0.13448f
C23771 DVDD.n20933 VSS 0.066473f
C23772 DVDD.n20934 VSS 0.007995f
C23773 DVDD.n20935 VSS 0.015989f
C23774 DVDD.n20936 VSS 0.015989f
C23775 DVDD.n20937 VSS 0.015989f
C23776 DVDD.n20938 VSS 0.015989f
C23777 DVDD.n20939 VSS 0.015989f
C23778 DVDD.n20940 VSS 0.015989f
C23779 DVDD.n20941 VSS 0.015989f
C23780 DVDD.n20942 VSS 0.015989f
C23781 DVDD.n20943 VSS 0.015989f
C23782 DVDD.n20944 VSS 0.015989f
C23783 DVDD.n20945 VSS 0.015989f
C23784 DVDD.n20946 VSS 0.015989f
C23785 DVDD.n20947 VSS 0.015989f
C23786 DVDD.n20948 VSS 0.007995f
C23787 DVDD.n20949 VSS 0.035267f
C23788 DVDD.t156 VSS 1.03157f
C23789 DVDD.n20950 VSS 0.035267f
C23790 DVDD.n20951 VSS 0.007995f
C23791 DVDD.n20952 VSS 0.015989f
C23792 DVDD.n20953 VSS 0.015989f
C23793 DVDD.n20954 VSS 0.015989f
C23794 DVDD.n20955 VSS 0.015989f
C23795 DVDD.n20956 VSS 0.015989f
C23796 DVDD.n20957 VSS 0.015989f
C23797 DVDD.n20958 VSS 0.015989f
C23798 DVDD.n20959 VSS 0.015989f
C23799 DVDD.n20960 VSS 0.015989f
C23800 DVDD.n20961 VSS 0.015989f
C23801 DVDD.n20962 VSS 0.015989f
C23802 DVDD.n20963 VSS 0.015989f
C23803 DVDD.n20964 VSS 0.015989f
C23804 DVDD.n20965 VSS 0.007995f
C23805 DVDD.n20966 VSS 0.066473f
C23806 DVDD.n20967 VSS 0.13448f
C23807 DVDD.n20968 VSS 0.096197f
C23808 DVDD.n20969 VSS 0.081946f
C23809 DVDD.n20970 VSS 0.064086f
C23810 DVDD.n20971 VSS 0.128866f
C23811 DVDD.n20972 VSS 0.096137f
C23812 DVDD.n20973 VSS 0.13448f
C23813 DVDD.n20974 VSS 0.596461f
C23814 DVDD.n20975 VSS 0.015989f
C23815 DVDD.n20976 VSS 0.015989f
C23816 DVDD.n20977 VSS 0.015989f
C23817 DVDD.n20978 VSS 0.617235f
C23818 DVDD.n20979 VSS 0.015989f
C23819 DVDD.n20980 VSS 0.015989f
C23820 DVDD.n20981 VSS 0.020374f
C23821 DVDD.n20982 VSS 0.553132f
C23822 DVDD.n20983 VSS 0.075212f
C23823 DVDD.n20984 VSS 0.02942f
C23824 DVDD.n20985 VSS 0.02942f
C23825 DVDD.n20986 VSS 0.02942f
C23826 DVDD.n20987 VSS 0.02942f
C23827 DVDD.n20988 VSS 0.02942f
C23828 DVDD.n20989 VSS 0.02942f
C23829 DVDD.n20991 VSS 0.02942f
C23830 DVDD.n20994 VSS 0.02942f
C23831 DVDD.n20997 VSS 0.02942f
C23832 DVDD.n21000 VSS 0.02942f
C23833 DVDD.n21003 VSS 0.02942f
C23834 DVDD.n21006 VSS 0.02942f
C23835 DVDD.n21009 VSS 0.02942f
C23836 DVDD.n21011 VSS 0.02942f
C23837 DVDD.n21012 VSS 0.553132f
C23838 DVDD.n21013 VSS 0.319382f
C23839 DVDD.n21014 VSS -0.09737f
C23840 DVDD.n21015 VSS 1.94148f
C23841 DVDD.n21016 VSS 1.35823f
C23842 DVDD.n21017 VSS 1.94148f
C23843 DVDD.n21018 VSS -0.09737f
C23844 DVDD.n21019 VSS 0.319382f
C23845 DVDD.n21020 VSS 0.02942f
C23846 DVDD.n21021 VSS 0.02942f
C23847 DVDD.n21022 VSS 0.02942f
C23848 DVDD.n21023 VSS 0.02942f
C23849 DVDD.n21024 VSS 0.02942f
C23850 DVDD.n21025 VSS 0.02942f
C23851 DVDD.n21027 VSS 0.02942f
C23852 DVDD.n21030 VSS 0.02942f
C23853 DVDD.n21033 VSS 0.02942f
C23854 DVDD.n21036 VSS 0.02942f
C23855 DVDD.n21039 VSS 0.02942f
C23856 DVDD.n21042 VSS 0.02942f
C23857 DVDD.n21044 VSS 0.02942f
C23858 DVDD.n21047 VSS 0.02942f
C23859 DVDD.n21048 VSS 0.553132f
C23860 DVDD.n21049 VSS 0.075212f
C23861 DVDD.n21050 VSS 0.075212f
C23862 DVDD.n21051 VSS 0.553132f
C23863 DVDD.n21052 VSS 0.553132f
C23864 DVDD.n21053 VSS 0.035267f
C23865 DVDD.t160 VSS 1.03157f
C23866 DVDD.n21054 VSS 0.035267f
C23867 DVDD.n21055 VSS 0.617235f
C23868 DVDD.n21056 VSS 0.015989f
C23869 DVDD.n21057 VSS 0.015989f
C23870 DVDD.n21058 VSS 0.040554f
C23871 DVDD.n21059 VSS 0.553132f
C23872 DVDD.n21061 VSS 0.02942f
C23873 DVDD.n21062 VSS 0.02942f
C23874 DVDD.n21063 VSS 0.02942f
C23875 DVDD.n21064 VSS 0.02942f
C23876 DVDD.n21065 VSS 0.02942f
C23877 DVDD.n21066 VSS 0.02942f
C23878 DVDD.n21068 VSS 0.02942f
C23879 DVDD.n21070 VSS 0.02942f
C23880 DVDD.n21072 VSS 0.02942f
C23881 DVDD.n21074 VSS 0.02942f
C23882 DVDD.n21076 VSS 0.02942f
C23883 DVDD.n21078 VSS 0.02942f
C23884 DVDD.n21080 VSS 0.02942f
C23885 DVDD.n21081 VSS 0.553132f
C23886 DVDD.n21082 VSS 0.064891f
C23887 DVDD.n21083 VSS 0.081946f
C23888 DVDD.n21088 VSS 0.064086f
C23889 DVDD.n21094 VSS 0.061379f
C23890 DVDD.n21095 VSS 0.064086f
C23891 DVDD.n21096 VSS 0.064086f
C23892 DVDD.n21097 VSS 0.064086f
C23893 DVDD.n21099 VSS 0.060476f
C23894 DVDD.n21100 VSS 0.055963f
C23895 DVDD.n21101 VSS 0.128173f
C23896 DVDD.n21102 VSS 0.055963f
C23897 DVDD.n21103 VSS 0.128173f
C23898 DVDD.n21104 VSS 0.128173f
C23899 DVDD.n21105 VSS 0.128173f
C23900 DVDD.n21106 VSS 0.128173f
C23901 DVDD.n21107 VSS 0.128173f
C23902 DVDD.n21108 VSS 0.055963f
C23903 DVDD.n21109 VSS 0.128173f
C23904 DVDD.n21110 VSS 0.055963f
C23905 DVDD.n21111 VSS 0.128173f
C23906 DVDD.n21112 VSS 0.055963f
C23907 DVDD.n21113 VSS 0.128173f
C23908 DVDD.n21114 VSS 0.055963f
C23909 DVDD.n21115 VSS 0.128173f
C23910 DVDD.n21116 VSS 0.128173f
C23911 DVDD.n21117 VSS 0.128173f
C23912 DVDD.n21118 VSS 0.128173f
C23913 DVDD.n21119 VSS 0.128173f
C23914 DVDD.n21120 VSS 0.128173f
C23915 DVDD.n21121 VSS 0.055963f
C23916 DVDD.n21122 VSS 0.128173f
C23917 DVDD.n21123 VSS 0.128173f
C23918 DVDD.n21124 VSS 0.055963f
C23919 DVDD.n21125 VSS 0.128173f
C23920 DVDD.n21126 VSS 0.055963f
C23921 DVDD.n21127 VSS 0.128173f
C23922 DVDD.n21128 VSS 0.055963f
C23923 DVDD.n21129 VSS 0.128173f
C23924 DVDD.n21130 VSS 0.055963f
C23925 DVDD.n21131 VSS 0.128173f
C23926 DVDD.n21132 VSS 0.128173f
C23927 DVDD.n21133 VSS 0.128173f
C23928 DVDD.n21134 VSS 0.055963f
C23929 DVDD.n21135 VSS 0.128173f
C23930 DVDD.n21136 VSS 0.055963f
C23931 DVDD.n21137 VSS 0.128173f
C23932 DVDD.n21138 VSS 0.128173f
C23933 DVDD.n21139 VSS 0.128173f
C23934 DVDD.n21140 VSS 0.128173f
C23935 DVDD.n21141 VSS 0.128173f
C23936 DVDD.n21142 VSS 0.055963f
C23937 DVDD.n21143 VSS 0.128173f
C23938 DVDD.n21144 VSS 0.055963f
C23939 DVDD.n21145 VSS 0.128173f
C23940 DVDD.n21146 VSS 0.128173f
C23941 DVDD.n21147 VSS 0.128173f
C23942 DVDD.n21148 VSS 0.128173f
C23943 DVDD.n21149 VSS 0.128173f
C23944 DVDD.n21150 VSS 0.128173f
C23945 DVDD.n21151 VSS 0.128173f
C23946 DVDD.n21152 VSS 0.128173f
C23947 DVDD.n21153 VSS 0.128173f
C23948 DVDD.n21154 VSS 0.128173f
C23949 DVDD.n21155 VSS 0.128173f
C23950 DVDD.n21156 VSS 0.128173f
C23951 DVDD.n21157 VSS 0.128173f
C23952 DVDD.n21158 VSS 0.128173f
C23953 DVDD.n21159 VSS 0.093873f
C23954 DVDD.n21160 VSS 0.128173f
C23955 DVDD.n21161 VSS 0.055963f
C23956 DVDD.n21162 VSS 0.128173f
C23957 DVDD.n21163 VSS 0.128173f
C23958 DVDD.n21164 VSS 0.128173f
C23959 DVDD.n21165 VSS 0.128173f
C23960 DVDD.n21166 VSS 0.128173f
C23961 DVDD.n21167 VSS 0.055963f
C23962 DVDD.n21168 VSS 0.128173f
C23963 DVDD.n21169 VSS 0.055963f
C23964 DVDD.n21170 VSS 0.128173f
C23965 DVDD.n21171 VSS 0.128173f
C23966 DVDD.n21172 VSS 0.128173f
C23967 DVDD.n21173 VSS 0.128173f
C23968 DVDD.n21174 VSS 0.128173f
C23969 DVDD.n21175 VSS 0.055963f
C23970 DVDD.n21176 VSS 0.128173f
C23971 DVDD.n21177 VSS 0.055963f
C23972 DVDD.n21178 VSS 0.128173f
C23973 DVDD.n21179 VSS 0.128173f
C23974 DVDD.n21180 VSS 0.128173f
C23975 DVDD.n21181 VSS 0.128173f
C23976 DVDD.n21182 VSS 0.128173f
C23977 DVDD.n21183 VSS 0.055963f
C23978 DVDD.n21184 VSS 0.064086f
C23979 DVDD.n21185 VSS 0.081946f
C23980 DVDD.n21186 VSS 0.064086f
C23981 DVDD.n21187 VSS 0.092068f
C23982 DVDD.n21188 VSS 0.128173f
C23983 DVDD.n21189 VSS 0.128173f
C23984 DVDD.n21190 VSS 0.128173f
C23985 DVDD.n21191 VSS 0.128173f
C23986 DVDD.n21192 VSS 0.128173f
C23987 DVDD.n21193 VSS 0.128173f
C23988 DVDD.n21194 VSS 0.055963f
C23989 DVDD.n21195 VSS 0.128173f
C23990 DVDD.n21196 VSS 0.055963f
C23991 DVDD.n21197 VSS 0.128173f
C23992 DVDD.n21198 VSS 0.128173f
C23993 DVDD.n21199 VSS 0.128173f
C23994 DVDD.n21200 VSS 0.128173f
C23995 DVDD.n21201 VSS 0.128173f
C23996 DVDD.n21202 VSS 0.055963f
C23997 DVDD.n21203 VSS 0.128173f
C23998 DVDD.n21204 VSS 0.055963f
C23999 DVDD.n21205 VSS 0.128173f
C24000 DVDD.n21206 VSS 0.128173f
C24001 DVDD.n21207 VSS 0.128173f
C24002 DVDD.n21208 VSS 0.128173f
C24003 DVDD.n21209 VSS 0.128173f
C24004 DVDD.n21210 VSS 0.055963f
C24005 DVDD.n21211 VSS 0.056865f
C24006 DVDD.n21212 VSS 0.081946f
C24007 DVDD.n21213 VSS 0.064086f
C24008 DVDD.n21214 VSS 1.37721f
C24009 DVDD.n21215 VSS 0.163891f
C24010 DVDD.n21216 VSS 0.124756f
C24011 DVDD.n21217 VSS 0.163891f
C24012 DVDD.n21218 VSS 0.035087f
C24013 DVDD.n21219 VSS 0.016634f
C24014 DVDD.n21220 VSS 0.124756f
C24015 DVDD.n21221 VSS 0.038113f
C24016 DVDD.n21222 VSS 0.151899f
C24017 DVDD.n21223 VSS 0.137328f
C24018 DVDD.n21224 VSS 0.11992f
C24019 DVDD.n21225 VSS 0.274656f
C24020 DVDD.n21226 VSS 0.209861f
C24021 DVDD.n21227 VSS 0.274656f
C24022 DVDD.n21228 VSS 0.261596f
C24023 DVDD.n21229 VSS 0.274656f
C24024 DVDD.n21230 VSS 0.780268f
C24025 DVDD.n21231 VSS 0.274656f
C24026 DVDD.n21232 VSS 0.11992f
C24027 DVDD.n21233 VSS 0.132493f
C24028 DVDD.n21234 VSS 0.163891f
C24029 DVDD.n21235 VSS 0.017666f
C24030 DVDD.n21236 VSS 0.015989f
C24031 DVDD.n21237 VSS 0.01831f
C24032 DVDD.n21238 VSS 0.015989f
C24033 DVDD.n21239 VSS 0.027981f
C24034 DVDD.n21240 VSS 0.036621f
C24035 DVDD.n21241 VSS 0.036621f
C24036 DVDD.n21242 VSS 0.103874f
C24037 DVDD.n21243 VSS 0.036621f
C24038 DVDD.n21244 VSS 0.036621f
C24039 DVDD.n21245 VSS 0.015989f
C24040 DVDD.n21246 VSS 0.036277f
C24041 DVDD.n21247 VSS 1.37721f
C24042 DVDD.n21248 VSS 0.272424f
C24043 DVDD.n21249 VSS 0.261596f
C24044 DVDD.n21250 VSS 0.274656f
C24045 DVDD.n21251 VSS 0.780268f
C24046 DVDD.n21252 VSS 0.274656f
C24047 DVDD.n21253 VSS 0.11992f
C24048 DVDD.n21254 VSS 0.137328f
C24049 DVDD.n21255 VSS 0.163891f
C24050 DVDD.n21256 VSS 0.163891f
C24051 DVDD.n21257 VSS 0.137328f
C24052 DVDD.n21258 VSS 0.163891f
C24053 DVDD.n21259 VSS 0.137328f
C24054 DVDD.n21260 VSS 0.151899f
C24055 DVDD.n21261 VSS 0.039504f
C24056 DVDD.n21262 VSS 0.034496f
C24057 DVDD.n21263 VSS 0.06037f
C24058 DVDD.n21264 VSS 0.079009f
C24059 DVDD.n21265 VSS 0.079009f
C24060 DVDD.n21266 VSS 0.225252f
C24061 DVDD.n21267 VSS 0.079009f
C24062 DVDD.n21268 VSS 0.079009f
C24063 DVDD.n21269 VSS 0.034496f
C24064 DVDD.n21270 VSS 0.078141f
C24065 DVDD.n21271 VSS 0.469785f
C24066 DVDD.n21272 VSS 1.20049f
C24067 DVDD.n21273 VSS 0.002548f
C24068 DVDD.n21274 VSS 0.003773f
C24069 DVDD.n21275 VSS 0.006035f
C24070 DVDD.n21276 VSS 0.852657f
C24071 DVDD.n21277 VSS 0.006035f
C24072 DVDD.n21278 VSS 0.003773f
C24073 DVDD.n21279 VSS 0.005096f
C24074 DVDD.n21280 VSS 0.005096f
C24075 DVDD.n21281 VSS 0.006035f
C24076 DVDD.n21282 VSS 0.710547f
C24077 DVDD.n21283 VSS 0.923711f
C24078 DVDD.n21284 VSS 0.006035f
C24079 DVDD.n21285 VSS 0.005096f
C24080 DVDD.n21286 VSS 0.005096f
C24081 DVDD.n21287 VSS 0.005096f
C24082 DVDD.n21288 VSS 0.006035f
C24083 DVDD.n21289 VSS 0.67502f
C24084 DVDD.n21290 VSS 0.006035f
C24085 DVDD.n21291 VSS 0.005096f
C24086 DVDD.n21292 VSS 0.005096f
C24087 DVDD.n21293 VSS 0.005096f
C24088 DVDD.n21294 VSS 0.006035f
C24089 DVDD.t71 VSS 0.461856f
C24090 DVDD.n21295 VSS 0.568438f
C24091 DVDD.n21296 VSS 0.006035f
C24092 DVDD.n21297 VSS 0.005096f
C24093 DVDD.n21298 VSS 0.005096f
C24094 DVDD.n21299 VSS 0.005096f
C24095 DVDD.n21300 VSS 0.006035f
C24096 DVDD.n21301 VSS 0.888184f
C24097 DVDD.n21302 VSS 0.006035f
C24098 DVDD.n21303 VSS 0.005096f
C24099 DVDD.n21304 VSS 0.005096f
C24100 DVDD.n21305 VSS 0.005096f
C24101 DVDD.n21306 VSS 0.006035f
C24102 DVDD.n21307 VSS 0.746075f
C24103 DVDD.n21308 VSS 0.923711f
C24104 DVDD.n21309 VSS 0.006035f
C24105 DVDD.n21310 VSS 0.005096f
C24106 DVDD.n21311 VSS 0.005096f
C24107 DVDD.n21312 VSS 0.005096f
C24108 DVDD.n21313 VSS 0.006035f
C24109 DVDD.n21314 VSS 0.639492f
C24110 DVDD.n21315 VSS 0.006035f
C24111 DVDD.n21316 VSS 0.005096f
C24112 DVDD.n21317 VSS 0.005096f
C24113 DVDD.n21318 VSS 0.005096f
C24114 DVDD.n21319 VSS 0.005096f
C24115 DVDD.n21320 VSS 0.006035f
C24116 DVDD.t65 VSS 0.461856f
C24117 DVDD.n21321 VSS 0.603965f
C24118 DVDD.n21322 VSS 0.006035f
C24119 DVDD.n21323 VSS 0.005096f
C24120 DVDD.n21324 VSS 0.005096f
C24121 DVDD.n21325 VSS 0.005096f
C24122 DVDD.n21326 VSS 0.005096f
C24123 DVDD.n21327 VSS 0.006035f
C24124 DVDD.n21328 VSS 0.003332f
C24125 DVDD.n21330 VSS 0.006035f
C24126 DVDD.n21331 VSS 0.134427f
C24127 DVDD.n21332 VSS 0.122822f
C24128 DVDD.n21333 VSS 0.034496f
C24129 DVDD.n21334 VSS 0.079009f
C24130 DVDD.n21335 VSS 0.079009f
C24131 DVDD.n21336 VSS 0.058144f
C24132 DVDD.n21337 VSS 0.079009f
C24133 DVDD.n21338 VSS 0.034496f
C24134 DVDD.n21339 VSS 0.11992f
C24135 DVDD.n21340 VSS 0.01831f
C24136 DVDD.n21341 VSS 0.02695f
C24137 DVDD.n21342 VSS 0.015989f
C24138 DVDD.n21343 VSS 0.036621f
C24139 DVDD.n21344 VSS 0.036964f
C24140 DVDD.n21345 VSS 0.016376f
C24141 DVDD.n21346 VSS 0.015989f
C24142 DVDD.n21347 VSS 0.036621f
C24143 DVDD.n21348 VSS 0.037194f
C24144 DVDD.n21349 VSS 0.105852f
C24145 DVDD.n21350 VSS 0.036621f
C24146 DVDD.n21351 VSS 0.036621f
C24147 DVDD.n21352 VSS 0.015989f
C24148 DVDD.n21353 VSS 0.01831f
C24149 DVDD.n21354 VSS 0.163891f
C24150 DVDD.n21355 VSS 0.137328f
C24151 DVDD.n21356 VSS 0.163891f
C24152 DVDD.n21357 VSS 0.137328f
C24153 DVDD.n21358 VSS 0.039504f
C24154 DVDD.n21359 VSS 0.151899f
C24155 DVDD.n21360 VSS 0.151899f
C24156 DVDD.n21361 VSS 0.039504f
C24157 DVDD.n21362 VSS 0.039504f
C24158 DVDD.n21363 VSS 0.034496f
C24159 DVDD.n21364 VSS 0.079009f
C24160 DVDD.n21365 VSS 0.229561f
C24161 DVDD.n21366 VSS 0.079206f
C24162 DVDD.n21367 VSS 0.079603f
C24163 DVDD.n21368 VSS 0.035331f
C24164 DVDD.n21369 VSS 0.142712f
C24165 DVDD.n21370 VSS 0.075949f
C24166 DVDD.n21371 VSS 0.002548f
C24167 DVDD.n21372 VSS 0.005096f
C24168 DVDD.n21374 VSS 0.006035f
C24169 DVDD.n21375 VSS 0.005096f
C24170 DVDD.n21377 VSS 0.006035f
C24171 DVDD.n21378 VSS 0.005096f
C24172 DVDD.n21380 VSS 0.006035f
C24173 DVDD.n21381 VSS 0.005096f
C24174 DVDD.n21383 VSS 0.006035f
C24175 DVDD.n21384 VSS 0.005096f
C24176 DVDD.n21386 VSS 0.006035f
C24177 DVDD.n21387 VSS 0.005096f
C24178 DVDD.n21389 VSS 0.006035f
C24179 DVDD.n21390 VSS 0.005096f
C24180 DVDD.n21392 VSS 0.006035f
C24181 DVDD.n21393 VSS 0.005096f
C24182 DVDD.n21395 VSS 0.006035f
C24183 DVDD.n21396 VSS 0.005096f
C24184 DVDD.n21398 VSS 0.006035f
C24185 DVDD.n21399 VSS 0.005096f
C24186 DVDD.n21401 VSS 0.006035f
C24187 DVDD.n21403 VSS 0.006035f
C24188 DVDD.n21404 VSS 0.006035f
C24189 DVDD.n21405 VSS 0.005096f
C24190 DVDD.n21406 VSS 0.005096f
C24191 DVDD.n21407 VSS 0.005096f
C24192 DVDD.n21408 VSS 0.006035f
C24193 DVDD.n21410 VSS 0.006035f
C24194 DVDD.n21411 VSS 0.006035f
C24195 DVDD.n21412 VSS 0.005096f
C24196 DVDD.n21413 VSS 0.005096f
C24197 DVDD.n21414 VSS 0.005096f
C24198 DVDD.n21415 VSS 0.006035f
C24199 DVDD.n21417 VSS 0.006035f
C24200 DVDD.n21418 VSS 0.006035f
C24201 DVDD.n21419 VSS 0.005096f
C24202 DVDD.n21420 VSS 0.005096f
C24203 DVDD.n21421 VSS 0.005096f
C24204 DVDD.n21422 VSS 0.006035f
C24205 DVDD.n21424 VSS 0.006035f
C24206 DVDD.n21425 VSS 0.006035f
C24207 DVDD.n21426 VSS 0.005096f
C24208 DVDD.n21427 VSS 0.005096f
C24209 DVDD.n21428 VSS 0.005096f
C24210 DVDD.n21429 VSS 0.006035f
C24211 DVDD.n21431 VSS 0.006035f
C24212 DVDD.n21432 VSS 0.006035f
C24213 DVDD.n21433 VSS 0.005096f
C24214 DVDD.n21434 VSS 0.005096f
C24215 DVDD.n21435 VSS 0.005096f
C24216 DVDD.n21436 VSS 0.006035f
C24217 DVDD.n21438 VSS 0.006035f
C24218 DVDD.n21439 VSS 0.006035f
C24219 DVDD.n21440 VSS 0.004581f
C24220 DVDD.n21441 VSS 0.081946f
C24221 DVDD.n21442 VSS 0.002548f
C24222 DVDD.n21443 VSS 0.003062f
C24223 DVDD.n21444 VSS 0.005096f
C24224 DVDD.n21445 VSS 0.006035f
C24225 DVDD.n21447 VSS 0.006035f
C24226 DVDD.n21448 VSS 0.006035f
C24227 DVDD.n21449 VSS 0.005096f
C24228 DVDD.n21450 VSS 0.005096f
C24229 DVDD.n21451 VSS 0.005096f
C24230 DVDD.n21452 VSS 0.006035f
C24231 DVDD.n21454 VSS 0.006035f
C24232 DVDD.n21455 VSS 0.006035f
C24233 DVDD.n21456 VSS 0.005096f
C24234 DVDD.n21457 VSS 0.005096f
C24235 DVDD.n21458 VSS 0.005096f
C24236 DVDD.n21459 VSS 0.006035f
C24237 DVDD.n21461 VSS 0.006035f
C24238 DVDD.n21462 VSS 0.006035f
C24239 DVDD.n21463 VSS 0.005096f
C24240 DVDD.n21464 VSS 0.005096f
C24241 DVDD.n21465 VSS 0.005096f
C24242 DVDD.n21466 VSS 0.006035f
C24243 DVDD.n21468 VSS 0.006035f
C24244 DVDD.n21469 VSS 0.006035f
C24245 DVDD.n21470 VSS 0.005096f
C24246 DVDD.n21471 VSS 0.005096f
C24247 DVDD.n21472 VSS 0.005096f
C24248 DVDD.n21473 VSS 0.006035f
C24249 DVDD.n21475 VSS 0.006035f
C24250 DVDD.n21476 VSS 0.006035f
C24251 DVDD.n21477 VSS 0.005096f
C24252 DVDD.n21478 VSS 0.005096f
C24253 DVDD.n21479 VSS 0.004312f
C24254 DVDD.n21480 VSS 0.006035f
C24255 DVDD.n21482 VSS 0.006035f
C24256 DVDD.n21483 VSS 0.006035f
C24257 DVDD.n21484 VSS 0.005096f
C24258 DVDD.n21485 VSS 0.005096f
C24259 DVDD.n21486 VSS 0.005096f
C24260 DVDD.n21487 VSS 0.006035f
C24261 DVDD.n21489 VSS 0.006035f
C24262 DVDD.n21490 VSS 0.006035f
C24263 DVDD.n21492 VSS 0.006035f
C24264 DVDD.n21493 VSS 0.005096f
C24265 DVDD.n21494 VSS 0.007098f
C24266 DVDD.n21495 VSS 0.005543f
C24267 DVDD.n21496 VSS 0.00618f
C24268 DVDD.n21497 VSS 1.14576f
C24269 DVDD.n21498 VSS 0.00618f
C24270 DVDD.n21499 VSS 0.008791f
C24271 DVDD.n21501 VSS 0.015142f
C24272 DVDD.n21502 VSS 0.015189f
C24273 DVDD.n21503 VSS 0.00362f
C24274 DVDD.n21504 VSS 0.014838f
C24275 DVDD.n21505 VSS 0.004802f
C24276 DVDD.n21506 VSS 0.006035f
C24277 DVDD.n21508 VSS 0.006035f
C24278 DVDD.n21509 VSS 0.006035f
C24279 DVDD.n21510 VSS 0.005096f
C24280 DVDD.n21511 VSS 0.005096f
C24281 DVDD.n21512 VSS 0.005096f
C24282 DVDD.n21513 VSS 0.006035f
C24283 DVDD.n21515 VSS 0.006035f
C24284 DVDD.n21516 VSS 0.006035f
C24285 DVDD.n21517 VSS 0.005096f
C24286 DVDD.n21518 VSS 0.005096f
C24287 DVDD.n21519 VSS 0.005096f
C24288 DVDD.n21520 VSS 0.006035f
C24289 DVDD.n21522 VSS 0.006035f
C24290 DVDD.n21523 VSS 0.006035f
C24291 DVDD.n21524 VSS 0.005096f
C24292 DVDD.n21525 VSS 0.005096f
C24293 DVDD.n21526 VSS 0.005096f
C24294 DVDD.n21527 VSS 0.006035f
C24295 DVDD.n21529 VSS 0.006035f
C24296 DVDD.n21530 VSS 0.006035f
C24297 DVDD.n21531 VSS 0.005096f
C24298 DVDD.n21532 VSS 0.005096f
C24299 DVDD.n21533 VSS 0.005096f
C24300 DVDD.n21534 VSS 0.006035f
C24301 DVDD.n21536 VSS 0.006035f
C24302 DVDD.n21537 VSS 0.006035f
C24303 DVDD.n21538 VSS 0.005096f
C24304 DVDD.n21539 VSS 0.005096f
C24305 DVDD.n21540 VSS 0.005096f
C24306 DVDD.n21541 VSS 0.006035f
C24307 DVDD.n21543 VSS 0.006035f
C24308 DVDD.n21544 VSS 0.006035f
C24309 DVDD.n21545 VSS 0.004581f
C24310 DVDD.n21546 VSS 0.005096f
C24311 DVDD.n21547 VSS 0.005096f
C24312 DVDD.n21548 VSS 0.006035f
C24313 DVDD.n21550 VSS 0.006035f
C24314 DVDD.n21551 VSS 0.006035f
C24315 DVDD.n21552 VSS 0.005096f
C24316 DVDD.n21553 VSS 0.005096f
C24317 DVDD.n21554 VSS 0.005096f
C24318 DVDD.n21555 VSS 0.006035f
C24319 DVDD.n21557 VSS 0.006035f
C24320 DVDD.n21558 VSS 0.006035f
C24321 DVDD.n21559 VSS 0.005096f
C24322 DVDD.n21560 VSS 0.005096f
C24323 DVDD.n21561 VSS 0.005096f
C24324 DVDD.n21562 VSS 0.006035f
C24325 DVDD.n21564 VSS 0.006035f
C24326 DVDD.n21565 VSS 0.006035f
C24327 DVDD.n21566 VSS 0.005096f
C24328 DVDD.n21567 VSS 0.005096f
C24329 DVDD.n21568 VSS 0.005096f
C24330 DVDD.n21569 VSS 0.006035f
C24331 DVDD.n21571 VSS 0.006035f
C24332 DVDD.n21572 VSS 0.006035f
C24333 DVDD.n21573 VSS 0.005096f
C24334 DVDD.n21574 VSS 0.005096f
C24335 DVDD.n21575 VSS 0.005096f
C24336 DVDD.n21576 VSS 0.006035f
C24337 DVDD.n21578 VSS 0.006035f
C24338 DVDD.n21579 VSS 0.006035f
C24339 DVDD.n21580 VSS 0.005096f
C24340 DVDD.n21581 VSS 0.005071f
C24341 DVDD.n21582 VSS 0.163891f
C24342 DVDD.n21583 VSS 0.163891f
C24343 DVDD.n21584 VSS 0.202124f
C24344 DVDD.n21585 VSS 0.11992f
C24345 DVDD.n21586 VSS 0.274656f
C24346 DVDD.n21587 VSS 0.274656f
C24347 DVDD.n21588 VSS 0.274656f
C24348 DVDD.n21589 VSS 0.274656f
C24349 DVDD.n21590 VSS 0.11992f
C24350 DVDD.n21591 VSS 0.11992f
C24351 DVDD.n21592 VSS 0.137328f
C24352 DVDD.n21593 VSS 0.163891f
C24353 DVDD.n21594 VSS 0.153978f
C24354 DVDD.n21595 VSS 0.081946f
C24355 DVDD.n21596 VSS 0.002548f
C24356 DVDD.n21597 VSS 0.002572f
C24357 DVDD.n21598 VSS 0.006035f
C24358 DVDD.n21600 VSS 0.006035f
C24359 DVDD.n21601 VSS 0.006035f
C24360 DVDD.n21602 VSS 0.005096f
C24361 DVDD.n21603 VSS 0.005096f
C24362 DVDD.n21604 VSS 0.005096f
C24363 DVDD.n21605 VSS 0.006035f
C24364 DVDD.n21607 VSS 0.006035f
C24365 DVDD.n21608 VSS 0.006035f
C24366 DVDD.n21609 VSS 0.005096f
C24367 DVDD.n21610 VSS 0.005096f
C24368 DVDD.n21611 VSS 0.005096f
C24369 DVDD.n21612 VSS 0.006035f
C24370 DVDD.n21614 VSS 0.006035f
C24371 DVDD.n21615 VSS 0.006035f
C24372 DVDD.n21616 VSS 0.005096f
C24373 DVDD.n21617 VSS 0.005096f
C24374 DVDD.n21618 VSS 0.005096f
C24375 DVDD.n21619 VSS 0.006035f
C24376 DVDD.n21621 VSS 0.006035f
C24377 DVDD.n21622 VSS 0.006035f
C24378 DVDD.n21623 VSS 0.005096f
C24379 DVDD.n21624 VSS 0.005096f
C24380 DVDD.n21625 VSS 0.005096f
C24381 DVDD.n21626 VSS 0.006035f
C24382 DVDD.n21628 VSS 0.006035f
C24383 DVDD.n21629 VSS 0.006035f
C24384 DVDD.n21630 VSS 0.005096f
C24385 DVDD.n21631 VSS 0.005096f
C24386 DVDD.n21632 VSS 0.005096f
C24387 DVDD.n21633 VSS 0.006035f
C24388 DVDD.n21635 VSS 0.006035f
C24389 DVDD.n21636 VSS 0.006035f
C24390 DVDD.n21637 VSS 0.005096f
C24391 DVDD.n21638 VSS 0.005096f
C24392 DVDD.n21639 VSS 0.005096f
C24393 DVDD.n21640 VSS 0.006035f
C24394 DVDD.n21642 VSS 0.006035f
C24395 DVDD.n21643 VSS 0.006035f
C24396 DVDD.n21644 VSS 0.002572f
C24397 DVDD.n21645 VSS 0.002548f
C24398 DVDD.n21646 VSS 0.081946f
C24399 DVDD.n21647 VSS 0.247819f
C24400 DVDD.n21648 VSS 0.134427f
C24401 DVDD.n21649 VSS 0.122822f
C24402 DVDD.n21650 VSS 0.153978f
C24403 DVDD.n21651 VSS 0.163891f
C24404 DVDD.n21652 VSS 0.137328f
C24405 DVDD.n21653 VSS 0.163891f
C24406 DVDD.n21654 VSS 0.137328f
C24407 DVDD.n21655 VSS 0.11992f
C24408 DVDD.n21656 VSS 0.274656f
C24409 DVDD.n21657 VSS 0.274656f
C24410 DVDD.n21658 VSS 0.274656f
C24411 DVDD.n21659 VSS 0.456471f
C24412 DVDD.n21660 VSS 0.456471f
C24413 DVDD.n21661 VSS 0.456471f
C24414 DVDD.n21662 VSS 0.11992f
C24415 DVDD.n21663 VSS 0.274656f
C24416 DVDD.n21664 VSS 0.274656f
C24417 DVDD.n21665 VSS 0.274656f
C24418 DVDD.n21666 VSS 0.202124f
C24419 DVDD.n21667 VSS 0.274656f
C24420 DVDD.n21668 VSS 0.274656f
C24421 DVDD.n21669 VSS 0.11992f
C24422 DVDD.n21670 VSS 0.137328f
C24423 DVDD.n21671 VSS 0.151899f
C24424 DVDD.n21672 VSS 0.151899f
C24425 DVDD.n21673 VSS 0.039504f
C24426 DVDD.n21674 VSS 0.034496f
C24427 DVDD.n21675 VSS 0.079009f
C24428 DVDD.n21676 VSS 0.058144f
C24429 DVDD.n21677 VSS 0.079009f
C24430 DVDD.n21678 VSS 0.229561f
C24431 DVDD.n21679 VSS 0.079009f
C24432 DVDD.n21680 VSS 0.079009f
C24433 DVDD.n21681 VSS 0.034496f
C24434 DVDD.n21682 VSS 0.035331f
C24435 DVDD.n21683 VSS 0.079603f
C24436 DVDD.n21684 VSS 0.296448f
C24437 DVDD.n21685 VSS 0.134427f
C24438 DVDD.n21686 VSS 0.319852f
C24439 DVDD.n21687 VSS 0.134427f
C24440 DVDD.n21688 VSS 0.122822f
C24441 DVDD.n21689 VSS 0.163891f
C24442 DVDD.n21690 VSS 0.163891f
C24443 DVDD.n21691 VSS 0.163891f
C24444 DVDD.n21692 VSS 0.137328f
C24445 DVDD.n21693 VSS 0.163891f
C24446 DVDD.n21694 VSS 0.01831f
C24447 DVDD.n21695 VSS 0.015989f
C24448 DVDD.n21696 VSS 0.036621f
C24449 DVDD.n21697 VSS 0.037178f
C24450 DVDD.n21698 VSS 0.105853f
C24451 DVDD.n21699 VSS 0.02695f
C24452 DVDD.n21700 VSS 0.036621f
C24453 DVDD.n21701 VSS 0.036621f
C24454 DVDD.n21702 VSS 0.015989f
C24455 DVDD.n21703 VSS 0.01831f
C24456 DVDD.n21704 VSS 0.163891f
C24457 DVDD.n21705 VSS 0.137328f
C24458 DVDD.n21706 VSS 0.11992f
C24459 DVDD.n21707 VSS 0.274656f
C24460 DVDD.n21708 VSS 0.274656f
C24461 DVDD.n21709 VSS 0.274656f
C24462 DVDD.n21710 VSS 0.274656f
C24463 DVDD.n21711 VSS 0.274656f
C24464 DVDD.n21712 VSS 0.456471f
C24465 DVDD.n21713 VSS 0.456471f
C24466 DVDD.n21714 VSS 0.456471f
C24467 DVDD.n21715 VSS 0.274656f
C24468 DVDD.n21716 VSS 0.274656f
C24469 DVDD.n21717 VSS 0.274656f
C24470 DVDD.n21718 VSS 0.274656f
C24471 DVDD.n21719 VSS 0.202124f
C24472 DVDD.n21720 VSS 0.202124f
C24473 DVDD.n21721 VSS 0.996184f
C24474 DVDD.n21722 VSS 0.06313f
C24475 DVDD.n21723 VSS 0.06313f
C24476 DVDD.n21724 VSS 0.085784f
C24477 DVDD.n21725 VSS 0.037455f
C24478 DVDD.n21726 VSS 0.042891f
C24479 DVDD.n21727 VSS 0.042891f
C24480 DVDD.n21728 VSS 0.037455f
C24481 DVDD.n21729 VSS 0.085784f
C24482 DVDD.n21730 VSS 0.248785f
C24483 DVDD.n21731 VSS 0.086386f
C24484 DVDD.n21732 VSS 0.0865f
C24485 DVDD.n21733 VSS 0.038361f
C24486 DVDD.n21734 VSS 0.142712f
C24487 DVDD.n21735 VSS 0.122822f
C24488 DVDD.n21736 VSS 0.134427f
C24489 DVDD.n21737 VSS 0.247819f
C24490 DVDD.n21738 VSS 0.134427f
C24491 DVDD.n21739 VSS 0.333649f
C24492 DVDD.n21740 VSS 0.333649f
C24493 DVDD.n21741 VSS 0.456471f
C24494 DVDD.n21742 VSS 0.456471f
C24495 DVDD.n21743 VSS 0.456471f
C24496 DVDD.n21744 VSS 0.274656f
C24497 DVDD.n21745 VSS 0.274656f
C24498 DVDD.n21746 VSS 0.202124f
C24499 DVDD.n21747 VSS 0.274656f
C24500 DVDD.n21748 VSS 0.274656f
C24501 DVDD.n21749 VSS 0.11992f
C24502 DVDD.n21750 VSS 0.274656f
C24503 DVDD.n21751 VSS 0.274656f
C24504 DVDD.n21752 VSS 0.11992f
C24505 DVDD.n21753 VSS 0.122822f
C24506 DVDD.n21754 VSS 0.163891f
C24507 DVDD.n21755 VSS 0.163891f
C24508 DVDD.n21756 VSS 0.163891f
C24509 DVDD.n21757 VSS 0.163891f
C24510 DVDD.n21758 VSS 0.137328f
C24511 DVDD.n21759 VSS 0.163891f
C24512 DVDD.n21760 VSS 0.137328f
C24513 DVDD.n21761 VSS 0.163891f
C24514 DVDD.n21762 VSS 0.163891f
C24515 DVDD.n21763 VSS 0.137328f
C24516 DVDD.n21764 VSS 0.037455f
C24517 DVDD.n21765 VSS 0.037455f
C24518 DVDD.n21766 VSS 0.042891f
C24519 DVDD.n21767 VSS 0.151899f
C24520 DVDD.n21768 VSS 0.151899f
C24521 DVDD.n21769 VSS 0.296448f
C24522 DVDD.n21770 VSS 0.086839f
C24523 DVDD.n21771 VSS 0.086037f
C24524 DVDD.n21772 VSS 0.248795f
C24525 DVDD.n21773 VSS 0.06313f
C24526 DVDD.n21774 VSS 0.085784f
C24527 DVDD.n21775 VSS 0.085784f
C24528 DVDD.n21776 VSS 0.037455f
C24529 DVDD.n21777 VSS 0.042891f
C24530 DVDD.n21778 VSS 0.151899f
C24531 DVDD.n21779 VSS 0.137328f
C24532 DVDD.n21780 VSS 0.151899f
C24533 DVDD.n21781 VSS 0.042891f
C24534 DVDD.n21782 VSS 0.085784f
C24535 DVDD.n21783 VSS 0.039569f
C24536 DVDD.n21784 VSS 0.084905f
C24537 DVDD.n21785 VSS 0.037455f
C24538 DVDD.n21786 VSS 0.041382f
C24539 DVDD.n21787 VSS 0.151899f
C24540 DVDD.n21788 VSS 0.124756f
C24541 DVDD.n21789 VSS 0.137328f
C24542 DVDD.n21790 VSS 0.137328f
C24543 DVDD.n21791 VSS 0.151899f
C24544 DVDD.n21792 VSS 0.081138f
C24545 DVDD.n21793 VSS 0.038965f
C24546 DVDD.n21794 VSS 0.085784f
C24547 DVDD.n21795 VSS 0.037455f
C24548 DVDD.n21796 VSS 0.037455f
C24549 DVDD.n21797 VSS 0.042891f
C24550 DVDD.n21798 VSS 0.151899f
C24551 DVDD.n21799 VSS 0.11992f
C24552 DVDD.n21800 VSS 0.163891f
C24553 DVDD.n21801 VSS 0.01831f
C24554 DVDD.n21802 VSS 0.11992f
C24555 DVDD.n21803 VSS 0.163891f
C24556 DVDD.n21804 VSS 0.132493f
C24557 DVDD.n21805 VSS 0.274656f
C24558 DVDD.n21806 VSS 0.440997f
C24559 DVDD.n21807 VSS 0.440997f
C24560 DVDD.n21808 VSS 0.325912f
C24561 DVDD.n21809 VSS 0.319852f
C24562 DVDD.n21810 VSS 0.11992f
C24563 DVDD.n21811 VSS 0.319852f
C24564 DVDD.n21812 VSS 0.036292f
C24565 DVDD.n21813 VSS 0.016634f
C24566 DVDD.n21814 VSS 0.163891f
C24567 DVDD.n21815 VSS 0.124756f
C24568 DVDD.n21816 VSS 0.01831f
C24569 DVDD.n21817 VSS 0.015989f
C24570 DVDD.n21818 VSS 0.036621f
C24571 DVDD.n21819 VSS 0.015989f
C24572 DVDD.n21820 VSS 0.027981f
C24573 DVDD.n21821 VSS 0.036621f
C24574 DVDD.n21822 VSS 0.035072f
C24575 DVDD.n21823 VSS 0.036621f
C24576 DVDD.n21824 VSS 0.103875f
C24577 DVDD.n21825 VSS 0.036621f
C24578 DVDD.n21826 VSS 0.015989f
C24579 DVDD.n21827 VSS 0.017666f
C24580 DVDD.n21828 VSS 0.163891f
C24581 DVDD.n21829 VSS 0.11992f
C24582 DVDD.n21830 VSS 0.137328f
C24583 DVDD.n21831 VSS 0.274656f
C24584 DVDD.n21832 VSS 0.209861f
C24585 DVDD.n21833 VSS 0.274656f
C24586 DVDD.n21834 VSS 0.440997f
C24587 DVDD.n21835 VSS 0.274656f
C24588 DVDD.n21836 VSS 0.11992f
C24589 DVDD.n21837 VSS 0.209861f
C24590 DVDD.n21838 VSS 0.11992f
C24591 DVDD.n21839 VSS 0.163891f
C24592 DVDD.n21840 VSS 0.01831f
C24593 DVDD.n21841 VSS 0.137328f
C24594 DVDD.n21842 VSS 0.017666f
C24595 DVDD.n21843 VSS 0.132493f
C24596 DVDD.n21844 VSS 0.036277f
C24597 DVDD.n21845 VSS 0.015989f
C24598 DVDD.n21846 VSS 0.036621f
C24599 DVDD.n21847 VSS 0.027981f
C24600 DVDD.n21848 VSS 0.01831f
C24601 DVDD.n21849 VSS 0.015989f
C24602 DVDD.n21850 VSS 0.036621f
C24603 DVDD.n21851 VSS 0.036621f
C24604 DVDD.n21852 VSS 0.103874f
C24605 DVDD.n21853 VSS 0.035087f
C24606 DVDD.n21854 VSS 0.036621f
C24607 DVDD.n21855 VSS 0.015989f
C24608 DVDD.n21856 VSS 0.016634f
C24609 DVDD.n21857 VSS 0.163891f
C24610 DVDD.n21858 VSS 0.319852f
C24611 DVDD.n21859 VSS 0.137328f
C24612 DVDD.n21860 VSS 0.11992f
C24613 DVDD.n21861 VSS 0.274656f
C24614 DVDD.n21862 VSS 0.209861f
C24615 DVDD.n21863 VSS 0.163891f
C24616 DVDD.n21864 VSS 0.163891f
C24617 DVDD.n21865 VSS 0.163891f
C24618 DVDD.n21866 VSS 0.137328f
C24619 DVDD.n21867 VSS 0.11992f
C24620 DVDD.n21868 VSS 0.274656f
C24621 DVDD.n21869 VSS 0.274656f
C24622 DVDD.n21870 VSS 0.274656f
C24623 DVDD.n21871 VSS 0.274656f
C24624 DVDD.n21872 VSS 0.274656f
C24625 DVDD.n21873 VSS 0.11992f
C24626 DVDD.n21874 VSS 0.124756f
C24627 DVDD.n21875 VSS 0.163891f
C24628 DVDD.n21876 VSS 0.132493f
C24629 DVDD.n21877 VSS 0.163891f
C24630 DVDD.n21878 VSS 0.163891f
C24631 DVDD.n21879 VSS 0.137328f
C24632 DVDD.n21880 VSS 0.11992f
C24633 DVDD.n21881 VSS 0.274656f
C24634 DVDD.n21882 VSS 0.274656f
C24635 DVDD.n21883 VSS 0.274656f
C24636 DVDD.n21884 VSS 0.274656f
C24637 DVDD.n21885 VSS 0.274656f
C24638 DVDD.n21886 VSS 0.440997f
C24639 DVDD.n21887 VSS 0.325912f
C24640 DVDD.n21888 VSS 0.325912f
C24641 DVDD.n21889 VSS 0.440997f
C24642 DVDD.n21890 VSS 0.440997f
C24643 DVDD.n21891 VSS 0.274656f
C24644 DVDD.n21892 VSS 0.274656f
C24645 DVDD.n21893 VSS 0.274656f
C24646 DVDD.n21894 VSS 0.274656f
C24647 DVDD.n21895 VSS 0.11992f
C24648 DVDD.n21896 VSS 0.041382f
C24649 DVDD.n21897 VSS 0.151899f
C24650 DVDD.n21898 VSS 0.132493f
C24651 DVDD.n21899 VSS 0.124756f
C24652 DVDD.n21900 VSS 0.163891f
C24653 DVDD.n21901 VSS 0.319852f
C24654 DVDD.n21902 VSS 0.137328f
C24655 DVDD.n21903 VSS 0.325912f
C24656 DVDD.n21904 VSS 0.440997f
C24657 DVDD.n21905 VSS 0.440997f
C24658 DVDD.n21906 VSS 0.274656f
C24659 DVDD.n21907 VSS 0.274656f
C24660 DVDD.n21908 VSS 0.274656f
C24661 DVDD.n21909 VSS 0.209861f
C24662 DVDD.n21910 VSS 0.274656f
C24663 DVDD.n21911 VSS 0.274656f
C24664 DVDD.n21912 VSS 0.11992f
C24665 DVDD.n21913 VSS 0.137328f
C24666 DVDD.n21914 VSS 0.163891f
C24667 DVDD.n21915 VSS 0.163891f
C24668 DVDD.n21916 VSS 0.137328f
C24669 DVDD.n21917 VSS 0.163891f
C24670 DVDD.n21918 VSS 0.137328f
C24671 DVDD.n21919 VSS 0.151899f
C24672 DVDD.n21920 VSS 0.042891f
C24673 DVDD.n21921 VSS 0.027184f
C24674 DVDD.n21922 VSS 0.055276f
C24675 DVDD.n21923 VSS 0.055276f
C24676 DVDD.n21924 VSS 0.085784f
C24677 DVDD.n21925 VSS 0.244133f
C24678 DVDD.n21926 VSS 0.085784f
C24679 DVDD.n21927 VSS 0.085784f
C24680 DVDD.n21928 VSS 0.037455f
C24681 DVDD.n21929 VSS 0.085223f
C24682 DVDD.n21930 VSS 0.296448f
C24683 DVDD.n21931 VSS 0.296448f
C24684 DVDD.n21932 VSS 0.151899f
C24685 DVDD.n21933 VSS 0.038965f
C24686 DVDD.n21934 VSS 0.037455f
C24687 DVDD.n21935 VSS 0.085784f
C24688 DVDD.n21936 VSS 0.081467f
C24689 DVDD.n21937 VSS 0.244123f
C24690 DVDD.n21938 VSS 0.068869f
C24691 DVDD.n21939 VSS 0.068869f
C24692 DVDD.n21940 VSS 0.03534f
C24693 DVDD.n21941 VSS 0.016915f
C24694 DVDD.n21942 VSS 0.151899f
C24695 DVDD.n21943 VSS 0.151899f
C24696 DVDD.n21944 VSS 0.992458f
C24697 DVDD.n21945 VSS 0.163891f
C24698 DVDD.n21946 VSS 0.137328f
C24699 DVDD.n21947 VSS 0.163891f
C24700 DVDD.n21948 VSS 0.163891f
C24701 DVDD.n21949 VSS 0.137328f
C24702 DVDD.n21950 VSS 0.163891f
C24703 DVDD.n21951 VSS 0.01831f
C24704 DVDD.n21952 VSS 0.015989f
C24705 DVDD.n21953 VSS 0.036621f
C24706 DVDD.n21954 VSS 0.036621f
C24707 DVDD.n21955 VSS 0.103874f
C24708 DVDD.n21956 VSS 0.035087f
C24709 DVDD.n21957 VSS 0.036621f
C24710 DVDD.n21958 VSS 0.015989f
C24711 DVDD.n21959 VSS 0.016634f
C24712 DVDD.n21960 VSS 0.163891f
C24713 DVDD.n21961 VSS 0.124756f
C24714 DVDD.n21962 VSS 0.163891f
C24715 DVDD.n21963 VSS 0.137328f
C24716 DVDD.n21964 VSS 0.319852f
C24717 DVDD.n21965 VSS 0.319852f
C24718 DVDD.n21966 VSS 0.137328f
C24719 DVDD.n21967 VSS 0.319852f
C24720 DVDD.n21968 VSS 0.036292f
C24721 DVDD.n21969 VSS 0.035072f
C24722 DVDD.n21970 VSS 0.036621f
C24723 DVDD.n21971 VSS 0.103875f
C24724 DVDD.n21972 VSS 0.036621f
C24725 DVDD.n21973 VSS 0.015989f
C24726 DVDD.n21974 VSS 0.017666f
C24727 DVDD.n21975 VSS 0.163891f
C24728 DVDD.n21976 VSS 0.132493f
C24729 DVDD.n21977 VSS 0.163891f
C24730 DVDD.n21978 VSS 0.137328f
C24731 DVDD.n21979 VSS 0.163891f
C24732 DVDD.n21980 VSS 0.163891f
C24733 DVDD.n21981 VSS 0.137328f
C24734 DVDD.n21982 VSS 0.163891f
C24735 DVDD.n21983 VSS 0.137328f
C24736 DVDD.n21984 VSS 0.163891f
C24737 DVDD.n21985 VSS 0.01831f
C24738 DVDD.n21986 VSS 0.11992f
C24739 DVDD.n21987 VSS 0.163891f
C24740 DVDD.n21988 VSS 0.11992f
C24741 DVDD.n21989 VSS 0.137328f
C24742 DVDD.n21990 VSS 0.151899f
C24743 DVDD.n21991 VSS 0.151899f
C24744 DVDD.n21992 VSS 0.034496f
C24745 DVDD.n21993 VSS 0.035331f
C24746 DVDD.n21994 VSS 0.079009f
C24747 DVDD.n21995 VSS 0.079603f
C24748 DVDD.n21996 VSS 0.058144f
C24749 DVDD.n21997 VSS 0.151899f
C24750 DVDD.n21998 VSS 0.039504f
C24751 DVDD.n21999 VSS 0.039504f
C24752 DVDD.n22000 VSS 0.034496f
C24753 DVDD.n22001 VSS 0.079009f
C24754 DVDD.n22002 VSS 0.079009f
C24755 DVDD.n22003 VSS 0.229561f
C24756 DVDD.n22004 VSS 0.079206f
C24757 DVDD.n22005 VSS 0.079009f
C24758 DVDD.n22006 VSS 0.034496f
C24759 DVDD.n22007 VSS 0.039504f
C24760 DVDD.n22008 VSS 0.151899f
C24761 DVDD.n22009 VSS 0.137328f
C24762 DVDD.n22010 VSS 0.015989f
C24763 DVDD.n22011 VSS 0.016376f
C24764 DVDD.n22012 VSS 0.036621f
C24765 DVDD.n22013 VSS 0.02695f
C24766 DVDD.n22014 VSS 0.01831f
C24767 DVDD.n22015 VSS 0.015989f
C24768 DVDD.n22016 VSS 0.036621f
C24769 DVDD.n22017 VSS 0.036621f
C24770 DVDD.n22018 VSS 0.105852f
C24771 DVDD.n22019 VSS 0.037194f
C24772 DVDD.n22020 VSS 0.036621f
C24773 DVDD.n22021 VSS 0.015989f
C24774 DVDD.n22022 VSS 0.01831f
C24775 DVDD.n22023 VSS 0.163891f
C24776 DVDD.n22024 VSS 0.137328f
C24777 DVDD.n22025 VSS 0.202124f
C24778 DVDD.n22026 VSS 0.274656f
C24779 DVDD.n22027 VSS 0.11992f
C24780 DVDD.n22028 VSS 0.274656f
C24781 DVDD.n22029 VSS 0.274656f
C24782 DVDD.n22030 VSS 0.795146f
C24783 DVDD.n22031 VSS 0.274656f
C24784 DVDD.n22032 VSS 0.11992f
C24785 DVDD.n22033 VSS 0.137328f
C24786 DVDD.n22034 VSS 0.163891f
C24787 DVDD.n22035 VSS 0.163891f
C24788 DVDD.n22036 VSS 0.137328f
C24789 DVDD.n22037 VSS 0.163891f
C24790 DVDD.n22038 VSS 0.163891f
C24791 DVDD.n22039 VSS 0.980062f
C24792 DVDD.n22040 VSS 0.06313f
C24793 DVDD.n22041 VSS 0.037455f
C24794 DVDD.n22042 VSS 0.037455f
C24795 DVDD.n22043 VSS 0.042891f
C24796 DVDD.n22044 VSS 0.151899f
C24797 DVDD.n22045 VSS 0.137328f
C24798 DVDD.n22046 VSS 0.163891f
C24799 DVDD.n22047 VSS 0.137328f
C24800 DVDD.n22048 VSS 0.163891f
C24801 DVDD.n22049 VSS 0.163891f
C24802 DVDD.n22050 VSS 0.163891f
C24803 DVDD.n22051 VSS 0.137328f
C24804 DVDD.n22052 VSS 0.11992f
C24805 DVDD.n22053 VSS 0.274656f
C24806 DVDD.n22054 VSS 0.795146f
C24807 DVDD.n22055 VSS 0.277343f
C24808 DVDD.n22056 VSS 0.277582f
C24809 DVDD.n22057 VSS 0.122822f
C24810 DVDD.n22058 VSS 0.122822f
C24811 DVDD.n22059 VSS 0.163891f
C24812 DVDD.n22060 VSS 0.163891f
C24813 DVDD.n22061 VSS 0.137328f
C24814 DVDD.n22062 VSS 0.151899f
C24815 DVDD.n22063 VSS 0.042891f
C24816 DVDD.n22064 VSS 0.037455f
C24817 DVDD.n22065 VSS 0.085784f
C24818 DVDD.n22066 VSS 0.248785f
C24819 DVDD.n22067 VSS 0.086386f
C24820 DVDD.n22068 VSS 0.0865f
C24821 DVDD.n22069 VSS 0.296448f
C24822 DVDD.n22071 VSS 0.064086f
C24823 DVDD.n22072 VSS 0.064086f
C24824 DVDD.n22073 VSS 0.057317f
C24825 DVDD.n22074 VSS 0.064086f
C24826 DVDD.n22076 VSS 0.062732f
C24827 DVDD.n22077 VSS 0.064086f
C24828 DVDD.n22078 VSS 0.064086f
C24829 DVDD.n22079 VSS 0.05145f
C24830 DVDD.n22086 VSS 0.058219f
C24831 DVDD.n22087 VSS 0.055963f
C24832 DVDD.n22088 VSS 0.589426f
C24833 DVDD.n22089 VSS 0.128173f
C24834 DVDD.n22090 VSS 0.055963f
C24835 DVDD.n22091 VSS 0.128173f
C24836 DVDD.n22092 VSS 0.128173f
C24837 DVDD.n22093 VSS 0.055963f
C24838 DVDD.n22094 VSS 0.128173f
C24839 DVDD.n22095 VSS 0.055963f
C24840 DVDD.n22096 VSS 0.128173f
C24841 DVDD.n22097 VSS 0.128173f
C24842 DVDD.n22098 VSS 0.128173f
C24843 DVDD.n22099 VSS 0.128173f
C24844 DVDD.n22100 VSS 0.055963f
C24845 DVDD.n22101 VSS 0.128173f
C24846 DVDD.n22102 VSS 0.055963f
C24847 DVDD.n22103 VSS 0.128173f
C24848 DVDD.n22104 VSS 0.055963f
C24849 DVDD.n22105 VSS 0.115536f
C24850 DVDD.n22106 VSS 0.128173f
C24851 DVDD.n22107 VSS 0.065892f
C24852 DVDD.n22108 VSS 0.076723f
C24853 DVDD.n22109 VSS 0.026627f
C24854 DVDD.n22114 VSS 0.064086f
C24855 DVDD.n22115 VSS 0.06183f
C24856 DVDD.n22116 VSS 0.055963f
C24857 DVDD.n22117 VSS 0.128173f
C24858 DVDD.n22118 VSS 0.159414f
C24859 DVDD.n22119 VSS 0.35687f
C24860 DVDD.n22120 VSS 0.37595f
C24861 DVDD.n22121 VSS 0.296448f
C24862 DVDD.n22122 VSS 0.064086f
C24863 DVDD.n22123 VSS 0.055963f
C24864 DVDD.n22124 VSS 0.128173f
C24865 DVDD.n22125 VSS 0.128173f
C24866 DVDD.n22126 VSS 0.128173f
C24867 DVDD.n22127 VSS 0.128173f
C24868 DVDD.n22128 VSS 0.128173f
C24869 DVDD.n22129 VSS 0.103351f
C24870 DVDD.n22130 VSS 0.128173f
C24871 DVDD.n22131 VSS 0.128173f
C24872 DVDD.n22132 VSS 0.128173f
C24873 DVDD.n22133 VSS 0.128173f
C24874 DVDD.n22134 VSS 0.128173f
C24875 DVDD.n22135 VSS 0.128173f
C24876 DVDD.n22136 VSS 0.128173f
C24877 DVDD.n22137 VSS 0.11012f
C24878 DVDD.n22138 VSS 0.064086f
C24879 DVDD.n22139 VSS 0.319852f
C24880 DVDD.n22140 VSS 0.064086f
C24881 DVDD.n22141 VSS 0.075821f
C24882 DVDD.n22142 VSS 0.128173f
C24883 DVDD.n22143 VSS 0.128173f
C24884 DVDD.n22144 VSS 0.128173f
C24885 DVDD.n22145 VSS 0.128173f
C24886 DVDD.n22146 VSS 0.128173f
C24887 DVDD.n22147 VSS 0.128173f
C24888 DVDD.n22148 VSS 0.128173f
C24889 DVDD.n22149 VSS 0.055963f
C24890 DVDD.n22150 VSS 0.128173f
C24891 DVDD.n22151 VSS 0.128173f
C24892 DVDD.n22152 VSS 0.128173f
C24893 DVDD.n22153 VSS 0.128173f
C24894 DVDD.n22154 VSS 0.128173f
C24895 DVDD.n22155 VSS 0.055963f
C24896 DVDD.n22156 VSS 0.062281f
C24897 DVDD.n22157 VSS 0.319852f
C24898 DVDD.n22158 VSS 0.064086f
C24899 DVDD.n22159 VSS 3.48797f
C24900 DVDD.n22160 VSS 0.064086f
C24901 DVDD.n22161 VSS 0.095678f
C24902 DVDD.n22162 VSS 0.128173f
C24903 DVDD.n22163 VSS 0.128173f
C24904 DVDD.n22164 VSS 0.128173f
C24905 DVDD.n22165 VSS 0.128173f
C24906 DVDD.n22166 VSS 0.128173f
C24907 DVDD.n22167 VSS 0.128173f
C24908 DVDD.n22168 VSS 0.128173f
C24909 DVDD.n22169 VSS 0.128173f
C24910 DVDD.n22170 VSS 0.128173f
C24911 DVDD.n22171 VSS 0.128173f
C24912 DVDD.n22172 VSS 0.128173f
C24913 DVDD.n22173 VSS 0.128173f
C24914 DVDD.n22174 VSS 0.128173f
C24915 DVDD.n22175 VSS 0.128173f
C24916 DVDD.n22176 VSS 0.128173f
C24917 DVDD.n22177 VSS 0.055963f
C24918 DVDD.n22178 VSS 0.061379f
C24919 DVDD.n22180 VSS 0.163891f
C24920 DVDD.n22181 VSS 0.064086f
C24921 DVDD.n22182 VSS 0.319852f
C24922 DVDD.n22183 VSS 0.319852f
C24923 DVDD.n22184 VSS 0.277582f
C24924 DVDD.n22185 VSS 0.319852f
C24925 DVDD.n22186 VSS 0.277582f
C24926 DVDD.n22187 VSS 0.277343f
C24927 DVDD.n22188 VSS 0.795146f
C24928 DVDD.n22189 VSS 0.274656f
C24929 DVDD.n22190 VSS 0.274656f
C24930 DVDD.n22191 VSS 0.202124f
C24931 DVDD.n22192 VSS 0.202124f
C24932 DVDD.n22193 VSS 0.99631f
C24933 DVDD.n22194 VSS 0.209861f
C24934 DVDD.n22195 VSS 0.274656f
C24935 DVDD.n22196 VSS 0.274656f
C24936 DVDD.n22197 VSS 0.274656f
C24937 DVDD.n22198 VSS 0.274656f
C24938 DVDD.n22199 VSS 0.274656f
C24939 DVDD.n22200 VSS 0.440997f
C24940 DVDD.n22201 VSS 0.440997f
C24941 DVDD.n22202 VSS 0.440997f
C24942 DVDD.n22203 VSS 0.274656f
C24943 DVDD.n22204 VSS 0.274656f
C24944 DVDD.n22205 VSS 0.274656f
C24945 DVDD.n22206 VSS 0.274656f
C24946 DVDD.n22207 VSS 0.209861f
C24947 DVDD.n22208 VSS 0.209861f
C24948 DVDD.n22209 VSS 0.757165f
C24949 DVDD.n22210 VSS 0.202124f
C24950 DVDD.n22211 VSS 0.274656f
C24951 DVDD.n22212 VSS 0.274656f
C24952 DVDD.n22213 VSS 0.274656f
C24953 DVDD.n22214 VSS 0.274656f
C24954 DVDD.n22215 VSS 0.274656f
C24955 DVDD.n22216 VSS 0.456471f
C24956 DVDD.n22217 VSS 0.456471f
C24957 DVDD.n22218 VSS 0.456471f
C24958 DVDD.n22219 VSS 0.274656f
C24959 DVDD.n22220 VSS 0.274656f
C24960 DVDD.n22221 VSS 0.274656f
C24961 DVDD.n22222 VSS 0.11992f
C24962 DVDD.n22223 VSS 0.137328f
C24963 DVDD.n22224 VSS 0.163891f
C24964 DVDD.n22225 VSS 0.163891f
C24965 DVDD.n22226 VSS 0.137328f
C24966 DVDD.n22227 VSS 0.151899f
C24967 DVDD.n22228 VSS 0.151899f
C24968 DVDD.n22229 VSS 0.979582f
C24969 DVDD.n22230 VSS 0.027184f
C24970 DVDD.n22231 VSS 0.055276f
C24971 DVDD.n22232 VSS 0.055276f
C24972 DVDD.n22233 VSS 0.085784f
C24973 DVDD.n22234 VSS 0.244123f
C24974 DVDD.n22235 VSS 0.085784f
C24975 DVDD.n22236 VSS 0.085784f
C24976 DVDD.n22237 VSS 0.037455f
C24977 DVDD.n22238 VSS 0.084905f
C24978 DVDD.n22239 VSS 0.469785f
C24979 DVDD.n22240 VSS 0.272424f
C24980 DVDD.n22241 VSS 1.37721f
C24981 DVDD.n22242 VSS 0.272424f
C24982 DVDD.n22243 VSS 1.37721f
C24983 DVDD.n22244 VSS 1.37721f
C24984 DVDD.n22246 VSS 0.163891f
C24985 DVDD.n22248 VSS 0.163891f
C24986 DVDD.n22250 VSS 0.163891f
C24987 DVDD.n22251 VSS 0.064086f
C24988 DVDD.n22252 VSS 0.081946f
C24989 DVDD.n22253 VSS 0.064086f
C24990 DVDD.n22254 VSS 0.055963f
C24991 DVDD.n22255 VSS 0.128173f
C24992 DVDD.n22256 VSS 0.128173f
C24993 DVDD.n22257 VSS 0.128173f
C24994 DVDD.n22258 VSS 0.128173f
C24995 DVDD.n22259 VSS 0.128173f
C24996 DVDD.n22260 VSS 0.090263f
C24997 DVDD.n22261 VSS 0.128173f
C24998 DVDD.n22262 VSS 0.128173f
C24999 DVDD.n22263 VSS 0.128173f
C25000 DVDD.n22264 VSS 0.128173f
C25001 DVDD.n22265 VSS 0.128173f
C25002 DVDD.n22266 VSS 0.128173f
C25003 DVDD.n22267 VSS 0.055963f
C25004 DVDD.n22268 VSS 0.128173f
C25005 DVDD.n22269 VSS 0.055963f
C25006 DVDD.n22270 VSS 0.128173f
C25007 DVDD.n22271 VSS 0.055963f
C25008 DVDD.n22272 VSS 0.128173f
C25009 DVDD.n22273 VSS 0.055963f
C25010 DVDD.n22274 VSS 0.055963f
C25011 DVDD.n22275 VSS 0.128173f
C25012 DVDD.n22276 VSS 0.128173f
C25013 DVDD.n22277 VSS 0.128173f
C25014 DVDD.n22278 VSS 0.128173f
C25015 DVDD.n22279 VSS 0.128173f
C25016 DVDD.n22280 VSS 0.055963f
C25017 DVDD.n22281 VSS 0.128173f
C25018 DVDD.n22282 VSS 0.055963f
C25019 DVDD.n22283 VSS 0.128173f
C25020 DVDD.n22284 VSS 0.128173f
C25021 DVDD.n22285 VSS 0.128173f
C25022 DVDD.n22286 VSS 0.128173f
C25023 DVDD.n22287 VSS 0.128173f
C25024 DVDD.n22288 VSS 0.055963f
C25025 DVDD.n22289 VSS 0.128173f
C25026 DVDD.n22290 VSS 0.055963f
C25027 DVDD.n22291 VSS 0.128173f
C25028 DVDD.n22292 VSS 0.128173f
C25029 DVDD.n22293 VSS 0.128173f
C25030 DVDD.n22294 VSS 0.128173f
C25031 DVDD.n22295 VSS 0.128173f
C25032 DVDD.n22296 VSS 0.055963f
C25033 DVDD.n22297 VSS 0.064086f
C25034 DVDD.n22298 VSS 0.081946f
C25035 DVDD.n22299 VSS 0.064086f
C25036 DVDD.n22300 VSS 0.055963f
C25037 DVDD.n22301 VSS 0.128173f
C25038 DVDD.n22302 VSS 0.128173f
C25039 DVDD.n22303 VSS 0.128173f
C25040 DVDD.n22304 VSS 0.128173f
C25041 DVDD.n22305 VSS 0.128173f
C25042 DVDD.n22306 VSS 0.128173f
C25043 DVDD.n22307 VSS 0.128173f
C25044 DVDD.n22308 VSS 0.128173f
C25045 DVDD.n22309 VSS 0.128173f
C25046 DVDD.n22310 VSS 0.128173f
C25047 DVDD.n22311 VSS 0.128173f
C25048 DVDD.n22312 VSS 0.128173f
C25049 DVDD.n22313 VSS 0.055963f
C25050 DVDD.n22314 VSS 0.128173f
C25051 DVDD.n22315 VSS 0.055963f
C25052 DVDD.n22316 VSS 0.128173f
C25053 DVDD.n22317 VSS 0.055963f
C25054 DVDD.n22318 VSS 0.115536f
C25055 DVDD.n22319 VSS 0.055963f
C25056 DVDD.n22320 VSS 0.128173f
C25057 DVDD.n22321 VSS 0.055963f
C25058 DVDD.n22322 VSS 0.128173f
C25059 DVDD.n22323 VSS 0.128173f
C25060 DVDD.n22324 VSS 0.128173f
C25061 DVDD.n22325 VSS 0.128173f
C25062 DVDD.n22326 VSS 0.128173f
C25063 DVDD.n22327 VSS 0.055963f
C25064 DVDD.n22328 VSS 0.128173f
C25065 DVDD.n22329 VSS 0.055963f
C25066 DVDD.n22330 VSS 0.128173f
C25067 DVDD.n22331 VSS 0.128173f
C25068 DVDD.n22332 VSS 0.128173f
C25069 DVDD.n22333 VSS 0.128173f
C25070 DVDD.n22334 VSS 0.128173f
C25071 DVDD.n22335 VSS 0.055963f
C25072 DVDD.n22337 VSS 0.115762f
C25073 DVDD.n22339 VSS 0.151899f
C25074 DVDD.n22341 VSS 0.151899f
C25075 DVDD.n22342 VSS 0.064086f
C25076 DVDD.n22343 VSS 0.112087f
C25077 DVDD.n22344 VSS 0.058219f
C25078 DVDD.n22345 VSS 0.055963f
C25079 DVDD.n22346 VSS 0.159421f
C25080 DVDD.n22347 VSS 0.35693f
C25081 DVDD.n22348 VSS 0.588875f
C25082 DVDD.n22349 VSS 0.065892f
C25083 DVDD.n22350 VSS 0.076723f
C25084 DVDD.n22351 VSS 0.026627f
C25085 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n0 VSS 5.86309f
C25086 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n1 VSS 4.42434f
C25087 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n2 VSS 3.51977f
C25088 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n3 VSS 4.29519f
C25089 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n4 VSS 4.3335f
C25090 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n5 VSS 3.51615f
C25091 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n6 VSS 4.28022f
C25092 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n7 VSS 12.436501f
C25093 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n8 VSS 3.63431f
C25094 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n9 VSS 4.29519f
C25095 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n10 VSS 0.533869f
C25096 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n11 VSS 0.430076f
C25097 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n12 VSS 3.55081f
C25098 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n13 VSS 0.482302f
C25099 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n14 VSS 0.657707f
C25100 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n15 VSS 0.63528f
C25101 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n16 VSS 0.482302f
C25102 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n17 VSS 6.15514f
C25103 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n18 VSS 0.43882f
C25104 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n19 VSS 0.262563f
C25105 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n20 VSS 0.219739f
C25106 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n21 VSS 0.262563f
C25107 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n22 VSS 0.262563f
C25108 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n23 VSS 0.262563f
C25109 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n24 VSS 0.262563f
C25110 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n25 VSS 0.262563f
C25111 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n26 VSS 0.262563f
C25112 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n27 VSS 0.262563f
C25113 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n28 VSS 0.197637f
C25114 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n29 VSS 0.262563f
C25115 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n30 VSS 0.153708f
C25116 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n31 VSS 0.262563f
C25117 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n32 VSS 0.262563f
C25118 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n33 VSS 0.262563f
C25119 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n34 VSS 0.262563f
C25120 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n35 VSS 0.262563f
C25121 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n36 VSS 0.262563f
C25122 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n37 VSS 0.262563f
C25123 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n38 VSS 0.241493f
C25124 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n39 VSS 0.504461f
C25125 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n40 VSS 3.62797f
C25126 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n41 VSS 0.262563f
C25127 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n42 VSS 0.262563f
C25128 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n43 VSS 0.219739f
C25129 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n44 VSS 0.262563f
C25130 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n45 VSS 0.262563f
C25131 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n46 VSS 0.262563f
C25132 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n47 VSS 0.262563f
C25133 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n48 VSS 0.262563f
C25134 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n49 VSS 0.262563f
C25135 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n50 VSS 0.262563f
C25136 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n51 VSS 0.197637f
C25137 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n52 VSS 0.262563f
C25138 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n53 VSS 0.153708f
C25139 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n54 VSS 0.262563f
C25140 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n55 VSS 0.262563f
C25141 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n56 VSS 0.262563f
C25142 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n57 VSS 0.262563f
C25143 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n58 VSS 0.262563f
C25144 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n59 VSS 0.262563f
C25145 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n60 VSS 0.504461f
C25146 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n61 VSS 0.241493f
C25147 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n62 VSS 3.64116f
C25148 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n63 VSS 0.43882f
C25149 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n64 VSS 0.262563f
C25150 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n65 VSS 0.219739f
C25151 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n66 VSS 0.262563f
C25152 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n67 VSS 0.262563f
C25153 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n68 VSS 0.262563f
C25154 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n69 VSS 0.262563f
C25155 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n70 VSS 0.262563f
C25156 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n71 VSS 0.262563f
C25157 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n72 VSS 0.262563f
C25158 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n73 VSS 0.197637f
C25159 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n74 VSS 0.262563f
C25160 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n75 VSS 0.153708f
C25161 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n76 VSS 0.262563f
C25162 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n77 VSS 0.262563f
C25163 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n78 VSS 0.262563f
C25164 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n79 VSS 0.262563f
C25165 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n80 VSS 0.262563f
C25166 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n81 VSS 0.262563f
C25167 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n82 VSS 0.262563f
C25168 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n83 VSS 0.241493f
C25169 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n84 VSS 2.13477f
C25170 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n85 VSS 3.62978f
C25171 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n86 VSS 3.77257f
C25172 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n87 VSS 0.43882f
C25173 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n88 VSS 3.7904f
C25174 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n89 VSS 3.77257f
C25175 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.t14 VSS 0.323661f
C25176 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n90 VSS 0.349909f
C25177 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n91 VSS 0.712344f
C25178 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.t10 VSS 0.323661f
C25179 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n92 VSS 0.349909f
C25180 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.t12 VSS 0.323661f
C25181 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n93 VSS 0.254768f
C25182 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.t16 VSS 0.323661f
C25183 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n94 VSS 0.349909f
C25184 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n95 VSS 0.349909f
C25185 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.t15 VSS 0.323661f
C25186 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n96 VSS 0.349909f
C25187 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.t8 VSS 0.323661f
C25188 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n97 VSS 0.349909f
C25189 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.t9 VSS 0.323661f
C25190 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n98 VSS 0.349909f
C25191 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.t7 VSS 0.323661f
C25192 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n99 VSS 0.349909f
C25193 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.t13 VSS 0.323661f
C25194 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.t5 VSS 0.882832f
C25195 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.t11 VSS 0.416732f
C25196 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.t6 VSS 0.079012f
C25197 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.t4 VSS 0.079012f
C25198 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n100 VSS 0.260778f
C25199 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.t1 VSS 0.242287f
C25200 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n101 VSS 0.127545f
C25201 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n102 VSS 0.220681f
C25202 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.t3 VSS 0.079012f
C25203 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n103 VSS 0.068218f
C25204 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.t51 VSS 2.15277f
C25205 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.t72 VSS 2.15277f
C25206 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.t57 VSS 2.15277f
C25207 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.t79 VSS 2.15277f
C25208 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.t67 VSS 2.15277f
C25209 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.t93 VSS 2.15277f
C25210 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.t52 VSS 2.15277f
C25211 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.t36 VSS 2.15277f
C25212 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.t62 VSS 2.15277f
C25213 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n104 VSS 1.17871f
C25214 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n105 VSS 1.21282f
C25215 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n106 VSS 1.21282f
C25216 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n107 VSS 1.21282f
C25217 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n108 VSS 1.21282f
C25218 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n109 VSS 1.21282f
C25219 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n110 VSS 1.21282f
C25220 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n111 VSS 1.21282f
C25221 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n112 VSS 2.35467f
C25222 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.t47 VSS 2.23656f
C25223 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n113 VSS 2.35467f
C25224 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n114 VSS 1.21282f
C25225 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n115 VSS 1.21282f
C25226 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n116 VSS 1.21282f
C25227 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n117 VSS 1.21282f
C25228 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n118 VSS 1.21282f
C25229 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n119 VSS 1.21282f
C25230 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n120 VSS 1.21282f
C25231 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n121 VSS 1.17871f
C25232 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.t86 VSS 2.15277f
C25233 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.t40 VSS 2.15277f
C25234 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.t78 VSS 2.15277f
C25235 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.t96 VSS 2.15277f
C25236 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.t65 VSS 2.15277f
C25237 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.t29 VSS 2.15277f
C25238 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.t61 VSS 2.15277f
C25239 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.t24 VSS 2.15277f
C25240 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.t50 VSS 2.15277f
C25241 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n122 VSS 1.17871f
C25242 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n123 VSS 1.21282f
C25243 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n124 VSS 1.21282f
C25244 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n125 VSS 1.21282f
C25245 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n126 VSS 1.21282f
C25246 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n127 VSS 1.21282f
C25247 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n128 VSS 1.21282f
C25248 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n129 VSS 1.21282f
C25249 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n130 VSS 2.35467f
C25250 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.t90 VSS 2.23656f
C25251 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n131 VSS 2.35467f
C25252 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n132 VSS 1.21282f
C25253 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n133 VSS 1.21282f
C25254 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n134 VSS 1.21282f
C25255 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n135 VSS 1.21282f
C25256 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n136 VSS 1.21282f
C25257 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n137 VSS 1.21282f
C25258 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n138 VSS 1.21282f
C25259 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n139 VSS 1.17871f
C25260 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n140 VSS 0.559014f
C25261 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n141 VSS 0.476663f
C25262 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.t95 VSS 2.15277f
C25263 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.t55 VSS 2.15277f
C25264 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.t22 VSS 2.15277f
C25265 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.t60 VSS 2.15277f
C25266 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.t68 VSS 2.15277f
C25267 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.t35 VSS 2.15277f
C25268 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.t76 VSS 2.15277f
C25269 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.t44 VSS 2.15277f
C25270 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.t87 VSS 2.15277f
C25271 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n142 VSS 1.17871f
C25272 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n143 VSS 1.21282f
C25273 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n144 VSS 1.21282f
C25274 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n145 VSS 1.21282f
C25275 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n146 VSS 1.21282f
C25276 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n147 VSS 1.21282f
C25277 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n148 VSS 1.21282f
C25278 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n149 VSS 1.21282f
C25279 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n150 VSS 2.35467f
C25280 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.t30 VSS 2.23656f
C25281 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n151 VSS 2.35467f
C25282 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n152 VSS 1.21282f
C25283 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n153 VSS 1.21282f
C25284 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n154 VSS 1.21282f
C25285 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n155 VSS 1.21282f
C25286 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n156 VSS 1.21282f
C25287 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n157 VSS 1.21282f
C25288 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n158 VSS 1.21282f
C25289 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n159 VSS 1.17871f
C25290 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.t45 VSS 2.15277f
C25291 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.t84 VSS 2.15277f
C25292 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.t59 VSS 2.15277f
C25293 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.t74 VSS 2.15277f
C25294 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.t49 VSS 2.15277f
C25295 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.t64 VSS 2.15277f
C25296 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.t27 VSS 2.15277f
C25297 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.t81 VSS 2.15277f
C25298 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.t19 VSS 2.15277f
C25299 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n160 VSS 1.17871f
C25300 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n161 VSS 1.21282f
C25301 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n162 VSS 1.21282f
C25302 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n163 VSS 1.21282f
C25303 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n164 VSS 1.21282f
C25304 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n165 VSS 1.21282f
C25305 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n166 VSS 1.21282f
C25306 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n167 VSS 1.21282f
C25307 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n168 VSS 2.35467f
C25308 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.t69 VSS 2.23656f
C25309 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n169 VSS 2.35467f
C25310 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n170 VSS 1.21282f
C25311 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n171 VSS 1.21282f
C25312 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n172 VSS 1.21282f
C25313 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n173 VSS 1.21282f
C25314 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n174 VSS 1.21282f
C25315 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n175 VSS 1.21282f
C25316 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n176 VSS 1.21282f
C25317 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n177 VSS 1.17871f
C25318 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n178 VSS 0.068218f
C25319 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n179 VSS 0.173781f
C25320 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n180 VSS 0.068218f
C25321 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.t38 VSS 2.15277f
C25322 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.t77 VSS 2.15277f
C25323 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.t23 VSS 2.15277f
C25324 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.t91 VSS 2.15277f
C25325 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.t33 VSS 2.15277f
C25326 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.t17 VSS 2.15277f
C25327 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.t39 VSS 2.15277f
C25328 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.t85 VSS 2.15277f
C25329 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.t66 VSS 2.15277f
C25330 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n181 VSS 1.17871f
C25331 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n182 VSS 1.21282f
C25332 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n183 VSS 1.21282f
C25333 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n184 VSS 1.21282f
C25334 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n185 VSS 1.21282f
C25335 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n186 VSS 1.21282f
C25336 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n187 VSS 1.21282f
C25337 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n188 VSS 1.21282f
C25338 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n189 VSS 2.35467f
C25339 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.t92 VSS 2.23656f
C25340 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n190 VSS 2.35467f
C25341 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n191 VSS 1.21282f
C25342 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n192 VSS 1.21282f
C25343 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n193 VSS 1.21282f
C25344 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n194 VSS 1.21282f
C25345 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n195 VSS 1.21282f
C25346 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n196 VSS 1.21282f
C25347 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n197 VSS 1.21282f
C25348 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n198 VSS 1.17871f
C25349 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.t71 VSS 2.15277f
C25350 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.t28 VSS 2.15277f
C25351 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.t43 VSS 2.15277f
C25352 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.t21 VSS 2.15277f
C25353 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.t58 VSS 2.15277f
C25354 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.t89 VSS 2.15277f
C25355 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.t48 VSS 2.15277f
C25356 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.t83 VSS 2.15277f
C25357 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.t42 VSS 2.15277f
C25358 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n199 VSS 1.17871f
C25359 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n200 VSS 1.21282f
C25360 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n201 VSS 1.21282f
C25361 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n202 VSS 1.21282f
C25362 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n203 VSS 1.21282f
C25363 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n204 VSS 1.21282f
C25364 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n205 VSS 1.21282f
C25365 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n206 VSS 1.21282f
C25366 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n207 VSS 2.35467f
C25367 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.t75 VSS 2.23656f
C25368 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n208 VSS 2.35467f
C25369 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n209 VSS 1.21282f
C25370 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n210 VSS 1.21282f
C25371 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n211 VSS 1.21282f
C25372 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n212 VSS 1.21282f
C25373 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n213 VSS 1.21282f
C25374 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n214 VSS 1.21282f
C25375 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n215 VSS 1.21282f
C25376 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n216 VSS 1.17871f
C25377 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n217 VSS 0.559014f
C25378 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n218 VSS 1.17871f
C25379 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.t34 VSS 2.15277f
C25380 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.t88 VSS 2.15277f
C25381 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.t26 VSS 2.15277f
C25382 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.t80 VSS 2.15277f
C25383 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.t18 VSS 2.15277f
C25384 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.t56 VSS 2.15277f
C25385 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.t31 VSS 2.15277f
C25386 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.t46 VSS 2.15277f
C25387 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.t25 VSS 2.15277f
C25388 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.t73 VSS 2.15277f
C25389 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.t41 VSS 2.15277f
C25390 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.t82 VSS 2.15277f
C25391 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.t53 VSS 2.15277f
C25392 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.t94 VSS 2.15277f
C25393 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.t54 VSS 2.15277f
C25394 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.t20 VSS 2.15277f
C25395 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.t63 VSS 2.15277f
C25396 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.t32 VSS 2.15277f
C25397 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n219 VSS 1.21282f
C25398 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n220 VSS 1.21282f
C25399 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n221 VSS 1.21282f
C25400 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n222 VSS 1.21282f
C25401 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n223 VSS 1.21282f
C25402 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n224 VSS 1.21282f
C25403 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n225 VSS 1.21282f
C25404 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n226 VSS 2.35467f
C25405 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.t70 VSS 2.23656f
C25406 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n227 VSS 2.35467f
C25407 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n228 VSS 1.21282f
C25408 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n229 VSS 1.21282f
C25409 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n230 VSS 1.21282f
C25410 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n231 VSS 1.21282f
C25411 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n232 VSS 1.21282f
C25412 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n233 VSS 1.21282f
C25413 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n234 VSS 1.21282f
C25414 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n235 VSS 1.17871f
C25415 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n236 VSS 0.068218f
C25416 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n237 VSS 1.17871f
C25417 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n238 VSS 1.21282f
C25418 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n239 VSS 1.21282f
C25419 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n240 VSS 1.21282f
C25420 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n241 VSS 1.21282f
C25421 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n242 VSS 1.21282f
C25422 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n243 VSS 1.21282f
C25423 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n244 VSS 1.21282f
C25424 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n245 VSS 2.35467f
C25425 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.t37 VSS 2.23656f
C25426 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n246 VSS 2.35467f
C25427 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n247 VSS 1.21282f
C25428 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n248 VSS 1.21282f
C25429 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n249 VSS 1.21282f
C25430 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n250 VSS 1.21282f
C25431 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n251 VSS 1.21282f
C25432 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n252 VSS 1.21282f
C25433 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n253 VSS 1.21282f
C25434 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n254 VSS 1.17871f
C25435 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n255 VSS 0.173781f
C25436 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n256 VSS 0.173781f
C25437 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n257 VSS 4.96058f
C25438 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.t2 VSS 0.079012f
C25439 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n258 VSS 0.158024f
C25440 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n259 VSS 0.239043f
C25441 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n260 VSS 0.518305f
C25442 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.t0 VSS 0.242287f
C25443 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_0.D.n261 VSS 0.127545f
C25444 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_1.D.n0 VSS 0.229397f
C25445 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_1.D.n1 VSS 2.54242f
C25446 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_1.D.t0 VSS 0.750086f
C25447 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_1.D.t2 VSS 2.78176f
C25448 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_1.D.t3 VSS 1.93087f
C25449 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_1.D.t1 VSS 0.747757f
C25450 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_1.D.t24 VSS 0.691125f
C25451 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_1.D.t32 VSS 0.626919f
C25452 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_1.D.n2 VSS 0.628841f
C25453 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_1.D.t22 VSS 0.626919f
C25454 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_1.D.n3 VSS 0.346524f
C25455 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_1.D.t11 VSS 0.691125f
C25456 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_1.D.t10 VSS 0.626919f
C25457 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_1.D.n4 VSS 0.628841f
C25458 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_1.D.t23 VSS 0.626919f
C25459 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_1.D.n5 VSS 0.346524f
C25460 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_1.D.t7 VSS 0.691125f
C25461 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_1.D.t21 VSS 0.626919f
C25462 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_1.D.n6 VSS 0.628841f
C25463 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_1.D.t31 VSS 0.626919f
C25464 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_1.D.n7 VSS 0.358436f
C25465 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_1.D.t9 VSS 0.626919f
C25466 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_1.D.n8 VSS 0.358436f
C25467 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_1.D.t20 VSS 0.626919f
C25468 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_1.D.n9 VSS 0.358436f
C25469 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_1.D.t27 VSS 0.626919f
C25470 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_1.D.n10 VSS 0.358436f
C25471 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_1.D.t4 VSS 0.626919f
C25472 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_1.D.n11 VSS 0.358436f
C25473 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_1.D.t12 VSS 0.626919f
C25474 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_1.D.n12 VSS 0.358436f
C25475 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_1.D.t25 VSS 0.626919f
C25476 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_1.D.n13 VSS 0.358436f
C25477 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_1.D.t29 VSS 0.626919f
C25478 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_1.D.n14 VSS 0.358436f
C25479 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_1.D.t14 VSS 0.626919f
C25480 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_1.D.n15 VSS 0.358436f
C25481 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_1.D.t15 VSS 0.626919f
C25482 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_1.D.n16 VSS 0.346524f
C25483 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_1.D.t19 VSS 0.691125f
C25484 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_1.D.t18 VSS 0.626919f
C25485 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_1.D.n17 VSS 0.628841f
C25486 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_1.D.t28 VSS 0.626919f
C25487 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_1.D.n18 VSS 0.358436f
C25488 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_1.D.t16 VSS 0.626919f
C25489 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_1.D.n19 VSS 0.358436f
C25490 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_1.D.t8 VSS 0.626919f
C25491 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_1.D.n20 VSS 0.358436f
C25492 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_1.D.t30 VSS 0.626919f
C25493 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_1.D.n21 VSS 0.358436f
C25494 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_1.D.t26 VSS 0.626919f
C25495 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_1.D.n22 VSS 0.358436f
C25496 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_1.D.t6 VSS 0.626919f
C25497 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_1.D.n23 VSS 0.358436f
C25498 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_1.D.t5 VSS 0.626919f
C25499 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_1.D.n24 VSS 0.358436f
C25500 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_1.D.t17 VSS 0.626919f
C25501 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_1.D.n25 VSS 0.358436f
C25502 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_1.D.t13 VSS 0.626919f
C25503 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_1.D.n26 VSS 0.358436f
C25504 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_1.D.t33 VSS 0.626919f
C25505 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/nmos_6p0_CDNS_406619531458_1.D.n27 VSS 0.346524f
.ends

