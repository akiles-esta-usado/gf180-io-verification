* NGSPICE file created from gf180mcu_fd_io__dvdd_flat.ext - technology: gf180mcuD

.subckt gf180mcu_fd_io__dvdd_flat VSS DVSS DVDD
X0 DVDD GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/pmos_6p0_CDNS_406619531456_0.D GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/pmos_6p0_CDNS_406619531455_0.D DVDD pfet_06v0 ad=1.3p pd=5.52u as=1.3p ps=5.52u w=5u l=0.7u
X1 DVDD GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/pmos_6p0_CDNS_406619531455_0.D DVSS DVSS nfet_06v0 ad=12.999999p pd=50.52u as=12.999999p ps=50.52u w=50u l=0.7u
X2 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/pmos_6p0_CDNS_406619531455_0.D GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/pmos_6p0_CDNS_406619531456_0.D DVDD DVDD pfet_06v0 ad=1.3p pd=5.52u as=1.3p ps=5.52u w=5u l=0.7u
X3 DVDD GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/pmos_6p0_CDNS_406619531455_0.D DVSS DVSS nfet_06v0 ad=12.999999p pd=50.52u as=12.999999p ps=50.52u w=50u l=0.7u
X4 DVDD GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/pmos_6p0_CDNS_406619531455_0.D DVSS DVSS nfet_06v0 ad=12.999999p pd=50.52u as=12.999999p ps=50.52u w=50u l=0.7u
X5 DVDD GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/pmos_6p0_CDNS_406619531456_0.D GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/pmos_6p0_CDNS_406619531455_0.D DVDD pfet_06v0 ad=1.3p pd=5.52u as=1.3p ps=5.52u w=5u l=0.7u
X6 DVDD GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/pmos_6p0_CDNS_406619531456_0.D GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/pmos_6p0_CDNS_406619531455_0.D DVDD pfet_06v0 ad=2.2p pd=10.879999u as=1.3p ps=5.52u w=5u l=0.7u
X7 DVSS GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/pmos_6p0_CDNS_406619531455_0.D DVDD DVSS nfet_06v0 ad=12.999999p pd=50.52u as=12.999999p ps=50.52u w=50u l=0.7u
X8 DVSS GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/pmos_6p0_CDNS_406619531455_0.D DVDD DVSS nfet_06v0 ad=12.999999p pd=50.52u as=12.999999p ps=50.52u w=50u l=0.7u
X9 DVSS GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/pmos_6p0_CDNS_406619531455_0.D DVDD DVSS nfet_06v0 ad=12.999999p pd=50.52u as=12.999999p ps=50.52u w=50u l=0.7u
X10 DVSS GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/pmos_6p0_CDNS_406619531455_0.D DVDD DVSS nfet_06v0 ad=12.999999p pd=50.52u as=12.999999p ps=50.52u w=50u l=0.7u
X11 DVSS GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/pmos_6p0_CDNS_406619531455_0.D DVDD DVSS nfet_06v0 ad=12.999999p pd=50.52u as=12.999999p ps=50.52u w=50u l=0.7u
X12 DVDD DVSS cap_nmos_06v0 c_width=15u c_length=15u
X13 DVDD GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/pmos_6p0_CDNS_406619531455_0.D DVSS DVSS nfet_06v0 ad=12.999999p pd=50.52u as=12.999999p ps=50.52u w=50u l=0.7u
X14 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/pmos_6p0_CDNS_406619531456_0.D GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/pmos_6p0_CDNS_406619531452_0.D DVDD DVDD pfet_06v0 ad=2.2p pd=10.879999u as=1.3p ps=5.52u w=5u l=0.7u
X15 DVDD GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/pmos_6p0_CDNS_406619531455_0.D DVSS DVSS nfet_06v0 ad=12.999999p pd=50.52u as=12.999999p ps=50.52u w=50u l=0.7u
X16 DVDD GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/pmos_6p0_CDNS_406619531455_0.D DVSS DVSS nfet_06v0 ad=12.999999p pd=50.52u as=12.999999p ps=50.52u w=50u l=0.7u
X17 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/pmos_6p0_CDNS_406619531455_0.D GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/pmos_6p0_CDNS_406619531456_0.D DVDD DVDD pfet_06v0 ad=1.3p pd=5.52u as=1.3p ps=5.52u w=5u l=0.7u
X18 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/pmos_6p0_CDNS_406619531455_0.D GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/pmos_6p0_CDNS_406619531456_0.D DVDD DVDD pfet_06v0 ad=1.3p pd=5.52u as=1.3p ps=5.52u w=5u l=0.7u
X19 DVSS GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/pmos_6p0_CDNS_406619531455_0.D DVDD DVSS nfet_06v0 ad=12.999999p pd=50.52u as=12.999999p ps=50.52u w=50u l=0.7u
X20 DVSS GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/pmos_6p0_CDNS_406619531455_0.D DVDD DVSS nfet_06v0 ad=12.999999p pd=50.52u as=12.999999p ps=50.52u w=50u l=0.7u
X21 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/comp018green_esd_rc_v5p0_0.ppolyf_u_CDNS_406619531453_1.MINUS GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/comp018green_esd_rc_v5p0_0.ppolyf_u_CDNS_406619531453_0.PLUS DVDD ppolyf_u r_width=0.8u r_length=63.854996u
X22 DVDD GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/pmos_6p0_CDNS_406619531455_0.D DVSS DVSS nfet_06v0 ad=21.999998p pd=0.10088m as=12.999999p ps=50.52u w=50u l=0.7u
X23 DVDD GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/comp018green_esd_rc_v5p0_0.VRC GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/pmos_6p0_CDNS_406619531452_0.D DVDD pfet_06v0 ad=1.3p pd=5.52u as=1.3p ps=5.52u w=5u l=0.7u
X24 DVDD GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/pmos_6p0_CDNS_406619531455_0.D DVSS DVSS nfet_06v0 ad=12.999999p pd=50.52u as=12.999999p ps=50.52u w=50u l=0.7u
D0 DVSS DVDD diode_nd2ps_06v0 pj=82u area=40p
X25 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/pmos_6p0_CDNS_406619531452_0.D GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/comp018green_esd_rc_v5p0_0.VRC DVDD DVDD pfet_06v0 ad=1.3p pd=5.52u as=1.3p ps=5.52u w=5u l=0.7u
X26 DVSS GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/pmos_6p0_CDNS_406619531455_0.D DVDD DVSS nfet_06v0 ad=12.999999p pd=50.52u as=12.999999p ps=50.52u w=50u l=0.7u
X27 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/comp018green_esd_rc_v5p0_0.ppolyf_u_CDNS_406619531453_5.MINUS GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/comp018green_esd_rc_v5p0_0.ppolyf_u_CDNS_406619531453_3.PLUS DVDD ppolyf_u r_width=0.8u r_length=63.854996u
X28 DVSS GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/pmos_6p0_CDNS_406619531455_0.D DVDD DVSS nfet_06v0 ad=12.999999p pd=50.52u as=12.999999p ps=50.52u w=50u l=0.7u
X29 DVDD DVSS cap_nmos_06v0 c_width=15u c_length=15u
X30 DVDD DVSS cap_nmos_06v0 c_width=15u c_length=15u
X31 DVSS GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/pmos_6p0_CDNS_406619531456_0.D GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/pmos_6p0_CDNS_406619531455_0.D DVSS nfet_06v0 ad=1.3p pd=5.52u as=1.3p ps=5.52u w=5u l=0.7u
X32 DVDD GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/pmos_6p0_CDNS_406619531455_0.D DVSS DVSS nfet_06v0 ad=12.999999p pd=50.52u as=12.999999p ps=50.52u w=50u l=0.7u
X33 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/pmos_6p0_CDNS_406619531455_0.D GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/pmos_6p0_CDNS_406619531456_0.D DVSS DVSS nfet_06v0 ad=1.3p pd=5.52u as=1.3p ps=5.52u w=5u l=0.7u
X34 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/comp018green_esd_rc_v5p0_0.ppolyf_u_CDNS_406619531453_2.MINUS GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/comp018green_esd_rc_v5p0_0.ppolyf_u_CDNS_406619531453_4.PLUS DVDD ppolyf_u r_width=0.8u r_length=63.854996u
X35 DVDD GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/pmos_6p0_CDNS_406619531455_0.D DVSS DVSS nfet_06v0 ad=12.999999p pd=50.52u as=12.999999p ps=50.52u w=50u l=0.7u
X36 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/pmos_6p0_CDNS_406619531455_0.D GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/pmos_6p0_CDNS_406619531456_0.D DVDD DVDD pfet_06v0 ad=1.3p pd=5.52u as=1.3p ps=5.52u w=5u l=0.7u
X37 DVDD GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/pmos_6p0_CDNS_406619531455_0.D DVSS DVSS nfet_06v0 ad=12.999999p pd=50.52u as=12.999999p ps=50.52u w=50u l=0.7u
X38 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/pmos_6p0_CDNS_406619531452_0.D GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/comp018green_esd_rc_v5p0_0.VRC DVSS DVSS nfet_06v0 ad=2.2p pd=10.879999u as=2.2p ps=10.879999u w=5u l=0.7u
X39 DVSS GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/pmos_6p0_CDNS_406619531455_0.D DVDD DVSS nfet_06v0 ad=12.999999p pd=50.52u as=21.999998p ps=0.10088m w=50u l=0.7u
X40 DVSS GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/pmos_6p0_CDNS_406619531455_0.D DVDD DVSS nfet_06v0 ad=12.999999p pd=50.52u as=12.999999p ps=50.52u w=50u l=0.7u
X41 DVSS GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/pmos_6p0_CDNS_406619531455_0.D DVDD DVSS nfet_06v0 ad=12.999999p pd=50.52u as=12.999999p ps=50.52u w=50u l=0.7u
X42 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/pmos_6p0_CDNS_406619531456_0.D GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/pmos_6p0_CDNS_406619531452_0.D DVSS DVSS nfet_06v0 ad=1.3p pd=5.52u as=2.2p ps=10.879999u w=5u l=0.7u
X43 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/pmos_6p0_CDNS_406619531455_0.D GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/pmos_6p0_CDNS_406619531456_0.D DVDD DVDD pfet_06v0 ad=1.3p pd=5.52u as=1.3p ps=5.52u w=5u l=0.7u
X44 DVSS GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/pmos_6p0_CDNS_406619531455_0.D DVDD DVSS nfet_06v0 ad=12.999999p pd=50.52u as=12.999999p ps=50.52u w=50u l=0.7u
X45 DVSS GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/pmos_6p0_CDNS_406619531452_0.D GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/pmos_6p0_CDNS_406619531456_0.D DVSS nfet_06v0 ad=1.3p pd=5.52u as=1.3p ps=5.52u w=5u l=0.7u
X46 DVDD GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/pmos_6p0_CDNS_406619531455_0.D DVSS DVSS nfet_06v0 ad=12.999999p pd=50.52u as=12.999999p ps=50.52u w=50u l=0.7u
X47 DVDD GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/pmos_6p0_CDNS_406619531456_0.D GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/pmos_6p0_CDNS_406619531455_0.D DVDD pfet_06v0 ad=1.3p pd=5.52u as=1.3p ps=5.52u w=5u l=0.7u
X48 DVDD GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/pmos_6p0_CDNS_406619531455_0.D DVSS DVSS nfet_06v0 ad=12.999999p pd=50.52u as=12.999999p ps=50.52u w=50u l=0.7u
X49 DVDD GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/pmos_6p0_CDNS_406619531455_0.D DVSS DVSS nfet_06v0 ad=12.999999p pd=50.52u as=12.999999p ps=50.52u w=50u l=0.7u
X50 DVDD GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/pmos_6p0_CDNS_406619531455_0.D DVSS DVSS nfet_06v0 ad=12.999999p pd=50.52u as=12.999999p ps=50.52u w=50u l=0.7u
X51 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/pmos_6p0_CDNS_406619531455_0.D GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/pmos_6p0_CDNS_406619531456_0.D DVDD DVDD pfet_06v0 ad=1.3p pd=5.52u as=1.3p ps=5.52u w=5u l=0.7u
X52 DVDD GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/pmos_6p0_CDNS_406619531455_0.D DVSS DVSS nfet_06v0 ad=12.999999p pd=50.52u as=12.999999p ps=50.52u w=50u l=0.7u
X53 DVDD GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/pmos_6p0_CDNS_406619531456_0.D GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/pmos_6p0_CDNS_406619531455_0.D DVDD pfet_06v0 ad=1.3p pd=5.52u as=1.3p ps=5.52u w=5u l=0.7u
X54 DVSS GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/pmos_6p0_CDNS_406619531455_0.D DVDD DVSS nfet_06v0 ad=12.999999p pd=50.52u as=12.999999p ps=50.52u w=50u l=0.7u
X55 DVDD GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/pmos_6p0_CDNS_406619531455_0.D DVSS DVSS nfet_06v0 ad=21.999998p pd=0.10088m as=12.999999p ps=50.52u w=50u l=0.7u
X56 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/comp018green_esd_rc_v5p0_0.VRC DVSS cap_nmos_06v0 c_width=25u c_length=10u
X57 DVDD GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/pmos_6p0_CDNS_406619531455_0.D DVSS DVSS nfet_06v0 ad=12.999999p pd=50.52u as=12.999999p ps=50.52u w=50u l=0.7u
X58 DVDD GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/pmos_6p0_CDNS_406619531456_0.D GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/pmos_6p0_CDNS_406619531455_0.D DVDD pfet_06v0 ad=1.3p pd=5.52u as=1.3p ps=5.52u w=5u l=0.7u
X59 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/comp018green_esd_rc_v5p0_0.VRC GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/comp018green_esd_rc_v5p0_0.ppolyf_u_CDNS_406619531453_0.PLUS DVDD ppolyf_u r_width=0.8u r_length=63.854996u
X60 DVDD GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/pmos_6p0_CDNS_406619531455_0.D DVSS DVSS nfet_06v0 ad=12.999999p pd=50.52u as=12.999999p ps=50.52u w=50u l=0.7u
X61 DVDD GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/pmos_6p0_CDNS_406619531456_0.D GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/pmos_6p0_CDNS_406619531455_0.D DVDD pfet_06v0 ad=1.3p pd=5.52u as=1.3p ps=5.52u w=5u l=0.7u
X62 DVDD GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/pmos_6p0_CDNS_406619531455_0.D DVSS DVSS nfet_06v0 ad=12.999999p pd=50.52u as=12.999999p ps=50.52u w=50u l=0.7u
X63 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/comp018green_esd_rc_v5p0_0.VRC DVSS cap_nmos_06v0 c_width=25u c_length=10u
X64 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/pmos_6p0_CDNS_406619531455_0.D GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/pmos_6p0_CDNS_406619531456_0.D DVDD DVDD pfet_06v0 ad=1.3p pd=5.52u as=2.2p ps=10.879999u w=5u l=0.7u
X65 DVSS GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/pmos_6p0_CDNS_406619531455_0.D DVDD DVSS nfet_06v0 ad=12.999999p pd=50.52u as=12.999999p ps=50.52u w=50u l=0.7u
X66 DVSS GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/pmos_6p0_CDNS_406619531455_0.D DVDD DVSS nfet_06v0 ad=12.999999p pd=50.52u as=12.999999p ps=50.52u w=50u l=0.7u
X67 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/comp018green_esd_rc_v5p0_0.VRC DVSS cap_nmos_06v0 c_width=25u c_length=10u
X68 DVDD GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/pmos_6p0_CDNS_406619531456_0.D GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/pmos_6p0_CDNS_406619531455_0.D DVDD pfet_06v0 ad=1.3p pd=5.52u as=1.3p ps=5.52u w=5u l=0.7u
X69 DVDD GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/pmos_6p0_CDNS_406619531455_0.D DVSS DVSS nfet_06v0 ad=12.999999p pd=50.52u as=12.999999p ps=50.52u w=50u l=0.7u
X70 DVDD GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/pmos_6p0_CDNS_406619531455_0.D DVSS DVSS nfet_06v0 ad=12.999999p pd=50.52u as=12.999999p ps=50.52u w=50u l=0.7u
X71 DVDD GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/pmos_6p0_CDNS_406619531455_0.D DVSS DVSS nfet_06v0 ad=12.999999p pd=50.52u as=12.999999p ps=50.52u w=50u l=0.7u
X72 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/pmos_6p0_CDNS_406619531455_0.D GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/pmos_6p0_CDNS_406619531456_0.D DVDD DVDD pfet_06v0 ad=1.3p pd=5.52u as=1.3p ps=5.52u w=5u l=0.7u
X73 DVSS GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/pmos_6p0_CDNS_406619531456_0.D GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/pmos_6p0_CDNS_406619531455_0.D DVSS nfet_06v0 ad=1.3p pd=5.52u as=1.3p ps=5.52u w=5u l=0.7u
X74 DVSS GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/pmos_6p0_CDNS_406619531455_0.D DVDD DVSS nfet_06v0 ad=12.999999p pd=50.52u as=12.999999p ps=50.52u w=50u l=0.7u
X75 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/pmos_6p0_CDNS_406619531455_0.D GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/pmos_6p0_CDNS_406619531456_0.D DVSS DVSS nfet_06v0 ad=1.3p pd=5.52u as=1.3p ps=5.52u w=5u l=0.7u
X76 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/comp018green_esd_rc_v5p0_0.ppolyf_u_CDNS_406619531453_3.MINUS GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/comp018green_esd_rc_v5p0_0.ppolyf_u_CDNS_406619531453_3.PLUS DVDD ppolyf_u r_width=0.8u r_length=63.854996u
X77 DVSS GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/pmos_6p0_CDNS_406619531455_0.D DVDD DVSS nfet_06v0 ad=12.999999p pd=50.52u as=12.999999p ps=50.52u w=50u l=0.7u
X78 DVDD GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/pmos_6p0_CDNS_406619531455_0.D DVSS DVSS nfet_06v0 ad=12.999999p pd=50.52u as=12.999999p ps=50.52u w=50u l=0.7u
X79 DVSS GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/pmos_6p0_CDNS_406619531456_0.D GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/pmos_6p0_CDNS_406619531455_0.D DVSS nfet_06v0 ad=2.2p pd=10.879999u as=1.3p ps=5.52u w=5u l=0.7u
X80 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/comp018green_esd_rc_v5p0_0.ppolyf_u_CDNS_406619531453_4.MINUS GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/comp018green_esd_rc_v5p0_0.ppolyf_u_CDNS_406619531453_4.PLUS DVDD ppolyf_u r_width=0.8u r_length=63.854996u
X81 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/comp018green_esd_rc_v5p0_0.VRC DVSS cap_nmos_06v0 c_width=25u c_length=10u
X82 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/comp018green_esd_rc_v5p0_0.VRC DVSS cap_nmos_06v0 c_width=25u c_length=10u
X83 DVDD GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/pmos_6p0_CDNS_406619531452_0.D GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/pmos_6p0_CDNS_406619531456_0.D DVDD pfet_06v0 ad=1.3p pd=5.52u as=1.3p ps=5.52u w=5u l=0.7u
X84 DVDD GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/pmos_6p0_CDNS_406619531455_0.D DVSS DVSS nfet_06v0 ad=12.999999p pd=50.52u as=12.999999p ps=50.52u w=50u l=0.7u
X85 DVDD GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/pmos_6p0_CDNS_406619531455_0.D DVSS DVSS nfet_06v0 ad=12.999999p pd=50.52u as=12.999999p ps=50.52u w=50u l=0.7u
X86 DVDD GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/pmos_6p0_CDNS_406619531455_0.D DVSS DVSS nfet_06v0 ad=12.999999p pd=50.52u as=12.999999p ps=50.52u w=50u l=0.7u
X87 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/comp018green_esd_rc_v5p0_0.ppolyf_u_CDNS_406619531453_4.MINUS GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/comp018green_esd_rc_v5p0_0.ppolyf_u_CDNS_406619531453_5.PLUS DVDD ppolyf_u r_width=0.8u r_length=63.854996u
X88 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/pmos_6p0_CDNS_406619531456_0.D GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/pmos_6p0_CDNS_406619531452_0.D DVDD DVDD pfet_06v0 ad=1.3p pd=5.52u as=1.3p ps=5.52u w=5u l=0.7u
X89 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/pmos_6p0_CDNS_406619531456_0.D GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/pmos_6p0_CDNS_406619531452_0.D DVSS DVSS nfet_06v0 ad=1.3p pd=5.52u as=1.3p ps=5.52u w=5u l=0.7u
X90 DVSS GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/pmos_6p0_CDNS_406619531455_0.D DVDD DVSS nfet_06v0 ad=12.999999p pd=50.52u as=12.999999p ps=50.52u w=50u l=0.7u
X91 DVSS GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/pmos_6p0_CDNS_406619531452_0.D GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/pmos_6p0_CDNS_406619531456_0.D DVSS nfet_06v0 ad=1.3p pd=5.52u as=1.3p ps=5.52u w=5u l=0.7u
X92 DVDD GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/pmos_6p0_CDNS_406619531456_0.D GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/pmos_6p0_CDNS_406619531455_0.D DVDD pfet_06v0 ad=1.3p pd=5.52u as=1.3p ps=5.52u w=5u l=0.7u
X93 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/comp018green_esd_rc_v5p0_0.VRC DVSS cap_nmos_06v0 c_width=25u c_length=10u
X94 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/comp018green_esd_rc_v5p0_0.VRC DVSS cap_nmos_06v0 c_width=25u c_length=10u
X95 DVDD GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/pmos_6p0_CDNS_406619531455_0.D DVSS DVSS nfet_06v0 ad=12.999999p pd=50.52u as=12.999999p ps=50.52u w=50u l=0.7u
X96 DVSS GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/pmos_6p0_CDNS_406619531455_0.D DVDD DVSS nfet_06v0 ad=12.999999p pd=50.52u as=12.999999p ps=50.52u w=50u l=0.7u
X97 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/pmos_6p0_CDNS_406619531455_0.D GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/pmos_6p0_CDNS_406619531456_0.D DVDD DVDD pfet_06v0 ad=1.3p pd=5.52u as=1.3p ps=5.52u w=5u l=0.7u
X98 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/pmos_6p0_CDNS_406619531455_0.D GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/pmos_6p0_CDNS_406619531456_0.D DVDD DVDD pfet_06v0 ad=1.3p pd=5.52u as=1.3p ps=5.52u w=5u l=0.7u
X99 DVDD GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/pmos_6p0_CDNS_406619531455_0.D DVSS DVSS nfet_06v0 ad=12.999999p pd=50.52u as=12.999999p ps=50.52u w=50u l=0.7u
X100 DVSS GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/pmos_6p0_CDNS_406619531455_0.D DVDD DVSS nfet_06v0 ad=12.999999p pd=50.52u as=12.999999p ps=50.52u w=50u l=0.7u
X101 DVSS GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/pmos_6p0_CDNS_406619531455_0.D DVDD DVSS nfet_06v0 ad=12.999999p pd=50.52u as=12.999999p ps=50.52u w=50u l=0.7u
X102 DVDD GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/comp018green_esd_rc_v5p0_0.ppolyf_u_CDNS_406619531453_2.PLUS DVDD ppolyf_u r_width=0.8u r_length=63.854996u
X103 DVSS GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/pmos_6p0_CDNS_406619531455_0.D DVDD DVSS nfet_06v0 ad=12.999999p pd=50.52u as=12.999999p ps=50.52u w=50u l=0.7u
X104 DVSS GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/pmos_6p0_CDNS_406619531455_0.D DVDD DVSS nfet_06v0 ad=12.999999p pd=50.52u as=21.999998p ps=0.10088m w=50u l=0.7u
X105 DVDD GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/pmos_6p0_CDNS_406619531455_0.D DVSS DVSS nfet_06v0 ad=21.999998p pd=0.10088m as=12.999999p ps=50.52u w=50u l=0.7u
X106 DVDD GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/pmos_6p0_CDNS_406619531455_0.D DVSS DVSS nfet_06v0 ad=12.999999p pd=50.52u as=12.999999p ps=50.52u w=50u l=0.7u
D1 DVSS DVDD diode_nd2ps_06v0 pj=82u area=40p
X107 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/comp018green_esd_rc_v5p0_0.VRC DVSS cap_nmos_06v0 c_width=25u c_length=10u
X108 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/pmos_6p0_CDNS_406619531455_0.D GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/pmos_6p0_CDNS_406619531456_0.D DVDD DVDD pfet_06v0 ad=1.3p pd=5.52u as=1.3p ps=5.52u w=5u l=0.7u
X109 DVDD GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/pmos_6p0_CDNS_406619531455_0.D DVSS DVSS nfet_06v0 ad=12.999999p pd=50.52u as=12.999999p ps=50.52u w=50u l=0.7u
X110 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/pmos_6p0_CDNS_406619531455_0.D GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/pmos_6p0_CDNS_406619531456_0.D DVDD DVDD pfet_06v0 ad=1.3p pd=5.52u as=1.3p ps=5.52u w=5u l=0.7u
X111 DVSS GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/pmos_6p0_CDNS_406619531455_0.D DVDD DVSS nfet_06v0 ad=12.999999p pd=50.52u as=12.999999p ps=50.52u w=50u l=0.7u
X112 DVSS GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/pmos_6p0_CDNS_406619531455_0.D DVDD DVSS nfet_06v0 ad=12.999999p pd=50.52u as=12.999999p ps=50.52u w=50u l=0.7u
D2 DVSS DVDD diode_nd2ps_06v0 pj=82u area=40p
X113 DVDD GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/pmos_6p0_CDNS_406619531456_0.D GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/pmos_6p0_CDNS_406619531455_0.D DVDD pfet_06v0 ad=1.3p pd=5.52u as=1.3p ps=5.52u w=5u l=0.7u
X114 DVSS GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/pmos_6p0_CDNS_406619531455_0.D DVDD DVSS nfet_06v0 ad=12.999999p pd=50.52u as=21.999998p ps=0.10088m w=50u l=0.7u
X115 DVSS GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/pmos_6p0_CDNS_406619531455_0.D DVDD DVSS nfet_06v0 ad=12.999999p pd=50.52u as=12.999999p ps=50.52u w=50u l=0.7u
X116 DVDD GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/pmos_6p0_CDNS_406619531456_0.D GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/pmos_6p0_CDNS_406619531455_0.D DVDD pfet_06v0 ad=1.3p pd=5.52u as=1.3p ps=5.52u w=5u l=0.7u
X117 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/comp018green_esd_rc_v5p0_0.ppolyf_u_CDNS_406619531453_3.MINUS GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/comp018green_esd_rc_v5p0_0.ppolyf_u_CDNS_406619531453_1.PLUS DVDD ppolyf_u r_width=0.8u r_length=63.854996u
X118 DVDD GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/pmos_6p0_CDNS_406619531455_0.D DVSS DVSS nfet_06v0 ad=12.999999p pd=50.52u as=12.999999p ps=50.52u w=50u l=0.7u
X119 DVDD GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/pmos_6p0_CDNS_406619531455_0.D DVSS DVSS nfet_06v0 ad=12.999999p pd=50.52u as=12.999999p ps=50.52u w=50u l=0.7u
X120 DVDD GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/pmos_6p0_CDNS_406619531455_0.D DVSS DVSS nfet_06v0 ad=12.999999p pd=50.52u as=12.999999p ps=50.52u w=50u l=0.7u
X121 DVDD DVSS cap_nmos_06v0 c_width=15u c_length=15u
X122 DVSS GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/pmos_6p0_CDNS_406619531455_0.D DVDD DVSS nfet_06v0 ad=12.999999p pd=50.52u as=12.999999p ps=50.52u w=50u l=0.7u
X123 DVSS GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/pmos_6p0_CDNS_406619531455_0.D DVDD DVSS nfet_06v0 ad=12.999999p pd=50.52u as=12.999999p ps=50.52u w=50u l=0.7u
X124 DVSS GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/pmos_6p0_CDNS_406619531455_0.D DVDD DVSS nfet_06v0 ad=12.999999p pd=50.52u as=12.999999p ps=50.52u w=50u l=0.7u
X125 DVSS GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/pmos_6p0_CDNS_406619531455_0.D DVDD DVSS nfet_06v0 ad=12.999999p pd=50.52u as=12.999999p ps=50.52u w=50u l=0.7u
X126 DVSS GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/pmos_6p0_CDNS_406619531455_0.D DVDD DVSS nfet_06v0 ad=12.999999p pd=50.52u as=12.999999p ps=50.52u w=50u l=0.7u
X127 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/comp018green_esd_rc_v5p0_0.ppolyf_u_CDNS_406619531453_1.MINUS GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/comp018green_esd_rc_v5p0_0.ppolyf_u_CDNS_406619531453_1.PLUS DVDD ppolyf_u r_width=0.8u r_length=63.854996u
X128 DVDD GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/pmos_6p0_CDNS_406619531455_0.D DVSS DVSS nfet_06v0 ad=12.999999p pd=50.52u as=12.999999p ps=50.52u w=50u l=0.7u
X129 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/pmos_6p0_CDNS_406619531456_0.D GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/pmos_6p0_CDNS_406619531452_0.D DVSS DVSS nfet_06v0 ad=1.3p pd=5.52u as=1.3p ps=5.52u w=5u l=0.7u
X130 DVDD GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/pmos_6p0_CDNS_406619531455_0.D DVSS DVSS nfet_06v0 ad=12.999999p pd=50.52u as=12.999999p ps=50.52u w=50u l=0.7u
X131 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/comp018green_esd_rc_v5p0_0.ppolyf_u_CDNS_406619531453_5.MINUS GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/comp018green_esd_rc_v5p0_0.ppolyf_u_CDNS_406619531453_5.PLUS DVDD ppolyf_u r_width=0.8u r_length=63.854996u
X132 DVSS GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/pmos_6p0_CDNS_406619531455_0.D DVDD DVSS nfet_06v0 ad=12.999999p pd=50.52u as=12.999999p ps=50.52u w=50u l=0.7u
D3 DVSS DVDD diode_nd2ps_06v0 pj=82u area=40p
X133 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/pmos_6p0_CDNS_406619531455_0.D GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/pmos_6p0_CDNS_406619531456_0.D DVSS DVSS nfet_06v0 ad=1.3p pd=5.52u as=1.3p ps=5.52u w=5u l=0.7u
X134 DVDD GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/comp018green_esd_rc_v5p0_0.VRC GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/pmos_6p0_CDNS_406619531452_0.D DVDD pfet_06v0 ad=1.3p pd=5.52u as=1.3p ps=5.52u w=5u l=0.7u
X135 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/pmos_6p0_CDNS_406619531452_0.D GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/comp018green_esd_rc_v5p0_0.VRC DVDD DVDD pfet_06v0 ad=1.3p pd=5.52u as=2.2p ps=10.879999u w=5u l=0.7u
X136 DVSS GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/pmos_6p0_CDNS_406619531455_0.D DVDD DVSS nfet_06v0 ad=12.999999p pd=50.52u as=12.999999p ps=50.52u w=50u l=0.7u
X137 DVSS GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/pmos_6p0_CDNS_406619531455_0.D DVDD DVSS nfet_06v0 ad=12.999999p pd=50.52u as=12.999999p ps=50.52u w=50u l=0.7u
X138 DVSS GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/pmos_6p0_CDNS_406619531455_0.D DVDD DVSS nfet_06v0 ad=12.999999p pd=50.52u as=21.999998p ps=0.10088m w=50u l=0.7u
X139 GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/comp018green_esd_rc_v5p0_0.ppolyf_u_CDNS_406619531453_2.MINUS GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/comp018green_esd_rc_v5p0_0.ppolyf_u_CDNS_406619531453_2.PLUS DVDD ppolyf_u r_width=0.8u r_length=63.854996u
X140 DVDD GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/pmos_6p0_CDNS_406619531455_0.D DVSS DVSS nfet_06v0 ad=12.999999p pd=50.52u as=12.999999p ps=50.52u w=50u l=0.7u
X141 DVSS GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/pmos_6p0_CDNS_406619531452_0.D GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/pmos_6p0_CDNS_406619531456_0.D DVSS nfet_06v0 ad=1.3p pd=5.52u as=1.3p ps=5.52u w=5u l=0.7u
X142 DVDD GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/pmos_6p0_CDNS_406619531455_0.D DVSS DVSS nfet_06v0 ad=21.999998p pd=0.10088m as=12.999999p ps=50.52u w=50u l=0.7u
X143 DVDD GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/pmos_6p0_CDNS_406619531455_0.D DVSS DVSS nfet_06v0 ad=12.999999p pd=50.52u as=12.999999p ps=50.52u w=50u l=0.7u
X144 DVDD GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/pmos_6p0_CDNS_406619531456_0.D GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/pmos_6p0_CDNS_406619531455_0.D DVDD pfet_06v0 ad=1.3p pd=5.52u as=1.3p ps=5.52u w=5u l=0.7u
X145 DVSS GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/pmos_6p0_CDNS_406619531455_0.D DVDD DVSS nfet_06v0 ad=12.999999p pd=50.52u as=12.999999p ps=50.52u w=50u l=0.7u
X146 DVSS GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/pmos_6p0_CDNS_406619531455_0.D DVDD DVSS nfet_06v0 ad=12.999999p pd=50.52u as=12.999999p ps=50.52u w=50u l=0.7u
X147 DVSS GF_NI_DVDD_BASE_0.comp018green_esd_clamp_v5p0_DVDD_0/pmos_6p0_CDNS_406619531455_0.D DVDD DVSS nfet_06v0 ad=12.999999p pd=50.52u as=12.999999p ps=50.52u w=50u l=0.7u
.ends

